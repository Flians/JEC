/*

c5315:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jdff: 3034
	jand: 605
	jor: 419

Summary:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jdff: 3034
	jand: 605
	jor: 419

The maximum logic level gap of any gate:
	c5315: 21
*/

module rf_c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1157;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[1:0] w_G1_2;
	wire[2:0] w_G4_0;
	wire[1:0] w_G4_1;
	wire[1:0] w_G11_0;
	wire[1:0] w_G14_0;
	wire[1:0] w_G17_0;
	wire[1:0] w_G20_0;
	wire[1:0] w_G37_0;
	wire[1:0] w_G40_0;
	wire[1:0] w_G43_0;
	wire[1:0] w_G46_0;
	wire[1:0] w_G49_0;
	wire[1:0] w_G54_0;
	wire[1:0] w_G61_0;
	wire[1:0] w_G64_0;
	wire[1:0] w_G67_0;
	wire[1:0] w_G70_0;
	wire[1:0] w_G73_0;
	wire[1:0] w_G76_0;
	wire[1:0] w_G91_0;
	wire[1:0] w_G100_0;
	wire[1:0] w_G103_0;
	wire[1:0] w_G106_0;
	wire[1:0] w_G109_0;
	wire[1:0] w_G123_0;
	wire[1:0] w_G132_0;
	wire[2:0] w_G137_0;
	wire[2:0] w_G137_1;
	wire[2:0] w_G137_2;
	wire[2:0] w_G137_3;
	wire[2:0] w_G137_4;
	wire[2:0] w_G137_5;
	wire[2:0] w_G137_6;
	wire[2:0] w_G137_7;
	wire[2:0] w_G137_8;
	wire[1:0] w_G137_9;
	wire[2:0] w_G141_0;
	wire[2:0] w_G141_1;
	wire[2:0] w_G141_2;
	wire[1:0] w_G146_0;
	wire[1:0] w_G149_0;
	wire[1:0] w_G152_0;
	wire[1:0] w_G155_0;
	wire[1:0] w_G158_0;
	wire[1:0] w_G161_0;
	wire[1:0] w_G164_0;
	wire[1:0] w_G167_0;
	wire[1:0] w_G170_0;
	wire[1:0] w_G173_0;
	wire[1:0] w_G182_0;
	wire[1:0] w_G185_0;
	wire[1:0] w_G188_0;
	wire[1:0] w_G191_0;
	wire[1:0] w_G194_0;
	wire[1:0] w_G197_0;
	wire[1:0] w_G200_0;
	wire[1:0] w_G203_0;
	wire[2:0] w_G206_0;
	wire[2:0] w_G210_0;
	wire[2:0] w_G210_1;
	wire[2:0] w_G210_2;
	wire[2:0] w_G218_0;
	wire[2:0] w_G218_1;
	wire[2:0] w_G218_2;
	wire[2:0] w_G226_0;
	wire[2:0] w_G226_1;
	wire[2:0] w_G226_2;
	wire[2:0] w_G234_0;
	wire[2:0] w_G234_1;
	wire[1:0] w_G234_2;
	wire[2:0] w_G242_0;
	wire[2:0] w_G242_1;
	wire[1:0] w_G245_0;
	wire[2:0] w_G248_0;
	wire[2:0] w_G248_1;
	wire[2:0] w_G248_2;
	wire[2:0] w_G248_3;
	wire[2:0] w_G248_4;
	wire[1:0] w_G248_5;
	wire[2:0] w_G251_0;
	wire[2:0] w_G251_1;
	wire[2:0] w_G251_2;
	wire[2:0] w_G251_3;
	wire[2:0] w_G251_4;
	wire[2:0] w_G254_0;
	wire[2:0] w_G254_1;
	wire[2:0] w_G257_0;
	wire[2:0] w_G257_1;
	wire[2:0] w_G257_2;
	wire[2:0] w_G265_0;
	wire[2:0] w_G265_1;
	wire[1:0] w_G265_2;
	wire[2:0] w_G273_0;
	wire[2:0] w_G273_1;
	wire[2:0] w_G273_2;
	wire[1:0] w_G280_0;
	wire[2:0] w_G281_0;
	wire[2:0] w_G281_1;
	wire[1:0] w_G281_2;
	wire[1:0] w_G289_0;
	wire[2:0] w_G293_0;
	wire[2:0] w_G299_0;
	wire[2:0] w_G302_0;
	wire[2:0] w_G308_0;
	wire[2:0] w_G308_1;
	wire[2:0] w_G316_0;
	wire[2:0] w_G316_1;
	wire[2:0] w_G324_0;
	wire[2:0] w_G324_1;
	wire[1:0] w_G331_0;
	wire[2:0] w_G332_0;
	wire[2:0] w_G332_1;
	wire[2:0] w_G332_2;
	wire[2:0] w_G332_3;
	wire[2:0] w_G332_4;
	wire[2:0] w_G335_0;
	wire[2:0] w_G335_1;
	wire[2:0] w_G335_2;
	wire[2:0] w_G335_3;
	wire[1:0] w_G335_4;
	wire[2:0] w_G341_0;
	wire[2:0] w_G341_1;
	wire[2:0] w_G341_2;
	wire[1:0] w_G348_0;
	wire[2:0] w_G351_0;
	wire[2:0] w_G351_1;
	wire[2:0] w_G351_2;
	wire[1:0] w_G358_0;
	wire[2:0] w_G361_0;
	wire[1:0] w_G369_0;
	wire[2:0] w_G374_0;
	wire[2:0] w_G389_0;
	wire[2:0] w_G400_0;
	wire[1:0] w_G400_1;
	wire[2:0] w_G411_0;
	wire[2:0] w_G422_0;
	wire[2:0] w_G422_1;
	wire[1:0] w_G422_2;
	wire[2:0] w_G435_0;
	wire[2:0] w_G435_1;
	wire[2:0] w_G446_0;
	wire[2:0] w_G446_1;
	wire[2:0] w_G457_0;
	wire[2:0] w_G457_1;
	wire[1:0] w_G457_2;
	wire[2:0] w_G468_0;
	wire[2:0] w_G468_1;
	wire[2:0] w_G479_0;
	wire[1:0] w_G479_1;
	wire[2:0] w_G490_0;
	wire[2:0] w_G490_1;
	wire[2:0] w_G503_0;
	wire[2:0] w_G503_1;
	wire[2:0] w_G514_0;
	wire[1:0] w_G514_1;
	wire[2:0] w_G523_0;
	wire[1:0] w_G523_1;
	wire[2:0] w_G534_0;
	wire[2:0] w_G534_1;
	wire[2:0] w_G545_0;
	wire[2:0] w_G549_0;
	wire[1:0] w_G552_0;
	wire[1:0] w_G559_0;
	wire[1:0] w_G562_0;
	wire[2:0] w_G1497_0;
	wire[2:0] w_G1689_0;
	wire[2:0] w_G1690_0;
	wire[2:0] w_G1691_0;
	wire[2:0] w_G1694_0;
	wire[2:0] w_G2174_0;
	wire[2:0] w_G2358_0;
	wire[2:0] w_G2358_1;
	wire[2:0] w_G2358_2;
	wire[1:0] w_G3173_0;
	wire[2:0] w_G3546_0;
	wire[2:0] w_G3546_1;
	wire[2:0] w_G3546_2;
	wire[2:0] w_G3546_3;
	wire[2:0] w_G3546_4;
	wire[1:0] w_G3546_5;
	wire[2:0] w_G3548_0;
	wire[2:0] w_G3548_1;
	wire[2:0] w_G3548_2;
	wire[2:0] w_G3548_3;
	wire[2:0] w_G3548_4;
	wire[1:0] w_G3552_0;
	wire[1:0] w_G3717_0;
	wire[2:0] w_G3724_0;
	wire[2:0] w_G4087_0;
	wire[2:0] w_G4088_0;
	wire[2:0] w_G4089_0;
	wire[2:0] w_G4090_0;
	wire[2:0] w_G4091_0;
	wire[2:0] w_G4091_1;
	wire[2:0] w_G4091_2;
	wire[2:0] w_G4092_0;
	wire[2:0] w_G4092_1;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G600_0;
	wire G600_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G611_0;
	wire G611_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire[2:0] w_G809_0;
	wire[2:0] w_G809_1;
	wire[2:0] w_G809_2;
	wire[1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G1000_0;
	wire G1000_fa_;
	wire w_G826_0;
	wire G826_fa_;
	wire w_G828_0;
	wire G828_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G867_0;
	wire G867_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire[1:0] w_n316_0;
	wire[1:0] w_n318_0;
	wire[2:0] w_n326_0;
	wire[2:0] w_n326_1;
	wire[1:0] w_n326_2;
	wire[1:0] w_n333_0;
	wire[1:0] w_n336_0;
	wire[1:0] w_n360_0;
	wire[1:0] w_n362_0;
	wire[2:0] w_n366_0;
	wire[2:0] w_n366_1;
	wire[2:0] w_n366_2;
	wire[2:0] w_n366_3;
	wire[2:0] w_n366_4;
	wire[2:0] w_n368_0;
	wire[2:0] w_n368_1;
	wire[2:0] w_n368_2;
	wire[2:0] w_n368_3;
	wire[2:0] w_n368_4;
	wire[1:0] w_n368_5;
	wire[2:0] w_n372_0;
	wire[1:0] w_n373_0;
	wire[2:0] w_n383_0;
	wire[2:0] w_n385_0;
	wire[2:0] w_n385_1;
	wire[2:0] w_n386_0;
	wire[2:0] w_n386_1;
	wire[2:0] w_n386_2;
	wire[2:0] w_n386_3;
	wire[2:0] w_n386_4;
	wire[2:0] w_n388_0;
	wire[2:0] w_n388_1;
	wire[2:0] w_n389_0;
	wire[2:0] w_n389_1;
	wire[2:0] w_n389_2;
	wire[2:0] w_n389_3;
	wire[2:0] w_n389_4;
	wire[1:0] w_n397_0;
	wire[2:0] w_n398_0;
	wire[2:0] w_n401_0;
	wire[2:0] w_n402_0;
	wire[2:0] w_n402_1;
	wire[1:0] w_n402_2;
	wire[1:0] w_n403_0;
	wire[2:0] w_n405_0;
	wire[2:0] w_n405_1;
	wire[1:0] w_n405_2;
	wire[1:0] w_n407_0;
	wire[1:0] w_n408_0;
	wire[2:0] w_n410_0;
	wire[1:0] w_n410_1;
	wire[1:0] w_n414_0;
	wire[1:0] w_n416_0;
	wire[2:0] w_n419_0;
	wire[2:0] w_n424_0;
	wire[2:0] w_n424_1;
	wire[1:0] w_n424_2;
	wire[1:0] w_n426_0;
	wire[1:0] w_n434_0;
	wire[2:0] w_n435_0;
	wire[2:0] w_n435_1;
	wire[2:0] w_n437_0;
	wire[2:0] w_n437_1;
	wire[1:0] w_n445_0;
	wire[2:0] w_n449_0;
	wire[2:0] w_n449_1;
	wire[2:0] w_n451_0;
	wire[1:0] w_n451_1;
	wire[1:0] w_n459_0;
	wire[2:0] w_n460_0;
	wire[2:0] w_n460_1;
	wire[2:0] w_n462_0;
	wire[1:0] w_n470_0;
	wire[2:0] w_n471_0;
	wire[1:0] w_n471_1;
	wire[2:0] w_n473_0;
	wire[2:0] w_n473_1;
	wire[1:0] w_n481_0;
	wire[2:0] w_n484_0;
	wire[1:0] w_n484_1;
	wire[2:0] w_n486_0;
	wire[1:0] w_n486_1;
	wire[1:0] w_n494_0;
	wire[2:0] w_n495_0;
	wire[2:0] w_n495_1;
	wire[2:0] w_n497_0;
	wire[1:0] w_n497_1;
	wire[1:0] w_n505_0;
	wire[2:0] w_n507_0;
	wire[1:0] w_n507_1;
	wire[1:0] w_n509_0;
	wire[1:0] w_n517_0;
	wire[2:0] w_n518_0;
	wire[1:0] w_n518_1;
	wire[2:0] w_n528_0;
	wire[2:0] w_n530_0;
	wire[1:0] w_n530_1;
	wire[1:0] w_n532_0;
	wire[1:0] w_n540_0;
	wire[2:0] w_n541_0;
	wire[1:0] w_n541_1;
	wire[1:0] w_n543_0;
	wire[1:0] w_n551_0;
	wire[2:0] w_n556_0;
	wire[2:0] w_n556_1;
	wire[2:0] w_n556_2;
	wire[2:0] w_n556_3;
	wire[2:0] w_n556_4;
	wire[1:0] w_n556_5;
	wire[2:0] w_n560_0;
	wire[1:0] w_n560_1;
	wire[2:0] w_n561_0;
	wire[1:0] w_n562_0;
	wire[2:0] w_n566_0;
	wire[2:0] w_n567_0;
	wire[1:0] w_n567_1;
	wire[1:0] w_n569_0;
	wire[1:0] w_n570_0;
	wire[2:0] w_n571_0;
	wire[1:0] w_n571_1;
	wire[2:0] w_n572_0;
	wire[2:0] w_n574_0;
	wire[2:0] w_n577_0;
	wire[2:0] w_n578_0;
	wire[2:0] w_n582_0;
	wire[1:0] w_n582_1;
	wire[2:0] w_n583_0;
	wire[1:0] w_n583_1;
	wire[1:0] w_n585_0;
	wire[2:0] w_n587_0;
	wire[1:0] w_n587_1;
	wire[2:0] w_n590_0;
	wire[1:0] w_n590_1;
	wire[1:0] w_n591_0;
	wire[2:0] w_n595_0;
	wire[1:0] w_n595_1;
	wire[2:0] w_n596_0;
	wire[2:0] w_n600_0;
	wire[1:0] w_n600_1;
	wire[1:0] w_n601_0;
	wire[2:0] w_n604_0;
	wire[2:0] w_n605_0;
	wire[2:0] w_n605_1;
	wire[2:0] w_n605_2;
	wire[2:0] w_n607_0;
	wire[2:0] w_n609_0;
	wire[2:0] w_n609_1;
	wire[2:0] w_n609_2;
	wire[2:0] w_n609_3;
	wire[2:0] w_n609_4;
	wire[2:0] w_n609_5;
	wire[2:0] w_n613_0;
	wire[2:0] w_n614_0;
	wire[2:0] w_n614_1;
	wire[1:0] w_n614_2;
	wire[2:0] w_n617_0;
	wire[1:0] w_n617_1;
	wire[2:0] w_n618_0;
	wire[1:0] w_n618_1;
	wire[2:0] w_n621_0;
	wire[2:0] w_n621_1;
	wire[1:0] w_n621_2;
	wire[2:0] w_n622_0;
	wire[1:0] w_n622_1;
	wire[1:0] w_n623_0;
	wire[2:0] w_n624_0;
	wire[2:0] w_n624_1;
	wire[2:0] w_n625_0;
	wire[2:0] w_n628_0;
	wire[2:0] w_n629_0;
	wire[1:0] w_n631_0;
	wire[2:0] w_n633_0;
	wire[1:0] w_n633_1;
	wire[2:0] w_n636_0;
	wire[1:0] w_n636_1;
	wire[2:0] w_n640_0;
	wire[2:0] w_n640_1;
	wire[1:0] w_n641_0;
	wire[1:0] w_n642_0;
	wire[2:0] w_n645_0;
	wire[2:0] w_n646_0;
	wire[2:0] w_n649_0;
	wire[1:0] w_n649_1;
	wire[1:0] w_n650_0;
	wire[2:0] w_n651_0;
	wire[1:0] w_n651_1;
	wire[1:0] w_n652_0;
	wire[1:0] w_n661_0;
	wire[1:0] w_n671_0;
	wire[1:0] w_n677_0;
	wire[1:0] w_n678_0;
	wire[1:0] w_n679_0;
	wire[1:0] w_n680_0;
	wire[2:0] w_n681_0;
	wire[2:0] w_n681_1;
	wire[1:0] w_n681_2;
	wire[1:0] w_n682_0;
	wire[2:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[2:0] w_n691_0;
	wire[2:0] w_n693_0;
	wire[2:0] w_n696_0;
	wire[1:0] w_n697_0;
	wire[1:0] w_n700_0;
	wire[1:0] w_n702_0;
	wire[2:0] w_n703_0;
	wire[1:0] w_n705_0;
	wire[1:0] w_n706_0;
	wire[2:0] w_n707_0;
	wire[1:0] w_n709_0;
	wire[1:0] w_n716_0;
	wire[2:0] w_n717_0;
	wire[1:0] w_n720_0;
	wire[2:0] w_n721_0;
	wire[1:0] w_n723_0;
	wire[1:0] w_n726_0;
	wire[2:0] w_n727_0;
	wire[2:0] w_n729_0;
	wire[1:0] w_n729_1;
	wire[2:0] w_n732_0;
	wire[1:0] w_n733_0;
	wire[1:0] w_n735_0;
	wire[1:0] w_n736_0;
	wire[2:0] w_n739_0;
	wire[1:0] w_n739_1;
	wire[1:0] w_n740_0;
	wire[1:0] w_n741_0;
	wire[1:0] w_n742_0;
	wire[2:0] w_n744_0;
	wire[2:0] w_n744_1;
	wire[2:0] w_n746_0;
	wire[2:0] w_n746_1;
	wire[2:0] w_n747_0;
	wire[2:0] w_n747_1;
	wire[2:0] w_n747_2;
	wire[2:0] w_n747_3;
	wire[2:0] w_n748_0;
	wire[2:0] w_n748_1;
	wire[2:0] w_n748_2;
	wire[2:0] w_n748_3;
	wire[1:0] w_n748_4;
	wire[2:0] w_n750_0;
	wire[1:0] w_n750_1;
	wire[2:0] w_n751_0;
	wire[2:0] w_n751_1;
	wire[1:0] w_n751_2;
	wire[2:0] w_n753_0;
	wire[2:0] w_n753_1;
	wire[2:0] w_n753_2;
	wire[2:0] w_n753_3;
	wire[2:0] w_n753_4;
	wire[2:0] w_n753_5;
	wire[2:0] w_n753_6;
	wire[2:0] w_n753_7;
	wire[1:0] w_n753_8;
	wire[1:0] w_n759_0;
	wire[1:0] w_n760_0;
	wire[1:0] w_n761_0;
	wire[2:0] w_n765_0;
	wire[2:0] w_n765_1;
	wire[2:0] w_n765_2;
	wire[2:0] w_n765_3;
	wire[2:0] w_n765_4;
	wire[2:0] w_n765_5;
	wire[1:0] w_n771_0;
	wire[1:0] w_n779_0;
	wire[2:0] w_n781_0;
	wire[2:0] w_n783_0;
	wire[1:0] w_n783_1;
	wire[1:0] w_n786_0;
	wire[1:0] w_n787_0;
	wire[2:0] w_n789_0;
	wire[2:0] w_n791_0;
	wire[1:0] w_n791_1;
	wire[1:0] w_n792_0;
	wire[2:0] w_n793_0;
	wire[2:0] w_n793_1;
	wire[2:0] w_n793_2;
	wire[2:0] w_n793_3;
	wire[1:0] w_n793_4;
	wire[2:0] w_n795_0;
	wire[1:0] w_n795_1;
	wire[1:0] w_n796_0;
	wire[2:0] w_n797_0;
	wire[2:0] w_n797_1;
	wire[2:0] w_n797_2;
	wire[2:0] w_n797_3;
	wire[1:0] w_n797_4;
	wire[2:0] w_n799_0;
	wire[2:0] w_n799_1;
	wire[2:0] w_n799_2;
	wire[2:0] w_n799_3;
	wire[1:0] w_n799_4;
	wire[2:0] w_n801_0;
	wire[2:0] w_n801_1;
	wire[2:0] w_n801_2;
	wire[2:0] w_n801_3;
	wire[1:0] w_n801_4;
	wire[2:0] w_n806_0;
	wire[1:0] w_n809_0;
	wire[1:0] w_n819_0;
	wire[1:0] w_n821_0;
	wire[2:0] w_n828_0;
	wire[1:0] w_n829_0;
	wire[1:0] w_n832_0;
	wire[1:0] w_n839_0;
	wire[2:0] w_n840_0;
	wire[2:0] w_n840_1;
	wire[2:0] w_n840_2;
	wire[2:0] w_n840_3;
	wire[1:0] w_n840_4;
	wire[1:0] w_n842_0;
	wire[2:0] w_n843_0;
	wire[2:0] w_n843_1;
	wire[2:0] w_n843_2;
	wire[2:0] w_n843_3;
	wire[1:0] w_n843_4;
	wire[2:0] w_n845_0;
	wire[2:0] w_n845_1;
	wire[2:0] w_n845_2;
	wire[2:0] w_n845_3;
	wire[1:0] w_n845_4;
	wire[2:0] w_n847_0;
	wire[2:0] w_n847_1;
	wire[2:0] w_n847_2;
	wire[2:0] w_n847_3;
	wire[1:0] w_n847_4;
	wire[1:0] w_n853_0;
	wire[1:0] w_n855_0;
	wire[1:0] w_n856_0;
	wire[1:0] w_n857_0;
	wire[1:0] w_n859_0;
	wire[1:0] w_n862_0;
	wire[1:0] w_n869_0;
	wire[1:0] w_n877_0;
	wire[1:0] w_n879_0;
	wire[1:0] w_n881_0;
	wire[1:0] w_n892_0;
	wire[1:0] w_n914_0;
	wire[1:0] w_n928_0;
	wire[2:0] w_n930_0;
	wire[1:0] w_n932_0;
	wire[2:0] w_n936_0;
	wire[1:0] w_n938_0;
	wire[1:0] w_n941_0;
	wire[1:0] w_n943_0;
	wire[1:0] w_n944_0;
	wire[1:0] w_n946_0;
	wire[2:0] w_n948_0;
	wire[1:0] w_n953_0;
	wire[1:0] w_n954_0;
	wire[1:0] w_n968_0;
	wire[1:0] w_n971_0;
	wire[1:0] w_n972_0;
	wire[1:0] w_n973_0;
	wire[1:0] w_n984_0;
	wire[2:0] w_n985_0;
	wire[2:0] w_n985_1;
	wire[2:0] w_n985_2;
	wire[2:0] w_n985_3;
	wire[1:0] w_n985_4;
	wire[1:0] w_n987_0;
	wire[2:0] w_n988_0;
	wire[2:0] w_n988_1;
	wire[2:0] w_n988_2;
	wire[2:0] w_n988_3;
	wire[1:0] w_n988_4;
	wire[2:0] w_n990_0;
	wire[2:0] w_n990_1;
	wire[2:0] w_n990_2;
	wire[2:0] w_n990_3;
	wire[1:0] w_n990_4;
	wire[2:0] w_n992_0;
	wire[2:0] w_n992_1;
	wire[2:0] w_n992_2;
	wire[2:0] w_n992_3;
	wire[1:0] w_n992_4;
	wire[1:0] w_n998_0;
	wire[2:0] w_n999_0;
	wire[2:0] w_n999_1;
	wire[2:0] w_n999_2;
	wire[2:0] w_n999_3;
	wire[1:0] w_n999_4;
	wire[1:0] w_n1001_0;
	wire[2:0] w_n1002_0;
	wire[2:0] w_n1002_1;
	wire[2:0] w_n1002_2;
	wire[2:0] w_n1002_3;
	wire[1:0] w_n1002_4;
	wire[2:0] w_n1004_0;
	wire[2:0] w_n1004_1;
	wire[2:0] w_n1004_2;
	wire[2:0] w_n1004_3;
	wire[1:0] w_n1004_4;
	wire[2:0] w_n1006_0;
	wire[2:0] w_n1006_1;
	wire[2:0] w_n1006_2;
	wire[2:0] w_n1006_3;
	wire[1:0] w_n1006_4;
	wire[2:0] w_n1012_0;
	wire[1:0] w_n1012_1;
	wire[2:0] w_n1014_0;
	wire[1:0] w_n1014_1;
	wire[2:0] w_n1021_0;
	wire[1:0] w_n1021_1;
	wire[2:0] w_n1023_0;
	wire[1:0] w_n1023_1;
	wire[2:0] w_n1030_0;
	wire[1:0] w_n1030_1;
	wire[2:0] w_n1032_0;
	wire[1:0] w_n1032_1;
	wire[2:0] w_n1039_0;
	wire[1:0] w_n1039_1;
	wire[2:0] w_n1041_0;
	wire[1:0] w_n1041_1;
	wire[1:0] w_n1142_0;
	wire[1:0] w_n1151_0;
	wire[2:0] w_n1163_0;
	wire[2:0] w_n1163_1;
	wire[2:0] w_n1197_0;
	wire[2:0] w_n1197_1;
	wire[2:0] w_n1205_0;
	wire[2:0] w_n1205_1;
	wire[2:0] w_n1235_0;
	wire[1:0] w_n1235_1;
	wire[2:0] w_n1242_0;
	wire[1:0] w_n1242_1;
	wire[2:0] w_n1244_0;
	wire[1:0] w_n1244_1;
	wire[2:0] w_n1251_0;
	wire[1:0] w_n1251_1;
	wire[2:0] w_n1253_0;
	wire[1:0] w_n1253_1;
	wire[1:0] w_n1358_0;
	wire[1:0] w_n1383_0;
	wire[1:0] w_n1391_0;
	wire[1:0] w_n1394_0;
	wire[1:0] w_n1398_0;
	wire[1:0] w_n1399_0;
	wire[1:0] w_n1409_0;
	wire[1:0] w_n1410_0;
	wire[1:0] w_n1411_0;
	wire[1:0] w_n1421_0;
	wire[1:0] w_n1425_0;
	wire[1:0] w_n1434_0;
	wire[1:0] w_n1438_0;
	wire[1:0] w_n1445_0;
	wire[1:0] w_n1446_0;
	wire[1:0] w_n1447_0;
	wire[1:0] w_n1452_0;
	wire[1:0] w_n1494_0;
	wire[1:0] w_n1533_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1545_0;
	wire[1:0] w_n1553_0;
	wire[1:0] w_n1555_0;
	wire[1:0] w_n1560_0;
	wire[1:0] w_n1568_0;
	wire[1:0] w_n1591_0;
	wire[1:0] w_n1597_0;
	wire[2:0] w_n1601_0;
	wire[1:0] w_n1602_0;
	wire[1:0] w_n1609_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1624_0;
	wire[1:0] w_n1629_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1634_0;
	wire w_dff_B_RzBELWjC6_1;
	wire w_dff_B_JWqUGSMZ8_0;
	wire w_dff_B_ptZ81eDE6_1;
	wire w_dff_B_OAjlNXEo5_1;
	wire w_dff_B_FWUboPEb9_2;
	wire w_dff_B_8DrVy7Dt6_1;
	wire w_dff_B_bHJaaGt51_1;
	wire w_dff_B_qX6aa1gp2_0;
	wire w_dff_B_3tVcDugs0_1;
	wire w_dff_B_HADBglPu0_0;
	wire w_dff_A_9C0pgMBL7_0;
	wire w_dff_A_C3bV5UDH8_0;
	wire w_dff_A_kXzyRFoB3_0;
	wire w_dff_A_Q4mVXVSm9_0;
	wire w_dff_A_ZObNW4Ey2_1;
	wire w_dff_A_B86FrkrD4_1;
	wire w_dff_A_COhjQtNa9_1;
	wire w_dff_A_IVtEBFxm4_1;
	wire w_dff_B_vFmQ5TlV0_1;
	wire w_dff_B_YDEUWMNi4_0;
	wire w_dff_B_f2fpSkCN8_1;
	wire w_dff_B_wmy6YsLa3_0;
	wire w_dff_A_ZxugpCx67_1;
	wire w_dff_A_DrQHCVWM3_1;
	wire w_dff_A_PvaVoCTq9_1;
	wire w_dff_A_TiUCt4UZ9_1;
	wire w_dff_A_gN7N4X8q9_2;
	wire w_dff_A_mg8gFpYf6_2;
	wire w_dff_A_WTy7MJiF3_2;
	wire w_dff_A_c4hnKAkf8_2;
	wire w_dff_B_iKaawZhP2_1;
	wire w_dff_B_kgDrTsHG1_1;
	wire w_dff_B_k2BhBUC50_1;
	wire w_dff_B_uaqFFGz90_2;
	wire w_dff_B_fWpcCLRF3_2;
	wire w_dff_B_eHWaVUCs6_2;
	wire w_dff_B_ukggaXHx1_2;
	wire w_dff_B_QishoWLg1_2;
	wire w_dff_B_mOqa1OGg6_2;
	wire w_dff_B_ZSLKpmE55_2;
	wire w_dff_B_R69B89aU0_2;
	wire w_dff_B_HG903BB55_2;
	wire w_dff_A_OW39dcyk1_0;
	wire w_dff_A_GtpwQz4h7_0;
	wire w_dff_A_ZXz8anXH0_0;
	wire w_dff_A_xsnU0FGa5_0;
	wire w_dff_A_yUFgaqvw7_0;
	wire w_dff_A_hirtmZVm7_0;
	wire w_dff_B_mKOBTZB24_0;
	wire w_dff_B_2lQ0J8dv0_0;
	wire w_dff_B_uiqNtDor1_0;
	wire w_dff_B_ic366AMP9_0;
	wire w_dff_B_o5YSYmXM7_0;
	wire w_dff_B_YP1E7uEv8_0;
	wire w_dff_B_0LWkBtLA4_0;
	wire w_dff_B_RWa4FnYE8_0;
	wire w_dff_B_4EWw5jV12_0;
	wire w_dff_B_BaO8iXGJ0_0;
	wire w_dff_B_VpSRf2wQ8_0;
	wire w_dff_B_dXMUhcYZ7_0;
	wire w_dff_B_YzYh7TTY3_0;
	wire w_dff_B_k9iDq4bf2_0;
	wire w_dff_B_umkbvgcF8_0;
	wire w_dff_B_gMOCBXgU4_0;
	wire w_dff_B_7rs07MRI9_0;
	wire w_dff_B_KdGRFTnr7_0;
	wire w_dff_B_x0AhPXlO8_0;
	wire w_dff_B_9prtjbAa3_0;
	wire w_dff_B_HzcAlp7l2_0;
	wire w_dff_B_gMxSx6Ho5_0;
	wire w_dff_B_ca9zya6x5_0;
	wire w_dff_B_gpB42W571_0;
	wire w_dff_B_H2TjMq3a0_0;
	wire w_dff_B_AMDlZ77B5_0;
	wire w_dff_B_0wHZ84El8_1;
	wire w_dff_B_3UTEDciD9_0;
	wire w_dff_B_0wMPxvlQ4_0;
	wire w_dff_B_II81o4S52_0;
	wire w_dff_B_nptmKkUZ1_0;
	wire w_dff_B_2hotGX0c9_0;
	wire w_dff_B_nDnBkqnF8_0;
	wire w_dff_B_4pV60Ame4_0;
	wire w_dff_B_IDIr9lHx6_0;
	wire w_dff_B_GUp9kupK6_0;
	wire w_dff_B_o8EYHMOg5_0;
	wire w_dff_B_7HyvhXRI1_0;
	wire w_dff_B_8rz9pWQc7_0;
	wire w_dff_B_Q3Wm8lkY8_0;
	wire w_dff_A_PB21WzYN0_0;
	wire w_dff_A_6OXAzj3g5_0;
	wire w_dff_A_2DuL7SYO4_0;
	wire w_dff_A_gCDMYwaD2_0;
	wire w_dff_A_ueYTv5xU0_0;
	wire w_dff_A_M8ldEAB83_0;
	wire w_dff_A_3leGPe2H6_0;
	wire w_dff_A_0aM3uvZb7_0;
	wire w_dff_A_jkpXis341_0;
	wire w_dff_A_lU0dF5Bv0_0;
	wire w_dff_A_mwdpgRYx4_0;
	wire w_dff_A_ekywUrWf7_0;
	wire w_dff_A_mkqb6dMC3_0;
	wire w_dff_A_T2sGO75z4_0;
	wire w_dff_A_rNTfHfPH9_0;
	wire w_dff_B_O8lDN2Ov1_0;
	wire w_dff_B_fwOQSZm62_0;
	wire w_dff_B_icSoDn673_0;
	wire w_dff_B_YGzhREhr9_0;
	wire w_dff_B_4USECAa41_0;
	wire w_dff_B_Pn8onG5L1_0;
	wire w_dff_B_PooRPk5o2_0;
	wire w_dff_B_iOivrpSl1_0;
	wire w_dff_B_fIDJAEzU8_0;
	wire w_dff_B_S4DsBMNP4_0;
	wire w_dff_B_0qEmyr9a0_0;
	wire w_dff_B_26fQGdqr6_0;
	wire w_dff_B_qyYTazVA2_0;
	wire w_dff_B_yWOP5syg3_0;
	wire w_dff_B_tiZsxCVD0_0;
	wire w_dff_B_YIK1oPkM0_0;
	wire w_dff_B_cYoiz19V4_0;
	wire w_dff_B_xZN0ED6Q6_0;
	wire w_dff_B_PC2KF1KL5_0;
	wire w_dff_B_3VDSy90D4_0;
	wire w_dff_B_7x1yOwOB6_0;
	wire w_dff_B_6f2NhJRQ0_0;
	wire w_dff_B_DWLt45xz0_0;
	wire w_dff_B_jAtPmFYd6_0;
	wire w_dff_B_2sCn4Gkj0_0;
	wire w_dff_B_kRNEjy8b1_0;
	wire w_dff_B_DEOkiNkd0_0;
	wire w_dff_B_c4SzRoxO9_0;
	wire w_dff_B_eehwCpWg4_0;
	wire w_dff_B_Lylrgo3b1_0;
	wire w_dff_A_iXVDWhc73_1;
	wire w_dff_A_flohxssd4_1;
	wire w_dff_A_tAJ90iUP1_2;
	wire w_dff_A_wjNf8aSE5_2;
	wire w_dff_A_IjFKvcOz3_2;
	wire w_dff_A_km2ZL4Gp9_2;
	wire w_dff_A_JeyMDLcV1_1;
	wire w_dff_A_U2G2gjC92_2;
	wire w_dff_A_bGOD6Vfc2_2;
	wire w_dff_B_WLJDP7aX5_0;
	wire w_dff_B_hyVEFCOX6_0;
	wire w_dff_B_bp8oz2Yp3_0;
	wire w_dff_B_SV85jtcn9_0;
	wire w_dff_B_NcgEUrkH8_0;
	wire w_dff_B_0FqPBkLi0_0;
	wire w_dff_B_H9MgKrMR1_0;
	wire w_dff_B_4vtpxsRP6_0;
	wire w_dff_B_n19WXVD79_0;
	wire w_dff_B_ML3hLjTP6_0;
	wire w_dff_B_DUNvPQbT4_0;
	wire w_dff_B_TmxpdT241_0;
	wire w_dff_B_1xC9NPUj3_0;
	wire w_dff_A_UFT1gAXt4_0;
	wire w_dff_A_SLDxeEnB5_0;
	wire w_dff_A_nvwh3Ayz7_0;
	wire w_dff_A_BlE8r4On6_0;
	wire w_dff_A_YAPHpsN59_0;
	wire w_dff_A_89UIB3AV2_0;
	wire w_dff_A_f5jDzHUl3_0;
	wire w_dff_A_Dn6AKhlp1_0;
	wire w_dff_A_V2AWPLil1_0;
	wire w_dff_A_NEcVzGTV4_0;
	wire w_dff_A_V9dJ05ZL2_0;
	wire w_dff_A_5g7Q5P4u8_0;
	wire w_dff_A_SODyiXzN0_0;
	wire w_dff_A_JpJbzvPb0_0;
	wire w_dff_A_fxS3wW5c0_0;
	wire w_dff_B_QY6h3Pf56_0;
	wire w_dff_B_9s8bNhxA6_0;
	wire w_dff_B_EXUBk9iq9_0;
	wire w_dff_B_bvpstB1Y4_0;
	wire w_dff_B_HME17iCn7_0;
	wire w_dff_B_pbUwHfwR9_0;
	wire w_dff_B_kmZmkbn24_0;
	wire w_dff_B_rGgHRLoE1_0;
	wire w_dff_B_lHVgOqDK4_0;
	wire w_dff_B_uIX37U5y7_0;
	wire w_dff_B_JMXQfCuI4_0;
	wire w_dff_B_COsA15oz2_0;
	wire w_dff_B_1oV735lj2_0;
	wire w_dff_B_Bw4APaHX1_0;
	wire w_dff_B_L4X6iy017_0;
	wire w_dff_B_jLJQThCl5_0;
	wire w_dff_B_VkH9BJvj3_0;
	wire w_dff_B_c8FW5eSL9_0;
	wire w_dff_B_o0NNZpMN0_0;
	wire w_dff_B_Ye1H5Dwo8_0;
	wire w_dff_B_TCuaHdYd2_0;
	wire w_dff_B_l7mRFPEA2_0;
	wire w_dff_B_VtPGMql03_0;
	wire w_dff_B_mqzvoDyA5_0;
	wire w_dff_B_MhN27Q6f9_0;
	wire w_dff_B_2W4kTnps9_0;
	wire w_dff_B_2eOnCZPV5_0;
	wire w_dff_B_hdNBlLk22_0;
	wire w_dff_B_2HS9pGTJ6_0;
	wire w_dff_B_CotwCRay0_0;
	wire w_dff_A_alt0yisF4_1;
	wire w_dff_A_j2B9s7A08_1;
	wire w_dff_A_imaJQpu46_2;
	wire w_dff_A_UWynk47f2_2;
	wire w_dff_A_WuBffQWu7_2;
	wire w_dff_A_HIp2utQk6_2;
	wire w_dff_A_2ZX1RZLv2_1;
	wire w_dff_A_NejeZ81z2_2;
	wire w_dff_A_lkHYSTEn1_2;
	wire w_dff_B_5PjVobUQ4_0;
	wire w_dff_B_I1otXkx41_0;
	wire w_dff_B_bDqmygbW1_0;
	wire w_dff_B_yJnZLiSd8_0;
	wire w_dff_B_bB0Sr1Gj6_0;
	wire w_dff_B_QZeE7Yp02_0;
	wire w_dff_B_5xzEO4Rc1_0;
	wire w_dff_B_ziWQ1k7Z5_0;
	wire w_dff_B_VByOyEj53_0;
	wire w_dff_B_DziEf5Bx5_0;
	wire w_dff_B_Zo5WcvMW7_0;
	wire w_dff_B_kZVqFo4l3_0;
	wire w_dff_B_3ID8azaP2_0;
	wire w_dff_A_4APADHfG0_0;
	wire w_dff_A_jcdf759Q8_0;
	wire w_dff_A_rKq1Rlm87_0;
	wire w_dff_A_a8eUjuHY3_0;
	wire w_dff_A_0vywOJOq4_0;
	wire w_dff_A_9yAP0nK09_0;
	wire w_dff_A_SOjh66Ht0_0;
	wire w_dff_A_UpiIgfVy1_0;
	wire w_dff_A_fsVXSeFl0_0;
	wire w_dff_A_cy8CQDxH4_0;
	wire w_dff_A_zzzPEC1N0_0;
	wire w_dff_A_964eO37u6_0;
	wire w_dff_A_4kvJzyfI4_0;
	wire w_dff_A_KlEHEaxs4_0;
	wire w_dff_A_H1Eerfff1_0;
	wire w_dff_B_n8QyPZdT5_0;
	wire w_dff_B_J89I7pNR6_0;
	wire w_dff_B_AjhPezaV8_0;
	wire w_dff_B_hl0GFvEU1_0;
	wire w_dff_B_59bO7vdM3_0;
	wire w_dff_B_5A4vBxa52_0;
	wire w_dff_B_gBCqngKc3_0;
	wire w_dff_B_mFkarUnK7_0;
	wire w_dff_B_mVA8vvvh4_0;
	wire w_dff_B_QUZvArLB3_0;
	wire w_dff_B_dZoSkuxT9_0;
	wire w_dff_B_qiUae91M4_0;
	wire w_dff_B_mUnvMIsE0_0;
	wire w_dff_B_e6Alg1Mr6_0;
	wire w_dff_B_GoOfclq14_0;
	wire w_dff_B_w8BDqJrV8_0;
	wire w_dff_B_hmhDHuWd3_0;
	wire w_dff_B_oCB45nCt6_0;
	wire w_dff_B_Wb3Mxokv3_0;
	wire w_dff_A_OlofKs7A9_0;
	wire w_dff_A_bREHY6Oa2_2;
	wire w_dff_A_eOWBWetz2_2;
	wire w_dff_A_jpqL0GFx2_2;
	wire w_dff_A_WB8BAewC6_2;
	wire w_dff_B_8LNnabtE7_0;
	wire w_dff_B_6w2Kod5f0_0;
	wire w_dff_B_hmWfcwRY6_0;
	wire w_dff_B_rr7bKtVM8_0;
	wire w_dff_B_WuTUTdSS1_0;
	wire w_dff_B_6HsbXZa65_0;
	wire w_dff_B_i1eWqLSa7_0;
	wire w_dff_B_G396cFwj5_0;
	wire w_dff_B_0EXkct223_0;
	wire w_dff_B_laPSel7d8_0;
	wire w_dff_B_3mQ230dl9_0;
	wire w_dff_A_uDFr2mIy1_0;
	wire w_dff_A_AYsweUT61_0;
	wire w_dff_A_gVcqTXIN4_0;
	wire w_dff_A_vx7I6ae47_0;
	wire w_dff_A_d1pj2AEB0_1;
	wire w_dff_A_WOHbjGuG2_1;
	wire w_dff_A_qna2aV5G5_0;
	wire w_dff_A_GmbTiMEO1_0;
	wire w_dff_A_XxnP5lNH6_1;
	wire w_dff_B_wJYACATe1_0;
	wire w_dff_B_7JyMLTIr8_0;
	wire w_dff_B_eEsi5fVW9_0;
	wire w_dff_B_It73lj5j5_0;
	wire w_dff_B_yIlIV1J45_0;
	wire w_dff_B_plmtYHbb9_0;
	wire w_dff_B_l5u8Te2Z8_0;
	wire w_dff_B_8UNPt5Sv4_0;
	wire w_dff_B_oozMzcuF2_0;
	wire w_dff_B_6lvN3kSY0_0;
	wire w_dff_B_eNv3ff9E1_0;
	wire w_dff_B_AVJI1IGX1_0;
	wire w_dff_B_YhCP3RJR5_0;
	wire w_dff_A_qID4WNNU8_0;
	wire w_dff_A_2EyN7qET1_0;
	wire w_dff_A_7pCpBBN39_0;
	wire w_dff_A_frxi9byD9_0;
	wire w_dff_A_PIR7mxAp2_0;
	wire w_dff_A_Hz0GPvP20_0;
	wire w_dff_A_2nH0GZxE3_0;
	wire w_dff_B_dznslKDQ1_0;
	wire w_dff_B_bJrgIGLC4_0;
	wire w_dff_B_CDdEo12k0_0;
	wire w_dff_B_tPZA7zsE2_0;
	wire w_dff_B_xwxKc0KW7_0;
	wire w_dff_B_hhbfhIuz9_0;
	wire w_dff_A_6kLcD7zL4_0;
	wire w_dff_A_fyRQIDpf3_0;
	wire w_dff_A_M7r3Zzt85_0;
	wire w_dff_A_EvWzUAqm3_0;
	wire w_dff_A_iWtviGMz6_0;
	wire w_dff_A_N4bFkALy3_0;
	wire w_dff_A_51Bj5kf34_0;
	wire w_dff_A_pgXuwcnj2_0;
	wire w_dff_B_7VAQKTC95_0;
	wire w_dff_B_NdJPE4XP6_0;
	wire w_dff_B_NqLTbuqA7_0;
	wire w_dff_B_b2l72KXE0_0;
	wire w_dff_B_puZNNBTg3_0;
	wire w_dff_B_bqrvePcn8_0;
	wire w_dff_B_eR5ExF3L0_0;
	wire w_dff_B_q3KNssiL8_0;
	wire w_dff_B_HqQAKbo35_0;
	wire w_dff_A_hLumddvH0_0;
	wire w_dff_A_FcZ1TBoQ8_1;
	wire w_dff_A_Yt9IkgeX9_1;
	wire w_dff_A_A7acxXNr1_1;
	wire w_dff_A_VV06EGpu8_1;
	wire w_dff_A_A2z92gkD7_2;
	wire w_dff_A_dScTuOOL0_2;
	wire w_dff_A_trArhmMH5_0;
	wire w_dff_A_WX7dlkav2_0;
	wire w_dff_A_JFdvwC3B2_0;
	wire w_dff_A_j8iNbbck6_0;
	wire w_dff_A_DDdwYcRt3_1;
	wire w_dff_A_eilzWOxb9_1;
	wire w_dff_A_vkpMb6d29_1;
	wire w_dff_A_0Jc3Av869_1;
	wire w_dff_B_Ui3Wbu158_0;
	wire w_dff_B_iRjXtJ673_0;
	wire w_dff_B_vx82K3jn8_0;
	wire w_dff_B_0JvGJIpZ7_0;
	wire w_dff_B_r3oxkau82_0;
	wire w_dff_B_uAxXgHkX8_0;
	wire w_dff_B_zeKLxmuS2_0;
	wire w_dff_B_zUKjxpJd9_0;
	wire w_dff_B_gtojMpQM8_0;
	wire w_dff_B_xyY6mh8V6_0;
	wire w_dff_B_fUVttPHp4_0;
	wire w_dff_B_WuXpcJCp9_0;
	wire w_dff_A_ePj6LctY5_0;
	wire w_dff_A_erJPVHtM0_0;
	wire w_dff_A_mqkXTEC06_0;
	wire w_dff_A_QWQ1DtKV1_0;
	wire w_dff_A_6GtY2fWE3_0;
	wire w_dff_A_NBhpaSKd4_0;
	wire w_dff_B_u7wzn8vO0_0;
	wire w_dff_B_cVsXPlA27_0;
	wire w_dff_B_Ov8xtgzA0_0;
	wire w_dff_B_NJ97wETJ8_0;
	wire w_dff_B_BFfsGoj11_0;
	wire w_dff_B_VY4PXC7P1_0;
	wire w_dff_B_Nc3HHK5z7_0;
	wire w_dff_B_jdsmzO9M8_0;
	wire w_dff_B_1x5XozI66_0;
	wire w_dff_B_1JQcsZdo7_0;
	wire w_dff_B_HC3u8Yfs7_0;
	wire w_dff_A_AnsKQqqE0_0;
	wire w_dff_A_xLxi7wiR3_0;
	wire w_dff_A_UnNXMQmK4_0;
	wire w_dff_A_Lx5GNs0P4_0;
	wire w_dff_A_iJuM50qB6_1;
	wire w_dff_A_xd58JnAC1_1;
	wire w_dff_B_MFpA3PmB1_0;
	wire w_dff_B_h24csGr33_0;
	wire w_dff_B_7bd266Fo3_0;
	wire w_dff_B_8e3r9I3s4_0;
	wire w_dff_B_WIS3tm177_0;
	wire w_dff_B_edJd0PSN8_1;
	wire w_dff_B_PFUI3WGK3_1;
	wire w_dff_B_HBotJQtt4_1;
	wire w_dff_B_YCA7qrw44_1;
	wire w_dff_B_w6uc7q442_1;
	wire w_dff_A_eEVCHfL63_2;
	wire w_dff_A_TYG6RqQH6_2;
	wire w_dff_A_BOUseHkY4_2;
	wire w_dff_A_pQVO2DnM4_2;
	wire w_dff_B_7Ckizk8O9_3;
	wire w_dff_B_5L8eXvRX9_3;
	wire w_dff_A_SbDorVq62_1;
	wire w_dff_A_jFHnAu0m2_1;
	wire w_dff_A_zbrVtRZs8_2;
	wire w_dff_A_aGlFT7kQ1_2;
	wire w_dff_A_Xd5ZtYE87_2;
	wire w_dff_A_hufhjLzc9_2;
	wire w_dff_A_srgj378l7_0;
	wire w_dff_A_J3xX0R6e9_0;
	wire w_dff_A_63C5xwlS3_1;
	wire w_dff_B_0MxfRhmf0_0;
	wire w_dff_B_ZRRdUf0t4_0;
	wire w_dff_B_Ad1FpN0L5_0;
	wire w_dff_B_0MQe6lWW1_0;
	wire w_dff_B_oo6W34xP8_0;
	wire w_dff_B_Ja4dFN6o6_0;
	wire w_dff_B_7lV4R1GT0_0;
	wire w_dff_B_Ylw5k3Sn7_0;
	wire w_dff_B_rvqpqrK55_0;
	wire w_dff_B_iPMnBdR27_0;
	wire w_dff_B_DC1GyhgS8_0;
	wire w_dff_B_JCS4xw4h9_0;
	wire w_dff_B_0IB2FlBJ4_1;
	wire w_dff_B_h5U9nSjY9_1;
	wire w_dff_B_yZnwq2mo7_1;
	wire w_dff_B_p7z6dGUC4_1;
	wire w_dff_B_pBkP35yK1_1;
	wire w_dff_B_6brFvEQp9_1;
	wire w_dff_B_MKXPRiIA4_0;
	wire w_dff_B_MSBtCVXB7_0;
	wire w_dff_B_cX4bX2wC5_0;
	wire w_dff_B_u3e0XFcK3_0;
	wire w_dff_B_Zh2vVE8k0_0;
	wire w_dff_B_xAj5UnQL7_0;
	wire w_dff_B_IOXXKdlo9_0;
	wire w_dff_B_6pfDf5zb1_0;
	wire w_dff_B_xgbodGGy8_0;
	wire w_dff_B_r6MnnN211_0;
	wire w_dff_B_TIgTC8974_0;
	wire w_dff_B_PyZvP6qq3_0;
	wire w_dff_B_SsieJO0D3_0;
	wire w_dff_B_c9zkGq5W6_0;
	wire w_dff_B_qi0isgWG9_0;
	wire w_dff_B_mGPgZ6e00_0;
	wire w_dff_A_ZpDx0m9G7_0;
	wire w_dff_A_SdFcJZea0_0;
	wire w_dff_A_eb7nZeEv0_0;
	wire w_dff_A_S9FFe9xl5_0;
	wire w_dff_A_dqGPOkbq0_0;
	wire w_dff_A_DfsfmLgO2_0;
	wire w_dff_A_URXsBbbI2_0;
	wire w_dff_A_dxTqvqTy7_0;
	wire w_dff_A_AFd7f6Rv8_0;
	wire w_dff_A_lcN9nOVf8_0;
	wire w_dff_A_xdHQU8AK9_0;
	wire w_dff_A_wAknh2uT2_0;
	wire w_dff_A_W3xZVqvd4_0;
	wire w_dff_B_wozXgap33_2;
	wire w_dff_B_9FQwUB159_2;
	wire w_dff_B_06mJDRfX3_2;
	wire w_dff_B_eyaGwMpD4_1;
	wire w_dff_B_ABuABlaC9_0;
	wire w_dff_B_nZg96tG07_0;
	wire w_dff_B_KhItkqzk3_0;
	wire w_dff_A_Ie9xyNkC3_0;
	wire w_dff_A_xUU0Go5l4_0;
	wire w_dff_B_dS2amFQa1_1;
	wire w_dff_B_plUzJaFz2_1;
	wire w_dff_B_sllcrRqo5_1;
	wire w_dff_B_QTcJ8GD28_0;
	wire w_dff_B_Xa60deEF0_1;
	wire w_dff_A_F5GbhCwJ8_0;
	wire w_dff_A_k1WEk1cg5_0;
	wire w_dff_A_g2qvW19T6_0;
	wire w_dff_B_EotxGwAx0_0;
	wire w_dff_B_iTkLQcMp7_0;
	wire w_dff_B_rdP2cBpa7_0;
	wire w_dff_B_mHxqDbkI9_0;
	wire w_dff_B_dydXWkAG1_0;
	wire w_dff_B_cNIQDl6x0_0;
	wire w_dff_B_hC8IRBhE2_0;
	wire w_dff_B_wMdryTNs7_0;
	wire w_dff_B_tSRR7OHY0_0;
	wire w_dff_B_eQlnZ8Qu4_0;
	wire w_dff_B_HoKMSo2h1_0;
	wire w_dff_B_Cx6fu5b54_0;
	wire w_dff_B_Mhreckzp8_0;
	wire w_dff_B_vUORmcoW8_0;
	wire w_dff_B_s4r1RweA3_0;
	wire w_dff_B_q1B1dQ8c0_0;
	wire w_dff_B_ENRx4VdZ0_0;
	wire w_dff_B_8dfXrwUE8_0;
	wire w_dff_B_2pSBb1It8_0;
	wire w_dff_B_nn2TNj9B1_0;
	wire w_dff_B_XSuppEvn0_0;
	wire w_dff_B_LUp4y5Es7_0;
	wire w_dff_B_rIokX5MD0_0;
	wire w_dff_B_WJz1cW5s9_0;
	wire w_dff_B_M1ugVF4f8_0;
	wire w_dff_B_HJI0caO23_0;
	wire w_dff_B_cTn7yaGx3_0;
	wire w_dff_B_mfFp6fPu3_0;
	wire w_dff_B_DoSfxQP35_0;
	wire w_dff_B_74honPYO8_0;
	wire w_dff_B_x6LEa6qZ5_0;
	wire w_dff_B_1P5ecuwR7_0;
	wire w_dff_B_PvSL4RGA3_0;
	wire w_dff_B_b4hchHMT6_0;
	wire w_dff_B_jEu3uKf42_0;
	wire w_dff_B_N0FrtKqe5_0;
	wire w_dff_B_mS3eU0v09_0;
	wire w_dff_B_JS06cY6x5_0;
	wire w_dff_B_00goqtmS8_0;
	wire w_dff_B_3SBlXBzr3_0;
	wire w_dff_B_cMs4zbZn3_0;
	wire w_dff_B_n1GR9eCH5_0;
	wire w_dff_B_QRYJSOMe6_0;
	wire w_dff_B_5ktwBSEr4_0;
	wire w_dff_B_R2YyRbre9_0;
	wire w_dff_B_0PBvX6cm9_0;
	wire w_dff_B_dKlhZPq20_0;
	wire w_dff_B_1Us2ToPD9_0;
	wire w_dff_B_LH6IW6O59_0;
	wire w_dff_B_QDtKQf1m5_0;
	wire w_dff_B_C9N0WaPe6_0;
	wire w_dff_B_0snA5S6R4_0;
	wire w_dff_B_fayqID8R3_0;
	wire w_dff_B_RM4lGBpA6_0;
	wire w_dff_B_2YJFvSrb2_0;
	wire w_dff_B_Bbhvj9oR7_0;
	wire w_dff_B_gppSaH1L6_0;
	wire w_dff_B_migT0Gto1_0;
	wire w_dff_B_nMECjpHA2_0;
	wire w_dff_B_0DyUbfF35_0;
	wire w_dff_B_c7B0cfh38_0;
	wire w_dff_B_fqtFCQS57_0;
	wire w_dff_B_QXjM2iX20_0;
	wire w_dff_B_sQDB2RRH4_0;
	wire w_dff_B_HLbwSYic4_0;
	wire w_dff_B_AEJFMYQM6_0;
	wire w_dff_A_5qNoMRjg8_2;
	wire w_dff_B_CNQBkg7b9_0;
	wire w_dff_B_vc34ktVE2_0;
	wire w_dff_B_KRdhPSbg3_0;
	wire w_dff_B_TtdLE9hd2_0;
	wire w_dff_B_ruwOShWD6_0;
	wire w_dff_B_cyu3NbDF3_0;
	wire w_dff_B_FUk0zazF8_0;
	wire w_dff_B_T2qaG3YU5_0;
	wire w_dff_B_exC4SqlK1_0;
	wire w_dff_B_VzWR4oNC5_0;
	wire w_dff_B_no18nUS60_0;
	wire w_dff_B_RalU1xJW2_0;
	wire w_dff_B_VrJ1q9iA0_0;
	wire w_dff_B_1n95tzUM9_0;
	wire w_dff_B_KgDYaSie1_0;
	wire w_dff_B_lwEbFgj60_0;
	wire w_dff_B_Gkg6xUWo8_0;
	wire w_dff_B_GqIl0CA70_0;
	wire w_dff_B_3joDtvDu4_0;
	wire w_dff_B_IUhWtjRK8_0;
	wire w_dff_B_hl0ZoUVV2_0;
	wire w_dff_B_aY2qJ7Uj7_0;
	wire w_dff_B_bG8jNRRN5_0;
	wire w_dff_B_BuaV49N24_0;
	wire w_dff_B_bQcKaRrB8_0;
	wire w_dff_B_6lcXngbE4_0;
	wire w_dff_B_2glnAwbx2_0;
	wire w_dff_B_DzuMuKFa3_0;
	wire w_dff_B_AppQ0ae82_0;
	wire w_dff_B_6vpdyqyI3_0;
	wire w_dff_B_q4CWaEu15_0;
	wire w_dff_B_YoO9hlOX4_0;
	wire w_dff_B_DTuPXmxO9_0;
	wire w_dff_B_igmCWPGS9_0;
	wire w_dff_B_ezbEN3bN9_0;
	wire w_dff_B_iXRED5V68_0;
	wire w_dff_B_zItBIIjr8_0;
	wire w_dff_B_nmIXI8LO8_0;
	wire w_dff_B_pN6pqK9c2_0;
	wire w_dff_B_ufYIeoxd5_0;
	wire w_dff_B_QgVjl2Fm4_0;
	wire w_dff_B_AT4Ksb5E8_0;
	wire w_dff_B_gQBlGxro9_0;
	wire w_dff_B_bvJjKRG98_0;
	wire w_dff_B_pPT8A5wd8_0;
	wire w_dff_B_6GmiaF7s2_0;
	wire w_dff_B_E8rqHHnu5_0;
	wire w_dff_A_gYn5Hg3Q0_2;
	wire w_dff_B_iNXZlW3r2_0;
	wire w_dff_B_3y4FPi4V0_0;
	wire w_dff_B_PXcxPdDC5_0;
	wire w_dff_B_viHkD6KI0_0;
	wire w_dff_B_1S0oTDmG0_0;
	wire w_dff_B_jAVwv1X53_0;
	wire w_dff_B_d1yc9kdY1_0;
	wire w_dff_B_GCeIe2qI6_0;
	wire w_dff_B_IeY6iOT53_0;
	wire w_dff_B_u8gcdKr60_0;
	wire w_dff_B_kraurtIm3_0;
	wire w_dff_B_LWL3Bvv69_0;
	wire w_dff_B_wucsWPP73_0;
	wire w_dff_B_QrDz30uT0_0;
	wire w_dff_B_Qel3kc1U0_0;
	wire w_dff_B_LuOho6Yf9_0;
	wire w_dff_B_rA7zrRTu0_0;
	wire w_dff_B_HqvYioco9_0;
	wire w_dff_B_BVNuGsYc6_0;
	wire w_dff_B_DwTJcZbn1_0;
	wire w_dff_B_vHm2o6g43_0;
	wire w_dff_B_cHcW2Ou94_0;
	wire w_dff_B_2Mh2Rxch6_0;
	wire w_dff_B_Qbcn8qdw5_0;
	wire w_dff_B_PECfEeY57_0;
	wire w_dff_B_LZ01Pdfs7_0;
	wire w_dff_B_cgEPQjgE8_0;
	wire w_dff_B_nACt00vD2_0;
	wire w_dff_B_Io3g9NpZ5_0;
	wire w_dff_B_ivEV8khi6_0;
	wire w_dff_A_FNWn3Sj62_0;
	wire w_dff_A_ijzbJFWI3_0;
	wire w_dff_A_tq1U0GGZ5_0;
	wire w_dff_A_eaCfkIxx1_0;
	wire w_dff_A_aTLt1TvC9_0;
	wire w_dff_A_gnvf12y66_1;
	wire w_dff_B_fIhC1bEs2_0;
	wire w_dff_B_55U8fgP86_0;
	wire w_dff_B_aFEG09Le2_0;
	wire w_dff_B_pwyNGTQH1_0;
	wire w_dff_B_YEozEZos9_0;
	wire w_dff_B_05XECJyc3_0;
	wire w_dff_B_o7snKGUJ2_0;
	wire w_dff_B_TqTnbU8u1_0;
	wire w_dff_B_gMtFwqZE5_0;
	wire w_dff_B_UMhhWcBC5_0;
	wire w_dff_B_tzW2bO0a6_0;
	wire w_dff_B_X6DAxqdc9_0;
	wire w_dff_B_QQPVuDjs5_0;
	wire w_dff_B_0UfmfBky0_0;
	wire w_dff_B_AkQAFKTD6_0;
	wire w_dff_B_7cxBKTql8_0;
	wire w_dff_B_kPihtcfq0_0;
	wire w_dff_B_MJjWQueo0_0;
	wire w_dff_B_7gBuS4RL1_0;
	wire w_dff_B_nXjjKyHT1_0;
	wire w_dff_B_uZHh1tCw2_0;
	wire w_dff_B_fNoYMSYB2_0;
	wire w_dff_B_tNelqQ8X3_0;
	wire w_dff_B_P5L4WvUp8_0;
	wire w_dff_B_U6ciIMBv3_0;
	wire w_dff_B_evhXXUnD4_0;
	wire w_dff_B_ZQzU5vwe6_0;
	wire w_dff_B_k97cFn8n1_0;
	wire w_dff_B_QzoUBXs07_0;
	wire w_dff_B_rCYqDyRv0_0;
	wire w_dff_B_uh6p67i63_0;
	wire w_dff_B_yNQ5VDmC3_0;
	wire w_dff_A_cDTlSNpc6_0;
	wire w_dff_A_FloPqlkm3_1;
	wire w_dff_B_zBPvyyCS1_0;
	wire w_dff_B_jlFY93gi6_0;
	wire w_dff_B_k0rNrJ1c2_0;
	wire w_dff_B_4TKULP6y5_0;
	wire w_dff_B_2WrTKrlo8_0;
	wire w_dff_B_kl7zVGTp8_0;
	wire w_dff_B_YQ8XrtVg8_0;
	wire w_dff_B_gjucRhre0_0;
	wire w_dff_B_8J3MSDqz3_0;
	wire w_dff_B_aTGJZAjK2_0;
	wire w_dff_B_nhHj1Imt5_0;
	wire w_dff_B_JvpRnzoU2_0;
	wire w_dff_B_4dMPYloV4_0;
	wire w_dff_B_U5aV58BB3_0;
	wire w_dff_B_p4k3zeD80_0;
	wire w_dff_B_m67jEMao4_0;
	wire w_dff_B_2MPKNbl66_0;
	wire w_dff_A_qJgKLL8u9_0;
	wire w_dff_B_XJpeDObO3_0;
	wire w_dff_B_cL2PpUl82_0;
	wire w_dff_B_qb506v3Z0_0;
	wire w_dff_B_eRsD4t8b1_0;
	wire w_dff_B_jAwzG7nk6_0;
	wire w_dff_B_9rJZOjZh9_0;
	wire w_dff_B_n1AFnr4Q8_0;
	wire w_dff_B_uV5UYMyO3_0;
	wire w_dff_B_zeMpWe9z5_0;
	wire w_dff_B_vrDX8wic6_0;
	wire w_dff_B_r4UYfseN6_0;
	wire w_dff_B_PVzfH2SY9_0;
	wire w_dff_B_4AVRx9sL0_0;
	wire w_dff_B_BnKnPaLt8_0;
	wire w_dff_B_Mup6Tlwp7_0;
	wire w_dff_B_5SouL8NG9_0;
	wire w_dff_B_NYlbQWSk9_0;
	wire w_dff_B_NCa3gi3n0_0;
	wire w_dff_B_AI5BY90G9_0;
	wire w_dff_B_ZJieQwOd0_0;
	wire w_dff_B_kYWpZLDo2_0;
	wire w_dff_B_gjvM1czA5_0;
	wire w_dff_B_klsYbLLS0_0;
	wire w_dff_B_8UP3HyQ55_0;
	wire w_dff_B_8p6gElg63_0;
	wire w_dff_B_4P8f9Ny66_0;
	wire w_dff_B_jYHSEWlK0_0;
	wire w_dff_B_9CvpiysM6_0;
	wire w_dff_B_TsASmaCN8_0;
	wire w_dff_B_qE1TCVdM7_0;
	wire w_dff_B_6ISH0d4T1_0;
	wire w_dff_B_gGCs0xl34_0;
	wire w_dff_B_8chnMslM1_0;
	wire w_dff_B_zoiRCATK0_0;
	wire w_dff_B_2cVd1BrQ8_0;
	wire w_dff_B_plECz23Q3_0;
	wire w_dff_B_FwmdaOID9_0;
	wire w_dff_B_RKNmEgFa5_0;
	wire w_dff_B_EPlXEoKE7_0;
	wire w_dff_B_fyySlzZz8_0;
	wire w_dff_B_Gc2x3gDv4_0;
	wire w_dff_B_rv5iWwR70_0;
	wire w_dff_B_Q2jbklSd2_0;
	wire w_dff_B_FmE9Q68m8_0;
	wire w_dff_B_8UL0vcXR7_0;
	wire w_dff_B_GQE5kjLi0_0;
	wire w_dff_B_y0ZNfa0L1_0;
	wire w_dff_B_ilB1twKe4_0;
	wire w_dff_B_aB83t4lO5_0;
	wire w_dff_B_h7shaPp49_0;
	wire w_dff_A_bR1HbHEC2_1;
	wire w_dff_B_Md8tmAYG5_1;
	wire w_dff_B_JEw2LQZI4_1;
	wire w_dff_B_3XOpD3QT0_1;
	wire w_dff_B_regfi3Nb9_1;
	wire w_dff_B_ulL4W7kF5_1;
	wire w_dff_B_jtnHOeD41_1;
	wire w_dff_B_GMeH9Gjj8_1;
	wire w_dff_B_rDtJ97Wr4_1;
	wire w_dff_B_NchFnFQt8_1;
	wire w_dff_B_0Kif5Asu6_1;
	wire w_dff_B_ax1g88iu3_0;
	wire w_dff_B_K9lTEUfB1_0;
	wire w_dff_B_tgkvf8EM9_0;
	wire w_dff_B_73hCfHj40_0;
	wire w_dff_B_LhRFzZDx7_0;
	wire w_dff_B_8SbfsnlG3_0;
	wire w_dff_B_DMvDLERm5_0;
	wire w_dff_B_LfujWgXt4_0;
	wire w_dff_B_AfdXMorj6_0;
	wire w_dff_B_EMQrR9uk0_0;
	wire w_dff_B_AasOB3Pe0_0;
	wire w_dff_B_TBQjZteW8_0;
	wire w_dff_B_7f7NxTVv0_0;
	wire w_dff_B_sobignSw7_0;
	wire w_dff_B_TNP94jqn5_0;
	wire w_dff_B_7nkid9JF1_0;
	wire w_dff_B_msqNHctB7_0;
	wire w_dff_B_KVGJjC7d6_0;
	wire w_dff_B_07dPEegx8_0;
	wire w_dff_B_STWy7eZy0_0;
	wire w_dff_B_zDvnauw57_0;
	wire w_dff_B_M8A39Fs55_0;
	wire w_dff_B_ubpiBd992_0;
	wire w_dff_B_hQaZzNId4_0;
	wire w_dff_B_uZmqZvfC6_0;
	wire w_dff_B_b1F8kxF96_0;
	wire w_dff_B_7Ql7B85O2_0;
	wire w_dff_A_qKPaqswS4_0;
	wire w_dff_A_oWjaihkA6_1;
	wire w_dff_A_jocxXTXK8_0;
	wire w_dff_A_QabQwMds8_1;
	wire w_dff_A_GlLFU3d46_0;
	wire w_dff_A_GWW1Se4x3_0;
	wire w_dff_A_CwvoGdPP4_0;
	wire w_dff_A_DVMP496W0_0;
	wire w_dff_A_iq7Ngik62_0;
	wire w_dff_A_7iSlBHLh0_1;
	wire w_dff_A_FmSL0BLO9_1;
	wire w_dff_A_hGgPQXpz4_1;
	wire w_dff_A_W4dugbOG9_1;
	wire w_dff_A_PtzTfacB8_1;
	wire w_dff_A_UZnqtXha6_1;
	wire w_dff_B_ztWMvnCi3_0;
	wire w_dff_B_i9BkSOeO2_0;
	wire w_dff_B_K6lqkOYs0_0;
	wire w_dff_B_wtCgTdzf5_0;
	wire w_dff_B_x24JaxCH9_0;
	wire w_dff_B_c0flpRF76_0;
	wire w_dff_B_BEpWc7Ml2_0;
	wire w_dff_B_CL9tZ6D97_0;
	wire w_dff_B_yXl9WjRb8_0;
	wire w_dff_B_lAWTE3J57_0;
	wire w_dff_B_C9oS9cZS5_0;
	wire w_dff_B_7JEv4aTO8_0;
	wire w_dff_B_myWQJ2y58_0;
	wire w_dff_B_ailZ8pec2_0;
	wire w_dff_B_QcyVKDaF5_0;
	wire w_dff_B_UkYxzIAK4_0;
	wire w_dff_B_Ll5YcClR3_0;
	wire w_dff_B_1wGWBeyi0_0;
	wire w_dff_B_6102vNKn3_0;
	wire w_dff_B_javK3lxR8_0;
	wire w_dff_B_0OJJpXqw0_0;
	wire w_dff_B_WIsIyD9v8_0;
	wire w_dff_B_jsCtqBh03_0;
	wire w_dff_B_VnT4vukm2_0;
	wire w_dff_B_BNbcHZR40_0;
	wire w_dff_B_2z7KQv9V0_0;
	wire w_dff_B_WfaJa27F4_0;
	wire w_dff_B_80mx3hGy4_0;
	wire w_dff_B_3RTyat0o0_0;
	wire w_dff_B_E5a09JiM7_0;
	wire w_dff_B_b8gTI8kT6_0;
	wire w_dff_B_jdigdjsC9_0;
	wire w_dff_B_UKNgXBOI0_0;
	wire w_dff_B_6RQQT2QQ7_0;
	wire w_dff_A_9IVKEkEa9_0;
	wire w_dff_A_ajFVRjMK4_0;
	wire w_dff_A_gHNU9yhO6_0;
	wire w_dff_A_bhsedOfo1_0;
	wire w_dff_A_b5O4umPe7_0;
	wire w_dff_A_7VdwYuTi0_0;
	wire w_dff_A_mdUzwDUP4_0;
	wire w_dff_B_USQKzslP9_1;
	wire w_dff_B_KMgMnI7B3_1;
	wire w_dff_B_UnAVtBLJ5_1;
	wire w_dff_B_jXurijec5_1;
	wire w_dff_B_Ujp1Wrmx9_1;
	wire w_dff_B_LOmY5tsq4_1;
	wire w_dff_B_h9gUpSve0_1;
	wire w_dff_B_70ZbSBTX3_1;
	wire w_dff_B_HwQpfLCs0_1;
	wire w_dff_B_Wj5Eu4qw1_1;
	wire w_dff_B_kthcHHMA1_1;
	wire w_dff_B_hPwYu4Mw4_1;
	wire w_dff_B_aIS0yRux6_1;
	wire w_dff_B_RO05wpNx0_1;
	wire w_dff_B_v3kV7VdB5_1;
	wire w_dff_B_KP5xW9d20_1;
	wire w_dff_B_swx7ICbF7_1;
	wire w_dff_B_KIBYLFHW4_1;
	wire w_dff_B_EcgkE7Vz6_1;
	wire w_dff_B_liJr58Gv3_1;
	wire w_dff_B_tOD8Gnln8_1;
	wire w_dff_B_v8CpiGlj6_1;
	wire w_dff_B_AGoGd4HH0_1;
	wire w_dff_B_vu1PC1aU6_1;
	wire w_dff_B_d5C077gz9_1;
	wire w_dff_B_LeTPWCFM4_1;
	wire w_dff_B_fKpBDmCz7_1;
	wire w_dff_B_DeftKvjS2_1;
	wire w_dff_B_bn9wfamB6_1;
	wire w_dff_B_6EXBxlqf7_1;
	wire w_dff_B_6phi5lZD8_1;
	wire w_dff_B_04OXJUHx2_1;
	wire w_dff_B_PZtoP8qq6_1;
	wire w_dff_B_cMYxrKRs6_1;
	wire w_dff_B_rVQQE3yR9_1;
	wire w_dff_B_myWxgLJO3_1;
	wire w_dff_B_IWjoElcz7_1;
	wire w_dff_B_aFV8wzDx3_1;
	wire w_dff_B_15hlmeCz0_0;
	wire w_dff_B_Mqf5ubJI2_0;
	wire w_dff_B_mhDj21vY9_0;
	wire w_dff_B_gHqZyo5M7_0;
	wire w_dff_B_6e6B1n8h3_0;
	wire w_dff_B_0QVzKUlI6_0;
	wire w_dff_B_A4W80aMP3_0;
	wire w_dff_B_pUvIAmOp9_0;
	wire w_dff_B_RZc1oA6Y5_0;
	wire w_dff_B_HInz9TbG4_0;
	wire w_dff_B_HTo36Pef8_0;
	wire w_dff_B_TpL66Lr31_0;
	wire w_dff_B_ZyIjFXTA6_0;
	wire w_dff_B_qMi1Wg3H9_0;
	wire w_dff_B_sozDVgp64_0;
	wire w_dff_B_2ckhzU1K5_0;
	wire w_dff_B_qd0F33eQ0_0;
	wire w_dff_B_3LrkiBDe3_0;
	wire w_dff_B_vgKwEqZe7_0;
	wire w_dff_A_BK9DTSEo1_1;
	wire w_dff_A_XkEeD6U12_1;
	wire w_dff_A_550Je7HB8_1;
	wire w_dff_A_qSYZXzx47_1;
	wire w_dff_A_erIcdBdF1_1;
	wire w_dff_A_xoV0igcO0_1;
	wire w_dff_A_1ncj9mPS5_1;
	wire w_dff_A_IKqy2qAP1_1;
	wire w_dff_A_d56hPKNM7_1;
	wire w_dff_A_cjfv5gIw6_1;
	wire w_dff_A_bPPu9Tme4_1;
	wire w_dff_A_ymqvpjQT3_1;
	wire w_dff_A_A0CkILy93_1;
	wire w_dff_A_BXunqfwI6_1;
	wire w_dff_A_ywngHWxn3_2;
	wire w_dff_A_lhgl286T7_2;
	wire w_dff_A_j9Srvw5M9_2;
	wire w_dff_A_2j0g19Jd4_2;
	wire w_dff_A_KCpLv8PW7_2;
	wire w_dff_A_dxrN5TwR8_2;
	wire w_dff_A_DxVstlTq2_2;
	wire w_dff_A_NBfNvf6M3_2;
	wire w_dff_A_vZFeOSNe6_2;
	wire w_dff_A_o2tyTjap4_2;
	wire w_dff_A_URiRgjP36_1;
	wire w_dff_A_brXW6BiL6_1;
	wire w_dff_A_syESiIjk9_1;
	wire w_dff_A_7fLkCLQR7_1;
	wire w_dff_A_HqXYa5SV1_1;
	wire w_dff_A_kYvtkn6Q2_1;
	wire w_dff_A_fAEBuU884_1;
	wire w_dff_A_0gVQfX8d2_1;
	wire w_dff_A_wnyp9gVQ4_1;
	wire w_dff_A_aH6KF7Li9_1;
	wire w_dff_A_OTsvVIaB8_1;
	wire w_dff_A_GB2w0Nnn0_2;
	wire w_dff_B_r4tGmRXW1_3;
	wire w_dff_B_DQimDwlC9_3;
	wire w_dff_B_NUKKHghL4_3;
	wire w_dff_B_zkAyo6es1_3;
	wire w_dff_B_yBgG9BUT3_3;
	wire w_dff_B_YIZo3wIt3_3;
	wire w_dff_B_Cfafl5Uw9_0;
	wire w_dff_B_1D3tNEbH5_0;
	wire w_dff_B_T25pqIU90_0;
	wire w_dff_B_e3Z69bgo0_0;
	wire w_dff_B_mi6ossYj6_0;
	wire w_dff_B_M2eGyQQH9_0;
	wire w_dff_B_crkvjXU33_0;
	wire w_dff_B_PXaCXsGn0_0;
	wire w_dff_B_Q96U06dn2_0;
	wire w_dff_B_JwB8c2Id0_0;
	wire w_dff_B_vsJHQTFH3_0;
	wire w_dff_B_rTmzJXWY9_0;
	wire w_dff_B_uz2v2gJP5_0;
	wire w_dff_B_Ki1C5p8s9_0;
	wire w_dff_B_dtxE527h8_0;
	wire w_dff_B_Dq1ziY9a4_0;
	wire w_dff_B_WDVpWqM91_0;
	wire w_dff_B_U695gRXs2_0;
	wire w_dff_B_e5vsVdSQ9_0;
	wire w_dff_A_faJqbZCj9_1;
	wire w_dff_A_hDhfidel2_1;
	wire w_dff_A_cd3zl5239_1;
	wire w_dff_A_wT0kuPVf2_1;
	wire w_dff_A_DdZi7buT0_1;
	wire w_dff_A_Dt55PWry9_1;
	wire w_dff_A_CO8St1YS9_1;
	wire w_dff_A_m2S8yrAU7_1;
	wire w_dff_A_JbvicfCw8_1;
	wire w_dff_A_9UsFVfnC9_1;
	wire w_dff_A_z0St6chz6_1;
	wire w_dff_A_gXaqboLV4_1;
	wire w_dff_A_7D589fGb6_1;
	wire w_dff_A_z7biw8aO7_1;
	wire w_dff_A_kmdKYBFs7_2;
	wire w_dff_A_NLfBXjRI9_2;
	wire w_dff_A_6BhN392g9_2;
	wire w_dff_A_tT0ww60T9_2;
	wire w_dff_A_v1pKFrwK2_2;
	wire w_dff_A_GhHJEumA4_2;
	wire w_dff_A_HxdeZnw21_2;
	wire w_dff_A_s2EadMFx9_2;
	wire w_dff_A_AtRqkxFK9_2;
	wire w_dff_A_O4GArnQ14_2;
	wire w_dff_A_h7NcRlSa2_1;
	wire w_dff_A_0CI0HYfu6_1;
	wire w_dff_A_7qNmDIMF2_1;
	wire w_dff_A_lTT1lmQx8_1;
	wire w_dff_A_Lm2jK0k00_1;
	wire w_dff_A_k3Mg6Bdz5_1;
	wire w_dff_A_426JwAvx2_1;
	wire w_dff_A_tdIr1GZD7_1;
	wire w_dff_A_fW4zbuyv3_1;
	wire w_dff_A_2nYDDVP93_1;
	wire w_dff_A_0idNOgO82_1;
	wire w_dff_A_mxYrmpWq2_2;
	wire w_dff_B_yKeoj2Oi7_3;
	wire w_dff_B_rcgxDbXG3_3;
	wire w_dff_B_30fadAIL9_3;
	wire w_dff_B_4vRaUZrI7_3;
	wire w_dff_B_qIwBJaZA5_3;
	wire w_dff_B_nbEnGORg5_3;
	wire w_dff_B_Xoebksbe1_1;
	wire w_dff_B_mXHIPi7r6_0;
	wire w_dff_B_lOF0kPk27_0;
	wire w_dff_B_PyGoNv9p6_0;
	wire w_dff_B_ludczpeP3_0;
	wire w_dff_B_3OlqcsDz3_0;
	wire w_dff_B_jJrx93m36_0;
	wire w_dff_B_b1uaOjDS4_0;
	wire w_dff_B_N9payxge5_0;
	wire w_dff_B_wHRzwpWI8_0;
	wire w_dff_B_4tHvCdM24_0;
	wire w_dff_B_AwFToQub6_0;
	wire w_dff_B_Rud5IheJ3_0;
	wire w_dff_B_Tylp1GK25_0;
	wire w_dff_B_4oj8cpEW1_0;
	wire w_dff_B_VWeBcbz51_0;
	wire w_dff_B_KxkvSA1o5_0;
	wire w_dff_B_V9uOycli7_0;
	wire w_dff_B_bVZczMbx8_0;
	wire w_dff_B_8n3vo7RB0_1;
	wire w_dff_B_h88qhk292_1;
	wire w_dff_B_N3mal6mu1_1;
	wire w_dff_B_aucyYDED9_1;
	wire w_dff_B_7yJ48Wmp3_1;
	wire w_dff_B_pqxQBoJZ4_1;
	wire w_dff_B_dLr0mNqu5_1;
	wire w_dff_B_ImSWn67M3_1;
	wire w_dff_B_KU9aBWNF6_1;
	wire w_dff_B_n4c1XlKr5_1;
	wire w_dff_B_bRad8Ntl3_1;
	wire w_dff_B_sywqYdfQ3_1;
	wire w_dff_B_HQJVhmfY9_1;
	wire w_dff_B_MQAqoOmp5_1;
	wire w_dff_B_Po53HvDG2_1;
	wire w_dff_B_YY6E9Tr81_1;
	wire w_dff_B_IMCEMDY18_1;
	wire w_dff_B_auoXWo6O9_1;
	wire w_dff_B_e33LovgP0_1;
	wire w_dff_B_ddURQ7Dr9_1;
	wire w_dff_B_GksMrAHL7_0;
	wire w_dff_B_SKtUkjFX0_0;
	wire w_dff_B_lXl8u2807_0;
	wire w_dff_B_JlAfKRAv1_0;
	wire w_dff_B_VxsxfR1i8_0;
	wire w_dff_B_ZymxUA9Z4_0;
	wire w_dff_B_rTnONUwH8_0;
	wire w_dff_B_Og2fEFdx8_0;
	wire w_dff_B_5v2nRLVr1_0;
	wire w_dff_B_58IJzkPx7_0;
	wire w_dff_B_mfk3XKas0_0;
	wire w_dff_B_nqUp5bem5_0;
	wire w_dff_B_AkmkdL2U3_0;
	wire w_dff_B_0J3oHaDB2_0;
	wire w_dff_B_5GFmOFuN7_0;
	wire w_dff_B_8nt7m9RE2_0;
	wire w_dff_B_5WhggEDT5_0;
	wire w_dff_B_5W8CGx180_0;
	wire w_dff_B_zkO0tHSn5_1;
	wire w_dff_B_I25RDzZ94_1;
	wire w_dff_B_BXLNxTsJ5_1;
	wire w_dff_B_PdTixlrW5_1;
	wire w_dff_B_5EXA678H7_1;
	wire w_dff_B_lLdSiesg9_1;
	wire w_dff_B_lkYcCaAH7_1;
	wire w_dff_B_ZAdAPF8j4_1;
	wire w_dff_B_Q9bXY9iO6_1;
	wire w_dff_B_hIoZZVs60_1;
	wire w_dff_B_92wjE9lL0_1;
	wire w_dff_B_JC9ErbD70_1;
	wire w_dff_B_ZrC4OjzC0_1;
	wire w_dff_B_3XgyYXZy4_1;
	wire w_dff_B_bM6IEAfH0_1;
	wire w_dff_B_egznxpg66_1;
	wire w_dff_B_8iwuC1d94_1;
	wire w_dff_B_Jv6B9aF50_1;
	wire w_dff_B_bZbagBGo7_1;
	wire w_dff_B_sZtMb9X57_0;
	wire w_dff_B_MeOL8bvJ5_0;
	wire w_dff_B_s5lFu9w62_0;
	wire w_dff_B_1lp7X9HY6_0;
	wire w_dff_B_YZFR1aXT5_0;
	wire w_dff_B_pJbITUhM1_0;
	wire w_dff_B_ndNDPUJj3_0;
	wire w_dff_B_FnEFXOok1_0;
	wire w_dff_B_RLSgYVnb4_0;
	wire w_dff_B_7TivSpXc5_0;
	wire w_dff_B_98cSCAkM7_0;
	wire w_dff_B_QUkMZbLA4_0;
	wire w_dff_B_UymDJ8TM2_0;
	wire w_dff_B_8neHo7o57_0;
	wire w_dff_B_sVCac5ow6_0;
	wire w_dff_B_mKIAvnbD5_0;
	wire w_dff_B_aj220N9X9_0;
	wire w_dff_B_xBJkETM87_0;
	wire w_dff_B_turOlrt26_0;
	wire w_dff_B_6bZxOr787_1;
	wire w_dff_B_9siOO4ek5_1;
	wire w_dff_B_mOMU5UYN2_1;
	wire w_dff_B_yTRY5S2l2_1;
	wire w_dff_B_dhj9MhGd1_1;
	wire w_dff_B_VJgNpd3v5_1;
	wire w_dff_A_5N9tgYEO1_1;
	wire w_dff_B_5zaBbffg4_1;
	wire w_dff_B_GGZBohVy0_1;
	wire w_dff_B_pV08APgv4_1;
	wire w_dff_B_g1A5T19g6_1;
	wire w_dff_B_rMH6wThe5_1;
	wire w_dff_B_Wb2gv5YS1_1;
	wire w_dff_B_B963ehN05_1;
	wire w_dff_B_LtgTD4Ez4_1;
	wire w_dff_B_zRcmY1Ug2_1;
	wire w_dff_B_LLiJKrcD2_1;
	wire w_dff_B_jNf0BP9R3_0;
	wire w_dff_B_fKpEoIgw7_0;
	wire w_dff_A_nCygsGsv6_1;
	wire w_dff_A_9u0yrDq81_1;
	wire w_dff_A_e0btWtwj6_1;
	wire w_dff_B_wzRzGDvU7_0;
	wire w_dff_B_EeCOdrtz7_1;
	wire w_dff_B_fYc4TshO6_1;
	wire w_dff_B_qUs1wJ4M1_1;
	wire w_dff_B_iHtukHpL5_1;
	wire w_dff_B_fUbz4NVr5_1;
	wire w_dff_B_qbgis4aG8_1;
	wire w_dff_B_5e9lLEwP3_1;
	wire w_dff_B_jkjH0v9K4_1;
	wire w_dff_B_zScbqlEf1_1;
	wire w_dff_B_Yymp456X4_1;
	wire w_dff_B_l9yYNM3y7_1;
	wire w_dff_B_02WrUaWC2_1;
	wire w_dff_B_LzQJJeCb3_1;
	wire w_dff_B_fm3FDxps1_1;
	wire w_dff_B_IJO3eluU6_1;
	wire w_dff_B_8XP8jZ1L9_1;
	wire w_dff_B_2Lkh4R635_1;
	wire w_dff_B_VoHCHtBi5_0;
	wire w_dff_A_RzFfuChi6_0;
	wire w_dff_A_H3ScOOKu0_0;
	wire w_dff_A_x8XgfZtr4_0;
	wire w_dff_B_Zfy0bBXR1_1;
	wire w_dff_A_6A7OUpET3_1;
	wire w_dff_A_5DQrxhTw1_1;
	wire w_dff_A_mIDnUMUY1_1;
	wire w_dff_A_E4Rsaesr7_1;
	wire w_dff_A_f8jnsMYH5_1;
	wire w_dff_A_bsUiUq3R8_1;
	wire w_dff_A_yiHJB6z70_2;
	wire w_dff_A_A0PVhH983_2;
	wire w_dff_B_kpcoNTEd7_2;
	wire w_dff_B_tXUJF08v1_2;
	wire w_dff_B_6eRvWGTO2_2;
	wire w_dff_B_lWDXr2Zo0_2;
	wire w_dff_B_Xv9pZukw0_2;
	wire w_dff_B_AtfNQjRJ0_2;
	wire w_dff_B_mechHiC69_2;
	wire w_dff_B_6D9HwHrJ2_2;
	wire w_dff_B_hcZWEMPy7_2;
	wire w_dff_A_Txqjbibg9_1;
	wire w_dff_A_Zzfl8d7n6_1;
	wire w_dff_A_fVfHPFEl1_1;
	wire w_dff_A_oTy64uHq9_1;
	wire w_dff_A_1TEmmUns4_1;
	wire w_dff_A_4Pe0hfd69_1;
	wire w_dff_A_0pVFSIYZ0_1;
	wire w_dff_A_QVo1U4UG6_1;
	wire w_dff_A_PHILE3gA2_1;
	wire w_dff_A_rTKPoJwV1_1;
	wire w_dff_A_fwg9U8jF2_1;
	wire w_dff_A_ylRM2eMt7_1;
	wire w_dff_A_mtdFSZKM7_1;
	wire w_dff_A_VzvL9tk17_1;
	wire w_dff_A_6l12njUS4_2;
	wire w_dff_A_wDmslZSH7_0;
	wire w_dff_A_fBeSBzmf9_0;
	wire w_dff_A_gRmMcFN92_0;
	wire w_dff_A_NzKBFKV83_0;
	wire w_dff_A_naENVEYz1_0;
	wire w_dff_A_QC4rYQS22_0;
	wire w_dff_A_715MGgWo7_0;
	wire w_dff_A_dNhsUvwf9_0;
	wire w_dff_A_TqAmVVtt4_0;
	wire w_dff_A_7YHxvuJ43_0;
	wire w_dff_A_w4ia18uG3_0;
	wire w_dff_A_sXYZBzkT3_0;
	wire w_dff_B_z6nn5o6q1_1;
	wire w_dff_B_ZxZfcKbg4_0;
	wire w_dff_B_d9hPlEia5_0;
	wire w_dff_B_1mqFA4Qc4_0;
	wire w_dff_B_r0NRFXqF2_0;
	wire w_dff_B_gZekIbB44_0;
	wire w_dff_B_jwnaOYvi6_0;
	wire w_dff_B_r2Z0Yv1L6_0;
	wire w_dff_B_jPkWfscm1_0;
	wire w_dff_B_Gpxjw03t9_0;
	wire w_dff_A_o6Ok0uWN0_0;
	wire w_dff_A_g1iU1Asj6_0;
	wire w_dff_A_yhM1GGPX8_0;
	wire w_dff_A_W3AJjpbZ6_1;
	wire w_dff_A_PrVgnCwx1_1;
	wire w_dff_A_a62VI9RO2_1;
	wire w_dff_A_QCo5rrFG2_0;
	wire w_dff_A_41iniY6v3_2;
	wire w_dff_A_Gxmw2GQZ2_0;
	wire w_dff_B_LnF8sMbi2_1;
	wire w_dff_B_BIiJJkwU9_1;
	wire w_dff_B_xyxYBYEl9_1;
	wire w_dff_B_VreztqLC8_1;
	wire w_dff_B_YAseiAYS2_1;
	wire w_dff_B_qNVll6yt7_1;
	wire w_dff_B_Tc99gfYc0_1;
	wire w_dff_B_BqxP2BEn1_1;
	wire w_dff_B_OzkxPolt3_1;
	wire w_dff_B_8rssqo1N2_1;
	wire w_dff_B_xpRPAu6s1_1;
	wire w_dff_B_eHJf75vv5_1;
	wire w_dff_B_GfqzFmgf1_1;
	wire w_dff_B_Oe513zkN7_1;
	wire w_dff_B_Q7B98Heb2_1;
	wire w_dff_A_OEnd0fHr7_0;
	wire w_dff_A_uK0Xd9Vt0_0;
	wire w_dff_A_GyvaTXiS2_1;
	wire w_dff_A_GqrbQujp2_1;
	wire w_dff_A_c9idzpQo8_1;
	wire w_dff_A_QMAibGF28_1;
	wire w_dff_A_YxPcOlQR0_1;
	wire w_dff_A_4MaBBqXA9_1;
	wire w_dff_A_ezdLpXPg4_1;
	wire w_dff_A_Ufs7lqJq2_1;
	wire w_dff_A_nsxbk5Go9_1;
	wire w_dff_A_5xlRuwxL9_2;
	wire w_dff_A_o3ibLdIi1_2;
	wire w_dff_A_NNKvvsPr7_0;
	wire w_dff_A_KSXrmRRr3_0;
	wire w_dff_A_HJLLE2YR5_0;
	wire w_dff_B_gz6R6oVC8_2;
	wire w_dff_B_tExL2pd21_2;
	wire w_dff_B_s79O3IVw3_2;
	wire w_dff_B_pTRwyhQr3_2;
	wire w_dff_B_acY2Vds50_2;
	wire w_dff_B_kQjNf0Ez3_2;
	wire w_dff_B_vIR1s6d80_2;
	wire w_dff_B_FjLdEi1b4_2;
	wire w_dff_B_0ZaLwdyt5_2;
	wire w_dff_B_nVuEXnZw3_2;
	wire w_dff_B_8utvpYlG1_2;
	wire w_dff_B_U0al0I6L3_2;
	wire w_dff_B_hdSSqI6c3_2;
	wire w_dff_B_gkIOj6l26_2;
	wire w_dff_B_Iwg9H4X03_2;
	wire w_dff_B_f2i64VtA7_2;
	wire w_dff_B_71eaoaDk3_2;
	wire w_dff_B_5t5qpv1I5_2;
	wire w_dff_B_vHwQew9u1_2;
	wire w_dff_B_wzPkVA5E0_2;
	wire w_dff_B_BTqCJAI29_2;
	wire w_dff_B_aSJdigHj0_2;
	wire w_dff_B_yotyiVqZ9_2;
	wire w_dff_B_eJRdOaJC4_2;
	wire w_dff_A_L8i6nSmj8_1;
	wire w_dff_A_nC8NIUml7_0;
	wire w_dff_A_BY1mYJK41_0;
	wire w_dff_A_b73VTaDF7_0;
	wire w_dff_A_UyijAhBH0_0;
	wire w_dff_A_sNYrpXW42_0;
	wire w_dff_A_zWDWptYv9_0;
	wire w_dff_A_8R0OgeLw1_0;
	wire w_dff_A_1HEAJ2Rf5_0;
	wire w_dff_A_0HRkchec2_0;
	wire w_dff_A_RyHajLb78_0;
	wire w_dff_A_iePnse2A4_0;
	wire w_dff_A_w85hnXY70_0;
	wire w_dff_A_bkZH3Xcz7_0;
	wire w_dff_A_rz6xaLAj5_0;
	wire w_dff_A_OGwDk4DX4_0;
	wire w_dff_A_ixQCzRUg9_0;
	wire w_dff_A_LhOp4ex32_0;
	wire w_dff_A_32OQkVZa1_0;
	wire w_dff_A_G9K6tBZ61_0;
	wire w_dff_A_D4IT5YDC8_0;
	wire w_dff_A_reQRNsTe7_0;
	wire w_dff_A_tehqSbla9_0;
	wire w_dff_A_2UR8aYlw4_0;
	wire w_dff_A_SctOiIYD5_0;
	wire w_dff_A_iAL19hqC7_0;
	wire w_dff_A_xzFbqVFy4_1;
	wire w_dff_A_mdeFull68_0;
	wire w_dff_A_qpTcncIA8_0;
	wire w_dff_A_G9ZYLKqt8_0;
	wire w_dff_A_VBu5CG410_0;
	wire w_dff_A_9u2UjhkD7_0;
	wire w_dff_A_r8IzaxXH4_0;
	wire w_dff_A_HASDwZ0E1_0;
	wire w_dff_A_GB8Aja8V0_0;
	wire w_dff_A_QMsyAdqG1_0;
	wire w_dff_A_Z9WzIFaZ6_0;
	wire w_dff_A_93yMKHsq2_0;
	wire w_dff_A_chYaKOcK7_0;
	wire w_dff_A_HCo5tBmy8_0;
	wire w_dff_A_mWZCSMJ39_0;
	wire w_dff_A_9Qa2rzvi7_0;
	wire w_dff_A_mogR2yJN6_0;
	wire w_dff_A_G3WcGPul8_0;
	wire w_dff_A_FqgHiXhR5_0;
	wire w_dff_A_WlktV3d53_0;
	wire w_dff_A_s3zZi4AZ3_0;
	wire w_dff_A_GmDXqLHv5_0;
	wire w_dff_A_xpQ2pYsZ3_0;
	wire w_dff_A_O0a02aXr0_0;
	wire w_dff_A_lotCgd6q8_0;
	wire w_dff_A_kNLoaKsm3_0;
	wire w_dff_A_MwhKPAJt6_1;
	wire w_dff_A_8DSwKiPK5_0;
	wire w_dff_A_YDBqf7dz2_0;
	wire w_dff_A_3OkWTd0k6_0;
	wire w_dff_A_9GEjySGP9_0;
	wire w_dff_A_6L2J0ckt4_0;
	wire w_dff_A_d7O9XkWb9_0;
	wire w_dff_A_YkeI5BVx7_0;
	wire w_dff_A_bEXsGrKu1_0;
	wire w_dff_A_6sDJd9sI2_0;
	wire w_dff_A_0DwipA3O4_0;
	wire w_dff_A_zYuQYnx05_0;
	wire w_dff_A_aT5uoKTe2_0;
	wire w_dff_A_HovGehEh4_0;
	wire w_dff_A_2awL2d8H3_0;
	wire w_dff_A_B2zJ4YEZ0_0;
	wire w_dff_A_uvOoS5l04_0;
	wire w_dff_A_KjUKImIS3_0;
	wire w_dff_A_WHok27LG9_0;
	wire w_dff_A_OL4y1KYB5_0;
	wire w_dff_A_wFIdRpWy9_0;
	wire w_dff_A_EAmQGzpo5_0;
	wire w_dff_A_OAfYR3df3_0;
	wire w_dff_A_iFBZSlSi9_0;
	wire w_dff_A_oThtbLix2_0;
	wire w_dff_A_umplgO0A1_0;
	wire w_dff_A_qxuufKM28_1;
	wire w_dff_A_B7dVYRKr2_0;
	wire w_dff_A_tnOYKNRe1_0;
	wire w_dff_A_eKUyWfJJ8_0;
	wire w_dff_A_ilHvDOjW2_0;
	wire w_dff_A_3a6uZq8s0_0;
	wire w_dff_A_rFnpqvyo8_0;
	wire w_dff_A_v5QSkWTu4_0;
	wire w_dff_A_YnAczJ0q1_0;
	wire w_dff_A_XpSlgmas0_0;
	wire w_dff_A_adib1pqi5_0;
	wire w_dff_A_Y5NX0GwP9_0;
	wire w_dff_A_bS02rXEU1_0;
	wire w_dff_A_ozBu0WPf3_0;
	wire w_dff_A_0LK8BBPg1_0;
	wire w_dff_A_r4RY1TO81_0;
	wire w_dff_A_yEwhhbqh6_0;
	wire w_dff_A_x9vz4WlQ1_0;
	wire w_dff_A_AaxuenLJ6_0;
	wire w_dff_A_NtormZjw0_0;
	wire w_dff_A_fiIeZXGv0_0;
	wire w_dff_A_sC1YFJpX2_0;
	wire w_dff_A_Vyb4M1o19_0;
	wire w_dff_A_gQpL75o37_0;
	wire w_dff_A_JtZ3ZgxX8_0;
	wire w_dff_A_bSb3TJii9_1;
	wire w_dff_A_o3ZVTnGo1_0;
	wire w_dff_A_Ob7uzYGM3_0;
	wire w_dff_A_Kyo6X4tZ2_0;
	wire w_dff_A_XqtPLVJt3_0;
	wire w_dff_A_vOj6XkBM0_0;
	wire w_dff_A_SY02V9pO7_0;
	wire w_dff_A_0309OFbp7_0;
	wire w_dff_A_2sBjf7r18_0;
	wire w_dff_A_62MvLBeq7_0;
	wire w_dff_A_eEo3fZPx2_0;
	wire w_dff_A_BczQ3AWs6_0;
	wire w_dff_A_iw4eHbsx8_0;
	wire w_dff_A_3zl7JXeM4_0;
	wire w_dff_A_DZSzWZbQ3_0;
	wire w_dff_A_VBEpL0Q74_0;
	wire w_dff_A_ShwZ0unR9_0;
	wire w_dff_A_zRVTRC1R6_0;
	wire w_dff_A_Epg5lDUC8_0;
	wire w_dff_A_ka3hEXUS8_0;
	wire w_dff_A_ozr4ErDd0_0;
	wire w_dff_A_A3ImSNKF3_0;
	wire w_dff_A_eLft2fKP0_0;
	wire w_dff_A_Utc5zoXZ0_0;
	wire w_dff_A_KWTBCgkk7_0;
	wire w_dff_A_1FoVNhmo2_1;
	wire w_dff_A_EqblviLa4_0;
	wire w_dff_A_x4dS4KNm3_0;
	wire w_dff_A_hxWnKqoD4_0;
	wire w_dff_A_Wk4Ua9No1_0;
	wire w_dff_A_IfJBLCrn5_0;
	wire w_dff_A_Hi1DSY4q7_0;
	wire w_dff_A_VN4bPgD34_0;
	wire w_dff_A_QFRhVDnB1_0;
	wire w_dff_A_a6f3iM4m2_0;
	wire w_dff_A_zM1NMrti9_0;
	wire w_dff_A_JknuqsQ69_0;
	wire w_dff_A_LsD8gn9B6_0;
	wire w_dff_A_gYXmfC4y0_0;
	wire w_dff_A_FYUnYbAd7_0;
	wire w_dff_A_xXXvQaTo4_0;
	wire w_dff_A_jmcsJKy64_0;
	wire w_dff_A_UzYq3r1H0_0;
	wire w_dff_A_LnHxCXJN1_0;
	wire w_dff_A_Y4Qr51QY6_0;
	wire w_dff_A_BjHHcAUc2_0;
	wire w_dff_A_eEV9Abv68_0;
	wire w_dff_A_Y17b1LG46_0;
	wire w_dff_A_ItoGbDu54_0;
	wire w_dff_A_FSHB2BVx2_0;
	wire w_dff_A_5HCiJFb58_1;
	wire w_dff_A_xrcT79jh6_0;
	wire w_dff_A_cSNY9F118_0;
	wire w_dff_A_tZ4QfeYo2_0;
	wire w_dff_A_xMth6Vab5_0;
	wire w_dff_A_k72Yj2Ya3_0;
	wire w_dff_A_YBrByc0o2_0;
	wire w_dff_A_zEBEAsmK3_0;
	wire w_dff_A_grbhomvc9_0;
	wire w_dff_A_qYBpGPHq2_0;
	wire w_dff_A_ucFCkGzM2_0;
	wire w_dff_A_hakhRnzV9_0;
	wire w_dff_A_n0IMI8yt8_0;
	wire w_dff_A_QXgVB1VL2_0;
	wire w_dff_A_dKeolqRn3_0;
	wire w_dff_A_3I87KtaD1_0;
	wire w_dff_A_MqNN865V1_0;
	wire w_dff_A_ty9njzzq6_0;
	wire w_dff_A_jYMPg27r9_0;
	wire w_dff_A_FxqWgxyw8_0;
	wire w_dff_A_YJvCoOxH3_0;
	wire w_dff_A_HDhPVR4P6_0;
	wire w_dff_A_ue5fVz9Y1_0;
	wire w_dff_A_hx8webFW0_0;
	wire w_dff_A_vStQhvT93_0;
	wire w_dff_A_aQkG8FTE9_1;
	wire w_dff_A_yECJxp9H1_0;
	wire w_dff_A_H1xXD0rB6_0;
	wire w_dff_A_zYHP0WZh3_0;
	wire w_dff_A_uenPKdjy2_0;
	wire w_dff_A_F42ENXhK8_0;
	wire w_dff_A_CWHT7mns5_0;
	wire w_dff_A_wKd1hncY2_0;
	wire w_dff_A_0cuR7wp02_0;
	wire w_dff_A_pyZpVygc5_0;
	wire w_dff_A_DfJK21kO9_0;
	wire w_dff_A_vVjsGcHC3_0;
	wire w_dff_A_Mq5LqRSY2_0;
	wire w_dff_A_r7wCzyxi5_0;
	wire w_dff_A_arbtq3m29_0;
	wire w_dff_A_vXx1Mv7l5_0;
	wire w_dff_A_oJshd60A7_0;
	wire w_dff_A_wxZOrlqw9_0;
	wire w_dff_A_Tc8TjFDV1_0;
	wire w_dff_A_9XjoMj7o2_0;
	wire w_dff_A_dpQPqRNB4_0;
	wire w_dff_A_r9dDJkmY5_0;
	wire w_dff_A_RioAGGVx9_0;
	wire w_dff_A_siWcFYow7_0;
	wire w_dff_A_ucmJ6k8S5_0;
	wire w_dff_A_gr7tdRmi6_1;
	wire w_dff_A_hBn5ttdH3_0;
	wire w_dff_A_gDl5Fn464_0;
	wire w_dff_A_Ve6aCRAt1_0;
	wire w_dff_A_aWUn4EZ20_0;
	wire w_dff_A_NLzJa5X31_0;
	wire w_dff_A_jVfIlE819_0;
	wire w_dff_A_hQJdSSje8_0;
	wire w_dff_A_ONpbsbqp3_0;
	wire w_dff_A_swmwDC7v6_0;
	wire w_dff_A_9xAhxXP04_0;
	wire w_dff_A_MqvQPcUc6_0;
	wire w_dff_A_gI361zfA6_0;
	wire w_dff_A_IapgDGrg0_0;
	wire w_dff_A_81dyt1Uy2_0;
	wire w_dff_A_RRZIrERw8_0;
	wire w_dff_A_oZToYoLD5_0;
	wire w_dff_A_a78YLMOZ7_0;
	wire w_dff_A_WQaws6Ie6_0;
	wire w_dff_A_OcsYoPst5_0;
	wire w_dff_A_rtFC0nVv9_0;
	wire w_dff_A_LGPgYbvx0_0;
	wire w_dff_A_nnq9LSC41_0;
	wire w_dff_A_4etVxjX29_0;
	wire w_dff_A_oVV3ENCY3_0;
	wire w_dff_A_OUjptODI7_1;
	wire w_dff_A_plwWFb4D4_0;
	wire w_dff_A_b7aZoJ4a6_0;
	wire w_dff_A_URFVMIDc3_0;
	wire w_dff_A_McK0uXlW5_0;
	wire w_dff_A_i5qE0GQn1_0;
	wire w_dff_A_POdY9Rtj7_0;
	wire w_dff_A_6dNJKmMS2_0;
	wire w_dff_A_Yln3uv1E0_0;
	wire w_dff_A_4bv8kuBe7_0;
	wire w_dff_A_masqWA0e1_0;
	wire w_dff_A_nMyXoepL7_0;
	wire w_dff_A_NvlA8NfG9_0;
	wire w_dff_A_dqIuYJhf9_0;
	wire w_dff_A_d8sPpaa22_0;
	wire w_dff_A_pCTziFrW5_0;
	wire w_dff_A_NddNnJEM5_0;
	wire w_dff_A_lmun7lGa6_0;
	wire w_dff_A_gfvOh1a45_0;
	wire w_dff_A_qUjReKbK7_0;
	wire w_dff_A_oO653SGZ4_0;
	wire w_dff_A_N4EMP4Qv4_0;
	wire w_dff_A_16pNIE2M8_0;
	wire w_dff_A_A1ul20vT2_0;
	wire w_dff_A_IttKCy8j5_0;
	wire w_dff_A_FJjvtOnm3_1;
	wire w_dff_A_YSYzDgDs9_0;
	wire w_dff_A_xMWjtSNp1_0;
	wire w_dff_A_yKytuZkK8_0;
	wire w_dff_A_chnn2FVy3_0;
	wire w_dff_A_hSLVk3pN7_0;
	wire w_dff_A_KvJrlhri3_0;
	wire w_dff_A_46m0Oqh99_0;
	wire w_dff_A_y7Mq608C2_0;
	wire w_dff_A_xVLCQ4Ec3_0;
	wire w_dff_A_fyj0MEvt2_0;
	wire w_dff_A_ysNRlxUY1_0;
	wire w_dff_A_zsvlQMd40_0;
	wire w_dff_A_vy9FQOrt1_0;
	wire w_dff_A_pzE5bXhX1_0;
	wire w_dff_A_hZRFcWxc3_0;
	wire w_dff_A_24ox9GgO9_0;
	wire w_dff_A_S2ARY1D45_0;
	wire w_dff_A_rovhe0RP3_0;
	wire w_dff_A_aRQobSYC4_0;
	wire w_dff_A_zTDctRW94_0;
	wire w_dff_A_1ZrL74WM5_0;
	wire w_dff_A_lwp0zlzh8_0;
	wire w_dff_A_y6xwCR5I3_0;
	wire w_dff_A_NhO4xXpN6_0;
	wire w_dff_A_HPCQADGE6_1;
	wire w_dff_A_aLCa9vOG5_0;
	wire w_dff_A_NDprfOMW5_0;
	wire w_dff_A_ESlHrX7O2_0;
	wire w_dff_A_8yHfk8Mw6_0;
	wire w_dff_A_QKp91s2h2_0;
	wire w_dff_A_L0ThTLBV3_0;
	wire w_dff_A_G7Zt6O8T7_0;
	wire w_dff_A_hgnZjgYK5_0;
	wire w_dff_A_SfblFLUk0_0;
	wire w_dff_A_64hgeVf47_0;
	wire w_dff_A_ETNdEqhN5_0;
	wire w_dff_A_zbdnEx7K1_0;
	wire w_dff_A_22EscIR99_0;
	wire w_dff_A_a8aItw0v3_0;
	wire w_dff_A_5kpXoC1t2_0;
	wire w_dff_A_EHeaxokn1_0;
	wire w_dff_A_wZR2sSl97_0;
	wire w_dff_A_NavXcQAt2_0;
	wire w_dff_A_lhIPVIyD9_0;
	wire w_dff_A_f03qnhYt6_0;
	wire w_dff_A_b7yAy11t3_0;
	wire w_dff_A_KvEh6WsY7_0;
	wire w_dff_A_OmK0mBkb3_0;
	wire w_dff_A_2svKVKTn5_0;
	wire w_dff_A_Tx7LCMRQ4_2;
	wire w_dff_A_14kAUU5Z8_0;
	wire w_dff_A_tOR2rClx1_0;
	wire w_dff_A_8tKSUArA0_0;
	wire w_dff_A_O4WH3Moz6_0;
	wire w_dff_A_qAHQIeSR5_0;
	wire w_dff_A_8R6gCynq5_0;
	wire w_dff_A_GAQ4nw440_0;
	wire w_dff_A_otVRNlBZ3_0;
	wire w_dff_A_GVJYovpm6_0;
	wire w_dff_A_ba9wSJl45_0;
	wire w_dff_A_zwwR4PAW8_0;
	wire w_dff_A_Y94x4yeA1_0;
	wire w_dff_A_Oklqd7mC8_0;
	wire w_dff_A_5kEttWOO0_0;
	wire w_dff_A_jRwE7Bb38_0;
	wire w_dff_A_Fxwxn6190_0;
	wire w_dff_A_Nwbfqv7e6_0;
	wire w_dff_A_IUMgHBSb2_0;
	wire w_dff_A_6RVcPaFp7_0;
	wire w_dff_A_b9U8rvN75_0;
	wire w_dff_A_nOvPMse80_0;
	wire w_dff_A_Y4c4Oc1T8_0;
	wire w_dff_A_Ogr1fN703_0;
	wire w_dff_A_VG6Z7uxI3_0;
	wire w_dff_A_4t5qomYy6_1;
	wire w_dff_A_JglmjN1Z4_0;
	wire w_dff_A_ccemzdBD0_0;
	wire w_dff_A_aCyYX4Zv1_0;
	wire w_dff_A_WfZ5zNkY2_0;
	wire w_dff_A_ZoDMpAIF7_0;
	wire w_dff_A_RPbtjc4T1_0;
	wire w_dff_A_yNyL1sjl9_0;
	wire w_dff_A_vP5aHVhj6_0;
	wire w_dff_A_LvHLTHhK7_0;
	wire w_dff_A_dA07wt589_0;
	wire w_dff_A_b8fij2VU1_0;
	wire w_dff_A_HZaXf0B80_0;
	wire w_dff_A_ntKySZrP0_0;
	wire w_dff_A_arLOqNh44_0;
	wire w_dff_A_rlY5AMvy7_0;
	wire w_dff_A_tve4drrI3_0;
	wire w_dff_A_iiRJTXmZ6_0;
	wire w_dff_A_LRxqIdLm7_0;
	wire w_dff_A_9NSZLUZQ9_0;
	wire w_dff_A_vc2SNTHS3_0;
	wire w_dff_A_f4EUHqpe8_0;
	wire w_dff_A_vZyTu1z64_0;
	wire w_dff_A_xcBrXdKy1_0;
	wire w_dff_A_0ppt8fdD7_0;
	wire w_dff_A_f8vZYw3H0_1;
	wire w_dff_A_yBdxMWK71_0;
	wire w_dff_A_vN1cUOXQ7_0;
	wire w_dff_A_7JvcQmRO2_0;
	wire w_dff_A_nDuukRtl4_0;
	wire w_dff_A_rKIDSq7L0_0;
	wire w_dff_A_1mCManc11_0;
	wire w_dff_A_fBWVuOqo5_0;
	wire w_dff_A_CKKeH1dR4_0;
	wire w_dff_A_3K8EO7L29_0;
	wire w_dff_A_1tByP6EO5_0;
	wire w_dff_A_yCCE39p71_0;
	wire w_dff_A_wMWEL7dG6_0;
	wire w_dff_A_pTEvlNLI1_0;
	wire w_dff_A_cJcdngc56_0;
	wire w_dff_A_rlQvqZ9v0_0;
	wire w_dff_A_BPeS75Ta9_0;
	wire w_dff_A_F4V4fGZr8_0;
	wire w_dff_A_rGqMNOaA1_0;
	wire w_dff_A_cpvzZGOd5_0;
	wire w_dff_A_MtZUFIL39_0;
	wire w_dff_A_EUW4a9A54_0;
	wire w_dff_A_zeWAjc868_0;
	wire w_dff_A_7gTExLR42_0;
	wire w_dff_A_8T28QgsW3_0;
	wire w_dff_A_BdUBaggz8_1;
	wire w_dff_A_Iyz5s8VD6_0;
	wire w_dff_A_rJa9VwBA8_0;
	wire w_dff_A_QVPeiX7F6_0;
	wire w_dff_A_qhyRiV6p2_0;
	wire w_dff_A_nf3YsK3B5_0;
	wire w_dff_A_vHtItjyK8_0;
	wire w_dff_A_QAtxzspg8_0;
	wire w_dff_A_VsD6A8DB1_0;
	wire w_dff_A_zqBjAU7L5_0;
	wire w_dff_A_6iaFECpC8_0;
	wire w_dff_A_1dBIaVfv0_0;
	wire w_dff_A_la3wU6Ia6_0;
	wire w_dff_A_UhXVFHhA6_0;
	wire w_dff_A_aSed0eb27_0;
	wire w_dff_A_YbUCoBjD5_0;
	wire w_dff_A_LRApCwlo7_0;
	wire w_dff_A_2N5mlHuM8_0;
	wire w_dff_A_9Y56wAhA6_0;
	wire w_dff_A_XszV9iEO3_0;
	wire w_dff_A_n3Rrntqs8_0;
	wire w_dff_A_u3IPBKOP0_0;
	wire w_dff_A_aKAfical2_0;
	wire w_dff_A_AybOmuZK5_0;
	wire w_dff_A_luNwuZrr4_0;
	wire w_dff_A_O7dZoQl30_1;
	wire w_dff_A_V1Tcj7mQ9_0;
	wire w_dff_A_3Pi8NwzR5_0;
	wire w_dff_A_OXFg8ti32_0;
	wire w_dff_A_F5iUhkOb8_0;
	wire w_dff_A_wzrhIHIU7_0;
	wire w_dff_A_oSXYUSXL2_0;
	wire w_dff_A_eVhtiyi51_0;
	wire w_dff_A_UAzuIQyo6_0;
	wire w_dff_A_N0pLwbjx8_0;
	wire w_dff_A_PLXJVj9Y1_0;
	wire w_dff_A_BxwhdICT1_0;
	wire w_dff_A_kP9unsOF2_0;
	wire w_dff_A_20PUEmxL3_0;
	wire w_dff_A_ejkMAAZs3_0;
	wire w_dff_A_dCApbI2O4_0;
	wire w_dff_A_aU1wrsgp7_0;
	wire w_dff_A_jQsRCO0U5_0;
	wire w_dff_A_nXIB78Kc9_0;
	wire w_dff_A_kYEm73el2_0;
	wire w_dff_A_1PRRtXaw3_0;
	wire w_dff_A_HobxA5Cj0_0;
	wire w_dff_A_B0gsQ4BK5_0;
	wire w_dff_A_GiycBwh69_0;
	wire w_dff_A_qkA4Mohq0_0;
	wire w_dff_A_A73KRriC2_2;
	wire w_dff_A_QHRYgLdv8_0;
	wire w_dff_A_4LsF9tOB4_0;
	wire w_dff_A_hCGA9hfk1_0;
	wire w_dff_A_5FvsBG0u8_0;
	wire w_dff_A_dKeRzE1w3_0;
	wire w_dff_A_gHQSSUmJ3_0;
	wire w_dff_A_t3MjPj938_0;
	wire w_dff_A_tZ0GWu3a2_0;
	wire w_dff_A_gLu1sFFu8_0;
	wire w_dff_A_qqsvjRxu1_0;
	wire w_dff_A_tC2Pwm532_0;
	wire w_dff_A_2uffUFaM1_0;
	wire w_dff_A_O6e1pLXQ9_0;
	wire w_dff_A_7cT1evW32_0;
	wire w_dff_A_z1RjZZO91_0;
	wire w_dff_A_YijuYlJI4_0;
	wire w_dff_A_8FDWZXzS1_0;
	wire w_dff_A_Nuw0kKu89_0;
	wire w_dff_A_6TvhlGT81_0;
	wire w_dff_A_B4UaiNhs6_0;
	wire w_dff_A_UHQVVD6z6_0;
	wire w_dff_A_Ok9DwsHL7_0;
	wire w_dff_A_b9BxmFUo9_0;
	wire w_dff_A_EItsgsMe4_0;
	wire w_dff_A_qRvqPe0K0_2;
	wire w_dff_A_D7KvJIcy7_0;
	wire w_dff_A_DaslA0fS3_0;
	wire w_dff_A_3QGzizf21_0;
	wire w_dff_A_tsk0zT4j5_0;
	wire w_dff_A_gduYHa7o0_0;
	wire w_dff_A_DvSzl4zs3_0;
	wire w_dff_A_v50RVdLI0_0;
	wire w_dff_A_orj4xZUA5_0;
	wire w_dff_A_rh5tpSUG7_0;
	wire w_dff_A_I0CqYIGO7_0;
	wire w_dff_A_4wdrDtqJ4_0;
	wire w_dff_A_Mxse4G6a9_0;
	wire w_dff_A_Cx8DkS5H3_0;
	wire w_dff_A_eBnPuevc3_0;
	wire w_dff_A_uROkI5549_0;
	wire w_dff_A_bdmvwmqG5_0;
	wire w_dff_A_YfhpMKSF4_0;
	wire w_dff_A_66Mgpz6z8_0;
	wire w_dff_A_CfEES1kc0_0;
	wire w_dff_A_4ab1mCmT7_0;
	wire w_dff_A_jGYyayqq1_0;
	wire w_dff_A_qjFC11q62_0;
	wire w_dff_A_sdlJCghR9_0;
	wire w_dff_A_hpXzg0xe9_2;
	wire w_dff_A_TWtoqQQE9_0;
	wire w_dff_A_ngK5VdIU5_0;
	wire w_dff_A_G65L7igr6_0;
	wire w_dff_A_nlB2Z9oG0_0;
	wire w_dff_A_SeMPnqRd8_0;
	wire w_dff_A_jBQt9ucz5_0;
	wire w_dff_A_ubcbUSwX4_0;
	wire w_dff_A_zlTo5ASg6_0;
	wire w_dff_A_ppqfRdBU7_0;
	wire w_dff_A_WB1f71cN7_0;
	wire w_dff_A_leGahstU2_0;
	wire w_dff_A_UOCkYlVC0_0;
	wire w_dff_A_TXicrlqP7_0;
	wire w_dff_A_7AJTUEqQ3_0;
	wire w_dff_A_LMJS409g4_0;
	wire w_dff_A_QR8GrEX93_0;
	wire w_dff_A_sDua6Qoj6_0;
	wire w_dff_A_G2eDTmua9_0;
	wire w_dff_A_w8qi5ew93_0;
	wire w_dff_A_Eeoy4mWu5_0;
	wire w_dff_A_l9LU6LYt1_0;
	wire w_dff_A_2gjwdEwy1_0;
	wire w_dff_A_V33cnRmT1_0;
	wire w_dff_A_ViUahs343_1;
	wire w_dff_A_iooO0VpB8_0;
	wire w_dff_A_GqFfNTRm6_0;
	wire w_dff_A_DIAmK1Gj2_0;
	wire w_dff_A_l58GALg67_0;
	wire w_dff_A_VwiD7fc74_0;
	wire w_dff_A_jQ7aw5Ve5_0;
	wire w_dff_A_ZXp10W1O4_0;
	wire w_dff_A_TLzDrl8S1_0;
	wire w_dff_A_x4LqO9DE2_0;
	wire w_dff_A_Q5EXAufB1_0;
	wire w_dff_A_FubuaEPB5_0;
	wire w_dff_A_mq4gRUuZ2_0;
	wire w_dff_A_DalA584P0_0;
	wire w_dff_A_SvTN4RbA8_0;
	wire w_dff_A_v4muk1iP9_0;
	wire w_dff_A_c7zLx6yB7_0;
	wire w_dff_A_tprq0Hsr1_0;
	wire w_dff_A_aNegmzWn2_0;
	wire w_dff_A_M0CC1hHB9_0;
	wire w_dff_A_j82XPKqP0_0;
	wire w_dff_A_jXyNHNnt2_0;
	wire w_dff_A_6ayynWL57_0;
	wire w_dff_A_QBe88BDj7_0;
	wire w_dff_A_sj71NC4V1_1;
	wire w_dff_A_u8QhvmQL6_0;
	wire w_dff_A_18pQDlkp1_0;
	wire w_dff_A_zNK6xxn77_0;
	wire w_dff_A_YN3cziQw5_0;
	wire w_dff_A_Bpgxn6Dk3_0;
	wire w_dff_A_RY7KrXhu6_0;
	wire w_dff_A_XBvdImye8_0;
	wire w_dff_A_Zcu60hBh6_0;
	wire w_dff_A_jumul6F60_0;
	wire w_dff_A_KpG0jdCq9_0;
	wire w_dff_A_rx8Hxp1C9_0;
	wire w_dff_A_lD9JQRWf1_0;
	wire w_dff_A_yvK7Q4Cv6_0;
	wire w_dff_A_eICuoqTu9_0;
	wire w_dff_A_kWXSdlQl2_0;
	wire w_dff_A_Yr1dCKCl0_0;
	wire w_dff_A_PugyfsXq2_0;
	wire w_dff_A_KFSqPgz87_0;
	wire w_dff_A_palNUYEn7_0;
	wire w_dff_A_B5b7hgEZ1_0;
	wire w_dff_A_FFtnOU926_0;
	wire w_dff_A_NPFPFwoX6_0;
	wire w_dff_A_hlJLiJZ32_0;
	wire w_dff_A_T4XgKpFB1_0;
	wire w_dff_A_lBK96Nf12_0;
	wire w_dff_A_HaCj6xuk2_1;
	wire w_dff_A_Do4ByAWj8_0;
	wire w_dff_A_pEXzaAKn9_0;
	wire w_dff_A_LneWEKAY7_0;
	wire w_dff_A_eDcx02rZ3_0;
	wire w_dff_A_Bxoy26mD0_0;
	wire w_dff_A_s6as2Cm73_0;
	wire w_dff_A_Xo2Jylnz4_0;
	wire w_dff_A_MoZ7CPFV7_0;
	wire w_dff_A_3m05lXNH2_0;
	wire w_dff_A_epk0eIWO1_0;
	wire w_dff_A_GLoXhBjM3_0;
	wire w_dff_A_SwNnoWVC5_0;
	wire w_dff_A_GDDK4qB99_0;
	wire w_dff_A_UlkBzqS80_0;
	wire w_dff_A_RjcBw8jC4_0;
	wire w_dff_A_NDF14ZRB0_0;
	wire w_dff_A_4NIJGMTk7_0;
	wire w_dff_A_p0ja5tRh9_0;
	wire w_dff_A_XQSXx6Ub9_0;
	wire w_dff_A_RKpPEadB9_0;
	wire w_dff_A_7SHw5ATD8_0;
	wire w_dff_A_6Khi0dL85_0;
	wire w_dff_A_s42y9RX06_0;
	wire w_dff_A_nuSZYBV88_0;
	wire w_dff_A_Y3MnGbpo4_0;
	wire w_dff_A_n3PHt2IB0_1;
	wire w_dff_A_bslqJ3iy3_0;
	wire w_dff_A_lwbjCbjp8_0;
	wire w_dff_A_5A6w6emc4_0;
	wire w_dff_A_ssXT6xpk9_0;
	wire w_dff_A_dCNjHbkt8_0;
	wire w_dff_A_5pspdUro8_0;
	wire w_dff_A_qdlZwsXj9_0;
	wire w_dff_A_CI3UD1XA2_0;
	wire w_dff_A_BIuxpNiH4_0;
	wire w_dff_A_ypZiefm88_0;
	wire w_dff_A_nD5N2UIu4_0;
	wire w_dff_A_YcznuUwt2_0;
	wire w_dff_A_CVAGcaXa1_0;
	wire w_dff_A_n09Nnwt84_0;
	wire w_dff_A_pfBjQgUp0_0;
	wire w_dff_A_6DapTIE14_0;
	wire w_dff_A_oZW4B5QZ4_0;
	wire w_dff_A_bUsUSjIn0_0;
	wire w_dff_A_EA4aZZpD4_0;
	wire w_dff_A_xj2oHy7A8_0;
	wire w_dff_A_urw1ziEL2_0;
	wire w_dff_A_nKjh5oZt2_0;
	wire w_dff_A_FILaSPKv5_0;
	wire w_dff_A_KI8CJEtM4_0;
	wire w_dff_A_9FnmD0E05_0;
	wire w_dff_A_Gx44yVSc7_1;
	wire w_dff_A_kfethRvJ8_0;
	wire w_dff_A_wNrtEa7B8_0;
	wire w_dff_A_aXEvXYaV5_0;
	wire w_dff_A_61Yjs9Fi8_0;
	wire w_dff_A_JlmwLIQT2_0;
	wire w_dff_A_fong6TIP8_0;
	wire w_dff_A_4MXegcaY7_0;
	wire w_dff_A_Q55zYvG36_0;
	wire w_dff_A_GXKKp3W53_0;
	wire w_dff_A_tZpmmXVc1_0;
	wire w_dff_A_75xU5udf0_0;
	wire w_dff_A_fMTdgve52_0;
	wire w_dff_A_jwNI3Ic87_0;
	wire w_dff_A_8r6bQmHS7_0;
	wire w_dff_A_IZb8XFCE9_0;
	wire w_dff_A_Nfs7hVum7_0;
	wire w_dff_A_xvxoChTQ2_0;
	wire w_dff_A_ySY0MIM84_0;
	wire w_dff_A_BmZI0J9D9_0;
	wire w_dff_A_cG0Ai9um9_0;
	wire w_dff_A_TZDqMABz9_0;
	wire w_dff_A_qdRxkQvC4_0;
	wire w_dff_A_VCRbQayE6_0;
	wire w_dff_A_MIiA93gJ4_0;
	wire w_dff_A_4HnryNRv4_0;
	wire w_dff_A_omMcWl0V5_1;
	wire w_dff_A_tRwaXqEU9_0;
	wire w_dff_A_ACf52F0F0_0;
	wire w_dff_A_W5kvFPZr5_0;
	wire w_dff_A_uzBXmwV79_0;
	wire w_dff_A_hMjOgwuS1_0;
	wire w_dff_A_nh3uSt8b6_0;
	wire w_dff_A_759wugz15_0;
	wire w_dff_A_zyIDLgoI3_0;
	wire w_dff_A_MnNdpAUC3_0;
	wire w_dff_A_crKFmxLn0_0;
	wire w_dff_A_lzMNu7TQ3_0;
	wire w_dff_A_y47jTir70_0;
	wire w_dff_A_2NXNj62p0_0;
	wire w_dff_A_TJn0iHql8_0;
	wire w_dff_A_nWBDILmJ2_0;
	wire w_dff_A_tds29IkS8_0;
	wire w_dff_A_bXJ5YoBX1_0;
	wire w_dff_A_LzUIwyaC7_0;
	wire w_dff_A_gGxr83iC6_0;
	wire w_dff_A_IlIOQTTt9_0;
	wire w_dff_A_FfXLtBh03_0;
	wire w_dff_A_QDHA37He2_0;
	wire w_dff_A_TxLsiOcT8_0;
	wire w_dff_A_TVUS04Wy4_0;
	wire w_dff_A_bw4nEjLL6_0;
	wire w_dff_A_KkjYaiEQ9_1;
	wire w_dff_A_37rmaHFS4_0;
	wire w_dff_A_iAvk41Do5_0;
	wire w_dff_A_CGg2NHQu7_0;
	wire w_dff_A_BUorYZW25_0;
	wire w_dff_A_l1iMm9iP7_0;
	wire w_dff_A_3eQzTXUd7_0;
	wire w_dff_A_Au4ouYjb2_0;
	wire w_dff_A_Hnnb46RA5_0;
	wire w_dff_A_u0FIKi8D7_0;
	wire w_dff_A_98jx0DKn8_0;
	wire w_dff_A_GQsBvA5B7_0;
	wire w_dff_A_Trn5Sxqr3_0;
	wire w_dff_A_KAHbB80g2_0;
	wire w_dff_A_BVxY8GzL7_0;
	wire w_dff_A_Srngh5hg1_0;
	wire w_dff_A_gJnKQ1gH6_0;
	wire w_dff_A_13zGVZPW0_0;
	wire w_dff_A_PA6JAdQw6_0;
	wire w_dff_A_lkMTwbdw2_0;
	wire w_dff_A_Uz3M34Jx7_0;
	wire w_dff_A_6WIGjWsv7_0;
	wire w_dff_A_kgYb3Kz07_0;
	wire w_dff_A_7zLEWMT62_0;
	wire w_dff_A_xHjP5IS19_0;
	wire w_dff_A_TeUGITqX2_2;
	wire w_dff_A_ZCWtzJSQ0_0;
	wire w_dff_A_FB0ppcoU5_0;
	wire w_dff_A_dprZnLz11_0;
	wire w_dff_A_Rz8X0FA01_0;
	wire w_dff_A_GMOGhMJd9_0;
	wire w_dff_A_UlIXDjWl3_0;
	wire w_dff_A_r09MFtEO1_0;
	wire w_dff_A_BIZe2Idh7_0;
	wire w_dff_A_pSDFP8IT6_0;
	wire w_dff_A_GuPYyWVO8_0;
	wire w_dff_A_3qr1ixEV8_0;
	wire w_dff_A_XfhO3DZo7_0;
	wire w_dff_A_fGRjIBvF9_0;
	wire w_dff_A_P83KR6rp4_0;
	wire w_dff_A_3IKFuf0c0_0;
	wire w_dff_A_EFgaN5sF1_0;
	wire w_dff_A_XnDof0qX9_0;
	wire w_dff_A_VgPj72L81_0;
	wire w_dff_A_Y4mUHlXV0_0;
	wire w_dff_A_Sur98lIL2_0;
	wire w_dff_A_hv8wnq873_0;
	wire w_dff_A_3P1pUxhw8_0;
	wire w_dff_A_j3HNxQs77_2;
	wire w_dff_A_Ts6Jurkj7_0;
	wire w_dff_A_nK0AWwSp4_0;
	wire w_dff_A_2UtaPUNn0_0;
	wire w_dff_A_A2bSnDeh5_0;
	wire w_dff_A_xnDITRUY1_0;
	wire w_dff_A_pmuwjlej6_0;
	wire w_dff_A_sqWnpmwm9_0;
	wire w_dff_A_RrO9wq0O9_0;
	wire w_dff_A_G5CRzuJP7_0;
	wire w_dff_A_vQDry5gr4_0;
	wire w_dff_A_Z1Q08JJD2_0;
	wire w_dff_A_TFX58myf6_0;
	wire w_dff_A_iJbLTe5r2_0;
	wire w_dff_A_77SJkW3d7_0;
	wire w_dff_A_HDs3TPly7_0;
	wire w_dff_A_PHcTUTMS3_0;
	wire w_dff_A_X8316fVC6_0;
	wire w_dff_A_9angCHJB9_0;
	wire w_dff_A_gaDTap2v7_0;
	wire w_dff_A_avJB5NEK5_0;
	wire w_dff_A_gNvvd1LB5_0;
	wire w_dff_A_XdcOMGSy6_0;
	wire w_dff_A_BV1QvbK34_0;
	wire w_dff_A_souf8wzQ9_1;
	wire w_dff_A_sohbHvtO3_0;
	wire w_dff_A_1hlssLp53_0;
	wire w_dff_A_56rwGcC02_0;
	wire w_dff_A_cNgu48bF9_0;
	wire w_dff_A_8I3ladya6_0;
	wire w_dff_A_XMMLbFry8_0;
	wire w_dff_A_dTQuhFCU0_0;
	wire w_dff_A_eoLUDWS09_0;
	wire w_dff_A_SsN5C4260_0;
	wire w_dff_A_Va0eIH452_0;
	wire w_dff_A_zTDQF9uP0_0;
	wire w_dff_A_qMzMVPyK5_0;
	wire w_dff_A_SKNZPdFB0_0;
	wire w_dff_A_hRGfadrq8_0;
	wire w_dff_A_yqKAlLtL1_0;
	wire w_dff_A_CT5Xi9Sc4_0;
	wire w_dff_A_Tu7SSuAh3_0;
	wire w_dff_A_tWKfunQL0_0;
	wire w_dff_A_FMxVe5KS4_0;
	wire w_dff_A_TUaljnmm9_0;
	wire w_dff_A_NYjwMUd90_0;
	wire w_dff_A_xYxAgG1G7_0;
	wire w_dff_A_VXAjTzj17_0;
	wire w_dff_A_hJTCLf5r2_0;
	wire w_dff_A_iRIb9Db31_0;
	wire w_dff_A_ezKNDcPo0_1;
	wire w_dff_A_kTjnUn804_0;
	wire w_dff_A_ypujY40A4_0;
	wire w_dff_A_OsNx4ymZ7_0;
	wire w_dff_A_8zcrnIHL0_0;
	wire w_dff_A_YOUzHR8T8_0;
	wire w_dff_A_OCLBUumw8_0;
	wire w_dff_A_NJjdlZkG5_0;
	wire w_dff_A_eOvvMheU8_0;
	wire w_dff_A_eLgRBT7h4_0;
	wire w_dff_A_Wvf1Pxkn8_0;
	wire w_dff_A_lnqTQAeb4_0;
	wire w_dff_A_CuEQSgoi6_0;
	wire w_dff_A_nfTbMoVz2_0;
	wire w_dff_A_NDjX91AQ8_0;
	wire w_dff_A_zFNT25fk3_0;
	wire w_dff_A_Da44n6E71_0;
	wire w_dff_A_pFs9W2I26_0;
	wire w_dff_A_ANyzpBGA6_0;
	wire w_dff_A_Zx3Z1ZgQ9_0;
	wire w_dff_A_uHNbxmZ29_0;
	wire w_dff_A_QUweVljw1_0;
	wire w_dff_A_TGETJrkQ3_0;
	wire w_dff_A_GbRv2wqN1_0;
	wire w_dff_A_RTci2qEH8_0;
	wire w_dff_A_8gEV0b435_0;
	wire w_dff_A_FmBKNEEe6_1;
	wire w_dff_A_uHjSMvx90_0;
	wire w_dff_A_MtrizcXo7_0;
	wire w_dff_A_JHPeRswh6_0;
	wire w_dff_A_s2Wbzplc0_0;
	wire w_dff_A_9xtsbFfg2_0;
	wire w_dff_A_4niLbNtt5_0;
	wire w_dff_A_I3ZjgZK78_0;
	wire w_dff_A_SXGMLNcz5_0;
	wire w_dff_A_FZoCUiy34_0;
	wire w_dff_A_yap5GLYK3_0;
	wire w_dff_A_gyNZpwcy1_0;
	wire w_dff_A_en156vvS4_0;
	wire w_dff_A_AfeoRSEh3_0;
	wire w_dff_A_x8giCt9r2_0;
	wire w_dff_A_dRtqPKuB3_0;
	wire w_dff_A_pFqz7zf01_0;
	wire w_dff_A_hz3Cv4bT7_0;
	wire w_dff_A_YzRnybzk7_0;
	wire w_dff_A_rqQ9f4I73_0;
	wire w_dff_A_eTohmUmJ5_0;
	wire w_dff_A_tlembwPc2_0;
	wire w_dff_A_oynZh5sH8_0;
	wire w_dff_A_7NQSHuoH9_0;
	wire w_dff_A_7qS01c9g8_0;
	wire w_dff_A_8itBNWBZ5_0;
	wire w_dff_A_nZRgG5262_1;
	wire w_dff_A_n0DEsO647_0;
	wire w_dff_A_NxA3MFIe6_0;
	wire w_dff_A_Bxlv6EiW3_0;
	wire w_dff_A_EMW9azd01_0;
	wire w_dff_A_Sbput8P13_0;
	wire w_dff_A_u7iNuL7L9_0;
	wire w_dff_A_7r5mLf335_0;
	wire w_dff_A_oTyKjcqZ7_0;
	wire w_dff_A_BkCOtPlg8_0;
	wire w_dff_A_u9XL9JiD6_0;
	wire w_dff_A_Qd88GtDw2_0;
	wire w_dff_A_LftG2yA64_0;
	wire w_dff_A_ZuijdhyB5_0;
	wire w_dff_A_i2dPcf8c3_0;
	wire w_dff_A_1v6fKkZt6_0;
	wire w_dff_A_SsNQQLZ38_0;
	wire w_dff_A_M4wsOCKc6_0;
	wire w_dff_A_1kPZT8yf6_0;
	wire w_dff_A_f0tGfCn38_0;
	wire w_dff_A_irplmtP10_0;
	wire w_dff_A_UU2y8qZI4_0;
	wire w_dff_A_WDG89NpS6_0;
	wire w_dff_A_lSmUJkuW6_0;
	wire w_dff_A_sRiGetB06_0;
	wire w_dff_A_p9zxiRJd1_0;
	wire w_dff_A_eXIkQR0I3_1;
	wire w_dff_A_LU4KLaQz4_0;
	wire w_dff_A_kXyhF1CE8_0;
	wire w_dff_A_nY08GLQu3_0;
	wire w_dff_A_ZFvPONps7_0;
	wire w_dff_A_cajAvpJP8_0;
	wire w_dff_A_Om81QiMW5_0;
	wire w_dff_A_N6G5mIwj7_0;
	wire w_dff_A_sYLLraH33_0;
	wire w_dff_A_n8riWIWi9_0;
	wire w_dff_A_GcRCZb8I2_0;
	wire w_dff_A_2G98fjIZ7_0;
	wire w_dff_A_jz2AJcTg0_0;
	wire w_dff_A_QWZmy7Hx4_0;
	wire w_dff_A_33uK8JQk4_0;
	wire w_dff_A_mGRRoOep8_0;
	wire w_dff_A_MxJ6BjHc7_0;
	wire w_dff_A_GX7WeA8R7_0;
	wire w_dff_A_wpCDQzop7_0;
	wire w_dff_A_PDL2VOF95_0;
	wire w_dff_A_ZDLqX4uF2_0;
	wire w_dff_A_u8bgHKvf1_0;
	wire w_dff_A_dGBChYzy0_0;
	wire w_dff_A_FG7jujTQ9_0;
	wire w_dff_A_RC6yfMHf3_0;
	wire w_dff_A_envOpYwf6_0;
	wire w_dff_A_KMUkwXSO1_1;
	wire w_dff_A_89a6khRD5_0;
	wire w_dff_A_t7KoX3Mz3_0;
	wire w_dff_A_UNcfpJRv2_0;
	wire w_dff_A_iab2UFPQ0_0;
	wire w_dff_A_uYkEWure5_0;
	wire w_dff_A_F3iC9brH9_0;
	wire w_dff_A_HUxslvW57_0;
	wire w_dff_A_xp9gBtPA6_0;
	wire w_dff_A_mEcvr3lh2_0;
	wire w_dff_A_uf2sLu1l1_0;
	wire w_dff_A_4Wsui3iD7_0;
	wire w_dff_A_yx5CXPkn7_0;
	wire w_dff_A_ZdgZX82D2_0;
	wire w_dff_A_y5NJj0W41_0;
	wire w_dff_A_4nWin5EN5_0;
	wire w_dff_A_JYYNbSlL3_0;
	wire w_dff_A_rkXzrh7J8_0;
	wire w_dff_A_3BXvPA8k1_0;
	wire w_dff_A_eTTwXyHP5_0;
	wire w_dff_A_MX4lXgeB5_0;
	wire w_dff_A_13nVuEtI9_0;
	wire w_dff_A_RkqjJyFY5_0;
	wire w_dff_A_8jLSMEHM0_0;
	wire w_dff_A_OYwj7SfF3_0;
	wire w_dff_A_he6umlfr2_2;
	wire w_dff_A_sexO35Lf7_0;
	wire w_dff_A_AgcW8LBO0_0;
	wire w_dff_A_mMV86RFB5_0;
	wire w_dff_A_ty5sv9pU7_0;
	wire w_dff_A_lnJ1U2dA9_0;
	wire w_dff_A_cwO910r85_0;
	wire w_dff_A_6ymS5dNn5_0;
	wire w_dff_A_CIgUKtGE0_0;
	wire w_dff_A_mvMVnw3A7_0;
	wire w_dff_A_WMlCXaE18_0;
	wire w_dff_A_V7Iw77Eo1_0;
	wire w_dff_A_6gkHl4Gz2_0;
	wire w_dff_A_gxIXcJuF4_0;
	wire w_dff_A_HjMMdCrg9_0;
	wire w_dff_A_fszR8mFn5_0;
	wire w_dff_A_hXjQTx3Z5_0;
	wire w_dff_A_wBdsQp144_0;
	wire w_dff_A_iSippFl31_0;
	wire w_dff_A_sDAWGRxa1_0;
	wire w_dff_A_23BfwigB4_0;
	wire w_dff_A_rNopzjx29_0;
	wire w_dff_A_NGvHq2GN5_2;
	wire w_dff_A_vNm62C9x0_0;
	wire w_dff_A_vcZGSRff3_0;
	wire w_dff_A_vKDY7iSK7_0;
	wire w_dff_A_nMlA0hMx5_0;
	wire w_dff_A_YAOJots17_0;
	wire w_dff_A_PAUk9OZU5_0;
	wire w_dff_A_ryMEEiyR5_0;
	wire w_dff_A_l0XSivFZ6_0;
	wire w_dff_A_VV8wepkk8_0;
	wire w_dff_A_8u3yfmOK5_0;
	wire w_dff_A_dVh5TqkM3_0;
	wire w_dff_A_Pqxdr7IE9_0;
	wire w_dff_A_4AChNxay2_0;
	wire w_dff_A_C150Q0tt3_0;
	wire w_dff_A_9N38gbhl7_0;
	wire w_dff_A_0mBXMIi36_0;
	wire w_dff_A_wh0uLp1j0_0;
	wire w_dff_A_pOdBPloB2_0;
	wire w_dff_A_BTQsVohP9_0;
	wire w_dff_A_7Dqc6S1E0_0;
	wire w_dff_A_d6dtyzNd9_0;
	wire w_dff_A_uUv6KBve7_2;
	wire w_dff_A_EewyZC9F5_0;
	wire w_dff_A_VyOlxq200_0;
	wire w_dff_A_ufqK6YQZ5_0;
	wire w_dff_A_AstLLh6v8_0;
	wire w_dff_A_Rfi9z38C6_0;
	wire w_dff_A_g0742VEN5_0;
	wire w_dff_A_YeRBJudE5_0;
	wire w_dff_A_r96IHjct1_0;
	wire w_dff_A_p7ShS8qT7_0;
	wire w_dff_A_KvcXPd341_0;
	wire w_dff_A_tN0ZeT0k5_0;
	wire w_dff_A_rqYdR5fk6_0;
	wire w_dff_A_THHISChu1_0;
	wire w_dff_A_lXoB0zgw1_0;
	wire w_dff_A_IY7JPQEK2_0;
	wire w_dff_A_UYODEuev1_0;
	wire w_dff_A_uVaMD4Ke5_0;
	wire w_dff_A_KMrbPvDL8_0;
	wire w_dff_A_EjvmdIYi6_0;
	wire w_dff_A_gogDgxR12_0;
	wire w_dff_A_Zo98GRJt8_0;
	wire w_dff_A_AJ2uePYK9_2;
	wire w_dff_A_9nfbdfoe2_0;
	wire w_dff_A_PZbiJtIr9_0;
	wire w_dff_A_cIx3DeVm6_0;
	wire w_dff_A_svPrc4Ps7_0;
	wire w_dff_A_WWGGyxbn3_0;
	wire w_dff_A_4zeLb0rg3_0;
	wire w_dff_A_Nyo9VvHv1_0;
	wire w_dff_A_e3D1hQGu9_0;
	wire w_dff_A_NhqbKtqH8_0;
	wire w_dff_A_Nztr2vP84_0;
	wire w_dff_A_hsgqY5G03_0;
	wire w_dff_A_Xq7WlHVc4_0;
	wire w_dff_A_ghgonSyV3_0;
	wire w_dff_A_nfWjngP05_0;
	wire w_dff_A_EmvpCxco3_0;
	wire w_dff_A_nERXVkdJ8_0;
	wire w_dff_A_aPRijR0j0_0;
	wire w_dff_A_faV913vR9_0;
	wire w_dff_A_tJjvZw6A3_0;
	wire w_dff_A_d4dY939z5_0;
	wire w_dff_A_VjaejBQp5_0;
	wire w_dff_A_eBx9In5N7_0;
	wire w_dff_A_GFQkePVS7_2;
	wire w_dff_A_IuSSsg0Y5_0;
	wire w_dff_A_K5eCaWLY0_0;
	wire w_dff_A_yV3IbMqT1_0;
	wire w_dff_A_PhUHrHOZ7_0;
	wire w_dff_A_86xheCjg3_0;
	wire w_dff_A_MvYWYMLm1_0;
	wire w_dff_A_afGqxUSh5_0;
	wire w_dff_A_29OzCClW3_0;
	wire w_dff_A_xPfzRuKI6_0;
	wire w_dff_A_i3he0eTn3_0;
	wire w_dff_A_FBinRMAB2_0;
	wire w_dff_A_s9NQpRPR7_0;
	wire w_dff_A_qsIl0uKV7_0;
	wire w_dff_A_YAR7DUGh4_0;
	wire w_dff_A_xnnGLDJX7_0;
	wire w_dff_A_TuGhBZeR4_0;
	wire w_dff_A_XmFxiQdh2_0;
	wire w_dff_A_NVDhUuzE8_0;
	wire w_dff_A_2FCebLD21_0;
	wire w_dff_A_KaQOO7I14_0;
	wire w_dff_A_ws6qj8t84_2;
	wire w_dff_A_015pBpAd3_0;
	wire w_dff_A_OyNego9h7_0;
	wire w_dff_A_EqMQ4B6w1_0;
	wire w_dff_A_LdP7p3BV4_0;
	wire w_dff_A_6oMK9IOl0_0;
	wire w_dff_A_tjrGxKfB4_0;
	wire w_dff_A_z2q3Y7aL0_0;
	wire w_dff_A_NdQf38A18_0;
	wire w_dff_A_8imp4K072_0;
	wire w_dff_A_qQleIalw2_0;
	wire w_dff_A_HcjAf0SE6_0;
	wire w_dff_A_7YkBhXD80_0;
	wire w_dff_A_3zOfexpy2_0;
	wire w_dff_A_jq9AWYos0_0;
	wire w_dff_A_icRQlaTT8_0;
	wire w_dff_A_T92Cjpfb7_0;
	wire w_dff_A_4gYHMlAg4_0;
	wire w_dff_A_kbRzr4z37_0;
	wire w_dff_A_w7CZ9g636_0;
	wire w_dff_A_WfSr0u5T5_0;
	wire w_dff_A_JaHo8t0x7_2;
	wire w_dff_A_dIzQhL2j5_0;
	wire w_dff_A_ZvrQpCfx1_0;
	wire w_dff_A_V2esmU2Z2_0;
	wire w_dff_A_NaYIGfTX9_0;
	wire w_dff_A_UjMM8cGS7_0;
	wire w_dff_A_IlGHhJde7_0;
	wire w_dff_A_v6NsRYfv4_0;
	wire w_dff_A_bHbZaIgZ1_0;
	wire w_dff_A_lqN2WGM14_0;
	wire w_dff_A_jyyJPsk94_0;
	wire w_dff_A_6wu7qkfH2_0;
	wire w_dff_A_lHcTP5hU3_0;
	wire w_dff_A_3j7EJt0w8_0;
	wire w_dff_A_vXu0IyyP8_0;
	wire w_dff_A_x9rn4HH10_0;
	wire w_dff_A_OOPfshA13_0;
	wire w_dff_A_XT5aZqsB6_0;
	wire w_dff_A_duFMRqfy3_0;
	wire w_dff_A_p7YBxnct8_0;
	wire w_dff_A_3zglwhZp4_0;
	wire w_dff_A_bWD9Wu3L6_2;
	wire w_dff_A_egedGTJ07_0;
	wire w_dff_A_JygkQk1H6_0;
	wire w_dff_A_Lzy4S0Fj9_0;
	wire w_dff_A_n7pbn32l1_0;
	wire w_dff_A_C1JZcZK63_0;
	wire w_dff_A_Iat9NUY51_0;
	wire w_dff_A_N2p1n2bt4_0;
	wire w_dff_A_9TcUCaah0_0;
	wire w_dff_A_JvxMqBwD5_0;
	wire w_dff_A_RGvKg6k77_0;
	wire w_dff_A_onUMk9qV1_0;
	wire w_dff_A_sXd9QkmX8_0;
	wire w_dff_A_G2JjN1e75_0;
	wire w_dff_A_YNuWrXEO2_0;
	wire w_dff_A_qKhKx99B7_0;
	wire w_dff_A_YrSPJqTx1_0;
	wire w_dff_A_ON6UoYrD8_0;
	wire w_dff_A_BIfRkML18_0;
	wire w_dff_A_UrCQuzzc8_0;
	wire w_dff_A_hqxELb3E2_0;
	wire w_dff_A_xzIOgP9N0_2;
	wire w_dff_A_qtp2Zvl69_0;
	wire w_dff_A_tcxHJBT64_0;
	wire w_dff_A_fTmQci600_0;
	wire w_dff_A_zp8MIT2P7_0;
	wire w_dff_A_NkCSW3o55_0;
	wire w_dff_A_5z7rmwx18_0;
	wire w_dff_A_ryEFsn1F1_0;
	wire w_dff_A_TOGoBy9I1_0;
	wire w_dff_A_4FNNIWn95_0;
	wire w_dff_A_cxr9omFl3_0;
	wire w_dff_A_EPombFkj9_0;
	wire w_dff_A_nbJAbxhj8_0;
	wire w_dff_A_KwAFMWfm1_0;
	wire w_dff_A_vZP2OyaB3_0;
	wire w_dff_A_n81M39BH6_0;
	wire w_dff_A_nfvfRpeA3_0;
	wire w_dff_A_zRJ957kz3_2;
	wire w_dff_A_eJFULSEg9_0;
	wire w_dff_A_sf6JQtNE6_0;
	wire w_dff_A_y9QQgcGv4_0;
	wire w_dff_A_KxERmOrj0_0;
	wire w_dff_A_ZQ6MBruf4_0;
	wire w_dff_A_ljvutjJj6_0;
	wire w_dff_A_rFhpsRjl1_0;
	wire w_dff_A_qbzp1b9S9_0;
	wire w_dff_A_pPTsB0Vw1_0;
	wire w_dff_A_xBHpKUf87_0;
	wire w_dff_A_7yyuQvP80_0;
	wire w_dff_A_qQ24Hh9Q0_0;
	wire w_dff_A_OXYQVFwB5_0;
	wire w_dff_A_Tx7pZEYF5_0;
	wire w_dff_A_XXE4mgvB2_0;
	wire w_dff_A_3OQY6HDV2_0;
	wire w_dff_A_hKGz8qj65_2;
	wire w_dff_A_j6UBRRzF3_0;
	wire w_dff_A_wkuCNJ3M2_0;
	wire w_dff_A_NARCoohC0_0;
	wire w_dff_A_zyEip4tR0_0;
	wire w_dff_A_FPzSBU0J1_0;
	wire w_dff_A_C87JJzYi4_0;
	wire w_dff_A_NPoU0ZkM2_0;
	wire w_dff_A_6R3G86rj1_0;
	wire w_dff_A_3ItQFBkA7_0;
	wire w_dff_A_GsfTw6EV4_0;
	wire w_dff_A_LoKY0wd96_0;
	wire w_dff_A_c3XjQSlA5_0;
	wire w_dff_A_PZkWU55K1_0;
	wire w_dff_A_bIRRAvyk5_0;
	wire w_dff_A_CvoF0cw43_2;
	wire w_dff_A_DnFb1OsR6_0;
	wire w_dff_A_ropaRYC16_0;
	wire w_dff_A_zx6cagAZ3_0;
	wire w_dff_A_mnxyhXD91_0;
	wire w_dff_A_sOroxrfW4_0;
	wire w_dff_A_W8JoGkbB8_0;
	wire w_dff_A_Erdnakmx7_0;
	wire w_dff_A_fPdeymrQ6_0;
	wire w_dff_A_9tuJvtRw3_0;
	wire w_dff_A_8la4g7xV9_0;
	wire w_dff_A_38uRb4FB7_0;
	wire w_dff_A_iTXTnXOr7_0;
	wire w_dff_A_pRS8QfrQ9_0;
	wire w_dff_A_RrFlHIi41_0;
	wire w_dff_A_XN60dkC87_0;
	wire w_dff_A_Sz51mRe62_0;
	wire w_dff_A_VtM4hs6P0_2;
	wire w_dff_A_3zCBu4vo4_0;
	wire w_dff_A_TPdnABiS4_0;
	wire w_dff_A_By7JXafK2_0;
	wire w_dff_A_plpcEgRW6_0;
	wire w_dff_A_12BWs4LY1_0;
	wire w_dff_A_capNGH7F3_0;
	wire w_dff_A_qTvV0HAi9_0;
	wire w_dff_A_TbGJumbf8_0;
	wire w_dff_A_evBqJTV83_0;
	wire w_dff_A_pkH8XC9j1_0;
	wire w_dff_A_OcIZUuSL6_0;
	wire w_dff_A_81D5i6Vu8_0;
	wire w_dff_A_oWJNu1ep4_0;
	wire w_dff_A_5CkQLVEd2_0;
	wire w_dff_A_3g0Gxo518_0;
	wire w_dff_A_yBeqkK3y9_0;
	wire w_dff_A_tughExAl8_2;
	wire w_dff_A_ffPO6mIn1_0;
	wire w_dff_A_czdf2fEN5_0;
	wire w_dff_A_l7WpYvAV6_0;
	wire w_dff_A_YVKVgraS4_0;
	wire w_dff_A_Hczlb0RS4_0;
	wire w_dff_A_4lOsBLii7_0;
	wire w_dff_A_EEjO3bnx3_0;
	wire w_dff_A_VMSzwsEh6_0;
	wire w_dff_A_onJo3shw3_0;
	wire w_dff_A_1vlwOEM77_0;
	wire w_dff_A_eWvLJsfQ7_0;
	wire w_dff_A_2nzI1wQl5_0;
	wire w_dff_A_ra7phtSO1_0;
	wire w_dff_A_qJuZHddv4_0;
	wire w_dff_A_gwSMvLaq9_1;
	wire w_dff_A_40XfPXOS1_0;
	wire w_dff_A_jgLQuiM91_0;
	wire w_dff_A_h6R6veJV8_0;
	wire w_dff_A_8bO67LWI0_0;
	wire w_dff_A_JMNeqgL47_0;
	wire w_dff_A_YQK5lujo8_0;
	wire w_dff_A_ZTU1AUDK6_0;
	wire w_dff_A_h3ptnhXD5_0;
	wire w_dff_A_eva45roY5_0;
	wire w_dff_A_zWGAw06Y1_0;
	wire w_dff_A_3C5ScsxO7_0;
	wire w_dff_A_W1Lie4tp9_0;
	wire w_dff_A_7FKntTBz6_0;
	wire w_dff_A_t8OrPUSl5_0;
	wire w_dff_A_XNeGWqrB2_0;
	wire w_dff_A_drHtD34t4_0;
	wire w_dff_A_LBgFRq4P6_0;
	wire w_dff_A_40x3LFmT8_0;
	wire w_dff_A_TRxscYJQ9_0;
	wire w_dff_A_FQB1xfgN4_0;
	wire w_dff_A_ByIlIlBF7_1;
	wire w_dff_A_1fjAoNQt7_0;
	wire w_dff_A_yXhwmdtn3_0;
	wire w_dff_A_Deg2164w2_0;
	wire w_dff_A_noa6RaVy0_0;
	wire w_dff_A_DQG24vuE2_0;
	wire w_dff_A_d1i08bp22_0;
	wire w_dff_A_izEHIz1J5_0;
	wire w_dff_A_RCgnpovW7_0;
	wire w_dff_A_nn7kXtBx3_0;
	wire w_dff_A_kzNCJH836_0;
	wire w_dff_A_lmWg2PGX7_0;
	wire w_dff_A_Ek1LmCHy2_0;
	wire w_dff_A_cUWurIMW4_0;
	wire w_dff_A_kfCCRjIW9_0;
	wire w_dff_A_1Y1BBiEM8_0;
	wire w_dff_A_Dn8KA3kl9_0;
	wire w_dff_A_779Jtbhz6_0;
	wire w_dff_A_Jr3op34A3_0;
	wire w_dff_A_1TSZgapw6_0;
	wire w_dff_A_EPZ5jgC17_0;
	wire w_dff_A_svarlViU6_2;
	wire w_dff_A_CgGqpF836_0;
	wire w_dff_A_NMg4pjqI3_0;
	wire w_dff_A_6yfJuldK0_0;
	wire w_dff_A_PV4zbMzR9_0;
	wire w_dff_A_RIoTzfc38_0;
	wire w_dff_A_waHd4PJK8_0;
	wire w_dff_A_dcll5poU7_0;
	wire w_dff_A_BUpZESyO3_0;
	wire w_dff_A_R79aHdUu8_0;
	wire w_dff_A_WcT5831S3_0;
	wire w_dff_A_VbhswlOh8_0;
	wire w_dff_A_RURQqRW80_2;
	wire w_dff_A_gaijMJHj4_0;
	wire w_dff_A_EOaFZLwC3_0;
	wire w_dff_A_kZDFzEJi7_0;
	wire w_dff_A_G2tpAyLK6_0;
	wire w_dff_A_YUh8VSiC0_0;
	wire w_dff_A_sxFqwfWM4_0;
	wire w_dff_A_48QXFV8i3_0;
	wire w_dff_A_n1RyJHH69_0;
	wire w_dff_A_gNYiTFhq3_0;
	wire w_dff_A_wUMRnsvn6_0;
	wire w_dff_A_hMXyVOhu2_0;
	wire w_dff_A_xNiLG5rl1_2;
	wire w_dff_A_eLEZesFI3_0;
	wire w_dff_A_fX2CMInd4_0;
	wire w_dff_A_YXwtDJSN6_0;
	wire w_dff_A_OJCfiZg33_0;
	wire w_dff_A_ljoRMatz8_0;
	wire w_dff_A_uZNefROj7_0;
	wire w_dff_A_D6VtxZDf1_0;
	wire w_dff_A_30YzxlNw4_0;
	wire w_dff_A_mWntxtlV6_0;
	wire w_dff_A_2yVoIHCO8_0;
	wire w_dff_A_GU3Y6RPS4_0;
	wire w_dff_A_ePXT8ufG1_2;
	wire w_dff_A_z0Jec8un6_0;
	wire w_dff_A_8QYV5llE3_0;
	wire w_dff_A_SqtgFKu97_0;
	wire w_dff_A_GVGw5AXK7_0;
	wire w_dff_A_HBLn7Tfs9_0;
	wire w_dff_A_B0zSvSYp4_0;
	wire w_dff_A_BcDV8OsJ0_0;
	wire w_dff_A_GRimIAkU9_0;
	wire w_dff_A_srliIiHF8_0;
	wire w_dff_A_KCNV2Rsn3_0;
	wire w_dff_A_3jyohAHz4_0;
	wire w_dff_A_RYzzMdAy5_1;
	wire w_dff_A_FTpbQIZu1_0;
	wire w_dff_A_g6uo8kvg5_0;
	wire w_dff_A_VIJkmWqd7_0;
	wire w_dff_A_6TS5PpXV2_0;
	wire w_dff_A_gd5GNGdK7_0;
	wire w_dff_A_DNLsY7me4_0;
	wire w_dff_A_DDZHHVvW1_0;
	wire w_dff_A_AWAQaOAL0_0;
	wire w_dff_A_jzN1owR77_0;
	wire w_dff_A_NLwQEubE8_0;
	wire w_dff_A_g6X9JLKu1_0;
	wire w_dff_A_wyNgCw4k0_0;
	wire w_dff_A_iYCXIxq65_0;
	wire w_dff_A_3XKw3vF77_0;
	wire w_dff_A_ATk9Yafj6_0;
	wire w_dff_A_jgTXMd1D3_0;
	wire w_dff_A_UYBiSPz62_0;
	wire w_dff_A_BXewrYB48_0;
	wire w_dff_A_E3YaYj4k1_1;
	wire w_dff_A_GaVWyCWi6_0;
	wire w_dff_A_6RANbNUR6_0;
	wire w_dff_A_APKok7Mx8_0;
	wire w_dff_A_dToRJRTv6_0;
	wire w_dff_A_DPKrV4l86_0;
	wire w_dff_A_CA9LWPdx7_0;
	wire w_dff_A_U0qeOcNV5_0;
	wire w_dff_A_b1jmlzFU5_0;
	wire w_dff_A_lV6tL9Hb7_0;
	wire w_dff_A_7fxiZP2l2_0;
	wire w_dff_A_talPBM797_0;
	wire w_dff_A_3ojc82UW1_0;
	wire w_dff_A_98adCmWY7_0;
	wire w_dff_A_2JDsfYhm0_0;
	wire w_dff_A_vNzLAaKh6_0;
	wire w_dff_A_79Yqd6rA2_0;
	wire w_dff_A_ttEH5mM63_0;
	wire w_dff_A_A4wx6Pyj7_1;
	wire w_dff_A_x68XK9Bu2_0;
	wire w_dff_A_stzO46h05_0;
	wire w_dff_A_7XYiZ6wc2_0;
	wire w_dff_A_fvTuBpcE8_0;
	wire w_dff_A_b2KY147M0_0;
	wire w_dff_A_XXLaziDU4_0;
	wire w_dff_A_Nb9BxdPP4_0;
	wire w_dff_A_2E9AXDMD2_0;
	wire w_dff_A_FXggS7873_0;
	wire w_dff_A_a1WpbsJ89_0;
	wire w_dff_A_3oDDxfvV7_0;
	wire w_dff_A_Ff62aGNT9_0;
	wire w_dff_A_FdUActS05_0;
	wire w_dff_A_9NCUS5xc5_0;
	wire w_dff_A_NI5tmFbJ7_0;
	wire w_dff_A_GDeeSVIW2_0;
	wire w_dff_A_xa8ghJdf6_0;
	wire w_dff_A_FnIaWamW8_1;
	wire w_dff_A_LuPtvtwU1_0;
	wire w_dff_A_AXYs8PUz4_0;
	wire w_dff_A_FKcJVPB64_0;
	wire w_dff_A_KVT10t0a9_0;
	wire w_dff_A_lBqJxuSC9_0;
	wire w_dff_A_A5K3ofS42_0;
	wire w_dff_A_rihHI8OF6_2;
	wire w_dff_A_eeI1Jxay0_0;
	wire w_dff_A_OID7a4sf6_0;
	wire w_dff_A_55xCm2xS7_0;
	wire w_dff_A_bOqR8A041_0;
	wire w_dff_A_8O4T1LoU1_0;
	wire w_dff_A_HZEnsD2K1_0;
	wire w_dff_A_hlx3HPY17_0;
	wire w_dff_A_xrxJ6JMc9_0;
	wire w_dff_A_gKWlEoYD7_0;
	wire w_dff_A_ao8qu1wi5_0;
	wire w_dff_A_rjySDON30_0;
	wire w_dff_A_ryfqMpwG1_0;
	wire w_dff_A_Ccq3ENsc4_0;
	wire w_dff_A_FVQW5aGI6_0;
	wire w_dff_A_uwSrejso2_1;
	wire w_dff_A_qnVcuwuj1_0;
	wire w_dff_A_nx1js3GU7_0;
	wire w_dff_A_VyItlWFG2_0;
	wire w_dff_A_WxS5WOep8_0;
	wire w_dff_A_bsHJIzgf4_0;
	wire w_dff_A_SjmwnRyf1_0;
	wire w_dff_A_8LZyY8y66_0;
	wire w_dff_A_tgDbKMGN3_0;
	wire w_dff_A_0kykd7A99_0;
	wire w_dff_A_WxpaqE778_0;
	wire w_dff_A_FyKjELc89_0;
	wire w_dff_A_aPDiXqIJ5_1;
	wire w_dff_A_jNaqojDm6_0;
	wire w_dff_A_W2K8uwQ28_0;
	wire w_dff_A_eC56YHPc0_0;
	wire w_dff_A_jvbCF3kw6_0;
	wire w_dff_A_gPnaKhCS8_0;
	wire w_dff_A_5o62JWbn0_0;
	wire w_dff_A_3y4AB5eA4_0;
	wire w_dff_A_9AJ9G0cl9_0;
	wire w_dff_A_i4oXyeDj5_0;
	wire w_dff_A_I23kZXU87_0;
	wire w_dff_A_l5dGryT81_0;
	wire w_dff_A_LZdknmCY0_0;
	wire w_dff_A_u1r3E6Lz7_0;
	wire w_dff_A_oZ7aU2kK3_1;
	wire w_dff_A_uPCk3orv8_0;
	wire w_dff_A_E3loVfFT8_0;
	wire w_dff_A_a4aICiYl3_0;
	wire w_dff_A_bWO7ZxzZ0_0;
	wire w_dff_A_iElLYdJA5_0;
	wire w_dff_A_sCfjvzOF9_0;
	wire w_dff_A_u2rWZShp9_0;
	wire w_dff_A_ZqTfgCM72_0;
	wire w_dff_A_7XkPEuzN8_0;
	wire w_dff_A_EiyyASsV5_0;
	wire w_dff_A_beys8m2r1_0;
	wire w_dff_A_iVwUzesP6_0;
	wire w_dff_A_g0bV30pU2_0;
	wire w_dff_A_SyfuU3iZ7_0;
	wire w_dff_A_1ouZPPoB1_0;
	wire w_dff_A_89q19c2f0_2;
	wire w_dff_A_Ypvo3d9D6_0;
	wire w_dff_A_14VL949c5_0;
	wire w_dff_A_K739I5T62_0;
	wire w_dff_A_5m158jww1_0;
	wire w_dff_A_yx4Be42c0_0;
	wire w_dff_A_IzKVrTnF2_0;
	wire w_dff_A_NkjrtaDa3_0;
	wire w_dff_A_p2ptYhKI1_0;
	wire w_dff_A_nUA2XqSZ3_0;
	wire w_dff_A_SsrVvxOi9_0;
	wire w_dff_A_WefwJ0vb9_0;
	wire w_dff_A_tBWTraNr8_0;
	wire w_dff_A_K2ITEvA84_0;
	wire w_dff_A_q5P2WgGR7_0;
	wire w_dff_A_FEyi87VO8_1;
	wire w_dff_A_g4BCbAGH7_0;
	wire w_dff_A_wjhtsViz9_0;
	wire w_dff_A_xARsMCBG9_0;
	wire w_dff_A_0Z21CPDY7_0;
	wire w_dff_A_czH35Aou9_0;
	wire w_dff_A_Sb4LqZoM2_0;
	wire w_dff_A_48AlIWm59_0;
	wire w_dff_A_43Z0e5Zk7_0;
	wire w_dff_A_IpvMKZ2f3_0;
	wire w_dff_A_tbRIqskU5_1;
	wire w_dff_A_jMFEEjMW7_0;
	wire w_dff_A_H7hzk3cm5_0;
	wire w_dff_A_s6bBg3Zs0_0;
	wire w_dff_A_YldWtFF73_0;
	wire w_dff_A_vv40dYLN9_0;
	wire w_dff_A_FaAOVuM28_0;
	wire w_dff_A_xNzHx3ek6_0;
	wire w_dff_A_EnZ2ah4O2_0;
	wire w_dff_A_bYz1awt74_0;
	wire w_dff_A_COjP7ukv2_0;
	wire w_dff_A_XU7UePSo6_0;
	wire w_dff_A_mfZM6VHe2_1;
	wire w_dff_A_2Z2QYpFd4_0;
	wire w_dff_A_DeUiF1kp8_0;
	wire w_dff_A_IyahUs1U7_0;
	wire w_dff_A_nT7nrwXk7_0;
	wire w_dff_A_VPe2t4FT5_0;
	wire w_dff_A_vp1eqQtn9_0;
	wire w_dff_A_owdiU8qH9_0;
	wire w_dff_A_G8uOQpYS1_0;
	wire w_dff_A_5GlFC2W62_0;
	wire w_dff_A_Dop3JM336_0;
	wire w_dff_A_Yk4AJPXb0_0;
	wire w_dff_A_BnLjLJI84_0;
	wire w_dff_A_znHZByz42_1;
	wire w_dff_A_bkWzsQ1I4_0;
	wire w_dff_A_sQWx8T7X6_0;
	wire w_dff_A_XxRApIf52_0;
	wire w_dff_A_A1KtQVro2_0;
	wire w_dff_A_fIrn3unf0_0;
	wire w_dff_A_oCaCzonU1_0;
	wire w_dff_A_0oIqhyer7_0;
	wire w_dff_A_LI6TumCQ7_0;
	wire w_dff_A_JGhTj1ON6_0;
	wire w_dff_A_1WWVbI2O2_0;
	wire w_dff_A_BLXfFyri2_0;
	wire w_dff_A_DqE5aA3t1_0;
	wire w_dff_A_uUU8ObDp9_0;
	wire w_dff_A_DRK3FxjO7_1;
	wire w_dff_A_LdVKKNJk3_0;
	wire w_dff_A_vPBu5CHI5_0;
	wire w_dff_A_d5Y9Q4os1_0;
	wire w_dff_A_rifLNMZb9_0;
	wire w_dff_A_tXLLOhGW7_0;
	wire w_dff_A_fFGPrXvU8_0;
	wire w_dff_A_tqFdZqy68_0;
	wire w_dff_A_Y8W3ZcjZ7_0;
	wire w_dff_A_jD3nV72H4_0;
	wire w_dff_A_edx1i5tO4_0;
	wire w_dff_A_P0Pt5xk05_0;
	wire w_dff_A_246iYMQa6_0;
	wire w_dff_A_rLiQtCLX5_0;
	wire w_dff_A_MGmmWgBm1_0;
	wire w_dff_A_rOj99gq84_0;
	wire w_dff_A_hEiH5Yli0_0;
	wire w_dff_A_BMw7y2Ba7_1;
	wire w_dff_A_85Zvejto0_0;
	wire w_dff_A_xEBOynEa0_0;
	wire w_dff_A_XWd0Ya9Q3_0;
	wire w_dff_A_9HGnU0W98_0;
	wire w_dff_A_TGUJ1Fp62_0;
	wire w_dff_A_i2aa1icl5_0;
	wire w_dff_A_9rCsXmKf0_0;
	wire w_dff_A_y5ERnFou8_0;
	wire w_dff_A_twHqRVW34_0;
	wire w_dff_A_wl96eY8Y5_0;
	wire w_dff_A_oD8hCD429_0;
	wire w_dff_A_GcBTACSu1_0;
	wire w_dff_A_kgLVwoGE1_0;
	wire w_dff_A_qDdY1JAL2_0;
	wire w_dff_A_5iNAJwdU9_0;
	wire w_dff_A_B3HaQMSk3_0;
	wire w_dff_A_u6GuB5Nt4_0;
	wire w_dff_A_TjcllJTG9_0;
	wire w_dff_A_Fwk1ch9u3_2;
	wire w_dff_A_o8oOY3LR4_0;
	wire w_dff_A_AjGncHWn6_0;
	wire w_dff_A_RqljxeTi6_0;
	wire w_dff_A_igU8JoqH3_0;
	wire w_dff_A_Z53KL96c4_2;
	wire w_dff_A_5mJ2m0Ek4_0;
	wire w_dff_A_gpkqj7kl2_0;
	wire w_dff_A_v8GOvxvW2_0;
	wire w_dff_A_D3bAE0a97_0;
	wire w_dff_A_RBfckbjc4_0;
	wire w_dff_A_gmvIMtBQ3_0;
	wire w_dff_A_uf72IVJc7_0;
	wire w_dff_A_D17Lvw550_2;
	wire w_dff_A_Nl0vYpIb0_0;
	wire w_dff_A_EZFQrtM53_0;
	wire w_dff_A_TqrqK8yW0_0;
	wire w_dff_A_43TVzXho1_0;
	wire w_dff_A_GFDcnW2p4_0;
	wire w_dff_A_9wvA3qCw4_0;
	wire w_dff_A_n31SPELV6_0;
	wire w_dff_A_jIjvrTmC1_0;
	wire w_dff_A_BSvfZcAU7_0;
	wire w_dff_A_nwXmLbGK1_0;
	wire w_dff_A_8uShcWI16_0;
	wire w_dff_A_B2yupq7I3_0;
	wire w_dff_A_b8A31Ifd6_0;
	wire w_dff_A_vv4HfquM5_2;
	wire w_dff_A_KkjXm6oy9_0;
	wire w_dff_A_b7qG6Eah3_0;
	wire w_dff_A_dFXod8zO7_0;
	wire w_dff_A_FFtiDZHx9_0;
	wire w_dff_A_Hhjb7vcS3_0;
	wire w_dff_A_s6hIwy4Y9_0;
	wire w_dff_A_hFTaZZPg3_0;
	wire w_dff_A_p0oUpqlK1_0;
	wire w_dff_A_RAhw5FkQ9_0;
	wire w_dff_A_YryeKUfV2_0;
	wire w_dff_A_JdqdH2V45_0;
	wire w_dff_A_ugyEBPjS9_0;
	wire w_dff_A_CseCJxZM2_0;
	wire w_dff_A_4Kw7kf7E8_2;
	wire w_dff_A_q03HGYQX7_0;
	wire w_dff_A_k2zxiMXj1_0;
	wire w_dff_A_i8B80i0D0_0;
	wire w_dff_A_sPy6G2BC2_0;
	wire w_dff_A_KtRbgIqS5_0;
	wire w_dff_A_Rx4OdOu72_0;
	wire w_dff_A_J3ukU9lO6_2;
	wire w_dff_A_bPu5C7j15_0;
	wire w_dff_A_6WgIFvcY2_0;
	wire w_dff_A_1hRwUTZd1_0;
	wire w_dff_A_jREYj0yz0_0;
	wire w_dff_A_fb5Ztfsv2_0;
	wire w_dff_A_JQIK37c57_0;
	wire w_dff_A_UPgCFFjT2_0;
	wire w_dff_A_cas8e2kd0_0;
	wire w_dff_A_olIlU6Rz9_2;
	wire w_dff_A_KgngQVaW4_0;
	wire w_dff_A_zy7EuiiC8_0;
	wire w_dff_A_2VAYShV77_0;
	wire w_dff_A_sHQIN9RV8_0;
	wire w_dff_A_YfEFb6rC7_0;
	wire w_dff_A_8hvyRWUh6_0;
	wire w_dff_A_ziAl6mkq0_0;
	wire w_dff_A_ZdHL2U0N9_0;
	wire w_dff_A_5qZihNdj5_0;
	wire w_dff_A_4jmLlBEL6_2;
	wire w_dff_A_K7dGq1W42_0;
	wire w_dff_A_78ErQpbl6_0;
	wire w_dff_A_oiP58vZN1_0;
	wire w_dff_A_MBacnCiC5_0;
	wire w_dff_A_TbjA9WKO4_0;
	wire w_dff_A_bZcxRaf15_0;
	wire w_dff_A_BTPkT3Ar5_0;
	wire w_dff_A_P5kiD42M5_0;
	wire w_dff_A_UVRF8aHg7_0;
	wire w_dff_A_YA4PgFku5_0;
	wire w_dff_A_AoLkuKZ61_2;
	wire w_dff_A_ylw4dDrN6_0;
	wire w_dff_A_Xdd7ok6a8_0;
	wire w_dff_A_54dByUgn2_0;
	wire w_dff_A_wFhZF4Ua8_0;
	wire w_dff_A_lFjcVmsP9_0;
	wire w_dff_A_pG7puxD84_0;
	wire w_dff_A_YAvYkCbM4_2;
	wire w_dff_A_NP1UhJWR0_0;
	wire w_dff_A_xmFAMjXS1_0;
	wire w_dff_A_wl6vBbvG5_0;
	wire w_dff_A_n9OBKh7T0_0;
	wire w_dff_A_VYZunaUg1_0;
	wire w_dff_A_KFNQHDik9_0;
	wire w_dff_A_UCB5aFk39_0;
	wire w_dff_A_HgVkLhSQ4_0;
	wire w_dff_A_DSdWtge17_2;
	wire w_dff_A_OKCOEJBq8_0;
	wire w_dff_A_R4F0qpPw9_0;
	wire w_dff_A_MeOEPxwg2_0;
	wire w_dff_A_ldtHwkm14_0;
	wire w_dff_A_BM0TILL55_0;
	wire w_dff_A_09sC8z2F0_0;
	wire w_dff_A_SEI4HRti9_0;
	wire w_dff_A_0KaDLOvR8_0;
	wire w_dff_A_8z21HOci0_0;
	wire w_dff_A_8xMKGdES8_2;
	wire w_dff_A_AGXVRCXs4_0;
	wire w_dff_A_nfZXKJYC6_0;
	wire w_dff_A_9iL3PPUR3_0;
	wire w_dff_A_phLtGnGA2_0;
	wire w_dff_A_IL80sVEE0_0;
	wire w_dff_A_EIST3LLL7_0;
	wire w_dff_A_QMTxobcq3_0;
	wire w_dff_A_8Cu09kgp5_0;
	wire w_dff_A_sJsXddFe9_0;
	wire w_dff_A_gtRm3smp8_0;
	wire w_dff_A_vpF12bp06_2;
	wire w_dff_A_94yHG7RF0_0;
	wire w_dff_A_hzy0GCaL9_0;
	wire w_dff_A_o1lTLpvY3_0;
	wire w_dff_A_N8RH7KoB4_0;
	wire w_dff_A_ptN1hIfg7_0;
	wire w_dff_A_f74DpKmn1_2;
	wire w_dff_A_stUBsX9Y3_0;
	wire w_dff_A_B0VYz8H04_0;
	wire w_dff_A_61KOlwvS7_0;
	wire w_dff_A_oMX9Z7mC0_0;
	wire w_dff_A_l9EQlrUr5_0;
	wire w_dff_A_CndLagRN3_0;
	wire w_dff_A_suQ69fZk6_0;
	wire w_dff_A_saarCmgb1_0;
	wire w_dff_A_ZeBcVuVL1_0;
	wire w_dff_A_E82YkNP98_2;
	wire w_dff_A_NiXddwT25_0;
	wire w_dff_A_yHork1d10_0;
	wire w_dff_A_bDHBIp0h1_0;
	wire w_dff_A_bMyTcRzc2_0;
	wire w_dff_A_XSMtrSdO4_0;
	wire w_dff_A_IKk72nFo2_0;
	wire w_dff_A_IzPlc5I72_0;
	wire w_dff_A_R2TdcyTO5_0;
	wire w_dff_A_IXXnVHd24_2;
	wire w_dff_A_JWVPPvce1_0;
	wire w_dff_A_7qBRIocz2_0;
	wire w_dff_A_N08CUWNV6_0;
	wire w_dff_A_ayycVdQ24_0;
	wire w_dff_A_wCdQqJ2e4_0;
	wire w_dff_A_VdDQx32P4_0;
	wire w_dff_A_hUoNM79V4_0;
	wire w_dff_A_D1HnF7sc8_2;
	wire w_dff_A_uDhLzK2H6_0;
	wire w_dff_A_zpmEnjqy5_0;
	wire w_dff_A_NgIu6MSO1_0;
	wire w_dff_A_BjGsCpof1_0;
	wire w_dff_A_Y8mCYuq03_0;
	wire w_dff_A_DeuY0TwH2_2;
	wire w_dff_A_uYU0wR1Y6_0;
	wire w_dff_A_2U6ZxD2y9_0;
	wire w_dff_A_zXGG6A3l3_0;
	wire w_dff_A_LVO1btpO5_0;
	wire w_dff_A_uSXEqGXQ0_0;
	wire w_dff_A_P6Iyrhfh6_0;
	wire w_dff_A_GBhKIpXW7_0;
	wire w_dff_A_nFhCDl725_0;
	wire w_dff_A_SW2DSLHN4_0;
	wire w_dff_A_tZp0S1964_2;
	wire w_dff_A_yXpZtutY9_0;
	wire w_dff_A_phIhrlIT6_0;
	wire w_dff_A_dIoFMkvd0_0;
	wire w_dff_A_ovASpoot4_0;
	wire w_dff_A_Jv8ZzEsr9_0;
	wire w_dff_A_OdjIXAnE5_0;
	wire w_dff_A_4U8VAeQc6_0;
	wire w_dff_A_rLkYxBE65_0;
	wire w_dff_A_zqQOhykr8_2;
	wire w_dff_A_RNMnEmSD7_0;
	wire w_dff_A_eBa1twq74_0;
	wire w_dff_A_LpVFuWwL7_0;
	wire w_dff_A_rvi8Gjiq1_0;
	wire w_dff_A_KhMthFUg3_0;
	wire w_dff_A_edT1prM79_0;
	wire w_dff_A_xKM4KbzX0_0;
	wire w_dff_A_YI0eKhC97_2;
	wire w_dff_A_ggvozNz20_0;
	wire w_dff_A_Fxtp3UOU7_0;
	wire w_dff_A_gNweMcxI6_0;
	wire w_dff_A_0MkrORxv9_0;
	wire w_dff_A_Yu4al2p14_2;
	wire w_dff_A_h1v9vGOI7_0;
	wire w_dff_A_UUWrqDDP6_0;
	wire w_dff_A_URLnBkPd3_0;
	wire w_dff_A_8OqOhb8R9_0;
	wire w_dff_A_XuJHswCl0_0;
	wire w_dff_A_lSebnpja3_0;
	wire w_dff_A_274ycebk5_0;
	wire w_dff_A_mUdzZVc44_0;
	wire w_dff_A_F0NuwJLN0_1;
	wire w_dff_A_pFZOshJI0_0;
	wire w_dff_A_Gzq185nm1_0;
	wire w_dff_A_60ocbiJO4_0;
	wire w_dff_A_fF6WKln45_0;
	wire w_dff_A_eohpnt6F6_1;
	wire w_dff_A_YGmloTLo6_0;
	wire w_dff_A_AcAIj35K0_0;
	wire w_dff_A_g2g6DWCU6_0;
	wire w_dff_A_G04pAWMR5_0;
	wire w_dff_A_YjWHI2wT6_0;
	wire w_dff_A_X6pQOWnC1_0;
	wire w_dff_A_vCiBwh1v3_0;
	wire w_dff_A_0qERABzF8_1;
	wire w_dff_A_uoxTgMsL9_0;
	wire w_dff_A_qzccYyi69_0;
	wire w_dff_A_cN1iB1Up1_0;
	wire w_dff_A_fiZoD7uK1_0;
	wire w_dff_A_BdgTRnEU4_0;
	wire w_dff_A_h5oOv5FZ8_0;
	wire w_dff_A_be7i5FF67_0;
	wire w_dff_A_ouuG4aRI7_1;
	wire w_dff_A_YE0QG9OJ6_0;
	wire w_dff_A_idd1QvNh1_0;
	wire w_dff_A_2nJ8TReo9_0;
	wire w_dff_A_CP5Ezoe12_0;
	wire w_dff_A_xdhtc1bk9_0;
	wire w_dff_A_cjnk1i2V4_0;
	wire w_dff_A_K6l5DGdU5_0;
	wire w_dff_A_XKSW6wSY4_0;
	wire w_dff_A_YmBmEb0r2_2;
	wire w_dff_A_9CSwpaIN3_0;
	wire w_dff_A_bBtz4Z1h2_0;
	wire w_dff_A_9f2imN564_0;
	wire w_dff_A_6ng2kMVn3_0;
	wire w_dff_A_JlYr2jNi4_0;
	wire w_dff_A_FwuVeJOo5_0;
	wire w_dff_A_znqiFMAL6_0;
	wire w_dff_A_twxvD3j61_0;
	wire w_dff_A_WNTOuDZt5_0;
	wire w_dff_A_kMvYQVCE4_0;
	wire w_dff_A_WtxT0LXO4_0;
	wire w_dff_A_qSKMrMZx9_0;
	wire w_dff_A_T9Ik5eot6_0;
	wire w_dff_A_udz9AGVI8_0;
	wire w_dff_A_vKV8Xpt58_0;
	wire w_dff_A_61pVhAxr4_1;
	wire w_dff_A_seXWpN1q0_0;
	wire w_dff_A_GpPQJ5n18_0;
	wire w_dff_A_clNs3gR33_0;
	wire w_dff_A_TCYtEEkG3_1;
	wire w_dff_A_FPGbjeBh2_0;
	wire w_dff_A_uqdmkj5g6_0;
	wire w_dff_A_M0ScsGu73_0;
	wire w_dff_A_4rUlnZbF1_0;
	wire w_dff_A_gLMnYhGz8_1;
	wire w_dff_A_kpCeFwp51_0;
	wire w_dff_A_nx0MMVWJ4_0;
	wire w_dff_A_KdvHlEDf7_0;
	wire w_dff_A_1Yh8oYJL3_0;
	wire w_dff_A_5vABDvfk0_0;
	wire w_dff_A_LThrxDie4_0;
	wire w_dff_A_p0X5p3Tl8_1;
	wire w_dff_A_NfrbBAt62_0;
	wire w_dff_A_XwmGzCL66_0;
	wire w_dff_A_SIzjbgeo5_0;
	wire w_dff_A_swZFf9zW1_0;
	wire w_dff_A_H9dev3Yc7_0;
	wire w_dff_A_Z5Z00TpU1_0;
	wire w_dff_A_TkidTaBr5_0;
	wire w_dff_A_NjJ1rGZa7_2;
	wire w_dff_A_iV3hby8N7_0;
	wire w_dff_A_pcos2Awu2_0;
	wire w_dff_A_AebEAUfu6_2;
	wire w_dff_A_CeuSNheH4_0;
	wire w_dff_A_PqBZ0Zbl1_0;
	wire w_dff_A_tP90ihO79_2;
	wire w_dff_A_qiwq2d6T7_0;
	wire w_dff_A_MO6P1RqA3_0;
	wire w_dff_A_PP9HAOUA6_0;
	wire w_dff_A_4CRHhEj26_2;
	wire w_dff_A_bJHdQplT0_0;
	wire w_dff_A_NGh9qX0l8_0;
	wire w_dff_A_Ko8nmzGj4_0;
	wire w_dff_A_7Y0fh7EU0_2;
	wire w_dff_A_1whWSXqV6_0;
	wire w_dff_A_VQ8RYErW9_0;
	wire w_dff_A_glMeisTk3_0;
	wire w_dff_A_QI885KOz2_0;
	wire w_dff_A_rFepXOn66_2;
	wire w_dff_A_IyhwQnPo8_0;
	wire w_dff_A_NIgJUmOK0_0;
	wire w_dff_A_HRJtcXab0_0;
	wire w_dff_A_WBcazqRS7_2;
	wire w_dff_A_17Zn9pqn1_0;
	wire w_dff_A_aV5rwXLd1_0;
	wire w_dff_A_8Lwqji8D4_0;
	wire w_dff_A_d2B7YkhN0_2;
	wire w_dff_A_EGtU07CN5_0;
	wire w_dff_A_FC8nWnbz8_0;
	wire w_dff_A_F4ap0ghy6_0;
	wire w_dff_A_CmABijxt0_0;
	wire w_dff_A_7YR1FAlA0_2;
	wire w_dff_A_qekfAvYc7_0;
	wire w_dff_A_lnddDsbh6_0;
	wire w_dff_A_dAjtFB3P0_0;
	wire w_dff_A_2lBg0wOi0_2;
	wire w_dff_A_HaWR7sXJ9_0;
	wire w_dff_A_kddjHfwT8_0;
	wire w_dff_A_hz6kOtRe3_2;
	wire w_dff_A_cKpcwRpm3_0;
	wire w_dff_A_xdlkBVQ79_0;
	wire w_dff_A_RrQzvuqd9_2;
	wire w_dff_A_ij4W11Rm5_0;
	wire w_dff_A_0wj4FSAV3_2;
	wire w_dff_A_D5XrwMvF1_0;
	wire w_dff_A_fwAv4NU81_0;
	wire w_dff_A_8iQwItBN6_0;
	wire w_dff_A_YzzF2G7s5_2;
	wire w_dff_A_pvim20DF8_0;
	wire w_dff_A_H80Avglf3_0;
	wire w_dff_A_o0JBYaTp4_2;
	wire w_dff_A_Hr8xD5Kc0_0;
	wire w_dff_A_MF5afOLJ9_0;
	wire w_dff_A_S3yRiD3O3_2;
	wire w_dff_A_vtmMt5Mp6_0;
	wire w_dff_A_WDxtKaJz2_2;
	wire w_dff_A_V6m1J4yy1_0;
	wire w_dff_A_r0HmbdrS9_0;
	wire w_dff_A_78VkBBwL2_0;
	wire w_dff_A_73tBNL023_2;
	wire w_dff_A_cWNtw4yV7_0;
	wire w_dff_A_XE5T6Wwp1_0;
	wire w_dff_A_WMXgV8dg7_0;
	wire w_dff_A_hMdQYkwo2_2;
	wire w_dff_A_IsWFdUh62_2;
	jnot g0000(.din(w_G545_0[2]),.dout(w_dff_A_qxuufKM28_1),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(G366),.dout(G600_fa_),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(w_dff_A_aQkG8FTE9_1),.clk(gclk));
	jnot g0005(.din(G338),.dout(G611_fa_),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(w_dff_A_Tx7LCMRQ4_2),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(w_dff_A_4t5qomYy6_1),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(w_dff_A_f8vZYw3H0_1),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(w_dff_A_BdUBaggz8_1),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(w_dff_A_O7dZoQl30_1),.clk(gclk));
	jand g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(w_dff_A_A73KRriC2_2),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_RzBELWjC6_1),.dout(w_dff_A_qRvqPe0K0_2),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jor g0016(.dina(w_dff_B_JWqUGSMZ8_0),.dinb(w_n316_0[1]),.dout(w_dff_A_hpXzg0xe9_2),.clk(gclk));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(w_dff_A_ViUahs343_1),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jor g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_),.clk(gclk));
	jor g0022(.dina(w_G809_3[1]),.dinb(w_dff_B_ptZ81eDE6_1),.dout(w_dff_A_TeUGITqX2_2),.clk(gclk));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jor g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330),.clk(gclk));
	jor g0030(.dina(n330),.dinb(w_dff_B_OAjlNXEo5_1),.dout(w_dff_A_he6umlfr2_2),.clk(gclk));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jor g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336),.clk(gclk));
	jor g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(w_dff_A_NGvHq2GN5_2),.clk(gclk));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jor g0038(.dina(w_G809_2[1]),.dinb(w_dff_B_8DrVy7Dt6_1),.dout(w_dff_A_AJ2uePYK9_2),.clk(gclk));
	jand g0039(.dina(w_n326_1[2]),.dinb(G24),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jor g0041(.dina(w_dff_B_qX6aa1gp2_0),.dinb(w_G809_2[0]),.dout(n342),.clk(gclk));
	jor g0042(.dina(n342),.dinb(w_dff_B_bHJaaGt51_1),.dout(n343),.clk(gclk));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(w_dff_A_GFQkePVS7_2),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(G26),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jor g0046(.dina(w_dff_B_HADBglPu0_0),.dinb(w_G809_1[2]),.dout(n347),.clk(gclk));
	jor g0047(.dina(n347),.dinb(w_dff_B_3tVcDugs0_1),.dout(n348),.clk(gclk));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(w_dff_A_ws6qj8t84_2),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(G79),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jor g0051(.dina(w_dff_B_YDEUWMNi4_0),.dinb(w_G809_1[1]),.dout(n352),.clk(gclk));
	jor g0052(.dina(n352),.dinb(w_dff_B_vFmQ5TlV0_1),.dout(n353),.clk(gclk));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(w_dff_A_JaHo8t0x7_2),.clk(gclk));
	jand g0054(.dina(w_n326_0[2]),.dinb(G82),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_G2358_0[2]),.dinb(G80),.dout(n356),.clk(gclk));
	jor g0056(.dina(w_dff_B_wmy6YsLa3_0),.dinb(w_G809_1[0]),.dout(n357),.clk(gclk));
	jor g0057(.dina(n357),.dinb(w_dff_B_f2fpSkCN8_1),.dout(n358),.clk(gclk));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(w_dff_A_bWD9Wu3L6_2),.clk(gclk));
	jnot g0059(.din(w_G308_1[2]),.dout(n360),.clk(gclk));
	jand g0060(.dina(w_n360_0[1]),.dinb(w_G251_4[2]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G479_1[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(w_G308_1[1]),.dinb(w_G248_5[1]),.dout(n363),.clk(gclk));
	jor g0063(.dina(n363),.dinb(w_n362_0[1]),.dout(n364),.clk(gclk));
	jor g0064(.dina(n364),.dinb(n361),.dout(n365),.clk(gclk));
	jnot g0065(.din(w_G254_1[2]),.dout(n366),.clk(gclk));
	jand g0066(.dina(w_n360_0[0]),.dinb(w_n366_4[2]),.dout(n367),.clk(gclk));
	jnot g0067(.din(w_G242_1[2]),.dout(n368),.clk(gclk));
	jand g0068(.dina(w_G308_1[0]),.dinb(w_n368_5[1]),.dout(n369),.clk(gclk));
	jor g0069(.dina(n369),.dinb(w_G479_1[0]),.dout(n370),.clk(gclk));
	jor g0070(.dina(n370),.dinb(n367),.dout(n371),.clk(gclk));
	jand g0071(.dina(n371),.dinb(n365),.dout(n372),.clk(gclk));
	jnot g0072(.din(w_G316_1[2]),.dout(n373),.clk(gclk));
	jand g0073(.dina(w_n373_0[1]),.dinb(w_G251_4[1]),.dout(n374),.clk(gclk));
	jnot g0074(.din(w_G490_1[2]),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_G316_1[1]),.dinb(w_G248_5[0]),.dout(n376),.clk(gclk));
	jor g0076(.dina(n376),.dinb(n375),.dout(n377),.clk(gclk));
	jor g0077(.dina(n377),.dinb(n374),.dout(n378),.clk(gclk));
	jand g0078(.dina(w_n373_0[0]),.dinb(w_n366_4[1]),.dout(n379),.clk(gclk));
	jand g0079(.dina(w_G316_1[0]),.dinb(w_n368_5[0]),.dout(n380),.clk(gclk));
	jor g0080(.dina(n380),.dinb(w_G490_1[1]),.dout(n381),.clk(gclk));
	jor g0081(.dina(n381),.dinb(n379),.dout(n382),.clk(gclk));
	jand g0082(.dina(n382),.dinb(n378),.dout(n383),.clk(gclk));
	jand g0083(.dina(w_n383_0[2]),.dinb(w_n372_0[2]),.dout(n384),.clk(gclk));
	jnot g0084(.din(w_G351_2[2]),.dout(n385),.clk(gclk));
	jnot g0085(.din(G3550),.dout(n386),.clk(gclk));
	jand g0086(.dina(w_n386_4[2]),.dinb(w_n385_1[2]),.dout(n387),.clk(gclk));
	jnot g0087(.din(w_G534_1[2]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G3552_0[1]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n389_4[2]),.dinb(w_G351_2[1]),.dout(n390),.clk(gclk));
	jor g0090(.dina(n390),.dinb(w_n388_1[2]),.dout(n391),.clk(gclk));
	jor g0091(.dina(n391),.dinb(n387),.dout(n392),.clk(gclk));
	jand g0092(.dina(w_G3548_4[2]),.dinb(w_n385_1[1]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3546_5[1]),.dinb(w_G351_2[0]),.dout(n394),.clk(gclk));
	jor g0094(.dina(n394),.dinb(w_G534_1[1]),.dout(n395),.clk(gclk));
	jor g0095(.dina(n395),.dinb(n393),.dout(n396),.clk(gclk));
	jand g0096(.dina(n396),.dinb(n392),.dout(n397),.clk(gclk));
	jnot g0097(.din(w_G293_0[2]),.dout(n398),.clk(gclk));
	jand g0098(.dina(w_n398_0[2]),.dinb(w_n366_4[0]),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G293_0[1]),.dinb(w_n368_4[2]),.dout(n400),.clk(gclk));
	jor g0100(.dina(n400),.dinb(n399),.dout(n401),.clk(gclk));
	jnot g0101(.din(w_G251_4[0]),.dout(n402),.clk(gclk));
	jnot g0102(.din(w_G302_0[2]),.dout(n403),.clk(gclk));
	jand g0103(.dina(w_n403_0[1]),.dinb(w_n402_2[1]),.dout(n404),.clk(gclk));
	jnot g0104(.din(w_G248_4[2]),.dout(n405),.clk(gclk));
	jand g0105(.dina(w_G302_0[1]),.dinb(w_n405_2[1]),.dout(n406),.clk(gclk));
	jor g0106(.dina(n406),.dinb(n404),.dout(n407),.clk(gclk));
	jnot g0107(.din(w_n407_0[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_n408_0[1]),.dinb(w_n401_0[2]),.dout(n409),.clk(gclk));
	jnot g0109(.din(w_G514_1[1]),.dout(n410),.clk(gclk));
	jnot g0110(.din(w_G3546_5[0]),.dout(n411),.clk(gclk));
	jand g0111(.dina(n411),.dinb(w_n410_1[1]),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G3552_0[0]),.dinb(w_G514_1[0]),.dout(n413),.clk(gclk));
	jor g0113(.dina(n413),.dinb(n412),.dout(n414),.clk(gclk));
	jnot g0114(.din(w_n414_0[1]),.dout(n415),.clk(gclk));
	jnot g0115(.din(w_G361_0[2]),.dout(n416),.clk(gclk));
	jand g0116(.dina(w_n416_0[1]),.dinb(w_n402_2[0]),.dout(n417),.clk(gclk));
	jand g0117(.dina(w_G361_0[1]),.dinb(w_n405_2[0]),.dout(n418),.clk(gclk));
	jor g0118(.dina(n418),.dinb(n417),.dout(n419),.clk(gclk));
	jnot g0119(.din(w_n419_0[2]),.dout(n420),.clk(gclk));
	jand g0120(.dina(n420),.dinb(n415),.dout(n421),.clk(gclk));
	jand g0121(.dina(n421),.dinb(n409),.dout(n422),.clk(gclk));
	jand g0122(.dina(n422),.dinb(w_n397_0[1]),.dout(n423),.clk(gclk));
	jnot g0123(.din(w_G324_1[2]),.dout(n424),.clk(gclk));
	jand g0124(.dina(w_n386_4[1]),.dinb(w_n424_2[1]),.dout(n425),.clk(gclk));
	jnot g0125(.din(w_G503_1[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_n389_4[1]),.dinb(w_G324_1[1]),.dout(n427),.clk(gclk));
	jor g0127(.dina(n427),.dinb(w_n426_0[1]),.dout(n428),.clk(gclk));
	jor g0128(.dina(n428),.dinb(n425),.dout(n429),.clk(gclk));
	jand g0129(.dina(w_G3548_4[1]),.dinb(w_n424_2[0]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G3546_4[2]),.dinb(w_G324_1[0]),.dout(n431),.clk(gclk));
	jor g0131(.dina(n431),.dinb(w_G503_1[1]),.dout(n432),.clk(gclk));
	jor g0132(.dina(n432),.dinb(n430),.dout(n433),.clk(gclk));
	jand g0133(.dina(n433),.dinb(n429),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G341_2[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n386_4[0]),.dinb(w_n435_1[2]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G523_1[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n389_4[0]),.dinb(w_G341_2[1]),.dout(n438),.clk(gclk));
	jor g0138(.dina(n438),.dinb(w_n437_1[2]),.dout(n439),.clk(gclk));
	jor g0139(.dina(n439),.dinb(n436),.dout(n440),.clk(gclk));
	jand g0140(.dina(w_G3548_4[0]),.dinb(w_n435_1[1]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3546_4[1]),.dinb(w_G341_2[0]),.dout(n442),.clk(gclk));
	jor g0142(.dina(n442),.dinb(w_G523_1[0]),.dout(n443),.clk(gclk));
	jor g0143(.dina(n443),.dinb(n441),.dout(n444),.clk(gclk));
	jand g0144(.dina(n444),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(w_n434_0[1]),.dout(n446),.clk(gclk));
	jand g0146(.dina(n446),.dinb(n423),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(w_dff_B_kgDrTsHG1_1),.dout(w_dff_A_xzIOgP9N0_2),.clk(gclk));
	jnot g0148(.din(w_G265_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n386_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G400_1[1]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n389_3[2]),.dinb(w_G265_2[0]),.dout(n452),.clk(gclk));
	jor g0152(.dina(n452),.dinb(w_n451_1[1]),.dout(n453),.clk(gclk));
	jor g0153(.dina(n453),.dinb(n450),.dout(n454),.clk(gclk));
	jand g0154(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3546_4[0]),.dinb(w_G265_1[2]),.dout(n456),.clk(gclk));
	jor g0156(.dina(n456),.dinb(w_G400_1[0]),.dout(n457),.clk(gclk));
	jor g0157(.dina(n457),.dinb(n455),.dout(n458),.clk(gclk));
	jand g0158(.dina(n458),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n386_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n389_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jor g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464),.clk(gclk));
	jor g0164(.dina(n464),.dinb(n461),.dout(n465),.clk(gclk));
	jand g0165(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n467),.clk(gclk));
	jor g0167(.dina(n467),.dinb(w_G435_1[1]),.dout(n468),.clk(gclk));
	jor g0168(.dina(n468),.dinb(n466),.dout(n469),.clk(gclk));
	jand g0169(.dina(n469),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G257_2[2]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n386_3[0]),.dinb(w_n471_1[1]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G389_0[2]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n389_3[0]),.dinb(w_G257_2[1]),.dout(n474),.clk(gclk));
	jor g0174(.dina(n474),.dinb(w_n473_1[2]),.dout(n475),.clk(gclk));
	jor g0175(.dina(n475),.dinb(n472),.dout(n476),.clk(gclk));
	jand g0176(.dina(w_G3548_3[0]),.dinb(w_n471_1[0]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3546_3[1]),.dinb(w_G257_2[0]),.dout(n478),.clk(gclk));
	jor g0178(.dina(n478),.dinb(w_G389_0[1]),.dout(n479),.clk(gclk));
	jor g0179(.dina(n479),.dinb(n477),.dout(n480),.clk(gclk));
	jand g0180(.dina(n480),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jand g0182(.dina(n482),.dinb(w_n459_0[1]),.dout(n483),.clk(gclk));
	jnot g0183(.din(w_G273_2[2]),.dout(n484),.clk(gclk));
	jand g0184(.dina(w_n386_2[2]),.dinb(w_n484_1[1]),.dout(n485),.clk(gclk));
	jnot g0185(.din(w_G411_0[2]),.dout(n486),.clk(gclk));
	jand g0186(.dina(w_n389_2[2]),.dinb(w_G273_2[1]),.dout(n487),.clk(gclk));
	jor g0187(.dina(n487),.dinb(w_n486_1[1]),.dout(n488),.clk(gclk));
	jor g0188(.dina(n488),.dinb(n485),.dout(n489),.clk(gclk));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n484_1[0]),.dout(n490),.clk(gclk));
	jand g0190(.dina(w_G3546_3[0]),.dinb(w_G273_2[0]),.dout(n491),.clk(gclk));
	jor g0191(.dina(n491),.dinb(w_G411_0[1]),.dout(n492),.clk(gclk));
	jor g0192(.dina(n492),.dinb(n490),.dout(n493),.clk(gclk));
	jand g0193(.dina(n493),.dinb(n489),.dout(n494),.clk(gclk));
	jnot g0194(.din(w_G281_2[1]),.dout(n495),.clk(gclk));
	jand g0195(.dina(w_n386_2[1]),.dinb(w_n495_1[2]),.dout(n496),.clk(gclk));
	jnot g0196(.din(w_G374_0[2]),.dout(n497),.clk(gclk));
	jand g0197(.dina(w_n389_2[1]),.dinb(w_G281_2[0]),.dout(n498),.clk(gclk));
	jor g0198(.dina(n498),.dinb(w_n497_1[1]),.dout(n499),.clk(gclk));
	jor g0199(.dina(n499),.dinb(n496),.dout(n500),.clk(gclk));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n495_1[1]),.dout(n501),.clk(gclk));
	jand g0201(.dina(w_G3546_2[2]),.dinb(w_G281_1[2]),.dout(n502),.clk(gclk));
	jor g0202(.dina(n502),.dinb(w_G374_0[1]),.dout(n503),.clk(gclk));
	jor g0203(.dina(n503),.dinb(n501),.dout(n504),.clk(gclk));
	jand g0204(.dina(n504),.dinb(n500),.dout(n505),.clk(gclk));
	jand g0205(.dina(w_n505_0[1]),.dinb(w_n494_0[1]),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[2]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n386_2[0]),.dinb(w_n507_1[1]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n389_2[0]),.dinb(w_G218_2[1]),.dout(n510),.clk(gclk));
	jor g0210(.dina(n510),.dinb(w_n509_0[1]),.dout(n511),.clk(gclk));
	jor g0211(.dina(n511),.dinb(n508),.dout(n512),.clk(gclk));
	jand g0212(.dina(w_G3548_2[0]),.dinb(w_n507_1[0]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3546_2[1]),.dinb(w_G218_2[0]),.dout(n514),.clk(gclk));
	jor g0214(.dina(n514),.dinb(w_G468_1[1]),.dout(n515),.clk(gclk));
	jor g0215(.dina(n515),.dinb(n513),.dout(n516),.clk(gclk));
	jand g0216(.dina(n516),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G206_0[2]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_G251_3[2]),.dinb(w_n518_1[1]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G446_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_G248_4[1]),.dinb(w_G206_0[1]),.dout(n521),.clk(gclk));
	jor g0221(.dina(n521),.dinb(n520),.dout(n522),.clk(gclk));
	jor g0222(.dina(n522),.dinb(n519),.dout(n523),.clk(gclk));
	jand g0223(.dina(w_n366_3[2]),.dinb(w_n518_1[0]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_n368_4[1]),.dinb(w_G206_0[0]),.dout(n525),.clk(gclk));
	jor g0225(.dina(n525),.dinb(w_G446_1[1]),.dout(n526),.clk(gclk));
	jor g0226(.dina(n526),.dinb(n524),.dout(n527),.clk(gclk));
	jand g0227(.dina(n527),.dinb(n523),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[2]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G226_2[2]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n386_1[2]),.dinb(w_n530_1[1]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G422_2[1]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n389_1[2]),.dinb(w_G226_2[1]),.dout(n533),.clk(gclk));
	jor g0233(.dina(n533),.dinb(w_n532_0[1]),.dout(n534),.clk(gclk));
	jor g0234(.dina(n534),.dinb(n531),.dout(n535),.clk(gclk));
	jand g0235(.dina(w_G3548_1[2]),.dinb(w_n530_1[0]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3546_2[0]),.dinb(w_G226_2[0]),.dout(n537),.clk(gclk));
	jor g0237(.dina(n537),.dinb(w_G422_2[0]),.dout(n538),.clk(gclk));
	jor g0238(.dina(n538),.dinb(n536),.dout(n539),.clk(gclk));
	jand g0239(.dina(n539),.dinb(n535),.dout(n540),.clk(gclk));
	jnot g0240(.din(w_G210_2[2]),.dout(n541),.clk(gclk));
	jand g0241(.dina(w_n386_1[1]),.dinb(w_n541_1[1]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G457_2[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_n389_1[1]),.dinb(w_G210_2[1]),.dout(n544),.clk(gclk));
	jor g0244(.dina(n544),.dinb(w_n543_0[1]),.dout(n545),.clk(gclk));
	jor g0245(.dina(n545),.dinb(n542),.dout(n546),.clk(gclk));
	jand g0246(.dina(w_G3548_1[1]),.dinb(w_n541_1[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_G3546_1[2]),.dinb(w_G210_2[0]),.dout(n548),.clk(gclk));
	jor g0248(.dina(n548),.dinb(w_G457_2[0]),.dout(n549),.clk(gclk));
	jor g0249(.dina(n549),.dinb(n547),.dout(n550),.clk(gclk));
	jand g0250(.dina(n550),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[1]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(n506),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_dff_B_k2BhBUC50_1),.dout(w_dff_A_zRJ957kz3_2),.clk(gclk));
	jnot g0255(.din(w_G335_4[1]),.dout(n556),.clk(gclk));
	jor g0256(.dina(w_n556_5[1]),.dinb(G241),.dout(n557),.clk(gclk));
	jand g0257(.dina(w_n556_5[0]),.dinb(w_n460_1[0]),.dout(n558),.clk(gclk));
	jnot g0258(.din(n558),.dout(n559),.clk(gclk));
	jand g0259(.dina(n559),.dinb(n557),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_1[1]),.dinb(w_G435_1[0]),.dout(n561),.clk(gclk));
	jnot g0261(.din(w_n561_0[2]),.dout(n562),.clk(gclk));
	jnot g0262(.din(G288),.dout(n563),.clk(gclk));
	jand g0263(.dina(w_G335_4[0]),.dinb(n563),.dout(n564),.clk(gclk));
	jand g0264(.dina(w_n556_4[2]),.dinb(w_n495_1[0]),.dout(n565),.clk(gclk));
	jor g0265(.dina(n565),.dinb(n564),.dout(n566),.clk(gclk));
	jxor g0266(.dina(w_n566_0[2]),.dinb(w_n497_1[0]),.dout(n567),.clk(gclk));
	jor g0267(.dina(w_n556_4[1]),.dinb(w_G280_0[1]),.dout(n568),.clk(gclk));
	jor g0268(.dina(w_G335_3[2]),.dinb(w_G273_1[2]),.dout(n569),.clk(gclk));
	jand g0269(.dina(w_n569_0[1]),.dinb(n568),.dout(n570),.clk(gclk));
	jxor g0270(.dina(w_n570_0[1]),.dinb(w_n486_1[0]),.dout(n571),.clk(gclk));
	jnot g0271(.din(w_n571_1[1]),.dout(n572),.clk(gclk));
	jand g0272(.dina(w_n572_0[2]),.dinb(w_n567_1[1]),.dout(n573),.clk(gclk));
	jnot g0273(.din(n573),.dout(n574),.clk(gclk));
	jor g0274(.dina(w_n556_4[0]),.dinb(G264),.dout(n575),.clk(gclk));
	jor g0275(.dina(w_G335_3[1]),.dinb(w_G257_1[2]),.dout(n576),.clk(gclk));
	jand g0276(.dina(n576),.dinb(n575),.dout(n577),.clk(gclk));
	jxor g0277(.dina(w_n577_0[2]),.dinb(w_n473_1[1]),.dout(n578),.clk(gclk));
	jnot g0278(.din(G272),.dout(n579),.clk(gclk));
	jand g0279(.dina(w_G335_3[0]),.dinb(n579),.dout(n580),.clk(gclk));
	jand g0280(.dina(w_n556_3[2]),.dinb(w_n449_1[0]),.dout(n581),.clk(gclk));
	jor g0281(.dina(n581),.dinb(n580),.dout(n582),.clk(gclk));
	jxor g0282(.dina(w_n582_1[1]),.dinb(w_G400_0[2]),.dout(n583),.clk(gclk));
	jor g0283(.dina(w_n583_1[1]),.dinb(w_n578_0[2]),.dout(n584),.clk(gclk));
	jor g0284(.dina(n584),.dinb(w_n574_0[2]),.dout(n585),.clk(gclk));
	jor g0285(.dina(w_n585_0[1]),.dinb(w_n562_0[1]),.dout(n586),.clk(gclk));
	jnot g0286(.din(n586),.dout(n587),.clk(gclk));
	jor g0287(.dina(w_n556_3[1]),.dinb(G217),.dout(n588),.clk(gclk));
	jor g0288(.dina(w_G335_2[2]),.dinb(w_G210_1[2]),.dout(n589),.clk(gclk));
	jand g0289(.dina(n589),.dinb(n588),.dout(n590),.clk(gclk));
	jxor g0290(.dina(w_n590_1[1]),.dinb(w_G457_1[2]),.dout(n591),.clk(gclk));
	jor g0291(.dina(w_n556_3[0]),.dinb(G209),.dout(n592),.clk(gclk));
	jand g0292(.dina(w_n556_2[2]),.dinb(w_n518_0[2]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jand g0294(.dina(n594),.dinb(n592),.dout(n595),.clk(gclk));
	jxor g0295(.dina(w_n595_1[1]),.dinb(w_G446_1[0]),.dout(n596),.clk(gclk));
	jand g0296(.dina(w_n596_0[2]),.dinb(w_n591_0[1]),.dout(n597),.clk(gclk));
	jor g0297(.dina(w_n556_2[1]),.dinb(G233),.dout(n598),.clk(gclk));
	jor g0298(.dina(w_G335_2[1]),.dinb(w_G226_1[2]),.dout(n599),.clk(gclk));
	jand g0299(.dina(n599),.dinb(n598),.dout(n600),.clk(gclk));
	jxor g0300(.dina(w_n600_1[1]),.dinb(w_G422_1[2]),.dout(n601),.clk(gclk));
	jor g0301(.dina(w_n556_2[0]),.dinb(G225),.dout(n602),.clk(gclk));
	jor g0302(.dina(w_G335_2[0]),.dinb(w_G218_1[2]),.dout(n603),.clk(gclk));
	jand g0303(.dina(n603),.dinb(n602),.dout(n604),.clk(gclk));
	jxor g0304(.dina(w_n604_0[2]),.dinb(w_G468_1[0]),.dout(n605),.clk(gclk));
	jand g0305(.dina(w_n605_2[2]),.dinb(w_n601_0[1]),.dout(n606),.clk(gclk));
	jand g0306(.dina(n606),.dinb(n597),.dout(n607),.clk(gclk));
	jand g0307(.dina(w_n607_0[2]),.dinb(w_n587_1[1]),.dout(w_dff_A_hKGz8qj65_2),.clk(gclk));
	jnot g0308(.din(w_G332_4[2]),.dout(n609),.clk(gclk));
	jor g0309(.dina(w_n609_5[2]),.dinb(w_G331_0[1]),.dout(n610),.clk(gclk));
	jand g0310(.dina(w_n609_5[1]),.dinb(w_n424_1[2]),.dout(n611),.clk(gclk));
	jnot g0311(.din(n611),.dout(n612),.clk(gclk));
	jand g0312(.dina(n612),.dinb(n610),.dout(n613),.clk(gclk));
	jxor g0313(.dina(w_n613_0[2]),.dinb(w_G503_1[0]),.dout(n614),.clk(gclk));
	jor g0314(.dina(w_G358_0[0]),.dinb(w_n609_5[0]),.dout(n615),.clk(gclk));
	jor g0315(.dina(w_G351_1[2]),.dinb(w_G332_4[1]),.dout(n616),.clk(gclk));
	jand g0316(.dina(n616),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_n388_1[1]),.dout(n618),.clk(gclk));
	jand g0318(.dina(w_G600_0),.dinb(w_G332_4[0]),.dout(n619),.clk(gclk));
	jand g0319(.dina(w_n416_0[0]),.dinb(w_n609_4[2]),.dout(n620),.clk(gclk));
	jor g0320(.dina(n620),.dinb(n619),.dout(n621),.clk(gclk));
	jnot g0321(.din(w_n621_2[1]),.dout(n622),.clk(gclk));
	jor g0322(.dina(w_n622_1[1]),.dinb(w_n618_1[1]),.dout(n623),.clk(gclk));
	jand g0323(.dina(w_G611_0),.dinb(w_G332_3[2]),.dout(n624),.clk(gclk));
	jxor g0324(.dina(w_n624_1[2]),.dinb(w_G514_0[2]),.dout(n625),.clk(gclk));
	jor g0325(.dina(w_G348_0[0]),.dinb(w_n609_4[1]),.dout(n626),.clk(gclk));
	jor g0326(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n627),.clk(gclk));
	jand g0327(.dina(n627),.dinb(n626),.dout(n628),.clk(gclk));
	jxor g0328(.dina(w_n628_0[2]),.dinb(w_n437_1[1]),.dout(n629),.clk(gclk));
	jor g0329(.dina(w_n629_0[2]),.dinb(w_n625_0[2]),.dout(n630),.clk(gclk));
	jor g0330(.dina(n630),.dinb(w_n623_0[1]),.dout(n631),.clk(gclk));
	jnot g0331(.din(w_n631_0[1]),.dout(n632),.clk(gclk));
	jand g0332(.dina(n632),.dinb(w_n614_2[1]),.dout(n633),.clk(gclk));
	jand g0333(.dina(w_G332_3[0]),.dinb(w_G593_0),.dout(n634),.clk(gclk));
	jand g0334(.dina(w_n609_4[0]),.dinb(w_n398_0[1]),.dout(n635),.clk(gclk));
	jor g0335(.dina(n635),.dinb(n634),.dout(n636),.clk(gclk));
	jor g0336(.dina(w_n609_3[2]),.dinb(G307),.dout(n637),.clk(gclk));
	jand g0337(.dina(w_n609_3[1]),.dinb(w_n403_0[0]),.dout(n638),.clk(gclk));
	jnot g0338(.din(n638),.dout(n639),.clk(gclk));
	jand g0339(.dina(n639),.dinb(n637),.dout(n640),.clk(gclk));
	jnot g0340(.din(w_n640_1[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n641_0[1]),.dinb(w_n636_1[1]),.dout(n642),.clk(gclk));
	jor g0342(.dina(w_n609_3[0]),.dinb(G315),.dout(n643),.clk(gclk));
	jor g0343(.dina(w_G332_2[2]),.dinb(w_G308_0[2]),.dout(n644),.clk(gclk));
	jand g0344(.dina(n644),.dinb(n643),.dout(n645),.clk(gclk));
	jxor g0345(.dina(w_n645_0[2]),.dinb(w_G479_0[2]),.dout(n646),.clk(gclk));
	jor g0346(.dina(w_n609_2[2]),.dinb(G323),.dout(n647),.clk(gclk));
	jor g0347(.dina(w_G332_2[1]),.dinb(w_G316_0[2]),.dout(n648),.clk(gclk));
	jand g0348(.dina(n648),.dinb(n647),.dout(n649),.clk(gclk));
	jxor g0349(.dina(w_n649_1[1]),.dinb(w_G490_1[0]),.dout(n650),.clk(gclk));
	jand g0350(.dina(w_n650_0[1]),.dinb(w_n646_0[2]),.dout(n651),.clk(gclk));
	jand g0351(.dina(w_n651_1[1]),.dinb(w_n642_0[1]),.dout(n652),.clk(gclk));
	jand g0352(.dina(w_n652_0[1]),.dinb(w_n633_1[1]),.dout(w_dff_A_CvoF0cw43_2),.clk(gclk));
	jxor g0353(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n654),.clk(gclk));
	jxor g0354(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n655),.clk(gclk));
	jxor g0355(.dina(n655),.dinb(n654),.dout(n656),.clk(gclk));
	jxor g0356(.dina(w_G369_0[1]),.dinb(w_G361_0[0]),.dout(n657),.clk(gclk));
	jxor g0357(.dina(n657),.dinb(w_n424_1[1]),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_G302_0[0]),.dinb(w_n398_0[0]),.dout(n659),.clk(gclk));
	jxor g0359(.dina(n659),.dinb(n658),.dout(n660),.clk(gclk));
	jxor g0360(.dina(n660),.dinb(n656),.dout(n661),.clk(gclk));
	jnot g0361(.din(w_n661_0[1]),.dout(w_dff_A_gwSMvLaq9_1),.clk(gclk));
	jxor g0362(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G273_1[1]),.dinb(w_G265_1[1]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(n663),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(n667),.dinb(n666),.dout(n668),.clk(gclk));
	jxor g0368(.dina(w_G210_1[1]),.dinb(w_n518_0[1]),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n668),.dout(n670),.clk(gclk));
	jxor g0370(.dina(n670),.dinb(n665),.dout(n671),.clk(gclk));
	jnot g0371(.din(w_n671_0[1]),.dout(w_dff_A_ByIlIlBF7_1),.clk(gclk));
	jnot g0372(.din(w_n560_1[0]),.dout(n673),.clk(gclk));
	jand g0373(.dina(n673),.dinb(w_n462_0[1]),.dout(n674),.clk(gclk));
	jnot g0374(.din(n674),.dout(n675),.clk(gclk));
	jand g0375(.dina(w_n560_0[2]),.dinb(w_G435_0[2]),.dout(n676),.clk(gclk));
	jnot g0376(.din(w_n577_0[1]),.dout(n677),.clk(gclk));
	jand g0377(.dina(w_n677_0[1]),.dinb(w_n473_1[0]),.dout(n678),.clk(gclk));
	jor g0378(.dina(w_n677_0[0]),.dinb(w_n473_0[2]),.dout(n679),.clk(gclk));
	jand g0379(.dina(w_n582_1[0]),.dinb(w_n451_1[0]),.dout(n680),.clk(gclk));
	jor g0380(.dina(w_n566_0[1]),.dinb(w_n497_0[2]),.dout(n681),.clk(gclk));
	jor g0381(.dina(w_n571_1[0]),.dinb(w_n681_2[1]),.dout(n682),.clk(gclk));
	jnot g0382(.din(w_G280_0[0]),.dout(n683),.clk(gclk));
	jand g0383(.dina(w_G335_1[2]),.dinb(n683),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n569_0[0]),.dout(n685),.clk(gclk));
	jor g0385(.dina(n685),.dinb(n684),.dout(n686),.clk(gclk));
	jor g0386(.dina(n686),.dinb(w_n486_0[2]),.dout(n687),.clk(gclk));
	jor g0387(.dina(w_n582_0[2]),.dinb(w_n451_0[2]),.dout(n688),.clk(gclk));
	jand g0388(.dina(n688),.dinb(w_n687_0[2]),.dout(n689),.clk(gclk));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n682_0[1]),.dout(n690),.clk(gclk));
	jor g0390(.dina(n690),.dinb(w_n680_0[1]),.dout(n691),.clk(gclk));
	jand g0391(.dina(w_n691_0[2]),.dinb(w_n679_0[1]),.dout(n692),.clk(gclk));
	jor g0392(.dina(n692),.dinb(w_n678_0[1]),.dout(n693),.clk(gclk));
	jnot g0393(.din(w_n693_0[2]),.dout(n694),.clk(gclk));
	jor g0394(.dina(n694),.dinb(n676),.dout(n695),.clk(gclk));
	jand g0395(.dina(n695),.dinb(n675),.dout(n696),.clk(gclk));
	jand g0396(.dina(w_n696_0[2]),.dinb(w_n607_0[1]),.dout(n697),.clk(gclk));
	jand g0397(.dina(w_n595_1[0]),.dinb(w_G446_0[2]),.dout(n698),.clk(gclk));
	jor g0398(.dina(w_n595_0[2]),.dinb(w_G446_0[1]),.dout(n699),.clk(gclk));
	jor g0399(.dina(w_n590_1[0]),.dinb(w_G457_1[1]),.dout(n700),.clk(gclk));
	jand g0400(.dina(w_n590_0[2]),.dinb(w_G457_1[0]),.dout(n701),.clk(gclk));
	jand g0401(.dina(w_n604_0[1]),.dinb(w_G468_0[2]),.dout(n702),.clk(gclk));
	jand g0402(.dina(w_n600_1[0]),.dinb(w_G422_1[1]),.dout(n703),.clk(gclk));
	jand g0403(.dina(w_n605_2[1]),.dinb(w_n703_0[2]),.dout(n704),.clk(gclk));
	jor g0404(.dina(n704),.dinb(w_n702_0[1]),.dout(n705),.clk(gclk));
	jor g0405(.dina(w_n705_0[1]),.dinb(n701),.dout(n706),.clk(gclk));
	jand g0406(.dina(w_n706_0[1]),.dinb(w_n700_0[1]),.dout(n707),.clk(gclk));
	jand g0407(.dina(w_n707_0[2]),.dinb(n699),.dout(n708),.clk(gclk));
	jor g0408(.dina(n708),.dinb(n698),.dout(n709),.clk(gclk));
	jor g0409(.dina(w_n709_0[1]),.dinb(w_n697_0[1]),.dout(w_dff_A_svarlViU6_2),.clk(gclk));
	jand g0410(.dina(w_n613_0[1]),.dinb(w_G503_0[2]),.dout(n711),.clk(gclk));
	jor g0411(.dina(w_n624_1[1]),.dinb(w_n410_1[0]),.dout(n712),.clk(gclk));
	jand g0412(.dina(w_n624_1[0]),.dinb(w_n410_0[2]),.dout(n713),.clk(gclk));
	jand g0413(.dina(w_G599_0),.dinb(w_G332_2[0]),.dout(n714),.clk(gclk));
	jand g0414(.dina(w_n435_1[0]),.dinb(w_n609_2[1]),.dout(n715),.clk(gclk));
	jor g0415(.dina(n715),.dinb(n714),.dout(n716),.clk(gclk));
	jand g0416(.dina(w_n716_0[1]),.dinb(w_n437_1[0]),.dout(n717),.clk(gclk));
	jand g0417(.dina(w_G612_0),.dinb(w_G332_1[2]),.dout(n718),.clk(gclk));
	jand g0418(.dina(w_n385_1[0]),.dinb(w_n609_2[0]),.dout(n719),.clk(gclk));
	jor g0419(.dina(n719),.dinb(n718),.dout(n720),.clk(gclk));
	jand g0420(.dina(w_n720_0[1]),.dinb(w_n388_1[0]),.dout(n721),.clk(gclk));
	jor g0421(.dina(w_n621_2[0]),.dinb(w_n721_0[2]),.dout(n722),.clk(gclk));
	jor g0422(.dina(w_n720_0[0]),.dinb(w_n388_0[2]),.dout(n723),.clk(gclk));
	jor g0423(.dina(w_n716_0[0]),.dinb(w_n437_0[2]),.dout(n724),.clk(gclk));
	jand g0424(.dina(n724),.dinb(w_n723_0[1]),.dout(n725),.clk(gclk));
	jand g0425(.dina(n725),.dinb(n722),.dout(n726),.clk(gclk));
	jor g0426(.dina(w_n726_0[1]),.dinb(w_n717_0[2]),.dout(n727),.clk(gclk));
	jor g0427(.dina(w_n727_0[2]),.dinb(w_dff_B_Q7B98Heb2_1),.dout(n728),.clk(gclk));
	jand g0428(.dina(n728),.dinb(w_dff_B_xpRPAu6s1_1),.dout(n729),.clk(gclk));
	jnot g0429(.din(w_n729_1[1]),.dout(n730),.clk(gclk));
	jand g0430(.dina(n730),.dinb(w_n614_2[0]),.dout(n731),.clk(gclk));
	jor g0431(.dina(n731),.dinb(w_dff_B_qNVll6yt7_1),.dout(n732),.clk(gclk));
	jand g0432(.dina(w_n732_0[2]),.dinb(w_n651_1[0]),.dout(n733),.clk(gclk));
	jnot g0433(.din(w_n642_0[0]),.dout(n734),.clk(gclk));
	jnot g0434(.din(w_n645_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[1]),.dinb(w_n362_0[0]),.dout(n736),.clk(gclk));
	jnot g0436(.din(w_n736_0[1]),.dout(n737),.clk(gclk));
	jand g0437(.dina(w_n645_0[0]),.dinb(w_G479_0[1]),.dout(n738),.clk(gclk));
	jand g0438(.dina(w_n649_1[0]),.dinb(w_G490_0[2]),.dout(n739),.clk(gclk));
	jor g0439(.dina(w_n739_1[1]),.dinb(n738),.dout(n740),.clk(gclk));
	jand g0440(.dina(w_n740_0[1]),.dinb(n737),.dout(n741),.clk(gclk));
	jor g0441(.dina(w_n741_0[1]),.dinb(n734),.dout(n742),.clk(gclk));
	jor g0442(.dina(w_n742_0[1]),.dinb(w_n733_0[1]),.dout(w_dff_A_RURQqRW80_2),.clk(gclk));
	jnot g0443(.din(w_G54_0[1]),.dout(n744),.clk(gclk));
	jxor g0444(.dina(w_n621_1[2]),.dinb(w_n744_1[2]),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_G4092_1[2]),.dout(n746),.clk(gclk));
	jand g0446(.dina(w_n746_1[2]),.dinb(w_G4091_2[2]),.dout(n747),.clk(gclk));
	jnot g0447(.din(w_n747_3[2]),.dout(n748),.clk(gclk));
	jor g0448(.dina(w_n748_4[1]),.dinb(n745),.dout(n749),.clk(gclk));
	jnot g0449(.din(w_G4091_2[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n746_1[1]),.dinb(w_n750_1[1]),.dout(n751),.clk(gclk));
	jand g0451(.dina(w_n751_2[1]),.dinb(w_n419_0[1]),.dout(n752),.clk(gclk));
	jand g0452(.dina(w_G4092_1[1]),.dinb(w_n750_1[0]),.dout(n753),.clk(gclk));
	jand g0453(.dina(w_n753_8[1]),.dinb(G131),.dout(n754),.clk(gclk));
	jor g0454(.dina(n754),.dinb(n752),.dout(n755),.clk(gclk));
	jnot g0455(.din(n755),.dout(n756),.clk(gclk));
	jand g0456(.dina(n756),.dinb(w_dff_B_0wHZ84El8_1),.dout(G822_fa_),.clk(gclk));
	jnot g0457(.din(w_n618_1[0]),.dout(n758),.clk(gclk));
	jand g0458(.dina(w_n621_1[1]),.dinb(w_n744_1[1]),.dout(n759),.clk(gclk));
	jnot g0459(.din(w_n759_0[1]),.dout(n760),.clk(gclk));
	jand g0460(.dina(w_n760_0[1]),.dinb(n758),.dout(n761),.clk(gclk));
	jand g0461(.dina(w_n759_0[0]),.dinb(w_n618_0[2]),.dout(n762),.clk(gclk));
	jor g0462(.dina(n762),.dinb(w_n748_4[0]),.dout(n763),.clk(gclk));
	jor g0463(.dina(n763),.dinb(w_n761_0[1]),.dout(n764),.clk(gclk));
	jnot g0464(.din(w_n751_2[0]),.dout(n765),.clk(gclk));
	jor g0465(.dina(w_n765_5[2]),.dinb(w_n397_0[0]),.dout(n766),.clk(gclk));
	jand g0466(.dina(w_n753_8[0]),.dinb(G129),.dout(n767),.clk(gclk));
	jnot g0467(.din(n767),.dout(n768),.clk(gclk));
	jand g0468(.dina(n768),.dinb(n766),.dout(n769),.clk(gclk));
	jand g0469(.dina(n769),.dinb(n764),.dout(G838_fa_),.clk(gclk));
	jxor g0470(.dina(w_n567_1[0]),.dinb(w_G4_1[1]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n771_0[1]),.dinb(w_n747_3[1]),.dout(n772),.clk(gclk));
	jnot g0472(.din(n772),.dout(n773),.clk(gclk));
	jor g0473(.dina(w_n765_5[1]),.dinb(w_n505_0[0]),.dout(n774),.clk(gclk));
	jand g0474(.dina(w_n753_7[2]),.dinb(G117),.dout(n775),.clk(gclk));
	jnot g0475(.din(n775),.dout(n776),.clk(gclk));
	jand g0476(.dina(n776),.dinb(n774),.dout(n777),.clk(gclk));
	jand g0477(.dina(n777),.dinb(n773),.dout(G861_fa_),.clk(gclk));
	jnot g0478(.din(w_n636_1[0]),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n633_1[0]),.dinb(w_G54_0[0]),.dout(n780),.clk(gclk));
	jor g0480(.dina(w_dff_B_6RQQT2QQ7_0),.dinb(w_n732_0[1]),.dout(n781),.clk(gclk));
	jand g0481(.dina(w_n781_0[2]),.dinb(w_n651_0[2]),.dout(n782),.clk(gclk));
	jor g0482(.dina(n782),.dinb(w_n741_0[0]),.dout(n783),.clk(gclk));
	jnot g0483(.din(w_n783_1[1]),.dout(n784),.clk(gclk));
	jor g0484(.dina(n784),.dinb(w_n779_0[1]),.dout(n785),.clk(gclk));
	jxor g0485(.dina(w_n640_1[1]),.dinb(w_n779_0[0]),.dout(n786),.clk(gclk));
	jnot g0486(.din(w_n786_0[1]),.dout(n787),.clk(gclk));
	jor g0487(.dina(w_n787_0[1]),.dinb(w_n783_1[0]),.dout(n788),.clk(gclk));
	jand g0488(.dina(w_dff_B_b8gTI8kT6_0),.dinb(n785),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n789_0[2]),.dout(w_dff_A_FnIaWamW8_1),.clk(gclk));
	jnot g0490(.din(w_G861_0),.dout(n791),.clk(gclk));
	jnot g0491(.din(w_G4087_0[2]),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_G4088_0[2]),.dinb(w_n792_0[1]),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n793_4[1]),.dinb(w_n791_1[1]),.dout(n794),.clk(gclk));
	jnot g0494(.din(w_G822_0),.dout(n795),.clk(gclk));
	jnot g0495(.din(w_G4088_0[1]),.dout(n796),.clk(gclk));
	jand g0496(.dina(w_n796_0[1]),.dinb(w_n792_0[0]),.dout(n797),.clk(gclk));
	jand g0497(.dina(w_n797_4[1]),.dinb(w_n795_1[1]),.dout(n798),.clk(gclk));
	jand g0498(.dina(w_n796_0[0]),.dinb(w_G4087_0[1]),.dout(n799),.clk(gclk));
	jand g0499(.dina(w_n799_4[1]),.dinb(w_G11_0[1]),.dout(n800),.clk(gclk));
	jand g0500(.dina(w_G4088_0[0]),.dinb(w_G4087_0[0]),.dout(n801),.clk(gclk));
	jand g0501(.dina(w_n801_4[1]),.dinb(w_G61_0[1]),.dout(n802),.clk(gclk));
	jor g0502(.dina(n802),.dinb(n800),.dout(n803),.clk(gclk));
	jor g0503(.dina(w_dff_B_o5YSYmXM7_0),.dinb(n798),.dout(n804),.clk(gclk));
	jor g0504(.dina(n804),.dinb(n794),.dout(w_dff_A_rihHI8OF6_2),.clk(gclk));
	jand g0505(.dina(w_n729_1[0]),.dinb(w_n631_0[0]),.dout(n806),.clk(gclk));
	jand g0506(.dina(w_n729_0[2]),.dinb(w_n744_1[0]),.dout(n807),.clk(gclk));
	jor g0507(.dina(n807),.dinb(w_n806_0[2]),.dout(n808),.clk(gclk));
	jxor g0508(.dina(n808),.dinb(w_n614_1[2]),.dout(n809),.clk(gclk));
	jor g0509(.dina(w_n809_0[1]),.dinb(w_n748_3[2]),.dout(n810),.clk(gclk));
	jor g0510(.dina(w_n765_5[0]),.dinb(w_n434_0[0]),.dout(n811),.clk(gclk));
	jand g0511(.dina(w_n753_7[1]),.dinb(G52),.dout(n812),.clk(gclk));
	jnot g0512(.din(n812),.dout(n813),.clk(gclk));
	jand g0513(.dina(n813),.dinb(n811),.dout(n814),.clk(gclk));
	jand g0514(.dina(w_dff_B_hhbfhIuz9_0),.dinb(n810),.dout(G832_fa_),.clk(gclk));
	jnot g0515(.din(w_n625_0[1]),.dout(n816),.clk(gclk));
	jand g0516(.dina(w_n727_0[1]),.dinb(w_n744_0[2]),.dout(n817),.clk(gclk));
	jand g0517(.dina(w_n726_0[0]),.dinb(w_n623_0[0]),.dout(n818),.clk(gclk));
	jor g0518(.dina(n818),.dinb(w_n717_0[1]),.dout(n819),.clk(gclk));
	jor g0519(.dina(w_n819_0[1]),.dinb(n817),.dout(n820),.clk(gclk));
	jxor g0520(.dina(n820),.dinb(w_dff_B_w6uc7q442_1),.dout(n821),.clk(gclk));
	jor g0521(.dina(w_n821_0[1]),.dinb(w_n748_3[1]),.dout(n822),.clk(gclk));
	jand g0522(.dina(w_n751_1[2]),.dinb(w_n414_0[0]),.dout(n823),.clk(gclk));
	jand g0523(.dina(w_n753_7[0]),.dinb(G130),.dout(n824),.clk(gclk));
	jor g0524(.dina(n824),.dinb(n823),.dout(n825),.clk(gclk));
	jnot g0525(.din(n825),.dout(n826),.clk(gclk));
	jand g0526(.dina(w_dff_B_WIS3tm177_0),.dinb(n822),.dout(G834_fa_),.clk(gclk));
	jor g0527(.dina(w_n617_1[0]),.dinb(w_G534_1[0]),.dout(n828),.clk(gclk));
	jand g0528(.dina(w_n617_0[2]),.dinb(w_G534_0[2]),.dout(n829),.clk(gclk));
	jor g0529(.dina(w_n760_0[0]),.dinb(w_n829_0[1]),.dout(n830),.clk(gclk));
	jand g0530(.dina(n830),.dinb(w_n828_0[2]),.dout(n831),.clk(gclk));
	jxor g0531(.dina(n831),.dinb(w_n629_0[1]),.dout(n832),.clk(gclk));
	jor g0532(.dina(w_n832_0[1]),.dinb(w_n748_3[0]),.dout(n833),.clk(gclk));
	jor g0533(.dina(w_n765_4[2]),.dinb(w_n445_0[0]),.dout(n834),.clk(gclk));
	jand g0534(.dina(w_n753_6[2]),.dinb(G119),.dout(n835),.clk(gclk));
	jnot g0535(.din(n835),.dout(n836),.clk(gclk));
	jand g0536(.dina(n836),.dinb(n834),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_dff_B_WuXpcJCp9_0),.dinb(n833),.dout(G836_fa_),.clk(gclk));
	jnot g0538(.din(w_G4090_0[2]),.dout(n839),.clk(gclk));
	jand g0539(.dina(w_n839_0[1]),.dinb(w_G4089_0[2]),.dout(n840),.clk(gclk));
	jand g0540(.dina(w_n840_4[1]),.dinb(w_n791_1[0]),.dout(n841),.clk(gclk));
	jnot g0541(.din(w_G4089_0[1]),.dout(n842),.clk(gclk));
	jand g0542(.dina(w_n839_0[0]),.dinb(w_n842_0[1]),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n843_4[1]),.dinb(w_n795_1[0]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_G4090_0[1]),.dinb(w_n842_0[0]),.dout(n845),.clk(gclk));
	jand g0545(.dina(w_n845_4[1]),.dinb(w_G11_0[0]),.dout(n846),.clk(gclk));
	jand g0546(.dina(w_G4090_0[0]),.dinb(w_G4089_0[0]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_4[1]),.dinb(w_G61_0[0]),.dout(n848),.clk(gclk));
	jor g0548(.dina(n848),.dinb(n846),.dout(n849),.clk(gclk));
	jor g0549(.dina(w_dff_B_BaO8iXGJ0_0),.dinb(n844),.dout(n850),.clk(gclk));
	jor g0550(.dina(n850),.dinb(n841),.dout(w_dff_A_89q19c2f0_2),.clk(gclk));
	jnot g0551(.din(w_n678_0[0]),.dout(n852),.clk(gclk));
	jnot g0552(.din(w_n679_0[0]),.dout(n853),.clk(gclk));
	jor g0553(.dina(w_n583_1[0]),.dinb(w_n574_0[1]),.dout(n854),.clk(gclk));
	jand g0554(.dina(n854),.dinb(w_n691_0[1]),.dout(n855),.clk(gclk));
	jnot g0555(.din(w_n855_0[1]),.dout(n856),.clk(gclk));
	jnot g0556(.din(w_n691_0[0]),.dout(n857),.clk(gclk));
	jor g0557(.dina(w_n857_0[1]),.dinb(w_G4_1[0]),.dout(n858),.clk(gclk));
	jand g0558(.dina(n858),.dinb(w_n856_0[1]),.dout(n859),.clk(gclk));
	jor g0559(.dina(w_n859_0[1]),.dinb(w_n853_0[1]),.dout(n860),.clk(gclk));
	jand g0560(.dina(n860),.dinb(n852),.dout(n861),.clk(gclk));
	jxor g0561(.dina(n861),.dinb(w_n562_0[0]),.dout(n862),.clk(gclk));
	jor g0562(.dina(w_n862_0[1]),.dinb(w_n748_2[2]),.dout(n863),.clk(gclk));
	jor g0563(.dina(w_n765_4[1]),.dinb(w_n470_0[0]),.dout(n864),.clk(gclk));
	jand g0564(.dina(w_n753_6[1]),.dinb(G122),.dout(n865),.clk(gclk));
	jnot g0565(.din(n865),.dout(n866),.clk(gclk));
	jand g0566(.dina(n866),.dinb(n864),.dout(n867),.clk(gclk));
	jand g0567(.dina(n867),.dinb(n863),.dout(G871_fa_),.clk(gclk));
	jxor g0568(.dina(w_n859_0[0]),.dinb(w_n578_0[1]),.dout(n869),.clk(gclk));
	jor g0569(.dina(w_n869_0[1]),.dinb(w_n748_2[1]),.dout(n870),.clk(gclk));
	jor g0570(.dina(w_n765_4[0]),.dinb(w_n481_0[0]),.dout(n871),.clk(gclk));
	jand g0571(.dina(w_n753_6[0]),.dinb(G128),.dout(n872),.clk(gclk));
	jnot g0572(.din(n872),.dout(n873),.clk(gclk));
	jand g0573(.dina(n873),.dinb(n871),.dout(n874),.clk(gclk));
	jand g0574(.dina(n874),.dinb(n870),.dout(G873_fa_),.clk(gclk));
	jand g0575(.dina(w_n567_0[2]),.dinb(w_G4_0[2]),.dout(n876),.clk(gclk));
	jnot g0576(.din(n876),.dout(n877),.clk(gclk));
	jand g0577(.dina(w_n877_0[1]),.dinb(w_n681_2[0]),.dout(n878),.clk(gclk));
	jor g0578(.dina(n878),.dinb(w_n571_0[2]),.dout(n879),.clk(gclk));
	jand g0579(.dina(w_n879_0[1]),.dinb(w_n687_0[1]),.dout(n880),.clk(gclk));
	jxor g0580(.dina(n880),.dinb(w_n583_0[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n881_0[1]),.dinb(w_n747_3[0]),.dout(n882),.clk(gclk));
	jnot g0582(.din(n882),.dout(n883),.clk(gclk));
	jor g0583(.dina(w_n765_3[2]),.dinb(w_n459_0[0]),.dout(n884),.clk(gclk));
	jand g0584(.dina(w_n753_5[2]),.dinb(G127),.dout(n885),.clk(gclk));
	jnot g0585(.din(n885),.dout(n886),.clk(gclk));
	jand g0586(.dina(n886),.dinb(n884),.dout(n887),.clk(gclk));
	jand g0587(.dina(n887),.dinb(n883),.dout(G875_fa_),.clk(gclk));
	jand g0588(.dina(w_n571_0[1]),.dinb(w_n681_1[2]),.dout(n889),.clk(gclk));
	jand g0589(.dina(n889),.dinb(w_n877_0[0]),.dout(n890),.clk(gclk));
	jnot g0590(.din(n890),.dout(n891),.clk(gclk));
	jand g0591(.dina(n891),.dinb(w_n879_0[0]),.dout(n892),.clk(gclk));
	jand g0592(.dina(w_n892_0[1]),.dinb(w_n747_2[2]),.dout(n893),.clk(gclk));
	jnot g0593(.din(n893),.dout(n894),.clk(gclk));
	jor g0594(.dina(w_n765_3[1]),.dinb(w_n494_0[0]),.dout(n895),.clk(gclk));
	jand g0595(.dina(w_n753_5[1]),.dinb(G126),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jand g0597(.dina(n897),.dinb(n895),.dout(n898),.clk(gclk));
	jand g0598(.dina(n898),.dinb(n894),.dout(G877_fa_),.clk(gclk));
	jxor g0599(.dina(w_n649_0[2]),.dinb(w_n735_0[0]),.dout(n900),.clk(gclk));
	jxor g0600(.dina(n900),.dinb(w_n786_0[0]),.dout(n901),.clk(gclk));
	jxor g0601(.dina(n901),.dinb(w_n621_1[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_G369_0[0]),.dinb(w_n609_1[2]),.dout(n903),.clk(gclk));
	jand g0603(.dina(G372),.dinb(w_G332_1[1]),.dout(n904),.clk(gclk));
	jor g0604(.dina(n904),.dinb(n903),.dout(n905),.clk(gclk));
	jxor g0605(.dina(n905),.dinb(w_n617_0[1]),.dout(n906),.clk(gclk));
	jxor g0606(.dina(n906),.dinb(w_n628_0[1]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_G331_0[0]),.dout(n908),.clk(gclk));
	jand g0608(.dina(w_n624_0[2]),.dinb(w_dff_B_Xa60deEF0_1),.dout(n909),.clk(gclk));
	jnot g0609(.din(w_n624_0[1]),.dout(n910),.clk(gclk));
	jand g0610(.dina(w_dff_B_QTcJ8GD28_0),.dinb(w_n613_0[0]),.dout(n911),.clk(gclk));
	jor g0611(.dina(n911),.dinb(w_dff_B_sllcrRqo5_1),.dout(n912),.clk(gclk));
	jxor g0612(.dina(n912),.dinb(w_dff_B_dS2amFQa1_1),.dout(n913),.clk(gclk));
	jxor g0613(.dina(n913),.dinb(n902),.dout(n914),.clk(gclk));
	jnot g0614(.din(w_n914_0[1]),.dout(w_dff_A_DRK3FxjO7_1),.clk(gclk));
	jxor g0615(.dina(w_n577_0[0]),.dinb(w_n566_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n582_0[1]),.dinb(w_n570_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(n917),.dinb(n916),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_n590_0[1]),.dout(n919),.clk(gclk));
	jand g0619(.dina(w_n556_1[2]),.dinb(w_G289_0[0]),.dout(n920),.clk(gclk));
	jand g0620(.dina(w_G335_1[1]),.dinb(G292),.dout(n921),.clk(gclk));
	jor g0621(.dina(n921),.dinb(n920),.dout(n922),.clk(gclk));
	jxor g0622(.dina(n922),.dinb(w_n600_0[2]),.dout(n923),.clk(gclk));
	jxor g0623(.dina(n923),.dinb(w_n560_0[1]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n604_0[0]),.dinb(w_n595_0[1]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jxor g0626(.dina(n926),.dinb(n919),.dout(G1000_fa_),.clk(gclk));
	jnot g0627(.din(w_n596_0[1]),.dout(n928),.clk(gclk));
	jnot g0628(.din(w_n707_0[1]),.dout(n929),.clk(gclk));
	jnot g0629(.din(w_n700_0[0]),.dout(n930),.clk(gclk));
	jnot g0630(.din(w_n605_2[0]),.dout(n931),.clk(gclk));
	jnot g0631(.din(w_n601_0[0]),.dout(n932),.clk(gclk));
	jnot g0632(.din(w_n696_0[1]),.dout(n933),.clk(gclk));
	jand g0633(.dina(w_n587_1[0]),.dinb(w_G4_0[1]),.dout(n934),.clk(gclk));
	jnot g0634(.din(n934),.dout(n935),.clk(gclk));
	jand g0635(.dina(n935),.dinb(n933),.dout(n936),.clk(gclk));
	jor g0636(.dina(w_n936_0[2]),.dinb(w_n932_0[1]),.dout(n937),.clk(gclk));
	jor g0637(.dina(n937),.dinb(n931),.dout(n938),.clk(gclk));
	jor g0638(.dina(w_n938_0[1]),.dinb(w_n930_0[2]),.dout(n939),.clk(gclk));
	jand g0639(.dina(n939),.dinb(n929),.dout(n940),.clk(gclk));
	jxor g0640(.dina(n940),.dinb(w_n928_0[1]),.dout(n941),.clk(gclk));
	jnot g0641(.din(w_n941_0[1]),.dout(n942),.clk(gclk));
	jnot g0642(.din(w_n591_0[0]),.dout(n943),.clk(gclk));
	jnot g0643(.din(w_n705_0[0]),.dout(n944),.clk(gclk));
	jand g0644(.dina(w_n938_0[0]),.dinb(w_n944_0[1]),.dout(n945),.clk(gclk));
	jxor g0645(.dina(n945),.dinb(w_n943_0[1]),.dout(n946),.clk(gclk));
	jnot g0646(.din(w_n946_0[1]),.dout(n947),.clk(gclk));
	jor g0647(.dina(w_n600_0[1]),.dinb(w_G422_1[0]),.dout(n948),.clk(gclk));
	jnot g0648(.din(w_n948_0[2]),.dout(n949),.clk(gclk));
	jnot g0649(.din(w_n703_0[1]),.dout(n950),.clk(gclk));
	jand g0650(.dina(w_n936_0[1]),.dinb(n950),.dout(n951),.clk(gclk));
	jor g0651(.dina(n951),.dinb(n949),.dout(n952),.clk(gclk));
	jxor g0652(.dina(n952),.dinb(w_n605_1[2]),.dout(n953),.clk(gclk));
	jxor g0653(.dina(w_n936_0[0]),.dinb(w_n932_0[0]),.dout(n954),.clk(gclk));
	jnot g0654(.din(w_n954_0[1]),.dout(n955),.clk(gclk));
	jnot g0655(.din(w_n881_0[0]),.dout(n956),.clk(gclk));
	jnot g0656(.din(w_n771_0[0]),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n892_0[0]),.dout(n958),.clk(gclk));
	jand g0658(.dina(n958),.dinb(n957),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(n956),.dout(n960),.clk(gclk));
	jand g0660(.dina(n960),.dinb(w_n869_0[0]),.dout(n961),.clk(gclk));
	jand g0661(.dina(n961),.dinb(w_n862_0[0]),.dout(n962),.clk(gclk));
	jand g0662(.dina(n962),.dinb(n955),.dout(n963),.clk(gclk));
	jand g0663(.dina(n963),.dinb(w_n953_0[1]),.dout(n964),.clk(gclk));
	jand g0664(.dina(n964),.dinb(n947),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(n942),.dout(w_dff_A_Fwk1ch9u3_2),.clk(gclk));
	jnot g0666(.din(w_n646_0[1]),.dout(n967),.clk(gclk));
	jor g0667(.dina(w_n649_0[1]),.dinb(w_G490_0[1]),.dout(n968),.clk(gclk));
	jor g0668(.dina(w_n781_0[1]),.dinb(w_n739_1[0]),.dout(n969),.clk(gclk));
	jand g0669(.dina(n969),.dinb(w_n968_0[1]),.dout(n970),.clk(gclk));
	jxor g0670(.dina(n970),.dinb(w_dff_B_0Kif5Asu6_1),.dout(n971),.clk(gclk));
	jxor g0671(.dina(w_n783_0[2]),.dinb(w_n640_1[0]),.dout(n972),.clk(gclk));
	jxor g0672(.dina(w_n781_0[0]),.dinb(w_n650_0[0]),.dout(n973),.clk(gclk));
	jnot g0673(.din(w_n973_0[1]),.dout(n974),.clk(gclk));
	jor g0674(.dina(w_n621_0[2]),.dinb(w_n744_0[1]),.dout(n975),.clk(gclk));
	jand g0675(.dina(n975),.dinb(w_n636_0[2]),.dout(n976),.clk(gclk));
	jand g0676(.dina(w_dff_B_gMOCBXgU4_0),.dinb(w_n761_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(w_dff_B_umkbvgcF8_0),.dinb(w_n832_0[0]),.dout(n978),.clk(gclk));
	jand g0678(.dina(w_dff_B_k9iDq4bf2_0),.dinb(w_n821_0[0]),.dout(n979),.clk(gclk));
	jand g0679(.dina(w_dff_B_YzYh7TTY3_0),.dinb(w_n809_0[0]),.dout(n980),.clk(gclk));
	jand g0680(.dina(w_dff_B_dXMUhcYZ7_0),.dinb(n974),.dout(n981),.clk(gclk));
	jand g0681(.dina(n981),.dinb(w_n972_0[1]),.dout(n982),.clk(gclk));
	jand g0682(.dina(n982),.dinb(w_n971_0[1]),.dout(w_dff_A_Z53KL96c4_2),.clk(gclk));
	jnot g0683(.din(w_G1690_0[2]),.dout(n984),.clk(gclk));
	jand g0684(.dina(w_n984_0[1]),.dinb(w_G1689_0[2]),.dout(n985),.clk(gclk));
	jand g0685(.dina(w_n985_4[1]),.dinb(w_n791_0[2]),.dout(n986),.clk(gclk));
	jnot g0686(.din(w_G1689_0[1]),.dout(n987),.clk(gclk));
	jand g0687(.dina(w_n984_0[0]),.dinb(w_n987_0[1]),.dout(n988),.clk(gclk));
	jand g0688(.dina(w_n988_4[1]),.dinb(w_n795_0[2]),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_G1690_0[1]),.dinb(w_n987_0[0]),.dout(n990),.clk(gclk));
	jand g0690(.dina(w_n990_4[1]),.dinb(w_G182_0[1]),.dout(n991),.clk(gclk));
	jand g0691(.dina(w_G1690_0[0]),.dinb(w_G1689_0[0]),.dout(n992),.clk(gclk));
	jand g0692(.dina(w_n992_4[1]),.dinb(w_G185_0[1]),.dout(n993),.clk(gclk));
	jor g0693(.dina(n993),.dinb(n991),.dout(n994),.clk(gclk));
	jor g0694(.dina(w_dff_B_HzcAlp7l2_0),.dinb(n989),.dout(n995),.clk(gclk));
	jor g0695(.dina(n995),.dinb(n986),.dout(n996),.clk(gclk));
	jand g0696(.dina(n996),.dinb(w_G137_9[1]),.dout(w_dff_A_D17Lvw550_2),.clk(gclk));
	jnot g0697(.din(w_G1694_0[2]),.dout(n998),.clk(gclk));
	jand g0698(.dina(w_n998_0[1]),.dinb(w_G1691_0[2]),.dout(n999),.clk(gclk));
	jand g0699(.dina(w_n999_4[1]),.dinb(w_n791_0[1]),.dout(n1000),.clk(gclk));
	jnot g0700(.din(w_G1691_0[1]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_n998_0[0]),.dinb(w_n1001_0[1]),.dout(n1002),.clk(gclk));
	jand g0702(.dina(w_n1002_4[1]),.dinb(w_n795_0[1]),.dout(n1003),.clk(gclk));
	jand g0703(.dina(w_G1694_0[1]),.dinb(w_n1001_0[0]),.dout(n1004),.clk(gclk));
	jand g0704(.dina(w_n1004_4[1]),.dinb(w_G182_0[0]),.dout(n1005),.clk(gclk));
	jand g0705(.dina(w_G1694_0[0]),.dinb(w_G1691_0[0]),.dout(n1006),.clk(gclk));
	jand g0706(.dina(w_n1006_4[1]),.dinb(w_G185_0[0]),.dout(n1007),.clk(gclk));
	jor g0707(.dina(n1007),.dinb(n1005),.dout(n1008),.clk(gclk));
	jor g0708(.dina(w_dff_B_AMDlZ77B5_0),.dinb(n1003),.dout(n1009),.clk(gclk));
	jor g0709(.dina(n1009),.dinb(n1000),.dout(n1010),.clk(gclk));
	jand g0710(.dina(n1010),.dinb(w_G137_9[0]),.dout(w_dff_A_vv4HfquM5_2),.clk(gclk));
	jnot g0711(.din(w_G871_0),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_1[1]),.dinb(w_n793_4[0]),.dout(n1013),.clk(gclk));
	jnot g0713(.din(w_G832_0),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_1[1]),.dinb(w_n797_4[0]),.dout(n1015),.clk(gclk));
	jand g0715(.dina(w_n799_4[0]),.dinb(w_G43_0[1]),.dout(n1016),.clk(gclk));
	jand g0716(.dina(w_n801_4[0]),.dinb(w_G37_0[1]),.dout(n1017),.clk(gclk));
	jor g0717(.dina(n1017),.dinb(n1016),.dout(n1018),.clk(gclk));
	jor g0718(.dina(w_dff_B_Q3Wm8lkY8_0),.dinb(n1015),.dout(n1019),.clk(gclk));
	jor g0719(.dina(w_dff_B_3UTEDciD9_0),.dinb(n1013),.dout(w_dff_A_4Kw7kf7E8_2),.clk(gclk));
	jnot g0720(.din(w_G873_0),.dout(n1021),.clk(gclk));
	jand g0721(.dina(w_n1021_1[1]),.dinb(w_n793_3[2]),.dout(n1022),.clk(gclk));
	jnot g0722(.din(w_G834_0),.dout(n1023),.clk(gclk));
	jand g0723(.dina(w_n1023_1[1]),.dinb(w_n797_3[2]),.dout(n1024),.clk(gclk));
	jand g0724(.dina(w_n799_3[2]),.dinb(w_G76_0[1]),.dout(n1025),.clk(gclk));
	jand g0725(.dina(w_n801_3[2]),.dinb(w_G20_0[1]),.dout(n1026),.clk(gclk));
	jor g0726(.dina(n1026),.dinb(n1025),.dout(n1027),.clk(gclk));
	jor g0727(.dina(w_dff_B_0qEmyr9a0_0),.dinb(n1024),.dout(n1028),.clk(gclk));
	jor g0728(.dina(w_dff_B_O8lDN2Ov1_0),.dinb(n1022),.dout(w_dff_A_J3ukU9lO6_2),.clk(gclk));
	jnot g0729(.din(w_G875_0),.dout(n1030),.clk(gclk));
	jand g0730(.dina(w_n1030_1[1]),.dinb(w_n793_3[1]),.dout(n1031),.clk(gclk));
	jnot g0731(.din(w_G836_0),.dout(n1032),.clk(gclk));
	jand g0732(.dina(w_n1032_1[1]),.dinb(w_n797_3[1]),.dout(n1033),.clk(gclk));
	jand g0733(.dina(w_n799_3[1]),.dinb(w_G73_0[1]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(w_n801_3[1]),.dinb(w_G17_0[1]),.dout(n1035),.clk(gclk));
	jor g0735(.dina(n1035),.dinb(n1034),.dout(n1036),.clk(gclk));
	jor g0736(.dina(w_dff_B_7x1yOwOB6_0),.dinb(n1033),.dout(n1037),.clk(gclk));
	jor g0737(.dina(w_dff_B_qyYTazVA2_0),.dinb(n1031),.dout(w_dff_A_olIlU6Rz9_2),.clk(gclk));
	jnot g0738(.din(w_G877_0),.dout(n1039),.clk(gclk));
	jand g0739(.dina(w_n1039_1[1]),.dinb(w_n793_3[0]),.dout(n1040),.clk(gclk));
	jnot g0740(.din(w_G838_0),.dout(n1041),.clk(gclk));
	jand g0741(.dina(w_n797_3[0]),.dinb(w_n1041_1[1]),.dout(n1042),.clk(gclk));
	jand g0742(.dina(w_n799_3[0]),.dinb(w_G67_0[1]),.dout(n1043),.clk(gclk));
	jand g0743(.dina(w_n801_3[0]),.dinb(w_G70_0[1]),.dout(n1044),.clk(gclk));
	jor g0744(.dina(n1044),.dinb(n1043),.dout(n1045),.clk(gclk));
	jor g0745(.dina(w_dff_B_Lylrgo3b1_0),.dinb(n1042),.dout(n1046),.clk(gclk));
	jor g0746(.dina(w_dff_B_jAtPmFYd6_0),.dinb(n1040),.dout(w_dff_A_4jmLlBEL6_2),.clk(gclk));
	jand g0747(.dina(w_n1012_1[0]),.dinb(w_n840_4[0]),.dout(n1048),.clk(gclk));
	jand g0748(.dina(w_n843_4[0]),.dinb(w_n1014_1[0]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(w_n845_4[0]),.dinb(w_G43_0[0]),.dout(n1050),.clk(gclk));
	jand g0750(.dina(w_n847_4[0]),.dinb(w_G37_0[0]),.dout(n1051),.clk(gclk));
	jor g0751(.dina(n1051),.dinb(n1050),.dout(n1052),.clk(gclk));
	jor g0752(.dina(w_dff_B_1xC9NPUj3_0),.dinb(n1049),.dout(n1053),.clk(gclk));
	jor g0753(.dina(w_dff_B_WLJDP7aX5_0),.dinb(n1048),.dout(w_dff_A_AoLkuKZ61_2),.clk(gclk));
	jand g0754(.dina(w_n1021_1[0]),.dinb(w_n840_3[2]),.dout(n1055),.clk(gclk));
	jand g0755(.dina(w_n843_3[2]),.dinb(w_n1023_1[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(w_n845_3[2]),.dinb(w_G76_0[0]),.dout(n1057),.clk(gclk));
	jand g0757(.dina(w_n847_3[2]),.dinb(w_G20_0[0]),.dout(n1058),.clk(gclk));
	jor g0758(.dina(n1058),.dinb(n1057),.dout(n1059),.clk(gclk));
	jor g0759(.dina(w_dff_B_JMXQfCuI4_0),.dinb(n1056),.dout(n1060),.clk(gclk));
	jor g0760(.dina(w_dff_B_QY6h3Pf56_0),.dinb(n1055),.dout(w_dff_A_YAvYkCbM4_2),.clk(gclk));
	jand g0761(.dina(w_n1030_1[0]),.dinb(w_n840_3[1]),.dout(n1062),.clk(gclk));
	jand g0762(.dina(w_n843_3[1]),.dinb(w_n1032_1[0]),.dout(n1063),.clk(gclk));
	jand g0763(.dina(w_n845_3[1]),.dinb(w_G73_0[0]),.dout(n1064),.clk(gclk));
	jand g0764(.dina(w_n847_3[1]),.dinb(w_G17_0[0]),.dout(n1065),.clk(gclk));
	jor g0765(.dina(n1065),.dinb(n1064),.dout(n1066),.clk(gclk));
	jor g0766(.dina(w_dff_B_TCuaHdYd2_0),.dinb(n1063),.dout(n1067),.clk(gclk));
	jor g0767(.dina(w_dff_B_1oV735lj2_0),.dinb(n1062),.dout(w_dff_A_DSdWtge17_2),.clk(gclk));
	jand g0768(.dina(w_n1039_1[0]),.dinb(w_n840_3[0]),.dout(n1069),.clk(gclk));
	jand g0769(.dina(w_n843_3[0]),.dinb(w_n1041_1[0]),.dout(n1070),.clk(gclk));
	jand g0770(.dina(w_n845_3[0]),.dinb(w_G67_0[0]),.dout(n1071),.clk(gclk));
	jand g0771(.dina(w_n847_3[0]),.dinb(w_G70_0[0]),.dout(n1072),.clk(gclk));
	jor g0772(.dina(n1072),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0773(.dina(w_dff_B_CotwCRay0_0),.dinb(n1070),.dout(n1074),.clk(gclk));
	jor g0774(.dina(w_dff_B_mqzvoDyA5_0),.dinb(n1069),.dout(w_dff_A_8xMKGdES8_2),.clk(gclk));
	jand g0775(.dina(w_n985_4[0]),.dinb(w_n1012_0[2]),.dout(n1076),.clk(gclk));
	jand g0776(.dina(w_n988_4[0]),.dinb(w_n1014_0[2]),.dout(n1077),.clk(gclk));
	jand g0777(.dina(w_n990_4[0]),.dinb(w_G200_0[1]),.dout(n1078),.clk(gclk));
	jand g0778(.dina(w_n992_4[0]),.dinb(w_G170_0[1]),.dout(n1079),.clk(gclk));
	jor g0779(.dina(n1079),.dinb(n1078),.dout(n1080),.clk(gclk));
	jor g0780(.dina(w_dff_B_3ID8azaP2_0),.dinb(n1077),.dout(n1081),.clk(gclk));
	jor g0781(.dina(w_dff_B_5PjVobUQ4_0),.dinb(n1076),.dout(n1082),.clk(gclk));
	jand g0782(.dina(n1082),.dinb(w_G137_8[2]),.dout(w_dff_A_vpF12bp06_2),.clk(gclk));
	jand g0783(.dina(w_n985_3[2]),.dinb(w_n1039_0[2]),.dout(n1084),.clk(gclk));
	jand g0784(.dina(w_n988_3[2]),.dinb(w_n1041_0[2]),.dout(n1085),.clk(gclk));
	jand g0785(.dina(w_n990_3[2]),.dinb(w_G188_0[1]),.dout(n1086),.clk(gclk));
	jand g0786(.dina(w_n992_3[2]),.dinb(w_G158_0[1]),.dout(n1087),.clk(gclk));
	jor g0787(.dina(n1087),.dinb(n1086),.dout(n1088),.clk(gclk));
	jor g0788(.dina(w_dff_B_mVA8vvvh4_0),.dinb(n1085),.dout(n1089),.clk(gclk));
	jor g0789(.dina(w_dff_B_AjhPezaV8_0),.dinb(n1084),.dout(n1090),.clk(gclk));
	jand g0790(.dina(n1090),.dinb(w_G137_8[1]),.dout(w_dff_A_f74DpKmn1_2),.clk(gclk));
	jand g0791(.dina(w_n985_3[1]),.dinb(w_n1030_0[2]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(w_n988_3[1]),.dinb(w_n1032_0[2]),.dout(n1093),.clk(gclk));
	jand g0793(.dina(w_n990_3[1]),.dinb(w_G155_0[1]),.dout(n1094),.clk(gclk));
	jand g0794(.dina(w_n992_3[1]),.dinb(w_G152_0[1]),.dout(n1095),.clk(gclk));
	jor g0795(.dina(n1095),.dinb(n1094),.dout(n1096),.clk(gclk));
	jor g0796(.dina(w_dff_B_Wb3Mxokv3_0),.dinb(n1093),.dout(n1097),.clk(gclk));
	jor g0797(.dina(w_dff_B_dZoSkuxT9_0),.dinb(n1092),.dout(n1098),.clk(gclk));
	jand g0798(.dina(n1098),.dinb(w_G137_8[0]),.dout(w_dff_A_E82YkNP98_2),.clk(gclk));
	jand g0799(.dina(w_n985_3[0]),.dinb(w_n1021_0[2]),.dout(n1100),.clk(gclk));
	jand g0800(.dina(w_n988_3[0]),.dinb(w_n1023_0[2]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(w_n990_3[0]),.dinb(w_G149_0[1]),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n992_3[0]),.dinb(w_G146_0[1]),.dout(n1103),.clk(gclk));
	jor g0803(.dina(n1103),.dinb(n1102),.dout(n1104),.clk(gclk));
	jor g0804(.dina(w_dff_B_3mQ230dl9_0),.dinb(n1101),.dout(n1105),.clk(gclk));
	jor g0805(.dina(w_dff_B_8LNnabtE7_0),.dinb(n1100),.dout(n1106),.clk(gclk));
	jand g0806(.dina(n1106),.dinb(w_G137_7[2]),.dout(w_dff_A_IXXnVHd24_2),.clk(gclk));
	jand g0807(.dina(w_n999_4[0]),.dinb(w_n1012_0[1]),.dout(n1108),.clk(gclk));
	jand g0808(.dina(w_n1002_4[0]),.dinb(w_n1014_0[1]),.dout(n1109),.clk(gclk));
	jand g0809(.dina(w_n1004_4[0]),.dinb(w_G200_0[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(w_n1006_4[0]),.dinb(w_G170_0[0]),.dout(n1111),.clk(gclk));
	jor g0811(.dina(n1111),.dinb(n1110),.dout(n1112),.clk(gclk));
	jor g0812(.dina(w_dff_B_YhCP3RJR5_0),.dinb(n1109),.dout(n1113),.clk(gclk));
	jor g0813(.dina(w_dff_B_wJYACATe1_0),.dinb(n1108),.dout(n1114),.clk(gclk));
	jand g0814(.dina(n1114),.dinb(w_G137_7[1]),.dout(w_dff_A_D1HnF7sc8_2),.clk(gclk));
	jand g0815(.dina(w_n999_3[2]),.dinb(w_n1039_0[1]),.dout(n1116),.clk(gclk));
	jand g0816(.dina(w_n1002_3[2]),.dinb(w_n1041_0[1]),.dout(n1117),.clk(gclk));
	jand g0817(.dina(w_n1004_3[2]),.dinb(w_G188_0[0]),.dout(n1118),.clk(gclk));
	jand g0818(.dina(w_n1006_3[2]),.dinb(w_G158_0[0]),.dout(n1119),.clk(gclk));
	jor g0819(.dina(n1119),.dinb(n1118),.dout(n1120),.clk(gclk));
	jor g0820(.dina(w_dff_B_HqQAKbo35_0),.dinb(n1117),.dout(n1121),.clk(gclk));
	jor g0821(.dina(w_dff_B_NqLTbuqA7_0),.dinb(n1116),.dout(n1122),.clk(gclk));
	jand g0822(.dina(n1122),.dinb(w_G137_7[0]),.dout(w_dff_A_DeuY0TwH2_2),.clk(gclk));
	jand g0823(.dina(w_n999_3[1]),.dinb(w_n1030_0[1]),.dout(n1124),.clk(gclk));
	jand g0824(.dina(w_n1002_3[1]),.dinb(w_n1032_0[1]),.dout(n1125),.clk(gclk));
	jand g0825(.dina(w_n1004_3[1]),.dinb(w_G155_0[0]),.dout(n1126),.clk(gclk));
	jand g0826(.dina(w_n1006_3[1]),.dinb(w_G152_0[0]),.dout(n1127),.clk(gclk));
	jor g0827(.dina(n1127),.dinb(n1126),.dout(n1128),.clk(gclk));
	jor g0828(.dina(w_dff_B_xyY6mh8V6_0),.dinb(n1125),.dout(n1129),.clk(gclk));
	jor g0829(.dina(w_dff_B_iRjXtJ673_0),.dinb(n1124),.dout(n1130),.clk(gclk));
	jand g0830(.dina(n1130),.dinb(w_G137_6[2]),.dout(w_dff_A_tZp0S1964_2),.clk(gclk));
	jand g0831(.dina(w_n999_3[0]),.dinb(w_n1021_0[1]),.dout(n1132),.clk(gclk));
	jand g0832(.dina(w_n1002_3[0]),.dinb(w_n1023_0[1]),.dout(n1133),.clk(gclk));
	jand g0833(.dina(w_n1004_3[0]),.dinb(w_G149_0[0]),.dout(n1134),.clk(gclk));
	jand g0834(.dina(w_n1006_3[0]),.dinb(w_G146_0[0]),.dout(n1135),.clk(gclk));
	jor g0835(.dina(n1135),.dinb(n1134),.dout(n1136),.clk(gclk));
	jor g0836(.dina(w_dff_B_HC3u8Yfs7_0),.dinb(n1133),.dout(n1137),.clk(gclk));
	jor g0837(.dina(w_dff_B_u7wzn8vO0_0),.dinb(n1132),.dout(n1138),.clk(gclk));
	jand g0838(.dina(n1138),.dinb(w_G137_6[1]),.dout(w_dff_A_zqQOhykr8_2),.clk(gclk));
	jand g0839(.dina(w_n789_0[1]),.dinb(w_G3724_0[2]),.dout(n1140),.clk(gclk));
	jnot g0840(.din(w_G3717_0[1]),.dout(n1141),.clk(gclk));
	jnot g0841(.din(w_G3724_0[1]),.dout(n1142),.clk(gclk));
	jand g0842(.dina(w_n1142_0[1]),.dinb(w_G123_0[1]),.dout(n1143),.clk(gclk));
	jor g0843(.dina(n1143),.dinb(n1141),.dout(n1144),.clk(gclk));
	jor g0844(.dina(w_dff_B_mGPgZ6e00_0),.dinb(n1140),.dout(n1145),.clk(gclk));
	jnot g0845(.din(G135),.dout(n1146),.clk(gclk));
	jnot g0846(.din(G4115),.dout(n1147),.clk(gclk));
	jor g0847(.dina(n1147),.dinb(n1146),.dout(n1148),.clk(gclk));
	jxor g0848(.dina(w_n636_0[1]),.dinb(w_G132_0[1]),.dout(n1149),.clk(gclk));
	jand g0849(.dina(n1149),.dinb(w_G3724_0[0]),.dout(n1150),.clk(gclk));
	jnot g0850(.din(w_n401_0[1]),.dout(n1151),.clk(gclk));
	jand g0851(.dina(w_n1151_0[1]),.dinb(w_n1142_0[0]),.dout(n1152),.clk(gclk));
	jor g0852(.dina(n1152),.dinb(w_G3717_0[0]),.dout(n1153),.clk(gclk));
	jor g0853(.dina(n1153),.dinb(w_dff_B_6brFvEQp9_1),.dout(n1154),.clk(gclk));
	jand g0854(.dina(n1154),.dinb(w_dff_B_pBkP35yK1_1),.dout(n1155),.clk(gclk));
	jand g0855(.dina(w_dff_B_JCS4xw4h9_0),.dinb(n1145),.dout(w_dff_A_YI0eKhC97_2),.clk(gclk));
	jor g0856(.dina(w_n783_0[1]),.dinb(w_n640_0[2]),.dout(n1157),.clk(gclk));
	jxor g0857(.dina(n1157),.dinb(w_G132_0[0]),.dout(w_dff_A_Yu4al2p14_2),.clk(gclk));
	jand g0858(.dina(w_n789_0[0]),.dinb(w_n747_2[1]),.dout(n1159),.clk(gclk));
	jand g0859(.dina(w_n753_5[0]),.dinb(w_G123_0[0]),.dout(n1160),.clk(gclk));
	jand g0860(.dina(w_n751_1[1]),.dinb(w_n1151_0[0]),.dout(n1161),.clk(gclk));
	jor g0861(.dina(n1161),.dinb(n1160),.dout(n1162),.clk(gclk));
	jor g0862(.dina(w_dff_B_E5a09JiM7_0),.dinb(n1159),.dout(n1163),.clk(gclk));
	jnot g0863(.din(w_n1163_1[2]),.dout(w_dff_A_F0NuwJLN0_1),.clk(gclk));
	jor g0864(.dina(w_n972_0[0]),.dinb(w_n748_2[0]),.dout(n1165),.clk(gclk));
	jand g0865(.dina(w_n751_1[0]),.dinb(w_n407_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n753_4[2]),.dinb(G121),.dout(n1167),.clk(gclk));
	jor g0867(.dina(n1167),.dinb(n1166),.dout(n1168),.clk(gclk));
	jnot g0868(.din(n1168),.dout(n1169),.clk(gclk));
	jand g0869(.dina(w_dff_B_7Ql7B85O2_0),.dinb(n1165),.dout(G826_fa_),.clk(gclk));
	jor g0870(.dina(w_n971_0[0]),.dinb(w_n748_1[2]),.dout(n1171),.clk(gclk));
	jor g0871(.dina(w_n765_3[0]),.dinb(w_n372_0[1]),.dout(n1172),.clk(gclk));
	jand g0872(.dina(w_n753_4[1]),.dinb(G116),.dout(n1173),.clk(gclk));
	jnot g0873(.din(n1173),.dout(n1174),.clk(gclk));
	jand g0874(.dina(n1174),.dinb(n1172),.dout(n1175),.clk(gclk));
	jand g0875(.dina(w_dff_B_h7shaPp49_0),.dinb(n1171),.dout(G828_fa_),.clk(gclk));
	jand g0876(.dina(w_n973_0[0]),.dinb(w_n747_2[0]),.dout(n1177),.clk(gclk));
	jnot g0877(.din(n1177),.dout(n1178),.clk(gclk));
	jor g0878(.dina(w_n765_2[2]),.dinb(w_n383_0[1]),.dout(n1179),.clk(gclk));
	jand g0879(.dina(w_n753_4[0]),.dinb(G112),.dout(n1180),.clk(gclk));
	jnot g0880(.din(n1180),.dout(n1181),.clk(gclk));
	jand g0881(.dina(n1181),.dinb(n1179),.dout(n1182),.clk(gclk));
	jand g0882(.dina(w_dff_B_8UP3HyQ55_0),.dinb(n1178),.dout(G830_fa_),.clk(gclk));
	jnot g0883(.din(w_G1000_0),.dout(n1184),.clk(gclk));
	jand g0884(.dina(w_G559_0[0]),.dinb(w_G245_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(n1185),.dinb(w_n318_0[0]),.dout(n1186),.clk(gclk));
	jand g0886(.dina(n1186),.dinb(w_G601_0),.dout(n1187),.clk(gclk));
	jand g0887(.dina(w_dff_B_KhItkqzk3_0),.dinb(w_n661_0[0]),.dout(n1188),.clk(gclk));
	jand g0888(.dina(n1188),.dinb(w_n671_0[0]),.dout(n1189),.clk(gclk));
	jand g0889(.dina(w_dff_B_nZg96tG07_0),.dinb(w_n914_0[0]),.dout(n1190),.clk(gclk));
	jand g0890(.dina(n1190),.dinb(w_dff_B_eyaGwMpD4_1),.dout(w_dff_A_YmBmEb0r2_2),.clk(gclk));
	jand g0891(.dina(w_n941_0[0]),.dinb(w_n747_1[2]),.dout(n1192),.clk(gclk));
	jnot g0892(.din(w_n528_0[1]),.dout(n1193),.clk(gclk));
	jand g0893(.dina(w_n751_0[2]),.dinb(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_n753_3[2]),.dinb(G115),.dout(n1195),.clk(gclk));
	jor g0895(.dina(n1195),.dinb(n1194),.dout(n1196),.clk(gclk));
	jor g0896(.dina(n1196),.dinb(n1192),.dout(n1197),.clk(gclk));
	jnot g0897(.din(w_n1197_1[2]),.dout(w_dff_A_61pVhAxr4_1),.clk(gclk));
	jand g0898(.dina(w_n946_0[0]),.dinb(w_n747_1[1]),.dout(n1199),.clk(gclk));
	jor g0899(.dina(w_n765_2[1]),.dinb(w_n551_0[0]),.dout(n1200),.clk(gclk));
	jand g0900(.dina(w_n753_3[1]),.dinb(G114),.dout(n1201),.clk(gclk));
	jnot g0901(.din(n1201),.dout(n1202),.clk(gclk));
	jand g0902(.dina(n1202),.dinb(n1200),.dout(n1203),.clk(gclk));
	jnot g0903(.din(n1203),.dout(n1204),.clk(gclk));
	jor g0904(.dina(n1204),.dinb(n1199),.dout(n1205),.clk(gclk));
	jnot g0905(.din(w_n1205_1[2]),.dout(w_dff_A_TCYtEEkG3_1),.clk(gclk));
	jor g0906(.dina(w_n953_0[0]),.dinb(w_n748_1[1]),.dout(n1207),.clk(gclk));
	jor g0907(.dina(w_n765_2[0]),.dinb(w_n517_0[0]),.dout(n1208),.clk(gclk));
	jand g0908(.dina(w_n753_3[0]),.dinb(G53),.dout(n1209),.clk(gclk));
	jnot g0909(.din(n1209),.dout(n1210),.clk(gclk));
	jand g0910(.dina(n1210),.dinb(n1208),.dout(n1211),.clk(gclk));
	jand g0911(.dina(n1211),.dinb(n1207),.dout(G867_fa_),.clk(gclk));
	jand g0912(.dina(w_n954_0[0]),.dinb(w_n747_1[0]),.dout(n1213),.clk(gclk));
	jnot g0913(.din(n1213),.dout(n1214),.clk(gclk));
	jor g0914(.dina(w_n765_1[2]),.dinb(w_n540_0[0]),.dout(n1215),.clk(gclk));
	jand g0915(.dina(w_n753_2[2]),.dinb(G113),.dout(n1216),.clk(gclk));
	jnot g0916(.din(n1216),.dout(n1217),.clk(gclk));
	jand g0917(.dina(n1217),.dinb(n1215),.dout(n1218),.clk(gclk));
	jand g0918(.dina(n1218),.dinb(n1214),.dout(G869_fa_),.clk(gclk));
	jand g0919(.dina(w_n1197_1[1]),.dinb(w_n840_2[2]),.dout(n1220),.clk(gclk));
	jand g0920(.dina(w_n1163_1[1]),.dinb(w_n843_2[2]),.dout(n1221),.clk(gclk));
	jand g0921(.dina(w_n845_2[2]),.dinb(w_G109_0[1]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(w_n847_2[2]),.dinb(w_G106_0[1]),.dout(n1223),.clk(gclk));
	jor g0923(.dina(n1223),.dinb(n1222),.dout(n1224),.clk(gclk));
	jor g0924(.dina(w_dff_B_ENRx4VdZ0_0),.dinb(n1221),.dout(n1225),.clk(gclk));
	jor g0925(.dina(n1225),.dinb(n1220),.dout(w_dff_A_NjJ1rGZa7_2),.clk(gclk));
	jand g0926(.dina(w_n1197_1[0]),.dinb(w_n793_2[2]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_n1163_1[0]),.dinb(w_n797_2[2]),.dout(n1228),.clk(gclk));
	jand g0928(.dina(w_n799_2[2]),.dinb(w_G109_0[0]),.dout(n1229),.clk(gclk));
	jand g0929(.dina(w_n801_2[2]),.dinb(w_G106_0[0]),.dout(n1230),.clk(gclk));
	jor g0930(.dina(n1230),.dinb(n1229),.dout(n1231),.clk(gclk));
	jor g0931(.dina(w_dff_B_b4hchHMT6_0),.dinb(n1228),.dout(n1232),.clk(gclk));
	jor g0932(.dina(n1232),.dinb(n1227),.dout(w_dff_A_AebEAUfu6_2),.clk(gclk));
	jand g0933(.dina(w_n1205_1[1]),.dinb(w_n793_2[1]),.dout(n1234),.clk(gclk));
	jnot g0934(.din(w_G826_0),.dout(n1235),.clk(gclk));
	jand g0935(.dina(w_n1235_1[1]),.dinb(w_n797_2[1]),.dout(n1236),.clk(gclk));
	jand g0936(.dina(w_n799_2[1]),.dinb(w_G46_0[1]),.dout(n1237),.clk(gclk));
	jand g0937(.dina(w_n801_2[1]),.dinb(w_G49_0[1]),.dout(n1238),.clk(gclk));
	jor g0938(.dina(n1238),.dinb(n1237),.dout(n1239),.clk(gclk));
	jor g0939(.dina(w_dff_B_QDtKQf1m5_0),.dinb(n1236),.dout(n1240),.clk(gclk));
	jor g0940(.dina(n1240),.dinb(n1234),.dout(w_dff_A_tP90ihO79_2),.clk(gclk));
	jnot g0941(.din(w_G867_0),.dout(n1242),.clk(gclk));
	jand g0942(.dina(w_n1242_1[1]),.dinb(w_n793_2[0]),.dout(n1243),.clk(gclk));
	jnot g0943(.din(w_G828_0),.dout(n1244),.clk(gclk));
	jand g0944(.dina(w_n1244_1[1]),.dinb(w_n797_2[0]),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n799_2[0]),.dinb(w_G100_0[1]),.dout(n1246),.clk(gclk));
	jand g0946(.dina(w_n801_2[0]),.dinb(w_G103_0[1]),.dout(n1247),.clk(gclk));
	jor g0947(.dina(n1247),.dinb(n1246),.dout(n1248),.clk(gclk));
	jor g0948(.dina(w_dff_B_AEJFMYQM6_0),.dinb(n1245),.dout(n1249),.clk(gclk));
	jor g0949(.dina(n1249),.dinb(n1243),.dout(w_dff_A_4CRHhEj26_2),.clk(gclk));
	jnot g0950(.din(w_G869_0),.dout(n1251),.clk(gclk));
	jand g0951(.dina(w_n1251_1[1]),.dinb(w_n793_1[2]),.dout(n1252),.clk(gclk));
	jnot g0952(.din(w_G830_0),.dout(n1253),.clk(gclk));
	jand g0953(.dina(w_n1253_1[1]),.dinb(w_n797_1[2]),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n799_1[2]),.dinb(w_G91_0[1]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n801_1[2]),.dinb(w_G40_0[1]),.dout(n1256),.clk(gclk));
	jor g0956(.dina(n1256),.dinb(n1255),.dout(n1257),.clk(gclk));
	jor g0957(.dina(w_dff_B_KgDYaSie1_0),.dinb(n1254),.dout(n1258),.clk(gclk));
	jor g0958(.dina(n1258),.dinb(n1252),.dout(w_dff_A_7Y0fh7EU0_2),.clk(gclk));
	jand g0959(.dina(w_n1205_1[0]),.dinb(w_n840_2[1]),.dout(n1260),.clk(gclk));
	jand g0960(.dina(w_n1235_1[0]),.dinb(w_n843_2[1]),.dout(n1261),.clk(gclk));
	jand g0961(.dina(w_n845_2[1]),.dinb(w_G46_0[0]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(w_n847_2[1]),.dinb(w_G49_0[0]),.dout(n1263),.clk(gclk));
	jor g0963(.dina(n1263),.dinb(n1262),.dout(n1264),.clk(gclk));
	jor g0964(.dina(w_dff_B_q4CWaEu15_0),.dinb(n1261),.dout(n1265),.clk(gclk));
	jor g0965(.dina(n1265),.dinb(n1260),.dout(w_dff_A_rFepXOn66_2),.clk(gclk));
	jand g0966(.dina(w_n1242_1[0]),.dinb(w_n840_2[0]),.dout(n1267),.clk(gclk));
	jand g0967(.dina(w_n1244_1[0]),.dinb(w_n843_2[0]),.dout(n1268),.clk(gclk));
	jand g0968(.dina(w_n845_2[0]),.dinb(w_G100_0[0]),.dout(n1269),.clk(gclk));
	jand g0969(.dina(w_n847_2[0]),.dinb(w_G103_0[0]),.dout(n1270),.clk(gclk));
	jor g0970(.dina(n1270),.dinb(n1269),.dout(n1271),.clk(gclk));
	jor g0971(.dina(w_dff_B_E8rqHHnu5_0),.dinb(n1268),.dout(n1272),.clk(gclk));
	jor g0972(.dina(n1272),.dinb(n1267),.dout(w_dff_A_WBcazqRS7_2),.clk(gclk));
	jand g0973(.dina(w_n1251_1[0]),.dinb(w_n840_1[2]),.dout(n1274),.clk(gclk));
	jand g0974(.dina(w_n1253_1[0]),.dinb(w_n843_1[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(w_n845_1[2]),.dinb(w_G91_0[0]),.dout(n1276),.clk(gclk));
	jand g0976(.dina(w_n847_1[2]),.dinb(w_G40_0[0]),.dout(n1277),.clk(gclk));
	jor g0977(.dina(n1277),.dinb(n1276),.dout(n1278),.clk(gclk));
	jor g0978(.dina(w_dff_B_Qel3kc1U0_0),.dinb(n1275),.dout(n1279),.clk(gclk));
	jor g0979(.dina(n1279),.dinb(n1274),.dout(w_dff_A_d2B7YkhN0_2),.clk(gclk));
	jand g0980(.dina(w_n1251_0[2]),.dinb(w_n985_2[2]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(w_n1253_0[2]),.dinb(w_n988_2[2]),.dout(n1282),.clk(gclk));
	jand g0982(.dina(w_n990_2[2]),.dinb(w_G203_0[1]),.dout(n1283),.clk(gclk));
	jand g0983(.dina(w_n992_2[2]),.dinb(w_G173_0[1]),.dout(n1284),.clk(gclk));
	jor g0984(.dina(n1284),.dinb(n1283),.dout(n1285),.clk(gclk));
	jor g0985(.dina(w_dff_B_ivEV8khi6_0),.dinb(n1282),.dout(n1286),.clk(gclk));
	jor g0986(.dina(n1286),.dinb(n1281),.dout(n1287),.clk(gclk));
	jand g0987(.dina(n1287),.dinb(w_G137_6[0]),.dout(w_dff_A_7YR1FAlA0_2),.clk(gclk));
	jand g0988(.dina(w_n1242_0[2]),.dinb(w_n985_2[1]),.dout(n1289),.clk(gclk));
	jand g0989(.dina(w_n1244_0[2]),.dinb(w_n988_2[1]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(w_n990_2[1]),.dinb(w_G197_0[1]),.dout(n1291),.clk(gclk));
	jand g0991(.dina(w_n992_2[1]),.dinb(w_G167_0[1]),.dout(n1292),.clk(gclk));
	jor g0992(.dina(n1292),.dinb(n1291),.dout(n1293),.clk(gclk));
	jor g0993(.dina(w_dff_B_7cxBKTql8_0),.dinb(n1290),.dout(n1294),.clk(gclk));
	jor g0994(.dina(n1294),.dinb(n1289),.dout(n1295),.clk(gclk));
	jand g0995(.dina(n1295),.dinb(w_G137_5[2]),.dout(w_dff_A_2lBg0wOi0_2),.clk(gclk));
	jand g0996(.dina(w_n1205_0[2]),.dinb(w_n985_2[0]),.dout(n1297),.clk(gclk));
	jand g0997(.dina(w_n1235_0[2]),.dinb(w_n988_2[0]),.dout(n1298),.clk(gclk));
	jand g0998(.dina(w_n990_2[0]),.dinb(w_G194_0[1]),.dout(n1299),.clk(gclk));
	jand g0999(.dina(w_n992_2[0]),.dinb(w_G164_0[1]),.dout(n1300),.clk(gclk));
	jor g1000(.dina(n1300),.dinb(n1299),.dout(n1301),.clk(gclk));
	jor g1001(.dina(w_dff_B_yNQ5VDmC3_0),.dinb(n1298),.dout(n1302),.clk(gclk));
	jor g1002(.dina(n1302),.dinb(n1297),.dout(n1303),.clk(gclk));
	jand g1003(.dina(n1303),.dinb(w_G137_5[1]),.dout(w_dff_A_hz6kOtRe3_2),.clk(gclk));
	jand g1004(.dina(w_n1197_0[2]),.dinb(w_n985_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(w_n1163_0[2]),.dinb(w_n988_1[2]),.dout(n1306),.clk(gclk));
	jand g1006(.dina(w_n990_1[2]),.dinb(w_G191_0[1]),.dout(n1307),.clk(gclk));
	jand g1007(.dina(w_n992_1[2]),.dinb(w_G161_0[1]),.dout(n1308),.clk(gclk));
	jor g1008(.dina(n1308),.dinb(n1307),.dout(n1309),.clk(gclk));
	jor g1009(.dina(w_dff_B_2MPKNbl66_0),.dinb(n1306),.dout(n1310),.clk(gclk));
	jor g1010(.dina(n1310),.dinb(n1305),.dout(n1311),.clk(gclk));
	jand g1011(.dina(n1311),.dinb(w_G137_5[0]),.dout(w_dff_A_RrQzvuqd9_2),.clk(gclk));
	jand g1012(.dina(w_n1251_0[1]),.dinb(w_n999_2[2]),.dout(n1313),.clk(gclk));
	jand g1013(.dina(w_n1253_0[1]),.dinb(w_n1002_2[2]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(w_n1004_2[2]),.dinb(w_G203_0[0]),.dout(n1315),.clk(gclk));
	jand g1015(.dina(w_n1006_2[2]),.dinb(w_G173_0[0]),.dout(n1316),.clk(gclk));
	jor g1016(.dina(n1316),.dinb(n1315),.dout(n1317),.clk(gclk));
	jor g1017(.dina(w_dff_B_Mup6Tlwp7_0),.dinb(n1314),.dout(n1318),.clk(gclk));
	jor g1018(.dina(n1318),.dinb(n1313),.dout(n1319),.clk(gclk));
	jand g1019(.dina(n1319),.dinb(w_G137_4[2]),.dout(w_dff_A_0wj4FSAV3_2),.clk(gclk));
	jand g1020(.dina(w_n1242_0[1]),.dinb(w_n999_2[1]),.dout(n1321),.clk(gclk));
	jand g1021(.dina(w_n1244_0[1]),.dinb(w_n1002_2[1]),.dout(n1322),.clk(gclk));
	jand g1022(.dina(w_n1004_2[1]),.dinb(w_G197_0[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(w_n1006_2[1]),.dinb(w_G167_0[0]),.dout(n1324),.clk(gclk));
	jor g1024(.dina(n1324),.dinb(n1323),.dout(n1325),.clk(gclk));
	jor g1025(.dina(w_dff_B_fyySlzZz8_0),.dinb(n1322),.dout(n1326),.clk(gclk));
	jor g1026(.dina(n1326),.dinb(n1321),.dout(n1327),.clk(gclk));
	jand g1027(.dina(n1327),.dinb(w_G137_4[1]),.dout(w_dff_A_YzzF2G7s5_2),.clk(gclk));
	jand g1028(.dina(w_n1205_0[1]),.dinb(w_n999_2[0]),.dout(n1329),.clk(gclk));
	jand g1029(.dina(w_n1235_0[1]),.dinb(w_n1002_2[0]),.dout(n1330),.clk(gclk));
	jand g1030(.dina(w_n1004_2[0]),.dinb(w_G194_0[0]),.dout(n1331),.clk(gclk));
	jand g1031(.dina(w_n1006_2[0]),.dinb(w_G164_0[0]),.dout(n1332),.clk(gclk));
	jor g1032(.dina(n1332),.dinb(n1331),.dout(n1333),.clk(gclk));
	jor g1033(.dina(w_dff_B_7nkid9JF1_0),.dinb(n1330),.dout(n1334),.clk(gclk));
	jor g1034(.dina(n1334),.dinb(n1329),.dout(n1335),.clk(gclk));
	jand g1035(.dina(n1335),.dinb(w_G137_4[0]),.dout(w_dff_A_o0JBYaTp4_2),.clk(gclk));
	jand g1036(.dina(w_n1197_0[1]),.dinb(w_n999_1[2]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(w_n1163_0[1]),.dinb(w_n1002_1[2]),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n1004_1[2]),.dinb(w_G191_0[0]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n1006_1[2]),.dinb(w_G161_0[0]),.dout(n1340),.clk(gclk));
	jor g1040(.dina(n1340),.dinb(n1339),.dout(n1341),.clk(gclk));
	jor g1041(.dina(w_dff_B_Ll5YcClR3_0),.dinb(n1338),.dout(n1342),.clk(gclk));
	jor g1042(.dina(n1342),.dinb(n1337),.dout(n1343),.clk(gclk));
	jand g1043(.dina(n1343),.dinb(w_G137_3[2]),.dout(w_dff_A_S3yRiD3O3_2),.clk(gclk));
	jor g1044(.dina(w_G4091_2[0]),.dinb(G120),.dout(n1345),.clk(gclk));
	jand g1045(.dina(w_n435_0[2]),.dinb(w_G251_3[1]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1347),.clk(gclk));
	jor g1047(.dina(n1347),.dinb(w_n437_0[1]),.dout(n1348),.clk(gclk));
	jor g1048(.dina(n1348),.dinb(n1346),.dout(n1349),.clk(gclk));
	jand g1049(.dina(w_n435_0[1]),.dinb(w_n366_3[1]),.dout(n1350),.clk(gclk));
	jand g1050(.dina(w_G341_0[2]),.dinb(w_n368_4[0]),.dout(n1351),.clk(gclk));
	jor g1051(.dina(n1351),.dinb(w_G523_0[2]),.dout(n1352),.clk(gclk));
	jor g1052(.dina(n1352),.dinb(n1350),.dout(n1353),.clk(gclk));
	jand g1053(.dina(n1353),.dinb(n1349),.dout(n1354),.clk(gclk));
	jxor g1054(.dina(w_n408_0[0]),.dinb(w_n401_0[0]),.dout(n1355),.clk(gclk));
	jxor g1055(.dina(w_n383_0[0]),.dinb(w_n372_0[0]),.dout(n1356),.clk(gclk));
	jxor g1056(.dina(n1356),.dinb(n1355),.dout(n1357),.clk(gclk));
	jxor g1057(.dina(n1357),.dinb(n1354),.dout(n1358),.clk(gclk));
	jnot g1058(.din(w_n1358_0[1]),.dout(n1359),.clk(gclk));
	jor g1059(.dina(w_n410_0[1]),.dinb(w_G248_3[2]),.dout(n1360),.clk(gclk));
	jor g1060(.dina(w_G514_0[1]),.dinb(w_n368_3[2]),.dout(n1361),.clk(gclk));
	jand g1061(.dina(n1361),.dinb(n1360),.dout(n1362),.clk(gclk));
	jxor g1062(.dina(n1362),.dinb(w_n419_0[0]),.dout(n1363),.clk(gclk));
	jor g1063(.dina(w_G351_1[0]),.dinb(w_n402_1[2]),.dout(n1364),.clk(gclk));
	jor g1064(.dina(w_n385_0[2]),.dinb(w_n405_1[2]),.dout(n1365),.clk(gclk));
	jand g1065(.dina(n1365),.dinb(w_G534_0[1]),.dout(n1366),.clk(gclk));
	jand g1066(.dina(n1366),.dinb(n1364),.dout(n1367),.clk(gclk));
	jor g1067(.dina(w_G351_0[2]),.dinb(w_G254_1[1]),.dout(n1368),.clk(gclk));
	jor g1068(.dina(w_n385_0[1]),.dinb(w_G242_1[1]),.dout(n1369),.clk(gclk));
	jand g1069(.dina(n1369),.dinb(w_n388_0[1]),.dout(n1370),.clk(gclk));
	jand g1070(.dina(n1370),.dinb(n1368),.dout(n1371),.clk(gclk));
	jor g1071(.dina(n1371),.dinb(n1367),.dout(n1372),.clk(gclk));
	jand g1072(.dina(w_n424_1[0]),.dinb(w_G251_3[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(w_G324_0[2]),.dinb(w_G248_3[1]),.dout(n1374),.clk(gclk));
	jor g1074(.dina(n1374),.dinb(w_n426_0[0]),.dout(n1375),.clk(gclk));
	jor g1075(.dina(n1375),.dinb(n1373),.dout(n1376),.clk(gclk));
	jand g1076(.dina(w_n424_0[2]),.dinb(w_n366_3[0]),.dout(n1377),.clk(gclk));
	jand g1077(.dina(w_G324_0[1]),.dinb(w_n368_3[1]),.dout(n1378),.clk(gclk));
	jor g1078(.dina(n1378),.dinb(w_G503_0[1]),.dout(n1379),.clk(gclk));
	jor g1079(.dina(n1379),.dinb(n1377),.dout(n1380),.clk(gclk));
	jand g1080(.dina(n1380),.dinb(n1376),.dout(n1381),.clk(gclk));
	jxor g1081(.dina(n1381),.dinb(n1372),.dout(n1382),.clk(gclk));
	jxor g1082(.dina(n1382),.dinb(n1363),.dout(n1383),.clk(gclk));
	jnot g1083(.din(w_n1383_0[1]),.dout(n1384),.clk(gclk));
	jand g1084(.dina(w_n1383_0[0]),.dinb(n1359),.dout(n1385),.clk(gclk));
	jor g1085(.dina(n1385),.dinb(w_G4091_1[2]),.dout(n1386),.clk(gclk));
	jor g1086(.dina(n1345),.dinb(w_n746_1[0]),.dout(n1388),.clk(gclk));
	jand g1087(.dina(n1384),.dinb(w_n1358_0[0]),.dout(n1389),.clk(gclk));
	jor g1088(.dina(n1386),.dinb(n1389),.dout(n1390),.clk(gclk));
	jand g1089(.dina(n1390),.dinb(w_n746_0[2]),.dout(n1391),.clk(gclk));
	jnot g1090(.din(w_n1391_0[1]),.dout(n1392),.clk(gclk));
	jand g1091(.dina(w_n633_0[2]),.dinb(w_G2174_0[2]),.dout(n1393),.clk(gclk));
	jor g1092(.dina(w_dff_B_Gpxjw03t9_0),.dinb(w_n732_0[0]),.dout(n1394),.clk(gclk));
	jand g1093(.dina(w_n736_0[0]),.dinb(w_n640_0[1]),.dout(n1395),.clk(gclk));
	jor g1094(.dina(w_n740_0[0]),.dinb(w_n641_0[0]),.dout(n1396),.clk(gclk));
	jand g1095(.dina(n1396),.dinb(w_n646_0[0]),.dout(n1397),.clk(gclk));
	jor g1096(.dina(n1397),.dinb(n1395),.dout(n1398),.clk(gclk));
	jnot g1097(.din(w_n1398_0[1]),.dout(n1399),.clk(gclk));
	jand g1098(.dina(w_n1399_0[1]),.dinb(w_n739_0[2]),.dout(n1400),.clk(gclk));
	jnot g1099(.din(w_n739_0[1]),.dout(n1401),.clk(gclk));
	jand g1100(.dina(w_n1398_0[0]),.dinb(n1401),.dout(n1402),.clk(gclk));
	jor g1101(.dina(n1402),.dinb(w_n651_0[1]),.dout(n1403),.clk(gclk));
	jor g1102(.dina(n1403),.dinb(n1400),.dout(n1404),.clk(gclk));
	jand g1103(.dina(w_dff_B_jwnaOYvi6_0),.dinb(w_n1394_0[1]),.dout(n1405),.clk(gclk));
	jnot g1104(.din(w_n1394_0[0]),.dout(n1406),.clk(gclk));
	jxor g1105(.dina(w_n1399_0[0]),.dinb(w_n968_0[0]),.dout(n1407),.clk(gclk));
	jand g1106(.dina(w_dff_B_r0NRFXqF2_0),.dinb(n1406),.dout(n1408),.clk(gclk));
	jor g1107(.dina(n1408),.dinb(w_dff_B_z6nn5o6q1_1),.dout(n1409),.clk(gclk));
	jnot g1108(.din(w_n1409_0[1]),.dout(n1410),.clk(gclk));
	jxor g1109(.dina(w_n629_0[0]),.dinb(w_n625_0[0]),.dout(n1411),.clk(gclk));
	jnot g1110(.din(w_n1411_0[1]),.dout(n1412),.clk(gclk));
	jxor g1111(.dina(w_n806_0[1]),.dinb(w_n828_0[1]),.dout(n1413),.clk(gclk));
	jnot g1112(.din(w_n614_1[1]),.dout(n1414),.clk(gclk));
	jnot g1113(.din(w_n717_0[0]),.dout(n1415),.clk(gclk));
	jand g1114(.dina(w_n622_1[0]),.dinb(w_n828_0[0]),.dout(n1416),.clk(gclk));
	jand g1115(.dina(w_n628_0[0]),.dinb(w_G523_0[1]),.dout(n1417),.clk(gclk));
	jor g1116(.dina(n1417),.dinb(w_n829_0[0]),.dout(n1418),.clk(gclk));
	jor g1117(.dina(n1418),.dinb(n1416),.dout(n1419),.clk(gclk));
	jand g1118(.dina(n1419),.dinb(w_dff_B_Zfy0bBXR1_1),.dout(n1420),.clk(gclk));
	jxor g1119(.dina(w_n622_0[2]),.dinb(w_n618_0[1]),.dout(n1421),.clk(gclk));
	jnot g1120(.din(w_n1421_0[1]),.dout(n1422),.clk(gclk));
	jor g1121(.dina(w_dff_B_VoHCHtBi5_0),.dinb(n1420),.dout(n1423),.clk(gclk));
	jor g1122(.dina(w_n1421_0[0]),.dinb(w_n819_0[0]),.dout(n1424),.clk(gclk));
	jand g1123(.dina(n1424),.dinb(w_dff_B_2Lkh4R635_1),.dout(n1425),.clk(gclk));
	jxor g1124(.dina(w_n1425_0[1]),.dinb(w_dff_B_8XP8jZ1L9_1),.dout(n1426),.clk(gclk));
	jand g1125(.dina(n1426),.dinb(n1413),.dout(n1427),.clk(gclk));
	jnot g1126(.din(w_G2174_0[1]),.dout(n1428),.clk(gclk));
	jxor g1127(.dina(w_n806_0[0]),.dinb(w_n721_0[1]),.dout(n1429),.clk(gclk));
	jxor g1128(.dina(w_n1425_0[0]),.dinb(w_n614_1[0]),.dout(n1430),.clk(gclk));
	jand g1129(.dina(n1430),.dinb(n1429),.dout(n1431),.clk(gclk));
	jor g1130(.dina(n1431),.dinb(w_dff_B_02WrUaWC2_1),.dout(n1432),.clk(gclk));
	jor g1131(.dina(n1432),.dinb(w_dff_B_EeCOdrtz7_1),.dout(n1433),.clk(gclk));
	jxor g1132(.dina(w_n729_0[1]),.dinb(w_n614_0[2]),.dout(n1434),.clk(gclk));
	jnot g1133(.din(w_n1434_0[1]),.dout(n1435),.clk(gclk));
	jor g1134(.dina(w_n622_0[1]),.dinb(w_n721_0[0]),.dout(n1436),.clk(gclk));
	jand g1135(.dina(n1436),.dinb(w_n723_0[0]),.dout(n1437),.clk(gclk));
	jxor g1136(.dina(w_dff_B_wzRzGDvU7_0),.dinb(w_n727_0[0]),.dout(n1438),.clk(gclk));
	jand g1137(.dina(w_n1438_0[1]),.dinb(n1435),.dout(n1439),.clk(gclk));
	jnot g1138(.din(w_n1438_0[0]),.dout(n1440),.clk(gclk));
	jand g1139(.dina(w_dff_B_fKpEoIgw7_0),.dinb(w_n1434_0[0]),.dout(n1441),.clk(gclk));
	jor g1140(.dina(n1441),.dinb(w_G2174_0[0]),.dout(n1442),.clk(gclk));
	jor g1141(.dina(n1442),.dinb(n1439),.dout(n1443),.clk(gclk));
	jand g1142(.dina(w_dff_B_jNf0BP9R3_0),.dinb(n1433),.dout(n1444),.clk(gclk));
	jxor g1143(.dina(n1444),.dinb(w_n787_0[0]),.dout(n1445),.clk(gclk));
	jxor g1144(.dina(w_n1445_0[1]),.dinb(w_dff_B_LLiJKrcD2_1),.dout(n1446),.clk(gclk));
	jor g1145(.dina(w_n1446_0[1]),.dinb(w_n1410_0[1]),.dout(n1447),.clk(gclk));
	jxor g1146(.dina(w_n1445_0[0]),.dinb(w_n1411_0[0]),.dout(n1448),.clk(gclk));
	jor g1147(.dina(n1448),.dinb(w_n1409_0[0]),.dout(n1449),.clk(gclk));
	jand g1148(.dina(n1449),.dinb(w_G4091_1[1]),.dout(n1450),.clk(gclk));
	jand g1149(.dina(n1450),.dinb(w_n1447_0[1]),.dout(n1451),.clk(gclk));
	jor g1150(.dina(n1451),.dinb(w_dff_B_VJgNpd3v5_1),.dout(n1452),.clk(gclk));
	jand g1151(.dina(w_n1452_0[1]),.dinb(w_dff_B_EcgkE7Vz6_1),.dout(w_dff_A_WDxtKaJz2_2),.clk(gclk));
	jor g1152(.dina(w_G4091_1[0]),.dinb(G118),.dout(n1454),.clk(gclk));
	jand g1153(.dina(w_G251_2[2]),.dinb(w_n460_0[2]),.dout(n1455),.clk(gclk));
	jand g1154(.dina(w_G248_3[0]),.dinb(w_G234_1[0]),.dout(n1456),.clk(gclk));
	jor g1155(.dina(n1456),.dinb(w_n462_0[0]),.dout(n1457),.clk(gclk));
	jor g1156(.dina(n1457),.dinb(n1455),.dout(n1458),.clk(gclk));
	jand g1157(.dina(w_n366_2[2]),.dinb(w_n460_0[1]),.dout(n1459),.clk(gclk));
	jand g1158(.dina(w_n368_3[0]),.dinb(w_G234_0[2]),.dout(n1460),.clk(gclk));
	jor g1159(.dina(n1460),.dinb(w_G435_0[1]),.dout(n1461),.clk(gclk));
	jor g1160(.dina(n1461),.dinb(n1459),.dout(n1462),.clk(gclk));
	jand g1161(.dina(n1462),.dinb(n1458),.dout(n1463),.clk(gclk));
	jor g1162(.dina(w_n402_1[1]),.dinb(w_G226_1[0]),.dout(n1464),.clk(gclk));
	jor g1163(.dina(w_n405_1[1]),.dinb(w_n530_0[2]),.dout(n1465),.clk(gclk));
	jand g1164(.dina(n1465),.dinb(w_G422_0[2]),.dout(n1466),.clk(gclk));
	jand g1165(.dina(n1466),.dinb(n1464),.dout(n1467),.clk(gclk));
	jor g1166(.dina(w_G254_1[0]),.dinb(w_G226_0[2]),.dout(n1468),.clk(gclk));
	jor g1167(.dina(w_G242_1[0]),.dinb(w_n530_0[1]),.dout(n1469),.clk(gclk));
	jand g1168(.dina(n1469),.dinb(w_n532_0[0]),.dout(n1470),.clk(gclk));
	jand g1169(.dina(n1470),.dinb(n1468),.dout(n1471),.clk(gclk));
	jor g1170(.dina(n1471),.dinb(n1467),.dout(n1472),.clk(gclk));
	jxor g1171(.dina(n1472),.dinb(w_n528_0[0]),.dout(n1473),.clk(gclk));
	jor g1172(.dina(w_n402_1[0]),.dinb(w_G218_1[0]),.dout(n1474),.clk(gclk));
	jor g1173(.dina(w_n405_1[0]),.dinb(w_n507_0[2]),.dout(n1475),.clk(gclk));
	jand g1174(.dina(n1475),.dinb(w_G468_0[1]),.dout(n1476),.clk(gclk));
	jand g1175(.dina(n1476),.dinb(n1474),.dout(n1477),.clk(gclk));
	jor g1176(.dina(w_G254_0[2]),.dinb(w_G218_0[2]),.dout(n1478),.clk(gclk));
	jor g1177(.dina(w_G242_0[2]),.dinb(w_n507_0[1]),.dout(n1479),.clk(gclk));
	jand g1178(.dina(n1479),.dinb(w_n509_0[0]),.dout(n1480),.clk(gclk));
	jand g1179(.dina(n1480),.dinb(n1478),.dout(n1481),.clk(gclk));
	jor g1180(.dina(n1481),.dinb(n1477),.dout(n1482),.clk(gclk));
	jand g1181(.dina(w_G251_2[1]),.dinb(w_n541_0[2]),.dout(n1483),.clk(gclk));
	jand g1182(.dina(w_G248_2[2]),.dinb(w_G210_1[0]),.dout(n1484),.clk(gclk));
	jor g1183(.dina(n1484),.dinb(w_n543_0[0]),.dout(n1485),.clk(gclk));
	jor g1184(.dina(n1485),.dinb(n1483),.dout(n1486),.clk(gclk));
	jand g1185(.dina(w_n366_2[1]),.dinb(w_n541_0[1]),.dout(n1487),.clk(gclk));
	jand g1186(.dina(w_n368_2[2]),.dinb(w_G210_0[2]),.dout(n1488),.clk(gclk));
	jor g1187(.dina(n1488),.dinb(w_G457_0[2]),.dout(n1489),.clk(gclk));
	jor g1188(.dina(n1489),.dinb(n1487),.dout(n1490),.clk(gclk));
	jand g1189(.dina(n1490),.dinb(n1486),.dout(n1491),.clk(gclk));
	jxor g1190(.dina(n1491),.dinb(n1482),.dout(n1492),.clk(gclk));
	jxor g1191(.dina(n1492),.dinb(n1473),.dout(n1493),.clk(gclk));
	jxor g1192(.dina(n1493),.dinb(n1463),.dout(n1494),.clk(gclk));
	jand g1193(.dina(w_n495_0[2]),.dinb(w_G251_2[0]),.dout(n1495),.clk(gclk));
	jand g1194(.dina(w_G281_1[0]),.dinb(w_G248_2[1]),.dout(n1496),.clk(gclk));
	jor g1195(.dina(n1496),.dinb(w_n497_0[1]),.dout(n1497),.clk(gclk));
	jor g1196(.dina(n1497),.dinb(n1495),.dout(n1498),.clk(gclk));
	jand g1197(.dina(w_n495_0[1]),.dinb(w_n366_2[0]),.dout(n1499),.clk(gclk));
	jand g1198(.dina(w_G281_0[2]),.dinb(w_n368_2[1]),.dout(n1500),.clk(gclk));
	jor g1199(.dina(n1500),.dinb(w_G374_0[0]),.dout(n1501),.clk(gclk));
	jor g1200(.dina(n1501),.dinb(n1499),.dout(n1502),.clk(gclk));
	jand g1201(.dina(n1502),.dinb(n1498),.dout(n1503),.clk(gclk));
	jand g1202(.dina(w_n449_0[2]),.dinb(w_G251_1[2]),.dout(n1504),.clk(gclk));
	jand g1203(.dina(w_G265_1[0]),.dinb(w_G248_2[0]),.dout(n1505),.clk(gclk));
	jor g1204(.dina(n1505),.dinb(w_n451_0[1]),.dout(n1506),.clk(gclk));
	jor g1205(.dina(n1506),.dinb(n1504),.dout(n1507),.clk(gclk));
	jand g1206(.dina(w_n449_0[1]),.dinb(w_n366_1[2]),.dout(n1508),.clk(gclk));
	jand g1207(.dina(w_G265_0[2]),.dinb(w_n368_2[0]),.dout(n1509),.clk(gclk));
	jor g1208(.dina(n1509),.dinb(w_G400_0[1]),.dout(n1510),.clk(gclk));
	jor g1209(.dina(n1510),.dinb(n1508),.dout(n1511),.clk(gclk));
	jand g1210(.dina(n1511),.dinb(n1507),.dout(n1512),.clk(gclk));
	jxor g1211(.dina(n1512),.dinb(n1503),.dout(n1513),.clk(gclk));
	jor g1212(.dina(w_G257_1[0]),.dinb(w_n402_0[2]),.dout(n1514),.clk(gclk));
	jor g1213(.dina(w_n471_0[2]),.dinb(w_n405_0[2]),.dout(n1515),.clk(gclk));
	jand g1214(.dina(n1515),.dinb(w_G389_0[0]),.dout(n1516),.clk(gclk));
	jand g1215(.dina(n1516),.dinb(n1514),.dout(n1517),.clk(gclk));
	jor g1216(.dina(w_G257_0[2]),.dinb(w_G254_0[1]),.dout(n1518),.clk(gclk));
	jor g1217(.dina(w_n471_0[1]),.dinb(w_G242_0[1]),.dout(n1519),.clk(gclk));
	jand g1218(.dina(n1519),.dinb(w_n473_0[1]),.dout(n1520),.clk(gclk));
	jand g1219(.dina(n1520),.dinb(n1518),.dout(n1521),.clk(gclk));
	jor g1220(.dina(n1521),.dinb(n1517),.dout(n1522),.clk(gclk));
	jand g1221(.dina(w_n484_0[2]),.dinb(w_G251_1[1]),.dout(n1523),.clk(gclk));
	jand g1222(.dina(w_G273_1[0]),.dinb(w_G248_1[2]),.dout(n1524),.clk(gclk));
	jor g1223(.dina(n1524),.dinb(w_n486_0[1]),.dout(n1525),.clk(gclk));
	jor g1224(.dina(n1525),.dinb(n1523),.dout(n1526),.clk(gclk));
	jand g1225(.dina(w_n484_0[1]),.dinb(w_n366_1[1]),.dout(n1527),.clk(gclk));
	jand g1226(.dina(w_G273_0[2]),.dinb(w_n368_1[2]),.dout(n1528),.clk(gclk));
	jor g1227(.dina(n1528),.dinb(w_G411_0[0]),.dout(n1529),.clk(gclk));
	jor g1228(.dina(n1529),.dinb(n1527),.dout(n1530),.clk(gclk));
	jand g1229(.dina(n1530),.dinb(n1526),.dout(n1531),.clk(gclk));
	jxor g1230(.dina(n1531),.dinb(n1522),.dout(n1532),.clk(gclk));
	jxor g1231(.dina(n1532),.dinb(n1513),.dout(n1533),.clk(gclk));
	jand g1232(.dina(w_n1533_0[1]),.dinb(w_n1494_0[1]),.dout(n1534),.clk(gclk));
	jnot g1233(.din(n1534),.dout(n1535),.clk(gclk));
	jor g1234(.dina(w_n1533_0[0]),.dinb(w_n1494_0[0]),.dout(n1536),.clk(gclk));
	jand g1235(.dina(n1536),.dinb(w_n750_0[2]),.dout(n1537),.clk(gclk));
	jand g1236(.dina(n1537),.dinb(n1535),.dout(n1538),.clk(gclk));
	jor g1237(.dina(n1454),.dinb(w_n746_0[1]),.dout(n1539),.clk(gclk));
	jor g1238(.dina(n1538),.dinb(w_G4092_1[0]),.dout(n1540),.clk(gclk));
	jxor g1239(.dina(w_n583_0[1]),.dinb(w_n578_0[0]),.dout(n1541),.clk(gclk));
	jxor g1240(.dina(n1541),.dinb(w_n943_0[0]),.dout(n1542),.clk(gclk));
	jnot g1241(.din(n1542),.dout(n1543),.clk(gclk));
	jand g1242(.dina(w_n587_0[2]),.dinb(w_G1497_0[2]),.dout(n1544),.clk(gclk));
	jor g1243(.dina(n1544),.dinb(w_n696_0[0]),.dout(n1545),.clk(gclk));
	jnot g1244(.din(w_n1545_0[1]),.dout(n1546),.clk(gclk));
	jor g1245(.dina(w_n944_0[0]),.dinb(w_n930_0[1]),.dout(n1547),.clk(gclk));
	jand g1246(.dina(n1547),.dinb(w_n706_0[0]),.dout(n1548),.clk(gclk));
	jxor g1247(.dina(n1548),.dinb(w_n928_0[0]),.dout(n1549),.clk(gclk));
	jxor g1248(.dina(w_n605_1[1]),.dinb(w_n948_0[1]),.dout(n1550),.clk(gclk));
	jxor g1249(.dina(n1550),.dinb(n1549),.dout(n1551),.clk(gclk));
	jand g1250(.dina(n1551),.dinb(n1546),.dout(n1552),.clk(gclk));
	jxor g1251(.dina(w_n605_1[0]),.dinb(w_n703_0[0]),.dout(n1553),.clk(gclk));
	jand g1252(.dina(w_n605_0[2]),.dinb(w_n948_0[0]),.dout(n1554),.clk(gclk));
	jor g1253(.dina(n1554),.dinb(w_n702_0[0]),.dout(n1555),.clk(gclk));
	jnot g1254(.din(w_n1555_0[1]),.dout(n1556),.clk(gclk));
	jor g1255(.dina(n1556),.dinb(w_n930_0[0]),.dout(n1557),.clk(gclk));
	jor g1256(.dina(w_n1555_0[0]),.dinb(w_n707_0[0]),.dout(n1558),.clk(gclk));
	jand g1257(.dina(n1558),.dinb(n1557),.dout(n1559),.clk(gclk));
	jxor g1258(.dina(n1559),.dinb(w_n596_0[0]),.dout(n1560),.clk(gclk));
	jand g1259(.dina(w_n1560_0[1]),.dinb(w_n1553_0[1]),.dout(n1561),.clk(gclk));
	jnot g1260(.din(n1561),.dout(n1562),.clk(gclk));
	jor g1261(.dina(w_n1560_0[0]),.dinb(w_n1553_0[0]),.dout(n1563),.clk(gclk));
	jand g1262(.dina(n1563),.dinb(w_n1545_0[0]),.dout(n1564),.clk(gclk));
	jand g1263(.dina(n1564),.dinb(n1562),.dout(n1565),.clk(gclk));
	jor g1264(.dina(n1565),.dinb(n1552),.dout(n1566),.clk(gclk));
	jnot g1265(.din(w_G1497_0[1]),.dout(n1567),.clk(gclk));
	jand g1266(.dina(w_n682_0[0]),.dinb(w_n687_0[0]),.dout(n1568),.clk(gclk));
	jand g1267(.dina(w_n1568_0[1]),.dinb(w_n574_0[0]),.dout(n1569),.clk(gclk));
	jxor g1268(.dina(n1569),.dinb(w_n561_0[1]),.dout(n1570),.clk(gclk));
	jxor g1269(.dina(w_n572_0[1]),.dinb(w_n681_1[1]),.dout(n1571),.clk(gclk));
	jor g1270(.dina(w_n856_0[0]),.dinb(w_n853_0[0]),.dout(n1572),.clk(gclk));
	jand g1271(.dina(w_n693_0[1]),.dinb(w_n585_0[0]),.dout(n1573),.clk(gclk));
	jor g1272(.dina(n1573),.dinb(w_n855_0[0]),.dout(n1574),.clk(gclk));
	jand g1273(.dina(n1574),.dinb(n1572),.dout(n1575),.clk(gclk));
	jxor g1274(.dina(n1575),.dinb(n1571),.dout(n1576),.clk(gclk));
	jxor g1275(.dina(n1576),.dinb(n1570),.dout(n1577),.clk(gclk));
	jor g1276(.dina(n1577),.dinb(n1567),.dout(n1578),.clk(gclk));
	jxor g1277(.dina(w_n693_0[0]),.dinb(w_n572_0[0]),.dout(n1579),.clk(gclk));
	jor g1278(.dina(w_n857_0[0]),.dinb(w_n681_1[0]),.dout(n1580),.clk(gclk));
	jnot g1279(.din(w_n681_0[2]),.dout(n1581),.clk(gclk));
	jor g1280(.dina(w_n680_0[0]),.dinb(n1581),.dout(n1582),.clk(gclk));
	jor g1281(.dina(n1582),.dinb(w_n689_0[0]),.dout(n1583),.clk(gclk));
	jxor g1282(.dina(n1583),.dinb(w_n567_0[1]),.dout(n1584),.clk(gclk));
	jand g1283(.dina(n1584),.dinb(n1580),.dout(n1585),.clk(gclk));
	jxor g1284(.dina(w_n1568_0[0]),.dinb(w_n561_0[0]),.dout(n1586),.clk(gclk));
	jxor g1285(.dina(n1586),.dinb(n1585),.dout(n1587),.clk(gclk));
	jxor g1286(.dina(n1587),.dinb(n1579),.dout(n1588),.clk(gclk));
	jor g1287(.dina(n1588),.dinb(w_G1497_0[0]),.dout(n1589),.clk(gclk));
	jand g1288(.dina(n1589),.dinb(n1578),.dout(n1590),.clk(gclk));
	jxor g1289(.dina(n1590),.dinb(n1566),.dout(n1591),.clk(gclk));
	jand g1290(.dina(w_n1591_0[1]),.dinb(w_n1543_0[1]),.dout(n1592),.clk(gclk));
	jnot g1291(.din(n1592),.dout(n1593),.clk(gclk));
	jor g1292(.dina(w_n1591_0[0]),.dinb(w_n1543_0[0]),.dout(n1594),.clk(gclk));
	jand g1293(.dina(n1594),.dinb(w_G4091_0[2]),.dout(n1595),.clk(gclk));
	jand g1294(.dina(n1595),.dinb(n1593),.dout(n1596),.clk(gclk));
	jor g1295(.dina(n1596),.dinb(n1540),.dout(n1597),.clk(gclk));
	jand g1296(.dina(w_n1597_0[1]),.dinb(w_dff_B_aFV8wzDx3_1),.dout(w_dff_A_73tBNL023_2),.clk(gclk));
	jand g1297(.dina(w_G4092_0[2]),.dinb(G97),.dout(n1599),.clk(gclk));
	jnot g1298(.din(n1599),.dout(n1600),.clk(gclk));
	jand g1299(.dina(n1600),.dinb(w_n1597_0[0]),.dout(n1601),.clk(gclk));
	jnot g1300(.din(w_n1601_0[2]),.dout(n1602),.clk(gclk));
	jand g1301(.dina(w_n1602_0[1]),.dinb(w_n793_1[1]),.dout(n1603),.clk(gclk));
	jnot g1302(.din(w_n1447_0[0]),.dout(n1604),.clk(gclk));
	jand g1303(.dina(w_n1446_0[0]),.dinb(w_n1410_0[0]),.dout(n1605),.clk(gclk));
	jor g1304(.dina(n1605),.dinb(w_n750_0[1]),.dout(n1606),.clk(gclk));
	jor g1305(.dina(n1606),.dinb(n1604),.dout(n1607),.clk(gclk));
	jand g1306(.dina(n1607),.dinb(w_n1391_0[0]),.dout(n1608),.clk(gclk));
	jand g1307(.dina(w_G4092_0[1]),.dinb(G94),.dout(n1609),.clk(gclk));
	jor g1308(.dina(w_n1609_0[1]),.dinb(n1608),.dout(n1610),.clk(gclk));
	jand g1309(.dina(w_n1610_0[1]),.dinb(w_n797_1[1]),.dout(n1611),.clk(gclk));
	jand g1310(.dina(w_n799_1[1]),.dinb(w_G14_0[1]),.dout(n1612),.clk(gclk));
	jand g1311(.dina(w_n801_1[1]),.dinb(w_G64_0[1]),.dout(n1613),.clk(gclk));
	jor g1312(.dina(n1613),.dinb(n1612),.dout(n1614),.clk(gclk));
	jor g1313(.dina(w_dff_B_vgKwEqZe7_0),.dinb(n1611),.dout(n1615),.clk(gclk));
	jor g1314(.dina(n1615),.dinb(n1603),.dout(w_dff_A_hMdQYkwo2_2),.clk(gclk));
	jand g1315(.dina(w_n1602_0[0]),.dinb(w_n840_1[1]),.dout(n1617),.clk(gclk));
	jand g1316(.dina(w_n1610_0[0]),.dinb(w_n843_1[1]),.dout(n1618),.clk(gclk));
	jand g1317(.dina(w_n845_1[1]),.dinb(w_G14_0[0]),.dout(n1619),.clk(gclk));
	jand g1318(.dina(w_n847_1[1]),.dinb(w_G64_0[0]),.dout(n1620),.clk(gclk));
	jor g1319(.dina(n1620),.dinb(n1619),.dout(n1621),.clk(gclk));
	jor g1320(.dina(w_dff_B_e5vsVdSQ9_0),.dinb(n1618),.dout(n1622),.clk(gclk));
	jor g1321(.dina(n1622),.dinb(n1617),.dout(w_dff_A_IsWFdUh62_2),.clk(gclk));
	jnot g1322(.din(w_G137_3[1]),.dout(n1624),.clk(gclk));
	jnot g1323(.din(w_n985_1[1]),.dout(n1625),.clk(gclk));
	jor g1324(.dina(w_n1601_0[1]),.dinb(n1625),.dout(n1626),.clk(gclk));
	jnot g1325(.din(w_n988_1[1]),.dout(n1627),.clk(gclk));
	jnot g1326(.din(w_n1609_0[0]),.dout(n1628),.clk(gclk));
	jand g1327(.dina(w_dff_B_turOlrt26_0),.dinb(w_n1452_0[0]),.dout(n1629),.clk(gclk));
	jor g1328(.dina(w_n1629_0[1]),.dinb(w_dff_B_e33LovgP0_1),.dout(n1630),.clk(gclk));
	jnot g1329(.din(G179),.dout(n1631),.clk(gclk));
	jnot g1330(.din(w_n992_1[1]),.dout(n1632),.clk(gclk));
	jor g1331(.dina(n1632),.dinb(w_n1631_0[1]),.dout(n1633),.clk(gclk));
	jnot g1332(.din(G176),.dout(n1634),.clk(gclk));
	jnot g1333(.din(w_n990_1[1]),.dout(n1635),.clk(gclk));
	jor g1334(.dina(n1635),.dinb(w_n1634_0[1]),.dout(n1636),.clk(gclk));
	jand g1335(.dina(n1636),.dinb(n1633),.dout(n1637),.clk(gclk));
	jand g1336(.dina(w_dff_B_bVZczMbx8_0),.dinb(n1630),.dout(n1638),.clk(gclk));
	jand g1337(.dina(n1638),.dinb(w_dff_B_Xoebksbe1_1),.dout(n1639),.clk(gclk));
	jor g1338(.dina(n1639),.dinb(w_n1624_0[1]),.dout(G658),.clk(gclk));
	jnot g1339(.din(w_n999_1[1]),.dout(n1641),.clk(gclk));
	jor g1340(.dina(w_n1601_0[0]),.dinb(n1641),.dout(n1642),.clk(gclk));
	jnot g1341(.din(w_n1002_1[1]),.dout(n1643),.clk(gclk));
	jor g1342(.dina(w_n1629_0[0]),.dinb(w_dff_B_bZbagBGo7_1),.dout(n1644),.clk(gclk));
	jnot g1343(.din(w_n1006_1[1]),.dout(n1645),.clk(gclk));
	jor g1344(.dina(n1645),.dinb(w_n1631_0[0]),.dout(n1646),.clk(gclk));
	jnot g1345(.din(w_n1004_1[1]),.dout(n1647),.clk(gclk));
	jor g1346(.dina(n1647),.dinb(w_n1634_0[0]),.dout(n1648),.clk(gclk));
	jand g1347(.dina(n1648),.dinb(n1646),.dout(n1649),.clk(gclk));
	jand g1348(.dina(w_dff_B_5W8CGx180_0),.dinb(n1644),.dout(n1650),.clk(gclk));
	jand g1349(.dina(n1650),.dinb(w_dff_B_ddURQ7Dr9_1),.dout(n1651),.clk(gclk));
	jor g1350(.dina(n1651),.dinb(w_n1624_0[0]),.dout(G690),.clk(gclk));
	jdff g1351(.din(w_G141_1[0]),.dout(w_dff_A_L8i6nSmj8_1));
	jdff g1352(.din(w_G293_0[0]),.dout(w_dff_A_xzFbqVFy4_1));
	jdff g1353(.din(w_G3173_0[0]),.dout(w_dff_A_MwhKPAJt6_1));
	jnot g1354(.din(w_G545_0[1]),.dout(w_dff_A_gr7tdRmi6_1),.clk(gclk));
	jnot g1355(.din(w_G545_0[0]),.dout(w_dff_A_OUjptODI7_1),.clk(gclk));
	jdff g1356(.din(w_G137_3[0]),.dout(w_dff_A_sj71NC4V1_1));
	jdff g1357(.din(w_G141_0[2]),.dout(w_dff_A_HaCj6xuk2_1));
	jdff g1358(.din(w_G1_2[0]),.dout(w_dff_A_n3PHt2IB0_1));
	jdff g1359(.din(w_G549_0[1]),.dout(w_dff_A_Gx44yVSc7_1));
	jdff g1360(.din(w_G299_0[1]),.dout(w_dff_A_omMcWl0V5_1));
	jnot g1361(.din(w_G549_0[0]),.dout(w_dff_A_KkjYaiEQ9_1),.clk(gclk));
	jdff g1362(.din(w_G1_1[2]),.dout(w_dff_A_souf8wzQ9_1));
	jdff g1363(.din(w_G1_1[1]),.dout(w_dff_A_ezKNDcPo0_1));
	jdff g1364(.din(w_G1_1[0]),.dout(w_dff_A_FmBKNEEe6_1));
	jdff g1365(.din(w_G1_0[2]),.dout(w_dff_A_nZRgG5262_1));
	jdff g1366(.din(w_G299_0[0]),.dout(w_dff_A_eXIkQR0I3_1));
	jor g1367(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(w_dff_A_uUv6KBve7_2),.clk(gclk));
	jand g1368(.dina(w_n652_0[0]),.dinb(w_n633_0[1]),.dout(w_dff_A_VtM4hs6P0_2),.clk(gclk));
	jand g1369(.dina(w_n607_0[0]),.dinb(w_n587_0[1]),.dout(w_dff_A_tughExAl8_2),.clk(gclk));
	jor g1370(.dina(w_n709_0[0]),.dinb(w_n697_0[0]),.dout(w_dff_A_xNiLG5rl1_2),.clk(gclk));
	jor g1371(.dina(w_n742_0[0]),.dinb(w_n733_0[0]),.dout(w_dff_A_ePXT8ufG1_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_G4_0[1]),.doutc(w_G4_0[2]),.din(G4));
	jspl jspl_w_G4_1(.douta(w_G4_1[0]),.doutb(w_G4_1[1]),.din(w_G4_0[0]));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(G11));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(G14));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(G17));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(G20));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(G37));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(G40));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(G43));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(G46));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(G49));
	jspl jspl_w_G54_0(.douta(w_G54_0[0]),.doutb(w_G54_0[1]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(G61));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(G64));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(G67));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(G70));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(G73));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(G76));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(G91));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(G100));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(G103));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(G106));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(G109));
	jspl jspl_w_G123_0(.douta(w_G123_0[0]),.doutb(w_G123_0[1]),.din(G123));
	jspl jspl_w_G132_0(.douta(w_dff_A_W3xZVqvd4_0),.doutb(w_G132_0[1]),.din(w_dff_B_06mJDRfX3_2));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_iq7Ngik62_0),.doutb(w_dff_A_UZnqtXha6_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_j8iNbbck6_0),.doutb(w_dff_A_0Jc3Av869_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_G137_3[2]),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_dff_A_jocxXTXK8_0),.doutb(w_dff_A_QabQwMds8_1),.doutc(w_G137_4[2]),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_dff_A_qJgKLL8u9_0),.doutb(w_G137_5[1]),.doutc(w_G137_5[2]),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_aTLt1TvC9_0),.doutb(w_dff_A_gnvf12y66_1),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_VV06EGpu8_1),.doutc(w_dff_A_dScTuOOL0_2),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_dff_A_OlofKs7A9_0),.doutb(w_G137_8[1]),.doutc(w_dff_A_WB8BAewC6_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_G137_9[0]),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_TiUCt4UZ9_1),.doutc(w_dff_A_c4hnKAkf8_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_Q4mVXVSm9_0),.doutb(w_dff_A_IVtEBFxm4_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(G146));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(G149));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(G152));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(G155));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(G158));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(G161));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(G164));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(G167));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(G170));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(G173));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(G182));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(G185));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(G188));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(G191));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(G194));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(G197));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(G200));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(G203));
	jspl3 jspl3_w_G206_0(.douta(w_G206_0[0]),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_G210_0[2]),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_G210_1[1]),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl3 jspl3_w_G210_2(.douta(w_G210_2[0]),.doutb(w_G210_2[1]),.doutc(w_G210_2[2]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_G218_1[0]),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl3 jspl3_w_G218_2(.douta(w_G218_2[0]),.doutb(w_G218_2[1]),.doutc(w_G218_2[2]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_G226_0[2]),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_G226_1[0]),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G226_2(.douta(w_G226_2[0]),.doutb(w_G226_2[1]),.doutc(w_G226_2[2]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_G234_0[2]),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_G234_2[0]),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_G242_0[1]),.doutc(w_G242_0[2]),.din(G242));
	jspl3 jspl3_w_G242_1(.douta(w_G242_1[0]),.doutb(w_G242_1[1]),.doutc(w_G242_1[2]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_G245_0[0]),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_G248_3[2]),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl jspl_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_G251_0[1]),.doutc(w_G251_0[2]),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_G251_1[0]),.doutb(w_G251_1[1]),.doutc(w_G251_1[2]),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_G251_4[1]),.doutc(w_G251_4[2]),.din(w_G251_1[0]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl3 jspl3_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.doutc(w_G254_1[2]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_G257_0[2]),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_G257_1[0]),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G257_2(.douta(w_G257_2[0]),.doutb(w_G257_2[1]),.doutc(w_G257_2[2]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_G265_0[2]),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_G265_1[1]),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl jspl_w_G265_2(.douta(w_G265_2[0]),.doutb(w_G265_2[1]),.din(w_G265_0[1]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_G273_0[2]),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_G273_1[1]),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl3 jspl3_w_G273_2(.douta(w_G273_2[0]),.doutb(w_G273_2[1]),.doutc(w_G273_2[2]),.din(w_G273_0[1]));
	jspl jspl_w_G280_0(.douta(w_G280_0[0]),.doutb(w_G280_0[1]),.din(G280));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_G281_0[2]),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_G281_2[0]),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_G289_0[0]),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_G293_0[1]),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_G302_0[0]),.doutb(w_G302_0[1]),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_G308_1[0]),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_G316_0[2]),.din(G316));
	jspl3 jspl3_w_G316_1(.douta(w_G316_1[0]),.doutb(w_G316_1[1]),.doutc(w_G316_1[2]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_G324_0[1]),.doutc(w_G324_0[2]),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_G324_1[1]),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_G331_0[1]),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_G332_1[1]),.doutc(w_G332_1[2]),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_G332_2[0]),.doutb(w_G332_2[1]),.doutc(w_G332_2[2]),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_G332_3[0]),.doutb(w_G332_3[1]),.doutc(w_G332_3[2]),.din(w_G332_0[2]));
	jspl3 jspl3_w_G332_4(.douta(w_G332_4[0]),.doutb(w_G332_4[1]),.doutc(w_G332_4[2]),.din(w_G332_1[0]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl3 jspl3_w_G335_1(.douta(w_G335_1[0]),.doutb(w_G335_1[1]),.doutc(w_G335_1[2]),.din(w_G335_0[0]));
	jspl3 jspl3_w_G335_2(.douta(w_G335_2[0]),.doutb(w_G335_2[1]),.doutc(w_G335_2[2]),.din(w_G335_0[1]));
	jspl3 jspl3_w_G335_3(.douta(w_G335_3[0]),.doutb(w_G335_3[1]),.doutc(w_G335_3[2]),.din(w_G335_0[2]));
	jspl jspl_w_G335_4(.douta(w_G335_4[0]),.doutb(w_G335_4[1]),.din(w_G335_1[0]));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_G341_0[2]),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_G341_2[1]),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_G348_0[0]),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_G351_0[2]),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_G351_1[0]),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_G351_2[1]),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_G358_0[0]),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_G361_0[1]),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G369_0(.douta(w_G369_0[0]),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_G374_0[0]),.doutb(w_G374_0[1]),.doutc(w_G374_0[2]),.din(G374));
	jspl3 jspl3_w_G389_0(.douta(w_G389_0[0]),.doutb(w_G389_0[1]),.doutc(w_G389_0[2]),.din(G389));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_G400_0[1]),.doutc(w_G400_0[2]),.din(G400));
	jspl jspl_w_G400_1(.douta(w_G400_1[0]),.doutb(w_G400_1[1]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_G411_0[0]),.doutb(w_G411_0[1]),.doutc(w_G411_0[2]),.din(G411));
	jspl3 jspl3_w_G422_0(.douta(w_G422_0[0]),.doutb(w_G422_0[1]),.doutc(w_G422_0[2]),.din(G422));
	jspl3 jspl3_w_G422_1(.douta(w_G422_1[0]),.doutb(w_G422_1[1]),.doutc(w_G422_1[2]),.din(w_G422_0[0]));
	jspl jspl_w_G422_2(.douta(w_G422_2[0]),.doutb(w_G422_2[1]),.din(w_G422_0[1]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_G435_0[1]),.doutc(w_G435_0[2]),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_G435_1[0]),.doutb(w_G435_1[1]),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_G446_0[1]),.doutc(w_G446_0[2]),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_G446_1[0]),.doutb(w_G446_1[1]),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_G457_0[0]),.doutb(w_G457_0[1]),.doutc(w_G457_0[2]),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_G457_1[0]),.doutb(w_G457_1[1]),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl jspl_w_G457_2(.douta(w_G457_2[0]),.doutb(w_G457_2[1]),.din(w_G457_0[1]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_G468_0[1]),.doutc(w_G468_0[2]),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_G468_1[0]),.doutb(w_G468_1[1]),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_G479_0[0]),.doutb(w_G479_0[1]),.doutc(w_G479_0[2]),.din(G479));
	jspl jspl_w_G479_1(.douta(w_G479_1[0]),.doutb(w_G479_1[1]),.din(w_G479_0[0]));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_G490_0[1]),.doutc(w_G490_0[2]),.din(G490));
	jspl3 jspl3_w_G490_1(.douta(w_G490_1[0]),.doutb(w_G490_1[1]),.doutc(w_G490_1[2]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_G503_0[0]),.doutb(w_G503_0[1]),.doutc(w_G503_0[2]),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_G503_1[0]),.doutb(w_G503_1[1]),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl3 jspl3_w_G514_0(.douta(w_G514_0[0]),.doutb(w_G514_0[1]),.doutc(w_G514_0[2]),.din(G514));
	jspl jspl_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.din(w_G514_0[0]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_G523_0[1]),.doutc(w_G523_0[2]),.din(G523));
	jspl jspl_w_G523_1(.douta(w_G523_1[0]),.doutb(w_G523_1[1]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_G534_0[0]),.doutb(w_G534_0[1]),.doutc(w_G534_0[2]),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_G534_1[0]),.doutb(w_G534_1[1]),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_G559_0[0]),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_G1497_0[0]),.doutb(w_G1497_0[1]),.doutc(w_G1497_0[2]),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_G1689_0[1]),.doutc(w_G1689_0[2]),.din(G1689));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_G1690_0[1]),.doutc(w_G1690_0[2]),.din(G1690));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_G1691_0[1]),.doutc(w_G1691_0[2]),.din(G1691));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_G1694_0[1]),.doutc(w_G1694_0[2]),.din(G1694));
	jspl3 jspl3_w_G2174_0(.douta(w_G2174_0[0]),.doutb(w_G2174_0[1]),.doutc(w_G2174_0[2]),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_G2358_2[0]),.doutb(w_G2358_2[1]),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(G3548));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_G3717_0[0]),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_G3724_0[0]),.doutb(w_G3724_0[1]),.doutc(w_G3724_0[2]),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_G4087_0[1]),.doutc(w_G4087_0[2]),.din(G4087));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_G4088_0[2]),.din(G4088));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_G4089_0[2]),.din(G4089));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_G4090_0[1]),.doutc(w_G4090_0[2]),.din(G4090));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_G4091_0[1]),.doutc(w_G4091_0[2]),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_G4091_1[0]),.doutb(w_G4091_1[1]),.doutc(w_G4091_1[2]),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_G4091_2[0]),.doutb(w_G4091_2[1]),.doutc(w_G4091_2[2]),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_G4092_0[1]),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_G4092_1[0]),.doutb(w_G4092_1[1]),.doutc(w_G4092_1[2]),.din(w_G4092_0[0]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(w_dff_A_bSb3TJii9_1),.din(G599_fa_));
	jspl jspl_w_G600_0(.douta(w_G600_0),.doutb(w_dff_A_1FoVNhmo2_1),.din(G600_fa_));
	jspl jspl_w_G601_0(.douta(w_dff_A_Ie9xyNkC3_0),.doutb(w_dff_A_5HCiJFb58_1),.din(G601_fa_));
	jspl jspl_w_G611_0(.douta(w_G611_0),.doutb(w_dff_A_FJjvtOnm3_1),.din(G611_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(w_dff_A_HPCQADGE6_1),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_G809_1[0]),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_G809_2[2]),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_G809_3[0]),.doutb(w_G809_3[1]),.doutc(w_dff_A_j3HNxQs77_2),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(w_dff_A_KMUkwXSO1_1),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(w_dff_A_RYzzMdAy5_1),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(w_dff_A_E3YaYj4k1_1),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(w_dff_A_A4wx6Pyj7_1),.din(G861_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(w_dff_A_uwSrejso2_1),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(w_dff_A_aPDiXqIJ5_1),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(w_dff_A_oZ7aU2kK3_1),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(w_dff_A_FEyi87VO8_1),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(w_dff_A_tbRIqskU5_1),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(w_dff_A_mfZM6VHe2_1),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(w_dff_A_znHZByz42_1),.din(G877_fa_));
	jspl jspl_w_G1000_0(.douta(w_G1000_0),.doutb(w_dff_A_BMw7y2Ba7_1),.din(G1000_fa_));
	jspl jspl_w_G826_0(.douta(w_G826_0),.doutb(w_dff_A_eohpnt6F6_1),.din(G826_fa_));
	jspl jspl_w_G828_0(.douta(w_G828_0),.doutb(w_dff_A_0qERABzF8_1),.din(G828_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(w_dff_A_ouuG4aRI7_1),.din(G830_fa_));
	jspl jspl_w_G867_0(.douta(w_G867_0),.doutb(w_dff_A_gLMnYhGz8_1),.din(G867_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(w_dff_A_p0X5p3Tl8_1),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(w_dff_B_FWUboPEb9_2));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n366_2(.douta(w_n366_2[0]),.doutb(w_n366_2[1]),.doutc(w_n366_2[2]),.din(w_n366_0[1]));
	jspl3 jspl3_w_n366_3(.douta(w_n366_3[0]),.doutb(w_n366_3[1]),.doutc(w_n366_3[2]),.din(w_n366_0[2]));
	jspl3 jspl3_w_n366_4(.douta(w_n366_4[0]),.doutb(w_n366_4[1]),.doutc(w_n366_4[2]),.din(w_n366_1[0]));
	jspl3 jspl3_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.doutc(w_n368_0[2]),.din(n368));
	jspl3 jspl3_w_n368_1(.douta(w_n368_1[0]),.doutb(w_n368_1[1]),.doutc(w_n368_1[2]),.din(w_n368_0[0]));
	jspl3 jspl3_w_n368_2(.douta(w_n368_2[0]),.doutb(w_n368_2[1]),.doutc(w_n368_2[2]),.din(w_n368_0[1]));
	jspl3 jspl3_w_n368_3(.douta(w_n368_3[0]),.doutb(w_n368_3[1]),.doutc(w_n368_3[2]),.din(w_n368_0[2]));
	jspl3 jspl3_w_n368_4(.douta(w_n368_4[0]),.doutb(w_n368_4[1]),.doutc(w_n368_4[2]),.din(w_n368_1[0]));
	jspl jspl_w_n368_5(.douta(w_n368_5[0]),.doutb(w_n368_5[1]),.din(w_n368_1[1]));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.doutc(w_n372_0[2]),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl3 jspl3_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.doutc(w_n385_1[2]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n386_1(.douta(w_n386_1[0]),.doutb(w_n386_1[1]),.doutc(w_n386_1[2]),.din(w_n386_0[0]));
	jspl3 jspl3_w_n386_2(.douta(w_n386_2[0]),.doutb(w_n386_2[1]),.doutc(w_n386_2[2]),.din(w_n386_0[1]));
	jspl3 jspl3_w_n386_3(.douta(w_n386_3[0]),.doutb(w_n386_3[1]),.doutc(w_n386_3[2]),.din(w_n386_0[2]));
	jspl3 jspl3_w_n386_4(.douta(w_n386_4[0]),.doutb(w_n386_4[1]),.doutc(w_n386_4[2]),.din(w_n386_1[0]));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_n388_0[2]),.din(n388));
	jspl3 jspl3_w_n388_1(.douta(w_n388_1[0]),.doutb(w_n388_1[1]),.doutc(w_n388_1[2]),.din(w_n388_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_n389_0[2]),.din(n389));
	jspl3 jspl3_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.doutc(w_n389_1[2]),.din(w_n389_0[0]));
	jspl3 jspl3_w_n389_2(.douta(w_n389_2[0]),.doutb(w_n389_2[1]),.doutc(w_n389_2[2]),.din(w_n389_0[1]));
	jspl3 jspl3_w_n389_3(.douta(w_n389_3[0]),.doutb(w_n389_3[1]),.doutc(w_n389_3[2]),.din(w_n389_0[2]));
	jspl3 jspl3_w_n389_4(.douta(w_n389_4[0]),.doutb(w_n389_4[1]),.doutc(w_n389_4[2]),.din(w_n389_1[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl3 jspl3_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.doutc(w_n398_0[2]),.din(n398));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n402_1(.douta(w_n402_1[0]),.doutb(w_n402_1[1]),.doutc(w_n402_1[2]),.din(w_n402_0[0]));
	jspl jspl_w_n402_2(.douta(w_n402_2[0]),.doutb(w_n402_2[1]),.din(w_n402_0[1]));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl3 jspl3_w_n405_1(.douta(w_n405_1[0]),.doutb(w_n405_1[1]),.doutc(w_n405_1[2]),.din(w_n405_0[0]));
	jspl jspl_w_n405_2(.douta(w_n405_2[0]),.doutb(w_n405_2[1]),.din(w_n405_0[1]));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_n410_0[2]),.din(n410));
	jspl jspl_w_n410_1(.douta(w_n410_1[0]),.doutb(w_n410_1[1]),.din(w_n410_0[0]));
	jspl jspl_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.din(n414));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(n416));
	jspl3 jspl3_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.doutc(w_n419_0[2]),.din(n419));
	jspl3 jspl3_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.doutc(w_n424_0[2]),.din(n424));
	jspl3 jspl3_w_n424_1(.douta(w_n424_1[0]),.doutb(w_n424_1[1]),.doutc(w_n424_1[2]),.din(w_n424_0[0]));
	jspl jspl_w_n424_2(.douta(w_n424_2[0]),.doutb(w_n424_2[1]),.din(w_n424_0[1]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl3 jspl3_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.doutc(w_n437_0[2]),.din(n437));
	jspl3 jspl3_w_n437_1(.douta(w_n437_1[0]),.doutb(w_n437_1[1]),.doutc(w_n437_1[2]),.din(w_n437_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_n451_0[0]),.doutb(w_n451_0[1]),.doutc(w_n451_0[2]),.din(n451));
	jspl jspl_w_n451_1(.douta(w_n451_1[0]),.doutb(w_n451_1[1]),.din(w_n451_0[0]));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl jspl_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.doutc(w_n473_0[2]),.din(n473));
	jspl3 jspl3_w_n473_1(.douta(w_n473_1[0]),.doutb(w_n473_1[1]),.doutc(w_n473_1[2]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.doutc(w_n484_0[2]),.din(n484));
	jspl jspl_w_n484_1(.douta(w_n484_1[0]),.doutb(w_n484_1[1]),.din(w_n484_0[0]));
	jspl3 jspl3_w_n486_0(.douta(w_n486_0[0]),.doutb(w_n486_0[1]),.doutc(w_n486_0[2]),.din(n486));
	jspl jspl_w_n486_1(.douta(w_n486_1[0]),.doutb(w_n486_1[1]),.din(w_n486_0[0]));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl3 jspl3_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.doutc(w_n495_0[2]),.din(n495));
	jspl3 jspl3_w_n495_1(.douta(w_n495_1[0]),.doutb(w_n495_1[1]),.doutc(w_n495_1[2]),.din(w_n495_0[0]));
	jspl3 jspl3_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.doutc(w_n497_0[2]),.din(n497));
	jspl jspl_w_n497_1(.douta(w_n497_1[0]),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl jspl_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.din(w_n507_0[0]));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(n509));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl jspl_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.doutc(w_n528_0[2]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl jspl_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.din(w_n530_0[0]));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(n532));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl3 jspl3_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.doutc(w_n541_0[2]),.din(n541));
	jspl jspl_w_n541_1(.douta(w_n541_1[0]),.doutb(w_n541_1[1]),.din(w_n541_0[0]));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl jspl_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl jspl_w_n560_1(.douta(w_n560_1[0]),.doutb(w_n560_1[1]),.din(w_n560_0[0]));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n567_1(.douta(w_n567_1[0]),.doutb(w_n567_1[1]),.din(w_n567_0[0]));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.din(n569));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_n571_0[2]),.din(n571));
	jspl jspl_w_n571_1(.douta(w_n571_1[0]),.doutb(w_n571_1[1]),.din(w_n571_0[0]));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.doutc(w_n577_0[2]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.doutc(w_n578_0[2]),.din(n578));
	jspl3 jspl3_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.doutc(w_n582_0[2]),.din(n582));
	jspl jspl_w_n582_1(.douta(w_n582_1[0]),.doutb(w_n582_1[1]),.din(w_n582_0[0]));
	jspl3 jspl3_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.doutc(w_n583_0[2]),.din(n583));
	jspl jspl_w_n583_1(.douta(w_n583_1[0]),.doutb(w_n583_1[1]),.din(w_n583_0[0]));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.doutc(w_n587_0[2]),.din(n587));
	jspl jspl_w_n587_1(.douta(w_n587_1[0]),.doutb(w_n587_1[1]),.din(w_n587_0[0]));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.doutc(w_n590_0[2]),.din(n590));
	jspl jspl_w_n590_1(.douta(w_n590_1[0]),.doutb(w_n590_1[1]),.din(w_n590_0[0]));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.doutc(w_n595_0[2]),.din(n595));
	jspl jspl_w_n595_1(.douta(w_n595_1[0]),.doutb(w_n595_1[1]),.din(w_n595_0[0]));
	jspl3 jspl3_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl3 jspl3_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.doutc(w_n600_0[2]),.din(n600));
	jspl jspl_w_n600_1(.douta(w_n600_1[0]),.doutb(w_n600_1[1]),.din(w_n600_0[0]));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl3 jspl3_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.doutc(w_n604_0[2]),.din(n604));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_n605_1[2]),.din(w_n605_0[0]));
	jspl3 jspl3_w_n605_2(.douta(w_n605_2[0]),.doutb(w_n605_2[1]),.doutc(w_n605_2[2]),.din(w_n605_0[1]));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.doutc(w_n607_0[2]),.din(n607));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n609_1(.douta(w_n609_1[0]),.doutb(w_n609_1[1]),.doutc(w_n609_1[2]),.din(w_n609_0[0]));
	jspl3 jspl3_w_n609_2(.douta(w_n609_2[0]),.doutb(w_n609_2[1]),.doutc(w_n609_2[2]),.din(w_n609_0[1]));
	jspl3 jspl3_w_n609_3(.douta(w_n609_3[0]),.doutb(w_n609_3[1]),.doutc(w_n609_3[2]),.din(w_n609_0[2]));
	jspl3 jspl3_w_n609_4(.douta(w_n609_4[0]),.doutb(w_n609_4[1]),.doutc(w_n609_4[2]),.din(w_n609_1[0]));
	jspl3 jspl3_w_n609_5(.douta(w_n609_5[0]),.doutb(w_n609_5[1]),.doutc(w_n609_5[2]),.din(w_n609_1[1]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.doutc(w_n614_0[2]),.din(n614));
	jspl3 jspl3_w_n614_1(.douta(w_n614_1[0]),.doutb(w_n614_1[1]),.doutc(w_n614_1[2]),.din(w_n614_0[0]));
	jspl jspl_w_n614_2(.douta(w_dff_A_HJLLE2YR5_0),.doutb(w_n614_2[1]),.din(w_n614_0[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl jspl_w_n618_1(.douta(w_n618_1[0]),.doutb(w_n618_1[1]),.din(w_n618_0[0]));
	jspl3 jspl3_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.doutc(w_n621_0[2]),.din(n621));
	jspl3 jspl3_w_n621_1(.douta(w_dff_A_g2qvW19T6_0),.doutb(w_n621_1[1]),.doutc(w_n621_1[2]),.din(w_n621_0[0]));
	jspl jspl_w_n621_2(.douta(w_dff_A_uK0Xd9Vt0_0),.doutb(w_n621_2[1]),.din(w_n621_0[1]));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_n622_0[2]),.din(n622));
	jspl jspl_w_n622_1(.douta(w_n622_1[0]),.doutb(w_n622_1[1]),.din(w_n622_0[0]));
	jspl jspl_w_n623_0(.douta(w_dff_A_Gxmw2GQZ2_0),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.doutc(w_n624_0[2]),.din(n624));
	jspl3 jspl3_w_n624_1(.douta(w_n624_1[0]),.doutb(w_n624_1[1]),.doutc(w_n624_1[2]),.din(w_n624_0[0]));
	jspl3 jspl3_w_n625_0(.douta(w_dff_A_QCo5rrFG2_0),.doutb(w_n625_0[1]),.doutc(w_dff_A_41iniY6v3_2),.din(n625));
	jspl3 jspl3_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.doutc(w_n628_0[2]),.din(n628));
	jspl3 jspl3_w_n629_0(.douta(w_n629_0[0]),.doutb(w_dff_A_a62VI9RO2_1),.doutc(w_n629_0[2]),.din(n629));
	jspl jspl_w_n631_0(.douta(w_dff_A_yhM1GGPX8_0),.doutb(w_n631_0[1]),.din(n631));
	jspl3 jspl3_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.doutc(w_n633_0[2]),.din(n633));
	jspl jspl_w_n633_1(.douta(w_n633_1[0]),.doutb(w_n633_1[1]),.din(w_n633_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_dff_A_6l12njUS4_2),.din(n636));
	jspl jspl_w_n636_1(.douta(w_n636_1[0]),.doutb(w_dff_A_VzvL9tk17_1),.din(w_n636_0[0]));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.doutc(w_n645_0[2]),.din(n645));
	jspl3 jspl3_w_n646_0(.douta(w_n646_0[0]),.doutb(w_n646_0[1]),.doutc(w_n646_0[2]),.din(n646));
	jspl3 jspl3_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.doutc(w_n649_0[2]),.din(n649));
	jspl jspl_w_n649_1(.douta(w_n649_1[0]),.doutb(w_n649_1[1]),.din(w_n649_0[0]));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.doutc(w_n651_0[2]),.din(n651));
	jspl jspl_w_n651_1(.douta(w_dff_A_hirtmZVm7_0),.doutb(w_n651_1[1]),.din(w_n651_0[0]));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(w_dff_B_uaqFFGz90_2));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl jspl_w_n671_0(.douta(w_dff_A_xUU0Go5l4_0),.doutb(w_n671_0[1]),.din(n671));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.din(n679));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl3 jspl3_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.doutc(w_n681_0[2]),.din(n681));
	jspl3 jspl3_w_n681_1(.douta(w_n681_1[0]),.doutb(w_n681_1[1]),.doutc(w_n681_1[2]),.din(w_n681_0[0]));
	jspl jspl_w_n681_2(.douta(w_n681_2[0]),.doutb(w_n681_2[1]),.din(w_n681_0[1]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl3 jspl3_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.doutc(w_n687_0[2]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl3 jspl3_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.doutc(w_n691_0[2]),.din(n691));
	jspl3 jspl3_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.doutc(w_n693_0[2]),.din(n693));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.doutc(w_n696_0[2]),.din(n696));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_n700_0[1]),.din(n700));
	jspl jspl_w_n702_0(.douta(w_n702_0[0]),.doutb(w_n702_0[1]),.din(n702));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.doutc(w_n707_0[2]),.din(n707));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(w_dff_B_ukggaXHx1_2));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_dff_A_nsxbk5Go9_1),.doutc(w_dff_A_o3ibLdIi1_2),.din(n717));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl3 jspl3_w_n721_0(.douta(w_n721_0[0]),.doutb(w_dff_A_4MaBBqXA9_1),.doutc(w_n721_0[2]),.din(n721));
	jspl jspl_w_n723_0(.douta(w_dff_A_OEnd0fHr7_0),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl3 jspl3_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.doutc(w_n727_0[2]),.din(n727));
	jspl3 jspl3_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.doutc(w_n729_0[2]),.din(n729));
	jspl jspl_w_n729_1(.douta(w_n729_1[0]),.doutb(w_n729_1[1]),.din(w_n729_0[0]));
	jspl3 jspl3_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.doutc(w_n732_0[2]),.din(n732));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.din(n735));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl3 jspl3_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.doutc(w_n739_0[2]),.din(n739));
	jspl jspl_w_n739_1(.douta(w_n739_1[0]),.doutb(w_n739_1[1]),.din(w_n739_0[0]));
	jspl jspl_w_n740_0(.douta(w_n740_0[0]),.doutb(w_n740_0[1]),.din(n740));
	jspl jspl_w_n741_0(.douta(w_dff_A_mdUzwDUP4_0),.doutb(w_n741_0[1]),.din(n741));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(w_dff_B_HG903BB55_2));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_dff_A_pQVO2DnM4_2),.din(w_dff_B_5L8eXvRX9_3));
	jspl3 jspl3_w_n744_1(.douta(w_dff_A_NBhpaSKd4_0),.doutb(w_n744_1[1]),.doutc(w_n744_1[2]),.din(w_n744_0[0]));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.doutc(w_n746_0[2]),.din(n746));
	jspl3 jspl3_w_n746_1(.douta(w_n746_1[0]),.doutb(w_n746_1[1]),.doutc(w_n746_1[2]),.din(w_n746_0[0]));
	jspl3 jspl3_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.doutc(w_n747_0[2]),.din(n747));
	jspl3 jspl3_w_n747_1(.douta(w_n747_1[0]),.doutb(w_n747_1[1]),.doutc(w_n747_1[2]),.din(w_n747_0[0]));
	jspl3 jspl3_w_n747_2(.douta(w_n747_2[0]),.doutb(w_n747_2[1]),.doutc(w_n747_2[2]),.din(w_n747_0[1]));
	jspl3 jspl3_w_n747_3(.douta(w_n747_3[0]),.doutb(w_n747_3[1]),.doutc(w_n747_3[2]),.din(w_n747_0[2]));
	jspl3 jspl3_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.doutc(w_n748_0[2]),.din(n748));
	jspl3 jspl3_w_n748_1(.douta(w_n748_1[0]),.doutb(w_n748_1[1]),.doutc(w_n748_1[2]),.din(w_n748_0[0]));
	jspl3 jspl3_w_n748_2(.douta(w_n748_2[0]),.doutb(w_n748_2[1]),.doutc(w_n748_2[2]),.din(w_n748_0[1]));
	jspl3 jspl3_w_n748_3(.douta(w_n748_3[0]),.doutb(w_dff_A_jFHnAu0m2_1),.doutc(w_dff_A_hufhjLzc9_2),.din(w_n748_0[2]));
	jspl jspl_w_n748_4(.douta(w_dff_A_hLumddvH0_0),.doutb(w_n748_4[1]),.din(w_n748_1[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.doutc(w_n750_0[2]),.din(n750));
	jspl jspl_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n751_0(.douta(w_n751_0[0]),.doutb(w_n751_0[1]),.doutc(w_n751_0[2]),.din(n751));
	jspl3 jspl3_w_n751_1(.douta(w_n751_1[0]),.doutb(w_n751_1[1]),.doutc(w_n751_1[2]),.din(w_n751_0[0]));
	jspl jspl_w_n751_2(.douta(w_n751_2[0]),.doutb(w_n751_2[1]),.din(w_n751_0[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.doutc(w_n753_0[2]),.din(n753));
	jspl3 jspl3_w_n753_1(.douta(w_n753_1[0]),.doutb(w_n753_1[1]),.doutc(w_n753_1[2]),.din(w_n753_0[0]));
	jspl3 jspl3_w_n753_2(.douta(w_n753_2[0]),.doutb(w_n753_2[1]),.doutc(w_n753_2[2]),.din(w_n753_0[1]));
	jspl3 jspl3_w_n753_3(.douta(w_n753_3[0]),.doutb(w_n753_3[1]),.doutc(w_n753_3[2]),.din(w_n753_0[2]));
	jspl3 jspl3_w_n753_4(.douta(w_n753_4[0]),.doutb(w_n753_4[1]),.doutc(w_n753_4[2]),.din(w_n753_1[0]));
	jspl3 jspl3_w_n753_5(.douta(w_n753_5[0]),.doutb(w_n753_5[1]),.doutc(w_n753_5[2]),.din(w_n753_1[1]));
	jspl3 jspl3_w_n753_6(.douta(w_n753_6[0]),.doutb(w_n753_6[1]),.doutc(w_n753_6[2]),.din(w_n753_1[2]));
	jspl3 jspl3_w_n753_7(.douta(w_n753_7[0]),.doutb(w_n753_7[1]),.doutc(w_n753_7[2]),.din(w_n753_2[0]));
	jspl jspl_w_n753_8(.douta(w_n753_8[0]),.doutb(w_n753_8[1]),.din(w_n753_2[1]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.din(n761));
	jspl3 jspl3_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.doutc(w_n765_0[2]),.din(n765));
	jspl3 jspl3_w_n765_1(.douta(w_n765_1[0]),.doutb(w_n765_1[1]),.doutc(w_n765_1[2]),.din(w_n765_0[0]));
	jspl3 jspl3_w_n765_2(.douta(w_n765_2[0]),.doutb(w_n765_2[1]),.doutc(w_n765_2[2]),.din(w_n765_0[1]));
	jspl3 jspl3_w_n765_3(.douta(w_n765_3[0]),.doutb(w_n765_3[1]),.doutc(w_n765_3[2]),.din(w_n765_0[2]));
	jspl3 jspl3_w_n765_4(.douta(w_n765_4[0]),.doutb(w_n765_4[1]),.doutc(w_n765_4[2]),.din(w_n765_1[0]));
	jspl3 jspl3_w_n765_5(.douta(w_n765_5[0]),.doutb(w_n765_5[1]),.doutc(w_n765_5[2]),.din(w_n765_1[1]));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_dff_A_ylRM2eMt7_1),.din(n779));
	jspl3 jspl3_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.doutc(w_n781_0[2]),.din(n781));
	jspl3 jspl3_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.doutc(w_n783_0[2]),.din(n783));
	jspl jspl_w_n783_1(.douta(w_n783_1[0]),.doutb(w_n783_1[1]),.din(w_n783_0[0]));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_hcZWEMPy7_2));
	jspl3 jspl3_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.doutc(w_n789_0[2]),.din(n789));
	jspl3 jspl3_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.doutc(w_n791_0[2]),.din(n791));
	jspl jspl_w_n791_1(.douta(w_n791_1[0]),.doutb(w_n791_1[1]),.din(w_n791_0[0]));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl3 jspl3_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.doutc(w_n793_0[2]),.din(n793));
	jspl3 jspl3_w_n793_1(.douta(w_n793_1[0]),.doutb(w_n793_1[1]),.doutc(w_n793_1[2]),.din(w_n793_0[0]));
	jspl3 jspl3_w_n793_2(.douta(w_n793_2[0]),.doutb(w_n793_2[1]),.doutc(w_n793_2[2]),.din(w_n793_0[1]));
	jspl3 jspl3_w_n793_3(.douta(w_n793_3[0]),.doutb(w_dff_A_JeyMDLcV1_1),.doutc(w_dff_A_bGOD6Vfc2_2),.din(w_n793_0[2]));
	jspl jspl_w_n793_4(.douta(w_dff_A_rNTfHfPH9_0),.doutb(w_n793_4[1]),.din(w_n793_1[0]));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_dff_A_OTsvVIaB8_1),.doutc(w_dff_A_GB2w0Nnn0_2),.din(w_dff_B_YIZo3wIt3_3));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_dff_A_BXunqfwI6_1),.doutc(w_dff_A_o2tyTjap4_2),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_dff_A_5qNoMRjg8_2),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_n797_3[0]),.doutb(w_dff_A_flohxssd4_1),.doutc(w_dff_A_km2ZL4Gp9_2),.din(w_n797_0[2]));
	jspl jspl_w_n797_4(.douta(w_dff_A_3leGPe2H6_0),.doutb(w_n797_4[1]),.din(w_n797_1[0]));
	jspl3 jspl3_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.doutc(w_n799_0[2]),.din(n799));
	jspl3 jspl3_w_n799_1(.douta(w_n799_1[0]),.doutb(w_n799_1[1]),.doutc(w_n799_1[2]),.din(w_n799_0[0]));
	jspl3 jspl3_w_n799_2(.douta(w_n799_2[0]),.doutb(w_n799_2[1]),.doutc(w_n799_2[2]),.din(w_n799_0[1]));
	jspl3 jspl3_w_n799_3(.douta(w_n799_3[0]),.doutb(w_n799_3[1]),.doutc(w_n799_3[2]),.din(w_n799_0[2]));
	jspl jspl_w_n799_4(.douta(w_n799_4[0]),.doutb(w_n799_4[1]),.din(w_n799_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl3 jspl3_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.doutc(w_n801_1[2]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n801_2(.douta(w_n801_2[0]),.doutb(w_n801_2[1]),.doutc(w_n801_2[2]),.din(w_n801_0[1]));
	jspl3 jspl3_w_n801_3(.douta(w_n801_3[0]),.doutb(w_n801_3[1]),.doutc(w_n801_3[2]),.din(w_n801_0[2]));
	jspl jspl_w_n801_4(.douta(w_n801_4[0]),.doutb(w_n801_4[1]),.din(w_n801_1[0]));
	jspl3 jspl3_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.doutc(w_n806_0[2]),.din(n806));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(n821));
	jspl3 jspl3_w_n828_0(.douta(w_n828_0[0]),.doutb(w_dff_A_bsUiUq3R8_1),.doutc(w_dff_A_A0PVhH983_2),.din(n828));
	jspl jspl_w_n829_0(.douta(w_n829_0[0]),.doutb(w_n829_0[1]),.din(n829));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl3 jspl3_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.doutc(w_n840_0[2]),.din(n840));
	jspl3 jspl3_w_n840_1(.douta(w_n840_1[0]),.doutb(w_n840_1[1]),.doutc(w_n840_1[2]),.din(w_n840_0[0]));
	jspl3 jspl3_w_n840_2(.douta(w_n840_2[0]),.doutb(w_n840_2[1]),.doutc(w_n840_2[2]),.din(w_n840_0[1]));
	jspl3 jspl3_w_n840_3(.douta(w_n840_3[0]),.doutb(w_dff_A_2ZX1RZLv2_1),.doutc(w_dff_A_lkHYSTEn1_2),.din(w_n840_0[2]));
	jspl jspl_w_n840_4(.douta(w_dff_A_fxS3wW5c0_0),.doutb(w_n840_4[1]),.din(w_n840_1[0]));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(n842));
	jspl3 jspl3_w_n843_0(.douta(w_n843_0[0]),.doutb(w_dff_A_0idNOgO82_1),.doutc(w_dff_A_mxYrmpWq2_2),.din(w_dff_B_nbEnGORg5_3));
	jspl3 jspl3_w_n843_1(.douta(w_n843_1[0]),.doutb(w_dff_A_z7biw8aO7_1),.doutc(w_dff_A_O4GArnQ14_2),.din(w_n843_0[0]));
	jspl3 jspl3_w_n843_2(.douta(w_n843_2[0]),.doutb(w_n843_2[1]),.doutc(w_dff_A_gYn5Hg3Q0_2),.din(w_n843_0[1]));
	jspl3 jspl3_w_n843_3(.douta(w_n843_3[0]),.doutb(w_dff_A_j2B9s7A08_1),.doutc(w_dff_A_HIp2utQk6_2),.din(w_n843_0[2]));
	jspl jspl_w_n843_4(.douta(w_dff_A_f5jDzHUl3_0),.doutb(w_n843_4[1]),.din(w_n843_1[0]));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.doutc(w_n845_0[2]),.din(n845));
	jspl3 jspl3_w_n845_1(.douta(w_n845_1[0]),.doutb(w_n845_1[1]),.doutc(w_n845_1[2]),.din(w_n845_0[0]));
	jspl3 jspl3_w_n845_2(.douta(w_n845_2[0]),.doutb(w_n845_2[1]),.doutc(w_n845_2[2]),.din(w_n845_0[1]));
	jspl3 jspl3_w_n845_3(.douta(w_n845_3[0]),.doutb(w_n845_3[1]),.doutc(w_n845_3[2]),.din(w_n845_0[2]));
	jspl jspl_w_n845_4(.douta(w_n845_4[0]),.doutb(w_n845_4[1]),.din(w_n845_1[0]));
	jspl3 jspl3_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.doutc(w_n847_0[2]),.din(n847));
	jspl3 jspl3_w_n847_1(.douta(w_n847_1[0]),.doutb(w_n847_1[1]),.doutc(w_n847_1[2]),.din(w_n847_0[0]));
	jspl3 jspl3_w_n847_2(.douta(w_n847_2[0]),.doutb(w_n847_2[1]),.doutc(w_n847_2[2]),.din(w_n847_0[1]));
	jspl3 jspl3_w_n847_3(.douta(w_n847_3[0]),.doutb(w_n847_3[1]),.doutc(w_n847_3[2]),.din(w_n847_0[2]));
	jspl jspl_w_n847_4(.douta(w_n847_4[0]),.doutb(w_n847_4[1]),.din(w_n847_1[0]));
	jspl jspl_w_n853_0(.douta(w_n853_0[0]),.doutb(w_n853_0[1]),.din(n853));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(n857));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(n862));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.din(n877));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n928_0(.douta(w_n928_0[0]),.doutb(w_n928_0[1]),.din(n928));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_n930_0[2]),.din(n930));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl3 jspl3_w_n936_0(.douta(w_n936_0[0]),.doutb(w_n936_0[1]),.doutc(w_n936_0[2]),.din(n936));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(n938));
	jspl jspl_w_n941_0(.douta(w_n941_0[0]),.doutb(w_n941_0[1]),.din(n941));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_n943_0[1]),.din(n943));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(n944));
	jspl jspl_w_n946_0(.douta(w_n946_0[0]),.doutb(w_n946_0[1]),.din(n946));
	jspl3 jspl3_w_n948_0(.douta(w_n948_0[0]),.doutb(w_n948_0[1]),.doutc(w_n948_0[2]),.din(n948));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n968_0(.douta(w_n968_0[0]),.doutb(w_n968_0[1]),.din(n968));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_dff_A_bR1HbHEC2_1),.din(n971));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.din(n973));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl3 jspl3_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.doutc(w_n985_0[2]),.din(n985));
	jspl3 jspl3_w_n985_1(.douta(w_n985_1[0]),.doutb(w_n985_1[1]),.doutc(w_n985_1[2]),.din(w_n985_0[0]));
	jspl3 jspl3_w_n985_2(.douta(w_n985_2[0]),.doutb(w_n985_2[1]),.doutc(w_n985_2[2]),.din(w_n985_0[1]));
	jspl3 jspl3_w_n985_3(.douta(w_dff_A_GmbTiMEO1_0),.doutb(w_dff_A_XxnP5lNH6_1),.doutc(w_n985_3[2]),.din(w_n985_0[2]));
	jspl jspl_w_n985_4(.douta(w_dff_A_H1Eerfff1_0),.doutb(w_n985_4[1]),.din(w_n985_1[0]));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.doutc(w_n988_0[2]),.din(n988));
	jspl3 jspl3_w_n988_1(.douta(w_n988_1[0]),.doutb(w_n988_1[1]),.doutc(w_n988_1[2]),.din(w_n988_0[0]));
	jspl3 jspl3_w_n988_2(.douta(w_dff_A_cDTlSNpc6_0),.doutb(w_dff_A_FloPqlkm3_1),.doutc(w_n988_2[2]),.din(w_n988_0[1]));
	jspl3 jspl3_w_n988_3(.douta(w_dff_A_vx7I6ae47_0),.doutb(w_dff_A_WOHbjGuG2_1),.doutc(w_n988_3[2]),.din(w_n988_0[2]));
	jspl jspl_w_n988_4(.douta(w_dff_A_SOjh66Ht0_0),.doutb(w_n988_4[1]),.din(w_n988_1[0]));
	jspl3 jspl3_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.doutc(w_n990_0[2]),.din(n990));
	jspl3 jspl3_w_n990_1(.douta(w_n990_1[0]),.doutb(w_n990_1[1]),.doutc(w_n990_1[2]),.din(w_n990_0[0]));
	jspl3 jspl3_w_n990_2(.douta(w_n990_2[0]),.doutb(w_n990_2[1]),.doutc(w_n990_2[2]),.din(w_n990_0[1]));
	jspl3 jspl3_w_n990_3(.douta(w_n990_3[0]),.doutb(w_n990_3[1]),.doutc(w_n990_3[2]),.din(w_n990_0[2]));
	jspl jspl_w_n990_4(.douta(w_n990_4[0]),.doutb(w_n990_4[1]),.din(w_n990_1[0]));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl3 jspl3_w_n992_1(.douta(w_n992_1[0]),.doutb(w_n992_1[1]),.doutc(w_n992_1[2]),.din(w_n992_0[0]));
	jspl3 jspl3_w_n992_2(.douta(w_n992_2[0]),.doutb(w_n992_2[1]),.doutc(w_n992_2[2]),.din(w_n992_0[1]));
	jspl3 jspl3_w_n992_3(.douta(w_n992_3[0]),.doutb(w_n992_3[1]),.doutc(w_n992_3[2]),.din(w_n992_0[2]));
	jspl jspl_w_n992_4(.douta(w_n992_4[0]),.doutb(w_n992_4[1]),.din(w_n992_1[0]));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.doutc(w_n999_0[2]),.din(n999));
	jspl3 jspl3_w_n999_1(.douta(w_n999_1[0]),.doutb(w_n999_1[1]),.doutc(w_n999_1[2]),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_n999_2[0]),.doutb(w_n999_2[1]),.doutc(w_n999_2[2]),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_dff_A_J3xX0R6e9_0),.doutb(w_dff_A_63C5xwlS3_1),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl jspl_w_n999_4(.douta(w_dff_A_pgXuwcnj2_0),.doutb(w_n999_4[1]),.din(w_n999_1[0]));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.doutc(w_n1002_0[2]),.din(n1002));
	jspl3 jspl3_w_n1002_1(.douta(w_n1002_1[0]),.doutb(w_n1002_1[1]),.doutc(w_n1002_1[2]),.din(w_n1002_0[0]));
	jspl3 jspl3_w_n1002_2(.douta(w_dff_A_qKPaqswS4_0),.doutb(w_dff_A_oWjaihkA6_1),.doutc(w_n1002_2[2]),.din(w_n1002_0[1]));
	jspl3 jspl3_w_n1002_3(.douta(w_dff_A_Lx5GNs0P4_0),.doutb(w_dff_A_xd58JnAC1_1),.doutc(w_n1002_3[2]),.din(w_n1002_0[2]));
	jspl jspl_w_n1002_4(.douta(w_dff_A_2nH0GZxE3_0),.doutb(w_n1002_4[1]),.din(w_n1002_1[0]));
	jspl3 jspl3_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.doutc(w_n1004_0[2]),.din(n1004));
	jspl3 jspl3_w_n1004_1(.douta(w_n1004_1[0]),.doutb(w_n1004_1[1]),.doutc(w_n1004_1[2]),.din(w_n1004_0[0]));
	jspl3 jspl3_w_n1004_2(.douta(w_n1004_2[0]),.doutb(w_n1004_2[1]),.doutc(w_n1004_2[2]),.din(w_n1004_0[1]));
	jspl3 jspl3_w_n1004_3(.douta(w_n1004_3[0]),.doutb(w_n1004_3[1]),.doutc(w_n1004_3[2]),.din(w_n1004_0[2]));
	jspl jspl_w_n1004_4(.douta(w_n1004_4[0]),.doutb(w_n1004_4[1]),.din(w_n1004_1[0]));
	jspl3 jspl3_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.doutc(w_n1006_0[2]),.din(n1006));
	jspl3 jspl3_w_n1006_1(.douta(w_n1006_1[0]),.doutb(w_n1006_1[1]),.doutc(w_n1006_1[2]),.din(w_n1006_0[0]));
	jspl3 jspl3_w_n1006_2(.douta(w_n1006_2[0]),.doutb(w_n1006_2[1]),.doutc(w_n1006_2[2]),.din(w_n1006_0[1]));
	jspl3 jspl3_w_n1006_3(.douta(w_n1006_3[0]),.doutb(w_n1006_3[1]),.doutc(w_n1006_3[2]),.din(w_n1006_0[2]));
	jspl jspl_w_n1006_4(.douta(w_n1006_4[0]),.doutb(w_n1006_4[1]),.din(w_n1006_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl jspl_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl jspl_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.doutc(w_n1023_0[2]),.din(n1023));
	jspl jspl_w_n1023_1(.douta(w_n1023_1[0]),.doutb(w_n1023_1[1]),.din(w_n1023_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.doutc(w_n1039_0[2]),.din(n1039));
	jspl jspl_w_n1039_1(.douta(w_n1039_1[0]),.doutb(w_n1039_1[1]),.din(w_n1039_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl jspl_w_n1142_0(.douta(w_n1142_0[0]),.doutb(w_n1142_0[1]),.din(n1142));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(n1151));
	jspl3 jspl3_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.doutc(w_n1163_0[2]),.din(n1163));
	jspl3 jspl3_w_n1163_1(.douta(w_n1163_1[0]),.doutb(w_n1163_1[1]),.doutc(w_n1163_1[2]),.din(w_n1163_0[0]));
	jspl3 jspl3_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.doutc(w_n1197_0[2]),.din(n1197));
	jspl3 jspl3_w_n1197_1(.douta(w_n1197_1[0]),.doutb(w_n1197_1[1]),.doutc(w_n1197_1[2]),.din(w_n1197_0[0]));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.doutc(w_n1235_0[2]),.din(n1235));
	jspl jspl_w_n1235_1(.douta(w_n1235_1[0]),.doutb(w_n1235_1[1]),.din(w_n1235_0[0]));
	jspl3 jspl3_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.doutc(w_n1242_0[2]),.din(n1242));
	jspl jspl_w_n1242_1(.douta(w_n1242_1[0]),.doutb(w_n1242_1[1]),.din(w_n1242_0[0]));
	jspl3 jspl3_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.doutc(w_n1244_0[2]),.din(n1244));
	jspl jspl_w_n1244_1(.douta(w_n1244_1[0]),.doutb(w_n1244_1[1]),.din(w_n1244_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl jspl_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.doutc(w_n1253_0[2]),.din(n1253));
	jspl jspl_w_n1253_1(.douta(w_n1253_1[0]),.doutb(w_n1253_1[1]),.din(w_n1253_0[0]));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.din(n1383));
	jspl jspl_w_n1391_0(.douta(w_n1391_0[0]),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(n1399));
	jspl jspl_w_n1409_0(.douta(w_dff_A_sXYZBzkT3_0),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(n1410));
	jspl jspl_w_n1411_0(.douta(w_dff_A_w4ia18uG3_0),.doutb(w_n1411_0[1]),.din(n1411));
	jspl jspl_w_n1421_0(.douta(w_dff_A_x8XgfZtr4_0),.doutb(w_n1421_0[1]),.din(n1421));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_dff_A_e0btWtwj6_1),.din(n1438));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_dff_A_5N9tgYEO1_1),.din(n1447));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(n1494));
	jspl jspl_w_n1533_0(.douta(w_n1533_0[0]),.doutb(w_n1533_0[1]),.din(n1533));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(n1553));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_n1568_0[1]),.din(n1568));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(n1597));
	jspl3 jspl3_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.doutc(w_n1601_0[2]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.din(w_dff_B_eJRdOaJC4_2));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(n1631));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(n1634));
	jdff dff_B_RzBELWjC6_1(.din(G136),.dout(w_dff_B_RzBELWjC6_1),.clk(gclk));
	jdff dff_B_JWqUGSMZ8_0(.din(G2824),.dout(w_dff_B_JWqUGSMZ8_0),.clk(gclk));
	jdff dff_B_ptZ81eDE6_1(.din(n320),.dout(w_dff_B_ptZ81eDE6_1),.clk(gclk));
	jdff dff_B_OAjlNXEo5_1(.din(n327),.dout(w_dff_B_OAjlNXEo5_1),.clk(gclk));
	jdff dff_B_FWUboPEb9_2(.din(n333),.dout(w_dff_B_FWUboPEb9_2),.clk(gclk));
	jdff dff_B_8DrVy7Dt6_1(.din(n338),.dout(w_dff_B_8DrVy7Dt6_1),.clk(gclk));
	jdff dff_B_bHJaaGt51_1(.din(n340),.dout(w_dff_B_bHJaaGt51_1),.clk(gclk));
	jdff dff_B_qX6aa1gp2_0(.din(n341),.dout(w_dff_B_qX6aa1gp2_0),.clk(gclk));
	jdff dff_B_3tVcDugs0_1(.din(n345),.dout(w_dff_B_3tVcDugs0_1),.clk(gclk));
	jdff dff_B_HADBglPu0_0(.din(n346),.dout(w_dff_B_HADBglPu0_0),.clk(gclk));
	jdff dff_A_9C0pgMBL7_0(.dout(w_G141_2[0]),.din(w_dff_A_9C0pgMBL7_0),.clk(gclk));
	jdff dff_A_C3bV5UDH8_0(.dout(w_dff_A_9C0pgMBL7_0),.din(w_dff_A_C3bV5UDH8_0),.clk(gclk));
	jdff dff_A_kXzyRFoB3_0(.dout(w_dff_A_C3bV5UDH8_0),.din(w_dff_A_kXzyRFoB3_0),.clk(gclk));
	jdff dff_A_Q4mVXVSm9_0(.dout(w_dff_A_kXzyRFoB3_0),.din(w_dff_A_Q4mVXVSm9_0),.clk(gclk));
	jdff dff_A_ZObNW4Ey2_1(.dout(w_G141_2[1]),.din(w_dff_A_ZObNW4Ey2_1),.clk(gclk));
	jdff dff_A_B86FrkrD4_1(.dout(w_dff_A_ZObNW4Ey2_1),.din(w_dff_A_B86FrkrD4_1),.clk(gclk));
	jdff dff_A_COhjQtNa9_1(.dout(w_dff_A_B86FrkrD4_1),.din(w_dff_A_COhjQtNa9_1),.clk(gclk));
	jdff dff_A_IVtEBFxm4_1(.dout(w_dff_A_COhjQtNa9_1),.din(w_dff_A_IVtEBFxm4_1),.clk(gclk));
	jdff dff_B_vFmQ5TlV0_1(.din(n350),.dout(w_dff_B_vFmQ5TlV0_1),.clk(gclk));
	jdff dff_B_YDEUWMNi4_0(.din(n351),.dout(w_dff_B_YDEUWMNi4_0),.clk(gclk));
	jdff dff_B_f2fpSkCN8_1(.din(n355),.dout(w_dff_B_f2fpSkCN8_1),.clk(gclk));
	jdff dff_B_wmy6YsLa3_0(.din(n356),.dout(w_dff_B_wmy6YsLa3_0),.clk(gclk));
	jdff dff_A_ZxugpCx67_1(.dout(w_G141_1[1]),.din(w_dff_A_ZxugpCx67_1),.clk(gclk));
	jdff dff_A_DrQHCVWM3_1(.dout(w_dff_A_ZxugpCx67_1),.din(w_dff_A_DrQHCVWM3_1),.clk(gclk));
	jdff dff_A_PvaVoCTq9_1(.dout(w_dff_A_DrQHCVWM3_1),.din(w_dff_A_PvaVoCTq9_1),.clk(gclk));
	jdff dff_A_TiUCt4UZ9_1(.dout(w_dff_A_PvaVoCTq9_1),.din(w_dff_A_TiUCt4UZ9_1),.clk(gclk));
	jdff dff_A_gN7N4X8q9_2(.dout(w_G141_1[2]),.din(w_dff_A_gN7N4X8q9_2),.clk(gclk));
	jdff dff_A_mg8gFpYf6_2(.dout(w_dff_A_gN7N4X8q9_2),.din(w_dff_A_mg8gFpYf6_2),.clk(gclk));
	jdff dff_A_WTy7MJiF3_2(.dout(w_dff_A_mg8gFpYf6_2),.din(w_dff_A_WTy7MJiF3_2),.clk(gclk));
	jdff dff_A_c4hnKAkf8_2(.dout(w_dff_A_WTy7MJiF3_2),.din(w_dff_A_c4hnKAkf8_2),.clk(gclk));
	jdff dff_B_iKaawZhP2_1(.din(n384),.dout(w_dff_B_iKaawZhP2_1),.clk(gclk));
	jdff dff_B_kgDrTsHG1_1(.din(w_dff_B_iKaawZhP2_1),.dout(w_dff_B_kgDrTsHG1_1),.clk(gclk));
	jdff dff_B_k2BhBUC50_1(.din(n483),.dout(w_dff_B_k2BhBUC50_1),.clk(gclk));
	jdff dff_B_uaqFFGz90_2(.din(n652),.dout(w_dff_B_uaqFFGz90_2),.clk(gclk));
	jdff dff_B_fWpcCLRF3_2(.din(n709),.dout(w_dff_B_fWpcCLRF3_2),.clk(gclk));
	jdff dff_B_eHWaVUCs6_2(.din(w_dff_B_fWpcCLRF3_2),.dout(w_dff_B_eHWaVUCs6_2),.clk(gclk));
	jdff dff_B_ukggaXHx1_2(.din(w_dff_B_eHWaVUCs6_2),.dout(w_dff_B_ukggaXHx1_2),.clk(gclk));
	jdff dff_B_QishoWLg1_2(.din(n742),.dout(w_dff_B_QishoWLg1_2),.clk(gclk));
	jdff dff_B_mOqa1OGg6_2(.din(w_dff_B_QishoWLg1_2),.dout(w_dff_B_mOqa1OGg6_2),.clk(gclk));
	jdff dff_B_ZSLKpmE55_2(.din(w_dff_B_mOqa1OGg6_2),.dout(w_dff_B_ZSLKpmE55_2),.clk(gclk));
	jdff dff_B_R69B89aU0_2(.din(w_dff_B_ZSLKpmE55_2),.dout(w_dff_B_R69B89aU0_2),.clk(gclk));
	jdff dff_B_HG903BB55_2(.din(w_dff_B_R69B89aU0_2),.dout(w_dff_B_HG903BB55_2),.clk(gclk));
	jdff dff_A_OW39dcyk1_0(.dout(w_n651_1[0]),.din(w_dff_A_OW39dcyk1_0),.clk(gclk));
	jdff dff_A_GtpwQz4h7_0(.dout(w_dff_A_OW39dcyk1_0),.din(w_dff_A_GtpwQz4h7_0),.clk(gclk));
	jdff dff_A_ZXz8anXH0_0(.dout(w_dff_A_GtpwQz4h7_0),.din(w_dff_A_ZXz8anXH0_0),.clk(gclk));
	jdff dff_A_xsnU0FGa5_0(.dout(w_dff_A_ZXz8anXH0_0),.din(w_dff_A_xsnU0FGa5_0),.clk(gclk));
	jdff dff_A_yUFgaqvw7_0(.dout(w_dff_A_xsnU0FGa5_0),.din(w_dff_A_yUFgaqvw7_0),.clk(gclk));
	jdff dff_A_hirtmZVm7_0(.dout(w_dff_A_yUFgaqvw7_0),.din(w_dff_A_hirtmZVm7_0),.clk(gclk));
	jdff dff_B_mKOBTZB24_0(.din(n803),.dout(w_dff_B_mKOBTZB24_0),.clk(gclk));
	jdff dff_B_2lQ0J8dv0_0(.din(w_dff_B_mKOBTZB24_0),.dout(w_dff_B_2lQ0J8dv0_0),.clk(gclk));
	jdff dff_B_uiqNtDor1_0(.din(w_dff_B_2lQ0J8dv0_0),.dout(w_dff_B_uiqNtDor1_0),.clk(gclk));
	jdff dff_B_ic366AMP9_0(.din(w_dff_B_uiqNtDor1_0),.dout(w_dff_B_ic366AMP9_0),.clk(gclk));
	jdff dff_B_o5YSYmXM7_0(.din(w_dff_B_ic366AMP9_0),.dout(w_dff_B_o5YSYmXM7_0),.clk(gclk));
	jdff dff_B_YP1E7uEv8_0(.din(n849),.dout(w_dff_B_YP1E7uEv8_0),.clk(gclk));
	jdff dff_B_0LWkBtLA4_0(.din(w_dff_B_YP1E7uEv8_0),.dout(w_dff_B_0LWkBtLA4_0),.clk(gclk));
	jdff dff_B_RWa4FnYE8_0(.din(w_dff_B_0LWkBtLA4_0),.dout(w_dff_B_RWa4FnYE8_0),.clk(gclk));
	jdff dff_B_4EWw5jV12_0(.din(w_dff_B_RWa4FnYE8_0),.dout(w_dff_B_4EWw5jV12_0),.clk(gclk));
	jdff dff_B_BaO8iXGJ0_0(.din(w_dff_B_4EWw5jV12_0),.dout(w_dff_B_BaO8iXGJ0_0),.clk(gclk));
	jdff dff_B_VpSRf2wQ8_0(.din(n980),.dout(w_dff_B_VpSRf2wQ8_0),.clk(gclk));
	jdff dff_B_dXMUhcYZ7_0(.din(w_dff_B_VpSRf2wQ8_0),.dout(w_dff_B_dXMUhcYZ7_0),.clk(gclk));
	jdff dff_B_YzYh7TTY3_0(.din(n979),.dout(w_dff_B_YzYh7TTY3_0),.clk(gclk));
	jdff dff_B_k9iDq4bf2_0(.din(n978),.dout(w_dff_B_k9iDq4bf2_0),.clk(gclk));
	jdff dff_B_umkbvgcF8_0(.din(n977),.dout(w_dff_B_umkbvgcF8_0),.clk(gclk));
	jdff dff_B_gMOCBXgU4_0(.din(n976),.dout(w_dff_B_gMOCBXgU4_0),.clk(gclk));
	jdff dff_B_7rs07MRI9_0(.din(n994),.dout(w_dff_B_7rs07MRI9_0),.clk(gclk));
	jdff dff_B_KdGRFTnr7_0(.din(w_dff_B_7rs07MRI9_0),.dout(w_dff_B_KdGRFTnr7_0),.clk(gclk));
	jdff dff_B_x0AhPXlO8_0(.din(w_dff_B_KdGRFTnr7_0),.dout(w_dff_B_x0AhPXlO8_0),.clk(gclk));
	jdff dff_B_9prtjbAa3_0(.din(w_dff_B_x0AhPXlO8_0),.dout(w_dff_B_9prtjbAa3_0),.clk(gclk));
	jdff dff_B_HzcAlp7l2_0(.din(w_dff_B_9prtjbAa3_0),.dout(w_dff_B_HzcAlp7l2_0),.clk(gclk));
	jdff dff_B_gMxSx6Ho5_0(.din(n1008),.dout(w_dff_B_gMxSx6Ho5_0),.clk(gclk));
	jdff dff_B_ca9zya6x5_0(.din(w_dff_B_gMxSx6Ho5_0),.dout(w_dff_B_ca9zya6x5_0),.clk(gclk));
	jdff dff_B_gpB42W571_0(.din(w_dff_B_ca9zya6x5_0),.dout(w_dff_B_gpB42W571_0),.clk(gclk));
	jdff dff_B_H2TjMq3a0_0(.din(w_dff_B_gpB42W571_0),.dout(w_dff_B_H2TjMq3a0_0),.clk(gclk));
	jdff dff_B_AMDlZ77B5_0(.din(w_dff_B_H2TjMq3a0_0),.dout(w_dff_B_AMDlZ77B5_0),.clk(gclk));
	jdff dff_B_0wHZ84El8_1(.din(n749),.dout(w_dff_B_0wHZ84El8_1),.clk(gclk));
	jdff dff_B_3UTEDciD9_0(.din(n1019),.dout(w_dff_B_3UTEDciD9_0),.clk(gclk));
	jdff dff_B_0wMPxvlQ4_0(.din(n1018),.dout(w_dff_B_0wMPxvlQ4_0),.clk(gclk));
	jdff dff_B_II81o4S52_0(.din(w_dff_B_0wMPxvlQ4_0),.dout(w_dff_B_II81o4S52_0),.clk(gclk));
	jdff dff_B_nptmKkUZ1_0(.din(w_dff_B_II81o4S52_0),.dout(w_dff_B_nptmKkUZ1_0),.clk(gclk));
	jdff dff_B_2hotGX0c9_0(.din(w_dff_B_nptmKkUZ1_0),.dout(w_dff_B_2hotGX0c9_0),.clk(gclk));
	jdff dff_B_nDnBkqnF8_0(.din(w_dff_B_2hotGX0c9_0),.dout(w_dff_B_nDnBkqnF8_0),.clk(gclk));
	jdff dff_B_4pV60Ame4_0(.din(w_dff_B_nDnBkqnF8_0),.dout(w_dff_B_4pV60Ame4_0),.clk(gclk));
	jdff dff_B_IDIr9lHx6_0(.din(w_dff_B_4pV60Ame4_0),.dout(w_dff_B_IDIr9lHx6_0),.clk(gclk));
	jdff dff_B_GUp9kupK6_0(.din(w_dff_B_IDIr9lHx6_0),.dout(w_dff_B_GUp9kupK6_0),.clk(gclk));
	jdff dff_B_o8EYHMOg5_0(.din(w_dff_B_GUp9kupK6_0),.dout(w_dff_B_o8EYHMOg5_0),.clk(gclk));
	jdff dff_B_7HyvhXRI1_0(.din(w_dff_B_o8EYHMOg5_0),.dout(w_dff_B_7HyvhXRI1_0),.clk(gclk));
	jdff dff_B_8rz9pWQc7_0(.din(w_dff_B_7HyvhXRI1_0),.dout(w_dff_B_8rz9pWQc7_0),.clk(gclk));
	jdff dff_B_Q3Wm8lkY8_0(.din(w_dff_B_8rz9pWQc7_0),.dout(w_dff_B_Q3Wm8lkY8_0),.clk(gclk));
	jdff dff_A_PB21WzYN0_0(.dout(w_n797_4[0]),.din(w_dff_A_PB21WzYN0_0),.clk(gclk));
	jdff dff_A_6OXAzj3g5_0(.dout(w_dff_A_PB21WzYN0_0),.din(w_dff_A_6OXAzj3g5_0),.clk(gclk));
	jdff dff_A_2DuL7SYO4_0(.dout(w_dff_A_6OXAzj3g5_0),.din(w_dff_A_2DuL7SYO4_0),.clk(gclk));
	jdff dff_A_gCDMYwaD2_0(.dout(w_dff_A_2DuL7SYO4_0),.din(w_dff_A_gCDMYwaD2_0),.clk(gclk));
	jdff dff_A_ueYTv5xU0_0(.dout(w_dff_A_gCDMYwaD2_0),.din(w_dff_A_ueYTv5xU0_0),.clk(gclk));
	jdff dff_A_M8ldEAB83_0(.dout(w_dff_A_ueYTv5xU0_0),.din(w_dff_A_M8ldEAB83_0),.clk(gclk));
	jdff dff_A_3leGPe2H6_0(.dout(w_dff_A_M8ldEAB83_0),.din(w_dff_A_3leGPe2H6_0),.clk(gclk));
	jdff dff_A_0aM3uvZb7_0(.dout(w_n793_4[0]),.din(w_dff_A_0aM3uvZb7_0),.clk(gclk));
	jdff dff_A_jkpXis341_0(.dout(w_dff_A_0aM3uvZb7_0),.din(w_dff_A_jkpXis341_0),.clk(gclk));
	jdff dff_A_lU0dF5Bv0_0(.dout(w_dff_A_jkpXis341_0),.din(w_dff_A_lU0dF5Bv0_0),.clk(gclk));
	jdff dff_A_mwdpgRYx4_0(.dout(w_dff_A_lU0dF5Bv0_0),.din(w_dff_A_mwdpgRYx4_0),.clk(gclk));
	jdff dff_A_ekywUrWf7_0(.dout(w_dff_A_mwdpgRYx4_0),.din(w_dff_A_ekywUrWf7_0),.clk(gclk));
	jdff dff_A_mkqb6dMC3_0(.dout(w_dff_A_ekywUrWf7_0),.din(w_dff_A_mkqb6dMC3_0),.clk(gclk));
	jdff dff_A_T2sGO75z4_0(.dout(w_dff_A_mkqb6dMC3_0),.din(w_dff_A_T2sGO75z4_0),.clk(gclk));
	jdff dff_A_rNTfHfPH9_0(.dout(w_dff_A_T2sGO75z4_0),.din(w_dff_A_rNTfHfPH9_0),.clk(gclk));
	jdff dff_B_O8lDN2Ov1_0(.din(n1028),.dout(w_dff_B_O8lDN2Ov1_0),.clk(gclk));
	jdff dff_B_fwOQSZm62_0(.din(n1027),.dout(w_dff_B_fwOQSZm62_0),.clk(gclk));
	jdff dff_B_icSoDn673_0(.din(w_dff_B_fwOQSZm62_0),.dout(w_dff_B_icSoDn673_0),.clk(gclk));
	jdff dff_B_YGzhREhr9_0(.din(w_dff_B_icSoDn673_0),.dout(w_dff_B_YGzhREhr9_0),.clk(gclk));
	jdff dff_B_4USECAa41_0(.din(w_dff_B_YGzhREhr9_0),.dout(w_dff_B_4USECAa41_0),.clk(gclk));
	jdff dff_B_Pn8onG5L1_0(.din(w_dff_B_4USECAa41_0),.dout(w_dff_B_Pn8onG5L1_0),.clk(gclk));
	jdff dff_B_PooRPk5o2_0(.din(w_dff_B_Pn8onG5L1_0),.dout(w_dff_B_PooRPk5o2_0),.clk(gclk));
	jdff dff_B_iOivrpSl1_0(.din(w_dff_B_PooRPk5o2_0),.dout(w_dff_B_iOivrpSl1_0),.clk(gclk));
	jdff dff_B_fIDJAEzU8_0(.din(w_dff_B_iOivrpSl1_0),.dout(w_dff_B_fIDJAEzU8_0),.clk(gclk));
	jdff dff_B_S4DsBMNP4_0(.din(w_dff_B_fIDJAEzU8_0),.dout(w_dff_B_S4DsBMNP4_0),.clk(gclk));
	jdff dff_B_0qEmyr9a0_0(.din(w_dff_B_S4DsBMNP4_0),.dout(w_dff_B_0qEmyr9a0_0),.clk(gclk));
	jdff dff_B_26fQGdqr6_0(.din(n1037),.dout(w_dff_B_26fQGdqr6_0),.clk(gclk));
	jdff dff_B_qyYTazVA2_0(.din(w_dff_B_26fQGdqr6_0),.dout(w_dff_B_qyYTazVA2_0),.clk(gclk));
	jdff dff_B_yWOP5syg3_0(.din(n1036),.dout(w_dff_B_yWOP5syg3_0),.clk(gclk));
	jdff dff_B_tiZsxCVD0_0(.din(w_dff_B_yWOP5syg3_0),.dout(w_dff_B_tiZsxCVD0_0),.clk(gclk));
	jdff dff_B_YIK1oPkM0_0(.din(w_dff_B_tiZsxCVD0_0),.dout(w_dff_B_YIK1oPkM0_0),.clk(gclk));
	jdff dff_B_cYoiz19V4_0(.din(w_dff_B_YIK1oPkM0_0),.dout(w_dff_B_cYoiz19V4_0),.clk(gclk));
	jdff dff_B_xZN0ED6Q6_0(.din(w_dff_B_cYoiz19V4_0),.dout(w_dff_B_xZN0ED6Q6_0),.clk(gclk));
	jdff dff_B_PC2KF1KL5_0(.din(w_dff_B_xZN0ED6Q6_0),.dout(w_dff_B_PC2KF1KL5_0),.clk(gclk));
	jdff dff_B_3VDSy90D4_0(.din(w_dff_B_PC2KF1KL5_0),.dout(w_dff_B_3VDSy90D4_0),.clk(gclk));
	jdff dff_B_7x1yOwOB6_0(.din(w_dff_B_3VDSy90D4_0),.dout(w_dff_B_7x1yOwOB6_0),.clk(gclk));
	jdff dff_B_6f2NhJRQ0_0(.din(n1046),.dout(w_dff_B_6f2NhJRQ0_0),.clk(gclk));
	jdff dff_B_DWLt45xz0_0(.din(w_dff_B_6f2NhJRQ0_0),.dout(w_dff_B_DWLt45xz0_0),.clk(gclk));
	jdff dff_B_jAtPmFYd6_0(.din(w_dff_B_DWLt45xz0_0),.dout(w_dff_B_jAtPmFYd6_0),.clk(gclk));
	jdff dff_B_2sCn4Gkj0_0(.din(n1045),.dout(w_dff_B_2sCn4Gkj0_0),.clk(gclk));
	jdff dff_B_kRNEjy8b1_0(.din(w_dff_B_2sCn4Gkj0_0),.dout(w_dff_B_kRNEjy8b1_0),.clk(gclk));
	jdff dff_B_DEOkiNkd0_0(.din(w_dff_B_kRNEjy8b1_0),.dout(w_dff_B_DEOkiNkd0_0),.clk(gclk));
	jdff dff_B_c4SzRoxO9_0(.din(w_dff_B_DEOkiNkd0_0),.dout(w_dff_B_c4SzRoxO9_0),.clk(gclk));
	jdff dff_B_eehwCpWg4_0(.din(w_dff_B_c4SzRoxO9_0),.dout(w_dff_B_eehwCpWg4_0),.clk(gclk));
	jdff dff_B_Lylrgo3b1_0(.din(w_dff_B_eehwCpWg4_0),.dout(w_dff_B_Lylrgo3b1_0),.clk(gclk));
	jdff dff_A_iXVDWhc73_1(.dout(w_n797_3[1]),.din(w_dff_A_iXVDWhc73_1),.clk(gclk));
	jdff dff_A_flohxssd4_1(.dout(w_dff_A_iXVDWhc73_1),.din(w_dff_A_flohxssd4_1),.clk(gclk));
	jdff dff_A_tAJ90iUP1_2(.dout(w_n797_3[2]),.din(w_dff_A_tAJ90iUP1_2),.clk(gclk));
	jdff dff_A_wjNf8aSE5_2(.dout(w_dff_A_tAJ90iUP1_2),.din(w_dff_A_wjNf8aSE5_2),.clk(gclk));
	jdff dff_A_IjFKvcOz3_2(.dout(w_dff_A_wjNf8aSE5_2),.din(w_dff_A_IjFKvcOz3_2),.clk(gclk));
	jdff dff_A_km2ZL4Gp9_2(.dout(w_dff_A_IjFKvcOz3_2),.din(w_dff_A_km2ZL4Gp9_2),.clk(gclk));
	jdff dff_A_JeyMDLcV1_1(.dout(w_n793_3[1]),.din(w_dff_A_JeyMDLcV1_1),.clk(gclk));
	jdff dff_A_U2G2gjC92_2(.dout(w_n793_3[2]),.din(w_dff_A_U2G2gjC92_2),.clk(gclk));
	jdff dff_A_bGOD6Vfc2_2(.dout(w_dff_A_U2G2gjC92_2),.din(w_dff_A_bGOD6Vfc2_2),.clk(gclk));
	jdff dff_B_WLJDP7aX5_0(.din(n1053),.dout(w_dff_B_WLJDP7aX5_0),.clk(gclk));
	jdff dff_B_hyVEFCOX6_0(.din(n1052),.dout(w_dff_B_hyVEFCOX6_0),.clk(gclk));
	jdff dff_B_bp8oz2Yp3_0(.din(w_dff_B_hyVEFCOX6_0),.dout(w_dff_B_bp8oz2Yp3_0),.clk(gclk));
	jdff dff_B_SV85jtcn9_0(.din(w_dff_B_bp8oz2Yp3_0),.dout(w_dff_B_SV85jtcn9_0),.clk(gclk));
	jdff dff_B_NcgEUrkH8_0(.din(w_dff_B_SV85jtcn9_0),.dout(w_dff_B_NcgEUrkH8_0),.clk(gclk));
	jdff dff_B_0FqPBkLi0_0(.din(w_dff_B_NcgEUrkH8_0),.dout(w_dff_B_0FqPBkLi0_0),.clk(gclk));
	jdff dff_B_H9MgKrMR1_0(.din(w_dff_B_0FqPBkLi0_0),.dout(w_dff_B_H9MgKrMR1_0),.clk(gclk));
	jdff dff_B_4vtpxsRP6_0(.din(w_dff_B_H9MgKrMR1_0),.dout(w_dff_B_4vtpxsRP6_0),.clk(gclk));
	jdff dff_B_n19WXVD79_0(.din(w_dff_B_4vtpxsRP6_0),.dout(w_dff_B_n19WXVD79_0),.clk(gclk));
	jdff dff_B_ML3hLjTP6_0(.din(w_dff_B_n19WXVD79_0),.dout(w_dff_B_ML3hLjTP6_0),.clk(gclk));
	jdff dff_B_DUNvPQbT4_0(.din(w_dff_B_ML3hLjTP6_0),.dout(w_dff_B_DUNvPQbT4_0),.clk(gclk));
	jdff dff_B_TmxpdT241_0(.din(w_dff_B_DUNvPQbT4_0),.dout(w_dff_B_TmxpdT241_0),.clk(gclk));
	jdff dff_B_1xC9NPUj3_0(.din(w_dff_B_TmxpdT241_0),.dout(w_dff_B_1xC9NPUj3_0),.clk(gclk));
	jdff dff_A_UFT1gAXt4_0(.dout(w_n843_4[0]),.din(w_dff_A_UFT1gAXt4_0),.clk(gclk));
	jdff dff_A_SLDxeEnB5_0(.dout(w_dff_A_UFT1gAXt4_0),.din(w_dff_A_SLDxeEnB5_0),.clk(gclk));
	jdff dff_A_nvwh3Ayz7_0(.dout(w_dff_A_SLDxeEnB5_0),.din(w_dff_A_nvwh3Ayz7_0),.clk(gclk));
	jdff dff_A_BlE8r4On6_0(.dout(w_dff_A_nvwh3Ayz7_0),.din(w_dff_A_BlE8r4On6_0),.clk(gclk));
	jdff dff_A_YAPHpsN59_0(.dout(w_dff_A_BlE8r4On6_0),.din(w_dff_A_YAPHpsN59_0),.clk(gclk));
	jdff dff_A_89UIB3AV2_0(.dout(w_dff_A_YAPHpsN59_0),.din(w_dff_A_89UIB3AV2_0),.clk(gclk));
	jdff dff_A_f5jDzHUl3_0(.dout(w_dff_A_89UIB3AV2_0),.din(w_dff_A_f5jDzHUl3_0),.clk(gclk));
	jdff dff_A_Dn6AKhlp1_0(.dout(w_n840_4[0]),.din(w_dff_A_Dn6AKhlp1_0),.clk(gclk));
	jdff dff_A_V2AWPLil1_0(.dout(w_dff_A_Dn6AKhlp1_0),.din(w_dff_A_V2AWPLil1_0),.clk(gclk));
	jdff dff_A_NEcVzGTV4_0(.dout(w_dff_A_V2AWPLil1_0),.din(w_dff_A_NEcVzGTV4_0),.clk(gclk));
	jdff dff_A_V9dJ05ZL2_0(.dout(w_dff_A_NEcVzGTV4_0),.din(w_dff_A_V9dJ05ZL2_0),.clk(gclk));
	jdff dff_A_5g7Q5P4u8_0(.dout(w_dff_A_V9dJ05ZL2_0),.din(w_dff_A_5g7Q5P4u8_0),.clk(gclk));
	jdff dff_A_SODyiXzN0_0(.dout(w_dff_A_5g7Q5P4u8_0),.din(w_dff_A_SODyiXzN0_0),.clk(gclk));
	jdff dff_A_JpJbzvPb0_0(.dout(w_dff_A_SODyiXzN0_0),.din(w_dff_A_JpJbzvPb0_0),.clk(gclk));
	jdff dff_A_fxS3wW5c0_0(.dout(w_dff_A_JpJbzvPb0_0),.din(w_dff_A_fxS3wW5c0_0),.clk(gclk));
	jdff dff_B_QY6h3Pf56_0(.din(n1060),.dout(w_dff_B_QY6h3Pf56_0),.clk(gclk));
	jdff dff_B_9s8bNhxA6_0(.din(n1059),.dout(w_dff_B_9s8bNhxA6_0),.clk(gclk));
	jdff dff_B_EXUBk9iq9_0(.din(w_dff_B_9s8bNhxA6_0),.dout(w_dff_B_EXUBk9iq9_0),.clk(gclk));
	jdff dff_B_bvpstB1Y4_0(.din(w_dff_B_EXUBk9iq9_0),.dout(w_dff_B_bvpstB1Y4_0),.clk(gclk));
	jdff dff_B_HME17iCn7_0(.din(w_dff_B_bvpstB1Y4_0),.dout(w_dff_B_HME17iCn7_0),.clk(gclk));
	jdff dff_B_pbUwHfwR9_0(.din(w_dff_B_HME17iCn7_0),.dout(w_dff_B_pbUwHfwR9_0),.clk(gclk));
	jdff dff_B_kmZmkbn24_0(.din(w_dff_B_pbUwHfwR9_0),.dout(w_dff_B_kmZmkbn24_0),.clk(gclk));
	jdff dff_B_rGgHRLoE1_0(.din(w_dff_B_kmZmkbn24_0),.dout(w_dff_B_rGgHRLoE1_0),.clk(gclk));
	jdff dff_B_lHVgOqDK4_0(.din(w_dff_B_rGgHRLoE1_0),.dout(w_dff_B_lHVgOqDK4_0),.clk(gclk));
	jdff dff_B_uIX37U5y7_0(.din(w_dff_B_lHVgOqDK4_0),.dout(w_dff_B_uIX37U5y7_0),.clk(gclk));
	jdff dff_B_JMXQfCuI4_0(.din(w_dff_B_uIX37U5y7_0),.dout(w_dff_B_JMXQfCuI4_0),.clk(gclk));
	jdff dff_B_COsA15oz2_0(.din(n1067),.dout(w_dff_B_COsA15oz2_0),.clk(gclk));
	jdff dff_B_1oV735lj2_0(.din(w_dff_B_COsA15oz2_0),.dout(w_dff_B_1oV735lj2_0),.clk(gclk));
	jdff dff_B_Bw4APaHX1_0(.din(n1066),.dout(w_dff_B_Bw4APaHX1_0),.clk(gclk));
	jdff dff_B_L4X6iy017_0(.din(w_dff_B_Bw4APaHX1_0),.dout(w_dff_B_L4X6iy017_0),.clk(gclk));
	jdff dff_B_jLJQThCl5_0(.din(w_dff_B_L4X6iy017_0),.dout(w_dff_B_jLJQThCl5_0),.clk(gclk));
	jdff dff_B_VkH9BJvj3_0(.din(w_dff_B_jLJQThCl5_0),.dout(w_dff_B_VkH9BJvj3_0),.clk(gclk));
	jdff dff_B_c8FW5eSL9_0(.din(w_dff_B_VkH9BJvj3_0),.dout(w_dff_B_c8FW5eSL9_0),.clk(gclk));
	jdff dff_B_o0NNZpMN0_0(.din(w_dff_B_c8FW5eSL9_0),.dout(w_dff_B_o0NNZpMN0_0),.clk(gclk));
	jdff dff_B_Ye1H5Dwo8_0(.din(w_dff_B_o0NNZpMN0_0),.dout(w_dff_B_Ye1H5Dwo8_0),.clk(gclk));
	jdff dff_B_TCuaHdYd2_0(.din(w_dff_B_Ye1H5Dwo8_0),.dout(w_dff_B_TCuaHdYd2_0),.clk(gclk));
	jdff dff_B_l7mRFPEA2_0(.din(n1074),.dout(w_dff_B_l7mRFPEA2_0),.clk(gclk));
	jdff dff_B_VtPGMql03_0(.din(w_dff_B_l7mRFPEA2_0),.dout(w_dff_B_VtPGMql03_0),.clk(gclk));
	jdff dff_B_mqzvoDyA5_0(.din(w_dff_B_VtPGMql03_0),.dout(w_dff_B_mqzvoDyA5_0),.clk(gclk));
	jdff dff_B_MhN27Q6f9_0(.din(n1073),.dout(w_dff_B_MhN27Q6f9_0),.clk(gclk));
	jdff dff_B_2W4kTnps9_0(.din(w_dff_B_MhN27Q6f9_0),.dout(w_dff_B_2W4kTnps9_0),.clk(gclk));
	jdff dff_B_2eOnCZPV5_0(.din(w_dff_B_2W4kTnps9_0),.dout(w_dff_B_2eOnCZPV5_0),.clk(gclk));
	jdff dff_B_hdNBlLk22_0(.din(w_dff_B_2eOnCZPV5_0),.dout(w_dff_B_hdNBlLk22_0),.clk(gclk));
	jdff dff_B_2HS9pGTJ6_0(.din(w_dff_B_hdNBlLk22_0),.dout(w_dff_B_2HS9pGTJ6_0),.clk(gclk));
	jdff dff_B_CotwCRay0_0(.din(w_dff_B_2HS9pGTJ6_0),.dout(w_dff_B_CotwCRay0_0),.clk(gclk));
	jdff dff_A_alt0yisF4_1(.dout(w_n843_3[1]),.din(w_dff_A_alt0yisF4_1),.clk(gclk));
	jdff dff_A_j2B9s7A08_1(.dout(w_dff_A_alt0yisF4_1),.din(w_dff_A_j2B9s7A08_1),.clk(gclk));
	jdff dff_A_imaJQpu46_2(.dout(w_n843_3[2]),.din(w_dff_A_imaJQpu46_2),.clk(gclk));
	jdff dff_A_UWynk47f2_2(.dout(w_dff_A_imaJQpu46_2),.din(w_dff_A_UWynk47f2_2),.clk(gclk));
	jdff dff_A_WuBffQWu7_2(.dout(w_dff_A_UWynk47f2_2),.din(w_dff_A_WuBffQWu7_2),.clk(gclk));
	jdff dff_A_HIp2utQk6_2(.dout(w_dff_A_WuBffQWu7_2),.din(w_dff_A_HIp2utQk6_2),.clk(gclk));
	jdff dff_A_2ZX1RZLv2_1(.dout(w_n840_3[1]),.din(w_dff_A_2ZX1RZLv2_1),.clk(gclk));
	jdff dff_A_NejeZ81z2_2(.dout(w_n840_3[2]),.din(w_dff_A_NejeZ81z2_2),.clk(gclk));
	jdff dff_A_lkHYSTEn1_2(.dout(w_dff_A_NejeZ81z2_2),.din(w_dff_A_lkHYSTEn1_2),.clk(gclk));
	jdff dff_B_5PjVobUQ4_0(.din(n1081),.dout(w_dff_B_5PjVobUQ4_0),.clk(gclk));
	jdff dff_B_I1otXkx41_0(.din(n1080),.dout(w_dff_B_I1otXkx41_0),.clk(gclk));
	jdff dff_B_bDqmygbW1_0(.din(w_dff_B_I1otXkx41_0),.dout(w_dff_B_bDqmygbW1_0),.clk(gclk));
	jdff dff_B_yJnZLiSd8_0(.din(w_dff_B_bDqmygbW1_0),.dout(w_dff_B_yJnZLiSd8_0),.clk(gclk));
	jdff dff_B_bB0Sr1Gj6_0(.din(w_dff_B_yJnZLiSd8_0),.dout(w_dff_B_bB0Sr1Gj6_0),.clk(gclk));
	jdff dff_B_QZeE7Yp02_0(.din(w_dff_B_bB0Sr1Gj6_0),.dout(w_dff_B_QZeE7Yp02_0),.clk(gclk));
	jdff dff_B_5xzEO4Rc1_0(.din(w_dff_B_QZeE7Yp02_0),.dout(w_dff_B_5xzEO4Rc1_0),.clk(gclk));
	jdff dff_B_ziWQ1k7Z5_0(.din(w_dff_B_5xzEO4Rc1_0),.dout(w_dff_B_ziWQ1k7Z5_0),.clk(gclk));
	jdff dff_B_VByOyEj53_0(.din(w_dff_B_ziWQ1k7Z5_0),.dout(w_dff_B_VByOyEj53_0),.clk(gclk));
	jdff dff_B_DziEf5Bx5_0(.din(w_dff_B_VByOyEj53_0),.dout(w_dff_B_DziEf5Bx5_0),.clk(gclk));
	jdff dff_B_Zo5WcvMW7_0(.din(w_dff_B_DziEf5Bx5_0),.dout(w_dff_B_Zo5WcvMW7_0),.clk(gclk));
	jdff dff_B_kZVqFo4l3_0(.din(w_dff_B_Zo5WcvMW7_0),.dout(w_dff_B_kZVqFo4l3_0),.clk(gclk));
	jdff dff_B_3ID8azaP2_0(.din(w_dff_B_kZVqFo4l3_0),.dout(w_dff_B_3ID8azaP2_0),.clk(gclk));
	jdff dff_A_4APADHfG0_0(.dout(w_n988_4[0]),.din(w_dff_A_4APADHfG0_0),.clk(gclk));
	jdff dff_A_jcdf759Q8_0(.dout(w_dff_A_4APADHfG0_0),.din(w_dff_A_jcdf759Q8_0),.clk(gclk));
	jdff dff_A_rKq1Rlm87_0(.dout(w_dff_A_jcdf759Q8_0),.din(w_dff_A_rKq1Rlm87_0),.clk(gclk));
	jdff dff_A_a8eUjuHY3_0(.dout(w_dff_A_rKq1Rlm87_0),.din(w_dff_A_a8eUjuHY3_0),.clk(gclk));
	jdff dff_A_0vywOJOq4_0(.dout(w_dff_A_a8eUjuHY3_0),.din(w_dff_A_0vywOJOq4_0),.clk(gclk));
	jdff dff_A_9yAP0nK09_0(.dout(w_dff_A_0vywOJOq4_0),.din(w_dff_A_9yAP0nK09_0),.clk(gclk));
	jdff dff_A_SOjh66Ht0_0(.dout(w_dff_A_9yAP0nK09_0),.din(w_dff_A_SOjh66Ht0_0),.clk(gclk));
	jdff dff_A_UpiIgfVy1_0(.dout(w_n985_4[0]),.din(w_dff_A_UpiIgfVy1_0),.clk(gclk));
	jdff dff_A_fsVXSeFl0_0(.dout(w_dff_A_UpiIgfVy1_0),.din(w_dff_A_fsVXSeFl0_0),.clk(gclk));
	jdff dff_A_cy8CQDxH4_0(.dout(w_dff_A_fsVXSeFl0_0),.din(w_dff_A_cy8CQDxH4_0),.clk(gclk));
	jdff dff_A_zzzPEC1N0_0(.dout(w_dff_A_cy8CQDxH4_0),.din(w_dff_A_zzzPEC1N0_0),.clk(gclk));
	jdff dff_A_964eO37u6_0(.dout(w_dff_A_zzzPEC1N0_0),.din(w_dff_A_964eO37u6_0),.clk(gclk));
	jdff dff_A_4kvJzyfI4_0(.dout(w_dff_A_964eO37u6_0),.din(w_dff_A_4kvJzyfI4_0),.clk(gclk));
	jdff dff_A_KlEHEaxs4_0(.dout(w_dff_A_4kvJzyfI4_0),.din(w_dff_A_KlEHEaxs4_0),.clk(gclk));
	jdff dff_A_H1Eerfff1_0(.dout(w_dff_A_KlEHEaxs4_0),.din(w_dff_A_H1Eerfff1_0),.clk(gclk));
	jdff dff_B_n8QyPZdT5_0(.din(n1089),.dout(w_dff_B_n8QyPZdT5_0),.clk(gclk));
	jdff dff_B_J89I7pNR6_0(.din(w_dff_B_n8QyPZdT5_0),.dout(w_dff_B_J89I7pNR6_0),.clk(gclk));
	jdff dff_B_AjhPezaV8_0(.din(w_dff_B_J89I7pNR6_0),.dout(w_dff_B_AjhPezaV8_0),.clk(gclk));
	jdff dff_B_hl0GFvEU1_0(.din(n1088),.dout(w_dff_B_hl0GFvEU1_0),.clk(gclk));
	jdff dff_B_59bO7vdM3_0(.din(w_dff_B_hl0GFvEU1_0),.dout(w_dff_B_59bO7vdM3_0),.clk(gclk));
	jdff dff_B_5A4vBxa52_0(.din(w_dff_B_59bO7vdM3_0),.dout(w_dff_B_5A4vBxa52_0),.clk(gclk));
	jdff dff_B_gBCqngKc3_0(.din(w_dff_B_5A4vBxa52_0),.dout(w_dff_B_gBCqngKc3_0),.clk(gclk));
	jdff dff_B_mFkarUnK7_0(.din(w_dff_B_gBCqngKc3_0),.dout(w_dff_B_mFkarUnK7_0),.clk(gclk));
	jdff dff_B_mVA8vvvh4_0(.din(w_dff_B_mFkarUnK7_0),.dout(w_dff_B_mVA8vvvh4_0),.clk(gclk));
	jdff dff_B_QUZvArLB3_0(.din(n1097),.dout(w_dff_B_QUZvArLB3_0),.clk(gclk));
	jdff dff_B_dZoSkuxT9_0(.din(w_dff_B_QUZvArLB3_0),.dout(w_dff_B_dZoSkuxT9_0),.clk(gclk));
	jdff dff_B_qiUae91M4_0(.din(n1096),.dout(w_dff_B_qiUae91M4_0),.clk(gclk));
	jdff dff_B_mUnvMIsE0_0(.din(w_dff_B_qiUae91M4_0),.dout(w_dff_B_mUnvMIsE0_0),.clk(gclk));
	jdff dff_B_e6Alg1Mr6_0(.din(w_dff_B_mUnvMIsE0_0),.dout(w_dff_B_e6Alg1Mr6_0),.clk(gclk));
	jdff dff_B_GoOfclq14_0(.din(w_dff_B_e6Alg1Mr6_0),.dout(w_dff_B_GoOfclq14_0),.clk(gclk));
	jdff dff_B_w8BDqJrV8_0(.din(w_dff_B_GoOfclq14_0),.dout(w_dff_B_w8BDqJrV8_0),.clk(gclk));
	jdff dff_B_hmhDHuWd3_0(.din(w_dff_B_w8BDqJrV8_0),.dout(w_dff_B_hmhDHuWd3_0),.clk(gclk));
	jdff dff_B_oCB45nCt6_0(.din(w_dff_B_hmhDHuWd3_0),.dout(w_dff_B_oCB45nCt6_0),.clk(gclk));
	jdff dff_B_Wb3Mxokv3_0(.din(w_dff_B_oCB45nCt6_0),.dout(w_dff_B_Wb3Mxokv3_0),.clk(gclk));
	jdff dff_A_OlofKs7A9_0(.dout(w_G137_8[0]),.din(w_dff_A_OlofKs7A9_0),.clk(gclk));
	jdff dff_A_bREHY6Oa2_2(.dout(w_G137_8[2]),.din(w_dff_A_bREHY6Oa2_2),.clk(gclk));
	jdff dff_A_eOWBWetz2_2(.dout(w_dff_A_bREHY6Oa2_2),.din(w_dff_A_eOWBWetz2_2),.clk(gclk));
	jdff dff_A_jpqL0GFx2_2(.dout(w_dff_A_eOWBWetz2_2),.din(w_dff_A_jpqL0GFx2_2),.clk(gclk));
	jdff dff_A_WB8BAewC6_2(.dout(w_dff_A_jpqL0GFx2_2),.din(w_dff_A_WB8BAewC6_2),.clk(gclk));
	jdff dff_B_8LNnabtE7_0(.din(n1105),.dout(w_dff_B_8LNnabtE7_0),.clk(gclk));
	jdff dff_B_6w2Kod5f0_0(.din(n1104),.dout(w_dff_B_6w2Kod5f0_0),.clk(gclk));
	jdff dff_B_hmWfcwRY6_0(.din(w_dff_B_6w2Kod5f0_0),.dout(w_dff_B_hmWfcwRY6_0),.clk(gclk));
	jdff dff_B_rr7bKtVM8_0(.din(w_dff_B_hmWfcwRY6_0),.dout(w_dff_B_rr7bKtVM8_0),.clk(gclk));
	jdff dff_B_WuTUTdSS1_0(.din(w_dff_B_rr7bKtVM8_0),.dout(w_dff_B_WuTUTdSS1_0),.clk(gclk));
	jdff dff_B_6HsbXZa65_0(.din(w_dff_B_WuTUTdSS1_0),.dout(w_dff_B_6HsbXZa65_0),.clk(gclk));
	jdff dff_B_i1eWqLSa7_0(.din(w_dff_B_6HsbXZa65_0),.dout(w_dff_B_i1eWqLSa7_0),.clk(gclk));
	jdff dff_B_G396cFwj5_0(.din(w_dff_B_i1eWqLSa7_0),.dout(w_dff_B_G396cFwj5_0),.clk(gclk));
	jdff dff_B_0EXkct223_0(.din(w_dff_B_G396cFwj5_0),.dout(w_dff_B_0EXkct223_0),.clk(gclk));
	jdff dff_B_laPSel7d8_0(.din(w_dff_B_0EXkct223_0),.dout(w_dff_B_laPSel7d8_0),.clk(gclk));
	jdff dff_B_3mQ230dl9_0(.din(w_dff_B_laPSel7d8_0),.dout(w_dff_B_3mQ230dl9_0),.clk(gclk));
	jdff dff_A_uDFr2mIy1_0(.dout(w_n988_3[0]),.din(w_dff_A_uDFr2mIy1_0),.clk(gclk));
	jdff dff_A_AYsweUT61_0(.dout(w_dff_A_uDFr2mIy1_0),.din(w_dff_A_AYsweUT61_0),.clk(gclk));
	jdff dff_A_gVcqTXIN4_0(.dout(w_dff_A_AYsweUT61_0),.din(w_dff_A_gVcqTXIN4_0),.clk(gclk));
	jdff dff_A_vx7I6ae47_0(.dout(w_dff_A_gVcqTXIN4_0),.din(w_dff_A_vx7I6ae47_0),.clk(gclk));
	jdff dff_A_d1pj2AEB0_1(.dout(w_n988_3[1]),.din(w_dff_A_d1pj2AEB0_1),.clk(gclk));
	jdff dff_A_WOHbjGuG2_1(.dout(w_dff_A_d1pj2AEB0_1),.din(w_dff_A_WOHbjGuG2_1),.clk(gclk));
	jdff dff_A_qna2aV5G5_0(.dout(w_n985_3[0]),.din(w_dff_A_qna2aV5G5_0),.clk(gclk));
	jdff dff_A_GmbTiMEO1_0(.dout(w_dff_A_qna2aV5G5_0),.din(w_dff_A_GmbTiMEO1_0),.clk(gclk));
	jdff dff_A_XxnP5lNH6_1(.dout(w_n985_3[1]),.din(w_dff_A_XxnP5lNH6_1),.clk(gclk));
	jdff dff_B_wJYACATe1_0(.din(n1113),.dout(w_dff_B_wJYACATe1_0),.clk(gclk));
	jdff dff_B_7JyMLTIr8_0(.din(n1112),.dout(w_dff_B_7JyMLTIr8_0),.clk(gclk));
	jdff dff_B_eEsi5fVW9_0(.din(w_dff_B_7JyMLTIr8_0),.dout(w_dff_B_eEsi5fVW9_0),.clk(gclk));
	jdff dff_B_It73lj5j5_0(.din(w_dff_B_eEsi5fVW9_0),.dout(w_dff_B_It73lj5j5_0),.clk(gclk));
	jdff dff_B_yIlIV1J45_0(.din(w_dff_B_It73lj5j5_0),.dout(w_dff_B_yIlIV1J45_0),.clk(gclk));
	jdff dff_B_plmtYHbb9_0(.din(w_dff_B_yIlIV1J45_0),.dout(w_dff_B_plmtYHbb9_0),.clk(gclk));
	jdff dff_B_l5u8Te2Z8_0(.din(w_dff_B_plmtYHbb9_0),.dout(w_dff_B_l5u8Te2Z8_0),.clk(gclk));
	jdff dff_B_8UNPt5Sv4_0(.din(w_dff_B_l5u8Te2Z8_0),.dout(w_dff_B_8UNPt5Sv4_0),.clk(gclk));
	jdff dff_B_oozMzcuF2_0(.din(w_dff_B_8UNPt5Sv4_0),.dout(w_dff_B_oozMzcuF2_0),.clk(gclk));
	jdff dff_B_6lvN3kSY0_0(.din(w_dff_B_oozMzcuF2_0),.dout(w_dff_B_6lvN3kSY0_0),.clk(gclk));
	jdff dff_B_eNv3ff9E1_0(.din(w_dff_B_6lvN3kSY0_0),.dout(w_dff_B_eNv3ff9E1_0),.clk(gclk));
	jdff dff_B_AVJI1IGX1_0(.din(w_dff_B_eNv3ff9E1_0),.dout(w_dff_B_AVJI1IGX1_0),.clk(gclk));
	jdff dff_B_YhCP3RJR5_0(.din(w_dff_B_AVJI1IGX1_0),.dout(w_dff_B_YhCP3RJR5_0),.clk(gclk));
	jdff dff_A_qID4WNNU8_0(.dout(w_n1002_4[0]),.din(w_dff_A_qID4WNNU8_0),.clk(gclk));
	jdff dff_A_2EyN7qET1_0(.dout(w_dff_A_qID4WNNU8_0),.din(w_dff_A_2EyN7qET1_0),.clk(gclk));
	jdff dff_A_7pCpBBN39_0(.dout(w_dff_A_2EyN7qET1_0),.din(w_dff_A_7pCpBBN39_0),.clk(gclk));
	jdff dff_A_frxi9byD9_0(.dout(w_dff_A_7pCpBBN39_0),.din(w_dff_A_frxi9byD9_0),.clk(gclk));
	jdff dff_A_PIR7mxAp2_0(.dout(w_dff_A_frxi9byD9_0),.din(w_dff_A_PIR7mxAp2_0),.clk(gclk));
	jdff dff_A_Hz0GPvP20_0(.dout(w_dff_A_PIR7mxAp2_0),.din(w_dff_A_Hz0GPvP20_0),.clk(gclk));
	jdff dff_A_2nH0GZxE3_0(.dout(w_dff_A_Hz0GPvP20_0),.din(w_dff_A_2nH0GZxE3_0),.clk(gclk));
	jdff dff_B_dznslKDQ1_0(.din(n814),.dout(w_dff_B_dznslKDQ1_0),.clk(gclk));
	jdff dff_B_bJrgIGLC4_0(.din(w_dff_B_dznslKDQ1_0),.dout(w_dff_B_bJrgIGLC4_0),.clk(gclk));
	jdff dff_B_CDdEo12k0_0(.din(w_dff_B_bJrgIGLC4_0),.dout(w_dff_B_CDdEo12k0_0),.clk(gclk));
	jdff dff_B_tPZA7zsE2_0(.din(w_dff_B_CDdEo12k0_0),.dout(w_dff_B_tPZA7zsE2_0),.clk(gclk));
	jdff dff_B_xwxKc0KW7_0(.din(w_dff_B_tPZA7zsE2_0),.dout(w_dff_B_xwxKc0KW7_0),.clk(gclk));
	jdff dff_B_hhbfhIuz9_0(.din(w_dff_B_xwxKc0KW7_0),.dout(w_dff_B_hhbfhIuz9_0),.clk(gclk));
	jdff dff_A_6kLcD7zL4_0(.dout(w_n999_4[0]),.din(w_dff_A_6kLcD7zL4_0),.clk(gclk));
	jdff dff_A_fyRQIDpf3_0(.dout(w_dff_A_6kLcD7zL4_0),.din(w_dff_A_fyRQIDpf3_0),.clk(gclk));
	jdff dff_A_M7r3Zzt85_0(.dout(w_dff_A_fyRQIDpf3_0),.din(w_dff_A_M7r3Zzt85_0),.clk(gclk));
	jdff dff_A_EvWzUAqm3_0(.dout(w_dff_A_M7r3Zzt85_0),.din(w_dff_A_EvWzUAqm3_0),.clk(gclk));
	jdff dff_A_iWtviGMz6_0(.dout(w_dff_A_EvWzUAqm3_0),.din(w_dff_A_iWtviGMz6_0),.clk(gclk));
	jdff dff_A_N4bFkALy3_0(.dout(w_dff_A_iWtviGMz6_0),.din(w_dff_A_N4bFkALy3_0),.clk(gclk));
	jdff dff_A_51Bj5kf34_0(.dout(w_dff_A_N4bFkALy3_0),.din(w_dff_A_51Bj5kf34_0),.clk(gclk));
	jdff dff_A_pgXuwcnj2_0(.dout(w_dff_A_51Bj5kf34_0),.din(w_dff_A_pgXuwcnj2_0),.clk(gclk));
	jdff dff_B_7VAQKTC95_0(.din(n1121),.dout(w_dff_B_7VAQKTC95_0),.clk(gclk));
	jdff dff_B_NdJPE4XP6_0(.din(w_dff_B_7VAQKTC95_0),.dout(w_dff_B_NdJPE4XP6_0),.clk(gclk));
	jdff dff_B_NqLTbuqA7_0(.din(w_dff_B_NdJPE4XP6_0),.dout(w_dff_B_NqLTbuqA7_0),.clk(gclk));
	jdff dff_B_b2l72KXE0_0(.din(n1120),.dout(w_dff_B_b2l72KXE0_0),.clk(gclk));
	jdff dff_B_puZNNBTg3_0(.din(w_dff_B_b2l72KXE0_0),.dout(w_dff_B_puZNNBTg3_0),.clk(gclk));
	jdff dff_B_bqrvePcn8_0(.din(w_dff_B_puZNNBTg3_0),.dout(w_dff_B_bqrvePcn8_0),.clk(gclk));
	jdff dff_B_eR5ExF3L0_0(.din(w_dff_B_bqrvePcn8_0),.dout(w_dff_B_eR5ExF3L0_0),.clk(gclk));
	jdff dff_B_q3KNssiL8_0(.din(w_dff_B_eR5ExF3L0_0),.dout(w_dff_B_q3KNssiL8_0),.clk(gclk));
	jdff dff_B_HqQAKbo35_0(.din(w_dff_B_q3KNssiL8_0),.dout(w_dff_B_HqQAKbo35_0),.clk(gclk));
	jdff dff_A_hLumddvH0_0(.dout(w_n748_4[0]),.din(w_dff_A_hLumddvH0_0),.clk(gclk));
	jdff dff_A_FcZ1TBoQ8_1(.dout(w_G137_7[1]),.din(w_dff_A_FcZ1TBoQ8_1),.clk(gclk));
	jdff dff_A_Yt9IkgeX9_1(.dout(w_dff_A_FcZ1TBoQ8_1),.din(w_dff_A_Yt9IkgeX9_1),.clk(gclk));
	jdff dff_A_A7acxXNr1_1(.dout(w_dff_A_Yt9IkgeX9_1),.din(w_dff_A_A7acxXNr1_1),.clk(gclk));
	jdff dff_A_VV06EGpu8_1(.dout(w_dff_A_A7acxXNr1_1),.din(w_dff_A_VV06EGpu8_1),.clk(gclk));
	jdff dff_A_A2z92gkD7_2(.dout(w_G137_7[2]),.din(w_dff_A_A2z92gkD7_2),.clk(gclk));
	jdff dff_A_dScTuOOL0_2(.dout(w_dff_A_A2z92gkD7_2),.din(w_dff_A_dScTuOOL0_2),.clk(gclk));
	jdff dff_A_trArhmMH5_0(.dout(w_G137_2[0]),.din(w_dff_A_trArhmMH5_0),.clk(gclk));
	jdff dff_A_WX7dlkav2_0(.dout(w_dff_A_trArhmMH5_0),.din(w_dff_A_WX7dlkav2_0),.clk(gclk));
	jdff dff_A_JFdvwC3B2_0(.dout(w_dff_A_WX7dlkav2_0),.din(w_dff_A_JFdvwC3B2_0),.clk(gclk));
	jdff dff_A_j8iNbbck6_0(.dout(w_dff_A_JFdvwC3B2_0),.din(w_dff_A_j8iNbbck6_0),.clk(gclk));
	jdff dff_A_DDdwYcRt3_1(.dout(w_G137_2[1]),.din(w_dff_A_DDdwYcRt3_1),.clk(gclk));
	jdff dff_A_eilzWOxb9_1(.dout(w_dff_A_DDdwYcRt3_1),.din(w_dff_A_eilzWOxb9_1),.clk(gclk));
	jdff dff_A_vkpMb6d29_1(.dout(w_dff_A_eilzWOxb9_1),.din(w_dff_A_vkpMb6d29_1),.clk(gclk));
	jdff dff_A_0Jc3Av869_1(.dout(w_dff_A_vkpMb6d29_1),.din(w_dff_A_0Jc3Av869_1),.clk(gclk));
	jdff dff_B_Ui3Wbu158_0(.din(n1129),.dout(w_dff_B_Ui3Wbu158_0),.clk(gclk));
	jdff dff_B_iRjXtJ673_0(.din(w_dff_B_Ui3Wbu158_0),.dout(w_dff_B_iRjXtJ673_0),.clk(gclk));
	jdff dff_B_vx82K3jn8_0(.din(n1128),.dout(w_dff_B_vx82K3jn8_0),.clk(gclk));
	jdff dff_B_0JvGJIpZ7_0(.din(w_dff_B_vx82K3jn8_0),.dout(w_dff_B_0JvGJIpZ7_0),.clk(gclk));
	jdff dff_B_r3oxkau82_0(.din(w_dff_B_0JvGJIpZ7_0),.dout(w_dff_B_r3oxkau82_0),.clk(gclk));
	jdff dff_B_uAxXgHkX8_0(.din(w_dff_B_r3oxkau82_0),.dout(w_dff_B_uAxXgHkX8_0),.clk(gclk));
	jdff dff_B_zeKLxmuS2_0(.din(w_dff_B_uAxXgHkX8_0),.dout(w_dff_B_zeKLxmuS2_0),.clk(gclk));
	jdff dff_B_zUKjxpJd9_0(.din(w_dff_B_zeKLxmuS2_0),.dout(w_dff_B_zUKjxpJd9_0),.clk(gclk));
	jdff dff_B_gtojMpQM8_0(.din(w_dff_B_zUKjxpJd9_0),.dout(w_dff_B_gtojMpQM8_0),.clk(gclk));
	jdff dff_B_xyY6mh8V6_0(.din(w_dff_B_gtojMpQM8_0),.dout(w_dff_B_xyY6mh8V6_0),.clk(gclk));
	jdff dff_B_fUVttPHp4_0(.din(n837),.dout(w_dff_B_fUVttPHp4_0),.clk(gclk));
	jdff dff_B_WuXpcJCp9_0(.din(w_dff_B_fUVttPHp4_0),.dout(w_dff_B_WuXpcJCp9_0),.clk(gclk));
	jdff dff_A_ePj6LctY5_0(.dout(w_n744_1[0]),.din(w_dff_A_ePj6LctY5_0),.clk(gclk));
	jdff dff_A_erJPVHtM0_0(.dout(w_dff_A_ePj6LctY5_0),.din(w_dff_A_erJPVHtM0_0),.clk(gclk));
	jdff dff_A_mqkXTEC06_0(.dout(w_dff_A_erJPVHtM0_0),.din(w_dff_A_mqkXTEC06_0),.clk(gclk));
	jdff dff_A_QWQ1DtKV1_0(.dout(w_dff_A_mqkXTEC06_0),.din(w_dff_A_QWQ1DtKV1_0),.clk(gclk));
	jdff dff_A_6GtY2fWE3_0(.dout(w_dff_A_QWQ1DtKV1_0),.din(w_dff_A_6GtY2fWE3_0),.clk(gclk));
	jdff dff_A_NBhpaSKd4_0(.dout(w_dff_A_6GtY2fWE3_0),.din(w_dff_A_NBhpaSKd4_0),.clk(gclk));
	jdff dff_B_u7wzn8vO0_0(.din(n1137),.dout(w_dff_B_u7wzn8vO0_0),.clk(gclk));
	jdff dff_B_cVsXPlA27_0(.din(n1136),.dout(w_dff_B_cVsXPlA27_0),.clk(gclk));
	jdff dff_B_Ov8xtgzA0_0(.din(w_dff_B_cVsXPlA27_0),.dout(w_dff_B_Ov8xtgzA0_0),.clk(gclk));
	jdff dff_B_NJ97wETJ8_0(.din(w_dff_B_Ov8xtgzA0_0),.dout(w_dff_B_NJ97wETJ8_0),.clk(gclk));
	jdff dff_B_BFfsGoj11_0(.din(w_dff_B_NJ97wETJ8_0),.dout(w_dff_B_BFfsGoj11_0),.clk(gclk));
	jdff dff_B_VY4PXC7P1_0(.din(w_dff_B_BFfsGoj11_0),.dout(w_dff_B_VY4PXC7P1_0),.clk(gclk));
	jdff dff_B_Nc3HHK5z7_0(.din(w_dff_B_VY4PXC7P1_0),.dout(w_dff_B_Nc3HHK5z7_0),.clk(gclk));
	jdff dff_B_jdsmzO9M8_0(.din(w_dff_B_Nc3HHK5z7_0),.dout(w_dff_B_jdsmzO9M8_0),.clk(gclk));
	jdff dff_B_1x5XozI66_0(.din(w_dff_B_jdsmzO9M8_0),.dout(w_dff_B_1x5XozI66_0),.clk(gclk));
	jdff dff_B_1JQcsZdo7_0(.din(w_dff_B_1x5XozI66_0),.dout(w_dff_B_1JQcsZdo7_0),.clk(gclk));
	jdff dff_B_HC3u8Yfs7_0(.din(w_dff_B_1JQcsZdo7_0),.dout(w_dff_B_HC3u8Yfs7_0),.clk(gclk));
	jdff dff_A_AnsKQqqE0_0(.dout(w_n1002_3[0]),.din(w_dff_A_AnsKQqqE0_0),.clk(gclk));
	jdff dff_A_xLxi7wiR3_0(.dout(w_dff_A_AnsKQqqE0_0),.din(w_dff_A_xLxi7wiR3_0),.clk(gclk));
	jdff dff_A_UnNXMQmK4_0(.dout(w_dff_A_xLxi7wiR3_0),.din(w_dff_A_UnNXMQmK4_0),.clk(gclk));
	jdff dff_A_Lx5GNs0P4_0(.dout(w_dff_A_UnNXMQmK4_0),.din(w_dff_A_Lx5GNs0P4_0),.clk(gclk));
	jdff dff_A_iJuM50qB6_1(.dout(w_n1002_3[1]),.din(w_dff_A_iJuM50qB6_1),.clk(gclk));
	jdff dff_A_xd58JnAC1_1(.dout(w_dff_A_iJuM50qB6_1),.din(w_dff_A_xd58JnAC1_1),.clk(gclk));
	jdff dff_B_MFpA3PmB1_0(.din(n826),.dout(w_dff_B_MFpA3PmB1_0),.clk(gclk));
	jdff dff_B_h24csGr33_0(.din(w_dff_B_MFpA3PmB1_0),.dout(w_dff_B_h24csGr33_0),.clk(gclk));
	jdff dff_B_7bd266Fo3_0(.din(w_dff_B_h24csGr33_0),.dout(w_dff_B_7bd266Fo3_0),.clk(gclk));
	jdff dff_B_8e3r9I3s4_0(.din(w_dff_B_7bd266Fo3_0),.dout(w_dff_B_8e3r9I3s4_0),.clk(gclk));
	jdff dff_B_WIS3tm177_0(.din(w_dff_B_8e3r9I3s4_0),.dout(w_dff_B_WIS3tm177_0),.clk(gclk));
	jdff dff_B_edJd0PSN8_1(.din(n816),.dout(w_dff_B_edJd0PSN8_1),.clk(gclk));
	jdff dff_B_PFUI3WGK3_1(.din(w_dff_B_edJd0PSN8_1),.dout(w_dff_B_PFUI3WGK3_1),.clk(gclk));
	jdff dff_B_HBotJQtt4_1(.din(w_dff_B_PFUI3WGK3_1),.dout(w_dff_B_HBotJQtt4_1),.clk(gclk));
	jdff dff_B_YCA7qrw44_1(.din(w_dff_B_HBotJQtt4_1),.dout(w_dff_B_YCA7qrw44_1),.clk(gclk));
	jdff dff_B_w6uc7q442_1(.din(w_dff_B_YCA7qrw44_1),.dout(w_dff_B_w6uc7q442_1),.clk(gclk));
	jdff dff_A_eEVCHfL63_2(.dout(w_n744_0[2]),.din(w_dff_A_eEVCHfL63_2),.clk(gclk));
	jdff dff_A_TYG6RqQH6_2(.dout(w_dff_A_eEVCHfL63_2),.din(w_dff_A_TYG6RqQH6_2),.clk(gclk));
	jdff dff_A_BOUseHkY4_2(.dout(w_dff_A_TYG6RqQH6_2),.din(w_dff_A_BOUseHkY4_2),.clk(gclk));
	jdff dff_A_pQVO2DnM4_2(.dout(w_dff_A_BOUseHkY4_2),.din(w_dff_A_pQVO2DnM4_2),.clk(gclk));
	jdff dff_B_7Ckizk8O9_3(.din(n744),.dout(w_dff_B_7Ckizk8O9_3),.clk(gclk));
	jdff dff_B_5L8eXvRX9_3(.din(w_dff_B_7Ckizk8O9_3),.dout(w_dff_B_5L8eXvRX9_3),.clk(gclk));
	jdff dff_A_SbDorVq62_1(.dout(w_n748_3[1]),.din(w_dff_A_SbDorVq62_1),.clk(gclk));
	jdff dff_A_jFHnAu0m2_1(.dout(w_dff_A_SbDorVq62_1),.din(w_dff_A_jFHnAu0m2_1),.clk(gclk));
	jdff dff_A_zbrVtRZs8_2(.dout(w_n748_3[2]),.din(w_dff_A_zbrVtRZs8_2),.clk(gclk));
	jdff dff_A_aGlFT7kQ1_2(.dout(w_dff_A_zbrVtRZs8_2),.din(w_dff_A_aGlFT7kQ1_2),.clk(gclk));
	jdff dff_A_Xd5ZtYE87_2(.dout(w_dff_A_aGlFT7kQ1_2),.din(w_dff_A_Xd5ZtYE87_2),.clk(gclk));
	jdff dff_A_hufhjLzc9_2(.dout(w_dff_A_Xd5ZtYE87_2),.din(w_dff_A_hufhjLzc9_2),.clk(gclk));
	jdff dff_A_srgj378l7_0(.dout(w_n999_3[0]),.din(w_dff_A_srgj378l7_0),.clk(gclk));
	jdff dff_A_J3xX0R6e9_0(.dout(w_dff_A_srgj378l7_0),.din(w_dff_A_J3xX0R6e9_0),.clk(gclk));
	jdff dff_A_63C5xwlS3_1(.dout(w_n999_3[1]),.din(w_dff_A_63C5xwlS3_1),.clk(gclk));
	jdff dff_B_0MxfRhmf0_0(.din(n1155),.dout(w_dff_B_0MxfRhmf0_0),.clk(gclk));
	jdff dff_B_ZRRdUf0t4_0(.din(w_dff_B_0MxfRhmf0_0),.dout(w_dff_B_ZRRdUf0t4_0),.clk(gclk));
	jdff dff_B_Ad1FpN0L5_0(.din(w_dff_B_ZRRdUf0t4_0),.dout(w_dff_B_Ad1FpN0L5_0),.clk(gclk));
	jdff dff_B_0MQe6lWW1_0(.din(w_dff_B_Ad1FpN0L5_0),.dout(w_dff_B_0MQe6lWW1_0),.clk(gclk));
	jdff dff_B_oo6W34xP8_0(.din(w_dff_B_0MQe6lWW1_0),.dout(w_dff_B_oo6W34xP8_0),.clk(gclk));
	jdff dff_B_Ja4dFN6o6_0(.din(w_dff_B_oo6W34xP8_0),.dout(w_dff_B_Ja4dFN6o6_0),.clk(gclk));
	jdff dff_B_7lV4R1GT0_0(.din(w_dff_B_Ja4dFN6o6_0),.dout(w_dff_B_7lV4R1GT0_0),.clk(gclk));
	jdff dff_B_Ylw5k3Sn7_0(.din(w_dff_B_7lV4R1GT0_0),.dout(w_dff_B_Ylw5k3Sn7_0),.clk(gclk));
	jdff dff_B_rvqpqrK55_0(.din(w_dff_B_Ylw5k3Sn7_0),.dout(w_dff_B_rvqpqrK55_0),.clk(gclk));
	jdff dff_B_iPMnBdR27_0(.din(w_dff_B_rvqpqrK55_0),.dout(w_dff_B_iPMnBdR27_0),.clk(gclk));
	jdff dff_B_DC1GyhgS8_0(.din(w_dff_B_iPMnBdR27_0),.dout(w_dff_B_DC1GyhgS8_0),.clk(gclk));
	jdff dff_B_JCS4xw4h9_0(.din(w_dff_B_DC1GyhgS8_0),.dout(w_dff_B_JCS4xw4h9_0),.clk(gclk));
	jdff dff_B_0IB2FlBJ4_1(.din(n1148),.dout(w_dff_B_0IB2FlBJ4_1),.clk(gclk));
	jdff dff_B_h5U9nSjY9_1(.din(w_dff_B_0IB2FlBJ4_1),.dout(w_dff_B_h5U9nSjY9_1),.clk(gclk));
	jdff dff_B_yZnwq2mo7_1(.din(w_dff_B_h5U9nSjY9_1),.dout(w_dff_B_yZnwq2mo7_1),.clk(gclk));
	jdff dff_B_p7z6dGUC4_1(.din(w_dff_B_yZnwq2mo7_1),.dout(w_dff_B_p7z6dGUC4_1),.clk(gclk));
	jdff dff_B_pBkP35yK1_1(.din(w_dff_B_p7z6dGUC4_1),.dout(w_dff_B_pBkP35yK1_1),.clk(gclk));
	jdff dff_B_6brFvEQp9_1(.din(n1150),.dout(w_dff_B_6brFvEQp9_1),.clk(gclk));
	jdff dff_B_MKXPRiIA4_0(.din(n1144),.dout(w_dff_B_MKXPRiIA4_0),.clk(gclk));
	jdff dff_B_MSBtCVXB7_0(.din(w_dff_B_MKXPRiIA4_0),.dout(w_dff_B_MSBtCVXB7_0),.clk(gclk));
	jdff dff_B_cX4bX2wC5_0(.din(w_dff_B_MSBtCVXB7_0),.dout(w_dff_B_cX4bX2wC5_0),.clk(gclk));
	jdff dff_B_u3e0XFcK3_0(.din(w_dff_B_cX4bX2wC5_0),.dout(w_dff_B_u3e0XFcK3_0),.clk(gclk));
	jdff dff_B_Zh2vVE8k0_0(.din(w_dff_B_u3e0XFcK3_0),.dout(w_dff_B_Zh2vVE8k0_0),.clk(gclk));
	jdff dff_B_xAj5UnQL7_0(.din(w_dff_B_Zh2vVE8k0_0),.dout(w_dff_B_xAj5UnQL7_0),.clk(gclk));
	jdff dff_B_IOXXKdlo9_0(.din(w_dff_B_xAj5UnQL7_0),.dout(w_dff_B_IOXXKdlo9_0),.clk(gclk));
	jdff dff_B_6pfDf5zb1_0(.din(w_dff_B_IOXXKdlo9_0),.dout(w_dff_B_6pfDf5zb1_0),.clk(gclk));
	jdff dff_B_xgbodGGy8_0(.din(w_dff_B_6pfDf5zb1_0),.dout(w_dff_B_xgbodGGy8_0),.clk(gclk));
	jdff dff_B_r6MnnN211_0(.din(w_dff_B_xgbodGGy8_0),.dout(w_dff_B_r6MnnN211_0),.clk(gclk));
	jdff dff_B_TIgTC8974_0(.din(w_dff_B_r6MnnN211_0),.dout(w_dff_B_TIgTC8974_0),.clk(gclk));
	jdff dff_B_PyZvP6qq3_0(.din(w_dff_B_TIgTC8974_0),.dout(w_dff_B_PyZvP6qq3_0),.clk(gclk));
	jdff dff_B_SsieJO0D3_0(.din(w_dff_B_PyZvP6qq3_0),.dout(w_dff_B_SsieJO0D3_0),.clk(gclk));
	jdff dff_B_c9zkGq5W6_0(.din(w_dff_B_SsieJO0D3_0),.dout(w_dff_B_c9zkGq5W6_0),.clk(gclk));
	jdff dff_B_qi0isgWG9_0(.din(w_dff_B_c9zkGq5W6_0),.dout(w_dff_B_qi0isgWG9_0),.clk(gclk));
	jdff dff_B_mGPgZ6e00_0(.din(w_dff_B_qi0isgWG9_0),.dout(w_dff_B_mGPgZ6e00_0),.clk(gclk));
	jdff dff_A_ZpDx0m9G7_0(.dout(w_G132_0[0]),.din(w_dff_A_ZpDx0m9G7_0),.clk(gclk));
	jdff dff_A_SdFcJZea0_0(.dout(w_dff_A_ZpDx0m9G7_0),.din(w_dff_A_SdFcJZea0_0),.clk(gclk));
	jdff dff_A_eb7nZeEv0_0(.dout(w_dff_A_SdFcJZea0_0),.din(w_dff_A_eb7nZeEv0_0),.clk(gclk));
	jdff dff_A_S9FFe9xl5_0(.dout(w_dff_A_eb7nZeEv0_0),.din(w_dff_A_S9FFe9xl5_0),.clk(gclk));
	jdff dff_A_dqGPOkbq0_0(.dout(w_dff_A_S9FFe9xl5_0),.din(w_dff_A_dqGPOkbq0_0),.clk(gclk));
	jdff dff_A_DfsfmLgO2_0(.dout(w_dff_A_dqGPOkbq0_0),.din(w_dff_A_DfsfmLgO2_0),.clk(gclk));
	jdff dff_A_URXsBbbI2_0(.dout(w_dff_A_DfsfmLgO2_0),.din(w_dff_A_URXsBbbI2_0),.clk(gclk));
	jdff dff_A_dxTqvqTy7_0(.dout(w_dff_A_URXsBbbI2_0),.din(w_dff_A_dxTqvqTy7_0),.clk(gclk));
	jdff dff_A_AFd7f6Rv8_0(.dout(w_dff_A_dxTqvqTy7_0),.din(w_dff_A_AFd7f6Rv8_0),.clk(gclk));
	jdff dff_A_lcN9nOVf8_0(.dout(w_dff_A_AFd7f6Rv8_0),.din(w_dff_A_lcN9nOVf8_0),.clk(gclk));
	jdff dff_A_xdHQU8AK9_0(.dout(w_dff_A_lcN9nOVf8_0),.din(w_dff_A_xdHQU8AK9_0),.clk(gclk));
	jdff dff_A_wAknh2uT2_0(.dout(w_dff_A_xdHQU8AK9_0),.din(w_dff_A_wAknh2uT2_0),.clk(gclk));
	jdff dff_A_W3xZVqvd4_0(.dout(w_dff_A_wAknh2uT2_0),.din(w_dff_A_W3xZVqvd4_0),.clk(gclk));
	jdff dff_B_wozXgap33_2(.din(G132),.dout(w_dff_B_wozXgap33_2),.clk(gclk));
	jdff dff_B_9FQwUB159_2(.din(w_dff_B_wozXgap33_2),.dout(w_dff_B_9FQwUB159_2),.clk(gclk));
	jdff dff_B_06mJDRfX3_2(.din(w_dff_B_9FQwUB159_2),.dout(w_dff_B_06mJDRfX3_2),.clk(gclk));
	jdff dff_B_eyaGwMpD4_1(.din(n1184),.dout(w_dff_B_eyaGwMpD4_1),.clk(gclk));
	jdff dff_B_ABuABlaC9_0(.din(n1189),.dout(w_dff_B_ABuABlaC9_0),.clk(gclk));
	jdff dff_B_nZg96tG07_0(.din(w_dff_B_ABuABlaC9_0),.dout(w_dff_B_nZg96tG07_0),.clk(gclk));
	jdff dff_B_KhItkqzk3_0(.din(n1187),.dout(w_dff_B_KhItkqzk3_0),.clk(gclk));
	jdff dff_A_Ie9xyNkC3_0(.dout(w_G601_0),.din(w_dff_A_Ie9xyNkC3_0),.clk(gclk));
	jdff dff_A_xUU0Go5l4_0(.dout(w_n671_0[0]),.din(w_dff_A_xUU0Go5l4_0),.clk(gclk));
	jdff dff_B_dS2amFQa1_1(.din(n907),.dout(w_dff_B_dS2amFQa1_1),.clk(gclk));
	jdff dff_B_plUzJaFz2_1(.din(n909),.dout(w_dff_B_plUzJaFz2_1),.clk(gclk));
	jdff dff_B_sllcrRqo5_1(.din(w_dff_B_plUzJaFz2_1),.dout(w_dff_B_sllcrRqo5_1),.clk(gclk));
	jdff dff_B_QTcJ8GD28_0(.din(n910),.dout(w_dff_B_QTcJ8GD28_0),.clk(gclk));
	jdff dff_B_Xa60deEF0_1(.din(n908),.dout(w_dff_B_Xa60deEF0_1),.clk(gclk));
	jdff dff_A_F5GbhCwJ8_0(.dout(w_n621_1[0]),.din(w_dff_A_F5GbhCwJ8_0),.clk(gclk));
	jdff dff_A_k1WEk1cg5_0(.dout(w_dff_A_F5GbhCwJ8_0),.din(w_dff_A_k1WEk1cg5_0),.clk(gclk));
	jdff dff_A_g2qvW19T6_0(.dout(w_dff_A_k1WEk1cg5_0),.din(w_dff_A_g2qvW19T6_0),.clk(gclk));
	jdff dff_B_EotxGwAx0_0(.din(n1224),.dout(w_dff_B_EotxGwAx0_0),.clk(gclk));
	jdff dff_B_iTkLQcMp7_0(.din(w_dff_B_EotxGwAx0_0),.dout(w_dff_B_iTkLQcMp7_0),.clk(gclk));
	jdff dff_B_rdP2cBpa7_0(.din(w_dff_B_iTkLQcMp7_0),.dout(w_dff_B_rdP2cBpa7_0),.clk(gclk));
	jdff dff_B_mHxqDbkI9_0(.din(w_dff_B_rdP2cBpa7_0),.dout(w_dff_B_mHxqDbkI9_0),.clk(gclk));
	jdff dff_B_dydXWkAG1_0(.din(w_dff_B_mHxqDbkI9_0),.dout(w_dff_B_dydXWkAG1_0),.clk(gclk));
	jdff dff_B_cNIQDl6x0_0(.din(w_dff_B_dydXWkAG1_0),.dout(w_dff_B_cNIQDl6x0_0),.clk(gclk));
	jdff dff_B_hC8IRBhE2_0(.din(w_dff_B_cNIQDl6x0_0),.dout(w_dff_B_hC8IRBhE2_0),.clk(gclk));
	jdff dff_B_wMdryTNs7_0(.din(w_dff_B_hC8IRBhE2_0),.dout(w_dff_B_wMdryTNs7_0),.clk(gclk));
	jdff dff_B_tSRR7OHY0_0(.din(w_dff_B_wMdryTNs7_0),.dout(w_dff_B_tSRR7OHY0_0),.clk(gclk));
	jdff dff_B_eQlnZ8Qu4_0(.din(w_dff_B_tSRR7OHY0_0),.dout(w_dff_B_eQlnZ8Qu4_0),.clk(gclk));
	jdff dff_B_HoKMSo2h1_0(.din(w_dff_B_eQlnZ8Qu4_0),.dout(w_dff_B_HoKMSo2h1_0),.clk(gclk));
	jdff dff_B_Cx6fu5b54_0(.din(w_dff_B_HoKMSo2h1_0),.dout(w_dff_B_Cx6fu5b54_0),.clk(gclk));
	jdff dff_B_Mhreckzp8_0(.din(w_dff_B_Cx6fu5b54_0),.dout(w_dff_B_Mhreckzp8_0),.clk(gclk));
	jdff dff_B_vUORmcoW8_0(.din(w_dff_B_Mhreckzp8_0),.dout(w_dff_B_vUORmcoW8_0),.clk(gclk));
	jdff dff_B_s4r1RweA3_0(.din(w_dff_B_vUORmcoW8_0),.dout(w_dff_B_s4r1RweA3_0),.clk(gclk));
	jdff dff_B_q1B1dQ8c0_0(.din(w_dff_B_s4r1RweA3_0),.dout(w_dff_B_q1B1dQ8c0_0),.clk(gclk));
	jdff dff_B_ENRx4VdZ0_0(.din(w_dff_B_q1B1dQ8c0_0),.dout(w_dff_B_ENRx4VdZ0_0),.clk(gclk));
	jdff dff_B_8dfXrwUE8_0(.din(n1231),.dout(w_dff_B_8dfXrwUE8_0),.clk(gclk));
	jdff dff_B_2pSBb1It8_0(.din(w_dff_B_8dfXrwUE8_0),.dout(w_dff_B_2pSBb1It8_0),.clk(gclk));
	jdff dff_B_nn2TNj9B1_0(.din(w_dff_B_2pSBb1It8_0),.dout(w_dff_B_nn2TNj9B1_0),.clk(gclk));
	jdff dff_B_XSuppEvn0_0(.din(w_dff_B_nn2TNj9B1_0),.dout(w_dff_B_XSuppEvn0_0),.clk(gclk));
	jdff dff_B_LUp4y5Es7_0(.din(w_dff_B_XSuppEvn0_0),.dout(w_dff_B_LUp4y5Es7_0),.clk(gclk));
	jdff dff_B_rIokX5MD0_0(.din(w_dff_B_LUp4y5Es7_0),.dout(w_dff_B_rIokX5MD0_0),.clk(gclk));
	jdff dff_B_WJz1cW5s9_0(.din(w_dff_B_rIokX5MD0_0),.dout(w_dff_B_WJz1cW5s9_0),.clk(gclk));
	jdff dff_B_M1ugVF4f8_0(.din(w_dff_B_WJz1cW5s9_0),.dout(w_dff_B_M1ugVF4f8_0),.clk(gclk));
	jdff dff_B_HJI0caO23_0(.din(w_dff_B_M1ugVF4f8_0),.dout(w_dff_B_HJI0caO23_0),.clk(gclk));
	jdff dff_B_cTn7yaGx3_0(.din(w_dff_B_HJI0caO23_0),.dout(w_dff_B_cTn7yaGx3_0),.clk(gclk));
	jdff dff_B_mfFp6fPu3_0(.din(w_dff_B_cTn7yaGx3_0),.dout(w_dff_B_mfFp6fPu3_0),.clk(gclk));
	jdff dff_B_DoSfxQP35_0(.din(w_dff_B_mfFp6fPu3_0),.dout(w_dff_B_DoSfxQP35_0),.clk(gclk));
	jdff dff_B_74honPYO8_0(.din(w_dff_B_DoSfxQP35_0),.dout(w_dff_B_74honPYO8_0),.clk(gclk));
	jdff dff_B_x6LEa6qZ5_0(.din(w_dff_B_74honPYO8_0),.dout(w_dff_B_x6LEa6qZ5_0),.clk(gclk));
	jdff dff_B_1P5ecuwR7_0(.din(w_dff_B_x6LEa6qZ5_0),.dout(w_dff_B_1P5ecuwR7_0),.clk(gclk));
	jdff dff_B_PvSL4RGA3_0(.din(w_dff_B_1P5ecuwR7_0),.dout(w_dff_B_PvSL4RGA3_0),.clk(gclk));
	jdff dff_B_b4hchHMT6_0(.din(w_dff_B_PvSL4RGA3_0),.dout(w_dff_B_b4hchHMT6_0),.clk(gclk));
	jdff dff_B_jEu3uKf42_0(.din(n1239),.dout(w_dff_B_jEu3uKf42_0),.clk(gclk));
	jdff dff_B_N0FrtKqe5_0(.din(w_dff_B_jEu3uKf42_0),.dout(w_dff_B_N0FrtKqe5_0),.clk(gclk));
	jdff dff_B_mS3eU0v09_0(.din(w_dff_B_N0FrtKqe5_0),.dout(w_dff_B_mS3eU0v09_0),.clk(gclk));
	jdff dff_B_JS06cY6x5_0(.din(w_dff_B_mS3eU0v09_0),.dout(w_dff_B_JS06cY6x5_0),.clk(gclk));
	jdff dff_B_00goqtmS8_0(.din(w_dff_B_JS06cY6x5_0),.dout(w_dff_B_00goqtmS8_0),.clk(gclk));
	jdff dff_B_3SBlXBzr3_0(.din(w_dff_B_00goqtmS8_0),.dout(w_dff_B_3SBlXBzr3_0),.clk(gclk));
	jdff dff_B_cMs4zbZn3_0(.din(w_dff_B_3SBlXBzr3_0),.dout(w_dff_B_cMs4zbZn3_0),.clk(gclk));
	jdff dff_B_n1GR9eCH5_0(.din(w_dff_B_cMs4zbZn3_0),.dout(w_dff_B_n1GR9eCH5_0),.clk(gclk));
	jdff dff_B_QRYJSOMe6_0(.din(w_dff_B_n1GR9eCH5_0),.dout(w_dff_B_QRYJSOMe6_0),.clk(gclk));
	jdff dff_B_5ktwBSEr4_0(.din(w_dff_B_QRYJSOMe6_0),.dout(w_dff_B_5ktwBSEr4_0),.clk(gclk));
	jdff dff_B_R2YyRbre9_0(.din(w_dff_B_5ktwBSEr4_0),.dout(w_dff_B_R2YyRbre9_0),.clk(gclk));
	jdff dff_B_0PBvX6cm9_0(.din(w_dff_B_R2YyRbre9_0),.dout(w_dff_B_0PBvX6cm9_0),.clk(gclk));
	jdff dff_B_dKlhZPq20_0(.din(w_dff_B_0PBvX6cm9_0),.dout(w_dff_B_dKlhZPq20_0),.clk(gclk));
	jdff dff_B_1Us2ToPD9_0(.din(w_dff_B_dKlhZPq20_0),.dout(w_dff_B_1Us2ToPD9_0),.clk(gclk));
	jdff dff_B_LH6IW6O59_0(.din(w_dff_B_1Us2ToPD9_0),.dout(w_dff_B_LH6IW6O59_0),.clk(gclk));
	jdff dff_B_QDtKQf1m5_0(.din(w_dff_B_LH6IW6O59_0),.dout(w_dff_B_QDtKQf1m5_0),.clk(gclk));
	jdff dff_B_C9N0WaPe6_0(.din(n1248),.dout(w_dff_B_C9N0WaPe6_0),.clk(gclk));
	jdff dff_B_0snA5S6R4_0(.din(w_dff_B_C9N0WaPe6_0),.dout(w_dff_B_0snA5S6R4_0),.clk(gclk));
	jdff dff_B_fayqID8R3_0(.din(w_dff_B_0snA5S6R4_0),.dout(w_dff_B_fayqID8R3_0),.clk(gclk));
	jdff dff_B_RM4lGBpA6_0(.din(w_dff_B_fayqID8R3_0),.dout(w_dff_B_RM4lGBpA6_0),.clk(gclk));
	jdff dff_B_2YJFvSrb2_0(.din(w_dff_B_RM4lGBpA6_0),.dout(w_dff_B_2YJFvSrb2_0),.clk(gclk));
	jdff dff_B_Bbhvj9oR7_0(.din(w_dff_B_2YJFvSrb2_0),.dout(w_dff_B_Bbhvj9oR7_0),.clk(gclk));
	jdff dff_B_gppSaH1L6_0(.din(w_dff_B_Bbhvj9oR7_0),.dout(w_dff_B_gppSaH1L6_0),.clk(gclk));
	jdff dff_B_migT0Gto1_0(.din(w_dff_B_gppSaH1L6_0),.dout(w_dff_B_migT0Gto1_0),.clk(gclk));
	jdff dff_B_nMECjpHA2_0(.din(w_dff_B_migT0Gto1_0),.dout(w_dff_B_nMECjpHA2_0),.clk(gclk));
	jdff dff_B_0DyUbfF35_0(.din(w_dff_B_nMECjpHA2_0),.dout(w_dff_B_0DyUbfF35_0),.clk(gclk));
	jdff dff_B_c7B0cfh38_0(.din(w_dff_B_0DyUbfF35_0),.dout(w_dff_B_c7B0cfh38_0),.clk(gclk));
	jdff dff_B_fqtFCQS57_0(.din(w_dff_B_c7B0cfh38_0),.dout(w_dff_B_fqtFCQS57_0),.clk(gclk));
	jdff dff_B_QXjM2iX20_0(.din(w_dff_B_fqtFCQS57_0),.dout(w_dff_B_QXjM2iX20_0),.clk(gclk));
	jdff dff_B_sQDB2RRH4_0(.din(w_dff_B_QXjM2iX20_0),.dout(w_dff_B_sQDB2RRH4_0),.clk(gclk));
	jdff dff_B_HLbwSYic4_0(.din(w_dff_B_sQDB2RRH4_0),.dout(w_dff_B_HLbwSYic4_0),.clk(gclk));
	jdff dff_B_AEJFMYQM6_0(.din(w_dff_B_HLbwSYic4_0),.dout(w_dff_B_AEJFMYQM6_0),.clk(gclk));
	jdff dff_A_5qNoMRjg8_2(.dout(w_n797_2[2]),.din(w_dff_A_5qNoMRjg8_2),.clk(gclk));
	jdff dff_B_CNQBkg7b9_0(.din(n1257),.dout(w_dff_B_CNQBkg7b9_0),.clk(gclk));
	jdff dff_B_vc34ktVE2_0(.din(w_dff_B_CNQBkg7b9_0),.dout(w_dff_B_vc34ktVE2_0),.clk(gclk));
	jdff dff_B_KRdhPSbg3_0(.din(w_dff_B_vc34ktVE2_0),.dout(w_dff_B_KRdhPSbg3_0),.clk(gclk));
	jdff dff_B_TtdLE9hd2_0(.din(w_dff_B_KRdhPSbg3_0),.dout(w_dff_B_TtdLE9hd2_0),.clk(gclk));
	jdff dff_B_ruwOShWD6_0(.din(w_dff_B_TtdLE9hd2_0),.dout(w_dff_B_ruwOShWD6_0),.clk(gclk));
	jdff dff_B_cyu3NbDF3_0(.din(w_dff_B_ruwOShWD6_0),.dout(w_dff_B_cyu3NbDF3_0),.clk(gclk));
	jdff dff_B_FUk0zazF8_0(.din(w_dff_B_cyu3NbDF3_0),.dout(w_dff_B_FUk0zazF8_0),.clk(gclk));
	jdff dff_B_T2qaG3YU5_0(.din(w_dff_B_FUk0zazF8_0),.dout(w_dff_B_T2qaG3YU5_0),.clk(gclk));
	jdff dff_B_exC4SqlK1_0(.din(w_dff_B_T2qaG3YU5_0),.dout(w_dff_B_exC4SqlK1_0),.clk(gclk));
	jdff dff_B_VzWR4oNC5_0(.din(w_dff_B_exC4SqlK1_0),.dout(w_dff_B_VzWR4oNC5_0),.clk(gclk));
	jdff dff_B_no18nUS60_0(.din(w_dff_B_VzWR4oNC5_0),.dout(w_dff_B_no18nUS60_0),.clk(gclk));
	jdff dff_B_RalU1xJW2_0(.din(w_dff_B_no18nUS60_0),.dout(w_dff_B_RalU1xJW2_0),.clk(gclk));
	jdff dff_B_VrJ1q9iA0_0(.din(w_dff_B_RalU1xJW2_0),.dout(w_dff_B_VrJ1q9iA0_0),.clk(gclk));
	jdff dff_B_1n95tzUM9_0(.din(w_dff_B_VrJ1q9iA0_0),.dout(w_dff_B_1n95tzUM9_0),.clk(gclk));
	jdff dff_B_KgDYaSie1_0(.din(w_dff_B_1n95tzUM9_0),.dout(w_dff_B_KgDYaSie1_0),.clk(gclk));
	jdff dff_B_lwEbFgj60_0(.din(n1264),.dout(w_dff_B_lwEbFgj60_0),.clk(gclk));
	jdff dff_B_Gkg6xUWo8_0(.din(w_dff_B_lwEbFgj60_0),.dout(w_dff_B_Gkg6xUWo8_0),.clk(gclk));
	jdff dff_B_GqIl0CA70_0(.din(w_dff_B_Gkg6xUWo8_0),.dout(w_dff_B_GqIl0CA70_0),.clk(gclk));
	jdff dff_B_3joDtvDu4_0(.din(w_dff_B_GqIl0CA70_0),.dout(w_dff_B_3joDtvDu4_0),.clk(gclk));
	jdff dff_B_IUhWtjRK8_0(.din(w_dff_B_3joDtvDu4_0),.dout(w_dff_B_IUhWtjRK8_0),.clk(gclk));
	jdff dff_B_hl0ZoUVV2_0(.din(w_dff_B_IUhWtjRK8_0),.dout(w_dff_B_hl0ZoUVV2_0),.clk(gclk));
	jdff dff_B_aY2qJ7Uj7_0(.din(w_dff_B_hl0ZoUVV2_0),.dout(w_dff_B_aY2qJ7Uj7_0),.clk(gclk));
	jdff dff_B_bG8jNRRN5_0(.din(w_dff_B_aY2qJ7Uj7_0),.dout(w_dff_B_bG8jNRRN5_0),.clk(gclk));
	jdff dff_B_BuaV49N24_0(.din(w_dff_B_bG8jNRRN5_0),.dout(w_dff_B_BuaV49N24_0),.clk(gclk));
	jdff dff_B_bQcKaRrB8_0(.din(w_dff_B_BuaV49N24_0),.dout(w_dff_B_bQcKaRrB8_0),.clk(gclk));
	jdff dff_B_6lcXngbE4_0(.din(w_dff_B_bQcKaRrB8_0),.dout(w_dff_B_6lcXngbE4_0),.clk(gclk));
	jdff dff_B_2glnAwbx2_0(.din(w_dff_B_6lcXngbE4_0),.dout(w_dff_B_2glnAwbx2_0),.clk(gclk));
	jdff dff_B_DzuMuKFa3_0(.din(w_dff_B_2glnAwbx2_0),.dout(w_dff_B_DzuMuKFa3_0),.clk(gclk));
	jdff dff_B_AppQ0ae82_0(.din(w_dff_B_DzuMuKFa3_0),.dout(w_dff_B_AppQ0ae82_0),.clk(gclk));
	jdff dff_B_6vpdyqyI3_0(.din(w_dff_B_AppQ0ae82_0),.dout(w_dff_B_6vpdyqyI3_0),.clk(gclk));
	jdff dff_B_q4CWaEu15_0(.din(w_dff_B_6vpdyqyI3_0),.dout(w_dff_B_q4CWaEu15_0),.clk(gclk));
	jdff dff_B_YoO9hlOX4_0(.din(n1271),.dout(w_dff_B_YoO9hlOX4_0),.clk(gclk));
	jdff dff_B_DTuPXmxO9_0(.din(w_dff_B_YoO9hlOX4_0),.dout(w_dff_B_DTuPXmxO9_0),.clk(gclk));
	jdff dff_B_igmCWPGS9_0(.din(w_dff_B_DTuPXmxO9_0),.dout(w_dff_B_igmCWPGS9_0),.clk(gclk));
	jdff dff_B_ezbEN3bN9_0(.din(w_dff_B_igmCWPGS9_0),.dout(w_dff_B_ezbEN3bN9_0),.clk(gclk));
	jdff dff_B_iXRED5V68_0(.din(w_dff_B_ezbEN3bN9_0),.dout(w_dff_B_iXRED5V68_0),.clk(gclk));
	jdff dff_B_zItBIIjr8_0(.din(w_dff_B_iXRED5V68_0),.dout(w_dff_B_zItBIIjr8_0),.clk(gclk));
	jdff dff_B_nmIXI8LO8_0(.din(w_dff_B_zItBIIjr8_0),.dout(w_dff_B_nmIXI8LO8_0),.clk(gclk));
	jdff dff_B_pN6pqK9c2_0(.din(w_dff_B_nmIXI8LO8_0),.dout(w_dff_B_pN6pqK9c2_0),.clk(gclk));
	jdff dff_B_ufYIeoxd5_0(.din(w_dff_B_pN6pqK9c2_0),.dout(w_dff_B_ufYIeoxd5_0),.clk(gclk));
	jdff dff_B_QgVjl2Fm4_0(.din(w_dff_B_ufYIeoxd5_0),.dout(w_dff_B_QgVjl2Fm4_0),.clk(gclk));
	jdff dff_B_AT4Ksb5E8_0(.din(w_dff_B_QgVjl2Fm4_0),.dout(w_dff_B_AT4Ksb5E8_0),.clk(gclk));
	jdff dff_B_gQBlGxro9_0(.din(w_dff_B_AT4Ksb5E8_0),.dout(w_dff_B_gQBlGxro9_0),.clk(gclk));
	jdff dff_B_bvJjKRG98_0(.din(w_dff_B_gQBlGxro9_0),.dout(w_dff_B_bvJjKRG98_0),.clk(gclk));
	jdff dff_B_pPT8A5wd8_0(.din(w_dff_B_bvJjKRG98_0),.dout(w_dff_B_pPT8A5wd8_0),.clk(gclk));
	jdff dff_B_6GmiaF7s2_0(.din(w_dff_B_pPT8A5wd8_0),.dout(w_dff_B_6GmiaF7s2_0),.clk(gclk));
	jdff dff_B_E8rqHHnu5_0(.din(w_dff_B_6GmiaF7s2_0),.dout(w_dff_B_E8rqHHnu5_0),.clk(gclk));
	jdff dff_A_gYn5Hg3Q0_2(.dout(w_n843_2[2]),.din(w_dff_A_gYn5Hg3Q0_2),.clk(gclk));
	jdff dff_B_iNXZlW3r2_0(.din(n1278),.dout(w_dff_B_iNXZlW3r2_0),.clk(gclk));
	jdff dff_B_3y4FPi4V0_0(.din(w_dff_B_iNXZlW3r2_0),.dout(w_dff_B_3y4FPi4V0_0),.clk(gclk));
	jdff dff_B_PXcxPdDC5_0(.din(w_dff_B_3y4FPi4V0_0),.dout(w_dff_B_PXcxPdDC5_0),.clk(gclk));
	jdff dff_B_viHkD6KI0_0(.din(w_dff_B_PXcxPdDC5_0),.dout(w_dff_B_viHkD6KI0_0),.clk(gclk));
	jdff dff_B_1S0oTDmG0_0(.din(w_dff_B_viHkD6KI0_0),.dout(w_dff_B_1S0oTDmG0_0),.clk(gclk));
	jdff dff_B_jAVwv1X53_0(.din(w_dff_B_1S0oTDmG0_0),.dout(w_dff_B_jAVwv1X53_0),.clk(gclk));
	jdff dff_B_d1yc9kdY1_0(.din(w_dff_B_jAVwv1X53_0),.dout(w_dff_B_d1yc9kdY1_0),.clk(gclk));
	jdff dff_B_GCeIe2qI6_0(.din(w_dff_B_d1yc9kdY1_0),.dout(w_dff_B_GCeIe2qI6_0),.clk(gclk));
	jdff dff_B_IeY6iOT53_0(.din(w_dff_B_GCeIe2qI6_0),.dout(w_dff_B_IeY6iOT53_0),.clk(gclk));
	jdff dff_B_u8gcdKr60_0(.din(w_dff_B_IeY6iOT53_0),.dout(w_dff_B_u8gcdKr60_0),.clk(gclk));
	jdff dff_B_kraurtIm3_0(.din(w_dff_B_u8gcdKr60_0),.dout(w_dff_B_kraurtIm3_0),.clk(gclk));
	jdff dff_B_LWL3Bvv69_0(.din(w_dff_B_kraurtIm3_0),.dout(w_dff_B_LWL3Bvv69_0),.clk(gclk));
	jdff dff_B_wucsWPP73_0(.din(w_dff_B_LWL3Bvv69_0),.dout(w_dff_B_wucsWPP73_0),.clk(gclk));
	jdff dff_B_QrDz30uT0_0(.din(w_dff_B_wucsWPP73_0),.dout(w_dff_B_QrDz30uT0_0),.clk(gclk));
	jdff dff_B_Qel3kc1U0_0(.din(w_dff_B_QrDz30uT0_0),.dout(w_dff_B_Qel3kc1U0_0),.clk(gclk));
	jdff dff_B_LuOho6Yf9_0(.din(n1285),.dout(w_dff_B_LuOho6Yf9_0),.clk(gclk));
	jdff dff_B_rA7zrRTu0_0(.din(w_dff_B_LuOho6Yf9_0),.dout(w_dff_B_rA7zrRTu0_0),.clk(gclk));
	jdff dff_B_HqvYioco9_0(.din(w_dff_B_rA7zrRTu0_0),.dout(w_dff_B_HqvYioco9_0),.clk(gclk));
	jdff dff_B_BVNuGsYc6_0(.din(w_dff_B_HqvYioco9_0),.dout(w_dff_B_BVNuGsYc6_0),.clk(gclk));
	jdff dff_B_DwTJcZbn1_0(.din(w_dff_B_BVNuGsYc6_0),.dout(w_dff_B_DwTJcZbn1_0),.clk(gclk));
	jdff dff_B_vHm2o6g43_0(.din(w_dff_B_DwTJcZbn1_0),.dout(w_dff_B_vHm2o6g43_0),.clk(gclk));
	jdff dff_B_cHcW2Ou94_0(.din(w_dff_B_vHm2o6g43_0),.dout(w_dff_B_cHcW2Ou94_0),.clk(gclk));
	jdff dff_B_2Mh2Rxch6_0(.din(w_dff_B_cHcW2Ou94_0),.dout(w_dff_B_2Mh2Rxch6_0),.clk(gclk));
	jdff dff_B_Qbcn8qdw5_0(.din(w_dff_B_2Mh2Rxch6_0),.dout(w_dff_B_Qbcn8qdw5_0),.clk(gclk));
	jdff dff_B_PECfEeY57_0(.din(w_dff_B_Qbcn8qdw5_0),.dout(w_dff_B_PECfEeY57_0),.clk(gclk));
	jdff dff_B_LZ01Pdfs7_0(.din(w_dff_B_PECfEeY57_0),.dout(w_dff_B_LZ01Pdfs7_0),.clk(gclk));
	jdff dff_B_cgEPQjgE8_0(.din(w_dff_B_LZ01Pdfs7_0),.dout(w_dff_B_cgEPQjgE8_0),.clk(gclk));
	jdff dff_B_nACt00vD2_0(.din(w_dff_B_cgEPQjgE8_0),.dout(w_dff_B_nACt00vD2_0),.clk(gclk));
	jdff dff_B_Io3g9NpZ5_0(.din(w_dff_B_nACt00vD2_0),.dout(w_dff_B_Io3g9NpZ5_0),.clk(gclk));
	jdff dff_B_ivEV8khi6_0(.din(w_dff_B_Io3g9NpZ5_0),.dout(w_dff_B_ivEV8khi6_0),.clk(gclk));
	jdff dff_A_FNWn3Sj62_0(.dout(w_G137_6[0]),.din(w_dff_A_FNWn3Sj62_0),.clk(gclk));
	jdff dff_A_ijzbJFWI3_0(.dout(w_dff_A_FNWn3Sj62_0),.din(w_dff_A_ijzbJFWI3_0),.clk(gclk));
	jdff dff_A_tq1U0GGZ5_0(.dout(w_dff_A_ijzbJFWI3_0),.din(w_dff_A_tq1U0GGZ5_0),.clk(gclk));
	jdff dff_A_eaCfkIxx1_0(.dout(w_dff_A_tq1U0GGZ5_0),.din(w_dff_A_eaCfkIxx1_0),.clk(gclk));
	jdff dff_A_aTLt1TvC9_0(.dout(w_dff_A_eaCfkIxx1_0),.din(w_dff_A_aTLt1TvC9_0),.clk(gclk));
	jdff dff_A_gnvf12y66_1(.dout(w_G137_6[1]),.din(w_dff_A_gnvf12y66_1),.clk(gclk));
	jdff dff_B_fIhC1bEs2_0(.din(n1293),.dout(w_dff_B_fIhC1bEs2_0),.clk(gclk));
	jdff dff_B_55U8fgP86_0(.din(w_dff_B_fIhC1bEs2_0),.dout(w_dff_B_55U8fgP86_0),.clk(gclk));
	jdff dff_B_aFEG09Le2_0(.din(w_dff_B_55U8fgP86_0),.dout(w_dff_B_aFEG09Le2_0),.clk(gclk));
	jdff dff_B_pwyNGTQH1_0(.din(w_dff_B_aFEG09Le2_0),.dout(w_dff_B_pwyNGTQH1_0),.clk(gclk));
	jdff dff_B_YEozEZos9_0(.din(w_dff_B_pwyNGTQH1_0),.dout(w_dff_B_YEozEZos9_0),.clk(gclk));
	jdff dff_B_05XECJyc3_0(.din(w_dff_B_YEozEZos9_0),.dout(w_dff_B_05XECJyc3_0),.clk(gclk));
	jdff dff_B_o7snKGUJ2_0(.din(w_dff_B_05XECJyc3_0),.dout(w_dff_B_o7snKGUJ2_0),.clk(gclk));
	jdff dff_B_TqTnbU8u1_0(.din(w_dff_B_o7snKGUJ2_0),.dout(w_dff_B_TqTnbU8u1_0),.clk(gclk));
	jdff dff_B_gMtFwqZE5_0(.din(w_dff_B_TqTnbU8u1_0),.dout(w_dff_B_gMtFwqZE5_0),.clk(gclk));
	jdff dff_B_UMhhWcBC5_0(.din(w_dff_B_gMtFwqZE5_0),.dout(w_dff_B_UMhhWcBC5_0),.clk(gclk));
	jdff dff_B_tzW2bO0a6_0(.din(w_dff_B_UMhhWcBC5_0),.dout(w_dff_B_tzW2bO0a6_0),.clk(gclk));
	jdff dff_B_X6DAxqdc9_0(.din(w_dff_B_tzW2bO0a6_0),.dout(w_dff_B_X6DAxqdc9_0),.clk(gclk));
	jdff dff_B_QQPVuDjs5_0(.din(w_dff_B_X6DAxqdc9_0),.dout(w_dff_B_QQPVuDjs5_0),.clk(gclk));
	jdff dff_B_0UfmfBky0_0(.din(w_dff_B_QQPVuDjs5_0),.dout(w_dff_B_0UfmfBky0_0),.clk(gclk));
	jdff dff_B_AkQAFKTD6_0(.din(w_dff_B_0UfmfBky0_0),.dout(w_dff_B_AkQAFKTD6_0),.clk(gclk));
	jdff dff_B_7cxBKTql8_0(.din(w_dff_B_AkQAFKTD6_0),.dout(w_dff_B_7cxBKTql8_0),.clk(gclk));
	jdff dff_B_kPihtcfq0_0(.din(n1301),.dout(w_dff_B_kPihtcfq0_0),.clk(gclk));
	jdff dff_B_MJjWQueo0_0(.din(w_dff_B_kPihtcfq0_0),.dout(w_dff_B_MJjWQueo0_0),.clk(gclk));
	jdff dff_B_7gBuS4RL1_0(.din(w_dff_B_MJjWQueo0_0),.dout(w_dff_B_7gBuS4RL1_0),.clk(gclk));
	jdff dff_B_nXjjKyHT1_0(.din(w_dff_B_7gBuS4RL1_0),.dout(w_dff_B_nXjjKyHT1_0),.clk(gclk));
	jdff dff_B_uZHh1tCw2_0(.din(w_dff_B_nXjjKyHT1_0),.dout(w_dff_B_uZHh1tCw2_0),.clk(gclk));
	jdff dff_B_fNoYMSYB2_0(.din(w_dff_B_uZHh1tCw2_0),.dout(w_dff_B_fNoYMSYB2_0),.clk(gclk));
	jdff dff_B_tNelqQ8X3_0(.din(w_dff_B_fNoYMSYB2_0),.dout(w_dff_B_tNelqQ8X3_0),.clk(gclk));
	jdff dff_B_P5L4WvUp8_0(.din(w_dff_B_tNelqQ8X3_0),.dout(w_dff_B_P5L4WvUp8_0),.clk(gclk));
	jdff dff_B_U6ciIMBv3_0(.din(w_dff_B_P5L4WvUp8_0),.dout(w_dff_B_U6ciIMBv3_0),.clk(gclk));
	jdff dff_B_evhXXUnD4_0(.din(w_dff_B_U6ciIMBv3_0),.dout(w_dff_B_evhXXUnD4_0),.clk(gclk));
	jdff dff_B_ZQzU5vwe6_0(.din(w_dff_B_evhXXUnD4_0),.dout(w_dff_B_ZQzU5vwe6_0),.clk(gclk));
	jdff dff_B_k97cFn8n1_0(.din(w_dff_B_ZQzU5vwe6_0),.dout(w_dff_B_k97cFn8n1_0),.clk(gclk));
	jdff dff_B_QzoUBXs07_0(.din(w_dff_B_k97cFn8n1_0),.dout(w_dff_B_QzoUBXs07_0),.clk(gclk));
	jdff dff_B_rCYqDyRv0_0(.din(w_dff_B_QzoUBXs07_0),.dout(w_dff_B_rCYqDyRv0_0),.clk(gclk));
	jdff dff_B_uh6p67i63_0(.din(w_dff_B_rCYqDyRv0_0),.dout(w_dff_B_uh6p67i63_0),.clk(gclk));
	jdff dff_B_yNQ5VDmC3_0(.din(w_dff_B_uh6p67i63_0),.dout(w_dff_B_yNQ5VDmC3_0),.clk(gclk));
	jdff dff_A_cDTlSNpc6_0(.dout(w_n988_2[0]),.din(w_dff_A_cDTlSNpc6_0),.clk(gclk));
	jdff dff_A_FloPqlkm3_1(.dout(w_n988_2[1]),.din(w_dff_A_FloPqlkm3_1),.clk(gclk));
	jdff dff_B_zBPvyyCS1_0(.din(n1309),.dout(w_dff_B_zBPvyyCS1_0),.clk(gclk));
	jdff dff_B_jlFY93gi6_0(.din(w_dff_B_zBPvyyCS1_0),.dout(w_dff_B_jlFY93gi6_0),.clk(gclk));
	jdff dff_B_k0rNrJ1c2_0(.din(w_dff_B_jlFY93gi6_0),.dout(w_dff_B_k0rNrJ1c2_0),.clk(gclk));
	jdff dff_B_4TKULP6y5_0(.din(w_dff_B_k0rNrJ1c2_0),.dout(w_dff_B_4TKULP6y5_0),.clk(gclk));
	jdff dff_B_2WrTKrlo8_0(.din(w_dff_B_4TKULP6y5_0),.dout(w_dff_B_2WrTKrlo8_0),.clk(gclk));
	jdff dff_B_kl7zVGTp8_0(.din(w_dff_B_2WrTKrlo8_0),.dout(w_dff_B_kl7zVGTp8_0),.clk(gclk));
	jdff dff_B_YQ8XrtVg8_0(.din(w_dff_B_kl7zVGTp8_0),.dout(w_dff_B_YQ8XrtVg8_0),.clk(gclk));
	jdff dff_B_gjucRhre0_0(.din(w_dff_B_YQ8XrtVg8_0),.dout(w_dff_B_gjucRhre0_0),.clk(gclk));
	jdff dff_B_8J3MSDqz3_0(.din(w_dff_B_gjucRhre0_0),.dout(w_dff_B_8J3MSDqz3_0),.clk(gclk));
	jdff dff_B_aTGJZAjK2_0(.din(w_dff_B_8J3MSDqz3_0),.dout(w_dff_B_aTGJZAjK2_0),.clk(gclk));
	jdff dff_B_nhHj1Imt5_0(.din(w_dff_B_aTGJZAjK2_0),.dout(w_dff_B_nhHj1Imt5_0),.clk(gclk));
	jdff dff_B_JvpRnzoU2_0(.din(w_dff_B_nhHj1Imt5_0),.dout(w_dff_B_JvpRnzoU2_0),.clk(gclk));
	jdff dff_B_4dMPYloV4_0(.din(w_dff_B_JvpRnzoU2_0),.dout(w_dff_B_4dMPYloV4_0),.clk(gclk));
	jdff dff_B_U5aV58BB3_0(.din(w_dff_B_4dMPYloV4_0),.dout(w_dff_B_U5aV58BB3_0),.clk(gclk));
	jdff dff_B_p4k3zeD80_0(.din(w_dff_B_U5aV58BB3_0),.dout(w_dff_B_p4k3zeD80_0),.clk(gclk));
	jdff dff_B_m67jEMao4_0(.din(w_dff_B_p4k3zeD80_0),.dout(w_dff_B_m67jEMao4_0),.clk(gclk));
	jdff dff_B_2MPKNbl66_0(.din(w_dff_B_m67jEMao4_0),.dout(w_dff_B_2MPKNbl66_0),.clk(gclk));
	jdff dff_A_qJgKLL8u9_0(.dout(w_G137_5[0]),.din(w_dff_A_qJgKLL8u9_0),.clk(gclk));
	jdff dff_B_XJpeDObO3_0(.din(n1317),.dout(w_dff_B_XJpeDObO3_0),.clk(gclk));
	jdff dff_B_cL2PpUl82_0(.din(w_dff_B_XJpeDObO3_0),.dout(w_dff_B_cL2PpUl82_0),.clk(gclk));
	jdff dff_B_qb506v3Z0_0(.din(w_dff_B_cL2PpUl82_0),.dout(w_dff_B_qb506v3Z0_0),.clk(gclk));
	jdff dff_B_eRsD4t8b1_0(.din(w_dff_B_qb506v3Z0_0),.dout(w_dff_B_eRsD4t8b1_0),.clk(gclk));
	jdff dff_B_jAwzG7nk6_0(.din(w_dff_B_eRsD4t8b1_0),.dout(w_dff_B_jAwzG7nk6_0),.clk(gclk));
	jdff dff_B_9rJZOjZh9_0(.din(w_dff_B_jAwzG7nk6_0),.dout(w_dff_B_9rJZOjZh9_0),.clk(gclk));
	jdff dff_B_n1AFnr4Q8_0(.din(w_dff_B_9rJZOjZh9_0),.dout(w_dff_B_n1AFnr4Q8_0),.clk(gclk));
	jdff dff_B_uV5UYMyO3_0(.din(w_dff_B_n1AFnr4Q8_0),.dout(w_dff_B_uV5UYMyO3_0),.clk(gclk));
	jdff dff_B_zeMpWe9z5_0(.din(w_dff_B_uV5UYMyO3_0),.dout(w_dff_B_zeMpWe9z5_0),.clk(gclk));
	jdff dff_B_vrDX8wic6_0(.din(w_dff_B_zeMpWe9z5_0),.dout(w_dff_B_vrDX8wic6_0),.clk(gclk));
	jdff dff_B_r4UYfseN6_0(.din(w_dff_B_vrDX8wic6_0),.dout(w_dff_B_r4UYfseN6_0),.clk(gclk));
	jdff dff_B_PVzfH2SY9_0(.din(w_dff_B_r4UYfseN6_0),.dout(w_dff_B_PVzfH2SY9_0),.clk(gclk));
	jdff dff_B_4AVRx9sL0_0(.din(w_dff_B_PVzfH2SY9_0),.dout(w_dff_B_4AVRx9sL0_0),.clk(gclk));
	jdff dff_B_BnKnPaLt8_0(.din(w_dff_B_4AVRx9sL0_0),.dout(w_dff_B_BnKnPaLt8_0),.clk(gclk));
	jdff dff_B_Mup6Tlwp7_0(.din(w_dff_B_BnKnPaLt8_0),.dout(w_dff_B_Mup6Tlwp7_0),.clk(gclk));
	jdff dff_B_5SouL8NG9_0(.din(n1182),.dout(w_dff_B_5SouL8NG9_0),.clk(gclk));
	jdff dff_B_NYlbQWSk9_0(.din(w_dff_B_5SouL8NG9_0),.dout(w_dff_B_NYlbQWSk9_0),.clk(gclk));
	jdff dff_B_NCa3gi3n0_0(.din(w_dff_B_NYlbQWSk9_0),.dout(w_dff_B_NCa3gi3n0_0),.clk(gclk));
	jdff dff_B_AI5BY90G9_0(.din(w_dff_B_NCa3gi3n0_0),.dout(w_dff_B_AI5BY90G9_0),.clk(gclk));
	jdff dff_B_ZJieQwOd0_0(.din(w_dff_B_AI5BY90G9_0),.dout(w_dff_B_ZJieQwOd0_0),.clk(gclk));
	jdff dff_B_kYWpZLDo2_0(.din(w_dff_B_ZJieQwOd0_0),.dout(w_dff_B_kYWpZLDo2_0),.clk(gclk));
	jdff dff_B_gjvM1czA5_0(.din(w_dff_B_kYWpZLDo2_0),.dout(w_dff_B_gjvM1czA5_0),.clk(gclk));
	jdff dff_B_klsYbLLS0_0(.din(w_dff_B_gjvM1czA5_0),.dout(w_dff_B_klsYbLLS0_0),.clk(gclk));
	jdff dff_B_8UP3HyQ55_0(.din(w_dff_B_klsYbLLS0_0),.dout(w_dff_B_8UP3HyQ55_0),.clk(gclk));
	jdff dff_B_8p6gElg63_0(.din(n1325),.dout(w_dff_B_8p6gElg63_0),.clk(gclk));
	jdff dff_B_4P8f9Ny66_0(.din(w_dff_B_8p6gElg63_0),.dout(w_dff_B_4P8f9Ny66_0),.clk(gclk));
	jdff dff_B_jYHSEWlK0_0(.din(w_dff_B_4P8f9Ny66_0),.dout(w_dff_B_jYHSEWlK0_0),.clk(gclk));
	jdff dff_B_9CvpiysM6_0(.din(w_dff_B_jYHSEWlK0_0),.dout(w_dff_B_9CvpiysM6_0),.clk(gclk));
	jdff dff_B_TsASmaCN8_0(.din(w_dff_B_9CvpiysM6_0),.dout(w_dff_B_TsASmaCN8_0),.clk(gclk));
	jdff dff_B_qE1TCVdM7_0(.din(w_dff_B_TsASmaCN8_0),.dout(w_dff_B_qE1TCVdM7_0),.clk(gclk));
	jdff dff_B_6ISH0d4T1_0(.din(w_dff_B_qE1TCVdM7_0),.dout(w_dff_B_6ISH0d4T1_0),.clk(gclk));
	jdff dff_B_gGCs0xl34_0(.din(w_dff_B_6ISH0d4T1_0),.dout(w_dff_B_gGCs0xl34_0),.clk(gclk));
	jdff dff_B_8chnMslM1_0(.din(w_dff_B_gGCs0xl34_0),.dout(w_dff_B_8chnMslM1_0),.clk(gclk));
	jdff dff_B_zoiRCATK0_0(.din(w_dff_B_8chnMslM1_0),.dout(w_dff_B_zoiRCATK0_0),.clk(gclk));
	jdff dff_B_2cVd1BrQ8_0(.din(w_dff_B_zoiRCATK0_0),.dout(w_dff_B_2cVd1BrQ8_0),.clk(gclk));
	jdff dff_B_plECz23Q3_0(.din(w_dff_B_2cVd1BrQ8_0),.dout(w_dff_B_plECz23Q3_0),.clk(gclk));
	jdff dff_B_FwmdaOID9_0(.din(w_dff_B_plECz23Q3_0),.dout(w_dff_B_FwmdaOID9_0),.clk(gclk));
	jdff dff_B_RKNmEgFa5_0(.din(w_dff_B_FwmdaOID9_0),.dout(w_dff_B_RKNmEgFa5_0),.clk(gclk));
	jdff dff_B_EPlXEoKE7_0(.din(w_dff_B_RKNmEgFa5_0),.dout(w_dff_B_EPlXEoKE7_0),.clk(gclk));
	jdff dff_B_fyySlzZz8_0(.din(w_dff_B_EPlXEoKE7_0),.dout(w_dff_B_fyySlzZz8_0),.clk(gclk));
	jdff dff_B_Gc2x3gDv4_0(.din(n1175),.dout(w_dff_B_Gc2x3gDv4_0),.clk(gclk));
	jdff dff_B_rv5iWwR70_0(.din(w_dff_B_Gc2x3gDv4_0),.dout(w_dff_B_rv5iWwR70_0),.clk(gclk));
	jdff dff_B_Q2jbklSd2_0(.din(w_dff_B_rv5iWwR70_0),.dout(w_dff_B_Q2jbklSd2_0),.clk(gclk));
	jdff dff_B_FmE9Q68m8_0(.din(w_dff_B_Q2jbklSd2_0),.dout(w_dff_B_FmE9Q68m8_0),.clk(gclk));
	jdff dff_B_8UL0vcXR7_0(.din(w_dff_B_FmE9Q68m8_0),.dout(w_dff_B_8UL0vcXR7_0),.clk(gclk));
	jdff dff_B_GQE5kjLi0_0(.din(w_dff_B_8UL0vcXR7_0),.dout(w_dff_B_GQE5kjLi0_0),.clk(gclk));
	jdff dff_B_y0ZNfa0L1_0(.din(w_dff_B_GQE5kjLi0_0),.dout(w_dff_B_y0ZNfa0L1_0),.clk(gclk));
	jdff dff_B_ilB1twKe4_0(.din(w_dff_B_y0ZNfa0L1_0),.dout(w_dff_B_ilB1twKe4_0),.clk(gclk));
	jdff dff_B_aB83t4lO5_0(.din(w_dff_B_ilB1twKe4_0),.dout(w_dff_B_aB83t4lO5_0),.clk(gclk));
	jdff dff_B_h7shaPp49_0(.din(w_dff_B_aB83t4lO5_0),.dout(w_dff_B_h7shaPp49_0),.clk(gclk));
	jdff dff_A_bR1HbHEC2_1(.dout(w_n971_0[1]),.din(w_dff_A_bR1HbHEC2_1),.clk(gclk));
	jdff dff_B_Md8tmAYG5_1(.din(n967),.dout(w_dff_B_Md8tmAYG5_1),.clk(gclk));
	jdff dff_B_JEw2LQZI4_1(.din(w_dff_B_Md8tmAYG5_1),.dout(w_dff_B_JEw2LQZI4_1),.clk(gclk));
	jdff dff_B_3XOpD3QT0_1(.din(w_dff_B_JEw2LQZI4_1),.dout(w_dff_B_3XOpD3QT0_1),.clk(gclk));
	jdff dff_B_regfi3Nb9_1(.din(w_dff_B_3XOpD3QT0_1),.dout(w_dff_B_regfi3Nb9_1),.clk(gclk));
	jdff dff_B_ulL4W7kF5_1(.din(w_dff_B_regfi3Nb9_1),.dout(w_dff_B_ulL4W7kF5_1),.clk(gclk));
	jdff dff_B_jtnHOeD41_1(.din(w_dff_B_ulL4W7kF5_1),.dout(w_dff_B_jtnHOeD41_1),.clk(gclk));
	jdff dff_B_GMeH9Gjj8_1(.din(w_dff_B_jtnHOeD41_1),.dout(w_dff_B_GMeH9Gjj8_1),.clk(gclk));
	jdff dff_B_rDtJ97Wr4_1(.din(w_dff_B_GMeH9Gjj8_1),.dout(w_dff_B_rDtJ97Wr4_1),.clk(gclk));
	jdff dff_B_NchFnFQt8_1(.din(w_dff_B_rDtJ97Wr4_1),.dout(w_dff_B_NchFnFQt8_1),.clk(gclk));
	jdff dff_B_0Kif5Asu6_1(.din(w_dff_B_NchFnFQt8_1),.dout(w_dff_B_0Kif5Asu6_1),.clk(gclk));
	jdff dff_B_ax1g88iu3_0(.din(n1333),.dout(w_dff_B_ax1g88iu3_0),.clk(gclk));
	jdff dff_B_K9lTEUfB1_0(.din(w_dff_B_ax1g88iu3_0),.dout(w_dff_B_K9lTEUfB1_0),.clk(gclk));
	jdff dff_B_tgkvf8EM9_0(.din(w_dff_B_K9lTEUfB1_0),.dout(w_dff_B_tgkvf8EM9_0),.clk(gclk));
	jdff dff_B_73hCfHj40_0(.din(w_dff_B_tgkvf8EM9_0),.dout(w_dff_B_73hCfHj40_0),.clk(gclk));
	jdff dff_B_LhRFzZDx7_0(.din(w_dff_B_73hCfHj40_0),.dout(w_dff_B_LhRFzZDx7_0),.clk(gclk));
	jdff dff_B_8SbfsnlG3_0(.din(w_dff_B_LhRFzZDx7_0),.dout(w_dff_B_8SbfsnlG3_0),.clk(gclk));
	jdff dff_B_DMvDLERm5_0(.din(w_dff_B_8SbfsnlG3_0),.dout(w_dff_B_DMvDLERm5_0),.clk(gclk));
	jdff dff_B_LfujWgXt4_0(.din(w_dff_B_DMvDLERm5_0),.dout(w_dff_B_LfujWgXt4_0),.clk(gclk));
	jdff dff_B_AfdXMorj6_0(.din(w_dff_B_LfujWgXt4_0),.dout(w_dff_B_AfdXMorj6_0),.clk(gclk));
	jdff dff_B_EMQrR9uk0_0(.din(w_dff_B_AfdXMorj6_0),.dout(w_dff_B_EMQrR9uk0_0),.clk(gclk));
	jdff dff_B_AasOB3Pe0_0(.din(w_dff_B_EMQrR9uk0_0),.dout(w_dff_B_AasOB3Pe0_0),.clk(gclk));
	jdff dff_B_TBQjZteW8_0(.din(w_dff_B_AasOB3Pe0_0),.dout(w_dff_B_TBQjZteW8_0),.clk(gclk));
	jdff dff_B_7f7NxTVv0_0(.din(w_dff_B_TBQjZteW8_0),.dout(w_dff_B_7f7NxTVv0_0),.clk(gclk));
	jdff dff_B_sobignSw7_0(.din(w_dff_B_7f7NxTVv0_0),.dout(w_dff_B_sobignSw7_0),.clk(gclk));
	jdff dff_B_TNP94jqn5_0(.din(w_dff_B_sobignSw7_0),.dout(w_dff_B_TNP94jqn5_0),.clk(gclk));
	jdff dff_B_7nkid9JF1_0(.din(w_dff_B_TNP94jqn5_0),.dout(w_dff_B_7nkid9JF1_0),.clk(gclk));
	jdff dff_B_msqNHctB7_0(.din(n1169),.dout(w_dff_B_msqNHctB7_0),.clk(gclk));
	jdff dff_B_KVGJjC7d6_0(.din(w_dff_B_msqNHctB7_0),.dout(w_dff_B_KVGJjC7d6_0),.clk(gclk));
	jdff dff_B_07dPEegx8_0(.din(w_dff_B_KVGJjC7d6_0),.dout(w_dff_B_07dPEegx8_0),.clk(gclk));
	jdff dff_B_STWy7eZy0_0(.din(w_dff_B_07dPEegx8_0),.dout(w_dff_B_STWy7eZy0_0),.clk(gclk));
	jdff dff_B_zDvnauw57_0(.din(w_dff_B_STWy7eZy0_0),.dout(w_dff_B_zDvnauw57_0),.clk(gclk));
	jdff dff_B_M8A39Fs55_0(.din(w_dff_B_zDvnauw57_0),.dout(w_dff_B_M8A39Fs55_0),.clk(gclk));
	jdff dff_B_ubpiBd992_0(.din(w_dff_B_M8A39Fs55_0),.dout(w_dff_B_ubpiBd992_0),.clk(gclk));
	jdff dff_B_hQaZzNId4_0(.din(w_dff_B_ubpiBd992_0),.dout(w_dff_B_hQaZzNId4_0),.clk(gclk));
	jdff dff_B_uZmqZvfC6_0(.din(w_dff_B_hQaZzNId4_0),.dout(w_dff_B_uZmqZvfC6_0),.clk(gclk));
	jdff dff_B_b1F8kxF96_0(.din(w_dff_B_uZmqZvfC6_0),.dout(w_dff_B_b1F8kxF96_0),.clk(gclk));
	jdff dff_B_7Ql7B85O2_0(.din(w_dff_B_b1F8kxF96_0),.dout(w_dff_B_7Ql7B85O2_0),.clk(gclk));
	jdff dff_A_qKPaqswS4_0(.dout(w_n1002_2[0]),.din(w_dff_A_qKPaqswS4_0),.clk(gclk));
	jdff dff_A_oWjaihkA6_1(.dout(w_n1002_2[1]),.din(w_dff_A_oWjaihkA6_1),.clk(gclk));
	jdff dff_A_jocxXTXK8_0(.dout(w_G137_4[0]),.din(w_dff_A_jocxXTXK8_0),.clk(gclk));
	jdff dff_A_QabQwMds8_1(.dout(w_G137_4[1]),.din(w_dff_A_QabQwMds8_1),.clk(gclk));
	jdff dff_A_GlLFU3d46_0(.dout(w_G137_1[0]),.din(w_dff_A_GlLFU3d46_0),.clk(gclk));
	jdff dff_A_GWW1Se4x3_0(.dout(w_dff_A_GlLFU3d46_0),.din(w_dff_A_GWW1Se4x3_0),.clk(gclk));
	jdff dff_A_CwvoGdPP4_0(.dout(w_dff_A_GWW1Se4x3_0),.din(w_dff_A_CwvoGdPP4_0),.clk(gclk));
	jdff dff_A_DVMP496W0_0(.dout(w_dff_A_CwvoGdPP4_0),.din(w_dff_A_DVMP496W0_0),.clk(gclk));
	jdff dff_A_iq7Ngik62_0(.dout(w_dff_A_DVMP496W0_0),.din(w_dff_A_iq7Ngik62_0),.clk(gclk));
	jdff dff_A_7iSlBHLh0_1(.dout(w_G137_1[1]),.din(w_dff_A_7iSlBHLh0_1),.clk(gclk));
	jdff dff_A_FmSL0BLO9_1(.dout(w_dff_A_7iSlBHLh0_1),.din(w_dff_A_FmSL0BLO9_1),.clk(gclk));
	jdff dff_A_hGgPQXpz4_1(.dout(w_dff_A_FmSL0BLO9_1),.din(w_dff_A_hGgPQXpz4_1),.clk(gclk));
	jdff dff_A_W4dugbOG9_1(.dout(w_dff_A_hGgPQXpz4_1),.din(w_dff_A_W4dugbOG9_1),.clk(gclk));
	jdff dff_A_PtzTfacB8_1(.dout(w_dff_A_W4dugbOG9_1),.din(w_dff_A_PtzTfacB8_1),.clk(gclk));
	jdff dff_A_UZnqtXha6_1(.dout(w_dff_A_PtzTfacB8_1),.din(w_dff_A_UZnqtXha6_1),.clk(gclk));
	jdff dff_B_ztWMvnCi3_0(.din(n1341),.dout(w_dff_B_ztWMvnCi3_0),.clk(gclk));
	jdff dff_B_i9BkSOeO2_0(.din(w_dff_B_ztWMvnCi3_0),.dout(w_dff_B_i9BkSOeO2_0),.clk(gclk));
	jdff dff_B_K6lqkOYs0_0(.din(w_dff_B_i9BkSOeO2_0),.dout(w_dff_B_K6lqkOYs0_0),.clk(gclk));
	jdff dff_B_wtCgTdzf5_0(.din(w_dff_B_K6lqkOYs0_0),.dout(w_dff_B_wtCgTdzf5_0),.clk(gclk));
	jdff dff_B_x24JaxCH9_0(.din(w_dff_B_wtCgTdzf5_0),.dout(w_dff_B_x24JaxCH9_0),.clk(gclk));
	jdff dff_B_c0flpRF76_0(.din(w_dff_B_x24JaxCH9_0),.dout(w_dff_B_c0flpRF76_0),.clk(gclk));
	jdff dff_B_BEpWc7Ml2_0(.din(w_dff_B_c0flpRF76_0),.dout(w_dff_B_BEpWc7Ml2_0),.clk(gclk));
	jdff dff_B_CL9tZ6D97_0(.din(w_dff_B_BEpWc7Ml2_0),.dout(w_dff_B_CL9tZ6D97_0),.clk(gclk));
	jdff dff_B_yXl9WjRb8_0(.din(w_dff_B_CL9tZ6D97_0),.dout(w_dff_B_yXl9WjRb8_0),.clk(gclk));
	jdff dff_B_lAWTE3J57_0(.din(w_dff_B_yXl9WjRb8_0),.dout(w_dff_B_lAWTE3J57_0),.clk(gclk));
	jdff dff_B_C9oS9cZS5_0(.din(w_dff_B_lAWTE3J57_0),.dout(w_dff_B_C9oS9cZS5_0),.clk(gclk));
	jdff dff_B_7JEv4aTO8_0(.din(w_dff_B_C9oS9cZS5_0),.dout(w_dff_B_7JEv4aTO8_0),.clk(gclk));
	jdff dff_B_myWQJ2y58_0(.din(w_dff_B_7JEv4aTO8_0),.dout(w_dff_B_myWQJ2y58_0),.clk(gclk));
	jdff dff_B_ailZ8pec2_0(.din(w_dff_B_myWQJ2y58_0),.dout(w_dff_B_ailZ8pec2_0),.clk(gclk));
	jdff dff_B_QcyVKDaF5_0(.din(w_dff_B_ailZ8pec2_0),.dout(w_dff_B_QcyVKDaF5_0),.clk(gclk));
	jdff dff_B_UkYxzIAK4_0(.din(w_dff_B_QcyVKDaF5_0),.dout(w_dff_B_UkYxzIAK4_0),.clk(gclk));
	jdff dff_B_Ll5YcClR3_0(.din(w_dff_B_UkYxzIAK4_0),.dout(w_dff_B_Ll5YcClR3_0),.clk(gclk));
	jdff dff_B_1wGWBeyi0_0(.din(n1162),.dout(w_dff_B_1wGWBeyi0_0),.clk(gclk));
	jdff dff_B_6102vNKn3_0(.din(w_dff_B_1wGWBeyi0_0),.dout(w_dff_B_6102vNKn3_0),.clk(gclk));
	jdff dff_B_javK3lxR8_0(.din(w_dff_B_6102vNKn3_0),.dout(w_dff_B_javK3lxR8_0),.clk(gclk));
	jdff dff_B_0OJJpXqw0_0(.din(w_dff_B_javK3lxR8_0),.dout(w_dff_B_0OJJpXqw0_0),.clk(gclk));
	jdff dff_B_WIsIyD9v8_0(.din(w_dff_B_0OJJpXqw0_0),.dout(w_dff_B_WIsIyD9v8_0),.clk(gclk));
	jdff dff_B_jsCtqBh03_0(.din(w_dff_B_WIsIyD9v8_0),.dout(w_dff_B_jsCtqBh03_0),.clk(gclk));
	jdff dff_B_VnT4vukm2_0(.din(w_dff_B_jsCtqBh03_0),.dout(w_dff_B_VnT4vukm2_0),.clk(gclk));
	jdff dff_B_BNbcHZR40_0(.din(w_dff_B_VnT4vukm2_0),.dout(w_dff_B_BNbcHZR40_0),.clk(gclk));
	jdff dff_B_2z7KQv9V0_0(.din(w_dff_B_BNbcHZR40_0),.dout(w_dff_B_2z7KQv9V0_0),.clk(gclk));
	jdff dff_B_WfaJa27F4_0(.din(w_dff_B_2z7KQv9V0_0),.dout(w_dff_B_WfaJa27F4_0),.clk(gclk));
	jdff dff_B_80mx3hGy4_0(.din(w_dff_B_WfaJa27F4_0),.dout(w_dff_B_80mx3hGy4_0),.clk(gclk));
	jdff dff_B_3RTyat0o0_0(.din(w_dff_B_80mx3hGy4_0),.dout(w_dff_B_3RTyat0o0_0),.clk(gclk));
	jdff dff_B_E5a09JiM7_0(.din(w_dff_B_3RTyat0o0_0),.dout(w_dff_B_E5a09JiM7_0),.clk(gclk));
	jdff dff_B_b8gTI8kT6_0(.din(n788),.dout(w_dff_B_b8gTI8kT6_0),.clk(gclk));
	jdff dff_B_jdigdjsC9_0(.din(n780),.dout(w_dff_B_jdigdjsC9_0),.clk(gclk));
	jdff dff_B_UKNgXBOI0_0(.din(w_dff_B_jdigdjsC9_0),.dout(w_dff_B_UKNgXBOI0_0),.clk(gclk));
	jdff dff_B_6RQQT2QQ7_0(.din(w_dff_B_UKNgXBOI0_0),.dout(w_dff_B_6RQQT2QQ7_0),.clk(gclk));
	jdff dff_A_9IVKEkEa9_0(.dout(w_n741_0[0]),.din(w_dff_A_9IVKEkEa9_0),.clk(gclk));
	jdff dff_A_ajFVRjMK4_0(.dout(w_dff_A_9IVKEkEa9_0),.din(w_dff_A_ajFVRjMK4_0),.clk(gclk));
	jdff dff_A_gHNU9yhO6_0(.dout(w_dff_A_ajFVRjMK4_0),.din(w_dff_A_gHNU9yhO6_0),.clk(gclk));
	jdff dff_A_bhsedOfo1_0(.dout(w_dff_A_gHNU9yhO6_0),.din(w_dff_A_bhsedOfo1_0),.clk(gclk));
	jdff dff_A_b5O4umPe7_0(.dout(w_dff_A_bhsedOfo1_0),.din(w_dff_A_b5O4umPe7_0),.clk(gclk));
	jdff dff_A_7VdwYuTi0_0(.dout(w_dff_A_b5O4umPe7_0),.din(w_dff_A_7VdwYuTi0_0),.clk(gclk));
	jdff dff_A_mdUzwDUP4_0(.dout(w_dff_A_7VdwYuTi0_0),.din(w_dff_A_mdUzwDUP4_0),.clk(gclk));
	jdff dff_B_USQKzslP9_1(.din(n1388),.dout(w_dff_B_USQKzslP9_1),.clk(gclk));
	jdff dff_B_KMgMnI7B3_1(.din(w_dff_B_USQKzslP9_1),.dout(w_dff_B_KMgMnI7B3_1),.clk(gclk));
	jdff dff_B_UnAVtBLJ5_1(.din(w_dff_B_KMgMnI7B3_1),.dout(w_dff_B_UnAVtBLJ5_1),.clk(gclk));
	jdff dff_B_jXurijec5_1(.din(w_dff_B_UnAVtBLJ5_1),.dout(w_dff_B_jXurijec5_1),.clk(gclk));
	jdff dff_B_Ujp1Wrmx9_1(.din(w_dff_B_jXurijec5_1),.dout(w_dff_B_Ujp1Wrmx9_1),.clk(gclk));
	jdff dff_B_LOmY5tsq4_1(.din(w_dff_B_Ujp1Wrmx9_1),.dout(w_dff_B_LOmY5tsq4_1),.clk(gclk));
	jdff dff_B_h9gUpSve0_1(.din(w_dff_B_LOmY5tsq4_1),.dout(w_dff_B_h9gUpSve0_1),.clk(gclk));
	jdff dff_B_70ZbSBTX3_1(.din(w_dff_B_h9gUpSve0_1),.dout(w_dff_B_70ZbSBTX3_1),.clk(gclk));
	jdff dff_B_HwQpfLCs0_1(.din(w_dff_B_70ZbSBTX3_1),.dout(w_dff_B_HwQpfLCs0_1),.clk(gclk));
	jdff dff_B_Wj5Eu4qw1_1(.din(w_dff_B_HwQpfLCs0_1),.dout(w_dff_B_Wj5Eu4qw1_1),.clk(gclk));
	jdff dff_B_kthcHHMA1_1(.din(w_dff_B_Wj5Eu4qw1_1),.dout(w_dff_B_kthcHHMA1_1),.clk(gclk));
	jdff dff_B_hPwYu4Mw4_1(.din(w_dff_B_kthcHHMA1_1),.dout(w_dff_B_hPwYu4Mw4_1),.clk(gclk));
	jdff dff_B_aIS0yRux6_1(.din(w_dff_B_hPwYu4Mw4_1),.dout(w_dff_B_aIS0yRux6_1),.clk(gclk));
	jdff dff_B_RO05wpNx0_1(.din(w_dff_B_aIS0yRux6_1),.dout(w_dff_B_RO05wpNx0_1),.clk(gclk));
	jdff dff_B_v3kV7VdB5_1(.din(w_dff_B_RO05wpNx0_1),.dout(w_dff_B_v3kV7VdB5_1),.clk(gclk));
	jdff dff_B_KP5xW9d20_1(.din(w_dff_B_v3kV7VdB5_1),.dout(w_dff_B_KP5xW9d20_1),.clk(gclk));
	jdff dff_B_swx7ICbF7_1(.din(w_dff_B_KP5xW9d20_1),.dout(w_dff_B_swx7ICbF7_1),.clk(gclk));
	jdff dff_B_KIBYLFHW4_1(.din(w_dff_B_swx7ICbF7_1),.dout(w_dff_B_KIBYLFHW4_1),.clk(gclk));
	jdff dff_B_EcgkE7Vz6_1(.din(w_dff_B_KIBYLFHW4_1),.dout(w_dff_B_EcgkE7Vz6_1),.clk(gclk));
	jdff dff_B_liJr58Gv3_1(.din(n1539),.dout(w_dff_B_liJr58Gv3_1),.clk(gclk));
	jdff dff_B_tOD8Gnln8_1(.din(w_dff_B_liJr58Gv3_1),.dout(w_dff_B_tOD8Gnln8_1),.clk(gclk));
	jdff dff_B_v8CpiGlj6_1(.din(w_dff_B_tOD8Gnln8_1),.dout(w_dff_B_v8CpiGlj6_1),.clk(gclk));
	jdff dff_B_AGoGd4HH0_1(.din(w_dff_B_v8CpiGlj6_1),.dout(w_dff_B_AGoGd4HH0_1),.clk(gclk));
	jdff dff_B_vu1PC1aU6_1(.din(w_dff_B_AGoGd4HH0_1),.dout(w_dff_B_vu1PC1aU6_1),.clk(gclk));
	jdff dff_B_d5C077gz9_1(.din(w_dff_B_vu1PC1aU6_1),.dout(w_dff_B_d5C077gz9_1),.clk(gclk));
	jdff dff_B_LeTPWCFM4_1(.din(w_dff_B_d5C077gz9_1),.dout(w_dff_B_LeTPWCFM4_1),.clk(gclk));
	jdff dff_B_fKpBDmCz7_1(.din(w_dff_B_LeTPWCFM4_1),.dout(w_dff_B_fKpBDmCz7_1),.clk(gclk));
	jdff dff_B_DeftKvjS2_1(.din(w_dff_B_fKpBDmCz7_1),.dout(w_dff_B_DeftKvjS2_1),.clk(gclk));
	jdff dff_B_bn9wfamB6_1(.din(w_dff_B_DeftKvjS2_1),.dout(w_dff_B_bn9wfamB6_1),.clk(gclk));
	jdff dff_B_6EXBxlqf7_1(.din(w_dff_B_bn9wfamB6_1),.dout(w_dff_B_6EXBxlqf7_1),.clk(gclk));
	jdff dff_B_6phi5lZD8_1(.din(w_dff_B_6EXBxlqf7_1),.dout(w_dff_B_6phi5lZD8_1),.clk(gclk));
	jdff dff_B_04OXJUHx2_1(.din(w_dff_B_6phi5lZD8_1),.dout(w_dff_B_04OXJUHx2_1),.clk(gclk));
	jdff dff_B_PZtoP8qq6_1(.din(w_dff_B_04OXJUHx2_1),.dout(w_dff_B_PZtoP8qq6_1),.clk(gclk));
	jdff dff_B_cMYxrKRs6_1(.din(w_dff_B_PZtoP8qq6_1),.dout(w_dff_B_cMYxrKRs6_1),.clk(gclk));
	jdff dff_B_rVQQE3yR9_1(.din(w_dff_B_cMYxrKRs6_1),.dout(w_dff_B_rVQQE3yR9_1),.clk(gclk));
	jdff dff_B_myWxgLJO3_1(.din(w_dff_B_rVQQE3yR9_1),.dout(w_dff_B_myWxgLJO3_1),.clk(gclk));
	jdff dff_B_IWjoElcz7_1(.din(w_dff_B_myWxgLJO3_1),.dout(w_dff_B_IWjoElcz7_1),.clk(gclk));
	jdff dff_B_aFV8wzDx3_1(.din(w_dff_B_IWjoElcz7_1),.dout(w_dff_B_aFV8wzDx3_1),.clk(gclk));
	jdff dff_B_15hlmeCz0_0(.din(n1614),.dout(w_dff_B_15hlmeCz0_0),.clk(gclk));
	jdff dff_B_Mqf5ubJI2_0(.din(w_dff_B_15hlmeCz0_0),.dout(w_dff_B_Mqf5ubJI2_0),.clk(gclk));
	jdff dff_B_mhDj21vY9_0(.din(w_dff_B_Mqf5ubJI2_0),.dout(w_dff_B_mhDj21vY9_0),.clk(gclk));
	jdff dff_B_gHqZyo5M7_0(.din(w_dff_B_mhDj21vY9_0),.dout(w_dff_B_gHqZyo5M7_0),.clk(gclk));
	jdff dff_B_6e6B1n8h3_0(.din(w_dff_B_gHqZyo5M7_0),.dout(w_dff_B_6e6B1n8h3_0),.clk(gclk));
	jdff dff_B_0QVzKUlI6_0(.din(w_dff_B_6e6B1n8h3_0),.dout(w_dff_B_0QVzKUlI6_0),.clk(gclk));
	jdff dff_B_A4W80aMP3_0(.din(w_dff_B_0QVzKUlI6_0),.dout(w_dff_B_A4W80aMP3_0),.clk(gclk));
	jdff dff_B_pUvIAmOp9_0(.din(w_dff_B_A4W80aMP3_0),.dout(w_dff_B_pUvIAmOp9_0),.clk(gclk));
	jdff dff_B_RZc1oA6Y5_0(.din(w_dff_B_pUvIAmOp9_0),.dout(w_dff_B_RZc1oA6Y5_0),.clk(gclk));
	jdff dff_B_HInz9TbG4_0(.din(w_dff_B_RZc1oA6Y5_0),.dout(w_dff_B_HInz9TbG4_0),.clk(gclk));
	jdff dff_B_HTo36Pef8_0(.din(w_dff_B_HInz9TbG4_0),.dout(w_dff_B_HTo36Pef8_0),.clk(gclk));
	jdff dff_B_TpL66Lr31_0(.din(w_dff_B_HTo36Pef8_0),.dout(w_dff_B_TpL66Lr31_0),.clk(gclk));
	jdff dff_B_ZyIjFXTA6_0(.din(w_dff_B_TpL66Lr31_0),.dout(w_dff_B_ZyIjFXTA6_0),.clk(gclk));
	jdff dff_B_qMi1Wg3H9_0(.din(w_dff_B_ZyIjFXTA6_0),.dout(w_dff_B_qMi1Wg3H9_0),.clk(gclk));
	jdff dff_B_sozDVgp64_0(.din(w_dff_B_qMi1Wg3H9_0),.dout(w_dff_B_sozDVgp64_0),.clk(gclk));
	jdff dff_B_2ckhzU1K5_0(.din(w_dff_B_sozDVgp64_0),.dout(w_dff_B_2ckhzU1K5_0),.clk(gclk));
	jdff dff_B_qd0F33eQ0_0(.din(w_dff_B_2ckhzU1K5_0),.dout(w_dff_B_qd0F33eQ0_0),.clk(gclk));
	jdff dff_B_3LrkiBDe3_0(.din(w_dff_B_qd0F33eQ0_0),.dout(w_dff_B_3LrkiBDe3_0),.clk(gclk));
	jdff dff_B_vgKwEqZe7_0(.din(w_dff_B_3LrkiBDe3_0),.dout(w_dff_B_vgKwEqZe7_0),.clk(gclk));
	jdff dff_A_BK9DTSEo1_1(.dout(w_n797_1[1]),.din(w_dff_A_BK9DTSEo1_1),.clk(gclk));
	jdff dff_A_XkEeD6U12_1(.dout(w_dff_A_BK9DTSEo1_1),.din(w_dff_A_XkEeD6U12_1),.clk(gclk));
	jdff dff_A_550Je7HB8_1(.dout(w_dff_A_XkEeD6U12_1),.din(w_dff_A_550Je7HB8_1),.clk(gclk));
	jdff dff_A_qSYZXzx47_1(.dout(w_dff_A_550Je7HB8_1),.din(w_dff_A_qSYZXzx47_1),.clk(gclk));
	jdff dff_A_erIcdBdF1_1(.dout(w_dff_A_qSYZXzx47_1),.din(w_dff_A_erIcdBdF1_1),.clk(gclk));
	jdff dff_A_xoV0igcO0_1(.dout(w_dff_A_erIcdBdF1_1),.din(w_dff_A_xoV0igcO0_1),.clk(gclk));
	jdff dff_A_1ncj9mPS5_1(.dout(w_dff_A_xoV0igcO0_1),.din(w_dff_A_1ncj9mPS5_1),.clk(gclk));
	jdff dff_A_IKqy2qAP1_1(.dout(w_dff_A_1ncj9mPS5_1),.din(w_dff_A_IKqy2qAP1_1),.clk(gclk));
	jdff dff_A_d56hPKNM7_1(.dout(w_dff_A_IKqy2qAP1_1),.din(w_dff_A_d56hPKNM7_1),.clk(gclk));
	jdff dff_A_cjfv5gIw6_1(.dout(w_dff_A_d56hPKNM7_1),.din(w_dff_A_cjfv5gIw6_1),.clk(gclk));
	jdff dff_A_bPPu9Tme4_1(.dout(w_dff_A_cjfv5gIw6_1),.din(w_dff_A_bPPu9Tme4_1),.clk(gclk));
	jdff dff_A_ymqvpjQT3_1(.dout(w_dff_A_bPPu9Tme4_1),.din(w_dff_A_ymqvpjQT3_1),.clk(gclk));
	jdff dff_A_A0CkILy93_1(.dout(w_dff_A_ymqvpjQT3_1),.din(w_dff_A_A0CkILy93_1),.clk(gclk));
	jdff dff_A_BXunqfwI6_1(.dout(w_dff_A_A0CkILy93_1),.din(w_dff_A_BXunqfwI6_1),.clk(gclk));
	jdff dff_A_ywngHWxn3_2(.dout(w_n797_1[2]),.din(w_dff_A_ywngHWxn3_2),.clk(gclk));
	jdff dff_A_lhgl286T7_2(.dout(w_dff_A_ywngHWxn3_2),.din(w_dff_A_lhgl286T7_2),.clk(gclk));
	jdff dff_A_j9Srvw5M9_2(.dout(w_dff_A_lhgl286T7_2),.din(w_dff_A_j9Srvw5M9_2),.clk(gclk));
	jdff dff_A_2j0g19Jd4_2(.dout(w_dff_A_j9Srvw5M9_2),.din(w_dff_A_2j0g19Jd4_2),.clk(gclk));
	jdff dff_A_KCpLv8PW7_2(.dout(w_dff_A_2j0g19Jd4_2),.din(w_dff_A_KCpLv8PW7_2),.clk(gclk));
	jdff dff_A_dxrN5TwR8_2(.dout(w_dff_A_KCpLv8PW7_2),.din(w_dff_A_dxrN5TwR8_2),.clk(gclk));
	jdff dff_A_DxVstlTq2_2(.dout(w_dff_A_dxrN5TwR8_2),.din(w_dff_A_DxVstlTq2_2),.clk(gclk));
	jdff dff_A_NBfNvf6M3_2(.dout(w_dff_A_DxVstlTq2_2),.din(w_dff_A_NBfNvf6M3_2),.clk(gclk));
	jdff dff_A_vZFeOSNe6_2(.dout(w_dff_A_NBfNvf6M3_2),.din(w_dff_A_vZFeOSNe6_2),.clk(gclk));
	jdff dff_A_o2tyTjap4_2(.dout(w_dff_A_vZFeOSNe6_2),.din(w_dff_A_o2tyTjap4_2),.clk(gclk));
	jdff dff_A_URiRgjP36_1(.dout(w_n797_0[1]),.din(w_dff_A_URiRgjP36_1),.clk(gclk));
	jdff dff_A_brXW6BiL6_1(.dout(w_dff_A_URiRgjP36_1),.din(w_dff_A_brXW6BiL6_1),.clk(gclk));
	jdff dff_A_syESiIjk9_1(.dout(w_dff_A_brXW6BiL6_1),.din(w_dff_A_syESiIjk9_1),.clk(gclk));
	jdff dff_A_7fLkCLQR7_1(.dout(w_dff_A_syESiIjk9_1),.din(w_dff_A_7fLkCLQR7_1),.clk(gclk));
	jdff dff_A_HqXYa5SV1_1(.dout(w_dff_A_7fLkCLQR7_1),.din(w_dff_A_HqXYa5SV1_1),.clk(gclk));
	jdff dff_A_kYvtkn6Q2_1(.dout(w_dff_A_HqXYa5SV1_1),.din(w_dff_A_kYvtkn6Q2_1),.clk(gclk));
	jdff dff_A_fAEBuU884_1(.dout(w_dff_A_kYvtkn6Q2_1),.din(w_dff_A_fAEBuU884_1),.clk(gclk));
	jdff dff_A_0gVQfX8d2_1(.dout(w_dff_A_fAEBuU884_1),.din(w_dff_A_0gVQfX8d2_1),.clk(gclk));
	jdff dff_A_wnyp9gVQ4_1(.dout(w_dff_A_0gVQfX8d2_1),.din(w_dff_A_wnyp9gVQ4_1),.clk(gclk));
	jdff dff_A_aH6KF7Li9_1(.dout(w_dff_A_wnyp9gVQ4_1),.din(w_dff_A_aH6KF7Li9_1),.clk(gclk));
	jdff dff_A_OTsvVIaB8_1(.dout(w_dff_A_aH6KF7Li9_1),.din(w_dff_A_OTsvVIaB8_1),.clk(gclk));
	jdff dff_A_GB2w0Nnn0_2(.dout(w_n797_0[2]),.din(w_dff_A_GB2w0Nnn0_2),.clk(gclk));
	jdff dff_B_r4tGmRXW1_3(.din(n797),.dout(w_dff_B_r4tGmRXW1_3),.clk(gclk));
	jdff dff_B_DQimDwlC9_3(.din(w_dff_B_r4tGmRXW1_3),.dout(w_dff_B_DQimDwlC9_3),.clk(gclk));
	jdff dff_B_NUKKHghL4_3(.din(w_dff_B_DQimDwlC9_3),.dout(w_dff_B_NUKKHghL4_3),.clk(gclk));
	jdff dff_B_zkAyo6es1_3(.din(w_dff_B_NUKKHghL4_3),.dout(w_dff_B_zkAyo6es1_3),.clk(gclk));
	jdff dff_B_yBgG9BUT3_3(.din(w_dff_B_zkAyo6es1_3),.dout(w_dff_B_yBgG9BUT3_3),.clk(gclk));
	jdff dff_B_YIZo3wIt3_3(.din(w_dff_B_yBgG9BUT3_3),.dout(w_dff_B_YIZo3wIt3_3),.clk(gclk));
	jdff dff_B_Cfafl5Uw9_0(.din(n1621),.dout(w_dff_B_Cfafl5Uw9_0),.clk(gclk));
	jdff dff_B_1D3tNEbH5_0(.din(w_dff_B_Cfafl5Uw9_0),.dout(w_dff_B_1D3tNEbH5_0),.clk(gclk));
	jdff dff_B_T25pqIU90_0(.din(w_dff_B_1D3tNEbH5_0),.dout(w_dff_B_T25pqIU90_0),.clk(gclk));
	jdff dff_B_e3Z69bgo0_0(.din(w_dff_B_T25pqIU90_0),.dout(w_dff_B_e3Z69bgo0_0),.clk(gclk));
	jdff dff_B_mi6ossYj6_0(.din(w_dff_B_e3Z69bgo0_0),.dout(w_dff_B_mi6ossYj6_0),.clk(gclk));
	jdff dff_B_M2eGyQQH9_0(.din(w_dff_B_mi6ossYj6_0),.dout(w_dff_B_M2eGyQQH9_0),.clk(gclk));
	jdff dff_B_crkvjXU33_0(.din(w_dff_B_M2eGyQQH9_0),.dout(w_dff_B_crkvjXU33_0),.clk(gclk));
	jdff dff_B_PXaCXsGn0_0(.din(w_dff_B_crkvjXU33_0),.dout(w_dff_B_PXaCXsGn0_0),.clk(gclk));
	jdff dff_B_Q96U06dn2_0(.din(w_dff_B_PXaCXsGn0_0),.dout(w_dff_B_Q96U06dn2_0),.clk(gclk));
	jdff dff_B_JwB8c2Id0_0(.din(w_dff_B_Q96U06dn2_0),.dout(w_dff_B_JwB8c2Id0_0),.clk(gclk));
	jdff dff_B_vsJHQTFH3_0(.din(w_dff_B_JwB8c2Id0_0),.dout(w_dff_B_vsJHQTFH3_0),.clk(gclk));
	jdff dff_B_rTmzJXWY9_0(.din(w_dff_B_vsJHQTFH3_0),.dout(w_dff_B_rTmzJXWY9_0),.clk(gclk));
	jdff dff_B_uz2v2gJP5_0(.din(w_dff_B_rTmzJXWY9_0),.dout(w_dff_B_uz2v2gJP5_0),.clk(gclk));
	jdff dff_B_Ki1C5p8s9_0(.din(w_dff_B_uz2v2gJP5_0),.dout(w_dff_B_Ki1C5p8s9_0),.clk(gclk));
	jdff dff_B_dtxE527h8_0(.din(w_dff_B_Ki1C5p8s9_0),.dout(w_dff_B_dtxE527h8_0),.clk(gclk));
	jdff dff_B_Dq1ziY9a4_0(.din(w_dff_B_dtxE527h8_0),.dout(w_dff_B_Dq1ziY9a4_0),.clk(gclk));
	jdff dff_B_WDVpWqM91_0(.din(w_dff_B_Dq1ziY9a4_0),.dout(w_dff_B_WDVpWqM91_0),.clk(gclk));
	jdff dff_B_U695gRXs2_0(.din(w_dff_B_WDVpWqM91_0),.dout(w_dff_B_U695gRXs2_0),.clk(gclk));
	jdff dff_B_e5vsVdSQ9_0(.din(w_dff_B_U695gRXs2_0),.dout(w_dff_B_e5vsVdSQ9_0),.clk(gclk));
	jdff dff_A_faJqbZCj9_1(.dout(w_n843_1[1]),.din(w_dff_A_faJqbZCj9_1),.clk(gclk));
	jdff dff_A_hDhfidel2_1(.dout(w_dff_A_faJqbZCj9_1),.din(w_dff_A_hDhfidel2_1),.clk(gclk));
	jdff dff_A_cd3zl5239_1(.dout(w_dff_A_hDhfidel2_1),.din(w_dff_A_cd3zl5239_1),.clk(gclk));
	jdff dff_A_wT0kuPVf2_1(.dout(w_dff_A_cd3zl5239_1),.din(w_dff_A_wT0kuPVf2_1),.clk(gclk));
	jdff dff_A_DdZi7buT0_1(.dout(w_dff_A_wT0kuPVf2_1),.din(w_dff_A_DdZi7buT0_1),.clk(gclk));
	jdff dff_A_Dt55PWry9_1(.dout(w_dff_A_DdZi7buT0_1),.din(w_dff_A_Dt55PWry9_1),.clk(gclk));
	jdff dff_A_CO8St1YS9_1(.dout(w_dff_A_Dt55PWry9_1),.din(w_dff_A_CO8St1YS9_1),.clk(gclk));
	jdff dff_A_m2S8yrAU7_1(.dout(w_dff_A_CO8St1YS9_1),.din(w_dff_A_m2S8yrAU7_1),.clk(gclk));
	jdff dff_A_JbvicfCw8_1(.dout(w_dff_A_m2S8yrAU7_1),.din(w_dff_A_JbvicfCw8_1),.clk(gclk));
	jdff dff_A_9UsFVfnC9_1(.dout(w_dff_A_JbvicfCw8_1),.din(w_dff_A_9UsFVfnC9_1),.clk(gclk));
	jdff dff_A_z0St6chz6_1(.dout(w_dff_A_9UsFVfnC9_1),.din(w_dff_A_z0St6chz6_1),.clk(gclk));
	jdff dff_A_gXaqboLV4_1(.dout(w_dff_A_z0St6chz6_1),.din(w_dff_A_gXaqboLV4_1),.clk(gclk));
	jdff dff_A_7D589fGb6_1(.dout(w_dff_A_gXaqboLV4_1),.din(w_dff_A_7D589fGb6_1),.clk(gclk));
	jdff dff_A_z7biw8aO7_1(.dout(w_dff_A_7D589fGb6_1),.din(w_dff_A_z7biw8aO7_1),.clk(gclk));
	jdff dff_A_kmdKYBFs7_2(.dout(w_n843_1[2]),.din(w_dff_A_kmdKYBFs7_2),.clk(gclk));
	jdff dff_A_NLfBXjRI9_2(.dout(w_dff_A_kmdKYBFs7_2),.din(w_dff_A_NLfBXjRI9_2),.clk(gclk));
	jdff dff_A_6BhN392g9_2(.dout(w_dff_A_NLfBXjRI9_2),.din(w_dff_A_6BhN392g9_2),.clk(gclk));
	jdff dff_A_tT0ww60T9_2(.dout(w_dff_A_6BhN392g9_2),.din(w_dff_A_tT0ww60T9_2),.clk(gclk));
	jdff dff_A_v1pKFrwK2_2(.dout(w_dff_A_tT0ww60T9_2),.din(w_dff_A_v1pKFrwK2_2),.clk(gclk));
	jdff dff_A_GhHJEumA4_2(.dout(w_dff_A_v1pKFrwK2_2),.din(w_dff_A_GhHJEumA4_2),.clk(gclk));
	jdff dff_A_HxdeZnw21_2(.dout(w_dff_A_GhHJEumA4_2),.din(w_dff_A_HxdeZnw21_2),.clk(gclk));
	jdff dff_A_s2EadMFx9_2(.dout(w_dff_A_HxdeZnw21_2),.din(w_dff_A_s2EadMFx9_2),.clk(gclk));
	jdff dff_A_AtRqkxFK9_2(.dout(w_dff_A_s2EadMFx9_2),.din(w_dff_A_AtRqkxFK9_2),.clk(gclk));
	jdff dff_A_O4GArnQ14_2(.dout(w_dff_A_AtRqkxFK9_2),.din(w_dff_A_O4GArnQ14_2),.clk(gclk));
	jdff dff_A_h7NcRlSa2_1(.dout(w_n843_0[1]),.din(w_dff_A_h7NcRlSa2_1),.clk(gclk));
	jdff dff_A_0CI0HYfu6_1(.dout(w_dff_A_h7NcRlSa2_1),.din(w_dff_A_0CI0HYfu6_1),.clk(gclk));
	jdff dff_A_7qNmDIMF2_1(.dout(w_dff_A_0CI0HYfu6_1),.din(w_dff_A_7qNmDIMF2_1),.clk(gclk));
	jdff dff_A_lTT1lmQx8_1(.dout(w_dff_A_7qNmDIMF2_1),.din(w_dff_A_lTT1lmQx8_1),.clk(gclk));
	jdff dff_A_Lm2jK0k00_1(.dout(w_dff_A_lTT1lmQx8_1),.din(w_dff_A_Lm2jK0k00_1),.clk(gclk));
	jdff dff_A_k3Mg6Bdz5_1(.dout(w_dff_A_Lm2jK0k00_1),.din(w_dff_A_k3Mg6Bdz5_1),.clk(gclk));
	jdff dff_A_426JwAvx2_1(.dout(w_dff_A_k3Mg6Bdz5_1),.din(w_dff_A_426JwAvx2_1),.clk(gclk));
	jdff dff_A_tdIr1GZD7_1(.dout(w_dff_A_426JwAvx2_1),.din(w_dff_A_tdIr1GZD7_1),.clk(gclk));
	jdff dff_A_fW4zbuyv3_1(.dout(w_dff_A_tdIr1GZD7_1),.din(w_dff_A_fW4zbuyv3_1),.clk(gclk));
	jdff dff_A_2nYDDVP93_1(.dout(w_dff_A_fW4zbuyv3_1),.din(w_dff_A_2nYDDVP93_1),.clk(gclk));
	jdff dff_A_0idNOgO82_1(.dout(w_dff_A_2nYDDVP93_1),.din(w_dff_A_0idNOgO82_1),.clk(gclk));
	jdff dff_A_mxYrmpWq2_2(.dout(w_n843_0[2]),.din(w_dff_A_mxYrmpWq2_2),.clk(gclk));
	jdff dff_B_yKeoj2Oi7_3(.din(n843),.dout(w_dff_B_yKeoj2Oi7_3),.clk(gclk));
	jdff dff_B_rcgxDbXG3_3(.din(w_dff_B_yKeoj2Oi7_3),.dout(w_dff_B_rcgxDbXG3_3),.clk(gclk));
	jdff dff_B_30fadAIL9_3(.din(w_dff_B_rcgxDbXG3_3),.dout(w_dff_B_30fadAIL9_3),.clk(gclk));
	jdff dff_B_4vRaUZrI7_3(.din(w_dff_B_30fadAIL9_3),.dout(w_dff_B_4vRaUZrI7_3),.clk(gclk));
	jdff dff_B_qIwBJaZA5_3(.din(w_dff_B_4vRaUZrI7_3),.dout(w_dff_B_qIwBJaZA5_3),.clk(gclk));
	jdff dff_B_nbEnGORg5_3(.din(w_dff_B_qIwBJaZA5_3),.dout(w_dff_B_nbEnGORg5_3),.clk(gclk));
	jdff dff_B_Xoebksbe1_1(.din(n1626),.dout(w_dff_B_Xoebksbe1_1),.clk(gclk));
	jdff dff_B_mXHIPi7r6_0(.din(n1637),.dout(w_dff_B_mXHIPi7r6_0),.clk(gclk));
	jdff dff_B_lOF0kPk27_0(.din(w_dff_B_mXHIPi7r6_0),.dout(w_dff_B_lOF0kPk27_0),.clk(gclk));
	jdff dff_B_PyGoNv9p6_0(.din(w_dff_B_lOF0kPk27_0),.dout(w_dff_B_PyGoNv9p6_0),.clk(gclk));
	jdff dff_B_ludczpeP3_0(.din(w_dff_B_PyGoNv9p6_0),.dout(w_dff_B_ludczpeP3_0),.clk(gclk));
	jdff dff_B_3OlqcsDz3_0(.din(w_dff_B_ludczpeP3_0),.dout(w_dff_B_3OlqcsDz3_0),.clk(gclk));
	jdff dff_B_jJrx93m36_0(.din(w_dff_B_3OlqcsDz3_0),.dout(w_dff_B_jJrx93m36_0),.clk(gclk));
	jdff dff_B_b1uaOjDS4_0(.din(w_dff_B_jJrx93m36_0),.dout(w_dff_B_b1uaOjDS4_0),.clk(gclk));
	jdff dff_B_N9payxge5_0(.din(w_dff_B_b1uaOjDS4_0),.dout(w_dff_B_N9payxge5_0),.clk(gclk));
	jdff dff_B_wHRzwpWI8_0(.din(w_dff_B_N9payxge5_0),.dout(w_dff_B_wHRzwpWI8_0),.clk(gclk));
	jdff dff_B_4tHvCdM24_0(.din(w_dff_B_wHRzwpWI8_0),.dout(w_dff_B_4tHvCdM24_0),.clk(gclk));
	jdff dff_B_AwFToQub6_0(.din(w_dff_B_4tHvCdM24_0),.dout(w_dff_B_AwFToQub6_0),.clk(gclk));
	jdff dff_B_Rud5IheJ3_0(.din(w_dff_B_AwFToQub6_0),.dout(w_dff_B_Rud5IheJ3_0),.clk(gclk));
	jdff dff_B_Tylp1GK25_0(.din(w_dff_B_Rud5IheJ3_0),.dout(w_dff_B_Tylp1GK25_0),.clk(gclk));
	jdff dff_B_4oj8cpEW1_0(.din(w_dff_B_Tylp1GK25_0),.dout(w_dff_B_4oj8cpEW1_0),.clk(gclk));
	jdff dff_B_VWeBcbz51_0(.din(w_dff_B_4oj8cpEW1_0),.dout(w_dff_B_VWeBcbz51_0),.clk(gclk));
	jdff dff_B_KxkvSA1o5_0(.din(w_dff_B_VWeBcbz51_0),.dout(w_dff_B_KxkvSA1o5_0),.clk(gclk));
	jdff dff_B_V9uOycli7_0(.din(w_dff_B_KxkvSA1o5_0),.dout(w_dff_B_V9uOycli7_0),.clk(gclk));
	jdff dff_B_bVZczMbx8_0(.din(w_dff_B_V9uOycli7_0),.dout(w_dff_B_bVZczMbx8_0),.clk(gclk));
	jdff dff_B_8n3vo7RB0_1(.din(n1627),.dout(w_dff_B_8n3vo7RB0_1),.clk(gclk));
	jdff dff_B_h88qhk292_1(.din(w_dff_B_8n3vo7RB0_1),.dout(w_dff_B_h88qhk292_1),.clk(gclk));
	jdff dff_B_N3mal6mu1_1(.din(w_dff_B_h88qhk292_1),.dout(w_dff_B_N3mal6mu1_1),.clk(gclk));
	jdff dff_B_aucyYDED9_1(.din(w_dff_B_N3mal6mu1_1),.dout(w_dff_B_aucyYDED9_1),.clk(gclk));
	jdff dff_B_7yJ48Wmp3_1(.din(w_dff_B_aucyYDED9_1),.dout(w_dff_B_7yJ48Wmp3_1),.clk(gclk));
	jdff dff_B_pqxQBoJZ4_1(.din(w_dff_B_7yJ48Wmp3_1),.dout(w_dff_B_pqxQBoJZ4_1),.clk(gclk));
	jdff dff_B_dLr0mNqu5_1(.din(w_dff_B_pqxQBoJZ4_1),.dout(w_dff_B_dLr0mNqu5_1),.clk(gclk));
	jdff dff_B_ImSWn67M3_1(.din(w_dff_B_dLr0mNqu5_1),.dout(w_dff_B_ImSWn67M3_1),.clk(gclk));
	jdff dff_B_KU9aBWNF6_1(.din(w_dff_B_ImSWn67M3_1),.dout(w_dff_B_KU9aBWNF6_1),.clk(gclk));
	jdff dff_B_n4c1XlKr5_1(.din(w_dff_B_KU9aBWNF6_1),.dout(w_dff_B_n4c1XlKr5_1),.clk(gclk));
	jdff dff_B_bRad8Ntl3_1(.din(w_dff_B_n4c1XlKr5_1),.dout(w_dff_B_bRad8Ntl3_1),.clk(gclk));
	jdff dff_B_sywqYdfQ3_1(.din(w_dff_B_bRad8Ntl3_1),.dout(w_dff_B_sywqYdfQ3_1),.clk(gclk));
	jdff dff_B_HQJVhmfY9_1(.din(w_dff_B_sywqYdfQ3_1),.dout(w_dff_B_HQJVhmfY9_1),.clk(gclk));
	jdff dff_B_MQAqoOmp5_1(.din(w_dff_B_HQJVhmfY9_1),.dout(w_dff_B_MQAqoOmp5_1),.clk(gclk));
	jdff dff_B_Po53HvDG2_1(.din(w_dff_B_MQAqoOmp5_1),.dout(w_dff_B_Po53HvDG2_1),.clk(gclk));
	jdff dff_B_YY6E9Tr81_1(.din(w_dff_B_Po53HvDG2_1),.dout(w_dff_B_YY6E9Tr81_1),.clk(gclk));
	jdff dff_B_IMCEMDY18_1(.din(w_dff_B_YY6E9Tr81_1),.dout(w_dff_B_IMCEMDY18_1),.clk(gclk));
	jdff dff_B_auoXWo6O9_1(.din(w_dff_B_IMCEMDY18_1),.dout(w_dff_B_auoXWo6O9_1),.clk(gclk));
	jdff dff_B_e33LovgP0_1(.din(w_dff_B_auoXWo6O9_1),.dout(w_dff_B_e33LovgP0_1),.clk(gclk));
	jdff dff_B_ddURQ7Dr9_1(.din(n1642),.dout(w_dff_B_ddURQ7Dr9_1),.clk(gclk));
	jdff dff_B_GksMrAHL7_0(.din(n1649),.dout(w_dff_B_GksMrAHL7_0),.clk(gclk));
	jdff dff_B_SKtUkjFX0_0(.din(w_dff_B_GksMrAHL7_0),.dout(w_dff_B_SKtUkjFX0_0),.clk(gclk));
	jdff dff_B_lXl8u2807_0(.din(w_dff_B_SKtUkjFX0_0),.dout(w_dff_B_lXl8u2807_0),.clk(gclk));
	jdff dff_B_JlAfKRAv1_0(.din(w_dff_B_lXl8u2807_0),.dout(w_dff_B_JlAfKRAv1_0),.clk(gclk));
	jdff dff_B_VxsxfR1i8_0(.din(w_dff_B_JlAfKRAv1_0),.dout(w_dff_B_VxsxfR1i8_0),.clk(gclk));
	jdff dff_B_ZymxUA9Z4_0(.din(w_dff_B_VxsxfR1i8_0),.dout(w_dff_B_ZymxUA9Z4_0),.clk(gclk));
	jdff dff_B_rTnONUwH8_0(.din(w_dff_B_ZymxUA9Z4_0),.dout(w_dff_B_rTnONUwH8_0),.clk(gclk));
	jdff dff_B_Og2fEFdx8_0(.din(w_dff_B_rTnONUwH8_0),.dout(w_dff_B_Og2fEFdx8_0),.clk(gclk));
	jdff dff_B_5v2nRLVr1_0(.din(w_dff_B_Og2fEFdx8_0),.dout(w_dff_B_5v2nRLVr1_0),.clk(gclk));
	jdff dff_B_58IJzkPx7_0(.din(w_dff_B_5v2nRLVr1_0),.dout(w_dff_B_58IJzkPx7_0),.clk(gclk));
	jdff dff_B_mfk3XKas0_0(.din(w_dff_B_58IJzkPx7_0),.dout(w_dff_B_mfk3XKas0_0),.clk(gclk));
	jdff dff_B_nqUp5bem5_0(.din(w_dff_B_mfk3XKas0_0),.dout(w_dff_B_nqUp5bem5_0),.clk(gclk));
	jdff dff_B_AkmkdL2U3_0(.din(w_dff_B_nqUp5bem5_0),.dout(w_dff_B_AkmkdL2U3_0),.clk(gclk));
	jdff dff_B_0J3oHaDB2_0(.din(w_dff_B_AkmkdL2U3_0),.dout(w_dff_B_0J3oHaDB2_0),.clk(gclk));
	jdff dff_B_5GFmOFuN7_0(.din(w_dff_B_0J3oHaDB2_0),.dout(w_dff_B_5GFmOFuN7_0),.clk(gclk));
	jdff dff_B_8nt7m9RE2_0(.din(w_dff_B_5GFmOFuN7_0),.dout(w_dff_B_8nt7m9RE2_0),.clk(gclk));
	jdff dff_B_5WhggEDT5_0(.din(w_dff_B_8nt7m9RE2_0),.dout(w_dff_B_5WhggEDT5_0),.clk(gclk));
	jdff dff_B_5W8CGx180_0(.din(w_dff_B_5WhggEDT5_0),.dout(w_dff_B_5W8CGx180_0),.clk(gclk));
	jdff dff_B_zkO0tHSn5_1(.din(n1643),.dout(w_dff_B_zkO0tHSn5_1),.clk(gclk));
	jdff dff_B_I25RDzZ94_1(.din(w_dff_B_zkO0tHSn5_1),.dout(w_dff_B_I25RDzZ94_1),.clk(gclk));
	jdff dff_B_BXLNxTsJ5_1(.din(w_dff_B_I25RDzZ94_1),.dout(w_dff_B_BXLNxTsJ5_1),.clk(gclk));
	jdff dff_B_PdTixlrW5_1(.din(w_dff_B_BXLNxTsJ5_1),.dout(w_dff_B_PdTixlrW5_1),.clk(gclk));
	jdff dff_B_5EXA678H7_1(.din(w_dff_B_PdTixlrW5_1),.dout(w_dff_B_5EXA678H7_1),.clk(gclk));
	jdff dff_B_lLdSiesg9_1(.din(w_dff_B_5EXA678H7_1),.dout(w_dff_B_lLdSiesg9_1),.clk(gclk));
	jdff dff_B_lkYcCaAH7_1(.din(w_dff_B_lLdSiesg9_1),.dout(w_dff_B_lkYcCaAH7_1),.clk(gclk));
	jdff dff_B_ZAdAPF8j4_1(.din(w_dff_B_lkYcCaAH7_1),.dout(w_dff_B_ZAdAPF8j4_1),.clk(gclk));
	jdff dff_B_Q9bXY9iO6_1(.din(w_dff_B_ZAdAPF8j4_1),.dout(w_dff_B_Q9bXY9iO6_1),.clk(gclk));
	jdff dff_B_hIoZZVs60_1(.din(w_dff_B_Q9bXY9iO6_1),.dout(w_dff_B_hIoZZVs60_1),.clk(gclk));
	jdff dff_B_92wjE9lL0_1(.din(w_dff_B_hIoZZVs60_1),.dout(w_dff_B_92wjE9lL0_1),.clk(gclk));
	jdff dff_B_JC9ErbD70_1(.din(w_dff_B_92wjE9lL0_1),.dout(w_dff_B_JC9ErbD70_1),.clk(gclk));
	jdff dff_B_ZrC4OjzC0_1(.din(w_dff_B_JC9ErbD70_1),.dout(w_dff_B_ZrC4OjzC0_1),.clk(gclk));
	jdff dff_B_3XgyYXZy4_1(.din(w_dff_B_ZrC4OjzC0_1),.dout(w_dff_B_3XgyYXZy4_1),.clk(gclk));
	jdff dff_B_bM6IEAfH0_1(.din(w_dff_B_3XgyYXZy4_1),.dout(w_dff_B_bM6IEAfH0_1),.clk(gclk));
	jdff dff_B_egznxpg66_1(.din(w_dff_B_bM6IEAfH0_1),.dout(w_dff_B_egznxpg66_1),.clk(gclk));
	jdff dff_B_8iwuC1d94_1(.din(w_dff_B_egznxpg66_1),.dout(w_dff_B_8iwuC1d94_1),.clk(gclk));
	jdff dff_B_Jv6B9aF50_1(.din(w_dff_B_8iwuC1d94_1),.dout(w_dff_B_Jv6B9aF50_1),.clk(gclk));
	jdff dff_B_bZbagBGo7_1(.din(w_dff_B_Jv6B9aF50_1),.dout(w_dff_B_bZbagBGo7_1),.clk(gclk));
	jdff dff_B_sZtMb9X57_0(.din(n1628),.dout(w_dff_B_sZtMb9X57_0),.clk(gclk));
	jdff dff_B_MeOL8bvJ5_0(.din(w_dff_B_sZtMb9X57_0),.dout(w_dff_B_MeOL8bvJ5_0),.clk(gclk));
	jdff dff_B_s5lFu9w62_0(.din(w_dff_B_MeOL8bvJ5_0),.dout(w_dff_B_s5lFu9w62_0),.clk(gclk));
	jdff dff_B_1lp7X9HY6_0(.din(w_dff_B_s5lFu9w62_0),.dout(w_dff_B_1lp7X9HY6_0),.clk(gclk));
	jdff dff_B_YZFR1aXT5_0(.din(w_dff_B_1lp7X9HY6_0),.dout(w_dff_B_YZFR1aXT5_0),.clk(gclk));
	jdff dff_B_pJbITUhM1_0(.din(w_dff_B_YZFR1aXT5_0),.dout(w_dff_B_pJbITUhM1_0),.clk(gclk));
	jdff dff_B_ndNDPUJj3_0(.din(w_dff_B_pJbITUhM1_0),.dout(w_dff_B_ndNDPUJj3_0),.clk(gclk));
	jdff dff_B_FnEFXOok1_0(.din(w_dff_B_ndNDPUJj3_0),.dout(w_dff_B_FnEFXOok1_0),.clk(gclk));
	jdff dff_B_RLSgYVnb4_0(.din(w_dff_B_FnEFXOok1_0),.dout(w_dff_B_RLSgYVnb4_0),.clk(gclk));
	jdff dff_B_7TivSpXc5_0(.din(w_dff_B_RLSgYVnb4_0),.dout(w_dff_B_7TivSpXc5_0),.clk(gclk));
	jdff dff_B_98cSCAkM7_0(.din(w_dff_B_7TivSpXc5_0),.dout(w_dff_B_98cSCAkM7_0),.clk(gclk));
	jdff dff_B_QUkMZbLA4_0(.din(w_dff_B_98cSCAkM7_0),.dout(w_dff_B_QUkMZbLA4_0),.clk(gclk));
	jdff dff_B_UymDJ8TM2_0(.din(w_dff_B_QUkMZbLA4_0),.dout(w_dff_B_UymDJ8TM2_0),.clk(gclk));
	jdff dff_B_8neHo7o57_0(.din(w_dff_B_UymDJ8TM2_0),.dout(w_dff_B_8neHo7o57_0),.clk(gclk));
	jdff dff_B_sVCac5ow6_0(.din(w_dff_B_8neHo7o57_0),.dout(w_dff_B_sVCac5ow6_0),.clk(gclk));
	jdff dff_B_mKIAvnbD5_0(.din(w_dff_B_sVCac5ow6_0),.dout(w_dff_B_mKIAvnbD5_0),.clk(gclk));
	jdff dff_B_aj220N9X9_0(.din(w_dff_B_mKIAvnbD5_0),.dout(w_dff_B_aj220N9X9_0),.clk(gclk));
	jdff dff_B_xBJkETM87_0(.din(w_dff_B_aj220N9X9_0),.dout(w_dff_B_xBJkETM87_0),.clk(gclk));
	jdff dff_B_turOlrt26_0(.din(w_dff_B_xBJkETM87_0),.dout(w_dff_B_turOlrt26_0),.clk(gclk));
	jdff dff_B_6bZxOr787_1(.din(n1392),.dout(w_dff_B_6bZxOr787_1),.clk(gclk));
	jdff dff_B_9siOO4ek5_1(.din(w_dff_B_6bZxOr787_1),.dout(w_dff_B_9siOO4ek5_1),.clk(gclk));
	jdff dff_B_mOMU5UYN2_1(.din(w_dff_B_9siOO4ek5_1),.dout(w_dff_B_mOMU5UYN2_1),.clk(gclk));
	jdff dff_B_yTRY5S2l2_1(.din(w_dff_B_mOMU5UYN2_1),.dout(w_dff_B_yTRY5S2l2_1),.clk(gclk));
	jdff dff_B_dhj9MhGd1_1(.din(w_dff_B_yTRY5S2l2_1),.dout(w_dff_B_dhj9MhGd1_1),.clk(gclk));
	jdff dff_B_VJgNpd3v5_1(.din(w_dff_B_dhj9MhGd1_1),.dout(w_dff_B_VJgNpd3v5_1),.clk(gclk));
	jdff dff_A_5N9tgYEO1_1(.dout(w_n1447_0[1]),.din(w_dff_A_5N9tgYEO1_1),.clk(gclk));
	jdff dff_B_5zaBbffg4_1(.din(n1412),.dout(w_dff_B_5zaBbffg4_1),.clk(gclk));
	jdff dff_B_GGZBohVy0_1(.din(w_dff_B_5zaBbffg4_1),.dout(w_dff_B_GGZBohVy0_1),.clk(gclk));
	jdff dff_B_pV08APgv4_1(.din(w_dff_B_GGZBohVy0_1),.dout(w_dff_B_pV08APgv4_1),.clk(gclk));
	jdff dff_B_g1A5T19g6_1(.din(w_dff_B_pV08APgv4_1),.dout(w_dff_B_g1A5T19g6_1),.clk(gclk));
	jdff dff_B_rMH6wThe5_1(.din(w_dff_B_g1A5T19g6_1),.dout(w_dff_B_rMH6wThe5_1),.clk(gclk));
	jdff dff_B_Wb2gv5YS1_1(.din(w_dff_B_rMH6wThe5_1),.dout(w_dff_B_Wb2gv5YS1_1),.clk(gclk));
	jdff dff_B_B963ehN05_1(.din(w_dff_B_Wb2gv5YS1_1),.dout(w_dff_B_B963ehN05_1),.clk(gclk));
	jdff dff_B_LtgTD4Ez4_1(.din(w_dff_B_B963ehN05_1),.dout(w_dff_B_LtgTD4Ez4_1),.clk(gclk));
	jdff dff_B_zRcmY1Ug2_1(.din(w_dff_B_LtgTD4Ez4_1),.dout(w_dff_B_zRcmY1Ug2_1),.clk(gclk));
	jdff dff_B_LLiJKrcD2_1(.din(w_dff_B_zRcmY1Ug2_1),.dout(w_dff_B_LLiJKrcD2_1),.clk(gclk));
	jdff dff_B_jNf0BP9R3_0(.din(n1443),.dout(w_dff_B_jNf0BP9R3_0),.clk(gclk));
	jdff dff_B_fKpEoIgw7_0(.din(n1440),.dout(w_dff_B_fKpEoIgw7_0),.clk(gclk));
	jdff dff_A_nCygsGsv6_1(.dout(w_n1438_0[1]),.din(w_dff_A_nCygsGsv6_1),.clk(gclk));
	jdff dff_A_9u0yrDq81_1(.dout(w_dff_A_nCygsGsv6_1),.din(w_dff_A_9u0yrDq81_1),.clk(gclk));
	jdff dff_A_e0btWtwj6_1(.dout(w_dff_A_9u0yrDq81_1),.din(w_dff_A_e0btWtwj6_1),.clk(gclk));
	jdff dff_B_wzRzGDvU7_0(.din(n1437),.dout(w_dff_B_wzRzGDvU7_0),.clk(gclk));
	jdff dff_B_EeCOdrtz7_1(.din(n1427),.dout(w_dff_B_EeCOdrtz7_1),.clk(gclk));
	jdff dff_B_fYc4TshO6_1(.din(n1428),.dout(w_dff_B_fYc4TshO6_1),.clk(gclk));
	jdff dff_B_qUs1wJ4M1_1(.din(w_dff_B_fYc4TshO6_1),.dout(w_dff_B_qUs1wJ4M1_1),.clk(gclk));
	jdff dff_B_iHtukHpL5_1(.din(w_dff_B_qUs1wJ4M1_1),.dout(w_dff_B_iHtukHpL5_1),.clk(gclk));
	jdff dff_B_fUbz4NVr5_1(.din(w_dff_B_iHtukHpL5_1),.dout(w_dff_B_fUbz4NVr5_1),.clk(gclk));
	jdff dff_B_qbgis4aG8_1(.din(w_dff_B_fUbz4NVr5_1),.dout(w_dff_B_qbgis4aG8_1),.clk(gclk));
	jdff dff_B_5e9lLEwP3_1(.din(w_dff_B_qbgis4aG8_1),.dout(w_dff_B_5e9lLEwP3_1),.clk(gclk));
	jdff dff_B_jkjH0v9K4_1(.din(w_dff_B_5e9lLEwP3_1),.dout(w_dff_B_jkjH0v9K4_1),.clk(gclk));
	jdff dff_B_zScbqlEf1_1(.din(w_dff_B_jkjH0v9K4_1),.dout(w_dff_B_zScbqlEf1_1),.clk(gclk));
	jdff dff_B_Yymp456X4_1(.din(w_dff_B_zScbqlEf1_1),.dout(w_dff_B_Yymp456X4_1),.clk(gclk));
	jdff dff_B_l9yYNM3y7_1(.din(w_dff_B_Yymp456X4_1),.dout(w_dff_B_l9yYNM3y7_1),.clk(gclk));
	jdff dff_B_02WrUaWC2_1(.din(w_dff_B_l9yYNM3y7_1),.dout(w_dff_B_02WrUaWC2_1),.clk(gclk));
	jdff dff_B_LzQJJeCb3_1(.din(n1414),.dout(w_dff_B_LzQJJeCb3_1),.clk(gclk));
	jdff dff_B_fm3FDxps1_1(.din(w_dff_B_LzQJJeCb3_1),.dout(w_dff_B_fm3FDxps1_1),.clk(gclk));
	jdff dff_B_IJO3eluU6_1(.din(w_dff_B_fm3FDxps1_1),.dout(w_dff_B_IJO3eluU6_1),.clk(gclk));
	jdff dff_B_8XP8jZ1L9_1(.din(w_dff_B_IJO3eluU6_1),.dout(w_dff_B_8XP8jZ1L9_1),.clk(gclk));
	jdff dff_B_2Lkh4R635_1(.din(n1423),.dout(w_dff_B_2Lkh4R635_1),.clk(gclk));
	jdff dff_B_VoHCHtBi5_0(.din(n1422),.dout(w_dff_B_VoHCHtBi5_0),.clk(gclk));
	jdff dff_A_RzFfuChi6_0(.dout(w_n1421_0[0]),.din(w_dff_A_RzFfuChi6_0),.clk(gclk));
	jdff dff_A_H3ScOOKu0_0(.dout(w_dff_A_RzFfuChi6_0),.din(w_dff_A_H3ScOOKu0_0),.clk(gclk));
	jdff dff_A_x8XgfZtr4_0(.dout(w_dff_A_H3ScOOKu0_0),.din(w_dff_A_x8XgfZtr4_0),.clk(gclk));
	jdff dff_B_Zfy0bBXR1_1(.din(n1415),.dout(w_dff_B_Zfy0bBXR1_1),.clk(gclk));
	jdff dff_A_6A7OUpET3_1(.dout(w_n828_0[1]),.din(w_dff_A_6A7OUpET3_1),.clk(gclk));
	jdff dff_A_5DQrxhTw1_1(.dout(w_dff_A_6A7OUpET3_1),.din(w_dff_A_5DQrxhTw1_1),.clk(gclk));
	jdff dff_A_mIDnUMUY1_1(.dout(w_dff_A_5DQrxhTw1_1),.din(w_dff_A_mIDnUMUY1_1),.clk(gclk));
	jdff dff_A_E4Rsaesr7_1(.dout(w_dff_A_mIDnUMUY1_1),.din(w_dff_A_E4Rsaesr7_1),.clk(gclk));
	jdff dff_A_f8jnsMYH5_1(.dout(w_dff_A_E4Rsaesr7_1),.din(w_dff_A_f8jnsMYH5_1),.clk(gclk));
	jdff dff_A_bsUiUq3R8_1(.dout(w_dff_A_f8jnsMYH5_1),.din(w_dff_A_bsUiUq3R8_1),.clk(gclk));
	jdff dff_A_yiHJB6z70_2(.dout(w_n828_0[2]),.din(w_dff_A_yiHJB6z70_2),.clk(gclk));
	jdff dff_A_A0PVhH983_2(.dout(w_dff_A_yiHJB6z70_2),.din(w_dff_A_A0PVhH983_2),.clk(gclk));
	jdff dff_B_kpcoNTEd7_2(.din(n787),.dout(w_dff_B_kpcoNTEd7_2),.clk(gclk));
	jdff dff_B_tXUJF08v1_2(.din(w_dff_B_kpcoNTEd7_2),.dout(w_dff_B_tXUJF08v1_2),.clk(gclk));
	jdff dff_B_6eRvWGTO2_2(.din(w_dff_B_tXUJF08v1_2),.dout(w_dff_B_6eRvWGTO2_2),.clk(gclk));
	jdff dff_B_lWDXr2Zo0_2(.din(w_dff_B_6eRvWGTO2_2),.dout(w_dff_B_lWDXr2Zo0_2),.clk(gclk));
	jdff dff_B_Xv9pZukw0_2(.din(w_dff_B_lWDXr2Zo0_2),.dout(w_dff_B_Xv9pZukw0_2),.clk(gclk));
	jdff dff_B_AtfNQjRJ0_2(.din(w_dff_B_Xv9pZukw0_2),.dout(w_dff_B_AtfNQjRJ0_2),.clk(gclk));
	jdff dff_B_mechHiC69_2(.din(w_dff_B_AtfNQjRJ0_2),.dout(w_dff_B_mechHiC69_2),.clk(gclk));
	jdff dff_B_6D9HwHrJ2_2(.din(w_dff_B_mechHiC69_2),.dout(w_dff_B_6D9HwHrJ2_2),.clk(gclk));
	jdff dff_B_hcZWEMPy7_2(.din(w_dff_B_6D9HwHrJ2_2),.dout(w_dff_B_hcZWEMPy7_2),.clk(gclk));
	jdff dff_A_Txqjbibg9_1(.dout(w_n779_0[1]),.din(w_dff_A_Txqjbibg9_1),.clk(gclk));
	jdff dff_A_Zzfl8d7n6_1(.dout(w_dff_A_Txqjbibg9_1),.din(w_dff_A_Zzfl8d7n6_1),.clk(gclk));
	jdff dff_A_fVfHPFEl1_1(.dout(w_dff_A_Zzfl8d7n6_1),.din(w_dff_A_fVfHPFEl1_1),.clk(gclk));
	jdff dff_A_oTy64uHq9_1(.dout(w_dff_A_fVfHPFEl1_1),.din(w_dff_A_oTy64uHq9_1),.clk(gclk));
	jdff dff_A_1TEmmUns4_1(.dout(w_dff_A_oTy64uHq9_1),.din(w_dff_A_1TEmmUns4_1),.clk(gclk));
	jdff dff_A_4Pe0hfd69_1(.dout(w_dff_A_1TEmmUns4_1),.din(w_dff_A_4Pe0hfd69_1),.clk(gclk));
	jdff dff_A_0pVFSIYZ0_1(.dout(w_dff_A_4Pe0hfd69_1),.din(w_dff_A_0pVFSIYZ0_1),.clk(gclk));
	jdff dff_A_QVo1U4UG6_1(.dout(w_dff_A_0pVFSIYZ0_1),.din(w_dff_A_QVo1U4UG6_1),.clk(gclk));
	jdff dff_A_PHILE3gA2_1(.dout(w_dff_A_QVo1U4UG6_1),.din(w_dff_A_PHILE3gA2_1),.clk(gclk));
	jdff dff_A_rTKPoJwV1_1(.dout(w_dff_A_PHILE3gA2_1),.din(w_dff_A_rTKPoJwV1_1),.clk(gclk));
	jdff dff_A_fwg9U8jF2_1(.dout(w_dff_A_rTKPoJwV1_1),.din(w_dff_A_fwg9U8jF2_1),.clk(gclk));
	jdff dff_A_ylRM2eMt7_1(.dout(w_dff_A_fwg9U8jF2_1),.din(w_dff_A_ylRM2eMt7_1),.clk(gclk));
	jdff dff_A_mtdFSZKM7_1(.dout(w_n636_1[1]),.din(w_dff_A_mtdFSZKM7_1),.clk(gclk));
	jdff dff_A_VzvL9tk17_1(.dout(w_dff_A_mtdFSZKM7_1),.din(w_dff_A_VzvL9tk17_1),.clk(gclk));
	jdff dff_A_6l12njUS4_2(.dout(w_n636_0[2]),.din(w_dff_A_6l12njUS4_2),.clk(gclk));
	jdff dff_A_wDmslZSH7_0(.dout(w_n1411_0[0]),.din(w_dff_A_wDmslZSH7_0),.clk(gclk));
	jdff dff_A_fBeSBzmf9_0(.dout(w_dff_A_wDmslZSH7_0),.din(w_dff_A_fBeSBzmf9_0),.clk(gclk));
	jdff dff_A_gRmMcFN92_0(.dout(w_dff_A_fBeSBzmf9_0),.din(w_dff_A_gRmMcFN92_0),.clk(gclk));
	jdff dff_A_NzKBFKV83_0(.dout(w_dff_A_gRmMcFN92_0),.din(w_dff_A_NzKBFKV83_0),.clk(gclk));
	jdff dff_A_naENVEYz1_0(.dout(w_dff_A_NzKBFKV83_0),.din(w_dff_A_naENVEYz1_0),.clk(gclk));
	jdff dff_A_QC4rYQS22_0(.dout(w_dff_A_naENVEYz1_0),.din(w_dff_A_QC4rYQS22_0),.clk(gclk));
	jdff dff_A_715MGgWo7_0(.dout(w_dff_A_QC4rYQS22_0),.din(w_dff_A_715MGgWo7_0),.clk(gclk));
	jdff dff_A_dNhsUvwf9_0(.dout(w_dff_A_715MGgWo7_0),.din(w_dff_A_dNhsUvwf9_0),.clk(gclk));
	jdff dff_A_TqAmVVtt4_0(.dout(w_dff_A_dNhsUvwf9_0),.din(w_dff_A_TqAmVVtt4_0),.clk(gclk));
	jdff dff_A_7YHxvuJ43_0(.dout(w_dff_A_TqAmVVtt4_0),.din(w_dff_A_7YHxvuJ43_0),.clk(gclk));
	jdff dff_A_w4ia18uG3_0(.dout(w_dff_A_7YHxvuJ43_0),.din(w_dff_A_w4ia18uG3_0),.clk(gclk));
	jdff dff_A_sXYZBzkT3_0(.dout(w_n1409_0[0]),.din(w_dff_A_sXYZBzkT3_0),.clk(gclk));
	jdff dff_B_z6nn5o6q1_1(.din(n1405),.dout(w_dff_B_z6nn5o6q1_1),.clk(gclk));
	jdff dff_B_ZxZfcKbg4_0(.din(n1407),.dout(w_dff_B_ZxZfcKbg4_0),.clk(gclk));
	jdff dff_B_d9hPlEia5_0(.din(w_dff_B_ZxZfcKbg4_0),.dout(w_dff_B_d9hPlEia5_0),.clk(gclk));
	jdff dff_B_1mqFA4Qc4_0(.din(w_dff_B_d9hPlEia5_0),.dout(w_dff_B_1mqFA4Qc4_0),.clk(gclk));
	jdff dff_B_r0NRFXqF2_0(.din(w_dff_B_1mqFA4Qc4_0),.dout(w_dff_B_r0NRFXqF2_0),.clk(gclk));
	jdff dff_B_gZekIbB44_0(.din(n1404),.dout(w_dff_B_gZekIbB44_0),.clk(gclk));
	jdff dff_B_jwnaOYvi6_0(.din(w_dff_B_gZekIbB44_0),.dout(w_dff_B_jwnaOYvi6_0),.clk(gclk));
	jdff dff_B_r2Z0Yv1L6_0(.din(n1393),.dout(w_dff_B_r2Z0Yv1L6_0),.clk(gclk));
	jdff dff_B_jPkWfscm1_0(.din(w_dff_B_r2Z0Yv1L6_0),.dout(w_dff_B_jPkWfscm1_0),.clk(gclk));
	jdff dff_B_Gpxjw03t9_0(.din(w_dff_B_jPkWfscm1_0),.dout(w_dff_B_Gpxjw03t9_0),.clk(gclk));
	jdff dff_A_o6Ok0uWN0_0(.dout(w_n631_0[0]),.din(w_dff_A_o6Ok0uWN0_0),.clk(gclk));
	jdff dff_A_g1iU1Asj6_0(.dout(w_dff_A_o6Ok0uWN0_0),.din(w_dff_A_g1iU1Asj6_0),.clk(gclk));
	jdff dff_A_yhM1GGPX8_0(.dout(w_dff_A_g1iU1Asj6_0),.din(w_dff_A_yhM1GGPX8_0),.clk(gclk));
	jdff dff_A_W3AJjpbZ6_1(.dout(w_n629_0[1]),.din(w_dff_A_W3AJjpbZ6_1),.clk(gclk));
	jdff dff_A_PrVgnCwx1_1(.dout(w_dff_A_W3AJjpbZ6_1),.din(w_dff_A_PrVgnCwx1_1),.clk(gclk));
	jdff dff_A_a62VI9RO2_1(.dout(w_dff_A_PrVgnCwx1_1),.din(w_dff_A_a62VI9RO2_1),.clk(gclk));
	jdff dff_A_QCo5rrFG2_0(.dout(w_n625_0[0]),.din(w_dff_A_QCo5rrFG2_0),.clk(gclk));
	jdff dff_A_41iniY6v3_2(.dout(w_n625_0[2]),.din(w_dff_A_41iniY6v3_2),.clk(gclk));
	jdff dff_A_Gxmw2GQZ2_0(.dout(w_n623_0[0]),.din(w_dff_A_Gxmw2GQZ2_0),.clk(gclk));
	jdff dff_B_LnF8sMbi2_1(.din(n711),.dout(w_dff_B_LnF8sMbi2_1),.clk(gclk));
	jdff dff_B_BIiJJkwU9_1(.din(w_dff_B_LnF8sMbi2_1),.dout(w_dff_B_BIiJJkwU9_1),.clk(gclk));
	jdff dff_B_xyxYBYEl9_1(.din(w_dff_B_BIiJJkwU9_1),.dout(w_dff_B_xyxYBYEl9_1),.clk(gclk));
	jdff dff_B_VreztqLC8_1(.din(w_dff_B_xyxYBYEl9_1),.dout(w_dff_B_VreztqLC8_1),.clk(gclk));
	jdff dff_B_YAseiAYS2_1(.din(w_dff_B_VreztqLC8_1),.dout(w_dff_B_YAseiAYS2_1),.clk(gclk));
	jdff dff_B_qNVll6yt7_1(.din(w_dff_B_YAseiAYS2_1),.dout(w_dff_B_qNVll6yt7_1),.clk(gclk));
	jdff dff_B_Tc99gfYc0_1(.din(n712),.dout(w_dff_B_Tc99gfYc0_1),.clk(gclk));
	jdff dff_B_BqxP2BEn1_1(.din(w_dff_B_Tc99gfYc0_1),.dout(w_dff_B_BqxP2BEn1_1),.clk(gclk));
	jdff dff_B_OzkxPolt3_1(.din(w_dff_B_BqxP2BEn1_1),.dout(w_dff_B_OzkxPolt3_1),.clk(gclk));
	jdff dff_B_8rssqo1N2_1(.din(w_dff_B_OzkxPolt3_1),.dout(w_dff_B_8rssqo1N2_1),.clk(gclk));
	jdff dff_B_xpRPAu6s1_1(.din(w_dff_B_8rssqo1N2_1),.dout(w_dff_B_xpRPAu6s1_1),.clk(gclk));
	jdff dff_B_eHJf75vv5_1(.din(n713),.dout(w_dff_B_eHJf75vv5_1),.clk(gclk));
	jdff dff_B_GfqzFmgf1_1(.din(w_dff_B_eHJf75vv5_1),.dout(w_dff_B_GfqzFmgf1_1),.clk(gclk));
	jdff dff_B_Oe513zkN7_1(.din(w_dff_B_GfqzFmgf1_1),.dout(w_dff_B_Oe513zkN7_1),.clk(gclk));
	jdff dff_B_Q7B98Heb2_1(.din(w_dff_B_Oe513zkN7_1),.dout(w_dff_B_Q7B98Heb2_1),.clk(gclk));
	jdff dff_A_OEnd0fHr7_0(.dout(w_n723_0[0]),.din(w_dff_A_OEnd0fHr7_0),.clk(gclk));
	jdff dff_A_uK0Xd9Vt0_0(.dout(w_n621_2[0]),.din(w_dff_A_uK0Xd9Vt0_0),.clk(gclk));
	jdff dff_A_GyvaTXiS2_1(.dout(w_n721_0[1]),.din(w_dff_A_GyvaTXiS2_1),.clk(gclk));
	jdff dff_A_GqrbQujp2_1(.dout(w_dff_A_GyvaTXiS2_1),.din(w_dff_A_GqrbQujp2_1),.clk(gclk));
	jdff dff_A_c9idzpQo8_1(.dout(w_dff_A_GqrbQujp2_1),.din(w_dff_A_c9idzpQo8_1),.clk(gclk));
	jdff dff_A_QMAibGF28_1(.dout(w_dff_A_c9idzpQo8_1),.din(w_dff_A_QMAibGF28_1),.clk(gclk));
	jdff dff_A_YxPcOlQR0_1(.dout(w_dff_A_QMAibGF28_1),.din(w_dff_A_YxPcOlQR0_1),.clk(gclk));
	jdff dff_A_4MaBBqXA9_1(.dout(w_dff_A_YxPcOlQR0_1),.din(w_dff_A_4MaBBqXA9_1),.clk(gclk));
	jdff dff_A_ezdLpXPg4_1(.dout(w_n717_0[1]),.din(w_dff_A_ezdLpXPg4_1),.clk(gclk));
	jdff dff_A_Ufs7lqJq2_1(.dout(w_dff_A_ezdLpXPg4_1),.din(w_dff_A_Ufs7lqJq2_1),.clk(gclk));
	jdff dff_A_nsxbk5Go9_1(.dout(w_dff_A_Ufs7lqJq2_1),.din(w_dff_A_nsxbk5Go9_1),.clk(gclk));
	jdff dff_A_5xlRuwxL9_2(.dout(w_n717_0[2]),.din(w_dff_A_5xlRuwxL9_2),.clk(gclk));
	jdff dff_A_o3ibLdIi1_2(.dout(w_dff_A_5xlRuwxL9_2),.din(w_dff_A_o3ibLdIi1_2),.clk(gclk));
	jdff dff_A_NNKvvsPr7_0(.dout(w_n614_2[0]),.din(w_dff_A_NNKvvsPr7_0),.clk(gclk));
	jdff dff_A_KSXrmRRr3_0(.dout(w_dff_A_NNKvvsPr7_0),.din(w_dff_A_KSXrmRRr3_0),.clk(gclk));
	jdff dff_A_HJLLE2YR5_0(.dout(w_dff_A_KSXrmRRr3_0),.din(w_dff_A_HJLLE2YR5_0),.clk(gclk));
	jdff dff_B_gz6R6oVC8_2(.din(n1624),.dout(w_dff_B_gz6R6oVC8_2),.clk(gclk));
	jdff dff_B_tExL2pd21_2(.din(w_dff_B_gz6R6oVC8_2),.dout(w_dff_B_tExL2pd21_2),.clk(gclk));
	jdff dff_B_s79O3IVw3_2(.din(w_dff_B_tExL2pd21_2),.dout(w_dff_B_s79O3IVw3_2),.clk(gclk));
	jdff dff_B_pTRwyhQr3_2(.din(w_dff_B_s79O3IVw3_2),.dout(w_dff_B_pTRwyhQr3_2),.clk(gclk));
	jdff dff_B_acY2Vds50_2(.din(w_dff_B_pTRwyhQr3_2),.dout(w_dff_B_acY2Vds50_2),.clk(gclk));
	jdff dff_B_kQjNf0Ez3_2(.din(w_dff_B_acY2Vds50_2),.dout(w_dff_B_kQjNf0Ez3_2),.clk(gclk));
	jdff dff_B_vIR1s6d80_2(.din(w_dff_B_kQjNf0Ez3_2),.dout(w_dff_B_vIR1s6d80_2),.clk(gclk));
	jdff dff_B_FjLdEi1b4_2(.din(w_dff_B_vIR1s6d80_2),.dout(w_dff_B_FjLdEi1b4_2),.clk(gclk));
	jdff dff_B_0ZaLwdyt5_2(.din(w_dff_B_FjLdEi1b4_2),.dout(w_dff_B_0ZaLwdyt5_2),.clk(gclk));
	jdff dff_B_nVuEXnZw3_2(.din(w_dff_B_0ZaLwdyt5_2),.dout(w_dff_B_nVuEXnZw3_2),.clk(gclk));
	jdff dff_B_8utvpYlG1_2(.din(w_dff_B_nVuEXnZw3_2),.dout(w_dff_B_8utvpYlG1_2),.clk(gclk));
	jdff dff_B_U0al0I6L3_2(.din(w_dff_B_8utvpYlG1_2),.dout(w_dff_B_U0al0I6L3_2),.clk(gclk));
	jdff dff_B_hdSSqI6c3_2(.din(w_dff_B_U0al0I6L3_2),.dout(w_dff_B_hdSSqI6c3_2),.clk(gclk));
	jdff dff_B_gkIOj6l26_2(.din(w_dff_B_hdSSqI6c3_2),.dout(w_dff_B_gkIOj6l26_2),.clk(gclk));
	jdff dff_B_Iwg9H4X03_2(.din(w_dff_B_gkIOj6l26_2),.dout(w_dff_B_Iwg9H4X03_2),.clk(gclk));
	jdff dff_B_f2i64VtA7_2(.din(w_dff_B_Iwg9H4X03_2),.dout(w_dff_B_f2i64VtA7_2),.clk(gclk));
	jdff dff_B_71eaoaDk3_2(.din(w_dff_B_f2i64VtA7_2),.dout(w_dff_B_71eaoaDk3_2),.clk(gclk));
	jdff dff_B_5t5qpv1I5_2(.din(w_dff_B_71eaoaDk3_2),.dout(w_dff_B_5t5qpv1I5_2),.clk(gclk));
	jdff dff_B_vHwQew9u1_2(.din(w_dff_B_5t5qpv1I5_2),.dout(w_dff_B_vHwQew9u1_2),.clk(gclk));
	jdff dff_B_wzPkVA5E0_2(.din(w_dff_B_vHwQew9u1_2),.dout(w_dff_B_wzPkVA5E0_2),.clk(gclk));
	jdff dff_B_BTqCJAI29_2(.din(w_dff_B_wzPkVA5E0_2),.dout(w_dff_B_BTqCJAI29_2),.clk(gclk));
	jdff dff_B_aSJdigHj0_2(.din(w_dff_B_BTqCJAI29_2),.dout(w_dff_B_aSJdigHj0_2),.clk(gclk));
	jdff dff_B_yotyiVqZ9_2(.din(w_dff_B_aSJdigHj0_2),.dout(w_dff_B_yotyiVqZ9_2),.clk(gclk));
	jdff dff_B_eJRdOaJC4_2(.din(w_dff_B_yotyiVqZ9_2),.dout(w_dff_B_eJRdOaJC4_2),.clk(gclk));
	jdff dff_A_L8i6nSmj8_1(.dout(w_dff_A_nC8NIUml7_0),.din(w_dff_A_L8i6nSmj8_1),.clk(gclk));
	jdff dff_A_nC8NIUml7_0(.dout(w_dff_A_BY1mYJK41_0),.din(w_dff_A_nC8NIUml7_0),.clk(gclk));
	jdff dff_A_BY1mYJK41_0(.dout(w_dff_A_b73VTaDF7_0),.din(w_dff_A_BY1mYJK41_0),.clk(gclk));
	jdff dff_A_b73VTaDF7_0(.dout(w_dff_A_UyijAhBH0_0),.din(w_dff_A_b73VTaDF7_0),.clk(gclk));
	jdff dff_A_UyijAhBH0_0(.dout(w_dff_A_sNYrpXW42_0),.din(w_dff_A_UyijAhBH0_0),.clk(gclk));
	jdff dff_A_sNYrpXW42_0(.dout(w_dff_A_zWDWptYv9_0),.din(w_dff_A_sNYrpXW42_0),.clk(gclk));
	jdff dff_A_zWDWptYv9_0(.dout(w_dff_A_8R0OgeLw1_0),.din(w_dff_A_zWDWptYv9_0),.clk(gclk));
	jdff dff_A_8R0OgeLw1_0(.dout(w_dff_A_1HEAJ2Rf5_0),.din(w_dff_A_8R0OgeLw1_0),.clk(gclk));
	jdff dff_A_1HEAJ2Rf5_0(.dout(w_dff_A_0HRkchec2_0),.din(w_dff_A_1HEAJ2Rf5_0),.clk(gclk));
	jdff dff_A_0HRkchec2_0(.dout(w_dff_A_RyHajLb78_0),.din(w_dff_A_0HRkchec2_0),.clk(gclk));
	jdff dff_A_RyHajLb78_0(.dout(w_dff_A_iePnse2A4_0),.din(w_dff_A_RyHajLb78_0),.clk(gclk));
	jdff dff_A_iePnse2A4_0(.dout(w_dff_A_w85hnXY70_0),.din(w_dff_A_iePnse2A4_0),.clk(gclk));
	jdff dff_A_w85hnXY70_0(.dout(w_dff_A_bkZH3Xcz7_0),.din(w_dff_A_w85hnXY70_0),.clk(gclk));
	jdff dff_A_bkZH3Xcz7_0(.dout(w_dff_A_rz6xaLAj5_0),.din(w_dff_A_bkZH3Xcz7_0),.clk(gclk));
	jdff dff_A_rz6xaLAj5_0(.dout(w_dff_A_OGwDk4DX4_0),.din(w_dff_A_rz6xaLAj5_0),.clk(gclk));
	jdff dff_A_OGwDk4DX4_0(.dout(w_dff_A_ixQCzRUg9_0),.din(w_dff_A_OGwDk4DX4_0),.clk(gclk));
	jdff dff_A_ixQCzRUg9_0(.dout(w_dff_A_LhOp4ex32_0),.din(w_dff_A_ixQCzRUg9_0),.clk(gclk));
	jdff dff_A_LhOp4ex32_0(.dout(w_dff_A_32OQkVZa1_0),.din(w_dff_A_LhOp4ex32_0),.clk(gclk));
	jdff dff_A_32OQkVZa1_0(.dout(w_dff_A_G9K6tBZ61_0),.din(w_dff_A_32OQkVZa1_0),.clk(gclk));
	jdff dff_A_G9K6tBZ61_0(.dout(w_dff_A_D4IT5YDC8_0),.din(w_dff_A_G9K6tBZ61_0),.clk(gclk));
	jdff dff_A_D4IT5YDC8_0(.dout(w_dff_A_reQRNsTe7_0),.din(w_dff_A_D4IT5YDC8_0),.clk(gclk));
	jdff dff_A_reQRNsTe7_0(.dout(w_dff_A_tehqSbla9_0),.din(w_dff_A_reQRNsTe7_0),.clk(gclk));
	jdff dff_A_tehqSbla9_0(.dout(w_dff_A_2UR8aYlw4_0),.din(w_dff_A_tehqSbla9_0),.clk(gclk));
	jdff dff_A_2UR8aYlw4_0(.dout(w_dff_A_SctOiIYD5_0),.din(w_dff_A_2UR8aYlw4_0),.clk(gclk));
	jdff dff_A_SctOiIYD5_0(.dout(w_dff_A_iAL19hqC7_0),.din(w_dff_A_SctOiIYD5_0),.clk(gclk));
	jdff dff_A_iAL19hqC7_0(.dout(G144),.din(w_dff_A_iAL19hqC7_0),.clk(gclk));
	jdff dff_A_xzFbqVFy4_1(.dout(w_dff_A_mdeFull68_0),.din(w_dff_A_xzFbqVFy4_1),.clk(gclk));
	jdff dff_A_mdeFull68_0(.dout(w_dff_A_qpTcncIA8_0),.din(w_dff_A_mdeFull68_0),.clk(gclk));
	jdff dff_A_qpTcncIA8_0(.dout(w_dff_A_G9ZYLKqt8_0),.din(w_dff_A_qpTcncIA8_0),.clk(gclk));
	jdff dff_A_G9ZYLKqt8_0(.dout(w_dff_A_VBu5CG410_0),.din(w_dff_A_G9ZYLKqt8_0),.clk(gclk));
	jdff dff_A_VBu5CG410_0(.dout(w_dff_A_9u2UjhkD7_0),.din(w_dff_A_VBu5CG410_0),.clk(gclk));
	jdff dff_A_9u2UjhkD7_0(.dout(w_dff_A_r8IzaxXH4_0),.din(w_dff_A_9u2UjhkD7_0),.clk(gclk));
	jdff dff_A_r8IzaxXH4_0(.dout(w_dff_A_HASDwZ0E1_0),.din(w_dff_A_r8IzaxXH4_0),.clk(gclk));
	jdff dff_A_HASDwZ0E1_0(.dout(w_dff_A_GB8Aja8V0_0),.din(w_dff_A_HASDwZ0E1_0),.clk(gclk));
	jdff dff_A_GB8Aja8V0_0(.dout(w_dff_A_QMsyAdqG1_0),.din(w_dff_A_GB8Aja8V0_0),.clk(gclk));
	jdff dff_A_QMsyAdqG1_0(.dout(w_dff_A_Z9WzIFaZ6_0),.din(w_dff_A_QMsyAdqG1_0),.clk(gclk));
	jdff dff_A_Z9WzIFaZ6_0(.dout(w_dff_A_93yMKHsq2_0),.din(w_dff_A_Z9WzIFaZ6_0),.clk(gclk));
	jdff dff_A_93yMKHsq2_0(.dout(w_dff_A_chYaKOcK7_0),.din(w_dff_A_93yMKHsq2_0),.clk(gclk));
	jdff dff_A_chYaKOcK7_0(.dout(w_dff_A_HCo5tBmy8_0),.din(w_dff_A_chYaKOcK7_0),.clk(gclk));
	jdff dff_A_HCo5tBmy8_0(.dout(w_dff_A_mWZCSMJ39_0),.din(w_dff_A_HCo5tBmy8_0),.clk(gclk));
	jdff dff_A_mWZCSMJ39_0(.dout(w_dff_A_9Qa2rzvi7_0),.din(w_dff_A_mWZCSMJ39_0),.clk(gclk));
	jdff dff_A_9Qa2rzvi7_0(.dout(w_dff_A_mogR2yJN6_0),.din(w_dff_A_9Qa2rzvi7_0),.clk(gclk));
	jdff dff_A_mogR2yJN6_0(.dout(w_dff_A_G3WcGPul8_0),.din(w_dff_A_mogR2yJN6_0),.clk(gclk));
	jdff dff_A_G3WcGPul8_0(.dout(w_dff_A_FqgHiXhR5_0),.din(w_dff_A_G3WcGPul8_0),.clk(gclk));
	jdff dff_A_FqgHiXhR5_0(.dout(w_dff_A_WlktV3d53_0),.din(w_dff_A_FqgHiXhR5_0),.clk(gclk));
	jdff dff_A_WlktV3d53_0(.dout(w_dff_A_s3zZi4AZ3_0),.din(w_dff_A_WlktV3d53_0),.clk(gclk));
	jdff dff_A_s3zZi4AZ3_0(.dout(w_dff_A_GmDXqLHv5_0),.din(w_dff_A_s3zZi4AZ3_0),.clk(gclk));
	jdff dff_A_GmDXqLHv5_0(.dout(w_dff_A_xpQ2pYsZ3_0),.din(w_dff_A_GmDXqLHv5_0),.clk(gclk));
	jdff dff_A_xpQ2pYsZ3_0(.dout(w_dff_A_O0a02aXr0_0),.din(w_dff_A_xpQ2pYsZ3_0),.clk(gclk));
	jdff dff_A_O0a02aXr0_0(.dout(w_dff_A_lotCgd6q8_0),.din(w_dff_A_O0a02aXr0_0),.clk(gclk));
	jdff dff_A_lotCgd6q8_0(.dout(w_dff_A_kNLoaKsm3_0),.din(w_dff_A_lotCgd6q8_0),.clk(gclk));
	jdff dff_A_kNLoaKsm3_0(.dout(G298),.din(w_dff_A_kNLoaKsm3_0),.clk(gclk));
	jdff dff_A_MwhKPAJt6_1(.dout(w_dff_A_8DSwKiPK5_0),.din(w_dff_A_MwhKPAJt6_1),.clk(gclk));
	jdff dff_A_8DSwKiPK5_0(.dout(w_dff_A_YDBqf7dz2_0),.din(w_dff_A_8DSwKiPK5_0),.clk(gclk));
	jdff dff_A_YDBqf7dz2_0(.dout(w_dff_A_3OkWTd0k6_0),.din(w_dff_A_YDBqf7dz2_0),.clk(gclk));
	jdff dff_A_3OkWTd0k6_0(.dout(w_dff_A_9GEjySGP9_0),.din(w_dff_A_3OkWTd0k6_0),.clk(gclk));
	jdff dff_A_9GEjySGP9_0(.dout(w_dff_A_6L2J0ckt4_0),.din(w_dff_A_9GEjySGP9_0),.clk(gclk));
	jdff dff_A_6L2J0ckt4_0(.dout(w_dff_A_d7O9XkWb9_0),.din(w_dff_A_6L2J0ckt4_0),.clk(gclk));
	jdff dff_A_d7O9XkWb9_0(.dout(w_dff_A_YkeI5BVx7_0),.din(w_dff_A_d7O9XkWb9_0),.clk(gclk));
	jdff dff_A_YkeI5BVx7_0(.dout(w_dff_A_bEXsGrKu1_0),.din(w_dff_A_YkeI5BVx7_0),.clk(gclk));
	jdff dff_A_bEXsGrKu1_0(.dout(w_dff_A_6sDJd9sI2_0),.din(w_dff_A_bEXsGrKu1_0),.clk(gclk));
	jdff dff_A_6sDJd9sI2_0(.dout(w_dff_A_0DwipA3O4_0),.din(w_dff_A_6sDJd9sI2_0),.clk(gclk));
	jdff dff_A_0DwipA3O4_0(.dout(w_dff_A_zYuQYnx05_0),.din(w_dff_A_0DwipA3O4_0),.clk(gclk));
	jdff dff_A_zYuQYnx05_0(.dout(w_dff_A_aT5uoKTe2_0),.din(w_dff_A_zYuQYnx05_0),.clk(gclk));
	jdff dff_A_aT5uoKTe2_0(.dout(w_dff_A_HovGehEh4_0),.din(w_dff_A_aT5uoKTe2_0),.clk(gclk));
	jdff dff_A_HovGehEh4_0(.dout(w_dff_A_2awL2d8H3_0),.din(w_dff_A_HovGehEh4_0),.clk(gclk));
	jdff dff_A_2awL2d8H3_0(.dout(w_dff_A_B2zJ4YEZ0_0),.din(w_dff_A_2awL2d8H3_0),.clk(gclk));
	jdff dff_A_B2zJ4YEZ0_0(.dout(w_dff_A_uvOoS5l04_0),.din(w_dff_A_B2zJ4YEZ0_0),.clk(gclk));
	jdff dff_A_uvOoS5l04_0(.dout(w_dff_A_KjUKImIS3_0),.din(w_dff_A_uvOoS5l04_0),.clk(gclk));
	jdff dff_A_KjUKImIS3_0(.dout(w_dff_A_WHok27LG9_0),.din(w_dff_A_KjUKImIS3_0),.clk(gclk));
	jdff dff_A_WHok27LG9_0(.dout(w_dff_A_OL4y1KYB5_0),.din(w_dff_A_WHok27LG9_0),.clk(gclk));
	jdff dff_A_OL4y1KYB5_0(.dout(w_dff_A_wFIdRpWy9_0),.din(w_dff_A_OL4y1KYB5_0),.clk(gclk));
	jdff dff_A_wFIdRpWy9_0(.dout(w_dff_A_EAmQGzpo5_0),.din(w_dff_A_wFIdRpWy9_0),.clk(gclk));
	jdff dff_A_EAmQGzpo5_0(.dout(w_dff_A_OAfYR3df3_0),.din(w_dff_A_EAmQGzpo5_0),.clk(gclk));
	jdff dff_A_OAfYR3df3_0(.dout(w_dff_A_iFBZSlSi9_0),.din(w_dff_A_OAfYR3df3_0),.clk(gclk));
	jdff dff_A_iFBZSlSi9_0(.dout(w_dff_A_oThtbLix2_0),.din(w_dff_A_iFBZSlSi9_0),.clk(gclk));
	jdff dff_A_oThtbLix2_0(.dout(w_dff_A_umplgO0A1_0),.din(w_dff_A_oThtbLix2_0),.clk(gclk));
	jdff dff_A_umplgO0A1_0(.dout(G973),.din(w_dff_A_umplgO0A1_0),.clk(gclk));
	jdff dff_A_qxuufKM28_1(.dout(w_dff_A_B7dVYRKr2_0),.din(w_dff_A_qxuufKM28_1),.clk(gclk));
	jdff dff_A_B7dVYRKr2_0(.dout(w_dff_A_tnOYKNRe1_0),.din(w_dff_A_B7dVYRKr2_0),.clk(gclk));
	jdff dff_A_tnOYKNRe1_0(.dout(w_dff_A_eKUyWfJJ8_0),.din(w_dff_A_tnOYKNRe1_0),.clk(gclk));
	jdff dff_A_eKUyWfJJ8_0(.dout(w_dff_A_ilHvDOjW2_0),.din(w_dff_A_eKUyWfJJ8_0),.clk(gclk));
	jdff dff_A_ilHvDOjW2_0(.dout(w_dff_A_3a6uZq8s0_0),.din(w_dff_A_ilHvDOjW2_0),.clk(gclk));
	jdff dff_A_3a6uZq8s0_0(.dout(w_dff_A_rFnpqvyo8_0),.din(w_dff_A_3a6uZq8s0_0),.clk(gclk));
	jdff dff_A_rFnpqvyo8_0(.dout(w_dff_A_v5QSkWTu4_0),.din(w_dff_A_rFnpqvyo8_0),.clk(gclk));
	jdff dff_A_v5QSkWTu4_0(.dout(w_dff_A_YnAczJ0q1_0),.din(w_dff_A_v5QSkWTu4_0),.clk(gclk));
	jdff dff_A_YnAczJ0q1_0(.dout(w_dff_A_XpSlgmas0_0),.din(w_dff_A_YnAczJ0q1_0),.clk(gclk));
	jdff dff_A_XpSlgmas0_0(.dout(w_dff_A_adib1pqi5_0),.din(w_dff_A_XpSlgmas0_0),.clk(gclk));
	jdff dff_A_adib1pqi5_0(.dout(w_dff_A_Y5NX0GwP9_0),.din(w_dff_A_adib1pqi5_0),.clk(gclk));
	jdff dff_A_Y5NX0GwP9_0(.dout(w_dff_A_bS02rXEU1_0),.din(w_dff_A_Y5NX0GwP9_0),.clk(gclk));
	jdff dff_A_bS02rXEU1_0(.dout(w_dff_A_ozBu0WPf3_0),.din(w_dff_A_bS02rXEU1_0),.clk(gclk));
	jdff dff_A_ozBu0WPf3_0(.dout(w_dff_A_0LK8BBPg1_0),.din(w_dff_A_ozBu0WPf3_0),.clk(gclk));
	jdff dff_A_0LK8BBPg1_0(.dout(w_dff_A_r4RY1TO81_0),.din(w_dff_A_0LK8BBPg1_0),.clk(gclk));
	jdff dff_A_r4RY1TO81_0(.dout(w_dff_A_yEwhhbqh6_0),.din(w_dff_A_r4RY1TO81_0),.clk(gclk));
	jdff dff_A_yEwhhbqh6_0(.dout(w_dff_A_x9vz4WlQ1_0),.din(w_dff_A_yEwhhbqh6_0),.clk(gclk));
	jdff dff_A_x9vz4WlQ1_0(.dout(w_dff_A_AaxuenLJ6_0),.din(w_dff_A_x9vz4WlQ1_0),.clk(gclk));
	jdff dff_A_AaxuenLJ6_0(.dout(w_dff_A_NtormZjw0_0),.din(w_dff_A_AaxuenLJ6_0),.clk(gclk));
	jdff dff_A_NtormZjw0_0(.dout(w_dff_A_fiIeZXGv0_0),.din(w_dff_A_NtormZjw0_0),.clk(gclk));
	jdff dff_A_fiIeZXGv0_0(.dout(w_dff_A_sC1YFJpX2_0),.din(w_dff_A_fiIeZXGv0_0),.clk(gclk));
	jdff dff_A_sC1YFJpX2_0(.dout(w_dff_A_Vyb4M1o19_0),.din(w_dff_A_sC1YFJpX2_0),.clk(gclk));
	jdff dff_A_Vyb4M1o19_0(.dout(w_dff_A_gQpL75o37_0),.din(w_dff_A_Vyb4M1o19_0),.clk(gclk));
	jdff dff_A_gQpL75o37_0(.dout(w_dff_A_JtZ3ZgxX8_0),.din(w_dff_A_gQpL75o37_0),.clk(gclk));
	jdff dff_A_JtZ3ZgxX8_0(.dout(G594),.din(w_dff_A_JtZ3ZgxX8_0),.clk(gclk));
	jdff dff_A_bSb3TJii9_1(.dout(w_dff_A_o3ZVTnGo1_0),.din(w_dff_A_bSb3TJii9_1),.clk(gclk));
	jdff dff_A_o3ZVTnGo1_0(.dout(w_dff_A_Ob7uzYGM3_0),.din(w_dff_A_o3ZVTnGo1_0),.clk(gclk));
	jdff dff_A_Ob7uzYGM3_0(.dout(w_dff_A_Kyo6X4tZ2_0),.din(w_dff_A_Ob7uzYGM3_0),.clk(gclk));
	jdff dff_A_Kyo6X4tZ2_0(.dout(w_dff_A_XqtPLVJt3_0),.din(w_dff_A_Kyo6X4tZ2_0),.clk(gclk));
	jdff dff_A_XqtPLVJt3_0(.dout(w_dff_A_vOj6XkBM0_0),.din(w_dff_A_XqtPLVJt3_0),.clk(gclk));
	jdff dff_A_vOj6XkBM0_0(.dout(w_dff_A_SY02V9pO7_0),.din(w_dff_A_vOj6XkBM0_0),.clk(gclk));
	jdff dff_A_SY02V9pO7_0(.dout(w_dff_A_0309OFbp7_0),.din(w_dff_A_SY02V9pO7_0),.clk(gclk));
	jdff dff_A_0309OFbp7_0(.dout(w_dff_A_2sBjf7r18_0),.din(w_dff_A_0309OFbp7_0),.clk(gclk));
	jdff dff_A_2sBjf7r18_0(.dout(w_dff_A_62MvLBeq7_0),.din(w_dff_A_2sBjf7r18_0),.clk(gclk));
	jdff dff_A_62MvLBeq7_0(.dout(w_dff_A_eEo3fZPx2_0),.din(w_dff_A_62MvLBeq7_0),.clk(gclk));
	jdff dff_A_eEo3fZPx2_0(.dout(w_dff_A_BczQ3AWs6_0),.din(w_dff_A_eEo3fZPx2_0),.clk(gclk));
	jdff dff_A_BczQ3AWs6_0(.dout(w_dff_A_iw4eHbsx8_0),.din(w_dff_A_BczQ3AWs6_0),.clk(gclk));
	jdff dff_A_iw4eHbsx8_0(.dout(w_dff_A_3zl7JXeM4_0),.din(w_dff_A_iw4eHbsx8_0),.clk(gclk));
	jdff dff_A_3zl7JXeM4_0(.dout(w_dff_A_DZSzWZbQ3_0),.din(w_dff_A_3zl7JXeM4_0),.clk(gclk));
	jdff dff_A_DZSzWZbQ3_0(.dout(w_dff_A_VBEpL0Q74_0),.din(w_dff_A_DZSzWZbQ3_0),.clk(gclk));
	jdff dff_A_VBEpL0Q74_0(.dout(w_dff_A_ShwZ0unR9_0),.din(w_dff_A_VBEpL0Q74_0),.clk(gclk));
	jdff dff_A_ShwZ0unR9_0(.dout(w_dff_A_zRVTRC1R6_0),.din(w_dff_A_ShwZ0unR9_0),.clk(gclk));
	jdff dff_A_zRVTRC1R6_0(.dout(w_dff_A_Epg5lDUC8_0),.din(w_dff_A_zRVTRC1R6_0),.clk(gclk));
	jdff dff_A_Epg5lDUC8_0(.dout(w_dff_A_ka3hEXUS8_0),.din(w_dff_A_Epg5lDUC8_0),.clk(gclk));
	jdff dff_A_ka3hEXUS8_0(.dout(w_dff_A_ozr4ErDd0_0),.din(w_dff_A_ka3hEXUS8_0),.clk(gclk));
	jdff dff_A_ozr4ErDd0_0(.dout(w_dff_A_A3ImSNKF3_0),.din(w_dff_A_ozr4ErDd0_0),.clk(gclk));
	jdff dff_A_A3ImSNKF3_0(.dout(w_dff_A_eLft2fKP0_0),.din(w_dff_A_A3ImSNKF3_0),.clk(gclk));
	jdff dff_A_eLft2fKP0_0(.dout(w_dff_A_Utc5zoXZ0_0),.din(w_dff_A_eLft2fKP0_0),.clk(gclk));
	jdff dff_A_Utc5zoXZ0_0(.dout(w_dff_A_KWTBCgkk7_0),.din(w_dff_A_Utc5zoXZ0_0),.clk(gclk));
	jdff dff_A_KWTBCgkk7_0(.dout(G599),.din(w_dff_A_KWTBCgkk7_0),.clk(gclk));
	jdff dff_A_1FoVNhmo2_1(.dout(w_dff_A_EqblviLa4_0),.din(w_dff_A_1FoVNhmo2_1),.clk(gclk));
	jdff dff_A_EqblviLa4_0(.dout(w_dff_A_x4dS4KNm3_0),.din(w_dff_A_EqblviLa4_0),.clk(gclk));
	jdff dff_A_x4dS4KNm3_0(.dout(w_dff_A_hxWnKqoD4_0),.din(w_dff_A_x4dS4KNm3_0),.clk(gclk));
	jdff dff_A_hxWnKqoD4_0(.dout(w_dff_A_Wk4Ua9No1_0),.din(w_dff_A_hxWnKqoD4_0),.clk(gclk));
	jdff dff_A_Wk4Ua9No1_0(.dout(w_dff_A_IfJBLCrn5_0),.din(w_dff_A_Wk4Ua9No1_0),.clk(gclk));
	jdff dff_A_IfJBLCrn5_0(.dout(w_dff_A_Hi1DSY4q7_0),.din(w_dff_A_IfJBLCrn5_0),.clk(gclk));
	jdff dff_A_Hi1DSY4q7_0(.dout(w_dff_A_VN4bPgD34_0),.din(w_dff_A_Hi1DSY4q7_0),.clk(gclk));
	jdff dff_A_VN4bPgD34_0(.dout(w_dff_A_QFRhVDnB1_0),.din(w_dff_A_VN4bPgD34_0),.clk(gclk));
	jdff dff_A_QFRhVDnB1_0(.dout(w_dff_A_a6f3iM4m2_0),.din(w_dff_A_QFRhVDnB1_0),.clk(gclk));
	jdff dff_A_a6f3iM4m2_0(.dout(w_dff_A_zM1NMrti9_0),.din(w_dff_A_a6f3iM4m2_0),.clk(gclk));
	jdff dff_A_zM1NMrti9_0(.dout(w_dff_A_JknuqsQ69_0),.din(w_dff_A_zM1NMrti9_0),.clk(gclk));
	jdff dff_A_JknuqsQ69_0(.dout(w_dff_A_LsD8gn9B6_0),.din(w_dff_A_JknuqsQ69_0),.clk(gclk));
	jdff dff_A_LsD8gn9B6_0(.dout(w_dff_A_gYXmfC4y0_0),.din(w_dff_A_LsD8gn9B6_0),.clk(gclk));
	jdff dff_A_gYXmfC4y0_0(.dout(w_dff_A_FYUnYbAd7_0),.din(w_dff_A_gYXmfC4y0_0),.clk(gclk));
	jdff dff_A_FYUnYbAd7_0(.dout(w_dff_A_xXXvQaTo4_0),.din(w_dff_A_FYUnYbAd7_0),.clk(gclk));
	jdff dff_A_xXXvQaTo4_0(.dout(w_dff_A_jmcsJKy64_0),.din(w_dff_A_xXXvQaTo4_0),.clk(gclk));
	jdff dff_A_jmcsJKy64_0(.dout(w_dff_A_UzYq3r1H0_0),.din(w_dff_A_jmcsJKy64_0),.clk(gclk));
	jdff dff_A_UzYq3r1H0_0(.dout(w_dff_A_LnHxCXJN1_0),.din(w_dff_A_UzYq3r1H0_0),.clk(gclk));
	jdff dff_A_LnHxCXJN1_0(.dout(w_dff_A_Y4Qr51QY6_0),.din(w_dff_A_LnHxCXJN1_0),.clk(gclk));
	jdff dff_A_Y4Qr51QY6_0(.dout(w_dff_A_BjHHcAUc2_0),.din(w_dff_A_Y4Qr51QY6_0),.clk(gclk));
	jdff dff_A_BjHHcAUc2_0(.dout(w_dff_A_eEV9Abv68_0),.din(w_dff_A_BjHHcAUc2_0),.clk(gclk));
	jdff dff_A_eEV9Abv68_0(.dout(w_dff_A_Y17b1LG46_0),.din(w_dff_A_eEV9Abv68_0),.clk(gclk));
	jdff dff_A_Y17b1LG46_0(.dout(w_dff_A_ItoGbDu54_0),.din(w_dff_A_Y17b1LG46_0),.clk(gclk));
	jdff dff_A_ItoGbDu54_0(.dout(w_dff_A_FSHB2BVx2_0),.din(w_dff_A_ItoGbDu54_0),.clk(gclk));
	jdff dff_A_FSHB2BVx2_0(.dout(G600),.din(w_dff_A_FSHB2BVx2_0),.clk(gclk));
	jdff dff_A_5HCiJFb58_1(.dout(w_dff_A_xrcT79jh6_0),.din(w_dff_A_5HCiJFb58_1),.clk(gclk));
	jdff dff_A_xrcT79jh6_0(.dout(w_dff_A_cSNY9F118_0),.din(w_dff_A_xrcT79jh6_0),.clk(gclk));
	jdff dff_A_cSNY9F118_0(.dout(w_dff_A_tZ4QfeYo2_0),.din(w_dff_A_cSNY9F118_0),.clk(gclk));
	jdff dff_A_tZ4QfeYo2_0(.dout(w_dff_A_xMth6Vab5_0),.din(w_dff_A_tZ4QfeYo2_0),.clk(gclk));
	jdff dff_A_xMth6Vab5_0(.dout(w_dff_A_k72Yj2Ya3_0),.din(w_dff_A_xMth6Vab5_0),.clk(gclk));
	jdff dff_A_k72Yj2Ya3_0(.dout(w_dff_A_YBrByc0o2_0),.din(w_dff_A_k72Yj2Ya3_0),.clk(gclk));
	jdff dff_A_YBrByc0o2_0(.dout(w_dff_A_zEBEAsmK3_0),.din(w_dff_A_YBrByc0o2_0),.clk(gclk));
	jdff dff_A_zEBEAsmK3_0(.dout(w_dff_A_grbhomvc9_0),.din(w_dff_A_zEBEAsmK3_0),.clk(gclk));
	jdff dff_A_grbhomvc9_0(.dout(w_dff_A_qYBpGPHq2_0),.din(w_dff_A_grbhomvc9_0),.clk(gclk));
	jdff dff_A_qYBpGPHq2_0(.dout(w_dff_A_ucFCkGzM2_0),.din(w_dff_A_qYBpGPHq2_0),.clk(gclk));
	jdff dff_A_ucFCkGzM2_0(.dout(w_dff_A_hakhRnzV9_0),.din(w_dff_A_ucFCkGzM2_0),.clk(gclk));
	jdff dff_A_hakhRnzV9_0(.dout(w_dff_A_n0IMI8yt8_0),.din(w_dff_A_hakhRnzV9_0),.clk(gclk));
	jdff dff_A_n0IMI8yt8_0(.dout(w_dff_A_QXgVB1VL2_0),.din(w_dff_A_n0IMI8yt8_0),.clk(gclk));
	jdff dff_A_QXgVB1VL2_0(.dout(w_dff_A_dKeolqRn3_0),.din(w_dff_A_QXgVB1VL2_0),.clk(gclk));
	jdff dff_A_dKeolqRn3_0(.dout(w_dff_A_3I87KtaD1_0),.din(w_dff_A_dKeolqRn3_0),.clk(gclk));
	jdff dff_A_3I87KtaD1_0(.dout(w_dff_A_MqNN865V1_0),.din(w_dff_A_3I87KtaD1_0),.clk(gclk));
	jdff dff_A_MqNN865V1_0(.dout(w_dff_A_ty9njzzq6_0),.din(w_dff_A_MqNN865V1_0),.clk(gclk));
	jdff dff_A_ty9njzzq6_0(.dout(w_dff_A_jYMPg27r9_0),.din(w_dff_A_ty9njzzq6_0),.clk(gclk));
	jdff dff_A_jYMPg27r9_0(.dout(w_dff_A_FxqWgxyw8_0),.din(w_dff_A_jYMPg27r9_0),.clk(gclk));
	jdff dff_A_FxqWgxyw8_0(.dout(w_dff_A_YJvCoOxH3_0),.din(w_dff_A_FxqWgxyw8_0),.clk(gclk));
	jdff dff_A_YJvCoOxH3_0(.dout(w_dff_A_HDhPVR4P6_0),.din(w_dff_A_YJvCoOxH3_0),.clk(gclk));
	jdff dff_A_HDhPVR4P6_0(.dout(w_dff_A_ue5fVz9Y1_0),.din(w_dff_A_HDhPVR4P6_0),.clk(gclk));
	jdff dff_A_ue5fVz9Y1_0(.dout(w_dff_A_hx8webFW0_0),.din(w_dff_A_ue5fVz9Y1_0),.clk(gclk));
	jdff dff_A_hx8webFW0_0(.dout(w_dff_A_vStQhvT93_0),.din(w_dff_A_hx8webFW0_0),.clk(gclk));
	jdff dff_A_vStQhvT93_0(.dout(G601),.din(w_dff_A_vStQhvT93_0),.clk(gclk));
	jdff dff_A_aQkG8FTE9_1(.dout(w_dff_A_yECJxp9H1_0),.din(w_dff_A_aQkG8FTE9_1),.clk(gclk));
	jdff dff_A_yECJxp9H1_0(.dout(w_dff_A_H1xXD0rB6_0),.din(w_dff_A_yECJxp9H1_0),.clk(gclk));
	jdff dff_A_H1xXD0rB6_0(.dout(w_dff_A_zYHP0WZh3_0),.din(w_dff_A_H1xXD0rB6_0),.clk(gclk));
	jdff dff_A_zYHP0WZh3_0(.dout(w_dff_A_uenPKdjy2_0),.din(w_dff_A_zYHP0WZh3_0),.clk(gclk));
	jdff dff_A_uenPKdjy2_0(.dout(w_dff_A_F42ENXhK8_0),.din(w_dff_A_uenPKdjy2_0),.clk(gclk));
	jdff dff_A_F42ENXhK8_0(.dout(w_dff_A_CWHT7mns5_0),.din(w_dff_A_F42ENXhK8_0),.clk(gclk));
	jdff dff_A_CWHT7mns5_0(.dout(w_dff_A_wKd1hncY2_0),.din(w_dff_A_CWHT7mns5_0),.clk(gclk));
	jdff dff_A_wKd1hncY2_0(.dout(w_dff_A_0cuR7wp02_0),.din(w_dff_A_wKd1hncY2_0),.clk(gclk));
	jdff dff_A_0cuR7wp02_0(.dout(w_dff_A_pyZpVygc5_0),.din(w_dff_A_0cuR7wp02_0),.clk(gclk));
	jdff dff_A_pyZpVygc5_0(.dout(w_dff_A_DfJK21kO9_0),.din(w_dff_A_pyZpVygc5_0),.clk(gclk));
	jdff dff_A_DfJK21kO9_0(.dout(w_dff_A_vVjsGcHC3_0),.din(w_dff_A_DfJK21kO9_0),.clk(gclk));
	jdff dff_A_vVjsGcHC3_0(.dout(w_dff_A_Mq5LqRSY2_0),.din(w_dff_A_vVjsGcHC3_0),.clk(gclk));
	jdff dff_A_Mq5LqRSY2_0(.dout(w_dff_A_r7wCzyxi5_0),.din(w_dff_A_Mq5LqRSY2_0),.clk(gclk));
	jdff dff_A_r7wCzyxi5_0(.dout(w_dff_A_arbtq3m29_0),.din(w_dff_A_r7wCzyxi5_0),.clk(gclk));
	jdff dff_A_arbtq3m29_0(.dout(w_dff_A_vXx1Mv7l5_0),.din(w_dff_A_arbtq3m29_0),.clk(gclk));
	jdff dff_A_vXx1Mv7l5_0(.dout(w_dff_A_oJshd60A7_0),.din(w_dff_A_vXx1Mv7l5_0),.clk(gclk));
	jdff dff_A_oJshd60A7_0(.dout(w_dff_A_wxZOrlqw9_0),.din(w_dff_A_oJshd60A7_0),.clk(gclk));
	jdff dff_A_wxZOrlqw9_0(.dout(w_dff_A_Tc8TjFDV1_0),.din(w_dff_A_wxZOrlqw9_0),.clk(gclk));
	jdff dff_A_Tc8TjFDV1_0(.dout(w_dff_A_9XjoMj7o2_0),.din(w_dff_A_Tc8TjFDV1_0),.clk(gclk));
	jdff dff_A_9XjoMj7o2_0(.dout(w_dff_A_dpQPqRNB4_0),.din(w_dff_A_9XjoMj7o2_0),.clk(gclk));
	jdff dff_A_dpQPqRNB4_0(.dout(w_dff_A_r9dDJkmY5_0),.din(w_dff_A_dpQPqRNB4_0),.clk(gclk));
	jdff dff_A_r9dDJkmY5_0(.dout(w_dff_A_RioAGGVx9_0),.din(w_dff_A_r9dDJkmY5_0),.clk(gclk));
	jdff dff_A_RioAGGVx9_0(.dout(w_dff_A_siWcFYow7_0),.din(w_dff_A_RioAGGVx9_0),.clk(gclk));
	jdff dff_A_siWcFYow7_0(.dout(w_dff_A_ucmJ6k8S5_0),.din(w_dff_A_siWcFYow7_0),.clk(gclk));
	jdff dff_A_ucmJ6k8S5_0(.dout(G602),.din(w_dff_A_ucmJ6k8S5_0),.clk(gclk));
	jdff dff_A_gr7tdRmi6_1(.dout(w_dff_A_hBn5ttdH3_0),.din(w_dff_A_gr7tdRmi6_1),.clk(gclk));
	jdff dff_A_hBn5ttdH3_0(.dout(w_dff_A_gDl5Fn464_0),.din(w_dff_A_hBn5ttdH3_0),.clk(gclk));
	jdff dff_A_gDl5Fn464_0(.dout(w_dff_A_Ve6aCRAt1_0),.din(w_dff_A_gDl5Fn464_0),.clk(gclk));
	jdff dff_A_Ve6aCRAt1_0(.dout(w_dff_A_aWUn4EZ20_0),.din(w_dff_A_Ve6aCRAt1_0),.clk(gclk));
	jdff dff_A_aWUn4EZ20_0(.dout(w_dff_A_NLzJa5X31_0),.din(w_dff_A_aWUn4EZ20_0),.clk(gclk));
	jdff dff_A_NLzJa5X31_0(.dout(w_dff_A_jVfIlE819_0),.din(w_dff_A_NLzJa5X31_0),.clk(gclk));
	jdff dff_A_jVfIlE819_0(.dout(w_dff_A_hQJdSSje8_0),.din(w_dff_A_jVfIlE819_0),.clk(gclk));
	jdff dff_A_hQJdSSje8_0(.dout(w_dff_A_ONpbsbqp3_0),.din(w_dff_A_hQJdSSje8_0),.clk(gclk));
	jdff dff_A_ONpbsbqp3_0(.dout(w_dff_A_swmwDC7v6_0),.din(w_dff_A_ONpbsbqp3_0),.clk(gclk));
	jdff dff_A_swmwDC7v6_0(.dout(w_dff_A_9xAhxXP04_0),.din(w_dff_A_swmwDC7v6_0),.clk(gclk));
	jdff dff_A_9xAhxXP04_0(.dout(w_dff_A_MqvQPcUc6_0),.din(w_dff_A_9xAhxXP04_0),.clk(gclk));
	jdff dff_A_MqvQPcUc6_0(.dout(w_dff_A_gI361zfA6_0),.din(w_dff_A_MqvQPcUc6_0),.clk(gclk));
	jdff dff_A_gI361zfA6_0(.dout(w_dff_A_IapgDGrg0_0),.din(w_dff_A_gI361zfA6_0),.clk(gclk));
	jdff dff_A_IapgDGrg0_0(.dout(w_dff_A_81dyt1Uy2_0),.din(w_dff_A_IapgDGrg0_0),.clk(gclk));
	jdff dff_A_81dyt1Uy2_0(.dout(w_dff_A_RRZIrERw8_0),.din(w_dff_A_81dyt1Uy2_0),.clk(gclk));
	jdff dff_A_RRZIrERw8_0(.dout(w_dff_A_oZToYoLD5_0),.din(w_dff_A_RRZIrERw8_0),.clk(gclk));
	jdff dff_A_oZToYoLD5_0(.dout(w_dff_A_a78YLMOZ7_0),.din(w_dff_A_oZToYoLD5_0),.clk(gclk));
	jdff dff_A_a78YLMOZ7_0(.dout(w_dff_A_WQaws6Ie6_0),.din(w_dff_A_a78YLMOZ7_0),.clk(gclk));
	jdff dff_A_WQaws6Ie6_0(.dout(w_dff_A_OcsYoPst5_0),.din(w_dff_A_WQaws6Ie6_0),.clk(gclk));
	jdff dff_A_OcsYoPst5_0(.dout(w_dff_A_rtFC0nVv9_0),.din(w_dff_A_OcsYoPst5_0),.clk(gclk));
	jdff dff_A_rtFC0nVv9_0(.dout(w_dff_A_LGPgYbvx0_0),.din(w_dff_A_rtFC0nVv9_0),.clk(gclk));
	jdff dff_A_LGPgYbvx0_0(.dout(w_dff_A_nnq9LSC41_0),.din(w_dff_A_LGPgYbvx0_0),.clk(gclk));
	jdff dff_A_nnq9LSC41_0(.dout(w_dff_A_4etVxjX29_0),.din(w_dff_A_nnq9LSC41_0),.clk(gclk));
	jdff dff_A_4etVxjX29_0(.dout(w_dff_A_oVV3ENCY3_0),.din(w_dff_A_4etVxjX29_0),.clk(gclk));
	jdff dff_A_oVV3ENCY3_0(.dout(G603),.din(w_dff_A_oVV3ENCY3_0),.clk(gclk));
	jdff dff_A_OUjptODI7_1(.dout(w_dff_A_plwWFb4D4_0),.din(w_dff_A_OUjptODI7_1),.clk(gclk));
	jdff dff_A_plwWFb4D4_0(.dout(w_dff_A_b7aZoJ4a6_0),.din(w_dff_A_plwWFb4D4_0),.clk(gclk));
	jdff dff_A_b7aZoJ4a6_0(.dout(w_dff_A_URFVMIDc3_0),.din(w_dff_A_b7aZoJ4a6_0),.clk(gclk));
	jdff dff_A_URFVMIDc3_0(.dout(w_dff_A_McK0uXlW5_0),.din(w_dff_A_URFVMIDc3_0),.clk(gclk));
	jdff dff_A_McK0uXlW5_0(.dout(w_dff_A_i5qE0GQn1_0),.din(w_dff_A_McK0uXlW5_0),.clk(gclk));
	jdff dff_A_i5qE0GQn1_0(.dout(w_dff_A_POdY9Rtj7_0),.din(w_dff_A_i5qE0GQn1_0),.clk(gclk));
	jdff dff_A_POdY9Rtj7_0(.dout(w_dff_A_6dNJKmMS2_0),.din(w_dff_A_POdY9Rtj7_0),.clk(gclk));
	jdff dff_A_6dNJKmMS2_0(.dout(w_dff_A_Yln3uv1E0_0),.din(w_dff_A_6dNJKmMS2_0),.clk(gclk));
	jdff dff_A_Yln3uv1E0_0(.dout(w_dff_A_4bv8kuBe7_0),.din(w_dff_A_Yln3uv1E0_0),.clk(gclk));
	jdff dff_A_4bv8kuBe7_0(.dout(w_dff_A_masqWA0e1_0),.din(w_dff_A_4bv8kuBe7_0),.clk(gclk));
	jdff dff_A_masqWA0e1_0(.dout(w_dff_A_nMyXoepL7_0),.din(w_dff_A_masqWA0e1_0),.clk(gclk));
	jdff dff_A_nMyXoepL7_0(.dout(w_dff_A_NvlA8NfG9_0),.din(w_dff_A_nMyXoepL7_0),.clk(gclk));
	jdff dff_A_NvlA8NfG9_0(.dout(w_dff_A_dqIuYJhf9_0),.din(w_dff_A_NvlA8NfG9_0),.clk(gclk));
	jdff dff_A_dqIuYJhf9_0(.dout(w_dff_A_d8sPpaa22_0),.din(w_dff_A_dqIuYJhf9_0),.clk(gclk));
	jdff dff_A_d8sPpaa22_0(.dout(w_dff_A_pCTziFrW5_0),.din(w_dff_A_d8sPpaa22_0),.clk(gclk));
	jdff dff_A_pCTziFrW5_0(.dout(w_dff_A_NddNnJEM5_0),.din(w_dff_A_pCTziFrW5_0),.clk(gclk));
	jdff dff_A_NddNnJEM5_0(.dout(w_dff_A_lmun7lGa6_0),.din(w_dff_A_NddNnJEM5_0),.clk(gclk));
	jdff dff_A_lmun7lGa6_0(.dout(w_dff_A_gfvOh1a45_0),.din(w_dff_A_lmun7lGa6_0),.clk(gclk));
	jdff dff_A_gfvOh1a45_0(.dout(w_dff_A_qUjReKbK7_0),.din(w_dff_A_gfvOh1a45_0),.clk(gclk));
	jdff dff_A_qUjReKbK7_0(.dout(w_dff_A_oO653SGZ4_0),.din(w_dff_A_qUjReKbK7_0),.clk(gclk));
	jdff dff_A_oO653SGZ4_0(.dout(w_dff_A_N4EMP4Qv4_0),.din(w_dff_A_oO653SGZ4_0),.clk(gclk));
	jdff dff_A_N4EMP4Qv4_0(.dout(w_dff_A_16pNIE2M8_0),.din(w_dff_A_N4EMP4Qv4_0),.clk(gclk));
	jdff dff_A_16pNIE2M8_0(.dout(w_dff_A_A1ul20vT2_0),.din(w_dff_A_16pNIE2M8_0),.clk(gclk));
	jdff dff_A_A1ul20vT2_0(.dout(w_dff_A_IttKCy8j5_0),.din(w_dff_A_A1ul20vT2_0),.clk(gclk));
	jdff dff_A_IttKCy8j5_0(.dout(G604),.din(w_dff_A_IttKCy8j5_0),.clk(gclk));
	jdff dff_A_FJjvtOnm3_1(.dout(w_dff_A_YSYzDgDs9_0),.din(w_dff_A_FJjvtOnm3_1),.clk(gclk));
	jdff dff_A_YSYzDgDs9_0(.dout(w_dff_A_xMWjtSNp1_0),.din(w_dff_A_YSYzDgDs9_0),.clk(gclk));
	jdff dff_A_xMWjtSNp1_0(.dout(w_dff_A_yKytuZkK8_0),.din(w_dff_A_xMWjtSNp1_0),.clk(gclk));
	jdff dff_A_yKytuZkK8_0(.dout(w_dff_A_chnn2FVy3_0),.din(w_dff_A_yKytuZkK8_0),.clk(gclk));
	jdff dff_A_chnn2FVy3_0(.dout(w_dff_A_hSLVk3pN7_0),.din(w_dff_A_chnn2FVy3_0),.clk(gclk));
	jdff dff_A_hSLVk3pN7_0(.dout(w_dff_A_KvJrlhri3_0),.din(w_dff_A_hSLVk3pN7_0),.clk(gclk));
	jdff dff_A_KvJrlhri3_0(.dout(w_dff_A_46m0Oqh99_0),.din(w_dff_A_KvJrlhri3_0),.clk(gclk));
	jdff dff_A_46m0Oqh99_0(.dout(w_dff_A_y7Mq608C2_0),.din(w_dff_A_46m0Oqh99_0),.clk(gclk));
	jdff dff_A_y7Mq608C2_0(.dout(w_dff_A_xVLCQ4Ec3_0),.din(w_dff_A_y7Mq608C2_0),.clk(gclk));
	jdff dff_A_xVLCQ4Ec3_0(.dout(w_dff_A_fyj0MEvt2_0),.din(w_dff_A_xVLCQ4Ec3_0),.clk(gclk));
	jdff dff_A_fyj0MEvt2_0(.dout(w_dff_A_ysNRlxUY1_0),.din(w_dff_A_fyj0MEvt2_0),.clk(gclk));
	jdff dff_A_ysNRlxUY1_0(.dout(w_dff_A_zsvlQMd40_0),.din(w_dff_A_ysNRlxUY1_0),.clk(gclk));
	jdff dff_A_zsvlQMd40_0(.dout(w_dff_A_vy9FQOrt1_0),.din(w_dff_A_zsvlQMd40_0),.clk(gclk));
	jdff dff_A_vy9FQOrt1_0(.dout(w_dff_A_pzE5bXhX1_0),.din(w_dff_A_vy9FQOrt1_0),.clk(gclk));
	jdff dff_A_pzE5bXhX1_0(.dout(w_dff_A_hZRFcWxc3_0),.din(w_dff_A_pzE5bXhX1_0),.clk(gclk));
	jdff dff_A_hZRFcWxc3_0(.dout(w_dff_A_24ox9GgO9_0),.din(w_dff_A_hZRFcWxc3_0),.clk(gclk));
	jdff dff_A_24ox9GgO9_0(.dout(w_dff_A_S2ARY1D45_0),.din(w_dff_A_24ox9GgO9_0),.clk(gclk));
	jdff dff_A_S2ARY1D45_0(.dout(w_dff_A_rovhe0RP3_0),.din(w_dff_A_S2ARY1D45_0),.clk(gclk));
	jdff dff_A_rovhe0RP3_0(.dout(w_dff_A_aRQobSYC4_0),.din(w_dff_A_rovhe0RP3_0),.clk(gclk));
	jdff dff_A_aRQobSYC4_0(.dout(w_dff_A_zTDctRW94_0),.din(w_dff_A_aRQobSYC4_0),.clk(gclk));
	jdff dff_A_zTDctRW94_0(.dout(w_dff_A_1ZrL74WM5_0),.din(w_dff_A_zTDctRW94_0),.clk(gclk));
	jdff dff_A_1ZrL74WM5_0(.dout(w_dff_A_lwp0zlzh8_0),.din(w_dff_A_1ZrL74WM5_0),.clk(gclk));
	jdff dff_A_lwp0zlzh8_0(.dout(w_dff_A_y6xwCR5I3_0),.din(w_dff_A_lwp0zlzh8_0),.clk(gclk));
	jdff dff_A_y6xwCR5I3_0(.dout(w_dff_A_NhO4xXpN6_0),.din(w_dff_A_y6xwCR5I3_0),.clk(gclk));
	jdff dff_A_NhO4xXpN6_0(.dout(G611),.din(w_dff_A_NhO4xXpN6_0),.clk(gclk));
	jdff dff_A_HPCQADGE6_1(.dout(w_dff_A_aLCa9vOG5_0),.din(w_dff_A_HPCQADGE6_1),.clk(gclk));
	jdff dff_A_aLCa9vOG5_0(.dout(w_dff_A_NDprfOMW5_0),.din(w_dff_A_aLCa9vOG5_0),.clk(gclk));
	jdff dff_A_NDprfOMW5_0(.dout(w_dff_A_ESlHrX7O2_0),.din(w_dff_A_NDprfOMW5_0),.clk(gclk));
	jdff dff_A_ESlHrX7O2_0(.dout(w_dff_A_8yHfk8Mw6_0),.din(w_dff_A_ESlHrX7O2_0),.clk(gclk));
	jdff dff_A_8yHfk8Mw6_0(.dout(w_dff_A_QKp91s2h2_0),.din(w_dff_A_8yHfk8Mw6_0),.clk(gclk));
	jdff dff_A_QKp91s2h2_0(.dout(w_dff_A_L0ThTLBV3_0),.din(w_dff_A_QKp91s2h2_0),.clk(gclk));
	jdff dff_A_L0ThTLBV3_0(.dout(w_dff_A_G7Zt6O8T7_0),.din(w_dff_A_L0ThTLBV3_0),.clk(gclk));
	jdff dff_A_G7Zt6O8T7_0(.dout(w_dff_A_hgnZjgYK5_0),.din(w_dff_A_G7Zt6O8T7_0),.clk(gclk));
	jdff dff_A_hgnZjgYK5_0(.dout(w_dff_A_SfblFLUk0_0),.din(w_dff_A_hgnZjgYK5_0),.clk(gclk));
	jdff dff_A_SfblFLUk0_0(.dout(w_dff_A_64hgeVf47_0),.din(w_dff_A_SfblFLUk0_0),.clk(gclk));
	jdff dff_A_64hgeVf47_0(.dout(w_dff_A_ETNdEqhN5_0),.din(w_dff_A_64hgeVf47_0),.clk(gclk));
	jdff dff_A_ETNdEqhN5_0(.dout(w_dff_A_zbdnEx7K1_0),.din(w_dff_A_ETNdEqhN5_0),.clk(gclk));
	jdff dff_A_zbdnEx7K1_0(.dout(w_dff_A_22EscIR99_0),.din(w_dff_A_zbdnEx7K1_0),.clk(gclk));
	jdff dff_A_22EscIR99_0(.dout(w_dff_A_a8aItw0v3_0),.din(w_dff_A_22EscIR99_0),.clk(gclk));
	jdff dff_A_a8aItw0v3_0(.dout(w_dff_A_5kpXoC1t2_0),.din(w_dff_A_a8aItw0v3_0),.clk(gclk));
	jdff dff_A_5kpXoC1t2_0(.dout(w_dff_A_EHeaxokn1_0),.din(w_dff_A_5kpXoC1t2_0),.clk(gclk));
	jdff dff_A_EHeaxokn1_0(.dout(w_dff_A_wZR2sSl97_0),.din(w_dff_A_EHeaxokn1_0),.clk(gclk));
	jdff dff_A_wZR2sSl97_0(.dout(w_dff_A_NavXcQAt2_0),.din(w_dff_A_wZR2sSl97_0),.clk(gclk));
	jdff dff_A_NavXcQAt2_0(.dout(w_dff_A_lhIPVIyD9_0),.din(w_dff_A_NavXcQAt2_0),.clk(gclk));
	jdff dff_A_lhIPVIyD9_0(.dout(w_dff_A_f03qnhYt6_0),.din(w_dff_A_lhIPVIyD9_0),.clk(gclk));
	jdff dff_A_f03qnhYt6_0(.dout(w_dff_A_b7yAy11t3_0),.din(w_dff_A_f03qnhYt6_0),.clk(gclk));
	jdff dff_A_b7yAy11t3_0(.dout(w_dff_A_KvEh6WsY7_0),.din(w_dff_A_b7yAy11t3_0),.clk(gclk));
	jdff dff_A_KvEh6WsY7_0(.dout(w_dff_A_OmK0mBkb3_0),.din(w_dff_A_KvEh6WsY7_0),.clk(gclk));
	jdff dff_A_OmK0mBkb3_0(.dout(w_dff_A_2svKVKTn5_0),.din(w_dff_A_OmK0mBkb3_0),.clk(gclk));
	jdff dff_A_2svKVKTn5_0(.dout(G612),.din(w_dff_A_2svKVKTn5_0),.clk(gclk));
	jdff dff_A_Tx7LCMRQ4_2(.dout(w_dff_A_14kAUU5Z8_0),.din(w_dff_A_Tx7LCMRQ4_2),.clk(gclk));
	jdff dff_A_14kAUU5Z8_0(.dout(w_dff_A_tOR2rClx1_0),.din(w_dff_A_14kAUU5Z8_0),.clk(gclk));
	jdff dff_A_tOR2rClx1_0(.dout(w_dff_A_8tKSUArA0_0),.din(w_dff_A_tOR2rClx1_0),.clk(gclk));
	jdff dff_A_8tKSUArA0_0(.dout(w_dff_A_O4WH3Moz6_0),.din(w_dff_A_8tKSUArA0_0),.clk(gclk));
	jdff dff_A_O4WH3Moz6_0(.dout(w_dff_A_qAHQIeSR5_0),.din(w_dff_A_O4WH3Moz6_0),.clk(gclk));
	jdff dff_A_qAHQIeSR5_0(.dout(w_dff_A_8R6gCynq5_0),.din(w_dff_A_qAHQIeSR5_0),.clk(gclk));
	jdff dff_A_8R6gCynq5_0(.dout(w_dff_A_GAQ4nw440_0),.din(w_dff_A_8R6gCynq5_0),.clk(gclk));
	jdff dff_A_GAQ4nw440_0(.dout(w_dff_A_otVRNlBZ3_0),.din(w_dff_A_GAQ4nw440_0),.clk(gclk));
	jdff dff_A_otVRNlBZ3_0(.dout(w_dff_A_GVJYovpm6_0),.din(w_dff_A_otVRNlBZ3_0),.clk(gclk));
	jdff dff_A_GVJYovpm6_0(.dout(w_dff_A_ba9wSJl45_0),.din(w_dff_A_GVJYovpm6_0),.clk(gclk));
	jdff dff_A_ba9wSJl45_0(.dout(w_dff_A_zwwR4PAW8_0),.din(w_dff_A_ba9wSJl45_0),.clk(gclk));
	jdff dff_A_zwwR4PAW8_0(.dout(w_dff_A_Y94x4yeA1_0),.din(w_dff_A_zwwR4PAW8_0),.clk(gclk));
	jdff dff_A_Y94x4yeA1_0(.dout(w_dff_A_Oklqd7mC8_0),.din(w_dff_A_Y94x4yeA1_0),.clk(gclk));
	jdff dff_A_Oklqd7mC8_0(.dout(w_dff_A_5kEttWOO0_0),.din(w_dff_A_Oklqd7mC8_0),.clk(gclk));
	jdff dff_A_5kEttWOO0_0(.dout(w_dff_A_jRwE7Bb38_0),.din(w_dff_A_5kEttWOO0_0),.clk(gclk));
	jdff dff_A_jRwE7Bb38_0(.dout(w_dff_A_Fxwxn6190_0),.din(w_dff_A_jRwE7Bb38_0),.clk(gclk));
	jdff dff_A_Fxwxn6190_0(.dout(w_dff_A_Nwbfqv7e6_0),.din(w_dff_A_Fxwxn6190_0),.clk(gclk));
	jdff dff_A_Nwbfqv7e6_0(.dout(w_dff_A_IUMgHBSb2_0),.din(w_dff_A_Nwbfqv7e6_0),.clk(gclk));
	jdff dff_A_IUMgHBSb2_0(.dout(w_dff_A_6RVcPaFp7_0),.din(w_dff_A_IUMgHBSb2_0),.clk(gclk));
	jdff dff_A_6RVcPaFp7_0(.dout(w_dff_A_b9U8rvN75_0),.din(w_dff_A_6RVcPaFp7_0),.clk(gclk));
	jdff dff_A_b9U8rvN75_0(.dout(w_dff_A_nOvPMse80_0),.din(w_dff_A_b9U8rvN75_0),.clk(gclk));
	jdff dff_A_nOvPMse80_0(.dout(w_dff_A_Y4c4Oc1T8_0),.din(w_dff_A_nOvPMse80_0),.clk(gclk));
	jdff dff_A_Y4c4Oc1T8_0(.dout(w_dff_A_Ogr1fN703_0),.din(w_dff_A_Y4c4Oc1T8_0),.clk(gclk));
	jdff dff_A_Ogr1fN703_0(.dout(w_dff_A_VG6Z7uxI3_0),.din(w_dff_A_Ogr1fN703_0),.clk(gclk));
	jdff dff_A_VG6Z7uxI3_0(.dout(G810),.din(w_dff_A_VG6Z7uxI3_0),.clk(gclk));
	jdff dff_A_4t5qomYy6_1(.dout(w_dff_A_JglmjN1Z4_0),.din(w_dff_A_4t5qomYy6_1),.clk(gclk));
	jdff dff_A_JglmjN1Z4_0(.dout(w_dff_A_ccemzdBD0_0),.din(w_dff_A_JglmjN1Z4_0),.clk(gclk));
	jdff dff_A_ccemzdBD0_0(.dout(w_dff_A_aCyYX4Zv1_0),.din(w_dff_A_ccemzdBD0_0),.clk(gclk));
	jdff dff_A_aCyYX4Zv1_0(.dout(w_dff_A_WfZ5zNkY2_0),.din(w_dff_A_aCyYX4Zv1_0),.clk(gclk));
	jdff dff_A_WfZ5zNkY2_0(.dout(w_dff_A_ZoDMpAIF7_0),.din(w_dff_A_WfZ5zNkY2_0),.clk(gclk));
	jdff dff_A_ZoDMpAIF7_0(.dout(w_dff_A_RPbtjc4T1_0),.din(w_dff_A_ZoDMpAIF7_0),.clk(gclk));
	jdff dff_A_RPbtjc4T1_0(.dout(w_dff_A_yNyL1sjl9_0),.din(w_dff_A_RPbtjc4T1_0),.clk(gclk));
	jdff dff_A_yNyL1sjl9_0(.dout(w_dff_A_vP5aHVhj6_0),.din(w_dff_A_yNyL1sjl9_0),.clk(gclk));
	jdff dff_A_vP5aHVhj6_0(.dout(w_dff_A_LvHLTHhK7_0),.din(w_dff_A_vP5aHVhj6_0),.clk(gclk));
	jdff dff_A_LvHLTHhK7_0(.dout(w_dff_A_dA07wt589_0),.din(w_dff_A_LvHLTHhK7_0),.clk(gclk));
	jdff dff_A_dA07wt589_0(.dout(w_dff_A_b8fij2VU1_0),.din(w_dff_A_dA07wt589_0),.clk(gclk));
	jdff dff_A_b8fij2VU1_0(.dout(w_dff_A_HZaXf0B80_0),.din(w_dff_A_b8fij2VU1_0),.clk(gclk));
	jdff dff_A_HZaXf0B80_0(.dout(w_dff_A_ntKySZrP0_0),.din(w_dff_A_HZaXf0B80_0),.clk(gclk));
	jdff dff_A_ntKySZrP0_0(.dout(w_dff_A_arLOqNh44_0),.din(w_dff_A_ntKySZrP0_0),.clk(gclk));
	jdff dff_A_arLOqNh44_0(.dout(w_dff_A_rlY5AMvy7_0),.din(w_dff_A_arLOqNh44_0),.clk(gclk));
	jdff dff_A_rlY5AMvy7_0(.dout(w_dff_A_tve4drrI3_0),.din(w_dff_A_rlY5AMvy7_0),.clk(gclk));
	jdff dff_A_tve4drrI3_0(.dout(w_dff_A_iiRJTXmZ6_0),.din(w_dff_A_tve4drrI3_0),.clk(gclk));
	jdff dff_A_iiRJTXmZ6_0(.dout(w_dff_A_LRxqIdLm7_0),.din(w_dff_A_iiRJTXmZ6_0),.clk(gclk));
	jdff dff_A_LRxqIdLm7_0(.dout(w_dff_A_9NSZLUZQ9_0),.din(w_dff_A_LRxqIdLm7_0),.clk(gclk));
	jdff dff_A_9NSZLUZQ9_0(.dout(w_dff_A_vc2SNTHS3_0),.din(w_dff_A_9NSZLUZQ9_0),.clk(gclk));
	jdff dff_A_vc2SNTHS3_0(.dout(w_dff_A_f4EUHqpe8_0),.din(w_dff_A_vc2SNTHS3_0),.clk(gclk));
	jdff dff_A_f4EUHqpe8_0(.dout(w_dff_A_vZyTu1z64_0),.din(w_dff_A_f4EUHqpe8_0),.clk(gclk));
	jdff dff_A_vZyTu1z64_0(.dout(w_dff_A_xcBrXdKy1_0),.din(w_dff_A_vZyTu1z64_0),.clk(gclk));
	jdff dff_A_xcBrXdKy1_0(.dout(w_dff_A_0ppt8fdD7_0),.din(w_dff_A_xcBrXdKy1_0),.clk(gclk));
	jdff dff_A_0ppt8fdD7_0(.dout(G848),.din(w_dff_A_0ppt8fdD7_0),.clk(gclk));
	jdff dff_A_f8vZYw3H0_1(.dout(w_dff_A_yBdxMWK71_0),.din(w_dff_A_f8vZYw3H0_1),.clk(gclk));
	jdff dff_A_yBdxMWK71_0(.dout(w_dff_A_vN1cUOXQ7_0),.din(w_dff_A_yBdxMWK71_0),.clk(gclk));
	jdff dff_A_vN1cUOXQ7_0(.dout(w_dff_A_7JvcQmRO2_0),.din(w_dff_A_vN1cUOXQ7_0),.clk(gclk));
	jdff dff_A_7JvcQmRO2_0(.dout(w_dff_A_nDuukRtl4_0),.din(w_dff_A_7JvcQmRO2_0),.clk(gclk));
	jdff dff_A_nDuukRtl4_0(.dout(w_dff_A_rKIDSq7L0_0),.din(w_dff_A_nDuukRtl4_0),.clk(gclk));
	jdff dff_A_rKIDSq7L0_0(.dout(w_dff_A_1mCManc11_0),.din(w_dff_A_rKIDSq7L0_0),.clk(gclk));
	jdff dff_A_1mCManc11_0(.dout(w_dff_A_fBWVuOqo5_0),.din(w_dff_A_1mCManc11_0),.clk(gclk));
	jdff dff_A_fBWVuOqo5_0(.dout(w_dff_A_CKKeH1dR4_0),.din(w_dff_A_fBWVuOqo5_0),.clk(gclk));
	jdff dff_A_CKKeH1dR4_0(.dout(w_dff_A_3K8EO7L29_0),.din(w_dff_A_CKKeH1dR4_0),.clk(gclk));
	jdff dff_A_3K8EO7L29_0(.dout(w_dff_A_1tByP6EO5_0),.din(w_dff_A_3K8EO7L29_0),.clk(gclk));
	jdff dff_A_1tByP6EO5_0(.dout(w_dff_A_yCCE39p71_0),.din(w_dff_A_1tByP6EO5_0),.clk(gclk));
	jdff dff_A_yCCE39p71_0(.dout(w_dff_A_wMWEL7dG6_0),.din(w_dff_A_yCCE39p71_0),.clk(gclk));
	jdff dff_A_wMWEL7dG6_0(.dout(w_dff_A_pTEvlNLI1_0),.din(w_dff_A_wMWEL7dG6_0),.clk(gclk));
	jdff dff_A_pTEvlNLI1_0(.dout(w_dff_A_cJcdngc56_0),.din(w_dff_A_pTEvlNLI1_0),.clk(gclk));
	jdff dff_A_cJcdngc56_0(.dout(w_dff_A_rlQvqZ9v0_0),.din(w_dff_A_cJcdngc56_0),.clk(gclk));
	jdff dff_A_rlQvqZ9v0_0(.dout(w_dff_A_BPeS75Ta9_0),.din(w_dff_A_rlQvqZ9v0_0),.clk(gclk));
	jdff dff_A_BPeS75Ta9_0(.dout(w_dff_A_F4V4fGZr8_0),.din(w_dff_A_BPeS75Ta9_0),.clk(gclk));
	jdff dff_A_F4V4fGZr8_0(.dout(w_dff_A_rGqMNOaA1_0),.din(w_dff_A_F4V4fGZr8_0),.clk(gclk));
	jdff dff_A_rGqMNOaA1_0(.dout(w_dff_A_cpvzZGOd5_0),.din(w_dff_A_rGqMNOaA1_0),.clk(gclk));
	jdff dff_A_cpvzZGOd5_0(.dout(w_dff_A_MtZUFIL39_0),.din(w_dff_A_cpvzZGOd5_0),.clk(gclk));
	jdff dff_A_MtZUFIL39_0(.dout(w_dff_A_EUW4a9A54_0),.din(w_dff_A_MtZUFIL39_0),.clk(gclk));
	jdff dff_A_EUW4a9A54_0(.dout(w_dff_A_zeWAjc868_0),.din(w_dff_A_EUW4a9A54_0),.clk(gclk));
	jdff dff_A_zeWAjc868_0(.dout(w_dff_A_7gTExLR42_0),.din(w_dff_A_zeWAjc868_0),.clk(gclk));
	jdff dff_A_7gTExLR42_0(.dout(w_dff_A_8T28QgsW3_0),.din(w_dff_A_7gTExLR42_0),.clk(gclk));
	jdff dff_A_8T28QgsW3_0(.dout(G849),.din(w_dff_A_8T28QgsW3_0),.clk(gclk));
	jdff dff_A_BdUBaggz8_1(.dout(w_dff_A_Iyz5s8VD6_0),.din(w_dff_A_BdUBaggz8_1),.clk(gclk));
	jdff dff_A_Iyz5s8VD6_0(.dout(w_dff_A_rJa9VwBA8_0),.din(w_dff_A_Iyz5s8VD6_0),.clk(gclk));
	jdff dff_A_rJa9VwBA8_0(.dout(w_dff_A_QVPeiX7F6_0),.din(w_dff_A_rJa9VwBA8_0),.clk(gclk));
	jdff dff_A_QVPeiX7F6_0(.dout(w_dff_A_qhyRiV6p2_0),.din(w_dff_A_QVPeiX7F6_0),.clk(gclk));
	jdff dff_A_qhyRiV6p2_0(.dout(w_dff_A_nf3YsK3B5_0),.din(w_dff_A_qhyRiV6p2_0),.clk(gclk));
	jdff dff_A_nf3YsK3B5_0(.dout(w_dff_A_vHtItjyK8_0),.din(w_dff_A_nf3YsK3B5_0),.clk(gclk));
	jdff dff_A_vHtItjyK8_0(.dout(w_dff_A_QAtxzspg8_0),.din(w_dff_A_vHtItjyK8_0),.clk(gclk));
	jdff dff_A_QAtxzspg8_0(.dout(w_dff_A_VsD6A8DB1_0),.din(w_dff_A_QAtxzspg8_0),.clk(gclk));
	jdff dff_A_VsD6A8DB1_0(.dout(w_dff_A_zqBjAU7L5_0),.din(w_dff_A_VsD6A8DB1_0),.clk(gclk));
	jdff dff_A_zqBjAU7L5_0(.dout(w_dff_A_6iaFECpC8_0),.din(w_dff_A_zqBjAU7L5_0),.clk(gclk));
	jdff dff_A_6iaFECpC8_0(.dout(w_dff_A_1dBIaVfv0_0),.din(w_dff_A_6iaFECpC8_0),.clk(gclk));
	jdff dff_A_1dBIaVfv0_0(.dout(w_dff_A_la3wU6Ia6_0),.din(w_dff_A_1dBIaVfv0_0),.clk(gclk));
	jdff dff_A_la3wU6Ia6_0(.dout(w_dff_A_UhXVFHhA6_0),.din(w_dff_A_la3wU6Ia6_0),.clk(gclk));
	jdff dff_A_UhXVFHhA6_0(.dout(w_dff_A_aSed0eb27_0),.din(w_dff_A_UhXVFHhA6_0),.clk(gclk));
	jdff dff_A_aSed0eb27_0(.dout(w_dff_A_YbUCoBjD5_0),.din(w_dff_A_aSed0eb27_0),.clk(gclk));
	jdff dff_A_YbUCoBjD5_0(.dout(w_dff_A_LRApCwlo7_0),.din(w_dff_A_YbUCoBjD5_0),.clk(gclk));
	jdff dff_A_LRApCwlo7_0(.dout(w_dff_A_2N5mlHuM8_0),.din(w_dff_A_LRApCwlo7_0),.clk(gclk));
	jdff dff_A_2N5mlHuM8_0(.dout(w_dff_A_9Y56wAhA6_0),.din(w_dff_A_2N5mlHuM8_0),.clk(gclk));
	jdff dff_A_9Y56wAhA6_0(.dout(w_dff_A_XszV9iEO3_0),.din(w_dff_A_9Y56wAhA6_0),.clk(gclk));
	jdff dff_A_XszV9iEO3_0(.dout(w_dff_A_n3Rrntqs8_0),.din(w_dff_A_XszV9iEO3_0),.clk(gclk));
	jdff dff_A_n3Rrntqs8_0(.dout(w_dff_A_u3IPBKOP0_0),.din(w_dff_A_n3Rrntqs8_0),.clk(gclk));
	jdff dff_A_u3IPBKOP0_0(.dout(w_dff_A_aKAfical2_0),.din(w_dff_A_u3IPBKOP0_0),.clk(gclk));
	jdff dff_A_aKAfical2_0(.dout(w_dff_A_AybOmuZK5_0),.din(w_dff_A_aKAfical2_0),.clk(gclk));
	jdff dff_A_AybOmuZK5_0(.dout(w_dff_A_luNwuZrr4_0),.din(w_dff_A_AybOmuZK5_0),.clk(gclk));
	jdff dff_A_luNwuZrr4_0(.dout(G850),.din(w_dff_A_luNwuZrr4_0),.clk(gclk));
	jdff dff_A_O7dZoQl30_1(.dout(w_dff_A_V1Tcj7mQ9_0),.din(w_dff_A_O7dZoQl30_1),.clk(gclk));
	jdff dff_A_V1Tcj7mQ9_0(.dout(w_dff_A_3Pi8NwzR5_0),.din(w_dff_A_V1Tcj7mQ9_0),.clk(gclk));
	jdff dff_A_3Pi8NwzR5_0(.dout(w_dff_A_OXFg8ti32_0),.din(w_dff_A_3Pi8NwzR5_0),.clk(gclk));
	jdff dff_A_OXFg8ti32_0(.dout(w_dff_A_F5iUhkOb8_0),.din(w_dff_A_OXFg8ti32_0),.clk(gclk));
	jdff dff_A_F5iUhkOb8_0(.dout(w_dff_A_wzrhIHIU7_0),.din(w_dff_A_F5iUhkOb8_0),.clk(gclk));
	jdff dff_A_wzrhIHIU7_0(.dout(w_dff_A_oSXYUSXL2_0),.din(w_dff_A_wzrhIHIU7_0),.clk(gclk));
	jdff dff_A_oSXYUSXL2_0(.dout(w_dff_A_eVhtiyi51_0),.din(w_dff_A_oSXYUSXL2_0),.clk(gclk));
	jdff dff_A_eVhtiyi51_0(.dout(w_dff_A_UAzuIQyo6_0),.din(w_dff_A_eVhtiyi51_0),.clk(gclk));
	jdff dff_A_UAzuIQyo6_0(.dout(w_dff_A_N0pLwbjx8_0),.din(w_dff_A_UAzuIQyo6_0),.clk(gclk));
	jdff dff_A_N0pLwbjx8_0(.dout(w_dff_A_PLXJVj9Y1_0),.din(w_dff_A_N0pLwbjx8_0),.clk(gclk));
	jdff dff_A_PLXJVj9Y1_0(.dout(w_dff_A_BxwhdICT1_0),.din(w_dff_A_PLXJVj9Y1_0),.clk(gclk));
	jdff dff_A_BxwhdICT1_0(.dout(w_dff_A_kP9unsOF2_0),.din(w_dff_A_BxwhdICT1_0),.clk(gclk));
	jdff dff_A_kP9unsOF2_0(.dout(w_dff_A_20PUEmxL3_0),.din(w_dff_A_kP9unsOF2_0),.clk(gclk));
	jdff dff_A_20PUEmxL3_0(.dout(w_dff_A_ejkMAAZs3_0),.din(w_dff_A_20PUEmxL3_0),.clk(gclk));
	jdff dff_A_ejkMAAZs3_0(.dout(w_dff_A_dCApbI2O4_0),.din(w_dff_A_ejkMAAZs3_0),.clk(gclk));
	jdff dff_A_dCApbI2O4_0(.dout(w_dff_A_aU1wrsgp7_0),.din(w_dff_A_dCApbI2O4_0),.clk(gclk));
	jdff dff_A_aU1wrsgp7_0(.dout(w_dff_A_jQsRCO0U5_0),.din(w_dff_A_aU1wrsgp7_0),.clk(gclk));
	jdff dff_A_jQsRCO0U5_0(.dout(w_dff_A_nXIB78Kc9_0),.din(w_dff_A_jQsRCO0U5_0),.clk(gclk));
	jdff dff_A_nXIB78Kc9_0(.dout(w_dff_A_kYEm73el2_0),.din(w_dff_A_nXIB78Kc9_0),.clk(gclk));
	jdff dff_A_kYEm73el2_0(.dout(w_dff_A_1PRRtXaw3_0),.din(w_dff_A_kYEm73el2_0),.clk(gclk));
	jdff dff_A_1PRRtXaw3_0(.dout(w_dff_A_HobxA5Cj0_0),.din(w_dff_A_1PRRtXaw3_0),.clk(gclk));
	jdff dff_A_HobxA5Cj0_0(.dout(w_dff_A_B0gsQ4BK5_0),.din(w_dff_A_HobxA5Cj0_0),.clk(gclk));
	jdff dff_A_B0gsQ4BK5_0(.dout(w_dff_A_GiycBwh69_0),.din(w_dff_A_B0gsQ4BK5_0),.clk(gclk));
	jdff dff_A_GiycBwh69_0(.dout(w_dff_A_qkA4Mohq0_0),.din(w_dff_A_GiycBwh69_0),.clk(gclk));
	jdff dff_A_qkA4Mohq0_0(.dout(G851),.din(w_dff_A_qkA4Mohq0_0),.clk(gclk));
	jdff dff_A_A73KRriC2_2(.dout(w_dff_A_QHRYgLdv8_0),.din(w_dff_A_A73KRriC2_2),.clk(gclk));
	jdff dff_A_QHRYgLdv8_0(.dout(w_dff_A_4LsF9tOB4_0),.din(w_dff_A_QHRYgLdv8_0),.clk(gclk));
	jdff dff_A_4LsF9tOB4_0(.dout(w_dff_A_hCGA9hfk1_0),.din(w_dff_A_4LsF9tOB4_0),.clk(gclk));
	jdff dff_A_hCGA9hfk1_0(.dout(w_dff_A_5FvsBG0u8_0),.din(w_dff_A_hCGA9hfk1_0),.clk(gclk));
	jdff dff_A_5FvsBG0u8_0(.dout(w_dff_A_dKeRzE1w3_0),.din(w_dff_A_5FvsBG0u8_0),.clk(gclk));
	jdff dff_A_dKeRzE1w3_0(.dout(w_dff_A_gHQSSUmJ3_0),.din(w_dff_A_dKeRzE1w3_0),.clk(gclk));
	jdff dff_A_gHQSSUmJ3_0(.dout(w_dff_A_t3MjPj938_0),.din(w_dff_A_gHQSSUmJ3_0),.clk(gclk));
	jdff dff_A_t3MjPj938_0(.dout(w_dff_A_tZ0GWu3a2_0),.din(w_dff_A_t3MjPj938_0),.clk(gclk));
	jdff dff_A_tZ0GWu3a2_0(.dout(w_dff_A_gLu1sFFu8_0),.din(w_dff_A_tZ0GWu3a2_0),.clk(gclk));
	jdff dff_A_gLu1sFFu8_0(.dout(w_dff_A_qqsvjRxu1_0),.din(w_dff_A_gLu1sFFu8_0),.clk(gclk));
	jdff dff_A_qqsvjRxu1_0(.dout(w_dff_A_tC2Pwm532_0),.din(w_dff_A_qqsvjRxu1_0),.clk(gclk));
	jdff dff_A_tC2Pwm532_0(.dout(w_dff_A_2uffUFaM1_0),.din(w_dff_A_tC2Pwm532_0),.clk(gclk));
	jdff dff_A_2uffUFaM1_0(.dout(w_dff_A_O6e1pLXQ9_0),.din(w_dff_A_2uffUFaM1_0),.clk(gclk));
	jdff dff_A_O6e1pLXQ9_0(.dout(w_dff_A_7cT1evW32_0),.din(w_dff_A_O6e1pLXQ9_0),.clk(gclk));
	jdff dff_A_7cT1evW32_0(.dout(w_dff_A_z1RjZZO91_0),.din(w_dff_A_7cT1evW32_0),.clk(gclk));
	jdff dff_A_z1RjZZO91_0(.dout(w_dff_A_YijuYlJI4_0),.din(w_dff_A_z1RjZZO91_0),.clk(gclk));
	jdff dff_A_YijuYlJI4_0(.dout(w_dff_A_8FDWZXzS1_0),.din(w_dff_A_YijuYlJI4_0),.clk(gclk));
	jdff dff_A_8FDWZXzS1_0(.dout(w_dff_A_Nuw0kKu89_0),.din(w_dff_A_8FDWZXzS1_0),.clk(gclk));
	jdff dff_A_Nuw0kKu89_0(.dout(w_dff_A_6TvhlGT81_0),.din(w_dff_A_Nuw0kKu89_0),.clk(gclk));
	jdff dff_A_6TvhlGT81_0(.dout(w_dff_A_B4UaiNhs6_0),.din(w_dff_A_6TvhlGT81_0),.clk(gclk));
	jdff dff_A_B4UaiNhs6_0(.dout(w_dff_A_UHQVVD6z6_0),.din(w_dff_A_B4UaiNhs6_0),.clk(gclk));
	jdff dff_A_UHQVVD6z6_0(.dout(w_dff_A_Ok9DwsHL7_0),.din(w_dff_A_UHQVVD6z6_0),.clk(gclk));
	jdff dff_A_Ok9DwsHL7_0(.dout(w_dff_A_b9BxmFUo9_0),.din(w_dff_A_Ok9DwsHL7_0),.clk(gclk));
	jdff dff_A_b9BxmFUo9_0(.dout(w_dff_A_EItsgsMe4_0),.din(w_dff_A_b9BxmFUo9_0),.clk(gclk));
	jdff dff_A_EItsgsMe4_0(.dout(G634),.din(w_dff_A_EItsgsMe4_0),.clk(gclk));
	jdff dff_A_qRvqPe0K0_2(.dout(w_dff_A_D7KvJIcy7_0),.din(w_dff_A_qRvqPe0K0_2),.clk(gclk));
	jdff dff_A_D7KvJIcy7_0(.dout(w_dff_A_DaslA0fS3_0),.din(w_dff_A_D7KvJIcy7_0),.clk(gclk));
	jdff dff_A_DaslA0fS3_0(.dout(w_dff_A_3QGzizf21_0),.din(w_dff_A_DaslA0fS3_0),.clk(gclk));
	jdff dff_A_3QGzizf21_0(.dout(w_dff_A_tsk0zT4j5_0),.din(w_dff_A_3QGzizf21_0),.clk(gclk));
	jdff dff_A_tsk0zT4j5_0(.dout(w_dff_A_gduYHa7o0_0),.din(w_dff_A_tsk0zT4j5_0),.clk(gclk));
	jdff dff_A_gduYHa7o0_0(.dout(w_dff_A_DvSzl4zs3_0),.din(w_dff_A_gduYHa7o0_0),.clk(gclk));
	jdff dff_A_DvSzl4zs3_0(.dout(w_dff_A_v50RVdLI0_0),.din(w_dff_A_DvSzl4zs3_0),.clk(gclk));
	jdff dff_A_v50RVdLI0_0(.dout(w_dff_A_orj4xZUA5_0),.din(w_dff_A_v50RVdLI0_0),.clk(gclk));
	jdff dff_A_orj4xZUA5_0(.dout(w_dff_A_rh5tpSUG7_0),.din(w_dff_A_orj4xZUA5_0),.clk(gclk));
	jdff dff_A_rh5tpSUG7_0(.dout(w_dff_A_I0CqYIGO7_0),.din(w_dff_A_rh5tpSUG7_0),.clk(gclk));
	jdff dff_A_I0CqYIGO7_0(.dout(w_dff_A_4wdrDtqJ4_0),.din(w_dff_A_I0CqYIGO7_0),.clk(gclk));
	jdff dff_A_4wdrDtqJ4_0(.dout(w_dff_A_Mxse4G6a9_0),.din(w_dff_A_4wdrDtqJ4_0),.clk(gclk));
	jdff dff_A_Mxse4G6a9_0(.dout(w_dff_A_Cx8DkS5H3_0),.din(w_dff_A_Mxse4G6a9_0),.clk(gclk));
	jdff dff_A_Cx8DkS5H3_0(.dout(w_dff_A_eBnPuevc3_0),.din(w_dff_A_Cx8DkS5H3_0),.clk(gclk));
	jdff dff_A_eBnPuevc3_0(.dout(w_dff_A_uROkI5549_0),.din(w_dff_A_eBnPuevc3_0),.clk(gclk));
	jdff dff_A_uROkI5549_0(.dout(w_dff_A_bdmvwmqG5_0),.din(w_dff_A_uROkI5549_0),.clk(gclk));
	jdff dff_A_bdmvwmqG5_0(.dout(w_dff_A_YfhpMKSF4_0),.din(w_dff_A_bdmvwmqG5_0),.clk(gclk));
	jdff dff_A_YfhpMKSF4_0(.dout(w_dff_A_66Mgpz6z8_0),.din(w_dff_A_YfhpMKSF4_0),.clk(gclk));
	jdff dff_A_66Mgpz6z8_0(.dout(w_dff_A_CfEES1kc0_0),.din(w_dff_A_66Mgpz6z8_0),.clk(gclk));
	jdff dff_A_CfEES1kc0_0(.dout(w_dff_A_4ab1mCmT7_0),.din(w_dff_A_CfEES1kc0_0),.clk(gclk));
	jdff dff_A_4ab1mCmT7_0(.dout(w_dff_A_jGYyayqq1_0),.din(w_dff_A_4ab1mCmT7_0),.clk(gclk));
	jdff dff_A_jGYyayqq1_0(.dout(w_dff_A_qjFC11q62_0),.din(w_dff_A_jGYyayqq1_0),.clk(gclk));
	jdff dff_A_qjFC11q62_0(.dout(w_dff_A_sdlJCghR9_0),.din(w_dff_A_qjFC11q62_0),.clk(gclk));
	jdff dff_A_sdlJCghR9_0(.dout(G815),.din(w_dff_A_sdlJCghR9_0),.clk(gclk));
	jdff dff_A_hpXzg0xe9_2(.dout(w_dff_A_TWtoqQQE9_0),.din(w_dff_A_hpXzg0xe9_2),.clk(gclk));
	jdff dff_A_TWtoqQQE9_0(.dout(w_dff_A_ngK5VdIU5_0),.din(w_dff_A_TWtoqQQE9_0),.clk(gclk));
	jdff dff_A_ngK5VdIU5_0(.dout(w_dff_A_G65L7igr6_0),.din(w_dff_A_ngK5VdIU5_0),.clk(gclk));
	jdff dff_A_G65L7igr6_0(.dout(w_dff_A_nlB2Z9oG0_0),.din(w_dff_A_G65L7igr6_0),.clk(gclk));
	jdff dff_A_nlB2Z9oG0_0(.dout(w_dff_A_SeMPnqRd8_0),.din(w_dff_A_nlB2Z9oG0_0),.clk(gclk));
	jdff dff_A_SeMPnqRd8_0(.dout(w_dff_A_jBQt9ucz5_0),.din(w_dff_A_SeMPnqRd8_0),.clk(gclk));
	jdff dff_A_jBQt9ucz5_0(.dout(w_dff_A_ubcbUSwX4_0),.din(w_dff_A_jBQt9ucz5_0),.clk(gclk));
	jdff dff_A_ubcbUSwX4_0(.dout(w_dff_A_zlTo5ASg6_0),.din(w_dff_A_ubcbUSwX4_0),.clk(gclk));
	jdff dff_A_zlTo5ASg6_0(.dout(w_dff_A_ppqfRdBU7_0),.din(w_dff_A_zlTo5ASg6_0),.clk(gclk));
	jdff dff_A_ppqfRdBU7_0(.dout(w_dff_A_WB1f71cN7_0),.din(w_dff_A_ppqfRdBU7_0),.clk(gclk));
	jdff dff_A_WB1f71cN7_0(.dout(w_dff_A_leGahstU2_0),.din(w_dff_A_WB1f71cN7_0),.clk(gclk));
	jdff dff_A_leGahstU2_0(.dout(w_dff_A_UOCkYlVC0_0),.din(w_dff_A_leGahstU2_0),.clk(gclk));
	jdff dff_A_UOCkYlVC0_0(.dout(w_dff_A_TXicrlqP7_0),.din(w_dff_A_UOCkYlVC0_0),.clk(gclk));
	jdff dff_A_TXicrlqP7_0(.dout(w_dff_A_7AJTUEqQ3_0),.din(w_dff_A_TXicrlqP7_0),.clk(gclk));
	jdff dff_A_7AJTUEqQ3_0(.dout(w_dff_A_LMJS409g4_0),.din(w_dff_A_7AJTUEqQ3_0),.clk(gclk));
	jdff dff_A_LMJS409g4_0(.dout(w_dff_A_QR8GrEX93_0),.din(w_dff_A_LMJS409g4_0),.clk(gclk));
	jdff dff_A_QR8GrEX93_0(.dout(w_dff_A_sDua6Qoj6_0),.din(w_dff_A_QR8GrEX93_0),.clk(gclk));
	jdff dff_A_sDua6Qoj6_0(.dout(w_dff_A_G2eDTmua9_0),.din(w_dff_A_sDua6Qoj6_0),.clk(gclk));
	jdff dff_A_G2eDTmua9_0(.dout(w_dff_A_w8qi5ew93_0),.din(w_dff_A_G2eDTmua9_0),.clk(gclk));
	jdff dff_A_w8qi5ew93_0(.dout(w_dff_A_Eeoy4mWu5_0),.din(w_dff_A_w8qi5ew93_0),.clk(gclk));
	jdff dff_A_Eeoy4mWu5_0(.dout(w_dff_A_l9LU6LYt1_0),.din(w_dff_A_Eeoy4mWu5_0),.clk(gclk));
	jdff dff_A_l9LU6LYt1_0(.dout(w_dff_A_2gjwdEwy1_0),.din(w_dff_A_l9LU6LYt1_0),.clk(gclk));
	jdff dff_A_2gjwdEwy1_0(.dout(w_dff_A_V33cnRmT1_0),.din(w_dff_A_2gjwdEwy1_0),.clk(gclk));
	jdff dff_A_V33cnRmT1_0(.dout(G845),.din(w_dff_A_V33cnRmT1_0),.clk(gclk));
	jdff dff_A_ViUahs343_1(.dout(w_dff_A_iooO0VpB8_0),.din(w_dff_A_ViUahs343_1),.clk(gclk));
	jdff dff_A_iooO0VpB8_0(.dout(w_dff_A_GqFfNTRm6_0),.din(w_dff_A_iooO0VpB8_0),.clk(gclk));
	jdff dff_A_GqFfNTRm6_0(.dout(w_dff_A_DIAmK1Gj2_0),.din(w_dff_A_GqFfNTRm6_0),.clk(gclk));
	jdff dff_A_DIAmK1Gj2_0(.dout(w_dff_A_l58GALg67_0),.din(w_dff_A_DIAmK1Gj2_0),.clk(gclk));
	jdff dff_A_l58GALg67_0(.dout(w_dff_A_VwiD7fc74_0),.din(w_dff_A_l58GALg67_0),.clk(gclk));
	jdff dff_A_VwiD7fc74_0(.dout(w_dff_A_jQ7aw5Ve5_0),.din(w_dff_A_VwiD7fc74_0),.clk(gclk));
	jdff dff_A_jQ7aw5Ve5_0(.dout(w_dff_A_ZXp10W1O4_0),.din(w_dff_A_jQ7aw5Ve5_0),.clk(gclk));
	jdff dff_A_ZXp10W1O4_0(.dout(w_dff_A_TLzDrl8S1_0),.din(w_dff_A_ZXp10W1O4_0),.clk(gclk));
	jdff dff_A_TLzDrl8S1_0(.dout(w_dff_A_x4LqO9DE2_0),.din(w_dff_A_TLzDrl8S1_0),.clk(gclk));
	jdff dff_A_x4LqO9DE2_0(.dout(w_dff_A_Q5EXAufB1_0),.din(w_dff_A_x4LqO9DE2_0),.clk(gclk));
	jdff dff_A_Q5EXAufB1_0(.dout(w_dff_A_FubuaEPB5_0),.din(w_dff_A_Q5EXAufB1_0),.clk(gclk));
	jdff dff_A_FubuaEPB5_0(.dout(w_dff_A_mq4gRUuZ2_0),.din(w_dff_A_FubuaEPB5_0),.clk(gclk));
	jdff dff_A_mq4gRUuZ2_0(.dout(w_dff_A_DalA584P0_0),.din(w_dff_A_mq4gRUuZ2_0),.clk(gclk));
	jdff dff_A_DalA584P0_0(.dout(w_dff_A_SvTN4RbA8_0),.din(w_dff_A_DalA584P0_0),.clk(gclk));
	jdff dff_A_SvTN4RbA8_0(.dout(w_dff_A_v4muk1iP9_0),.din(w_dff_A_SvTN4RbA8_0),.clk(gclk));
	jdff dff_A_v4muk1iP9_0(.dout(w_dff_A_c7zLx6yB7_0),.din(w_dff_A_v4muk1iP9_0),.clk(gclk));
	jdff dff_A_c7zLx6yB7_0(.dout(w_dff_A_tprq0Hsr1_0),.din(w_dff_A_c7zLx6yB7_0),.clk(gclk));
	jdff dff_A_tprq0Hsr1_0(.dout(w_dff_A_aNegmzWn2_0),.din(w_dff_A_tprq0Hsr1_0),.clk(gclk));
	jdff dff_A_aNegmzWn2_0(.dout(w_dff_A_M0CC1hHB9_0),.din(w_dff_A_aNegmzWn2_0),.clk(gclk));
	jdff dff_A_M0CC1hHB9_0(.dout(w_dff_A_j82XPKqP0_0),.din(w_dff_A_M0CC1hHB9_0),.clk(gclk));
	jdff dff_A_j82XPKqP0_0(.dout(w_dff_A_jXyNHNnt2_0),.din(w_dff_A_j82XPKqP0_0),.clk(gclk));
	jdff dff_A_jXyNHNnt2_0(.dout(w_dff_A_6ayynWL57_0),.din(w_dff_A_jXyNHNnt2_0),.clk(gclk));
	jdff dff_A_6ayynWL57_0(.dout(w_dff_A_QBe88BDj7_0),.din(w_dff_A_6ayynWL57_0),.clk(gclk));
	jdff dff_A_QBe88BDj7_0(.dout(G847),.din(w_dff_A_QBe88BDj7_0),.clk(gclk));
	jdff dff_A_sj71NC4V1_1(.dout(w_dff_A_u8QhvmQL6_0),.din(w_dff_A_sj71NC4V1_1),.clk(gclk));
	jdff dff_A_u8QhvmQL6_0(.dout(w_dff_A_18pQDlkp1_0),.din(w_dff_A_u8QhvmQL6_0),.clk(gclk));
	jdff dff_A_18pQDlkp1_0(.dout(w_dff_A_zNK6xxn77_0),.din(w_dff_A_18pQDlkp1_0),.clk(gclk));
	jdff dff_A_zNK6xxn77_0(.dout(w_dff_A_YN3cziQw5_0),.din(w_dff_A_zNK6xxn77_0),.clk(gclk));
	jdff dff_A_YN3cziQw5_0(.dout(w_dff_A_Bpgxn6Dk3_0),.din(w_dff_A_YN3cziQw5_0),.clk(gclk));
	jdff dff_A_Bpgxn6Dk3_0(.dout(w_dff_A_RY7KrXhu6_0),.din(w_dff_A_Bpgxn6Dk3_0),.clk(gclk));
	jdff dff_A_RY7KrXhu6_0(.dout(w_dff_A_XBvdImye8_0),.din(w_dff_A_RY7KrXhu6_0),.clk(gclk));
	jdff dff_A_XBvdImye8_0(.dout(w_dff_A_Zcu60hBh6_0),.din(w_dff_A_XBvdImye8_0),.clk(gclk));
	jdff dff_A_Zcu60hBh6_0(.dout(w_dff_A_jumul6F60_0),.din(w_dff_A_Zcu60hBh6_0),.clk(gclk));
	jdff dff_A_jumul6F60_0(.dout(w_dff_A_KpG0jdCq9_0),.din(w_dff_A_jumul6F60_0),.clk(gclk));
	jdff dff_A_KpG0jdCq9_0(.dout(w_dff_A_rx8Hxp1C9_0),.din(w_dff_A_KpG0jdCq9_0),.clk(gclk));
	jdff dff_A_rx8Hxp1C9_0(.dout(w_dff_A_lD9JQRWf1_0),.din(w_dff_A_rx8Hxp1C9_0),.clk(gclk));
	jdff dff_A_lD9JQRWf1_0(.dout(w_dff_A_yvK7Q4Cv6_0),.din(w_dff_A_lD9JQRWf1_0),.clk(gclk));
	jdff dff_A_yvK7Q4Cv6_0(.dout(w_dff_A_eICuoqTu9_0),.din(w_dff_A_yvK7Q4Cv6_0),.clk(gclk));
	jdff dff_A_eICuoqTu9_0(.dout(w_dff_A_kWXSdlQl2_0),.din(w_dff_A_eICuoqTu9_0),.clk(gclk));
	jdff dff_A_kWXSdlQl2_0(.dout(w_dff_A_Yr1dCKCl0_0),.din(w_dff_A_kWXSdlQl2_0),.clk(gclk));
	jdff dff_A_Yr1dCKCl0_0(.dout(w_dff_A_PugyfsXq2_0),.din(w_dff_A_Yr1dCKCl0_0),.clk(gclk));
	jdff dff_A_PugyfsXq2_0(.dout(w_dff_A_KFSqPgz87_0),.din(w_dff_A_PugyfsXq2_0),.clk(gclk));
	jdff dff_A_KFSqPgz87_0(.dout(w_dff_A_palNUYEn7_0),.din(w_dff_A_KFSqPgz87_0),.clk(gclk));
	jdff dff_A_palNUYEn7_0(.dout(w_dff_A_B5b7hgEZ1_0),.din(w_dff_A_palNUYEn7_0),.clk(gclk));
	jdff dff_A_B5b7hgEZ1_0(.dout(w_dff_A_FFtnOU926_0),.din(w_dff_A_B5b7hgEZ1_0),.clk(gclk));
	jdff dff_A_FFtnOU926_0(.dout(w_dff_A_NPFPFwoX6_0),.din(w_dff_A_FFtnOU926_0),.clk(gclk));
	jdff dff_A_NPFPFwoX6_0(.dout(w_dff_A_hlJLiJZ32_0),.din(w_dff_A_NPFPFwoX6_0),.clk(gclk));
	jdff dff_A_hlJLiJZ32_0(.dout(w_dff_A_T4XgKpFB1_0),.din(w_dff_A_hlJLiJZ32_0),.clk(gclk));
	jdff dff_A_T4XgKpFB1_0(.dout(w_dff_A_lBK96Nf12_0),.din(w_dff_A_T4XgKpFB1_0),.clk(gclk));
	jdff dff_A_lBK96Nf12_0(.dout(G926),.din(w_dff_A_lBK96Nf12_0),.clk(gclk));
	jdff dff_A_HaCj6xuk2_1(.dout(w_dff_A_Do4ByAWj8_0),.din(w_dff_A_HaCj6xuk2_1),.clk(gclk));
	jdff dff_A_Do4ByAWj8_0(.dout(w_dff_A_pEXzaAKn9_0),.din(w_dff_A_Do4ByAWj8_0),.clk(gclk));
	jdff dff_A_pEXzaAKn9_0(.dout(w_dff_A_LneWEKAY7_0),.din(w_dff_A_pEXzaAKn9_0),.clk(gclk));
	jdff dff_A_LneWEKAY7_0(.dout(w_dff_A_eDcx02rZ3_0),.din(w_dff_A_LneWEKAY7_0),.clk(gclk));
	jdff dff_A_eDcx02rZ3_0(.dout(w_dff_A_Bxoy26mD0_0),.din(w_dff_A_eDcx02rZ3_0),.clk(gclk));
	jdff dff_A_Bxoy26mD0_0(.dout(w_dff_A_s6as2Cm73_0),.din(w_dff_A_Bxoy26mD0_0),.clk(gclk));
	jdff dff_A_s6as2Cm73_0(.dout(w_dff_A_Xo2Jylnz4_0),.din(w_dff_A_s6as2Cm73_0),.clk(gclk));
	jdff dff_A_Xo2Jylnz4_0(.dout(w_dff_A_MoZ7CPFV7_0),.din(w_dff_A_Xo2Jylnz4_0),.clk(gclk));
	jdff dff_A_MoZ7CPFV7_0(.dout(w_dff_A_3m05lXNH2_0),.din(w_dff_A_MoZ7CPFV7_0),.clk(gclk));
	jdff dff_A_3m05lXNH2_0(.dout(w_dff_A_epk0eIWO1_0),.din(w_dff_A_3m05lXNH2_0),.clk(gclk));
	jdff dff_A_epk0eIWO1_0(.dout(w_dff_A_GLoXhBjM3_0),.din(w_dff_A_epk0eIWO1_0),.clk(gclk));
	jdff dff_A_GLoXhBjM3_0(.dout(w_dff_A_SwNnoWVC5_0),.din(w_dff_A_GLoXhBjM3_0),.clk(gclk));
	jdff dff_A_SwNnoWVC5_0(.dout(w_dff_A_GDDK4qB99_0),.din(w_dff_A_SwNnoWVC5_0),.clk(gclk));
	jdff dff_A_GDDK4qB99_0(.dout(w_dff_A_UlkBzqS80_0),.din(w_dff_A_GDDK4qB99_0),.clk(gclk));
	jdff dff_A_UlkBzqS80_0(.dout(w_dff_A_RjcBw8jC4_0),.din(w_dff_A_UlkBzqS80_0),.clk(gclk));
	jdff dff_A_RjcBw8jC4_0(.dout(w_dff_A_NDF14ZRB0_0),.din(w_dff_A_RjcBw8jC4_0),.clk(gclk));
	jdff dff_A_NDF14ZRB0_0(.dout(w_dff_A_4NIJGMTk7_0),.din(w_dff_A_NDF14ZRB0_0),.clk(gclk));
	jdff dff_A_4NIJGMTk7_0(.dout(w_dff_A_p0ja5tRh9_0),.din(w_dff_A_4NIJGMTk7_0),.clk(gclk));
	jdff dff_A_p0ja5tRh9_0(.dout(w_dff_A_XQSXx6Ub9_0),.din(w_dff_A_p0ja5tRh9_0),.clk(gclk));
	jdff dff_A_XQSXx6Ub9_0(.dout(w_dff_A_RKpPEadB9_0),.din(w_dff_A_XQSXx6Ub9_0),.clk(gclk));
	jdff dff_A_RKpPEadB9_0(.dout(w_dff_A_7SHw5ATD8_0),.din(w_dff_A_RKpPEadB9_0),.clk(gclk));
	jdff dff_A_7SHw5ATD8_0(.dout(w_dff_A_6Khi0dL85_0),.din(w_dff_A_7SHw5ATD8_0),.clk(gclk));
	jdff dff_A_6Khi0dL85_0(.dout(w_dff_A_s42y9RX06_0),.din(w_dff_A_6Khi0dL85_0),.clk(gclk));
	jdff dff_A_s42y9RX06_0(.dout(w_dff_A_nuSZYBV88_0),.din(w_dff_A_s42y9RX06_0),.clk(gclk));
	jdff dff_A_nuSZYBV88_0(.dout(w_dff_A_Y3MnGbpo4_0),.din(w_dff_A_nuSZYBV88_0),.clk(gclk));
	jdff dff_A_Y3MnGbpo4_0(.dout(G923),.din(w_dff_A_Y3MnGbpo4_0),.clk(gclk));
	jdff dff_A_n3PHt2IB0_1(.dout(w_dff_A_bslqJ3iy3_0),.din(w_dff_A_n3PHt2IB0_1),.clk(gclk));
	jdff dff_A_bslqJ3iy3_0(.dout(w_dff_A_lwbjCbjp8_0),.din(w_dff_A_bslqJ3iy3_0),.clk(gclk));
	jdff dff_A_lwbjCbjp8_0(.dout(w_dff_A_5A6w6emc4_0),.din(w_dff_A_lwbjCbjp8_0),.clk(gclk));
	jdff dff_A_5A6w6emc4_0(.dout(w_dff_A_ssXT6xpk9_0),.din(w_dff_A_5A6w6emc4_0),.clk(gclk));
	jdff dff_A_ssXT6xpk9_0(.dout(w_dff_A_dCNjHbkt8_0),.din(w_dff_A_ssXT6xpk9_0),.clk(gclk));
	jdff dff_A_dCNjHbkt8_0(.dout(w_dff_A_5pspdUro8_0),.din(w_dff_A_dCNjHbkt8_0),.clk(gclk));
	jdff dff_A_5pspdUro8_0(.dout(w_dff_A_qdlZwsXj9_0),.din(w_dff_A_5pspdUro8_0),.clk(gclk));
	jdff dff_A_qdlZwsXj9_0(.dout(w_dff_A_CI3UD1XA2_0),.din(w_dff_A_qdlZwsXj9_0),.clk(gclk));
	jdff dff_A_CI3UD1XA2_0(.dout(w_dff_A_BIuxpNiH4_0),.din(w_dff_A_CI3UD1XA2_0),.clk(gclk));
	jdff dff_A_BIuxpNiH4_0(.dout(w_dff_A_ypZiefm88_0),.din(w_dff_A_BIuxpNiH4_0),.clk(gclk));
	jdff dff_A_ypZiefm88_0(.dout(w_dff_A_nD5N2UIu4_0),.din(w_dff_A_ypZiefm88_0),.clk(gclk));
	jdff dff_A_nD5N2UIu4_0(.dout(w_dff_A_YcznuUwt2_0),.din(w_dff_A_nD5N2UIu4_0),.clk(gclk));
	jdff dff_A_YcznuUwt2_0(.dout(w_dff_A_CVAGcaXa1_0),.din(w_dff_A_YcznuUwt2_0),.clk(gclk));
	jdff dff_A_CVAGcaXa1_0(.dout(w_dff_A_n09Nnwt84_0),.din(w_dff_A_CVAGcaXa1_0),.clk(gclk));
	jdff dff_A_n09Nnwt84_0(.dout(w_dff_A_pfBjQgUp0_0),.din(w_dff_A_n09Nnwt84_0),.clk(gclk));
	jdff dff_A_pfBjQgUp0_0(.dout(w_dff_A_6DapTIE14_0),.din(w_dff_A_pfBjQgUp0_0),.clk(gclk));
	jdff dff_A_6DapTIE14_0(.dout(w_dff_A_oZW4B5QZ4_0),.din(w_dff_A_6DapTIE14_0),.clk(gclk));
	jdff dff_A_oZW4B5QZ4_0(.dout(w_dff_A_bUsUSjIn0_0),.din(w_dff_A_oZW4B5QZ4_0),.clk(gclk));
	jdff dff_A_bUsUSjIn0_0(.dout(w_dff_A_EA4aZZpD4_0),.din(w_dff_A_bUsUSjIn0_0),.clk(gclk));
	jdff dff_A_EA4aZZpD4_0(.dout(w_dff_A_xj2oHy7A8_0),.din(w_dff_A_EA4aZZpD4_0),.clk(gclk));
	jdff dff_A_xj2oHy7A8_0(.dout(w_dff_A_urw1ziEL2_0),.din(w_dff_A_xj2oHy7A8_0),.clk(gclk));
	jdff dff_A_urw1ziEL2_0(.dout(w_dff_A_nKjh5oZt2_0),.din(w_dff_A_urw1ziEL2_0),.clk(gclk));
	jdff dff_A_nKjh5oZt2_0(.dout(w_dff_A_FILaSPKv5_0),.din(w_dff_A_nKjh5oZt2_0),.clk(gclk));
	jdff dff_A_FILaSPKv5_0(.dout(w_dff_A_KI8CJEtM4_0),.din(w_dff_A_FILaSPKv5_0),.clk(gclk));
	jdff dff_A_KI8CJEtM4_0(.dout(w_dff_A_9FnmD0E05_0),.din(w_dff_A_KI8CJEtM4_0),.clk(gclk));
	jdff dff_A_9FnmD0E05_0(.dout(G921),.din(w_dff_A_9FnmD0E05_0),.clk(gclk));
	jdff dff_A_Gx44yVSc7_1(.dout(w_dff_A_kfethRvJ8_0),.din(w_dff_A_Gx44yVSc7_1),.clk(gclk));
	jdff dff_A_kfethRvJ8_0(.dout(w_dff_A_wNrtEa7B8_0),.din(w_dff_A_kfethRvJ8_0),.clk(gclk));
	jdff dff_A_wNrtEa7B8_0(.dout(w_dff_A_aXEvXYaV5_0),.din(w_dff_A_wNrtEa7B8_0),.clk(gclk));
	jdff dff_A_aXEvXYaV5_0(.dout(w_dff_A_61Yjs9Fi8_0),.din(w_dff_A_aXEvXYaV5_0),.clk(gclk));
	jdff dff_A_61Yjs9Fi8_0(.dout(w_dff_A_JlmwLIQT2_0),.din(w_dff_A_61Yjs9Fi8_0),.clk(gclk));
	jdff dff_A_JlmwLIQT2_0(.dout(w_dff_A_fong6TIP8_0),.din(w_dff_A_JlmwLIQT2_0),.clk(gclk));
	jdff dff_A_fong6TIP8_0(.dout(w_dff_A_4MXegcaY7_0),.din(w_dff_A_fong6TIP8_0),.clk(gclk));
	jdff dff_A_4MXegcaY7_0(.dout(w_dff_A_Q55zYvG36_0),.din(w_dff_A_4MXegcaY7_0),.clk(gclk));
	jdff dff_A_Q55zYvG36_0(.dout(w_dff_A_GXKKp3W53_0),.din(w_dff_A_Q55zYvG36_0),.clk(gclk));
	jdff dff_A_GXKKp3W53_0(.dout(w_dff_A_tZpmmXVc1_0),.din(w_dff_A_GXKKp3W53_0),.clk(gclk));
	jdff dff_A_tZpmmXVc1_0(.dout(w_dff_A_75xU5udf0_0),.din(w_dff_A_tZpmmXVc1_0),.clk(gclk));
	jdff dff_A_75xU5udf0_0(.dout(w_dff_A_fMTdgve52_0),.din(w_dff_A_75xU5udf0_0),.clk(gclk));
	jdff dff_A_fMTdgve52_0(.dout(w_dff_A_jwNI3Ic87_0),.din(w_dff_A_fMTdgve52_0),.clk(gclk));
	jdff dff_A_jwNI3Ic87_0(.dout(w_dff_A_8r6bQmHS7_0),.din(w_dff_A_jwNI3Ic87_0),.clk(gclk));
	jdff dff_A_8r6bQmHS7_0(.dout(w_dff_A_IZb8XFCE9_0),.din(w_dff_A_8r6bQmHS7_0),.clk(gclk));
	jdff dff_A_IZb8XFCE9_0(.dout(w_dff_A_Nfs7hVum7_0),.din(w_dff_A_IZb8XFCE9_0),.clk(gclk));
	jdff dff_A_Nfs7hVum7_0(.dout(w_dff_A_xvxoChTQ2_0),.din(w_dff_A_Nfs7hVum7_0),.clk(gclk));
	jdff dff_A_xvxoChTQ2_0(.dout(w_dff_A_ySY0MIM84_0),.din(w_dff_A_xvxoChTQ2_0),.clk(gclk));
	jdff dff_A_ySY0MIM84_0(.dout(w_dff_A_BmZI0J9D9_0),.din(w_dff_A_ySY0MIM84_0),.clk(gclk));
	jdff dff_A_BmZI0J9D9_0(.dout(w_dff_A_cG0Ai9um9_0),.din(w_dff_A_BmZI0J9D9_0),.clk(gclk));
	jdff dff_A_cG0Ai9um9_0(.dout(w_dff_A_TZDqMABz9_0),.din(w_dff_A_cG0Ai9um9_0),.clk(gclk));
	jdff dff_A_TZDqMABz9_0(.dout(w_dff_A_qdRxkQvC4_0),.din(w_dff_A_TZDqMABz9_0),.clk(gclk));
	jdff dff_A_qdRxkQvC4_0(.dout(w_dff_A_VCRbQayE6_0),.din(w_dff_A_qdRxkQvC4_0),.clk(gclk));
	jdff dff_A_VCRbQayE6_0(.dout(w_dff_A_MIiA93gJ4_0),.din(w_dff_A_VCRbQayE6_0),.clk(gclk));
	jdff dff_A_MIiA93gJ4_0(.dout(w_dff_A_4HnryNRv4_0),.din(w_dff_A_MIiA93gJ4_0),.clk(gclk));
	jdff dff_A_4HnryNRv4_0(.dout(G892),.din(w_dff_A_4HnryNRv4_0),.clk(gclk));
	jdff dff_A_omMcWl0V5_1(.dout(w_dff_A_tRwaXqEU9_0),.din(w_dff_A_omMcWl0V5_1),.clk(gclk));
	jdff dff_A_tRwaXqEU9_0(.dout(w_dff_A_ACf52F0F0_0),.din(w_dff_A_tRwaXqEU9_0),.clk(gclk));
	jdff dff_A_ACf52F0F0_0(.dout(w_dff_A_W5kvFPZr5_0),.din(w_dff_A_ACf52F0F0_0),.clk(gclk));
	jdff dff_A_W5kvFPZr5_0(.dout(w_dff_A_uzBXmwV79_0),.din(w_dff_A_W5kvFPZr5_0),.clk(gclk));
	jdff dff_A_uzBXmwV79_0(.dout(w_dff_A_hMjOgwuS1_0),.din(w_dff_A_uzBXmwV79_0),.clk(gclk));
	jdff dff_A_hMjOgwuS1_0(.dout(w_dff_A_nh3uSt8b6_0),.din(w_dff_A_hMjOgwuS1_0),.clk(gclk));
	jdff dff_A_nh3uSt8b6_0(.dout(w_dff_A_759wugz15_0),.din(w_dff_A_nh3uSt8b6_0),.clk(gclk));
	jdff dff_A_759wugz15_0(.dout(w_dff_A_zyIDLgoI3_0),.din(w_dff_A_759wugz15_0),.clk(gclk));
	jdff dff_A_zyIDLgoI3_0(.dout(w_dff_A_MnNdpAUC3_0),.din(w_dff_A_zyIDLgoI3_0),.clk(gclk));
	jdff dff_A_MnNdpAUC3_0(.dout(w_dff_A_crKFmxLn0_0),.din(w_dff_A_MnNdpAUC3_0),.clk(gclk));
	jdff dff_A_crKFmxLn0_0(.dout(w_dff_A_lzMNu7TQ3_0),.din(w_dff_A_crKFmxLn0_0),.clk(gclk));
	jdff dff_A_lzMNu7TQ3_0(.dout(w_dff_A_y47jTir70_0),.din(w_dff_A_lzMNu7TQ3_0),.clk(gclk));
	jdff dff_A_y47jTir70_0(.dout(w_dff_A_2NXNj62p0_0),.din(w_dff_A_y47jTir70_0),.clk(gclk));
	jdff dff_A_2NXNj62p0_0(.dout(w_dff_A_TJn0iHql8_0),.din(w_dff_A_2NXNj62p0_0),.clk(gclk));
	jdff dff_A_TJn0iHql8_0(.dout(w_dff_A_nWBDILmJ2_0),.din(w_dff_A_TJn0iHql8_0),.clk(gclk));
	jdff dff_A_nWBDILmJ2_0(.dout(w_dff_A_tds29IkS8_0),.din(w_dff_A_nWBDILmJ2_0),.clk(gclk));
	jdff dff_A_tds29IkS8_0(.dout(w_dff_A_bXJ5YoBX1_0),.din(w_dff_A_tds29IkS8_0),.clk(gclk));
	jdff dff_A_bXJ5YoBX1_0(.dout(w_dff_A_LzUIwyaC7_0),.din(w_dff_A_bXJ5YoBX1_0),.clk(gclk));
	jdff dff_A_LzUIwyaC7_0(.dout(w_dff_A_gGxr83iC6_0),.din(w_dff_A_LzUIwyaC7_0),.clk(gclk));
	jdff dff_A_gGxr83iC6_0(.dout(w_dff_A_IlIOQTTt9_0),.din(w_dff_A_gGxr83iC6_0),.clk(gclk));
	jdff dff_A_IlIOQTTt9_0(.dout(w_dff_A_FfXLtBh03_0),.din(w_dff_A_IlIOQTTt9_0),.clk(gclk));
	jdff dff_A_FfXLtBh03_0(.dout(w_dff_A_QDHA37He2_0),.din(w_dff_A_FfXLtBh03_0),.clk(gclk));
	jdff dff_A_QDHA37He2_0(.dout(w_dff_A_TxLsiOcT8_0),.din(w_dff_A_QDHA37He2_0),.clk(gclk));
	jdff dff_A_TxLsiOcT8_0(.dout(w_dff_A_TVUS04Wy4_0),.din(w_dff_A_TxLsiOcT8_0),.clk(gclk));
	jdff dff_A_TVUS04Wy4_0(.dout(w_dff_A_bw4nEjLL6_0),.din(w_dff_A_TVUS04Wy4_0),.clk(gclk));
	jdff dff_A_bw4nEjLL6_0(.dout(G887),.din(w_dff_A_bw4nEjLL6_0),.clk(gclk));
	jdff dff_A_KkjYaiEQ9_1(.dout(w_dff_A_37rmaHFS4_0),.din(w_dff_A_KkjYaiEQ9_1),.clk(gclk));
	jdff dff_A_37rmaHFS4_0(.dout(w_dff_A_iAvk41Do5_0),.din(w_dff_A_37rmaHFS4_0),.clk(gclk));
	jdff dff_A_iAvk41Do5_0(.dout(w_dff_A_CGg2NHQu7_0),.din(w_dff_A_iAvk41Do5_0),.clk(gclk));
	jdff dff_A_CGg2NHQu7_0(.dout(w_dff_A_BUorYZW25_0),.din(w_dff_A_CGg2NHQu7_0),.clk(gclk));
	jdff dff_A_BUorYZW25_0(.dout(w_dff_A_l1iMm9iP7_0),.din(w_dff_A_BUorYZW25_0),.clk(gclk));
	jdff dff_A_l1iMm9iP7_0(.dout(w_dff_A_3eQzTXUd7_0),.din(w_dff_A_l1iMm9iP7_0),.clk(gclk));
	jdff dff_A_3eQzTXUd7_0(.dout(w_dff_A_Au4ouYjb2_0),.din(w_dff_A_3eQzTXUd7_0),.clk(gclk));
	jdff dff_A_Au4ouYjb2_0(.dout(w_dff_A_Hnnb46RA5_0),.din(w_dff_A_Au4ouYjb2_0),.clk(gclk));
	jdff dff_A_Hnnb46RA5_0(.dout(w_dff_A_u0FIKi8D7_0),.din(w_dff_A_Hnnb46RA5_0),.clk(gclk));
	jdff dff_A_u0FIKi8D7_0(.dout(w_dff_A_98jx0DKn8_0),.din(w_dff_A_u0FIKi8D7_0),.clk(gclk));
	jdff dff_A_98jx0DKn8_0(.dout(w_dff_A_GQsBvA5B7_0),.din(w_dff_A_98jx0DKn8_0),.clk(gclk));
	jdff dff_A_GQsBvA5B7_0(.dout(w_dff_A_Trn5Sxqr3_0),.din(w_dff_A_GQsBvA5B7_0),.clk(gclk));
	jdff dff_A_Trn5Sxqr3_0(.dout(w_dff_A_KAHbB80g2_0),.din(w_dff_A_Trn5Sxqr3_0),.clk(gclk));
	jdff dff_A_KAHbB80g2_0(.dout(w_dff_A_BVxY8GzL7_0),.din(w_dff_A_KAHbB80g2_0),.clk(gclk));
	jdff dff_A_BVxY8GzL7_0(.dout(w_dff_A_Srngh5hg1_0),.din(w_dff_A_BVxY8GzL7_0),.clk(gclk));
	jdff dff_A_Srngh5hg1_0(.dout(w_dff_A_gJnKQ1gH6_0),.din(w_dff_A_Srngh5hg1_0),.clk(gclk));
	jdff dff_A_gJnKQ1gH6_0(.dout(w_dff_A_13zGVZPW0_0),.din(w_dff_A_gJnKQ1gH6_0),.clk(gclk));
	jdff dff_A_13zGVZPW0_0(.dout(w_dff_A_PA6JAdQw6_0),.din(w_dff_A_13zGVZPW0_0),.clk(gclk));
	jdff dff_A_PA6JAdQw6_0(.dout(w_dff_A_lkMTwbdw2_0),.din(w_dff_A_PA6JAdQw6_0),.clk(gclk));
	jdff dff_A_lkMTwbdw2_0(.dout(w_dff_A_Uz3M34Jx7_0),.din(w_dff_A_lkMTwbdw2_0),.clk(gclk));
	jdff dff_A_Uz3M34Jx7_0(.dout(w_dff_A_6WIGjWsv7_0),.din(w_dff_A_Uz3M34Jx7_0),.clk(gclk));
	jdff dff_A_6WIGjWsv7_0(.dout(w_dff_A_kgYb3Kz07_0),.din(w_dff_A_6WIGjWsv7_0),.clk(gclk));
	jdff dff_A_kgYb3Kz07_0(.dout(w_dff_A_7zLEWMT62_0),.din(w_dff_A_kgYb3Kz07_0),.clk(gclk));
	jdff dff_A_7zLEWMT62_0(.dout(w_dff_A_xHjP5IS19_0),.din(w_dff_A_7zLEWMT62_0),.clk(gclk));
	jdff dff_A_xHjP5IS19_0(.dout(G606),.din(w_dff_A_xHjP5IS19_0),.clk(gclk));
	jdff dff_A_TeUGITqX2_2(.dout(w_dff_A_ZCWtzJSQ0_0),.din(w_dff_A_TeUGITqX2_2),.clk(gclk));
	jdff dff_A_ZCWtzJSQ0_0(.dout(w_dff_A_FB0ppcoU5_0),.din(w_dff_A_ZCWtzJSQ0_0),.clk(gclk));
	jdff dff_A_FB0ppcoU5_0(.dout(w_dff_A_dprZnLz11_0),.din(w_dff_A_FB0ppcoU5_0),.clk(gclk));
	jdff dff_A_dprZnLz11_0(.dout(w_dff_A_Rz8X0FA01_0),.din(w_dff_A_dprZnLz11_0),.clk(gclk));
	jdff dff_A_Rz8X0FA01_0(.dout(w_dff_A_GMOGhMJd9_0),.din(w_dff_A_Rz8X0FA01_0),.clk(gclk));
	jdff dff_A_GMOGhMJd9_0(.dout(w_dff_A_UlIXDjWl3_0),.din(w_dff_A_GMOGhMJd9_0),.clk(gclk));
	jdff dff_A_UlIXDjWl3_0(.dout(w_dff_A_r09MFtEO1_0),.din(w_dff_A_UlIXDjWl3_0),.clk(gclk));
	jdff dff_A_r09MFtEO1_0(.dout(w_dff_A_BIZe2Idh7_0),.din(w_dff_A_r09MFtEO1_0),.clk(gclk));
	jdff dff_A_BIZe2Idh7_0(.dout(w_dff_A_pSDFP8IT6_0),.din(w_dff_A_BIZe2Idh7_0),.clk(gclk));
	jdff dff_A_pSDFP8IT6_0(.dout(w_dff_A_GuPYyWVO8_0),.din(w_dff_A_pSDFP8IT6_0),.clk(gclk));
	jdff dff_A_GuPYyWVO8_0(.dout(w_dff_A_3qr1ixEV8_0),.din(w_dff_A_GuPYyWVO8_0),.clk(gclk));
	jdff dff_A_3qr1ixEV8_0(.dout(w_dff_A_XfhO3DZo7_0),.din(w_dff_A_3qr1ixEV8_0),.clk(gclk));
	jdff dff_A_XfhO3DZo7_0(.dout(w_dff_A_fGRjIBvF9_0),.din(w_dff_A_XfhO3DZo7_0),.clk(gclk));
	jdff dff_A_fGRjIBvF9_0(.dout(w_dff_A_P83KR6rp4_0),.din(w_dff_A_fGRjIBvF9_0),.clk(gclk));
	jdff dff_A_P83KR6rp4_0(.dout(w_dff_A_3IKFuf0c0_0),.din(w_dff_A_P83KR6rp4_0),.clk(gclk));
	jdff dff_A_3IKFuf0c0_0(.dout(w_dff_A_EFgaN5sF1_0),.din(w_dff_A_3IKFuf0c0_0),.clk(gclk));
	jdff dff_A_EFgaN5sF1_0(.dout(w_dff_A_XnDof0qX9_0),.din(w_dff_A_EFgaN5sF1_0),.clk(gclk));
	jdff dff_A_XnDof0qX9_0(.dout(w_dff_A_VgPj72L81_0),.din(w_dff_A_XnDof0qX9_0),.clk(gclk));
	jdff dff_A_VgPj72L81_0(.dout(w_dff_A_Y4mUHlXV0_0),.din(w_dff_A_VgPj72L81_0),.clk(gclk));
	jdff dff_A_Y4mUHlXV0_0(.dout(w_dff_A_Sur98lIL2_0),.din(w_dff_A_Y4mUHlXV0_0),.clk(gclk));
	jdff dff_A_Sur98lIL2_0(.dout(w_dff_A_hv8wnq873_0),.din(w_dff_A_Sur98lIL2_0),.clk(gclk));
	jdff dff_A_hv8wnq873_0(.dout(w_dff_A_3P1pUxhw8_0),.din(w_dff_A_hv8wnq873_0),.clk(gclk));
	jdff dff_A_3P1pUxhw8_0(.dout(G656),.din(w_dff_A_3P1pUxhw8_0),.clk(gclk));
	jdff dff_A_j3HNxQs77_2(.dout(w_dff_A_Ts6Jurkj7_0),.din(w_dff_A_j3HNxQs77_2),.clk(gclk));
	jdff dff_A_Ts6Jurkj7_0(.dout(w_dff_A_nK0AWwSp4_0),.din(w_dff_A_Ts6Jurkj7_0),.clk(gclk));
	jdff dff_A_nK0AWwSp4_0(.dout(w_dff_A_2UtaPUNn0_0),.din(w_dff_A_nK0AWwSp4_0),.clk(gclk));
	jdff dff_A_2UtaPUNn0_0(.dout(w_dff_A_A2bSnDeh5_0),.din(w_dff_A_2UtaPUNn0_0),.clk(gclk));
	jdff dff_A_A2bSnDeh5_0(.dout(w_dff_A_xnDITRUY1_0),.din(w_dff_A_A2bSnDeh5_0),.clk(gclk));
	jdff dff_A_xnDITRUY1_0(.dout(w_dff_A_pmuwjlej6_0),.din(w_dff_A_xnDITRUY1_0),.clk(gclk));
	jdff dff_A_pmuwjlej6_0(.dout(w_dff_A_sqWnpmwm9_0),.din(w_dff_A_pmuwjlej6_0),.clk(gclk));
	jdff dff_A_sqWnpmwm9_0(.dout(w_dff_A_RrO9wq0O9_0),.din(w_dff_A_sqWnpmwm9_0),.clk(gclk));
	jdff dff_A_RrO9wq0O9_0(.dout(w_dff_A_G5CRzuJP7_0),.din(w_dff_A_RrO9wq0O9_0),.clk(gclk));
	jdff dff_A_G5CRzuJP7_0(.dout(w_dff_A_vQDry5gr4_0),.din(w_dff_A_G5CRzuJP7_0),.clk(gclk));
	jdff dff_A_vQDry5gr4_0(.dout(w_dff_A_Z1Q08JJD2_0),.din(w_dff_A_vQDry5gr4_0),.clk(gclk));
	jdff dff_A_Z1Q08JJD2_0(.dout(w_dff_A_TFX58myf6_0),.din(w_dff_A_Z1Q08JJD2_0),.clk(gclk));
	jdff dff_A_TFX58myf6_0(.dout(w_dff_A_iJbLTe5r2_0),.din(w_dff_A_TFX58myf6_0),.clk(gclk));
	jdff dff_A_iJbLTe5r2_0(.dout(w_dff_A_77SJkW3d7_0),.din(w_dff_A_iJbLTe5r2_0),.clk(gclk));
	jdff dff_A_77SJkW3d7_0(.dout(w_dff_A_HDs3TPly7_0),.din(w_dff_A_77SJkW3d7_0),.clk(gclk));
	jdff dff_A_HDs3TPly7_0(.dout(w_dff_A_PHcTUTMS3_0),.din(w_dff_A_HDs3TPly7_0),.clk(gclk));
	jdff dff_A_PHcTUTMS3_0(.dout(w_dff_A_X8316fVC6_0),.din(w_dff_A_PHcTUTMS3_0),.clk(gclk));
	jdff dff_A_X8316fVC6_0(.dout(w_dff_A_9angCHJB9_0),.din(w_dff_A_X8316fVC6_0),.clk(gclk));
	jdff dff_A_9angCHJB9_0(.dout(w_dff_A_gaDTap2v7_0),.din(w_dff_A_9angCHJB9_0),.clk(gclk));
	jdff dff_A_gaDTap2v7_0(.dout(w_dff_A_avJB5NEK5_0),.din(w_dff_A_gaDTap2v7_0),.clk(gclk));
	jdff dff_A_avJB5NEK5_0(.dout(w_dff_A_gNvvd1LB5_0),.din(w_dff_A_avJB5NEK5_0),.clk(gclk));
	jdff dff_A_gNvvd1LB5_0(.dout(w_dff_A_XdcOMGSy6_0),.din(w_dff_A_gNvvd1LB5_0),.clk(gclk));
	jdff dff_A_XdcOMGSy6_0(.dout(w_dff_A_BV1QvbK34_0),.din(w_dff_A_XdcOMGSy6_0),.clk(gclk));
	jdff dff_A_BV1QvbK34_0(.dout(G809),.din(w_dff_A_BV1QvbK34_0),.clk(gclk));
	jdff dff_A_souf8wzQ9_1(.dout(w_dff_A_sohbHvtO3_0),.din(w_dff_A_souf8wzQ9_1),.clk(gclk));
	jdff dff_A_sohbHvtO3_0(.dout(w_dff_A_1hlssLp53_0),.din(w_dff_A_sohbHvtO3_0),.clk(gclk));
	jdff dff_A_1hlssLp53_0(.dout(w_dff_A_56rwGcC02_0),.din(w_dff_A_1hlssLp53_0),.clk(gclk));
	jdff dff_A_56rwGcC02_0(.dout(w_dff_A_cNgu48bF9_0),.din(w_dff_A_56rwGcC02_0),.clk(gclk));
	jdff dff_A_cNgu48bF9_0(.dout(w_dff_A_8I3ladya6_0),.din(w_dff_A_cNgu48bF9_0),.clk(gclk));
	jdff dff_A_8I3ladya6_0(.dout(w_dff_A_XMMLbFry8_0),.din(w_dff_A_8I3ladya6_0),.clk(gclk));
	jdff dff_A_XMMLbFry8_0(.dout(w_dff_A_dTQuhFCU0_0),.din(w_dff_A_XMMLbFry8_0),.clk(gclk));
	jdff dff_A_dTQuhFCU0_0(.dout(w_dff_A_eoLUDWS09_0),.din(w_dff_A_dTQuhFCU0_0),.clk(gclk));
	jdff dff_A_eoLUDWS09_0(.dout(w_dff_A_SsN5C4260_0),.din(w_dff_A_eoLUDWS09_0),.clk(gclk));
	jdff dff_A_SsN5C4260_0(.dout(w_dff_A_Va0eIH452_0),.din(w_dff_A_SsN5C4260_0),.clk(gclk));
	jdff dff_A_Va0eIH452_0(.dout(w_dff_A_zTDQF9uP0_0),.din(w_dff_A_Va0eIH452_0),.clk(gclk));
	jdff dff_A_zTDQF9uP0_0(.dout(w_dff_A_qMzMVPyK5_0),.din(w_dff_A_zTDQF9uP0_0),.clk(gclk));
	jdff dff_A_qMzMVPyK5_0(.dout(w_dff_A_SKNZPdFB0_0),.din(w_dff_A_qMzMVPyK5_0),.clk(gclk));
	jdff dff_A_SKNZPdFB0_0(.dout(w_dff_A_hRGfadrq8_0),.din(w_dff_A_SKNZPdFB0_0),.clk(gclk));
	jdff dff_A_hRGfadrq8_0(.dout(w_dff_A_yqKAlLtL1_0),.din(w_dff_A_hRGfadrq8_0),.clk(gclk));
	jdff dff_A_yqKAlLtL1_0(.dout(w_dff_A_CT5Xi9Sc4_0),.din(w_dff_A_yqKAlLtL1_0),.clk(gclk));
	jdff dff_A_CT5Xi9Sc4_0(.dout(w_dff_A_Tu7SSuAh3_0),.din(w_dff_A_CT5Xi9Sc4_0),.clk(gclk));
	jdff dff_A_Tu7SSuAh3_0(.dout(w_dff_A_tWKfunQL0_0),.din(w_dff_A_Tu7SSuAh3_0),.clk(gclk));
	jdff dff_A_tWKfunQL0_0(.dout(w_dff_A_FMxVe5KS4_0),.din(w_dff_A_tWKfunQL0_0),.clk(gclk));
	jdff dff_A_FMxVe5KS4_0(.dout(w_dff_A_TUaljnmm9_0),.din(w_dff_A_FMxVe5KS4_0),.clk(gclk));
	jdff dff_A_TUaljnmm9_0(.dout(w_dff_A_NYjwMUd90_0),.din(w_dff_A_TUaljnmm9_0),.clk(gclk));
	jdff dff_A_NYjwMUd90_0(.dout(w_dff_A_xYxAgG1G7_0),.din(w_dff_A_NYjwMUd90_0),.clk(gclk));
	jdff dff_A_xYxAgG1G7_0(.dout(w_dff_A_VXAjTzj17_0),.din(w_dff_A_xYxAgG1G7_0),.clk(gclk));
	jdff dff_A_VXAjTzj17_0(.dout(w_dff_A_hJTCLf5r2_0),.din(w_dff_A_VXAjTzj17_0),.clk(gclk));
	jdff dff_A_hJTCLf5r2_0(.dout(w_dff_A_iRIb9Db31_0),.din(w_dff_A_hJTCLf5r2_0),.clk(gclk));
	jdff dff_A_iRIb9Db31_0(.dout(G993),.din(w_dff_A_iRIb9Db31_0),.clk(gclk));
	jdff dff_A_ezKNDcPo0_1(.dout(w_dff_A_kTjnUn804_0),.din(w_dff_A_ezKNDcPo0_1),.clk(gclk));
	jdff dff_A_kTjnUn804_0(.dout(w_dff_A_ypujY40A4_0),.din(w_dff_A_kTjnUn804_0),.clk(gclk));
	jdff dff_A_ypujY40A4_0(.dout(w_dff_A_OsNx4ymZ7_0),.din(w_dff_A_ypujY40A4_0),.clk(gclk));
	jdff dff_A_OsNx4ymZ7_0(.dout(w_dff_A_8zcrnIHL0_0),.din(w_dff_A_OsNx4ymZ7_0),.clk(gclk));
	jdff dff_A_8zcrnIHL0_0(.dout(w_dff_A_YOUzHR8T8_0),.din(w_dff_A_8zcrnIHL0_0),.clk(gclk));
	jdff dff_A_YOUzHR8T8_0(.dout(w_dff_A_OCLBUumw8_0),.din(w_dff_A_YOUzHR8T8_0),.clk(gclk));
	jdff dff_A_OCLBUumw8_0(.dout(w_dff_A_NJjdlZkG5_0),.din(w_dff_A_OCLBUumw8_0),.clk(gclk));
	jdff dff_A_NJjdlZkG5_0(.dout(w_dff_A_eOvvMheU8_0),.din(w_dff_A_NJjdlZkG5_0),.clk(gclk));
	jdff dff_A_eOvvMheU8_0(.dout(w_dff_A_eLgRBT7h4_0),.din(w_dff_A_eOvvMheU8_0),.clk(gclk));
	jdff dff_A_eLgRBT7h4_0(.dout(w_dff_A_Wvf1Pxkn8_0),.din(w_dff_A_eLgRBT7h4_0),.clk(gclk));
	jdff dff_A_Wvf1Pxkn8_0(.dout(w_dff_A_lnqTQAeb4_0),.din(w_dff_A_Wvf1Pxkn8_0),.clk(gclk));
	jdff dff_A_lnqTQAeb4_0(.dout(w_dff_A_CuEQSgoi6_0),.din(w_dff_A_lnqTQAeb4_0),.clk(gclk));
	jdff dff_A_CuEQSgoi6_0(.dout(w_dff_A_nfTbMoVz2_0),.din(w_dff_A_CuEQSgoi6_0),.clk(gclk));
	jdff dff_A_nfTbMoVz2_0(.dout(w_dff_A_NDjX91AQ8_0),.din(w_dff_A_nfTbMoVz2_0),.clk(gclk));
	jdff dff_A_NDjX91AQ8_0(.dout(w_dff_A_zFNT25fk3_0),.din(w_dff_A_NDjX91AQ8_0),.clk(gclk));
	jdff dff_A_zFNT25fk3_0(.dout(w_dff_A_Da44n6E71_0),.din(w_dff_A_zFNT25fk3_0),.clk(gclk));
	jdff dff_A_Da44n6E71_0(.dout(w_dff_A_pFs9W2I26_0),.din(w_dff_A_Da44n6E71_0),.clk(gclk));
	jdff dff_A_pFs9W2I26_0(.dout(w_dff_A_ANyzpBGA6_0),.din(w_dff_A_pFs9W2I26_0),.clk(gclk));
	jdff dff_A_ANyzpBGA6_0(.dout(w_dff_A_Zx3Z1ZgQ9_0),.din(w_dff_A_ANyzpBGA6_0),.clk(gclk));
	jdff dff_A_Zx3Z1ZgQ9_0(.dout(w_dff_A_uHNbxmZ29_0),.din(w_dff_A_Zx3Z1ZgQ9_0),.clk(gclk));
	jdff dff_A_uHNbxmZ29_0(.dout(w_dff_A_QUweVljw1_0),.din(w_dff_A_uHNbxmZ29_0),.clk(gclk));
	jdff dff_A_QUweVljw1_0(.dout(w_dff_A_TGETJrkQ3_0),.din(w_dff_A_QUweVljw1_0),.clk(gclk));
	jdff dff_A_TGETJrkQ3_0(.dout(w_dff_A_GbRv2wqN1_0),.din(w_dff_A_TGETJrkQ3_0),.clk(gclk));
	jdff dff_A_GbRv2wqN1_0(.dout(w_dff_A_RTci2qEH8_0),.din(w_dff_A_GbRv2wqN1_0),.clk(gclk));
	jdff dff_A_RTci2qEH8_0(.dout(w_dff_A_8gEV0b435_0),.din(w_dff_A_RTci2qEH8_0),.clk(gclk));
	jdff dff_A_8gEV0b435_0(.dout(G978),.din(w_dff_A_8gEV0b435_0),.clk(gclk));
	jdff dff_A_FmBKNEEe6_1(.dout(w_dff_A_uHjSMvx90_0),.din(w_dff_A_FmBKNEEe6_1),.clk(gclk));
	jdff dff_A_uHjSMvx90_0(.dout(w_dff_A_MtrizcXo7_0),.din(w_dff_A_uHjSMvx90_0),.clk(gclk));
	jdff dff_A_MtrizcXo7_0(.dout(w_dff_A_JHPeRswh6_0),.din(w_dff_A_MtrizcXo7_0),.clk(gclk));
	jdff dff_A_JHPeRswh6_0(.dout(w_dff_A_s2Wbzplc0_0),.din(w_dff_A_JHPeRswh6_0),.clk(gclk));
	jdff dff_A_s2Wbzplc0_0(.dout(w_dff_A_9xtsbFfg2_0),.din(w_dff_A_s2Wbzplc0_0),.clk(gclk));
	jdff dff_A_9xtsbFfg2_0(.dout(w_dff_A_4niLbNtt5_0),.din(w_dff_A_9xtsbFfg2_0),.clk(gclk));
	jdff dff_A_4niLbNtt5_0(.dout(w_dff_A_I3ZjgZK78_0),.din(w_dff_A_4niLbNtt5_0),.clk(gclk));
	jdff dff_A_I3ZjgZK78_0(.dout(w_dff_A_SXGMLNcz5_0),.din(w_dff_A_I3ZjgZK78_0),.clk(gclk));
	jdff dff_A_SXGMLNcz5_0(.dout(w_dff_A_FZoCUiy34_0),.din(w_dff_A_SXGMLNcz5_0),.clk(gclk));
	jdff dff_A_FZoCUiy34_0(.dout(w_dff_A_yap5GLYK3_0),.din(w_dff_A_FZoCUiy34_0),.clk(gclk));
	jdff dff_A_yap5GLYK3_0(.dout(w_dff_A_gyNZpwcy1_0),.din(w_dff_A_yap5GLYK3_0),.clk(gclk));
	jdff dff_A_gyNZpwcy1_0(.dout(w_dff_A_en156vvS4_0),.din(w_dff_A_gyNZpwcy1_0),.clk(gclk));
	jdff dff_A_en156vvS4_0(.dout(w_dff_A_AfeoRSEh3_0),.din(w_dff_A_en156vvS4_0),.clk(gclk));
	jdff dff_A_AfeoRSEh3_0(.dout(w_dff_A_x8giCt9r2_0),.din(w_dff_A_AfeoRSEh3_0),.clk(gclk));
	jdff dff_A_x8giCt9r2_0(.dout(w_dff_A_dRtqPKuB3_0),.din(w_dff_A_x8giCt9r2_0),.clk(gclk));
	jdff dff_A_dRtqPKuB3_0(.dout(w_dff_A_pFqz7zf01_0),.din(w_dff_A_dRtqPKuB3_0),.clk(gclk));
	jdff dff_A_pFqz7zf01_0(.dout(w_dff_A_hz3Cv4bT7_0),.din(w_dff_A_pFqz7zf01_0),.clk(gclk));
	jdff dff_A_hz3Cv4bT7_0(.dout(w_dff_A_YzRnybzk7_0),.din(w_dff_A_hz3Cv4bT7_0),.clk(gclk));
	jdff dff_A_YzRnybzk7_0(.dout(w_dff_A_rqQ9f4I73_0),.din(w_dff_A_YzRnybzk7_0),.clk(gclk));
	jdff dff_A_rqQ9f4I73_0(.dout(w_dff_A_eTohmUmJ5_0),.din(w_dff_A_rqQ9f4I73_0),.clk(gclk));
	jdff dff_A_eTohmUmJ5_0(.dout(w_dff_A_tlembwPc2_0),.din(w_dff_A_eTohmUmJ5_0),.clk(gclk));
	jdff dff_A_tlembwPc2_0(.dout(w_dff_A_oynZh5sH8_0),.din(w_dff_A_tlembwPc2_0),.clk(gclk));
	jdff dff_A_oynZh5sH8_0(.dout(w_dff_A_7NQSHuoH9_0),.din(w_dff_A_oynZh5sH8_0),.clk(gclk));
	jdff dff_A_7NQSHuoH9_0(.dout(w_dff_A_7qS01c9g8_0),.din(w_dff_A_7NQSHuoH9_0),.clk(gclk));
	jdff dff_A_7qS01c9g8_0(.dout(w_dff_A_8itBNWBZ5_0),.din(w_dff_A_7qS01c9g8_0),.clk(gclk));
	jdff dff_A_8itBNWBZ5_0(.dout(G949),.din(w_dff_A_8itBNWBZ5_0),.clk(gclk));
	jdff dff_A_nZRgG5262_1(.dout(w_dff_A_n0DEsO647_0),.din(w_dff_A_nZRgG5262_1),.clk(gclk));
	jdff dff_A_n0DEsO647_0(.dout(w_dff_A_NxA3MFIe6_0),.din(w_dff_A_n0DEsO647_0),.clk(gclk));
	jdff dff_A_NxA3MFIe6_0(.dout(w_dff_A_Bxlv6EiW3_0),.din(w_dff_A_NxA3MFIe6_0),.clk(gclk));
	jdff dff_A_Bxlv6EiW3_0(.dout(w_dff_A_EMW9azd01_0),.din(w_dff_A_Bxlv6EiW3_0),.clk(gclk));
	jdff dff_A_EMW9azd01_0(.dout(w_dff_A_Sbput8P13_0),.din(w_dff_A_EMW9azd01_0),.clk(gclk));
	jdff dff_A_Sbput8P13_0(.dout(w_dff_A_u7iNuL7L9_0),.din(w_dff_A_Sbput8P13_0),.clk(gclk));
	jdff dff_A_u7iNuL7L9_0(.dout(w_dff_A_7r5mLf335_0),.din(w_dff_A_u7iNuL7L9_0),.clk(gclk));
	jdff dff_A_7r5mLf335_0(.dout(w_dff_A_oTyKjcqZ7_0),.din(w_dff_A_7r5mLf335_0),.clk(gclk));
	jdff dff_A_oTyKjcqZ7_0(.dout(w_dff_A_BkCOtPlg8_0),.din(w_dff_A_oTyKjcqZ7_0),.clk(gclk));
	jdff dff_A_BkCOtPlg8_0(.dout(w_dff_A_u9XL9JiD6_0),.din(w_dff_A_BkCOtPlg8_0),.clk(gclk));
	jdff dff_A_u9XL9JiD6_0(.dout(w_dff_A_Qd88GtDw2_0),.din(w_dff_A_u9XL9JiD6_0),.clk(gclk));
	jdff dff_A_Qd88GtDw2_0(.dout(w_dff_A_LftG2yA64_0),.din(w_dff_A_Qd88GtDw2_0),.clk(gclk));
	jdff dff_A_LftG2yA64_0(.dout(w_dff_A_ZuijdhyB5_0),.din(w_dff_A_LftG2yA64_0),.clk(gclk));
	jdff dff_A_ZuijdhyB5_0(.dout(w_dff_A_i2dPcf8c3_0),.din(w_dff_A_ZuijdhyB5_0),.clk(gclk));
	jdff dff_A_i2dPcf8c3_0(.dout(w_dff_A_1v6fKkZt6_0),.din(w_dff_A_i2dPcf8c3_0),.clk(gclk));
	jdff dff_A_1v6fKkZt6_0(.dout(w_dff_A_SsNQQLZ38_0),.din(w_dff_A_1v6fKkZt6_0),.clk(gclk));
	jdff dff_A_SsNQQLZ38_0(.dout(w_dff_A_M4wsOCKc6_0),.din(w_dff_A_SsNQQLZ38_0),.clk(gclk));
	jdff dff_A_M4wsOCKc6_0(.dout(w_dff_A_1kPZT8yf6_0),.din(w_dff_A_M4wsOCKc6_0),.clk(gclk));
	jdff dff_A_1kPZT8yf6_0(.dout(w_dff_A_f0tGfCn38_0),.din(w_dff_A_1kPZT8yf6_0),.clk(gclk));
	jdff dff_A_f0tGfCn38_0(.dout(w_dff_A_irplmtP10_0),.din(w_dff_A_f0tGfCn38_0),.clk(gclk));
	jdff dff_A_irplmtP10_0(.dout(w_dff_A_UU2y8qZI4_0),.din(w_dff_A_irplmtP10_0),.clk(gclk));
	jdff dff_A_UU2y8qZI4_0(.dout(w_dff_A_WDG89NpS6_0),.din(w_dff_A_UU2y8qZI4_0),.clk(gclk));
	jdff dff_A_WDG89NpS6_0(.dout(w_dff_A_lSmUJkuW6_0),.din(w_dff_A_WDG89NpS6_0),.clk(gclk));
	jdff dff_A_lSmUJkuW6_0(.dout(w_dff_A_sRiGetB06_0),.din(w_dff_A_lSmUJkuW6_0),.clk(gclk));
	jdff dff_A_sRiGetB06_0(.dout(w_dff_A_p9zxiRJd1_0),.din(w_dff_A_sRiGetB06_0),.clk(gclk));
	jdff dff_A_p9zxiRJd1_0(.dout(G939),.din(w_dff_A_p9zxiRJd1_0),.clk(gclk));
	jdff dff_A_eXIkQR0I3_1(.dout(w_dff_A_LU4KLaQz4_0),.din(w_dff_A_eXIkQR0I3_1),.clk(gclk));
	jdff dff_A_LU4KLaQz4_0(.dout(w_dff_A_kXyhF1CE8_0),.din(w_dff_A_LU4KLaQz4_0),.clk(gclk));
	jdff dff_A_kXyhF1CE8_0(.dout(w_dff_A_nY08GLQu3_0),.din(w_dff_A_kXyhF1CE8_0),.clk(gclk));
	jdff dff_A_nY08GLQu3_0(.dout(w_dff_A_ZFvPONps7_0),.din(w_dff_A_nY08GLQu3_0),.clk(gclk));
	jdff dff_A_ZFvPONps7_0(.dout(w_dff_A_cajAvpJP8_0),.din(w_dff_A_ZFvPONps7_0),.clk(gclk));
	jdff dff_A_cajAvpJP8_0(.dout(w_dff_A_Om81QiMW5_0),.din(w_dff_A_cajAvpJP8_0),.clk(gclk));
	jdff dff_A_Om81QiMW5_0(.dout(w_dff_A_N6G5mIwj7_0),.din(w_dff_A_Om81QiMW5_0),.clk(gclk));
	jdff dff_A_N6G5mIwj7_0(.dout(w_dff_A_sYLLraH33_0),.din(w_dff_A_N6G5mIwj7_0),.clk(gclk));
	jdff dff_A_sYLLraH33_0(.dout(w_dff_A_n8riWIWi9_0),.din(w_dff_A_sYLLraH33_0),.clk(gclk));
	jdff dff_A_n8riWIWi9_0(.dout(w_dff_A_GcRCZb8I2_0),.din(w_dff_A_n8riWIWi9_0),.clk(gclk));
	jdff dff_A_GcRCZb8I2_0(.dout(w_dff_A_2G98fjIZ7_0),.din(w_dff_A_GcRCZb8I2_0),.clk(gclk));
	jdff dff_A_2G98fjIZ7_0(.dout(w_dff_A_jz2AJcTg0_0),.din(w_dff_A_2G98fjIZ7_0),.clk(gclk));
	jdff dff_A_jz2AJcTg0_0(.dout(w_dff_A_QWZmy7Hx4_0),.din(w_dff_A_jz2AJcTg0_0),.clk(gclk));
	jdff dff_A_QWZmy7Hx4_0(.dout(w_dff_A_33uK8JQk4_0),.din(w_dff_A_QWZmy7Hx4_0),.clk(gclk));
	jdff dff_A_33uK8JQk4_0(.dout(w_dff_A_mGRRoOep8_0),.din(w_dff_A_33uK8JQk4_0),.clk(gclk));
	jdff dff_A_mGRRoOep8_0(.dout(w_dff_A_MxJ6BjHc7_0),.din(w_dff_A_mGRRoOep8_0),.clk(gclk));
	jdff dff_A_MxJ6BjHc7_0(.dout(w_dff_A_GX7WeA8R7_0),.din(w_dff_A_MxJ6BjHc7_0),.clk(gclk));
	jdff dff_A_GX7WeA8R7_0(.dout(w_dff_A_wpCDQzop7_0),.din(w_dff_A_GX7WeA8R7_0),.clk(gclk));
	jdff dff_A_wpCDQzop7_0(.dout(w_dff_A_PDL2VOF95_0),.din(w_dff_A_wpCDQzop7_0),.clk(gclk));
	jdff dff_A_PDL2VOF95_0(.dout(w_dff_A_ZDLqX4uF2_0),.din(w_dff_A_PDL2VOF95_0),.clk(gclk));
	jdff dff_A_ZDLqX4uF2_0(.dout(w_dff_A_u8bgHKvf1_0),.din(w_dff_A_ZDLqX4uF2_0),.clk(gclk));
	jdff dff_A_u8bgHKvf1_0(.dout(w_dff_A_dGBChYzy0_0),.din(w_dff_A_u8bgHKvf1_0),.clk(gclk));
	jdff dff_A_dGBChYzy0_0(.dout(w_dff_A_FG7jujTQ9_0),.din(w_dff_A_dGBChYzy0_0),.clk(gclk));
	jdff dff_A_FG7jujTQ9_0(.dout(w_dff_A_RC6yfMHf3_0),.din(w_dff_A_FG7jujTQ9_0),.clk(gclk));
	jdff dff_A_RC6yfMHf3_0(.dout(w_dff_A_envOpYwf6_0),.din(w_dff_A_RC6yfMHf3_0),.clk(gclk));
	jdff dff_A_envOpYwf6_0(.dout(G889),.din(w_dff_A_envOpYwf6_0),.clk(gclk));
	jdff dff_A_KMUkwXSO1_1(.dout(w_dff_A_89a6khRD5_0),.din(w_dff_A_KMUkwXSO1_1),.clk(gclk));
	jdff dff_A_89a6khRD5_0(.dout(w_dff_A_t7KoX3Mz3_0),.din(w_dff_A_89a6khRD5_0),.clk(gclk));
	jdff dff_A_t7KoX3Mz3_0(.dout(w_dff_A_UNcfpJRv2_0),.din(w_dff_A_t7KoX3Mz3_0),.clk(gclk));
	jdff dff_A_UNcfpJRv2_0(.dout(w_dff_A_iab2UFPQ0_0),.din(w_dff_A_UNcfpJRv2_0),.clk(gclk));
	jdff dff_A_iab2UFPQ0_0(.dout(w_dff_A_uYkEWure5_0),.din(w_dff_A_iab2UFPQ0_0),.clk(gclk));
	jdff dff_A_uYkEWure5_0(.dout(w_dff_A_F3iC9brH9_0),.din(w_dff_A_uYkEWure5_0),.clk(gclk));
	jdff dff_A_F3iC9brH9_0(.dout(w_dff_A_HUxslvW57_0),.din(w_dff_A_F3iC9brH9_0),.clk(gclk));
	jdff dff_A_HUxslvW57_0(.dout(w_dff_A_xp9gBtPA6_0),.din(w_dff_A_HUxslvW57_0),.clk(gclk));
	jdff dff_A_xp9gBtPA6_0(.dout(w_dff_A_mEcvr3lh2_0),.din(w_dff_A_xp9gBtPA6_0),.clk(gclk));
	jdff dff_A_mEcvr3lh2_0(.dout(w_dff_A_uf2sLu1l1_0),.din(w_dff_A_mEcvr3lh2_0),.clk(gclk));
	jdff dff_A_uf2sLu1l1_0(.dout(w_dff_A_4Wsui3iD7_0),.din(w_dff_A_uf2sLu1l1_0),.clk(gclk));
	jdff dff_A_4Wsui3iD7_0(.dout(w_dff_A_yx5CXPkn7_0),.din(w_dff_A_4Wsui3iD7_0),.clk(gclk));
	jdff dff_A_yx5CXPkn7_0(.dout(w_dff_A_ZdgZX82D2_0),.din(w_dff_A_yx5CXPkn7_0),.clk(gclk));
	jdff dff_A_ZdgZX82D2_0(.dout(w_dff_A_y5NJj0W41_0),.din(w_dff_A_ZdgZX82D2_0),.clk(gclk));
	jdff dff_A_y5NJj0W41_0(.dout(w_dff_A_4nWin5EN5_0),.din(w_dff_A_y5NJj0W41_0),.clk(gclk));
	jdff dff_A_4nWin5EN5_0(.dout(w_dff_A_JYYNbSlL3_0),.din(w_dff_A_4nWin5EN5_0),.clk(gclk));
	jdff dff_A_JYYNbSlL3_0(.dout(w_dff_A_rkXzrh7J8_0),.din(w_dff_A_JYYNbSlL3_0),.clk(gclk));
	jdff dff_A_rkXzrh7J8_0(.dout(w_dff_A_3BXvPA8k1_0),.din(w_dff_A_rkXzrh7J8_0),.clk(gclk));
	jdff dff_A_3BXvPA8k1_0(.dout(w_dff_A_eTTwXyHP5_0),.din(w_dff_A_3BXvPA8k1_0),.clk(gclk));
	jdff dff_A_eTTwXyHP5_0(.dout(w_dff_A_MX4lXgeB5_0),.din(w_dff_A_eTTwXyHP5_0),.clk(gclk));
	jdff dff_A_MX4lXgeB5_0(.dout(w_dff_A_13nVuEtI9_0),.din(w_dff_A_MX4lXgeB5_0),.clk(gclk));
	jdff dff_A_13nVuEtI9_0(.dout(w_dff_A_RkqjJyFY5_0),.din(w_dff_A_13nVuEtI9_0),.clk(gclk));
	jdff dff_A_RkqjJyFY5_0(.dout(w_dff_A_8jLSMEHM0_0),.din(w_dff_A_RkqjJyFY5_0),.clk(gclk));
	jdff dff_A_8jLSMEHM0_0(.dout(w_dff_A_OYwj7SfF3_0),.din(w_dff_A_8jLSMEHM0_0),.clk(gclk));
	jdff dff_A_OYwj7SfF3_0(.dout(G593),.din(w_dff_A_OYwj7SfF3_0),.clk(gclk));
	jdff dff_A_he6umlfr2_2(.dout(w_dff_A_sexO35Lf7_0),.din(w_dff_A_he6umlfr2_2),.clk(gclk));
	jdff dff_A_sexO35Lf7_0(.dout(w_dff_A_AgcW8LBO0_0),.din(w_dff_A_sexO35Lf7_0),.clk(gclk));
	jdff dff_A_AgcW8LBO0_0(.dout(w_dff_A_mMV86RFB5_0),.din(w_dff_A_AgcW8LBO0_0),.clk(gclk));
	jdff dff_A_mMV86RFB5_0(.dout(w_dff_A_ty5sv9pU7_0),.din(w_dff_A_mMV86RFB5_0),.clk(gclk));
	jdff dff_A_ty5sv9pU7_0(.dout(w_dff_A_lnJ1U2dA9_0),.din(w_dff_A_ty5sv9pU7_0),.clk(gclk));
	jdff dff_A_lnJ1U2dA9_0(.dout(w_dff_A_cwO910r85_0),.din(w_dff_A_lnJ1U2dA9_0),.clk(gclk));
	jdff dff_A_cwO910r85_0(.dout(w_dff_A_6ymS5dNn5_0),.din(w_dff_A_cwO910r85_0),.clk(gclk));
	jdff dff_A_6ymS5dNn5_0(.dout(w_dff_A_CIgUKtGE0_0),.din(w_dff_A_6ymS5dNn5_0),.clk(gclk));
	jdff dff_A_CIgUKtGE0_0(.dout(w_dff_A_mvMVnw3A7_0),.din(w_dff_A_CIgUKtGE0_0),.clk(gclk));
	jdff dff_A_mvMVnw3A7_0(.dout(w_dff_A_WMlCXaE18_0),.din(w_dff_A_mvMVnw3A7_0),.clk(gclk));
	jdff dff_A_WMlCXaE18_0(.dout(w_dff_A_V7Iw77Eo1_0),.din(w_dff_A_WMlCXaE18_0),.clk(gclk));
	jdff dff_A_V7Iw77Eo1_0(.dout(w_dff_A_6gkHl4Gz2_0),.din(w_dff_A_V7Iw77Eo1_0),.clk(gclk));
	jdff dff_A_6gkHl4Gz2_0(.dout(w_dff_A_gxIXcJuF4_0),.din(w_dff_A_6gkHl4Gz2_0),.clk(gclk));
	jdff dff_A_gxIXcJuF4_0(.dout(w_dff_A_HjMMdCrg9_0),.din(w_dff_A_gxIXcJuF4_0),.clk(gclk));
	jdff dff_A_HjMMdCrg9_0(.dout(w_dff_A_fszR8mFn5_0),.din(w_dff_A_HjMMdCrg9_0),.clk(gclk));
	jdff dff_A_fszR8mFn5_0(.dout(w_dff_A_hXjQTx3Z5_0),.din(w_dff_A_fszR8mFn5_0),.clk(gclk));
	jdff dff_A_hXjQTx3Z5_0(.dout(w_dff_A_wBdsQp144_0),.din(w_dff_A_hXjQTx3Z5_0),.clk(gclk));
	jdff dff_A_wBdsQp144_0(.dout(w_dff_A_iSippFl31_0),.din(w_dff_A_wBdsQp144_0),.clk(gclk));
	jdff dff_A_iSippFl31_0(.dout(w_dff_A_sDAWGRxa1_0),.din(w_dff_A_iSippFl31_0),.clk(gclk));
	jdff dff_A_sDAWGRxa1_0(.dout(w_dff_A_23BfwigB4_0),.din(w_dff_A_sDAWGRxa1_0),.clk(gclk));
	jdff dff_A_23BfwigB4_0(.dout(w_dff_A_rNopzjx29_0),.din(w_dff_A_23BfwigB4_0),.clk(gclk));
	jdff dff_A_rNopzjx29_0(.dout(G636),.din(w_dff_A_rNopzjx29_0),.clk(gclk));
	jdff dff_A_NGvHq2GN5_2(.dout(w_dff_A_vNm62C9x0_0),.din(w_dff_A_NGvHq2GN5_2),.clk(gclk));
	jdff dff_A_vNm62C9x0_0(.dout(w_dff_A_vcZGSRff3_0),.din(w_dff_A_vNm62C9x0_0),.clk(gclk));
	jdff dff_A_vcZGSRff3_0(.dout(w_dff_A_vKDY7iSK7_0),.din(w_dff_A_vcZGSRff3_0),.clk(gclk));
	jdff dff_A_vKDY7iSK7_0(.dout(w_dff_A_nMlA0hMx5_0),.din(w_dff_A_vKDY7iSK7_0),.clk(gclk));
	jdff dff_A_nMlA0hMx5_0(.dout(w_dff_A_YAOJots17_0),.din(w_dff_A_nMlA0hMx5_0),.clk(gclk));
	jdff dff_A_YAOJots17_0(.dout(w_dff_A_PAUk9OZU5_0),.din(w_dff_A_YAOJots17_0),.clk(gclk));
	jdff dff_A_PAUk9OZU5_0(.dout(w_dff_A_ryMEEiyR5_0),.din(w_dff_A_PAUk9OZU5_0),.clk(gclk));
	jdff dff_A_ryMEEiyR5_0(.dout(w_dff_A_l0XSivFZ6_0),.din(w_dff_A_ryMEEiyR5_0),.clk(gclk));
	jdff dff_A_l0XSivFZ6_0(.dout(w_dff_A_VV8wepkk8_0),.din(w_dff_A_l0XSivFZ6_0),.clk(gclk));
	jdff dff_A_VV8wepkk8_0(.dout(w_dff_A_8u3yfmOK5_0),.din(w_dff_A_VV8wepkk8_0),.clk(gclk));
	jdff dff_A_8u3yfmOK5_0(.dout(w_dff_A_dVh5TqkM3_0),.din(w_dff_A_8u3yfmOK5_0),.clk(gclk));
	jdff dff_A_dVh5TqkM3_0(.dout(w_dff_A_Pqxdr7IE9_0),.din(w_dff_A_dVh5TqkM3_0),.clk(gclk));
	jdff dff_A_Pqxdr7IE9_0(.dout(w_dff_A_4AChNxay2_0),.din(w_dff_A_Pqxdr7IE9_0),.clk(gclk));
	jdff dff_A_4AChNxay2_0(.dout(w_dff_A_C150Q0tt3_0),.din(w_dff_A_4AChNxay2_0),.clk(gclk));
	jdff dff_A_C150Q0tt3_0(.dout(w_dff_A_9N38gbhl7_0),.din(w_dff_A_C150Q0tt3_0),.clk(gclk));
	jdff dff_A_9N38gbhl7_0(.dout(w_dff_A_0mBXMIi36_0),.din(w_dff_A_9N38gbhl7_0),.clk(gclk));
	jdff dff_A_0mBXMIi36_0(.dout(w_dff_A_wh0uLp1j0_0),.din(w_dff_A_0mBXMIi36_0),.clk(gclk));
	jdff dff_A_wh0uLp1j0_0(.dout(w_dff_A_pOdBPloB2_0),.din(w_dff_A_wh0uLp1j0_0),.clk(gclk));
	jdff dff_A_pOdBPloB2_0(.dout(w_dff_A_BTQsVohP9_0),.din(w_dff_A_pOdBPloB2_0),.clk(gclk));
	jdff dff_A_BTQsVohP9_0(.dout(w_dff_A_7Dqc6S1E0_0),.din(w_dff_A_BTQsVohP9_0),.clk(gclk));
	jdff dff_A_7Dqc6S1E0_0(.dout(w_dff_A_d6dtyzNd9_0),.din(w_dff_A_7Dqc6S1E0_0),.clk(gclk));
	jdff dff_A_d6dtyzNd9_0(.dout(G704),.din(w_dff_A_d6dtyzNd9_0),.clk(gclk));
	jdff dff_A_uUv6KBve7_2(.dout(w_dff_A_EewyZC9F5_0),.din(w_dff_A_uUv6KBve7_2),.clk(gclk));
	jdff dff_A_EewyZC9F5_0(.dout(w_dff_A_VyOlxq200_0),.din(w_dff_A_EewyZC9F5_0),.clk(gclk));
	jdff dff_A_VyOlxq200_0(.dout(w_dff_A_ufqK6YQZ5_0),.din(w_dff_A_VyOlxq200_0),.clk(gclk));
	jdff dff_A_ufqK6YQZ5_0(.dout(w_dff_A_AstLLh6v8_0),.din(w_dff_A_ufqK6YQZ5_0),.clk(gclk));
	jdff dff_A_AstLLh6v8_0(.dout(w_dff_A_Rfi9z38C6_0),.din(w_dff_A_AstLLh6v8_0),.clk(gclk));
	jdff dff_A_Rfi9z38C6_0(.dout(w_dff_A_g0742VEN5_0),.din(w_dff_A_Rfi9z38C6_0),.clk(gclk));
	jdff dff_A_g0742VEN5_0(.dout(w_dff_A_YeRBJudE5_0),.din(w_dff_A_g0742VEN5_0),.clk(gclk));
	jdff dff_A_YeRBJudE5_0(.dout(w_dff_A_r96IHjct1_0),.din(w_dff_A_YeRBJudE5_0),.clk(gclk));
	jdff dff_A_r96IHjct1_0(.dout(w_dff_A_p7ShS8qT7_0),.din(w_dff_A_r96IHjct1_0),.clk(gclk));
	jdff dff_A_p7ShS8qT7_0(.dout(w_dff_A_KvcXPd341_0),.din(w_dff_A_p7ShS8qT7_0),.clk(gclk));
	jdff dff_A_KvcXPd341_0(.dout(w_dff_A_tN0ZeT0k5_0),.din(w_dff_A_KvcXPd341_0),.clk(gclk));
	jdff dff_A_tN0ZeT0k5_0(.dout(w_dff_A_rqYdR5fk6_0),.din(w_dff_A_tN0ZeT0k5_0),.clk(gclk));
	jdff dff_A_rqYdR5fk6_0(.dout(w_dff_A_THHISChu1_0),.din(w_dff_A_rqYdR5fk6_0),.clk(gclk));
	jdff dff_A_THHISChu1_0(.dout(w_dff_A_lXoB0zgw1_0),.din(w_dff_A_THHISChu1_0),.clk(gclk));
	jdff dff_A_lXoB0zgw1_0(.dout(w_dff_A_IY7JPQEK2_0),.din(w_dff_A_lXoB0zgw1_0),.clk(gclk));
	jdff dff_A_IY7JPQEK2_0(.dout(w_dff_A_UYODEuev1_0),.din(w_dff_A_IY7JPQEK2_0),.clk(gclk));
	jdff dff_A_UYODEuev1_0(.dout(w_dff_A_uVaMD4Ke5_0),.din(w_dff_A_UYODEuev1_0),.clk(gclk));
	jdff dff_A_uVaMD4Ke5_0(.dout(w_dff_A_KMrbPvDL8_0),.din(w_dff_A_uVaMD4Ke5_0),.clk(gclk));
	jdff dff_A_KMrbPvDL8_0(.dout(w_dff_A_EjvmdIYi6_0),.din(w_dff_A_KMrbPvDL8_0),.clk(gclk));
	jdff dff_A_EjvmdIYi6_0(.dout(w_dff_A_gogDgxR12_0),.din(w_dff_A_EjvmdIYi6_0),.clk(gclk));
	jdff dff_A_gogDgxR12_0(.dout(w_dff_A_Zo98GRJt8_0),.din(w_dff_A_gogDgxR12_0),.clk(gclk));
	jdff dff_A_Zo98GRJt8_0(.dout(G717),.din(w_dff_A_Zo98GRJt8_0),.clk(gclk));
	jdff dff_A_AJ2uePYK9_2(.dout(w_dff_A_9nfbdfoe2_0),.din(w_dff_A_AJ2uePYK9_2),.clk(gclk));
	jdff dff_A_9nfbdfoe2_0(.dout(w_dff_A_PZbiJtIr9_0),.din(w_dff_A_9nfbdfoe2_0),.clk(gclk));
	jdff dff_A_PZbiJtIr9_0(.dout(w_dff_A_cIx3DeVm6_0),.din(w_dff_A_PZbiJtIr9_0),.clk(gclk));
	jdff dff_A_cIx3DeVm6_0(.dout(w_dff_A_svPrc4Ps7_0),.din(w_dff_A_cIx3DeVm6_0),.clk(gclk));
	jdff dff_A_svPrc4Ps7_0(.dout(w_dff_A_WWGGyxbn3_0),.din(w_dff_A_svPrc4Ps7_0),.clk(gclk));
	jdff dff_A_WWGGyxbn3_0(.dout(w_dff_A_4zeLb0rg3_0),.din(w_dff_A_WWGGyxbn3_0),.clk(gclk));
	jdff dff_A_4zeLb0rg3_0(.dout(w_dff_A_Nyo9VvHv1_0),.din(w_dff_A_4zeLb0rg3_0),.clk(gclk));
	jdff dff_A_Nyo9VvHv1_0(.dout(w_dff_A_e3D1hQGu9_0),.din(w_dff_A_Nyo9VvHv1_0),.clk(gclk));
	jdff dff_A_e3D1hQGu9_0(.dout(w_dff_A_NhqbKtqH8_0),.din(w_dff_A_e3D1hQGu9_0),.clk(gclk));
	jdff dff_A_NhqbKtqH8_0(.dout(w_dff_A_Nztr2vP84_0),.din(w_dff_A_NhqbKtqH8_0),.clk(gclk));
	jdff dff_A_Nztr2vP84_0(.dout(w_dff_A_hsgqY5G03_0),.din(w_dff_A_Nztr2vP84_0),.clk(gclk));
	jdff dff_A_hsgqY5G03_0(.dout(w_dff_A_Xq7WlHVc4_0),.din(w_dff_A_hsgqY5G03_0),.clk(gclk));
	jdff dff_A_Xq7WlHVc4_0(.dout(w_dff_A_ghgonSyV3_0),.din(w_dff_A_Xq7WlHVc4_0),.clk(gclk));
	jdff dff_A_ghgonSyV3_0(.dout(w_dff_A_nfWjngP05_0),.din(w_dff_A_ghgonSyV3_0),.clk(gclk));
	jdff dff_A_nfWjngP05_0(.dout(w_dff_A_EmvpCxco3_0),.din(w_dff_A_nfWjngP05_0),.clk(gclk));
	jdff dff_A_EmvpCxco3_0(.dout(w_dff_A_nERXVkdJ8_0),.din(w_dff_A_EmvpCxco3_0),.clk(gclk));
	jdff dff_A_nERXVkdJ8_0(.dout(w_dff_A_aPRijR0j0_0),.din(w_dff_A_nERXVkdJ8_0),.clk(gclk));
	jdff dff_A_aPRijR0j0_0(.dout(w_dff_A_faV913vR9_0),.din(w_dff_A_aPRijR0j0_0),.clk(gclk));
	jdff dff_A_faV913vR9_0(.dout(w_dff_A_tJjvZw6A3_0),.din(w_dff_A_faV913vR9_0),.clk(gclk));
	jdff dff_A_tJjvZw6A3_0(.dout(w_dff_A_d4dY939z5_0),.din(w_dff_A_tJjvZw6A3_0),.clk(gclk));
	jdff dff_A_d4dY939z5_0(.dout(w_dff_A_VjaejBQp5_0),.din(w_dff_A_d4dY939z5_0),.clk(gclk));
	jdff dff_A_VjaejBQp5_0(.dout(w_dff_A_eBx9In5N7_0),.din(w_dff_A_VjaejBQp5_0),.clk(gclk));
	jdff dff_A_eBx9In5N7_0(.dout(G820),.din(w_dff_A_eBx9In5N7_0),.clk(gclk));
	jdff dff_A_GFQkePVS7_2(.dout(w_dff_A_IuSSsg0Y5_0),.din(w_dff_A_GFQkePVS7_2),.clk(gclk));
	jdff dff_A_IuSSsg0Y5_0(.dout(w_dff_A_K5eCaWLY0_0),.din(w_dff_A_IuSSsg0Y5_0),.clk(gclk));
	jdff dff_A_K5eCaWLY0_0(.dout(w_dff_A_yV3IbMqT1_0),.din(w_dff_A_K5eCaWLY0_0),.clk(gclk));
	jdff dff_A_yV3IbMqT1_0(.dout(w_dff_A_PhUHrHOZ7_0),.din(w_dff_A_yV3IbMqT1_0),.clk(gclk));
	jdff dff_A_PhUHrHOZ7_0(.dout(w_dff_A_86xheCjg3_0),.din(w_dff_A_PhUHrHOZ7_0),.clk(gclk));
	jdff dff_A_86xheCjg3_0(.dout(w_dff_A_MvYWYMLm1_0),.din(w_dff_A_86xheCjg3_0),.clk(gclk));
	jdff dff_A_MvYWYMLm1_0(.dout(w_dff_A_afGqxUSh5_0),.din(w_dff_A_MvYWYMLm1_0),.clk(gclk));
	jdff dff_A_afGqxUSh5_0(.dout(w_dff_A_29OzCClW3_0),.din(w_dff_A_afGqxUSh5_0),.clk(gclk));
	jdff dff_A_29OzCClW3_0(.dout(w_dff_A_xPfzRuKI6_0),.din(w_dff_A_29OzCClW3_0),.clk(gclk));
	jdff dff_A_xPfzRuKI6_0(.dout(w_dff_A_i3he0eTn3_0),.din(w_dff_A_xPfzRuKI6_0),.clk(gclk));
	jdff dff_A_i3he0eTn3_0(.dout(w_dff_A_FBinRMAB2_0),.din(w_dff_A_i3he0eTn3_0),.clk(gclk));
	jdff dff_A_FBinRMAB2_0(.dout(w_dff_A_s9NQpRPR7_0),.din(w_dff_A_FBinRMAB2_0),.clk(gclk));
	jdff dff_A_s9NQpRPR7_0(.dout(w_dff_A_qsIl0uKV7_0),.din(w_dff_A_s9NQpRPR7_0),.clk(gclk));
	jdff dff_A_qsIl0uKV7_0(.dout(w_dff_A_YAR7DUGh4_0),.din(w_dff_A_qsIl0uKV7_0),.clk(gclk));
	jdff dff_A_YAR7DUGh4_0(.dout(w_dff_A_xnnGLDJX7_0),.din(w_dff_A_YAR7DUGh4_0),.clk(gclk));
	jdff dff_A_xnnGLDJX7_0(.dout(w_dff_A_TuGhBZeR4_0),.din(w_dff_A_xnnGLDJX7_0),.clk(gclk));
	jdff dff_A_TuGhBZeR4_0(.dout(w_dff_A_XmFxiQdh2_0),.din(w_dff_A_TuGhBZeR4_0),.clk(gclk));
	jdff dff_A_XmFxiQdh2_0(.dout(w_dff_A_NVDhUuzE8_0),.din(w_dff_A_XmFxiQdh2_0),.clk(gclk));
	jdff dff_A_NVDhUuzE8_0(.dout(w_dff_A_2FCebLD21_0),.din(w_dff_A_NVDhUuzE8_0),.clk(gclk));
	jdff dff_A_2FCebLD21_0(.dout(w_dff_A_KaQOO7I14_0),.din(w_dff_A_2FCebLD21_0),.clk(gclk));
	jdff dff_A_KaQOO7I14_0(.dout(G639),.din(w_dff_A_KaQOO7I14_0),.clk(gclk));
	jdff dff_A_ws6qj8t84_2(.dout(w_dff_A_015pBpAd3_0),.din(w_dff_A_ws6qj8t84_2),.clk(gclk));
	jdff dff_A_015pBpAd3_0(.dout(w_dff_A_OyNego9h7_0),.din(w_dff_A_015pBpAd3_0),.clk(gclk));
	jdff dff_A_OyNego9h7_0(.dout(w_dff_A_EqMQ4B6w1_0),.din(w_dff_A_OyNego9h7_0),.clk(gclk));
	jdff dff_A_EqMQ4B6w1_0(.dout(w_dff_A_LdP7p3BV4_0),.din(w_dff_A_EqMQ4B6w1_0),.clk(gclk));
	jdff dff_A_LdP7p3BV4_0(.dout(w_dff_A_6oMK9IOl0_0),.din(w_dff_A_LdP7p3BV4_0),.clk(gclk));
	jdff dff_A_6oMK9IOl0_0(.dout(w_dff_A_tjrGxKfB4_0),.din(w_dff_A_6oMK9IOl0_0),.clk(gclk));
	jdff dff_A_tjrGxKfB4_0(.dout(w_dff_A_z2q3Y7aL0_0),.din(w_dff_A_tjrGxKfB4_0),.clk(gclk));
	jdff dff_A_z2q3Y7aL0_0(.dout(w_dff_A_NdQf38A18_0),.din(w_dff_A_z2q3Y7aL0_0),.clk(gclk));
	jdff dff_A_NdQf38A18_0(.dout(w_dff_A_8imp4K072_0),.din(w_dff_A_NdQf38A18_0),.clk(gclk));
	jdff dff_A_8imp4K072_0(.dout(w_dff_A_qQleIalw2_0),.din(w_dff_A_8imp4K072_0),.clk(gclk));
	jdff dff_A_qQleIalw2_0(.dout(w_dff_A_HcjAf0SE6_0),.din(w_dff_A_qQleIalw2_0),.clk(gclk));
	jdff dff_A_HcjAf0SE6_0(.dout(w_dff_A_7YkBhXD80_0),.din(w_dff_A_HcjAf0SE6_0),.clk(gclk));
	jdff dff_A_7YkBhXD80_0(.dout(w_dff_A_3zOfexpy2_0),.din(w_dff_A_7YkBhXD80_0),.clk(gclk));
	jdff dff_A_3zOfexpy2_0(.dout(w_dff_A_jq9AWYos0_0),.din(w_dff_A_3zOfexpy2_0),.clk(gclk));
	jdff dff_A_jq9AWYos0_0(.dout(w_dff_A_icRQlaTT8_0),.din(w_dff_A_jq9AWYos0_0),.clk(gclk));
	jdff dff_A_icRQlaTT8_0(.dout(w_dff_A_T92Cjpfb7_0),.din(w_dff_A_icRQlaTT8_0),.clk(gclk));
	jdff dff_A_T92Cjpfb7_0(.dout(w_dff_A_4gYHMlAg4_0),.din(w_dff_A_T92Cjpfb7_0),.clk(gclk));
	jdff dff_A_4gYHMlAg4_0(.dout(w_dff_A_kbRzr4z37_0),.din(w_dff_A_4gYHMlAg4_0),.clk(gclk));
	jdff dff_A_kbRzr4z37_0(.dout(w_dff_A_w7CZ9g636_0),.din(w_dff_A_kbRzr4z37_0),.clk(gclk));
	jdff dff_A_w7CZ9g636_0(.dout(w_dff_A_WfSr0u5T5_0),.din(w_dff_A_w7CZ9g636_0),.clk(gclk));
	jdff dff_A_WfSr0u5T5_0(.dout(G673),.din(w_dff_A_WfSr0u5T5_0),.clk(gclk));
	jdff dff_A_JaHo8t0x7_2(.dout(w_dff_A_dIzQhL2j5_0),.din(w_dff_A_JaHo8t0x7_2),.clk(gclk));
	jdff dff_A_dIzQhL2j5_0(.dout(w_dff_A_ZvrQpCfx1_0),.din(w_dff_A_dIzQhL2j5_0),.clk(gclk));
	jdff dff_A_ZvrQpCfx1_0(.dout(w_dff_A_V2esmU2Z2_0),.din(w_dff_A_ZvrQpCfx1_0),.clk(gclk));
	jdff dff_A_V2esmU2Z2_0(.dout(w_dff_A_NaYIGfTX9_0),.din(w_dff_A_V2esmU2Z2_0),.clk(gclk));
	jdff dff_A_NaYIGfTX9_0(.dout(w_dff_A_UjMM8cGS7_0),.din(w_dff_A_NaYIGfTX9_0),.clk(gclk));
	jdff dff_A_UjMM8cGS7_0(.dout(w_dff_A_IlGHhJde7_0),.din(w_dff_A_UjMM8cGS7_0),.clk(gclk));
	jdff dff_A_IlGHhJde7_0(.dout(w_dff_A_v6NsRYfv4_0),.din(w_dff_A_IlGHhJde7_0),.clk(gclk));
	jdff dff_A_v6NsRYfv4_0(.dout(w_dff_A_bHbZaIgZ1_0),.din(w_dff_A_v6NsRYfv4_0),.clk(gclk));
	jdff dff_A_bHbZaIgZ1_0(.dout(w_dff_A_lqN2WGM14_0),.din(w_dff_A_bHbZaIgZ1_0),.clk(gclk));
	jdff dff_A_lqN2WGM14_0(.dout(w_dff_A_jyyJPsk94_0),.din(w_dff_A_lqN2WGM14_0),.clk(gclk));
	jdff dff_A_jyyJPsk94_0(.dout(w_dff_A_6wu7qkfH2_0),.din(w_dff_A_jyyJPsk94_0),.clk(gclk));
	jdff dff_A_6wu7qkfH2_0(.dout(w_dff_A_lHcTP5hU3_0),.din(w_dff_A_6wu7qkfH2_0),.clk(gclk));
	jdff dff_A_lHcTP5hU3_0(.dout(w_dff_A_3j7EJt0w8_0),.din(w_dff_A_lHcTP5hU3_0),.clk(gclk));
	jdff dff_A_3j7EJt0w8_0(.dout(w_dff_A_vXu0IyyP8_0),.din(w_dff_A_3j7EJt0w8_0),.clk(gclk));
	jdff dff_A_vXu0IyyP8_0(.dout(w_dff_A_x9rn4HH10_0),.din(w_dff_A_vXu0IyyP8_0),.clk(gclk));
	jdff dff_A_x9rn4HH10_0(.dout(w_dff_A_OOPfshA13_0),.din(w_dff_A_x9rn4HH10_0),.clk(gclk));
	jdff dff_A_OOPfshA13_0(.dout(w_dff_A_XT5aZqsB6_0),.din(w_dff_A_OOPfshA13_0),.clk(gclk));
	jdff dff_A_XT5aZqsB6_0(.dout(w_dff_A_duFMRqfy3_0),.din(w_dff_A_XT5aZqsB6_0),.clk(gclk));
	jdff dff_A_duFMRqfy3_0(.dout(w_dff_A_p7YBxnct8_0),.din(w_dff_A_duFMRqfy3_0),.clk(gclk));
	jdff dff_A_p7YBxnct8_0(.dout(w_dff_A_3zglwhZp4_0),.din(w_dff_A_p7YBxnct8_0),.clk(gclk));
	jdff dff_A_3zglwhZp4_0(.dout(G707),.din(w_dff_A_3zglwhZp4_0),.clk(gclk));
	jdff dff_A_bWD9Wu3L6_2(.dout(w_dff_A_egedGTJ07_0),.din(w_dff_A_bWD9Wu3L6_2),.clk(gclk));
	jdff dff_A_egedGTJ07_0(.dout(w_dff_A_JygkQk1H6_0),.din(w_dff_A_egedGTJ07_0),.clk(gclk));
	jdff dff_A_JygkQk1H6_0(.dout(w_dff_A_Lzy4S0Fj9_0),.din(w_dff_A_JygkQk1H6_0),.clk(gclk));
	jdff dff_A_Lzy4S0Fj9_0(.dout(w_dff_A_n7pbn32l1_0),.din(w_dff_A_Lzy4S0Fj9_0),.clk(gclk));
	jdff dff_A_n7pbn32l1_0(.dout(w_dff_A_C1JZcZK63_0),.din(w_dff_A_n7pbn32l1_0),.clk(gclk));
	jdff dff_A_C1JZcZK63_0(.dout(w_dff_A_Iat9NUY51_0),.din(w_dff_A_C1JZcZK63_0),.clk(gclk));
	jdff dff_A_Iat9NUY51_0(.dout(w_dff_A_N2p1n2bt4_0),.din(w_dff_A_Iat9NUY51_0),.clk(gclk));
	jdff dff_A_N2p1n2bt4_0(.dout(w_dff_A_9TcUCaah0_0),.din(w_dff_A_N2p1n2bt4_0),.clk(gclk));
	jdff dff_A_9TcUCaah0_0(.dout(w_dff_A_JvxMqBwD5_0),.din(w_dff_A_9TcUCaah0_0),.clk(gclk));
	jdff dff_A_JvxMqBwD5_0(.dout(w_dff_A_RGvKg6k77_0),.din(w_dff_A_JvxMqBwD5_0),.clk(gclk));
	jdff dff_A_RGvKg6k77_0(.dout(w_dff_A_onUMk9qV1_0),.din(w_dff_A_RGvKg6k77_0),.clk(gclk));
	jdff dff_A_onUMk9qV1_0(.dout(w_dff_A_sXd9QkmX8_0),.din(w_dff_A_onUMk9qV1_0),.clk(gclk));
	jdff dff_A_sXd9QkmX8_0(.dout(w_dff_A_G2JjN1e75_0),.din(w_dff_A_sXd9QkmX8_0),.clk(gclk));
	jdff dff_A_G2JjN1e75_0(.dout(w_dff_A_YNuWrXEO2_0),.din(w_dff_A_G2JjN1e75_0),.clk(gclk));
	jdff dff_A_YNuWrXEO2_0(.dout(w_dff_A_qKhKx99B7_0),.din(w_dff_A_YNuWrXEO2_0),.clk(gclk));
	jdff dff_A_qKhKx99B7_0(.dout(w_dff_A_YrSPJqTx1_0),.din(w_dff_A_qKhKx99B7_0),.clk(gclk));
	jdff dff_A_YrSPJqTx1_0(.dout(w_dff_A_ON6UoYrD8_0),.din(w_dff_A_YrSPJqTx1_0),.clk(gclk));
	jdff dff_A_ON6UoYrD8_0(.dout(w_dff_A_BIfRkML18_0),.din(w_dff_A_ON6UoYrD8_0),.clk(gclk));
	jdff dff_A_BIfRkML18_0(.dout(w_dff_A_UrCQuzzc8_0),.din(w_dff_A_BIfRkML18_0),.clk(gclk));
	jdff dff_A_UrCQuzzc8_0(.dout(w_dff_A_hqxELb3E2_0),.din(w_dff_A_UrCQuzzc8_0),.clk(gclk));
	jdff dff_A_hqxELb3E2_0(.dout(G715),.din(w_dff_A_hqxELb3E2_0),.clk(gclk));
	jdff dff_A_xzIOgP9N0_2(.dout(w_dff_A_qtp2Zvl69_0),.din(w_dff_A_xzIOgP9N0_2),.clk(gclk));
	jdff dff_A_qtp2Zvl69_0(.dout(w_dff_A_tcxHJBT64_0),.din(w_dff_A_qtp2Zvl69_0),.clk(gclk));
	jdff dff_A_tcxHJBT64_0(.dout(w_dff_A_fTmQci600_0),.din(w_dff_A_tcxHJBT64_0),.clk(gclk));
	jdff dff_A_fTmQci600_0(.dout(w_dff_A_zp8MIT2P7_0),.din(w_dff_A_fTmQci600_0),.clk(gclk));
	jdff dff_A_zp8MIT2P7_0(.dout(w_dff_A_NkCSW3o55_0),.din(w_dff_A_zp8MIT2P7_0),.clk(gclk));
	jdff dff_A_NkCSW3o55_0(.dout(w_dff_A_5z7rmwx18_0),.din(w_dff_A_NkCSW3o55_0),.clk(gclk));
	jdff dff_A_5z7rmwx18_0(.dout(w_dff_A_ryEFsn1F1_0),.din(w_dff_A_5z7rmwx18_0),.clk(gclk));
	jdff dff_A_ryEFsn1F1_0(.dout(w_dff_A_TOGoBy9I1_0),.din(w_dff_A_ryEFsn1F1_0),.clk(gclk));
	jdff dff_A_TOGoBy9I1_0(.dout(w_dff_A_4FNNIWn95_0),.din(w_dff_A_TOGoBy9I1_0),.clk(gclk));
	jdff dff_A_4FNNIWn95_0(.dout(w_dff_A_cxr9omFl3_0),.din(w_dff_A_4FNNIWn95_0),.clk(gclk));
	jdff dff_A_cxr9omFl3_0(.dout(w_dff_A_EPombFkj9_0),.din(w_dff_A_cxr9omFl3_0),.clk(gclk));
	jdff dff_A_EPombFkj9_0(.dout(w_dff_A_nbJAbxhj8_0),.din(w_dff_A_EPombFkj9_0),.clk(gclk));
	jdff dff_A_nbJAbxhj8_0(.dout(w_dff_A_KwAFMWfm1_0),.din(w_dff_A_nbJAbxhj8_0),.clk(gclk));
	jdff dff_A_KwAFMWfm1_0(.dout(w_dff_A_vZP2OyaB3_0),.din(w_dff_A_KwAFMWfm1_0),.clk(gclk));
	jdff dff_A_vZP2OyaB3_0(.dout(w_dff_A_n81M39BH6_0),.din(w_dff_A_vZP2OyaB3_0),.clk(gclk));
	jdff dff_A_n81M39BH6_0(.dout(w_dff_A_nfvfRpeA3_0),.din(w_dff_A_n81M39BH6_0),.clk(gclk));
	jdff dff_A_nfvfRpeA3_0(.dout(G598),.din(w_dff_A_nfvfRpeA3_0),.clk(gclk));
	jdff dff_A_zRJ957kz3_2(.dout(w_dff_A_eJFULSEg9_0),.din(w_dff_A_zRJ957kz3_2),.clk(gclk));
	jdff dff_A_eJFULSEg9_0(.dout(w_dff_A_sf6JQtNE6_0),.din(w_dff_A_eJFULSEg9_0),.clk(gclk));
	jdff dff_A_sf6JQtNE6_0(.dout(w_dff_A_y9QQgcGv4_0),.din(w_dff_A_sf6JQtNE6_0),.clk(gclk));
	jdff dff_A_y9QQgcGv4_0(.dout(w_dff_A_KxERmOrj0_0),.din(w_dff_A_y9QQgcGv4_0),.clk(gclk));
	jdff dff_A_KxERmOrj0_0(.dout(w_dff_A_ZQ6MBruf4_0),.din(w_dff_A_KxERmOrj0_0),.clk(gclk));
	jdff dff_A_ZQ6MBruf4_0(.dout(w_dff_A_ljvutjJj6_0),.din(w_dff_A_ZQ6MBruf4_0),.clk(gclk));
	jdff dff_A_ljvutjJj6_0(.dout(w_dff_A_rFhpsRjl1_0),.din(w_dff_A_ljvutjJj6_0),.clk(gclk));
	jdff dff_A_rFhpsRjl1_0(.dout(w_dff_A_qbzp1b9S9_0),.din(w_dff_A_rFhpsRjl1_0),.clk(gclk));
	jdff dff_A_qbzp1b9S9_0(.dout(w_dff_A_pPTsB0Vw1_0),.din(w_dff_A_qbzp1b9S9_0),.clk(gclk));
	jdff dff_A_pPTsB0Vw1_0(.dout(w_dff_A_xBHpKUf87_0),.din(w_dff_A_pPTsB0Vw1_0),.clk(gclk));
	jdff dff_A_xBHpKUf87_0(.dout(w_dff_A_7yyuQvP80_0),.din(w_dff_A_xBHpKUf87_0),.clk(gclk));
	jdff dff_A_7yyuQvP80_0(.dout(w_dff_A_qQ24Hh9Q0_0),.din(w_dff_A_7yyuQvP80_0),.clk(gclk));
	jdff dff_A_qQ24Hh9Q0_0(.dout(w_dff_A_OXYQVFwB5_0),.din(w_dff_A_qQ24Hh9Q0_0),.clk(gclk));
	jdff dff_A_OXYQVFwB5_0(.dout(w_dff_A_Tx7pZEYF5_0),.din(w_dff_A_OXYQVFwB5_0),.clk(gclk));
	jdff dff_A_Tx7pZEYF5_0(.dout(w_dff_A_XXE4mgvB2_0),.din(w_dff_A_Tx7pZEYF5_0),.clk(gclk));
	jdff dff_A_XXE4mgvB2_0(.dout(w_dff_A_3OQY6HDV2_0),.din(w_dff_A_XXE4mgvB2_0),.clk(gclk));
	jdff dff_A_3OQY6HDV2_0(.dout(G610),.din(w_dff_A_3OQY6HDV2_0),.clk(gclk));
	jdff dff_A_hKGz8qj65_2(.dout(w_dff_A_j6UBRRzF3_0),.din(w_dff_A_hKGz8qj65_2),.clk(gclk));
	jdff dff_A_j6UBRRzF3_0(.dout(w_dff_A_wkuCNJ3M2_0),.din(w_dff_A_j6UBRRzF3_0),.clk(gclk));
	jdff dff_A_wkuCNJ3M2_0(.dout(w_dff_A_NARCoohC0_0),.din(w_dff_A_wkuCNJ3M2_0),.clk(gclk));
	jdff dff_A_NARCoohC0_0(.dout(w_dff_A_zyEip4tR0_0),.din(w_dff_A_NARCoohC0_0),.clk(gclk));
	jdff dff_A_zyEip4tR0_0(.dout(w_dff_A_FPzSBU0J1_0),.din(w_dff_A_zyEip4tR0_0),.clk(gclk));
	jdff dff_A_FPzSBU0J1_0(.dout(w_dff_A_C87JJzYi4_0),.din(w_dff_A_FPzSBU0J1_0),.clk(gclk));
	jdff dff_A_C87JJzYi4_0(.dout(w_dff_A_NPoU0ZkM2_0),.din(w_dff_A_C87JJzYi4_0),.clk(gclk));
	jdff dff_A_NPoU0ZkM2_0(.dout(w_dff_A_6R3G86rj1_0),.din(w_dff_A_NPoU0ZkM2_0),.clk(gclk));
	jdff dff_A_6R3G86rj1_0(.dout(w_dff_A_3ItQFBkA7_0),.din(w_dff_A_6R3G86rj1_0),.clk(gclk));
	jdff dff_A_3ItQFBkA7_0(.dout(w_dff_A_GsfTw6EV4_0),.din(w_dff_A_3ItQFBkA7_0),.clk(gclk));
	jdff dff_A_GsfTw6EV4_0(.dout(w_dff_A_LoKY0wd96_0),.din(w_dff_A_GsfTw6EV4_0),.clk(gclk));
	jdff dff_A_LoKY0wd96_0(.dout(w_dff_A_c3XjQSlA5_0),.din(w_dff_A_LoKY0wd96_0),.clk(gclk));
	jdff dff_A_c3XjQSlA5_0(.dout(w_dff_A_PZkWU55K1_0),.din(w_dff_A_c3XjQSlA5_0),.clk(gclk));
	jdff dff_A_PZkWU55K1_0(.dout(w_dff_A_bIRRAvyk5_0),.din(w_dff_A_PZkWU55K1_0),.clk(gclk));
	jdff dff_A_bIRRAvyk5_0(.dout(G588),.din(w_dff_A_bIRRAvyk5_0),.clk(gclk));
	jdff dff_A_CvoF0cw43_2(.dout(w_dff_A_DnFb1OsR6_0),.din(w_dff_A_CvoF0cw43_2),.clk(gclk));
	jdff dff_A_DnFb1OsR6_0(.dout(w_dff_A_ropaRYC16_0),.din(w_dff_A_DnFb1OsR6_0),.clk(gclk));
	jdff dff_A_ropaRYC16_0(.dout(w_dff_A_zx6cagAZ3_0),.din(w_dff_A_ropaRYC16_0),.clk(gclk));
	jdff dff_A_zx6cagAZ3_0(.dout(w_dff_A_mnxyhXD91_0),.din(w_dff_A_zx6cagAZ3_0),.clk(gclk));
	jdff dff_A_mnxyhXD91_0(.dout(w_dff_A_sOroxrfW4_0),.din(w_dff_A_mnxyhXD91_0),.clk(gclk));
	jdff dff_A_sOroxrfW4_0(.dout(w_dff_A_W8JoGkbB8_0),.din(w_dff_A_sOroxrfW4_0),.clk(gclk));
	jdff dff_A_W8JoGkbB8_0(.dout(w_dff_A_Erdnakmx7_0),.din(w_dff_A_W8JoGkbB8_0),.clk(gclk));
	jdff dff_A_Erdnakmx7_0(.dout(w_dff_A_fPdeymrQ6_0),.din(w_dff_A_Erdnakmx7_0),.clk(gclk));
	jdff dff_A_fPdeymrQ6_0(.dout(w_dff_A_9tuJvtRw3_0),.din(w_dff_A_fPdeymrQ6_0),.clk(gclk));
	jdff dff_A_9tuJvtRw3_0(.dout(w_dff_A_8la4g7xV9_0),.din(w_dff_A_9tuJvtRw3_0),.clk(gclk));
	jdff dff_A_8la4g7xV9_0(.dout(w_dff_A_38uRb4FB7_0),.din(w_dff_A_8la4g7xV9_0),.clk(gclk));
	jdff dff_A_38uRb4FB7_0(.dout(w_dff_A_iTXTnXOr7_0),.din(w_dff_A_38uRb4FB7_0),.clk(gclk));
	jdff dff_A_iTXTnXOr7_0(.dout(w_dff_A_pRS8QfrQ9_0),.din(w_dff_A_iTXTnXOr7_0),.clk(gclk));
	jdff dff_A_pRS8QfrQ9_0(.dout(w_dff_A_RrFlHIi41_0),.din(w_dff_A_pRS8QfrQ9_0),.clk(gclk));
	jdff dff_A_RrFlHIi41_0(.dout(w_dff_A_XN60dkC87_0),.din(w_dff_A_RrFlHIi41_0),.clk(gclk));
	jdff dff_A_XN60dkC87_0(.dout(w_dff_A_Sz51mRe62_0),.din(w_dff_A_XN60dkC87_0),.clk(gclk));
	jdff dff_A_Sz51mRe62_0(.dout(G615),.din(w_dff_A_Sz51mRe62_0),.clk(gclk));
	jdff dff_A_VtM4hs6P0_2(.dout(w_dff_A_3zCBu4vo4_0),.din(w_dff_A_VtM4hs6P0_2),.clk(gclk));
	jdff dff_A_3zCBu4vo4_0(.dout(w_dff_A_TPdnABiS4_0),.din(w_dff_A_3zCBu4vo4_0),.clk(gclk));
	jdff dff_A_TPdnABiS4_0(.dout(w_dff_A_By7JXafK2_0),.din(w_dff_A_TPdnABiS4_0),.clk(gclk));
	jdff dff_A_By7JXafK2_0(.dout(w_dff_A_plpcEgRW6_0),.din(w_dff_A_By7JXafK2_0),.clk(gclk));
	jdff dff_A_plpcEgRW6_0(.dout(w_dff_A_12BWs4LY1_0),.din(w_dff_A_plpcEgRW6_0),.clk(gclk));
	jdff dff_A_12BWs4LY1_0(.dout(w_dff_A_capNGH7F3_0),.din(w_dff_A_12BWs4LY1_0),.clk(gclk));
	jdff dff_A_capNGH7F3_0(.dout(w_dff_A_qTvV0HAi9_0),.din(w_dff_A_capNGH7F3_0),.clk(gclk));
	jdff dff_A_qTvV0HAi9_0(.dout(w_dff_A_TbGJumbf8_0),.din(w_dff_A_qTvV0HAi9_0),.clk(gclk));
	jdff dff_A_TbGJumbf8_0(.dout(w_dff_A_evBqJTV83_0),.din(w_dff_A_TbGJumbf8_0),.clk(gclk));
	jdff dff_A_evBqJTV83_0(.dout(w_dff_A_pkH8XC9j1_0),.din(w_dff_A_evBqJTV83_0),.clk(gclk));
	jdff dff_A_pkH8XC9j1_0(.dout(w_dff_A_OcIZUuSL6_0),.din(w_dff_A_pkH8XC9j1_0),.clk(gclk));
	jdff dff_A_OcIZUuSL6_0(.dout(w_dff_A_81D5i6Vu8_0),.din(w_dff_A_OcIZUuSL6_0),.clk(gclk));
	jdff dff_A_81D5i6Vu8_0(.dout(w_dff_A_oWJNu1ep4_0),.din(w_dff_A_81D5i6Vu8_0),.clk(gclk));
	jdff dff_A_oWJNu1ep4_0(.dout(w_dff_A_5CkQLVEd2_0),.din(w_dff_A_oWJNu1ep4_0),.clk(gclk));
	jdff dff_A_5CkQLVEd2_0(.dout(w_dff_A_3g0Gxo518_0),.din(w_dff_A_5CkQLVEd2_0),.clk(gclk));
	jdff dff_A_3g0Gxo518_0(.dout(w_dff_A_yBeqkK3y9_0),.din(w_dff_A_3g0Gxo518_0),.clk(gclk));
	jdff dff_A_yBeqkK3y9_0(.dout(G626),.din(w_dff_A_yBeqkK3y9_0),.clk(gclk));
	jdff dff_A_tughExAl8_2(.dout(w_dff_A_ffPO6mIn1_0),.din(w_dff_A_tughExAl8_2),.clk(gclk));
	jdff dff_A_ffPO6mIn1_0(.dout(w_dff_A_czdf2fEN5_0),.din(w_dff_A_ffPO6mIn1_0),.clk(gclk));
	jdff dff_A_czdf2fEN5_0(.dout(w_dff_A_l7WpYvAV6_0),.din(w_dff_A_czdf2fEN5_0),.clk(gclk));
	jdff dff_A_l7WpYvAV6_0(.dout(w_dff_A_YVKVgraS4_0),.din(w_dff_A_l7WpYvAV6_0),.clk(gclk));
	jdff dff_A_YVKVgraS4_0(.dout(w_dff_A_Hczlb0RS4_0),.din(w_dff_A_YVKVgraS4_0),.clk(gclk));
	jdff dff_A_Hczlb0RS4_0(.dout(w_dff_A_4lOsBLii7_0),.din(w_dff_A_Hczlb0RS4_0),.clk(gclk));
	jdff dff_A_4lOsBLii7_0(.dout(w_dff_A_EEjO3bnx3_0),.din(w_dff_A_4lOsBLii7_0),.clk(gclk));
	jdff dff_A_EEjO3bnx3_0(.dout(w_dff_A_VMSzwsEh6_0),.din(w_dff_A_EEjO3bnx3_0),.clk(gclk));
	jdff dff_A_VMSzwsEh6_0(.dout(w_dff_A_onJo3shw3_0),.din(w_dff_A_VMSzwsEh6_0),.clk(gclk));
	jdff dff_A_onJo3shw3_0(.dout(w_dff_A_1vlwOEM77_0),.din(w_dff_A_onJo3shw3_0),.clk(gclk));
	jdff dff_A_1vlwOEM77_0(.dout(w_dff_A_eWvLJsfQ7_0),.din(w_dff_A_1vlwOEM77_0),.clk(gclk));
	jdff dff_A_eWvLJsfQ7_0(.dout(w_dff_A_2nzI1wQl5_0),.din(w_dff_A_eWvLJsfQ7_0),.clk(gclk));
	jdff dff_A_2nzI1wQl5_0(.dout(w_dff_A_ra7phtSO1_0),.din(w_dff_A_2nzI1wQl5_0),.clk(gclk));
	jdff dff_A_ra7phtSO1_0(.dout(w_dff_A_qJuZHddv4_0),.din(w_dff_A_ra7phtSO1_0),.clk(gclk));
	jdff dff_A_qJuZHddv4_0(.dout(G632),.din(w_dff_A_qJuZHddv4_0),.clk(gclk));
	jdff dff_A_gwSMvLaq9_1(.dout(w_dff_A_40XfPXOS1_0),.din(w_dff_A_gwSMvLaq9_1),.clk(gclk));
	jdff dff_A_40XfPXOS1_0(.dout(w_dff_A_jgLQuiM91_0),.din(w_dff_A_40XfPXOS1_0),.clk(gclk));
	jdff dff_A_jgLQuiM91_0(.dout(w_dff_A_h6R6veJV8_0),.din(w_dff_A_jgLQuiM91_0),.clk(gclk));
	jdff dff_A_h6R6veJV8_0(.dout(w_dff_A_8bO67LWI0_0),.din(w_dff_A_h6R6veJV8_0),.clk(gclk));
	jdff dff_A_8bO67LWI0_0(.dout(w_dff_A_JMNeqgL47_0),.din(w_dff_A_8bO67LWI0_0),.clk(gclk));
	jdff dff_A_JMNeqgL47_0(.dout(w_dff_A_YQK5lujo8_0),.din(w_dff_A_JMNeqgL47_0),.clk(gclk));
	jdff dff_A_YQK5lujo8_0(.dout(w_dff_A_ZTU1AUDK6_0),.din(w_dff_A_YQK5lujo8_0),.clk(gclk));
	jdff dff_A_ZTU1AUDK6_0(.dout(w_dff_A_h3ptnhXD5_0),.din(w_dff_A_ZTU1AUDK6_0),.clk(gclk));
	jdff dff_A_h3ptnhXD5_0(.dout(w_dff_A_eva45roY5_0),.din(w_dff_A_h3ptnhXD5_0),.clk(gclk));
	jdff dff_A_eva45roY5_0(.dout(w_dff_A_zWGAw06Y1_0),.din(w_dff_A_eva45roY5_0),.clk(gclk));
	jdff dff_A_zWGAw06Y1_0(.dout(w_dff_A_3C5ScsxO7_0),.din(w_dff_A_zWGAw06Y1_0),.clk(gclk));
	jdff dff_A_3C5ScsxO7_0(.dout(w_dff_A_W1Lie4tp9_0),.din(w_dff_A_3C5ScsxO7_0),.clk(gclk));
	jdff dff_A_W1Lie4tp9_0(.dout(w_dff_A_7FKntTBz6_0),.din(w_dff_A_W1Lie4tp9_0),.clk(gclk));
	jdff dff_A_7FKntTBz6_0(.dout(w_dff_A_t8OrPUSl5_0),.din(w_dff_A_7FKntTBz6_0),.clk(gclk));
	jdff dff_A_t8OrPUSl5_0(.dout(w_dff_A_XNeGWqrB2_0),.din(w_dff_A_t8OrPUSl5_0),.clk(gclk));
	jdff dff_A_XNeGWqrB2_0(.dout(w_dff_A_drHtD34t4_0),.din(w_dff_A_XNeGWqrB2_0),.clk(gclk));
	jdff dff_A_drHtD34t4_0(.dout(w_dff_A_LBgFRq4P6_0),.din(w_dff_A_drHtD34t4_0),.clk(gclk));
	jdff dff_A_LBgFRq4P6_0(.dout(w_dff_A_40x3LFmT8_0),.din(w_dff_A_LBgFRq4P6_0),.clk(gclk));
	jdff dff_A_40x3LFmT8_0(.dout(w_dff_A_TRxscYJQ9_0),.din(w_dff_A_40x3LFmT8_0),.clk(gclk));
	jdff dff_A_TRxscYJQ9_0(.dout(w_dff_A_FQB1xfgN4_0),.din(w_dff_A_TRxscYJQ9_0),.clk(gclk));
	jdff dff_A_FQB1xfgN4_0(.dout(G1002),.din(w_dff_A_FQB1xfgN4_0),.clk(gclk));
	jdff dff_A_ByIlIlBF7_1(.dout(w_dff_A_1fjAoNQt7_0),.din(w_dff_A_ByIlIlBF7_1),.clk(gclk));
	jdff dff_A_1fjAoNQt7_0(.dout(w_dff_A_yXhwmdtn3_0),.din(w_dff_A_1fjAoNQt7_0),.clk(gclk));
	jdff dff_A_yXhwmdtn3_0(.dout(w_dff_A_Deg2164w2_0),.din(w_dff_A_yXhwmdtn3_0),.clk(gclk));
	jdff dff_A_Deg2164w2_0(.dout(w_dff_A_noa6RaVy0_0),.din(w_dff_A_Deg2164w2_0),.clk(gclk));
	jdff dff_A_noa6RaVy0_0(.dout(w_dff_A_DQG24vuE2_0),.din(w_dff_A_noa6RaVy0_0),.clk(gclk));
	jdff dff_A_DQG24vuE2_0(.dout(w_dff_A_d1i08bp22_0),.din(w_dff_A_DQG24vuE2_0),.clk(gclk));
	jdff dff_A_d1i08bp22_0(.dout(w_dff_A_izEHIz1J5_0),.din(w_dff_A_d1i08bp22_0),.clk(gclk));
	jdff dff_A_izEHIz1J5_0(.dout(w_dff_A_RCgnpovW7_0),.din(w_dff_A_izEHIz1J5_0),.clk(gclk));
	jdff dff_A_RCgnpovW7_0(.dout(w_dff_A_nn7kXtBx3_0),.din(w_dff_A_RCgnpovW7_0),.clk(gclk));
	jdff dff_A_nn7kXtBx3_0(.dout(w_dff_A_kzNCJH836_0),.din(w_dff_A_nn7kXtBx3_0),.clk(gclk));
	jdff dff_A_kzNCJH836_0(.dout(w_dff_A_lmWg2PGX7_0),.din(w_dff_A_kzNCJH836_0),.clk(gclk));
	jdff dff_A_lmWg2PGX7_0(.dout(w_dff_A_Ek1LmCHy2_0),.din(w_dff_A_lmWg2PGX7_0),.clk(gclk));
	jdff dff_A_Ek1LmCHy2_0(.dout(w_dff_A_cUWurIMW4_0),.din(w_dff_A_Ek1LmCHy2_0),.clk(gclk));
	jdff dff_A_cUWurIMW4_0(.dout(w_dff_A_kfCCRjIW9_0),.din(w_dff_A_cUWurIMW4_0),.clk(gclk));
	jdff dff_A_kfCCRjIW9_0(.dout(w_dff_A_1Y1BBiEM8_0),.din(w_dff_A_kfCCRjIW9_0),.clk(gclk));
	jdff dff_A_1Y1BBiEM8_0(.dout(w_dff_A_Dn8KA3kl9_0),.din(w_dff_A_1Y1BBiEM8_0),.clk(gclk));
	jdff dff_A_Dn8KA3kl9_0(.dout(w_dff_A_779Jtbhz6_0),.din(w_dff_A_Dn8KA3kl9_0),.clk(gclk));
	jdff dff_A_779Jtbhz6_0(.dout(w_dff_A_Jr3op34A3_0),.din(w_dff_A_779Jtbhz6_0),.clk(gclk));
	jdff dff_A_Jr3op34A3_0(.dout(w_dff_A_1TSZgapw6_0),.din(w_dff_A_Jr3op34A3_0),.clk(gclk));
	jdff dff_A_1TSZgapw6_0(.dout(w_dff_A_EPZ5jgC17_0),.din(w_dff_A_1TSZgapw6_0),.clk(gclk));
	jdff dff_A_EPZ5jgC17_0(.dout(G1004),.din(w_dff_A_EPZ5jgC17_0),.clk(gclk));
	jdff dff_A_svarlViU6_2(.dout(w_dff_A_CgGqpF836_0),.din(w_dff_A_svarlViU6_2),.clk(gclk));
	jdff dff_A_CgGqpF836_0(.dout(w_dff_A_NMg4pjqI3_0),.din(w_dff_A_CgGqpF836_0),.clk(gclk));
	jdff dff_A_NMg4pjqI3_0(.dout(w_dff_A_6yfJuldK0_0),.din(w_dff_A_NMg4pjqI3_0),.clk(gclk));
	jdff dff_A_6yfJuldK0_0(.dout(w_dff_A_PV4zbMzR9_0),.din(w_dff_A_6yfJuldK0_0),.clk(gclk));
	jdff dff_A_PV4zbMzR9_0(.dout(w_dff_A_RIoTzfc38_0),.din(w_dff_A_PV4zbMzR9_0),.clk(gclk));
	jdff dff_A_RIoTzfc38_0(.dout(w_dff_A_waHd4PJK8_0),.din(w_dff_A_RIoTzfc38_0),.clk(gclk));
	jdff dff_A_waHd4PJK8_0(.dout(w_dff_A_dcll5poU7_0),.din(w_dff_A_waHd4PJK8_0),.clk(gclk));
	jdff dff_A_dcll5poU7_0(.dout(w_dff_A_BUpZESyO3_0),.din(w_dff_A_dcll5poU7_0),.clk(gclk));
	jdff dff_A_BUpZESyO3_0(.dout(w_dff_A_R79aHdUu8_0),.din(w_dff_A_BUpZESyO3_0),.clk(gclk));
	jdff dff_A_R79aHdUu8_0(.dout(w_dff_A_WcT5831S3_0),.din(w_dff_A_R79aHdUu8_0),.clk(gclk));
	jdff dff_A_WcT5831S3_0(.dout(w_dff_A_VbhswlOh8_0),.din(w_dff_A_WcT5831S3_0),.clk(gclk));
	jdff dff_A_VbhswlOh8_0(.dout(G591),.din(w_dff_A_VbhswlOh8_0),.clk(gclk));
	jdff dff_A_RURQqRW80_2(.dout(w_dff_A_gaijMJHj4_0),.din(w_dff_A_RURQqRW80_2),.clk(gclk));
	jdff dff_A_gaijMJHj4_0(.dout(w_dff_A_EOaFZLwC3_0),.din(w_dff_A_gaijMJHj4_0),.clk(gclk));
	jdff dff_A_EOaFZLwC3_0(.dout(w_dff_A_kZDFzEJi7_0),.din(w_dff_A_EOaFZLwC3_0),.clk(gclk));
	jdff dff_A_kZDFzEJi7_0(.dout(w_dff_A_G2tpAyLK6_0),.din(w_dff_A_kZDFzEJi7_0),.clk(gclk));
	jdff dff_A_G2tpAyLK6_0(.dout(w_dff_A_YUh8VSiC0_0),.din(w_dff_A_G2tpAyLK6_0),.clk(gclk));
	jdff dff_A_YUh8VSiC0_0(.dout(w_dff_A_sxFqwfWM4_0),.din(w_dff_A_YUh8VSiC0_0),.clk(gclk));
	jdff dff_A_sxFqwfWM4_0(.dout(w_dff_A_48QXFV8i3_0),.din(w_dff_A_sxFqwfWM4_0),.clk(gclk));
	jdff dff_A_48QXFV8i3_0(.dout(w_dff_A_n1RyJHH69_0),.din(w_dff_A_48QXFV8i3_0),.clk(gclk));
	jdff dff_A_n1RyJHH69_0(.dout(w_dff_A_gNYiTFhq3_0),.din(w_dff_A_n1RyJHH69_0),.clk(gclk));
	jdff dff_A_gNYiTFhq3_0(.dout(w_dff_A_wUMRnsvn6_0),.din(w_dff_A_gNYiTFhq3_0),.clk(gclk));
	jdff dff_A_wUMRnsvn6_0(.dout(w_dff_A_hMXyVOhu2_0),.din(w_dff_A_wUMRnsvn6_0),.clk(gclk));
	jdff dff_A_hMXyVOhu2_0(.dout(G618),.din(w_dff_A_hMXyVOhu2_0),.clk(gclk));
	jdff dff_A_xNiLG5rl1_2(.dout(w_dff_A_eLEZesFI3_0),.din(w_dff_A_xNiLG5rl1_2),.clk(gclk));
	jdff dff_A_eLEZesFI3_0(.dout(w_dff_A_fX2CMInd4_0),.din(w_dff_A_eLEZesFI3_0),.clk(gclk));
	jdff dff_A_fX2CMInd4_0(.dout(w_dff_A_YXwtDJSN6_0),.din(w_dff_A_fX2CMInd4_0),.clk(gclk));
	jdff dff_A_YXwtDJSN6_0(.dout(w_dff_A_OJCfiZg33_0),.din(w_dff_A_YXwtDJSN6_0),.clk(gclk));
	jdff dff_A_OJCfiZg33_0(.dout(w_dff_A_ljoRMatz8_0),.din(w_dff_A_OJCfiZg33_0),.clk(gclk));
	jdff dff_A_ljoRMatz8_0(.dout(w_dff_A_uZNefROj7_0),.din(w_dff_A_ljoRMatz8_0),.clk(gclk));
	jdff dff_A_uZNefROj7_0(.dout(w_dff_A_D6VtxZDf1_0),.din(w_dff_A_uZNefROj7_0),.clk(gclk));
	jdff dff_A_D6VtxZDf1_0(.dout(w_dff_A_30YzxlNw4_0),.din(w_dff_A_D6VtxZDf1_0),.clk(gclk));
	jdff dff_A_30YzxlNw4_0(.dout(w_dff_A_mWntxtlV6_0),.din(w_dff_A_30YzxlNw4_0),.clk(gclk));
	jdff dff_A_mWntxtlV6_0(.dout(w_dff_A_2yVoIHCO8_0),.din(w_dff_A_mWntxtlV6_0),.clk(gclk));
	jdff dff_A_2yVoIHCO8_0(.dout(w_dff_A_GU3Y6RPS4_0),.din(w_dff_A_2yVoIHCO8_0),.clk(gclk));
	jdff dff_A_GU3Y6RPS4_0(.dout(G621),.din(w_dff_A_GU3Y6RPS4_0),.clk(gclk));
	jdff dff_A_ePXT8ufG1_2(.dout(w_dff_A_z0Jec8un6_0),.din(w_dff_A_ePXT8ufG1_2),.clk(gclk));
	jdff dff_A_z0Jec8un6_0(.dout(w_dff_A_8QYV5llE3_0),.din(w_dff_A_z0Jec8un6_0),.clk(gclk));
	jdff dff_A_8QYV5llE3_0(.dout(w_dff_A_SqtgFKu97_0),.din(w_dff_A_8QYV5llE3_0),.clk(gclk));
	jdff dff_A_SqtgFKu97_0(.dout(w_dff_A_GVGw5AXK7_0),.din(w_dff_A_SqtgFKu97_0),.clk(gclk));
	jdff dff_A_GVGw5AXK7_0(.dout(w_dff_A_HBLn7Tfs9_0),.din(w_dff_A_GVGw5AXK7_0),.clk(gclk));
	jdff dff_A_HBLn7Tfs9_0(.dout(w_dff_A_B0zSvSYp4_0),.din(w_dff_A_HBLn7Tfs9_0),.clk(gclk));
	jdff dff_A_B0zSvSYp4_0(.dout(w_dff_A_BcDV8OsJ0_0),.din(w_dff_A_B0zSvSYp4_0),.clk(gclk));
	jdff dff_A_BcDV8OsJ0_0(.dout(w_dff_A_GRimIAkU9_0),.din(w_dff_A_BcDV8OsJ0_0),.clk(gclk));
	jdff dff_A_GRimIAkU9_0(.dout(w_dff_A_srliIiHF8_0),.din(w_dff_A_GRimIAkU9_0),.clk(gclk));
	jdff dff_A_srliIiHF8_0(.dout(w_dff_A_KCNV2Rsn3_0),.din(w_dff_A_srliIiHF8_0),.clk(gclk));
	jdff dff_A_KCNV2Rsn3_0(.dout(w_dff_A_3jyohAHz4_0),.din(w_dff_A_KCNV2Rsn3_0),.clk(gclk));
	jdff dff_A_3jyohAHz4_0(.dout(G629),.din(w_dff_A_3jyohAHz4_0),.clk(gclk));
	jdff dff_A_RYzzMdAy5_1(.dout(w_dff_A_FTpbQIZu1_0),.din(w_dff_A_RYzzMdAy5_1),.clk(gclk));
	jdff dff_A_FTpbQIZu1_0(.dout(w_dff_A_g6uo8kvg5_0),.din(w_dff_A_FTpbQIZu1_0),.clk(gclk));
	jdff dff_A_g6uo8kvg5_0(.dout(w_dff_A_VIJkmWqd7_0),.din(w_dff_A_g6uo8kvg5_0),.clk(gclk));
	jdff dff_A_VIJkmWqd7_0(.dout(w_dff_A_6TS5PpXV2_0),.din(w_dff_A_VIJkmWqd7_0),.clk(gclk));
	jdff dff_A_6TS5PpXV2_0(.dout(w_dff_A_gd5GNGdK7_0),.din(w_dff_A_6TS5PpXV2_0),.clk(gclk));
	jdff dff_A_gd5GNGdK7_0(.dout(w_dff_A_DNLsY7me4_0),.din(w_dff_A_gd5GNGdK7_0),.clk(gclk));
	jdff dff_A_DNLsY7me4_0(.dout(w_dff_A_DDZHHVvW1_0),.din(w_dff_A_DNLsY7me4_0),.clk(gclk));
	jdff dff_A_DDZHHVvW1_0(.dout(w_dff_A_AWAQaOAL0_0),.din(w_dff_A_DDZHHVvW1_0),.clk(gclk));
	jdff dff_A_AWAQaOAL0_0(.dout(w_dff_A_jzN1owR77_0),.din(w_dff_A_AWAQaOAL0_0),.clk(gclk));
	jdff dff_A_jzN1owR77_0(.dout(w_dff_A_NLwQEubE8_0),.din(w_dff_A_jzN1owR77_0),.clk(gclk));
	jdff dff_A_NLwQEubE8_0(.dout(w_dff_A_g6X9JLKu1_0),.din(w_dff_A_NLwQEubE8_0),.clk(gclk));
	jdff dff_A_g6X9JLKu1_0(.dout(w_dff_A_wyNgCw4k0_0),.din(w_dff_A_g6X9JLKu1_0),.clk(gclk));
	jdff dff_A_wyNgCw4k0_0(.dout(w_dff_A_iYCXIxq65_0),.din(w_dff_A_wyNgCw4k0_0),.clk(gclk));
	jdff dff_A_iYCXIxq65_0(.dout(w_dff_A_3XKw3vF77_0),.din(w_dff_A_iYCXIxq65_0),.clk(gclk));
	jdff dff_A_3XKw3vF77_0(.dout(w_dff_A_ATk9Yafj6_0),.din(w_dff_A_3XKw3vF77_0),.clk(gclk));
	jdff dff_A_ATk9Yafj6_0(.dout(w_dff_A_jgTXMd1D3_0),.din(w_dff_A_ATk9Yafj6_0),.clk(gclk));
	jdff dff_A_jgTXMd1D3_0(.dout(w_dff_A_UYBiSPz62_0),.din(w_dff_A_jgTXMd1D3_0),.clk(gclk));
	jdff dff_A_UYBiSPz62_0(.dout(w_dff_A_BXewrYB48_0),.din(w_dff_A_UYBiSPz62_0),.clk(gclk));
	jdff dff_A_BXewrYB48_0(.dout(G822),.din(w_dff_A_BXewrYB48_0),.clk(gclk));
	jdff dff_A_E3YaYj4k1_1(.dout(w_dff_A_GaVWyCWi6_0),.din(w_dff_A_E3YaYj4k1_1),.clk(gclk));
	jdff dff_A_GaVWyCWi6_0(.dout(w_dff_A_6RANbNUR6_0),.din(w_dff_A_GaVWyCWi6_0),.clk(gclk));
	jdff dff_A_6RANbNUR6_0(.dout(w_dff_A_APKok7Mx8_0),.din(w_dff_A_6RANbNUR6_0),.clk(gclk));
	jdff dff_A_APKok7Mx8_0(.dout(w_dff_A_dToRJRTv6_0),.din(w_dff_A_APKok7Mx8_0),.clk(gclk));
	jdff dff_A_dToRJRTv6_0(.dout(w_dff_A_DPKrV4l86_0),.din(w_dff_A_dToRJRTv6_0),.clk(gclk));
	jdff dff_A_DPKrV4l86_0(.dout(w_dff_A_CA9LWPdx7_0),.din(w_dff_A_DPKrV4l86_0),.clk(gclk));
	jdff dff_A_CA9LWPdx7_0(.dout(w_dff_A_U0qeOcNV5_0),.din(w_dff_A_CA9LWPdx7_0),.clk(gclk));
	jdff dff_A_U0qeOcNV5_0(.dout(w_dff_A_b1jmlzFU5_0),.din(w_dff_A_U0qeOcNV5_0),.clk(gclk));
	jdff dff_A_b1jmlzFU5_0(.dout(w_dff_A_lV6tL9Hb7_0),.din(w_dff_A_b1jmlzFU5_0),.clk(gclk));
	jdff dff_A_lV6tL9Hb7_0(.dout(w_dff_A_7fxiZP2l2_0),.din(w_dff_A_lV6tL9Hb7_0),.clk(gclk));
	jdff dff_A_7fxiZP2l2_0(.dout(w_dff_A_talPBM797_0),.din(w_dff_A_7fxiZP2l2_0),.clk(gclk));
	jdff dff_A_talPBM797_0(.dout(w_dff_A_3ojc82UW1_0),.din(w_dff_A_talPBM797_0),.clk(gclk));
	jdff dff_A_3ojc82UW1_0(.dout(w_dff_A_98adCmWY7_0),.din(w_dff_A_3ojc82UW1_0),.clk(gclk));
	jdff dff_A_98adCmWY7_0(.dout(w_dff_A_2JDsfYhm0_0),.din(w_dff_A_98adCmWY7_0),.clk(gclk));
	jdff dff_A_2JDsfYhm0_0(.dout(w_dff_A_vNzLAaKh6_0),.din(w_dff_A_2JDsfYhm0_0),.clk(gclk));
	jdff dff_A_vNzLAaKh6_0(.dout(w_dff_A_79Yqd6rA2_0),.din(w_dff_A_vNzLAaKh6_0),.clk(gclk));
	jdff dff_A_79Yqd6rA2_0(.dout(w_dff_A_ttEH5mM63_0),.din(w_dff_A_79Yqd6rA2_0),.clk(gclk));
	jdff dff_A_ttEH5mM63_0(.dout(G838),.din(w_dff_A_ttEH5mM63_0),.clk(gclk));
	jdff dff_A_A4wx6Pyj7_1(.dout(w_dff_A_x68XK9Bu2_0),.din(w_dff_A_A4wx6Pyj7_1),.clk(gclk));
	jdff dff_A_x68XK9Bu2_0(.dout(w_dff_A_stzO46h05_0),.din(w_dff_A_x68XK9Bu2_0),.clk(gclk));
	jdff dff_A_stzO46h05_0(.dout(w_dff_A_7XYiZ6wc2_0),.din(w_dff_A_stzO46h05_0),.clk(gclk));
	jdff dff_A_7XYiZ6wc2_0(.dout(w_dff_A_fvTuBpcE8_0),.din(w_dff_A_7XYiZ6wc2_0),.clk(gclk));
	jdff dff_A_fvTuBpcE8_0(.dout(w_dff_A_b2KY147M0_0),.din(w_dff_A_fvTuBpcE8_0),.clk(gclk));
	jdff dff_A_b2KY147M0_0(.dout(w_dff_A_XXLaziDU4_0),.din(w_dff_A_b2KY147M0_0),.clk(gclk));
	jdff dff_A_XXLaziDU4_0(.dout(w_dff_A_Nb9BxdPP4_0),.din(w_dff_A_XXLaziDU4_0),.clk(gclk));
	jdff dff_A_Nb9BxdPP4_0(.dout(w_dff_A_2E9AXDMD2_0),.din(w_dff_A_Nb9BxdPP4_0),.clk(gclk));
	jdff dff_A_2E9AXDMD2_0(.dout(w_dff_A_FXggS7873_0),.din(w_dff_A_2E9AXDMD2_0),.clk(gclk));
	jdff dff_A_FXggS7873_0(.dout(w_dff_A_a1WpbsJ89_0),.din(w_dff_A_FXggS7873_0),.clk(gclk));
	jdff dff_A_a1WpbsJ89_0(.dout(w_dff_A_3oDDxfvV7_0),.din(w_dff_A_a1WpbsJ89_0),.clk(gclk));
	jdff dff_A_3oDDxfvV7_0(.dout(w_dff_A_Ff62aGNT9_0),.din(w_dff_A_3oDDxfvV7_0),.clk(gclk));
	jdff dff_A_Ff62aGNT9_0(.dout(w_dff_A_FdUActS05_0),.din(w_dff_A_Ff62aGNT9_0),.clk(gclk));
	jdff dff_A_FdUActS05_0(.dout(w_dff_A_9NCUS5xc5_0),.din(w_dff_A_FdUActS05_0),.clk(gclk));
	jdff dff_A_9NCUS5xc5_0(.dout(w_dff_A_NI5tmFbJ7_0),.din(w_dff_A_9NCUS5xc5_0),.clk(gclk));
	jdff dff_A_NI5tmFbJ7_0(.dout(w_dff_A_GDeeSVIW2_0),.din(w_dff_A_NI5tmFbJ7_0),.clk(gclk));
	jdff dff_A_GDeeSVIW2_0(.dout(w_dff_A_xa8ghJdf6_0),.din(w_dff_A_GDeeSVIW2_0),.clk(gclk));
	jdff dff_A_xa8ghJdf6_0(.dout(G861),.din(w_dff_A_xa8ghJdf6_0),.clk(gclk));
	jdff dff_A_FnIaWamW8_1(.dout(w_dff_A_LuPtvtwU1_0),.din(w_dff_A_FnIaWamW8_1),.clk(gclk));
	jdff dff_A_LuPtvtwU1_0(.dout(w_dff_A_AXYs8PUz4_0),.din(w_dff_A_LuPtvtwU1_0),.clk(gclk));
	jdff dff_A_AXYs8PUz4_0(.dout(w_dff_A_FKcJVPB64_0),.din(w_dff_A_AXYs8PUz4_0),.clk(gclk));
	jdff dff_A_FKcJVPB64_0(.dout(w_dff_A_KVT10t0a9_0),.din(w_dff_A_FKcJVPB64_0),.clk(gclk));
	jdff dff_A_KVT10t0a9_0(.dout(w_dff_A_lBqJxuSC9_0),.din(w_dff_A_KVT10t0a9_0),.clk(gclk));
	jdff dff_A_lBqJxuSC9_0(.dout(w_dff_A_A5K3ofS42_0),.din(w_dff_A_lBqJxuSC9_0),.clk(gclk));
	jdff dff_A_A5K3ofS42_0(.dout(G623),.din(w_dff_A_A5K3ofS42_0),.clk(gclk));
	jdff dff_A_rihHI8OF6_2(.dout(w_dff_A_eeI1Jxay0_0),.din(w_dff_A_rihHI8OF6_2),.clk(gclk));
	jdff dff_A_eeI1Jxay0_0(.dout(w_dff_A_OID7a4sf6_0),.din(w_dff_A_eeI1Jxay0_0),.clk(gclk));
	jdff dff_A_OID7a4sf6_0(.dout(w_dff_A_55xCm2xS7_0),.din(w_dff_A_OID7a4sf6_0),.clk(gclk));
	jdff dff_A_55xCm2xS7_0(.dout(w_dff_A_bOqR8A041_0),.din(w_dff_A_55xCm2xS7_0),.clk(gclk));
	jdff dff_A_bOqR8A041_0(.dout(w_dff_A_8O4T1LoU1_0),.din(w_dff_A_bOqR8A041_0),.clk(gclk));
	jdff dff_A_8O4T1LoU1_0(.dout(w_dff_A_HZEnsD2K1_0),.din(w_dff_A_8O4T1LoU1_0),.clk(gclk));
	jdff dff_A_HZEnsD2K1_0(.dout(w_dff_A_hlx3HPY17_0),.din(w_dff_A_HZEnsD2K1_0),.clk(gclk));
	jdff dff_A_hlx3HPY17_0(.dout(w_dff_A_xrxJ6JMc9_0),.din(w_dff_A_hlx3HPY17_0),.clk(gclk));
	jdff dff_A_xrxJ6JMc9_0(.dout(w_dff_A_gKWlEoYD7_0),.din(w_dff_A_xrxJ6JMc9_0),.clk(gclk));
	jdff dff_A_gKWlEoYD7_0(.dout(w_dff_A_ao8qu1wi5_0),.din(w_dff_A_gKWlEoYD7_0),.clk(gclk));
	jdff dff_A_ao8qu1wi5_0(.dout(w_dff_A_rjySDON30_0),.din(w_dff_A_ao8qu1wi5_0),.clk(gclk));
	jdff dff_A_rjySDON30_0(.dout(w_dff_A_ryfqMpwG1_0),.din(w_dff_A_rjySDON30_0),.clk(gclk));
	jdff dff_A_ryfqMpwG1_0(.dout(w_dff_A_Ccq3ENsc4_0),.din(w_dff_A_ryfqMpwG1_0),.clk(gclk));
	jdff dff_A_Ccq3ENsc4_0(.dout(w_dff_A_FVQW5aGI6_0),.din(w_dff_A_Ccq3ENsc4_0),.clk(gclk));
	jdff dff_A_FVQW5aGI6_0(.dout(G722),.din(w_dff_A_FVQW5aGI6_0),.clk(gclk));
	jdff dff_A_uwSrejso2_1(.dout(w_dff_A_qnVcuwuj1_0),.din(w_dff_A_uwSrejso2_1),.clk(gclk));
	jdff dff_A_qnVcuwuj1_0(.dout(w_dff_A_nx1js3GU7_0),.din(w_dff_A_qnVcuwuj1_0),.clk(gclk));
	jdff dff_A_nx1js3GU7_0(.dout(w_dff_A_VyItlWFG2_0),.din(w_dff_A_nx1js3GU7_0),.clk(gclk));
	jdff dff_A_VyItlWFG2_0(.dout(w_dff_A_WxS5WOep8_0),.din(w_dff_A_VyItlWFG2_0),.clk(gclk));
	jdff dff_A_WxS5WOep8_0(.dout(w_dff_A_bsHJIzgf4_0),.din(w_dff_A_WxS5WOep8_0),.clk(gclk));
	jdff dff_A_bsHJIzgf4_0(.dout(w_dff_A_SjmwnRyf1_0),.din(w_dff_A_bsHJIzgf4_0),.clk(gclk));
	jdff dff_A_SjmwnRyf1_0(.dout(w_dff_A_8LZyY8y66_0),.din(w_dff_A_SjmwnRyf1_0),.clk(gclk));
	jdff dff_A_8LZyY8y66_0(.dout(w_dff_A_tgDbKMGN3_0),.din(w_dff_A_8LZyY8y66_0),.clk(gclk));
	jdff dff_A_tgDbKMGN3_0(.dout(w_dff_A_0kykd7A99_0),.din(w_dff_A_tgDbKMGN3_0),.clk(gclk));
	jdff dff_A_0kykd7A99_0(.dout(w_dff_A_WxpaqE778_0),.din(w_dff_A_0kykd7A99_0),.clk(gclk));
	jdff dff_A_WxpaqE778_0(.dout(w_dff_A_FyKjELc89_0),.din(w_dff_A_WxpaqE778_0),.clk(gclk));
	jdff dff_A_FyKjELc89_0(.dout(G832),.din(w_dff_A_FyKjELc89_0),.clk(gclk));
	jdff dff_A_aPDiXqIJ5_1(.dout(w_dff_A_jNaqojDm6_0),.din(w_dff_A_aPDiXqIJ5_1),.clk(gclk));
	jdff dff_A_jNaqojDm6_0(.dout(w_dff_A_W2K8uwQ28_0),.din(w_dff_A_jNaqojDm6_0),.clk(gclk));
	jdff dff_A_W2K8uwQ28_0(.dout(w_dff_A_eC56YHPc0_0),.din(w_dff_A_W2K8uwQ28_0),.clk(gclk));
	jdff dff_A_eC56YHPc0_0(.dout(w_dff_A_jvbCF3kw6_0),.din(w_dff_A_eC56YHPc0_0),.clk(gclk));
	jdff dff_A_jvbCF3kw6_0(.dout(w_dff_A_gPnaKhCS8_0),.din(w_dff_A_jvbCF3kw6_0),.clk(gclk));
	jdff dff_A_gPnaKhCS8_0(.dout(w_dff_A_5o62JWbn0_0),.din(w_dff_A_gPnaKhCS8_0),.clk(gclk));
	jdff dff_A_5o62JWbn0_0(.dout(w_dff_A_3y4AB5eA4_0),.din(w_dff_A_5o62JWbn0_0),.clk(gclk));
	jdff dff_A_3y4AB5eA4_0(.dout(w_dff_A_9AJ9G0cl9_0),.din(w_dff_A_3y4AB5eA4_0),.clk(gclk));
	jdff dff_A_9AJ9G0cl9_0(.dout(w_dff_A_i4oXyeDj5_0),.din(w_dff_A_9AJ9G0cl9_0),.clk(gclk));
	jdff dff_A_i4oXyeDj5_0(.dout(w_dff_A_I23kZXU87_0),.din(w_dff_A_i4oXyeDj5_0),.clk(gclk));
	jdff dff_A_I23kZXU87_0(.dout(w_dff_A_l5dGryT81_0),.din(w_dff_A_I23kZXU87_0),.clk(gclk));
	jdff dff_A_l5dGryT81_0(.dout(w_dff_A_LZdknmCY0_0),.din(w_dff_A_l5dGryT81_0),.clk(gclk));
	jdff dff_A_LZdknmCY0_0(.dout(w_dff_A_u1r3E6Lz7_0),.din(w_dff_A_LZdknmCY0_0),.clk(gclk));
	jdff dff_A_u1r3E6Lz7_0(.dout(G834),.din(w_dff_A_u1r3E6Lz7_0),.clk(gclk));
	jdff dff_A_oZ7aU2kK3_1(.dout(w_dff_A_uPCk3orv8_0),.din(w_dff_A_oZ7aU2kK3_1),.clk(gclk));
	jdff dff_A_uPCk3orv8_0(.dout(w_dff_A_E3loVfFT8_0),.din(w_dff_A_uPCk3orv8_0),.clk(gclk));
	jdff dff_A_E3loVfFT8_0(.dout(w_dff_A_a4aICiYl3_0),.din(w_dff_A_E3loVfFT8_0),.clk(gclk));
	jdff dff_A_a4aICiYl3_0(.dout(w_dff_A_bWO7ZxzZ0_0),.din(w_dff_A_a4aICiYl3_0),.clk(gclk));
	jdff dff_A_bWO7ZxzZ0_0(.dout(w_dff_A_iElLYdJA5_0),.din(w_dff_A_bWO7ZxzZ0_0),.clk(gclk));
	jdff dff_A_iElLYdJA5_0(.dout(w_dff_A_sCfjvzOF9_0),.din(w_dff_A_iElLYdJA5_0),.clk(gclk));
	jdff dff_A_sCfjvzOF9_0(.dout(w_dff_A_u2rWZShp9_0),.din(w_dff_A_sCfjvzOF9_0),.clk(gclk));
	jdff dff_A_u2rWZShp9_0(.dout(w_dff_A_ZqTfgCM72_0),.din(w_dff_A_u2rWZShp9_0),.clk(gclk));
	jdff dff_A_ZqTfgCM72_0(.dout(w_dff_A_7XkPEuzN8_0),.din(w_dff_A_ZqTfgCM72_0),.clk(gclk));
	jdff dff_A_7XkPEuzN8_0(.dout(w_dff_A_EiyyASsV5_0),.din(w_dff_A_7XkPEuzN8_0),.clk(gclk));
	jdff dff_A_EiyyASsV5_0(.dout(w_dff_A_beys8m2r1_0),.din(w_dff_A_EiyyASsV5_0),.clk(gclk));
	jdff dff_A_beys8m2r1_0(.dout(w_dff_A_iVwUzesP6_0),.din(w_dff_A_beys8m2r1_0),.clk(gclk));
	jdff dff_A_iVwUzesP6_0(.dout(w_dff_A_g0bV30pU2_0),.din(w_dff_A_iVwUzesP6_0),.clk(gclk));
	jdff dff_A_g0bV30pU2_0(.dout(w_dff_A_SyfuU3iZ7_0),.din(w_dff_A_g0bV30pU2_0),.clk(gclk));
	jdff dff_A_SyfuU3iZ7_0(.dout(w_dff_A_1ouZPPoB1_0),.din(w_dff_A_SyfuU3iZ7_0),.clk(gclk));
	jdff dff_A_1ouZPPoB1_0(.dout(G836),.din(w_dff_A_1ouZPPoB1_0),.clk(gclk));
	jdff dff_A_89q19c2f0_2(.dout(w_dff_A_Ypvo3d9D6_0),.din(w_dff_A_89q19c2f0_2),.clk(gclk));
	jdff dff_A_Ypvo3d9D6_0(.dout(w_dff_A_14VL949c5_0),.din(w_dff_A_Ypvo3d9D6_0),.clk(gclk));
	jdff dff_A_14VL949c5_0(.dout(w_dff_A_K739I5T62_0),.din(w_dff_A_14VL949c5_0),.clk(gclk));
	jdff dff_A_K739I5T62_0(.dout(w_dff_A_5m158jww1_0),.din(w_dff_A_K739I5T62_0),.clk(gclk));
	jdff dff_A_5m158jww1_0(.dout(w_dff_A_yx4Be42c0_0),.din(w_dff_A_5m158jww1_0),.clk(gclk));
	jdff dff_A_yx4Be42c0_0(.dout(w_dff_A_IzKVrTnF2_0),.din(w_dff_A_yx4Be42c0_0),.clk(gclk));
	jdff dff_A_IzKVrTnF2_0(.dout(w_dff_A_NkjrtaDa3_0),.din(w_dff_A_IzKVrTnF2_0),.clk(gclk));
	jdff dff_A_NkjrtaDa3_0(.dout(w_dff_A_p2ptYhKI1_0),.din(w_dff_A_NkjrtaDa3_0),.clk(gclk));
	jdff dff_A_p2ptYhKI1_0(.dout(w_dff_A_nUA2XqSZ3_0),.din(w_dff_A_p2ptYhKI1_0),.clk(gclk));
	jdff dff_A_nUA2XqSZ3_0(.dout(w_dff_A_SsrVvxOi9_0),.din(w_dff_A_nUA2XqSZ3_0),.clk(gclk));
	jdff dff_A_SsrVvxOi9_0(.dout(w_dff_A_WefwJ0vb9_0),.din(w_dff_A_SsrVvxOi9_0),.clk(gclk));
	jdff dff_A_WefwJ0vb9_0(.dout(w_dff_A_tBWTraNr8_0),.din(w_dff_A_WefwJ0vb9_0),.clk(gclk));
	jdff dff_A_tBWTraNr8_0(.dout(w_dff_A_K2ITEvA84_0),.din(w_dff_A_tBWTraNr8_0),.clk(gclk));
	jdff dff_A_K2ITEvA84_0(.dout(w_dff_A_q5P2WgGR7_0),.din(w_dff_A_K2ITEvA84_0),.clk(gclk));
	jdff dff_A_q5P2WgGR7_0(.dout(G859),.din(w_dff_A_q5P2WgGR7_0),.clk(gclk));
	jdff dff_A_FEyi87VO8_1(.dout(w_dff_A_g4BCbAGH7_0),.din(w_dff_A_FEyi87VO8_1),.clk(gclk));
	jdff dff_A_g4BCbAGH7_0(.dout(w_dff_A_wjhtsViz9_0),.din(w_dff_A_g4BCbAGH7_0),.clk(gclk));
	jdff dff_A_wjhtsViz9_0(.dout(w_dff_A_xARsMCBG9_0),.din(w_dff_A_wjhtsViz9_0),.clk(gclk));
	jdff dff_A_xARsMCBG9_0(.dout(w_dff_A_0Z21CPDY7_0),.din(w_dff_A_xARsMCBG9_0),.clk(gclk));
	jdff dff_A_0Z21CPDY7_0(.dout(w_dff_A_czH35Aou9_0),.din(w_dff_A_0Z21CPDY7_0),.clk(gclk));
	jdff dff_A_czH35Aou9_0(.dout(w_dff_A_Sb4LqZoM2_0),.din(w_dff_A_czH35Aou9_0),.clk(gclk));
	jdff dff_A_Sb4LqZoM2_0(.dout(w_dff_A_48AlIWm59_0),.din(w_dff_A_Sb4LqZoM2_0),.clk(gclk));
	jdff dff_A_48AlIWm59_0(.dout(w_dff_A_43Z0e5Zk7_0),.din(w_dff_A_48AlIWm59_0),.clk(gclk));
	jdff dff_A_43Z0e5Zk7_0(.dout(w_dff_A_IpvMKZ2f3_0),.din(w_dff_A_43Z0e5Zk7_0),.clk(gclk));
	jdff dff_A_IpvMKZ2f3_0(.dout(G871),.din(w_dff_A_IpvMKZ2f3_0),.clk(gclk));
	jdff dff_A_tbRIqskU5_1(.dout(w_dff_A_jMFEEjMW7_0),.din(w_dff_A_tbRIqskU5_1),.clk(gclk));
	jdff dff_A_jMFEEjMW7_0(.dout(w_dff_A_H7hzk3cm5_0),.din(w_dff_A_jMFEEjMW7_0),.clk(gclk));
	jdff dff_A_H7hzk3cm5_0(.dout(w_dff_A_s6bBg3Zs0_0),.din(w_dff_A_H7hzk3cm5_0),.clk(gclk));
	jdff dff_A_s6bBg3Zs0_0(.dout(w_dff_A_YldWtFF73_0),.din(w_dff_A_s6bBg3Zs0_0),.clk(gclk));
	jdff dff_A_YldWtFF73_0(.dout(w_dff_A_vv40dYLN9_0),.din(w_dff_A_YldWtFF73_0),.clk(gclk));
	jdff dff_A_vv40dYLN9_0(.dout(w_dff_A_FaAOVuM28_0),.din(w_dff_A_vv40dYLN9_0),.clk(gclk));
	jdff dff_A_FaAOVuM28_0(.dout(w_dff_A_xNzHx3ek6_0),.din(w_dff_A_FaAOVuM28_0),.clk(gclk));
	jdff dff_A_xNzHx3ek6_0(.dout(w_dff_A_EnZ2ah4O2_0),.din(w_dff_A_xNzHx3ek6_0),.clk(gclk));
	jdff dff_A_EnZ2ah4O2_0(.dout(w_dff_A_bYz1awt74_0),.din(w_dff_A_EnZ2ah4O2_0),.clk(gclk));
	jdff dff_A_bYz1awt74_0(.dout(w_dff_A_COjP7ukv2_0),.din(w_dff_A_bYz1awt74_0),.clk(gclk));
	jdff dff_A_COjP7ukv2_0(.dout(w_dff_A_XU7UePSo6_0),.din(w_dff_A_COjP7ukv2_0),.clk(gclk));
	jdff dff_A_XU7UePSo6_0(.dout(G873),.din(w_dff_A_XU7UePSo6_0),.clk(gclk));
	jdff dff_A_mfZM6VHe2_1(.dout(w_dff_A_2Z2QYpFd4_0),.din(w_dff_A_mfZM6VHe2_1),.clk(gclk));
	jdff dff_A_2Z2QYpFd4_0(.dout(w_dff_A_DeUiF1kp8_0),.din(w_dff_A_2Z2QYpFd4_0),.clk(gclk));
	jdff dff_A_DeUiF1kp8_0(.dout(w_dff_A_IyahUs1U7_0),.din(w_dff_A_DeUiF1kp8_0),.clk(gclk));
	jdff dff_A_IyahUs1U7_0(.dout(w_dff_A_nT7nrwXk7_0),.din(w_dff_A_IyahUs1U7_0),.clk(gclk));
	jdff dff_A_nT7nrwXk7_0(.dout(w_dff_A_VPe2t4FT5_0),.din(w_dff_A_nT7nrwXk7_0),.clk(gclk));
	jdff dff_A_VPe2t4FT5_0(.dout(w_dff_A_vp1eqQtn9_0),.din(w_dff_A_VPe2t4FT5_0),.clk(gclk));
	jdff dff_A_vp1eqQtn9_0(.dout(w_dff_A_owdiU8qH9_0),.din(w_dff_A_vp1eqQtn9_0),.clk(gclk));
	jdff dff_A_owdiU8qH9_0(.dout(w_dff_A_G8uOQpYS1_0),.din(w_dff_A_owdiU8qH9_0),.clk(gclk));
	jdff dff_A_G8uOQpYS1_0(.dout(w_dff_A_5GlFC2W62_0),.din(w_dff_A_G8uOQpYS1_0),.clk(gclk));
	jdff dff_A_5GlFC2W62_0(.dout(w_dff_A_Dop3JM336_0),.din(w_dff_A_5GlFC2W62_0),.clk(gclk));
	jdff dff_A_Dop3JM336_0(.dout(w_dff_A_Yk4AJPXb0_0),.din(w_dff_A_Dop3JM336_0),.clk(gclk));
	jdff dff_A_Yk4AJPXb0_0(.dout(w_dff_A_BnLjLJI84_0),.din(w_dff_A_Yk4AJPXb0_0),.clk(gclk));
	jdff dff_A_BnLjLJI84_0(.dout(G875),.din(w_dff_A_BnLjLJI84_0),.clk(gclk));
	jdff dff_A_znHZByz42_1(.dout(w_dff_A_bkWzsQ1I4_0),.din(w_dff_A_znHZByz42_1),.clk(gclk));
	jdff dff_A_bkWzsQ1I4_0(.dout(w_dff_A_sQWx8T7X6_0),.din(w_dff_A_bkWzsQ1I4_0),.clk(gclk));
	jdff dff_A_sQWx8T7X6_0(.dout(w_dff_A_XxRApIf52_0),.din(w_dff_A_sQWx8T7X6_0),.clk(gclk));
	jdff dff_A_XxRApIf52_0(.dout(w_dff_A_A1KtQVro2_0),.din(w_dff_A_XxRApIf52_0),.clk(gclk));
	jdff dff_A_A1KtQVro2_0(.dout(w_dff_A_fIrn3unf0_0),.din(w_dff_A_A1KtQVro2_0),.clk(gclk));
	jdff dff_A_fIrn3unf0_0(.dout(w_dff_A_oCaCzonU1_0),.din(w_dff_A_fIrn3unf0_0),.clk(gclk));
	jdff dff_A_oCaCzonU1_0(.dout(w_dff_A_0oIqhyer7_0),.din(w_dff_A_oCaCzonU1_0),.clk(gclk));
	jdff dff_A_0oIqhyer7_0(.dout(w_dff_A_LI6TumCQ7_0),.din(w_dff_A_0oIqhyer7_0),.clk(gclk));
	jdff dff_A_LI6TumCQ7_0(.dout(w_dff_A_JGhTj1ON6_0),.din(w_dff_A_LI6TumCQ7_0),.clk(gclk));
	jdff dff_A_JGhTj1ON6_0(.dout(w_dff_A_1WWVbI2O2_0),.din(w_dff_A_JGhTj1ON6_0),.clk(gclk));
	jdff dff_A_1WWVbI2O2_0(.dout(w_dff_A_BLXfFyri2_0),.din(w_dff_A_1WWVbI2O2_0),.clk(gclk));
	jdff dff_A_BLXfFyri2_0(.dout(w_dff_A_DqE5aA3t1_0),.din(w_dff_A_BLXfFyri2_0),.clk(gclk));
	jdff dff_A_DqE5aA3t1_0(.dout(w_dff_A_uUU8ObDp9_0),.din(w_dff_A_DqE5aA3t1_0),.clk(gclk));
	jdff dff_A_uUU8ObDp9_0(.dout(G877),.din(w_dff_A_uUU8ObDp9_0),.clk(gclk));
	jdff dff_A_DRK3FxjO7_1(.dout(w_dff_A_LdVKKNJk3_0),.din(w_dff_A_DRK3FxjO7_1),.clk(gclk));
	jdff dff_A_LdVKKNJk3_0(.dout(w_dff_A_vPBu5CHI5_0),.din(w_dff_A_LdVKKNJk3_0),.clk(gclk));
	jdff dff_A_vPBu5CHI5_0(.dout(w_dff_A_d5Y9Q4os1_0),.din(w_dff_A_vPBu5CHI5_0),.clk(gclk));
	jdff dff_A_d5Y9Q4os1_0(.dout(w_dff_A_rifLNMZb9_0),.din(w_dff_A_d5Y9Q4os1_0),.clk(gclk));
	jdff dff_A_rifLNMZb9_0(.dout(w_dff_A_tXLLOhGW7_0),.din(w_dff_A_rifLNMZb9_0),.clk(gclk));
	jdff dff_A_tXLLOhGW7_0(.dout(w_dff_A_fFGPrXvU8_0),.din(w_dff_A_tXLLOhGW7_0),.clk(gclk));
	jdff dff_A_fFGPrXvU8_0(.dout(w_dff_A_tqFdZqy68_0),.din(w_dff_A_fFGPrXvU8_0),.clk(gclk));
	jdff dff_A_tqFdZqy68_0(.dout(w_dff_A_Y8W3ZcjZ7_0),.din(w_dff_A_tqFdZqy68_0),.clk(gclk));
	jdff dff_A_Y8W3ZcjZ7_0(.dout(w_dff_A_jD3nV72H4_0),.din(w_dff_A_Y8W3ZcjZ7_0),.clk(gclk));
	jdff dff_A_jD3nV72H4_0(.dout(w_dff_A_edx1i5tO4_0),.din(w_dff_A_jD3nV72H4_0),.clk(gclk));
	jdff dff_A_edx1i5tO4_0(.dout(w_dff_A_P0Pt5xk05_0),.din(w_dff_A_edx1i5tO4_0),.clk(gclk));
	jdff dff_A_P0Pt5xk05_0(.dout(w_dff_A_246iYMQa6_0),.din(w_dff_A_P0Pt5xk05_0),.clk(gclk));
	jdff dff_A_246iYMQa6_0(.dout(w_dff_A_rLiQtCLX5_0),.din(w_dff_A_246iYMQa6_0),.clk(gclk));
	jdff dff_A_rLiQtCLX5_0(.dout(w_dff_A_MGmmWgBm1_0),.din(w_dff_A_rLiQtCLX5_0),.clk(gclk));
	jdff dff_A_MGmmWgBm1_0(.dout(w_dff_A_rOj99gq84_0),.din(w_dff_A_MGmmWgBm1_0),.clk(gclk));
	jdff dff_A_rOj99gq84_0(.dout(w_dff_A_hEiH5Yli0_0),.din(w_dff_A_rOj99gq84_0),.clk(gclk));
	jdff dff_A_hEiH5Yli0_0(.dout(G998),.din(w_dff_A_hEiH5Yli0_0),.clk(gclk));
	jdff dff_A_BMw7y2Ba7_1(.dout(w_dff_A_85Zvejto0_0),.din(w_dff_A_BMw7y2Ba7_1),.clk(gclk));
	jdff dff_A_85Zvejto0_0(.dout(w_dff_A_xEBOynEa0_0),.din(w_dff_A_85Zvejto0_0),.clk(gclk));
	jdff dff_A_xEBOynEa0_0(.dout(w_dff_A_XWd0Ya9Q3_0),.din(w_dff_A_xEBOynEa0_0),.clk(gclk));
	jdff dff_A_XWd0Ya9Q3_0(.dout(w_dff_A_9HGnU0W98_0),.din(w_dff_A_XWd0Ya9Q3_0),.clk(gclk));
	jdff dff_A_9HGnU0W98_0(.dout(w_dff_A_TGUJ1Fp62_0),.din(w_dff_A_9HGnU0W98_0),.clk(gclk));
	jdff dff_A_TGUJ1Fp62_0(.dout(w_dff_A_i2aa1icl5_0),.din(w_dff_A_TGUJ1Fp62_0),.clk(gclk));
	jdff dff_A_i2aa1icl5_0(.dout(w_dff_A_9rCsXmKf0_0),.din(w_dff_A_i2aa1icl5_0),.clk(gclk));
	jdff dff_A_9rCsXmKf0_0(.dout(w_dff_A_y5ERnFou8_0),.din(w_dff_A_9rCsXmKf0_0),.clk(gclk));
	jdff dff_A_y5ERnFou8_0(.dout(w_dff_A_twHqRVW34_0),.din(w_dff_A_y5ERnFou8_0),.clk(gclk));
	jdff dff_A_twHqRVW34_0(.dout(w_dff_A_wl96eY8Y5_0),.din(w_dff_A_twHqRVW34_0),.clk(gclk));
	jdff dff_A_wl96eY8Y5_0(.dout(w_dff_A_oD8hCD429_0),.din(w_dff_A_wl96eY8Y5_0),.clk(gclk));
	jdff dff_A_oD8hCD429_0(.dout(w_dff_A_GcBTACSu1_0),.din(w_dff_A_oD8hCD429_0),.clk(gclk));
	jdff dff_A_GcBTACSu1_0(.dout(w_dff_A_kgLVwoGE1_0),.din(w_dff_A_GcBTACSu1_0),.clk(gclk));
	jdff dff_A_kgLVwoGE1_0(.dout(w_dff_A_qDdY1JAL2_0),.din(w_dff_A_kgLVwoGE1_0),.clk(gclk));
	jdff dff_A_qDdY1JAL2_0(.dout(w_dff_A_5iNAJwdU9_0),.din(w_dff_A_qDdY1JAL2_0),.clk(gclk));
	jdff dff_A_5iNAJwdU9_0(.dout(w_dff_A_B3HaQMSk3_0),.din(w_dff_A_5iNAJwdU9_0),.clk(gclk));
	jdff dff_A_B3HaQMSk3_0(.dout(w_dff_A_u6GuB5Nt4_0),.din(w_dff_A_B3HaQMSk3_0),.clk(gclk));
	jdff dff_A_u6GuB5Nt4_0(.dout(w_dff_A_TjcllJTG9_0),.din(w_dff_A_u6GuB5Nt4_0),.clk(gclk));
	jdff dff_A_TjcllJTG9_0(.dout(G1000),.din(w_dff_A_TjcllJTG9_0),.clk(gclk));
	jdff dff_A_Fwk1ch9u3_2(.dout(w_dff_A_o8oOY3LR4_0),.din(w_dff_A_Fwk1ch9u3_2),.clk(gclk));
	jdff dff_A_o8oOY3LR4_0(.dout(w_dff_A_AjGncHWn6_0),.din(w_dff_A_o8oOY3LR4_0),.clk(gclk));
	jdff dff_A_AjGncHWn6_0(.dout(w_dff_A_RqljxeTi6_0),.din(w_dff_A_AjGncHWn6_0),.clk(gclk));
	jdff dff_A_RqljxeTi6_0(.dout(w_dff_A_igU8JoqH3_0),.din(w_dff_A_RqljxeTi6_0),.clk(gclk));
	jdff dff_A_igU8JoqH3_0(.dout(G575),.din(w_dff_A_igU8JoqH3_0),.clk(gclk));
	jdff dff_A_Z53KL96c4_2(.dout(w_dff_A_5mJ2m0Ek4_0),.din(w_dff_A_Z53KL96c4_2),.clk(gclk));
	jdff dff_A_5mJ2m0Ek4_0(.dout(w_dff_A_gpkqj7kl2_0),.din(w_dff_A_5mJ2m0Ek4_0),.clk(gclk));
	jdff dff_A_gpkqj7kl2_0(.dout(w_dff_A_v8GOvxvW2_0),.din(w_dff_A_gpkqj7kl2_0),.clk(gclk));
	jdff dff_A_v8GOvxvW2_0(.dout(w_dff_A_D3bAE0a97_0),.din(w_dff_A_v8GOvxvW2_0),.clk(gclk));
	jdff dff_A_D3bAE0a97_0(.dout(w_dff_A_RBfckbjc4_0),.din(w_dff_A_D3bAE0a97_0),.clk(gclk));
	jdff dff_A_RBfckbjc4_0(.dout(w_dff_A_gmvIMtBQ3_0),.din(w_dff_A_RBfckbjc4_0),.clk(gclk));
	jdff dff_A_gmvIMtBQ3_0(.dout(w_dff_A_uf72IVJc7_0),.din(w_dff_A_gmvIMtBQ3_0),.clk(gclk));
	jdff dff_A_uf72IVJc7_0(.dout(G585),.din(w_dff_A_uf72IVJc7_0),.clk(gclk));
	jdff dff_A_D17Lvw550_2(.dout(w_dff_A_Nl0vYpIb0_0),.din(w_dff_A_D17Lvw550_2),.clk(gclk));
	jdff dff_A_Nl0vYpIb0_0(.dout(w_dff_A_EZFQrtM53_0),.din(w_dff_A_Nl0vYpIb0_0),.clk(gclk));
	jdff dff_A_EZFQrtM53_0(.dout(w_dff_A_TqrqK8yW0_0),.din(w_dff_A_EZFQrtM53_0),.clk(gclk));
	jdff dff_A_TqrqK8yW0_0(.dout(w_dff_A_43TVzXho1_0),.din(w_dff_A_TqrqK8yW0_0),.clk(gclk));
	jdff dff_A_43TVzXho1_0(.dout(w_dff_A_GFDcnW2p4_0),.din(w_dff_A_43TVzXho1_0),.clk(gclk));
	jdff dff_A_GFDcnW2p4_0(.dout(w_dff_A_9wvA3qCw4_0),.din(w_dff_A_GFDcnW2p4_0),.clk(gclk));
	jdff dff_A_9wvA3qCw4_0(.dout(w_dff_A_n31SPELV6_0),.din(w_dff_A_9wvA3qCw4_0),.clk(gclk));
	jdff dff_A_n31SPELV6_0(.dout(w_dff_A_jIjvrTmC1_0),.din(w_dff_A_n31SPELV6_0),.clk(gclk));
	jdff dff_A_jIjvrTmC1_0(.dout(w_dff_A_BSvfZcAU7_0),.din(w_dff_A_jIjvrTmC1_0),.clk(gclk));
	jdff dff_A_BSvfZcAU7_0(.dout(w_dff_A_nwXmLbGK1_0),.din(w_dff_A_BSvfZcAU7_0),.clk(gclk));
	jdff dff_A_nwXmLbGK1_0(.dout(w_dff_A_8uShcWI16_0),.din(w_dff_A_nwXmLbGK1_0),.clk(gclk));
	jdff dff_A_8uShcWI16_0(.dout(w_dff_A_B2yupq7I3_0),.din(w_dff_A_8uShcWI16_0),.clk(gclk));
	jdff dff_A_B2yupq7I3_0(.dout(w_dff_A_b8A31Ifd6_0),.din(w_dff_A_B2yupq7I3_0),.clk(gclk));
	jdff dff_A_b8A31Ifd6_0(.dout(G661),.din(w_dff_A_b8A31Ifd6_0),.clk(gclk));
	jdff dff_A_vv4HfquM5_2(.dout(w_dff_A_KkjXm6oy9_0),.din(w_dff_A_vv4HfquM5_2),.clk(gclk));
	jdff dff_A_KkjXm6oy9_0(.dout(w_dff_A_b7qG6Eah3_0),.din(w_dff_A_KkjXm6oy9_0),.clk(gclk));
	jdff dff_A_b7qG6Eah3_0(.dout(w_dff_A_dFXod8zO7_0),.din(w_dff_A_b7qG6Eah3_0),.clk(gclk));
	jdff dff_A_dFXod8zO7_0(.dout(w_dff_A_FFtiDZHx9_0),.din(w_dff_A_dFXod8zO7_0),.clk(gclk));
	jdff dff_A_FFtiDZHx9_0(.dout(w_dff_A_Hhjb7vcS3_0),.din(w_dff_A_FFtiDZHx9_0),.clk(gclk));
	jdff dff_A_Hhjb7vcS3_0(.dout(w_dff_A_s6hIwy4Y9_0),.din(w_dff_A_Hhjb7vcS3_0),.clk(gclk));
	jdff dff_A_s6hIwy4Y9_0(.dout(w_dff_A_hFTaZZPg3_0),.din(w_dff_A_s6hIwy4Y9_0),.clk(gclk));
	jdff dff_A_hFTaZZPg3_0(.dout(w_dff_A_p0oUpqlK1_0),.din(w_dff_A_hFTaZZPg3_0),.clk(gclk));
	jdff dff_A_p0oUpqlK1_0(.dout(w_dff_A_RAhw5FkQ9_0),.din(w_dff_A_p0oUpqlK1_0),.clk(gclk));
	jdff dff_A_RAhw5FkQ9_0(.dout(w_dff_A_YryeKUfV2_0),.din(w_dff_A_RAhw5FkQ9_0),.clk(gclk));
	jdff dff_A_YryeKUfV2_0(.dout(w_dff_A_JdqdH2V45_0),.din(w_dff_A_YryeKUfV2_0),.clk(gclk));
	jdff dff_A_JdqdH2V45_0(.dout(w_dff_A_ugyEBPjS9_0),.din(w_dff_A_JdqdH2V45_0),.clk(gclk));
	jdff dff_A_ugyEBPjS9_0(.dout(w_dff_A_CseCJxZM2_0),.din(w_dff_A_ugyEBPjS9_0),.clk(gclk));
	jdff dff_A_CseCJxZM2_0(.dout(G693),.din(w_dff_A_CseCJxZM2_0),.clk(gclk));
	jdff dff_A_4Kw7kf7E8_2(.dout(w_dff_A_q03HGYQX7_0),.din(w_dff_A_4Kw7kf7E8_2),.clk(gclk));
	jdff dff_A_q03HGYQX7_0(.dout(w_dff_A_k2zxiMXj1_0),.din(w_dff_A_q03HGYQX7_0),.clk(gclk));
	jdff dff_A_k2zxiMXj1_0(.dout(w_dff_A_i8B80i0D0_0),.din(w_dff_A_k2zxiMXj1_0),.clk(gclk));
	jdff dff_A_i8B80i0D0_0(.dout(w_dff_A_sPy6G2BC2_0),.din(w_dff_A_i8B80i0D0_0),.clk(gclk));
	jdff dff_A_sPy6G2BC2_0(.dout(w_dff_A_KtRbgIqS5_0),.din(w_dff_A_sPy6G2BC2_0),.clk(gclk));
	jdff dff_A_KtRbgIqS5_0(.dout(w_dff_A_Rx4OdOu72_0),.din(w_dff_A_KtRbgIqS5_0),.clk(gclk));
	jdff dff_A_Rx4OdOu72_0(.dout(G747),.din(w_dff_A_Rx4OdOu72_0),.clk(gclk));
	jdff dff_A_J3ukU9lO6_2(.dout(w_dff_A_bPu5C7j15_0),.din(w_dff_A_J3ukU9lO6_2),.clk(gclk));
	jdff dff_A_bPu5C7j15_0(.dout(w_dff_A_6WgIFvcY2_0),.din(w_dff_A_bPu5C7j15_0),.clk(gclk));
	jdff dff_A_6WgIFvcY2_0(.dout(w_dff_A_1hRwUTZd1_0),.din(w_dff_A_6WgIFvcY2_0),.clk(gclk));
	jdff dff_A_1hRwUTZd1_0(.dout(w_dff_A_jREYj0yz0_0),.din(w_dff_A_1hRwUTZd1_0),.clk(gclk));
	jdff dff_A_jREYj0yz0_0(.dout(w_dff_A_fb5Ztfsv2_0),.din(w_dff_A_jREYj0yz0_0),.clk(gclk));
	jdff dff_A_fb5Ztfsv2_0(.dout(w_dff_A_JQIK37c57_0),.din(w_dff_A_fb5Ztfsv2_0),.clk(gclk));
	jdff dff_A_JQIK37c57_0(.dout(w_dff_A_UPgCFFjT2_0),.din(w_dff_A_JQIK37c57_0),.clk(gclk));
	jdff dff_A_UPgCFFjT2_0(.dout(w_dff_A_cas8e2kd0_0),.din(w_dff_A_UPgCFFjT2_0),.clk(gclk));
	jdff dff_A_cas8e2kd0_0(.dout(G752),.din(w_dff_A_cas8e2kd0_0),.clk(gclk));
	jdff dff_A_olIlU6Rz9_2(.dout(w_dff_A_KgngQVaW4_0),.din(w_dff_A_olIlU6Rz9_2),.clk(gclk));
	jdff dff_A_KgngQVaW4_0(.dout(w_dff_A_zy7EuiiC8_0),.din(w_dff_A_KgngQVaW4_0),.clk(gclk));
	jdff dff_A_zy7EuiiC8_0(.dout(w_dff_A_2VAYShV77_0),.din(w_dff_A_zy7EuiiC8_0),.clk(gclk));
	jdff dff_A_2VAYShV77_0(.dout(w_dff_A_sHQIN9RV8_0),.din(w_dff_A_2VAYShV77_0),.clk(gclk));
	jdff dff_A_sHQIN9RV8_0(.dout(w_dff_A_YfEFb6rC7_0),.din(w_dff_A_sHQIN9RV8_0),.clk(gclk));
	jdff dff_A_YfEFb6rC7_0(.dout(w_dff_A_8hvyRWUh6_0),.din(w_dff_A_YfEFb6rC7_0),.clk(gclk));
	jdff dff_A_8hvyRWUh6_0(.dout(w_dff_A_ziAl6mkq0_0),.din(w_dff_A_8hvyRWUh6_0),.clk(gclk));
	jdff dff_A_ziAl6mkq0_0(.dout(w_dff_A_ZdHL2U0N9_0),.din(w_dff_A_ziAl6mkq0_0),.clk(gclk));
	jdff dff_A_ZdHL2U0N9_0(.dout(w_dff_A_5qZihNdj5_0),.din(w_dff_A_ZdHL2U0N9_0),.clk(gclk));
	jdff dff_A_5qZihNdj5_0(.dout(G757),.din(w_dff_A_5qZihNdj5_0),.clk(gclk));
	jdff dff_A_4jmLlBEL6_2(.dout(w_dff_A_K7dGq1W42_0),.din(w_dff_A_4jmLlBEL6_2),.clk(gclk));
	jdff dff_A_K7dGq1W42_0(.dout(w_dff_A_78ErQpbl6_0),.din(w_dff_A_K7dGq1W42_0),.clk(gclk));
	jdff dff_A_78ErQpbl6_0(.dout(w_dff_A_oiP58vZN1_0),.din(w_dff_A_78ErQpbl6_0),.clk(gclk));
	jdff dff_A_oiP58vZN1_0(.dout(w_dff_A_MBacnCiC5_0),.din(w_dff_A_oiP58vZN1_0),.clk(gclk));
	jdff dff_A_MBacnCiC5_0(.dout(w_dff_A_TbjA9WKO4_0),.din(w_dff_A_MBacnCiC5_0),.clk(gclk));
	jdff dff_A_TbjA9WKO4_0(.dout(w_dff_A_bZcxRaf15_0),.din(w_dff_A_TbjA9WKO4_0),.clk(gclk));
	jdff dff_A_bZcxRaf15_0(.dout(w_dff_A_BTPkT3Ar5_0),.din(w_dff_A_bZcxRaf15_0),.clk(gclk));
	jdff dff_A_BTPkT3Ar5_0(.dout(w_dff_A_P5kiD42M5_0),.din(w_dff_A_BTPkT3Ar5_0),.clk(gclk));
	jdff dff_A_P5kiD42M5_0(.dout(w_dff_A_UVRF8aHg7_0),.din(w_dff_A_P5kiD42M5_0),.clk(gclk));
	jdff dff_A_UVRF8aHg7_0(.dout(w_dff_A_YA4PgFku5_0),.din(w_dff_A_UVRF8aHg7_0),.clk(gclk));
	jdff dff_A_YA4PgFku5_0(.dout(G762),.din(w_dff_A_YA4PgFku5_0),.clk(gclk));
	jdff dff_A_AoLkuKZ61_2(.dout(w_dff_A_ylw4dDrN6_0),.din(w_dff_A_AoLkuKZ61_2),.clk(gclk));
	jdff dff_A_ylw4dDrN6_0(.dout(w_dff_A_Xdd7ok6a8_0),.din(w_dff_A_ylw4dDrN6_0),.clk(gclk));
	jdff dff_A_Xdd7ok6a8_0(.dout(w_dff_A_54dByUgn2_0),.din(w_dff_A_Xdd7ok6a8_0),.clk(gclk));
	jdff dff_A_54dByUgn2_0(.dout(w_dff_A_wFhZF4Ua8_0),.din(w_dff_A_54dByUgn2_0),.clk(gclk));
	jdff dff_A_wFhZF4Ua8_0(.dout(w_dff_A_lFjcVmsP9_0),.din(w_dff_A_wFhZF4Ua8_0),.clk(gclk));
	jdff dff_A_lFjcVmsP9_0(.dout(w_dff_A_pG7puxD84_0),.din(w_dff_A_lFjcVmsP9_0),.clk(gclk));
	jdff dff_A_pG7puxD84_0(.dout(G787),.din(w_dff_A_pG7puxD84_0),.clk(gclk));
	jdff dff_A_YAvYkCbM4_2(.dout(w_dff_A_NP1UhJWR0_0),.din(w_dff_A_YAvYkCbM4_2),.clk(gclk));
	jdff dff_A_NP1UhJWR0_0(.dout(w_dff_A_xmFAMjXS1_0),.din(w_dff_A_NP1UhJWR0_0),.clk(gclk));
	jdff dff_A_xmFAMjXS1_0(.dout(w_dff_A_wl6vBbvG5_0),.din(w_dff_A_xmFAMjXS1_0),.clk(gclk));
	jdff dff_A_wl6vBbvG5_0(.dout(w_dff_A_n9OBKh7T0_0),.din(w_dff_A_wl6vBbvG5_0),.clk(gclk));
	jdff dff_A_n9OBKh7T0_0(.dout(w_dff_A_VYZunaUg1_0),.din(w_dff_A_n9OBKh7T0_0),.clk(gclk));
	jdff dff_A_VYZunaUg1_0(.dout(w_dff_A_KFNQHDik9_0),.din(w_dff_A_VYZunaUg1_0),.clk(gclk));
	jdff dff_A_KFNQHDik9_0(.dout(w_dff_A_UCB5aFk39_0),.din(w_dff_A_KFNQHDik9_0),.clk(gclk));
	jdff dff_A_UCB5aFk39_0(.dout(w_dff_A_HgVkLhSQ4_0),.din(w_dff_A_UCB5aFk39_0),.clk(gclk));
	jdff dff_A_HgVkLhSQ4_0(.dout(G792),.din(w_dff_A_HgVkLhSQ4_0),.clk(gclk));
	jdff dff_A_DSdWtge17_2(.dout(w_dff_A_OKCOEJBq8_0),.din(w_dff_A_DSdWtge17_2),.clk(gclk));
	jdff dff_A_OKCOEJBq8_0(.dout(w_dff_A_R4F0qpPw9_0),.din(w_dff_A_OKCOEJBq8_0),.clk(gclk));
	jdff dff_A_R4F0qpPw9_0(.dout(w_dff_A_MeOEPxwg2_0),.din(w_dff_A_R4F0qpPw9_0),.clk(gclk));
	jdff dff_A_MeOEPxwg2_0(.dout(w_dff_A_ldtHwkm14_0),.din(w_dff_A_MeOEPxwg2_0),.clk(gclk));
	jdff dff_A_ldtHwkm14_0(.dout(w_dff_A_BM0TILL55_0),.din(w_dff_A_ldtHwkm14_0),.clk(gclk));
	jdff dff_A_BM0TILL55_0(.dout(w_dff_A_09sC8z2F0_0),.din(w_dff_A_BM0TILL55_0),.clk(gclk));
	jdff dff_A_09sC8z2F0_0(.dout(w_dff_A_SEI4HRti9_0),.din(w_dff_A_09sC8z2F0_0),.clk(gclk));
	jdff dff_A_SEI4HRti9_0(.dout(w_dff_A_0KaDLOvR8_0),.din(w_dff_A_SEI4HRti9_0),.clk(gclk));
	jdff dff_A_0KaDLOvR8_0(.dout(w_dff_A_8z21HOci0_0),.din(w_dff_A_0KaDLOvR8_0),.clk(gclk));
	jdff dff_A_8z21HOci0_0(.dout(G797),.din(w_dff_A_8z21HOci0_0),.clk(gclk));
	jdff dff_A_8xMKGdES8_2(.dout(w_dff_A_AGXVRCXs4_0),.din(w_dff_A_8xMKGdES8_2),.clk(gclk));
	jdff dff_A_AGXVRCXs4_0(.dout(w_dff_A_nfZXKJYC6_0),.din(w_dff_A_AGXVRCXs4_0),.clk(gclk));
	jdff dff_A_nfZXKJYC6_0(.dout(w_dff_A_9iL3PPUR3_0),.din(w_dff_A_nfZXKJYC6_0),.clk(gclk));
	jdff dff_A_9iL3PPUR3_0(.dout(w_dff_A_phLtGnGA2_0),.din(w_dff_A_9iL3PPUR3_0),.clk(gclk));
	jdff dff_A_phLtGnGA2_0(.dout(w_dff_A_IL80sVEE0_0),.din(w_dff_A_phLtGnGA2_0),.clk(gclk));
	jdff dff_A_IL80sVEE0_0(.dout(w_dff_A_EIST3LLL7_0),.din(w_dff_A_IL80sVEE0_0),.clk(gclk));
	jdff dff_A_EIST3LLL7_0(.dout(w_dff_A_QMTxobcq3_0),.din(w_dff_A_EIST3LLL7_0),.clk(gclk));
	jdff dff_A_QMTxobcq3_0(.dout(w_dff_A_8Cu09kgp5_0),.din(w_dff_A_QMTxobcq3_0),.clk(gclk));
	jdff dff_A_8Cu09kgp5_0(.dout(w_dff_A_sJsXddFe9_0),.din(w_dff_A_8Cu09kgp5_0),.clk(gclk));
	jdff dff_A_sJsXddFe9_0(.dout(w_dff_A_gtRm3smp8_0),.din(w_dff_A_sJsXddFe9_0),.clk(gclk));
	jdff dff_A_gtRm3smp8_0(.dout(G802),.din(w_dff_A_gtRm3smp8_0),.clk(gclk));
	jdff dff_A_vpF12bp06_2(.dout(w_dff_A_94yHG7RF0_0),.din(w_dff_A_vpF12bp06_2),.clk(gclk));
	jdff dff_A_94yHG7RF0_0(.dout(w_dff_A_hzy0GCaL9_0),.din(w_dff_A_94yHG7RF0_0),.clk(gclk));
	jdff dff_A_hzy0GCaL9_0(.dout(w_dff_A_o1lTLpvY3_0),.din(w_dff_A_hzy0GCaL9_0),.clk(gclk));
	jdff dff_A_o1lTLpvY3_0(.dout(w_dff_A_N8RH7KoB4_0),.din(w_dff_A_o1lTLpvY3_0),.clk(gclk));
	jdff dff_A_N8RH7KoB4_0(.dout(w_dff_A_ptN1hIfg7_0),.din(w_dff_A_N8RH7KoB4_0),.clk(gclk));
	jdff dff_A_ptN1hIfg7_0(.dout(G642),.din(w_dff_A_ptN1hIfg7_0),.clk(gclk));
	jdff dff_A_f74DpKmn1_2(.dout(w_dff_A_stUBsX9Y3_0),.din(w_dff_A_f74DpKmn1_2),.clk(gclk));
	jdff dff_A_stUBsX9Y3_0(.dout(w_dff_A_B0VYz8H04_0),.din(w_dff_A_stUBsX9Y3_0),.clk(gclk));
	jdff dff_A_B0VYz8H04_0(.dout(w_dff_A_61KOlwvS7_0),.din(w_dff_A_B0VYz8H04_0),.clk(gclk));
	jdff dff_A_61KOlwvS7_0(.dout(w_dff_A_oMX9Z7mC0_0),.din(w_dff_A_61KOlwvS7_0),.clk(gclk));
	jdff dff_A_oMX9Z7mC0_0(.dout(w_dff_A_l9EQlrUr5_0),.din(w_dff_A_oMX9Z7mC0_0),.clk(gclk));
	jdff dff_A_l9EQlrUr5_0(.dout(w_dff_A_CndLagRN3_0),.din(w_dff_A_l9EQlrUr5_0),.clk(gclk));
	jdff dff_A_CndLagRN3_0(.dout(w_dff_A_suQ69fZk6_0),.din(w_dff_A_CndLagRN3_0),.clk(gclk));
	jdff dff_A_suQ69fZk6_0(.dout(w_dff_A_saarCmgb1_0),.din(w_dff_A_suQ69fZk6_0),.clk(gclk));
	jdff dff_A_saarCmgb1_0(.dout(w_dff_A_ZeBcVuVL1_0),.din(w_dff_A_saarCmgb1_0),.clk(gclk));
	jdff dff_A_ZeBcVuVL1_0(.dout(G664),.din(w_dff_A_ZeBcVuVL1_0),.clk(gclk));
	jdff dff_A_E82YkNP98_2(.dout(w_dff_A_NiXddwT25_0),.din(w_dff_A_E82YkNP98_2),.clk(gclk));
	jdff dff_A_NiXddwT25_0(.dout(w_dff_A_yHork1d10_0),.din(w_dff_A_NiXddwT25_0),.clk(gclk));
	jdff dff_A_yHork1d10_0(.dout(w_dff_A_bDHBIp0h1_0),.din(w_dff_A_yHork1d10_0),.clk(gclk));
	jdff dff_A_bDHBIp0h1_0(.dout(w_dff_A_bMyTcRzc2_0),.din(w_dff_A_bDHBIp0h1_0),.clk(gclk));
	jdff dff_A_bMyTcRzc2_0(.dout(w_dff_A_XSMtrSdO4_0),.din(w_dff_A_bMyTcRzc2_0),.clk(gclk));
	jdff dff_A_XSMtrSdO4_0(.dout(w_dff_A_IKk72nFo2_0),.din(w_dff_A_XSMtrSdO4_0),.clk(gclk));
	jdff dff_A_IKk72nFo2_0(.dout(w_dff_A_IzPlc5I72_0),.din(w_dff_A_IKk72nFo2_0),.clk(gclk));
	jdff dff_A_IzPlc5I72_0(.dout(w_dff_A_R2TdcyTO5_0),.din(w_dff_A_IzPlc5I72_0),.clk(gclk));
	jdff dff_A_R2TdcyTO5_0(.dout(G667),.din(w_dff_A_R2TdcyTO5_0),.clk(gclk));
	jdff dff_A_IXXnVHd24_2(.dout(w_dff_A_JWVPPvce1_0),.din(w_dff_A_IXXnVHd24_2),.clk(gclk));
	jdff dff_A_JWVPPvce1_0(.dout(w_dff_A_7qBRIocz2_0),.din(w_dff_A_JWVPPvce1_0),.clk(gclk));
	jdff dff_A_7qBRIocz2_0(.dout(w_dff_A_N08CUWNV6_0),.din(w_dff_A_7qBRIocz2_0),.clk(gclk));
	jdff dff_A_N08CUWNV6_0(.dout(w_dff_A_ayycVdQ24_0),.din(w_dff_A_N08CUWNV6_0),.clk(gclk));
	jdff dff_A_ayycVdQ24_0(.dout(w_dff_A_wCdQqJ2e4_0),.din(w_dff_A_ayycVdQ24_0),.clk(gclk));
	jdff dff_A_wCdQqJ2e4_0(.dout(w_dff_A_VdDQx32P4_0),.din(w_dff_A_wCdQqJ2e4_0),.clk(gclk));
	jdff dff_A_VdDQx32P4_0(.dout(w_dff_A_hUoNM79V4_0),.din(w_dff_A_VdDQx32P4_0),.clk(gclk));
	jdff dff_A_hUoNM79V4_0(.dout(G670),.din(w_dff_A_hUoNM79V4_0),.clk(gclk));
	jdff dff_A_D1HnF7sc8_2(.dout(w_dff_A_uDhLzK2H6_0),.din(w_dff_A_D1HnF7sc8_2),.clk(gclk));
	jdff dff_A_uDhLzK2H6_0(.dout(w_dff_A_zpmEnjqy5_0),.din(w_dff_A_uDhLzK2H6_0),.clk(gclk));
	jdff dff_A_zpmEnjqy5_0(.dout(w_dff_A_NgIu6MSO1_0),.din(w_dff_A_zpmEnjqy5_0),.clk(gclk));
	jdff dff_A_NgIu6MSO1_0(.dout(w_dff_A_BjGsCpof1_0),.din(w_dff_A_NgIu6MSO1_0),.clk(gclk));
	jdff dff_A_BjGsCpof1_0(.dout(w_dff_A_Y8mCYuq03_0),.din(w_dff_A_BjGsCpof1_0),.clk(gclk));
	jdff dff_A_Y8mCYuq03_0(.dout(G676),.din(w_dff_A_Y8mCYuq03_0),.clk(gclk));
	jdff dff_A_DeuY0TwH2_2(.dout(w_dff_A_uYU0wR1Y6_0),.din(w_dff_A_DeuY0TwH2_2),.clk(gclk));
	jdff dff_A_uYU0wR1Y6_0(.dout(w_dff_A_2U6ZxD2y9_0),.din(w_dff_A_uYU0wR1Y6_0),.clk(gclk));
	jdff dff_A_2U6ZxD2y9_0(.dout(w_dff_A_zXGG6A3l3_0),.din(w_dff_A_2U6ZxD2y9_0),.clk(gclk));
	jdff dff_A_zXGG6A3l3_0(.dout(w_dff_A_LVO1btpO5_0),.din(w_dff_A_zXGG6A3l3_0),.clk(gclk));
	jdff dff_A_LVO1btpO5_0(.dout(w_dff_A_uSXEqGXQ0_0),.din(w_dff_A_LVO1btpO5_0),.clk(gclk));
	jdff dff_A_uSXEqGXQ0_0(.dout(w_dff_A_P6Iyrhfh6_0),.din(w_dff_A_uSXEqGXQ0_0),.clk(gclk));
	jdff dff_A_P6Iyrhfh6_0(.dout(w_dff_A_GBhKIpXW7_0),.din(w_dff_A_P6Iyrhfh6_0),.clk(gclk));
	jdff dff_A_GBhKIpXW7_0(.dout(w_dff_A_nFhCDl725_0),.din(w_dff_A_GBhKIpXW7_0),.clk(gclk));
	jdff dff_A_nFhCDl725_0(.dout(w_dff_A_SW2DSLHN4_0),.din(w_dff_A_nFhCDl725_0),.clk(gclk));
	jdff dff_A_SW2DSLHN4_0(.dout(G696),.din(w_dff_A_SW2DSLHN4_0),.clk(gclk));
	jdff dff_A_tZp0S1964_2(.dout(w_dff_A_yXpZtutY9_0),.din(w_dff_A_tZp0S1964_2),.clk(gclk));
	jdff dff_A_yXpZtutY9_0(.dout(w_dff_A_phIhrlIT6_0),.din(w_dff_A_yXpZtutY9_0),.clk(gclk));
	jdff dff_A_phIhrlIT6_0(.dout(w_dff_A_dIoFMkvd0_0),.din(w_dff_A_phIhrlIT6_0),.clk(gclk));
	jdff dff_A_dIoFMkvd0_0(.dout(w_dff_A_ovASpoot4_0),.din(w_dff_A_dIoFMkvd0_0),.clk(gclk));
	jdff dff_A_ovASpoot4_0(.dout(w_dff_A_Jv8ZzEsr9_0),.din(w_dff_A_ovASpoot4_0),.clk(gclk));
	jdff dff_A_Jv8ZzEsr9_0(.dout(w_dff_A_OdjIXAnE5_0),.din(w_dff_A_Jv8ZzEsr9_0),.clk(gclk));
	jdff dff_A_OdjIXAnE5_0(.dout(w_dff_A_4U8VAeQc6_0),.din(w_dff_A_OdjIXAnE5_0),.clk(gclk));
	jdff dff_A_4U8VAeQc6_0(.dout(w_dff_A_rLkYxBE65_0),.din(w_dff_A_4U8VAeQc6_0),.clk(gclk));
	jdff dff_A_rLkYxBE65_0(.dout(G699),.din(w_dff_A_rLkYxBE65_0),.clk(gclk));
	jdff dff_A_zqQOhykr8_2(.dout(w_dff_A_RNMnEmSD7_0),.din(w_dff_A_zqQOhykr8_2),.clk(gclk));
	jdff dff_A_RNMnEmSD7_0(.dout(w_dff_A_eBa1twq74_0),.din(w_dff_A_RNMnEmSD7_0),.clk(gclk));
	jdff dff_A_eBa1twq74_0(.dout(w_dff_A_LpVFuWwL7_0),.din(w_dff_A_eBa1twq74_0),.clk(gclk));
	jdff dff_A_LpVFuWwL7_0(.dout(w_dff_A_rvi8Gjiq1_0),.din(w_dff_A_LpVFuWwL7_0),.clk(gclk));
	jdff dff_A_rvi8Gjiq1_0(.dout(w_dff_A_KhMthFUg3_0),.din(w_dff_A_rvi8Gjiq1_0),.clk(gclk));
	jdff dff_A_KhMthFUg3_0(.dout(w_dff_A_edT1prM79_0),.din(w_dff_A_KhMthFUg3_0),.clk(gclk));
	jdff dff_A_edT1prM79_0(.dout(w_dff_A_xKM4KbzX0_0),.din(w_dff_A_edT1prM79_0),.clk(gclk));
	jdff dff_A_xKM4KbzX0_0(.dout(G702),.din(w_dff_A_xKM4KbzX0_0),.clk(gclk));
	jdff dff_A_YI0eKhC97_2(.dout(w_dff_A_ggvozNz20_0),.din(w_dff_A_YI0eKhC97_2),.clk(gclk));
	jdff dff_A_ggvozNz20_0(.dout(w_dff_A_Fxtp3UOU7_0),.din(w_dff_A_ggvozNz20_0),.clk(gclk));
	jdff dff_A_Fxtp3UOU7_0(.dout(w_dff_A_gNweMcxI6_0),.din(w_dff_A_Fxtp3UOU7_0),.clk(gclk));
	jdff dff_A_gNweMcxI6_0(.dout(w_dff_A_0MkrORxv9_0),.din(w_dff_A_gNweMcxI6_0),.clk(gclk));
	jdff dff_A_0MkrORxv9_0(.dout(G818),.din(w_dff_A_0MkrORxv9_0),.clk(gclk));
	jdff dff_A_Yu4al2p14_2(.dout(w_dff_A_h1v9vGOI7_0),.din(w_dff_A_Yu4al2p14_2),.clk(gclk));
	jdff dff_A_h1v9vGOI7_0(.dout(w_dff_A_UUWrqDDP6_0),.din(w_dff_A_h1v9vGOI7_0),.clk(gclk));
	jdff dff_A_UUWrqDDP6_0(.dout(w_dff_A_URLnBkPd3_0),.din(w_dff_A_UUWrqDDP6_0),.clk(gclk));
	jdff dff_A_URLnBkPd3_0(.dout(w_dff_A_8OqOhb8R9_0),.din(w_dff_A_URLnBkPd3_0),.clk(gclk));
	jdff dff_A_8OqOhb8R9_0(.dout(w_dff_A_XuJHswCl0_0),.din(w_dff_A_8OqOhb8R9_0),.clk(gclk));
	jdff dff_A_XuJHswCl0_0(.dout(w_dff_A_lSebnpja3_0),.din(w_dff_A_XuJHswCl0_0),.clk(gclk));
	jdff dff_A_lSebnpja3_0(.dout(w_dff_A_274ycebk5_0),.din(w_dff_A_lSebnpja3_0),.clk(gclk));
	jdff dff_A_274ycebk5_0(.dout(w_dff_A_mUdzZVc44_0),.din(w_dff_A_274ycebk5_0),.clk(gclk));
	jdff dff_A_mUdzZVc44_0(.dout(G813),.din(w_dff_A_mUdzZVc44_0),.clk(gclk));
	jdff dff_A_F0NuwJLN0_1(.dout(w_dff_A_pFZOshJI0_0),.din(w_dff_A_F0NuwJLN0_1),.clk(gclk));
	jdff dff_A_pFZOshJI0_0(.dout(w_dff_A_Gzq185nm1_0),.din(w_dff_A_pFZOshJI0_0),.clk(gclk));
	jdff dff_A_Gzq185nm1_0(.dout(w_dff_A_60ocbiJO4_0),.din(w_dff_A_Gzq185nm1_0),.clk(gclk));
	jdff dff_A_60ocbiJO4_0(.dout(w_dff_A_fF6WKln45_0),.din(w_dff_A_60ocbiJO4_0),.clk(gclk));
	jdff dff_A_fF6WKln45_0(.dout(G824),.din(w_dff_A_fF6WKln45_0),.clk(gclk));
	jdff dff_A_eohpnt6F6_1(.dout(w_dff_A_YGmloTLo6_0),.din(w_dff_A_eohpnt6F6_1),.clk(gclk));
	jdff dff_A_YGmloTLo6_0(.dout(w_dff_A_AcAIj35K0_0),.din(w_dff_A_YGmloTLo6_0),.clk(gclk));
	jdff dff_A_AcAIj35K0_0(.dout(w_dff_A_g2g6DWCU6_0),.din(w_dff_A_AcAIj35K0_0),.clk(gclk));
	jdff dff_A_g2g6DWCU6_0(.dout(w_dff_A_G04pAWMR5_0),.din(w_dff_A_g2g6DWCU6_0),.clk(gclk));
	jdff dff_A_G04pAWMR5_0(.dout(w_dff_A_YjWHI2wT6_0),.din(w_dff_A_G04pAWMR5_0),.clk(gclk));
	jdff dff_A_YjWHI2wT6_0(.dout(w_dff_A_X6pQOWnC1_0),.din(w_dff_A_YjWHI2wT6_0),.clk(gclk));
	jdff dff_A_X6pQOWnC1_0(.dout(w_dff_A_vCiBwh1v3_0),.din(w_dff_A_X6pQOWnC1_0),.clk(gclk));
	jdff dff_A_vCiBwh1v3_0(.dout(G826),.din(w_dff_A_vCiBwh1v3_0),.clk(gclk));
	jdff dff_A_0qERABzF8_1(.dout(w_dff_A_uoxTgMsL9_0),.din(w_dff_A_0qERABzF8_1),.clk(gclk));
	jdff dff_A_uoxTgMsL9_0(.dout(w_dff_A_qzccYyi69_0),.din(w_dff_A_uoxTgMsL9_0),.clk(gclk));
	jdff dff_A_qzccYyi69_0(.dout(w_dff_A_cN1iB1Up1_0),.din(w_dff_A_qzccYyi69_0),.clk(gclk));
	jdff dff_A_cN1iB1Up1_0(.dout(w_dff_A_fiZoD7uK1_0),.din(w_dff_A_cN1iB1Up1_0),.clk(gclk));
	jdff dff_A_fiZoD7uK1_0(.dout(w_dff_A_BdgTRnEU4_0),.din(w_dff_A_fiZoD7uK1_0),.clk(gclk));
	jdff dff_A_BdgTRnEU4_0(.dout(w_dff_A_h5oOv5FZ8_0),.din(w_dff_A_BdgTRnEU4_0),.clk(gclk));
	jdff dff_A_h5oOv5FZ8_0(.dout(w_dff_A_be7i5FF67_0),.din(w_dff_A_h5oOv5FZ8_0),.clk(gclk));
	jdff dff_A_be7i5FF67_0(.dout(G828),.din(w_dff_A_be7i5FF67_0),.clk(gclk));
	jdff dff_A_ouuG4aRI7_1(.dout(w_dff_A_YE0QG9OJ6_0),.din(w_dff_A_ouuG4aRI7_1),.clk(gclk));
	jdff dff_A_YE0QG9OJ6_0(.dout(w_dff_A_idd1QvNh1_0),.din(w_dff_A_YE0QG9OJ6_0),.clk(gclk));
	jdff dff_A_idd1QvNh1_0(.dout(w_dff_A_2nJ8TReo9_0),.din(w_dff_A_idd1QvNh1_0),.clk(gclk));
	jdff dff_A_2nJ8TReo9_0(.dout(w_dff_A_CP5Ezoe12_0),.din(w_dff_A_2nJ8TReo9_0),.clk(gclk));
	jdff dff_A_CP5Ezoe12_0(.dout(w_dff_A_xdhtc1bk9_0),.din(w_dff_A_CP5Ezoe12_0),.clk(gclk));
	jdff dff_A_xdhtc1bk9_0(.dout(w_dff_A_cjnk1i2V4_0),.din(w_dff_A_xdhtc1bk9_0),.clk(gclk));
	jdff dff_A_cjnk1i2V4_0(.dout(w_dff_A_K6l5DGdU5_0),.din(w_dff_A_cjnk1i2V4_0),.clk(gclk));
	jdff dff_A_K6l5DGdU5_0(.dout(w_dff_A_XKSW6wSY4_0),.din(w_dff_A_K6l5DGdU5_0),.clk(gclk));
	jdff dff_A_XKSW6wSY4_0(.dout(G830),.din(w_dff_A_XKSW6wSY4_0),.clk(gclk));
	jdff dff_A_YmBmEb0r2_2(.dout(w_dff_A_9CSwpaIN3_0),.din(w_dff_A_YmBmEb0r2_2),.clk(gclk));
	jdff dff_A_9CSwpaIN3_0(.dout(w_dff_A_bBtz4Z1h2_0),.din(w_dff_A_9CSwpaIN3_0),.clk(gclk));
	jdff dff_A_bBtz4Z1h2_0(.dout(w_dff_A_9f2imN564_0),.din(w_dff_A_bBtz4Z1h2_0),.clk(gclk));
	jdff dff_A_9f2imN564_0(.dout(w_dff_A_6ng2kMVn3_0),.din(w_dff_A_9f2imN564_0),.clk(gclk));
	jdff dff_A_6ng2kMVn3_0(.dout(w_dff_A_JlYr2jNi4_0),.din(w_dff_A_6ng2kMVn3_0),.clk(gclk));
	jdff dff_A_JlYr2jNi4_0(.dout(w_dff_A_FwuVeJOo5_0),.din(w_dff_A_JlYr2jNi4_0),.clk(gclk));
	jdff dff_A_FwuVeJOo5_0(.dout(w_dff_A_znqiFMAL6_0),.din(w_dff_A_FwuVeJOo5_0),.clk(gclk));
	jdff dff_A_znqiFMAL6_0(.dout(w_dff_A_twxvD3j61_0),.din(w_dff_A_znqiFMAL6_0),.clk(gclk));
	jdff dff_A_twxvD3j61_0(.dout(w_dff_A_WNTOuDZt5_0),.din(w_dff_A_twxvD3j61_0),.clk(gclk));
	jdff dff_A_WNTOuDZt5_0(.dout(w_dff_A_kMvYQVCE4_0),.din(w_dff_A_WNTOuDZt5_0),.clk(gclk));
	jdff dff_A_kMvYQVCE4_0(.dout(w_dff_A_WtxT0LXO4_0),.din(w_dff_A_kMvYQVCE4_0),.clk(gclk));
	jdff dff_A_WtxT0LXO4_0(.dout(w_dff_A_qSKMrMZx9_0),.din(w_dff_A_WtxT0LXO4_0),.clk(gclk));
	jdff dff_A_qSKMrMZx9_0(.dout(w_dff_A_T9Ik5eot6_0),.din(w_dff_A_qSKMrMZx9_0),.clk(gclk));
	jdff dff_A_T9Ik5eot6_0(.dout(w_dff_A_udz9AGVI8_0),.din(w_dff_A_T9Ik5eot6_0),.clk(gclk));
	jdff dff_A_udz9AGVI8_0(.dout(w_dff_A_vKV8Xpt58_0),.din(w_dff_A_udz9AGVI8_0),.clk(gclk));
	jdff dff_A_vKV8Xpt58_0(.dout(G854),.din(w_dff_A_vKV8Xpt58_0),.clk(gclk));
	jdff dff_A_61pVhAxr4_1(.dout(w_dff_A_seXWpN1q0_0),.din(w_dff_A_61pVhAxr4_1),.clk(gclk));
	jdff dff_A_seXWpN1q0_0(.dout(w_dff_A_GpPQJ5n18_0),.din(w_dff_A_seXWpN1q0_0),.clk(gclk));
	jdff dff_A_GpPQJ5n18_0(.dout(w_dff_A_clNs3gR33_0),.din(w_dff_A_GpPQJ5n18_0),.clk(gclk));
	jdff dff_A_clNs3gR33_0(.dout(G863),.din(w_dff_A_clNs3gR33_0),.clk(gclk));
	jdff dff_A_TCYtEEkG3_1(.dout(w_dff_A_FPGbjeBh2_0),.din(w_dff_A_TCYtEEkG3_1),.clk(gclk));
	jdff dff_A_FPGbjeBh2_0(.dout(w_dff_A_uqdmkj5g6_0),.din(w_dff_A_FPGbjeBh2_0),.clk(gclk));
	jdff dff_A_uqdmkj5g6_0(.dout(w_dff_A_M0ScsGu73_0),.din(w_dff_A_uqdmkj5g6_0),.clk(gclk));
	jdff dff_A_M0ScsGu73_0(.dout(w_dff_A_4rUlnZbF1_0),.din(w_dff_A_M0ScsGu73_0),.clk(gclk));
	jdff dff_A_4rUlnZbF1_0(.dout(G865),.din(w_dff_A_4rUlnZbF1_0),.clk(gclk));
	jdff dff_A_gLMnYhGz8_1(.dout(w_dff_A_kpCeFwp51_0),.din(w_dff_A_gLMnYhGz8_1),.clk(gclk));
	jdff dff_A_kpCeFwp51_0(.dout(w_dff_A_nx0MMVWJ4_0),.din(w_dff_A_kpCeFwp51_0),.clk(gclk));
	jdff dff_A_nx0MMVWJ4_0(.dout(w_dff_A_KdvHlEDf7_0),.din(w_dff_A_nx0MMVWJ4_0),.clk(gclk));
	jdff dff_A_KdvHlEDf7_0(.dout(w_dff_A_1Yh8oYJL3_0),.din(w_dff_A_KdvHlEDf7_0),.clk(gclk));
	jdff dff_A_1Yh8oYJL3_0(.dout(w_dff_A_5vABDvfk0_0),.din(w_dff_A_1Yh8oYJL3_0),.clk(gclk));
	jdff dff_A_5vABDvfk0_0(.dout(w_dff_A_LThrxDie4_0),.din(w_dff_A_5vABDvfk0_0),.clk(gclk));
	jdff dff_A_LThrxDie4_0(.dout(G867),.din(w_dff_A_LThrxDie4_0),.clk(gclk));
	jdff dff_A_p0X5p3Tl8_1(.dout(w_dff_A_NfrbBAt62_0),.din(w_dff_A_p0X5p3Tl8_1),.clk(gclk));
	jdff dff_A_NfrbBAt62_0(.dout(w_dff_A_XwmGzCL66_0),.din(w_dff_A_NfrbBAt62_0),.clk(gclk));
	jdff dff_A_XwmGzCL66_0(.dout(w_dff_A_SIzjbgeo5_0),.din(w_dff_A_XwmGzCL66_0),.clk(gclk));
	jdff dff_A_SIzjbgeo5_0(.dout(w_dff_A_swZFf9zW1_0),.din(w_dff_A_SIzjbgeo5_0),.clk(gclk));
	jdff dff_A_swZFf9zW1_0(.dout(w_dff_A_H9dev3Yc7_0),.din(w_dff_A_swZFf9zW1_0),.clk(gclk));
	jdff dff_A_H9dev3Yc7_0(.dout(w_dff_A_Z5Z00TpU1_0),.din(w_dff_A_H9dev3Yc7_0),.clk(gclk));
	jdff dff_A_Z5Z00TpU1_0(.dout(w_dff_A_TkidTaBr5_0),.din(w_dff_A_Z5Z00TpU1_0),.clk(gclk));
	jdff dff_A_TkidTaBr5_0(.dout(G869),.din(w_dff_A_TkidTaBr5_0),.clk(gclk));
	jdff dff_A_NjJ1rGZa7_2(.dout(w_dff_A_iV3hby8N7_0),.din(w_dff_A_NjJ1rGZa7_2),.clk(gclk));
	jdff dff_A_iV3hby8N7_0(.dout(w_dff_A_pcos2Awu2_0),.din(w_dff_A_iV3hby8N7_0),.clk(gclk));
	jdff dff_A_pcos2Awu2_0(.dout(G712),.din(w_dff_A_pcos2Awu2_0),.clk(gclk));
	jdff dff_A_AebEAUfu6_2(.dout(w_dff_A_CeuSNheH4_0),.din(w_dff_A_AebEAUfu6_2),.clk(gclk));
	jdff dff_A_CeuSNheH4_0(.dout(w_dff_A_PqBZ0Zbl1_0),.din(w_dff_A_CeuSNheH4_0),.clk(gclk));
	jdff dff_A_PqBZ0Zbl1_0(.dout(G727),.din(w_dff_A_PqBZ0Zbl1_0),.clk(gclk));
	jdff dff_A_tP90ihO79_2(.dout(w_dff_A_qiwq2d6T7_0),.din(w_dff_A_tP90ihO79_2),.clk(gclk));
	jdff dff_A_qiwq2d6T7_0(.dout(w_dff_A_MO6P1RqA3_0),.din(w_dff_A_qiwq2d6T7_0),.clk(gclk));
	jdff dff_A_MO6P1RqA3_0(.dout(w_dff_A_PP9HAOUA6_0),.din(w_dff_A_MO6P1RqA3_0),.clk(gclk));
	jdff dff_A_PP9HAOUA6_0(.dout(G732),.din(w_dff_A_PP9HAOUA6_0),.clk(gclk));
	jdff dff_A_4CRHhEj26_2(.dout(w_dff_A_bJHdQplT0_0),.din(w_dff_A_4CRHhEj26_2),.clk(gclk));
	jdff dff_A_bJHdQplT0_0(.dout(w_dff_A_NGh9qX0l8_0),.din(w_dff_A_bJHdQplT0_0),.clk(gclk));
	jdff dff_A_NGh9qX0l8_0(.dout(w_dff_A_Ko8nmzGj4_0),.din(w_dff_A_NGh9qX0l8_0),.clk(gclk));
	jdff dff_A_Ko8nmzGj4_0(.dout(G737),.din(w_dff_A_Ko8nmzGj4_0),.clk(gclk));
	jdff dff_A_7Y0fh7EU0_2(.dout(w_dff_A_1whWSXqV6_0),.din(w_dff_A_7Y0fh7EU0_2),.clk(gclk));
	jdff dff_A_1whWSXqV6_0(.dout(w_dff_A_VQ8RYErW9_0),.din(w_dff_A_1whWSXqV6_0),.clk(gclk));
	jdff dff_A_VQ8RYErW9_0(.dout(w_dff_A_glMeisTk3_0),.din(w_dff_A_VQ8RYErW9_0),.clk(gclk));
	jdff dff_A_glMeisTk3_0(.dout(w_dff_A_QI885KOz2_0),.din(w_dff_A_glMeisTk3_0),.clk(gclk));
	jdff dff_A_QI885KOz2_0(.dout(G742),.din(w_dff_A_QI885KOz2_0),.clk(gclk));
	jdff dff_A_rFepXOn66_2(.dout(w_dff_A_IyhwQnPo8_0),.din(w_dff_A_rFepXOn66_2),.clk(gclk));
	jdff dff_A_IyhwQnPo8_0(.dout(w_dff_A_NIgJUmOK0_0),.din(w_dff_A_IyhwQnPo8_0),.clk(gclk));
	jdff dff_A_NIgJUmOK0_0(.dout(w_dff_A_HRJtcXab0_0),.din(w_dff_A_NIgJUmOK0_0),.clk(gclk));
	jdff dff_A_HRJtcXab0_0(.dout(G772),.din(w_dff_A_HRJtcXab0_0),.clk(gclk));
	jdff dff_A_WBcazqRS7_2(.dout(w_dff_A_17Zn9pqn1_0),.din(w_dff_A_WBcazqRS7_2),.clk(gclk));
	jdff dff_A_17Zn9pqn1_0(.dout(w_dff_A_aV5rwXLd1_0),.din(w_dff_A_17Zn9pqn1_0),.clk(gclk));
	jdff dff_A_aV5rwXLd1_0(.dout(w_dff_A_8Lwqji8D4_0),.din(w_dff_A_aV5rwXLd1_0),.clk(gclk));
	jdff dff_A_8Lwqji8D4_0(.dout(G777),.din(w_dff_A_8Lwqji8D4_0),.clk(gclk));
	jdff dff_A_d2B7YkhN0_2(.dout(w_dff_A_EGtU07CN5_0),.din(w_dff_A_d2B7YkhN0_2),.clk(gclk));
	jdff dff_A_EGtU07CN5_0(.dout(w_dff_A_FC8nWnbz8_0),.din(w_dff_A_EGtU07CN5_0),.clk(gclk));
	jdff dff_A_FC8nWnbz8_0(.dout(w_dff_A_F4ap0ghy6_0),.din(w_dff_A_FC8nWnbz8_0),.clk(gclk));
	jdff dff_A_F4ap0ghy6_0(.dout(w_dff_A_CmABijxt0_0),.din(w_dff_A_F4ap0ghy6_0),.clk(gclk));
	jdff dff_A_CmABijxt0_0(.dout(G782),.din(w_dff_A_CmABijxt0_0),.clk(gclk));
	jdff dff_A_7YR1FAlA0_2(.dout(w_dff_A_qekfAvYc7_0),.din(w_dff_A_7YR1FAlA0_2),.clk(gclk));
	jdff dff_A_qekfAvYc7_0(.dout(w_dff_A_lnddDsbh6_0),.din(w_dff_A_qekfAvYc7_0),.clk(gclk));
	jdff dff_A_lnddDsbh6_0(.dout(w_dff_A_dAjtFB3P0_0),.din(w_dff_A_lnddDsbh6_0),.clk(gclk));
	jdff dff_A_dAjtFB3P0_0(.dout(G645),.din(w_dff_A_dAjtFB3P0_0),.clk(gclk));
	jdff dff_A_2lBg0wOi0_2(.dout(w_dff_A_HaWR7sXJ9_0),.din(w_dff_A_2lBg0wOi0_2),.clk(gclk));
	jdff dff_A_HaWR7sXJ9_0(.dout(w_dff_A_kddjHfwT8_0),.din(w_dff_A_HaWR7sXJ9_0),.clk(gclk));
	jdff dff_A_kddjHfwT8_0(.dout(G648),.din(w_dff_A_kddjHfwT8_0),.clk(gclk));
	jdff dff_A_hz6kOtRe3_2(.dout(w_dff_A_cKpcwRpm3_0),.din(w_dff_A_hz6kOtRe3_2),.clk(gclk));
	jdff dff_A_cKpcwRpm3_0(.dout(w_dff_A_xdlkBVQ79_0),.din(w_dff_A_cKpcwRpm3_0),.clk(gclk));
	jdff dff_A_xdlkBVQ79_0(.dout(G651),.din(w_dff_A_xdlkBVQ79_0),.clk(gclk));
	jdff dff_A_RrQzvuqd9_2(.dout(w_dff_A_ij4W11Rm5_0),.din(w_dff_A_RrQzvuqd9_2),.clk(gclk));
	jdff dff_A_ij4W11Rm5_0(.dout(G654),.din(w_dff_A_ij4W11Rm5_0),.clk(gclk));
	jdff dff_A_0wj4FSAV3_2(.dout(w_dff_A_D5XrwMvF1_0),.din(w_dff_A_0wj4FSAV3_2),.clk(gclk));
	jdff dff_A_D5XrwMvF1_0(.dout(w_dff_A_fwAv4NU81_0),.din(w_dff_A_D5XrwMvF1_0),.clk(gclk));
	jdff dff_A_fwAv4NU81_0(.dout(w_dff_A_8iQwItBN6_0),.din(w_dff_A_fwAv4NU81_0),.clk(gclk));
	jdff dff_A_8iQwItBN6_0(.dout(G679),.din(w_dff_A_8iQwItBN6_0),.clk(gclk));
	jdff dff_A_YzzF2G7s5_2(.dout(w_dff_A_pvim20DF8_0),.din(w_dff_A_YzzF2G7s5_2),.clk(gclk));
	jdff dff_A_pvim20DF8_0(.dout(w_dff_A_H80Avglf3_0),.din(w_dff_A_pvim20DF8_0),.clk(gclk));
	jdff dff_A_H80Avglf3_0(.dout(G682),.din(w_dff_A_H80Avglf3_0),.clk(gclk));
	jdff dff_A_o0JBYaTp4_2(.dout(w_dff_A_Hr8xD5Kc0_0),.din(w_dff_A_o0JBYaTp4_2),.clk(gclk));
	jdff dff_A_Hr8xD5Kc0_0(.dout(w_dff_A_MF5afOLJ9_0),.din(w_dff_A_Hr8xD5Kc0_0),.clk(gclk));
	jdff dff_A_MF5afOLJ9_0(.dout(G685),.din(w_dff_A_MF5afOLJ9_0),.clk(gclk));
	jdff dff_A_S3yRiD3O3_2(.dout(w_dff_A_vtmMt5Mp6_0),.din(w_dff_A_S3yRiD3O3_2),.clk(gclk));
	jdff dff_A_vtmMt5Mp6_0(.dout(G688),.din(w_dff_A_vtmMt5Mp6_0),.clk(gclk));
	jdff dff_A_WDxtKaJz2_2(.dout(w_dff_A_V6m1J4yy1_0),.din(w_dff_A_WDxtKaJz2_2),.clk(gclk));
	jdff dff_A_V6m1J4yy1_0(.dout(w_dff_A_r0HmbdrS9_0),.din(w_dff_A_V6m1J4yy1_0),.clk(gclk));
	jdff dff_A_r0HmbdrS9_0(.dout(w_dff_A_78VkBBwL2_0),.din(w_dff_A_r0HmbdrS9_0),.clk(gclk));
	jdff dff_A_78VkBBwL2_0(.dout(G843),.din(w_dff_A_78VkBBwL2_0),.clk(gclk));
	jdff dff_A_73tBNL023_2(.dout(w_dff_A_cWNtw4yV7_0),.din(w_dff_A_73tBNL023_2),.clk(gclk));
	jdff dff_A_cWNtw4yV7_0(.dout(w_dff_A_XE5T6Wwp1_0),.din(w_dff_A_cWNtw4yV7_0),.clk(gclk));
	jdff dff_A_XE5T6Wwp1_0(.dout(w_dff_A_WMXgV8dg7_0),.din(w_dff_A_XE5T6Wwp1_0),.clk(gclk));
	jdff dff_A_WMXgV8dg7_0(.dout(G882),.din(w_dff_A_WMXgV8dg7_0),.clk(gclk));
	jdff dff_A_hMdQYkwo2_2(.dout(G767),.din(w_dff_A_hMdQYkwo2_2),.clk(gclk));
	jdff dff_A_IsWFdUh62_2(.dout(G807),.din(w_dff_A_IsWFdUh62_2),.clk(gclk));
endmodule

