/*

c6288:
	jxor: 446
	jspl: 940
	jspl3: 260
	jnot: 330
	jdff: 8448
	jand: 683
	jor: 331

Summary:
	jxor: 446
	jspl: 940
	jspl3: 260
	jnot: 330
	jdff: 8448
	jand: 683
	jor: 331
*/

module c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G1gat_1;
	wire[2:0] w_G1gat_2;
	wire[2:0] w_G1gat_3;
	wire[2:0] w_G1gat_4;
	wire[2:0] w_G1gat_5;
	wire[2:0] w_G1gat_6;
	wire[1:0] w_G1gat_7;
	wire[2:0] w_G18gat_0;
	wire[2:0] w_G18gat_1;
	wire[2:0] w_G18gat_2;
	wire[2:0] w_G18gat_3;
	wire[2:0] w_G18gat_4;
	wire[2:0] w_G18gat_5;
	wire[2:0] w_G18gat_6;
	wire[2:0] w_G18gat_7;
	wire[2:0] w_G35gat_0;
	wire[2:0] w_G35gat_1;
	wire[2:0] w_G35gat_2;
	wire[2:0] w_G35gat_3;
	wire[2:0] w_G35gat_4;
	wire[2:0] w_G35gat_5;
	wire[2:0] w_G35gat_6;
	wire[2:0] w_G35gat_7;
	wire[2:0] w_G52gat_0;
	wire[2:0] w_G52gat_1;
	wire[2:0] w_G52gat_2;
	wire[2:0] w_G52gat_3;
	wire[2:0] w_G52gat_4;
	wire[2:0] w_G52gat_5;
	wire[2:0] w_G52gat_6;
	wire[2:0] w_G52gat_7;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G69gat_1;
	wire[2:0] w_G69gat_2;
	wire[2:0] w_G69gat_3;
	wire[2:0] w_G69gat_4;
	wire[2:0] w_G69gat_5;
	wire[2:0] w_G69gat_6;
	wire[1:0] w_G69gat_7;
	wire[2:0] w_G86gat_0;
	wire[2:0] w_G86gat_1;
	wire[2:0] w_G86gat_2;
	wire[2:0] w_G86gat_3;
	wire[2:0] w_G86gat_4;
	wire[2:0] w_G86gat_5;
	wire[2:0] w_G86gat_6;
	wire[1:0] w_G86gat_7;
	wire[2:0] w_G103gat_0;
	wire[2:0] w_G103gat_1;
	wire[2:0] w_G103gat_2;
	wire[2:0] w_G103gat_3;
	wire[2:0] w_G103gat_4;
	wire[2:0] w_G103gat_5;
	wire[2:0] w_G103gat_6;
	wire[1:0] w_G103gat_7;
	wire[2:0] w_G120gat_0;
	wire[2:0] w_G120gat_1;
	wire[2:0] w_G120gat_2;
	wire[2:0] w_G120gat_3;
	wire[2:0] w_G120gat_4;
	wire[2:0] w_G120gat_5;
	wire[2:0] w_G120gat_6;
	wire[1:0] w_G120gat_7;
	wire[2:0] w_G137gat_0;
	wire[2:0] w_G137gat_1;
	wire[2:0] w_G137gat_2;
	wire[2:0] w_G137gat_3;
	wire[2:0] w_G137gat_4;
	wire[2:0] w_G137gat_5;
	wire[2:0] w_G137gat_6;
	wire[1:0] w_G137gat_7;
	wire[2:0] w_G154gat_0;
	wire[2:0] w_G154gat_1;
	wire[2:0] w_G154gat_2;
	wire[2:0] w_G154gat_3;
	wire[2:0] w_G154gat_4;
	wire[2:0] w_G154gat_5;
	wire[2:0] w_G154gat_6;
	wire[1:0] w_G154gat_7;
	wire[2:0] w_G171gat_0;
	wire[2:0] w_G171gat_1;
	wire[2:0] w_G171gat_2;
	wire[2:0] w_G171gat_3;
	wire[2:0] w_G171gat_4;
	wire[2:0] w_G171gat_5;
	wire[2:0] w_G171gat_6;
	wire[1:0] w_G171gat_7;
	wire[2:0] w_G188gat_0;
	wire[2:0] w_G188gat_1;
	wire[2:0] w_G188gat_2;
	wire[2:0] w_G188gat_3;
	wire[2:0] w_G188gat_4;
	wire[2:0] w_G188gat_5;
	wire[2:0] w_G188gat_6;
	wire[1:0] w_G188gat_7;
	wire[2:0] w_G205gat_0;
	wire[2:0] w_G205gat_1;
	wire[2:0] w_G205gat_2;
	wire[2:0] w_G205gat_3;
	wire[2:0] w_G205gat_4;
	wire[2:0] w_G205gat_5;
	wire[2:0] w_G205gat_6;
	wire[1:0] w_G205gat_7;
	wire[2:0] w_G222gat_0;
	wire[2:0] w_G222gat_1;
	wire[2:0] w_G222gat_2;
	wire[2:0] w_G222gat_3;
	wire[2:0] w_G222gat_4;
	wire[2:0] w_G222gat_5;
	wire[2:0] w_G222gat_6;
	wire[1:0] w_G222gat_7;
	wire[2:0] w_G239gat_0;
	wire[2:0] w_G239gat_1;
	wire[2:0] w_G239gat_2;
	wire[2:0] w_G239gat_3;
	wire[2:0] w_G239gat_4;
	wire[2:0] w_G239gat_5;
	wire[2:0] w_G239gat_6;
	wire[1:0] w_G239gat_7;
	wire[2:0] w_G256gat_0;
	wire[2:0] w_G256gat_1;
	wire[2:0] w_G256gat_2;
	wire[2:0] w_G256gat_3;
	wire[2:0] w_G256gat_4;
	wire[2:0] w_G256gat_5;
	wire[2:0] w_G256gat_6;
	wire[1:0] w_G256gat_7;
	wire[2:0] w_G273gat_0;
	wire[2:0] w_G273gat_1;
	wire[2:0] w_G273gat_2;
	wire[2:0] w_G273gat_3;
	wire[2:0] w_G273gat_4;
	wire[2:0] w_G273gat_5;
	wire[2:0] w_G273gat_6;
	wire[2:0] w_G273gat_7;
	wire[2:0] w_G290gat_0;
	wire[2:0] w_G290gat_1;
	wire[2:0] w_G290gat_2;
	wire[2:0] w_G290gat_3;
	wire[2:0] w_G290gat_4;
	wire[2:0] w_G290gat_5;
	wire[2:0] w_G290gat_6;
	wire[2:0] w_G290gat_7;
	wire[2:0] w_G307gat_0;
	wire[2:0] w_G307gat_1;
	wire[2:0] w_G307gat_2;
	wire[2:0] w_G307gat_3;
	wire[2:0] w_G307gat_4;
	wire[2:0] w_G307gat_5;
	wire[2:0] w_G307gat_6;
	wire[2:0] w_G307gat_7;
	wire[2:0] w_G324gat_0;
	wire[2:0] w_G324gat_1;
	wire[2:0] w_G324gat_2;
	wire[2:0] w_G324gat_3;
	wire[2:0] w_G324gat_4;
	wire[2:0] w_G324gat_5;
	wire[2:0] w_G324gat_6;
	wire[1:0] w_G324gat_7;
	wire[2:0] w_G341gat_0;
	wire[2:0] w_G341gat_1;
	wire[2:0] w_G341gat_2;
	wire[2:0] w_G341gat_3;
	wire[2:0] w_G341gat_4;
	wire[2:0] w_G341gat_5;
	wire[2:0] w_G341gat_6;
	wire[1:0] w_G341gat_7;
	wire[2:0] w_G358gat_0;
	wire[2:0] w_G358gat_1;
	wire[2:0] w_G358gat_2;
	wire[2:0] w_G358gat_3;
	wire[2:0] w_G358gat_4;
	wire[2:0] w_G358gat_5;
	wire[2:0] w_G358gat_6;
	wire[1:0] w_G358gat_7;
	wire[2:0] w_G375gat_0;
	wire[2:0] w_G375gat_1;
	wire[2:0] w_G375gat_2;
	wire[2:0] w_G375gat_3;
	wire[2:0] w_G375gat_4;
	wire[2:0] w_G375gat_5;
	wire[2:0] w_G375gat_6;
	wire[1:0] w_G375gat_7;
	wire[2:0] w_G392gat_0;
	wire[2:0] w_G392gat_1;
	wire[2:0] w_G392gat_2;
	wire[2:0] w_G392gat_3;
	wire[2:0] w_G392gat_4;
	wire[2:0] w_G392gat_5;
	wire[2:0] w_G392gat_6;
	wire[1:0] w_G392gat_7;
	wire[2:0] w_G409gat_0;
	wire[2:0] w_G409gat_1;
	wire[2:0] w_G409gat_2;
	wire[2:0] w_G409gat_3;
	wire[2:0] w_G409gat_4;
	wire[2:0] w_G409gat_5;
	wire[2:0] w_G409gat_6;
	wire[1:0] w_G409gat_7;
	wire[2:0] w_G426gat_0;
	wire[2:0] w_G426gat_1;
	wire[2:0] w_G426gat_2;
	wire[2:0] w_G426gat_3;
	wire[2:0] w_G426gat_4;
	wire[2:0] w_G426gat_5;
	wire[2:0] w_G426gat_6;
	wire[1:0] w_G426gat_7;
	wire[2:0] w_G443gat_0;
	wire[2:0] w_G443gat_1;
	wire[2:0] w_G443gat_2;
	wire[2:0] w_G443gat_3;
	wire[2:0] w_G443gat_4;
	wire[2:0] w_G443gat_5;
	wire[2:0] w_G443gat_6;
	wire[1:0] w_G443gat_7;
	wire[2:0] w_G460gat_0;
	wire[2:0] w_G460gat_1;
	wire[2:0] w_G460gat_2;
	wire[2:0] w_G460gat_3;
	wire[2:0] w_G460gat_4;
	wire[2:0] w_G460gat_5;
	wire[2:0] w_G460gat_6;
	wire[1:0] w_G460gat_7;
	wire[2:0] w_G477gat_0;
	wire[2:0] w_G477gat_1;
	wire[2:0] w_G477gat_2;
	wire[2:0] w_G477gat_3;
	wire[2:0] w_G477gat_4;
	wire[2:0] w_G477gat_5;
	wire[2:0] w_G477gat_6;
	wire[1:0] w_G477gat_7;
	wire[2:0] w_G494gat_0;
	wire[2:0] w_G494gat_1;
	wire[2:0] w_G494gat_2;
	wire[2:0] w_G494gat_3;
	wire[2:0] w_G494gat_4;
	wire[2:0] w_G494gat_5;
	wire[2:0] w_G494gat_6;
	wire[1:0] w_G494gat_7;
	wire[2:0] w_G511gat_0;
	wire[2:0] w_G511gat_1;
	wire[2:0] w_G511gat_2;
	wire[2:0] w_G511gat_3;
	wire[2:0] w_G511gat_4;
	wire[2:0] w_G511gat_5;
	wire[2:0] w_G511gat_6;
	wire[1:0] w_G511gat_7;
	wire[2:0] w_G528gat_0;
	wire[2:0] w_G528gat_1;
	wire[2:0] w_G528gat_2;
	wire[2:0] w_G528gat_3;
	wire[2:0] w_G528gat_4;
	wire[2:0] w_G528gat_5;
	wire[2:0] w_G528gat_6;
	wire[1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire[1:0] w_n65_0;
	wire[1:0] w_n69_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n72_0;
	wire[1:0] w_n75_0;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[1:0] w_n81_0;
	wire[2:0] w_n82_0;
	wire[1:0] w_n82_1;
	wire[1:0] w_n84_0;
	wire[1:0] w_n85_0;
	wire[1:0] w_n87_0;
	wire[1:0] w_n89_0;
	wire[1:0] w_n93_0;
	wire[1:0] w_n94_0;
	wire[1:0] w_n96_0;
	wire[1:0] w_n99_0;
	wire[2:0] w_n100_0;
	wire[1:0] w_n100_1;
	wire[2:0] w_n101_0;
	wire[1:0] w_n103_0;
	wire[1:0] w_n104_0;
	wire[1:0] w_n107_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n110_0;
	wire[1:0] w_n115_0;
	wire[1:0] w_n116_0;
	wire[2:0] w_n126_0;
	wire[1:0] w_n128_0;
	wire[1:0] w_n129_0;
	wire[1:0] w_n130_0;
	wire[1:0] w_n131_0;
	wire[2:0] w_n132_0;
	wire[2:0] w_n133_0;
	wire[1:0] w_n138_0;
	wire[1:0] w_n139_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n142_0;
	wire[1:0] w_n143_0;
	wire[1:0] w_n145_0;
	wire[1:0] w_n150_0;
	wire[1:0] w_n151_0;
	wire[2:0] w_n156_0;
	wire[1:0] w_n158_0;
	wire[1:0] w_n163_0;
	wire[1:0] w_n165_0;
	wire[1:0] w_n166_0;
	wire[1:0] w_n168_0;
	wire[2:0] w_n169_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n172_0;
	wire[1:0] w_n174_0;
	wire[1:0] w_n175_0;
	wire[1:0] w_n176_0;
	wire[1:0] w_n177_0;
	wire[1:0] w_n178_0;
	wire[1:0] w_n180_0;
	wire[1:0] w_n181_0;
	wire[1:0] w_n183_0;
	wire[1:0] w_n188_0;
	wire[1:0] w_n189_0;
	wire[2:0] w_n194_0;
	wire[1:0] w_n196_0;
	wire[1:0] w_n199_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n207_0;
	wire[1:0] w_n209_0;
	wire[2:0] w_n210_0;
	wire[1:0] w_n210_1;
	wire[1:0] w_n213_0;
	wire[1:0] w_n215_0;
	wire[1:0] w_n216_0;
	wire[1:0] w_n217_0;
	wire[1:0] w_n218_0;
	wire[1:0] w_n219_0;
	wire[1:0] w_n220_0;
	wire[1:0] w_n221_0;
	wire[1:0] w_n223_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n226_0;
	wire[1:0] w_n231_0;
	wire[1:0] w_n232_0;
	wire[2:0] w_n237_0;
	wire[1:0] w_n239_0;
	wire[1:0] w_n242_0;
	wire[1:0] w_n244_0;
	wire[1:0] w_n247_0;
	wire[1:0] w_n249_0;
	wire[1:0] w_n252_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n255_0;
	wire[1:0] w_n257_0;
	wire[2:0] w_n258_0;
	wire[1:0] w_n259_0;
	wire[1:0] w_n261_0;
	wire[1:0] w_n264_0;
	wire[1:0] w_n265_0;
	wire[1:0] w_n266_0;
	wire[1:0] w_n267_0;
	wire[1:0] w_n268_0;
	wire[1:0] w_n269_0;
	wire[1:0] w_n270_0;
	wire[1:0] w_n271_0;
	wire[1:0] w_n272_0;
	wire[1:0] w_n274_0;
	wire[1:0] w_n275_0;
	wire[1:0] w_n277_0;
	wire[1:0] w_n282_0;
	wire[1:0] w_n283_0;
	wire[2:0] w_n288_0;
	wire[1:0] w_n290_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n295_0;
	wire[1:0] w_n298_0;
	wire[1:0] w_n300_0;
	wire[1:0] w_n303_0;
	wire[1:0] w_n305_0;
	wire[1:0] w_n308_0;
	wire[1:0] w_n310_0;
	wire[1:0] w_n311_0;
	wire[1:0] w_n313_0;
	wire[2:0] w_n314_0;
	wire[1:0] w_n315_0;
	wire[1:0] w_n317_0;
	wire[1:0] w_n320_0;
	wire[1:0] w_n321_0;
	wire[1:0] w_n322_0;
	wire[1:0] w_n323_0;
	wire[1:0] w_n324_0;
	wire[1:0] w_n325_0;
	wire[1:0] w_n326_0;
	wire[1:0] w_n327_0;
	wire[1:0] w_n328_0;
	wire[1:0] w_n329_0;
	wire[1:0] w_n330_0;
	wire[1:0] w_n332_0;
	wire[1:0] w_n333_0;
	wire[1:0] w_n335_0;
	wire[1:0] w_n340_0;
	wire[1:0] w_n341_0;
	wire[2:0] w_n346_0;
	wire[1:0] w_n348_0;
	wire[1:0] w_n351_0;
	wire[1:0] w_n353_0;
	wire[1:0] w_n356_0;
	wire[1:0] w_n358_0;
	wire[1:0] w_n361_0;
	wire[1:0] w_n363_0;
	wire[1:0] w_n366_0;
	wire[1:0] w_n368_0;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n373_0;
	wire[1:0] w_n375_0;
	wire[2:0] w_n376_0;
	wire[1:0] w_n377_0;
	wire[1:0] w_n380_0;
	wire[1:0] w_n382_0;
	wire[1:0] w_n383_0;
	wire[1:0] w_n384_0;
	wire[1:0] w_n385_0;
	wire[1:0] w_n386_0;
	wire[1:0] w_n387_0;
	wire[1:0] w_n388_0;
	wire[1:0] w_n389_0;
	wire[1:0] w_n390_0;
	wire[1:0] w_n391_0;
	wire[1:0] w_n392_0;
	wire[1:0] w_n393_0;
	wire[1:0] w_n394_0;
	wire[1:0] w_n396_0;
	wire[1:0] w_n397_0;
	wire[1:0] w_n399_0;
	wire[1:0] w_n404_0;
	wire[1:0] w_n405_0;
	wire[2:0] w_n410_0;
	wire[1:0] w_n412_0;
	wire[1:0] w_n415_0;
	wire[1:0] w_n417_0;
	wire[1:0] w_n420_0;
	wire[1:0] w_n422_0;
	wire[1:0] w_n425_0;
	wire[1:0] w_n427_0;
	wire[1:0] w_n430_0;
	wire[1:0] w_n432_0;
	wire[1:0] w_n435_0;
	wire[1:0] w_n437_0;
	wire[1:0] w_n441_0;
	wire[1:0] w_n442_0;
	wire[1:0] w_n443_0;
	wire[1:0] w_n445_0;
	wire[2:0] w_n446_0;
	wire[1:0] w_n447_0;
	wire[1:0] w_n450_0;
	wire[1:0] w_n452_0;
	wire[1:0] w_n453_0;
	wire[1:0] w_n454_0;
	wire[1:0] w_n455_0;
	wire[1:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[1:0] w_n458_0;
	wire[1:0] w_n459_0;
	wire[1:0] w_n460_0;
	wire[1:0] w_n461_0;
	wire[1:0] w_n462_0;
	wire[1:0] w_n463_0;
	wire[1:0] w_n464_0;
	wire[1:0] w_n465_0;
	wire[1:0] w_n466_0;
	wire[1:0] w_n468_0;
	wire[1:0] w_n469_0;
	wire[1:0] w_n471_0;
	wire[1:0] w_n476_0;
	wire[1:0] w_n477_0;
	wire[2:0] w_n482_0;
	wire[1:0] w_n484_0;
	wire[1:0] w_n487_0;
	wire[1:0] w_n489_0;
	wire[1:0] w_n492_0;
	wire[1:0] w_n494_0;
	wire[1:0] w_n497_0;
	wire[1:0] w_n499_0;
	wire[1:0] w_n502_0;
	wire[1:0] w_n504_0;
	wire[1:0] w_n507_0;
	wire[1:0] w_n509_0;
	wire[1:0] w_n512_0;
	wire[1:0] w_n514_0;
	wire[1:0] w_n518_0;
	wire[1:0] w_n519_0;
	wire[1:0] w_n520_0;
	wire[1:0] w_n522_0;
	wire[2:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n527_0;
	wire[1:0] w_n529_0;
	wire[1:0] w_n530_0;
	wire[1:0] w_n531_0;
	wire[1:0] w_n532_0;
	wire[1:0] w_n533_0;
	wire[1:0] w_n534_0;
	wire[1:0] w_n535_0;
	wire[1:0] w_n536_0;
	wire[1:0] w_n537_0;
	wire[1:0] w_n538_0;
	wire[1:0] w_n539_0;
	wire[1:0] w_n540_0;
	wire[1:0] w_n541_0;
	wire[1:0] w_n542_0;
	wire[1:0] w_n543_0;
	wire[1:0] w_n544_0;
	wire[1:0] w_n545_0;
	wire[1:0] w_n547_0;
	wire[1:0] w_n548_0;
	wire[1:0] w_n550_0;
	wire[1:0] w_n555_0;
	wire[1:0] w_n556_0;
	wire[2:0] w_n561_0;
	wire[1:0] w_n563_0;
	wire[1:0] w_n566_0;
	wire[1:0] w_n568_0;
	wire[1:0] w_n571_0;
	wire[1:0] w_n573_0;
	wire[1:0] w_n576_0;
	wire[1:0] w_n578_0;
	wire[1:0] w_n581_0;
	wire[1:0] w_n583_0;
	wire[1:0] w_n586_0;
	wire[1:0] w_n588_0;
	wire[1:0] w_n591_0;
	wire[1:0] w_n593_0;
	wire[1:0] w_n596_0;
	wire[1:0] w_n598_0;
	wire[1:0] w_n602_0;
	wire[1:0] w_n603_0;
	wire[1:0] w_n604_0;
	wire[1:0] w_n606_0;
	wire[2:0] w_n607_0;
	wire[1:0] w_n608_0;
	wire[1:0] w_n611_0;
	wire[1:0] w_n613_0;
	wire[1:0] w_n614_0;
	wire[1:0] w_n615_0;
	wire[1:0] w_n616_0;
	wire[1:0] w_n617_0;
	wire[1:0] w_n618_0;
	wire[1:0] w_n619_0;
	wire[1:0] w_n620_0;
	wire[1:0] w_n621_0;
	wire[1:0] w_n622_0;
	wire[1:0] w_n623_0;
	wire[1:0] w_n624_0;
	wire[1:0] w_n625_0;
	wire[1:0] w_n626_0;
	wire[1:0] w_n627_0;
	wire[1:0] w_n628_0;
	wire[1:0] w_n629_0;
	wire[1:0] w_n630_0;
	wire[1:0] w_n631_0;
	wire[1:0] w_n633_0;
	wire[1:0] w_n634_0;
	wire[1:0] w_n636_0;
	wire[1:0] w_n641_0;
	wire[1:0] w_n642_0;
	wire[2:0] w_n647_0;
	wire[1:0] w_n649_0;
	wire[1:0] w_n652_0;
	wire[1:0] w_n654_0;
	wire[1:0] w_n657_0;
	wire[1:0] w_n659_0;
	wire[1:0] w_n662_0;
	wire[1:0] w_n664_0;
	wire[1:0] w_n667_0;
	wire[1:0] w_n669_0;
	wire[1:0] w_n672_0;
	wire[1:0] w_n674_0;
	wire[1:0] w_n677_0;
	wire[1:0] w_n679_0;
	wire[1:0] w_n682_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n693_0;
	wire[1:0] w_n694_0;
	wire[2:0] w_n695_0;
	wire[1:0] w_n697_0;
	wire[2:0] w_n698_0;
	wire[1:0] w_n699_0;
	wire[1:0] w_n702_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n705_0;
	wire[1:0] w_n706_0;
	wire[1:0] w_n707_0;
	wire[1:0] w_n708_0;
	wire[1:0] w_n709_0;
	wire[1:0] w_n710_0;
	wire[1:0] w_n711_0;
	wire[1:0] w_n712_0;
	wire[1:0] w_n713_0;
	wire[1:0] w_n714_0;
	wire[1:0] w_n715_0;
	wire[1:0] w_n716_0;
	wire[1:0] w_n717_0;
	wire[1:0] w_n718_0;
	wire[1:0] w_n719_0;
	wire[1:0] w_n720_0;
	wire[1:0] w_n721_0;
	wire[1:0] w_n722_0;
	wire[1:0] w_n723_0;
	wire[1:0] w_n724_0;
	wire[1:0] w_n726_0;
	wire[1:0] w_n727_0;
	wire[1:0] w_n729_0;
	wire[1:0] w_n734_0;
	wire[1:0] w_n735_0;
	wire[2:0] w_n740_0;
	wire[1:0] w_n742_0;
	wire[1:0] w_n745_0;
	wire[1:0] w_n747_0;
	wire[1:0] w_n750_0;
	wire[1:0] w_n752_0;
	wire[1:0] w_n755_0;
	wire[1:0] w_n757_0;
	wire[1:0] w_n760_0;
	wire[1:0] w_n762_0;
	wire[1:0] w_n765_0;
	wire[1:0] w_n767_0;
	wire[1:0] w_n770_0;
	wire[1:0] w_n772_0;
	wire[1:0] w_n775_0;
	wire[1:0] w_n777_0;
	wire[1:0] w_n780_0;
	wire[1:0] w_n782_0;
	wire[1:0] w_n785_0;
	wire[1:0] w_n787_0;
	wire[1:0] w_n791_0;
	wire[1:0] w_n792_0;
	wire[1:0] w_n793_0;
	wire[1:0] w_n795_0;
	wire[2:0] w_n797_0;
	wire[1:0] w_n800_0;
	wire[1:0] w_n802_0;
	wire[1:0] w_n803_0;
	wire[1:0] w_n804_0;
	wire[1:0] w_n805_0;
	wire[1:0] w_n806_0;
	wire[1:0] w_n807_0;
	wire[1:0] w_n808_0;
	wire[1:0] w_n809_0;
	wire[1:0] w_n810_0;
	wire[1:0] w_n811_0;
	wire[1:0] w_n812_0;
	wire[1:0] w_n813_0;
	wire[1:0] w_n814_0;
	wire[1:0] w_n815_0;
	wire[1:0] w_n816_0;
	wire[1:0] w_n817_0;
	wire[1:0] w_n818_0;
	wire[1:0] w_n819_0;
	wire[1:0] w_n820_0;
	wire[1:0] w_n821_0;
	wire[1:0] w_n822_0;
	wire[1:0] w_n823_0;
	wire[1:0] w_n824_0;
	wire[1:0] w_n826_0;
	wire[1:0] w_n827_0;
	wire[1:0] w_n829_0;
	wire[1:0] w_n834_0;
	wire[1:0] w_n835_0;
	wire[1:0] w_n839_0;
	wire[1:0] w_n840_0;
	wire[2:0] w_n844_0;
	wire[1:0] w_n846_0;
	wire[1:0] w_n849_0;
	wire[1:0] w_n851_0;
	wire[1:0] w_n854_0;
	wire[1:0] w_n856_0;
	wire[1:0] w_n859_0;
	wire[1:0] w_n861_0;
	wire[1:0] w_n864_0;
	wire[1:0] w_n866_0;
	wire[1:0] w_n869_0;
	wire[1:0] w_n871_0;
	wire[1:0] w_n874_0;
	wire[1:0] w_n876_0;
	wire[1:0] w_n879_0;
	wire[1:0] w_n881_0;
	wire[1:0] w_n884_0;
	wire[1:0] w_n886_0;
	wire[1:0] w_n889_0;
	wire[1:0] w_n891_0;
	wire[1:0] w_n895_0;
	wire[1:0] w_n896_0;
	wire[1:0] w_n897_0;
	wire[1:0] w_n898_0;
	wire[1:0] w_n901_0;
	wire[1:0] w_n903_0;
	wire[1:0] w_n906_0;
	wire[1:0] w_n907_0;
	wire[1:0] w_n908_0;
	wire[1:0] w_n909_0;
	wire[1:0] w_n910_0;
	wire[1:0] w_n911_0;
	wire[1:0] w_n912_0;
	wire[1:0] w_n913_0;
	wire[1:0] w_n914_0;
	wire[1:0] w_n915_0;
	wire[1:0] w_n916_0;
	wire[1:0] w_n917_0;
	wire[1:0] w_n918_0;
	wire[1:0] w_n919_0;
	wire[1:0] w_n920_0;
	wire[1:0] w_n921_0;
	wire[1:0] w_n922_0;
	wire[1:0] w_n923_0;
	wire[1:0] w_n924_0;
	wire[1:0] w_n925_0;
	wire[1:0] w_n926_0;
	wire[2:0] w_n927_0;
	wire[1:0] w_n929_0;
	wire[1:0] w_n930_0;
	wire[1:0] w_n931_0;
	wire[1:0] w_n932_0;
	wire[1:0] w_n937_0;
	wire[1:0] w_n938_0;
	wire[2:0] w_n942_0;
	wire[1:0] w_n943_0;
	wire[1:0] w_n949_0;
	wire[1:0] w_n951_0;
	wire[1:0] w_n954_0;
	wire[1:0] w_n956_0;
	wire[1:0] w_n959_0;
	wire[1:0] w_n961_0;
	wire[1:0] w_n964_0;
	wire[1:0] w_n966_0;
	wire[1:0] w_n969_0;
	wire[1:0] w_n971_0;
	wire[1:0] w_n974_0;
	wire[1:0] w_n976_0;
	wire[1:0] w_n979_0;
	wire[1:0] w_n981_0;
	wire[1:0] w_n984_0;
	wire[1:0] w_n986_0;
	wire[1:0] w_n989_0;
	wire[1:0] w_n991_0;
	wire[1:0] w_n994_0;
	wire[1:0] w_n996_0;
	wire[1:0] w_n999_0;
	wire[1:0] w_n1001_0;
	wire[1:0] w_n1005_0;
	wire[1:0] w_n1006_0;
	wire[1:0] w_n1008_0;
	wire[1:0] w_n1009_0;
	wire[1:0] w_n1010_0;
	wire[1:0] w_n1011_0;
	wire[1:0] w_n1012_0;
	wire[1:0] w_n1013_0;
	wire[1:0] w_n1014_0;
	wire[1:0] w_n1015_0;
	wire[1:0] w_n1016_0;
	wire[1:0] w_n1017_0;
	wire[1:0] w_n1018_0;
	wire[1:0] w_n1019_0;
	wire[1:0] w_n1020_0;
	wire[1:0] w_n1021_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1023_0;
	wire[1:0] w_n1024_0;
	wire[1:0] w_n1025_0;
	wire[1:0] w_n1026_0;
	wire[1:0] w_n1027_0;
	wire[1:0] w_n1028_0;
	wire[1:0] w_n1029_0;
	wire[1:0] w_n1030_0;
	wire[1:0] w_n1031_0;
	wire[1:0] w_n1032_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1034_0;
	wire[1:0] w_n1035_0;
	wire[1:0] w_n1037_0;
	wire[1:0] w_n1039_0;
	wire[1:0] w_n1043_0;
	wire[1:0] w_n1044_0;
	wire[1:0] w_n1048_0;
	wire[1:0] w_n1049_0;
	wire[1:0] w_n1052_0;
	wire[1:0] w_n1054_0;
	wire[1:0] w_n1057_0;
	wire[1:0] w_n1059_0;
	wire[1:0] w_n1062_0;
	wire[1:0] w_n1064_0;
	wire[1:0] w_n1067_0;
	wire[1:0] w_n1069_0;
	wire[1:0] w_n1072_0;
	wire[1:0] w_n1074_0;
	wire[1:0] w_n1077_0;
	wire[1:0] w_n1079_0;
	wire[1:0] w_n1082_0;
	wire[1:0] w_n1084_0;
	wire[1:0] w_n1087_0;
	wire[1:0] w_n1089_0;
	wire[1:0] w_n1092_0;
	wire[1:0] w_n1094_0;
	wire[1:0] w_n1097_0;
	wire[1:0] w_n1099_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1103_0;
	wire[1:0] w_n1109_0;
	wire[1:0] w_n1110_0;
	wire[1:0] w_n1114_0;
	wire[1:0] w_n1115_0;
	wire[1:0] w_n1116_0;
	wire[1:0] w_n1117_0;
	wire[1:0] w_n1118_0;
	wire[1:0] w_n1119_0;
	wire[1:0] w_n1120_0;
	wire[1:0] w_n1121_0;
	wire[1:0] w_n1122_0;
	wire[1:0] w_n1123_0;
	wire[1:0] w_n1124_0;
	wire[1:0] w_n1125_0;
	wire[1:0] w_n1126_0;
	wire[1:0] w_n1127_0;
	wire[1:0] w_n1128_0;
	wire[1:0] w_n1129_0;
	wire[1:0] w_n1130_0;
	wire[1:0] w_n1131_0;
	wire[1:0] w_n1132_0;
	wire[1:0] w_n1133_0;
	wire[1:0] w_n1134_0;
	wire[1:0] w_n1135_0;
	wire[1:0] w_n1137_0;
	wire[1:0] w_n1138_0;
	wire[1:0] w_n1139_0;
	wire[1:0] w_n1140_0;
	wire[1:0] w_n1141_0;
	wire[1:0] w_n1147_0;
	wire[1:0] w_n1151_0;
	wire[1:0] w_n1152_0;
	wire[1:0] w_n1156_0;
	wire[1:0] w_n1158_0;
	wire[1:0] w_n1161_0;
	wire[1:0] w_n1163_0;
	wire[1:0] w_n1166_0;
	wire[1:0] w_n1168_0;
	wire[1:0] w_n1171_0;
	wire[1:0] w_n1173_0;
	wire[1:0] w_n1176_0;
	wire[1:0] w_n1178_0;
	wire[1:0] w_n1181_0;
	wire[1:0] w_n1183_0;
	wire[1:0] w_n1186_0;
	wire[1:0] w_n1188_0;
	wire[1:0] w_n1191_0;
	wire[1:0] w_n1193_0;
	wire[1:0] w_n1196_0;
	wire[1:0] w_n1198_0;
	wire[1:0] w_n1201_0;
	wire[1:0] w_n1203_0;
	wire[1:0] w_n1206_0;
	wire[1:0] w_n1207_0;
	wire[1:0] w_n1208_0;
	wire[1:0] w_n1210_0;
	wire[1:0] w_n1212_0;
	wire[1:0] w_n1213_0;
	wire[1:0] w_n1214_0;
	wire[1:0] w_n1215_0;
	wire[1:0] w_n1216_0;
	wire[1:0] w_n1217_0;
	wire[1:0] w_n1218_0;
	wire[1:0] w_n1219_0;
	wire[1:0] w_n1220_0;
	wire[1:0] w_n1221_0;
	wire[1:0] w_n1222_0;
	wire[1:0] w_n1223_0;
	wire[1:0] w_n1224_0;
	wire[1:0] w_n1225_0;
	wire[1:0] w_n1226_0;
	wire[1:0] w_n1227_0;
	wire[1:0] w_n1228_0;
	wire[1:0] w_n1229_0;
	wire[1:0] w_n1230_0;
	wire[1:0] w_n1231_0;
	wire[1:0] w_n1232_0;
	wire[1:0] w_n1234_0;
	wire[1:0] w_n1236_0;
	wire[1:0] w_n1237_0;
	wire[1:0] w_n1238_0;
	wire[1:0] w_n1244_0;
	wire[1:0] w_n1247_0;
	wire[1:0] w_n1248_0;
	wire[1:0] w_n1251_0;
	wire[1:0] w_n1253_0;
	wire[1:0] w_n1256_0;
	wire[1:0] w_n1258_0;
	wire[1:0] w_n1261_0;
	wire[1:0] w_n1263_0;
	wire[1:0] w_n1266_0;
	wire[1:0] w_n1268_0;
	wire[1:0] w_n1271_0;
	wire[1:0] w_n1273_0;
	wire[1:0] w_n1276_0;
	wire[1:0] w_n1278_0;
	wire[1:0] w_n1281_0;
	wire[1:0] w_n1283_0;
	wire[1:0] w_n1286_0;
	wire[1:0] w_n1288_0;
	wire[1:0] w_n1291_0;
	wire[1:0] w_n1293_0;
	wire[1:0] w_n1296_0;
	wire[1:0] w_n1297_0;
	wire[1:0] w_n1298_0;
	wire[1:0] w_n1301_0;
	wire[1:0] w_n1303_0;
	wire[1:0] w_n1304_0;
	wire[1:0] w_n1305_0;
	wire[1:0] w_n1306_0;
	wire[1:0] w_n1307_0;
	wire[1:0] w_n1308_0;
	wire[1:0] w_n1309_0;
	wire[1:0] w_n1310_0;
	wire[1:0] w_n1311_0;
	wire[1:0] w_n1312_0;
	wire[1:0] w_n1313_0;
	wire[1:0] w_n1314_0;
	wire[1:0] w_n1315_0;
	wire[1:0] w_n1316_0;
	wire[1:0] w_n1317_0;
	wire[1:0] w_n1318_0;
	wire[1:0] w_n1319_0;
	wire[1:0] w_n1320_0;
	wire[1:0] w_n1321_0;
	wire[1:0] w_n1322_0;
	wire[1:0] w_n1324_0;
	wire[1:0] w_n1325_0;
	wire[1:0] w_n1326_0;
	wire[1:0] w_n1332_0;
	wire[1:0] w_n1337_0;
	wire[1:0] w_n1338_0;
	wire[1:0] w_n1341_0;
	wire[1:0] w_n1343_0;
	wire[1:0] w_n1346_0;
	wire[1:0] w_n1348_0;
	wire[1:0] w_n1351_0;
	wire[1:0] w_n1353_0;
	wire[1:0] w_n1356_0;
	wire[1:0] w_n1358_0;
	wire[1:0] w_n1361_0;
	wire[1:0] w_n1363_0;
	wire[1:0] w_n1366_0;
	wire[1:0] w_n1368_0;
	wire[1:0] w_n1371_0;
	wire[1:0] w_n1373_0;
	wire[1:0] w_n1376_0;
	wire[1:0] w_n1378_0;
	wire[1:0] w_n1381_0;
	wire[1:0] w_n1382_0;
	wire[1:0] w_n1383_0;
	wire[1:0] w_n1386_0;
	wire[1:0] w_n1388_0;
	wire[1:0] w_n1389_0;
	wire[1:0] w_n1390_0;
	wire[1:0] w_n1391_0;
	wire[1:0] w_n1392_0;
	wire[1:0] w_n1393_0;
	wire[1:0] w_n1394_0;
	wire[1:0] w_n1395_0;
	wire[1:0] w_n1396_0;
	wire[1:0] w_n1397_0;
	wire[1:0] w_n1398_0;
	wire[1:0] w_n1399_0;
	wire[1:0] w_n1400_0;
	wire[1:0] w_n1401_0;
	wire[1:0] w_n1402_0;
	wire[1:0] w_n1403_0;
	wire[1:0] w_n1404_0;
	wire[1:0] w_n1405_0;
	wire[1:0] w_n1407_0;
	wire[1:0] w_n1409_0;
	wire[1:0] w_n1410_0;
	wire[1:0] w_n1415_0;
	wire[1:0] w_n1420_0;
	wire[1:0] w_n1421_0;
	wire[1:0] w_n1424_0;
	wire[1:0] w_n1426_0;
	wire[1:0] w_n1429_0;
	wire[1:0] w_n1431_0;
	wire[1:0] w_n1434_0;
	wire[1:0] w_n1436_0;
	wire[1:0] w_n1439_0;
	wire[1:0] w_n1441_0;
	wire[1:0] w_n1444_0;
	wire[1:0] w_n1446_0;
	wire[1:0] w_n1449_0;
	wire[1:0] w_n1451_0;
	wire[1:0] w_n1454_0;
	wire[1:0] w_n1456_0;
	wire[1:0] w_n1459_0;
	wire[1:0] w_n1460_0;
	wire[1:0] w_n1461_0;
	wire[1:0] w_n1464_0;
	wire[1:0] w_n1466_0;
	wire[1:0] w_n1467_0;
	wire[1:0] w_n1468_0;
	wire[1:0] w_n1469_0;
	wire[1:0] w_n1470_0;
	wire[1:0] w_n1471_0;
	wire[1:0] w_n1472_0;
	wire[1:0] w_n1473_0;
	wire[1:0] w_n1474_0;
	wire[1:0] w_n1475_0;
	wire[1:0] w_n1476_0;
	wire[1:0] w_n1477_0;
	wire[1:0] w_n1478_0;
	wire[1:0] w_n1479_0;
	wire[1:0] w_n1480_0;
	wire[1:0] w_n1481_0;
	wire[1:0] w_n1483_0;
	wire[1:0] w_n1485_0;
	wire[1:0] w_n1486_0;
	wire[1:0] w_n1491_0;
	wire[1:0] w_n1496_0;
	wire[1:0] w_n1497_0;
	wire[1:0] w_n1500_0;
	wire[1:0] w_n1502_0;
	wire[1:0] w_n1505_0;
	wire[1:0] w_n1507_0;
	wire[1:0] w_n1510_0;
	wire[1:0] w_n1512_0;
	wire[1:0] w_n1515_0;
	wire[1:0] w_n1517_0;
	wire[1:0] w_n1520_0;
	wire[1:0] w_n1522_0;
	wire[1:0] w_n1525_0;
	wire[1:0] w_n1527_0;
	wire[1:0] w_n1530_0;
	wire[1:0] w_n1531_0;
	wire[1:0] w_n1532_0;
	wire[1:0] w_n1535_0;
	wire[1:0] w_n1537_0;
	wire[1:0] w_n1538_0;
	wire[1:0] w_n1539_0;
	wire[1:0] w_n1540_0;
	wire[1:0] w_n1541_0;
	wire[1:0] w_n1542_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1544_0;
	wire[1:0] w_n1545_0;
	wire[1:0] w_n1546_0;
	wire[1:0] w_n1547_0;
	wire[1:0] w_n1548_0;
	wire[1:0] w_n1549_0;
	wire[1:0] w_n1550_0;
	wire[1:0] w_n1552_0;
	wire[1:0] w_n1554_0;
	wire[1:0] w_n1555_0;
	wire[1:0] w_n1560_0;
	wire[1:0] w_n1565_0;
	wire[1:0] w_n1566_0;
	wire[1:0] w_n1569_0;
	wire[1:0] w_n1571_0;
	wire[1:0] w_n1574_0;
	wire[1:0] w_n1576_0;
	wire[1:0] w_n1579_0;
	wire[1:0] w_n1581_0;
	wire[1:0] w_n1584_0;
	wire[1:0] w_n1586_0;
	wire[1:0] w_n1589_0;
	wire[1:0] w_n1591_0;
	wire[1:0] w_n1594_0;
	wire[1:0] w_n1595_0;
	wire[1:0] w_n1596_0;
	wire[1:0] w_n1599_0;
	wire[1:0] w_n1601_0;
	wire[1:0] w_n1602_0;
	wire[1:0] w_n1603_0;
	wire[1:0] w_n1604_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1606_0;
	wire[1:0] w_n1607_0;
	wire[1:0] w_n1608_0;
	wire[1:0] w_n1609_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1611_0;
	wire[1:0] w_n1612_0;
	wire[1:0] w_n1614_0;
	wire[1:0] w_n1616_0;
	wire[1:0] w_n1617_0;
	wire[1:0] w_n1622_0;
	wire[1:0] w_n1627_0;
	wire[1:0] w_n1628_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1633_0;
	wire[1:0] w_n1636_0;
	wire[1:0] w_n1638_0;
	wire[1:0] w_n1641_0;
	wire[1:0] w_n1643_0;
	wire[1:0] w_n1646_0;
	wire[1:0] w_n1648_0;
	wire[1:0] w_n1651_0;
	wire[1:0] w_n1652_0;
	wire[1:0] w_n1653_0;
	wire[1:0] w_n1656_0;
	wire[1:0] w_n1658_0;
	wire[1:0] w_n1659_0;
	wire[1:0] w_n1660_0;
	wire[1:0] w_n1661_0;
	wire[1:0] w_n1662_0;
	wire[1:0] w_n1663_0;
	wire[1:0] w_n1664_0;
	wire[1:0] w_n1665_0;
	wire[1:0] w_n1666_0;
	wire[1:0] w_n1667_0;
	wire[1:0] w_n1669_0;
	wire[1:0] w_n1671_0;
	wire[1:0] w_n1672_0;
	wire[1:0] w_n1677_0;
	wire[1:0] w_n1682_0;
	wire[1:0] w_n1684_0;
	wire[1:0] w_n1687_0;
	wire[1:0] w_n1689_0;
	wire[1:0] w_n1692_0;
	wire[1:0] w_n1694_0;
	wire[1:0] w_n1697_0;
	wire[1:0] w_n1699_0;
	wire[1:0] w_n1702_0;
	wire[1:0] w_n1703_0;
	wire[1:0] w_n1704_0;
	wire[1:0] w_n1707_0;
	wire[1:0] w_n1709_0;
	wire[1:0] w_n1710_0;
	wire[1:0] w_n1711_0;
	wire[1:0] w_n1712_0;
	wire[1:0] w_n1713_0;
	wire[1:0] w_n1714_0;
	wire[1:0] w_n1715_0;
	wire[1:0] w_n1716_0;
	wire[1:0] w_n1717_0;
	wire[1:0] w_n1719_0;
	wire[1:0] w_n1720_0;
	wire[1:0] w_n1725_0;
	wire[1:0] w_n1728_0;
	wire[1:0] w_n1730_0;
	wire[1:0] w_n1733_0;
	wire[1:0] w_n1735_0;
	wire[1:0] w_n1738_0;
	wire[1:0] w_n1740_0;
	wire[1:0] w_n1743_0;
	wire[1:0] w_n1744_0;
	wire[1:0] w_n1745_0;
	wire[1:0] w_n1748_0;
	wire[1:0] w_n1750_0;
	wire[1:0] w_n1751_0;
	wire[1:0] w_n1752_0;
	wire[1:0] w_n1753_0;
	wire[1:0] w_n1754_0;
	wire[1:0] w_n1755_0;
	wire[1:0] w_n1756_0;
	wire[1:0] w_n1757_0;
	wire[1:0] w_n1758_0;
	wire[1:0] w_n1765_0;
	wire[1:0] w_n1768_0;
	wire[1:0] w_n1770_0;
	wire[1:0] w_n1773_0;
	wire[1:0] w_n1775_0;
	wire[1:0] w_n1778_0;
	wire[1:0] w_n1779_0;
	wire[1:0] w_n1780_0;
	wire[1:0] w_n1783_0;
	wire[1:0] w_n1785_0;
	wire[1:0] w_n1786_0;
	wire[1:0] w_n1787_0;
	wire[1:0] w_n1788_0;
	wire[1:0] w_n1789_0;
	wire[1:0] w_n1790_0;
	wire[1:0] w_n1791_0;
	wire[1:0] w_n1798_0;
	wire[1:0] w_n1801_0;
	wire[1:0] w_n1803_0;
	wire[1:0] w_n1806_0;
	wire[1:0] w_n1807_0;
	wire[1:0] w_n1808_0;
	wire[1:0] w_n1811_0;
	wire[1:0] w_n1813_0;
	wire[1:0] w_n1814_0;
	wire[1:0] w_n1815_0;
	wire[1:0] w_n1816_0;
	wire[1:0] w_n1817_0;
	wire[1:0] w_n1824_0;
	wire[1:0] w_n1827_0;
	wire[1:0] w_n1828_0;
	wire[1:0] w_n1829_0;
	wire[1:0] w_n1832_0;
	wire[1:0] w_n1834_0;
	wire[1:0] w_n1835_0;
	wire[1:0] w_n1836_0;
	wire[1:0] w_n1838_0;
	wire[1:0] w_n1841_0;
	wire[1:0] w_n1848_0;
	wire[1:0] w_n1849_0;
	wire w_dff_B_FlnRawTX7_1;
	wire w_dff_B_wCMHpDOi5_1;
	wire w_dff_B_sdJfy7uL5_1;
	wire w_dff_B_STxbppBs3_1;
	wire w_dff_B_HbMs7I9A8_1;
	wire w_dff_B_60O3SjDB7_1;
	wire w_dff_B_ERxjwXja7_1;
	wire w_dff_B_0F0VZf8u2_1;
	wire w_dff_B_Lr8oXvTq9_1;
	wire w_dff_B_ilYyFsgQ3_1;
	wire w_dff_B_4iotCQpn5_1;
	wire w_dff_B_Zp5c4yA99_1;
	wire w_dff_B_rRivL0kd8_1;
	wire w_dff_B_SJSr3X7k5_1;
	wire w_dff_B_VvhWuhwe8_1;
	wire w_dff_B_aSgInQzn5_1;
	wire w_dff_B_IIVETUCY5_1;
	wire w_dff_B_O86EOvnT3_1;
	wire w_dff_B_Gufbg2BB4_1;
	wire w_dff_B_zjxJOgeN3_1;
	wire w_dff_B_gl7VcSe70_1;
	wire w_dff_B_oWExCNQ75_1;
	wire w_dff_B_vtS2lXxj3_1;
	wire w_dff_B_UbgYM5jy7_1;
	wire w_dff_B_T2EdSbCF4_1;
	wire w_dff_B_G9KAKXTI4_1;
	wire w_dff_B_BCjl6DfE9_1;
	wire w_dff_B_shKcgyAq3_1;
	wire w_dff_B_1fo167qq5_1;
	wire w_dff_B_DsEquqky4_1;
	wire w_dff_B_Iw9Bbdmu3_1;
	wire w_dff_B_4593GmyZ5_1;
	wire w_dff_B_8BOnlKVH7_1;
	wire w_dff_B_9sJ4FH923_1;
	wire w_dff_B_nEJzxkY00_1;
	wire w_dff_B_6Q1zjGBA2_1;
	wire w_dff_B_sLWALcqO7_1;
	wire w_dff_B_VGKpUuhp3_1;
	wire w_dff_B_SXvicOZ97_1;
	wire w_dff_B_8nFYkbrA6_1;
	wire w_dff_B_brptCj5c0_1;
	wire w_dff_B_R31P1xF99_1;
	wire w_dff_B_5oPOPCIv2_1;
	wire w_dff_B_MKZEa4wR8_1;
	wire w_dff_B_DBHOqC0l8_1;
	wire w_dff_B_B3Z3reUi3_1;
	wire w_dff_B_Ak2Bm4ee3_1;
	wire w_dff_B_3F6TGqKX7_1;
	wire w_dff_B_9fUtzQSP0_1;
	wire w_dff_B_wDHTkjfr6_1;
	wire w_dff_B_YCIsNlDY6_1;
	wire w_dff_B_whqYXsbT0_1;
	wire w_dff_B_S96bL5oT8_1;
	wire w_dff_B_EaGbqYTL1_1;
	wire w_dff_B_PI3bVm1B4_1;
	wire w_dff_B_qqi9RPW07_1;
	wire w_dff_B_dzhTTeFT2_1;
	wire w_dff_B_CuLD6BCu9_1;
	wire w_dff_B_cLVzMxuz2_1;
	wire w_dff_B_B2XPbEAQ1_1;
	wire w_dff_B_uO8pLFjw1_1;
	wire w_dff_B_m5IUpABs2_1;
	wire w_dff_B_dmF44GG68_1;
	wire w_dff_B_5gBjBoyz1_1;
	wire w_dff_B_u41Sj2Aq7_1;
	wire w_dff_B_wYKy2GAs8_1;
	wire w_dff_B_05xGj70w6_1;
	wire w_dff_B_ykSk5iGP3_1;
	wire w_dff_B_6aNrz2ZU6_1;
	wire w_dff_B_rVL77JfP0_1;
	wire w_dff_B_a2zzzpxG1_1;
	wire w_dff_B_0lqUBRAk6_1;
	wire w_dff_B_q0MGXqm38_1;
	wire w_dff_B_dsNivNOQ9_1;
	wire w_dff_B_Iwv3UNpM2_1;
	wire w_dff_B_2gRP9Kha2_1;
	wire w_dff_B_SbEy35GQ2_1;
	wire w_dff_B_MHas7a3Z4_1;
	wire w_dff_B_SsfSV83S3_1;
	wire w_dff_B_VJ4NDuJq5_1;
	wire w_dff_B_3xCvqsgU0_1;
	wire w_dff_B_Hvnz8wtV3_1;
	wire w_dff_B_GRHxvnvb1_1;
	wire w_dff_B_copsStCz9_1;
	wire w_dff_B_g54p5iyo6_1;
	wire w_dff_B_IaJhPYqY2_1;
	wire w_dff_B_kyPMqsYh0_1;
	wire w_dff_B_W6V02sKH1_1;
	wire w_dff_B_gzhWT1iK0_1;
	wire w_dff_B_AmtNKtQH0_1;
	wire w_dff_B_TNbf3rd33_1;
	wire w_dff_B_oH3KqGwB4_1;
	wire w_dff_B_wEIEdFzp5_1;
	wire w_dff_B_7QXIm5Yn0_1;
	wire w_dff_B_oYSEhs1h1_1;
	wire w_dff_B_NxNILxUd8_1;
	wire w_dff_B_cWchFx2B2_1;
	wire w_dff_B_Saglca3F8_1;
	wire w_dff_B_dyXn8XrA1_1;
	wire w_dff_B_ZbQhgMU97_1;
	wire w_dff_B_Aax07fdp0_1;
	wire w_dff_B_1vQ5ORq25_1;
	wire w_dff_B_CjQAJZ9z5_1;
	wire w_dff_B_ZE1xVrXg4_1;
	wire w_dff_B_Fa4hIdED2_1;
	wire w_dff_B_WUvc9dgb7_1;
	wire w_dff_B_h1ZqDlFJ3_1;
	wire w_dff_B_KFiCfCiN7_1;
	wire w_dff_B_c2Igsh980_1;
	wire w_dff_B_OXCMwMYx9_1;
	wire w_dff_B_Xs4uT3ic5_1;
	wire w_dff_B_UxQEuFzx7_1;
	wire w_dff_B_V23efQt70_1;
	wire w_dff_B_a2Q06y577_1;
	wire w_dff_B_p4C8DXdO9_1;
	wire w_dff_B_AlgJPJUD7_1;
	wire w_dff_B_piHzdoiB6_1;
	wire w_dff_B_twgeBedW1_1;
	wire w_dff_B_wxuHUL808_1;
	wire w_dff_B_EiKE7WDD1_1;
	wire w_dff_B_mcgllPVV0_1;
	wire w_dff_B_mi42vg061_1;
	wire w_dff_B_sylcrNYg0_1;
	wire w_dff_B_s9HluGJc9_1;
	wire w_dff_B_9oAPPFJD4_1;
	wire w_dff_B_r1BgwDeh7_1;
	wire w_dff_B_keb4xBe01_1;
	wire w_dff_B_PmQBQZJ82_1;
	wire w_dff_B_EXJ4tpse4_1;
	wire w_dff_B_XXn03XVt7_1;
	wire w_dff_B_L2Do306Q9_1;
	wire w_dff_B_bWAoU4x65_1;
	wire w_dff_B_ak3ovxsm3_1;
	wire w_dff_B_fK0Zv3Bt1_1;
	wire w_dff_B_zR2l0qQX4_1;
	wire w_dff_B_7vS8L6GY2_1;
	wire w_dff_B_gRLERNxY0_1;
	wire w_dff_B_qkHWLBlB4_1;
	wire w_dff_B_PybMpjAB1_1;
	wire w_dff_B_HFhK5X3L2_1;
	wire w_dff_B_kOkW5tSF7_1;
	wire w_dff_B_mkB5CaAJ5_1;
	wire w_dff_B_1HiSq3Lm1_1;
	wire w_dff_B_NBLTAN7Q0_1;
	wire w_dff_B_erQVcywS2_1;
	wire w_dff_B_NYGj0Y1o1_1;
	wire w_dff_B_IldXXGwX6_1;
	wire w_dff_B_QYrHQz6Q2_1;
	wire w_dff_B_ILTw8DYX2_1;
	wire w_dff_B_hjRQWfnk3_1;
	wire w_dff_B_A2p1NaP77_1;
	wire w_dff_B_sCTWq8G43_1;
	wire w_dff_B_yA6YbsKe0_1;
	wire w_dff_B_yT2TeJI65_1;
	wire w_dff_B_gZqqw59y5_1;
	wire w_dff_B_qcdJzEly7_1;
	wire w_dff_B_GSQHUgRC2_1;
	wire w_dff_B_OkR3p2hZ6_1;
	wire w_dff_B_fhJQTi3w3_1;
	wire w_dff_B_vdgutqrR8_1;
	wire w_dff_B_yHJfLbJI9_1;
	wire w_dff_B_SljHnOOY0_1;
	wire w_dff_B_lJKQxDEb3_1;
	wire w_dff_B_Wl3a5Hia0_1;
	wire w_dff_B_3Ry4I1MU7_1;
	wire w_dff_B_I7q5oAJW0_1;
	wire w_dff_B_ryj4xiuG5_1;
	wire w_dff_B_FkILoM930_1;
	wire w_dff_B_4OpwQnyS8_1;
	wire w_dff_B_BtFzJvlK8_1;
	wire w_dff_B_xevlMDq26_1;
	wire w_dff_B_DCzy1yr71_1;
	wire w_dff_B_ttirPb0p5_1;
	wire w_dff_B_V6OycExF9_1;
	wire w_dff_B_d4Dqqnfg6_1;
	wire w_dff_B_OwwZINRB0_1;
	wire w_dff_B_ktBhtVTz7_1;
	wire w_dff_B_RzNlVu1r1_1;
	wire w_dff_B_HLDLkxPu9_1;
	wire w_dff_B_gtQXxrHa1_1;
	wire w_dff_B_8aA5e3yu7_1;
	wire w_dff_B_6rM5mEZx0_1;
	wire w_dff_B_N1FIAjYu3_1;
	wire w_dff_B_uuZLULmc9_1;
	wire w_dff_B_y39mqIOx5_1;
	wire w_dff_B_N66UojaU8_1;
	wire w_dff_B_kzgJ6SHl0_1;
	wire w_dff_B_aW1bQlwx5_1;
	wire w_dff_B_DCsPMNPK1_1;
	wire w_dff_B_VPO3duGm6_1;
	wire w_dff_B_ObMTLEoV8_1;
	wire w_dff_B_yqQPOCkE4_1;
	wire w_dff_B_etbc91OF2_1;
	wire w_dff_B_BPzNYXxU8_1;
	wire w_dff_B_YRzLklgY1_1;
	wire w_dff_B_THBOFXCS7_1;
	wire w_dff_B_LwRIqg1o0_1;
	wire w_dff_B_wfSShkjz8_1;
	wire w_dff_B_ongBu5qs5_1;
	wire w_dff_B_sYEdVRJL3_1;
	wire w_dff_B_ZAAZaKp33_1;
	wire w_dff_B_WV6TQTm70_1;
	wire w_dff_B_IdOjdoJ26_1;
	wire w_dff_B_qw3yPsm44_1;
	wire w_dff_B_ZDiVBwSW1_1;
	wire w_dff_B_OYW74MFD7_1;
	wire w_dff_B_82QcN2bB2_1;
	wire w_dff_B_F9V7fWIk4_1;
	wire w_dff_B_y9UtJkD21_1;
	wire w_dff_B_kK36N8uP3_1;
	wire w_dff_B_ZEYgtjty0_1;
	wire w_dff_B_oqDz8hAC1_1;
	wire w_dff_B_unukIL8g8_1;
	wire w_dff_B_LNj8l2Mm3_1;
	wire w_dff_B_rpPXZwUs2_1;
	wire w_dff_B_sSMNNu0M6_1;
	wire w_dff_B_VbDqiQwg3_1;
	wire w_dff_B_ozUNbSNK1_1;
	wire w_dff_B_98Shzfw17_1;
	wire w_dff_B_2IY5qGhI4_1;
	wire w_dff_B_SLvFabNq4_1;
	wire w_dff_B_qxZSQcba9_1;
	wire w_dff_B_KJsQRmJY9_1;
	wire w_dff_B_Xn7QxX964_1;
	wire w_dff_B_mXNgArBm6_1;
	wire w_dff_B_x0SIfecO0_1;
	wire w_dff_B_3Pfl5ZEQ4_1;
	wire w_dff_B_m51UgDzc6_1;
	wire w_dff_B_XIa552yP9_1;
	wire w_dff_B_tzj67nvd6_1;
	wire w_dff_B_Nanzewwn2_1;
	wire w_dff_B_3yRAxRhV6_1;
	wire w_dff_B_DZXN19Ym3_1;
	wire w_dff_B_6XQ7hKEd0_1;
	wire w_dff_B_ckUrSzjC9_1;
	wire w_dff_B_gS1NIQse5_1;
	wire w_dff_B_X5qHLXuE6_1;
	wire w_dff_B_TsvRSnEh7_1;
	wire w_dff_B_FcIdlVHP6_1;
	wire w_dff_B_y53I3yOU9_1;
	wire w_dff_B_EY0OYSmp4_1;
	wire w_dff_B_gvARfhkR2_1;
	wire w_dff_B_NpKctRtW2_1;
	wire w_dff_B_0E9cUlez9_1;
	wire w_dff_B_ibRxwUPP8_1;
	wire w_dff_B_xs3BxYij3_1;
	wire w_dff_B_r8jvjtir1_1;
	wire w_dff_B_kaDOa3CU8_1;
	wire w_dff_B_BPW3frcf6_1;
	wire w_dff_B_7kNDhn4b4_1;
	wire w_dff_B_8ScdTIkO8_1;
	wire w_dff_B_zHPOdMG66_1;
	wire w_dff_B_nZJqR1a20_1;
	wire w_dff_B_XnphZwK74_1;
	wire w_dff_B_3voclOSs7_1;
	wire w_dff_B_O2kuxKOs0_1;
	wire w_dff_B_xpL578oA7_1;
	wire w_dff_B_USkmvQ2t4_1;
	wire w_dff_B_zIZtKdkO8_1;
	wire w_dff_B_REkL5Tur8_1;
	wire w_dff_B_XcsPeYpc6_1;
	wire w_dff_B_0xOEg74p3_1;
	wire w_dff_B_ONtpKoir0_1;
	wire w_dff_B_8OQ14b2L7_1;
	wire w_dff_B_G9KYFOPh5_1;
	wire w_dff_B_uQRYcA7X6_1;
	wire w_dff_B_kbomD1TL5_1;
	wire w_dff_B_ArfNz0o08_1;
	wire w_dff_B_T7YQxieu8_1;
	wire w_dff_B_3kBdBnNv0_1;
	wire w_dff_B_dCiJrYpe1_1;
	wire w_dff_B_dAEAkRyB1_1;
	wire w_dff_B_6MefftY48_1;
	wire w_dff_B_JKi06wMq4_1;
	wire w_dff_B_JezrVyNm5_1;
	wire w_dff_B_ebkeY8eE6_1;
	wire w_dff_B_1KXdIPwK7_1;
	wire w_dff_B_wG01vPSr8_1;
	wire w_dff_B_2qgeSkaM3_1;
	wire w_dff_B_3JBG7tbr1_1;
	wire w_dff_B_nImkeq1M7_1;
	wire w_dff_B_TkuOc68t9_1;
	wire w_dff_B_ZwTUEMLH1_1;
	wire w_dff_B_m7MKIcwi0_1;
	wire w_dff_B_DxUyB6ww3_1;
	wire w_dff_B_OfJVT3ax0_1;
	wire w_dff_B_eVLHXhof4_1;
	wire w_dff_B_0HGfBFmk8_1;
	wire w_dff_B_B7Ah3vti3_1;
	wire w_dff_B_tolJagxi0_1;
	wire w_dff_B_yfR3WOZH0_1;
	wire w_dff_B_ZD3T5Btk8_1;
	wire w_dff_B_eHHOcdQg9_1;
	wire w_dff_B_MzMZgsoR4_1;
	wire w_dff_B_zPTnjEN10_1;
	wire w_dff_B_9IgSwGIK9_1;
	wire w_dff_B_lBw163TE5_1;
	wire w_dff_B_bNjQ7o7w2_1;
	wire w_dff_B_7LdLhKzY1_1;
	wire w_dff_B_bKqTumec4_1;
	wire w_dff_B_FFdO61uq1_1;
	wire w_dff_B_HHMDA5zG7_1;
	wire w_dff_B_gyYYBCfy4_1;
	wire w_dff_B_wi7HRvc36_1;
	wire w_dff_B_el9pkpPi1_1;
	wire w_dff_B_llOe2NHT7_1;
	wire w_dff_B_cR8OxUy66_1;
	wire w_dff_B_ML6Af0WK5_1;
	wire w_dff_B_n7lek9Bk3_1;
	wire w_dff_B_6kHImbUL5_1;
	wire w_dff_B_1fYz7J8g3_1;
	wire w_dff_B_P2PIbB795_1;
	wire w_dff_B_BUerrUPW6_1;
	wire w_dff_B_IEBvoBpi7_1;
	wire w_dff_B_wqUt48lV2_1;
	wire w_dff_B_vHtlslYq7_1;
	wire w_dff_B_6qiNbwWT0_1;
	wire w_dff_B_dro4N5VE5_1;
	wire w_dff_B_4VsBXKE91_1;
	wire w_dff_B_Q0I7I8ae0_1;
	wire w_dff_B_xv0YMTVj1_1;
	wire w_dff_B_a1QxwmEr6_1;
	wire w_dff_B_PrYNMY7t2_1;
	wire w_dff_B_X7aRTx155_1;
	wire w_dff_B_2DeyiiQs4_1;
	wire w_dff_B_dYDUkzgO3_1;
	wire w_dff_B_VQNox5Wu7_1;
	wire w_dff_B_kik3iT5f1_1;
	wire w_dff_B_qG0HeMm17_1;
	wire w_dff_B_0R1rp4Wc2_1;
	wire w_dff_B_u11I65Fp8_0;
	wire w_dff_B_n0LX8HK47_1;
	wire w_dff_B_6ns2AneW4_1;
	wire w_dff_B_1koqxMBQ5_1;
	wire w_dff_B_dFS5DP7C6_1;
	wire w_dff_B_Z9aypmpx9_1;
	wire w_dff_B_eH4ngXJK0_1;
	wire w_dff_B_mk1sOs1A8_1;
	wire w_dff_B_9Cy1jNDN7_1;
	wire w_dff_B_LrXHFHu72_1;
	wire w_dff_B_iPdCQyZc7_1;
	wire w_dff_B_AOIVlaK13_1;
	wire w_dff_B_fjcqt6UR5_1;
	wire w_dff_B_CRQgdMGd2_1;
	wire w_dff_B_Bp1dfDng5_0;
	wire w_dff_B_z1qPUNpM0_0;
	wire w_dff_B_XCngyXQD0_0;
	wire w_dff_B_fZWO75Y52_0;
	wire w_dff_B_ZEjg1Ehh8_0;
	wire w_dff_B_JBwtRBqg2_0;
	wire w_dff_B_HrtTerQR4_0;
	wire w_dff_B_dJbWj8eF4_0;
	wire w_dff_B_SbVYbqqq7_0;
	wire w_dff_B_5mEyW3ZQ4_0;
	wire w_dff_B_3PRkUcnj7_0;
	wire w_dff_A_BJ4y7Wle8_0;
	wire w_dff_A_wh3y0wNg4_0;
	wire w_dff_A_rDD0R9Uk3_0;
	wire w_dff_A_y2g2Omgw0_0;
	wire w_dff_A_dIvK8EgK9_0;
	wire w_dff_A_OSycrRUc6_0;
	wire w_dff_A_GPXpLpwF7_0;
	wire w_dff_A_d5Ti3UEX0_0;
	wire w_dff_A_vhdZGHMM4_0;
	wire w_dff_A_vlFk7etE4_0;
	wire w_dff_A_eTZknVkp3_0;
	wire w_dff_A_S3oaBWKP4_0;
	wire w_dff_B_koBkdfDe4_1;
	wire w_dff_B_WOnb8SOF2_1;
	wire w_dff_B_nEuXBt0h1_2;
	wire w_dff_B_JOzWbBhU9_2;
	wire w_dff_B_fUgv6U4v4_2;
	wire w_dff_B_tHlkeFko2_2;
	wire w_dff_B_dqBnVESn8_2;
	wire w_dff_B_jgzWMh1h8_2;
	wire w_dff_B_9IqJ6khm4_2;
	wire w_dff_B_JMbEtx3p4_2;
	wire w_dff_B_F8Kl8dPW8_2;
	wire w_dff_B_CVcCcHL35_2;
	wire w_dff_B_bZEdkymb4_2;
	wire w_dff_B_IRnNEqf71_2;
	wire w_dff_B_YM5kcdg20_2;
	wire w_dff_B_8CZW2qvp4_2;
	wire w_dff_B_sNv1zJeD5_2;
	wire w_dff_B_k0K2nnHz3_2;
	wire w_dff_B_rb1w8U7q5_2;
	wire w_dff_B_sCXdE0Tt4_2;
	wire w_dff_B_HBTy6h9n8_2;
	wire w_dff_B_jBWqYXq38_2;
	wire w_dff_B_jujs5ISR1_2;
	wire w_dff_B_AT4jU38D8_2;
	wire w_dff_B_IqqRYEiy4_2;
	wire w_dff_B_2IVRv3ae7_2;
	wire w_dff_B_JdbAeKTF4_2;
	wire w_dff_B_NIdbV4B44_2;
	wire w_dff_B_yjSWPEpy6_2;
	wire w_dff_B_N3XxefAG9_2;
	wire w_dff_B_cepbRAYc7_2;
	wire w_dff_B_XCfK2yRO3_2;
	wire w_dff_B_8dlMRbOE5_2;
	wire w_dff_B_hyXwfLLg6_2;
	wire w_dff_B_hdxH3QjP6_2;
	wire w_dff_B_xAcshE6C9_2;
	wire w_dff_B_wZIRk25T4_2;
	wire w_dff_B_d9ARTDuk8_2;
	wire w_dff_B_tg4T8bQB5_2;
	wire w_dff_B_MsXe6ssV0_2;
	wire w_dff_B_z7R67VBi6_2;
	wire w_dff_B_I48V4YaI3_2;
	wire w_dff_B_nhlUiY0X9_2;
	wire w_dff_B_UCUluUy38_2;
	wire w_dff_B_6tHIm0Zj1_2;
	wire w_dff_B_fDrxW39B4_2;
	wire w_dff_B_zUhDUf382_2;
	wire w_dff_B_hdtmYOMd1_2;
	wire w_dff_B_HHIV3MQM1_2;
	wire w_dff_B_LRdvF6EQ6_2;
	wire w_dff_B_CVZWGe6c4_2;
	wire w_dff_B_x8EtMWeH1_2;
	wire w_dff_B_oaMw4zbH6_2;
	wire w_dff_B_hWBi9QTS3_2;
	wire w_dff_B_MsJNs49r5_2;
	wire w_dff_B_tB4TPbVH7_2;
	wire w_dff_B_rZzduNnC5_2;
	wire w_dff_B_lv8uBgJO8_2;
	wire w_dff_B_VapzC66b9_2;
	wire w_dff_B_JoxeLlV34_2;
	wire w_dff_B_Z8eS5z1F6_2;
	wire w_dff_B_ePcqAiRz6_2;
	wire w_dff_B_JnwV1ZWt8_1;
	wire w_dff_B_qXSxj49q2_1;
	wire w_dff_B_5CsEPWPS6_1;
	wire w_dff_B_GW4GZKY47_1;
	wire w_dff_B_xEw3p8Zd7_1;
	wire w_dff_B_qOxhTNHt7_1;
	wire w_dff_B_0JORbhdS1_1;
	wire w_dff_B_LM8C4jpA7_1;
	wire w_dff_B_Ehttn7093_1;
	wire w_dff_B_H66ywrZl3_1;
	wire w_dff_B_9BjyQurF6_1;
	wire w_dff_B_PYOtlqJO2_0;
	wire w_dff_B_vWoNWi672_0;
	wire w_dff_B_Yp3G70995_0;
	wire w_dff_B_aYeKkPR34_0;
	wire w_dff_B_8amJfuLy1_0;
	wire w_dff_B_Pk2uFOrX4_0;
	wire w_dff_B_OLgVuWOW8_0;
	wire w_dff_B_WYbEhz6C4_0;
	wire w_dff_B_fxyJUvnQ9_0;
	wire w_dff_B_qFQVdwG56_0;
	wire w_dff_A_nk87A8Dq2_1;
	wire w_dff_A_Mcdi5QNK0_1;
	wire w_dff_A_ghVWx5al9_1;
	wire w_dff_A_f6FrMDOM6_1;
	wire w_dff_A_akaDuShF5_1;
	wire w_dff_A_cFeDyn1d0_1;
	wire w_dff_A_WoOF1ovi5_1;
	wire w_dff_A_A7m0i16D3_1;
	wire w_dff_A_X8l1TA9i6_1;
	wire w_dff_A_75M4gMx63_1;
	wire w_dff_A_zIOHEaBV8_1;
	wire w_dff_B_YpfZXQss1_1;
	wire w_dff_B_ax82Dsdr0_1;
	wire w_dff_B_cm0kPttC7_1;
	wire w_dff_B_XE2IO5qy3_1;
	wire w_dff_B_OuOoZMZN4_1;
	wire w_dff_B_nnBCEnVs7_1;
	wire w_dff_B_6pROSCHP8_1;
	wire w_dff_B_2SBE1Oq47_1;
	wire w_dff_B_ehtuY3Tn8_1;
	wire w_dff_B_Gp4NQj3s2_1;
	wire w_dff_B_NQTZLS0q4_1;
	wire w_dff_B_4jBcN43r6_0;
	wire w_dff_B_CGkeXy6N7_0;
	wire w_dff_B_o3HO7RTu9_0;
	wire w_dff_B_Y1CNqHxN0_0;
	wire w_dff_B_C4VeJW8r2_0;
	wire w_dff_B_1CAcnE9l7_0;
	wire w_dff_B_vqAhaM5b6_0;
	wire w_dff_B_nGS1uDC61_0;
	wire w_dff_B_5sbpvJjw0_0;
	wire w_dff_B_EHataNLT3_0;
	wire w_dff_A_QE8AgDb75_1;
	wire w_dff_A_0mUsjU6w3_1;
	wire w_dff_A_aF4XfnDL2_1;
	wire w_dff_A_gbt5IOib1_1;
	wire w_dff_A_1oH8ZtIp1_1;
	wire w_dff_A_TBAGzUVs1_1;
	wire w_dff_A_FuYVuRKB3_1;
	wire w_dff_A_ncEp9u7e5_1;
	wire w_dff_A_XSva6HVo6_1;
	wire w_dff_A_lOHNcVEa5_1;
	wire w_dff_A_2B9FjQxb3_1;
	wire w_dff_B_i52lIxVR4_1;
	wire w_dff_B_Dr5ldv727_1;
	wire w_dff_B_lhzLMJYF4_1;
	wire w_dff_B_xbZ3ChDl6_1;
	wire w_dff_B_FhL4hDBK2_1;
	wire w_dff_B_48HKwAtk5_1;
	wire w_dff_B_jSK22BhL5_1;
	wire w_dff_B_P5IiImCZ2_1;
	wire w_dff_B_zAkpJhzv9_1;
	wire w_dff_B_An3zfZ9k7_1;
	wire w_dff_B_fdbJkxX72_1;
	wire w_dff_B_EiUK8CGZ9_0;
	wire w_dff_B_AytBTrla6_0;
	wire w_dff_B_HU5yLeRN6_0;
	wire w_dff_B_lFt0TUh56_0;
	wire w_dff_B_VhFZKmrQ3_0;
	wire w_dff_B_8uuVBiwE2_0;
	wire w_dff_B_PWajHzqd0_0;
	wire w_dff_B_Lcsf8UQD7_0;
	wire w_dff_B_U0J3qJw59_0;
	wire w_dff_B_tvgH6RWW3_0;
	wire w_dff_A_G0CghVSE2_1;
	wire w_dff_A_mXmWR6iq6_1;
	wire w_dff_A_eATnJKXS0_1;
	wire w_dff_A_5amLb5yT3_1;
	wire w_dff_A_geN1YJdJ8_1;
	wire w_dff_A_NcAAZBOy2_1;
	wire w_dff_A_zCvsgT2n8_1;
	wire w_dff_A_xaus8U144_1;
	wire w_dff_A_Fs5VNS545_1;
	wire w_dff_A_5J14Okyl9_1;
	wire w_dff_A_xi9bByvv3_1;
	wire w_dff_B_apthHD0e7_1;
	wire w_dff_B_3CNzG3aN4_1;
	wire w_dff_B_PzWddbZx0_1;
	wire w_dff_B_CITiLbRG3_1;
	wire w_dff_B_NmzAodJC2_1;
	wire w_dff_B_XNOh7ZWf3_1;
	wire w_dff_B_1LpawFoo9_1;
	wire w_dff_B_6YCGpQLP2_1;
	wire w_dff_B_Ohoibt1s9_1;
	wire w_dff_B_MvQb0VFd2_1;
	wire w_dff_B_yegT27uo2_1;
	wire w_dff_B_64NhoyK05_0;
	wire w_dff_B_d3hNrJBK0_0;
	wire w_dff_B_DrIMhhQN8_0;
	wire w_dff_B_vfYykq8t3_0;
	wire w_dff_B_mj6D7phu8_0;
	wire w_dff_B_2eSu4Mxe3_0;
	wire w_dff_B_tfxb9vAU6_0;
	wire w_dff_B_2tc02Oid4_0;
	wire w_dff_B_1UsXatsV3_0;
	wire w_dff_B_3nD9Myey6_0;
	wire w_dff_A_9mQsSc2g5_1;
	wire w_dff_A_Sjtr7ByO3_1;
	wire w_dff_A_IcP6V3Gg1_1;
	wire w_dff_A_6pYpxFGI2_1;
	wire w_dff_A_qTjsp5wm9_1;
	wire w_dff_A_vjUs6s9b9_1;
	wire w_dff_A_C7Mk18sD1_1;
	wire w_dff_A_fAbhAN8Z0_1;
	wire w_dff_A_oP21dmZr9_1;
	wire w_dff_A_KjjI57cC0_1;
	wire w_dff_A_E6PWdTsO3_1;
	wire w_dff_B_lH4AGOPK9_1;
	wire w_dff_B_pZCIYfz65_1;
	wire w_dff_B_aN1T8Bvq5_1;
	wire w_dff_B_drALFYzw0_1;
	wire w_dff_B_mqANwPTm8_1;
	wire w_dff_B_bzga3F7h5_1;
	wire w_dff_B_tmtsrMiO3_1;
	wire w_dff_B_JrbHG7JQ6_1;
	wire w_dff_B_D8UuVnSp3_1;
	wire w_dff_B_BIWYyO460_1;
	wire w_dff_B_Wq2Kv3s35_1;
	wire w_dff_B_rScQOwiB1_0;
	wire w_dff_B_wggJHljV9_0;
	wire w_dff_B_a9eyFLI59_0;
	wire w_dff_B_6mFfBnNw7_0;
	wire w_dff_B_ZNYORSge3_0;
	wire w_dff_B_50Jg3p789_0;
	wire w_dff_B_JD6PozWB6_0;
	wire w_dff_B_yb3ddDnU1_0;
	wire w_dff_B_apjOOWYS0_0;
	wire w_dff_A_ZBUv3hRO5_1;
	wire w_dff_A_fnYVZVd12_1;
	wire w_dff_A_CMyBLQ227_1;
	wire w_dff_A_3qhdM4hb1_1;
	wire w_dff_A_fKZfkly18_1;
	wire w_dff_A_sUQCH0aM0_1;
	wire w_dff_A_jWvFyAXy9_1;
	wire w_dff_A_9fOCJ18c2_1;
	wire w_dff_A_qbZioxW05_1;
	wire w_dff_A_HV3sCXwW3_1;
	wire w_dff_B_QrDZuXk75_1;
	wire w_dff_B_8U7dz88v0_1;
	wire w_dff_B_4eQubw3Y2_1;
	wire w_dff_B_EyYA1Y8n3_1;
	wire w_dff_B_vpjXqzBJ5_1;
	wire w_dff_B_v4zOHPYL9_1;
	wire w_dff_B_tGZy8yPl4_1;
	wire w_dff_B_ih7J4Yym1_1;
	wire w_dff_B_iHJZqq0E4_1;
	wire w_dff_B_Hczv6KUZ7_1;
	wire w_dff_B_60htQl7F3_0;
	wire w_dff_B_44xPq9ta6_0;
	wire w_dff_B_BZYUnd6j5_0;
	wire w_dff_B_ymnNBS8V3_0;
	wire w_dff_B_aCjEXt151_0;
	wire w_dff_B_vCJ1xMxt7_0;
	wire w_dff_B_pkYusNoI1_0;
	wire w_dff_B_a4Snyv5j7_0;
	wire w_dff_A_kte2a3xO4_1;
	wire w_dff_A_sJigHy9A3_1;
	wire w_dff_A_c8gRWP3l6_1;
	wire w_dff_A_WtoWpsNH6_1;
	wire w_dff_A_W4V3Bqox1_1;
	wire w_dff_A_4qbFL7Py8_1;
	wire w_dff_A_8jqlQjjl5_1;
	wire w_dff_A_rwhWemd01_1;
	wire w_dff_A_7o8BL2rh8_1;
	wire w_dff_B_WyKDqC1u0_1;
	wire w_dff_B_DSabBSQw0_1;
	wire w_dff_B_wYbgBOcU3_1;
	wire w_dff_B_7BPj9n451_1;
	wire w_dff_B_nQ2cNvO85_1;
	wire w_dff_B_OjKeyUXM1_1;
	wire w_dff_B_ctM5bRNX0_1;
	wire w_dff_B_j1GPd84g8_1;
	wire w_dff_B_qDT9jkU24_1;
	wire w_dff_B_9hYt5XTP8_1;
	wire w_dff_B_nxXT2Woi2_0;
	wire w_dff_B_5fQYakNd8_0;
	wire w_dff_B_IqNuwjlM2_0;
	wire w_dff_B_cWKUjQgH9_0;
	wire w_dff_B_7mwu9n2e0_0;
	wire w_dff_B_zY4VCRG69_0;
	wire w_dff_B_Nie2abV93_0;
	wire w_dff_B_JCTp6ct86_0;
	wire w_dff_A_Vm8e3S9c9_1;
	wire w_dff_A_LTLZkO4D4_1;
	wire w_dff_A_YNaUGyI08_1;
	wire w_dff_A_YdmhWq4o0_1;
	wire w_dff_A_aH0kG7nK6_1;
	wire w_dff_A_nkz9XtE07_1;
	wire w_dff_A_H7g02P1A2_1;
	wire w_dff_A_eDaLSKlu8_1;
	wire w_dff_A_IMnnVenA9_1;
	wire w_dff_B_n4RELTC35_1;
	wire w_dff_B_XgKRyzh94_1;
	wire w_dff_B_RhTGLby80_1;
	wire w_dff_B_ZRKTzA5T5_1;
	wire w_dff_B_BGWNLnmi0_1;
	wire w_dff_B_DP6C2C9o9_1;
	wire w_dff_B_LfiWfs5q6_1;
	wire w_dff_B_a8uOOsQh7_1;
	wire w_dff_B_kZXr2ywO9_0;
	wire w_dff_B_tfKKtK025_0;
	wire w_dff_B_SSCxDJ4F7_0;
	wire w_dff_B_nr4biGt38_0;
	wire w_dff_B_CZlildiN7_0;
	wire w_dff_B_vDfTjoF11_0;
	wire w_dff_A_b56HJCUi8_1;
	wire w_dff_A_qSmd7q688_1;
	wire w_dff_A_ZTURvvJv4_1;
	wire w_dff_A_qir4WC4H3_1;
	wire w_dff_A_qTk1zyAX2_1;
	wire w_dff_A_YdbMfr8e5_1;
	wire w_dff_A_GWaUef9G5_1;
	wire w_dff_B_USfsmGXm0_1;
	wire w_dff_B_lWRSwoYc0_1;
	wire w_dff_B_sdsv42lk8_1;
	wire w_dff_B_XQRFyYYN7_1;
	wire w_dff_B_HeOI2PSo2_1;
	wire w_dff_B_Ry5I1mhL5_1;
	wire w_dff_B_PspZc4QJ1_1;
	wire w_dff_B_mpPu7rD83_0;
	wire w_dff_B_i3HfL7z81_0;
	wire w_dff_B_NvseCO2M7_0;
	wire w_dff_B_veZRmBQf5_0;
	wire w_dff_B_l8h2kqKv1_0;
	wire w_dff_A_Tz4EQcmS4_1;
	wire w_dff_A_pLs5YupV5_1;
	wire w_dff_A_W3HsODiu8_1;
	wire w_dff_A_gtlsd8vm0_1;
	wire w_dff_A_ac1VM2QA6_1;
	wire w_dff_A_6OXjizs55_1;
	wire w_dff_B_tjKHlDfa3_1;
	wire w_dff_B_FKK0XW893_1;
	wire w_dff_B_9NEI6zxU5_1;
	wire w_dff_B_GTSAcAkx5_1;
	wire w_dff_B_J2ojcNg75_1;
	wire w_dff_B_G3MHIb661_1;
	wire w_dff_B_rgvWZtm54_0;
	wire w_dff_B_jazBqxMe8_0;
	wire w_dff_B_saUc9m3L0_0;
	wire w_dff_B_SJt7GV7E3_0;
	wire w_dff_A_teWPpJ3x2_1;
	wire w_dff_A_f3GD0nUL2_1;
	wire w_dff_A_BTauswms8_1;
	wire w_dff_A_IBuaDJlC0_1;
	wire w_dff_A_lgICghwQ9_1;
	wire w_dff_B_frxD2xVz1_1;
	wire w_dff_B_g5XiQJX29_1;
	wire w_dff_B_GlvTNpIt5_1;
	wire w_dff_A_mSqC7HeX1_0;
	wire w_dff_A_Fc4YPKTA5_0;
	wire w_dff_B_2vRuOUkq5_1;
	wire w_dff_A_YtIxMlso6_0;
	wire w_dff_B_jo2C4wSM4_1;
	wire w_dff_A_8iyxgJFi0_1;
	wire w_dff_B_sIVTiUs64_2;
	wire w_dff_B_byKfvmww9_1;
	wire w_dff_A_qNRg8aGX1_0;
	wire w_dff_A_JgXN2zTt1_0;
	wire w_dff_A_DfQ8exKU5_0;
	wire w_dff_A_XtxeZWxf2_0;
	wire w_dff_A_HCtayFC97_0;
	wire w_dff_A_80Tal6Wq3_0;
	wire w_dff_A_17tMaAR57_0;
	wire w_dff_A_UBTuDwGq1_0;
	wire w_dff_A_oUoOvbm24_0;
	wire w_dff_A_hBNQuMGh6_0;
	wire w_dff_A_ZYSSPDsR3_0;
	wire w_dff_A_lvVskOPa4_0;
	wire w_dff_A_sifpBE7k8_0;
	wire w_dff_A_RmpMzXNi0_0;
	wire w_dff_A_VO2i2IdE4_0;
	wire w_dff_A_GYSUPLGE8_0;
	wire w_dff_A_k1Zd2eOK2_0;
	wire w_dff_A_alQEwqyh8_0;
	wire w_dff_A_Lby3IRmd5_0;
	wire w_dff_A_STlUFQBE4_0;
	wire w_dff_A_CburmB6r4_0;
	wire w_dff_A_TwfLiWdX0_0;
	wire w_dff_A_phh4mHJV9_0;
	wire w_dff_A_5kSOOloa8_0;
	wire w_dff_A_nRGcuvUV7_0;
	wire w_dff_A_wMLIcOJV0_0;
	wire w_dff_A_AW3zlEQG8_0;
	wire w_dff_A_IHV4G6Sb8_0;
	wire w_dff_A_5b8AV0XN8_0;
	wire w_dff_A_DGqxklfv6_0;
	wire w_dff_A_MjMeCmeQ8_0;
	wire w_dff_A_KDIwBGNi1_0;
	wire w_dff_A_864cxI9s6_0;
	wire w_dff_A_PaXeYqjV7_0;
	wire w_dff_A_3xPJlGV88_0;
	wire w_dff_A_R6u16fb98_0;
	wire w_dff_A_tf8mc7TZ5_0;
	wire w_dff_A_vDJPMjFE9_0;
	wire w_dff_A_BvGu7WyE3_0;
	wire w_dff_A_h5l2llis0_0;
	wire w_dff_A_TvAQHO4q6_0;
	wire w_dff_A_xyr3zLB41_0;
	wire w_dff_A_lMon71Tu2_0;
	wire w_dff_A_kyZTZRFM8_0;
	wire w_dff_A_rPD8mdkc9_1;
	wire w_dff_B_WUFQEIHg0_1;
	wire w_dff_A_t3yutd8v3_0;
	wire w_dff_A_2IW4mItI8_0;
	wire w_dff_A_vlMTcgpY1_0;
	wire w_dff_A_fbo78wwa9_0;
	wire w_dff_A_4R9mg1Gv7_0;
	wire w_dff_A_vTHGO2To3_0;
	wire w_dff_A_jQ28pvgX0_0;
	wire w_dff_A_9q6bxR0N9_0;
	wire w_dff_A_Yahpox9g3_0;
	wire w_dff_A_RKyrTVUw0_0;
	wire w_dff_A_DrxZLU1J7_0;
	wire w_dff_A_drsOUfEZ3_0;
	wire w_dff_A_HuVd3Y6V7_0;
	wire w_dff_A_e74l0oWE2_0;
	wire w_dff_A_I04age3X6_0;
	wire w_dff_A_cnvKZSoj3_0;
	wire w_dff_A_rFllEZ7S9_0;
	wire w_dff_A_ArdhJ4v70_0;
	wire w_dff_A_t8FkTvUv5_0;
	wire w_dff_A_TIzXt2Qc1_0;
	wire w_dff_A_wcACY4Mm1_0;
	wire w_dff_A_9s1Sia4g4_0;
	wire w_dff_A_VMbvWN9B1_0;
	wire w_dff_A_es8PT67q7_0;
	wire w_dff_A_3tZjujnG8_0;
	wire w_dff_A_nKUHsgCu2_0;
	wire w_dff_A_XHaYsywL2_0;
	wire w_dff_A_mqhKkZ8E0_0;
	wire w_dff_A_4cySiSeH1_0;
	wire w_dff_A_HB7cFgzJ3_0;
	wire w_dff_A_hwbYGpQC2_0;
	wire w_dff_A_dCYxRYtA2_0;
	wire w_dff_A_rVwR51FL1_0;
	wire w_dff_A_5tASqAVF5_0;
	wire w_dff_A_UGPkjZmw0_0;
	wire w_dff_A_EvEAvwR46_0;
	wire w_dff_A_WMyZgvck7_0;
	wire w_dff_A_N6AoFGDw4_0;
	wire w_dff_A_ApnZFqMo9_0;
	wire w_dff_A_8Taggs821_0;
	wire w_dff_A_rg9oEtRT9_0;
	wire w_dff_A_HUmEwnRZ3_1;
	wire w_dff_B_3t9gZx5K6_1;
	wire w_dff_B_L7VvIAtI3_1;
	wire w_dff_B_okdm2yDn5_1;
	wire w_dff_B_vlaR4Psj6_1;
	wire w_dff_B_TsRoWXeD1_1;
	wire w_dff_B_L6p6CLBb1_1;
	wire w_dff_B_YiE75Lzf9_1;
	wire w_dff_B_2zV4ajEy0_1;
	wire w_dff_B_D5roRV2S7_1;
	wire w_dff_B_VLSOsmEX6_1;
	wire w_dff_B_8SXLJU0a1_1;
	wire w_dff_B_0hnHS7hT4_1;
	wire w_dff_B_MzaqPRWa0_1;
	wire w_dff_B_5dBb4DJN7_1;
	wire w_dff_B_bL39RRKl0_1;
	wire w_dff_B_SqYK75VZ2_1;
	wire w_dff_B_31AAucs20_1;
	wire w_dff_B_otlpwXtr3_1;
	wire w_dff_B_v6pmgBCp7_1;
	wire w_dff_B_B8LIxpM91_1;
	wire w_dff_B_JPKN5Tqy6_1;
	wire w_dff_B_HxKgMiqD4_1;
	wire w_dff_B_Scn7qKiP2_1;
	wire w_dff_B_HFWmZ27m9_1;
	wire w_dff_B_K3Nt58Zx1_1;
	wire w_dff_B_NTV7a2sP9_1;
	wire w_dff_B_sMCjv46i2_1;
	wire w_dff_B_VHZkwYA20_1;
	wire w_dff_B_sfJyiSy11_1;
	wire w_dff_B_G652oqZV7_1;
	wire w_dff_B_Kw3aQ7mJ5_1;
	wire w_dff_B_7HOgLgjF9_1;
	wire w_dff_B_2rB4suMf6_1;
	wire w_dff_B_Tt7ssnoQ1_1;
	wire w_dff_B_BAK52qaT6_1;
	wire w_dff_B_08Y2FHn92_1;
	wire w_dff_B_APixYkF69_1;
	wire w_dff_B_jxu3HVWu3_1;
	wire w_dff_A_3Se68il30_0;
	wire w_dff_A_qegC0KNM3_0;
	wire w_dff_A_T7PijzyN8_0;
	wire w_dff_A_U99S566E9_0;
	wire w_dff_A_a5F5TQay5_0;
	wire w_dff_A_gYHFqeoV4_0;
	wire w_dff_A_Ixnpqw4C1_0;
	wire w_dff_A_H5hEAAHK7_0;
	wire w_dff_A_tzzZlqe55_0;
	wire w_dff_A_gsbXq6Qo4_0;
	wire w_dff_A_Eiy7Uz6W0_0;
	wire w_dff_A_KtEIAcWO1_0;
	wire w_dff_A_CZOV7ISu0_0;
	wire w_dff_A_hom3Zi0f2_0;
	wire w_dff_A_I8A3ZDls4_0;
	wire w_dff_A_EAJPG4996_0;
	wire w_dff_A_O4TzIQaN9_0;
	wire w_dff_A_o6ONkrSf6_0;
	wire w_dff_A_3eR9Xw4o1_0;
	wire w_dff_A_7NH5S5IB5_0;
	wire w_dff_A_R7hFAMTz8_0;
	wire w_dff_A_Kish0dB56_0;
	wire w_dff_A_tsK7WZvd3_0;
	wire w_dff_A_xG60JkBl0_0;
	wire w_dff_A_mlHfyNgV3_0;
	wire w_dff_A_Rci0Molr9_0;
	wire w_dff_A_PVZvRimo4_0;
	wire w_dff_A_cag03PwF6_0;
	wire w_dff_A_j1DM6ePW0_0;
	wire w_dff_A_BQnAje3Q7_0;
	wire w_dff_A_NhyM3Bc79_0;
	wire w_dff_A_Unu0pAN28_0;
	wire w_dff_A_0kKlBQdF0_0;
	wire w_dff_A_BgfZlWBi2_0;
	wire w_dff_A_PDnNGCep8_0;
	wire w_dff_A_BRoNz3jn2_0;
	wire w_dff_A_14cqpYVj0_0;
	wire w_dff_A_iTXaZvbS8_0;
	wire w_dff_A_9NszZZ8G3_1;
	wire w_dff_B_lU9l0C5p5_1;
	wire w_dff_B_xrLqgSAx0_1;
	wire w_dff_B_monT6oy97_1;
	wire w_dff_B_Tyc6hKCI3_1;
	wire w_dff_B_vi922Aph6_1;
	wire w_dff_B_qvDo52W75_1;
	wire w_dff_B_noQNMYPZ2_1;
	wire w_dff_B_t80WDKL63_1;
	wire w_dff_B_OFx7J3Sg9_1;
	wire w_dff_B_oW5DSX7p3_1;
	wire w_dff_B_ueSlggYk1_1;
	wire w_dff_B_AqGEbTsd4_1;
	wire w_dff_B_ggtqc0Wz1_1;
	wire w_dff_B_6P39f6xr3_1;
	wire w_dff_B_3GqyIPiY7_1;
	wire w_dff_B_2bK0TQyd9_1;
	wire w_dff_B_eGtVeBXP3_1;
	wire w_dff_B_oR4LQKt69_1;
	wire w_dff_B_hB3YcFAy3_1;
	wire w_dff_B_VysaI1qI3_1;
	wire w_dff_B_eK0D9hSg1_1;
	wire w_dff_B_v5yPIENZ2_1;
	wire w_dff_B_WlQVzxEd2_1;
	wire w_dff_B_2puEdKtI9_1;
	wire w_dff_B_w4bNLSnL4_1;
	wire w_dff_B_05lzDWlB2_1;
	wire w_dff_B_OeihB6SH1_1;
	wire w_dff_B_BbmTrQTR7_1;
	wire w_dff_B_FqDt8CYB4_1;
	wire w_dff_B_LysVxLLV6_1;
	wire w_dff_B_Gh9WNbTS0_1;
	wire w_dff_B_oly3NsYK1_1;
	wire w_dff_B_VPvJsWGj0_1;
	wire w_dff_B_XsTpae6H8_1;
	wire w_dff_B_5vRFOpjz6_1;
	wire w_dff_A_28fmAf4M3_0;
	wire w_dff_A_gv55jvDa9_0;
	wire w_dff_A_mUVL712O0_0;
	wire w_dff_A_EVGLiU8n8_0;
	wire w_dff_A_lLe2K2uN4_0;
	wire w_dff_A_Q83hYziu9_0;
	wire w_dff_A_JhB8Y5r74_0;
	wire w_dff_A_YcPnmJBb5_0;
	wire w_dff_A_wwubtDUj4_0;
	wire w_dff_A_D94wLc9M4_0;
	wire w_dff_A_uwkHHHXP5_0;
	wire w_dff_A_ev3T4ELG1_0;
	wire w_dff_A_YbTiujcb2_0;
	wire w_dff_A_WsLhl5zJ4_0;
	wire w_dff_A_qeBLLR2w4_0;
	wire w_dff_A_2Fgg3fG85_0;
	wire w_dff_A_JDd2GKi55_0;
	wire w_dff_A_64SMlF383_0;
	wire w_dff_A_su2s0Tvr5_0;
	wire w_dff_A_aRAuyn407_0;
	wire w_dff_A_xA13lmIc0_0;
	wire w_dff_A_DTTdvm9I0_0;
	wire w_dff_A_PTgevmWC4_0;
	wire w_dff_A_NcbltGHV6_0;
	wire w_dff_A_kprWxV2v2_0;
	wire w_dff_A_sxDBOWrp1_0;
	wire w_dff_A_RSMlVI9d3_0;
	wire w_dff_A_HrUUWE7i2_0;
	wire w_dff_A_XE4UNfHk2_0;
	wire w_dff_A_Thmjh4gW0_0;
	wire w_dff_A_2rnCKYeo7_0;
	wire w_dff_A_juz2ebfG8_0;
	wire w_dff_A_WHW0Pjbg7_0;
	wire w_dff_A_qV0J2Adw5_0;
	wire w_dff_A_B7YqcfYP3_0;
	wire w_dff_A_VEujq0b56_1;
	wire w_dff_B_OJfJScoz0_1;
	wire w_dff_B_joy5pEiW6_1;
	wire w_dff_B_3DAOgqIv0_1;
	wire w_dff_B_YBPywL6Y7_1;
	wire w_dff_B_EnBhvp3R5_1;
	wire w_dff_B_C964AZh05_1;
	wire w_dff_B_hL3MVVJ48_1;
	wire w_dff_B_UVMXs8U84_1;
	wire w_dff_B_NilN6uRf9_1;
	wire w_dff_B_lrcE3rTO2_1;
	wire w_dff_B_OcEBqq0a0_1;
	wire w_dff_B_rGFg2lv54_1;
	wire w_dff_B_C98GHJac1_1;
	wire w_dff_B_SRazcrER0_1;
	wire w_dff_B_B5Mhl2501_1;
	wire w_dff_B_XCivvqJI1_1;
	wire w_dff_B_yzdRFT6X2_1;
	wire w_dff_B_8XdL0IZy2_1;
	wire w_dff_B_rd4GnHpT2_1;
	wire w_dff_B_GAred9fU3_1;
	wire w_dff_B_ScXbBoIh5_1;
	wire w_dff_B_CEfqVYqh2_1;
	wire w_dff_B_u2mvNLNg6_1;
	wire w_dff_B_rdiRkRYn2_1;
	wire w_dff_B_LFjcMIIR9_1;
	wire w_dff_B_qrdrG9vH9_1;
	wire w_dff_B_hA2MNSKg1_1;
	wire w_dff_B_paERo2nw3_1;
	wire w_dff_B_50uwYBqb8_1;
	wire w_dff_B_5bCHPLMj2_1;
	wire w_dff_B_roJGW98C6_1;
	wire w_dff_B_SiMRqYSP0_1;
	wire w_dff_A_TfVGntJz7_0;
	wire w_dff_A_cb660BSI2_0;
	wire w_dff_A_wsJKOmr06_0;
	wire w_dff_A_OarxkGwb9_0;
	wire w_dff_A_MJEZPcC65_0;
	wire w_dff_A_jE0oqnOV1_0;
	wire w_dff_A_NgTIrXBe0_0;
	wire w_dff_A_WOEk7TDI7_0;
	wire w_dff_A_ZwcKZ1oD1_0;
	wire w_dff_A_1KYVI5oj1_0;
	wire w_dff_A_q3sEG3wu9_0;
	wire w_dff_A_FECjCLY76_0;
	wire w_dff_A_VVB6rwfg3_0;
	wire w_dff_A_RgaFQV2E3_0;
	wire w_dff_A_V0BsDLNf3_0;
	wire w_dff_A_PHckNOMP3_0;
	wire w_dff_A_796bviRN4_0;
	wire w_dff_A_ha7oxkKw9_0;
	wire w_dff_A_fJfDg6ol7_0;
	wire w_dff_A_m6oYLtBJ3_0;
	wire w_dff_A_atYdfedi5_0;
	wire w_dff_A_iQ4PABgr5_0;
	wire w_dff_A_jrbihYW94_0;
	wire w_dff_A_VNghTjrV4_0;
	wire w_dff_A_uMVnOkCX0_0;
	wire w_dff_A_T6f6kl7h9_0;
	wire w_dff_A_G7SOcXHi1_0;
	wire w_dff_A_Wpkx4X1d1_0;
	wire w_dff_A_wON9vDc00_0;
	wire w_dff_A_pKmVraOf9_0;
	wire w_dff_A_ecIxD9CN5_0;
	wire w_dff_A_3ewd5nH07_0;
	wire w_dff_A_iE7a1jkd8_1;
	wire w_dff_B_SHXBKMV59_1;
	wire w_dff_B_KUkdH2Ek2_1;
	wire w_dff_B_jSczWzAw1_1;
	wire w_dff_B_e7XHIZua4_1;
	wire w_dff_B_oeIymY4S7_1;
	wire w_dff_B_qvpSU4mg0_1;
	wire w_dff_B_YCHuXqUO9_1;
	wire w_dff_B_Dlg3pveE8_1;
	wire w_dff_B_Y6Ph1RZp8_1;
	wire w_dff_B_7bbmL7kk0_1;
	wire w_dff_B_82q5e7au1_1;
	wire w_dff_B_0NGNH7rw5_1;
	wire w_dff_B_sb2qU9gS3_1;
	wire w_dff_B_ca2ebekT1_1;
	wire w_dff_B_WtQrNsz83_1;
	wire w_dff_B_DXAwpNOh7_1;
	wire w_dff_B_LYqCxyIv1_1;
	wire w_dff_B_0xslFham9_1;
	wire w_dff_B_BPA1vyTb9_1;
	wire w_dff_B_SKAL9PmQ0_1;
	wire w_dff_B_2CZqNCrI2_1;
	wire w_dff_B_12IyrgCF9_1;
	wire w_dff_B_cs4ZLtuU8_1;
	wire w_dff_B_ZgCJ9OWN6_1;
	wire w_dff_B_oXIPgjlU4_1;
	wire w_dff_B_rRGPNQS83_1;
	wire w_dff_B_SGNPYJPA7_1;
	wire w_dff_B_KRdIAUVx8_1;
	wire w_dff_B_AYmBTs4D8_1;
	wire w_dff_A_MsZw9eL00_0;
	wire w_dff_A_S9aX8mER4_0;
	wire w_dff_A_mhz7RFrQ9_0;
	wire w_dff_A_eOpELvlj0_0;
	wire w_dff_A_fncPAUtS0_0;
	wire w_dff_A_7CsSnZhN1_0;
	wire w_dff_A_nWL8wY5z6_0;
	wire w_dff_A_XvWY4woz7_0;
	wire w_dff_A_V5Yvs6a06_0;
	wire w_dff_A_aJmCCQqP3_0;
	wire w_dff_A_AF8J90EB8_0;
	wire w_dff_A_DrVyjojO3_0;
	wire w_dff_A_SZnW5jyC4_0;
	wire w_dff_A_Hput9qZ54_0;
	wire w_dff_A_DCA00LGs1_0;
	wire w_dff_A_ifkn9wne2_0;
	wire w_dff_A_rnapPzg55_0;
	wire w_dff_A_mbKfXsXN0_0;
	wire w_dff_A_LDsKEhHh2_0;
	wire w_dff_A_zzaQnLjh7_0;
	wire w_dff_A_ZYQKrtTy8_0;
	wire w_dff_A_XRk1wtlT0_0;
	wire w_dff_A_RXDF3Jaj7_0;
	wire w_dff_A_KkKty4pY6_0;
	wire w_dff_A_PW1IC8L31_0;
	wire w_dff_A_Pi5vtkFv3_0;
	wire w_dff_A_Cq33Vq0E9_0;
	wire w_dff_A_PPh594NK9_0;
	wire w_dff_A_pnmCap4I7_0;
	wire w_dff_A_JKTgIqrw1_1;
	wire w_dff_B_8tM1nnR65_1;
	wire w_dff_B_expECOPx3_1;
	wire w_dff_B_dGtnS4Ig9_1;
	wire w_dff_B_WZX3xJTF5_1;
	wire w_dff_B_AKeJy0H19_1;
	wire w_dff_B_0L4ounem3_1;
	wire w_dff_B_qNH2hI4z3_1;
	wire w_dff_B_qBuVi36n1_1;
	wire w_dff_B_mWMq3leq7_1;
	wire w_dff_B_JVaVW0bZ0_1;
	wire w_dff_B_wTJPMqFx7_1;
	wire w_dff_B_7NRFgcrF2_1;
	wire w_dff_B_ZrTlRkxe0_1;
	wire w_dff_B_fE8E5YMv9_1;
	wire w_dff_B_jxd1XQPV9_1;
	wire w_dff_B_xdaXtQ4L7_1;
	wire w_dff_B_BSxM0G4N5_1;
	wire w_dff_B_vos2f6LB7_1;
	wire w_dff_B_OpBSgC7a5_1;
	wire w_dff_B_gZP13rbP1_1;
	wire w_dff_B_UNG6iTBt4_1;
	wire w_dff_B_Ct6SxtCE4_1;
	wire w_dff_B_v9jalWxg6_1;
	wire w_dff_B_qUdHmnrM6_1;
	wire w_dff_B_5LHCkCEA4_1;
	wire w_dff_B_G8Fc5G387_1;
	wire w_dff_A_o0IdYv1X2_0;
	wire w_dff_A_41d7oRsv5_0;
	wire w_dff_A_YlLJb8ht6_0;
	wire w_dff_A_fFEXxIo36_0;
	wire w_dff_A_f37HOTUI0_0;
	wire w_dff_A_hB5TfpfO7_0;
	wire w_dff_A_U0MRCOKw7_0;
	wire w_dff_A_a49wjfty6_0;
	wire w_dff_A_ZDdbKGXc0_0;
	wire w_dff_A_pJp30FFi1_0;
	wire w_dff_A_tfuJ1Uo45_0;
	wire w_dff_A_l6USH4Oj8_0;
	wire w_dff_A_ic76lS2t2_0;
	wire w_dff_A_PLur7qtH0_0;
	wire w_dff_A_gN9wrMQX9_0;
	wire w_dff_A_dnwwuee63_0;
	wire w_dff_A_cpotRyDG6_0;
	wire w_dff_A_zRKrqAC58_0;
	wire w_dff_A_0tUIz5fG9_0;
	wire w_dff_A_Mtw9PDXq7_0;
	wire w_dff_A_9KWDlbn13_0;
	wire w_dff_A_A5AhjcCE6_0;
	wire w_dff_A_diIkPePp5_0;
	wire w_dff_A_Wb3qlsaT2_0;
	wire w_dff_A_RNesFzje9_0;
	wire w_dff_A_PEKduRXH7_0;
	wire w_dff_A_3CJq4Na68_1;
	wire w_dff_B_VrrZgCmV6_1;
	wire w_dff_B_mDYnHiFa7_1;
	wire w_dff_B_xohbVPTK9_1;
	wire w_dff_B_o7QfjYe32_1;
	wire w_dff_B_VbRvaQ872_1;
	wire w_dff_B_MjjmvXDn0_1;
	wire w_dff_B_e3iHZ4Zg2_1;
	wire w_dff_B_USundpJN9_1;
	wire w_dff_B_2WSZ42HF4_1;
	wire w_dff_B_GaVuTz163_1;
	wire w_dff_B_llBApBEW4_1;
	wire w_dff_B_BNOntGvT6_1;
	wire w_dff_B_aExB5qGr1_1;
	wire w_dff_B_Lwq3ozrN1_1;
	wire w_dff_B_diMeUvQl1_1;
	wire w_dff_B_CJGC58Sf0_1;
	wire w_dff_B_feXLolQg1_1;
	wire w_dff_B_Cy9ppjHU9_1;
	wire w_dff_B_Boy1qROf5_1;
	wire w_dff_B_aerMXmxU8_1;
	wire w_dff_B_zDDQiLEs8_1;
	wire w_dff_B_qyHnPJs31_1;
	wire w_dff_B_ibo5FJdy2_1;
	wire w_dff_A_MTGAcOxS8_0;
	wire w_dff_A_Dqlxau3C9_0;
	wire w_dff_A_ZyvMiqwv7_0;
	wire w_dff_A_AF5Godks4_0;
	wire w_dff_A_t49iNQX13_0;
	wire w_dff_A_Vou0topv5_0;
	wire w_dff_A_8V5MMddR3_0;
	wire w_dff_A_NDxk09Lm9_0;
	wire w_dff_A_3bqzTno87_0;
	wire w_dff_A_u740gv2z5_0;
	wire w_dff_A_JUX6K2h81_0;
	wire w_dff_A_qiFtbCbr5_0;
	wire w_dff_A_MPJ39nPw9_0;
	wire w_dff_A_1uLbwkqc1_0;
	wire w_dff_A_cnvrGUbq3_0;
	wire w_dff_A_66IuD3qm1_0;
	wire w_dff_A_vcHSnjrt3_0;
	wire w_dff_A_Xol5qGsh0_0;
	wire w_dff_A_Rs6q3HyB2_0;
	wire w_dff_A_7h3mI36C1_0;
	wire w_dff_A_GJNayBME6_0;
	wire w_dff_A_vIIkb0HD7_0;
	wire w_dff_A_WJYgSSeq1_0;
	wire w_dff_A_VidqzFNW6_1;
	wire w_dff_B_f0vyNdGs6_1;
	wire w_dff_B_JFgCKWVc8_1;
	wire w_dff_B_MvkArjkZ4_1;
	wire w_dff_B_QfVfJSCB6_1;
	wire w_dff_B_aWIF8es22_1;
	wire w_dff_B_ay02jxqo6_1;
	wire w_dff_B_dLsXYE3Z5_1;
	wire w_dff_B_zgHnO0sP7_1;
	wire w_dff_B_n4NTiLWU4_1;
	wire w_dff_B_9DF1XkZM9_1;
	wire w_dff_B_6VFewGtb1_1;
	wire w_dff_B_XspO4uMb3_1;
	wire w_dff_B_qyoP1Ca73_1;
	wire w_dff_B_6tf9Yp4V8_1;
	wire w_dff_B_qeR3ms464_1;
	wire w_dff_B_Z2TokshB1_1;
	wire w_dff_B_k3rcn5xi0_1;
	wire w_dff_B_YQ8XFpW90_1;
	wire w_dff_B_qwvf0gmh5_1;
	wire w_dff_B_zvFQplgs5_1;
	wire w_dff_A_DxyQf3yv1_0;
	wire w_dff_A_WGEYsVGX8_0;
	wire w_dff_A_McTraJS24_0;
	wire w_dff_A_sBNH4PME7_0;
	wire w_dff_A_sLsyXSrp2_0;
	wire w_dff_A_a2o728ux5_0;
	wire w_dff_A_uf9mn53k1_0;
	wire w_dff_A_mRaioLGc7_0;
	wire w_dff_A_YpSBvYFC1_0;
	wire w_dff_A_aAAURnAq8_0;
	wire w_dff_A_XCPjNbdl0_0;
	wire w_dff_A_gOyCnO5A1_0;
	wire w_dff_A_4L6LIz1d6_0;
	wire w_dff_A_PoUpHa9o8_0;
	wire w_dff_A_MtB7Ibou8_0;
	wire w_dff_A_slhcY3sp1_0;
	wire w_dff_A_8hqnuJXv0_0;
	wire w_dff_A_teltklyC2_0;
	wire w_dff_A_Nzpx970u6_0;
	wire w_dff_A_r7OMeDpp7_0;
	wire w_dff_A_uk6LQE8m1_1;
	wire w_dff_B_GXZScAZ97_1;
	wire w_dff_B_sNXOD5Te5_1;
	wire w_dff_B_mosPq6Iw7_1;
	wire w_dff_B_DmqVEt9h3_1;
	wire w_dff_B_WqQ9P0BI9_1;
	wire w_dff_B_tYMvDHjF9_1;
	wire w_dff_B_mYvwLHIE3_1;
	wire w_dff_B_jy7V7kH94_1;
	wire w_dff_B_nYSoaTrs1_1;
	wire w_dff_B_I7oXqdZX9_1;
	wire w_dff_B_xjCOxvEJ8_1;
	wire w_dff_B_A0SwQJBz2_1;
	wire w_dff_B_9neIFpWk8_1;
	wire w_dff_B_9kGByPrb8_1;
	wire w_dff_B_KNAIm56a4_1;
	wire w_dff_B_zlTyNM2h9_1;
	wire w_dff_B_0vmM2Dpk6_1;
	wire w_dff_A_RQoc8dDu3_0;
	wire w_dff_A_3UYvoCjL7_0;
	wire w_dff_A_JYJIqle31_0;
	wire w_dff_A_Zam404ga7_0;
	wire w_dff_A_xpaw3GIc3_0;
	wire w_dff_A_qtTvdTNd6_0;
	wire w_dff_A_b0WoWlA55_0;
	wire w_dff_A_ipcMJtvZ3_0;
	wire w_dff_A_lllFJPyA9_0;
	wire w_dff_A_NIXy8Lja8_0;
	wire w_dff_A_XuSvxjEP4_0;
	wire w_dff_A_evmWHlwv5_0;
	wire w_dff_A_sRkSva2B6_0;
	wire w_dff_A_s7YYj71d7_0;
	wire w_dff_A_eI7iRPhF5_0;
	wire w_dff_A_CKC3Yn8f7_0;
	wire w_dff_A_VZPaFjUV4_0;
	wire w_dff_A_jlM84O8q0_1;
	wire w_dff_B_zfuvNCQQ3_1;
	wire w_dff_B_bpvSJBRK9_1;
	wire w_dff_B_7oNspLiC5_1;
	wire w_dff_B_EEACuwh76_1;
	wire w_dff_B_Eu5engjA1_1;
	wire w_dff_B_vQnexihB6_1;
	wire w_dff_B_ILKNcXJf1_1;
	wire w_dff_B_nQtXH1jO1_1;
	wire w_dff_B_8ZTVRIvv5_1;
	wire w_dff_B_xxPN8qXu7_1;
	wire w_dff_B_MfqZ7y0c9_1;
	wire w_dff_B_u1ziF5763_1;
	wire w_dff_B_EHlu3dn94_1;
	wire w_dff_B_NiuiUYAR7_1;
	wire w_dff_A_3morTeKC0_0;
	wire w_dff_A_xHNVvKMT8_0;
	wire w_dff_A_nlkU3F5a8_0;
	wire w_dff_A_YRrVLZFO9_0;
	wire w_dff_A_aTQPuo2u3_0;
	wire w_dff_A_NBLHVlz99_0;
	wire w_dff_A_svvjYLuG6_0;
	wire w_dff_A_8VOR3zpj2_0;
	wire w_dff_A_ev0RHqGZ3_0;
	wire w_dff_A_wHYSETMK7_0;
	wire w_dff_A_VCuonMYy9_0;
	wire w_dff_A_mvCLfD9x0_0;
	wire w_dff_A_syDCTWfq5_0;
	wire w_dff_A_zXoueFPQ6_0;
	wire w_dff_A_t5eeBDnN5_1;
	wire w_dff_B_9xiLlT4y2_1;
	wire w_dff_B_9KRAEmbh7_1;
	wire w_dff_B_ggZTS0gd1_1;
	wire w_dff_B_4LKlCLrA7_1;
	wire w_dff_B_2R25WAQK8_1;
	wire w_dff_B_TppLyg4v4_1;
	wire w_dff_B_9nLxrKgD3_1;
	wire w_dff_B_sNuIyDiq9_1;
	wire w_dff_B_M5kAxx6I7_1;
	wire w_dff_B_owl5xRXF4_1;
	wire w_dff_B_2rxQ8rZv0_1;
	wire w_dff_A_OpndN7z58_0;
	wire w_dff_A_keAsB39M8_0;
	wire w_dff_A_gKgPIvD13_0;
	wire w_dff_A_4cydyGjc7_0;
	wire w_dff_A_udABFOUe6_0;
	wire w_dff_A_CCdgCSaS5_0;
	wire w_dff_A_YRpxcmXh3_0;
	wire w_dff_A_9KFj6Kic7_0;
	wire w_dff_A_fghwch2a5_0;
	wire w_dff_A_fswP8Brl5_0;
	wire w_dff_A_1tP4Ojsj6_0;
	wire w_dff_A_16lnEayP7_1;
	wire w_dff_B_ql0xxNOV8_1;
	wire w_dff_B_yEyi6Bcm2_1;
	wire w_dff_B_dByFWDg89_1;
	wire w_dff_B_3mjKI0g11_1;
	wire w_dff_B_bu9REvml5_1;
	wire w_dff_B_tmlWrp378_1;
	wire w_dff_B_WOKIVqPd1_1;
	wire w_dff_B_uBqySN0o4_1;
	wire w_dff_A_6Iqt84Uz8_0;
	wire w_dff_A_lkj7oKoR0_0;
	wire w_dff_A_RxECoBzC0_0;
	wire w_dff_A_RJrAcvEy5_0;
	wire w_dff_A_sMiz8vT45_0;
	wire w_dff_A_zR5A5U2s7_0;
	wire w_dff_A_ld20n9FH2_0;
	wire w_dff_A_3bc51pMd5_0;
	wire w_dff_A_CTRaqL9B3_1;
	wire w_dff_B_somNRr3K8_1;
	wire w_dff_B_3z8o40fg2_1;
	wire w_dff_B_pGbrx3Wv3_1;
	wire w_dff_B_5uOOUoA52_1;
	wire w_dff_B_3MngmSLX7_1;
	wire w_dff_B_8fabrxSB4_0;
	wire w_dff_A_DuRvFlYK3_0;
	wire w_dff_A_dzP8WDLp8_0;
	wire w_dff_A_XjuzOzbT6_0;
	wire w_dff_A_OePys8Kz6_0;
	wire w_dff_A_yQlDCY0r9_0;
	wire w_dff_A_jVSOrltG9_0;
	wire w_dff_A_qNtSau7H0_0;
	wire w_dff_A_Om9vCIER8_1;
	wire w_dff_B_rxFTLE6m4_1;
	wire w_dff_B_JeJeGQdS0_2;
	wire w_dff_B_eeC0TOx72_2;
	wire w_dff_B_EqNcRvMn0_2;
	wire w_dff_B_sd4iDbTu4_2;
	wire w_dff_B_4JqgDNrV1_2;
	wire w_dff_B_NhZ0ttCJ2_2;
	wire w_dff_B_u1Un5rHB2_2;
	wire w_dff_B_nI3qGxFd2_2;
	wire w_dff_B_HK9IvcZv5_2;
	wire w_dff_B_TY5MJ6X65_2;
	wire w_dff_B_KR9ir9qC3_2;
	wire w_dff_B_hwQDgPLZ3_2;
	wire w_dff_B_KBRszzhj2_2;
	wire w_dff_B_4yDbemdy3_2;
	wire w_dff_B_dU7Dbcac8_2;
	wire w_dff_B_aLJbCdnY1_2;
	wire w_dff_B_pZzzmzNk9_2;
	wire w_dff_B_jFmfJljb9_2;
	wire w_dff_B_y0ggQzps5_2;
	wire w_dff_B_WLtX5I5J0_2;
	wire w_dff_B_Px9ysO1c9_2;
	wire w_dff_B_2NAuces67_2;
	wire w_dff_B_oUs2DGfX2_2;
	wire w_dff_B_B2ynoS7N8_2;
	wire w_dff_B_Gv73NBPG9_2;
	wire w_dff_B_cGbWw0kq6_2;
	wire w_dff_B_hwS2Wrzm3_2;
	wire w_dff_B_T0DtvykX4_2;
	wire w_dff_B_BLzPcQXz2_2;
	wire w_dff_B_lCFiarFR4_2;
	wire w_dff_B_EtTf68cC0_2;
	wire w_dff_B_O675cwWI4_2;
	wire w_dff_B_w3paKbUS7_2;
	wire w_dff_B_4e2zvKBd8_2;
	wire w_dff_B_OsatqXEn2_2;
	wire w_dff_B_6gcFq2qZ4_2;
	wire w_dff_B_43cWqXcJ9_2;
	wire w_dff_B_XmiBbv9O8_2;
	wire w_dff_B_dbi9DG9r0_2;
	wire w_dff_B_cSCjdipF3_2;
	wire w_dff_B_iQbbHtVj4_2;
	wire w_dff_B_3iPC0LYk7_2;
	wire w_dff_B_xWKZTo7M7_2;
	wire w_dff_B_UgomcaYM9_2;
	wire w_dff_A_IYu9QDqv2_0;
	wire w_dff_B_9J9G5dhP3_1;
	wire w_dff_B_TA4DWdGV8_2;
	wire w_dff_B_CLklGeY05_2;
	wire w_dff_B_QyBjJ8Vn9_2;
	wire w_dff_B_wTBYR0hu4_2;
	wire w_dff_B_TfGXVdAR0_2;
	wire w_dff_B_YJqXvrmm9_2;
	wire w_dff_B_k0IZG2Hc4_2;
	wire w_dff_B_LMwbwHTU1_2;
	wire w_dff_B_UGMUiXF57_2;
	wire w_dff_B_AAgdIXzo4_2;
	wire w_dff_B_wKENF1XL0_2;
	wire w_dff_B_ZSJlHGs64_2;
	wire w_dff_B_j4xQdnXq2_2;
	wire w_dff_B_kmFz5Dci2_2;
	wire w_dff_B_sucw9Ygt1_2;
	wire w_dff_B_IfUz4ndu2_2;
	wire w_dff_B_qVy19lph5_2;
	wire w_dff_B_zly0R7qp5_2;
	wire w_dff_B_m7VVN3qx0_2;
	wire w_dff_B_lywSVzBg9_2;
	wire w_dff_B_SqR5ieOD9_2;
	wire w_dff_B_qCfP3pXC0_2;
	wire w_dff_B_Ge9IynTe0_2;
	wire w_dff_B_pHsg5nmV1_2;
	wire w_dff_B_PouuHYAR1_2;
	wire w_dff_B_2BO1y4Tc3_2;
	wire w_dff_B_hqLbpPmL6_2;
	wire w_dff_B_hMjNrgmF9_2;
	wire w_dff_B_A23ukn8M6_2;
	wire w_dff_B_NJyS9AiW9_2;
	wire w_dff_B_QYCS95NF0_2;
	wire w_dff_B_NdiLhKAS4_2;
	wire w_dff_B_E70GJp9W9_2;
	wire w_dff_B_rpYQZu1i4_2;
	wire w_dff_B_ffCQGSql1_2;
	wire w_dff_B_zNG8Nvgp8_2;
	wire w_dff_B_7pssP60b0_2;
	wire w_dff_B_m2SC6Q7j9_2;
	wire w_dff_B_yrfeAPaT5_2;
	wire w_dff_B_JqAG9UCb9_2;
	wire w_dff_B_wO10LduC0_2;
	wire w_dff_A_Oj2QZeXD0_1;
	wire w_dff_B_V0dPnTPX0_1;
	wire w_dff_B_Ji9pX2ES4_1;
	wire w_dff_B_0LUshjrx3_1;
	wire w_dff_B_T8rBcWFe3_1;
	wire w_dff_B_HRWhvgFq4_1;
	wire w_dff_B_fd6niYRp1_1;
	wire w_dff_B_xOW05q3B3_1;
	wire w_dff_B_DfFrf3BO6_1;
	wire w_dff_B_FzFgK3iN0_1;
	wire w_dff_B_UbiBswyu7_1;
	wire w_dff_B_DonOGi5j8_1;
	wire w_dff_B_DVlO2hi82_1;
	wire w_dff_B_sXy64Lbe9_1;
	wire w_dff_B_yA48ylDb6_1;
	wire w_dff_B_WqyKBDO63_1;
	wire w_dff_B_GEvAHh4Q7_1;
	wire w_dff_B_szhGWO7G2_1;
	wire w_dff_B_InNh9hGR3_1;
	wire w_dff_B_deOhBe0D3_1;
	wire w_dff_B_65BZeBJU7_1;
	wire w_dff_B_UTvbge8z0_1;
	wire w_dff_B_E2CMcfpL2_1;
	wire w_dff_B_HoBcODdq0_1;
	wire w_dff_B_xNpdHfJl8_1;
	wire w_dff_B_SJcwfZQ30_1;
	wire w_dff_B_p86gTzkp7_1;
	wire w_dff_B_wCHZHEGk1_1;
	wire w_dff_B_TwMEC49E3_1;
	wire w_dff_B_x1jdbZhI2_1;
	wire w_dff_B_4wxA6eZn4_1;
	wire w_dff_B_pxfrCFT81_1;
	wire w_dff_B_2zceQQ1i8_1;
	wire w_dff_B_9Lah1VMm0_1;
	wire w_dff_B_ASKlD0uT5_1;
	wire w_dff_B_Cb7Bv95w9_1;
	wire w_dff_B_xYDsoEwY9_1;
	wire w_dff_B_sNHx9GFp7_1;
	wire w_dff_B_HWRDEJIq8_1;
	wire w_dff_A_8Ls6SQMY1_0;
	wire w_dff_A_jOD8LKnJ0_0;
	wire w_dff_A_xBUhKTzQ8_0;
	wire w_dff_A_ibTJclNI9_0;
	wire w_dff_A_CQtyuUFf5_0;
	wire w_dff_A_k9P9u1CZ4_0;
	wire w_dff_A_hnt2NgWO6_0;
	wire w_dff_A_Sc62zVqh8_0;
	wire w_dff_A_3RBACpkU1_0;
	wire w_dff_A_zP82B3G82_0;
	wire w_dff_A_nIQTdYas5_0;
	wire w_dff_A_kHK3pD0g0_0;
	wire w_dff_A_LUAWhf7J4_0;
	wire w_dff_A_BTA1JJRI6_0;
	wire w_dff_A_NcKBC49r1_0;
	wire w_dff_A_U36aJKzV6_0;
	wire w_dff_A_LGM7CuMA1_0;
	wire w_dff_A_kX1Zn2fm0_0;
	wire w_dff_A_z5RbAXbL2_0;
	wire w_dff_A_9bIR5dQA7_0;
	wire w_dff_A_c3TXFA8I1_0;
	wire w_dff_A_fhBQCqvb4_0;
	wire w_dff_A_Gwt5aC6M9_0;
	wire w_dff_A_un2q7DOg9_0;
	wire w_dff_A_Fw41wDSs7_0;
	wire w_dff_A_gFL68rjQ3_0;
	wire w_dff_A_lJLprpNW4_0;
	wire w_dff_A_9muuIYZa4_0;
	wire w_dff_A_XDBXbmDU9_0;
	wire w_dff_A_zDsM3TAb9_0;
	wire w_dff_A_BtDzUKUL9_0;
	wire w_dff_A_W2ao1JDL2_0;
	wire w_dff_A_rZmwKjpC6_0;
	wire w_dff_A_FHz3OLs28_0;
	wire w_dff_A_P6mwVooE5_0;
	wire w_dff_A_udAcokyh0_0;
	wire w_dff_A_I6WCFdXQ7_0;
	wire w_dff_A_Bb9hNL731_0;
	wire w_dff_A_ykRVGLmZ7_0;
	wire w_dff_B_3XNwPl930_1;
	wire w_dff_A_V0al9raf3_0;
	wire w_dff_A_p7IMXphc6_0;
	wire w_dff_A_b2PrGeK75_0;
	wire w_dff_A_ok5d407S7_0;
	wire w_dff_A_5Zjy2mMT3_0;
	wire w_dff_A_zHP9eEiN3_0;
	wire w_dff_A_rUsxgoGb9_0;
	wire w_dff_A_UkVNKsnp5_0;
	wire w_dff_A_hzDffdzX1_0;
	wire w_dff_A_WcQP0GVk7_0;
	wire w_dff_A_kJPQVcKW1_0;
	wire w_dff_A_qhnUAuHw9_0;
	wire w_dff_A_oVsqIYz31_0;
	wire w_dff_A_5tCBRLI28_0;
	wire w_dff_A_LNjcHkWh6_0;
	wire w_dff_A_IM2OIQZE5_0;
	wire w_dff_A_F87PH2eY3_0;
	wire w_dff_A_3WGIdDBq0_0;
	wire w_dff_A_GXxg27Sd2_0;
	wire w_dff_A_swUgQyJJ3_0;
	wire w_dff_A_PP0Q3MYf6_0;
	wire w_dff_A_lWUYQwJa5_0;
	wire w_dff_A_XLGvzO3m2_0;
	wire w_dff_A_RCDgZQ4G3_0;
	wire w_dff_A_T5knTiQt4_0;
	wire w_dff_A_2I5mb8x68_0;
	wire w_dff_A_x7BSejfI0_0;
	wire w_dff_A_6fOqBFAZ8_0;
	wire w_dff_A_SueV4pZG8_0;
	wire w_dff_A_a24faCMM5_0;
	wire w_dff_A_oM5fdqOE2_0;
	wire w_dff_A_8D5ntETR4_0;
	wire w_dff_A_MBWUmYwd6_0;
	wire w_dff_A_s3ndbN176_0;
	wire w_dff_A_ovFp6XYL3_0;
	wire w_dff_A_hp903XOU7_0;
	wire w_dff_B_wsW7Faqe1_1;
	wire w_dff_A_dd4K6fuO5_0;
	wire w_dff_A_XpPiGr3x1_0;
	wire w_dff_A_yC0MeDY08_0;
	wire w_dff_A_cGGgTJYQ8_0;
	wire w_dff_A_ukmfKaNG1_0;
	wire w_dff_A_kV8hlzAE2_0;
	wire w_dff_A_8E0wrzOd7_0;
	wire w_dff_A_FGnF1Twi8_0;
	wire w_dff_A_8FWgaAg45_0;
	wire w_dff_A_3IbXwgMp1_0;
	wire w_dff_A_ZLevxzaJ1_0;
	wire w_dff_A_BgRLUtul7_0;
	wire w_dff_A_sg8rqorY3_0;
	wire w_dff_A_fa6nMazo9_0;
	wire w_dff_A_p5UHkiEQ0_0;
	wire w_dff_A_Ye9ch74A0_0;
	wire w_dff_A_spBK6mPB3_0;
	wire w_dff_A_oFRqVpEZ1_0;
	wire w_dff_A_FYQN9leY6_0;
	wire w_dff_A_OeR9mgBf7_0;
	wire w_dff_A_6IydYeZ35_0;
	wire w_dff_A_fpoXmepm6_0;
	wire w_dff_A_QailJnZE4_0;
	wire w_dff_A_PxFHXmx40_0;
	wire w_dff_A_CaQIVJYX8_0;
	wire w_dff_A_qSSv5qNJ3_0;
	wire w_dff_A_lztAnQVH3_0;
	wire w_dff_A_wLoomBFP2_0;
	wire w_dff_A_MoHgFzyH7_0;
	wire w_dff_A_m1KXgRUx1_0;
	wire w_dff_A_TP7SxmJx9_0;
	wire w_dff_A_V61aGOcA3_0;
	wire w_dff_A_8nZPzhWn0_0;
	wire w_dff_B_ceJJ1TqA2_1;
	wire w_dff_A_P6dJldKc0_0;
	wire w_dff_A_x6mkCbD29_0;
	wire w_dff_A_hvsux0TA0_0;
	wire w_dff_A_U6oKz77h8_0;
	wire w_dff_A_2qflyQ9V8_0;
	wire w_dff_A_r3vTuDxT8_0;
	wire w_dff_A_QKav6WDD9_0;
	wire w_dff_A_wotP33kW4_0;
	wire w_dff_A_FYhn0K6s0_0;
	wire w_dff_A_NEr2QcCr4_0;
	wire w_dff_A_fVHvH0Nz1_0;
	wire w_dff_A_W4O9bCZS5_0;
	wire w_dff_A_U8nw2nkM6_0;
	wire w_dff_A_oSDvXZGQ8_0;
	wire w_dff_A_QTqKNitV0_0;
	wire w_dff_A_nzcDwDXq8_0;
	wire w_dff_A_UDeiaAs46_0;
	wire w_dff_A_2y9Kiczx8_0;
	wire w_dff_A_rOYROLLh6_0;
	wire w_dff_A_Aoo1p9QS5_0;
	wire w_dff_A_5CtkRo1O9_0;
	wire w_dff_A_5KCFZhqS6_0;
	wire w_dff_A_XVNGvzzC1_0;
	wire w_dff_A_wyWBpMfD2_0;
	wire w_dff_A_2LZFltMa0_0;
	wire w_dff_A_YI0jEpQn0_0;
	wire w_dff_A_IyPEsJ6c7_0;
	wire w_dff_A_dFHcTdGH8_0;
	wire w_dff_A_CoUUaYe63_0;
	wire w_dff_A_OzxLbf6k9_0;
	wire w_dff_B_gogWROKv2_1;
	wire w_dff_A_v21n0fTZ4_0;
	wire w_dff_A_VILfCfRD9_0;
	wire w_dff_A_XKmlLdVR4_0;
	wire w_dff_A_x92JFB3l0_0;
	wire w_dff_A_pRdAAAwT4_0;
	wire w_dff_A_vKtNUfFu8_0;
	wire w_dff_A_lbrnj7yG3_0;
	wire w_dff_A_7y4nNyga7_0;
	wire w_dff_A_GbCvOvxI3_0;
	wire w_dff_A_sm1ugC7Q9_0;
	wire w_dff_A_BIg1jQKh9_0;
	wire w_dff_A_aK53XAkd9_0;
	wire w_dff_A_kUkYfGiZ6_0;
	wire w_dff_A_uHWkqcUh3_0;
	wire w_dff_A_C9NYpTyg8_0;
	wire w_dff_A_1ZSlr2KI2_0;
	wire w_dff_A_S7ZC8g7x1_0;
	wire w_dff_A_Qgvyx5An0_0;
	wire w_dff_A_2vqSeVJR0_0;
	wire w_dff_A_viXzDErQ3_0;
	wire w_dff_A_kpOJqIyM6_0;
	wire w_dff_A_oEz2Eta81_0;
	wire w_dff_A_bva2DfvG1_0;
	wire w_dff_A_DNk0Tqry6_0;
	wire w_dff_A_VuyPjDBI5_0;
	wire w_dff_A_QtvxpQdK0_0;
	wire w_dff_A_pvQlB12I5_0;
	wire w_dff_B_NRDAfc2w1_1;
	wire w_dff_A_EFaKOvSU7_0;
	wire w_dff_A_F9W2pI9J0_0;
	wire w_dff_A_MKkkEXvY5_0;
	wire w_dff_A_9wQh1g897_0;
	wire w_dff_A_pP0MZyNU7_0;
	wire w_dff_A_dafSOxb04_0;
	wire w_dff_A_SEhsINf50_0;
	wire w_dff_A_x5GVXpIL1_0;
	wire w_dff_A_SMUWz6sn9_0;
	wire w_dff_A_0MaEnKQ37_0;
	wire w_dff_A_uYojGnKC8_0;
	wire w_dff_A_7b83H1by4_0;
	wire w_dff_A_Ub93Ysst8_0;
	wire w_dff_A_yIPqrXrz2_0;
	wire w_dff_A_s33j0M6c0_0;
	wire w_dff_A_u8e92U088_0;
	wire w_dff_A_KjTGQSAi7_0;
	wire w_dff_A_Ohaj9CmS3_0;
	wire w_dff_A_wCqiOfDk2_0;
	wire w_dff_A_nek62cl68_0;
	wire w_dff_A_9rEGXyCu4_0;
	wire w_dff_A_M2X7AVgt9_0;
	wire w_dff_A_wwsr9i9c7_0;
	wire w_dff_A_kU40C3S38_0;
	wire w_dff_B_MxR0tMp03_1;
	wire w_dff_A_FLit4rH82_0;
	wire w_dff_A_mP77Y0bP5_0;
	wire w_dff_A_uxR7mQh25_0;
	wire w_dff_A_XD2yMGAe1_0;
	wire w_dff_A_92gyhUh10_0;
	wire w_dff_A_TmepH2FY5_0;
	wire w_dff_A_Pb1Ua0MB8_0;
	wire w_dff_A_8dbla37a9_0;
	wire w_dff_A_XYdVrmuR4_0;
	wire w_dff_A_430wvDOS2_0;
	wire w_dff_A_AxfoHPAD1_0;
	wire w_dff_A_bCANLyk59_0;
	wire w_dff_A_IQiOv7Kf8_0;
	wire w_dff_A_wHQKoMmj4_0;
	wire w_dff_A_TFEjcWnh6_0;
	wire w_dff_A_OBycHW4B6_0;
	wire w_dff_A_Tdsyh3pk5_0;
	wire w_dff_A_uUK32Z9q1_0;
	wire w_dff_A_DUFK8B177_0;
	wire w_dff_A_OPdTFdsX8_0;
	wire w_dff_A_iWTcsfKo0_0;
	wire w_dff_B_9jqgJuYA5_1;
	wire w_dff_A_gbicxs0O4_0;
	wire w_dff_A_cHAz5HE42_0;
	wire w_dff_A_RrNwHRsJ0_0;
	wire w_dff_A_SWr58CsJ3_0;
	wire w_dff_A_rl4DFSnm6_0;
	wire w_dff_A_vj842KFM7_0;
	wire w_dff_A_vs0t15Ym1_0;
	wire w_dff_A_9njqBmUc0_0;
	wire w_dff_A_fhxewFaJ4_0;
	wire w_dff_A_vtSVeODc7_0;
	wire w_dff_A_GNnBl4sc3_0;
	wire w_dff_A_g5m0mqt44_0;
	wire w_dff_A_pVJcJDce9_0;
	wire w_dff_A_Xe22HY7d1_0;
	wire w_dff_A_DIlmSFjG2_0;
	wire w_dff_A_Mbt6qhLF3_0;
	wire w_dff_A_jgurZwdt9_0;
	wire w_dff_A_6MqYMjVg1_0;
	wire w_dff_B_dAuOBgIL1_1;
	wire w_dff_A_xR1gWTJD2_0;
	wire w_dff_A_F0WIojUQ1_0;
	wire w_dff_A_640Skq8P8_0;
	wire w_dff_A_Nhn8XYwv4_0;
	wire w_dff_A_RFyH1kny0_0;
	wire w_dff_A_LrCsXBUG6_0;
	wire w_dff_A_DBQeq0Fo2_0;
	wire w_dff_A_9mbuu8nP3_0;
	wire w_dff_A_uy2i3tGS0_0;
	wire w_dff_A_eRscqzXf0_0;
	wire w_dff_A_7XGsQS204_0;
	wire w_dff_A_81lRWZBC6_0;
	wire w_dff_A_jTQmQ8Kn5_0;
	wire w_dff_A_ashIQI344_0;
	wire w_dff_A_DPpMOZQn6_0;
	wire w_dff_B_ScOtqCUR0_1;
	wire w_dff_A_pVE7kE5D0_0;
	wire w_dff_A_nXxWpgoZ6_0;
	wire w_dff_A_MbDdXnqq0_0;
	wire w_dff_A_4Vysn0yB1_0;
	wire w_dff_A_AaMmI03z0_0;
	wire w_dff_A_0wW5U7509_0;
	wire w_dff_A_lnPhx0Ix4_0;
	wire w_dff_A_Hmj2pzsU1_0;
	wire w_dff_A_VfvNn8Ru3_0;
	wire w_dff_A_lVMWhBhW4_0;
	wire w_dff_A_Npyp55tc1_0;
	wire w_dff_A_JG8iwnZG5_0;
	wire w_dff_B_6qB0mknv3_1;
	wire w_dff_A_JbFnYCS59_0;
	wire w_dff_A_i1TlMSzT1_0;
	wire w_dff_A_55wZ5YOo2_0;
	wire w_dff_A_LYe7BlVf2_0;
	wire w_dff_A_e6xyxHaw5_0;
	wire w_dff_A_RryRbKAU6_0;
	wire w_dff_A_zBfqEmkV3_0;
	wire w_dff_A_t8goGsCr9_0;
	wire w_dff_A_1LCq0UX68_0;
	wire w_dff_A_IGVxKSBU0_0;
	wire w_dff_A_zA7efneb1_0;
	wire w_dff_A_wzFeeiny6_1;
	wire w_dff_A_8wOEl3lt9_0;
	wire w_dff_A_gxb0Kmdb6_0;
	wire w_dff_A_LRuQbPIa4_0;
	wire w_dff_A_BmzAGfJI1_0;
	wire w_dff_A_o96JgnLg3_0;
	wire w_dff_A_GRJDodBM4_0;
	wire w_dff_A_ULikrVqh5_0;
	wire w_dff_B_GllUaxUV7_1;
	wire w_dff_A_2wtDOQkA6_1;
	wire w_dff_A_X3OPPVNu9_2;
	wire w_dff_A_isb7tLK02_2;
	wire w_dff_A_1qgBAHnM3_0;
	wire w_dff_B_BmLhtFuJ1_2;
	wire w_dff_B_ocyQzzZ21_2;
	wire w_dff_B_rlT6IMnw4_2;
	wire w_dff_B_S06AnL1I2_2;
	wire w_dff_B_GVqKwmtX8_2;
	wire w_dff_B_a2AGywqX0_2;
	wire w_dff_B_wPdW3wBw0_2;
	wire w_dff_B_FOn5djG20_2;
	wire w_dff_B_MuIMJzik6_2;
	wire w_dff_B_t4louVvR6_2;
	wire w_dff_B_8M1DNNVT9_2;
	wire w_dff_B_WMtLWxSR4_2;
	wire w_dff_B_D2hovTJA7_2;
	wire w_dff_B_AiX9Q5Fi9_2;
	wire w_dff_B_fxczt5X34_2;
	wire w_dff_B_HikhZ2YX1_2;
	wire w_dff_B_eaS9SxWf4_2;
	wire w_dff_B_ToWGlZ6L7_2;
	wire w_dff_B_XqaD1iUu4_2;
	wire w_dff_B_iMY4XgAd2_2;
	wire w_dff_B_ccy3aQBn2_2;
	wire w_dff_B_8mRcifVg1_2;
	wire w_dff_B_Vtzj9JXw7_2;
	wire w_dff_B_NgY4FC6y5_2;
	wire w_dff_B_jPjNxvub3_2;
	wire w_dff_B_jW6skY2Y9_2;
	wire w_dff_B_Mlb2ZzGS0_2;
	wire w_dff_B_0qcN5Jcl8_2;
	wire w_dff_B_02whfXKO2_2;
	wire w_dff_B_yii16jwC2_2;
	wire w_dff_B_hlyFtVtZ3_2;
	wire w_dff_B_Yx4TN7v45_2;
	wire w_dff_B_Sj6uyHAj9_2;
	wire w_dff_B_ODy9GZzg9_2;
	wire w_dff_B_N1ACvKMH5_2;
	wire w_dff_B_fl60HsEZ2_2;
	wire w_dff_B_pAuD7G3b6_2;
	wire w_dff_B_ErWk5laX0_2;
	wire w_dff_B_XZjISiha4_2;
	wire w_dff_B_UUXTOPCD8_2;
	wire w_dff_B_dHfnf7lJ6_2;
	wire w_dff_B_fFjd9uOZ2_2;
	wire w_dff_B_ttZn8Y1j7_2;
	wire w_dff_B_q4ru4Yif6_2;
	wire w_dff_B_aZrjLaUP2_2;
	wire w_dff_A_kLeTUCqx2_0;
	wire w_dff_B_UWPl9sBx1_1;
	wire w_dff_B_6VcU4rsP4_2;
	wire w_dff_B_xXkI68eK1_2;
	wire w_dff_B_j32ADvOg1_2;
	wire w_dff_B_apGrgngt8_2;
	wire w_dff_B_SbNGzs4J6_2;
	wire w_dff_B_03NIjkI52_2;
	wire w_dff_B_bCRIOj3k1_2;
	wire w_dff_B_C8OKsyJY5_2;
	wire w_dff_B_yFH92Y7X3_2;
	wire w_dff_B_LRDRYvPu5_2;
	wire w_dff_B_EROViqrh7_2;
	wire w_dff_B_TPUpIvki3_2;
	wire w_dff_B_DEg7uwmr2_2;
	wire w_dff_B_is3IUrvB0_2;
	wire w_dff_B_vWBpL7ha8_2;
	wire w_dff_B_jvzpxm137_2;
	wire w_dff_B_HSCV1UZj3_2;
	wire w_dff_B_kbidfiAl4_2;
	wire w_dff_B_FmCeQ5XW9_2;
	wire w_dff_B_hGAzrKfH0_2;
	wire w_dff_B_sRsis2oF1_2;
	wire w_dff_B_RrRBUQwa0_2;
	wire w_dff_B_JECTympL4_2;
	wire w_dff_B_UH5Pltlm0_2;
	wire w_dff_B_RsuIk8EJ6_2;
	wire w_dff_B_VBB7XORv4_2;
	wire w_dff_B_Mh2uFYUk4_2;
	wire w_dff_B_e2dKciYF1_2;
	wire w_dff_B_HW40Zgwk5_2;
	wire w_dff_B_hlq2KFZ66_2;
	wire w_dff_B_d1iyb83h8_2;
	wire w_dff_B_o4lWT9hn1_2;
	wire w_dff_B_jYBENLzS3_2;
	wire w_dff_B_L7mBxDtg2_2;
	wire w_dff_B_AcX11O4H3_2;
	wire w_dff_B_BtUbDKoU7_2;
	wire w_dff_B_wEF0KkXg4_2;
	wire w_dff_B_u2KJDh9v3_2;
	wire w_dff_B_wG1EELJS9_2;
	wire w_dff_B_C6GIKeOi4_2;
	wire w_dff_B_OlErDkei0_2;
	wire w_dff_A_rzHhCtPL6_1;
	wire w_dff_A_sfvkaepl4_0;
	wire w_dff_A_j09C3lLo8_0;
	wire w_dff_A_tHCBWyJb3_0;
	wire w_dff_A_55kyTyUN6_0;
	wire w_dff_A_NkHF0lWc3_0;
	wire w_dff_A_GL9lb41z9_0;
	wire w_dff_A_u5qBhXCf2_0;
	wire w_dff_A_Xurl298G2_0;
	wire w_dff_A_0r240fVN2_0;
	wire w_dff_A_iHrnoSBO6_0;
	wire w_dff_A_gRMC4qa37_0;
	wire w_dff_A_NiK3pdK10_0;
	wire w_dff_A_POaw8Ohg6_0;
	wire w_dff_A_ziWenKew8_0;
	wire w_dff_A_Z54ryrHP1_0;
	wire w_dff_A_DdlyYtEd5_0;
	wire w_dff_A_xmNPZfBT7_0;
	wire w_dff_A_axi8cN4E5_0;
	wire w_dff_A_neikj1IE3_0;
	wire w_dff_A_csYina3v8_0;
	wire w_dff_A_oW39yD0f9_0;
	wire w_dff_A_QbXBvsLp1_0;
	wire w_dff_A_ghnwqKhI1_0;
	wire w_dff_A_2LDLtKfd4_0;
	wire w_dff_A_I4C6SkdQ7_0;
	wire w_dff_A_ThYMcMxK0_0;
	wire w_dff_A_yfPUh4IJ2_0;
	wire w_dff_A_WCTDRuKu5_0;
	wire w_dff_A_XcFEmsJT1_0;
	wire w_dff_A_vNu79JpS6_0;
	wire w_dff_A_ImD6d5LR1_0;
	wire w_dff_A_OOiy5AA68_0;
	wire w_dff_A_E9MTsjz49_0;
	wire w_dff_A_nbq3ehR25_0;
	wire w_dff_A_NWSDKE085_0;
	wire w_dff_A_uKNqnDtx9_0;
	wire w_dff_A_8X035g628_0;
	wire w_dff_A_8g1bLN284_0;
	wire w_dff_A_3epEYrKA2_1;
	wire w_dff_A_axzWNOhv0_2;
	wire w_dff_B_KML9lAql1_1;
	wire w_dff_B_HMGSGBSP1_2;
	wire w_dff_B_viWuZVKu5_2;
	wire w_dff_B_2Ip3rDe58_2;
	wire w_dff_B_3f3pOnVF1_2;
	wire w_dff_B_E1cjXEZG9_2;
	wire w_dff_B_CgVBLYsv9_2;
	wire w_dff_B_ef0mOmRk2_2;
	wire w_dff_B_VPO8kEh80_2;
	wire w_dff_B_tnCHmtY43_2;
	wire w_dff_B_NFqTWkbm1_2;
	wire w_dff_B_4vm3ZSHt4_2;
	wire w_dff_B_jCJebprb0_2;
	wire w_dff_B_5g4GjFHb2_2;
	wire w_dff_B_GmQejb4D7_2;
	wire w_dff_B_tmAxVij19_2;
	wire w_dff_B_Eo0JXkHB4_2;
	wire w_dff_B_hnZ2YC053_2;
	wire w_dff_B_v4KJ7nUd5_2;
	wire w_dff_B_1fYsJQyi3_2;
	wire w_dff_B_Zo9Rq65i6_2;
	wire w_dff_B_DawQzYpX3_2;
	wire w_dff_B_ckZuosHW4_2;
	wire w_dff_B_HEYw3L3e2_2;
	wire w_dff_B_vwTgl1Pe5_2;
	wire w_dff_B_S3tY8KDi6_2;
	wire w_dff_B_orX2KXrt7_2;
	wire w_dff_B_m7CL91jd0_2;
	wire w_dff_B_exGLuhs23_2;
	wire w_dff_B_GVhOx6UT8_2;
	wire w_dff_B_thoognot0_2;
	wire w_dff_B_76CJ4OMI8_2;
	wire w_dff_B_vPIU9umq5_2;
	wire w_dff_B_t2YhdeBC0_2;
	wire w_dff_B_X2BvY5948_2;
	wire w_dff_B_0o7XpGAz9_2;
	wire w_dff_B_f52rD6cQ1_1;
	wire w_dff_B_Ez3ezwi98_2;
	wire w_dff_B_DsaySTek7_2;
	wire w_dff_B_pASD9vDS0_2;
	wire w_dff_B_i545mfNE5_2;
	wire w_dff_B_TEQPCNfb2_2;
	wire w_dff_B_QLoZTlQL2_2;
	wire w_dff_B_gXzPuCI46_2;
	wire w_dff_B_MZSskENs3_2;
	wire w_dff_B_EbkmuCLV9_2;
	wire w_dff_B_uRNj2x3J9_2;
	wire w_dff_B_GYlkhpAa9_2;
	wire w_dff_B_wQbd0lRN8_2;
	wire w_dff_B_5iSkpzgT3_2;
	wire w_dff_B_85IqjXRi8_2;
	wire w_dff_B_D8MWlv167_2;
	wire w_dff_B_qcfRUw7a2_2;
	wire w_dff_B_KnYwV7Ie8_2;
	wire w_dff_B_nY1BbMpL2_2;
	wire w_dff_B_xUBq8LUz9_2;
	wire w_dff_B_2L2fDyKB8_2;
	wire w_dff_B_mpkc6BD26_2;
	wire w_dff_B_fJUf09Y04_2;
	wire w_dff_B_aCiqBmLW9_2;
	wire w_dff_B_EhWBx6Cq5_2;
	wire w_dff_B_bwI9yltF0_2;
	wire w_dff_B_Cp9nh4yP6_2;
	wire w_dff_B_6KF8uVbC1_2;
	wire w_dff_B_Inpf2ij73_2;
	wire w_dff_B_asRicJ5x4_2;
	wire w_dff_B_KWMNtjam0_2;
	wire w_dff_B_69glCq6x7_2;
	wire w_dff_B_G3QqpJfF0_2;
	wire w_dff_B_X9AQeE1F8_1;
	wire w_dff_B_Srme0Lsp1_2;
	wire w_dff_B_MCA5sysm1_2;
	wire w_dff_B_JC33sl7w7_2;
	wire w_dff_B_MESuZzuJ8_2;
	wire w_dff_B_UYbyn5cS6_2;
	wire w_dff_B_0bZi3Wt47_2;
	wire w_dff_B_MV0H9icV7_2;
	wire w_dff_B_c9VWh5OX0_2;
	wire w_dff_B_rXITN77F3_2;
	wire w_dff_B_wUOv5E3n4_2;
	wire w_dff_B_wlul32NE4_2;
	wire w_dff_B_l6YuJYHl6_2;
	wire w_dff_B_MISHKE7b1_2;
	wire w_dff_B_tbDNQlhJ1_2;
	wire w_dff_B_6DlFXdW13_2;
	wire w_dff_B_jrn2BW7N3_2;
	wire w_dff_B_opw29W1Y4_2;
	wire w_dff_B_sKks8iMG7_2;
	wire w_dff_B_EAIjP8xk8_2;
	wire w_dff_B_ksWvyQwx3_2;
	wire w_dff_B_QcLFNgqx4_2;
	wire w_dff_B_A2PWGXGY4_2;
	wire w_dff_B_SKACZcwk2_2;
	wire w_dff_B_8Ade8wf23_2;
	wire w_dff_B_AiBGui6H6_2;
	wire w_dff_B_xZoxIi9v4_2;
	wire w_dff_B_bx3pvt1y4_2;
	wire w_dff_B_OO7HPbty9_2;
	wire w_dff_B_WD6Ur2R19_2;
	wire w_dff_B_zFuVlLZs2_1;
	wire w_dff_B_fWL7QoAV2_2;
	wire w_dff_B_NrMuFbNg8_2;
	wire w_dff_B_614uzick1_2;
	wire w_dff_B_1TKcZNRU7_2;
	wire w_dff_B_Ak6k3QKo9_2;
	wire w_dff_B_9s2dY15T7_2;
	wire w_dff_B_49VkbSUp9_2;
	wire w_dff_B_d6MHqYF23_2;
	wire w_dff_B_JeWNfWkH0_2;
	wire w_dff_B_srGNjmG24_2;
	wire w_dff_B_x9Ddx2Xm5_2;
	wire w_dff_B_3TTVyZJ61_2;
	wire w_dff_B_id4z2nxo8_2;
	wire w_dff_B_hOGl5MEE6_2;
	wire w_dff_B_dx61HIkF0_2;
	wire w_dff_B_EdzsSPAA7_2;
	wire w_dff_B_zarxGLFy5_2;
	wire w_dff_B_GnEUns0H7_2;
	wire w_dff_B_HvH16jII8_2;
	wire w_dff_B_VwjtGjNL9_2;
	wire w_dff_B_HUK9nZOo4_2;
	wire w_dff_B_RUlh8mkv9_2;
	wire w_dff_B_y449ZoZd7_2;
	wire w_dff_B_qTjIi8T84_2;
	wire w_dff_B_ukBH0eR21_2;
	wire w_dff_B_PlMEJB0o9_2;
	wire w_dff_B_cQqrFy9q4_1;
	wire w_dff_B_oGXZN2S17_2;
	wire w_dff_B_dcmPLmwV5_2;
	wire w_dff_B_OY363PeA3_2;
	wire w_dff_B_84f9GGzJ0_2;
	wire w_dff_B_wTdFwfpJ7_2;
	wire w_dff_B_afeorywH9_2;
	wire w_dff_B_qEeyTEU21_2;
	wire w_dff_B_hmjmKlc68_2;
	wire w_dff_B_hfJE7aeS1_2;
	wire w_dff_B_SEGgKQXj4_2;
	wire w_dff_B_YSbcQQLq3_2;
	wire w_dff_B_Z1dCurid3_2;
	wire w_dff_B_8nG992SQ6_2;
	wire w_dff_B_DupaHDwX9_2;
	wire w_dff_B_MrsWqR4A0_2;
	wire w_dff_B_DTPpgtrK7_2;
	wire w_dff_B_AqPc4pSF0_2;
	wire w_dff_B_AN0G1K7T0_2;
	wire w_dff_B_PPoL0E3m5_2;
	wire w_dff_B_bnRtv1O20_2;
	wire w_dff_B_5oHCXnj42_2;
	wire w_dff_B_vJ5JRxYC2_2;
	wire w_dff_B_Moc7km7x7_2;
	wire w_dff_B_vkyvK0Dy8_1;
	wire w_dff_B_YDiGq3YV8_2;
	wire w_dff_B_1fbf1D4U9_2;
	wire w_dff_B_OGMxSz1Z2_2;
	wire w_dff_B_1NxLQ00i4_2;
	wire w_dff_B_5onlD2pa3_2;
	wire w_dff_B_PQcHEGID9_2;
	wire w_dff_B_9CQLLmy53_2;
	wire w_dff_B_WSfaPRf54_2;
	wire w_dff_B_8IVexXC99_2;
	wire w_dff_B_CwI58KiC7_2;
	wire w_dff_B_1alBs9ag3_2;
	wire w_dff_B_sRYweDbj3_2;
	wire w_dff_B_gwIHCuXq4_2;
	wire w_dff_B_O8NHjyGe1_2;
	wire w_dff_B_tn5qo77Q2_2;
	wire w_dff_B_2qljnYKr5_2;
	wire w_dff_B_6lOs4cgo8_2;
	wire w_dff_B_ei6UQS5s0_2;
	wire w_dff_B_InpKIDaf8_2;
	wire w_dff_B_Cv00onWb5_2;
	wire w_dff_B_KohjZSWe6_1;
	wire w_dff_B_9RCnqk8y0_2;
	wire w_dff_B_kkfzAReT7_2;
	wire w_dff_B_8dxjvqVf7_2;
	wire w_dff_B_Ktm2YA779_2;
	wire w_dff_B_f58Lg4jI1_2;
	wire w_dff_B_3xP7YiDt0_2;
	wire w_dff_B_MjApJ2Ef2_2;
	wire w_dff_B_RYj4j7GR7_2;
	wire w_dff_B_JN8Rmjbu0_2;
	wire w_dff_B_Zwgq2YQn4_2;
	wire w_dff_B_Qvv4S3gL1_2;
	wire w_dff_B_tXkMbQqq4_2;
	wire w_dff_B_ItELkwND8_2;
	wire w_dff_B_7emjLOGz8_2;
	wire w_dff_B_San30miK3_2;
	wire w_dff_B_KvgfoixZ0_2;
	wire w_dff_B_otGOyUp50_2;
	wire w_dff_B_93cARDKC8_1;
	wire w_dff_B_0zxOQWab8_2;
	wire w_dff_B_NB1dVVAN1_2;
	wire w_dff_B_TY4KntTa0_2;
	wire w_dff_B_1uek05gj7_2;
	wire w_dff_B_nB2cmqc60_2;
	wire w_dff_B_BFGcQ4OJ9_2;
	wire w_dff_B_9pq8nSal8_2;
	wire w_dff_B_i2pGKpnn3_2;
	wire w_dff_B_XQCe5YRT3_2;
	wire w_dff_B_OlLvvtdM3_2;
	wire w_dff_B_ddhbREas5_2;
	wire w_dff_B_lDmu6JHi8_2;
	wire w_dff_B_z2IB3KoP5_2;
	wire w_dff_B_lNc23o2r7_2;
	wire w_dff_B_Q7T7t4QA3_1;
	wire w_dff_B_d10n6hdY6_2;
	wire w_dff_B_vwJ3UIP02_2;
	wire w_dff_B_kCJ6zncB5_2;
	wire w_dff_B_sQywHaUr9_2;
	wire w_dff_B_pbbOhqe95_2;
	wire w_dff_B_TdgP8NmY8_2;
	wire w_dff_B_fZMRQ7B03_2;
	wire w_dff_B_8WR5SiN83_2;
	wire w_dff_B_SWtnxoTH5_2;
	wire w_dff_B_SL8ZdoEa6_2;
	wire w_dff_B_BwpPDbDd4_2;
	wire w_dff_B_rb5e9BaE9_1;
	wire w_dff_B_93yd9Np29_2;
	wire w_dff_B_KNPyR0fw0_2;
	wire w_dff_B_VUCyno7I9_2;
	wire w_dff_B_ByoylkFx9_2;
	wire w_dff_B_FKoK8ueI5_2;
	wire w_dff_B_wHPEqHOf6_2;
	wire w_dff_B_6WHuhTtx4_2;
	wire w_dff_B_CZmZ4Z1s3_2;
	wire w_dff_B_C0xixdSd6_1;
	wire w_dff_B_CJuuASMf2_1;
	wire w_dff_B_TFIA9FbN7_2;
	wire w_dff_B_nx8LWBXN6_2;
	wire w_dff_B_7FwG0O9p1_2;
	wire w_dff_B_LmbkEhOm2_2;
	wire w_dff_A_kaDeBZSS5_1;
	wire w_dff_A_jIE5RpNV8_0;
	wire w_dff_A_wRGR6vxt7_0;
	wire w_dff_A_IqkzQ5Xs0_1;
	wire w_dff_A_iZRBN08a4_2;
	wire w_dff_A_Z0PxXlJi4_2;
	wire w_dff_B_urI1xCRA6_0;
	wire w_dff_A_9iBBkNyV8_1;
	wire w_dff_A_YmfkltVR9_1;
	wire w_dff_B_X81WlWxz2_1;
	wire w_dff_B_RMb7G1lh3_1;
	wire w_dff_B_jhpcgWXj2_2;
	wire w_dff_B_EcjBM6v66_2;
	wire w_dff_B_MzH7DKhg3_2;
	wire w_dff_B_uzJEh9QK8_2;
	wire w_dff_B_fwHIOZsQ5_2;
	wire w_dff_B_TzEie9ks1_2;
	wire w_dff_B_I9yRw00K5_2;
	wire w_dff_B_feK24Jrs0_2;
	wire w_dff_B_55uPTe7i2_2;
	wire w_dff_B_R1CqWste0_2;
	wire w_dff_B_09BZpA1C9_2;
	wire w_dff_B_s6E45NDp1_2;
	wire w_dff_B_UcicT4r90_2;
	wire w_dff_B_0oW87VPB8_2;
	wire w_dff_B_D2OBaIQS0_2;
	wire w_dff_B_wm7YZmGz4_2;
	wire w_dff_B_SqgLxptV8_2;
	wire w_dff_B_M49xPGwf2_2;
	wire w_dff_B_f6DXcH6h7_2;
	wire w_dff_B_0OHa1wGY5_2;
	wire w_dff_B_Hygmnn8X4_2;
	wire w_dff_B_5BfroobQ8_2;
	wire w_dff_B_gac5Wmuo4_2;
	wire w_dff_B_M0PEp5102_2;
	wire w_dff_B_3gsk11nK3_2;
	wire w_dff_B_rY1cNEMX2_2;
	wire w_dff_B_1vGEAePT3_2;
	wire w_dff_B_f3np73zH5_2;
	wire w_dff_B_iDjT3xKg4_2;
	wire w_dff_B_eNsimHCv9_2;
	wire w_dff_B_LQ0INL6c9_2;
	wire w_dff_B_x27H9P4l9_2;
	wire w_dff_B_oXeVwatv8_2;
	wire w_dff_B_qlOvGnHU8_2;
	wire w_dff_B_d7us3JCG8_2;
	wire w_dff_B_tZXwgX9O2_2;
	wire w_dff_B_ecgv8P0H5_2;
	wire w_dff_B_7SBnluyj4_2;
	wire w_dff_B_jCILsPOp8_2;
	wire w_dff_B_4UOyRuZP9_2;
	wire w_dff_B_dkaREQ6B8_2;
	wire w_dff_B_xiS8vVXY8_2;
	wire w_dff_B_mfTSQzP12_2;
	wire w_dff_B_6M2XYg5C5_2;
	wire w_dff_B_HyFIu3p40_2;
	wire w_dff_B_OFFb5aQu2_2;
	wire w_dff_B_QyiOm4660_2;
	wire w_dff_B_SnrhP7B65_1;
	wire w_dff_B_iNMnHjWV0_2;
	wire w_dff_B_5HjPxClh0_2;
	wire w_dff_B_OMV4n6lG3_2;
	wire w_dff_B_hXRvGQNO1_2;
	wire w_dff_B_0kH68DPw6_2;
	wire w_dff_B_15w2wBG63_2;
	wire w_dff_B_scZFHE220_2;
	wire w_dff_B_bmzkcFqB3_2;
	wire w_dff_B_FcHGVivP9_2;
	wire w_dff_B_T5T2sVXp3_2;
	wire w_dff_B_zuMkanZg0_2;
	wire w_dff_B_waRBfHkp0_2;
	wire w_dff_B_O2HnyURc9_2;
	wire w_dff_B_r8YJhsfO0_2;
	wire w_dff_B_0yELmqbw9_2;
	wire w_dff_B_uq6Sipvg6_2;
	wire w_dff_B_n2ALeWO01_2;
	wire w_dff_B_LUnbG5p03_2;
	wire w_dff_B_W1xe0KwH4_2;
	wire w_dff_B_6kZjZzGb6_2;
	wire w_dff_B_SNG295vV5_2;
	wire w_dff_B_gRNLXhAW7_2;
	wire w_dff_B_Rsmzu8z67_2;
	wire w_dff_B_wHxO7Paz8_2;
	wire w_dff_B_gRYISlmU2_2;
	wire w_dff_B_lLJ5ZAtj5_2;
	wire w_dff_B_3JQvdVkT6_2;
	wire w_dff_B_uWdZWg122_2;
	wire w_dff_B_6wqui3nG3_2;
	wire w_dff_B_FmUM072u5_2;
	wire w_dff_B_WbZHUZFl1_2;
	wire w_dff_B_Yf8cyQ189_2;
	wire w_dff_B_vJf8brBr6_2;
	wire w_dff_B_3xVWWNr32_2;
	wire w_dff_B_HXsqowzj6_2;
	wire w_dff_B_b2t2bj9c2_2;
	wire w_dff_B_xkpS3onQ1_2;
	wire w_dff_B_8F4401XA9_2;
	wire w_dff_B_3ys7jXIa3_2;
	wire w_dff_B_1D5F9tCx2_2;
	wire w_dff_B_1ePHcbk11_2;
	wire w_dff_B_AbRIsUjF5_2;
	wire w_dff_B_rdvUAVGU5_2;
	wire w_dff_B_meIcJku66_1;
	wire w_dff_B_eqQbwuD19_2;
	wire w_dff_B_7ZEhjk2q5_2;
	wire w_dff_B_Mhh4rQ9h0_2;
	wire w_dff_B_Ky6pV3WL6_2;
	wire w_dff_B_T0ZUg2d78_2;
	wire w_dff_B_DZX70JOu0_2;
	wire w_dff_B_iRPohZZU0_2;
	wire w_dff_B_k8TgaVrf1_2;
	wire w_dff_B_TRonZ1RH1_2;
	wire w_dff_B_nmb0H0LR2_2;
	wire w_dff_B_6PKRvAUd2_2;
	wire w_dff_B_NkxEajnw3_2;
	wire w_dff_B_02xyN4cw8_2;
	wire w_dff_B_ViQZTLPK3_2;
	wire w_dff_B_SUAiV7wt4_2;
	wire w_dff_B_QvBLEJa96_2;
	wire w_dff_B_sOd6C8IF1_2;
	wire w_dff_B_HmjaLFUn7_2;
	wire w_dff_B_9iBz9BZr0_2;
	wire w_dff_B_Br0IU2by3_2;
	wire w_dff_B_SLRbH0SZ3_2;
	wire w_dff_B_akP5Pr0z6_2;
	wire w_dff_B_i98bKQRl3_2;
	wire w_dff_B_sLw84q5N1_2;
	wire w_dff_B_oGgnWCGX6_2;
	wire w_dff_B_2hc1pEix2_2;
	wire w_dff_B_RizyaOpd5_2;
	wire w_dff_B_UmSXSHi78_2;
	wire w_dff_B_oSXyEGlP8_2;
	wire w_dff_B_PiAyqK7i8_2;
	wire w_dff_B_FGcdhoVp0_2;
	wire w_dff_B_QrRRimLK3_2;
	wire w_dff_B_o7DzriGY2_2;
	wire w_dff_B_pcx0bA3k5_2;
	wire w_dff_B_CmIl0sOT2_2;
	wire w_dff_B_D6a944kG4_2;
	wire w_dff_B_AHIF6KrI3_2;
	wire w_dff_B_m3dEVGtb0_2;
	wire w_dff_B_mILTqqt04_1;
	wire w_dff_B_stFAc2Bj6_2;
	wire w_dff_B_AJ5NI2ek9_2;
	wire w_dff_B_zgHu8R7O3_2;
	wire w_dff_B_V5qaQwey2_2;
	wire w_dff_B_ab4FaQyv0_2;
	wire w_dff_B_uJUWv9AP1_2;
	wire w_dff_B_bWnqCw5C6_2;
	wire w_dff_B_PaWFGgsD9_2;
	wire w_dff_B_8Rvi8o8v8_2;
	wire w_dff_B_8xmQrgpQ3_2;
	wire w_dff_B_NjSlqKvw5_2;
	wire w_dff_B_zKfxGX9u6_2;
	wire w_dff_B_uyj7bbH26_2;
	wire w_dff_B_Ix0kHojs9_2;
	wire w_dff_B_HiZ5F0NJ0_2;
	wire w_dff_B_qQjwxNPs8_2;
	wire w_dff_B_9mPjWmwy7_2;
	wire w_dff_B_PzFpS3aL9_2;
	wire w_dff_B_IW8xLLZV9_2;
	wire w_dff_B_tWWScgaR0_2;
	wire w_dff_B_QjwAqWEO9_2;
	wire w_dff_B_lztXbDZL0_2;
	wire w_dff_B_lO9uSmIZ2_2;
	wire w_dff_B_gM7O6HhC5_2;
	wire w_dff_B_YeQYBF960_2;
	wire w_dff_B_A404kjfF5_2;
	wire w_dff_B_WgbQywpY3_2;
	wire w_dff_B_SElweEU06_2;
	wire w_dff_B_6DmLUu9r0_2;
	wire w_dff_B_hEL1jvx86_2;
	wire w_dff_B_nn9nDP6E8_2;
	wire w_dff_B_FEd5SPu67_2;
	wire w_dff_B_QULM0WWm1_2;
	wire w_dff_B_jU74dILT4_2;
	wire w_dff_B_7XoFcijs1_2;
	wire w_dff_B_zyKCsiWb0_1;
	wire w_dff_B_We9Z8XBh8_2;
	wire w_dff_B_mdNiJjxS3_2;
	wire w_dff_B_p9xagXVH9_2;
	wire w_dff_B_9YjJxp4u5_2;
	wire w_dff_B_KYKnToLb7_2;
	wire w_dff_B_J254yehR8_2;
	wire w_dff_B_1XtR4fN54_2;
	wire w_dff_B_v1FinV3Y0_2;
	wire w_dff_B_vOF6JRXL2_2;
	wire w_dff_B_LsNQSsFU8_2;
	wire w_dff_B_mky0OAFw7_2;
	wire w_dff_B_qIioBpRo0_2;
	wire w_dff_B_1aYFacmk1_2;
	wire w_dff_B_JDyPD08J4_2;
	wire w_dff_B_RlB8V2kd5_2;
	wire w_dff_B_aqMNWGO69_2;
	wire w_dff_B_pUn6F2fF2_2;
	wire w_dff_B_2WaI5Fi15_2;
	wire w_dff_B_kKOUUeLy4_2;
	wire w_dff_B_xUUM9IQG0_2;
	wire w_dff_B_l4cFAL2j9_2;
	wire w_dff_B_OBvKMMPj5_2;
	wire w_dff_B_aAv4rUYN1_2;
	wire w_dff_B_xDnmvA5n8_2;
	wire w_dff_B_P0N2xsry4_2;
	wire w_dff_B_ejzxZOMW8_2;
	wire w_dff_B_lJscurRa6_2;
	wire w_dff_B_kBwr3cgl3_2;
	wire w_dff_B_8ASJgFOC1_2;
	wire w_dff_B_keIzBWij9_2;
	wire w_dff_B_98cUKTy00_2;
	wire w_dff_B_WcmNniVo7_2;
	wire w_dff_B_Jrwnh8Ov3_1;
	wire w_dff_B_f00ZAlqR5_2;
	wire w_dff_B_yqK1LtDd4_2;
	wire w_dff_B_nP5fgjlh6_2;
	wire w_dff_B_AX33OKgJ0_2;
	wire w_dff_B_oBrERymj0_2;
	wire w_dff_B_tp3C8vCo8_2;
	wire w_dff_B_XEShJlEV0_2;
	wire w_dff_B_uDKTL3zM7_2;
	wire w_dff_B_CGADboC25_2;
	wire w_dff_B_ji3YnJRP1_2;
	wire w_dff_B_Fk6tUKYK7_2;
	wire w_dff_B_gzq3zFZ36_2;
	wire w_dff_B_0pJMLwpF8_2;
	wire w_dff_B_1HH0YJwX0_2;
	wire w_dff_B_AdOsjWVc7_2;
	wire w_dff_B_n8hsLvsJ5_2;
	wire w_dff_B_bw8R6iq72_2;
	wire w_dff_B_8rQg8CkI4_2;
	wire w_dff_B_npgGVab36_2;
	wire w_dff_B_DHoi7CfD6_2;
	wire w_dff_B_Wlbn5PPV2_2;
	wire w_dff_B_ZtaRnt5t4_2;
	wire w_dff_B_PVi658TA6_2;
	wire w_dff_B_OX7rEuTv8_2;
	wire w_dff_B_wlGdNU8N8_2;
	wire w_dff_B_DwIRPnk66_2;
	wire w_dff_B_gRlJwIzp3_2;
	wire w_dff_B_YybAkBW14_2;
	wire w_dff_B_5HHz45KX0_2;
	wire w_dff_B_k3h97Z802_1;
	wire w_dff_B_Zhfs6oPJ0_2;
	wire w_dff_B_r4oaUgYX9_2;
	wire w_dff_B_pPeQXJGT4_2;
	wire w_dff_B_QulQVZjg9_2;
	wire w_dff_B_KOPuALy08_2;
	wire w_dff_B_adQbcNVJ6_2;
	wire w_dff_B_X32gJhcy3_2;
	wire w_dff_B_GiLNzKdD2_2;
	wire w_dff_B_KADIC0AV0_2;
	wire w_dff_B_VJ0LrDsJ5_2;
	wire w_dff_B_pbBzgsqh9_2;
	wire w_dff_B_ilkwgL9p6_2;
	wire w_dff_B_zpPXU2Yq2_2;
	wire w_dff_B_9Hw1d2E67_2;
	wire w_dff_B_ci6Xkj838_2;
	wire w_dff_B_T6ThZ1VN7_2;
	wire w_dff_B_efEoOrsF5_2;
	wire w_dff_B_1xQnkExC8_2;
	wire w_dff_B_4UzZik378_2;
	wire w_dff_B_LKVDHP0r2_2;
	wire w_dff_B_VtqfVqPy5_2;
	wire w_dff_B_ytQFanFC4_2;
	wire w_dff_B_oHZMPEqB3_2;
	wire w_dff_B_xayU2yD50_2;
	wire w_dff_B_DAT7my1X3_2;
	wire w_dff_B_YdHV0KgQ8_2;
	wire w_dff_B_1RE9BRv90_1;
	wire w_dff_B_1xrU55Ru8_2;
	wire w_dff_B_YaV28dQQ3_2;
	wire w_dff_B_Yjrc6gJ42_2;
	wire w_dff_B_Ukr3cB5x0_2;
	wire w_dff_B_ERwYQfkc0_2;
	wire w_dff_B_oQal8ZrF4_2;
	wire w_dff_B_usZwKi3J4_2;
	wire w_dff_B_bCqitPJ50_2;
	wire w_dff_B_2ZyK4bWL7_2;
	wire w_dff_B_7gN6gaJ66_2;
	wire w_dff_B_w8L7IhV79_2;
	wire w_dff_B_7KutKp0b0_2;
	wire w_dff_B_yT8tjpoK7_2;
	wire w_dff_B_uMs7yRyT9_2;
	wire w_dff_B_i2f7Y6Yv4_2;
	wire w_dff_B_AZdkpHa16_2;
	wire w_dff_B_QmRVezwg1_2;
	wire w_dff_B_kjwPxhGc7_2;
	wire w_dff_B_m4TgB3lK0_2;
	wire w_dff_B_gYPxl9zq4_2;
	wire w_dff_B_VWWjJVTc9_2;
	wire w_dff_B_vtYozoDN3_2;
	wire w_dff_B_Jjsyq7Hc5_2;
	wire w_dff_B_nNxqHRh25_1;
	wire w_dff_B_6FVp7wfK9_2;
	wire w_dff_B_uSVM9zp24_2;
	wire w_dff_B_ZbwXR7sd0_2;
	wire w_dff_B_GR5cHUbp3_2;
	wire w_dff_B_xBPaiVfs0_2;
	wire w_dff_B_wf3B6y9T1_2;
	wire w_dff_B_7yUhBR1v1_2;
	wire w_dff_B_u7qckrIH4_2;
	wire w_dff_B_GZEZDqxD6_2;
	wire w_dff_B_uTWclKZB0_2;
	wire w_dff_B_kuWK8RGY5_2;
	wire w_dff_B_y3VFfP5Q0_2;
	wire w_dff_B_gqIGHKLq7_2;
	wire w_dff_B_BJbuCKz14_2;
	wire w_dff_B_hEekkcA76_2;
	wire w_dff_B_3Yq3fpC63_2;
	wire w_dff_B_EQFCMH9U8_2;
	wire w_dff_B_Bpc4qT336_2;
	wire w_dff_B_YprPyH070_2;
	wire w_dff_B_g1o7SUW86_2;
	wire w_dff_B_Wnsct9yN9_1;
	wire w_dff_B_WLEthIES4_2;
	wire w_dff_B_JPVB1Lln7_2;
	wire w_dff_B_zoNuClxX2_2;
	wire w_dff_B_MCAlPrUI6_2;
	wire w_dff_B_MveQxUIh7_2;
	wire w_dff_B_0yqxMRmq8_2;
	wire w_dff_B_1uR6By4x2_2;
	wire w_dff_B_G9FjQpuX6_2;
	wire w_dff_B_pTXcbLj86_2;
	wire w_dff_B_13aWHWaf9_2;
	wire w_dff_B_5omikSVf3_2;
	wire w_dff_B_4TOZWLV17_2;
	wire w_dff_B_nZPCvxHK3_2;
	wire w_dff_B_rMH96HVO0_2;
	wire w_dff_B_Z3Zdxp6i2_2;
	wire w_dff_B_N8WbGEM79_2;
	wire w_dff_B_6D1veawk7_2;
	wire w_dff_B_ySOKwf7v3_1;
	wire w_dff_B_Bu5kDFb36_2;
	wire w_dff_B_1gvMluSc3_2;
	wire w_dff_B_pBCjjGPm9_2;
	wire w_dff_B_Dk3u8Pgi5_2;
	wire w_dff_B_IshrJwqg4_2;
	wire w_dff_B_PMtM9BMi8_2;
	wire w_dff_B_yRbYU5eQ1_2;
	wire w_dff_B_kpwSXUlE6_2;
	wire w_dff_B_O39suy319_2;
	wire w_dff_B_WArw8JPJ4_2;
	wire w_dff_B_uyBdwhtL5_2;
	wire w_dff_B_11zFcYfw0_2;
	wire w_dff_B_OiP437gK3_2;
	wire w_dff_B_XBXvx0H27_2;
	wire w_dff_B_iRswQ0ey1_1;
	wire w_dff_B_jcTjOypa2_2;
	wire w_dff_B_9JznZKBa8_2;
	wire w_dff_B_6dmY5Vls7_2;
	wire w_dff_B_4tL5MAtu1_2;
	wire w_dff_B_BF3tYk9g0_2;
	wire w_dff_B_bZvf2xlb5_2;
	wire w_dff_B_pZgW24Ge1_2;
	wire w_dff_B_NG9iA7hD7_2;
	wire w_dff_B_GD7v6uAu6_2;
	wire w_dff_B_oKHH0kyI4_2;
	wire w_dff_B_1ynuhIjH3_2;
	wire w_dff_B_15bCaxtq3_1;
	wire w_dff_B_PwWkD2i26_2;
	wire w_dff_B_QuL2VtNh3_2;
	wire w_dff_B_64nu832F7_2;
	wire w_dff_B_JFjJ9UwW9_2;
	wire w_dff_B_cktnGQw64_2;
	wire w_dff_B_3hfS6LpD7_2;
	wire w_dff_B_mfADympr8_2;
	wire w_dff_B_my4An37E2_2;
	wire w_dff_B_CnGC1LJ43_1;
	wire w_dff_B_WDlZjkOk6_0;
	wire w_dff_B_SzUfRClK4_2;
	wire w_dff_B_OIrHpVDL6_2;
	wire w_dff_B_BOnTrUgh6_2;
	wire w_dff_B_kzWq9imN9_2;
	wire w_dff_B_pFdws3C57_1;
	wire w_dff_A_WuclRIoY1_0;
	wire w_dff_A_dBh5L1BT2_0;
	wire w_dff_A_nybzF4DU4_1;
	wire w_dff_B_2M717mWW2_1;
	wire w_dff_B_LSlQbbUc4_2;
	wire w_dff_B_L7JheQjM9_2;
	wire w_dff_B_OooR60JJ8_2;
	wire w_dff_B_eh7Up9Fu0_2;
	wire w_dff_B_NV1Z95S91_2;
	wire w_dff_B_CHB7EotM9_2;
	wire w_dff_B_IxPt0z7L4_2;
	wire w_dff_B_knxtopdp1_2;
	wire w_dff_B_5hYVt8dC3_2;
	wire w_dff_B_CNUex1ct3_2;
	wire w_dff_B_LCopGGo09_2;
	wire w_dff_B_A6UB1nQT5_2;
	wire w_dff_B_7D7BeYab0_2;
	wire w_dff_B_AmGCKWCi0_2;
	wire w_dff_B_0w51Zm1m6_2;
	wire w_dff_B_U7wlVsm69_2;
	wire w_dff_B_M7oa6wst3_2;
	wire w_dff_B_LtiZDGRA0_2;
	wire w_dff_B_uMYL27yz2_2;
	wire w_dff_B_Us7xfdiy0_2;
	wire w_dff_B_CyVHJF063_2;
	wire w_dff_B_Prtpxoy29_2;
	wire w_dff_B_hesYcBQ25_2;
	wire w_dff_B_MSFfHjxj9_2;
	wire w_dff_B_ovwrTjgN8_2;
	wire w_dff_B_NIEcuV0g4_2;
	wire w_dff_B_6Q6vAWed1_2;
	wire w_dff_B_NVTlvgY32_2;
	wire w_dff_B_KoJIRmpW9_2;
	wire w_dff_B_Szg31fkN9_2;
	wire w_dff_B_mioyXxj12_2;
	wire w_dff_B_kf9bFCNS9_2;
	wire w_dff_B_eqosYD2w2_2;
	wire w_dff_B_Dmf6m8BR0_2;
	wire w_dff_B_N9Qi9z0Q9_2;
	wire w_dff_B_HpP7aRbU9_2;
	wire w_dff_B_b8e2FE217_2;
	wire w_dff_B_YexX2FXP8_2;
	wire w_dff_B_v1u9n2wh9_2;
	wire w_dff_B_IqiPKs9H6_2;
	wire w_dff_B_vkPk90SI4_2;
	wire w_dff_B_dRHV32lw6_2;
	wire w_dff_B_w4YMeVRn7_2;
	wire w_dff_B_gJ4jzwkt7_2;
	wire w_dff_B_0xiW4LK49_2;
	wire w_dff_B_Ee5XMWLf9_0;
	wire w_dff_A_w51f6fKg9_1;
	wire w_dff_B_xnCG75dL2_1;
	wire w_dff_B_53MaQN4X4_2;
	wire w_dff_B_KGanxDDu1_2;
	wire w_dff_B_Bs6gDwtV9_2;
	wire w_dff_B_ISeXTPpf9_2;
	wire w_dff_B_lWNKAr9w4_2;
	wire w_dff_B_GmAjXuqL2_2;
	wire w_dff_B_Mnrrvqfb6_2;
	wire w_dff_B_JUEOp0jP2_2;
	wire w_dff_B_d1KfKdJO8_2;
	wire w_dff_B_43ejrfAY0_2;
	wire w_dff_B_BjvUevhY5_2;
	wire w_dff_B_cnJSCd992_2;
	wire w_dff_B_jUgNDZPm7_2;
	wire w_dff_B_xcCmmGRM3_2;
	wire w_dff_B_Hmhlsa1h3_2;
	wire w_dff_B_QIkXkwcQ2_2;
	wire w_dff_B_jI0iw5Yv2_2;
	wire w_dff_B_93vMeepE7_2;
	wire w_dff_B_NskGbCXo3_2;
	wire w_dff_B_Q01G0jzX9_2;
	wire w_dff_B_zHH4s5XG7_2;
	wire w_dff_B_qKiqwGLP5_2;
	wire w_dff_B_NfEjddmh5_2;
	wire w_dff_B_9th4BbCO1_2;
	wire w_dff_B_DWX6gro16_2;
	wire w_dff_B_jvwO0Dk37_2;
	wire w_dff_B_yyvrSAqx6_2;
	wire w_dff_B_kJII4sUl3_2;
	wire w_dff_B_DCXxTNcP3_2;
	wire w_dff_B_FhfigvyI6_2;
	wire w_dff_B_gxHPoZ764_2;
	wire w_dff_B_uiGsonpX5_2;
	wire w_dff_B_jmigQF8R8_2;
	wire w_dff_B_1BkoRZqD4_2;
	wire w_dff_B_xJJ4MQxu6_2;
	wire w_dff_B_Af9XluMH3_2;
	wire w_dff_B_d0u4lOUS5_2;
	wire w_dff_B_eSchcl8v1_2;
	wire w_dff_B_Qs3PfOV91_2;
	wire w_dff_B_2ErB38d85_2;
	wire w_dff_B_mr1nHZhz7_2;
	wire w_dff_B_pNGp6yFR8_1;
	wire w_dff_B_T1ijMHX20_2;
	wire w_dff_B_wFZKOjKB2_2;
	wire w_dff_B_BbMdPf1Y1_2;
	wire w_dff_B_FpTDjBFC9_2;
	wire w_dff_B_BLBZhFu03_2;
	wire w_dff_B_4gbJmk3O4_2;
	wire w_dff_B_soxMN8Ja5_2;
	wire w_dff_B_oIvImuyX3_2;
	wire w_dff_B_Shfkdzxj6_2;
	wire w_dff_B_Fv119xlz5_2;
	wire w_dff_B_LIRzKSoi3_2;
	wire w_dff_B_ckSUSvKi3_2;
	wire w_dff_B_QX8ZCOEV9_2;
	wire w_dff_B_biCmIdwW5_2;
	wire w_dff_B_In7ss3oz2_2;
	wire w_dff_B_m9R1ue6B1_2;
	wire w_dff_B_jD5TeEdK8_2;
	wire w_dff_B_1tAT5HYP9_2;
	wire w_dff_B_w0lhWW4L0_2;
	wire w_dff_B_KaG9cDgs9_2;
	wire w_dff_B_t41gk4817_2;
	wire w_dff_B_RRKOLcpu0_2;
	wire w_dff_B_VPu0juO67_2;
	wire w_dff_B_sNgMEBVH1_2;
	wire w_dff_B_31fMGXW38_2;
	wire w_dff_B_ijDPh3q34_2;
	wire w_dff_B_5BWcjAtN8_2;
	wire w_dff_B_9gQurTIf8_2;
	wire w_dff_B_vHMpXA5p1_2;
	wire w_dff_B_C4hSN5h07_2;
	wire w_dff_B_i6Kh2RHd0_2;
	wire w_dff_B_6ZXrghi65_2;
	wire w_dff_B_a94EnyxS3_2;
	wire w_dff_B_1sUde2R02_2;
	wire w_dff_B_EMJpRulh7_2;
	wire w_dff_B_UPNvuDtc2_2;
	wire w_dff_B_e94QfI5g5_2;
	wire w_dff_B_5LD0MFNh0_2;
	wire w_dff_B_ECAasbK75_1;
	wire w_dff_B_Ke20WAPe4_2;
	wire w_dff_B_1XjXP9l55_2;
	wire w_dff_B_MMPIrmgd5_2;
	wire w_dff_B_uAyCDodE7_2;
	wire w_dff_B_c6lRLEDj9_2;
	wire w_dff_B_o0bpbOf17_2;
	wire w_dff_B_igfgnHTu4_2;
	wire w_dff_B_kNvsuaeZ6_2;
	wire w_dff_B_xy4bWwsH0_2;
	wire w_dff_B_EbQJL6L00_2;
	wire w_dff_B_cXD23sEV0_2;
	wire w_dff_B_lDxFzLCk0_2;
	wire w_dff_B_whBou9vE4_2;
	wire w_dff_B_QksqPF8d0_2;
	wire w_dff_B_u9vO1Nvb6_2;
	wire w_dff_B_J6XSEByu4_2;
	wire w_dff_B_oDqUxfck0_2;
	wire w_dff_B_tJIPaCUI7_2;
	wire w_dff_B_j86xvJXf7_2;
	wire w_dff_B_4N91gOOs5_2;
	wire w_dff_B_wVyFThKK2_2;
	wire w_dff_B_B1s2MeMh6_2;
	wire w_dff_B_rb2LQZfP5_2;
	wire w_dff_B_RqShlrS31_2;
	wire w_dff_B_1GESWonR3_2;
	wire w_dff_B_2Ar4nirw1_2;
	wire w_dff_B_6yqp78Sn4_2;
	wire w_dff_B_q1ZkHdQL5_2;
	wire w_dff_B_A9k3sJDT7_2;
	wire w_dff_B_0fyOtX0z4_2;
	wire w_dff_B_EkfVU8YA2_2;
	wire w_dff_B_ropKusnn7_2;
	wire w_dff_B_nEgpEXPa6_2;
	wire w_dff_B_KSl44vcR5_2;
	wire w_dff_B_n7NZzqfv9_2;
	wire w_dff_B_uw7NCiMR7_1;
	wire w_dff_B_KvSqF5Xf6_2;
	wire w_dff_B_zt9nszF87_2;
	wire w_dff_B_vrcl4GP45_2;
	wire w_dff_B_9IiAZcp32_2;
	wire w_dff_B_QYnN5lha2_2;
	wire w_dff_B_KrHSFf0N1_2;
	wire w_dff_B_o4bt0WnC5_2;
	wire w_dff_B_nJnovh7Y1_2;
	wire w_dff_B_iFBffaZp4_2;
	wire w_dff_B_FMGVtxxm0_2;
	wire w_dff_B_ZDhITpnG4_2;
	wire w_dff_B_fG6TlCOR6_2;
	wire w_dff_B_1DB1riyM5_2;
	wire w_dff_B_HBVtvih01_2;
	wire w_dff_B_SBkTADVc5_2;
	wire w_dff_B_gsO7nT6D4_2;
	wire w_dff_B_AKbNUzs42_2;
	wire w_dff_B_JPix2ID42_2;
	wire w_dff_B_NF7cbl9P3_2;
	wire w_dff_B_tIBo4Md27_2;
	wire w_dff_B_k7wjO0wN6_2;
	wire w_dff_B_ovyvEWee1_2;
	wire w_dff_B_X9jQoiQo6_2;
	wire w_dff_B_7BOU26IH7_2;
	wire w_dff_B_6yiJD5CE7_2;
	wire w_dff_B_Dyf31tXD6_2;
	wire w_dff_B_cGnUEqZN1_2;
	wire w_dff_B_TULUFHFB5_2;
	wire w_dff_B_mAr4DQtM5_2;
	wire w_dff_B_IzK4a4Es8_2;
	wire w_dff_B_hS6AMZ2m3_2;
	wire w_dff_B_y0ItLKzh4_2;
	wire w_dff_B_Dwps49C11_1;
	wire w_dff_B_LnBYv4ut4_2;
	wire w_dff_B_MRdZLkga7_2;
	wire w_dff_B_Qv2GJThw2_2;
	wire w_dff_B_AUs6zmqn3_2;
	wire w_dff_B_BgdQMJFT1_2;
	wire w_dff_B_4ATcdP1I6_2;
	wire w_dff_B_EPcGaCRJ9_2;
	wire w_dff_B_b9YLYGBa5_2;
	wire w_dff_B_VXtbv3575_2;
	wire w_dff_B_5riRUXIX6_2;
	wire w_dff_B_GYAY10FO0_2;
	wire w_dff_B_quLp7gEl4_2;
	wire w_dff_B_ygIfWRUg1_2;
	wire w_dff_B_M1W2GrJw3_2;
	wire w_dff_B_cXqLT28b1_2;
	wire w_dff_B_ZaJZXSuO1_2;
	wire w_dff_B_1cObaf4I7_2;
	wire w_dff_B_P6bPwYBd5_2;
	wire w_dff_B_k67Jsa5P8_2;
	wire w_dff_B_u9uXpZsG0_2;
	wire w_dff_B_WbeRbB8t3_2;
	wire w_dff_B_RDibWo8g7_2;
	wire w_dff_B_Ttu6j5n41_2;
	wire w_dff_B_mBkjRJXv2_2;
	wire w_dff_B_I9S76K1N0_2;
	wire w_dff_B_DtafXJMb0_2;
	wire w_dff_B_u96r5TEf0_2;
	wire w_dff_B_s1oEiOdU9_2;
	wire w_dff_B_sJWUG6142_2;
	wire w_dff_B_ZjSS2dJ77_1;
	wire w_dff_B_OovdVmMD9_2;
	wire w_dff_B_mbrfkRjZ6_2;
	wire w_dff_B_ph9WnQB71_2;
	wire w_dff_B_2hCHuFoX9_2;
	wire w_dff_B_jyrAqK5y4_2;
	wire w_dff_B_kFs4xjBA9_2;
	wire w_dff_B_P6mMWZoB0_2;
	wire w_dff_B_cIFSHJkA6_2;
	wire w_dff_B_5h9pYmoR2_2;
	wire w_dff_B_LWGaaqau1_2;
	wire w_dff_B_sTiLKptz2_2;
	wire w_dff_B_4QxDY0h17_2;
	wire w_dff_B_fs4NH9nC7_2;
	wire w_dff_B_gLHlhhrj7_2;
	wire w_dff_B_CzNupRbp4_2;
	wire w_dff_B_MdoKOw5Z7_2;
	wire w_dff_B_uM6XrG4b9_2;
	wire w_dff_B_1aPqaaPW2_2;
	wire w_dff_B_j7IJ6u3j3_2;
	wire w_dff_B_oaqFlQSI1_2;
	wire w_dff_B_oFe5B9XV2_2;
	wire w_dff_B_BwPWjQ027_2;
	wire w_dff_B_XFwmC7VM9_2;
	wire w_dff_B_5z3krZC54_2;
	wire w_dff_B_1yZeRs0z3_2;
	wire w_dff_B_wQdkmXAX3_2;
	wire w_dff_B_PxDcOGDe3_1;
	wire w_dff_B_JZ8SG1Fu1_2;
	wire w_dff_B_p8YDnsjB4_2;
	wire w_dff_B_zd57863Y5_2;
	wire w_dff_B_Ir1YAI7m4_2;
	wire w_dff_B_03C02Cah2_2;
	wire w_dff_B_yvtZqhmy4_2;
	wire w_dff_B_p8HTkv9f6_2;
	wire w_dff_B_dt2I0D6d6_2;
	wire w_dff_B_umRCVLAJ1_2;
	wire w_dff_B_7qArkClW9_2;
	wire w_dff_B_myxRQu1h0_2;
	wire w_dff_B_aurLMFSO6_2;
	wire w_dff_B_w5XKOL2x8_2;
	wire w_dff_B_t0ytvEDT6_2;
	wire w_dff_B_IiC9sOro1_2;
	wire w_dff_B_Z95Fs6UR2_2;
	wire w_dff_B_M4r6nRbe2_2;
	wire w_dff_B_vCcrBO4m3_2;
	wire w_dff_B_MoG9zz6F2_2;
	wire w_dff_B_bJtg3bdA2_2;
	wire w_dff_B_YnVZirDT9_2;
	wire w_dff_B_X1JJlNGf9_2;
	wire w_dff_B_TuOrFy6A8_2;
	wire w_dff_B_8DXc4VHP2_1;
	wire w_dff_B_oIsN6uep7_2;
	wire w_dff_B_Ih5CN3Tj0_2;
	wire w_dff_B_4kcX0mzb1_2;
	wire w_dff_B_ZvltgaRF3_2;
	wire w_dff_B_koZp7SGU2_2;
	wire w_dff_B_7kP5wfc11_2;
	wire w_dff_B_wR9LdgtU5_2;
	wire w_dff_B_1GTjPDU11_2;
	wire w_dff_B_AeK5lfvI7_2;
	wire w_dff_B_q0iyvY4j2_2;
	wire w_dff_B_zRi0fW0q7_2;
	wire w_dff_B_J2u2ttDO0_2;
	wire w_dff_B_bEtRwI3i2_2;
	wire w_dff_B_5LR6fvlK2_2;
	wire w_dff_B_pAFZ88CO8_2;
	wire w_dff_B_3rWeH4hL8_2;
	wire w_dff_B_J2hirTEo0_2;
	wire w_dff_B_vJKj6JTm9_2;
	wire w_dff_B_P90XYJTQ4_2;
	wire w_dff_B_dPQiGyWm2_2;
	wire w_dff_B_UeXsh9uZ9_1;
	wire w_dff_B_F82px3E89_2;
	wire w_dff_B_Br0cfbnG1_2;
	wire w_dff_B_pZrQ5QnB7_2;
	wire w_dff_B_q9BiA5k03_2;
	wire w_dff_B_LiQDsVnC5_2;
	wire w_dff_B_G0BU64Od8_2;
	wire w_dff_B_6rtVPpiT1_2;
	wire w_dff_B_2lvusSrS3_2;
	wire w_dff_B_gfQtg04x3_2;
	wire w_dff_B_wq79QjT70_2;
	wire w_dff_B_KViurxnT3_2;
	wire w_dff_B_lRr41Z7I0_2;
	wire w_dff_B_Q93eLLWX4_2;
	wire w_dff_B_IVnHvEPA5_2;
	wire w_dff_B_9IdZrWbO3_2;
	wire w_dff_B_bCkENo171_2;
	wire w_dff_B_joj2jMnZ3_2;
	wire w_dff_B_S3LDvzAM3_1;
	wire w_dff_B_GKexaLQJ6_2;
	wire w_dff_B_Z677QtdV3_2;
	wire w_dff_B_uVB1NLlq7_2;
	wire w_dff_B_Xk1LeGoS3_2;
	wire w_dff_B_wPG9Mjms5_2;
	wire w_dff_B_uIo3Bg5t1_2;
	wire w_dff_B_unD14ByA0_2;
	wire w_dff_B_P4FCEVZp9_2;
	wire w_dff_B_bPnAOKI30_2;
	wire w_dff_B_l01mquOU9_2;
	wire w_dff_B_7tYK5xUI4_2;
	wire w_dff_B_PA96h7SR8_2;
	wire w_dff_B_d7k18fMk7_2;
	wire w_dff_B_OSIDnEiA1_2;
	wire w_dff_B_OnsABkWv7_1;
	wire w_dff_B_1vjrn6XB0_2;
	wire w_dff_B_RVQJDNk02_2;
	wire w_dff_B_U01tVpCE9_2;
	wire w_dff_B_AZjQPbyp1_2;
	wire w_dff_B_pQJyU4jZ5_2;
	wire w_dff_B_alz9Qaub2_2;
	wire w_dff_B_qcvaPbNc8_2;
	wire w_dff_B_de23805L4_2;
	wire w_dff_B_G6F0HEmv0_2;
	wire w_dff_B_gwbk1L7D7_2;
	wire w_dff_B_in7sRfZw5_2;
	wire w_dff_B_OkUzAfi64_1;
	wire w_dff_B_uO7Gtbni9_2;
	wire w_dff_B_2YxeOzGf2_2;
	wire w_dff_B_iQHxFL9o1_2;
	wire w_dff_B_ObLDN0uT1_2;
	wire w_dff_B_GvXDFjLQ8_2;
	wire w_dff_B_cFWyPtRn7_2;
	wire w_dff_B_60eohaZi9_2;
	wire w_dff_B_2ccDlXr84_2;
	wire w_dff_B_f4uAbTBS5_1;
	wire w_dff_B_KeyIPZfW7_0;
	wire w_dff_B_ipChMsk04_2;
	wire w_dff_B_AIGDCwhD8_2;
	wire w_dff_B_zmvDwT8o8_2;
	wire w_dff_B_eL30RuV68_2;
	wire w_dff_B_x3G1lenS0_1;
	wire w_dff_A_ab6agvHO7_0;
	wire w_dff_A_SLtjRVKq4_0;
	wire w_dff_A_a8R000an1_0;
	wire w_dff_A_gZCz23As0_1;
	wire w_dff_B_Cngn24uH1_2;
	wire w_dff_B_3bupPnHd6_1;
	wire w_dff_B_aZ3jnh142_2;
	wire w_dff_B_vtqBcY7A7_2;
	wire w_dff_B_bmTkb4Q08_2;
	wire w_dff_B_8HMpiAWT9_2;
	wire w_dff_B_oxlVLBY17_2;
	wire w_dff_B_oJ57Udyv6_2;
	wire w_dff_B_tB2jw37h8_2;
	wire w_dff_B_dXUyMAfa5_2;
	wire w_dff_B_7U5BNE2h3_2;
	wire w_dff_B_vT7X76Rv3_2;
	wire w_dff_B_zny6G3B55_2;
	wire w_dff_B_mR0cDyN53_2;
	wire w_dff_B_2TyaRKCI0_2;
	wire w_dff_B_NJOjni0j8_2;
	wire w_dff_B_DRfNpyRh3_2;
	wire w_dff_B_GmYBuXMx6_2;
	wire w_dff_B_ob7u66dA5_2;
	wire w_dff_B_g1bXdf332_2;
	wire w_dff_B_xcT8Hw5A6_2;
	wire w_dff_B_JNoD57bK9_2;
	wire w_dff_B_P4IWm8Lw4_2;
	wire w_dff_B_t7xLGml19_2;
	wire w_dff_B_u2nNLLRN7_2;
	wire w_dff_B_h90Ymaf81_2;
	wire w_dff_B_RmhpkNBi2_2;
	wire w_dff_B_Cb2JB3eH4_2;
	wire w_dff_B_DlERetDA5_2;
	wire w_dff_B_AtO0RiFG2_2;
	wire w_dff_B_cPKFPiaE4_2;
	wire w_dff_B_5bqZ0WpY3_2;
	wire w_dff_B_p8vXaVt50_2;
	wire w_dff_B_kX8bOGQ94_2;
	wire w_dff_B_8lO6u5X73_2;
	wire w_dff_B_NvdEGkyk9_2;
	wire w_dff_B_xto9W2mR5_2;
	wire w_dff_B_vRuAq3F79_2;
	wire w_dff_B_OQkdBmkH5_2;
	wire w_dff_B_gBTA61rt3_2;
	wire w_dff_B_GYWVTZGF9_2;
	wire w_dff_B_fPrVdaRI2_2;
	wire w_dff_B_d3KbCPHj1_2;
	wire w_dff_B_0LAtOIli8_2;
	wire w_dff_B_Fn2HwZ4t2_2;
	wire w_dff_B_wfVjBIIC1_2;
	wire w_dff_B_1eQL6QIs8_2;
	wire w_dff_B_j079FCM32_1;
	wire w_dff_B_PI422c360_2;
	wire w_dff_B_0k1qYqts8_2;
	wire w_dff_B_n4X64WQn4_2;
	wire w_dff_B_fkPcQl4o1_2;
	wire w_dff_B_PpdQCT3Z0_2;
	wire w_dff_B_8hCRoQ5t5_2;
	wire w_dff_B_APuEXC5e9_2;
	wire w_dff_B_GbCPCTYz1_2;
	wire w_dff_B_K7jJE0Jy3_2;
	wire w_dff_B_3TK67x301_2;
	wire w_dff_B_v5NBp9iH1_2;
	wire w_dff_B_Y7fFNuvr6_2;
	wire w_dff_B_Eu5KtEvZ1_2;
	wire w_dff_B_aueFfBGV6_2;
	wire w_dff_B_tQZZZIRE0_2;
	wire w_dff_B_HQV4qQML0_2;
	wire w_dff_B_0fbb3tXx2_2;
	wire w_dff_B_1FHJatrq9_2;
	wire w_dff_B_vi3PR3DX7_2;
	wire w_dff_B_XuLUhRgw8_2;
	wire w_dff_B_Mvz7x8wc9_2;
	wire w_dff_B_zAgSOMbJ1_2;
	wire w_dff_B_LEZ89wzN3_2;
	wire w_dff_B_NOF0MlVd2_2;
	wire w_dff_B_gnkp2g2F3_2;
	wire w_dff_B_WhNPmtF40_2;
	wire w_dff_B_J0cWdLFq7_2;
	wire w_dff_B_cqEnRLDh7_2;
	wire w_dff_B_7MYw9aY48_2;
	wire w_dff_B_tb6suika7_2;
	wire w_dff_B_xXZRh6PY2_2;
	wire w_dff_B_TYtpAtfY6_2;
	wire w_dff_B_aN8JocuM8_2;
	wire w_dff_B_Vq5kSKGY4_2;
	wire w_dff_B_4gq6v1Mr3_2;
	wire w_dff_B_9AkKwsAe4_2;
	wire w_dff_B_POJg5BVq9_2;
	wire w_dff_B_uqq4h8726_2;
	wire w_dff_B_YfD2Hzhk8_2;
	wire w_dff_B_cOfaW6Mn8_2;
	wire w_dff_B_Ve6XuVT70_1;
	wire w_dff_B_nfOcNSbU3_2;
	wire w_dff_B_NTvImXe40_2;
	wire w_dff_B_QcKZOX7W0_2;
	wire w_dff_B_wmjLikGs7_2;
	wire w_dff_B_Pf16pe8T2_2;
	wire w_dff_B_UvhsvRMM4_2;
	wire w_dff_B_ojG4mz3I3_2;
	wire w_dff_B_SkndRomy4_2;
	wire w_dff_B_dVZpe6im1_2;
	wire w_dff_B_yT33qTN85_2;
	wire w_dff_B_uNT2z6zX7_2;
	wire w_dff_B_YL1NPOqU4_2;
	wire w_dff_B_uBnxwzTY1_2;
	wire w_dff_B_xGQWlKlm2_2;
	wire w_dff_B_z5IbGw5I9_2;
	wire w_dff_B_9YUShBSr9_2;
	wire w_dff_B_B6jRnsGT6_2;
	wire w_dff_B_X6eKo2i10_2;
	wire w_dff_B_lRAPt5F47_2;
	wire w_dff_B_4NuHBtki4_2;
	wire w_dff_B_Hstqz02F4_2;
	wire w_dff_B_7nDGbcRP0_2;
	wire w_dff_B_FxvLFpN11_2;
	wire w_dff_B_o8poyn7j6_2;
	wire w_dff_B_sm4MqfOX2_2;
	wire w_dff_B_Xl17A2n18_2;
	wire w_dff_B_9f07JttR6_2;
	wire w_dff_B_b9V4tXMK4_2;
	wire w_dff_B_HUBpYrcV2_2;
	wire w_dff_B_Ps0V7Caa8_2;
	wire w_dff_B_V2RoNlDE6_2;
	wire w_dff_B_sVCQM1Ir8_2;
	wire w_dff_B_mROPoYsL2_2;
	wire w_dff_B_h4CYYHiG5_2;
	wire w_dff_B_1PGqQiA23_2;
	wire w_dff_B_YpX0O3M52_2;
	wire w_dff_B_7O8tEm8a3_2;
	wire w_dff_B_tzPycaO79_1;
	wire w_dff_B_o2go5oBQ2_2;
	wire w_dff_B_7oH5w5b32_2;
	wire w_dff_B_7vc7kcyo9_2;
	wire w_dff_B_FX0QTQVc8_2;
	wire w_dff_B_3yEABLAK2_2;
	wire w_dff_B_EzfpCxNI3_2;
	wire w_dff_B_jeQIlDFF1_2;
	wire w_dff_B_FpXZ0RLg1_2;
	wire w_dff_B_mG9kDgzC6_2;
	wire w_dff_B_lZg8j7oV9_2;
	wire w_dff_B_gvRoVTrJ8_2;
	wire w_dff_B_Gn0TFo9s3_2;
	wire w_dff_B_LiQhnnfs6_2;
	wire w_dff_B_SLIBLd9q1_2;
	wire w_dff_B_2NbuIvYu0_2;
	wire w_dff_B_sAiHmYUk3_2;
	wire w_dff_B_3FM4j2vm9_2;
	wire w_dff_B_ItvwI4py1_2;
	wire w_dff_B_mDSpuFgx6_2;
	wire w_dff_B_FwMBvBaX3_2;
	wire w_dff_B_3yNBNeIM2_2;
	wire w_dff_B_HVNi8iDy8_2;
	wire w_dff_B_TFLqg0jh5_2;
	wire w_dff_B_0SAOxi2C2_2;
	wire w_dff_B_plDDwwII2_2;
	wire w_dff_B_ZxBJxJsb5_2;
	wire w_dff_B_5xG3zZT59_2;
	wire w_dff_B_ednsvzuj3_2;
	wire w_dff_B_bqNnc41A2_2;
	wire w_dff_B_NUxBqaob5_2;
	wire w_dff_B_WYutRZFW9_2;
	wire w_dff_B_4955CFnq5_2;
	wire w_dff_B_3jmo5Plu7_2;
	wire w_dff_B_jgMd85UI9_2;
	wire w_dff_B_5zfOOgKH1_1;
	wire w_dff_B_QIxohLxn2_2;
	wire w_dff_B_6hxwt7Fy4_2;
	wire w_dff_B_3XGwUPQP5_2;
	wire w_dff_B_G7giD9hq9_2;
	wire w_dff_B_xToTssDQ7_2;
	wire w_dff_B_e5iwbTld5_2;
	wire w_dff_B_Gph20BZe6_2;
	wire w_dff_B_hyqFPLER3_2;
	wire w_dff_B_lA07zuv24_2;
	wire w_dff_B_wxoAQ9ZA1_2;
	wire w_dff_B_ujlAmiKJ0_2;
	wire w_dff_B_sKJQqRI01_2;
	wire w_dff_B_PUwZJS0q9_2;
	wire w_dff_B_EvvaHqgi8_2;
	wire w_dff_B_XYBGXCFu3_2;
	wire w_dff_B_JNYZAVaS6_2;
	wire w_dff_B_tXoteiTe4_2;
	wire w_dff_B_9Dq2HxPU6_2;
	wire w_dff_B_jE9CHGHA6_2;
	wire w_dff_B_9eHXxFAx0_2;
	wire w_dff_B_o0Co45uI2_2;
	wire w_dff_B_84v3fYGE8_2;
	wire w_dff_B_VwQvWoxP5_2;
	wire w_dff_B_HMMxcNY57_2;
	wire w_dff_B_gE0BVxXE6_2;
	wire w_dff_B_Pf201PmX5_2;
	wire w_dff_B_CRxlwRcg9_2;
	wire w_dff_B_sSNVoSWM0_2;
	wire w_dff_B_5HPx6JnY1_2;
	wire w_dff_B_B1c5aMwc9_2;
	wire w_dff_B_vAKqYFTu3_2;
	wire w_dff_B_P0j1A7UR7_1;
	wire w_dff_B_OXIUOoLh4_2;
	wire w_dff_B_CmZbFzZh6_2;
	wire w_dff_B_z1UvYoPe3_2;
	wire w_dff_B_8zS91aOP5_2;
	wire w_dff_B_HaCrWVrX1_2;
	wire w_dff_B_uon66A4t7_2;
	wire w_dff_B_CAVtoGyb2_2;
	wire w_dff_B_d38Y6Adh0_2;
	wire w_dff_B_qRpnyxTx7_2;
	wire w_dff_B_0KhrJO591_2;
	wire w_dff_B_fYYc96mb7_2;
	wire w_dff_B_UAMoE8dV9_2;
	wire w_dff_B_fKhjjdYX9_2;
	wire w_dff_B_KrdBSDVd2_2;
	wire w_dff_B_7zN15ypl5_2;
	wire w_dff_B_QRhlHi2y5_2;
	wire w_dff_B_OZcXcJNC6_2;
	wire w_dff_B_xsb35Enf5_2;
	wire w_dff_B_iyTO8Kl67_2;
	wire w_dff_B_ManyWFd04_2;
	wire w_dff_B_o9S6mCbt4_2;
	wire w_dff_B_hMoX1NjO8_2;
	wire w_dff_B_M6S4EStO2_2;
	wire w_dff_B_hI21th195_2;
	wire w_dff_B_NjjlAV5p3_2;
	wire w_dff_B_wliBZn6i9_2;
	wire w_dff_B_Nhrj8v1l1_2;
	wire w_dff_B_dJ60ay428_2;
	wire w_dff_B_UDL5hThD3_1;
	wire w_dff_B_WYR6X4fS7_2;
	wire w_dff_B_1EiUASCF3_2;
	wire w_dff_B_wNJco7zY9_2;
	wire w_dff_B_5Cj3yCW42_2;
	wire w_dff_B_hT4hPMCR3_2;
	wire w_dff_B_vA6MhM9C2_2;
	wire w_dff_B_FIpGf8mP1_2;
	wire w_dff_B_MVsv0wPv0_2;
	wire w_dff_B_mg0O518l1_2;
	wire w_dff_B_kMt8oLOT1_2;
	wire w_dff_B_wSNUgtch3_2;
	wire w_dff_B_8y9ykXg09_2;
	wire w_dff_B_uKuqM9kx5_2;
	wire w_dff_B_XyAt3mok3_2;
	wire w_dff_B_dnhHSFST4_2;
	wire w_dff_B_5cpiIYba4_2;
	wire w_dff_B_NGJkUk2B5_2;
	wire w_dff_B_DWgZfIhi8_2;
	wire w_dff_B_qqAHShGX3_2;
	wire w_dff_B_DAyPCTnv6_2;
	wire w_dff_B_FfYx2GC76_2;
	wire w_dff_B_NpaD1rYU5_2;
	wire w_dff_B_9B3sKFAV5_2;
	wire w_dff_B_dn1IyzkQ2_2;
	wire w_dff_B_3UUv34cF6_2;
	wire w_dff_B_TCeNeTdF2_1;
	wire w_dff_B_QcUiI7CH3_2;
	wire w_dff_B_p0mKxhVA7_2;
	wire w_dff_B_Gzj7WSl15_2;
	wire w_dff_B_Sj4h1qfx0_2;
	wire w_dff_B_pkvnDbSG7_2;
	wire w_dff_B_PenXEBXB5_2;
	wire w_dff_B_GQXZorl61_2;
	wire w_dff_B_ifYq9zLr9_2;
	wire w_dff_B_6w5OLoTf3_2;
	wire w_dff_B_glB7C4ag2_2;
	wire w_dff_B_NV1kw4X71_2;
	wire w_dff_B_Yxm4oLyq7_2;
	wire w_dff_B_YqoqONaq2_2;
	wire w_dff_B_HYyigz4y9_2;
	wire w_dff_B_WMOHkmnw6_2;
	wire w_dff_B_30Lm1NbZ3_2;
	wire w_dff_B_ribJBYlS7_2;
	wire w_dff_B_z8FhWHer3_2;
	wire w_dff_B_67wGB1fs5_2;
	wire w_dff_B_oejDmRnQ4_2;
	wire w_dff_B_qWIwacVh8_2;
	wire w_dff_B_jReiZpSs1_2;
	wire w_dff_B_YElVKpLK0_1;
	wire w_dff_B_xlbZDUBi6_2;
	wire w_dff_B_kLXiJHaK5_2;
	wire w_dff_B_3MZieGVZ5_2;
	wire w_dff_B_nvGxiWNk0_2;
	wire w_dff_B_7SBpEuGF3_2;
	wire w_dff_B_WoGYCLPa6_2;
	wire w_dff_B_hfEpRZxv5_2;
	wire w_dff_B_04pQeXka8_2;
	wire w_dff_B_LTIjk67s1_2;
	wire w_dff_B_ZppctRjs8_2;
	wire w_dff_B_xCudkfpS0_2;
	wire w_dff_B_FAMxKb3Q8_2;
	wire w_dff_B_WbTqpJMO0_2;
	wire w_dff_B_gZhJ61136_2;
	wire w_dff_B_LbLHEl9s2_2;
	wire w_dff_B_WplqsmkK7_2;
	wire w_dff_B_cPkiZ6ip5_2;
	wire w_dff_B_KezsfKsU0_2;
	wire w_dff_B_UEsYEI8b8_2;
	wire w_dff_B_o79ldpKl3_1;
	wire w_dff_B_KLDDFsu83_2;
	wire w_dff_B_FpqF9WsI6_2;
	wire w_dff_B_jmIzYgfK4_2;
	wire w_dff_B_wtpiBXXw0_2;
	wire w_dff_B_u5QYdera1_2;
	wire w_dff_B_FQ9oS25q2_2;
	wire w_dff_B_PXb4sKmT7_2;
	wire w_dff_B_ctwbJgRX1_2;
	wire w_dff_B_HSQXpIsl9_2;
	wire w_dff_B_dlzBw1uu6_2;
	wire w_dff_B_8YaGXYWq7_2;
	wire w_dff_B_O5Pov7Hy9_2;
	wire w_dff_B_K0kHUNdJ1_2;
	wire w_dff_B_T5OkNbqd0_2;
	wire w_dff_B_ZlqvOwWy0_2;
	wire w_dff_B_2oiaiKTi4_2;
	wire w_dff_B_6jsqFIrz7_1;
	wire w_dff_B_u7E9BCYc3_2;
	wire w_dff_B_A3UpByrr6_2;
	wire w_dff_B_ECMFJSbV7_2;
	wire w_dff_B_97I8f5Tv9_2;
	wire w_dff_B_cbLYQat23_2;
	wire w_dff_B_VZbOWOIH8_2;
	wire w_dff_B_jCLVR2lx4_2;
	wire w_dff_B_HRevj4JV1_2;
	wire w_dff_B_B6d6QJdc7_2;
	wire w_dff_B_Q5eu5QZV0_2;
	wire w_dff_B_dNJb3Yeb1_2;
	wire w_dff_B_zIQaBel87_2;
	wire w_dff_B_ip1OYZXP2_2;
	wire w_dff_B_OxFG7zEq4_1;
	wire w_dff_B_IaqEn6cD0_2;
	wire w_dff_B_95LMWnMg1_2;
	wire w_dff_B_wScDON8r5_2;
	wire w_dff_B_gUmVQuXm4_2;
	wire w_dff_B_rqajqbQu9_2;
	wire w_dff_B_ksSQGzqn5_2;
	wire w_dff_B_r85wganR1_2;
	wire w_dff_B_TXbdvrH06_2;
	wire w_dff_B_QPOFtPMW1_2;
	wire w_dff_B_VkUFP3RP6_2;
	wire w_dff_B_io9CbdDf0_2;
	wire w_dff_B_FqnL9AwD9_1;
	wire w_dff_B_DYZfqvEo8_2;
	wire w_dff_B_HGKg3pE81_2;
	wire w_dff_B_X03eZoHQ5_2;
	wire w_dff_B_UPMDiGPW9_2;
	wire w_dff_B_cxJ5nufr4_2;
	wire w_dff_B_VSZnugCs8_2;
	wire w_dff_B_qiqaGBdF2_2;
	wire w_dff_B_GQJav8ev3_2;
	wire w_dff_B_Us5gRVrN8_1;
	wire w_dff_B_reSi97mk6_2;
	wire w_dff_B_plJwiYGs8_2;
	wire w_dff_B_kqNS9IRA6_2;
	wire w_dff_B_NxmFnLMh2_2;
	wire w_dff_B_ld0GMe2J5_1;
	wire w_dff_A_ihGef0np8_1;
	wire w_dff_A_UFdfwBAu8_2;
	wire w_dff_A_ME7jCby71_2;
	wire w_dff_B_a33fP2nu5_2;
	wire w_dff_B_ldfrfag78_1;
	wire w_dff_B_YopbOVgc0_2;
	wire w_dff_B_eWIuPVRh6_2;
	wire w_dff_B_GRDWU3Zx6_2;
	wire w_dff_B_0fyB5x247_2;
	wire w_dff_B_VLvMbGr95_2;
	wire w_dff_B_kDS3O4KO7_2;
	wire w_dff_B_06gyuQDf8_2;
	wire w_dff_B_31MFiyW06_2;
	wire w_dff_B_v2kQEH1V3_2;
	wire w_dff_B_hxE3nZQB8_2;
	wire w_dff_B_HBifSMOO0_2;
	wire w_dff_B_4C4RFaPW2_2;
	wire w_dff_B_wLYE6GuJ5_2;
	wire w_dff_B_9m9kf7zg4_2;
	wire w_dff_B_znXQe2J80_2;
	wire w_dff_B_teBCpntl9_2;
	wire w_dff_B_wicxiOmA5_2;
	wire w_dff_B_Zy60lVAV2_2;
	wire w_dff_B_lE6DP6rJ8_2;
	wire w_dff_B_aKSAEdNP7_2;
	wire w_dff_B_fSk7J3782_2;
	wire w_dff_B_pfO65SxL1_2;
	wire w_dff_B_8b1SmzKf6_2;
	wire w_dff_B_mJ85caAD8_2;
	wire w_dff_B_miI1PorH1_2;
	wire w_dff_B_HD7tQvOF1_2;
	wire w_dff_B_KbYHEZsq2_2;
	wire w_dff_B_WUSUN2y83_2;
	wire w_dff_B_zM5xh3Ux3_2;
	wire w_dff_B_gYXFpMN14_2;
	wire w_dff_B_2vbDUsx77_2;
	wire w_dff_B_yGgFNGF35_2;
	wire w_dff_B_Ae60r8WL9_2;
	wire w_dff_B_xHv7a9Jw2_2;
	wire w_dff_B_NtRzrdJq3_2;
	wire w_dff_B_8vEXte5I0_2;
	wire w_dff_B_P19jcpSz5_2;
	wire w_dff_B_6udUZmPU9_2;
	wire w_dff_B_D3CIDLky0_2;
	wire w_dff_B_xByME6L32_2;
	wire w_dff_B_VPP5cuBQ8_2;
	wire w_dff_B_gUpcipTp4_2;
	wire w_dff_B_vlb96aLX1_2;
	wire w_dff_B_FsrhkoL98_2;
	wire w_dff_B_hFQBophy3_2;
	wire w_dff_B_Vzsvtm4e3_2;
	wire w_dff_B_gMOD04LK8_1;
	wire w_dff_B_JPKKkgyZ2_2;
	wire w_dff_B_XI1hN6LU8_2;
	wire w_dff_B_OEp2csFP1_2;
	wire w_dff_B_zSLDlSjR2_2;
	wire w_dff_B_qroJzE191_2;
	wire w_dff_B_HPeq6HI29_2;
	wire w_dff_B_IHE6y6hl2_2;
	wire w_dff_B_TL7fwjhG1_2;
	wire w_dff_B_gnjlbvzi4_2;
	wire w_dff_B_wWluNzAv1_2;
	wire w_dff_B_G8Ao3u3H9_2;
	wire w_dff_B_fUqjQJOO1_2;
	wire w_dff_B_hbdkR3oi6_2;
	wire w_dff_B_iisJzLOF6_2;
	wire w_dff_B_rlV2Adwh7_2;
	wire w_dff_B_voFJmxMS9_2;
	wire w_dff_B_QBGxZDqj4_2;
	wire w_dff_B_GVEgjdkh0_2;
	wire w_dff_B_fiMewi637_2;
	wire w_dff_B_TnyTLXOj3_2;
	wire w_dff_B_tIBRf3oc1_2;
	wire w_dff_B_jeO4sf1y5_2;
	wire w_dff_B_9aiGenyJ0_2;
	wire w_dff_B_KgMIuiRv3_2;
	wire w_dff_B_maD6bYUp0_2;
	wire w_dff_B_E3hVxtbw5_2;
	wire w_dff_B_jnNrYOPt7_2;
	wire w_dff_B_mJSkHJbU7_2;
	wire w_dff_B_m3eRQ6ht4_2;
	wire w_dff_B_NkWAB6qo9_2;
	wire w_dff_B_6iqaITqX3_2;
	wire w_dff_B_Q6cPTMuz3_2;
	wire w_dff_B_Q72KRGlz9_2;
	wire w_dff_B_j9AdApCh5_2;
	wire w_dff_B_GEDCO0BG4_2;
	wire w_dff_B_MN5QEbox8_2;
	wire w_dff_B_faP0WOb70_2;
	wire w_dff_B_iNdENpZB7_2;
	wire w_dff_B_TcqLODSQ1_2;
	wire w_dff_B_uRxpRYjz2_2;
	wire w_dff_B_48lD1CKl9_2;
	wire w_dff_B_RZ68iGV39_1;
	wire w_dff_B_KFJiuq5N9_2;
	wire w_dff_B_0YKe3tCR5_2;
	wire w_dff_B_3rbb7qLk6_2;
	wire w_dff_B_sJUeJWGk0_2;
	wire w_dff_B_75jZM8Ny8_2;
	wire w_dff_B_djLFzpT95_2;
	wire w_dff_B_reFHK3Yc4_2;
	wire w_dff_B_BHvNkurK6_2;
	wire w_dff_B_kAeCw6A77_2;
	wire w_dff_B_pqociOfC7_2;
	wire w_dff_B_89rbMWGo2_2;
	wire w_dff_B_g7c2nQDA0_2;
	wire w_dff_B_rG3yH1Hq7_2;
	wire w_dff_B_liKv9Xwc3_2;
	wire w_dff_B_rY5h51Sy4_2;
	wire w_dff_B_L5JkQPZ33_2;
	wire w_dff_B_yU6BNIox6_2;
	wire w_dff_B_ko1uQX8q9_2;
	wire w_dff_B_94YFYyOb3_2;
	wire w_dff_B_cLWsJTfx5_2;
	wire w_dff_B_Nc7jlJOn1_2;
	wire w_dff_B_bpA98IQ31_2;
	wire w_dff_B_crlLbWCT1_2;
	wire w_dff_B_FbxaMjPy3_2;
	wire w_dff_B_2fl6Fxwo8_2;
	wire w_dff_B_TPbtqJO76_2;
	wire w_dff_B_V1Yo2WOt2_2;
	wire w_dff_B_6PHdLnga7_2;
	wire w_dff_B_cnaKGKw74_2;
	wire w_dff_B_236yhGDc5_2;
	wire w_dff_B_git90gTn4_2;
	wire w_dff_B_YFZr2Nw31_2;
	wire w_dff_B_npnLzxhn2_2;
	wire w_dff_B_AAQ7mzk81_2;
	wire w_dff_B_KMmU36vm5_2;
	wire w_dff_B_6zEDXQG32_2;
	wire w_dff_B_ftoLNtMu0_2;
	wire w_dff_B_WDf10k9W8_2;
	wire w_dff_B_ZI9ttziG9_1;
	wire w_dff_B_5H3rShpr7_2;
	wire w_dff_B_8VVajlqj1_2;
	wire w_dff_B_bAVnja4l2_2;
	wire w_dff_B_Uc6xRWYa9_2;
	wire w_dff_B_LRvRgw2j0_2;
	wire w_dff_B_xcJPdG8w2_2;
	wire w_dff_B_1bvD3nxm7_2;
	wire w_dff_B_ASBkdjsz7_2;
	wire w_dff_B_8I2C815e1_2;
	wire w_dff_B_z1QCF9jJ6_2;
	wire w_dff_B_nxCQ0w4O1_2;
	wire w_dff_B_JDDM5JJs7_2;
	wire w_dff_B_jGGTOKtQ5_2;
	wire w_dff_B_tsV8RmVd3_2;
	wire w_dff_B_lQjfcswZ6_2;
	wire w_dff_B_cO59nhhm8_2;
	wire w_dff_B_pyoOHU246_2;
	wire w_dff_B_mJlORRbv0_2;
	wire w_dff_B_SUStyfXp9_2;
	wire w_dff_B_bHfjIWcU9_2;
	wire w_dff_B_3NuufQ5J1_2;
	wire w_dff_B_u2X4psDd6_2;
	wire w_dff_B_2pH2f6uW9_2;
	wire w_dff_B_lwC2gSPs2_2;
	wire w_dff_B_fSBAsAr70_2;
	wire w_dff_B_3CeHHTiH2_2;
	wire w_dff_B_twBWysc17_2;
	wire w_dff_B_iZWSx8Ib7_2;
	wire w_dff_B_xu8kWeZT1_2;
	wire w_dff_B_YoSLBF7D6_2;
	wire w_dff_B_4X8NU8Ze6_2;
	wire w_dff_B_MrRiON2f2_2;
	wire w_dff_B_M13MTssq1_2;
	wire w_dff_B_iZoOIOJk2_2;
	wire w_dff_B_f2fXMfxO2_2;
	wire w_dff_B_h96iplJp8_1;
	wire w_dff_B_qf1KbyvZ9_2;
	wire w_dff_B_GiRXq2pD7_2;
	wire w_dff_B_sFXmxg8H3_2;
	wire w_dff_B_0yoVnBMw0_2;
	wire w_dff_B_RwYS4Orm3_2;
	wire w_dff_B_oIzowEBO4_2;
	wire w_dff_B_1m30Jtb47_2;
	wire w_dff_B_G3DM9bid2_2;
	wire w_dff_B_ko52E0RT1_2;
	wire w_dff_B_16dFWnR53_2;
	wire w_dff_B_wSzjwccF5_2;
	wire w_dff_B_YvuMUbEI9_2;
	wire w_dff_B_JFGP2rfe0_2;
	wire w_dff_B_17Hop5s74_2;
	wire w_dff_B_6ZYgppYs0_2;
	wire w_dff_B_w5Qj2VkR7_2;
	wire w_dff_B_p80WPCGv9_2;
	wire w_dff_B_IvxFYclK9_2;
	wire w_dff_B_83514W5S9_2;
	wire w_dff_B_gagttwTN8_2;
	wire w_dff_B_fagEDV9h5_2;
	wire w_dff_B_Wf05x0wK6_2;
	wire w_dff_B_AHPGsVDo8_2;
	wire w_dff_B_eImlIFJa4_2;
	wire w_dff_B_EQlOIpa20_2;
	wire w_dff_B_bTKE2vxA3_2;
	wire w_dff_B_dMcF30JL8_2;
	wire w_dff_B_XDxMHo5Z4_2;
	wire w_dff_B_rdtuf9CZ9_2;
	wire w_dff_B_UQtSHOaW8_2;
	wire w_dff_B_Ymx0eTka8_2;
	wire w_dff_B_K9MfCiiH9_2;
	wire w_dff_B_gKd82W6n2_1;
	wire w_dff_B_k0xdLmBg4_2;
	wire w_dff_B_VRLMVOOx8_2;
	wire w_dff_B_BRIZJtgZ4_2;
	wire w_dff_B_IkzqHC132_2;
	wire w_dff_B_tNdueXcE1_2;
	wire w_dff_B_ffOYEBMO4_2;
	wire w_dff_B_ESnLHkbH0_2;
	wire w_dff_B_FUYTKE2j4_2;
	wire w_dff_B_G8btJlP34_2;
	wire w_dff_B_k4qDj2Ga0_2;
	wire w_dff_B_BXDDCU8X4_2;
	wire w_dff_B_0rgr56EP8_2;
	wire w_dff_B_NgqsGmwE2_2;
	wire w_dff_B_lpKppnX52_2;
	wire w_dff_B_NiP8qZpS5_2;
	wire w_dff_B_uzvUZMxA4_2;
	wire w_dff_B_ZlbwXcYs5_2;
	wire w_dff_B_N01fWury7_2;
	wire w_dff_B_izJRony38_2;
	wire w_dff_B_tEBojRND8_2;
	wire w_dff_B_0hkuzV6i5_2;
	wire w_dff_B_dgR86CNW8_2;
	wire w_dff_B_zYhZMvND2_2;
	wire w_dff_B_FLVCCj0G8_2;
	wire w_dff_B_hAwQIO8k7_2;
	wire w_dff_B_cmJXqYMn6_2;
	wire w_dff_B_qeQMGMeM3_2;
	wire w_dff_B_U38vW7tC1_2;
	wire w_dff_B_hSUeKmrL0_2;
	wire w_dff_B_kCfO6Aus2_1;
	wire w_dff_B_PbN4Eizn7_2;
	wire w_dff_B_dwGTMwxF7_2;
	wire w_dff_B_cog3cDJ09_2;
	wire w_dff_B_PO7USqUY7_2;
	wire w_dff_B_4DxmM4Yi2_2;
	wire w_dff_B_fpKF7vWF4_2;
	wire w_dff_B_E6J55IHH9_2;
	wire w_dff_B_ptzncvBY9_2;
	wire w_dff_B_cyAbCoaC9_2;
	wire w_dff_B_bWapu2ob4_2;
	wire w_dff_B_7ry2q6NH6_2;
	wire w_dff_B_eP9fNeyA4_2;
	wire w_dff_B_eGQr13TS4_2;
	wire w_dff_B_OxZD4LAk5_2;
	wire w_dff_B_UBY4ksMm9_2;
	wire w_dff_B_tTd7OPdb0_2;
	wire w_dff_B_SHeUR4Sv5_2;
	wire w_dff_B_8eaMojvU9_2;
	wire w_dff_B_OUWETMbk1_2;
	wire w_dff_B_90v5L3Bz6_2;
	wire w_dff_B_xO9qI2a85_2;
	wire w_dff_B_EfJ9Vx9R3_2;
	wire w_dff_B_Rvcy1IOO3_2;
	wire w_dff_B_vIhzUtvF0_2;
	wire w_dff_B_ldwTfSl73_2;
	wire w_dff_B_bsFbhQmc0_2;
	wire w_dff_B_Nv9sc4k00_1;
	wire w_dff_B_J9T8q5a18_2;
	wire w_dff_B_ZbyGjajf2_2;
	wire w_dff_B_NUel66ar8_2;
	wire w_dff_B_TNfSqxTJ1_2;
	wire w_dff_B_OYSSLdlg7_2;
	wire w_dff_B_OeFb2pvZ6_2;
	wire w_dff_B_xiEhIQEO9_2;
	wire w_dff_B_GxzQNKvI3_2;
	wire w_dff_B_2rAVyXYa2_2;
	wire w_dff_B_9XTBTupQ8_2;
	wire w_dff_B_28YkXFdP4_2;
	wire w_dff_B_PPAgc3366_2;
	wire w_dff_B_NP0XiZvg9_2;
	wire w_dff_B_yDuHGVi34_2;
	wire w_dff_B_wj3lF2p25_2;
	wire w_dff_B_yJ5YPjel7_2;
	wire w_dff_B_rqKP1Z425_2;
	wire w_dff_B_h2d35uWt7_2;
	wire w_dff_B_5SmefWIh7_2;
	wire w_dff_B_8qpIUJ1q2_2;
	wire w_dff_B_WV1L8tsl5_2;
	wire w_dff_B_bB0kAjRn7_2;
	wire w_dff_B_jXm3dBaj8_2;
	wire w_dff_B_NfzOU8uG7_1;
	wire w_dff_B_UddFAk9F3_2;
	wire w_dff_B_aF20CRb32_2;
	wire w_dff_B_Mm38oxW87_2;
	wire w_dff_B_0AWD1DAx1_2;
	wire w_dff_B_j55uUv796_2;
	wire w_dff_B_zcBHRLik0_2;
	wire w_dff_B_a2gGLxfn6_2;
	wire w_dff_B_CODX0LgQ2_2;
	wire w_dff_B_KJRbJor27_2;
	wire w_dff_B_Zn7slPYZ7_2;
	wire w_dff_B_EGJCjpjA7_2;
	wire w_dff_B_alIpKFw52_2;
	wire w_dff_B_w5LNbcyV9_2;
	wire w_dff_B_983xOmMV2_2;
	wire w_dff_B_h8Q7jCOb0_2;
	wire w_dff_B_wGWHjVzP5_2;
	wire w_dff_B_eQ816E361_2;
	wire w_dff_B_C7wYALGK1_2;
	wire w_dff_B_aI2f7H149_2;
	wire w_dff_B_Ef4mkVVx3_2;
	wire w_dff_B_aS9WQCEK1_1;
	wire w_dff_B_XvBRwcpl7_2;
	wire w_dff_B_EHf0HZtO6_2;
	wire w_dff_B_FFe7cNla8_2;
	wire w_dff_B_5RicMekn8_2;
	wire w_dff_B_o3ALsuSM7_2;
	wire w_dff_B_Ctyu6zb89_2;
	wire w_dff_B_ccLgiHjv4_2;
	wire w_dff_B_CN69VyeF0_2;
	wire w_dff_B_jHP4GolN1_2;
	wire w_dff_B_7VzO5X2y9_2;
	wire w_dff_B_1zwhxOMR1_2;
	wire w_dff_B_dcc151WO0_2;
	wire w_dff_B_VGhdKhtI2_2;
	wire w_dff_B_YnkYjL2D3_2;
	wire w_dff_B_cs1K0E3V8_2;
	wire w_dff_B_lwA8I24v7_2;
	wire w_dff_B_fFbzYEDd7_2;
	wire w_dff_B_OlGt9Uuj4_1;
	wire w_dff_B_ukYQadji0_2;
	wire w_dff_B_W4KVTdUj5_2;
	wire w_dff_B_hxCJIC1i1_2;
	wire w_dff_B_YkFgylAc6_2;
	wire w_dff_B_azSjNYVm9_2;
	wire w_dff_B_nhe4O2Va9_2;
	wire w_dff_B_RpVEfoGQ7_2;
	wire w_dff_B_zH4DftIt4_2;
	wire w_dff_B_eCttojSS2_2;
	wire w_dff_B_dVKWTuVr6_2;
	wire w_dff_B_tAecjG1c2_2;
	wire w_dff_B_MQ9nJEQ77_2;
	wire w_dff_B_H8BgJNg37_2;
	wire w_dff_B_UOTUdhWY3_2;
	wire w_dff_B_g62wjsut6_1;
	wire w_dff_B_mofUbUYw9_2;
	wire w_dff_B_niybe1Iv7_2;
	wire w_dff_B_ZyESmRrZ5_2;
	wire w_dff_B_EPUifdh25_2;
	wire w_dff_B_rja1QFI06_2;
	wire w_dff_B_R8tjpMQq4_2;
	wire w_dff_B_vCFwQKYd9_2;
	wire w_dff_B_nzeE4d2Q3_2;
	wire w_dff_B_wzXhIDkY3_2;
	wire w_dff_B_YYVXrBV72_2;
	wire w_dff_B_wz3dzYdM9_2;
	wire w_dff_B_j6F4Nlxt6_2;
	wire w_dff_B_qL2BFsb78_1;
	wire w_dff_B_3Se7Sk4K0_2;
	wire w_dff_B_2osNilFo9_2;
	wire w_dff_B_xnS6lx2i0_2;
	wire w_dff_B_ehvJyKEo2_2;
	wire w_dff_B_AdIRERwX0_2;
	wire w_dff_B_OkaMSu4h5_2;
	wire w_dff_B_9r95EjvW0_2;
	wire w_dff_B_8bw6Fr9D8_1;
	wire w_dff_B_F4LgOeMa1_2;
	wire w_dff_B_Uly7U9a64_2;
	wire w_dff_B_Ytmx2Tpe3_2;
	wire w_dff_B_CpkB4cPl0_2;
	wire w_dff_B_COEn0i7q4_1;
	wire w_dff_A_aBDBlh6d9_0;
	wire w_dff_A_OWBOdTT50_1;
	wire w_dff_A_eBdNRukX7_1;
	wire w_dff_B_dNZdGybo7_1;
	wire w_dff_B_OaC6pXkf2_2;
	wire w_dff_B_bzQZHME51_2;
	wire w_dff_B_qjo4ML0j0_2;
	wire w_dff_B_lW6ummAk4_2;
	wire w_dff_B_HAMdJXqj4_2;
	wire w_dff_B_SP7WhHL67_2;
	wire w_dff_B_LaQCwOWy0_2;
	wire w_dff_B_14Xlus2t8_2;
	wire w_dff_B_xOSKmMFo8_2;
	wire w_dff_B_V5YreD3D5_2;
	wire w_dff_B_uvhoH1SS8_2;
	wire w_dff_B_f8BKMykT4_2;
	wire w_dff_B_zSr0kpJE8_2;
	wire w_dff_B_xZbkgrvL4_2;
	wire w_dff_B_dXkBzECY6_2;
	wire w_dff_B_yjUKA5dm2_2;
	wire w_dff_B_vZeAWra68_2;
	wire w_dff_B_eB5GVjmy3_2;
	wire w_dff_B_ZwGW23gW1_2;
	wire w_dff_B_0gVfbluu6_2;
	wire w_dff_B_eFVkGurk6_2;
	wire w_dff_B_XJM0d1OB9_2;
	wire w_dff_B_ouWZbJ9b9_2;
	wire w_dff_B_19cuWiUj1_2;
	wire w_dff_B_IvR2Vxpf3_2;
	wire w_dff_B_sAfgoOGC1_2;
	wire w_dff_B_oI9oCBLJ8_2;
	wire w_dff_B_GAGxHBL25_2;
	wire w_dff_B_57mQVH8X6_2;
	wire w_dff_B_Ahei8Xw10_2;
	wire w_dff_B_zNAtCrG97_2;
	wire w_dff_B_zG7eIA2k6_2;
	wire w_dff_B_WLeD4J7R0_2;
	wire w_dff_B_x1VE0BXf2_2;
	wire w_dff_B_3UDgbXl85_2;
	wire w_dff_B_w7r14DpS8_2;
	wire w_dff_B_TLOdqBCR5_2;
	wire w_dff_B_oqcAXjZY4_2;
	wire w_dff_B_WCVgGZJd3_2;
	wire w_dff_B_gxzjjlWO1_2;
	wire w_dff_B_JQKp7SRZ4_2;
	wire w_dff_B_dqZnbUCp3_2;
	wire w_dff_B_p47rBmF72_2;
	wire w_dff_B_rFbxQWOV3_2;
	wire w_dff_B_syuyrcj01_2;
	wire w_dff_B_p6FGVhTh7_2;
	wire w_dff_B_f5hCBJZx7_2;
	wire w_dff_B_rSxV2MYi3_0;
	wire w_dff_A_fK9qtCNH5_1;
	wire w_dff_B_pVRMKH112_1;
	wire w_dff_B_2s4yTaNW8_2;
	wire w_dff_B_339u2ylJ9_2;
	wire w_dff_B_pqbFETGt8_2;
	wire w_dff_B_NG2Kevfy5_2;
	wire w_dff_B_nlJtgKHu2_2;
	wire w_dff_B_LE3cqdHL7_2;
	wire w_dff_B_WfpD5SbF6_2;
	wire w_dff_B_LKhtnuhk3_2;
	wire w_dff_B_j0c0Kj3Y1_2;
	wire w_dff_B_njHtBhzj3_2;
	wire w_dff_B_kAtIHfPU9_2;
	wire w_dff_B_LHFPeuCu5_2;
	wire w_dff_B_5UO3cQxI7_2;
	wire w_dff_B_MspLqAmI8_2;
	wire w_dff_B_16qeeGLi6_2;
	wire w_dff_B_77yuZhVP2_2;
	wire w_dff_B_p5eHDbOQ4_2;
	wire w_dff_B_iPzakK8z5_2;
	wire w_dff_B_PcNY3Rs13_2;
	wire w_dff_B_a0ifAPls6_2;
	wire w_dff_B_IzEMmRMk8_2;
	wire w_dff_B_uDY1FGLF6_2;
	wire w_dff_B_YWYEcBk66_2;
	wire w_dff_B_Jzjomdso8_2;
	wire w_dff_B_BOFqJPvP0_2;
	wire w_dff_B_tBXtUiTt4_2;
	wire w_dff_B_U3lGBHK96_2;
	wire w_dff_B_oqA7mvpU6_2;
	wire w_dff_B_Wge6w4UP6_2;
	wire w_dff_B_TZBI3ML91_2;
	wire w_dff_B_e3m7vQf03_2;
	wire w_dff_B_l9h8n5uz4_2;
	wire w_dff_B_2smcDJBn8_2;
	wire w_dff_B_l5yMxhnj3_2;
	wire w_dff_B_S1eIQdOD7_2;
	wire w_dff_B_FWzn2Zgp8_2;
	wire w_dff_B_Gr5JGbmA5_2;
	wire w_dff_B_cMdYXuJ37_2;
	wire w_dff_B_HguAhdNx3_2;
	wire w_dff_B_6Sa4aOd89_2;
	wire w_dff_B_nEVlyori2_2;
	wire w_dff_B_Z9LoOTDA7_2;
	wire w_dff_B_8w6Vab4P0_2;
	wire w_dff_B_9e3ArnSM4_1;
	wire w_dff_B_XfwUtztd4_2;
	wire w_dff_B_ZYpPyd7D8_2;
	wire w_dff_B_o8JqlCPX7_2;
	wire w_dff_B_5PIcEdNX7_2;
	wire w_dff_B_omAJYMEv7_2;
	wire w_dff_B_Wasq2FvN5_2;
	wire w_dff_B_WscfOdyS2_2;
	wire w_dff_B_5KsJoTbB1_2;
	wire w_dff_B_Gu6FDvBM0_2;
	wire w_dff_B_AMrgHlco9_2;
	wire w_dff_B_jTrfBuMJ3_2;
	wire w_dff_B_s60lqEXF6_2;
	wire w_dff_B_tqwzxJFg1_2;
	wire w_dff_B_fBToE5Ig5_2;
	wire w_dff_B_KlosOtsY3_2;
	wire w_dff_B_EtYeH5jM2_2;
	wire w_dff_B_RDhSc2Hj0_2;
	wire w_dff_B_9CaG2y445_2;
	wire w_dff_B_zD1M4WBq9_2;
	wire w_dff_B_VCoDaFvr7_2;
	wire w_dff_B_qpvjGOiZ6_2;
	wire w_dff_B_p176txV42_2;
	wire w_dff_B_yH86lC9q1_2;
	wire w_dff_B_VxUcgy9p7_2;
	wire w_dff_B_e1u9NH2T7_2;
	wire w_dff_B_8ZXWSOco2_2;
	wire w_dff_B_Yslkd1rH1_2;
	wire w_dff_B_viwLNiED5_2;
	wire w_dff_B_oRVTyjUm3_2;
	wire w_dff_B_sOmRu7fn8_2;
	wire w_dff_B_ImAHvpZZ1_2;
	wire w_dff_B_dLpTrMyX5_2;
	wire w_dff_B_JtrT2PDz5_2;
	wire w_dff_B_2lOJk4B49_2;
	wire w_dff_B_nc1ovFbM5_2;
	wire w_dff_B_b28KNNQc0_2;
	wire w_dff_B_JBxP3dqb3_2;
	wire w_dff_B_e12GkItb2_2;
	wire w_dff_B_mTGVb2Y87_2;
	wire w_dff_B_wRhOut4q0_2;
	wire w_dff_B_HdN6e2QS5_1;
	wire w_dff_B_cfbh6X9D7_2;
	wire w_dff_B_pOT4qoYE9_2;
	wire w_dff_B_rjq7m8fe5_2;
	wire w_dff_B_MTuFUmnU5_2;
	wire w_dff_B_wvJP5jEF0_2;
	wire w_dff_B_Nk7tMNV87_2;
	wire w_dff_B_F9uI3vXr8_2;
	wire w_dff_B_9ESwFd571_2;
	wire w_dff_B_CTQr98h62_2;
	wire w_dff_B_O6Cj7JoH4_2;
	wire w_dff_B_ynsDrXfz9_2;
	wire w_dff_B_Uf3367ra5_2;
	wire w_dff_B_0af13xxu5_2;
	wire w_dff_B_Kw7vO2ZE4_2;
	wire w_dff_B_A50lyDmP1_2;
	wire w_dff_B_B12yDqG91_2;
	wire w_dff_B_5uO59pTn4_2;
	wire w_dff_B_gtldhGR49_2;
	wire w_dff_B_btLbHQG55_2;
	wire w_dff_B_jdCCI9yg0_2;
	wire w_dff_B_b3oEeMNT3_2;
	wire w_dff_B_rpLcmaKz7_2;
	wire w_dff_B_GIpjYGQf5_2;
	wire w_dff_B_4XeTKFQn7_2;
	wire w_dff_B_v6ceRsv35_2;
	wire w_dff_B_i8lKL3H85_2;
	wire w_dff_B_6EyYZzVG6_2;
	wire w_dff_B_zKpleKsM8_2;
	wire w_dff_B_X3hfhygc5_2;
	wire w_dff_B_9yGH2G2T3_2;
	wire w_dff_B_rqUVYrVU9_2;
	wire w_dff_B_HFkZRdSW2_2;
	wire w_dff_B_hv2AnX7z3_2;
	wire w_dff_B_djjgwTXb7_2;
	wire w_dff_B_Wx6OaocS6_2;
	wire w_dff_B_LczfR24N0_2;
	wire w_dff_B_iqP04Ira2_2;
	wire w_dff_B_z5RhBe3P9_1;
	wire w_dff_B_ahExX52R0_2;
	wire w_dff_B_v1RNsA6J9_2;
	wire w_dff_B_cJL8jU797_2;
	wire w_dff_B_eA16Gydg5_2;
	wire w_dff_B_HzZ6NIKZ0_2;
	wire w_dff_B_lIS2M8i35_2;
	wire w_dff_B_BlvSV2fL8_2;
	wire w_dff_B_IYhS2iSa6_2;
	wire w_dff_B_amg2TSHd5_2;
	wire w_dff_B_CBRTIi9H5_2;
	wire w_dff_B_9RfQCK361_2;
	wire w_dff_B_Y3ycp56H7_2;
	wire w_dff_B_UqpjfU9K1_2;
	wire w_dff_B_WerwZNX65_2;
	wire w_dff_B_XIXe867m6_2;
	wire w_dff_B_UiRo5sdd1_2;
	wire w_dff_B_NwydGrbz1_2;
	wire w_dff_B_YLDc6gkU2_2;
	wire w_dff_B_2N1Yr9ex1_2;
	wire w_dff_B_QXlBy0AW5_2;
	wire w_dff_B_P4ZlhUqU8_2;
	wire w_dff_B_leDsltOd6_2;
	wire w_dff_B_4oJiMfPy2_2;
	wire w_dff_B_SVfCfHwD8_2;
	wire w_dff_B_q3wKuDe99_2;
	wire w_dff_B_650xjR7n2_2;
	wire w_dff_B_Slrvo9Ty9_2;
	wire w_dff_B_89vM4sNl6_2;
	wire w_dff_B_pfgS2cDN7_2;
	wire w_dff_B_7mbIxNWX3_2;
	wire w_dff_B_xJj2QTNd3_2;
	wire w_dff_B_V0XZExdl1_2;
	wire w_dff_B_Za3PwOC99_2;
	wire w_dff_B_AvICfoV98_2;
	wire w_dff_B_gkznpBEf4_1;
	wire w_dff_B_Um5dOghd3_2;
	wire w_dff_B_H9E6PndJ4_2;
	wire w_dff_B_mLYq6oUH3_2;
	wire w_dff_B_qOMWTWBP5_2;
	wire w_dff_B_1whUBTFv3_2;
	wire w_dff_B_Mwfq03dg8_2;
	wire w_dff_B_srBU42iG0_2;
	wire w_dff_B_AKkFTaAY9_2;
	wire w_dff_B_hEVWqqtR3_2;
	wire w_dff_B_JmZnRLM25_2;
	wire w_dff_B_7jVS0mXv5_2;
	wire w_dff_B_UHmDUxO57_2;
	wire w_dff_B_CjtcbXPy7_2;
	wire w_dff_B_7lY1tv9g5_2;
	wire w_dff_B_WwvHEjaQ0_2;
	wire w_dff_B_snmFQfGG1_2;
	wire w_dff_B_qyeUTYx37_2;
	wire w_dff_B_uW37g5LN3_2;
	wire w_dff_B_equ5fY3g1_2;
	wire w_dff_B_cdQk5QfP5_2;
	wire w_dff_B_AviJSpvS3_2;
	wire w_dff_B_owY0euqi6_2;
	wire w_dff_B_yvbmzEOI3_2;
	wire w_dff_B_7E72KJj92_2;
	wire w_dff_B_vXbupGDE7_2;
	wire w_dff_B_LiKea8F97_2;
	wire w_dff_B_X3kIljoC4_2;
	wire w_dff_B_vRZtnJ3b7_2;
	wire w_dff_B_dlF8wpcl4_2;
	wire w_dff_B_QMuW436K2_2;
	wire w_dff_B_tK1POAiv8_2;
	wire w_dff_B_AWEkbpKd1_1;
	wire w_dff_B_5vBfRpeh4_2;
	wire w_dff_B_M2ILRsz14_2;
	wire w_dff_B_QjrNtuYS3_2;
	wire w_dff_B_kb4jkFpI7_2;
	wire w_dff_B_1RBGOdJH1_2;
	wire w_dff_B_enG3Nk1C4_2;
	wire w_dff_B_9gFfoXFU0_2;
	wire w_dff_B_ZFHIbfop4_2;
	wire w_dff_B_8SNUpDdJ0_2;
	wire w_dff_B_8EDZHkR78_2;
	wire w_dff_B_H52xUj512_2;
	wire w_dff_B_Hcx913mr2_2;
	wire w_dff_B_GJBaQ3Y26_2;
	wire w_dff_B_AXk6Rmex0_2;
	wire w_dff_B_tBAQOmxm2_2;
	wire w_dff_B_JwLdyZUt0_2;
	wire w_dff_B_2Uys5daT8_2;
	wire w_dff_B_VvDPI0nO7_2;
	wire w_dff_B_QAnNtVyB4_2;
	wire w_dff_B_fImbjnfv7_2;
	wire w_dff_B_193FPRAe6_2;
	wire w_dff_B_0XLaWxPT5_2;
	wire w_dff_B_gNZp66ua7_2;
	wire w_dff_B_uURC9QOx5_2;
	wire w_dff_B_Hywtq1Vt1_2;
	wire w_dff_B_VUUqCtZM2_2;
	wire w_dff_B_MjkJMhHw9_2;
	wire w_dff_B_BLi57DKT7_2;
	wire w_dff_B_qwmlGLoC7_1;
	wire w_dff_B_euHYX45B4_2;
	wire w_dff_B_A1z9AQnR1_2;
	wire w_dff_B_UejawuOu4_2;
	wire w_dff_B_qrnNWu0h4_2;
	wire w_dff_B_UN6E8hBU2_2;
	wire w_dff_B_GZc0UFjg3_2;
	wire w_dff_B_Sziofqbt8_2;
	wire w_dff_B_wP0DZBgY8_2;
	wire w_dff_B_yLXbKVKd0_2;
	wire w_dff_B_b3WXyUQe3_2;
	wire w_dff_B_sK9bpa6M6_2;
	wire w_dff_B_eQWzRKi33_2;
	wire w_dff_B_P6aWvTaA8_2;
	wire w_dff_B_qZmgXeD04_2;
	wire w_dff_B_rPhT8Vtk6_2;
	wire w_dff_B_LNrPLZp47_2;
	wire w_dff_B_tgrg1QM66_2;
	wire w_dff_B_PokZ6lb99_2;
	wire w_dff_B_1EwewgJP1_2;
	wire w_dff_B_rrtrXJzX3_2;
	wire w_dff_B_pzAnSdtX1_2;
	wire w_dff_B_UABLJ9ch4_2;
	wire w_dff_B_hWnCGiGP0_2;
	wire w_dff_B_Iell99iK5_2;
	wire w_dff_B_fIPyYPm37_2;
	wire w_dff_B_5qkz8cg51_1;
	wire w_dff_B_BoEwLXE98_2;
	wire w_dff_B_s3DLjG1M5_2;
	wire w_dff_B_72R1pmrG2_2;
	wire w_dff_B_N8CUq8oI7_2;
	wire w_dff_B_ZrPzR4LO1_2;
	wire w_dff_B_zOVgel6M8_2;
	wire w_dff_B_ooH9eEDJ8_2;
	wire w_dff_B_prHYvDcF8_2;
	wire w_dff_B_LoJzzz282_2;
	wire w_dff_B_KG9YTMnp0_2;
	wire w_dff_B_NPG4eW0u9_2;
	wire w_dff_B_sr5SH9mf4_2;
	wire w_dff_B_PYtNlISA0_2;
	wire w_dff_B_2noJLMqk7_2;
	wire w_dff_B_9NFdoTIe5_2;
	wire w_dff_B_Y3j9pDfy8_2;
	wire w_dff_B_kPVOvwrw1_2;
	wire w_dff_B_D2eo2n0s1_2;
	wire w_dff_B_jpcMik465_2;
	wire w_dff_B_Paijxd6A3_2;
	wire w_dff_B_Z8L1CnUT9_2;
	wire w_dff_B_WSBkRGqV8_2;
	wire w_dff_B_at4LAabB1_1;
	wire w_dff_B_xm9sL97L3_2;
	wire w_dff_B_IJM3OSEj6_2;
	wire w_dff_B_UaIeGqz83_2;
	wire w_dff_B_2PDd1dUx3_2;
	wire w_dff_B_diK9KQf09_2;
	wire w_dff_B_CgqCN6Ob6_2;
	wire w_dff_B_yrbs7l8d4_2;
	wire w_dff_B_apjji1UT0_2;
	wire w_dff_B_ek5MbE8t4_2;
	wire w_dff_B_A8GwERoR6_2;
	wire w_dff_B_llqUQRuw1_2;
	wire w_dff_B_RoFBmCux9_2;
	wire w_dff_B_B8SSFgt11_2;
	wire w_dff_B_h79TveDr7_2;
	wire w_dff_B_XsGsk21n0_2;
	wire w_dff_B_Hi2RD2N60_2;
	wire w_dff_B_wFOIOPRv5_2;
	wire w_dff_B_hsU6ID7L5_2;
	wire w_dff_B_wuzspgXl2_2;
	wire w_dff_B_7p28RDIn2_1;
	wire w_dff_B_IvhAtpny5_2;
	wire w_dff_B_ntUjpUV23_2;
	wire w_dff_B_aXQJ4Nol2_2;
	wire w_dff_B_F6eAuYKZ0_2;
	wire w_dff_B_Udhy0t6J0_2;
	wire w_dff_B_lmWiHY131_2;
	wire w_dff_B_OvqtrIH24_2;
	wire w_dff_B_Ai7eka4U2_2;
	wire w_dff_B_iLaE0e8Z1_2;
	wire w_dff_B_Inh5uVQS7_2;
	wire w_dff_B_EMq02nqV4_2;
	wire w_dff_B_KFImtiDl6_2;
	wire w_dff_B_tSfP3CgY5_2;
	wire w_dff_B_UlTiNIbn1_2;
	wire w_dff_B_KZqUSP9O5_2;
	wire w_dff_B_Y2egNx893_2;
	wire w_dff_B_31QFqtey6_1;
	wire w_dff_B_vP52Pb2a6_2;
	wire w_dff_B_1t8bvtjs3_2;
	wire w_dff_B_NrlT1bAy1_2;
	wire w_dff_B_Z9SNXE2q4_2;
	wire w_dff_B_WKUyCBj38_2;
	wire w_dff_B_LB8L9Yvo7_2;
	wire w_dff_B_p2RIrWX56_2;
	wire w_dff_B_pNC0CmEc3_2;
	wire w_dff_B_RyrqkUYe9_2;
	wire w_dff_B_zCXSiF3q7_2;
	wire w_dff_B_kAILsstx7_2;
	wire w_dff_B_c848xsSQ9_2;
	wire w_dff_B_upS3G5Yz1_2;
	wire w_dff_B_d1adPsZB7_1;
	wire w_dff_B_fw470LLj2_2;
	wire w_dff_B_6EfH1EH60_2;
	wire w_dff_B_9WPp3wtB4_2;
	wire w_dff_B_g4yDPvSI4_2;
	wire w_dff_B_6ZYf0Wku2_2;
	wire w_dff_B_nTiI5cAn6_2;
	wire w_dff_B_RKafCkak1_2;
	wire w_dff_B_qYiD3Cj93_2;
	wire w_dff_B_mJYNJxgE9_2;
	wire w_dff_B_hguGGLuJ8_2;
	wire w_dff_B_pOhTzdCH3_2;
	wire w_dff_B_oo7D6KYu1_1;
	wire w_dff_B_sjyUoo7r6_1;
	wire w_dff_B_miAtFRV98_1;
	wire w_dff_B_8EBzYBeb4_1;
	wire w_dff_B_NQ3EdVAi2_1;
	wire w_dff_B_Un0ukGf28_1;
	wire w_dff_B_WX9qKg549_0;
	wire w_dff_B_4BpUftWB8_0;
	wire w_dff_A_l59cnuZg1_0;
	wire w_dff_A_kSDZ4KsA5_0;
	wire w_dff_A_FNgLIZwm6_0;
	wire w_dff_B_qmu8Bjy34_1;
	wire w_dff_A_BCYGFEtJ4_0;
	wire w_dff_A_XTS216BY7_1;
	wire w_dff_A_TShp7RaZ3_1;
	wire w_dff_A_xGyqHUB36_1;
	wire w_dff_A_gzqnjVnz3_1;
	wire w_dff_A_vBbfU2UW7_1;
	wire w_dff_A_Fin152cb7_1;
	wire w_dff_A_AIO1wok05_1;
	wire w_dff_A_Fn4KLys41_1;
	wire w_dff_B_SRfgufy24_2;
	wire w_dff_B_eA7aoaMJ9_2;
	wire w_dff_B_sOht3dtF1_1;
	wire w_dff_B_7UQ2vDpt1_2;
	wire w_dff_B_huhSvj3r8_2;
	wire w_dff_B_871pwHoW0_2;
	wire w_dff_B_S5GWN62B7_2;
	wire w_dff_B_r78LakDc8_2;
	wire w_dff_B_tBkInLPj6_2;
	wire w_dff_B_XONPbD7x5_2;
	wire w_dff_B_xk9jNLee5_2;
	wire w_dff_B_h78Cr5E01_2;
	wire w_dff_B_qwMZolfl7_2;
	wire w_dff_B_jB0rlgym9_2;
	wire w_dff_B_PDPXy9p86_2;
	wire w_dff_B_IMQ55Fku5_2;
	wire w_dff_B_FqKH4nCt2_2;
	wire w_dff_B_LSj3fhoK4_2;
	wire w_dff_B_oLxYCPow6_2;
	wire w_dff_B_LRzd3Ust8_2;
	wire w_dff_B_38XKmR9x9_2;
	wire w_dff_B_7aqk4jRV4_2;
	wire w_dff_B_zkkDv3E37_2;
	wire w_dff_B_MdZXwrO87_2;
	wire w_dff_B_RWiWCDx43_2;
	wire w_dff_B_pfZ4jjN22_2;
	wire w_dff_B_5yxv7tkq0_2;
	wire w_dff_B_iI5Wie4t2_2;
	wire w_dff_B_W5IwKxo92_2;
	wire w_dff_B_xhY1LQaj5_2;
	wire w_dff_B_lCgs9Int7_2;
	wire w_dff_B_jUamT2Mz3_2;
	wire w_dff_B_UQbfboNu6_2;
	wire w_dff_B_hPou34aI7_2;
	wire w_dff_B_hwJ0obT02_2;
	wire w_dff_B_2AQTaIZL4_2;
	wire w_dff_B_0kuy7kFZ9_2;
	wire w_dff_B_Z6HkTEQZ8_2;
	wire w_dff_B_8aMgngwz9_2;
	wire w_dff_B_rvc7jwsb6_2;
	wire w_dff_B_oGK8bSH33_2;
	wire w_dff_B_InQRtAr46_2;
	wire w_dff_B_QnJnjJhi7_2;
	wire w_dff_B_QuMjzmJb6_2;
	wire w_dff_B_HpTYzOoU6_2;
	wire w_dff_B_tnFkS6LD3_2;
	wire w_dff_B_7nSIKhlr0_2;
	wire w_dff_B_H5P1Ru7E9_2;
	wire w_dff_B_x57F2QSf8_2;
	wire w_dff_B_NFOVWNVB8_2;
	wire w_dff_B_rwbfXufI7_1;
	wire w_dff_B_Mvf2yZgD3_2;
	wire w_dff_B_pQvDS6CJ8_2;
	wire w_dff_B_9isAehT03_2;
	wire w_dff_B_NPzyMXyw8_2;
	wire w_dff_B_JDaUb3UT0_2;
	wire w_dff_B_4HkQPYwG4_2;
	wire w_dff_B_wUAZFx8i3_2;
	wire w_dff_B_kqgyDSbB7_2;
	wire w_dff_B_WBU4xJDb6_2;
	wire w_dff_B_Txeyitlz0_2;
	wire w_dff_B_3gEGxFem4_2;
	wire w_dff_B_GagQk1B23_2;
	wire w_dff_B_K9MDhRgH9_2;
	wire w_dff_B_bVpb0vZx3_2;
	wire w_dff_B_ysoCoTuV6_2;
	wire w_dff_B_CjHb5NVu2_2;
	wire w_dff_B_zbeL8hEc1_2;
	wire w_dff_B_FqnPh0Ac3_2;
	wire w_dff_B_mEzzAhU84_2;
	wire w_dff_B_DHNhYu8h6_2;
	wire w_dff_B_jIlodVVD3_2;
	wire w_dff_B_NQEFVnjF8_2;
	wire w_dff_B_vXDTy26G7_2;
	wire w_dff_B_f3ccBAjS1_2;
	wire w_dff_B_DWNrcmau4_2;
	wire w_dff_B_GNGYj2926_2;
	wire w_dff_B_MhkjpI8u8_2;
	wire w_dff_B_m3iwztcT4_2;
	wire w_dff_B_yzcaKUmW1_2;
	wire w_dff_B_4o77uoY66_2;
	wire w_dff_B_JskkLIcq3_2;
	wire w_dff_B_ObfWJ0v77_2;
	wire w_dff_B_Z5x83MkA7_2;
	wire w_dff_B_0o0WE9rC9_2;
	wire w_dff_B_0eA6watc4_2;
	wire w_dff_B_dHiVH9Qm0_2;
	wire w_dff_B_18vL9vgB9_2;
	wire w_dff_B_oBmBB0qd8_2;
	wire w_dff_B_smj5HRXp3_2;
	wire w_dff_B_iAHRBxRd4_2;
	wire w_dff_B_9VX2uy3g5_2;
	wire w_dff_B_TV43XzgL1_2;
	wire w_dff_B_BwMT4r4s5_2;
	wire w_dff_B_XiSKkmLA7_1;
	wire w_dff_B_UFZsLjkw2_2;
	wire w_dff_B_OxU07TAa7_2;
	wire w_dff_B_b3kbwmDA4_2;
	wire w_dff_B_uzCmvRUr1_2;
	wire w_dff_B_Q3yPZTjQ0_2;
	wire w_dff_B_JtNrimHy7_2;
	wire w_dff_B_vHKvY9xx8_2;
	wire w_dff_B_LYmqUexy1_2;
	wire w_dff_B_nzXB5Axe0_2;
	wire w_dff_B_o0KuoGH45_2;
	wire w_dff_B_HrqJFEGP7_2;
	wire w_dff_B_vwEbBfa66_2;
	wire w_dff_B_j4FjnTbs3_2;
	wire w_dff_B_XTStYCP62_2;
	wire w_dff_B_lXXVWJKZ8_2;
	wire w_dff_B_d9bnuhPI1_2;
	wire w_dff_B_O00mVJWo6_2;
	wire w_dff_B_OmdAFn3f6_2;
	wire w_dff_B_QrG3MQFZ8_2;
	wire w_dff_B_PBiylGLt6_2;
	wire w_dff_B_UKFjPI116_2;
	wire w_dff_B_WuS5Uz2n7_2;
	wire w_dff_B_niOnAxFJ5_2;
	wire w_dff_B_v9QocWb95_2;
	wire w_dff_B_buf3OLjB7_2;
	wire w_dff_B_yRftY1Vk2_2;
	wire w_dff_B_onEH6jfg7_2;
	wire w_dff_B_tcI9A7fe1_2;
	wire w_dff_B_9mt8ZGc07_2;
	wire w_dff_B_Tslrz7OR0_2;
	wire w_dff_B_1OcW82H66_2;
	wire w_dff_B_1lC2vAhN2_2;
	wire w_dff_B_8Ds5zo293_2;
	wire w_dff_B_6eiamWys7_2;
	wire w_dff_B_C4rtvTfn2_2;
	wire w_dff_B_SjAAH8dP5_2;
	wire w_dff_B_cXN8GZMR2_2;
	wire w_dff_B_RFzc39rY8_2;
	wire w_dff_B_dZq68j420_2;
	wire w_dff_B_HDcp3aG34_2;
	wire w_dff_B_1JFEX1qQ4_1;
	wire w_dff_B_HZGu3cma2_2;
	wire w_dff_B_XNIyxbBy3_2;
	wire w_dff_B_I98fVVhP9_2;
	wire w_dff_B_ZSGFVfg87_2;
	wire w_dff_B_Q11PkA5z9_2;
	wire w_dff_B_oIDAby5q5_2;
	wire w_dff_B_qgDDOgEK5_2;
	wire w_dff_B_CmEJZYRf7_2;
	wire w_dff_B_AZQy3XSX2_2;
	wire w_dff_B_YHB9kQED6_2;
	wire w_dff_B_s7wvoDhq8_2;
	wire w_dff_B_vY3Anbyk1_2;
	wire w_dff_B_odDdmaQV4_2;
	wire w_dff_B_Wzpp64Y94_2;
	wire w_dff_B_L8OC3DjU9_2;
	wire w_dff_B_jIfNha519_2;
	wire w_dff_B_92Bf2roA2_2;
	wire w_dff_B_Sblvx5pt6_2;
	wire w_dff_B_dR5qpD550_2;
	wire w_dff_B_T8zy2mK06_2;
	wire w_dff_B_4wktHXKN7_2;
	wire w_dff_B_PXdDBign1_2;
	wire w_dff_B_ltelvjfZ1_2;
	wire w_dff_B_rdjL7JGq1_2;
	wire w_dff_B_bx2Zq2VQ7_2;
	wire w_dff_B_rSmeVuHS9_2;
	wire w_dff_B_FDqiVCnI7_2;
	wire w_dff_B_pq9IWWZu5_2;
	wire w_dff_B_33Z4DPbN0_2;
	wire w_dff_B_OjK0KNgq1_2;
	wire w_dff_B_L3eFov7W4_2;
	wire w_dff_B_b87Rd3sz6_2;
	wire w_dff_B_cSb3M2FH2_2;
	wire w_dff_B_ixZfKWQW1_2;
	wire w_dff_B_h44IoPU77_2;
	wire w_dff_B_4jwkYf7z2_2;
	wire w_dff_B_Fjw6Mauc8_2;
	wire w_dff_B_ckoJgik34_1;
	wire w_dff_B_BUzwAzmW1_2;
	wire w_dff_B_nhGAj5Hc6_2;
	wire w_dff_B_goePkZZT3_2;
	wire w_dff_B_LQsgcfT99_2;
	wire w_dff_B_xkuW47bO8_2;
	wire w_dff_B_ZXGmVv0z9_2;
	wire w_dff_B_L6EvGvoJ5_2;
	wire w_dff_B_TS6mNVD46_2;
	wire w_dff_B_jfFICcWr8_2;
	wire w_dff_B_R1sKQJhC0_2;
	wire w_dff_B_Ze2Ww4tU6_2;
	wire w_dff_B_BTBcaIhU8_2;
	wire w_dff_B_pt1L801d0_2;
	wire w_dff_B_OwH5Bnl94_2;
	wire w_dff_B_kUUqCF2v9_2;
	wire w_dff_B_1ezRevFb5_2;
	wire w_dff_B_7EaYkE927_2;
	wire w_dff_B_FkC94jJG1_2;
	wire w_dff_B_MRv00Cms0_2;
	wire w_dff_B_bRLP17tr7_2;
	wire w_dff_B_GVDXnYiT3_2;
	wire w_dff_B_tmmyJO6H8_2;
	wire w_dff_B_KCuZ7vS78_2;
	wire w_dff_B_8jOKard33_2;
	wire w_dff_B_I1ZoLuMB0_2;
	wire w_dff_B_CjplzZ6j5_2;
	wire w_dff_B_W94DCY7N9_2;
	wire w_dff_B_8IRTFaGX9_2;
	wire w_dff_B_T9Hi2CWP2_2;
	wire w_dff_B_vGJjGu0s8_2;
	wire w_dff_B_TRXvdSrD5_2;
	wire w_dff_B_rB5tgRum1_2;
	wire w_dff_B_eC9RpPVU6_2;
	wire w_dff_B_2UwdX7bc2_2;
	wire w_dff_B_q3cqk8wI7_1;
	wire w_dff_B_auwTIVFR1_2;
	wire w_dff_B_0DsliCtt0_2;
	wire w_dff_B_bkOpRP0e6_2;
	wire w_dff_B_LaTCcrM55_2;
	wire w_dff_B_8T85ZtNL2_2;
	wire w_dff_B_oJSSqais1_2;
	wire w_dff_B_nJvTM4YU0_2;
	wire w_dff_B_tYsAHgzx2_2;
	wire w_dff_B_DSTjxvUO3_2;
	wire w_dff_B_FGLdiDzD1_2;
	wire w_dff_B_5syXlhcn3_2;
	wire w_dff_B_PoHsGxcf9_2;
	wire w_dff_B_pdl2veQ49_2;
	wire w_dff_B_EgZqF5cf8_2;
	wire w_dff_B_PLN4BaHI4_2;
	wire w_dff_B_TcNQNQQ27_2;
	wire w_dff_B_ndL5Mfm68_2;
	wire w_dff_B_JDGjRaL27_2;
	wire w_dff_B_FUppF7bS9_2;
	wire w_dff_B_3IPEXlJ09_2;
	wire w_dff_B_URgeEkML7_2;
	wire w_dff_B_3AKeL1FL9_2;
	wire w_dff_B_SFaYoCVH2_2;
	wire w_dff_B_S4C5hUq79_2;
	wire w_dff_B_JqsryJaH7_2;
	wire w_dff_B_tlftLW2g3_2;
	wire w_dff_B_3tMK8PX95_2;
	wire w_dff_B_c44AnU8s7_2;
	wire w_dff_B_JVPyZeaB5_2;
	wire w_dff_B_xlGvVhf30_2;
	wire w_dff_B_dW6wxl6L3_2;
	wire w_dff_B_XgFFSGbv9_1;
	wire w_dff_B_2o09OKuV8_2;
	wire w_dff_B_zgYJ0pHr6_2;
	wire w_dff_B_nLOEvRYt2_2;
	wire w_dff_B_NCjfJO1t4_2;
	wire w_dff_B_4PD5ByvA2_2;
	wire w_dff_B_n8SZAGFl6_2;
	wire w_dff_B_rllWA5NL2_2;
	wire w_dff_B_1TlrS8Wi4_2;
	wire w_dff_B_4mXHrKEz8_2;
	wire w_dff_B_RiGlJB8F7_2;
	wire w_dff_B_7ErlvpRI7_2;
	wire w_dff_B_VGQaozw35_2;
	wire w_dff_B_iDcCYbTy9_2;
	wire w_dff_B_hFnnzyKg9_2;
	wire w_dff_B_36aCdQqs1_2;
	wire w_dff_B_zJWHwpmw2_2;
	wire w_dff_B_xu99mW7m6_2;
	wire w_dff_B_L9WJ1Hq10_2;
	wire w_dff_B_OzzuWtfr4_2;
	wire w_dff_B_eSSNZ9hf2_2;
	wire w_dff_B_0cSgwv064_2;
	wire w_dff_B_Yk2TGZCQ6_2;
	wire w_dff_B_MeEXKSJ12_2;
	wire w_dff_B_w7HHdtyQ2_2;
	wire w_dff_B_RWcd2X5d0_2;
	wire w_dff_B_Me1QunXb1_2;
	wire w_dff_B_YDUtoW4R7_2;
	wire w_dff_B_EisvOOA97_2;
	wire w_dff_B_UXKY7mn06_1;
	wire w_dff_B_8sgDm9NF2_2;
	wire w_dff_B_TBDdfDyR2_2;
	wire w_dff_B_r6JjjiU71_2;
	wire w_dff_B_XGovgof19_2;
	wire w_dff_B_Fo1XGixH7_2;
	wire w_dff_B_C9pKSjZ53_2;
	wire w_dff_B_BZ0JSpxN5_2;
	wire w_dff_B_JOaHNq4c1_2;
	wire w_dff_B_HfweC5BM9_2;
	wire w_dff_B_girXWb537_2;
	wire w_dff_B_wVH4Xcqz8_2;
	wire w_dff_B_3ZZ3Zrdy8_2;
	wire w_dff_B_MZzN1EZd7_2;
	wire w_dff_B_qwGsE8z64_2;
	wire w_dff_B_5DkLULiV4_2;
	wire w_dff_B_hNzpbAAV5_2;
	wire w_dff_B_hXs4bfJi6_2;
	wire w_dff_B_F1VjSATd5_2;
	wire w_dff_B_TwQghdDz1_2;
	wire w_dff_B_EtLqrdVo4_2;
	wire w_dff_B_xKke7LSc0_2;
	wire w_dff_B_IAYLx7mw7_2;
	wire w_dff_B_6dGQuVQ40_2;
	wire w_dff_B_g97xEijh0_2;
	wire w_dff_B_FNpHUw6v3_2;
	wire w_dff_B_hxo8JQPg8_1;
	wire w_dff_B_mYCkYm2d2_2;
	wire w_dff_B_VYQj7Cxz5_2;
	wire w_dff_B_fB3zviGM0_2;
	wire w_dff_B_5iPVPvLl8_2;
	wire w_dff_B_MveOTinn4_2;
	wire w_dff_B_Jz4oOYo95_2;
	wire w_dff_B_wHK2ikOq9_2;
	wire w_dff_B_I8Epqzad1_2;
	wire w_dff_B_qQDpREwL1_2;
	wire w_dff_B_FnVBqF0B2_2;
	wire w_dff_B_6G4OdG8v9_2;
	wire w_dff_B_RpOu18NR3_2;
	wire w_dff_B_AnvPfdSS4_2;
	wire w_dff_B_heKggPzN9_2;
	wire w_dff_B_YnvwImeh3_2;
	wire w_dff_B_hdgmBAZ34_2;
	wire w_dff_B_diaAH8yP6_2;
	wire w_dff_B_3LujCoJV6_2;
	wire w_dff_B_a4iW99d93_2;
	wire w_dff_B_CjApRlu04_2;
	wire w_dff_B_22rxImAM4_2;
	wire w_dff_B_znWFqW642_2;
	wire w_dff_B_7ThjlGih2_1;
	wire w_dff_B_XaOk3fSX7_2;
	wire w_dff_B_JO6KkWhK4_2;
	wire w_dff_B_lfY27dJP3_2;
	wire w_dff_B_jneRnVpk7_2;
	wire w_dff_B_yB8FO8Wb0_2;
	wire w_dff_B_fr8RiATb0_2;
	wire w_dff_B_droAkZxZ3_2;
	wire w_dff_B_CGHNnbgz0_2;
	wire w_dff_B_XRuruMet1_2;
	wire w_dff_B_UrkMKO8C4_2;
	wire w_dff_B_uZXURiRo4_2;
	wire w_dff_B_vK2tTix46_2;
	wire w_dff_B_JELBREoE1_2;
	wire w_dff_B_hi6wsLRV7_2;
	wire w_dff_B_EUHJQGSs1_2;
	wire w_dff_B_QlcaS6xt6_2;
	wire w_dff_B_CpTTwEOK3_2;
	wire w_dff_B_ikKPjnGQ6_2;
	wire w_dff_B_szXqKr1U5_2;
	wire w_dff_B_EHm0L3KP9_1;
	wire w_dff_B_HyrPJHJQ3_2;
	wire w_dff_B_GDAsc6sk7_2;
	wire w_dff_B_NDxrJoVg9_2;
	wire w_dff_B_SEvZthWw3_2;
	wire w_dff_B_EdB1Pe199_2;
	wire w_dff_B_GguUIXlm3_2;
	wire w_dff_B_U4KAo54S1_2;
	wire w_dff_B_K1waBADP9_2;
	wire w_dff_B_SWPEdXiK2_2;
	wire w_dff_B_9byeOhXv5_2;
	wire w_dff_B_Shz1Aqw69_2;
	wire w_dff_B_4e2VIIbb2_2;
	wire w_dff_B_oKTa9Z6e8_2;
	wire w_dff_B_PnGStDAv7_2;
	wire w_dff_B_k2iDG3JR1_2;
	wire w_dff_B_rnu65OlP0_2;
	wire w_dff_B_Y9MhPSzk2_1;
	wire w_dff_B_LIXcAc2O5_2;
	wire w_dff_B_mvFRcGWT2_2;
	wire w_dff_B_onSIMLQJ6_2;
	wire w_dff_B_z7hSY4bY5_2;
	wire w_dff_B_4T76rDuK2_2;
	wire w_dff_B_DlqGR35S1_2;
	wire w_dff_B_IYdwAWZH0_2;
	wire w_dff_B_ypl0N8wR2_2;
	wire w_dff_B_ZHpkIu0s7_2;
	wire w_dff_B_XLpWBxtc2_2;
	wire w_dff_B_hepGxWQP0_2;
	wire w_dff_B_NZTP6NYu9_2;
	wire w_dff_B_fZAO0HLr4_2;
	wire w_dff_B_9ghebZGk8_1;
	wire w_dff_B_lQCrSu5l7_2;
	wire w_dff_B_oIP1yoqL8_2;
	wire w_dff_B_IcS8Xf7q7_2;
	wire w_dff_B_VIutb0F06_2;
	wire w_dff_B_9QkdcicG0_2;
	wire w_dff_B_P5mEoDRL9_2;
	wire w_dff_B_IwPzVIZl5_2;
	wire w_dff_B_a0lQqF4h6_2;
	wire w_dff_B_ldFlnqha2_2;
	wire w_dff_B_2i1IVh7i6_2;
	wire w_dff_B_AaPrnNlc1_2;
	wire w_dff_B_8EbeydnL5_1;
	wire w_dff_B_ttxOODxp4_1;
	wire w_dff_B_SNA3vDRz5_1;
	wire w_dff_B_isjKHTxj5_1;
	wire w_dff_B_3ZRXdkm85_1;
	wire w_dff_B_qyNN8air7_1;
	wire w_dff_B_tFPh4Pe25_0;
	wire w_dff_B_RAreoxw01_0;
	wire w_dff_A_tAE24NYn6_0;
	wire w_dff_A_SiIxT2xb8_0;
	wire w_dff_A_1dQUkF5l2_0;
	wire w_dff_B_N7i4VHMt8_1;
	wire w_dff_A_vbg071tF9_0;
	wire w_dff_A_Wwcu4ipG4_1;
	wire w_dff_A_zMPDIusV4_1;
	wire w_dff_A_W4w189eW0_1;
	wire w_dff_A_a2mVrLoC1_1;
	wire w_dff_A_SrNpZSN95_1;
	wire w_dff_A_Dm8KbRbH0_1;
	wire w_dff_A_smyor4li1_1;
	wire w_dff_A_tRz3lwnQ9_1;
	wire w_dff_B_AsdTUFM99_2;
	wire w_dff_B_YpIpUHEK4_1;
	wire w_dff_B_PArHlcTp7_2;
	wire w_dff_B_qiwI0KSH8_2;
	wire w_dff_B_cKtvtclL9_2;
	wire w_dff_B_0LNSKlF92_2;
	wire w_dff_B_J4sxSRGO4_2;
	wire w_dff_B_z8U5FOiJ5_2;
	wire w_dff_B_dLOTGVoM0_2;
	wire w_dff_B_YlSTYzZj9_2;
	wire w_dff_B_JyIuXjHS8_2;
	wire w_dff_B_YgBJPPjW0_2;
	wire w_dff_B_Szt3aTFi8_2;
	wire w_dff_B_snRKwoe24_2;
	wire w_dff_B_MpW5awIF6_2;
	wire w_dff_B_FxxATGpD3_2;
	wire w_dff_B_amgqkloe2_2;
	wire w_dff_B_WsOKPWoK0_2;
	wire w_dff_B_PEQ2wayV7_2;
	wire w_dff_B_GVk2yZF33_2;
	wire w_dff_B_xDf3TU6n5_2;
	wire w_dff_B_GBlKSAWE9_2;
	wire w_dff_B_V03I3ieu8_2;
	wire w_dff_B_Sd3JDFYY6_2;
	wire w_dff_B_bZJ2N5px0_2;
	wire w_dff_B_AowOnzXc9_2;
	wire w_dff_B_dpQU4WUr3_2;
	wire w_dff_B_s3U6reL44_2;
	wire w_dff_B_P58tzSC07_2;
	wire w_dff_B_5lApa9jI1_2;
	wire w_dff_B_GKWVAdBZ3_2;
	wire w_dff_B_C6jXFXyJ4_2;
	wire w_dff_B_a83QJQJW7_2;
	wire w_dff_B_ImdX8alE0_2;
	wire w_dff_B_N5mzrMAR5_2;
	wire w_dff_B_SC5LjA8y3_2;
	wire w_dff_B_UaAiIiiB6_2;
	wire w_dff_B_ZEMXU4sU1_2;
	wire w_dff_B_r8ryJgr71_2;
	wire w_dff_B_ij2djt9q8_2;
	wire w_dff_B_If8Kb8MC5_2;
	wire w_dff_B_r4cU4sKg0_2;
	wire w_dff_B_i3zVcTM01_2;
	wire w_dff_B_4k1mpOB02_2;
	wire w_dff_B_wykz0jUS4_2;
	wire w_dff_B_4sxKzeg92_2;
	wire w_dff_B_VzGOJpHZ2_2;
	wire w_dff_B_ppU07i4X5_2;
	wire w_dff_B_SOd0D7wR4_2;
	wire w_dff_B_WUkWgVNA1_2;
	wire w_dff_B_okOZllCj2_2;
	wire w_dff_B_BpAGy5bV6_1;
	wire w_dff_A_Wswiurrn4_1;
	wire w_dff_B_5Zokezc54_1;
	wire w_dff_B_EII6tz7c4_2;
	wire w_dff_B_5iBeThyd4_2;
	wire w_dff_B_X06eB6e28_2;
	wire w_dff_B_0Q2tU6qi6_2;
	wire w_dff_B_rCvZpAjm5_2;
	wire w_dff_B_dXyaVulQ1_2;
	wire w_dff_B_FYtV1i0B1_2;
	wire w_dff_B_XEC6lTLt3_2;
	wire w_dff_B_ZMzzyrzm2_2;
	wire w_dff_B_kyp6GfXr6_2;
	wire w_dff_B_4vyHJ6G09_2;
	wire w_dff_B_5SOLiOdu3_2;
	wire w_dff_B_o1GIZ1Sd5_2;
	wire w_dff_B_3la8R4sz0_2;
	wire w_dff_B_hu7kdU4w6_2;
	wire w_dff_B_h07Pw2yX7_2;
	wire w_dff_B_9V2VZvxe5_2;
	wire w_dff_B_ASsZyJm94_2;
	wire w_dff_B_A9yI4gMT4_2;
	wire w_dff_B_u5Omsozp9_2;
	wire w_dff_B_yprUHcKH6_2;
	wire w_dff_B_s3PM9E6V0_2;
	wire w_dff_B_mBAHCuQW4_2;
	wire w_dff_B_wa7If9a09_2;
	wire w_dff_B_ZPzbgEgX5_2;
	wire w_dff_B_GGYKYHp36_2;
	wire w_dff_B_hki1wbsE5_2;
	wire w_dff_B_vSXcGfHH8_2;
	wire w_dff_B_gRcf7Shg7_2;
	wire w_dff_B_YUEU3PB34_2;
	wire w_dff_B_v7IBVsMS7_2;
	wire w_dff_B_jXEB89iI1_2;
	wire w_dff_B_4cQLnrIp3_2;
	wire w_dff_B_k2y5Llhv9_2;
	wire w_dff_B_jzle25lS0_2;
	wire w_dff_B_7j9wF6AW7_2;
	wire w_dff_B_rSElkkp40_2;
	wire w_dff_B_oMDpZC6N7_2;
	wire w_dff_B_nlzTKguN6_2;
	wire w_dff_B_tAEciqjq9_2;
	wire w_dff_B_yrwraxs34_2;
	wire w_dff_B_gOCfkhlM7_2;
	wire w_dff_B_SsRb6lpj6_2;
	wire w_dff_B_2R8NMV0v3_2;
	wire w_dff_B_pagIvr6A9_1;
	wire w_dff_B_TLuVNcfx0_2;
	wire w_dff_B_WRy6xeMn3_2;
	wire w_dff_B_91c7I6DH5_2;
	wire w_dff_B_aBp54Wtv4_2;
	wire w_dff_B_CODpvkFf0_2;
	wire w_dff_B_1iRxiGVT0_2;
	wire w_dff_B_vdQYW4Hw1_2;
	wire w_dff_B_reTqCqZp4_2;
	wire w_dff_B_voqJWS125_2;
	wire w_dff_B_yl3ejYsE6_2;
	wire w_dff_B_kjCn1hoO6_2;
	wire w_dff_B_yuqiEWKI0_2;
	wire w_dff_B_0HFGYiWl6_2;
	wire w_dff_B_oP3nAfxX5_2;
	wire w_dff_B_08jXME4B6_2;
	wire w_dff_B_GMloJzhW1_2;
	wire w_dff_B_pa8eGOHw3_2;
	wire w_dff_B_aGfszCib8_2;
	wire w_dff_B_B2uFpXqJ9_2;
	wire w_dff_B_h0qAKFFr9_2;
	wire w_dff_B_m71BTlAj1_2;
	wire w_dff_B_jamaZ3bo1_2;
	wire w_dff_B_Tc0hrw154_2;
	wire w_dff_B_WsdiyoMh8_2;
	wire w_dff_B_dJOOY7kP7_2;
	wire w_dff_B_tpVz6Gsm7_2;
	wire w_dff_B_55SGtvPf6_2;
	wire w_dff_B_AXwMpPAh1_2;
	wire w_dff_B_0zhgQm5e9_2;
	wire w_dff_B_3qGD6MkH2_2;
	wire w_dff_B_IUUhIEmi9_2;
	wire w_dff_B_jQqc8zqU4_2;
	wire w_dff_B_829tdbsk5_2;
	wire w_dff_B_DTEQhiTy4_2;
	wire w_dff_B_lzgvobre2_2;
	wire w_dff_B_JUoSF68r3_2;
	wire w_dff_B_XK4FhS402_2;
	wire w_dff_B_6mmEAo6i4_2;
	wire w_dff_B_4CzgkvPs3_2;
	wire w_dff_B_K41MyTbU4_1;
	wire w_dff_B_TyK5dQqj5_2;
	wire w_dff_B_arrXisRy6_2;
	wire w_dff_B_Zk13VLht1_2;
	wire w_dff_B_TW86E0Zv5_2;
	wire w_dff_B_9pVyEPLW4_2;
	wire w_dff_B_7s6xVT6I4_2;
	wire w_dff_B_0uIMJlZc9_2;
	wire w_dff_B_AEQteULq6_2;
	wire w_dff_B_mQgpQWQO8_2;
	wire w_dff_B_Du1S8MxW8_2;
	wire w_dff_B_snbtd5uG4_2;
	wire w_dff_B_R7HZpIr20_2;
	wire w_dff_B_QGdQG0sN8_2;
	wire w_dff_B_1JuYYxyY3_2;
	wire w_dff_B_69TUTZL13_2;
	wire w_dff_B_eWu280fD2_2;
	wire w_dff_B_OqfR5k8g6_2;
	wire w_dff_B_Sesxpo9h3_2;
	wire w_dff_B_ozzNEXzh1_2;
	wire w_dff_B_uDazpirA8_2;
	wire w_dff_B_L6QxvCDs1_2;
	wire w_dff_B_ThLEIJR14_2;
	wire w_dff_B_oo2V7gSP7_2;
	wire w_dff_B_eJ8H1CBG3_2;
	wire w_dff_B_SvzLXKei0_2;
	wire w_dff_B_kntGFaS84_2;
	wire w_dff_B_KCi92yq28_2;
	wire w_dff_B_mYEcX1I12_2;
	wire w_dff_B_LZNvlh2l6_2;
	wire w_dff_B_AmcbLqlN5_2;
	wire w_dff_B_avgG7PRt1_2;
	wire w_dff_B_cGP2vjTw7_2;
	wire w_dff_B_Qc3ocyp11_2;
	wire w_dff_B_6Xsy4sUD5_2;
	wire w_dff_B_O80VdUpm7_2;
	wire w_dff_B_itcEa49g7_2;
	wire w_dff_B_bYfsVfi42_2;
	wire w_dff_B_3ivT3rTn6_1;
	wire w_dff_B_flQf7tPn4_2;
	wire w_dff_B_56Pqgc8c1_2;
	wire w_dff_B_7dtkclOw9_2;
	wire w_dff_B_KlDK33Mf7_2;
	wire w_dff_B_eHFgj4Ve3_2;
	wire w_dff_B_d7Wy6wTi6_2;
	wire w_dff_B_D0d9A9qJ6_2;
	wire w_dff_B_P6mjiWLb0_2;
	wire w_dff_B_tBCFtUkA8_2;
	wire w_dff_B_FBTOGR5y4_2;
	wire w_dff_B_V34flryK0_2;
	wire w_dff_B_wdQgBuBB6_2;
	wire w_dff_B_Hgs3QckX9_2;
	wire w_dff_B_sc8IGDxq3_2;
	wire w_dff_B_MwTtwYIr2_2;
	wire w_dff_B_EyFblM9y6_2;
	wire w_dff_B_6MxbI05r8_2;
	wire w_dff_B_VVAKi3DV0_2;
	wire w_dff_B_hk35RDvd0_2;
	wire w_dff_B_PSrJARcw7_2;
	wire w_dff_B_owJ0xV6P1_2;
	wire w_dff_B_376C6p1S1_2;
	wire w_dff_B_tQNyFucx4_2;
	wire w_dff_B_Q4xVar3X0_2;
	wire w_dff_B_a2AdSJ5e5_2;
	wire w_dff_B_rJHnmdi38_2;
	wire w_dff_B_ZgWZNZGs6_2;
	wire w_dff_B_VkjFSMyx0_2;
	wire w_dff_B_mMgjSKlN0_2;
	wire w_dff_B_2cmTMOFd7_2;
	wire w_dff_B_ckOJNAx06_2;
	wire w_dff_B_Zvq4qjqE0_2;
	wire w_dff_B_5S7Cx1Wo0_2;
	wire w_dff_B_eRYndxZQ9_2;
	wire w_dff_B_r1QgCYWE8_1;
	wire w_dff_B_mAp5Wr2U3_2;
	wire w_dff_B_jZRyMvmh3_2;
	wire w_dff_B_xAe6ydeR9_2;
	wire w_dff_B_9EdJwgCh9_2;
	wire w_dff_B_vdzOl8vN5_2;
	wire w_dff_B_eqZXP6sM3_2;
	wire w_dff_B_4D0HCNlm1_2;
	wire w_dff_B_6UWdwD3b1_2;
	wire w_dff_B_JAXKTocg6_2;
	wire w_dff_B_38PoEDjK5_2;
	wire w_dff_B_FDHm8uDc8_2;
	wire w_dff_B_DER76iIo3_2;
	wire w_dff_B_8lS6xrSr4_2;
	wire w_dff_B_4XGQjpMt0_2;
	wire w_dff_B_tOyO4qrW9_2;
	wire w_dff_B_R1BRX1oa3_2;
	wire w_dff_B_l9io95j56_2;
	wire w_dff_B_U2nah3FP2_2;
	wire w_dff_B_ICOJaBic1_2;
	wire w_dff_B_u6t4UeYS9_2;
	wire w_dff_B_iyr9dA2w2_2;
	wire w_dff_B_Gc4LD6193_2;
	wire w_dff_B_PJB8swyl7_2;
	wire w_dff_B_W3BSKrt41_2;
	wire w_dff_B_nnKpUWXO7_2;
	wire w_dff_B_44aVBxuU2_2;
	wire w_dff_B_gllUJLha2_2;
	wire w_dff_B_JofmrGE47_2;
	wire w_dff_B_k60LU9g95_2;
	wire w_dff_B_kFyMKoK27_2;
	wire w_dff_B_bBFQ8uv53_2;
	wire w_dff_B_wagfIO683_1;
	wire w_dff_B_PdHUiMdJ8_2;
	wire w_dff_B_UpRxfvD89_2;
	wire w_dff_B_tkGe4RU20_2;
	wire w_dff_B_wczrDmUN1_2;
	wire w_dff_B_oBmvKOG43_2;
	wire w_dff_B_IEimpLLb4_2;
	wire w_dff_B_RiZfGMyU6_2;
	wire w_dff_B_dJafIPej1_2;
	wire w_dff_B_PA2s1AEB4_2;
	wire w_dff_B_3vqY1THw9_2;
	wire w_dff_B_1dOSfdRo8_2;
	wire w_dff_B_hWh6G7eG3_2;
	wire w_dff_B_LuGowNgP7_2;
	wire w_dff_B_hMAT3ppX4_2;
	wire w_dff_B_hN2Og05J4_2;
	wire w_dff_B_GFGmnGVU7_2;
	wire w_dff_B_D5IPn25S0_2;
	wire w_dff_B_vYPnYFYf5_2;
	wire w_dff_B_eN7zp82a4_2;
	wire w_dff_B_vb6Wdhxy4_2;
	wire w_dff_B_a0kRmkz70_2;
	wire w_dff_B_kQM9N60a5_2;
	wire w_dff_B_U7kB5AXn3_2;
	wire w_dff_B_PKA8kakU5_2;
	wire w_dff_B_1o7Vschu5_2;
	wire w_dff_B_BWgj89hY8_2;
	wire w_dff_B_IwuZxtfj9_2;
	wire w_dff_B_rFjJMvLB6_2;
	wire w_dff_B_xYPBzUfi5_1;
	wire w_dff_B_ZlQXV9LP0_2;
	wire w_dff_B_Oor7oGdn0_2;
	wire w_dff_B_Bh1fsua58_2;
	wire w_dff_B_Jf3z8ZEo1_2;
	wire w_dff_B_n9kziAFO6_2;
	wire w_dff_B_D5EpSTut7_2;
	wire w_dff_B_rsGyHwG74_2;
	wire w_dff_B_rvyRnOh60_2;
	wire w_dff_B_fuDwmqRr1_2;
	wire w_dff_B_Eq7Pr4C17_2;
	wire w_dff_B_IJ0O3Nk72_2;
	wire w_dff_B_KRvi5V9U8_2;
	wire w_dff_B_cukbiTFI2_2;
	wire w_dff_B_pHA1L4m16_2;
	wire w_dff_B_jWlWgwqZ9_2;
	wire w_dff_B_onhZauR79_2;
	wire w_dff_B_U8cur0Jw2_2;
	wire w_dff_B_jnn794fg4_2;
	wire w_dff_B_hxT1HbQd3_2;
	wire w_dff_B_Rv0JryFq4_2;
	wire w_dff_B_k4bGixr26_2;
	wire w_dff_B_7CKXMnQ41_2;
	wire w_dff_B_TsgmmHrT5_2;
	wire w_dff_B_czjghiQe6_2;
	wire w_dff_B_RuQq9Eub5_2;
	wire w_dff_B_pcewXHOL5_1;
	wire w_dff_B_V8XIUyyD9_2;
	wire w_dff_B_mnaP1wgb4_2;
	wire w_dff_B_Zedg13GE5_2;
	wire w_dff_B_D4JC1RTp0_2;
	wire w_dff_B_Xx2gwmqm1_2;
	wire w_dff_B_ZgY6m3Il0_2;
	wire w_dff_B_sgwBHFZn2_2;
	wire w_dff_B_gINrAaA18_2;
	wire w_dff_B_0GOtKah77_2;
	wire w_dff_B_XuSJ6VgI9_2;
	wire w_dff_B_gNIDXnNk7_2;
	wire w_dff_B_VPNAr3yf0_2;
	wire w_dff_B_zyNYa4Zf0_2;
	wire w_dff_B_lZ58jvSi3_2;
	wire w_dff_B_JvaKCZre8_2;
	wire w_dff_B_3vXwOkX01_2;
	wire w_dff_B_ixZqhkfJ8_2;
	wire w_dff_B_TaXcv2j70_2;
	wire w_dff_B_T7MIpknU2_2;
	wire w_dff_B_Dm1VWGbe4_2;
	wire w_dff_B_thbvFUV31_2;
	wire w_dff_B_ao4BY8oo8_2;
	wire w_dff_B_DZRvO2GV2_1;
	wire w_dff_B_tSSnxbXa8_2;
	wire w_dff_B_76t1DMNq6_2;
	wire w_dff_B_6zSNXt7N2_2;
	wire w_dff_B_fteipKbY6_2;
	wire w_dff_B_JfjY3Nog7_2;
	wire w_dff_B_KcNaJbXd4_2;
	wire w_dff_B_MDSMfXng6_2;
	wire w_dff_B_f6n8BLPv9_2;
	wire w_dff_B_3Wyhvwui8_2;
	wire w_dff_B_vvbHeEAI8_2;
	wire w_dff_B_SbSxcFOS3_2;
	wire w_dff_B_kZzSmu0J0_2;
	wire w_dff_B_vlvc2Jgj6_2;
	wire w_dff_B_konWLJGr2_2;
	wire w_dff_B_C7HhDz9u0_2;
	wire w_dff_B_izwclW5u7_2;
	wire w_dff_B_3BVpdZpE4_2;
	wire w_dff_B_DFyjm9Ys5_2;
	wire w_dff_B_pK0UmoXy1_2;
	wire w_dff_B_FCxt0qPm9_1;
	wire w_dff_B_b34qV6ic3_2;
	wire w_dff_B_4YiGYZGb6_2;
	wire w_dff_B_B8NqnJWJ9_2;
	wire w_dff_B_7HJiycvM3_2;
	wire w_dff_B_SzadATYM5_2;
	wire w_dff_B_it1ksGdT6_2;
	wire w_dff_B_RkngrY8w2_2;
	wire w_dff_B_iim0fEk80_2;
	wire w_dff_B_NEwVDMBL5_2;
	wire w_dff_B_UVljeYQg8_2;
	wire w_dff_B_vFP3rCBv2_2;
	wire w_dff_B_Quv42M9X6_2;
	wire w_dff_B_FYcs07zF6_2;
	wire w_dff_B_hh67WdTi6_2;
	wire w_dff_B_zmwDxNgR1_2;
	wire w_dff_B_ybKDPPf21_2;
	wire w_dff_B_GEBf26LN1_1;
	wire w_dff_B_tquyCFwV4_2;
	wire w_dff_B_eQMVtQdk8_2;
	wire w_dff_B_lE8BO4Ak8_2;
	wire w_dff_B_Z4DX1izX5_2;
	wire w_dff_B_tu2IuUGn9_2;
	wire w_dff_B_hmkxXFmX5_2;
	wire w_dff_B_N7Rujm9g6_2;
	wire w_dff_B_PMYZG2Gs1_2;
	wire w_dff_B_H6Hjpk5R6_2;
	wire w_dff_B_neCTmOi35_2;
	wire w_dff_B_6IlgLLGe7_2;
	wire w_dff_B_bFjrIidG9_2;
	wire w_dff_B_4IdKWKoN1_2;
	wire w_dff_B_cAHDlMdl3_1;
	wire w_dff_B_Tmwl9KId3_2;
	wire w_dff_B_kgt4KW890_2;
	wire w_dff_B_BH4dHiRb6_2;
	wire w_dff_B_2OqAu5By9_2;
	wire w_dff_B_tTRWVKnj0_2;
	wire w_dff_B_G2VAy9Qs4_2;
	wire w_dff_B_yZ9mZk8C6_2;
	wire w_dff_B_B6uDATif7_2;
	wire w_dff_B_9ozcuxUk2_2;
	wire w_dff_B_cHkEKdtp7_2;
	wire w_dff_B_pV3RM8kO6_2;
	wire w_dff_B_SSi1Nx618_1;
	wire w_dff_B_PWgDQNB48_1;
	wire w_dff_B_eEqzv1yO6_1;
	wire w_dff_B_NBSVDX3K8_1;
	wire w_dff_B_uawajdVm2_1;
	wire w_dff_B_nDYSgVV54_1;
	wire w_dff_B_1ZmkyheE0_0;
	wire w_dff_B_n7fgtk1y8_0;
	wire w_dff_A_OlbhUUiF2_0;
	wire w_dff_A_bUW1CBpB1_0;
	wire w_dff_A_ORLsOMXy6_0;
	wire w_dff_B_oQXcnDpm6_1;
	wire w_dff_A_TrtfMKBO0_0;
	wire w_dff_A_TiCADdSY4_1;
	wire w_dff_A_hDjMxZIc3_1;
	wire w_dff_A_TAdN2pcZ7_1;
	wire w_dff_A_TpDKr2Pl4_1;
	wire w_dff_A_q3D9U0OS2_1;
	wire w_dff_A_tlK2ukNF8_1;
	wire w_dff_A_fmims8R39_1;
	wire w_dff_A_rAkL1biL0_1;
	wire w_dff_B_ujHNKIta2_1;
	wire w_dff_A_KO0EuAWu9_1;
	wire w_dff_B_apJ5POHG4_1;
	wire w_dff_B_9xz2TAaz5_2;
	wire w_dff_B_osJnFlgF0_2;
	wire w_dff_B_oLKqF3Bw1_2;
	wire w_dff_B_q9exviJh9_2;
	wire w_dff_B_MbBfWPil6_2;
	wire w_dff_B_3CSI38gN1_2;
	wire w_dff_B_LjxN97AI1_2;
	wire w_dff_B_sdzPZ9Sw3_2;
	wire w_dff_B_CPsJ53rU2_2;
	wire w_dff_B_la46kmkC6_2;
	wire w_dff_B_Y1iJcdN41_2;
	wire w_dff_B_mtLx5q6a1_2;
	wire w_dff_B_QPk1gBoU5_2;
	wire w_dff_B_GUxVZLTq6_2;
	wire w_dff_B_HxGEV71P4_2;
	wire w_dff_B_UUFraiRB4_2;
	wire w_dff_B_Muyuscta5_2;
	wire w_dff_B_LZdvBhbe2_2;
	wire w_dff_B_l2uNAhBI8_2;
	wire w_dff_B_FcDlXBvW1_2;
	wire w_dff_B_3fxmqe3e9_2;
	wire w_dff_B_yho9OXWh9_2;
	wire w_dff_B_CBHIiu7x3_2;
	wire w_dff_B_F1Bx0yKk5_2;
	wire w_dff_B_e92sGs230_2;
	wire w_dff_B_DAIOBDHK2_2;
	wire w_dff_B_1ovJIxFL4_2;
	wire w_dff_B_SWDD36d69_2;
	wire w_dff_B_7LPw1nqW3_2;
	wire w_dff_B_HyHON5LR1_2;
	wire w_dff_B_Bvfy7t9D9_2;
	wire w_dff_B_En6pPMKo1_2;
	wire w_dff_B_o50OStId1_2;
	wire w_dff_B_3DSU8NNU4_2;
	wire w_dff_B_Bd7DnAjV1_2;
	wire w_dff_B_0Xxlr55z2_2;
	wire w_dff_B_mm9FWPiT4_2;
	wire w_dff_B_qFm6eFQb1_2;
	wire w_dff_B_w9Maiqfx9_2;
	wire w_dff_B_nHcQtLIw8_2;
	wire w_dff_B_N0VRdw9b2_2;
	wire w_dff_B_DSx5GGT06_2;
	wire w_dff_B_Qa1UIgWT5_2;
	wire w_dff_B_a1ZSYa9u1_2;
	wire w_dff_B_qhsrqwUt1_2;
	wire w_dff_B_XK2uILrM8_2;
	wire w_dff_B_2XFUkYcT6_2;
	wire w_dff_B_xiZ0u1Xr4_2;
	wire w_dff_B_Md1qSbaj1_2;
	wire w_dff_B_GZgJyiDF4_2;
	wire w_dff_B_rH54O8kr0_1;
	wire w_dff_B_k66MwJLp8_2;
	wire w_dff_B_bkeVVpIO9_2;
	wire w_dff_B_4pebG2L49_2;
	wire w_dff_B_J1VdQMTL7_2;
	wire w_dff_B_fb4IbUOw3_2;
	wire w_dff_B_FrA7bjqF2_2;
	wire w_dff_B_CovZDhnp4_2;
	wire w_dff_B_lrlDqXVL1_2;
	wire w_dff_B_psq5de8v6_2;
	wire w_dff_B_Vz4VUZNa6_2;
	wire w_dff_B_zZi9vpUJ3_2;
	wire w_dff_B_bei4QNnw6_2;
	wire w_dff_B_9PYZaKk22_2;
	wire w_dff_B_MACv1VX81_2;
	wire w_dff_B_bmuiqEK48_2;
	wire w_dff_B_RXpBW1OE1_2;
	wire w_dff_B_cMAqL4IR1_2;
	wire w_dff_B_UdPbB9rR5_2;
	wire w_dff_B_z6YKWQYh4_2;
	wire w_dff_B_B59K5Qmb4_2;
	wire w_dff_B_zl22vhKO1_2;
	wire w_dff_B_MD0eqtep3_2;
	wire w_dff_B_wtVkrcJt5_2;
	wire w_dff_B_K42KxeUG1_2;
	wire w_dff_B_9UR64zlS8_2;
	wire w_dff_B_pAWjWLdN1_2;
	wire w_dff_B_MRoQTFT48_2;
	wire w_dff_B_mMoH7CHO8_2;
	wire w_dff_B_xaz2qoEw2_2;
	wire w_dff_B_BwYFzB2s0_2;
	wire w_dff_B_1RZ1TZC06_2;
	wire w_dff_B_8vJGM7z75_2;
	wire w_dff_B_t9uBPWse6_2;
	wire w_dff_B_Zoo3vDB21_2;
	wire w_dff_B_Nge3wDfC4_2;
	wire w_dff_B_16v6yqL68_2;
	wire w_dff_B_qo7QaHEe8_2;
	wire w_dff_B_mJYvVkCf4_2;
	wire w_dff_B_0h7UaMMb7_2;
	wire w_dff_B_IAqsdOpI8_2;
	wire w_dff_B_CUFAMhhL3_2;
	wire w_dff_B_rxe1wSSc2_2;
	wire w_dff_B_YdhuBDJN6_2;
	wire w_dff_B_gLWcJpwC8_2;
	wire w_dff_B_vDxlcce85_2;
	wire w_dff_B_uIBjKJe90_2;
	wire w_dff_B_UDKKrrrV9_1;
	wire w_dff_B_bO1HDDwj3_2;
	wire w_dff_B_chIXy3lL2_2;
	wire w_dff_B_r3Gu3hpD8_2;
	wire w_dff_B_qpJxfoZs3_2;
	wire w_dff_B_NKy6GcsM3_2;
	wire w_dff_B_BxgWGTsK4_2;
	wire w_dff_B_BDbAN8D03_2;
	wire w_dff_B_WyaPA5Ay1_2;
	wire w_dff_B_rumB24580_2;
	wire w_dff_B_IoaFiZMh7_2;
	wire w_dff_B_3reBQm4S5_2;
	wire w_dff_B_hKVPuUGl2_2;
	wire w_dff_B_w2onzORz0_2;
	wire w_dff_B_Wu3zD1GT5_2;
	wire w_dff_B_3oRQ7EPQ5_2;
	wire w_dff_B_V2T2MCnd2_2;
	wire w_dff_B_D62z7zpH8_2;
	wire w_dff_B_xO1lNm0a8_2;
	wire w_dff_B_RcoLN56Y8_2;
	wire w_dff_B_9Sfyq3fq3_2;
	wire w_dff_B_GCtRIySl5_2;
	wire w_dff_B_Rxzq6Hj58_2;
	wire w_dff_B_MVwDUCoH2_2;
	wire w_dff_B_U4ZsiqT29_2;
	wire w_dff_B_21KJvFnr3_2;
	wire w_dff_B_HWFBSknv5_2;
	wire w_dff_B_f0A0QqQH0_2;
	wire w_dff_B_vjyf2qyx1_2;
	wire w_dff_B_QlaCx6Ry9_2;
	wire w_dff_B_UH0OclH40_2;
	wire w_dff_B_Q67uGzm68_2;
	wire w_dff_B_EaeVlffx3_2;
	wire w_dff_B_Onr2JCiq4_2;
	wire w_dff_B_waqcrjzC2_2;
	wire w_dff_B_jPtQqvO00_2;
	wire w_dff_B_noyzE1Lq2_2;
	wire w_dff_B_atTiopd40_2;
	wire w_dff_B_czSDJJiW8_2;
	wire w_dff_B_bAjjmrUk2_2;
	wire w_dff_B_HzXNkwGQ5_2;
	wire w_dff_B_ZP7WsaNU0_2;
	wire w_dff_B_diTzV2yZ9_2;
	wire w_dff_B_WXGUjXj40_1;
	wire w_dff_B_5ppg6Ajf3_2;
	wire w_dff_B_W7yAxnHD6_2;
	wire w_dff_B_5NqwLzV36_2;
	wire w_dff_B_CeGX5VUo4_2;
	wire w_dff_B_GHlkrBiz1_2;
	wire w_dff_B_OR7FTlHf7_2;
	wire w_dff_B_kSwtPMCL1_2;
	wire w_dff_B_mlEsU0SL2_2;
	wire w_dff_B_RwDcWrAK2_2;
	wire w_dff_B_h1NsZ8C62_2;
	wire w_dff_B_stCasSyO9_2;
	wire w_dff_B_KvRttgXt2_2;
	wire w_dff_B_FfBVZBr27_2;
	wire w_dff_B_0soXRjRa4_2;
	wire w_dff_B_z4tShkuq0_2;
	wire w_dff_B_Wmm1juw91_2;
	wire w_dff_B_4Uowic3k0_2;
	wire w_dff_B_S1lm61At7_2;
	wire w_dff_B_pChfuww06_2;
	wire w_dff_B_qgAKR1ne5_2;
	wire w_dff_B_SYWtNSKa2_2;
	wire w_dff_B_xd8kkPwt5_2;
	wire w_dff_B_LQgl3NRM4_2;
	wire w_dff_B_oyWHq5wA9_2;
	wire w_dff_B_bnUwPA7f9_2;
	wire w_dff_B_2sJRKZjp7_2;
	wire w_dff_B_grEGwFDf6_2;
	wire w_dff_B_L9PRyrWY3_2;
	wire w_dff_B_M7FDF4N17_2;
	wire w_dff_B_VI1Dtueh6_2;
	wire w_dff_B_Gnz4gFRi6_2;
	wire w_dff_B_seSrTjLh5_2;
	wire w_dff_B_aYfvuTza0_2;
	wire w_dff_B_LIo79Tfs1_2;
	wire w_dff_B_zHXtUCGX5_2;
	wire w_dff_B_Luf9Nf274_2;
	wire w_dff_B_vWEqRT4V1_2;
	wire w_dff_B_IcO8rX5a7_2;
	wire w_dff_B_dEwrKoGB5_1;
	wire w_dff_B_j5H20azp7_2;
	wire w_dff_B_F5wZsKrk6_2;
	wire w_dff_B_nw90zict1_2;
	wire w_dff_B_7vDRSFeR0_2;
	wire w_dff_B_wHzxIEBr5_2;
	wire w_dff_B_Mc71VNGq4_2;
	wire w_dff_B_oNbjh2yC5_2;
	wire w_dff_B_nGTDOzjN8_2;
	wire w_dff_B_taxqBUud3_2;
	wire w_dff_B_9yUfE9mN0_2;
	wire w_dff_B_elH7HKcZ1_2;
	wire w_dff_B_QeYhkzT07_2;
	wire w_dff_B_XnRU8dS32_2;
	wire w_dff_B_kuokYYNo3_2;
	wire w_dff_B_YDfAOY1p7_2;
	wire w_dff_B_veox868p9_2;
	wire w_dff_B_nvOSqB0B4_2;
	wire w_dff_B_7uh7XS7l9_2;
	wire w_dff_B_4BSMdsXu5_2;
	wire w_dff_B_LEs3JQ704_2;
	wire w_dff_B_pnvOZK6z4_2;
	wire w_dff_B_0ajzQRWW9_2;
	wire w_dff_B_6IVayNTO5_2;
	wire w_dff_B_j4aMwnCJ3_2;
	wire w_dff_B_IrdULxle6_2;
	wire w_dff_B_PlYmr6iJ2_2;
	wire w_dff_B_h2itkcX45_2;
	wire w_dff_B_kleeMFqW0_2;
	wire w_dff_B_wcWwAPLW3_2;
	wire w_dff_B_2AjHcWcm6_2;
	wire w_dff_B_9dZpEyNN0_2;
	wire w_dff_B_MiSq2gaE4_2;
	wire w_dff_B_Lm7RFGGj8_2;
	wire w_dff_B_6TwkF4Yo1_1;
	wire w_dff_B_svmI7hRn1_2;
	wire w_dff_B_RlCsqdxM7_2;
	wire w_dff_B_O6OPwk9x2_2;
	wire w_dff_B_ebBitJCz4_2;
	wire w_dff_B_WmmHSPAr8_2;
	wire w_dff_B_TIBZ03Xc2_2;
	wire w_dff_B_zG5oYa8T0_2;
	wire w_dff_B_N3keFv7v3_2;
	wire w_dff_B_nzvJ5CoE7_2;
	wire w_dff_B_uBSzNkwD9_2;
	wire w_dff_B_FFkodaBl1_2;
	wire w_dff_B_MtD9L4fq2_2;
	wire w_dff_B_wtNZsY9p5_2;
	wire w_dff_B_H4qA5dOq5_2;
	wire w_dff_B_imVBRHtE0_2;
	wire w_dff_B_20nZ7xzd7_2;
	wire w_dff_B_pIx08jGb9_2;
	wire w_dff_B_SIWUZzmW4_2;
	wire w_dff_B_Ub0zW7589_2;
	wire w_dff_B_QXuqqmhL8_2;
	wire w_dff_B_jzJVLdmV8_2;
	wire w_dff_B_2A2K6pco0_2;
	wire w_dff_B_Q6e4xXjn6_2;
	wire w_dff_B_pJ6jJO6X4_2;
	wire w_dff_B_Giaq3oEH5_2;
	wire w_dff_B_F1pyfHCD8_2;
	wire w_dff_B_LFCXrPL63_2;
	wire w_dff_B_OG3yEUGn6_2;
	wire w_dff_B_DeO4FRWO6_2;
	wire w_dff_B_vCLHSOEX6_2;
	wire w_dff_B_sSCut7rS2_2;
	wire w_dff_B_bemMx2d96_1;
	wire w_dff_B_4AC5pT9Q8_2;
	wire w_dff_B_28tN70Jt4_2;
	wire w_dff_B_XigzSZeI8_2;
	wire w_dff_B_7087JP5Z0_2;
	wire w_dff_B_FZvQ8w9q8_2;
	wire w_dff_B_ljSEm1H61_2;
	wire w_dff_B_YW2hYdpE4_2;
	wire w_dff_B_kMFhGTuv6_2;
	wire w_dff_B_aA8uHYOJ9_2;
	wire w_dff_B_a09USQzg9_2;
	wire w_dff_B_HlBs94x52_2;
	wire w_dff_B_RjlK8Ewe4_2;
	wire w_dff_B_0gwwOZZh3_2;
	wire w_dff_B_5b65wC8t8_2;
	wire w_dff_B_Aqt3R2jC1_2;
	wire w_dff_B_6rSPOryw7_2;
	wire w_dff_B_4sbSCeOV9_2;
	wire w_dff_B_Ucw76F171_2;
	wire w_dff_B_vfiwW1cI5_2;
	wire w_dff_B_BaPgsUkv8_2;
	wire w_dff_B_C0w1Xh9z6_2;
	wire w_dff_B_ySMyQfaL6_2;
	wire w_dff_B_xger0zA40_2;
	wire w_dff_B_2qLdy5R17_2;
	wire w_dff_B_7UwSXrye8_2;
	wire w_dff_B_7ol1otzE3_2;
	wire w_dff_B_MuvFa1BM3_2;
	wire w_dff_B_KrtcCkho1_2;
	wire w_dff_B_Mhl3G5ff3_1;
	wire w_dff_B_JF4915eS3_2;
	wire w_dff_B_jpfrmX392_2;
	wire w_dff_B_WGARxPBc3_2;
	wire w_dff_B_z25QBqam0_2;
	wire w_dff_B_o9T6pYs51_2;
	wire w_dff_B_90HNUajS3_2;
	wire w_dff_B_AzmHqcUH8_2;
	wire w_dff_B_RKOPdOCw7_2;
	wire w_dff_B_dQdVIRSe7_2;
	wire w_dff_B_EIJQmjBq7_2;
	wire w_dff_B_mHWjMcIl5_2;
	wire w_dff_B_3706xz309_2;
	wire w_dff_B_aXZB5NRb8_2;
	wire w_dff_B_9k1Sy2v61_2;
	wire w_dff_B_8OYUEyyz1_2;
	wire w_dff_B_jmNlidCd0_2;
	wire w_dff_B_0SJ0gnuq1_2;
	wire w_dff_B_yFFtZVHl8_2;
	wire w_dff_B_I4HaKqUQ0_2;
	wire w_dff_B_zZLvfhrD0_2;
	wire w_dff_B_NmKAB2KR4_2;
	wire w_dff_B_q5mlOs9c6_2;
	wire w_dff_B_IgJPhkhL0_2;
	wire w_dff_B_Qb35jaaX6_2;
	wire w_dff_B_26ORQgZm0_2;
	wire w_dff_B_y1QTgYa17_1;
	wire w_dff_B_3I0pdiAz6_2;
	wire w_dff_B_Qwey936N3_2;
	wire w_dff_B_BGGLXxHc5_2;
	wire w_dff_B_pdzRoFHZ1_2;
	wire w_dff_B_D8daikzJ5_2;
	wire w_dff_B_Wduch9Zu9_2;
	wire w_dff_B_92e2RsYI5_2;
	wire w_dff_B_9tTjV6HB5_2;
	wire w_dff_B_PhXhOdmP9_2;
	wire w_dff_B_gFxfOnAp5_2;
	wire w_dff_B_6VfZPh0A2_2;
	wire w_dff_B_DfHUZZgs5_2;
	wire w_dff_B_fRkCD2Mu6_2;
	wire w_dff_B_GGbfKkwR8_2;
	wire w_dff_B_yf7b5EYl3_2;
	wire w_dff_B_jGHlGI6w4_2;
	wire w_dff_B_47WLpT4Z0_2;
	wire w_dff_B_c259OeZs9_2;
	wire w_dff_B_9gvvRstr6_2;
	wire w_dff_B_ctAfkzK51_2;
	wire w_dff_B_E8f9MlnF1_2;
	wire w_dff_B_zGdvxZ9X5_2;
	wire w_dff_B_ITjObB5K9_1;
	wire w_dff_B_N7TCNxmV2_2;
	wire w_dff_B_6RLHAqst4_2;
	wire w_dff_B_weu18uus0_2;
	wire w_dff_B_dMckLTxl9_2;
	wire w_dff_B_YYehwJwc0_2;
	wire w_dff_B_GE8Zn5Oz5_2;
	wire w_dff_B_BhW9enfR8_2;
	wire w_dff_B_FtgXLwPf4_2;
	wire w_dff_B_2HUK1EPC7_2;
	wire w_dff_B_LIsFbDa67_2;
	wire w_dff_B_x61XG7fo3_2;
	wire w_dff_B_YdDsdxE02_2;
	wire w_dff_B_jY7xnavw9_2;
	wire w_dff_B_82ANAqHI4_2;
	wire w_dff_B_JLQenPXC9_2;
	wire w_dff_B_DaNXQWe25_2;
	wire w_dff_B_868EQ2Rv7_2;
	wire w_dff_B_ZWgEyIQa3_2;
	wire w_dff_B_CvCblr1X9_2;
	wire w_dff_B_UnQj650K1_1;
	wire w_dff_B_lSW0Sf5z8_2;
	wire w_dff_B_As7dHRBf6_2;
	wire w_dff_B_y7zUfQeL0_2;
	wire w_dff_B_q9xohqDe9_2;
	wire w_dff_B_7Ck9HBFN0_2;
	wire w_dff_B_5uZJCWtN4_2;
	wire w_dff_B_KK6Lbwbz1_2;
	wire w_dff_B_76jY0EUF1_2;
	wire w_dff_B_kM1yDmwx5_2;
	wire w_dff_B_nUDDhB3m6_2;
	wire w_dff_B_6C7m0p0u1_2;
	wire w_dff_B_FAL7FRdG4_2;
	wire w_dff_B_kOQqsB679_2;
	wire w_dff_B_AB5qckfb4_2;
	wire w_dff_B_iSePcQlc6_2;
	wire w_dff_B_r3cc26Gc8_2;
	wire w_dff_B_A83BQhCB9_1;
	wire w_dff_B_BTA1Y7983_2;
	wire w_dff_B_dod5aWcE3_2;
	wire w_dff_B_TEBdbmRm8_2;
	wire w_dff_B_HJa9TXUS7_2;
	wire w_dff_B_KBNOUwhS6_2;
	wire w_dff_B_WXsuBGhM2_2;
	wire w_dff_B_hIgtUtU92_2;
	wire w_dff_B_R8KQHlkm7_2;
	wire w_dff_B_uCaSF1VP0_2;
	wire w_dff_B_sAONswcD3_2;
	wire w_dff_B_hPr8WnV05_2;
	wire w_dff_B_AxSNxK3Y9_2;
	wire w_dff_B_RFXlgBXa0_2;
	wire w_dff_B_0sWTkjSX6_1;
	wire w_dff_B_Nw7rkneU4_2;
	wire w_dff_B_aX5oDOtj1_2;
	wire w_dff_B_gRw1XyA56_2;
	wire w_dff_B_ri45ITj27_2;
	wire w_dff_B_0SiDLvBJ1_2;
	wire w_dff_B_0WmB5jlO3_2;
	wire w_dff_B_q6eho9w43_2;
	wire w_dff_B_sMHNr9xq6_2;
	wire w_dff_B_3vDR8Cz34_2;
	wire w_dff_B_rAYZzfgx4_2;
	wire w_dff_B_zqjynpTp0_2;
	wire w_dff_B_f5CxgFtA9_1;
	wire w_dff_B_PdCCOk0H0_1;
	wire w_dff_B_ZcJnCOHM2_1;
	wire w_dff_B_3NgXzHpP7_1;
	wire w_dff_B_kZNmdq1V6_1;
	wire w_dff_B_1BovEjzp0_1;
	wire w_dff_B_PFpMQHd80_0;
	wire w_dff_B_oqDe2AjM2_0;
	wire w_dff_A_z98Y48qf6_0;
	wire w_dff_A_d6xTdqEj1_0;
	wire w_dff_A_p1ExIVA06_0;
	wire w_dff_B_TWlLduFk8_1;
	wire w_dff_A_okRv4hTg5_0;
	wire w_dff_A_DVRWxS9i3_1;
	wire w_dff_A_w7exM3Ua5_1;
	wire w_dff_A_LWJKdsaV1_1;
	wire w_dff_A_uvCOXY9n2_1;
	wire w_dff_A_Eai8yYZ14_1;
	wire w_dff_A_9Ad9Y1rS2_1;
	wire w_dff_A_rB9uUE8L9_1;
	wire w_dff_A_uAiNKDt00_1;
	wire w_dff_B_zTqoFgxU7_1;
	wire w_dff_A_9n7XV7sv6_1;
	wire w_dff_B_K1E8wuCf6_1;
	wire w_dff_B_SkQNsE0M6_2;
	wire w_dff_B_w3i1aKTt9_2;
	wire w_dff_B_hCIO0l0H0_2;
	wire w_dff_B_HUsAG0Bc3_2;
	wire w_dff_B_sDwQ91w46_2;
	wire w_dff_B_JuYwKgke5_2;
	wire w_dff_B_yZashIj38_2;
	wire w_dff_B_DWfgVCHX7_2;
	wire w_dff_B_Yc5Rit5X9_2;
	wire w_dff_B_aqevY56E3_2;
	wire w_dff_B_1izovzXb4_2;
	wire w_dff_B_xk8K3NKn4_2;
	wire w_dff_B_NW2TZ1SI7_2;
	wire w_dff_B_ow8MaT5U3_2;
	wire w_dff_B_ok1lrZg16_2;
	wire w_dff_B_YljKQU2P6_2;
	wire w_dff_B_YqoBb55R4_2;
	wire w_dff_B_ekYBECWE4_2;
	wire w_dff_B_vnu85MWu4_2;
	wire w_dff_B_KumHp6UV7_2;
	wire w_dff_B_G3nIlvgo2_2;
	wire w_dff_B_MY3V3YK05_2;
	wire w_dff_B_wgqfjphk6_2;
	wire w_dff_B_SQUwVAfB3_2;
	wire w_dff_B_6A4tvn5k5_2;
	wire w_dff_B_6P8tyPpl9_2;
	wire w_dff_B_J8XDlvFm4_2;
	wire w_dff_B_c7t0rdZN5_2;
	wire w_dff_B_hBHlLwk92_2;
	wire w_dff_B_1GkWyzn78_2;
	wire w_dff_B_JxF8Aspo5_2;
	wire w_dff_B_UvdGenDh4_2;
	wire w_dff_B_evC6RRMu9_2;
	wire w_dff_B_6FPuRBBm1_2;
	wire w_dff_B_MzHYpbmN9_2;
	wire w_dff_B_691UAJeL7_2;
	wire w_dff_B_VPRZIXJZ7_2;
	wire w_dff_B_DtWwtbae9_2;
	wire w_dff_B_flGWL8Yd0_2;
	wire w_dff_B_0b1gWJAs8_2;
	wire w_dff_B_aMeCVaG10_2;
	wire w_dff_B_AhiHYvNf7_2;
	wire w_dff_B_5uCvNK794_2;
	wire w_dff_B_Ha2VZqoK3_2;
	wire w_dff_B_usbleS4f2_2;
	wire w_dff_B_omIE2QMI7_2;
	wire w_dff_B_T22nB26N6_2;
	wire w_dff_B_Jky6HVNF1_2;
	wire w_dff_B_8qzRylMw2_2;
	wire w_dff_B_wLlSA1MN9_2;
	wire w_dff_B_YqZFdzjd8_2;
	wire w_dff_B_eWqtMJtR2_2;
	wire w_dff_B_tYvUEpmN3_1;
	wire w_dff_B_xjz1kvxf4_2;
	wire w_dff_B_UKazAOJP9_2;
	wire w_dff_B_QZTb955o4_2;
	wire w_dff_B_u8kKB4xi8_2;
	wire w_dff_B_WDQG8Xzs0_2;
	wire w_dff_B_PNBdtUvD7_2;
	wire w_dff_B_8RhFjxJJ7_2;
	wire w_dff_B_IQTDBg2f4_2;
	wire w_dff_B_ORLxoJ2g3_2;
	wire w_dff_B_uLUTfVXl5_2;
	wire w_dff_B_hcNAJMin2_2;
	wire w_dff_B_iAY9FUAB4_2;
	wire w_dff_B_bDhbvrd39_2;
	wire w_dff_B_Pz7ULMi99_2;
	wire w_dff_B_3duShExP0_2;
	wire w_dff_B_0bIIEBpI1_2;
	wire w_dff_B_nFbHJGNl0_2;
	wire w_dff_B_lwGAUJsl3_2;
	wire w_dff_B_BEXyloxr5_2;
	wire w_dff_B_wEf2Nuqw1_2;
	wire w_dff_B_GlXLRHWq2_2;
	wire w_dff_B_KRHJzMcj7_2;
	wire w_dff_B_gcwYpLyo3_2;
	wire w_dff_B_eQ0q6MuY7_2;
	wire w_dff_B_dENTBUA79_2;
	wire w_dff_B_3dOZS4Kg8_2;
	wire w_dff_B_dsDenCKx9_2;
	wire w_dff_B_RKUxxegn4_2;
	wire w_dff_B_znAGUxhz9_2;
	wire w_dff_B_Cif6COd73_2;
	wire w_dff_B_hJMqL0hB1_2;
	wire w_dff_B_4IzAYm0o3_2;
	wire w_dff_B_C2COPUGV2_2;
	wire w_dff_B_xHxTZdoA7_2;
	wire w_dff_B_FU12nnqy4_2;
	wire w_dff_B_K6mIsrgp0_2;
	wire w_dff_B_BRnou9A14_2;
	wire w_dff_B_Rq0sGR780_2;
	wire w_dff_B_V0WEGXW86_2;
	wire w_dff_B_CCNeJ2CH6_2;
	wire w_dff_B_pXd4sEYr6_2;
	wire w_dff_B_avZv5ACW8_2;
	wire w_dff_B_bexQZ2CP0_2;
	wire w_dff_B_X1U51X8C8_2;
	wire w_dff_B_fxO94WAp4_2;
	wire w_dff_B_2nJbfz1l7_2;
	wire w_dff_B_wWyQm1T04_2;
	wire w_dff_B_EzRe3tCe8_2;
	wire w_dff_B_JljeUlJQ0_1;
	wire w_dff_B_DBqr7t5P3_2;
	wire w_dff_B_M2vUMp7K1_2;
	wire w_dff_B_CpigqGl21_2;
	wire w_dff_B_WNmUCUVW1_2;
	wire w_dff_B_wAIm0fYC7_2;
	wire w_dff_B_bGz67cqn3_2;
	wire w_dff_B_gpBi5Byj0_2;
	wire w_dff_B_gzDQXrBx2_2;
	wire w_dff_B_BnwCrT4V8_2;
	wire w_dff_B_MZ78ol9p4_2;
	wire w_dff_B_64QAvVpK5_2;
	wire w_dff_B_T2tIO3I22_2;
	wire w_dff_B_Xk6LG3D73_2;
	wire w_dff_B_i1Z1PAty5_2;
	wire w_dff_B_6sv6gaOj2_2;
	wire w_dff_B_DAj1jKV31_2;
	wire w_dff_B_ZxYpR0Ov1_2;
	wire w_dff_B_yPsvRPbX9_2;
	wire w_dff_B_gcJvnEP77_2;
	wire w_dff_B_6GfsG9kL5_2;
	wire w_dff_B_07glfzRU9_2;
	wire w_dff_B_YDRyvsVQ5_2;
	wire w_dff_B_VJRMPvHG5_2;
	wire w_dff_B_Xk2AC1qs0_2;
	wire w_dff_B_X5ev7AnE6_2;
	wire w_dff_B_AKFIMH0n2_2;
	wire w_dff_B_RUUmnh4T6_2;
	wire w_dff_B_KEa06emA7_2;
	wire w_dff_B_xXSYyKvA2_2;
	wire w_dff_B_iI8u8BKe5_2;
	wire w_dff_B_UjUHYEMc3_2;
	wire w_dff_B_6bZtp23N2_2;
	wire w_dff_B_C2SozrwU2_2;
	wire w_dff_B_NFZfAwyU8_2;
	wire w_dff_B_WQKBUYiM7_2;
	wire w_dff_B_2Js7OGcF1_2;
	wire w_dff_B_2Q56mQTX6_2;
	wire w_dff_B_oirdcrNs4_2;
	wire w_dff_B_6e6IMxZ20_2;
	wire w_dff_B_NeaCHM014_2;
	wire w_dff_B_K1KHXBW88_2;
	wire w_dff_B_ChUkjOSL6_2;
	wire w_dff_B_dz0k26vB2_2;
	wire w_dff_B_tEmEHAdO5_2;
	wire w_dff_B_PuxHg3Gn7_1;
	wire w_dff_B_NiV5Ry3s4_2;
	wire w_dff_B_MbTDFteX9_2;
	wire w_dff_B_z9ZR1lCT3_2;
	wire w_dff_B_cBvxXdsU4_2;
	wire w_dff_B_cLGkST2x8_2;
	wire w_dff_B_Ut6etf7H3_2;
	wire w_dff_B_KA75vRZH2_2;
	wire w_dff_B_hhQWxWsW0_2;
	wire w_dff_B_g9cGFbmd5_2;
	wire w_dff_B_n4Th0laP3_2;
	wire w_dff_B_xuof9Mpq7_2;
	wire w_dff_B_7XlAPCrD7_2;
	wire w_dff_B_OAyvb5cV0_2;
	wire w_dff_B_jazKxcXp4_2;
	wire w_dff_B_Al86i8bD1_2;
	wire w_dff_B_AlLf2q5C1_2;
	wire w_dff_B_ZItTtAfd6_2;
	wire w_dff_B_JMKddtrc4_2;
	wire w_dff_B_ACa5mpu87_2;
	wire w_dff_B_SGuNUVAz9_2;
	wire w_dff_B_nZCvjOUe4_2;
	wire w_dff_B_7AFXXhwe9_2;
	wire w_dff_B_FLGJ8WNf6_2;
	wire w_dff_B_yLdseEDo5_2;
	wire w_dff_B_7057YDcd2_2;
	wire w_dff_B_y4Yu8g8X3_2;
	wire w_dff_B_Gl3NF1rb1_2;
	wire w_dff_B_e8DEKZqL1_2;
	wire w_dff_B_xqymBRys9_2;
	wire w_dff_B_wxedBgbg0_2;
	wire w_dff_B_2VWZ8N0X9_2;
	wire w_dff_B_LY4kAkbG8_2;
	wire w_dff_B_o6OC3ZCQ1_2;
	wire w_dff_B_XdqYoZuF3_2;
	wire w_dff_B_jAHP4GMu9_2;
	wire w_dff_B_NVPOjIt99_2;
	wire w_dff_B_iW66WLK87_2;
	wire w_dff_B_VEHPxe3j2_2;
	wire w_dff_B_Sddow3bz4_2;
	wire w_dff_B_LAskapZm5_2;
	wire w_dff_B_OAaZjvPj1_1;
	wire w_dff_B_YvArSvkU1_2;
	wire w_dff_B_9Amf4eFI1_2;
	wire w_dff_B_b1Yq46iO8_2;
	wire w_dff_B_PBDpsqR14_2;
	wire w_dff_B_dt0BS1H90_2;
	wire w_dff_B_tejImq9y6_2;
	wire w_dff_B_5dEDRGNQ8_2;
	wire w_dff_B_X2H6td5e5_2;
	wire w_dff_B_pTLxAzCZ9_2;
	wire w_dff_B_GDvjLGlX3_2;
	wire w_dff_B_EN1qjhzT2_2;
	wire w_dff_B_VmMD9niZ8_2;
	wire w_dff_B_a7geb3ul0_2;
	wire w_dff_B_6fKO13WA4_2;
	wire w_dff_B_ywRatiSP5_2;
	wire w_dff_B_HQ2tvnZ50_2;
	wire w_dff_B_QG5kuPBS3_2;
	wire w_dff_B_CD3OADq45_2;
	wire w_dff_B_zYpnQ2Ig0_2;
	wire w_dff_B_cEGvPtLY2_2;
	wire w_dff_B_oirJ4AZ60_2;
	wire w_dff_B_hGizR7cq6_2;
	wire w_dff_B_qJeZbiVS0_2;
	wire w_dff_B_SV8i3JPX5_2;
	wire w_dff_B_cDQJ7fM50_2;
	wire w_dff_B_P5cb6zY73_2;
	wire w_dff_B_vDXw7Xci5_2;
	wire w_dff_B_HqQiNcsV3_2;
	wire w_dff_B_acsSjEvN0_2;
	wire w_dff_B_hvPFtZkC6_2;
	wire w_dff_B_HciZw9o28_2;
	wire w_dff_B_xbllgv9y5_2;
	wire w_dff_B_hQ5NkmOB9_2;
	wire w_dff_B_jLRC9c199_2;
	wire w_dff_B_y9GIDU0I4_2;
	wire w_dff_B_uIocQ37G6_2;
	wire w_dff_B_ojVnhXCC2_1;
	wire w_dff_B_daI1jvuT4_2;
	wire w_dff_B_sAPYZK8Y7_2;
	wire w_dff_B_Gk4uQ0640_2;
	wire w_dff_B_LmAKy6Eo2_2;
	wire w_dff_B_QrPblEgJ0_2;
	wire w_dff_B_207anArg1_2;
	wire w_dff_B_pAbdW2I46_2;
	wire w_dff_B_zvHk8ibg3_2;
	wire w_dff_B_lFKr3KxZ5_2;
	wire w_dff_B_mlzJ81VE7_2;
	wire w_dff_B_jJcPbM4i2_2;
	wire w_dff_B_LrcQsu8Z2_2;
	wire w_dff_B_0GbhOBaB3_2;
	wire w_dff_B_9zDx6fE76_2;
	wire w_dff_B_ZaHYn9Kk4_2;
	wire w_dff_B_9ggUCfBK7_2;
	wire w_dff_B_zoZRn6Nl4_2;
	wire w_dff_B_469OYTAY2_2;
	wire w_dff_B_5e8tB98s3_2;
	wire w_dff_B_dBNHdffZ6_2;
	wire w_dff_B_THr6khAD3_2;
	wire w_dff_B_ybIgZP7g0_2;
	wire w_dff_B_uT77OrPm8_2;
	wire w_dff_B_smPQwfaU6_2;
	wire w_dff_B_bZB3Cq7N1_2;
	wire w_dff_B_BWDsVCAw7_2;
	wire w_dff_B_b1bbbxGR2_2;
	wire w_dff_B_QnheOsAk7_2;
	wire w_dff_B_EwS4Zgpp6_2;
	wire w_dff_B_bJddEd148_2;
	wire w_dff_B_StFokFFU0_2;
	wire w_dff_B_iLfpviWR0_2;
	wire w_dff_B_t0a1Cb0x2_1;
	wire w_dff_B_gbLdcTBz1_2;
	wire w_dff_B_3yPBi7Xl0_2;
	wire w_dff_B_zPcgEp8b9_2;
	wire w_dff_B_OCdsBj5S9_2;
	wire w_dff_B_J1YdYyb88_2;
	wire w_dff_B_RrPFprv53_2;
	wire w_dff_B_TWY3H4s41_2;
	wire w_dff_B_8b7HdJju7_2;
	wire w_dff_B_5szc8Lyv9_2;
	wire w_dff_B_5prMed0M1_2;
	wire w_dff_B_mSexEWmK2_2;
	wire w_dff_B_Q4r0viye4_2;
	wire w_dff_B_J71A9wNR8_2;
	wire w_dff_B_RDohniPh7_2;
	wire w_dff_B_lfFljG9L5_2;
	wire w_dff_B_lNOsGHfN4_2;
	wire w_dff_B_qH7mVeSB1_2;
	wire w_dff_B_k7UpXjk40_2;
	wire w_dff_B_gxkE9eGk8_2;
	wire w_dff_B_kTFSDjs02_2;
	wire w_dff_B_KIFSxei32_2;
	wire w_dff_B_lS8iLh7H7_2;
	wire w_dff_B_PQp5RMD44_2;
	wire w_dff_B_0uNv9ZCo7_2;
	wire w_dff_B_b2HnPl0F6_2;
	wire w_dff_B_aIE8N9OT4_2;
	wire w_dff_B_dOjXQLHZ1_2;
	wire w_dff_B_lW6ZkaRh0_1;
	wire w_dff_B_G26W0DGU8_2;
	wire w_dff_B_HgZ7q5jk5_2;
	wire w_dff_B_a5yJQUzD8_2;
	wire w_dff_B_o2BMIsvw4_2;
	wire w_dff_B_K93xpsFb6_2;
	wire w_dff_B_mcofuDX07_2;
	wire w_dff_B_dxjETRKv3_2;
	wire w_dff_B_HTWBfWzI0_2;
	wire w_dff_B_g9fWyUSA1_2;
	wire w_dff_B_uA1SB5e10_2;
	wire w_dff_B_MQj0Ym9K7_2;
	wire w_dff_B_aSg1ez8S6_2;
	wire w_dff_B_DvOTFCWY4_2;
	wire w_dff_B_e4OMPagk2_2;
	wire w_dff_B_94PG2yZX9_2;
	wire w_dff_B_z25d29tI2_2;
	wire w_dff_B_kxh2SXZf6_2;
	wire w_dff_B_bbKUNQuY0_2;
	wire w_dff_B_Hofe42hk7_2;
	wire w_dff_B_32zujJz23_2;
	wire w_dff_B_14Iop9Gf0_2;
	wire w_dff_B_VOZWeydZ5_2;
	wire w_dff_B_f1YkdpU64_2;
	wire w_dff_B_LPIVmATe5_2;
	wire w_dff_B_sajY995T2_2;
	wire w_dff_B_Mq3GucuZ0_1;
	wire w_dff_B_FGkQiYP45_2;
	wire w_dff_B_jjTzbVSN0_2;
	wire w_dff_B_GXxEVzKw7_2;
	wire w_dff_B_AGYJOGDB8_2;
	wire w_dff_B_FuCZzOor0_2;
	wire w_dff_B_2X6svhfX3_2;
	wire w_dff_B_EWTXv7YF9_2;
	wire w_dff_B_POKoi7GG1_2;
	wire w_dff_B_pNkfxMLZ1_2;
	wire w_dff_B_soEM9Kco3_2;
	wire w_dff_B_GBbWMwcr4_2;
	wire w_dff_B_f3q3hBLW0_2;
	wire w_dff_B_TOgBGkuo6_2;
	wire w_dff_B_xOL9zfQv9_2;
	wire w_dff_B_MbdUYURa1_2;
	wire w_dff_B_rYVRGUli5_2;
	wire w_dff_B_855Ns1t19_2;
	wire w_dff_B_bRXgNsFt9_2;
	wire w_dff_B_UeGESLzn7_2;
	wire w_dff_B_hBlHuSKQ7_2;
	wire w_dff_B_3zLaC3ht5_2;
	wire w_dff_B_ajak31ho7_2;
	wire w_dff_B_Qjvy0QeU2_1;
	wire w_dff_B_mUoqfXpb6_2;
	wire w_dff_B_I5ekQYDB4_2;
	wire w_dff_B_Vxpr2bKG5_2;
	wire w_dff_B_AGojQlLr7_2;
	wire w_dff_B_6ZQeAD4R5_2;
	wire w_dff_B_svxZVkm66_2;
	wire w_dff_B_MXek9y2s8_2;
	wire w_dff_B_7iQWFiJG2_2;
	wire w_dff_B_xRUPNnY77_2;
	wire w_dff_B_RWVtGkIZ4_2;
	wire w_dff_B_xtJpvz2c0_2;
	wire w_dff_B_VO0qJIZt6_2;
	wire w_dff_B_kv3EngaH2_2;
	wire w_dff_B_47QfcKSa2_2;
	wire w_dff_B_Xp8eM6Dc5_2;
	wire w_dff_B_vyo7kTGM4_2;
	wire w_dff_B_3YLVvh6J3_2;
	wire w_dff_B_W4qd8b791_2;
	wire w_dff_B_6X1GQTtL4_2;
	wire w_dff_B_P3kYKh2x3_1;
	wire w_dff_B_n9PjZANv1_2;
	wire w_dff_B_BaxYGzmB6_2;
	wire w_dff_B_Cltch9Dv1_2;
	wire w_dff_B_J7td25uE2_2;
	wire w_dff_B_W2wE3Ibc1_2;
	wire w_dff_B_tS8MYGS40_2;
	wire w_dff_B_HrDbt5qB8_2;
	wire w_dff_B_ICxvdQxH0_2;
	wire w_dff_B_W3Sw7jZn6_2;
	wire w_dff_B_0GcYqEDU9_2;
	wire w_dff_B_3IuKSbMU0_2;
	wire w_dff_B_Dqd4RCCR4_2;
	wire w_dff_B_4dUU2XSZ9_2;
	wire w_dff_B_oeuxeKZW7_2;
	wire w_dff_B_oOUT4ZHk3_2;
	wire w_dff_B_BmViWpj58_2;
	wire w_dff_B_SIoX6JBv3_1;
	wire w_dff_B_dzEnWlGx0_2;
	wire w_dff_B_Ry4equLn1_2;
	wire w_dff_B_kt5DRlV32_2;
	wire w_dff_B_ZSQoWJbJ6_2;
	wire w_dff_B_mVklfNNI6_2;
	wire w_dff_B_XHI14um30_2;
	wire w_dff_B_qtgCMpEG1_2;
	wire w_dff_B_3Ul1QpQD9_2;
	wire w_dff_B_udoSRypK6_2;
	wire w_dff_B_ufUGcuMS3_2;
	wire w_dff_B_d18ygHiN3_2;
	wire w_dff_B_WSaq7kmt7_2;
	wire w_dff_B_HJJXPDLJ1_2;
	wire w_dff_B_EybfvUYZ7_1;
	wire w_dff_B_t2PhiEwp8_2;
	wire w_dff_B_HawM9VKV6_2;
	wire w_dff_B_AcRAbhG65_2;
	wire w_dff_B_2vL1UFbj1_2;
	wire w_dff_B_xB3fdIPI6_2;
	wire w_dff_B_ESApYGXA1_2;
	wire w_dff_B_nSWEkW2E6_2;
	wire w_dff_B_PgfyodEI6_2;
	wire w_dff_B_khvspGQO6_2;
	wire w_dff_B_9Ib3rFrG2_2;
	wire w_dff_B_z0LSDmXY5_2;
	wire w_dff_B_7ooSOI542_1;
	wire w_dff_B_p4ZKqOaR0_1;
	wire w_dff_B_35davhdi4_1;
	wire w_dff_B_JTDIvzWL1_1;
	wire w_dff_B_mhpKh3z56_1;
	wire w_dff_B_AbMIWrjY2_1;
	wire w_dff_B_lewCl6F46_0;
	wire w_dff_B_FN4EiElf2_0;
	wire w_dff_A_LtKs6naQ4_0;
	wire w_dff_A_QmNirHTN5_0;
	wire w_dff_A_PuqeexTg5_0;
	wire w_dff_B_y9utSxa10_1;
	wire w_dff_A_NXNylrvi2_0;
	wire w_dff_A_L65x3gO94_1;
	wire w_dff_A_M9IiwrW08_1;
	wire w_dff_A_EGLeKxBN2_1;
	wire w_dff_A_TJuwWHQb8_1;
	wire w_dff_A_1A2Pl0kz0_1;
	wire w_dff_A_pp2KJSQw2_1;
	wire w_dff_A_UVrgwKqi2_1;
	wire w_dff_A_pFIzj7hA7_1;
	wire w_dff_B_YhTOozlg0_1;
	wire w_dff_A_forErhb54_1;
	wire w_dff_B_M3dpZsFI7_1;
	wire w_dff_B_0HaB0axa1_2;
	wire w_dff_B_7k4QvExD2_2;
	wire w_dff_B_ff95Fdir3_2;
	wire w_dff_B_TfongzZn7_2;
	wire w_dff_B_wZEHvA7F2_2;
	wire w_dff_B_pXmYulmf2_2;
	wire w_dff_B_hyAbOmRm7_2;
	wire w_dff_B_NdWtZAad5_2;
	wire w_dff_B_2EvYEiLO7_2;
	wire w_dff_B_P6BeF5Ic8_2;
	wire w_dff_B_3iyorYZv3_2;
	wire w_dff_B_ohECjMdP8_2;
	wire w_dff_B_vsmlhH618_2;
	wire w_dff_B_mhVZrwmK5_2;
	wire w_dff_B_26FmZxsk4_2;
	wire w_dff_B_FITgjqxD6_2;
	wire w_dff_B_SCjdpMpj2_2;
	wire w_dff_B_saCfgQqm9_2;
	wire w_dff_B_z8m9NxYF4_2;
	wire w_dff_B_t7lFsx1r8_2;
	wire w_dff_B_WC7aDjPC7_2;
	wire w_dff_B_YDzMMs3k4_2;
	wire w_dff_B_snInNUvF6_2;
	wire w_dff_B_Eb2mfGpu2_2;
	wire w_dff_B_C67XFGMj4_2;
	wire w_dff_B_Et0VyXD14_2;
	wire w_dff_B_ghyagT206_2;
	wire w_dff_B_1TcmJCxp3_2;
	wire w_dff_B_2pibV6v52_2;
	wire w_dff_B_37YNWjfG8_2;
	wire w_dff_B_P72XedN77_2;
	wire w_dff_B_xIP8GnzF5_2;
	wire w_dff_B_U5rJyya81_2;
	wire w_dff_B_Cgri6rUs1_2;
	wire w_dff_B_V3iVCQRR9_2;
	wire w_dff_B_xWmgI4ER5_2;
	wire w_dff_B_PUcZxIoQ2_2;
	wire w_dff_B_KtU4aUNN1_2;
	wire w_dff_B_mZCFkYAs3_2;
	wire w_dff_B_YqQupxO30_2;
	wire w_dff_B_GgZharOd3_2;
	wire w_dff_B_Tl8NSNbd4_2;
	wire w_dff_B_8l0m3WpH6_2;
	wire w_dff_B_tSfQJftd3_2;
	wire w_dff_B_X4Yd2b2h3_2;
	wire w_dff_B_JKWxCRqU5_2;
	wire w_dff_B_weWzC20v2_2;
	wire w_dff_B_qpOnFZqU3_2;
	wire w_dff_B_zLPUFKln0_2;
	wire w_dff_B_frcMyTb66_2;
	wire w_dff_B_XZ7ZVWWB7_2;
	wire w_dff_B_8MOyUki03_2;
	wire w_dff_B_ZmKqx6aG2_2;
	wire w_dff_B_LyBfnB659_2;
	wire w_dff_B_DfFTOkR05_1;
	wire w_dff_B_YRZNjY0L5_2;
	wire w_dff_B_gGnvlyNI1_2;
	wire w_dff_B_9RO4XDfu8_2;
	wire w_dff_B_XYGfNuor9_2;
	wire w_dff_B_89Mem6RN5_2;
	wire w_dff_B_vi1Xy4W39_2;
	wire w_dff_B_YgBCan3K2_2;
	wire w_dff_B_9BusRFDI9_2;
	wire w_dff_B_0lHoUBJZ3_2;
	wire w_dff_B_JlD1X6Zy2_2;
	wire w_dff_B_MgqiZD7h9_2;
	wire w_dff_B_CIluDLVX6_2;
	wire w_dff_B_SFCQgHe50_2;
	wire w_dff_B_YJjqGf9e7_2;
	wire w_dff_B_k43PoL7w5_2;
	wire w_dff_B_3QikwAPS3_2;
	wire w_dff_B_Dxm82Scn5_2;
	wire w_dff_B_Tne9fqnL2_2;
	wire w_dff_B_rZctT1pP5_2;
	wire w_dff_B_40kpmGss3_2;
	wire w_dff_B_Uer9rEWK1_2;
	wire w_dff_B_765oAwsF8_2;
	wire w_dff_B_1R5ZorMF6_2;
	wire w_dff_B_qkNxMDal8_2;
	wire w_dff_B_HA4bT9nV5_2;
	wire w_dff_B_oiooNBCM8_2;
	wire w_dff_B_J8sTyzIM5_2;
	wire w_dff_B_KMKTM12T8_2;
	wire w_dff_B_zIA0RoIn2_2;
	wire w_dff_B_C1AJAiKq3_2;
	wire w_dff_B_5fr6FxiB9_2;
	wire w_dff_B_U0TSpj3E9_2;
	wire w_dff_B_n5lHouWi7_2;
	wire w_dff_B_p4jnIHe76_2;
	wire w_dff_B_1Jf62CBt7_2;
	wire w_dff_B_Bq6k7Bc37_2;
	wire w_dff_B_DiRQqmv01_2;
	wire w_dff_B_H2XFhAhq2_2;
	wire w_dff_B_hKB2wtra9_2;
	wire w_dff_B_mfFIpu5e7_2;
	wire w_dff_B_Sd5nOAgD9_2;
	wire w_dff_B_olUqor7E8_2;
	wire w_dff_B_ESaHf6bM1_2;
	wire w_dff_B_EXBnntxx7_2;
	wire w_dff_B_WcLJcDnf9_2;
	wire w_dff_B_sfl1UaQe2_2;
	wire w_dff_B_N6P56TQY2_2;
	wire w_dff_B_3c4LTtp89_2;
	wire w_dff_B_jlXX2w2d4_2;
	wire w_dff_B_4bnrSVb15_2;
	wire w_dff_B_th8nxmQb1_1;
	wire w_dff_B_spksI4KI0_2;
	wire w_dff_B_gHoaugaJ5_2;
	wire w_dff_B_viVHGa2t2_2;
	wire w_dff_B_UdS3I12J1_2;
	wire w_dff_B_AOLr9xT47_2;
	wire w_dff_B_9NBuqUrL2_2;
	wire w_dff_B_cnniJind8_2;
	wire w_dff_B_Plx1KvFc4_2;
	wire w_dff_B_yCEQ6V7U7_2;
	wire w_dff_B_aKePuP7k2_2;
	wire w_dff_B_MkIVpLcQ4_2;
	wire w_dff_B_kDx8BLnU9_2;
	wire w_dff_B_6UEBJIhl9_2;
	wire w_dff_B_UtZSgd8F0_2;
	wire w_dff_B_OQMvVDlt5_2;
	wire w_dff_B_8YfpEEqJ8_2;
	wire w_dff_B_ga1HpFPy4_2;
	wire w_dff_B_YsuQS3bt7_2;
	wire w_dff_B_Kgw5zafA2_2;
	wire w_dff_B_mxnlupeJ6_2;
	wire w_dff_B_XCeZ6X786_2;
	wire w_dff_B_U7h8D77U3_2;
	wire w_dff_B_zGSSVDbV3_2;
	wire w_dff_B_4dFxaZsZ6_2;
	wire w_dff_B_dW2WJBGK4_2;
	wire w_dff_B_eBkrm5Sx6_2;
	wire w_dff_B_IbEw2Xca7_2;
	wire w_dff_B_5MXoy1wm3_2;
	wire w_dff_B_UWiHhwvR6_2;
	wire w_dff_B_vN9s1hvP2_2;
	wire w_dff_B_Ah8tPILE5_2;
	wire w_dff_B_Sml7fttA9_2;
	wire w_dff_B_3n7fR1TM1_2;
	wire w_dff_B_tCttBEOm2_2;
	wire w_dff_B_7lD3d9d15_2;
	wire w_dff_B_UAbuuPvg5_2;
	wire w_dff_B_5ePkDAKo5_2;
	wire w_dff_B_7UIwb4sd0_2;
	wire w_dff_B_rZ6uSX1I1_2;
	wire w_dff_B_bI1QfeL17_2;
	wire w_dff_B_QfTPBrKg4_2;
	wire w_dff_B_lxgyNDby2_2;
	wire w_dff_B_u1V6BJSX0_2;
	wire w_dff_B_mldm1BE82_2;
	wire w_dff_B_Eg9FkntX4_2;
	wire w_dff_B_j8LajU4o8_2;
	wire w_dff_B_lFIuXwu42_1;
	wire w_dff_B_Qs3ojZcJ0_2;
	wire w_dff_B_uIbXlQDa0_2;
	wire w_dff_B_dcBuCuRl6_2;
	wire w_dff_B_gsMoO4Be2_2;
	wire w_dff_B_PN9urS541_2;
	wire w_dff_B_RXGdaVUM3_2;
	wire w_dff_B_hFY1IdO71_2;
	wire w_dff_B_RhxEi5HN8_2;
	wire w_dff_B_Ml4x5f5j1_2;
	wire w_dff_B_LV5TmCsu1_2;
	wire w_dff_B_Zn7zUcSl6_2;
	wire w_dff_B_Bw97XVjD4_2;
	wire w_dff_B_PNa2N3v14_2;
	wire w_dff_B_rPT91Zz68_2;
	wire w_dff_B_6ESbXcw15_2;
	wire w_dff_B_lM21z01S2_2;
	wire w_dff_B_6VHY6elh1_2;
	wire w_dff_B_5QK2eMPN4_2;
	wire w_dff_B_AkX6FeFy1_2;
	wire w_dff_B_OmAPtIcb8_2;
	wire w_dff_B_3mOYujGQ7_2;
	wire w_dff_B_0oO0W1rO1_2;
	wire w_dff_B_4804Unir7_2;
	wire w_dff_B_QWZeIdVw4_2;
	wire w_dff_B_Zb6eP5zx5_2;
	wire w_dff_B_Mbfv9tEX3_2;
	wire w_dff_B_y14YbYYC8_2;
	wire w_dff_B_MEB5eMOl8_2;
	wire w_dff_B_UyIA1UxH8_2;
	wire w_dff_B_RlgI2S1y2_2;
	wire w_dff_B_gL60ooUd5_2;
	wire w_dff_B_LYVrfjo41_2;
	wire w_dff_B_ZbhGg4gX2_2;
	wire w_dff_B_td786v915_2;
	wire w_dff_B_iMPfI7pk1_2;
	wire w_dff_B_ZQWJoX5c6_2;
	wire w_dff_B_VD1PKCFu3_2;
	wire w_dff_B_WSo1ZvR09_2;
	wire w_dff_B_B3u1pvnC9_2;
	wire w_dff_B_oB3QjWB10_2;
	wire w_dff_B_pLG9O1LA0_2;
	wire w_dff_B_sWdREgKP8_2;
	wire w_dff_B_xk3vPnoh0_1;
	wire w_dff_B_uxfWC7P78_2;
	wire w_dff_B_GJib9xOZ1_2;
	wire w_dff_B_3ez7Cg612_2;
	wire w_dff_B_LG7u3Kno1_2;
	wire w_dff_B_v3wBOw1y6_2;
	wire w_dff_B_6e14Ipz25_2;
	wire w_dff_B_tpddZU6i5_2;
	wire w_dff_B_3aX0VfXz2_2;
	wire w_dff_B_kXJGuqJH4_2;
	wire w_dff_B_gHmvmxyR7_2;
	wire w_dff_B_7JAUW5HU3_2;
	wire w_dff_B_nlt359wa6_2;
	wire w_dff_B_Vrl86BMW7_2;
	wire w_dff_B_NKtHwobk8_2;
	wire w_dff_B_bUSfSCpp7_2;
	wire w_dff_B_97LlHUBV3_2;
	wire w_dff_B_rcHDfZcH4_2;
	wire w_dff_B_8hUEyB7o2_2;
	wire w_dff_B_0GY5Vt3I3_2;
	wire w_dff_B_Zo7e0ClY7_2;
	wire w_dff_B_x4TZboyO8_2;
	wire w_dff_B_mEol29mC6_2;
	wire w_dff_B_sP7jbFzi9_2;
	wire w_dff_B_jdlrES7f4_2;
	wire w_dff_B_FVRPTocC9_2;
	wire w_dff_B_A7NlLIC69_2;
	wire w_dff_B_DlUjNFQq2_2;
	wire w_dff_B_uTBzcYKo6_2;
	wire w_dff_B_7GTTzrjg5_2;
	wire w_dff_B_Hm5u2qJ15_2;
	wire w_dff_B_RrjHD4372_2;
	wire w_dff_B_f7wSfMtQ4_2;
	wire w_dff_B_s6n4OxjG2_2;
	wire w_dff_B_AG23YI9i6_2;
	wire w_dff_B_HjmzoJX10_2;
	wire w_dff_B_0QPLeRFa5_2;
	wire w_dff_B_OncjjOTl6_2;
	wire w_dff_B_nlDQTvOA9_2;
	wire w_dff_B_h6vcaayM6_1;
	wire w_dff_B_LN1KLsKG0_2;
	wire w_dff_B_EKv3aaBO9_2;
	wire w_dff_B_ih1LFmet0_2;
	wire w_dff_B_TE6bvH520_2;
	wire w_dff_B_jbA2pDBE3_2;
	wire w_dff_B_6GS2D6WL2_2;
	wire w_dff_B_bahWkaCj8_2;
	wire w_dff_B_P4I6i2BR0_2;
	wire w_dff_B_wmB8RHgA4_2;
	wire w_dff_B_8MtvksDq9_2;
	wire w_dff_B_9rkhLf1N1_2;
	wire w_dff_B_20zguyvu0_2;
	wire w_dff_B_eem8j2Qn0_2;
	wire w_dff_B_ytUTXs197_2;
	wire w_dff_B_0KZ9AP1K8_2;
	wire w_dff_B_0vm24MMq6_2;
	wire w_dff_B_XkyvqK3f5_2;
	wire w_dff_B_1opj1cZ63_2;
	wire w_dff_B_hpXRjjSe9_2;
	wire w_dff_B_43zgnGut4_2;
	wire w_dff_B_A9Ks2ZsT2_2;
	wire w_dff_B_DsWwJvHK1_2;
	wire w_dff_B_uBt2GzZg2_2;
	wire w_dff_B_0fsiTw3x3_2;
	wire w_dff_B_jFZNP46H3_2;
	wire w_dff_B_SWmWQhEh6_2;
	wire w_dff_B_n6F17ieo9_2;
	wire w_dff_B_bwYKO1Fa7_2;
	wire w_dff_B_vVJPDswb5_2;
	wire w_dff_B_nCC9fcAH6_2;
	wire w_dff_B_Q9418DGX7_2;
	wire w_dff_B_zHfX8UyQ3_2;
	wire w_dff_B_1Wmbdlxi2_2;
	wire w_dff_B_JFgwEwTC7_2;
	wire w_dff_B_9L9nGFxd7_1;
	wire w_dff_B_fav47N7a8_2;
	wire w_dff_B_vUEzVpX84_2;
	wire w_dff_B_mSeKqQ5c7_2;
	wire w_dff_B_yGvZgSGm0_2;
	wire w_dff_B_tzXtrQJ47_2;
	wire w_dff_B_fsYCljgR8_2;
	wire w_dff_B_zOUDat0H1_2;
	wire w_dff_B_XOJTIFOE6_2;
	wire w_dff_B_7v3WGehJ8_2;
	wire w_dff_B_zwNYJRdG9_2;
	wire w_dff_B_zM3snEyE4_2;
	wire w_dff_B_lL1Lr7pY7_2;
	wire w_dff_B_5C1maZMv7_2;
	wire w_dff_B_Hv9BOByu3_2;
	wire w_dff_B_TXexaVhe4_2;
	wire w_dff_B_8CUlMfc80_2;
	wire w_dff_B_ouH1gUc92_2;
	wire w_dff_B_h9PFo6nE5_2;
	wire w_dff_B_xdJXjwU11_2;
	wire w_dff_B_LKbqQDaE5_2;
	wire w_dff_B_eoHwu7zi4_2;
	wire w_dff_B_ib0wdVZA5_2;
	wire w_dff_B_kHLkJIBB8_2;
	wire w_dff_B_nTmDnv9l4_2;
	wire w_dff_B_rjZuGj266_2;
	wire w_dff_B_LE2cHTDX0_2;
	wire w_dff_B_R7eja0Cs2_2;
	wire w_dff_B_4NG8Ychw2_2;
	wire w_dff_B_1Nd5QAbS8_2;
	wire w_dff_B_hg36VsNB6_2;
	wire w_dff_B_oNsStTFp5_1;
	wire w_dff_B_oHmv5qXR6_2;
	wire w_dff_B_NZgkpkxH2_2;
	wire w_dff_B_rDQfFCGb5_2;
	wire w_dff_B_aCA50iKr5_2;
	wire w_dff_B_6k1sIwv72_2;
	wire w_dff_B_F22AP4UG6_2;
	wire w_dff_B_B0ucpamH0_2;
	wire w_dff_B_ZpIMM9nD3_2;
	wire w_dff_B_nrmH1mBP0_2;
	wire w_dff_B_yxFTUBzI4_2;
	wire w_dff_B_p6vil0Wl2_2;
	wire w_dff_B_cHaKcw4M2_2;
	wire w_dff_B_aogjyaBg9_2;
	wire w_dff_B_wtCTFTy29_2;
	wire w_dff_B_0i6o4roQ2_2;
	wire w_dff_B_DFu1ENa23_2;
	wire w_dff_B_kjPesmOp9_2;
	wire w_dff_B_Ytcb8UoX6_2;
	wire w_dff_B_OfeB5gDa3_2;
	wire w_dff_B_GLibKxEC7_2;
	wire w_dff_B_gYCGV48K5_2;
	wire w_dff_B_Ak3YZDbs5_2;
	wire w_dff_B_oMftZqqS6_2;
	wire w_dff_B_2PNucZHP1_2;
	wire w_dff_B_Dq6CTl2L9_2;
	wire w_dff_B_IYIt1woL4_2;
	wire w_dff_B_GJ7x2nk19_1;
	wire w_dff_B_YrNXONms6_2;
	wire w_dff_B_5ZG9u9ZI9_2;
	wire w_dff_B_1Ze3lasn0_2;
	wire w_dff_B_zSvF6KbM8_2;
	wire w_dff_B_YXlU9lrF2_2;
	wire w_dff_B_EPTjINBL6_2;
	wire w_dff_B_qaMRMaTs9_2;
	wire w_dff_B_OgC9dRfe4_2;
	wire w_dff_B_OcOJGZyC7_2;
	wire w_dff_B_BxtNQLdp8_2;
	wire w_dff_B_qgFBy6918_2;
	wire w_dff_B_n5GFp7w90_2;
	wire w_dff_B_8MBLqyIJ4_2;
	wire w_dff_B_HDEZdqV55_2;
	wire w_dff_B_SDJSmfqO0_2;
	wire w_dff_B_LXZwxnQa9_2;
	wire w_dff_B_3Q1D1rBf2_2;
	wire w_dff_B_pVFPtswd1_2;
	wire w_dff_B_w0kiJNFI2_2;
	wire w_dff_B_uVhiqHwO3_2;
	wire w_dff_B_sEnDKUqv7_2;
	wire w_dff_B_3ek4XcaU4_1;
	wire w_dff_B_lJ7C1RDt4_2;
	wire w_dff_B_FO3yi2lv8_2;
	wire w_dff_B_GUmy7p0p6_2;
	wire w_dff_B_DyutjSWN5_2;
	wire w_dff_B_MXBeQyFu9_2;
	wire w_dff_B_3A2UMLPS5_2;
	wire w_dff_B_EbZpbqqa4_2;
	wire w_dff_B_rL8qINCn0_2;
	wire w_dff_B_cvGRX6as8_2;
	wire w_dff_B_kUGaiZG37_2;
	wire w_dff_B_6eYryBY42_2;
	wire w_dff_B_0z6X96Rf4_2;
	wire w_dff_B_dpRxWuvB5_2;
	wire w_dff_B_CyniIOTJ5_2;
	wire w_dff_B_RyO1k4AJ4_2;
	wire w_dff_B_Nsh1AuaP6_2;
	wire w_dff_B_n59VXHVa0_2;
	wire w_dff_B_65EnfEbg5_2;
	wire w_dff_B_OSqXrNmC5_2;
	wire w_dff_B_AINmtyNJ6_1;
	wire w_dff_B_iK2mAFDW3_2;
	wire w_dff_B_PCD0TPj07_2;
	wire w_dff_B_b6276lxL4_2;
	wire w_dff_B_wTwB5vvR5_2;
	wire w_dff_B_eqJobM641_2;
	wire w_dff_B_V5uOjYkI2_2;
	wire w_dff_B_FWrQbHA09_2;
	wire w_dff_B_QpfJ0azY9_2;
	wire w_dff_B_2kAvn4pW1_2;
	wire w_dff_B_siEFPnIM9_2;
	wire w_dff_B_IwFsrmHY7_2;
	wire w_dff_B_4ZJQmA1u2_2;
	wire w_dff_B_Jyg6YH0c9_2;
	wire w_dff_B_2MCgcwcC5_2;
	wire w_dff_B_ZfiCaKEH3_2;
	wire w_dff_B_hQnr7CKb1_2;
	wire w_dff_B_tsN5TVO52_2;
	wire w_dff_B_9lRe7hy55_1;
	wire w_dff_B_1lJKtMc85_2;
	wire w_dff_B_jppu77Gt1_2;
	wire w_dff_B_LSv5OsKr9_2;
	wire w_dff_B_UFnpmM8a5_2;
	wire w_dff_B_mmUVITa76_2;
	wire w_dff_B_WAzqaay31_2;
	wire w_dff_B_3BPAC2gE2_2;
	wire w_dff_B_OPDbgvjk9_2;
	wire w_dff_B_gRQjQGh94_2;
	wire w_dff_B_pcqWMDNl5_2;
	wire w_dff_B_nFu9CEJG0_2;
	wire w_dff_B_23rRmjYY1_2;
	wire w_dff_B_FiJjNlFe1_2;
	wire w_dff_B_ok5zClye5_2;
	wire w_dff_B_aSMKxdg69_1;
	wire w_dff_B_mjik72bq7_2;
	wire w_dff_B_RY9mRFZd0_2;
	wire w_dff_B_xSHMoOkf1_2;
	wire w_dff_B_K0Lx7DLD7_2;
	wire w_dff_B_AeZXW2289_2;
	wire w_dff_B_QaVHFWPL4_2;
	wire w_dff_B_zaEV6AUQ7_2;
	wire w_dff_B_OSsHow5H5_2;
	wire w_dff_B_3FIpdvcG0_2;
	wire w_dff_B_tcFqXBI95_2;
	wire w_dff_B_43zDDGAx6_2;
	wire w_dff_B_CF3fq3pc5_2;
	wire w_dff_B_YfhrVjh72_1;
	wire w_dff_B_6849uQSw6_1;
	wire w_dff_B_wWYbSLJf7_1;
	wire w_dff_B_FFR5M8UT0_1;
	wire w_dff_B_xmythnXI6_1;
	wire w_dff_B_ewdCX36A1_1;
	wire w_dff_B_8judfUTY8_0;
	wire w_dff_B_d7N1ZYqq2_0;
	wire w_dff_A_l2pq6lHB9_0;
	wire w_dff_A_7YwHJFsi2_0;
	wire w_dff_A_CxS8Eef66_0;
	wire w_dff_B_zrpbKDpH7_1;
	wire w_dff_A_T2OwA3n83_0;
	wire w_dff_A_NGDQpmyY8_1;
	wire w_dff_A_45MFTm1j1_1;
	wire w_dff_A_d2Qncvh02_1;
	wire w_dff_A_U5mbdxMM8_1;
	wire w_dff_A_4LbXaeqt2_1;
	wire w_dff_A_fFWhP3vZ1_1;
	wire w_dff_A_evkcmivS0_1;
	wire w_dff_A_kO1gTAnV0_1;
	wire w_dff_B_jCAK1uKJ6_1;
	wire w_dff_B_m74SQWxQ6_1;
	wire w_dff_B_SykyZ5wE9_1;
	wire w_dff_B_CUxnaWaM1_2;
	wire w_dff_B_b28AAknA0_2;
	wire w_dff_B_2F6PUUyV0_2;
	wire w_dff_B_skppOEvw0_2;
	wire w_dff_B_qCm9mVjM7_2;
	wire w_dff_B_3XdIOSMc7_2;
	wire w_dff_B_BK5kXT6W0_2;
	wire w_dff_B_9FxtHGkt3_2;
	wire w_dff_B_YrICbcdI5_2;
	wire w_dff_B_8qfAlAIl3_2;
	wire w_dff_B_NVIIEGVa5_2;
	wire w_dff_B_iSr6Q6Ml7_2;
	wire w_dff_B_iSNbBS7X0_2;
	wire w_dff_B_iXZyuVYv1_2;
	wire w_dff_B_3v1zFld53_2;
	wire w_dff_B_t6yA3jm96_2;
	wire w_dff_B_eDKF1vgK6_2;
	wire w_dff_B_g0hTqjNL0_2;
	wire w_dff_B_KkZANGyg3_2;
	wire w_dff_B_S4c2Pgr29_2;
	wire w_dff_B_4NnsSIQ28_2;
	wire w_dff_B_YsQ2ps2v5_2;
	wire w_dff_B_OuqYkvnT0_2;
	wire w_dff_B_Tcb3BKtD3_2;
	wire w_dff_B_pqwEOZ3h2_2;
	wire w_dff_B_HOgzSMcM2_2;
	wire w_dff_B_FQ59q70x2_2;
	wire w_dff_B_yvBEuBC50_2;
	wire w_dff_B_oWrJkv4c0_2;
	wire w_dff_B_O1VL38gO8_2;
	wire w_dff_B_0b5JWE0C3_2;
	wire w_dff_B_JIkDY88H5_2;
	wire w_dff_B_PgwT66Ft0_2;
	wire w_dff_B_x1E0QGhx9_2;
	wire w_dff_B_ca5zKw4h8_2;
	wire w_dff_B_uzznCBdC5_2;
	wire w_dff_B_pBLwVpBR3_2;
	wire w_dff_B_2vBVMB5V7_2;
	wire w_dff_B_PAPhILIy3_2;
	wire w_dff_B_WRwiQj2L4_2;
	wire w_dff_B_EHldMUyZ4_2;
	wire w_dff_B_6pIPIOnR0_2;
	wire w_dff_B_xGLIlCo35_2;
	wire w_dff_B_6SDlchVF5_2;
	wire w_dff_B_QVJawq5M1_2;
	wire w_dff_B_33JjJkgE1_2;
	wire w_dff_B_xYrxdJeJ8_2;
	wire w_dff_B_zlYVAhuQ2_2;
	wire w_dff_B_UdVcBu1Y2_2;
	wire w_dff_B_GSay1yMy4_2;
	wire w_dff_B_uJDcT60q3_2;
	wire w_dff_B_Vl3RO6UD6_2;
	wire w_dff_B_ic6kJmWQ0_2;
	wire w_dff_B_o3w5aTvI6_2;
	wire w_dff_B_tS3OpCkK8_2;
	wire w_dff_B_JpaPDBvt5_2;
	wire w_dff_B_Io0C18lm3_2;
	wire w_dff_B_0JpSH0Ks5_2;
	wire w_dff_B_JcwB5xj55_2;
	wire w_dff_B_3XafXdoa3_2;
	wire w_dff_B_6eWBLgkO9_2;
	wire w_dff_B_zwOG9EMm1_2;
	wire w_dff_B_fAMpavzh5_2;
	wire w_dff_B_43CkqX3Q6_2;
	wire w_dff_B_Oajl5QBZ0_2;
	wire w_dff_B_XbSfiRoT2_2;
	wire w_dff_B_2JzFZOws9_2;
	wire w_dff_B_JUogRO798_2;
	wire w_dff_B_6BTKIP6a1_2;
	wire w_dff_B_9QV78O5O7_2;
	wire w_dff_B_UbrfE7eD8_2;
	wire w_dff_B_PxKKlXrO1_2;
	wire w_dff_B_OBCWGu427_2;
	wire w_dff_B_Ftt84J4K6_2;
	wire w_dff_B_kXcQg8lf6_2;
	wire w_dff_B_g5fyCOod0_2;
	wire w_dff_B_WAIpNcRT3_2;
	wire w_dff_B_yGZJ0dbg3_2;
	wire w_dff_B_5aPNFg957_2;
	wire w_dff_B_UWkzjN9W7_2;
	wire w_dff_B_P8ozYtQT3_2;
	wire w_dff_B_EGpFVIuC6_2;
	wire w_dff_B_8sVdXMeF4_2;
	wire w_dff_B_mLXGekro9_2;
	wire w_dff_B_e0aBAl9o2_2;
	wire w_dff_B_xbANQquN3_2;
	wire w_dff_B_YwtbcyEk0_2;
	wire w_dff_B_ezY8Qn7m3_2;
	wire w_dff_B_4hHymzK85_2;
	wire w_dff_B_0FiXl07T4_2;
	wire w_dff_B_gRthv1q88_2;
	wire w_dff_B_zw7zxnwg9_2;
	wire w_dff_B_jxC1T4AV6_2;
	wire w_dff_B_E2dozOxm0_2;
	wire w_dff_B_BSDbIl0Z8_2;
	wire w_dff_B_i3i2BuvJ5_2;
	wire w_dff_B_lqrZSR975_2;
	wire w_dff_B_LDhrNUaG9_2;
	wire w_dff_B_vblGXDUh3_2;
	wire w_dff_B_Vh7J7k9B3_2;
	wire w_dff_B_uGbOiL3U2_2;
	wire w_dff_B_nTSBBC977_2;
	wire w_dff_B_DxOxGhbg6_2;
	wire w_dff_B_A9ejUpU21_2;
	wire w_dff_B_w5EglXWf4_2;
	wire w_dff_B_yx5ZLr0Q9_2;
	wire w_dff_B_S3CfbWQj4_2;
	wire w_dff_B_3NNnZg2w2_2;
	wire w_dff_B_p8UVPiSB4_2;
	wire w_dff_B_eEHRC27B2_2;
	wire w_dff_B_mcyc9t8e2_2;
	wire w_dff_B_HAS1H0Vi8_2;
	wire w_dff_B_xBEtQaQ09_2;
	wire w_dff_B_LrVQ6VMx0_2;
	wire w_dff_A_PxkUvdjD5_1;
	wire w_dff_B_tNkfSlSJ7_1;
	wire w_dff_B_4dLvkYWc8_2;
	wire w_dff_B_sLQsfsQl0_2;
	wire w_dff_B_oTplcCrl8_2;
	wire w_dff_B_a6odMmZx5_2;
	wire w_dff_B_YUE9JYIw7_2;
	wire w_dff_B_scrNy5P06_2;
	wire w_dff_B_I1FQNfmj5_2;
	wire w_dff_B_VmxyKjzi0_2;
	wire w_dff_B_fsLTpXFY3_2;
	wire w_dff_B_7ZwsPFYy8_2;
	wire w_dff_B_qOoOHsiR9_2;
	wire w_dff_B_BbupKVlH9_2;
	wire w_dff_B_P1Ih1j6K5_2;
	wire w_dff_B_DgXScoMA0_2;
	wire w_dff_B_NmBS3vZW2_2;
	wire w_dff_B_Q77MKcYK8_2;
	wire w_dff_B_WuHLpyfd9_2;
	wire w_dff_B_lo6BSgHR0_2;
	wire w_dff_B_HqPjGSw55_2;
	wire w_dff_B_IYTCDilo3_2;
	wire w_dff_B_LJCdHRll0_2;
	wire w_dff_B_fZnb51im9_2;
	wire w_dff_B_cs7d5pUm3_2;
	wire w_dff_B_kNTNVw497_2;
	wire w_dff_B_uVOH9iV53_2;
	wire w_dff_B_pd8cr83u1_2;
	wire w_dff_B_x0ZdlwOg4_2;
	wire w_dff_B_dxU6Rwjq1_2;
	wire w_dff_B_0HHP96Ct3_2;
	wire w_dff_B_FnpccuzM3_2;
	wire w_dff_B_JYGUfNFJ6_2;
	wire w_dff_B_KQVbYU6k0_2;
	wire w_dff_B_0avmNBE58_2;
	wire w_dff_B_tQU9bh5X8_2;
	wire w_dff_B_td7Gawrf0_2;
	wire w_dff_B_BifjfJIz2_2;
	wire w_dff_B_LNtVcsYs7_2;
	wire w_dff_B_JATmf3Qr5_2;
	wire w_dff_B_909Y0NrD1_2;
	wire w_dff_B_DCHDFsZj8_2;
	wire w_dff_B_0XEov4yd9_2;
	wire w_dff_B_A0hF8aBU9_2;
	wire w_dff_B_ksdZnOE90_2;
	wire w_dff_B_47ZBgnGh9_2;
	wire w_dff_B_Orxy2JUP1_2;
	wire w_dff_B_tJgmbYCk6_2;
	wire w_dff_B_dHAPEObs9_2;
	wire w_dff_B_FQuRCi891_2;
	wire w_dff_B_Y3F4Ii1O1_2;
	wire w_dff_B_t2O9zU334_2;
	wire w_dff_B_IfzgHusX8_2;
	wire w_dff_B_GOI5AjxA5_2;
	wire w_dff_B_BqzcS7iz9_2;
	wire w_dff_B_B12W2YLo8_2;
	wire w_dff_B_BDl4KhBR6_2;
	wire w_dff_B_sZ0n4Hta5_1;
	wire w_dff_B_4SA924Xj6_1;
	wire w_dff_B_pYtGxsg74_2;
	wire w_dff_B_6wcyaKks7_2;
	wire w_dff_B_tYVFheJu1_2;
	wire w_dff_B_ZXdJCphm5_2;
	wire w_dff_B_SgtXfrKJ1_2;
	wire w_dff_B_JUgGGi8m3_2;
	wire w_dff_B_BWMXU5Od6_2;
	wire w_dff_B_gXZI6gMM4_2;
	wire w_dff_B_sqKFri9O2_2;
	wire w_dff_B_KHD8PpI99_2;
	wire w_dff_B_D5HvEX1H6_2;
	wire w_dff_B_1MsBVYxW1_2;
	wire w_dff_B_HP6jWg9P9_2;
	wire w_dff_B_OgEhbXF22_2;
	wire w_dff_B_HGZZxS0u1_2;
	wire w_dff_B_skp5RAy89_2;
	wire w_dff_B_AKnNt36s7_2;
	wire w_dff_B_0TDGUQG90_2;
	wire w_dff_B_FCnxYKVA8_2;
	wire w_dff_B_1o47LyxD5_2;
	wire w_dff_B_KbJkTd8h5_2;
	wire w_dff_B_gkWCoAB23_2;
	wire w_dff_B_UQmXc7to0_2;
	wire w_dff_B_4UTup3KZ6_2;
	wire w_dff_B_LhTZJTzn6_2;
	wire w_dff_B_4cS2J8M68_2;
	wire w_dff_B_M6rGNXHB9_2;
	wire w_dff_B_MGhtXBaN5_2;
	wire w_dff_B_68U2CJkr2_2;
	wire w_dff_B_ufurvf7s9_2;
	wire w_dff_B_XZPkNmnU2_2;
	wire w_dff_B_VCQI0V6X0_2;
	wire w_dff_B_ZKBNlK0a0_2;
	wire w_dff_B_UYT9ceN93_2;
	wire w_dff_B_FMCpWyC84_2;
	wire w_dff_B_5Z13YJdr9_2;
	wire w_dff_B_S1UFURAg6_2;
	wire w_dff_B_pVaxPmDY7_2;
	wire w_dff_B_ezxlfzdC5_2;
	wire w_dff_B_Rm2GF1Gd0_2;
	wire w_dff_B_q2uh49Nx8_2;
	wire w_dff_B_e6DDI9pT2_2;
	wire w_dff_B_90gFSyaO2_2;
	wire w_dff_B_L8DhqAQa1_2;
	wire w_dff_B_0THf7X6Y9_2;
	wire w_dff_B_CFuopNKt8_2;
	wire w_dff_B_eRw48RmR9_2;
	wire w_dff_B_gY0Fu8SE1_2;
	wire w_dff_B_dcPATMxg5_2;
	wire w_dff_B_daCfm07m0_2;
	wire w_dff_B_rgODx5oW3_2;
	wire w_dff_B_liKzinUN3_2;
	wire w_dff_B_BsaTgHYw4_2;
	wire w_dff_B_t1O6oKSq9_2;
	wire w_dff_B_ffSl9Cab9_2;
	wire w_dff_B_rGwecK6y3_2;
	wire w_dff_B_iePs9Un07_2;
	wire w_dff_B_P7LeVSks1_2;
	wire w_dff_B_X9bENC9z3_2;
	wire w_dff_B_Kpkcmpxd9_2;
	wire w_dff_B_f7Ms2toJ7_2;
	wire w_dff_B_9UUunrXK7_2;
	wire w_dff_B_1D2L7WHF8_2;
	wire w_dff_B_xflbiNQm5_2;
	wire w_dff_B_O8R6TIUu0_2;
	wire w_dff_B_YyY3S8tN5_2;
	wire w_dff_B_tac62QeS5_2;
	wire w_dff_B_1ZNPkkAa9_2;
	wire w_dff_B_mvwwcEob5_2;
	wire w_dff_B_XsPAtI5j4_2;
	wire w_dff_B_ym3FaRK93_2;
	wire w_dff_B_9VbxueTl5_2;
	wire w_dff_B_nxuuSiIL1_2;
	wire w_dff_B_FaGLtmmB8_2;
	wire w_dff_B_ziSHAdvN8_2;
	wire w_dff_B_bvhQ0Iwp7_2;
	wire w_dff_B_uSY1jnWt4_2;
	wire w_dff_B_VHF6EVyl6_2;
	wire w_dff_B_npCI8OJT0_2;
	wire w_dff_B_ag9mSPOG2_2;
	wire w_dff_B_IrtbiRLW6_2;
	wire w_dff_B_ddDhfMnS6_2;
	wire w_dff_B_J5JQUBGL5_2;
	wire w_dff_B_502FbmUk1_2;
	wire w_dff_B_x3i6euFo9_2;
	wire w_dff_B_7LY5gOsh0_2;
	wire w_dff_B_pfohpeQA2_2;
	wire w_dff_B_S3xA4Bdw5_2;
	wire w_dff_B_hanA9ou25_2;
	wire w_dff_B_zTIxwpjW0_2;
	wire w_dff_B_rQbUJ0ru3_2;
	wire w_dff_B_fwqoqcxC6_2;
	wire w_dff_B_2EmyCWth1_2;
	wire w_dff_B_ioHhMvB60_2;
	wire w_dff_B_qUrc4GBi7_2;
	wire w_dff_B_ktSeaH7l9_2;
	wire w_dff_B_hQUK7uvr6_2;
	wire w_dff_B_OU9X3bAu4_2;
	wire w_dff_B_HMeGfbQN8_2;
	wire w_dff_B_Cjs9p1UA5_2;
	wire w_dff_B_ZXGHL8ZM3_2;
	wire w_dff_B_zlajOHoB8_2;
	wire w_dff_B_ikPHQRGp4_2;
	wire w_dff_B_6EMyCyQB3_2;
	wire w_dff_B_MKqAvzv91_2;
	wire w_dff_B_cMF3AuPD1_2;
	wire w_dff_B_MHVvfctY5_2;
	wire w_dff_B_F4FHKNsW0_1;
	wire w_dff_B_7th5Eu8k8_2;
	wire w_dff_B_eNtQf8L76_2;
	wire w_dff_B_ezqvSYVZ6_2;
	wire w_dff_B_9fcBDFs02_2;
	wire w_dff_B_qsmmEwuc5_2;
	wire w_dff_B_tfyTaVAS2_2;
	wire w_dff_B_zOb538h45_2;
	wire w_dff_B_RJjmI3QK1_2;
	wire w_dff_B_EYDSJ1sE8_2;
	wire w_dff_B_DO0oLwq75_2;
	wire w_dff_B_CuyjJIYD9_2;
	wire w_dff_B_6ozzNfPh4_2;
	wire w_dff_B_7YzEt90d8_2;
	wire w_dff_B_Dxn49qfq0_2;
	wire w_dff_B_5GdsDPw96_2;
	wire w_dff_B_22QqtQ808_2;
	wire w_dff_B_RqYL07YI1_2;
	wire w_dff_B_aNcYWcOO0_2;
	wire w_dff_B_MXDMfUh82_2;
	wire w_dff_B_dj062R2L6_2;
	wire w_dff_B_FMniWWpY4_2;
	wire w_dff_B_gwBjsHvd8_2;
	wire w_dff_B_8Js46k7n8_2;
	wire w_dff_B_GxZMVNUd0_2;
	wire w_dff_B_Y1jUCgmY4_2;
	wire w_dff_B_VHOplYd21_2;
	wire w_dff_B_sqHp7r664_2;
	wire w_dff_B_FJfdvBIf9_2;
	wire w_dff_B_DoIa5PwG1_2;
	wire w_dff_B_zN4Rv6WV8_2;
	wire w_dff_B_CuONGkfX1_2;
	wire w_dff_B_cPwlPMfn0_2;
	wire w_dff_B_cDJhrIkx9_2;
	wire w_dff_B_Iw2lApEp2_2;
	wire w_dff_B_Jz6mZXIg2_2;
	wire w_dff_B_dXfV98yg9_2;
	wire w_dff_B_9KmcZ8cl8_2;
	wire w_dff_B_zbFxFGgO2_2;
	wire w_dff_B_vO8nQTRu6_2;
	wire w_dff_B_hsKuwM0e2_2;
	wire w_dff_B_O796C1Mu8_2;
	wire w_dff_B_UClX28LH5_2;
	wire w_dff_B_nldJQdoc6_2;
	wire w_dff_B_6XfxOawj1_2;
	wire w_dff_B_BtpAo8wy3_2;
	wire w_dff_B_8tKzbF3I9_2;
	wire w_dff_B_3KXoA0oy1_2;
	wire w_dff_B_6wMB7NcD8_2;
	wire w_dff_B_jmGBCNw90_2;
	wire w_dff_B_PSwzMt0B0_2;
	wire w_dff_B_D4NOgbEQ5_2;
	wire w_dff_B_oYaDfUxp0_1;
	wire w_dff_B_Zw6pdW2B7_1;
	wire w_dff_B_OV4LUR9w6_2;
	wire w_dff_B_7xVEc9Hf6_2;
	wire w_dff_B_9zawBzxn9_2;
	wire w_dff_B_MieYUYhc0_2;
	wire w_dff_B_z5ZvKtdP1_2;
	wire w_dff_B_B1iToAsH0_2;
	wire w_dff_B_5gUBTiEV8_2;
	wire w_dff_B_OuEIFy7O2_2;
	wire w_dff_B_Zm7Vb1ab6_2;
	wire w_dff_B_GOhfNCV89_2;
	wire w_dff_B_IRBZdozG4_2;
	wire w_dff_B_yN02whnS4_2;
	wire w_dff_B_RHotYsHB3_2;
	wire w_dff_B_aiTtJlBd0_2;
	wire w_dff_B_30NKNu9z1_2;
	wire w_dff_B_J9XBmAWz3_2;
	wire w_dff_B_KRdQabDh0_2;
	wire w_dff_B_8xt4TcaS7_2;
	wire w_dff_B_DdQebRkn8_2;
	wire w_dff_B_5ndfVFLi2_2;
	wire w_dff_B_EJRUeUsm9_2;
	wire w_dff_B_Rsr9SgWK7_2;
	wire w_dff_B_UgIiy5Kt6_2;
	wire w_dff_B_CU6wx5aF5_2;
	wire w_dff_B_bCX4Ajy76_2;
	wire w_dff_B_TMm5lXh39_2;
	wire w_dff_B_hrHhPy0U8_2;
	wire w_dff_B_VlUjF8JE3_2;
	wire w_dff_B_PG7edLz47_2;
	wire w_dff_B_YeZoBVpI3_2;
	wire w_dff_B_2vuAxxcz5_2;
	wire w_dff_B_Zo7pIShD4_2;
	wire w_dff_B_YM1UwXZe3_2;
	wire w_dff_B_XHW13VCe7_2;
	wire w_dff_B_O3ViLOwi6_2;
	wire w_dff_B_ZJrLVXEH9_2;
	wire w_dff_B_dwrjPAOO5_2;
	wire w_dff_B_KcxmlSch9_2;
	wire w_dff_B_PnhtiqsM1_2;
	wire w_dff_B_AXtIdQhT6_2;
	wire w_dff_B_xWAgze7w9_2;
	wire w_dff_B_ZJAz3KHS8_2;
	wire w_dff_B_e0XZZnYI7_2;
	wire w_dff_B_zLltfwQ73_2;
	wire w_dff_B_BqDVFM0I9_2;
	wire w_dff_B_YB20j6aj7_2;
	wire w_dff_B_pAwqq2H84_2;
	wire w_dff_B_Pk8E9oz23_2;
	wire w_dff_B_JbmMvYa28_2;
	wire w_dff_B_HLYmbXXu4_2;
	wire w_dff_B_Bbe2et671_2;
	wire w_dff_B_MP2LU5qv2_2;
	wire w_dff_B_bPL2csOe3_2;
	wire w_dff_B_KvEjsbWD6_2;
	wire w_dff_B_YUhrlVBC6_2;
	wire w_dff_B_jOefrOrM7_2;
	wire w_dff_B_9d3OhIBC0_2;
	wire w_dff_B_eKpd4oYH6_2;
	wire w_dff_B_080ijP9M4_2;
	wire w_dff_B_yCaNAeC87_2;
	wire w_dff_B_bKPjXg5E8_2;
	wire w_dff_B_F7Cnun5r4_2;
	wire w_dff_B_yKzMgUDd6_2;
	wire w_dff_B_fkr5epSt1_2;
	wire w_dff_B_pEXQ0zAK8_2;
	wire w_dff_B_DdwJof3h4_2;
	wire w_dff_B_Ry7Emped2_2;
	wire w_dff_B_ZvyBeOMc0_2;
	wire w_dff_B_er71KSAg2_2;
	wire w_dff_B_TU1ZtA7S9_2;
	wire w_dff_B_TTQ0rCYZ5_2;
	wire w_dff_B_eq8TzAIK3_2;
	wire w_dff_B_wg6UR4za2_2;
	wire w_dff_B_ovCrJYmZ1_2;
	wire w_dff_B_uXlVHjDb6_2;
	wire w_dff_B_A8I7fDO20_2;
	wire w_dff_B_iNxsZu442_2;
	wire w_dff_B_U8TTNHZv1_2;
	wire w_dff_B_JjzevDjA3_2;
	wire w_dff_B_LdtPjObD7_2;
	wire w_dff_B_aNEvkxOt6_2;
	wire w_dff_B_cGjC7Z618_2;
	wire w_dff_B_05Ha8Hq07_2;
	wire w_dff_B_JBoKDsAG6_2;
	wire w_dff_B_5LjpxmwP3_2;
	wire w_dff_B_TeoLBedL4_2;
	wire w_dff_B_owtTLooF9_2;
	wire w_dff_B_m1RR29ev5_2;
	wire w_dff_B_21nNhFmo1_2;
	wire w_dff_B_VCGXyKEd7_2;
	wire w_dff_B_kljDPrGO5_2;
	wire w_dff_B_Ug5oEP0f3_2;
	wire w_dff_B_RESDTSlx4_2;
	wire w_dff_B_I8mhd0fK9_2;
	wire w_dff_B_IXvPLQhX8_2;
	wire w_dff_B_KvOeL6FU1_2;
	wire w_dff_B_BG45Licz8_2;
	wire w_dff_B_BBmT6JTF2_2;
	wire w_dff_B_nodTVjh30_2;
	wire w_dff_B_L2SDGRk72_1;
	wire w_dff_B_ZWkI9xn98_2;
	wire w_dff_B_RvkAJ08B5_2;
	wire w_dff_B_VeZ4sR612_2;
	wire w_dff_B_T4b7XMC90_2;
	wire w_dff_B_ZTQaUEub6_2;
	wire w_dff_B_0ujpAZ0z9_2;
	wire w_dff_B_SL921Pt80_2;
	wire w_dff_B_Bg7uuIgI8_2;
	wire w_dff_B_Iv1CUzmx8_2;
	wire w_dff_B_yPcKFBWT3_2;
	wire w_dff_B_kUBVjpyw2_2;
	wire w_dff_B_c5rXOnPh5_2;
	wire w_dff_B_y2X4KWtG6_2;
	wire w_dff_B_qap6YxH67_2;
	wire w_dff_B_dkeqJFbi4_2;
	wire w_dff_B_iCjWJ5809_2;
	wire w_dff_B_0ahnppPY8_2;
	wire w_dff_B_mhG9EiKt7_2;
	wire w_dff_B_ourMqqw07_2;
	wire w_dff_B_1jzBeIjY9_2;
	wire w_dff_B_BuZnoyKm4_2;
	wire w_dff_B_xR8vUvqk4_2;
	wire w_dff_B_ZxSQhSYP7_2;
	wire w_dff_B_0b1WvJfR3_2;
	wire w_dff_B_ogytpNaq0_2;
	wire w_dff_B_Jv6k8U4S0_2;
	wire w_dff_B_iYbHOVF81_2;
	wire w_dff_B_mNivilHR3_2;
	wire w_dff_B_3Bxzm1gu5_2;
	wire w_dff_B_PNOtDNoa6_2;
	wire w_dff_B_V2T9ES6U0_2;
	wire w_dff_B_DxUyRIN37_2;
	wire w_dff_B_suJtMlCG3_2;
	wire w_dff_B_uvYZZWps6_2;
	wire w_dff_B_jOBpItFi5_2;
	wire w_dff_B_pFtKX6H66_2;
	wire w_dff_B_1cJgRuth6_2;
	wire w_dff_B_sGfhoS9A5_2;
	wire w_dff_B_A4o8wSGS5_2;
	wire w_dff_B_z8ukxAKN1_2;
	wire w_dff_B_udZwhBoH5_2;
	wire w_dff_B_Qx1bUMC01_2;
	wire w_dff_B_3VzIIUf90_2;
	wire w_dff_B_9Qkthlom1_2;
	wire w_dff_B_DQDjo2Hn4_2;
	wire w_dff_B_5NGm393O6_2;
	wire w_dff_B_3kFUTehD8_2;
	wire w_dff_B_QKVueGWt5_1;
	wire w_dff_B_UoYNGMjq0_1;
	wire w_dff_B_t5MPMgJ02_2;
	wire w_dff_B_lrW06qFI9_2;
	wire w_dff_B_EoIaXoH00_2;
	wire w_dff_B_GDcqgL9b0_2;
	wire w_dff_B_d1cknSAX0_2;
	wire w_dff_B_iJOkd3Pb9_2;
	wire w_dff_B_g7jpPLsb0_2;
	wire w_dff_B_LQOt9SSH5_2;
	wire w_dff_B_rIUQq1Mi8_2;
	wire w_dff_B_WrZtnV7W3_2;
	wire w_dff_B_1ckAXzvD5_2;
	wire w_dff_B_OiRVNyhP4_2;
	wire w_dff_B_FLveHS3u5_2;
	wire w_dff_B_ppEP7JEA1_2;
	wire w_dff_B_KiWTMxKC7_2;
	wire w_dff_B_dkqkfHcX3_2;
	wire w_dff_B_v0BD1dhP2_2;
	wire w_dff_B_vvUL2odx1_2;
	wire w_dff_B_xDkxHkET9_2;
	wire w_dff_B_DDfNJLV50_2;
	wire w_dff_B_yMK4XQrG6_2;
	wire w_dff_B_E7co62372_2;
	wire w_dff_B_Vs09CW373_2;
	wire w_dff_B_meUnrAjw7_2;
	wire w_dff_B_lnKdbOrZ5_2;
	wire w_dff_B_jEPxsSch6_2;
	wire w_dff_B_1UbQTLs96_2;
	wire w_dff_B_ulXr90JH4_2;
	wire w_dff_B_qB7fgw5D7_2;
	wire w_dff_B_Pey73YRh2_2;
	wire w_dff_B_FZG5XH1I7_2;
	wire w_dff_B_H98D4H0h5_2;
	wire w_dff_B_Xq2bfW3m3_2;
	wire w_dff_B_4wh0O9dz1_2;
	wire w_dff_B_SXKCb8oS9_2;
	wire w_dff_B_cwKLAzCP2_2;
	wire w_dff_B_4HbENNXZ3_2;
	wire w_dff_B_3BE3aLDE4_2;
	wire w_dff_B_Q4sWiyoZ0_2;
	wire w_dff_B_lVKF3b875_2;
	wire w_dff_B_38muVdk36_2;
	wire w_dff_B_yopqtJGK1_2;
	wire w_dff_B_jArYjGoD7_2;
	wire w_dff_B_kT7sBeMi1_2;
	wire w_dff_B_21mEbh8I0_2;
	wire w_dff_B_x71n1UtL6_2;
	wire w_dff_B_Xz6RaKpE9_2;
	wire w_dff_B_ZITUsOKo8_2;
	wire w_dff_B_TF8YGS6n8_2;
	wire w_dff_B_y0gQJKMr9_2;
	wire w_dff_B_A5VmTtr62_2;
	wire w_dff_B_srEb0CD73_2;
	wire w_dff_B_yIM3PIHa5_2;
	wire w_dff_B_bbPAVANc9_2;
	wire w_dff_B_NnziGxkV6_2;
	wire w_dff_B_Tu8GgzAT2_2;
	wire w_dff_B_pvbCDjg29_2;
	wire w_dff_B_jr9uTGXa7_2;
	wire w_dff_B_vsfo1Fp33_2;
	wire w_dff_B_rInyRAr98_2;
	wire w_dff_B_q34B6lAI9_2;
	wire w_dff_B_xXnwfbrR8_2;
	wire w_dff_B_bXNbAUji5_2;
	wire w_dff_B_Gh591ANM2_2;
	wire w_dff_B_3wibqupe7_2;
	wire w_dff_B_QHEbQg640_2;
	wire w_dff_B_uNs538Jp8_2;
	wire w_dff_B_pkx9ikNH4_2;
	wire w_dff_B_yiDogyUX2_2;
	wire w_dff_B_xYrUPg4e8_2;
	wire w_dff_B_jhDuClEt7_2;
	wire w_dff_B_ZAxmcxZr4_2;
	wire w_dff_B_KJJV1X3J4_2;
	wire w_dff_B_VDMfBjA53_2;
	wire w_dff_B_69J16IMU4_2;
	wire w_dff_B_YhxIyYQG3_2;
	wire w_dff_B_2K4ObXET2_2;
	wire w_dff_B_RqV1isF89_2;
	wire w_dff_B_xuQuZlGa8_2;
	wire w_dff_B_R4bdEiuo9_2;
	wire w_dff_B_6MT5HUZl8_2;
	wire w_dff_B_7p8E9svd4_2;
	wire w_dff_B_qOMa1gSn6_2;
	wire w_dff_B_RcHkkidg7_2;
	wire w_dff_B_g5tMIoOe7_2;
	wire w_dff_B_E2sHLCiD5_2;
	wire w_dff_B_g7pGMShE4_2;
	wire w_dff_B_IWFQQsI89_2;
	wire w_dff_B_N4xurE2H7_2;
	wire w_dff_B_ziA82jg42_2;
	wire w_dff_B_2E4qR4cc6_2;
	wire w_dff_B_4Bt6y4zt0_1;
	wire w_dff_B_99QiTFjo3_2;
	wire w_dff_B_puupNxe36_2;
	wire w_dff_B_gmfk8Z0c1_2;
	wire w_dff_B_55CQjVaE2_2;
	wire w_dff_B_YdQAmE2O8_2;
	wire w_dff_B_50zTlLwx8_2;
	wire w_dff_B_EbqiYn3y9_2;
	wire w_dff_B_XKTlDXUp7_2;
	wire w_dff_B_J9eUGxIC7_2;
	wire w_dff_B_upil0NRb5_2;
	wire w_dff_B_XQ00n42s0_2;
	wire w_dff_B_0N8rdUdi5_2;
	wire w_dff_B_op4gHcy56_2;
	wire w_dff_B_zBgIB6pW4_2;
	wire w_dff_B_P18SjuOx9_2;
	wire w_dff_B_8nVLgy2D1_2;
	wire w_dff_B_4UjSdbpg6_2;
	wire w_dff_B_H63wemc78_2;
	wire w_dff_B_TsuXj3H28_2;
	wire w_dff_B_6pSlz7uU4_2;
	wire w_dff_B_1RDq1Ei12_2;
	wire w_dff_B_N5vehd0F0_2;
	wire w_dff_B_smXfCofL7_2;
	wire w_dff_B_fGhviDAs9_2;
	wire w_dff_B_FkjDaoI48_2;
	wire w_dff_B_pTgCKzc72_2;
	wire w_dff_B_kFprMZUL1_2;
	wire w_dff_B_DylwgarZ7_2;
	wire w_dff_B_9Zoh5yMy3_2;
	wire w_dff_B_cQg39ptg1_2;
	wire w_dff_B_W8Se07348_2;
	wire w_dff_B_rTnB1yrs8_2;
	wire w_dff_B_4Lvv8VEr4_2;
	wire w_dff_B_2ELtoSym4_2;
	wire w_dff_B_2hmTYA1d8_2;
	wire w_dff_B_1oIU5lsy4_2;
	wire w_dff_B_8tnOjYpD1_2;
	wire w_dff_B_JFD7i89n1_2;
	wire w_dff_B_Zf8WhofN0_2;
	wire w_dff_B_tHwOVsXV7_2;
	wire w_dff_B_Y9t54LXk6_2;
	wire w_dff_B_mUrMKwmt8_2;
	wire w_dff_B_0DfkFQY61_2;
	wire w_dff_B_GFrhTRzC6_1;
	wire w_dff_B_6xgTCNBr0_1;
	wire w_dff_B_HtI17TAk1_2;
	wire w_dff_B_gAMR6wl58_2;
	wire w_dff_B_KVN4DUkP1_2;
	wire w_dff_B_XxjmFJb54_2;
	wire w_dff_B_v0lSXM3x3_2;
	wire w_dff_B_R7odIVcI1_2;
	wire w_dff_B_ng9zFUrw5_2;
	wire w_dff_B_RqejzdbV0_2;
	wire w_dff_B_HlUJwcvE6_2;
	wire w_dff_B_X7qDLgT79_2;
	wire w_dff_B_bwROm8Dp8_2;
	wire w_dff_B_jDmUArPP6_2;
	wire w_dff_B_z3cttkUb5_2;
	wire w_dff_B_FSJYm9Vn8_2;
	wire w_dff_B_gBK1f5QN1_2;
	wire w_dff_B_36taeYWU1_2;
	wire w_dff_B_NPRxi8OQ9_2;
	wire w_dff_B_buj56fGq6_2;
	wire w_dff_B_L0PTnb5n9_2;
	wire w_dff_B_VWSX9ZV76_2;
	wire w_dff_B_zQI3K1NZ0_2;
	wire w_dff_B_s7afqwyq1_2;
	wire w_dff_B_55siENpu6_2;
	wire w_dff_B_5LFHCW8g7_2;
	wire w_dff_B_Vl9j5ygu2_2;
	wire w_dff_B_u8IcZ4Sm7_2;
	wire w_dff_B_HgXMQ7ya9_2;
	wire w_dff_B_YgMHxllh6_2;
	wire w_dff_B_unGaVVXG1_2;
	wire w_dff_B_Vc7kbnJk1_2;
	wire w_dff_B_1Vbt5vQf8_2;
	wire w_dff_B_6BBe5St64_2;
	wire w_dff_B_3CEOJI8g6_2;
	wire w_dff_B_Cvpd7jbn4_2;
	wire w_dff_B_62vw1PCN2_2;
	wire w_dff_B_g9EhUTMJ3_2;
	wire w_dff_B_PBlEnHlZ2_2;
	wire w_dff_B_Zby2zGPG7_2;
	wire w_dff_B_uhgPa5op1_2;
	wire w_dff_B_GMBo0y002_2;
	wire w_dff_B_uKRD97Xl5_2;
	wire w_dff_B_uJrXNTd85_2;
	wire w_dff_B_pwbLZByw2_2;
	wire w_dff_B_NJqILe4L0_2;
	wire w_dff_B_Uwkfa8z69_2;
	wire w_dff_B_XUthNvBx5_2;
	wire w_dff_B_A0lD3kJz7_2;
	wire w_dff_B_am6QIkWZ5_2;
	wire w_dff_B_vSN9umEr5_2;
	wire w_dff_B_WuM1gtbH4_2;
	wire w_dff_B_OU1O8fij0_2;
	wire w_dff_B_ecMNIr6G1_2;
	wire w_dff_B_BOPwxFL67_2;
	wire w_dff_B_7HtFwwe50_2;
	wire w_dff_B_QEaLeHvU7_2;
	wire w_dff_B_fDy71Ei10_2;
	wire w_dff_B_PmBQaupu9_2;
	wire w_dff_B_srpOVKbr2_2;
	wire w_dff_B_fWM9lthE8_2;
	wire w_dff_B_3nJq1qak6_2;
	wire w_dff_B_JWO8f5rj0_2;
	wire w_dff_B_HMkCkOnn1_2;
	wire w_dff_B_rmpInCQi9_2;
	wire w_dff_B_5LcFkU4d1_2;
	wire w_dff_B_fy6DyESh8_2;
	wire w_dff_B_gGHflhEb5_2;
	wire w_dff_B_6pt5q2tr5_2;
	wire w_dff_B_61jeyu9q3_2;
	wire w_dff_B_GD17m7B46_2;
	wire w_dff_B_8XUYucIN7_2;
	wire w_dff_B_8BIw16mB0_2;
	wire w_dff_B_2Fduc4aY2_2;
	wire w_dff_B_821GBm5b2_2;
	wire w_dff_B_nSgVZuvB2_2;
	wire w_dff_B_THRcDXML9_2;
	wire w_dff_B_DxNT2And2_2;
	wire w_dff_B_UIQV9kfH2_2;
	wire w_dff_B_hqHSZuvW4_2;
	wire w_dff_B_UsfujUSL3_2;
	wire w_dff_B_QZeg2vO21_2;
	wire w_dff_B_RNw92S2o0_2;
	wire w_dff_B_Yf9oaDTh0_2;
	wire w_dff_B_jmMqyqcm9_2;
	wire w_dff_B_FYAmhI927_1;
	wire w_dff_B_hHjWGShV1_2;
	wire w_dff_B_UL9m2h943_2;
	wire w_dff_B_uK8eEL0y1_2;
	wire w_dff_B_qaujD78D0_2;
	wire w_dff_B_e6BIrDic3_2;
	wire w_dff_B_bz3w8n586_2;
	wire w_dff_B_ABBDbDiQ0_2;
	wire w_dff_B_g8wW0jOW5_2;
	wire w_dff_B_veUdx0l33_2;
	wire w_dff_B_jO3H6MLN1_2;
	wire w_dff_B_LYmXvikb1_2;
	wire w_dff_B_LOSSiULb0_2;
	wire w_dff_B_HERjnJit9_2;
	wire w_dff_B_bWRSBSn73_2;
	wire w_dff_B_GWqy7FtZ7_2;
	wire w_dff_B_C509QPgg1_2;
	wire w_dff_B_Fxb7o3wR7_2;
	wire w_dff_B_ruzmsfsF0_2;
	wire w_dff_B_LtLCSeUH3_2;
	wire w_dff_B_Slm2Hbcx8_2;
	wire w_dff_B_SbdBcWsb4_2;
	wire w_dff_B_36GZfrMK8_2;
	wire w_dff_B_3aPlP3zY3_2;
	wire w_dff_B_sdF3dOd54_2;
	wire w_dff_B_qByIQEVR2_2;
	wire w_dff_B_xdbSU1DA6_2;
	wire w_dff_B_nssK0Cdd5_2;
	wire w_dff_B_dNQoKXOx3_2;
	wire w_dff_B_0XHagwRG1_2;
	wire w_dff_B_erVG94Jm5_2;
	wire w_dff_B_O9iQwq537_2;
	wire w_dff_B_zzUhDKMB8_2;
	wire w_dff_B_3vAkFII14_2;
	wire w_dff_B_iRkRLu2k1_2;
	wire w_dff_B_CpE1fB8t3_2;
	wire w_dff_B_OHmUMgqe9_2;
	wire w_dff_B_Big0HdWt4_2;
	wire w_dff_B_nYaLSc6g8_2;
	wire w_dff_B_rQO4g00b5_2;
	wire w_dff_B_xNpPTo8O6_1;
	wire w_dff_B_Hrnhfkl04_1;
	wire w_dff_B_aiAv9iMA3_2;
	wire w_dff_B_4qQoKklD7_2;
	wire w_dff_B_ky0nFzQR3_2;
	wire w_dff_B_DXAkzDQ93_2;
	wire w_dff_B_DJToPCO48_2;
	wire w_dff_B_unAENyFN0_2;
	wire w_dff_B_33wbuzg13_2;
	wire w_dff_B_ZOilHMra3_2;
	wire w_dff_B_xqC0jtwH6_2;
	wire w_dff_B_cuglOGOZ2_2;
	wire w_dff_B_nK7loTJd2_2;
	wire w_dff_B_qMskERQP1_2;
	wire w_dff_B_NxqkiUSf0_2;
	wire w_dff_B_UqrGwyf40_2;
	wire w_dff_B_Nzw9a53j2_2;
	wire w_dff_B_hBXJ9mjI7_2;
	wire w_dff_B_Lan52Tx93_2;
	wire w_dff_B_TgLl0Zq53_2;
	wire w_dff_B_0VmyhUMs9_2;
	wire w_dff_B_yXudTNvo4_2;
	wire w_dff_B_1G4XNrYe0_2;
	wire w_dff_B_3kQhJqD36_2;
	wire w_dff_B_X89BGa8y1_2;
	wire w_dff_B_NMO1wSXk8_2;
	wire w_dff_B_ng0dt2gY4_2;
	wire w_dff_B_gGtKYGyA7_2;
	wire w_dff_B_xs93OViw3_2;
	wire w_dff_B_ckgbo0At9_2;
	wire w_dff_B_xuEFvlmC0_2;
	wire w_dff_B_ysxzvZzi7_2;
	wire w_dff_B_IN8DNn2W9_2;
	wire w_dff_B_uTHUNJco7_2;
	wire w_dff_B_MlXZxz3L3_2;
	wire w_dff_B_YR980bIB9_2;
	wire w_dff_B_7xWgjYg03_2;
	wire w_dff_B_4fxGLIjY0_2;
	wire w_dff_B_ahMLwZnv2_2;
	wire w_dff_B_DoWjBlSB7_2;
	wire w_dff_B_P2XHzwit2_2;
	wire w_dff_B_luz8iKn08_2;
	wire w_dff_B_i1p9MT3M9_2;
	wire w_dff_B_EGjfu9GG1_2;
	wire w_dff_B_0ZJYfDSc2_2;
	wire w_dff_B_zL4NKhxe8_2;
	wire w_dff_B_Ydpl4CyJ9_2;
	wire w_dff_B_DnFdFUol0_2;
	wire w_dff_B_MRjghXZe9_2;
	wire w_dff_B_IMoRia2E5_2;
	wire w_dff_B_O37zx7IJ9_2;
	wire w_dff_B_mst2NUll6_2;
	wire w_dff_B_h9AEQIZW8_2;
	wire w_dff_B_6pY2AjZt4_2;
	wire w_dff_B_otJtoaek1_2;
	wire w_dff_B_NHdx7Krz7_2;
	wire w_dff_B_JOO2VYIq7_2;
	wire w_dff_B_3NExsbid3_2;
	wire w_dff_B_Ky1UEWae1_2;
	wire w_dff_B_r2HUpSFV1_2;
	wire w_dff_B_Yln5KWxh8_2;
	wire w_dff_B_3U6QBMYZ3_2;
	wire w_dff_B_15MVkSzs4_2;
	wire w_dff_B_JYu6r52R4_2;
	wire w_dff_B_D5NHkI6b2_2;
	wire w_dff_B_cpcDl0Io7_2;
	wire w_dff_B_T2QZDKY06_2;
	wire w_dff_B_e9FP3Sq65_2;
	wire w_dff_B_s9AsVBm07_2;
	wire w_dff_B_auyUwOzI0_2;
	wire w_dff_B_TZbnHOKy5_2;
	wire w_dff_B_D7GJBkBS3_2;
	wire w_dff_B_Pk1qeRbR0_2;
	wire w_dff_B_iyL8tIMv1_2;
	wire w_dff_B_4MBxpGec8_2;
	wire w_dff_B_2q3rfz6I1_2;
	wire w_dff_B_NRAchYUb4_2;
	wire w_dff_B_WSfU75pS8_1;
	wire w_dff_B_9YqY937n1_2;
	wire w_dff_B_TW2XgW4e9_2;
	wire w_dff_B_YrWW2sWS9_2;
	wire w_dff_B_BZ5ZWk8T9_2;
	wire w_dff_B_dK7QjaNy4_2;
	wire w_dff_B_b49xwTzO0_2;
	wire w_dff_B_27NgSyOQ6_2;
	wire w_dff_B_TNSyfA4P2_2;
	wire w_dff_B_58Ra11ci7_2;
	wire w_dff_B_yvvCVGsR9_2;
	wire w_dff_B_IIAeljsp1_2;
	wire w_dff_B_T2OsNlBx2_2;
	wire w_dff_B_IIuxMkak0_2;
	wire w_dff_B_S4hAwUkp0_2;
	wire w_dff_B_Xx5hVm8c0_2;
	wire w_dff_B_q6150sBa4_2;
	wire w_dff_B_gGVaxCJh9_2;
	wire w_dff_B_7RVl3BZv2_2;
	wire w_dff_B_u3wzTDDL2_2;
	wire w_dff_B_qz7PjDcJ2_2;
	wire w_dff_B_8CZyNRgL3_2;
	wire w_dff_B_2mkUKDoB5_2;
	wire w_dff_B_Ej8lV7WY5_2;
	wire w_dff_B_AtOxWHWd8_2;
	wire w_dff_B_cADvcp5S9_2;
	wire w_dff_B_I6kc8B7O6_2;
	wire w_dff_B_el5nAwQ95_2;
	wire w_dff_B_1bqxx8AJ0_2;
	wire w_dff_B_xhKGldnU6_2;
	wire w_dff_B_knhMGzkE6_2;
	wire w_dff_B_vWwshD5o0_2;
	wire w_dff_B_W1Z4epbj6_2;
	wire w_dff_B_BNTCPf5U2_2;
	wire w_dff_B_RdvNckQa5_2;
	wire w_dff_B_8WbYio3T6_2;
	wire w_dff_B_wVC0Od8X5_1;
	wire w_dff_B_p0m5Rv4t8_1;
	wire w_dff_B_hsVj3i1c3_2;
	wire w_dff_B_ZT0dNhtU2_2;
	wire w_dff_B_GPC05KQe3_2;
	wire w_dff_B_BC8DyLQX1_2;
	wire w_dff_B_q7KhCkDr1_2;
	wire w_dff_B_fwS1yGYl4_2;
	wire w_dff_B_J07C6Oyn3_2;
	wire w_dff_B_6oAxxxwR9_2;
	wire w_dff_B_1Gq7FYcR8_2;
	wire w_dff_B_TEmXnqMZ0_2;
	wire w_dff_B_6hKH2YtQ9_2;
	wire w_dff_B_Z8QBaZt10_2;
	wire w_dff_B_KkWRe1nx5_2;
	wire w_dff_B_UfwHAyvR2_2;
	wire w_dff_B_9jJtGC1b4_2;
	wire w_dff_B_ml0YPfgJ6_2;
	wire w_dff_B_jU4cg11p9_2;
	wire w_dff_B_YJnKEkYz6_2;
	wire w_dff_B_mtI54M7h6_2;
	wire w_dff_B_kngdEsDq6_2;
	wire w_dff_B_2sg2GHlP5_2;
	wire w_dff_B_8WaSW2uw4_2;
	wire w_dff_B_qH1qv8SU0_2;
	wire w_dff_B_AMlJ2WeA6_2;
	wire w_dff_B_JvsFduZG8_2;
	wire w_dff_B_lABYoHf46_2;
	wire w_dff_B_AkWFt7wP1_2;
	wire w_dff_B_JUlQF8ek7_2;
	wire w_dff_B_uicXuqRs0_2;
	wire w_dff_B_KAfbg7po1_2;
	wire w_dff_B_E7J8dNYc1_2;
	wire w_dff_B_b1k1UvD19_2;
	wire w_dff_B_qzyA06vm8_2;
	wire w_dff_B_2kB1rdeo4_2;
	wire w_dff_B_i3kPQFn68_2;
	wire w_dff_B_rBbVVXzk3_2;
	wire w_dff_B_OLMdOwMG3_2;
	wire w_dff_B_b6NPsDK31_2;
	wire w_dff_B_ybw575GR9_2;
	wire w_dff_B_dy9kZaq41_2;
	wire w_dff_B_uwIXpi7K9_2;
	wire w_dff_B_cWXnl7XS5_2;
	wire w_dff_B_KTN1cKTp9_2;
	wire w_dff_B_x1cTF8kr4_2;
	wire w_dff_B_LeIqCTrk5_2;
	wire w_dff_B_vWCYQ6mF5_2;
	wire w_dff_B_PBmy3mMv5_2;
	wire w_dff_B_mQBbPX3g1_2;
	wire w_dff_B_f65ZQx3T4_2;
	wire w_dff_B_czRJXl6b0_2;
	wire w_dff_B_YzHV5fm95_2;
	wire w_dff_B_Dg4U9h9C8_2;
	wire w_dff_B_0PjPSnM23_2;
	wire w_dff_B_xJNoHB8o2_2;
	wire w_dff_B_Mr35CR9c0_2;
	wire w_dff_B_zV26xBQO9_2;
	wire w_dff_B_UTC1WjZF3_2;
	wire w_dff_B_LA4S2oE08_2;
	wire w_dff_B_fRWjaOCM8_2;
	wire w_dff_B_9kTK7JHq5_2;
	wire w_dff_B_O9MgvkTA0_2;
	wire w_dff_B_TKdnRh3l9_2;
	wire w_dff_B_E6ymctXg9_2;
	wire w_dff_B_09sY0hXy6_2;
	wire w_dff_B_5ocwuLjD9_2;
	wire w_dff_B_fpEPPbdR3_2;
	wire w_dff_B_DoJLaGXc5_2;
	wire w_dff_B_bBKY3IsN3_1;
	wire w_dff_B_S0E1Sgjj8_2;
	wire w_dff_B_ihIBvree0_2;
	wire w_dff_B_2iquHi9D1_2;
	wire w_dff_B_CzZ6HtAg6_2;
	wire w_dff_B_kKufEeyC7_2;
	wire w_dff_B_yTZrpuH99_2;
	wire w_dff_B_Bu3Tw3l13_2;
	wire w_dff_B_M18nt3R75_2;
	wire w_dff_B_D1fpOwLX2_2;
	wire w_dff_B_zmWh65cA3_2;
	wire w_dff_B_uxgOLdre9_2;
	wire w_dff_B_hWPQHs9E8_2;
	wire w_dff_B_HTuYlEEF3_2;
	wire w_dff_B_jrhrHsHm6_2;
	wire w_dff_B_BH59cvnu4_2;
	wire w_dff_B_omuUOhtQ2_2;
	wire w_dff_B_ODdj48S42_2;
	wire w_dff_B_kHniHcMu6_2;
	wire w_dff_B_WqFMNQPa6_2;
	wire w_dff_B_IG64Vhwe4_2;
	wire w_dff_B_FUQTqP3s7_2;
	wire w_dff_B_ppIssLh38_2;
	wire w_dff_B_7ujWo1wp4_2;
	wire w_dff_B_xnWLW3Hf4_2;
	wire w_dff_B_wAT6RGA13_2;
	wire w_dff_B_7AnPn6AK1_2;
	wire w_dff_B_cuNydATm6_2;
	wire w_dff_B_mry06MKl3_2;
	wire w_dff_B_B9OZct8I1_2;
	wire w_dff_B_EVsL6J9n5_2;
	wire w_dff_B_e01CU9l05_2;
	wire w_dff_B_dmn7JpAz0_1;
	wire w_dff_B_4Q00MYR71_1;
	wire w_dff_B_scurrzbR6_2;
	wire w_dff_B_fuhby7C86_2;
	wire w_dff_B_mDgyuTP89_2;
	wire w_dff_B_da6GawuY7_2;
	wire w_dff_B_QXIo7UYj7_2;
	wire w_dff_B_KQ1pBGtY2_2;
	wire w_dff_B_uOkudGRp9_2;
	wire w_dff_B_CzTm0Stv3_2;
	wire w_dff_B_cknq3JRn7_2;
	wire w_dff_B_ws6DwHoa7_2;
	wire w_dff_B_EQiyyne30_2;
	wire w_dff_B_4Vbre3vb8_2;
	wire w_dff_B_qy4THqZw2_2;
	wire w_dff_B_w5pch2gz4_2;
	wire w_dff_B_nH2gAAy46_2;
	wire w_dff_B_XLGlIs8w1_2;
	wire w_dff_B_7R8rTkqg7_2;
	wire w_dff_B_q1b0CAl68_2;
	wire w_dff_B_zPg8FF8V3_2;
	wire w_dff_B_6RPAaIEA7_2;
	wire w_dff_B_XmjSXXtT9_2;
	wire w_dff_B_SccjLZju5_2;
	wire w_dff_B_mmlEdfil5_2;
	wire w_dff_B_WRsAhEQ13_2;
	wire w_dff_B_ENUEjEXN2_2;
	wire w_dff_B_Zf4A8C0H6_2;
	wire w_dff_B_6MRi33Rv2_2;
	wire w_dff_B_HTirBmXv6_2;
	wire w_dff_B_9Wk412pn0_2;
	wire w_dff_B_grQkBCCC6_2;
	wire w_dff_B_te9FeiMN5_2;
	wire w_dff_B_qCGkUKpX2_2;
	wire w_dff_B_fYafNUsP7_2;
	wire w_dff_B_5a2WX4Mw9_2;
	wire w_dff_B_E8VE4UNc9_2;
	wire w_dff_B_MBIVnSCj8_2;
	wire w_dff_B_2vh6456A7_2;
	wire w_dff_B_xngfjrw92_2;
	wire w_dff_B_1GR3noE43_2;
	wire w_dff_B_bhIN0PzF4_2;
	wire w_dff_B_dDvhnWjM9_2;
	wire w_dff_B_U6fTCYAX7_2;
	wire w_dff_B_JT229aKv2_2;
	wire w_dff_B_XvQqza6q9_2;
	wire w_dff_B_czJwQZmA5_2;
	wire w_dff_B_0qeOyR0j8_2;
	wire w_dff_B_VY8LuFNI5_2;
	wire w_dff_B_x6QElvNv7_2;
	wire w_dff_B_I9Kzl9jC0_2;
	wire w_dff_B_rlqbqyq75_2;
	wire w_dff_B_8q8zOGDW6_2;
	wire w_dff_B_iRAklezC6_2;
	wire w_dff_B_YXSfQCqT9_2;
	wire w_dff_B_8uXW4JLO6_2;
	wire w_dff_B_9VziUF1K0_2;
	wire w_dff_B_sGHKFza19_2;
	wire w_dff_B_4tJZXsBh5_2;
	wire w_dff_B_BLj5OV3O9_2;
	wire w_dff_B_J0E8nPgL3_2;
	wire w_dff_B_LWNVmBBi8_1;
	wire w_dff_B_XIF0rP9a6_2;
	wire w_dff_B_lo71QW9n0_2;
	wire w_dff_B_aEbaNfxu6_2;
	wire w_dff_B_auFmes176_2;
	wire w_dff_B_74P68oUx6_2;
	wire w_dff_B_QPTXPFBP8_2;
	wire w_dff_B_Cs6xXPxZ2_2;
	wire w_dff_B_mRKdPi8a7_2;
	wire w_dff_B_Unfnpv300_2;
	wire w_dff_B_Nsz6DUQ24_2;
	wire w_dff_B_l39oDSQO8_2;
	wire w_dff_B_fJxi8moJ3_2;
	wire w_dff_B_vCFdGXyA6_2;
	wire w_dff_B_7ku762rr3_2;
	wire w_dff_B_1TRYjNuL0_2;
	wire w_dff_B_LQ5cLO5H0_2;
	wire w_dff_B_oj15eDZ95_2;
	wire w_dff_B_jwGDfejS6_2;
	wire w_dff_B_gfDtRAlj2_2;
	wire w_dff_B_ZyHxGm152_2;
	wire w_dff_B_WmQrnVJf4_2;
	wire w_dff_B_zKUzstGZ3_2;
	wire w_dff_B_DfpeIN7G4_2;
	wire w_dff_B_SLJ8rhx79_2;
	wire w_dff_B_d3ki5epJ3_2;
	wire w_dff_B_tnVmR1Is8_2;
	wire w_dff_B_jxzYtriR6_2;
	wire w_dff_B_MglutVNZ3_1;
	wire w_dff_B_CzlX2EJb3_1;
	wire w_dff_B_24lQ92Uj5_2;
	wire w_dff_B_VqePKXnN5_2;
	wire w_dff_B_luNLzTs68_2;
	wire w_dff_B_CfEQACIT1_2;
	wire w_dff_B_oU9vCJA57_2;
	wire w_dff_B_I5s5Yn1E4_2;
	wire w_dff_B_8DoLXLE22_2;
	wire w_dff_B_pEmF8jXS9_2;
	wire w_dff_B_bAkR8X8O4_2;
	wire w_dff_B_jn9Hd0rS2_2;
	wire w_dff_B_liOd6g2o0_2;
	wire w_dff_B_iCqlXK5G2_2;
	wire w_dff_B_KYStjnHp2_2;
	wire w_dff_B_svIlcXZ58_2;
	wire w_dff_B_ZyP1ffpY5_2;
	wire w_dff_B_iqVRy71S2_2;
	wire w_dff_B_je1NiQkl5_2;
	wire w_dff_B_JP53Soyp6_2;
	wire w_dff_B_zxRBowWI9_2;
	wire w_dff_B_45ysJ7Du6_2;
	wire w_dff_B_QHMbO7P43_2;
	wire w_dff_B_LzDVF6rA3_2;
	wire w_dff_B_cFXRF5md3_2;
	wire w_dff_B_20Kyx2j61_2;
	wire w_dff_B_92FKZmHE8_2;
	wire w_dff_B_1icfifE90_2;
	wire w_dff_B_Aem7Old88_2;
	wire w_dff_B_aw4v8y6v6_2;
	wire w_dff_B_cQGfxCNI5_2;
	wire w_dff_B_NiD73eUP4_2;
	wire w_dff_B_wKV4GvXD7_2;
	wire w_dff_B_WdkR7PEB2_2;
	wire w_dff_B_3lHCz7hc8_2;
	wire w_dff_B_MDjeQiY99_2;
	wire w_dff_B_I2zqQL898_2;
	wire w_dff_B_MI3Y3TUG8_2;
	wire w_dff_B_DccHJvuu3_2;
	wire w_dff_B_2Ss5OX0X1_2;
	wire w_dff_B_FtBqalmJ7_2;
	wire w_dff_B_XqVAPHix5_2;
	wire w_dff_B_ihROzAI25_2;
	wire w_dff_B_BGrJD9gu5_2;
	wire w_dff_B_mZxX5Rsn6_2;
	wire w_dff_B_srjii0rw8_2;
	wire w_dff_B_DuFglYDS0_2;
	wire w_dff_B_nAVRZE284_2;
	wire w_dff_B_CEhV7ef81_2;
	wire w_dff_B_wRiG9jvG0_2;
	wire w_dff_B_xncYHh4L1_2;
	wire w_dff_B_hYRIFJQP7_2;
	wire w_dff_B_eCwWw4tB1_2;
	wire w_dff_B_0k0xiUEN0_1;
	wire w_dff_B_dAFThpXq4_2;
	wire w_dff_B_aXsj5ag90_2;
	wire w_dff_B_UjqjOdZq3_2;
	wire w_dff_B_Fd2Zhzq67_2;
	wire w_dff_B_omlmCLLu2_2;
	wire w_dff_B_G5DPJV9X7_2;
	wire w_dff_B_hIU0b7953_2;
	wire w_dff_B_IxtO8r7g2_2;
	wire w_dff_B_eQnNQWVM4_2;
	wire w_dff_B_cWaK1ZaQ8_2;
	wire w_dff_B_uHwp6gUm2_2;
	wire w_dff_B_HcDL6hYO4_2;
	wire w_dff_B_6sKYNW9V3_2;
	wire w_dff_B_bPYMBBJD3_2;
	wire w_dff_B_fRCMW0K32_2;
	wire w_dff_B_04kN3zBI2_2;
	wire w_dff_B_aT2rmnRT5_2;
	wire w_dff_B_9jdbiOqK4_2;
	wire w_dff_B_H6KYvTQw7_2;
	wire w_dff_B_qZKyA1Ne3_2;
	wire w_dff_B_OJ5jeE0E4_2;
	wire w_dff_B_adR5r4CT0_2;
	wire w_dff_B_1jCtZI1E6_2;
	wire w_dff_B_CnGbuHTM8_1;
	wire w_dff_B_yvVQoDbq7_1;
	wire w_dff_B_WemccfOp4_2;
	wire w_dff_B_aQG8d6OU9_2;
	wire w_dff_B_OdQAZ9Am7_2;
	wire w_dff_B_MB6ov2St0_2;
	wire w_dff_B_d8dcbpx88_2;
	wire w_dff_B_ciU02CoR8_2;
	wire w_dff_B_ywrgHNzR9_2;
	wire w_dff_B_nstDVpDs8_2;
	wire w_dff_B_wlr0YWQL8_2;
	wire w_dff_B_RsW0tuP66_2;
	wire w_dff_B_3p1hX5M57_2;
	wire w_dff_B_XYhPx7PJ1_2;
	wire w_dff_B_KsAvWhQ68_2;
	wire w_dff_B_ZCZzxZ5k2_2;
	wire w_dff_B_oSPh2pBG4_2;
	wire w_dff_B_l9nU6ptR2_2;
	wire w_dff_B_F15NscN18_2;
	wire w_dff_B_Wo2KnIhZ1_2;
	wire w_dff_B_D9ArtEgt2_2;
	wire w_dff_B_1Mlva9xD5_2;
	wire w_dff_B_IPzQLyDL4_2;
	wire w_dff_B_7Zpip4VS2_2;
	wire w_dff_B_4Vnrbr6y4_2;
	wire w_dff_B_089zXg7m1_2;
	wire w_dff_B_DLpVpjLg4_2;
	wire w_dff_B_6Gjf5fC50_2;
	wire w_dff_B_7qitiaO06_2;
	wire w_dff_B_bS2gYdg69_2;
	wire w_dff_B_KlAJC3fs6_2;
	wire w_dff_B_xvjmtu9Y6_2;
	wire w_dff_B_lp3dBn8P0_2;
	wire w_dff_B_iahT1t9A2_2;
	wire w_dff_B_bZDlMVdR8_2;
	wire w_dff_B_IbroD1ny2_2;
	wire w_dff_B_MQCCYPdm0_2;
	wire w_dff_B_ruqNx9nc0_2;
	wire w_dff_B_vHUPRim29_2;
	wire w_dff_B_yffsoico2_2;
	wire w_dff_B_LIoIJQCz5_2;
	wire w_dff_B_ch5qPKIW8_2;
	wire w_dff_B_RlL0fRtE4_2;
	wire w_dff_B_k8Ala0aO3_2;
	wire w_dff_B_Dh6JNuk36_2;
	wire w_dff_B_qudcE3uE2_1;
	wire w_dff_B_iiRm5VJO6_2;
	wire w_dff_B_osfoBoGh4_2;
	wire w_dff_B_RNAiMMtZ9_2;
	wire w_dff_B_xn9o05H20_2;
	wire w_dff_B_Nz7ycwM99_2;
	wire w_dff_B_EXBJhQLh2_2;
	wire w_dff_B_uoYL7YAf0_2;
	wire w_dff_B_Kc9WJSp76_2;
	wire w_dff_B_Dvx2WFBE6_2;
	wire w_dff_B_o2JZBoql4_2;
	wire w_dff_B_ElPwNQEa3_2;
	wire w_dff_B_xuNH8mrY4_2;
	wire w_dff_B_GcsqxNbq7_2;
	wire w_dff_B_mYS8SCNT5_2;
	wire w_dff_B_X7AgxXXx9_2;
	wire w_dff_B_mUIbw0n03_2;
	wire w_dff_B_kmn7GrF83_2;
	wire w_dff_B_dye1D9Xh4_2;
	wire w_dff_B_zz2U9j7y4_2;
	wire w_dff_B_hzgYHQ3m3_1;
	wire w_dff_B_VUJ8kK6J4_1;
	wire w_dff_B_XUwPFccG1_2;
	wire w_dff_B_qDf8yzvU8_2;
	wire w_dff_B_YfFESv7Y2_2;
	wire w_dff_B_6hGqH0oQ4_2;
	wire w_dff_B_meMNprm84_2;
	wire w_dff_B_Eaa4tlWh8_2;
	wire w_dff_B_KMoxkrgq0_2;
	wire w_dff_B_Ux04TXkM2_2;
	wire w_dff_B_tGhiMtQG1_2;
	wire w_dff_B_1rwjxNxj5_2;
	wire w_dff_B_sOGu36Ju5_2;
	wire w_dff_B_cxoNxekd9_2;
	wire w_dff_B_euAX7Zcr6_2;
	wire w_dff_B_tSq8EBt09_2;
	wire w_dff_B_6O732Ypn7_2;
	wire w_dff_B_q0E3ocqJ8_2;
	wire w_dff_B_r6SG1ciY6_2;
	wire w_dff_B_oHPu7e6b0_2;
	wire w_dff_B_CwIFVtBx7_2;
	wire w_dff_B_ncpZs0IK5_2;
	wire w_dff_B_c4XT9CKg9_2;
	wire w_dff_B_mZOzL4Oo1_2;
	wire w_dff_B_q7o620Wi1_2;
	wire w_dff_B_wzOJCRbd9_2;
	wire w_dff_B_OVmNq2RK6_2;
	wire w_dff_B_2jbcJW0z1_2;
	wire w_dff_B_B1T78iHV5_2;
	wire w_dff_B_yBkBYxM09_2;
	wire w_dff_B_1zay1wks4_2;
	wire w_dff_B_gYPRlT7H4_2;
	wire w_dff_B_yY6qZYRD5_2;
	wire w_dff_B_hUt2ukSY0_2;
	wire w_dff_B_P0PV6YsP7_2;
	wire w_dff_B_l7vSSOB04_2;
	wire w_dff_B_gXAYdozV7_2;
	wire w_dff_B_3kYMEyRn3_1;
	wire w_dff_B_MWdZUw5y2_2;
	wire w_dff_B_LqlzNphT4_2;
	wire w_dff_B_nj9zwWel5_2;
	wire w_dff_B_hYDwZY0m3_2;
	wire w_dff_B_IDqj7peY7_2;
	wire w_dff_B_HQYJAkKg8_2;
	wire w_dff_B_qVhPU3vs7_2;
	wire w_dff_B_mBYEv04h1_2;
	wire w_dff_B_Ql9u6AKD5_2;
	wire w_dff_B_yxJc6eEw4_2;
	wire w_dff_B_SoV47NXv2_2;
	wire w_dff_B_TakxGcfK5_2;
	wire w_dff_B_OJf8jh5j0_2;
	wire w_dff_B_hAx1BpvH7_2;
	wire w_dff_B_n8FDE26z7_2;
	wire w_dff_B_DXKOYRm12_2;
	wire w_dff_B_915OFzsM2_2;
	wire w_dff_B_Qe6BCVrA4_2;
	wire w_dff_B_OwqyJRuL6_2;
	wire w_dff_B_UYvk1XaJ9_2;
	wire w_dff_B_63czp9M95_2;
	wire w_dff_B_PoIkLgfo5_2;
	wire w_dff_B_lJSoJzUj9_2;
	wire w_dff_B_jnyN9bbn6_2;
	wire w_dff_B_VyhTxvWP0_2;
	wire w_dff_B_fJPyw12V8_2;
	wire w_dff_B_TRYhdKbR3_2;
	wire w_dff_B_XgHBT7UW8_2;
	wire w_dff_B_98jFRaQa7_2;
	wire w_dff_B_nE0TC1Ml7_2;
	wire w_dff_B_FGJPNzIn4_2;
	wire w_dff_B_3faphIZx1_2;
	wire w_dff_B_CegCFhZV5_2;
	wire w_dff_B_XXuOwCFI6_2;
	wire w_dff_B_X4cpIIKq4_2;
	wire w_dff_B_SkwsX9Kf0_2;
	wire w_dff_B_ZALXm2qD7_2;
	wire w_dff_B_wisMNCrq6_2;
	wire w_dff_B_fmfsgtvM9_2;
	wire w_dff_B_WtDL9gqU3_2;
	wire w_dff_B_Xn6nswdx1_2;
	wire w_dff_B_ZkUGvUdg8_2;
	wire w_dff_B_XdgiEJGx6_1;
	wire w_dff_B_8ojOxZMk7_2;
	wire w_dff_B_KHBwC0mO7_2;
	wire w_dff_B_L9tymt2o7_2;
	wire w_dff_B_gCEoc0ok0_2;
	wire w_dff_B_MPxCxC8F7_2;
	wire w_dff_B_GkVu1s132_2;
	wire w_dff_B_81nsxWVJ6_2;
	wire w_dff_B_xftHJnTj0_2;
	wire w_dff_B_jdfI6LIz8_2;
	wire w_dff_B_WuLqmkvo0_2;
	wire w_dff_B_ZwivAUV38_2;
	wire w_dff_A_XIjrmA6j7_0;
	wire w_dff_A_RnJEbFAG9_0;
	wire w_dff_A_QejrMFgQ1_0;
	wire w_dff_B_BWx1odqe4_2;
	wire w_dff_B_hLKPFkcp0_1;
	wire w_dff_B_WKbR0yNr9_1;
	wire w_dff_B_2L9qJ39V7_1;
	wire w_dff_B_QyGA5kwr6_1;
	wire w_dff_B_2ajsOZOZ6_1;
	wire w_dff_B_Ey840Zsi9_1;
	wire w_dff_B_lNYAzxww7_1;
	wire w_dff_B_bNAI5svb2_1;
	wire w_dff_A_mVit9xwJ2_1;
	wire w_dff_A_AZd2pNcg9_1;
	wire w_dff_A_ZYScIdGK7_1;
	wire w_dff_A_RuE7Rnip8_1;
	wire w_dff_A_1rfP5BYn6_1;
	wire w_dff_A_j2WdFBsr8_1;
	wire w_dff_A_x4eBRqMp2_1;
	wire w_dff_B_OdCm1bZC7_2;
	wire w_dff_B_yuwvpGbi1_2;
	wire w_dff_B_CrfCmex16_2;
	wire w_dff_B_SLp8eusp2_2;
	wire w_dff_B_9k9VjoeR7_2;
	wire w_dff_B_1LKT2Gyp5_2;
	wire w_dff_B_70ZJ2Mv85_2;
	wire w_dff_B_B9mgERzy1_2;
	wire w_dff_B_HO2IAvlh3_2;
	wire w_dff_B_hwGPVRFa1_2;
	wire w_dff_B_dGU27aM66_1;
	wire w_dff_B_4bTIsIFD2_2;
	wire w_dff_B_63rqYGLh9_2;
	wire w_dff_B_TEqF3pxj1_2;
	wire w_dff_B_6SuRuAjx5_2;
	wire w_dff_B_yEBdZkIb7_2;
	wire w_dff_B_XFdW4tmv0_2;
	wire w_dff_B_DOlnnmWH3_2;
	wire w_dff_B_fFN9NgEZ6_2;
	wire w_dff_B_EqFFoG9E7_2;
	wire w_dff_B_gh7giJJg6_2;
	wire w_dff_B_CPHW86HD7_2;
	wire w_dff_B_dgeRzY9T7_2;
	wire w_dff_B_WsuEKtQ94_2;
	wire w_dff_A_QAVTmnh25_0;
	wire w_dff_A_uvHSWtwa2_0;
	wire w_dff_A_N9UzwRK64_0;
	wire w_dff_A_t44wiNYu7_0;
	wire w_dff_A_QHOwzUSP9_1;
	wire w_dff_A_3cWmQLSM5_1;
	wire w_dff_B_hDAG1rPw4_1;
	wire w_dff_B_ivgsdJ9S8_1;
	wire w_dff_B_Y0XRAVZb6_1;
	wire w_dff_B_debJB5Lr6_1;
	wire w_dff_B_EWZpWhAQ7_1;
	wire w_dff_A_l0fFdRyQ1_0;
	wire w_dff_A_EHBpv6gX8_0;
	wire w_dff_A_UYrp90wJ3_0;
	wire w_dff_A_H5gxb2DF1_0;
	wire w_dff_A_zqS5QNMI5_0;
	wire w_dff_A_WbOULxLr1_0;
	wire w_dff_B_Ycy7sUPW7_2;
	wire w_dff_A_3d3NyK4D6_1;
	wire w_dff_A_GAtiqGUf0_1;
	wire w_dff_A_Rese1iCp1_1;
	wire w_dff_A_L2EGjFho3_1;
	wire w_dff_A_QgymNIau6_1;
	wire w_dff_A_qLYUvskc7_1;
	wire w_dff_A_sPfUjL1l8_0;
	wire w_dff_A_NE2GPuAv3_0;
	wire w_dff_A_PShVza2c8_0;
	wire w_dff_A_0zm7ulG42_0;
	wire w_dff_A_j5VviUPL2_0;
	wire w_dff_A_tTC9FYLk4_0;
	wire w_dff_A_eAwVwr0k7_0;
	wire w_dff_A_74UJSTH11_0;
	wire w_dff_A_64C90BHz5_0;
	wire w_dff_A_mrCsYqBD2_0;
	wire w_dff_A_ol9UgZWG4_0;
	wire w_dff_A_9flp1qGQ0_0;
	wire w_dff_A_t283ZKbl5_0;
	wire w_dff_A_Ha7xGOky4_0;
	wire w_dff_A_6uhpB0TI7_0;
	wire w_dff_A_FvP308hJ6_0;
	wire w_dff_A_1ibXjjTB8_0;
	wire w_dff_A_C57Ap0IH4_0;
	wire w_dff_A_Q46xReL81_0;
	wire w_dff_A_GwArLYlx8_0;
	wire w_dff_A_j4xyXNnf3_0;
	wire w_dff_A_7ISzBbUm8_0;
	wire w_dff_A_NRZdd1iT2_0;
	wire w_dff_A_oxjuRczw8_0;
	wire w_dff_A_HH0UcsaP7_0;
	wire w_dff_A_Jy3zRvlp3_0;
	wire w_dff_A_ja392aA08_0;
	wire w_dff_A_7QTZYZG49_0;
	wire w_dff_A_kjOKyZAa7_0;
	wire w_dff_A_jb79drfl2_0;
	wire w_dff_A_dkvrzT458_0;
	wire w_dff_A_qkk441TT3_0;
	wire w_dff_A_yWZ5wtNx4_0;
	wire w_dff_A_yUhV3XZu0_0;
	wire w_dff_A_T8KygEKp3_0;
	wire w_dff_A_QZHR3Mel1_0;
	wire w_dff_A_5Xdqzr8V9_0;
	wire w_dff_A_GcQnaqOF9_0;
	wire w_dff_A_AW643vpz2_0;
	wire w_dff_A_BOEsfZn71_0;
	wire w_dff_A_quydwrrO7_0;
	wire w_dff_A_lXfelNFT5_0;
	wire w_dff_A_Manmdn8F2_0;
	wire w_dff_A_Xuv4eNEh6_0;
	wire w_dff_A_mj5JHtcG4_0;
	wire w_dff_A_lr5i5jJ84_0;
	wire w_dff_A_0g0SfOiE8_0;
	wire w_dff_A_nuRitZCD0_0;
	wire w_dff_A_kAkSPkP93_0;
	wire w_dff_A_Up5xdlKm4_0;
	wire w_dff_A_d5qXlybP4_0;
	wire w_dff_A_mHEjEAwr8_0;
	wire w_dff_A_wiBrkzwd7_0;
	wire w_dff_A_QiXHZho40_0;
	wire w_dff_A_twFiy3y93_0;
	wire w_dff_A_qcCVN0BH5_0;
	wire w_dff_A_SlszP6vW7_0;
	wire w_dff_A_78x6wCWu6_0;
	wire w_dff_A_3lSMzqo55_0;
	wire w_dff_A_BLmCA7UH9_0;
	wire w_dff_A_uZLHxEEa3_0;
	wire w_dff_A_FSmdya4s2_0;
	wire w_dff_A_nyYDZOFl4_0;
	wire w_dff_A_q6O22de35_0;
	wire w_dff_A_hAS4SyhA4_0;
	wire w_dff_A_eDbKs2iV5_0;
	wire w_dff_A_ozHjHBjO1_0;
	wire w_dff_A_aRO1PoMv3_0;
	wire w_dff_A_iSJBwK9L3_0;
	wire w_dff_A_c7m5qKbU6_0;
	wire w_dff_A_mWuGthc55_0;
	wire w_dff_A_OStBu9fY9_0;
	wire w_dff_A_yTWRKoSS5_0;
	wire w_dff_A_cGgknGSv6_0;
	wire w_dff_A_oHlkIbp78_2;
	wire w_dff_A_Ioca4err9_0;
	wire w_dff_A_lpOZ5Fvf1_0;
	wire w_dff_A_LFXldfUV3_0;
	wire w_dff_A_xOJhOIUo9_0;
	wire w_dff_A_j22KwikW4_0;
	wire w_dff_A_pfopnZP06_0;
	wire w_dff_A_ICeAF8Rv5_0;
	wire w_dff_A_ZQbp5s5K0_0;
	wire w_dff_A_YlHX0BwN2_0;
	wire w_dff_A_ETy9gqGD1_0;
	wire w_dff_A_tezJ3UVG9_0;
	wire w_dff_A_nDsct10I7_0;
	wire w_dff_A_pkxGh6lD7_0;
	wire w_dff_A_IoOVz7to6_0;
	wire w_dff_A_ffVc2a3L0_0;
	wire w_dff_A_GpB6YlP24_0;
	wire w_dff_A_jT9aZRKk7_0;
	wire w_dff_A_5PaOZazT8_0;
	wire w_dff_A_wseCQdZJ7_0;
	wire w_dff_A_ViE1QtRD1_0;
	wire w_dff_A_aYFLuSr96_0;
	wire w_dff_A_YoHzFePB3_0;
	wire w_dff_A_3YhlgYa31_0;
	wire w_dff_A_fQwfeTq67_0;
	wire w_dff_A_a55hHrgC9_0;
	wire w_dff_A_YmbmVZ1Y5_0;
	wire w_dff_A_noCuUxlZ2_0;
	wire w_dff_A_6uwxm9735_0;
	wire w_dff_A_M1eDYs1t8_0;
	wire w_dff_A_ZLrn5UZR6_0;
	wire w_dff_A_jlMQbcnx0_0;
	wire w_dff_A_FI99FQIq5_0;
	wire w_dff_A_PY7d6QfG4_0;
	wire w_dff_A_MsWnJVJo1_0;
	wire w_dff_A_HlLZehqt3_0;
	wire w_dff_A_lpba5pzq6_0;
	wire w_dff_A_swV9s9Hu1_0;
	wire w_dff_A_isf6Pk4w8_0;
	wire w_dff_A_54BANchH9_0;
	wire w_dff_A_uBzSb6rx4_0;
	wire w_dff_A_gm0HgLDu1_0;
	wire w_dff_A_hcXpsd3A4_0;
	wire w_dff_A_JTFCEfen1_0;
	wire w_dff_A_IjNHmEwA4_0;
	wire w_dff_A_jtOqDm0C1_0;
	wire w_dff_A_QjAaaF7K9_0;
	wire w_dff_A_8GVQLnTP6_0;
	wire w_dff_A_Vjrix28J7_0;
	wire w_dff_A_cuvBx6Za0_0;
	wire w_dff_A_47q9H7HX8_0;
	wire w_dff_A_H6AhyeRT7_0;
	wire w_dff_A_PKpdpdsd9_0;
	wire w_dff_A_hD7rAjk38_0;
	wire w_dff_A_KthuUe4o7_0;
	wire w_dff_A_1IAF9V465_0;
	wire w_dff_A_rXU0VyyZ5_0;
	wire w_dff_A_WUe1CLaf3_0;
	wire w_dff_A_ngZ23UFr9_0;
	wire w_dff_A_Cc4exuqA1_0;
	wire w_dff_A_otkrwkU45_0;
	wire w_dff_A_dpU3uiMi9_0;
	wire w_dff_A_Lz5bU8Ya3_0;
	wire w_dff_A_KhCeDE7y0_0;
	wire w_dff_A_JE5APblT2_0;
	wire w_dff_A_3fHyx1Jv4_0;
	wire w_dff_A_9WSXcsoI9_0;
	wire w_dff_A_CrqKC3nq1_0;
	wire w_dff_A_CMHjCS0L6_0;
	wire w_dff_A_Ice4I31p7_0;
	wire w_dff_A_fpu40RXS1_0;
	wire w_dff_A_2GRSyJqq1_0;
	wire w_dff_A_vs4kgBu57_2;
	wire w_dff_A_vt4Y2m9N4_0;
	wire w_dff_A_tdJLxAiP5_0;
	wire w_dff_A_ysaXoF5z7_0;
	wire w_dff_A_yb9lUVjw4_0;
	wire w_dff_A_DZ3QFxdG1_0;
	wire w_dff_A_IKsb1xaL8_0;
	wire w_dff_A_X4Tjeb5v1_0;
	wire w_dff_A_LdUcYung7_0;
	wire w_dff_A_UcmHguER2_0;
	wire w_dff_A_72XggFCi2_0;
	wire w_dff_A_BDzujJga3_0;
	wire w_dff_A_Ws06adqW6_0;
	wire w_dff_A_8aQeNKaS1_0;
	wire w_dff_A_eej1nWK37_0;
	wire w_dff_A_3zS0AzMv2_0;
	wire w_dff_A_NpqL8I028_0;
	wire w_dff_A_wavaedhY7_0;
	wire w_dff_A_Rqw8Vh8i6_0;
	wire w_dff_A_WHQiO8fC0_0;
	wire w_dff_A_7uDrAlfu4_0;
	wire w_dff_A_qmfrpfF93_0;
	wire w_dff_A_KH2RYoTc0_0;
	wire w_dff_A_TyYzH7Uv2_0;
	wire w_dff_A_KfMod0ct7_0;
	wire w_dff_A_BVjaDU2z8_0;
	wire w_dff_A_umMVj3Sw2_0;
	wire w_dff_A_8XdyYXqr5_0;
	wire w_dff_A_FdIxDJKN6_0;
	wire w_dff_A_uAXBNBkM6_0;
	wire w_dff_A_XC0zWnLJ8_0;
	wire w_dff_A_u5SMg9nV2_0;
	wire w_dff_A_jKEUbQ1I1_0;
	wire w_dff_A_CDJ35Hec5_0;
	wire w_dff_A_lJ68NMyc3_0;
	wire w_dff_A_QVMWhmzb5_0;
	wire w_dff_A_oFYx4XUi9_0;
	wire w_dff_A_VzovCNYm7_0;
	wire w_dff_A_kUCaB2we9_0;
	wire w_dff_A_K0Ilz7YP0_0;
	wire w_dff_A_AlwT8s9K8_0;
	wire w_dff_A_8bn5XCZH8_0;
	wire w_dff_A_SJntTOgD2_0;
	wire w_dff_A_N7hK5Ywo5_0;
	wire w_dff_A_V1IkvfIo0_0;
	wire w_dff_A_C8vVumad3_0;
	wire w_dff_A_aB2V1atm8_0;
	wire w_dff_A_pIu8zC9C4_0;
	wire w_dff_A_1ItMPxZD5_0;
	wire w_dff_A_nFjwKY4e4_0;
	wire w_dff_A_7ylqROtw0_0;
	wire w_dff_A_vReCnBqg2_0;
	wire w_dff_A_wRKgzkYP8_0;
	wire w_dff_A_ykqs3oh58_0;
	wire w_dff_A_UBa2lvoL8_0;
	wire w_dff_A_f6GTBfjN3_0;
	wire w_dff_A_WpFZOaXU6_0;
	wire w_dff_A_R1PDDnD57_0;
	wire w_dff_A_yuUlPWbi8_0;
	wire w_dff_A_oPpAL3Eb8_0;
	wire w_dff_A_YOEyE2Ft4_0;
	wire w_dff_A_ymDkE7QA9_0;
	wire w_dff_A_PcpGoIOS7_0;
	wire w_dff_A_GVHM0wzS0_0;
	wire w_dff_A_DPLpEJdk3_0;
	wire w_dff_A_h4nhCUpe5_0;
	wire w_dff_A_jFUWWvbN5_0;
	wire w_dff_A_X2qNxCpV7_0;
	wire w_dff_A_ot49Qtx87_0;
	wire w_dff_A_D1J7lZ8S1_2;
	wire w_dff_A_5VdlFGQX8_0;
	wire w_dff_A_11uqXQUt4_0;
	wire w_dff_A_z0hbwh0k0_0;
	wire w_dff_A_5Ea3pvvn7_0;
	wire w_dff_A_3MSpyuVM9_0;
	wire w_dff_A_NPlD3U850_0;
	wire w_dff_A_aY6hHetZ2_0;
	wire w_dff_A_AYeoMJMa5_0;
	wire w_dff_A_DOvmNg326_0;
	wire w_dff_A_KIgKS7ex0_0;
	wire w_dff_A_dPOfIh3R4_0;
	wire w_dff_A_xxd3ghpm2_0;
	wire w_dff_A_4fX1ZjQL2_0;
	wire w_dff_A_9pAvsRqz4_0;
	wire w_dff_A_x6XmJUgp0_0;
	wire w_dff_A_gu6RG1KW0_0;
	wire w_dff_A_XcB9VRBe6_0;
	wire w_dff_A_SiOvmyOY5_0;
	wire w_dff_A_N8pYPSn50_0;
	wire w_dff_A_yjZxB4u51_0;
	wire w_dff_A_7kkk1XYh7_0;
	wire w_dff_A_IHH1p1JI5_0;
	wire w_dff_A_LziHCwwI2_0;
	wire w_dff_A_VQMpyaCL4_0;
	wire w_dff_A_qZ43ZVAg2_0;
	wire w_dff_A_ia4uFhAI3_0;
	wire w_dff_A_JBgWHlnm6_0;
	wire w_dff_A_jrHgQmEH5_0;
	wire w_dff_A_Ol8FOpdB8_0;
	wire w_dff_A_Ipo92fHW3_0;
	wire w_dff_A_XnBgPrZf6_0;
	wire w_dff_A_qGfGdB2L8_0;
	wire w_dff_A_MwnirlbD0_0;
	wire w_dff_A_ZFFw6czc6_0;
	wire w_dff_A_m4Ze4Ssf3_0;
	wire w_dff_A_ATdCIE9I0_0;
	wire w_dff_A_mTZKJUhg0_0;
	wire w_dff_A_1ylxeht97_0;
	wire w_dff_A_11aitGHD7_0;
	wire w_dff_A_NhXWoq7n7_0;
	wire w_dff_A_jGAapAjR2_0;
	wire w_dff_A_R34ICqlN3_0;
	wire w_dff_A_56vmJzb38_0;
	wire w_dff_A_floHRrHw9_0;
	wire w_dff_A_a6CXb8Ng1_0;
	wire w_dff_A_UYKcMncX9_0;
	wire w_dff_A_WRmRh7vK6_0;
	wire w_dff_A_ATRCgMXG2_0;
	wire w_dff_A_g6OSqU0P0_0;
	wire w_dff_A_4mTXAxGe0_0;
	wire w_dff_A_BvAqLBDM8_0;
	wire w_dff_A_vd4bv5001_0;
	wire w_dff_A_RDzJZCix4_0;
	wire w_dff_A_sZKMNCFf6_0;
	wire w_dff_A_rgER3r5x9_0;
	wire w_dff_A_CQLc17Wd1_0;
	wire w_dff_A_agLNOFAh4_0;
	wire w_dff_A_auIuwebJ2_0;
	wire w_dff_A_NjVTGFQ62_0;
	wire w_dff_A_Vzs7Oa837_0;
	wire w_dff_A_7D3sDAAy3_0;
	wire w_dff_A_9gn8rMLL5_0;
	wire w_dff_A_nWwozueN8_0;
	wire w_dff_A_TmBQdEiT0_0;
	wire w_dff_A_C7GbskCZ8_0;
	wire w_dff_A_PldpzvGS2_2;
	wire w_dff_A_QaN4hjlH1_0;
	wire w_dff_A_ux1XDO1D5_0;
	wire w_dff_A_VVd3iCVb6_0;
	wire w_dff_A_BiukFx9j7_0;
	wire w_dff_A_PDAsfrc99_0;
	wire w_dff_A_GSIKqZTW5_0;
	wire w_dff_A_dIJmV9rb3_0;
	wire w_dff_A_cwgYcYzE4_0;
	wire w_dff_A_hOtfK5E33_0;
	wire w_dff_A_1pHepJP47_0;
	wire w_dff_A_BpE9rstO0_0;
	wire w_dff_A_QXxbKmvC7_0;
	wire w_dff_A_U2ceAQvx6_0;
	wire w_dff_A_TK3rNgCK0_0;
	wire w_dff_A_EMGVVePw8_0;
	wire w_dff_A_WTfNUG740_0;
	wire w_dff_A_HHJvtuQG2_0;
	wire w_dff_A_1AZotT3V1_0;
	wire w_dff_A_uZp04kMa4_0;
	wire w_dff_A_2Qd176o97_0;
	wire w_dff_A_Pg0ws8P03_0;
	wire w_dff_A_98A75F9Z1_0;
	wire w_dff_A_zKruO8ht1_0;
	wire w_dff_A_vvt1aiZm5_0;
	wire w_dff_A_I1tgTuJy7_0;
	wire w_dff_A_y0RZYSPV7_0;
	wire w_dff_A_jxl0YOe47_0;
	wire w_dff_A_4k0oDl9z6_0;
	wire w_dff_A_tNSDqPDw4_0;
	wire w_dff_A_D1MbQm2I7_0;
	wire w_dff_A_PIlN1MBS3_0;
	wire w_dff_A_8CeeJWxV9_0;
	wire w_dff_A_9hxGB0Dr6_0;
	wire w_dff_A_7j24TzSO2_0;
	wire w_dff_A_ZrqnpYrO6_0;
	wire w_dff_A_NUuKzZNk9_0;
	wire w_dff_A_1osgNuPS4_0;
	wire w_dff_A_XtUBurmn0_0;
	wire w_dff_A_nCOAkcvA3_0;
	wire w_dff_A_OfAwnrYR2_0;
	wire w_dff_A_OfdBXbLF8_0;
	wire w_dff_A_eH0MGLK35_0;
	wire w_dff_A_whbKx2wh6_0;
	wire w_dff_A_5RoUYWqt7_0;
	wire w_dff_A_MfljODPt6_0;
	wire w_dff_A_Mv7MkqSf1_0;
	wire w_dff_A_spk3HlPx2_0;
	wire w_dff_A_59u8j0E63_0;
	wire w_dff_A_FsmbLvpH8_0;
	wire w_dff_A_T2n6wKPW0_0;
	wire w_dff_A_Jh2YMt7n6_0;
	wire w_dff_A_w9IxogiP3_0;
	wire w_dff_A_x22pA9Dg2_0;
	wire w_dff_A_Nn3xoHwg4_0;
	wire w_dff_A_iOplehm90_0;
	wire w_dff_A_SzGz9iH07_0;
	wire w_dff_A_wjnyXDYZ8_0;
	wire w_dff_A_lgjC48jg0_0;
	wire w_dff_A_ivBOeMVc6_0;
	wire w_dff_A_Su5wLHVe0_0;
	wire w_dff_A_B3yINSX60_0;
	wire w_dff_A_W3AJC9D04_0;
	wire w_dff_A_YL90IabU6_2;
	wire w_dff_A_hSbn9xYI2_0;
	wire w_dff_A_CVqIS5yc9_0;
	wire w_dff_A_8s2g5Me99_0;
	wire w_dff_A_TC7gfXnH7_0;
	wire w_dff_A_JjI8d8YY3_0;
	wire w_dff_A_etQJDmiQ9_0;
	wire w_dff_A_NbObjnJx2_0;
	wire w_dff_A_Up1xVSlF6_0;
	wire w_dff_A_dbZUezcG7_0;
	wire w_dff_A_EdVkP9cB3_0;
	wire w_dff_A_uDtCIdfn4_0;
	wire w_dff_A_cjIiqBUC8_0;
	wire w_dff_A_rjrB2rRP7_0;
	wire w_dff_A_pPMhbB8H3_0;
	wire w_dff_A_yVEumW7h3_0;
	wire w_dff_A_LYwKI1nT2_0;
	wire w_dff_A_DFMR8NpH6_0;
	wire w_dff_A_n3H0GgbP7_0;
	wire w_dff_A_WEIjJbIZ9_0;
	wire w_dff_A_bJL5Zpll8_0;
	wire w_dff_A_QvRfJ2HN2_0;
	wire w_dff_A_W6CIbonm3_0;
	wire w_dff_A_DoZteobw0_0;
	wire w_dff_A_7B6PW1H97_0;
	wire w_dff_A_Glb9PYKR3_0;
	wire w_dff_A_SWu8MAQi4_0;
	wire w_dff_A_ik55kIAn4_0;
	wire w_dff_A_OA7tcb1Q1_0;
	wire w_dff_A_Pp6EtWCg9_0;
	wire w_dff_A_JOacAFEL0_0;
	wire w_dff_A_taAlJBcR7_0;
	wire w_dff_A_FlVssQCe7_0;
	wire w_dff_A_okKLQTvm0_0;
	wire w_dff_A_8nvJZ0Vo1_0;
	wire w_dff_A_XsgQDMbk5_0;
	wire w_dff_A_F6EzjnPa6_0;
	wire w_dff_A_nDBPpSMl6_0;
	wire w_dff_A_n6jdrTl05_0;
	wire w_dff_A_2AYU47VH7_0;
	wire w_dff_A_lITkqGhi2_0;
	wire w_dff_A_mPJxec0m8_0;
	wire w_dff_A_PydP6ym81_0;
	wire w_dff_A_7B3GncZN1_0;
	wire w_dff_A_lUPKBMOB1_0;
	wire w_dff_A_71TYRVaG3_0;
	wire w_dff_A_Vr0tPljX2_0;
	wire w_dff_A_D7G1jR538_0;
	wire w_dff_A_zcL5PmoR3_0;
	wire w_dff_A_KQUOWqSc1_0;
	wire w_dff_A_KMp0WJip0_0;
	wire w_dff_A_3y1YA1Oa6_0;
	wire w_dff_A_ly3ySnyv7_0;
	wire w_dff_A_WXDRqHZG4_0;
	wire w_dff_A_msLZBPmv9_0;
	wire w_dff_A_P1l6Dv7z1_0;
	wire w_dff_A_gzUGqGrS0_0;
	wire w_dff_A_kv8RO6a14_0;
	wire w_dff_A_p1jXc0CU5_0;
	wire w_dff_A_3pnN2caj1_0;
	wire w_dff_A_ML3PYmGw6_2;
	wire w_dff_A_k3hbTgbw1_0;
	wire w_dff_A_7gMWKem29_0;
	wire w_dff_A_OVagVgzt8_0;
	wire w_dff_A_EQk1N8XE8_0;
	wire w_dff_A_o5UxAA9t6_0;
	wire w_dff_A_4owISbqM2_0;
	wire w_dff_A_ifry3w2J0_0;
	wire w_dff_A_19QwWR2D4_0;
	wire w_dff_A_Sz3kEFaI4_0;
	wire w_dff_A_8sPxZoJ60_0;
	wire w_dff_A_OCHEaoC98_0;
	wire w_dff_A_H6QVTEWY3_0;
	wire w_dff_A_zaog7Hqm6_0;
	wire w_dff_A_IJpfjMiy3_0;
	wire w_dff_A_DUwSHHoa4_0;
	wire w_dff_A_ry5I9gVV6_0;
	wire w_dff_A_COyi6Itd1_0;
	wire w_dff_A_yiq7gymJ9_0;
	wire w_dff_A_eZsxtNCc5_0;
	wire w_dff_A_ocRW2mOu0_0;
	wire w_dff_A_f0w3GwGQ1_0;
	wire w_dff_A_NdPr0yb54_0;
	wire w_dff_A_wm2ibPjd5_0;
	wire w_dff_A_h9W6Xg6G7_0;
	wire w_dff_A_P5ZI6iMN3_0;
	wire w_dff_A_t2s8Yrtq2_0;
	wire w_dff_A_1nzIiqnE1_0;
	wire w_dff_A_d4HTecqI3_0;
	wire w_dff_A_fk4qrDBu0_0;
	wire w_dff_A_ox2hGdUL6_0;
	wire w_dff_A_VnKYrr3r1_0;
	wire w_dff_A_v7AsgOaS8_0;
	wire w_dff_A_J0SWVODD8_0;
	wire w_dff_A_VjGxIN4R5_0;
	wire w_dff_A_8jbEMAUT0_0;
	wire w_dff_A_59W2UrYY3_0;
	wire w_dff_A_bMnUCCrQ0_0;
	wire w_dff_A_kKZM6Pi90_0;
	wire w_dff_A_CgrReBRv0_0;
	wire w_dff_A_7Icgqo6H8_0;
	wire w_dff_A_iNriN8iw9_0;
	wire w_dff_A_9hdkHlNi4_0;
	wire w_dff_A_Ok6iiI9m3_0;
	wire w_dff_A_wI49MFMv7_0;
	wire w_dff_A_A47xoUlP6_0;
	wire w_dff_A_asAKRf9w1_0;
	wire w_dff_A_XtuG2nkg8_0;
	wire w_dff_A_kTzuItIH0_0;
	wire w_dff_A_kcLgxgPP7_0;
	wire w_dff_A_4HfSNL7E7_0;
	wire w_dff_A_bhTdnMuf2_0;
	wire w_dff_A_mV8wK1155_0;
	wire w_dff_A_ePVaFnM57_0;
	wire w_dff_A_SpgU20S39_0;
	wire w_dff_A_GPpo5IbF2_0;
	wire w_dff_A_F81vDXYA9_0;
	wire w_dff_A_p8CWdcT47_2;
	wire w_dff_A_vIN3fXLZ2_0;
	wire w_dff_A_murdQeTr3_0;
	wire w_dff_A_qyRBVjgt4_0;
	wire w_dff_A_UWdhPYhA8_0;
	wire w_dff_A_Zc4eXUwU6_0;
	wire w_dff_A_Mc8Wha1q2_0;
	wire w_dff_A_VsphuY9H5_0;
	wire w_dff_A_HX2q0STK3_0;
	wire w_dff_A_8mvjjQ8w0_0;
	wire w_dff_A_bqESm2l63_0;
	wire w_dff_A_5Nl4WnvC9_0;
	wire w_dff_A_ykxwu6cd3_0;
	wire w_dff_A_lhpgddm69_0;
	wire w_dff_A_CWkLmZ9f6_0;
	wire w_dff_A_a0rjBk531_0;
	wire w_dff_A_2iedVuis6_0;
	wire w_dff_A_2GNJRJN49_0;
	wire w_dff_A_ENcapxbA2_0;
	wire w_dff_A_E7uQrMF42_0;
	wire w_dff_A_3xiSwC5F9_0;
	wire w_dff_A_svNWcnZz2_0;
	wire w_dff_A_6rhR35bC2_0;
	wire w_dff_A_n736qRW58_0;
	wire w_dff_A_9ixB6Oj44_0;
	wire w_dff_A_TSPdbDcl6_0;
	wire w_dff_A_EOI67Sd87_0;
	wire w_dff_A_BSHQMDeF5_0;
	wire w_dff_A_dku6XVqK9_0;
	wire w_dff_A_4IISccVA9_0;
	wire w_dff_A_vCWreVNQ1_0;
	wire w_dff_A_7blmHrjB1_0;
	wire w_dff_A_a6ZhVuG86_0;
	wire w_dff_A_WmshASpB0_0;
	wire w_dff_A_eviCvvc00_0;
	wire w_dff_A_vvNLWVY49_0;
	wire w_dff_A_2uH30iFi9_0;
	wire w_dff_A_73Jy1lAO5_0;
	wire w_dff_A_IWyQhmTp6_0;
	wire w_dff_A_QGZRqCOG2_0;
	wire w_dff_A_O2pv5VvY8_0;
	wire w_dff_A_5kDnpyuh7_0;
	wire w_dff_A_4bAvnC9u7_0;
	wire w_dff_A_CSfaVj1b3_0;
	wire w_dff_A_j2OmXIcK8_0;
	wire w_dff_A_nSO9w3xe7_0;
	wire w_dff_A_uzzkA84e1_0;
	wire w_dff_A_1EyFcUot8_0;
	wire w_dff_A_wMQ1QNGZ9_0;
	wire w_dff_A_BA22Zhw80_0;
	wire w_dff_A_qM72JduN4_0;
	wire w_dff_A_0iRaUxIe4_0;
	wire w_dff_A_c7RE4A0A9_0;
	wire w_dff_A_5JwUzXPA2_0;
	wire w_dff_A_aV8fpFrx0_2;
	wire w_dff_A_0U1eS1Nh1_0;
	wire w_dff_A_XciRZcPX6_0;
	wire w_dff_A_dNsXdzoD6_0;
	wire w_dff_A_DF4r45PI4_0;
	wire w_dff_A_6ib9vVbp3_0;
	wire w_dff_A_QbC4MRD40_0;
	wire w_dff_A_rllvemIL9_0;
	wire w_dff_A_cmiqokas9_0;
	wire w_dff_A_0aT3jov38_0;
	wire w_dff_A_Xjz9riNF7_0;
	wire w_dff_A_wZ7XgEnk5_0;
	wire w_dff_A_jvj58AaU0_0;
	wire w_dff_A_WGrBtmzJ3_0;
	wire w_dff_A_qrnMsTzN6_0;
	wire w_dff_A_IXZ4RphD5_0;
	wire w_dff_A_nDQT0Bqm9_0;
	wire w_dff_A_7DxEEq538_0;
	wire w_dff_A_VMbF0QFq1_0;
	wire w_dff_A_0h7Rnq0j9_0;
	wire w_dff_A_tObv25cz7_0;
	wire w_dff_A_edY2CSKo7_0;
	wire w_dff_A_rcOxops84_0;
	wire w_dff_A_1XIZFMrL2_0;
	wire w_dff_A_DecREavl0_0;
	wire w_dff_A_ZnuiK6Me8_0;
	wire w_dff_A_V9Z3Fxt27_0;
	wire w_dff_A_XGxsuKCA0_0;
	wire w_dff_A_jSFjKJnA5_0;
	wire w_dff_A_OBHTPb8G3_0;
	wire w_dff_A_hrMPtjRC3_0;
	wire w_dff_A_BEbtPiKp7_0;
	wire w_dff_A_fuPxVhmE3_0;
	wire w_dff_A_sxaPDRBN3_0;
	wire w_dff_A_FIHiv3Lw1_0;
	wire w_dff_A_nYZZPLxt4_0;
	wire w_dff_A_HKSJ8cgS3_0;
	wire w_dff_A_oefFO2oq7_0;
	wire w_dff_A_kywkKTac8_0;
	wire w_dff_A_u6LAQU9n0_0;
	wire w_dff_A_qyUEWSpa9_0;
	wire w_dff_A_nVfuuVEZ5_0;
	wire w_dff_A_y3Mg9dp28_0;
	wire w_dff_A_EJNd4H0Z3_0;
	wire w_dff_A_MvZc0U2H5_0;
	wire w_dff_A_R8zNVeUO6_0;
	wire w_dff_A_S69efoHJ6_0;
	wire w_dff_A_vYthnCn77_0;
	wire w_dff_A_dRhvuoNw9_0;
	wire w_dff_A_nk5z5N5r8_0;
	wire w_dff_A_9vRoFg8j0_0;
	wire w_dff_A_xLPUpw6m3_2;
	wire w_dff_A_QK12NJAC1_0;
	wire w_dff_A_QcGeXnrj0_0;
	wire w_dff_A_odvBaEmS8_0;
	wire w_dff_A_78ghDAb57_0;
	wire w_dff_A_OQNNHVWy1_0;
	wire w_dff_A_GMTVX1TR2_0;
	wire w_dff_A_f5UPQVK13_0;
	wire w_dff_A_DcUF1SkU7_0;
	wire w_dff_A_UtNgAUgX5_0;
	wire w_dff_A_khITjU2X8_0;
	wire w_dff_A_i0QThDGl5_0;
	wire w_dff_A_Y6p5te3r2_0;
	wire w_dff_A_dMnp0QqG2_0;
	wire w_dff_A_3em5remO9_0;
	wire w_dff_A_7GrAzDZs5_0;
	wire w_dff_A_Q0WNY1Xl4_0;
	wire w_dff_A_JL52Oqix5_0;
	wire w_dff_A_nuzg1xGW4_0;
	wire w_dff_A_RCarGdSy2_0;
	wire w_dff_A_K5rHSPpA1_0;
	wire w_dff_A_HHMFfhmR4_0;
	wire w_dff_A_S6AS7W723_0;
	wire w_dff_A_zZNXjYWQ1_0;
	wire w_dff_A_0Pawiz2H8_0;
	wire w_dff_A_ZOqTnZRI1_0;
	wire w_dff_A_frzqTFQU7_0;
	wire w_dff_A_ztZV15So3_0;
	wire w_dff_A_zRR3ME1v8_0;
	wire w_dff_A_YlS9cwIT6_0;
	wire w_dff_A_RtBY4bb97_0;
	wire w_dff_A_CVak30a55_0;
	wire w_dff_A_AwjAA4Kz2_0;
	wire w_dff_A_q6EBBycg5_0;
	wire w_dff_A_YQ6ZgHCP2_0;
	wire w_dff_A_l6TnnlmD7_0;
	wire w_dff_A_zLhYjaVg5_0;
	wire w_dff_A_r6EIwhAa1_0;
	wire w_dff_A_XYCROZpX6_0;
	wire w_dff_A_3n2ABVn97_0;
	wire w_dff_A_N2Jlv2Hl5_0;
	wire w_dff_A_1xRXt6jg0_0;
	wire w_dff_A_N3chEZbv8_0;
	wire w_dff_A_5XDC8Sma9_0;
	wire w_dff_A_9pOJfBB00_0;
	wire w_dff_A_APiTgBJb5_0;
	wire w_dff_A_ZVkuoleY1_0;
	wire w_dff_A_GgZyM2mP0_0;
	wire w_dff_A_0FjbwSqr7_2;
	wire w_dff_A_v2NlOv3r7_0;
	wire w_dff_A_vXtYIMoI8_0;
	wire w_dff_A_fWjPS95U8_0;
	wire w_dff_A_shWmwZ4i6_0;
	wire w_dff_A_vAk4AwuO0_0;
	wire w_dff_A_j3ZrDR6t3_0;
	wire w_dff_A_Ovwf8QUQ8_0;
	wire w_dff_A_Nf3Q58to4_0;
	wire w_dff_A_UrFSKH9n3_0;
	wire w_dff_A_BURDr2196_0;
	wire w_dff_A_ujZTwe5P2_0;
	wire w_dff_A_ugvHRZPQ8_0;
	wire w_dff_A_ptqPrW0t5_0;
	wire w_dff_A_D3V15u9R0_0;
	wire w_dff_A_10xftJvC4_0;
	wire w_dff_A_3jvctEhx4_0;
	wire w_dff_A_Sd4w4de37_0;
	wire w_dff_A_SUDhWvOt1_0;
	wire w_dff_A_ACkv5MI83_0;
	wire w_dff_A_AkXJFaCi0_0;
	wire w_dff_A_DcwAzE9I1_0;
	wire w_dff_A_BjJMKzPh1_0;
	wire w_dff_A_Wri9CrDy5_0;
	wire w_dff_A_fPcFWY5b5_0;
	wire w_dff_A_xf7iYQEE1_0;
	wire w_dff_A_hJst8t655_0;
	wire w_dff_A_66b8KN7Z9_0;
	wire w_dff_A_pfcZH3Ke6_0;
	wire w_dff_A_vdcsjvKF9_0;
	wire w_dff_A_QBNhy4Oo8_0;
	wire w_dff_A_i518BMWU1_0;
	wire w_dff_A_eGRyYK2v9_0;
	wire w_dff_A_RBsEs5yg9_0;
	wire w_dff_A_gxPcKutd1_0;
	wire w_dff_A_y5PqvIz20_0;
	wire w_dff_A_ZXblgs8T7_0;
	wire w_dff_A_MA85Bv5N4_0;
	wire w_dff_A_2Bp2y0Eh2_0;
	wire w_dff_A_pNyLUNaN5_0;
	wire w_dff_A_ifPUox836_0;
	wire w_dff_A_Vl8klQJT9_0;
	wire w_dff_A_PjwROmtr7_0;
	wire w_dff_A_5jvpmlY93_0;
	wire w_dff_A_2zTuU5tl4_0;
	wire w_dff_A_TjdGLRLw9_2;
	wire w_dff_A_a6dW4Wnh8_0;
	wire w_dff_A_NpRxMuo52_0;
	wire w_dff_A_c6flYkow7_0;
	wire w_dff_A_sCc4a96U6_0;
	wire w_dff_A_AwwDDlC17_0;
	wire w_dff_A_CiHco9fX7_0;
	wire w_dff_A_NzwOd8pu2_0;
	wire w_dff_A_Z41jJ2T81_0;
	wire w_dff_A_wWAq8bYL9_0;
	wire w_dff_A_1I6dMjJc0_0;
	wire w_dff_A_jGxsFTrn7_0;
	wire w_dff_A_y5wssT002_0;
	wire w_dff_A_vphPzTZF8_0;
	wire w_dff_A_Dg5TWWQc3_0;
	wire w_dff_A_Hjs7E3516_0;
	wire w_dff_A_r2bio3nM9_0;
	wire w_dff_A_FL9yVWlF8_0;
	wire w_dff_A_8R3uGzBw0_0;
	wire w_dff_A_tk7jAMRt0_0;
	wire w_dff_A_ADSz6GLN9_0;
	wire w_dff_A_e6UcSutJ9_0;
	wire w_dff_A_SQ0a9nQC3_0;
	wire w_dff_A_9nhDXwj06_0;
	wire w_dff_A_Md4bjF6Z9_0;
	wire w_dff_A_yMqzClJm9_0;
	wire w_dff_A_P2YcLkYv7_0;
	wire w_dff_A_wDcNvaE75_0;
	wire w_dff_A_zEjC8w5T5_0;
	wire w_dff_A_9NlEIUAy3_0;
	wire w_dff_A_SxsaFq6y8_0;
	wire w_dff_A_Bp11NYbI2_0;
	wire w_dff_A_1KgPX6CE6_0;
	wire w_dff_A_0ZrandTC4_0;
	wire w_dff_A_7bRrsiQk5_0;
	wire w_dff_A_SJq5fYCH5_0;
	wire w_dff_A_gvGWBQZQ6_0;
	wire w_dff_A_e7Ks6Wl86_0;
	wire w_dff_A_BZDT2QZj6_0;
	wire w_dff_A_0UNyN9CL2_0;
	wire w_dff_A_u4mEd3e62_0;
	wire w_dff_A_p1R9qLD41_0;
	wire w_dff_A_n39HOqln6_2;
	wire w_dff_A_PXYOGhAB5_0;
	wire w_dff_A_ccvQQc4W1_0;
	wire w_dff_A_v3OSxPsP3_0;
	wire w_dff_A_KrXAkzbj4_0;
	wire w_dff_A_QnyWjelI2_0;
	wire w_dff_A_cQwWQltv2_0;
	wire w_dff_A_JMQ0IoUh4_0;
	wire w_dff_A_DGbuDETQ3_0;
	wire w_dff_A_MGG4IEfF1_0;
	wire w_dff_A_KeSUoF4c3_0;
	wire w_dff_A_XUReLZzE0_0;
	wire w_dff_A_I3tK6U1N1_0;
	wire w_dff_A_GuwBZFwr8_0;
	wire w_dff_A_9eXdsHEP1_0;
	wire w_dff_A_UMpSS8Q03_0;
	wire w_dff_A_Pp0sLBA62_0;
	wire w_dff_A_skNgviXu7_0;
	wire w_dff_A_xTBEM8Fr0_0;
	wire w_dff_A_ysDfatWY2_0;
	wire w_dff_A_sIBXIBgh7_0;
	wire w_dff_A_D0BStk2N7_0;
	wire w_dff_A_O6fynBIh5_0;
	wire w_dff_A_ZrEvEVVm9_0;
	wire w_dff_A_KrVUD9wZ5_0;
	wire w_dff_A_3rmwHDer8_0;
	wire w_dff_A_ZM4Q09M85_0;
	wire w_dff_A_RLjrw6mG7_0;
	wire w_dff_A_7viF9eR54_0;
	wire w_dff_A_dQrwwRV21_0;
	wire w_dff_A_Oc7eU37c1_0;
	wire w_dff_A_TjjslqyG7_0;
	wire w_dff_A_s4eG32rq3_0;
	wire w_dff_A_tgEVvcUC2_0;
	wire w_dff_A_TojyohDe3_0;
	wire w_dff_A_bjCIdwKR9_0;
	wire w_dff_A_XPmKIEMU6_0;
	wire w_dff_A_eEbg3W3c2_0;
	wire w_dff_A_UmDYDhTC6_0;
	wire w_dff_A_WSl0EIyE8_2;
	wire w_dff_A_xitS8AkT0_0;
	wire w_dff_A_BSxvz88n7_0;
	wire w_dff_A_LSoJSI6f1_0;
	wire w_dff_A_DGL0CW8y4_0;
	wire w_dff_A_oTDyi2rv0_0;
	wire w_dff_A_Y4euN9vd1_0;
	wire w_dff_A_INVqkSpx5_0;
	wire w_dff_A_f2eq9Zt65_0;
	wire w_dff_A_lqJ6VHIA4_0;
	wire w_dff_A_a7SqyRw98_0;
	wire w_dff_A_N0SmX26K4_0;
	wire w_dff_A_BVmziCF87_0;
	wire w_dff_A_wRb2ybTo8_0;
	wire w_dff_A_HBEf2gIx4_0;
	wire w_dff_A_x3jQrAfc2_0;
	wire w_dff_A_RYrsZBUM6_0;
	wire w_dff_A_qKJwP7Kc2_0;
	wire w_dff_A_OrKjtW3x1_0;
	wire w_dff_A_A9mUCM720_0;
	wire w_dff_A_QmJ8Ul4Y6_0;
	wire w_dff_A_T9F5kV4w5_0;
	wire w_dff_A_4aa6IcZh6_0;
	wire w_dff_A_86YsFzoF3_0;
	wire w_dff_A_RvU0rqpO0_0;
	wire w_dff_A_zREhpBw31_0;
	wire w_dff_A_7yGCrpIi9_0;
	wire w_dff_A_L3I894qR8_0;
	wire w_dff_A_6FNDU8F08_0;
	wire w_dff_A_JZbZCbVK2_0;
	wire w_dff_A_lZbtv4Dn2_0;
	wire w_dff_A_xjQqyAC48_0;
	wire w_dff_A_NXVTaOIn1_0;
	wire w_dff_A_Arr6ZWbq3_0;
	wire w_dff_A_UEa5lEg98_0;
	wire w_dff_A_AgN3q7uf2_0;
	wire w_dff_A_ZhxLR9C13_2;
	wire w_dff_A_9WX7sZQQ7_0;
	wire w_dff_A_Ba3QuFnW3_0;
	wire w_dff_A_kWVBo9Cp2_0;
	wire w_dff_A_lqVv0DfJ7_0;
	wire w_dff_A_ZeDiL4Ar9_0;
	wire w_dff_A_JMvNQLNs0_0;
	wire w_dff_A_MzjB351A9_0;
	wire w_dff_A_CpuYyrwR5_0;
	wire w_dff_A_v7UpYvVh4_0;
	wire w_dff_A_YOXKoh117_0;
	wire w_dff_A_C6uF63eD0_0;
	wire w_dff_A_wvJpvDsk0_0;
	wire w_dff_A_dwkQyt1l6_0;
	wire w_dff_A_StsFwRK94_0;
	wire w_dff_A_njdFfX3w3_0;
	wire w_dff_A_Ozixgr5S6_0;
	wire w_dff_A_nG3rHP5V2_0;
	wire w_dff_A_ZJdGLJYx9_0;
	wire w_dff_A_clh1lQBc8_0;
	wire w_dff_A_B1DojI7m5_0;
	wire w_dff_A_zOwrnuid2_0;
	wire w_dff_A_TRer6PZN2_0;
	wire w_dff_A_F5ym6srX2_0;
	wire w_dff_A_SxJqZXzi3_0;
	wire w_dff_A_hmBfOyWc5_0;
	wire w_dff_A_xIqKHLJc8_0;
	wire w_dff_A_EAKZ0q5X5_0;
	wire w_dff_A_Rc7ncFnQ7_0;
	wire w_dff_A_qJOfDy521_0;
	wire w_dff_A_pzyh0SBC4_0;
	wire w_dff_A_XtjlzGCk4_0;
	wire w_dff_A_32zRcKXp9_0;
	wire w_dff_A_RiGNgq0v5_2;
	wire w_dff_A_BRaODm1z6_0;
	wire w_dff_A_y6YdgwjN3_0;
	wire w_dff_A_sA3CfVXX8_0;
	wire w_dff_A_nMnbmvvI1_0;
	wire w_dff_A_sQlvJgaY8_0;
	wire w_dff_A_uoPjVtxN1_0;
	wire w_dff_A_7yrMR0ab4_0;
	wire w_dff_A_VTEG6IL61_0;
	wire w_dff_A_4Uxi5dxr4_0;
	wire w_dff_A_YeTiCmJM6_0;
	wire w_dff_A_XEOHnWHI5_0;
	wire w_dff_A_mYFAKh8B8_0;
	wire w_dff_A_2Rl10XbI4_0;
	wire w_dff_A_8PSniu2M8_0;
	wire w_dff_A_WvLuzetH5_0;
	wire w_dff_A_7rhpeM8U9_0;
	wire w_dff_A_H6GXloK48_0;
	wire w_dff_A_m2SXRMYS6_0;
	wire w_dff_A_dP2cDpOZ9_0;
	wire w_dff_A_Ziz6r9ml4_0;
	wire w_dff_A_f8EEHrxG9_0;
	wire w_dff_A_IoTughCQ0_0;
	wire w_dff_A_akKqVMdM8_0;
	wire w_dff_A_pMCnnbfu9_0;
	wire w_dff_A_CWhxHb8s9_0;
	wire w_dff_A_i6BPHUvn5_0;
	wire w_dff_A_B2W53vBp3_0;
	wire w_dff_A_AjyUEPaL0_0;
	wire w_dff_A_4BgyMPAM4_0;
	wire w_dff_A_YCRvBVIi5_2;
	wire w_dff_A_HhMXcIse2_0;
	wire w_dff_A_k2PgIPBi0_0;
	wire w_dff_A_wJHW178i5_0;
	wire w_dff_A_KtLN4ZB32_0;
	wire w_dff_A_3ikgKnXR2_0;
	wire w_dff_A_UyHNsjUb8_0;
	wire w_dff_A_7S8vQGny7_0;
	wire w_dff_A_uqCEpxMI5_0;
	wire w_dff_A_Tlcq6KGg6_0;
	wire w_dff_A_vKU23z184_0;
	wire w_dff_A_IgztpfZa8_0;
	wire w_dff_A_uoBjILui7_0;
	wire w_dff_A_Cb9Hg85J4_0;
	wire w_dff_A_6akwj2CO0_0;
	wire w_dff_A_bS45ZKch5_0;
	wire w_dff_A_5dZKLWRO0_0;
	wire w_dff_A_3e9fCXZc2_0;
	wire w_dff_A_EH0zUNSa3_0;
	wire w_dff_A_jsneHnAm8_0;
	wire w_dff_A_sjZouKhD0_0;
	wire w_dff_A_4cBQzAk47_0;
	wire w_dff_A_9HaDc8zY5_0;
	wire w_dff_A_EQhHENGU5_0;
	wire w_dff_A_cHkLUQnw4_0;
	wire w_dff_A_4hAR9USW3_0;
	wire w_dff_A_ZJWPtwWd1_0;
	wire w_dff_A_cO1UaNWW3_0;
	wire w_dff_A_3j1PEYfK3_2;
	wire w_dff_A_sO9qh7Ax4_0;
	wire w_dff_A_GhHGmgVn7_0;
	wire w_dff_A_BrBtDBV98_0;
	wire w_dff_A_j3J5GqAj0_0;
	wire w_dff_A_av1uvVys2_0;
	wire w_dff_A_XaX95qps8_0;
	wire w_dff_A_mktdfFWU4_0;
	wire w_dff_A_kr2eQAx83_0;
	wire w_dff_A_BLsqHu6k6_0;
	wire w_dff_A_c6yqcFoO5_0;
	wire w_dff_A_khXknZXq3_0;
	wire w_dff_A_DEbtyCtf3_0;
	wire w_dff_A_h7t1cluU1_0;
	wire w_dff_A_jPpR8efA0_0;
	wire w_dff_A_rFk65SJ82_0;
	wire w_dff_A_wjJBQDJX9_0;
	wire w_dff_A_25khai6V3_0;
	wire w_dff_A_kQdSDMHx2_0;
	wire w_dff_A_TKnrswjf5_0;
	wire w_dff_A_k0T0mM0J9_0;
	wire w_dff_A_3ltsmNx67_0;
	wire w_dff_A_Z9Ci4EUj9_0;
	wire w_dff_A_SBKcqrin0_0;
	wire w_dff_A_tfMGGzxj6_0;
	wire w_dff_A_Se8Tumc06_0;
	wire w_dff_A_qleo09kn4_2;
	wire w_dff_A_lCBBv9QO2_0;
	wire w_dff_A_TtyIYZh40_0;
	wire w_dff_A_RfM33e8G2_0;
	wire w_dff_A_LWO1MQ7j5_0;
	wire w_dff_A_VlMxCanH3_0;
	wire w_dff_A_s1UldOVh1_0;
	wire w_dff_A_7EA0wUEj3_0;
	wire w_dff_A_XRwueToC5_0;
	wire w_dff_A_87h3UxEH1_0;
	wire w_dff_A_WtGHggMp3_0;
	wire w_dff_A_6GAAc6RP9_0;
	wire w_dff_A_NlVlxsS29_0;
	wire w_dff_A_qEFfAEZq2_0;
	wire w_dff_A_KAjV3HxG2_0;
	wire w_dff_A_zhSAuQKB4_0;
	wire w_dff_A_4lAkaNN30_0;
	wire w_dff_A_mHHFsiDr7_0;
	wire w_dff_A_JCOnup5O1_0;
	wire w_dff_A_EScLjh3c1_0;
	wire w_dff_A_KK68eYoc4_0;
	wire w_dff_A_A3dIK2xS6_0;
	wire w_dff_A_Adjwx5WL4_0;
	wire w_dff_A_zdxO5D4b5_0;
	wire w_dff_A_hsHi8AYr0_0;
	wire w_dff_A_Mg1X7kYi3_2;
	wire w_dff_A_2qyJRMkA9_0;
	wire w_dff_A_BvZPiXOZ1_0;
	wire w_dff_A_TvY2d2tY5_0;
	wire w_dff_A_7R5GOZxK4_0;
	wire w_dff_A_ATA3UeNa2_0;
	wire w_dff_A_NLanNwY27_0;
	wire w_dff_A_RfXxmmml3_0;
	wire w_dff_A_Y6LGIcFt5_0;
	wire w_dff_A_IHAPyJVP3_0;
	wire w_dff_A_dJ6Fhpld1_0;
	wire w_dff_A_JHshYPrD9_0;
	wire w_dff_A_seeCy2Kh2_0;
	wire w_dff_A_nhVTJuWH6_0;
	wire w_dff_A_H0NHJC9x9_0;
	wire w_dff_A_A8G9NNRv7_0;
	wire w_dff_A_FY8nLnZF1_0;
	wire w_dff_A_WMQTWhBY1_0;
	wire w_dff_A_76rm7cOk5_0;
	wire w_dff_A_OBMLu1gw6_0;
	wire w_dff_A_botBkKyD1_0;
	wire w_dff_A_HxraTx742_0;
	wire w_dff_A_iv5Ka1kQ3_0;
	wire w_dff_A_CwhZzTZn9_2;
	wire w_dff_A_tbPRJOkG3_0;
	wire w_dff_A_XslWL3Q60_0;
	wire w_dff_A_p12QtY3W0_0;
	wire w_dff_A_GAJ89qqD4_0;
	wire w_dff_A_tZIVaVvy3_0;
	wire w_dff_A_Rvp6YINZ0_0;
	wire w_dff_A_eeohvE6f8_0;
	wire w_dff_A_pWRahA418_0;
	wire w_dff_A_l0gaW0P47_0;
	wire w_dff_A_GfyRGFpY7_0;
	wire w_dff_A_ekRWmT9K0_0;
	wire w_dff_A_zo52ntwV2_0;
	wire w_dff_A_jqpPCvAa8_0;
	wire w_dff_A_LftrWyT60_0;
	wire w_dff_A_HbxrLCr01_0;
	wire w_dff_A_LCDLV67j8_0;
	wire w_dff_A_SJ9EuBEv5_0;
	wire w_dff_A_h5UXlaAh7_0;
	wire w_dff_A_1sC049pU4_0;
	wire w_dff_A_5mAlZ4cm9_0;
	wire w_dff_A_6Ai86vBq2_2;
	wire w_dff_A_a1VLTSCQ7_0;
	wire w_dff_A_IRgXpY0P6_0;
	wire w_dff_A_qDronPmb3_0;
	wire w_dff_A_FZN0y7y06_0;
	wire w_dff_A_O4Lpzdwo0_0;
	wire w_dff_A_XJFN3vim8_0;
	wire w_dff_A_Q4HwkHwE8_0;
	wire w_dff_A_w9looatv2_0;
	wire w_dff_A_dMMYrJ129_0;
	wire w_dff_A_xJTKLktf7_0;
	wire w_dff_A_6wb2kHls0_0;
	wire w_dff_A_EEPKoRtu3_0;
	wire w_dff_A_SLmZPEzj6_0;
	wire w_dff_A_0wp4JsRD2_0;
	wire w_dff_A_NecOSmkM1_0;
	wire w_dff_A_6a1JAple9_0;
	wire w_dff_A_GHovIGQH4_0;
	wire w_dff_A_gprhUM183_0;
	wire w_dff_A_L32hW2LS1_2;
	wire w_dff_A_iBoSeqZ20_0;
	wire w_dff_A_R1ARCxDp7_0;
	wire w_dff_A_FXDStuyO8_0;
	wire w_dff_A_cYNaAvBj0_0;
	wire w_dff_A_jUExLUyv5_0;
	wire w_dff_A_71jGEFgd5_0;
	wire w_dff_A_s4THd8ww1_0;
	wire w_dff_A_4PPJga7z6_0;
	wire w_dff_A_m6g3Z6dN4_0;
	wire w_dff_A_Fvialyc24_0;
	wire w_dff_A_S9UxOVWJ3_0;
	wire w_dff_A_XN0ANblW1_0;
	wire w_dff_A_Vf4sA6Ky9_0;
	wire w_dff_A_UqpThG0K5_0;
	wire w_dff_A_ID7eH4Lh0_0;
	wire w_dff_A_q9MdTBve0_0;
	wire w_dff_A_U4vuyFKf9_2;
	wire w_dff_A_1EfTJIz48_0;
	wire w_dff_A_ZD3ppNsg2_0;
	wire w_dff_A_dqws9YBK7_0;
	wire w_dff_A_hUuoMGJp2_0;
	wire w_dff_A_9fFbRT7h1_0;
	wire w_dff_A_3EUl0YvF1_0;
	wire w_dff_A_HoHzlm9f1_0;
	wire w_dff_A_8WCLFQ7O6_0;
	wire w_dff_A_tdvirqIT9_0;
	wire w_dff_A_ll3i0FjZ5_0;
	wire w_dff_A_EE7XoC5N7_0;
	wire w_dff_A_rsW6fxGB1_0;
	wire w_dff_A_gYBEpimB0_0;
	wire w_dff_A_0f26mPQq5_0;
	wire w_dff_A_nROzBrc79_2;
	wire w_dff_A_1vMYkrXz2_0;
	wire w_dff_A_XcRWpCha5_0;
	wire w_dff_A_y2jtvMmp1_0;
	wire w_dff_A_D9PLMhrS7_0;
	wire w_dff_A_O7AZxJAF0_0;
	wire w_dff_A_JpOTPatm4_0;
	wire w_dff_A_U3alkdkB6_0;
	wire w_dff_A_aBjB7jI41_0;
	wire w_dff_A_SaEu00Pt2_0;
	wire w_dff_A_DZtfkPET7_0;
	wire w_dff_A_Lj47b4v46_0;
	wire w_dff_A_rjdUdsfB2_0;
	wire w_dff_A_Hct20z8J2_2;
	wire w_dff_A_2UwWnLJQ9_0;
	wire w_dff_A_35PE9aVP0_0;
	wire w_dff_A_rlxzxRmH2_0;
	wire w_dff_A_kRC3yNG81_0;
	wire w_dff_A_ikuaTzLq8_0;
	wire w_dff_A_Nu0umgT08_0;
	wire w_dff_A_9Vrmr2321_0;
	wire w_dff_A_NjidA3oc1_0;
	wire w_dff_A_1mrt8IqO9_0;
	wire w_dff_A_alY01VwI7_0;
	wire w_dff_A_48KSIqDl5_2;
	wire w_dff_A_asVgSdPS4_0;
	wire w_dff_A_o8KvXOaC8_0;
	wire w_dff_A_mVAHhzcV7_0;
	wire w_dff_A_0WIRGioh0_0;
	wire w_dff_A_Xnt55Kve0_0;
	wire w_dff_A_ig11lh6X4_0;
	wire w_dff_A_YU1PYqp05_0;
	wire w_dff_A_pJpFmTC08_0;
	wire w_dff_A_uIbrthHL5_2;
	wire w_dff_A_nvLQ7oa05_0;
	wire w_dff_A_qEEUoxZz6_0;
	wire w_dff_A_e706UnFA6_0;
	wire w_dff_A_Wcb4ODzY8_0;
	wire w_dff_A_UOVXcXQh8_0;
	wire w_dff_A_XgkLyMkz7_0;
	wire w_dff_A_UUSXDR6i6_2;
	wire w_dff_A_uBwifqyv9_0;
	wire w_dff_A_oQ1DY9T72_0;
	wire w_dff_A_IQ7iIc6H0_0;
	wire w_dff_A_BKciDslk4_0;
	wire w_dff_A_zwUMdALK2_2;
	wire w_dff_A_xozSZBXo9_0;
	wire w_dff_A_odSiYtK84_0;
	wire w_dff_A_KQCoHiXA8_2;
	jand g0000(.dina(w_G273gat_7[2]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G273gat_7[1]),.dinb(w_G18gat_7[2]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_G290gat_7[2]),.dinb(w_G1gat_7[0]),.dout(n66),.clk(gclk));
	jor g0003(.dina(n66),.dinb(w_n65_0[1]),.dout(n67),.clk(gclk));
	jand g0004(.dina(w_G290gat_7[1]),.dinb(w_G18gat_7[1]),.dout(n68),.clk(gclk));
	jand g0005(.dina(n68),.dinb(w_G545gat_0),.dout(n69),.clk(gclk));
	jnot g0006(.din(w_n69_0[1]),.dout(n70),.clk(gclk));
	jand g0007(.dina(w_n70_0[1]),.dinb(w_dff_B_FlnRawTX7_1),.dout(w_dff_A_oHlkIbp78_2),.clk(gclk));
	jand g0008(.dina(w_G307gat_7[2]),.dinb(w_G1gat_6[2]),.dout(n72),.clk(gclk));
	jnot g0009(.din(w_n72_0[1]),.dout(n73),.clk(gclk));
	jnot g0010(.din(w_G18gat_7[0]),.dout(n74),.clk(gclk));
	jnot g0011(.din(w_G290gat_7[0]),.dout(n75),.clk(gclk));
	jor g0012(.dina(w_n75_0[1]),.dinb(n74),.dout(n76),.clk(gclk));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G273gat_7[0]),.dout(n78),.clk(gclk));
	jor g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79),.clk(gclk));
	jand g0016(.dina(n79),.dinb(n76),.dout(n80),.clk(gclk));
	jand g0017(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jand g0018(.dina(w_n81_0[1]),.dinb(w_n65_0[0]),.dout(n82),.clk(gclk));
	jor g0019(.dina(w_n82_1[1]),.dinb(n80),.dout(n83),.clk(gclk));
	jand g0020(.dina(n83),.dinb(w_n70_0[0]),.dout(n84),.clk(gclk));
	jnot g0021(.din(w_n82_1[0]),.dout(n85),.clk(gclk));
	jand g0022(.dina(w_n85_0[1]),.dinb(w_n69_0[0]),.dout(n86),.clk(gclk));
	jor g0023(.dina(w_dff_B_8fabrxSB4_0),.dinb(w_n84_0[1]),.dout(n87),.clk(gclk));
	jxor g0024(.dina(w_n87_0[1]),.dinb(w_dff_B_HbMs7I9A8_1),.dout(w_dff_A_vs4kgBu57_2),.clk(gclk));
	jand g0025(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n89),.clk(gclk));
	jnot g0026(.din(w_n89_0[1]),.dout(n90),.clk(gclk));
	jnot g0027(.din(w_n84_0[0]),.dout(n91),.clk(gclk));
	jor g0028(.dina(w_n87_0[0]),.dinb(w_n72_0[0]),.dout(n92),.clk(gclk));
	jand g0029(.dina(n92),.dinb(w_dff_B_3MngmSLX7_1),.dout(n93),.clk(gclk));
	jand g0030(.dina(w_G307gat_7[1]),.dinb(w_G18gat_6[2]),.dout(n94),.clk(gclk));
	jnot g0031(.din(w_n94_0[1]),.dout(n95),.clk(gclk));
	jand g0032(.dina(w_G273gat_6[2]),.dinb(w_G52gat_7[2]),.dout(n96),.clk(gclk));
	jor g0033(.dina(w_n96_0[1]),.dinb(w_n81_0[0]),.dout(n97),.clk(gclk));
	jand g0034(.dina(w_G273gat_6[1]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G290gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jand g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100),.clk(gclk));
	jnot g0037(.din(w_n100_1[1]),.dout(n101),.clk(gclk));
	jand g0038(.dina(w_n101_0[2]),.dinb(w_dff_B_GllUaxUV7_1),.dout(n102),.clk(gclk));
	jor g0039(.dina(n102),.dinb(w_n82_0[2]),.dout(n103),.clk(gclk));
	jand g0040(.dina(w_n101_0[1]),.dinb(w_n82_0[1]),.dout(n104),.clk(gclk));
	jnot g0041(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jand g0042(.dina(n105),.dinb(w_n103_0[1]),.dout(n106),.clk(gclk));
	jxor g0043(.dina(n106),.dinb(w_dff_B_5uOOUoA52_1),.dout(n107),.clk(gclk));
	jxor g0044(.dina(w_n107_0[1]),.dinb(w_n93_0[1]),.dout(n108),.clk(gclk));
	jxor g0045(.dina(w_n108_0[1]),.dinb(w_dff_B_Zp5c4yA99_1),.dout(w_dff_A_D1J7lZ8S1_2),.clk(gclk));
	jand g0046(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n110),.clk(gclk));
	jnot g0047(.din(w_n110_0[1]),.dout(n111),.clk(gclk));
	jnot g0048(.din(w_n107_0[0]),.dout(n112),.clk(gclk));
	jor g0049(.dina(n112),.dinb(w_n93_0[0]),.dout(n113),.clk(gclk));
	jor g0050(.dina(w_n108_0[0]),.dinb(w_n89_0[0]),.dout(n114),.clk(gclk));
	jand g0051(.dina(n114),.dinb(w_dff_B_uBqySN0o4_1),.dout(n115),.clk(gclk));
	jand g0052(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n116),.clk(gclk));
	jnot g0053(.din(w_n116_0[1]),.dout(n117),.clk(gclk));
	jor g0054(.dina(w_n75_0[0]),.dinb(w_n77_0[0]),.dout(n118),.clk(gclk));
	jnot g0055(.din(w_G52gat_7[0]),.dout(n119),.clk(gclk));
	jor g0056(.dina(w_n78_0[0]),.dinb(n119),.dout(n120),.clk(gclk));
	jand g0057(.dina(n120),.dinb(n118),.dout(n121),.clk(gclk));
	jor g0058(.dina(w_n100_1[0]),.dinb(n121),.dout(n122),.clk(gclk));
	jand g0059(.dina(n122),.dinb(w_n85_0[0]),.dout(n123),.clk(gclk));
	jor g0060(.dina(w_n104_0[0]),.dinb(n123),.dout(n124),.clk(gclk));
	jor g0061(.dina(n124),.dinb(w_n94_0[0]),.dout(n125),.clk(gclk));
	jand g0062(.dina(n125),.dinb(w_n103_0[0]),.dout(n126),.clk(gclk));
	jand g0063(.dina(w_G307gat_7[0]),.dinb(w_G35gat_6[2]),.dout(n127),.clk(gclk));
	jnot g0064(.din(n127),.dout(n128),.clk(gclk));
	jand g0065(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[1]),.dout(n129),.clk(gclk));
	jor g0066(.dina(w_n129_0[1]),.dinb(w_n99_0[0]),.dout(n130),.clk(gclk));
	jand g0067(.dina(w_G290gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n131),.clk(gclk));
	jand g0068(.dina(w_n131_0[1]),.dinb(w_n96_0[0]),.dout(n132),.clk(gclk));
	jnot g0069(.din(w_n132_0[2]),.dout(n133),.clk(gclk));
	jand g0070(.dina(w_n133_0[2]),.dinb(w_n130_0[1]),.dout(n134),.clk(gclk));
	jor g0071(.dina(n134),.dinb(w_n100_0[2]),.dout(n135),.clk(gclk));
	jand g0072(.dina(w_n133_0[1]),.dinb(w_n100_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(n136),.dout(n137),.clk(gclk));
	jand g0074(.dina(n137),.dinb(n135),.dout(n138),.clk(gclk));
	jxor g0075(.dina(w_n138_0[1]),.dinb(w_n128_0[1]),.dout(n139),.clk(gclk));
	jnot g0076(.din(w_n139_0[1]),.dout(n140),.clk(gclk));
	jxor g0077(.dina(w_n140_0[1]),.dinb(w_n126_0[2]),.dout(n141),.clk(gclk));
	jxor g0078(.dina(n141),.dinb(w_dff_B_WOKIVqPd1_1),.dout(n142),.clk(gclk));
	jxor g0079(.dina(w_n142_0[1]),.dinb(w_n115_0[1]),.dout(n143),.clk(gclk));
	jxor g0080(.dina(w_n143_0[1]),.dinb(w_dff_B_oWExCNQ75_1),.dout(w_dff_A_PldpzvGS2_2),.clk(gclk));
	jand g0081(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n145),.clk(gclk));
	jnot g0082(.din(w_n145_0[1]),.dout(n146),.clk(gclk));
	jnot g0083(.din(w_n142_0[0]),.dout(n147),.clk(gclk));
	jor g0084(.dina(n147),.dinb(w_n115_0[0]),.dout(n148),.clk(gclk));
	jor g0085(.dina(w_n143_0[0]),.dinb(w_n110_0[0]),.dout(n149),.clk(gclk));
	jand g0086(.dina(n149),.dinb(w_dff_B_2rxQ8rZv0_1),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n151),.clk(gclk));
	jnot g0088(.din(w_n151_0[1]),.dout(n152),.clk(gclk));
	jor g0089(.dina(w_n140_0[0]),.dinb(w_n126_0[1]),.dout(n153),.clk(gclk));
	jxor g0090(.dina(w_n139_0[0]),.dinb(w_n126_0[0]),.dout(n154),.clk(gclk));
	jor g0091(.dina(n154),.dinb(w_n116_0[0]),.dout(n155),.clk(gclk));
	jand g0092(.dina(n155),.dinb(w_dff_B_6qB0mknv3_1),.dout(n156),.clk(gclk));
	jand g0093(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n157),.clk(gclk));
	jnot g0094(.din(n157),.dout(n158),.clk(gclk));
	jnot g0095(.din(w_n130_0[0]),.dout(n159),.clk(gclk));
	jor g0096(.dina(w_n132_0[1]),.dinb(n159),.dout(n160),.clk(gclk));
	jand g0097(.dina(n160),.dinb(w_n101_0[0]),.dout(n161),.clk(gclk));
	jand g0098(.dina(w_n138_0[0]),.dinb(w_n128_0[0]),.dout(n162),.clk(gclk));
	jor g0099(.dina(n162),.dinb(w_dff_B_CJuuASMf2_1),.dout(n163),.clk(gclk));
	jand g0100(.dina(w_G307gat_6[2]),.dinb(w_G52gat_6[2]),.dout(n164),.clk(gclk));
	jnot g0101(.din(n164),.dout(n165),.clk(gclk));
	jand g0102(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n166),.clk(gclk));
	jor g0103(.dina(w_n166_0[1]),.dinb(w_n131_0[0]),.dout(n167),.clk(gclk));
	jand g0104(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n168),.clk(gclk));
	jand g0105(.dina(w_n168_0[1]),.dinb(w_n129_0[0]),.dout(n169),.clk(gclk));
	jnot g0106(.din(w_n169_0[2]),.dout(n170),.clk(gclk));
	jand g0107(.dina(w_n170_0[1]),.dinb(w_dff_B_pFdws3C57_1),.dout(n171),.clk(gclk));
	jor g0108(.dina(n171),.dinb(w_n132_0[0]),.dout(n172),.clk(gclk));
	jor g0109(.dina(w_n169_0[1]),.dinb(w_n133_0[0]),.dout(n173),.clk(gclk));
	jand g0110(.dina(w_dff_B_WDlZjkOk6_0),.dinb(w_n172_0[1]),.dout(n174),.clk(gclk));
	jxor g0111(.dina(w_n174_0[1]),.dinb(w_n165_0[1]),.dout(n175),.clk(gclk));
	jxor g0112(.dina(w_n175_0[1]),.dinb(w_n163_0[1]),.dout(n176),.clk(gclk));
	jxor g0113(.dina(w_n176_0[1]),.dinb(w_n158_0[1]),.dout(n177),.clk(gclk));
	jnot g0114(.din(w_n177_0[1]),.dout(n178),.clk(gclk));
	jxor g0115(.dina(w_n178_0[1]),.dinb(w_n156_0[2]),.dout(n179),.clk(gclk));
	jxor g0116(.dina(n179),.dinb(w_dff_B_owl5xRXF4_1),.dout(n180),.clk(gclk));
	jxor g0117(.dina(w_n180_0[1]),.dinb(w_n150_0[1]),.dout(n181),.clk(gclk));
	jxor g0118(.dina(w_n181_0[1]),.dinb(w_dff_B_nEJzxkY00_1),.dout(w_dff_A_YL90IabU6_2),.clk(gclk));
	jand g0119(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n183),.clk(gclk));
	jnot g0120(.din(w_n183_0[1]),.dout(n184),.clk(gclk));
	jnot g0121(.din(w_n180_0[0]),.dout(n185),.clk(gclk));
	jor g0122(.dina(n185),.dinb(w_n150_0[0]),.dout(n186),.clk(gclk));
	jor g0123(.dina(w_n181_0[0]),.dinb(w_n145_0[0]),.dout(n187),.clk(gclk));
	jand g0124(.dina(n187),.dinb(w_dff_B_NiuiUYAR7_1),.dout(n188),.clk(gclk));
	jand g0125(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n189),.clk(gclk));
	jnot g0126(.din(w_n189_0[1]),.dout(n190),.clk(gclk));
	jor g0127(.dina(w_n178_0[0]),.dinb(w_n156_0[1]),.dout(n191),.clk(gclk));
	jxor g0128(.dina(w_n177_0[0]),.dinb(w_n156_0[0]),.dout(n192),.clk(gclk));
	jor g0129(.dina(n192),.dinb(w_n151_0[0]),.dout(n193),.clk(gclk));
	jand g0130(.dina(n193),.dinb(w_dff_B_ScOtqCUR0_1),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n195),.clk(gclk));
	jnot g0132(.din(n195),.dout(n196),.clk(gclk));
	jand g0133(.dina(w_n175_0[0]),.dinb(w_n163_0[0]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_n176_0[0]),.dinb(w_n158_0[0]),.dout(n198),.clk(gclk));
	jor g0135(.dina(n198),.dinb(w_dff_B_rb5e9BaE9_1),.dout(n199),.clk(gclk));
	jand g0136(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n200),.clk(gclk));
	jnot g0137(.din(n200),.dout(n201),.clk(gclk));
	jnot g0138(.din(w_n172_0[0]),.dout(n202),.clk(gclk));
	jand g0139(.dina(w_n174_0[0]),.dinb(w_n165_0[0]),.dout(n203),.clk(gclk));
	jor g0140(.dina(n203),.dinb(w_dff_B_CnGC1LJ43_1),.dout(n204),.clk(gclk));
	jand g0141(.dina(w_G307gat_6[1]),.dinb(w_G69gat_6[2]),.dout(n205),.clk(gclk));
	jnot g0142(.din(n205),.dout(n206),.clk(gclk));
	jand g0143(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n207),.clk(gclk));
	jor g0144(.dina(w_n207_0[1]),.dinb(w_n168_0[0]),.dout(n208),.clk(gclk));
	jand g0145(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n209),.clk(gclk));
	jand g0146(.dina(w_n209_0[1]),.dinb(w_n166_0[0]),.dout(n210),.clk(gclk));
	jnot g0147(.din(w_n210_1[1]),.dout(n211),.clk(gclk));
	jand g0148(.dina(n211),.dinb(w_dff_B_x3G1lenS0_1),.dout(n212),.clk(gclk));
	jor g0149(.dina(n212),.dinb(w_n169_0[0]),.dout(n213),.clk(gclk));
	jor g0150(.dina(w_n210_1[0]),.dinb(w_n170_0[0]),.dout(n214),.clk(gclk));
	jand g0151(.dina(w_dff_B_KeyIPZfW7_0),.dinb(w_n213_0[1]),.dout(n215),.clk(gclk));
	jxor g0152(.dina(w_n215_0[1]),.dinb(w_n206_0[1]),.dout(n216),.clk(gclk));
	jxor g0153(.dina(w_n216_0[1]),.dinb(w_n204_0[1]),.dout(n217),.clk(gclk));
	jxor g0154(.dina(w_n217_0[1]),.dinb(w_n201_0[1]),.dout(n218),.clk(gclk));
	jxor g0155(.dina(w_n218_0[1]),.dinb(w_n199_0[1]),.dout(n219),.clk(gclk));
	jxor g0156(.dina(w_n219_0[1]),.dinb(w_n196_0[1]),.dout(n220),.clk(gclk));
	jnot g0157(.din(w_n220_0[1]),.dout(n221),.clk(gclk));
	jxor g0158(.dina(w_n221_0[1]),.dinb(w_n194_0[2]),.dout(n222),.clk(gclk));
	jxor g0159(.dina(n222),.dinb(w_dff_B_EHlu3dn94_1),.dout(n223),.clk(gclk));
	jxor g0160(.dina(w_n223_0[1]),.dinb(w_n188_0[1]),.dout(n224),.clk(gclk));
	jxor g0161(.dina(w_n224_0[1]),.dinb(w_dff_B_YCIsNlDY6_1),.dout(w_dff_A_ML3PYmGw6_2),.clk(gclk));
	jand g0162(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n226),.clk(gclk));
	jnot g0163(.din(w_n226_0[1]),.dout(n227),.clk(gclk));
	jnot g0164(.din(w_n223_0[0]),.dout(n228),.clk(gclk));
	jor g0165(.dina(n228),.dinb(w_n188_0[0]),.dout(n229),.clk(gclk));
	jor g0166(.dina(w_n224_0[0]),.dinb(w_n183_0[0]),.dout(n230),.clk(gclk));
	jand g0167(.dina(n230),.dinb(w_dff_B_0vmM2Dpk6_1),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n232),.clk(gclk));
	jnot g0169(.din(w_n232_0[1]),.dout(n233),.clk(gclk));
	jor g0170(.dina(w_n221_0[0]),.dinb(w_n194_0[1]),.dout(n234),.clk(gclk));
	jxor g0171(.dina(w_n220_0[0]),.dinb(w_n194_0[0]),.dout(n235),.clk(gclk));
	jor g0172(.dina(n235),.dinb(w_n189_0[0]),.dout(n236),.clk(gclk));
	jand g0173(.dina(n236),.dinb(w_dff_B_dAuOBgIL1_1),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n238),.clk(gclk));
	jnot g0175(.din(n238),.dout(n239),.clk(gclk));
	jand g0176(.dina(w_n218_0[0]),.dinb(w_n199_0[0]),.dout(n240),.clk(gclk));
	jand g0177(.dina(w_n219_0[0]),.dinb(w_n196_0[0]),.dout(n241),.clk(gclk));
	jor g0178(.dina(n241),.dinb(w_dff_B_Q7T7t4QA3_1),.dout(n242),.clk(gclk));
	jand g0179(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(n243),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_n216_0[0]),.dinb(w_n204_0[0]),.dout(n245),.clk(gclk));
	jand g0182(.dina(w_n217_0[0]),.dinb(w_n201_0[0]),.dout(n246),.clk(gclk));
	jor g0183(.dina(n246),.dinb(w_dff_B_15bCaxtq3_1),.dout(n247),.clk(gclk));
	jand g0184(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n248),.clk(gclk));
	jnot g0185(.din(n248),.dout(n249),.clk(gclk));
	jnot g0186(.din(w_n213_0[0]),.dout(n250),.clk(gclk));
	jand g0187(.dina(w_n215_0[0]),.dinb(w_n206_0[0]),.dout(n251),.clk(gclk));
	jor g0188(.dina(n251),.dinb(w_dff_B_f4uAbTBS5_1),.dout(n252),.clk(gclk));
	jand g0189(.dina(w_G307gat_6[0]),.dinb(w_G86gat_6[2]),.dout(n253),.clk(gclk));
	jnot g0190(.din(n253),.dout(n254),.clk(gclk));
	jand g0191(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n255),.clk(gclk));
	jor g0192(.dina(w_n255_0[1]),.dinb(w_n209_0[0]),.dout(n256),.clk(gclk));
	jand g0193(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n257),.clk(gclk));
	jand g0194(.dina(w_n257_0[1]),.dinb(w_n207_0[0]),.dout(n258),.clk(gclk));
	jnot g0195(.din(w_n258_0[2]),.dout(n259),.clk(gclk));
	jand g0196(.dina(w_n259_0[1]),.dinb(w_dff_B_ld0GMe2J5_1),.dout(n260),.clk(gclk));
	jor g0197(.dina(n260),.dinb(w_n210_0[2]),.dout(n261),.clk(gclk));
	jand g0198(.dina(w_n259_0[0]),.dinb(w_n210_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(n262),.dout(n263),.clk(gclk));
	jand g0200(.dina(n263),.dinb(w_n261_0[1]),.dout(n264),.clk(gclk));
	jxor g0201(.dina(w_n264_0[1]),.dinb(w_n254_0[1]),.dout(n265),.clk(gclk));
	jxor g0202(.dina(w_n265_0[1]),.dinb(w_n252_0[1]),.dout(n266),.clk(gclk));
	jxor g0203(.dina(w_n266_0[1]),.dinb(w_n249_0[1]),.dout(n267),.clk(gclk));
	jxor g0204(.dina(w_n267_0[1]),.dinb(w_n247_0[1]),.dout(n268),.clk(gclk));
	jxor g0205(.dina(w_n268_0[1]),.dinb(w_n244_0[1]),.dout(n269),.clk(gclk));
	jxor g0206(.dina(w_n269_0[1]),.dinb(w_n242_0[1]),.dout(n270),.clk(gclk));
	jxor g0207(.dina(w_n270_0[1]),.dinb(w_n239_0[1]),.dout(n271),.clk(gclk));
	jnot g0208(.din(w_n271_0[1]),.dout(n272),.clk(gclk));
	jxor g0209(.dina(w_n272_0[1]),.dinb(w_n237_0[2]),.dout(n273),.clk(gclk));
	jxor g0210(.dina(n273),.dinb(w_dff_B_zlTyNM2h9_1),.dout(n274),.clk(gclk));
	jxor g0211(.dina(w_n274_0[1]),.dinb(w_n231_0[1]),.dout(n275),.clk(gclk));
	jxor g0212(.dina(w_n275_0[1]),.dinb(w_dff_B_rVL77JfP0_1),.dout(w_dff_A_p8CWdcT47_2),.clk(gclk));
	jand g0213(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n277),.clk(gclk));
	jnot g0214(.din(w_n277_0[1]),.dout(n278),.clk(gclk));
	jnot g0215(.din(w_n274_0[0]),.dout(n279),.clk(gclk));
	jor g0216(.dina(n279),.dinb(w_n231_0[0]),.dout(n280),.clk(gclk));
	jor g0217(.dina(w_n275_0[0]),.dinb(w_n226_0[0]),.dout(n281),.clk(gclk));
	jand g0218(.dina(n281),.dinb(w_dff_B_zvFQplgs5_1),.dout(n282),.clk(gclk));
	jand g0219(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(w_n283_0[1]),.dout(n284),.clk(gclk));
	jor g0221(.dina(w_n272_0[0]),.dinb(w_n237_0[1]),.dout(n285),.clk(gclk));
	jxor g0222(.dina(w_n271_0[0]),.dinb(w_n237_0[0]),.dout(n286),.clk(gclk));
	jor g0223(.dina(n286),.dinb(w_n232_0[0]),.dout(n287),.clk(gclk));
	jand g0224(.dina(n287),.dinb(w_dff_B_9jqgJuYA5_1),.dout(n288),.clk(gclk));
	jand g0225(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n289),.clk(gclk));
	jnot g0226(.din(n289),.dout(n290),.clk(gclk));
	jand g0227(.dina(w_n269_0[0]),.dinb(w_n242_0[0]),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n270_0[0]),.dinb(w_n239_0[0]),.dout(n292),.clk(gclk));
	jor g0229(.dina(n292),.dinb(w_dff_B_93cARDKC8_1),.dout(n293),.clk(gclk));
	jand g0230(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_n267_0[0]),.dinb(w_n247_0[0]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n268_0[0]),.dinb(w_n244_0[0]),.dout(n297),.clk(gclk));
	jor g0234(.dina(n297),.dinb(w_dff_B_iRswQ0ey1_1),.dout(n298),.clk(gclk));
	jand g0235(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n299),.clk(gclk));
	jnot g0236(.din(n299),.dout(n300),.clk(gclk));
	jand g0237(.dina(w_n265_0[0]),.dinb(w_n252_0[0]),.dout(n301),.clk(gclk));
	jand g0238(.dina(w_n266_0[0]),.dinb(w_n249_0[0]),.dout(n302),.clk(gclk));
	jor g0239(.dina(n302),.dinb(w_dff_B_OkUzAfi64_1),.dout(n303),.clk(gclk));
	jand g0240(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n304),.clk(gclk));
	jnot g0241(.din(n304),.dout(n305),.clk(gclk));
	jnot g0242(.din(w_n261_0[0]),.dout(n306),.clk(gclk));
	jand g0243(.dina(w_n264_0[0]),.dinb(w_n254_0[0]),.dout(n307),.clk(gclk));
	jor g0244(.dina(n307),.dinb(w_dff_B_Us5gRVrN8_1),.dout(n308),.clk(gclk));
	jand g0245(.dina(w_G307gat_5[2]),.dinb(w_G103gat_6[2]),.dout(n309),.clk(gclk));
	jnot g0246(.din(n309),.dout(n310),.clk(gclk));
	jand g0247(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n311),.clk(gclk));
	jor g0248(.dina(w_n311_0[1]),.dinb(w_n257_0[0]),.dout(n312),.clk(gclk));
	jand g0249(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n313),.clk(gclk));
	jand g0250(.dina(w_n313_0[1]),.dinb(w_n255_0[0]),.dout(n314),.clk(gclk));
	jnot g0251(.din(w_n314_0[2]),.dout(n315),.clk(gclk));
	jand g0252(.dina(w_n315_0[1]),.dinb(w_dff_B_COEn0i7q4_1),.dout(n316),.clk(gclk));
	jor g0253(.dina(n316),.dinb(w_n258_0[1]),.dout(n317),.clk(gclk));
	jand g0254(.dina(w_n315_0[0]),.dinb(w_n258_0[0]),.dout(n318),.clk(gclk));
	jnot g0255(.din(n318),.dout(n319),.clk(gclk));
	jand g0256(.dina(n319),.dinb(w_n317_0[1]),.dout(n320),.clk(gclk));
	jxor g0257(.dina(w_n320_0[1]),.dinb(w_n310_0[1]),.dout(n321),.clk(gclk));
	jxor g0258(.dina(w_n321_0[1]),.dinb(w_n308_0[1]),.dout(n322),.clk(gclk));
	jxor g0259(.dina(w_n322_0[1]),.dinb(w_n305_0[1]),.dout(n323),.clk(gclk));
	jxor g0260(.dina(w_n323_0[1]),.dinb(w_n303_0[1]),.dout(n324),.clk(gclk));
	jxor g0261(.dina(w_n324_0[1]),.dinb(w_n300_0[1]),.dout(n325),.clk(gclk));
	jxor g0262(.dina(w_n325_0[1]),.dinb(w_n298_0[1]),.dout(n326),.clk(gclk));
	jxor g0263(.dina(w_n326_0[1]),.dinb(w_n295_0[1]),.dout(n327),.clk(gclk));
	jxor g0264(.dina(w_n327_0[1]),.dinb(w_n293_0[1]),.dout(n328),.clk(gclk));
	jxor g0265(.dina(w_n328_0[1]),.dinb(w_n290_0[1]),.dout(n329),.clk(gclk));
	jnot g0266(.din(w_n329_0[1]),.dout(n330),.clk(gclk));
	jxor g0267(.dina(w_n330_0[1]),.dinb(w_n288_0[2]),.dout(n331),.clk(gclk));
	jxor g0268(.dina(n331),.dinb(w_dff_B_qwvf0gmh5_1),.dout(n332),.clk(gclk));
	jxor g0269(.dina(w_n332_0[1]),.dinb(w_n282_0[1]),.dout(n333),.clk(gclk));
	jxor g0270(.dina(w_n333_0[1]),.dinb(w_dff_B_oH3KqGwB4_1),.dout(w_dff_A_aV8fpFrx0_2),.clk(gclk));
	jand g0271(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n335),.clk(gclk));
	jnot g0272(.din(w_n335_0[1]),.dout(n336),.clk(gclk));
	jnot g0273(.din(w_n332_0[0]),.dout(n337),.clk(gclk));
	jor g0274(.dina(n337),.dinb(w_n282_0[0]),.dout(n338),.clk(gclk));
	jor g0275(.dina(w_n333_0[0]),.dinb(w_n277_0[0]),.dout(n339),.clk(gclk));
	jand g0276(.dina(n339),.dinb(w_dff_B_ibo5FJdy2_1),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n341),.clk(gclk));
	jnot g0278(.din(w_n341_0[1]),.dout(n342),.clk(gclk));
	jor g0279(.dina(w_n330_0[0]),.dinb(w_n288_0[1]),.dout(n343),.clk(gclk));
	jxor g0280(.dina(w_n329_0[0]),.dinb(w_n288_0[0]),.dout(n344),.clk(gclk));
	jor g0281(.dina(n344),.dinb(w_n283_0[0]),.dout(n345),.clk(gclk));
	jand g0282(.dina(n345),.dinb(w_dff_B_MxR0tMp03_1),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n347),.clk(gclk));
	jnot g0284(.din(n347),.dout(n348),.clk(gclk));
	jand g0285(.dina(w_n327_0[0]),.dinb(w_n293_0[0]),.dout(n349),.clk(gclk));
	jand g0286(.dina(w_n328_0[0]),.dinb(w_n290_0[0]),.dout(n350),.clk(gclk));
	jor g0287(.dina(n350),.dinb(w_dff_B_KohjZSWe6_1),.dout(n351),.clk(gclk));
	jand g0288(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n352),.clk(gclk));
	jnot g0289(.din(n352),.dout(n353),.clk(gclk));
	jand g0290(.dina(w_n325_0[0]),.dinb(w_n298_0[0]),.dout(n354),.clk(gclk));
	jand g0291(.dina(w_n326_0[0]),.dinb(w_n295_0[0]),.dout(n355),.clk(gclk));
	jor g0292(.dina(n355),.dinb(w_dff_B_ySOKwf7v3_1),.dout(n356),.clk(gclk));
	jand g0293(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n357),.clk(gclk));
	jnot g0294(.din(n357),.dout(n358),.clk(gclk));
	jand g0295(.dina(w_n323_0[0]),.dinb(w_n303_0[0]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_n324_0[0]),.dinb(w_n300_0[0]),.dout(n360),.clk(gclk));
	jor g0297(.dina(n360),.dinb(w_dff_B_OnsABkWv7_1),.dout(n361),.clk(gclk));
	jand g0298(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n362),.clk(gclk));
	jnot g0299(.din(n362),.dout(n363),.clk(gclk));
	jand g0300(.dina(w_n321_0[0]),.dinb(w_n308_0[0]),.dout(n364),.clk(gclk));
	jand g0301(.dina(w_n322_0[0]),.dinb(w_n305_0[0]),.dout(n365),.clk(gclk));
	jor g0302(.dina(n365),.dinb(w_dff_B_FqnL9AwD9_1),.dout(n366),.clk(gclk));
	jand g0303(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n367),.clk(gclk));
	jnot g0304(.din(n367),.dout(n368),.clk(gclk));
	jnot g0305(.din(w_n317_0[0]),.dout(n369),.clk(gclk));
	jand g0306(.dina(w_n320_0[0]),.dinb(w_n310_0[0]),.dout(n370),.clk(gclk));
	jor g0307(.dina(n370),.dinb(w_dff_B_8bw6Fr9D8_1),.dout(n371),.clk(gclk));
	jand g0308(.dina(w_G307gat_5[1]),.dinb(w_G120gat_6[2]),.dout(n372),.clk(gclk));
	jand g0309(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n373),.clk(gclk));
	jor g0310(.dina(w_n373_0[1]),.dinb(w_n313_0[0]),.dout(n374),.clk(gclk));
	jand g0311(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n375),.clk(gclk));
	jand g0312(.dina(w_n375_0[1]),.dinb(w_n311_0[0]),.dout(n376),.clk(gclk));
	jnot g0313(.din(w_n376_0[2]),.dout(n377),.clk(gclk));
	jand g0314(.dina(w_n377_0[1]),.dinb(w_dff_B_qmu8Bjy34_1),.dout(n378),.clk(gclk));
	jor g0315(.dina(n378),.dinb(w_n314_0[1]),.dout(n379),.clk(gclk));
	jnot g0316(.din(n379),.dout(n380),.clk(gclk));
	jand g0317(.dina(w_n377_0[0]),.dinb(w_n314_0[0]),.dout(n381),.clk(gclk));
	jor g0318(.dina(w_dff_B_4BpUftWB8_0),.dinb(w_n380_0[1]),.dout(n382),.clk(gclk));
	jxor g0319(.dina(w_n382_0[1]),.dinb(w_n372_0[1]),.dout(n383),.clk(gclk));
	jxor g0320(.dina(w_n383_0[1]),.dinb(w_n371_0[1]),.dout(n384),.clk(gclk));
	jxor g0321(.dina(w_n384_0[1]),.dinb(w_n368_0[1]),.dout(n385),.clk(gclk));
	jxor g0322(.dina(w_n385_0[1]),.dinb(w_n366_0[1]),.dout(n386),.clk(gclk));
	jxor g0323(.dina(w_n386_0[1]),.dinb(w_n363_0[1]),.dout(n387),.clk(gclk));
	jxor g0324(.dina(w_n387_0[1]),.dinb(w_n361_0[1]),.dout(n388),.clk(gclk));
	jxor g0325(.dina(w_n388_0[1]),.dinb(w_n358_0[1]),.dout(n389),.clk(gclk));
	jxor g0326(.dina(w_n389_0[1]),.dinb(w_n356_0[1]),.dout(n390),.clk(gclk));
	jxor g0327(.dina(w_n390_0[1]),.dinb(w_n353_0[1]),.dout(n391),.clk(gclk));
	jxor g0328(.dina(w_n391_0[1]),.dinb(w_n351_0[1]),.dout(n392),.clk(gclk));
	jxor g0329(.dina(w_n392_0[1]),.dinb(w_n348_0[1]),.dout(n393),.clk(gclk));
	jnot g0330(.din(w_n393_0[1]),.dout(n394),.clk(gclk));
	jxor g0331(.dina(w_n394_0[1]),.dinb(w_n346_0[2]),.dout(n395),.clk(gclk));
	jxor g0332(.dina(n395),.dinb(w_dff_B_qyHnPJs31_1),.dout(n396),.clk(gclk));
	jxor g0333(.dina(w_n396_0[1]),.dinb(w_n340_0[1]),.dout(n397),.clk(gclk));
	jxor g0334(.dina(w_n397_0[1]),.dinb(w_dff_B_piHzdoiB6_1),.dout(w_dff_A_xLPUpw6m3_2),.clk(gclk));
	jand g0335(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n399),.clk(gclk));
	jnot g0336(.din(w_n399_0[1]),.dout(n400),.clk(gclk));
	jnot g0337(.din(w_n396_0[0]),.dout(n401),.clk(gclk));
	jor g0338(.dina(n401),.dinb(w_n340_0[0]),.dout(n402),.clk(gclk));
	jor g0339(.dina(w_n397_0[0]),.dinb(w_n335_0[0]),.dout(n403),.clk(gclk));
	jand g0340(.dina(n403),.dinb(w_dff_B_G8Fc5G387_1),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n405),.clk(gclk));
	jnot g0342(.din(w_n405_0[1]),.dout(n406),.clk(gclk));
	jor g0343(.dina(w_n394_0[0]),.dinb(w_n346_0[1]),.dout(n407),.clk(gclk));
	jxor g0344(.dina(w_n393_0[0]),.dinb(w_n346_0[0]),.dout(n408),.clk(gclk));
	jor g0345(.dina(n408),.dinb(w_n341_0[0]),.dout(n409),.clk(gclk));
	jand g0346(.dina(n409),.dinb(w_dff_B_NRDAfc2w1_1),.dout(n410),.clk(gclk));
	jand g0347(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n411),.clk(gclk));
	jnot g0348(.din(n411),.dout(n412),.clk(gclk));
	jand g0349(.dina(w_n391_0[0]),.dinb(w_n351_0[0]),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n392_0[0]),.dinb(w_n348_0[0]),.dout(n414),.clk(gclk));
	jor g0351(.dina(n414),.dinb(w_dff_B_vkyvK0Dy8_1),.dout(n415),.clk(gclk));
	jand g0352(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n416),.clk(gclk));
	jnot g0353(.din(n416),.dout(n417),.clk(gclk));
	jand g0354(.dina(w_n389_0[0]),.dinb(w_n356_0[0]),.dout(n418),.clk(gclk));
	jand g0355(.dina(w_n390_0[0]),.dinb(w_n353_0[0]),.dout(n419),.clk(gclk));
	jor g0356(.dina(n419),.dinb(w_dff_B_Wnsct9yN9_1),.dout(n420),.clk(gclk));
	jand g0357(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n421),.clk(gclk));
	jnot g0358(.din(n421),.dout(n422),.clk(gclk));
	jand g0359(.dina(w_n387_0[0]),.dinb(w_n361_0[0]),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_n388_0[0]),.dinb(w_n358_0[0]),.dout(n424),.clk(gclk));
	jor g0361(.dina(n424),.dinb(w_dff_B_S3LDvzAM3_1),.dout(n425),.clk(gclk));
	jand g0362(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n426),.clk(gclk));
	jnot g0363(.din(n426),.dout(n427),.clk(gclk));
	jand g0364(.dina(w_n385_0[0]),.dinb(w_n366_0[0]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_n386_0[0]),.dinb(w_n363_0[0]),.dout(n429),.clk(gclk));
	jor g0366(.dina(n429),.dinb(w_dff_B_OxFG7zEq4_1),.dout(n430),.clk(gclk));
	jand g0367(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n431),.clk(gclk));
	jnot g0368(.din(n431),.dout(n432),.clk(gclk));
	jand g0369(.dina(w_n383_0[0]),.dinb(w_n371_0[0]),.dout(n433),.clk(gclk));
	jand g0370(.dina(w_n384_0[0]),.dinb(w_n368_0[0]),.dout(n434),.clk(gclk));
	jor g0371(.dina(n434),.dinb(w_dff_B_qL2BFsb78_1),.dout(n435),.clk(gclk));
	jand g0372(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n436),.clk(gclk));
	jnot g0373(.din(n436),.dout(n437),.clk(gclk));
	jnot g0374(.din(w_n372_0[0]),.dout(n438),.clk(gclk));
	jnot g0375(.din(w_n382_0[0]),.dout(n439),.clk(gclk));
	jand g0376(.dina(n439),.dinb(w_dff_B_Un0ukGf28_1),.dout(n440),.clk(gclk));
	jor g0377(.dina(n440),.dinb(w_n380_0[0]),.dout(n441),.clk(gclk));
	jand g0378(.dina(w_G307gat_5[0]),.dinb(w_G137gat_6[2]),.dout(n442),.clk(gclk));
	jand g0379(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n443),.clk(gclk));
	jor g0380(.dina(w_n443_0[1]),.dinb(w_n375_0[0]),.dout(n444),.clk(gclk));
	jand g0381(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n445),.clk(gclk));
	jand g0382(.dina(w_n445_0[1]),.dinb(w_n373_0[0]),.dout(n446),.clk(gclk));
	jnot g0383(.din(w_n446_0[2]),.dout(n447),.clk(gclk));
	jand g0384(.dina(w_n447_0[1]),.dinb(w_dff_B_N7i4VHMt8_1),.dout(n448),.clk(gclk));
	jor g0385(.dina(n448),.dinb(w_n376_0[1]),.dout(n449),.clk(gclk));
	jnot g0386(.din(n449),.dout(n450),.clk(gclk));
	jand g0387(.dina(w_n447_0[0]),.dinb(w_n376_0[0]),.dout(n451),.clk(gclk));
	jor g0388(.dina(w_dff_B_RAreoxw01_0),.dinb(w_n450_0[1]),.dout(n452),.clk(gclk));
	jxor g0389(.dina(w_n452_0[1]),.dinb(w_n442_0[1]),.dout(n453),.clk(gclk));
	jxor g0390(.dina(w_n453_0[1]),.dinb(w_n441_0[1]),.dout(n454),.clk(gclk));
	jxor g0391(.dina(w_n454_0[1]),.dinb(w_n437_0[1]),.dout(n455),.clk(gclk));
	jxor g0392(.dina(w_n455_0[1]),.dinb(w_n435_0[1]),.dout(n456),.clk(gclk));
	jxor g0393(.dina(w_n456_0[1]),.dinb(w_n432_0[1]),.dout(n457),.clk(gclk));
	jxor g0394(.dina(w_n457_0[1]),.dinb(w_n430_0[1]),.dout(n458),.clk(gclk));
	jxor g0395(.dina(w_n458_0[1]),.dinb(w_n427_0[1]),.dout(n459),.clk(gclk));
	jxor g0396(.dina(w_n459_0[1]),.dinb(w_n425_0[1]),.dout(n460),.clk(gclk));
	jxor g0397(.dina(w_n460_0[1]),.dinb(w_n422_0[1]),.dout(n461),.clk(gclk));
	jxor g0398(.dina(w_n461_0[1]),.dinb(w_n420_0[1]),.dout(n462),.clk(gclk));
	jxor g0399(.dina(w_n462_0[1]),.dinb(w_n417_0[1]),.dout(n463),.clk(gclk));
	jxor g0400(.dina(w_n463_0[1]),.dinb(w_n415_0[1]),.dout(n464),.clk(gclk));
	jxor g0401(.dina(w_n464_0[1]),.dinb(w_n412_0[1]),.dout(n465),.clk(gclk));
	jnot g0402(.din(w_n465_0[1]),.dout(n466),.clk(gclk));
	jxor g0403(.dina(w_n466_0[1]),.dinb(w_n410_0[2]),.dout(n467),.clk(gclk));
	jxor g0404(.dina(n467),.dinb(w_dff_B_5LHCkCEA4_1),.dout(n468),.clk(gclk));
	jxor g0405(.dina(w_n468_0[1]),.dinb(w_n404_0[1]),.dout(n469),.clk(gclk));
	jxor g0406(.dina(w_n469_0[1]),.dinb(w_dff_B_erQVcywS2_1),.dout(w_dff_A_0FjbwSqr7_2),.clk(gclk));
	jand g0407(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n471),.clk(gclk));
	jnot g0408(.din(w_n471_0[1]),.dout(n472),.clk(gclk));
	jnot g0409(.din(w_n468_0[0]),.dout(n473),.clk(gclk));
	jor g0410(.dina(n473),.dinb(w_n404_0[0]),.dout(n474),.clk(gclk));
	jor g0411(.dina(w_n469_0[0]),.dinb(w_n399_0[0]),.dout(n475),.clk(gclk));
	jand g0412(.dina(n475),.dinb(w_dff_B_AYmBTs4D8_1),.dout(n476),.clk(gclk));
	jand g0413(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n477),.clk(gclk));
	jnot g0414(.din(w_n477_0[1]),.dout(n478),.clk(gclk));
	jor g0415(.dina(w_n466_0[0]),.dinb(w_n410_0[1]),.dout(n479),.clk(gclk));
	jxor g0416(.dina(w_n465_0[0]),.dinb(w_n410_0[0]),.dout(n480),.clk(gclk));
	jor g0417(.dina(n480),.dinb(w_n405_0[0]),.dout(n481),.clk(gclk));
	jand g0418(.dina(n481),.dinb(w_dff_B_gogWROKv2_1),.dout(n482),.clk(gclk));
	jand g0419(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n463_0[0]),.dinb(w_n415_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n464_0[0]),.dinb(w_n412_0[0]),.dout(n486),.clk(gclk));
	jor g0423(.dina(n486),.dinb(w_dff_B_cQqrFy9q4_1),.dout(n487),.clk(gclk));
	jand g0424(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n461_0[0]),.dinb(w_n420_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n462_0[0]),.dinb(w_n417_0[0]),.dout(n491),.clk(gclk));
	jor g0428(.dina(n491),.dinb(w_dff_B_nNxqHRh25_1),.dout(n492),.clk(gclk));
	jand g0429(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jand g0431(.dina(w_n459_0[0]),.dinb(w_n425_0[0]),.dout(n495),.clk(gclk));
	jand g0432(.dina(w_n460_0[0]),.dinb(w_n422_0[0]),.dout(n496),.clk(gclk));
	jor g0433(.dina(n496),.dinb(w_dff_B_UeXsh9uZ9_1),.dout(n497),.clk(gclk));
	jand g0434(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_n457_0[0]),.dinb(w_n430_0[0]),.dout(n500),.clk(gclk));
	jand g0437(.dina(w_n458_0[0]),.dinb(w_n427_0[0]),.dout(n501),.clk(gclk));
	jor g0438(.dina(n501),.dinb(w_dff_B_6jsqFIrz7_1),.dout(n502),.clk(gclk));
	jand g0439(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n503),.clk(gclk));
	jnot g0440(.din(n503),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_n455_0[0]),.dinb(w_n435_0[0]),.dout(n505),.clk(gclk));
	jand g0442(.dina(w_n456_0[0]),.dinb(w_n432_0[0]),.dout(n506),.clk(gclk));
	jor g0443(.dina(n506),.dinb(w_dff_B_g62wjsut6_1),.dout(n507),.clk(gclk));
	jand g0444(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n508),.clk(gclk));
	jnot g0445(.din(n508),.dout(n509),.clk(gclk));
	jand g0446(.dina(w_n453_0[0]),.dinb(w_n441_0[0]),.dout(n510),.clk(gclk));
	jand g0447(.dina(w_n454_0[0]),.dinb(w_n437_0[0]),.dout(n511),.clk(gclk));
	jor g0448(.dina(n511),.dinb(w_dff_B_d1adPsZB7_1),.dout(n512),.clk(gclk));
	jand g0449(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n513),.clk(gclk));
	jnot g0450(.din(n513),.dout(n514),.clk(gclk));
	jnot g0451(.din(w_n442_0[0]),.dout(n515),.clk(gclk));
	jnot g0452(.din(w_n452_0[0]),.dout(n516),.clk(gclk));
	jand g0453(.dina(n516),.dinb(w_dff_B_qyNN8air7_1),.dout(n517),.clk(gclk));
	jor g0454(.dina(n517),.dinb(w_n450_0[0]),.dout(n518),.clk(gclk));
	jand g0455(.dina(w_G307gat_4[2]),.dinb(w_G154gat_6[2]),.dout(n519),.clk(gclk));
	jand g0456(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n520),.clk(gclk));
	jor g0457(.dina(w_n520_0[1]),.dinb(w_n445_0[0]),.dout(n521),.clk(gclk));
	jand g0458(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n522),.clk(gclk));
	jand g0459(.dina(w_n522_0[1]),.dinb(w_n443_0[0]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[2]),.dout(n524),.clk(gclk));
	jand g0461(.dina(w_n524_0[1]),.dinb(w_dff_B_oQXcnDpm6_1),.dout(n525),.clk(gclk));
	jor g0462(.dina(n525),.dinb(w_n446_0[1]),.dout(n526),.clk(gclk));
	jnot g0463(.din(n526),.dout(n527),.clk(gclk));
	jand g0464(.dina(w_n524_0[0]),.dinb(w_n446_0[0]),.dout(n528),.clk(gclk));
	jor g0465(.dina(w_dff_B_n7fgtk1y8_0),.dinb(w_n527_0[1]),.dout(n529),.clk(gclk));
	jxor g0466(.dina(w_n529_0[1]),.dinb(w_n519_0[1]),.dout(n530),.clk(gclk));
	jxor g0467(.dina(w_n530_0[1]),.dinb(w_n518_0[1]),.dout(n531),.clk(gclk));
	jxor g0468(.dina(w_n531_0[1]),.dinb(w_n514_0[1]),.dout(n532),.clk(gclk));
	jxor g0469(.dina(w_n532_0[1]),.dinb(w_n512_0[1]),.dout(n533),.clk(gclk));
	jxor g0470(.dina(w_n533_0[1]),.dinb(w_n509_0[1]),.dout(n534),.clk(gclk));
	jxor g0471(.dina(w_n534_0[1]),.dinb(w_n507_0[1]),.dout(n535),.clk(gclk));
	jxor g0472(.dina(w_n535_0[1]),.dinb(w_n504_0[1]),.dout(n536),.clk(gclk));
	jxor g0473(.dina(w_n536_0[1]),.dinb(w_n502_0[1]),.dout(n537),.clk(gclk));
	jxor g0474(.dina(w_n537_0[1]),.dinb(w_n499_0[1]),.dout(n538),.clk(gclk));
	jxor g0475(.dina(w_n538_0[1]),.dinb(w_n497_0[1]),.dout(n539),.clk(gclk));
	jxor g0476(.dina(w_n539_0[1]),.dinb(w_n494_0[1]),.dout(n540),.clk(gclk));
	jxor g0477(.dina(w_n540_0[1]),.dinb(w_n492_0[1]),.dout(n541),.clk(gclk));
	jxor g0478(.dina(w_n541_0[1]),.dinb(w_n489_0[1]),.dout(n542),.clk(gclk));
	jxor g0479(.dina(w_n542_0[1]),.dinb(w_n487_0[1]),.dout(n543),.clk(gclk));
	jxor g0480(.dina(w_n543_0[1]),.dinb(w_n484_0[1]),.dout(n544),.clk(gclk));
	jnot g0481(.din(w_n544_0[1]),.dout(n545),.clk(gclk));
	jxor g0482(.dina(w_n545_0[1]),.dinb(w_n482_0[2]),.dout(n546),.clk(gclk));
	jxor g0483(.dina(n546),.dinb(w_dff_B_KRdIAUVx8_1),.dout(n547),.clk(gclk));
	jxor g0484(.dina(w_n547_0[1]),.dinb(w_n476_0[1]),.dout(n548),.clk(gclk));
	jxor g0485(.dina(w_n548_0[1]),.dinb(w_dff_B_OwwZINRB0_1),.dout(w_dff_A_TjdGLRLw9_2),.clk(gclk));
	jand g0486(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n550),.clk(gclk));
	jnot g0487(.din(w_n550_0[1]),.dout(n551),.clk(gclk));
	jnot g0488(.din(w_n547_0[0]),.dout(n552),.clk(gclk));
	jor g0489(.dina(n552),.dinb(w_n476_0[0]),.dout(n553),.clk(gclk));
	jor g0490(.dina(w_n548_0[0]),.dinb(w_n471_0[0]),.dout(n554),.clk(gclk));
	jand g0491(.dina(n554),.dinb(w_dff_B_SiMRqYSP0_1),.dout(n555),.clk(gclk));
	jand g0492(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n556),.clk(gclk));
	jnot g0493(.din(w_n556_0[1]),.dout(n557),.clk(gclk));
	jor g0494(.dina(w_n545_0[0]),.dinb(w_n482_0[1]),.dout(n558),.clk(gclk));
	jxor g0495(.dina(w_n544_0[0]),.dinb(w_n482_0[0]),.dout(n559),.clk(gclk));
	jor g0496(.dina(n559),.dinb(w_n477_0[0]),.dout(n560),.clk(gclk));
	jand g0497(.dina(n560),.dinb(w_dff_B_ceJJ1TqA2_1),.dout(n561),.clk(gclk));
	jand g0498(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n562),.clk(gclk));
	jnot g0499(.din(n562),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n542_0[0]),.dinb(w_n487_0[0]),.dout(n564),.clk(gclk));
	jand g0501(.dina(w_n543_0[0]),.dinb(w_n484_0[0]),.dout(n565),.clk(gclk));
	jor g0502(.dina(n565),.dinb(w_dff_B_zFuVlLZs2_1),.dout(n566),.clk(gclk));
	jand g0503(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n567),.clk(gclk));
	jnot g0504(.din(n567),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n540_0[0]),.dinb(w_n492_0[0]),.dout(n569),.clk(gclk));
	jand g0506(.dina(w_n541_0[0]),.dinb(w_n489_0[0]),.dout(n570),.clk(gclk));
	jor g0507(.dina(n570),.dinb(w_dff_B_1RE9BRv90_1),.dout(n571),.clk(gclk));
	jand g0508(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n572),.clk(gclk));
	jnot g0509(.din(n572),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n538_0[0]),.dinb(w_n497_0[0]),.dout(n574),.clk(gclk));
	jand g0511(.dina(w_n539_0[0]),.dinb(w_n494_0[0]),.dout(n575),.clk(gclk));
	jor g0512(.dina(n575),.dinb(w_dff_B_8DXc4VHP2_1),.dout(n576),.clk(gclk));
	jand g0513(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n577),.clk(gclk));
	jnot g0514(.din(n577),.dout(n578),.clk(gclk));
	jand g0515(.dina(w_n536_0[0]),.dinb(w_n502_0[0]),.dout(n579),.clk(gclk));
	jand g0516(.dina(w_n537_0[0]),.dinb(w_n499_0[0]),.dout(n580),.clk(gclk));
	jor g0517(.dina(n580),.dinb(w_dff_B_o79ldpKl3_1),.dout(n581),.clk(gclk));
	jand g0518(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n582),.clk(gclk));
	jnot g0519(.din(n582),.dout(n583),.clk(gclk));
	jand g0520(.dina(w_n534_0[0]),.dinb(w_n507_0[0]),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_n535_0[0]),.dinb(w_n504_0[0]),.dout(n585),.clk(gclk));
	jor g0522(.dina(n585),.dinb(w_dff_B_OlGt9Uuj4_1),.dout(n586),.clk(gclk));
	jand g0523(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n587),.clk(gclk));
	jnot g0524(.din(n587),.dout(n588),.clk(gclk));
	jand g0525(.dina(w_n532_0[0]),.dinb(w_n512_0[0]),.dout(n589),.clk(gclk));
	jand g0526(.dina(w_n533_0[0]),.dinb(w_n509_0[0]),.dout(n590),.clk(gclk));
	jor g0527(.dina(n590),.dinb(w_dff_B_31QFqtey6_1),.dout(n591),.clk(gclk));
	jand g0528(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n592),.clk(gclk));
	jnot g0529(.din(n592),.dout(n593),.clk(gclk));
	jand g0530(.dina(w_n530_0[0]),.dinb(w_n518_0[0]),.dout(n594),.clk(gclk));
	jand g0531(.dina(w_n531_0[0]),.dinb(w_n514_0[0]),.dout(n595),.clk(gclk));
	jor g0532(.dina(n595),.dinb(w_dff_B_9ghebZGk8_1),.dout(n596),.clk(gclk));
	jand g0533(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n597),.clk(gclk));
	jnot g0534(.din(n597),.dout(n598),.clk(gclk));
	jnot g0535(.din(w_n519_0[0]),.dout(n599),.clk(gclk));
	jnot g0536(.din(w_n529_0[0]),.dout(n600),.clk(gclk));
	jand g0537(.dina(n600),.dinb(w_dff_B_nDYSgVV54_1),.dout(n601),.clk(gclk));
	jor g0538(.dina(n601),.dinb(w_n527_0[0]),.dout(n602),.clk(gclk));
	jand g0539(.dina(w_G307gat_4[1]),.dinb(w_G171gat_6[2]),.dout(n603),.clk(gclk));
	jand g0540(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n604),.clk(gclk));
	jor g0541(.dina(w_n604_0[1]),.dinb(w_n522_0[0]),.dout(n605),.clk(gclk));
	jand g0542(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n606),.clk(gclk));
	jand g0543(.dina(w_n606_0[1]),.dinb(w_n520_0[0]),.dout(n607),.clk(gclk));
	jnot g0544(.din(w_n607_0[2]),.dout(n608),.clk(gclk));
	jand g0545(.dina(w_n608_0[1]),.dinb(w_dff_B_TWlLduFk8_1),.dout(n609),.clk(gclk));
	jor g0546(.dina(n609),.dinb(w_n523_0[1]),.dout(n610),.clk(gclk));
	jnot g0547(.din(n610),.dout(n611),.clk(gclk));
	jand g0548(.dina(w_n608_0[0]),.dinb(w_n523_0[0]),.dout(n612),.clk(gclk));
	jor g0549(.dina(w_dff_B_oqDe2AjM2_0),.dinb(w_n611_0[1]),.dout(n613),.clk(gclk));
	jxor g0550(.dina(w_n613_0[1]),.dinb(w_n603_0[1]),.dout(n614),.clk(gclk));
	jxor g0551(.dina(w_n614_0[1]),.dinb(w_n602_0[1]),.dout(n615),.clk(gclk));
	jxor g0552(.dina(w_n615_0[1]),.dinb(w_n598_0[1]),.dout(n616),.clk(gclk));
	jxor g0553(.dina(w_n616_0[1]),.dinb(w_n596_0[1]),.dout(n617),.clk(gclk));
	jxor g0554(.dina(w_n617_0[1]),.dinb(w_n593_0[1]),.dout(n618),.clk(gclk));
	jxor g0555(.dina(w_n618_0[1]),.dinb(w_n591_0[1]),.dout(n619),.clk(gclk));
	jxor g0556(.dina(w_n619_0[1]),.dinb(w_n588_0[1]),.dout(n620),.clk(gclk));
	jxor g0557(.dina(w_n620_0[1]),.dinb(w_n586_0[1]),.dout(n621),.clk(gclk));
	jxor g0558(.dina(w_n621_0[1]),.dinb(w_n583_0[1]),.dout(n622),.clk(gclk));
	jxor g0559(.dina(w_n622_0[1]),.dinb(w_n581_0[1]),.dout(n623),.clk(gclk));
	jxor g0560(.dina(w_n623_0[1]),.dinb(w_n578_0[1]),.dout(n624),.clk(gclk));
	jxor g0561(.dina(w_n624_0[1]),.dinb(w_n576_0[1]),.dout(n625),.clk(gclk));
	jxor g0562(.dina(w_n625_0[1]),.dinb(w_n573_0[1]),.dout(n626),.clk(gclk));
	jxor g0563(.dina(w_n626_0[1]),.dinb(w_n571_0[1]),.dout(n627),.clk(gclk));
	jxor g0564(.dina(w_n627_0[1]),.dinb(w_n568_0[1]),.dout(n628),.clk(gclk));
	jxor g0565(.dina(w_n628_0[1]),.dinb(w_n566_0[1]),.dout(n629),.clk(gclk));
	jxor g0566(.dina(w_n629_0[1]),.dinb(w_n563_0[1]),.dout(n630),.clk(gclk));
	jnot g0567(.din(w_n630_0[1]),.dout(n631),.clk(gclk));
	jxor g0568(.dina(w_n631_0[1]),.dinb(w_n561_0[2]),.dout(n632),.clk(gclk));
	jxor g0569(.dina(n632),.dinb(w_dff_B_roJGW98C6_1),.dout(n633),.clk(gclk));
	jxor g0570(.dina(w_n633_0[1]),.dinb(w_n555_0[1]),.dout(n634),.clk(gclk));
	jxor g0571(.dina(w_n634_0[1]),.dinb(w_dff_B_kK36N8uP3_1),.dout(w_dff_A_n39HOqln6_2),.clk(gclk));
	jand g0572(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n636),.clk(gclk));
	jnot g0573(.din(w_n636_0[1]),.dout(n637),.clk(gclk));
	jnot g0574(.din(w_n633_0[0]),.dout(n638),.clk(gclk));
	jor g0575(.dina(n638),.dinb(w_n555_0[0]),.dout(n639),.clk(gclk));
	jor g0576(.dina(w_n634_0[0]),.dinb(w_n550_0[0]),.dout(n640),.clk(gclk));
	jand g0577(.dina(n640),.dinb(w_dff_B_5vRFOpjz6_1),.dout(n641),.clk(gclk));
	jand g0578(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n642),.clk(gclk));
	jnot g0579(.din(w_n642_0[1]),.dout(n643),.clk(gclk));
	jor g0580(.dina(w_n631_0[0]),.dinb(w_n561_0[1]),.dout(n644),.clk(gclk));
	jxor g0581(.dina(w_n630_0[0]),.dinb(w_n561_0[0]),.dout(n645),.clk(gclk));
	jor g0582(.dina(n645),.dinb(w_n556_0[0]),.dout(n646),.clk(gclk));
	jand g0583(.dina(n646),.dinb(w_dff_B_wsW7Faqe1_1),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n648),.clk(gclk));
	jnot g0585(.din(n648),.dout(n649),.clk(gclk));
	jand g0586(.dina(w_n628_0[0]),.dinb(w_n566_0[0]),.dout(n650),.clk(gclk));
	jand g0587(.dina(w_n629_0[0]),.dinb(w_n563_0[0]),.dout(n651),.clk(gclk));
	jor g0588(.dina(n651),.dinb(w_dff_B_X9AQeE1F8_1),.dout(n652),.clk(gclk));
	jand g0589(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n653),.clk(gclk));
	jnot g0590(.din(n653),.dout(n654),.clk(gclk));
	jand g0591(.dina(w_n626_0[0]),.dinb(w_n571_0[0]),.dout(n655),.clk(gclk));
	jand g0592(.dina(w_n627_0[0]),.dinb(w_n568_0[0]),.dout(n656),.clk(gclk));
	jor g0593(.dina(n656),.dinb(w_dff_B_k3h97Z802_1),.dout(n657),.clk(gclk));
	jand g0594(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n658),.clk(gclk));
	jnot g0595(.din(n658),.dout(n659),.clk(gclk));
	jand g0596(.dina(w_n624_0[0]),.dinb(w_n576_0[0]),.dout(n660),.clk(gclk));
	jand g0597(.dina(w_n625_0[0]),.dinb(w_n573_0[0]),.dout(n661),.clk(gclk));
	jor g0598(.dina(n661),.dinb(w_dff_B_PxDcOGDe3_1),.dout(n662),.clk(gclk));
	jand g0599(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n663),.clk(gclk));
	jnot g0600(.din(n663),.dout(n664),.clk(gclk));
	jand g0601(.dina(w_n622_0[0]),.dinb(w_n581_0[0]),.dout(n665),.clk(gclk));
	jand g0602(.dina(w_n623_0[0]),.dinb(w_n578_0[0]),.dout(n666),.clk(gclk));
	jor g0603(.dina(n666),.dinb(w_dff_B_YElVKpLK0_1),.dout(n667),.clk(gclk));
	jand g0604(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n668),.clk(gclk));
	jnot g0605(.din(n668),.dout(n669),.clk(gclk));
	jand g0606(.dina(w_n620_0[0]),.dinb(w_n586_0[0]),.dout(n670),.clk(gclk));
	jand g0607(.dina(w_n621_0[0]),.dinb(w_n583_0[0]),.dout(n671),.clk(gclk));
	jor g0608(.dina(n671),.dinb(w_dff_B_aS9WQCEK1_1),.dout(n672),.clk(gclk));
	jand g0609(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_n618_0[0]),.dinb(w_n591_0[0]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n619_0[0]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jor g0613(.dina(n676),.dinb(w_dff_B_7p28RDIn2_1),.dout(n677),.clk(gclk));
	jand g0614(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n678),.clk(gclk));
	jnot g0615(.din(n678),.dout(n679),.clk(gclk));
	jand g0616(.dina(w_n616_0[0]),.dinb(w_n596_0[0]),.dout(n680),.clk(gclk));
	jand g0617(.dina(w_n617_0[0]),.dinb(w_n593_0[0]),.dout(n681),.clk(gclk));
	jor g0618(.dina(n681),.dinb(w_dff_B_Y9MhPSzk2_1),.dout(n682),.clk(gclk));
	jand g0619(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n683),.clk(gclk));
	jnot g0620(.din(n683),.dout(n684),.clk(gclk));
	jand g0621(.dina(w_n614_0[0]),.dinb(w_n602_0[0]),.dout(n685),.clk(gclk));
	jand g0622(.dina(w_n615_0[0]),.dinb(w_n598_0[0]),.dout(n686),.clk(gclk));
	jor g0623(.dina(n686),.dinb(w_dff_B_cAHDlMdl3_1),.dout(n687),.clk(gclk));
	jand g0624(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n688),.clk(gclk));
	jnot g0625(.din(n688),.dout(n689),.clk(gclk));
	jnot g0626(.din(w_n603_0[0]),.dout(n690),.clk(gclk));
	jnot g0627(.din(w_n613_0[0]),.dout(n691),.clk(gclk));
	jand g0628(.dina(n691),.dinb(w_dff_B_1BovEjzp0_1),.dout(n692),.clk(gclk));
	jor g0629(.dina(n692),.dinb(w_n611_0[0]),.dout(n693),.clk(gclk));
	jand g0630(.dina(w_G307gat_4[0]),.dinb(w_G188gat_6[2]),.dout(n694),.clk(gclk));
	jand g0631(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n695),.clk(gclk));
	jor g0632(.dina(w_n695_0[2]),.dinb(w_n606_0[0]),.dout(n696),.clk(gclk));
	jand g0633(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n697),.clk(gclk));
	jand g0634(.dina(w_n697_0[1]),.dinb(w_n604_0[0]),.dout(n698),.clk(gclk));
	jnot g0635(.din(w_n698_0[2]),.dout(n699),.clk(gclk));
	jand g0636(.dina(w_n699_0[1]),.dinb(w_dff_B_y9utSxa10_1),.dout(n700),.clk(gclk));
	jor g0637(.dina(n700),.dinb(w_n607_0[1]),.dout(n701),.clk(gclk));
	jnot g0638(.din(n701),.dout(n702),.clk(gclk));
	jand g0639(.dina(w_n699_0[0]),.dinb(w_n607_0[0]),.dout(n703),.clk(gclk));
	jor g0640(.dina(w_dff_B_FN4EiElf2_0),.dinb(w_n702_0[1]),.dout(n704),.clk(gclk));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_n694_0[1]),.dout(n705),.clk(gclk));
	jxor g0642(.dina(w_n705_0[1]),.dinb(w_n693_0[1]),.dout(n706),.clk(gclk));
	jxor g0643(.dina(w_n706_0[1]),.dinb(w_n689_0[1]),.dout(n707),.clk(gclk));
	jxor g0644(.dina(w_n707_0[1]),.dinb(w_n687_0[1]),.dout(n708),.clk(gclk));
	jxor g0645(.dina(w_n708_0[1]),.dinb(w_n684_0[1]),.dout(n709),.clk(gclk));
	jxor g0646(.dina(w_n709_0[1]),.dinb(w_n682_0[1]),.dout(n710),.clk(gclk));
	jxor g0647(.dina(w_n710_0[1]),.dinb(w_n679_0[1]),.dout(n711),.clk(gclk));
	jxor g0648(.dina(w_n711_0[1]),.dinb(w_n677_0[1]),.dout(n712),.clk(gclk));
	jxor g0649(.dina(w_n712_0[1]),.dinb(w_n674_0[1]),.dout(n713),.clk(gclk));
	jxor g0650(.dina(w_n713_0[1]),.dinb(w_n672_0[1]),.dout(n714),.clk(gclk));
	jxor g0651(.dina(w_n714_0[1]),.dinb(w_n669_0[1]),.dout(n715),.clk(gclk));
	jxor g0652(.dina(w_n715_0[1]),.dinb(w_n667_0[1]),.dout(n716),.clk(gclk));
	jxor g0653(.dina(w_n716_0[1]),.dinb(w_n664_0[1]),.dout(n717),.clk(gclk));
	jxor g0654(.dina(w_n717_0[1]),.dinb(w_n662_0[1]),.dout(n718),.clk(gclk));
	jxor g0655(.dina(w_n718_0[1]),.dinb(w_n659_0[1]),.dout(n719),.clk(gclk));
	jxor g0656(.dina(w_n719_0[1]),.dinb(w_n657_0[1]),.dout(n720),.clk(gclk));
	jxor g0657(.dina(w_n720_0[1]),.dinb(w_n654_0[1]),.dout(n721),.clk(gclk));
	jxor g0658(.dina(w_n721_0[1]),.dinb(w_n652_0[1]),.dout(n722),.clk(gclk));
	jxor g0659(.dina(w_n722_0[1]),.dinb(w_n649_0[1]),.dout(n723),.clk(gclk));
	jnot g0660(.din(w_n723_0[1]),.dout(n724),.clk(gclk));
	jxor g0661(.dina(w_n724_0[1]),.dinb(w_n647_0[2]),.dout(n725),.clk(gclk));
	jxor g0662(.dina(n725),.dinb(w_dff_B_XsTpae6H8_1),.dout(n726),.clk(gclk));
	jxor g0663(.dina(w_n726_0[1]),.dinb(w_n641_0[1]),.dout(n727),.clk(gclk));
	jxor g0664(.dina(w_n727_0[1]),.dinb(w_dff_B_r8jvjtir1_1),.dout(w_dff_A_WSl0EIyE8_2),.clk(gclk));
	jand g0665(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n729),.clk(gclk));
	jnot g0666(.din(w_n729_0[1]),.dout(n730),.clk(gclk));
	jnot g0667(.din(w_n726_0[0]),.dout(n731),.clk(gclk));
	jor g0668(.dina(n731),.dinb(w_n641_0[0]),.dout(n732),.clk(gclk));
	jor g0669(.dina(w_n727_0[0]),.dinb(w_n636_0[0]),.dout(n733),.clk(gclk));
	jand g0670(.dina(n733),.dinb(w_dff_B_jxu3HVWu3_1),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n735),.clk(gclk));
	jnot g0672(.din(w_n735_0[1]),.dout(n736),.clk(gclk));
	jor g0673(.dina(w_n724_0[0]),.dinb(w_n647_0[1]),.dout(n737),.clk(gclk));
	jxor g0674(.dina(w_n723_0[0]),.dinb(w_n647_0[0]),.dout(n738),.clk(gclk));
	jor g0675(.dina(n738),.dinb(w_n642_0[0]),.dout(n739),.clk(gclk));
	jand g0676(.dina(n739),.dinb(w_dff_B_3XNwPl930_1),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n741),.clk(gclk));
	jnot g0678(.din(n741),.dout(n742),.clk(gclk));
	jand g0679(.dina(w_n721_0[0]),.dinb(w_n652_0[0]),.dout(n743),.clk(gclk));
	jand g0680(.dina(w_n722_0[0]),.dinb(w_n649_0[0]),.dout(n744),.clk(gclk));
	jor g0681(.dina(n744),.dinb(w_dff_B_f52rD6cQ1_1),.dout(n745),.clk(gclk));
	jand g0682(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n746),.clk(gclk));
	jnot g0683(.din(n746),.dout(n747),.clk(gclk));
	jand g0684(.dina(w_n719_0[0]),.dinb(w_n657_0[0]),.dout(n748),.clk(gclk));
	jand g0685(.dina(w_n720_0[0]),.dinb(w_n654_0[0]),.dout(n749),.clk(gclk));
	jor g0686(.dina(n749),.dinb(w_dff_B_Jrwnh8Ov3_1),.dout(n750),.clk(gclk));
	jand g0687(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n751),.clk(gclk));
	jnot g0688(.din(n751),.dout(n752),.clk(gclk));
	jand g0689(.dina(w_n717_0[0]),.dinb(w_n662_0[0]),.dout(n753),.clk(gclk));
	jand g0690(.dina(w_n718_0[0]),.dinb(w_n659_0[0]),.dout(n754),.clk(gclk));
	jor g0691(.dina(n754),.dinb(w_dff_B_ZjSS2dJ77_1),.dout(n755),.clk(gclk));
	jand g0692(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n756),.clk(gclk));
	jnot g0693(.din(n756),.dout(n757),.clk(gclk));
	jand g0694(.dina(w_n715_0[0]),.dinb(w_n667_0[0]),.dout(n758),.clk(gclk));
	jand g0695(.dina(w_n716_0[0]),.dinb(w_n664_0[0]),.dout(n759),.clk(gclk));
	jor g0696(.dina(n759),.dinb(w_dff_B_TCeNeTdF2_1),.dout(n760),.clk(gclk));
	jand g0697(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n761),.clk(gclk));
	jnot g0698(.din(n761),.dout(n762),.clk(gclk));
	jand g0699(.dina(w_n713_0[0]),.dinb(w_n672_0[0]),.dout(n763),.clk(gclk));
	jand g0700(.dina(w_n714_0[0]),.dinb(w_n669_0[0]),.dout(n764),.clk(gclk));
	jor g0701(.dina(n764),.dinb(w_dff_B_NfzOU8uG7_1),.dout(n765),.clk(gclk));
	jand g0702(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(w_n711_0[0]),.dinb(w_n677_0[0]),.dout(n768),.clk(gclk));
	jand g0705(.dina(w_n712_0[0]),.dinb(w_n674_0[0]),.dout(n769),.clk(gclk));
	jor g0706(.dina(n769),.dinb(w_dff_B_at4LAabB1_1),.dout(n770),.clk(gclk));
	jand g0707(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n771),.clk(gclk));
	jnot g0708(.din(n771),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n709_0[0]),.dinb(w_n682_0[0]),.dout(n773),.clk(gclk));
	jand g0710(.dina(w_n710_0[0]),.dinb(w_n679_0[0]),.dout(n774),.clk(gclk));
	jor g0711(.dina(n774),.dinb(w_dff_B_EHm0L3KP9_1),.dout(n775),.clk(gclk));
	jand g0712(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n776),.clk(gclk));
	jnot g0713(.din(n776),.dout(n777),.clk(gclk));
	jand g0714(.dina(w_n707_0[0]),.dinb(w_n687_0[0]),.dout(n778),.clk(gclk));
	jand g0715(.dina(w_n708_0[0]),.dinb(w_n684_0[0]),.dout(n779),.clk(gclk));
	jor g0716(.dina(n779),.dinb(w_dff_B_GEBf26LN1_1),.dout(n780),.clk(gclk));
	jand g0717(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n781),.clk(gclk));
	jnot g0718(.din(n781),.dout(n782),.clk(gclk));
	jand g0719(.dina(w_n705_0[0]),.dinb(w_n693_0[0]),.dout(n783),.clk(gclk));
	jand g0720(.dina(w_n706_0[0]),.dinb(w_n689_0[0]),.dout(n784),.clk(gclk));
	jor g0721(.dina(n784),.dinb(w_dff_B_0sWTkjSX6_1),.dout(n785),.clk(gclk));
	jand g0722(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n786),.clk(gclk));
	jnot g0723(.din(n786),.dout(n787),.clk(gclk));
	jnot g0724(.din(w_n694_0[0]),.dout(n788),.clk(gclk));
	jnot g0725(.din(w_n704_0[0]),.dout(n789),.clk(gclk));
	jand g0726(.dina(n789),.dinb(w_dff_B_AbMIWrjY2_1),.dout(n790),.clk(gclk));
	jor g0727(.dina(n790),.dinb(w_n702_0[0]),.dout(n791),.clk(gclk));
	jand g0728(.dina(w_G307gat_3[2]),.dinb(w_G205gat_6[2]),.dout(n792),.clk(gclk));
	jand g0729(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n793),.clk(gclk));
	jor g0730(.dina(w_n793_0[1]),.dinb(w_n697_0[0]),.dout(n794),.clk(gclk));
	jand g0731(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n795),.clk(gclk));
	jand g0732(.dina(w_n795_0[1]),.dinb(w_n695_0[1]),.dout(n796),.clk(gclk));
	jnot g0733(.din(n796),.dout(n797),.clk(gclk));
	jand g0734(.dina(w_n797_0[2]),.dinb(w_dff_B_zrpbKDpH7_1),.dout(n798),.clk(gclk));
	jor g0735(.dina(n798),.dinb(w_n698_0[1]),.dout(n799),.clk(gclk));
	jnot g0736(.din(n799),.dout(n800),.clk(gclk));
	jand g0737(.dina(w_n797_0[1]),.dinb(w_n698_0[0]),.dout(n801),.clk(gclk));
	jor g0738(.dina(w_dff_B_d7N1ZYqq2_0),.dinb(w_n800_0[1]),.dout(n802),.clk(gclk));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n792_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_n791_0[1]),.dout(n804),.clk(gclk));
	jxor g0741(.dina(w_n804_0[1]),.dinb(w_n787_0[1]),.dout(n805),.clk(gclk));
	jxor g0742(.dina(w_n805_0[1]),.dinb(w_n785_0[1]),.dout(n806),.clk(gclk));
	jxor g0743(.dina(w_n806_0[1]),.dinb(w_n782_0[1]),.dout(n807),.clk(gclk));
	jxor g0744(.dina(w_n807_0[1]),.dinb(w_n780_0[1]),.dout(n808),.clk(gclk));
	jxor g0745(.dina(w_n808_0[1]),.dinb(w_n777_0[1]),.dout(n809),.clk(gclk));
	jxor g0746(.dina(w_n809_0[1]),.dinb(w_n775_0[1]),.dout(n810),.clk(gclk));
	jxor g0747(.dina(w_n810_0[1]),.dinb(w_n772_0[1]),.dout(n811),.clk(gclk));
	jxor g0748(.dina(w_n811_0[1]),.dinb(w_n770_0[1]),.dout(n812),.clk(gclk));
	jxor g0749(.dina(w_n812_0[1]),.dinb(w_n767_0[1]),.dout(n813),.clk(gclk));
	jxor g0750(.dina(w_n813_0[1]),.dinb(w_n765_0[1]),.dout(n814),.clk(gclk));
	jxor g0751(.dina(w_n814_0[1]),.dinb(w_n762_0[1]),.dout(n815),.clk(gclk));
	jxor g0752(.dina(w_n815_0[1]),.dinb(w_n760_0[1]),.dout(n816),.clk(gclk));
	jxor g0753(.dina(w_n816_0[1]),.dinb(w_n757_0[1]),.dout(n817),.clk(gclk));
	jxor g0754(.dina(w_n817_0[1]),.dinb(w_n755_0[1]),.dout(n818),.clk(gclk));
	jxor g0755(.dina(w_n818_0[1]),.dinb(w_n752_0[1]),.dout(n819),.clk(gclk));
	jxor g0756(.dina(w_n819_0[1]),.dinb(w_n750_0[1]),.dout(n820),.clk(gclk));
	jxor g0757(.dina(w_n820_0[1]),.dinb(w_n747_0[1]),.dout(n821),.clk(gclk));
	jxor g0758(.dina(w_n821_0[1]),.dinb(w_n745_0[1]),.dout(n822),.clk(gclk));
	jxor g0759(.dina(w_n822_0[1]),.dinb(w_n742_0[1]),.dout(n823),.clk(gclk));
	jnot g0760(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jxor g0761(.dina(w_n824_0[1]),.dinb(w_n740_0[2]),.dout(n825),.clk(gclk));
	jxor g0762(.dina(n825),.dinb(w_dff_B_APixYkF69_1),.dout(n826),.clk(gclk));
	jxor g0763(.dina(w_n826_0[1]),.dinb(w_n734_0[1]),.dout(n827),.clk(gclk));
	jxor g0764(.dina(w_n827_0[1]),.dinb(w_dff_B_eVLHXhof4_1),.dout(w_dff_A_ZhxLR9C13_2),.clk(gclk));
	jand g0765(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n829),.clk(gclk));
	jnot g0766(.din(w_n829_0[1]),.dout(n830),.clk(gclk));
	jnot g0767(.din(w_n826_0[0]),.dout(n831),.clk(gclk));
	jor g0768(.dina(n831),.dinb(w_n734_0[0]),.dout(n832),.clk(gclk));
	jor g0769(.dina(w_n827_0[0]),.dinb(w_n729_0[0]),.dout(n833),.clk(gclk));
	jand g0770(.dina(n833),.dinb(w_dff_B_WUFQEIHg0_1),.dout(n834),.clk(gclk));
	jand g0771(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n835),.clk(gclk));
	jor g0772(.dina(w_n824_0[0]),.dinb(w_n740_0[1]),.dout(n836),.clk(gclk));
	jxor g0773(.dina(w_n823_0[0]),.dinb(w_n740_0[0]),.dout(n837),.clk(gclk));
	jor g0774(.dina(n837),.dinb(w_n735_0[0]),.dout(n838),.clk(gclk));
	jand g0775(.dina(n838),.dinb(w_dff_B_HWRDEJIq8_1),.dout(n839),.clk(gclk));
	jand g0776(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n840),.clk(gclk));
	jnot g0777(.din(w_n840_0[1]),.dout(n841),.clk(gclk));
	jand g0778(.dina(w_n821_0[0]),.dinb(w_n745_0[0]),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n822_0[0]),.dinb(w_n742_0[0]),.dout(n843),.clk(gclk));
	jor g0780(.dina(n843),.dinb(w_dff_B_KML9lAql1_1),.dout(n844),.clk(gclk));
	jand g0781(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n845),.clk(gclk));
	jnot g0782(.din(n845),.dout(n846),.clk(gclk));
	jand g0783(.dina(w_n819_0[0]),.dinb(w_n750_0[0]),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n820_0[0]),.dinb(w_n747_0[0]),.dout(n848),.clk(gclk));
	jor g0785(.dina(n848),.dinb(w_dff_B_zyKCsiWb0_1),.dout(n849),.clk(gclk));
	jand g0786(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n850),.clk(gclk));
	jnot g0787(.din(n850),.dout(n851),.clk(gclk));
	jand g0788(.dina(w_n817_0[0]),.dinb(w_n755_0[0]),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n818_0[0]),.dinb(w_n752_0[0]),.dout(n853),.clk(gclk));
	jor g0790(.dina(n853),.dinb(w_dff_B_Dwps49C11_1),.dout(n854),.clk(gclk));
	jand g0791(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n855),.clk(gclk));
	jnot g0792(.din(n855),.dout(n856),.clk(gclk));
	jand g0793(.dina(w_n815_0[0]),.dinb(w_n760_0[0]),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n816_0[0]),.dinb(w_n757_0[0]),.dout(n858),.clk(gclk));
	jor g0795(.dina(n858),.dinb(w_dff_B_UDL5hThD3_1),.dout(n859),.clk(gclk));
	jand g0796(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n860),.clk(gclk));
	jnot g0797(.din(n860),.dout(n861),.clk(gclk));
	jand g0798(.dina(w_n813_0[0]),.dinb(w_n765_0[0]),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n814_0[0]),.dinb(w_n762_0[0]),.dout(n863),.clk(gclk));
	jor g0800(.dina(n863),.dinb(w_dff_B_Nv9sc4k00_1),.dout(n864),.clk(gclk));
	jand g0801(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n865),.clk(gclk));
	jnot g0802(.din(n865),.dout(n866),.clk(gclk));
	jand g0803(.dina(w_n811_0[0]),.dinb(w_n770_0[0]),.dout(n867),.clk(gclk));
	jand g0804(.dina(w_n812_0[0]),.dinb(w_n767_0[0]),.dout(n868),.clk(gclk));
	jor g0805(.dina(n868),.dinb(w_dff_B_5qkz8cg51_1),.dout(n869),.clk(gclk));
	jand g0806(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n870),.clk(gclk));
	jnot g0807(.din(n870),.dout(n871),.clk(gclk));
	jand g0808(.dina(w_n809_0[0]),.dinb(w_n775_0[0]),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_n810_0[0]),.dinb(w_n772_0[0]),.dout(n873),.clk(gclk));
	jor g0810(.dina(n873),.dinb(w_dff_B_7ThjlGih2_1),.dout(n874),.clk(gclk));
	jand g0811(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n875),.clk(gclk));
	jnot g0812(.din(n875),.dout(n876),.clk(gclk));
	jand g0813(.dina(w_n807_0[0]),.dinb(w_n780_0[0]),.dout(n877),.clk(gclk));
	jand g0814(.dina(w_n808_0[0]),.dinb(w_n777_0[0]),.dout(n878),.clk(gclk));
	jor g0815(.dina(n878),.dinb(w_dff_B_FCxt0qPm9_1),.dout(n879),.clk(gclk));
	jand g0816(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n880),.clk(gclk));
	jnot g0817(.din(n880),.dout(n881),.clk(gclk));
	jand g0818(.dina(w_n805_0[0]),.dinb(w_n785_0[0]),.dout(n882),.clk(gclk));
	jand g0819(.dina(w_n806_0[0]),.dinb(w_n782_0[0]),.dout(n883),.clk(gclk));
	jor g0820(.dina(n883),.dinb(w_dff_B_A83BQhCB9_1),.dout(n884),.clk(gclk));
	jand g0821(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n885),.clk(gclk));
	jnot g0822(.din(n885),.dout(n886),.clk(gclk));
	jand g0823(.dina(w_n803_0[0]),.dinb(w_n791_0[0]),.dout(n887),.clk(gclk));
	jand g0824(.dina(w_n804_0[0]),.dinb(w_n787_0[0]),.dout(n888),.clk(gclk));
	jor g0825(.dina(n888),.dinb(w_dff_B_EybfvUYZ7_1),.dout(n889),.clk(gclk));
	jand g0826(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n890),.clk(gclk));
	jnot g0827(.din(n890),.dout(n891),.clk(gclk));
	jnot g0828(.din(w_n792_0[0]),.dout(n892),.clk(gclk));
	jnot g0829(.din(w_n802_0[0]),.dout(n893),.clk(gclk));
	jand g0830(.dina(n893),.dinb(w_dff_B_ewdCX36A1_1),.dout(n894),.clk(gclk));
	jor g0831(.dina(n894),.dinb(w_n800_0[0]),.dout(n895),.clk(gclk));
	jand g0832(.dina(w_G307gat_3[1]),.dinb(w_G222gat_6[2]),.dout(n896),.clk(gclk));
	jnot g0833(.din(w_n795_0[0]),.dout(n897),.clk(gclk));
	jand g0834(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n898),.clk(gclk));
	jand g0835(.dina(w_n898_0[1]),.dinb(w_n897_0[1]),.dout(n899),.clk(gclk));
	jnot g0836(.din(n899),.dout(n900),.clk(gclk));
	jor g0837(.dina(w_n898_0[0]),.dinb(w_n897_0[0]),.dout(n901),.clk(gclk));
	jand g0838(.dina(w_n901_0[1]),.dinb(w_n797_0[0]),.dout(n902),.clk(gclk));
	jand g0839(.dina(n902),.dinb(n900),.dout(n903),.clk(gclk));
	jnot g0840(.din(w_n901_0[0]),.dout(n904),.clk(gclk));
	jand g0841(.dina(n904),.dinb(w_n695_0[0]),.dout(n905),.clk(gclk));
	jor g0842(.dina(n905),.dinb(w_n903_0[1]),.dout(n906),.clk(gclk));
	jxor g0843(.dina(w_n906_0[1]),.dinb(w_n896_0[1]),.dout(n907),.clk(gclk));
	jxor g0844(.dina(w_n907_0[1]),.dinb(w_n895_0[1]),.dout(n908),.clk(gclk));
	jxor g0845(.dina(w_n908_0[1]),.dinb(w_n891_0[1]),.dout(n909),.clk(gclk));
	jxor g0846(.dina(w_n909_0[1]),.dinb(w_n889_0[1]),.dout(n910),.clk(gclk));
	jxor g0847(.dina(w_n910_0[1]),.dinb(w_n886_0[1]),.dout(n911),.clk(gclk));
	jxor g0848(.dina(w_n911_0[1]),.dinb(w_n884_0[1]),.dout(n912),.clk(gclk));
	jxor g0849(.dina(w_n912_0[1]),.dinb(w_n881_0[1]),.dout(n913),.clk(gclk));
	jxor g0850(.dina(w_n913_0[1]),.dinb(w_n879_0[1]),.dout(n914),.clk(gclk));
	jxor g0851(.dina(w_n914_0[1]),.dinb(w_n876_0[1]),.dout(n915),.clk(gclk));
	jxor g0852(.dina(w_n915_0[1]),.dinb(w_n874_0[1]),.dout(n916),.clk(gclk));
	jxor g0853(.dina(w_n916_0[1]),.dinb(w_n871_0[1]),.dout(n917),.clk(gclk));
	jxor g0854(.dina(w_n917_0[1]),.dinb(w_n869_0[1]),.dout(n918),.clk(gclk));
	jxor g0855(.dina(w_n918_0[1]),.dinb(w_n866_0[1]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(w_n919_0[1]),.dinb(w_n864_0[1]),.dout(n920),.clk(gclk));
	jxor g0857(.dina(w_n920_0[1]),.dinb(w_n861_0[1]),.dout(n921),.clk(gclk));
	jxor g0858(.dina(w_n921_0[1]),.dinb(w_n859_0[1]),.dout(n922),.clk(gclk));
	jxor g0859(.dina(w_n922_0[1]),.dinb(w_n856_0[1]),.dout(n923),.clk(gclk));
	jxor g0860(.dina(w_n923_0[1]),.dinb(w_n854_0[1]),.dout(n924),.clk(gclk));
	jxor g0861(.dina(w_n924_0[1]),.dinb(w_n851_0[1]),.dout(n925),.clk(gclk));
	jxor g0862(.dina(w_n925_0[1]),.dinb(w_n849_0[1]),.dout(n926),.clk(gclk));
	jxor g0863(.dina(w_n926_0[1]),.dinb(w_n846_0[1]),.dout(n927),.clk(gclk));
	jxor g0864(.dina(w_n927_0[2]),.dinb(w_n844_0[2]),.dout(n928),.clk(gclk));
	jxor g0865(.dina(n928),.dinb(w_dff_B_sNHx9GFp7_1),.dout(n929),.clk(gclk));
	jxor g0866(.dina(w_n929_0[1]),.dinb(w_n839_0[1]),.dout(n930),.clk(gclk));
	jxor g0867(.dina(w_n930_0[1]),.dinb(w_n835_0[1]),.dout(n931),.clk(gclk));
	jxor g0868(.dina(w_n931_0[1]),.dinb(w_n834_0[1]),.dout(n932),.clk(gclk));
	jxor g0869(.dina(w_n932_0[1]),.dinb(w_dff_B_0R1rp4Wc2_1),.dout(w_dff_A_RiGNgq0v5_2),.clk(gclk));
	jnot g0870(.din(w_n931_0[0]),.dout(n934),.clk(gclk));
	jor g0871(.dina(n934),.dinb(w_n834_0[0]),.dout(n935),.clk(gclk));
	jor g0872(.dina(w_n932_0[0]),.dinb(w_n829_0[0]),.dout(n936),.clk(gclk));
	jand g0873(.dina(n936),.dinb(w_dff_B_byKfvmww9_1),.dout(n937),.clk(gclk));
	jand g0874(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n938),.clk(gclk));
	jnot g0875(.din(w_n929_0[0]),.dout(n939),.clk(gclk));
	jor g0876(.dina(n939),.dinb(w_n839_0[0]),.dout(n940),.clk(gclk));
	jor g0877(.dina(w_n930_0[0]),.dinb(w_n835_0[0]),.dout(n941),.clk(gclk));
	jand g0878(.dina(n941),.dinb(w_dff_B_9J9G5dhP3_1),.dout(n942),.clk(gclk));
	jand g0879(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n943),.clk(gclk));
	jand g0880(.dina(w_n927_0[1]),.dinb(w_n844_0[1]),.dout(n944),.clk(gclk));
	jnot g0881(.din(n944),.dout(n945),.clk(gclk));
	jnot g0882(.din(w_n927_0[0]),.dout(n946),.clk(gclk));
	jxor g0883(.dina(n946),.dinb(w_n844_0[0]),.dout(n947),.clk(gclk));
	jor g0884(.dina(n947),.dinb(w_n840_0[0]),.dout(n948),.clk(gclk));
	jand g0885(.dina(n948),.dinb(n945),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n950),.clk(gclk));
	jnot g0887(.din(n950),.dout(n951),.clk(gclk));
	jand g0888(.dina(w_n925_0[0]),.dinb(w_n849_0[0]),.dout(n952),.clk(gclk));
	jand g0889(.dina(w_n926_0[0]),.dinb(w_n846_0[0]),.dout(n953),.clk(gclk));
	jor g0890(.dina(n953),.dinb(w_dff_B_mILTqqt04_1),.dout(n954),.clk(gclk));
	jand g0891(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n955),.clk(gclk));
	jnot g0892(.din(n955),.dout(n956),.clk(gclk));
	jand g0893(.dina(w_n923_0[0]),.dinb(w_n854_0[0]),.dout(n957),.clk(gclk));
	jand g0894(.dina(w_n924_0[0]),.dinb(w_n851_0[0]),.dout(n958),.clk(gclk));
	jor g0895(.dina(n958),.dinb(w_dff_B_uw7NCiMR7_1),.dout(n959),.clk(gclk));
	jand g0896(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n960),.clk(gclk));
	jnot g0897(.din(n960),.dout(n961),.clk(gclk));
	jand g0898(.dina(w_n921_0[0]),.dinb(w_n859_0[0]),.dout(n962),.clk(gclk));
	jand g0899(.dina(w_n922_0[0]),.dinb(w_n856_0[0]),.dout(n963),.clk(gclk));
	jor g0900(.dina(n963),.dinb(w_dff_B_P0j1A7UR7_1),.dout(n964),.clk(gclk));
	jand g0901(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n965),.clk(gclk));
	jnot g0902(.din(n965),.dout(n966),.clk(gclk));
	jand g0903(.dina(w_n919_0[0]),.dinb(w_n864_0[0]),.dout(n967),.clk(gclk));
	jand g0904(.dina(w_n920_0[0]),.dinb(w_n861_0[0]),.dout(n968),.clk(gclk));
	jor g0905(.dina(n968),.dinb(w_dff_B_kCfO6Aus2_1),.dout(n969),.clk(gclk));
	jand g0906(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n970),.clk(gclk));
	jnot g0907(.din(n970),.dout(n971),.clk(gclk));
	jand g0908(.dina(w_n917_0[0]),.dinb(w_n869_0[0]),.dout(n972),.clk(gclk));
	jand g0909(.dina(w_n918_0[0]),.dinb(w_n866_0[0]),.dout(n973),.clk(gclk));
	jor g0910(.dina(n973),.dinb(w_dff_B_qwmlGLoC7_1),.dout(n974),.clk(gclk));
	jand g0911(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(w_n915_0[0]),.dinb(w_n874_0[0]),.dout(n977),.clk(gclk));
	jand g0914(.dina(w_n916_0[0]),.dinb(w_n871_0[0]),.dout(n978),.clk(gclk));
	jor g0915(.dina(n978),.dinb(w_dff_B_hxo8JQPg8_1),.dout(n979),.clk(gclk));
	jand g0916(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n980),.clk(gclk));
	jnot g0917(.din(n980),.dout(n981),.clk(gclk));
	jand g0918(.dina(w_n913_0[0]),.dinb(w_n879_0[0]),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_n914_0[0]),.dinb(w_n876_0[0]),.dout(n983),.clk(gclk));
	jor g0920(.dina(n983),.dinb(w_dff_B_DZRvO2GV2_1),.dout(n984),.clk(gclk));
	jand g0921(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n985),.clk(gclk));
	jnot g0922(.din(n985),.dout(n986),.clk(gclk));
	jand g0923(.dina(w_n911_0[0]),.dinb(w_n884_0[0]),.dout(n987),.clk(gclk));
	jand g0924(.dina(w_n912_0[0]),.dinb(w_n881_0[0]),.dout(n988),.clk(gclk));
	jor g0925(.dina(n988),.dinb(w_dff_B_UnQj650K1_1),.dout(n989),.clk(gclk));
	jand g0926(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n990),.clk(gclk));
	jnot g0927(.din(n990),.dout(n991),.clk(gclk));
	jand g0928(.dina(w_n909_0[0]),.dinb(w_n889_0[0]),.dout(n992),.clk(gclk));
	jand g0929(.dina(w_n910_0[0]),.dinb(w_n886_0[0]),.dout(n993),.clk(gclk));
	jor g0930(.dina(n993),.dinb(w_dff_B_SIoX6JBv3_1),.dout(n994),.clk(gclk));
	jand g0931(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n995),.clk(gclk));
	jnot g0932(.din(n995),.dout(n996),.clk(gclk));
	jand g0933(.dina(w_n907_0[0]),.dinb(w_n895_0[0]),.dout(n997),.clk(gclk));
	jand g0934(.dina(w_n908_0[0]),.dinb(w_n891_0[0]),.dout(n998),.clk(gclk));
	jor g0935(.dina(n998),.dinb(w_dff_B_aSMKxdg69_1),.dout(n999),.clk(gclk));
	jand g0936(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n1000),.clk(gclk));
	jnot g0937(.din(n1000),.dout(n1001),.clk(gclk));
	jnot g0938(.din(w_n896_0[0]),.dout(n1002),.clk(gclk));
	jnot g0939(.din(w_n906_0[0]),.dout(n1003),.clk(gclk));
	jand g0940(.dina(n1003),.dinb(w_dff_B_EWZpWhAQ7_1),.dout(n1004),.clk(gclk));
	jor g0941(.dina(n1004),.dinb(w_n903_0[0]),.dout(n1005),.clk(gclk));
	jand g0942(.dina(w_G307gat_3[0]),.dinb(w_G239gat_6[2]),.dout(n1006),.clk(gclk));
	jand g0943(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n1007),.clk(gclk));
	jnot g0944(.din(n1007),.dout(n1008),.clk(gclk));
	jor g0945(.dina(w_n1008_0[1]),.dinb(w_n793_0[0]),.dout(n1009),.clk(gclk));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n1006_0[1]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(w_n1010_0[1]),.dinb(w_n1005_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n1001_0[1]),.dout(n1012),.clk(gclk));
	jxor g0949(.dina(w_n1012_0[1]),.dinb(w_n999_0[1]),.dout(n1013),.clk(gclk));
	jxor g0950(.dina(w_n1013_0[1]),.dinb(w_n996_0[1]),.dout(n1014),.clk(gclk));
	jxor g0951(.dina(w_n1014_0[1]),.dinb(w_n994_0[1]),.dout(n1015),.clk(gclk));
	jxor g0952(.dina(w_n1015_0[1]),.dinb(w_n991_0[1]),.dout(n1016),.clk(gclk));
	jxor g0953(.dina(w_n1016_0[1]),.dinb(w_n989_0[1]),.dout(n1017),.clk(gclk));
	jxor g0954(.dina(w_n1017_0[1]),.dinb(w_n986_0[1]),.dout(n1018),.clk(gclk));
	jxor g0955(.dina(w_n1018_0[1]),.dinb(w_n984_0[1]),.dout(n1019),.clk(gclk));
	jxor g0956(.dina(w_n1019_0[1]),.dinb(w_n981_0[1]),.dout(n1020),.clk(gclk));
	jxor g0957(.dina(w_n1020_0[1]),.dinb(w_n979_0[1]),.dout(n1021),.clk(gclk));
	jxor g0958(.dina(w_n1021_0[1]),.dinb(w_n976_0[1]),.dout(n1022),.clk(gclk));
	jxor g0959(.dina(w_n1022_0[1]),.dinb(w_n974_0[1]),.dout(n1023),.clk(gclk));
	jxor g0960(.dina(w_n1023_0[1]),.dinb(w_n971_0[1]),.dout(n1024),.clk(gclk));
	jxor g0961(.dina(w_n1024_0[1]),.dinb(w_n969_0[1]),.dout(n1025),.clk(gclk));
	jxor g0962(.dina(w_n1025_0[1]),.dinb(w_n966_0[1]),.dout(n1026),.clk(gclk));
	jxor g0963(.dina(w_n1026_0[1]),.dinb(w_n964_0[1]),.dout(n1027),.clk(gclk));
	jxor g0964(.dina(w_n1027_0[1]),.dinb(w_n961_0[1]),.dout(n1028),.clk(gclk));
	jxor g0965(.dina(w_n1028_0[1]),.dinb(w_n959_0[1]),.dout(n1029),.clk(gclk));
	jxor g0966(.dina(w_n1029_0[1]),.dinb(w_n956_0[1]),.dout(n1030),.clk(gclk));
	jxor g0967(.dina(w_n1030_0[1]),.dinb(w_n954_0[1]),.dout(n1031),.clk(gclk));
	jxor g0968(.dina(w_n1031_0[1]),.dinb(w_n951_0[1]),.dout(n1032),.clk(gclk));
	jxor g0969(.dina(w_n1032_0[1]),.dinb(w_n949_0[1]),.dout(n1033),.clk(gclk));
	jxor g0970(.dina(w_n1033_0[1]),.dinb(w_n943_0[1]),.dout(n1034),.clk(gclk));
	jnot g0971(.din(w_n1034_0[1]),.dout(n1035),.clk(gclk));
	jxor g0972(.dina(w_n1035_0[1]),.dinb(w_n942_0[2]),.dout(n1036),.clk(gclk));
	jxor g0973(.dina(n1036),.dinb(w_n938_0[1]),.dout(n1037),.clk(gclk));
	jxor g0974(.dina(w_n1037_0[1]),.dinb(w_n937_0[1]),.dout(w_dff_A_YCRvBVIi5_2),.clk(gclk));
	jand g0975(.dina(w_n1037_0[0]),.dinb(w_n937_0[0]),.dout(n1039),.clk(gclk));
	jor g0976(.dina(w_n1035_0[0]),.dinb(w_n942_0[1]),.dout(n1040),.clk(gclk));
	jxor g0977(.dina(w_n1034_0[0]),.dinb(w_n942_0[0]),.dout(n1041),.clk(gclk));
	jor g0978(.dina(n1041),.dinb(w_n938_0[0]),.dout(n1042),.clk(gclk));
	jand g0979(.dina(n1042),.dinb(w_dff_B_rxFTLE6m4_1),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1044),.clk(gclk));
	jnot g0981(.din(w_n1032_0[0]),.dout(n1045),.clk(gclk));
	jor g0982(.dina(n1045),.dinb(w_n949_0[0]),.dout(n1046),.clk(gclk));
	jor g0983(.dina(w_n1033_0[0]),.dinb(w_n943_0[0]),.dout(n1047),.clk(gclk));
	jand g0984(.dina(n1047),.dinb(w_dff_B_UWPl9sBx1_1),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n1030_0[0]),.dinb(w_n954_0[0]),.dout(n1050),.clk(gclk));
	jand g0987(.dina(w_n1031_0[0]),.dinb(w_n951_0[0]),.dout(n1051),.clk(gclk));
	jor g0988(.dina(n1051),.dinb(w_dff_B_meIcJku66_1),.dout(n1052),.clk(gclk));
	jand g0989(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1053),.clk(gclk));
	jnot g0990(.din(n1053),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n1028_0[0]),.dinb(w_n959_0[0]),.dout(n1055),.clk(gclk));
	jand g0992(.dina(w_n1029_0[0]),.dinb(w_n956_0[0]),.dout(n1056),.clk(gclk));
	jor g0993(.dina(n1056),.dinb(w_dff_B_ECAasbK75_1),.dout(n1057),.clk(gclk));
	jand g0994(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1058),.clk(gclk));
	jnot g0995(.din(n1058),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n1026_0[0]),.dinb(w_n964_0[0]),.dout(n1060),.clk(gclk));
	jand g0997(.dina(w_n1027_0[0]),.dinb(w_n961_0[0]),.dout(n1061),.clk(gclk));
	jor g0998(.dina(n1061),.dinb(w_dff_B_5zfOOgKH1_1),.dout(n1062),.clk(gclk));
	jand g0999(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1063),.clk(gclk));
	jnot g1000(.din(n1063),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n1024_0[0]),.dinb(w_n969_0[0]),.dout(n1065),.clk(gclk));
	jand g1002(.dina(w_n1025_0[0]),.dinb(w_n966_0[0]),.dout(n1066),.clk(gclk));
	jor g1003(.dina(n1066),.dinb(w_dff_B_gKd82W6n2_1),.dout(n1067),.clk(gclk));
	jand g1004(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1068),.clk(gclk));
	jnot g1005(.din(n1068),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n1022_0[0]),.dinb(w_n974_0[0]),.dout(n1070),.clk(gclk));
	jand g1007(.dina(w_n1023_0[0]),.dinb(w_n971_0[0]),.dout(n1071),.clk(gclk));
	jor g1008(.dina(n1071),.dinb(w_dff_B_AWEkbpKd1_1),.dout(n1072),.clk(gclk));
	jand g1009(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1073),.clk(gclk));
	jnot g1010(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n1020_0[0]),.dinb(w_n979_0[0]),.dout(n1075),.clk(gclk));
	jand g1012(.dina(w_n1021_0[0]),.dinb(w_n976_0[0]),.dout(n1076),.clk(gclk));
	jor g1013(.dina(n1076),.dinb(w_dff_B_UXKY7mn06_1),.dout(n1077),.clk(gclk));
	jand g1014(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1078),.clk(gclk));
	jnot g1015(.din(n1078),.dout(n1079),.clk(gclk));
	jand g1016(.dina(w_n1018_0[0]),.dinb(w_n984_0[0]),.dout(n1080),.clk(gclk));
	jand g1017(.dina(w_n1019_0[0]),.dinb(w_n981_0[0]),.dout(n1081),.clk(gclk));
	jor g1018(.dina(n1081),.dinb(w_dff_B_pcewXHOL5_1),.dout(n1082),.clk(gclk));
	jand g1019(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1083),.clk(gclk));
	jnot g1020(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1021(.dina(w_n1016_0[0]),.dinb(w_n989_0[0]),.dout(n1085),.clk(gclk));
	jand g1022(.dina(w_n1017_0[0]),.dinb(w_n986_0[0]),.dout(n1086),.clk(gclk));
	jor g1023(.dina(n1086),.dinb(w_dff_B_ITjObB5K9_1),.dout(n1087),.clk(gclk));
	jand g1024(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1088),.clk(gclk));
	jnot g1025(.din(n1088),.dout(n1089),.clk(gclk));
	jand g1026(.dina(w_n1014_0[0]),.dinb(w_n994_0[0]),.dout(n1090),.clk(gclk));
	jand g1027(.dina(w_n1015_0[0]),.dinb(w_n991_0[0]),.dout(n1091),.clk(gclk));
	jor g1028(.dina(n1091),.dinb(w_dff_B_P3kYKh2x3_1),.dout(n1092),.clk(gclk));
	jand g1029(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1093),.clk(gclk));
	jnot g1030(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1031(.dina(w_n1012_0[0]),.dinb(w_n999_0[0]),.dout(n1095),.clk(gclk));
	jand g1032(.dina(w_n1013_0[0]),.dinb(w_n996_0[0]),.dout(n1096),.clk(gclk));
	jor g1033(.dina(n1096),.dinb(w_dff_B_9lRe7hy55_1),.dout(n1097),.clk(gclk));
	jand g1034(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1098),.clk(gclk));
	jnot g1035(.din(n1098),.dout(n1099),.clk(gclk));
	jand g1036(.dina(w_n1010_0[0]),.dinb(w_n1005_0[0]),.dout(n1100),.clk(gclk));
	jand g1037(.dina(w_n1011_0[0]),.dinb(w_n1001_0[0]),.dout(n1101),.clk(gclk));
	jor g1038(.dina(n1101),.dinb(w_dff_B_dGU27aM66_1),.dout(n1102),.clk(gclk));
	jand g1039(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1103),.clk(gclk));
	jand g1040(.dina(w_G307gat_2[2]),.dinb(w_G256gat_6[2]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(w_n1006_0[0]),.dout(n1105),.clk(gclk));
	jnot g1042(.din(w_n1009_0[0]),.dout(n1106),.clk(gclk));
	jand g1043(.dina(n1106),.dinb(w_dff_B_bNAI5svb2_1),.dout(n1107),.clk(gclk));
	jor g1044(.dina(n1107),.dinb(w_n1008_0[0]),.dout(n1108),.clk(gclk));
	jnot g1045(.din(n1108),.dout(n1109),.clk(gclk));
	jor g1046(.dina(w_n1109_0[1]),.dinb(w_dff_B_Ey840Zsi9_1),.dout(n1110),.clk(gclk));
	jand g1047(.dina(w_n1109_0[0]),.dinb(w_G307gat_2[1]),.dout(n1111),.clk(gclk));
	jnot g1048(.din(n1111),.dout(n1112),.clk(gclk));
	jand g1049(.dina(n1112),.dinb(w_n1110_0[1]),.dout(n1113),.clk(gclk));
	jnot g1050(.din(n1113),.dout(n1114),.clk(gclk));
	jxor g1051(.dina(w_n1114_0[1]),.dinb(w_n1103_0[1]),.dout(n1115),.clk(gclk));
	jxor g1052(.dina(w_n1115_0[1]),.dinb(w_n1102_0[1]),.dout(n1116),.clk(gclk));
	jxor g1053(.dina(w_n1116_0[1]),.dinb(w_n1099_0[1]),.dout(n1117),.clk(gclk));
	jxor g1054(.dina(w_n1117_0[1]),.dinb(w_n1097_0[1]),.dout(n1118),.clk(gclk));
	jxor g1055(.dina(w_n1118_0[1]),.dinb(w_n1094_0[1]),.dout(n1119),.clk(gclk));
	jxor g1056(.dina(w_n1119_0[1]),.dinb(w_n1092_0[1]),.dout(n1120),.clk(gclk));
	jxor g1057(.dina(w_n1120_0[1]),.dinb(w_n1089_0[1]),.dout(n1121),.clk(gclk));
	jxor g1058(.dina(w_n1121_0[1]),.dinb(w_n1087_0[1]),.dout(n1122),.clk(gclk));
	jxor g1059(.dina(w_n1122_0[1]),.dinb(w_n1084_0[1]),.dout(n1123),.clk(gclk));
	jxor g1060(.dina(w_n1123_0[1]),.dinb(w_n1082_0[1]),.dout(n1124),.clk(gclk));
	jxor g1061(.dina(w_n1124_0[1]),.dinb(w_n1079_0[1]),.dout(n1125),.clk(gclk));
	jxor g1062(.dina(w_n1125_0[1]),.dinb(w_n1077_0[1]),.dout(n1126),.clk(gclk));
	jxor g1063(.dina(w_n1126_0[1]),.dinb(w_n1074_0[1]),.dout(n1127),.clk(gclk));
	jxor g1064(.dina(w_n1127_0[1]),.dinb(w_n1072_0[1]),.dout(n1128),.clk(gclk));
	jxor g1065(.dina(w_n1128_0[1]),.dinb(w_n1069_0[1]),.dout(n1129),.clk(gclk));
	jxor g1066(.dina(w_n1129_0[1]),.dinb(w_n1067_0[1]),.dout(n1130),.clk(gclk));
	jxor g1067(.dina(w_n1130_0[1]),.dinb(w_n1064_0[1]),.dout(n1131),.clk(gclk));
	jxor g1068(.dina(w_n1131_0[1]),.dinb(w_n1062_0[1]),.dout(n1132),.clk(gclk));
	jxor g1069(.dina(w_n1132_0[1]),.dinb(w_n1059_0[1]),.dout(n1133),.clk(gclk));
	jxor g1070(.dina(w_n1133_0[1]),.dinb(w_n1057_0[1]),.dout(n1134),.clk(gclk));
	jxor g1071(.dina(w_n1134_0[1]),.dinb(w_n1054_0[1]),.dout(n1135),.clk(gclk));
	jxor g1072(.dina(w_n1135_0[1]),.dinb(w_n1052_0[1]),.dout(n1136),.clk(gclk));
	jnot g1073(.din(n1136),.dout(n1137),.clk(gclk));
	jxor g1074(.dina(w_n1137_0[1]),.dinb(w_n1049_0[1]),.dout(n1138),.clk(gclk));
	jxor g1075(.dina(w_n1138_0[1]),.dinb(w_n1048_0[1]),.dout(n1139),.clk(gclk));
	jxor g1076(.dina(w_n1139_0[1]),.dinb(w_n1044_0[1]),.dout(n1140),.clk(gclk));
	jxor g1077(.dina(w_n1140_0[1]),.dinb(w_n1043_0[1]),.dout(n1141),.clk(gclk));
	jnot g1078(.din(w_n1141_0[1]),.dout(n1142),.clk(gclk));
	jxor g1079(.dina(n1142),.dinb(w_n1039_0[1]),.dout(w_dff_A_3j1PEYfK3_2),.clk(gclk));
	jnot g1080(.din(w_n1140_0[0]),.dout(n1144),.clk(gclk));
	jor g1081(.dina(n1144),.dinb(w_n1043_0[0]),.dout(n1145),.clk(gclk));
	jor g1082(.dina(w_n1141_0[0]),.dinb(w_n1039_0[0]),.dout(n1146),.clk(gclk));
	jand g1083(.dina(n1146),.dinb(w_dff_B_jo2C4wSM4_1),.dout(n1147),.clk(gclk));
	jnot g1084(.din(w_n1138_0[0]),.dout(n1148),.clk(gclk));
	jor g1085(.dina(n1148),.dinb(w_n1048_0[0]),.dout(n1149),.clk(gclk));
	jor g1086(.dina(w_n1139_0[0]),.dinb(w_n1044_0[0]),.dout(n1150),.clk(gclk));
	jand g1087(.dina(n1150),.dinb(n1149),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1135_0[0]),.dinb(w_n1052_0[0]),.dout(n1153),.clk(gclk));
	jnot g1090(.din(n1153),.dout(n1154),.clk(gclk));
	jor g1091(.dina(w_n1137_0[0]),.dinb(w_n1049_0[0]),.dout(n1155),.clk(gclk));
	jand g1092(.dina(n1155),.dinb(w_dff_B_SnrhP7B65_1),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1157),.clk(gclk));
	jnot g1094(.din(n1157),.dout(n1158),.clk(gclk));
	jand g1095(.dina(w_n1133_0[0]),.dinb(w_n1057_0[0]),.dout(n1159),.clk(gclk));
	jand g1096(.dina(w_n1134_0[0]),.dinb(w_n1054_0[0]),.dout(n1160),.clk(gclk));
	jor g1097(.dina(n1160),.dinb(w_dff_B_pNGp6yFR8_1),.dout(n1161),.clk(gclk));
	jand g1098(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1162),.clk(gclk));
	jnot g1099(.din(n1162),.dout(n1163),.clk(gclk));
	jand g1100(.dina(w_n1131_0[0]),.dinb(w_n1062_0[0]),.dout(n1164),.clk(gclk));
	jand g1101(.dina(w_n1132_0[0]),.dinb(w_n1059_0[0]),.dout(n1165),.clk(gclk));
	jor g1102(.dina(n1165),.dinb(w_dff_B_tzPycaO79_1),.dout(n1166),.clk(gclk));
	jand g1103(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1167),.clk(gclk));
	jnot g1104(.din(n1167),.dout(n1168),.clk(gclk));
	jand g1105(.dina(w_n1129_0[0]),.dinb(w_n1067_0[0]),.dout(n1169),.clk(gclk));
	jand g1106(.dina(w_n1130_0[0]),.dinb(w_n1064_0[0]),.dout(n1170),.clk(gclk));
	jor g1107(.dina(n1170),.dinb(w_dff_B_h96iplJp8_1),.dout(n1171),.clk(gclk));
	jand g1108(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1172),.clk(gclk));
	jnot g1109(.din(n1172),.dout(n1173),.clk(gclk));
	jand g1110(.dina(w_n1127_0[0]),.dinb(w_n1072_0[0]),.dout(n1174),.clk(gclk));
	jand g1111(.dina(w_n1128_0[0]),.dinb(w_n1069_0[0]),.dout(n1175),.clk(gclk));
	jor g1112(.dina(n1175),.dinb(w_dff_B_gkznpBEf4_1),.dout(n1176),.clk(gclk));
	jand g1113(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1177),.clk(gclk));
	jnot g1114(.din(n1177),.dout(n1178),.clk(gclk));
	jand g1115(.dina(w_n1125_0[0]),.dinb(w_n1077_0[0]),.dout(n1179),.clk(gclk));
	jand g1116(.dina(w_n1126_0[0]),.dinb(w_n1074_0[0]),.dout(n1180),.clk(gclk));
	jor g1117(.dina(n1180),.dinb(w_dff_B_XgFFSGbv9_1),.dout(n1181),.clk(gclk));
	jand g1118(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1182),.clk(gclk));
	jnot g1119(.din(n1182),.dout(n1183),.clk(gclk));
	jand g1120(.dina(w_n1123_0[0]),.dinb(w_n1082_0[0]),.dout(n1184),.clk(gclk));
	jand g1121(.dina(w_n1124_0[0]),.dinb(w_n1079_0[0]),.dout(n1185),.clk(gclk));
	jor g1122(.dina(n1185),.dinb(w_dff_B_xYPBzUfi5_1),.dout(n1186),.clk(gclk));
	jand g1123(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1187),.clk(gclk));
	jnot g1124(.din(n1187),.dout(n1188),.clk(gclk));
	jand g1125(.dina(w_n1121_0[0]),.dinb(w_n1087_0[0]),.dout(n1189),.clk(gclk));
	jand g1126(.dina(w_n1122_0[0]),.dinb(w_n1084_0[0]),.dout(n1190),.clk(gclk));
	jor g1127(.dina(n1190),.dinb(w_dff_B_y1QTgYa17_1),.dout(n1191),.clk(gclk));
	jand g1128(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1192),.clk(gclk));
	jnot g1129(.din(n1192),.dout(n1193),.clk(gclk));
	jand g1130(.dina(w_n1119_0[0]),.dinb(w_n1092_0[0]),.dout(n1194),.clk(gclk));
	jand g1131(.dina(w_n1120_0[0]),.dinb(w_n1089_0[0]),.dout(n1195),.clk(gclk));
	jor g1132(.dina(n1195),.dinb(w_dff_B_Qjvy0QeU2_1),.dout(n1196),.clk(gclk));
	jand g1133(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1197),.clk(gclk));
	jnot g1134(.din(n1197),.dout(n1198),.clk(gclk));
	jand g1135(.dina(w_n1117_0[0]),.dinb(w_n1097_0[0]),.dout(n1199),.clk(gclk));
	jand g1136(.dina(w_n1118_0[0]),.dinb(w_n1094_0[0]),.dout(n1200),.clk(gclk));
	jor g1137(.dina(n1200),.dinb(w_dff_B_AINmtyNJ6_1),.dout(n1201),.clk(gclk));
	jand g1138(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jand g1140(.dina(w_n1115_0[0]),.dinb(w_n1102_0[0]),.dout(n1204),.clk(gclk));
	jand g1141(.dina(w_n1116_0[0]),.dinb(w_n1099_0[0]),.dout(n1205),.clk(gclk));
	jor g1142(.dina(n1205),.dinb(w_dff_B_XdgiEJGx6_1),.dout(n1206),.clk(gclk));
	jand g1143(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1207),.clk(gclk));
	jand g1144(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1208),.clk(gclk));
	jor g1145(.dina(w_n1114_0[0]),.dinb(w_n1103_0[0]),.dout(n1209),.clk(gclk));
	jand g1146(.dina(n1209),.dinb(w_n1110_0[0]),.dout(n1210),.clk(gclk));
	jxor g1147(.dina(w_n1210_0[1]),.dinb(w_n1208_0[1]),.dout(n1211),.clk(gclk));
	jnot g1148(.din(n1211),.dout(n1212),.clk(gclk));
	jxor g1149(.dina(w_n1212_0[1]),.dinb(w_n1207_0[1]),.dout(n1213),.clk(gclk));
	jxor g1150(.dina(w_n1213_0[1]),.dinb(w_n1206_0[1]),.dout(n1214),.clk(gclk));
	jxor g1151(.dina(w_n1214_0[1]),.dinb(w_n1203_0[1]),.dout(n1215),.clk(gclk));
	jxor g1152(.dina(w_n1215_0[1]),.dinb(w_n1201_0[1]),.dout(n1216),.clk(gclk));
	jxor g1153(.dina(w_n1216_0[1]),.dinb(w_n1198_0[1]),.dout(n1217),.clk(gclk));
	jxor g1154(.dina(w_n1217_0[1]),.dinb(w_n1196_0[1]),.dout(n1218),.clk(gclk));
	jxor g1155(.dina(w_n1218_0[1]),.dinb(w_n1193_0[1]),.dout(n1219),.clk(gclk));
	jxor g1156(.dina(w_n1219_0[1]),.dinb(w_n1191_0[1]),.dout(n1220),.clk(gclk));
	jxor g1157(.dina(w_n1220_0[1]),.dinb(w_n1188_0[1]),.dout(n1221),.clk(gclk));
	jxor g1158(.dina(w_n1221_0[1]),.dinb(w_n1186_0[1]),.dout(n1222),.clk(gclk));
	jxor g1159(.dina(w_n1222_0[1]),.dinb(w_n1183_0[1]),.dout(n1223),.clk(gclk));
	jxor g1160(.dina(w_n1223_0[1]),.dinb(w_n1181_0[1]),.dout(n1224),.clk(gclk));
	jxor g1161(.dina(w_n1224_0[1]),.dinb(w_n1178_0[1]),.dout(n1225),.clk(gclk));
	jxor g1162(.dina(w_n1225_0[1]),.dinb(w_n1176_0[1]),.dout(n1226),.clk(gclk));
	jxor g1163(.dina(w_n1226_0[1]),.dinb(w_n1173_0[1]),.dout(n1227),.clk(gclk));
	jxor g1164(.dina(w_n1227_0[1]),.dinb(w_n1171_0[1]),.dout(n1228),.clk(gclk));
	jxor g1165(.dina(w_n1228_0[1]),.dinb(w_n1168_0[1]),.dout(n1229),.clk(gclk));
	jxor g1166(.dina(w_n1229_0[1]),.dinb(w_n1166_0[1]),.dout(n1230),.clk(gclk));
	jxor g1167(.dina(w_n1230_0[1]),.dinb(w_n1163_0[1]),.dout(n1231),.clk(gclk));
	jxor g1168(.dina(w_n1231_0[1]),.dinb(w_n1161_0[1]),.dout(n1232),.clk(gclk));
	jxor g1169(.dina(w_n1232_0[1]),.dinb(w_n1158_0[1]),.dout(n1233),.clk(gclk));
	jnot g1170(.din(n1233),.dout(n1234),.clk(gclk));
	jxor g1171(.dina(w_n1234_0[1]),.dinb(w_n1156_0[1]),.dout(n1235),.clk(gclk));
	jnot g1172(.din(n1235),.dout(n1236),.clk(gclk));
	jxor g1173(.dina(w_n1236_0[1]),.dinb(w_n1152_0[1]),.dout(n1237),.clk(gclk));
	jxor g1174(.dina(w_n1237_0[1]),.dinb(w_n1151_0[1]),.dout(n1238),.clk(gclk));
	jnot g1175(.din(w_n1238_0[1]),.dout(n1239),.clk(gclk));
	jxor g1176(.dina(n1239),.dinb(w_n1147_0[1]),.dout(w_dff_A_qleo09kn4_2),.clk(gclk));
	jnot g1177(.din(w_n1237_0[0]),.dout(n1241),.clk(gclk));
	jor g1178(.dina(n1241),.dinb(w_n1151_0[0]),.dout(n1242),.clk(gclk));
	jor g1179(.dina(w_n1238_0[0]),.dinb(w_n1147_0[0]),.dout(n1243),.clk(gclk));
	jand g1180(.dina(n1243),.dinb(w_dff_B_2vRuOUkq5_1),.dout(n1244),.clk(gclk));
	jor g1181(.dina(w_n1234_0[0]),.dinb(w_n1156_0[0]),.dout(n1245),.clk(gclk));
	jor g1182(.dina(w_n1236_0[0]),.dinb(w_n1152_0[0]),.dout(n1246),.clk(gclk));
	jand g1183(.dina(n1246),.dinb(w_dff_B_RMb7G1lh3_1),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1231_0[0]),.dinb(w_n1161_0[0]),.dout(n1249),.clk(gclk));
	jand g1186(.dina(w_n1232_0[0]),.dinb(w_n1158_0[0]),.dout(n1250),.clk(gclk));
	jor g1187(.dina(n1250),.dinb(w_dff_B_xnCG75dL2_1),.dout(n1251),.clk(gclk));
	jand g1188(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1252),.clk(gclk));
	jnot g1189(.din(n1252),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1229_0[0]),.dinb(w_n1166_0[0]),.dout(n1254),.clk(gclk));
	jand g1191(.dina(w_n1230_0[0]),.dinb(w_n1163_0[0]),.dout(n1255),.clk(gclk));
	jor g1192(.dina(n1255),.dinb(w_dff_B_Ve6XuVT70_1),.dout(n1256),.clk(gclk));
	jand g1193(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1257),.clk(gclk));
	jnot g1194(.din(n1257),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1227_0[0]),.dinb(w_n1171_0[0]),.dout(n1259),.clk(gclk));
	jand g1196(.dina(w_n1228_0[0]),.dinb(w_n1168_0[0]),.dout(n1260),.clk(gclk));
	jor g1197(.dina(n1260),.dinb(w_dff_B_ZI9ttziG9_1),.dout(n1261),.clk(gclk));
	jand g1198(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1262),.clk(gclk));
	jnot g1199(.din(n1262),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1225_0[0]),.dinb(w_n1176_0[0]),.dout(n1264),.clk(gclk));
	jand g1201(.dina(w_n1226_0[0]),.dinb(w_n1173_0[0]),.dout(n1265),.clk(gclk));
	jor g1202(.dina(n1265),.dinb(w_dff_B_z5RhBe3P9_1),.dout(n1266),.clk(gclk));
	jand g1203(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1267),.clk(gclk));
	jnot g1204(.din(n1267),.dout(n1268),.clk(gclk));
	jand g1205(.dina(w_n1223_0[0]),.dinb(w_n1181_0[0]),.dout(n1269),.clk(gclk));
	jand g1206(.dina(w_n1224_0[0]),.dinb(w_n1178_0[0]),.dout(n1270),.clk(gclk));
	jor g1207(.dina(n1270),.dinb(w_dff_B_q3cqk8wI7_1),.dout(n1271),.clk(gclk));
	jand g1208(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1272),.clk(gclk));
	jnot g1209(.din(n1272),.dout(n1273),.clk(gclk));
	jand g1210(.dina(w_n1221_0[0]),.dinb(w_n1186_0[0]),.dout(n1274),.clk(gclk));
	jand g1211(.dina(w_n1222_0[0]),.dinb(w_n1183_0[0]),.dout(n1275),.clk(gclk));
	jor g1212(.dina(n1275),.dinb(w_dff_B_wagfIO683_1),.dout(n1276),.clk(gclk));
	jand g1213(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1277),.clk(gclk));
	jnot g1214(.din(n1277),.dout(n1278),.clk(gclk));
	jand g1215(.dina(w_n1219_0[0]),.dinb(w_n1191_0[0]),.dout(n1279),.clk(gclk));
	jand g1216(.dina(w_n1220_0[0]),.dinb(w_n1188_0[0]),.dout(n1280),.clk(gclk));
	jor g1217(.dina(n1280),.dinb(w_dff_B_Mhl3G5ff3_1),.dout(n1281),.clk(gclk));
	jand g1218(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1282),.clk(gclk));
	jnot g1219(.din(n1282),.dout(n1283),.clk(gclk));
	jand g1220(.dina(w_n1217_0[0]),.dinb(w_n1196_0[0]),.dout(n1284),.clk(gclk));
	jand g1221(.dina(w_n1218_0[0]),.dinb(w_n1193_0[0]),.dout(n1285),.clk(gclk));
	jor g1222(.dina(n1285),.dinb(w_dff_B_Mq3GucuZ0_1),.dout(n1286),.clk(gclk));
	jand g1223(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1287),.clk(gclk));
	jnot g1224(.din(n1287),.dout(n1288),.clk(gclk));
	jand g1225(.dina(w_n1215_0[0]),.dinb(w_n1201_0[0]),.dout(n1289),.clk(gclk));
	jand g1226(.dina(w_n1216_0[0]),.dinb(w_n1198_0[0]),.dout(n1290),.clk(gclk));
	jor g1227(.dina(n1290),.dinb(w_dff_B_3ek4XcaU4_1),.dout(n1291),.clk(gclk));
	jand g1228(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jand g1230(.dina(w_n1213_0[0]),.dinb(w_n1206_0[0]),.dout(n1294),.clk(gclk));
	jand g1231(.dina(w_n1214_0[0]),.dinb(w_n1203_0[0]),.dout(n1295),.clk(gclk));
	jor g1232(.dina(n1295),.dinb(w_dff_B_3kYMEyRn3_1),.dout(n1296),.clk(gclk));
	jand g1233(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1297),.clk(gclk));
	jand g1234(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1298),.clk(gclk));
	jor g1235(.dina(w_n1210_0[0]),.dinb(w_n1208_0[0]),.dout(n1299),.clk(gclk));
	jor g1236(.dina(w_n1212_0[0]),.dinb(w_n1207_0[0]),.dout(n1300),.clk(gclk));
	jand g1237(.dina(n1300),.dinb(w_dff_B_VUJ8kK6J4_1),.dout(n1301),.clk(gclk));
	jxor g1238(.dina(w_n1301_0[1]),.dinb(w_n1298_0[1]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(n1302),.dout(n1303),.clk(gclk));
	jxor g1240(.dina(w_n1303_0[1]),.dinb(w_n1297_0[1]),.dout(n1304),.clk(gclk));
	jxor g1241(.dina(w_n1304_0[1]),.dinb(w_n1296_0[1]),.dout(n1305),.clk(gclk));
	jxor g1242(.dina(w_n1305_0[1]),.dinb(w_n1293_0[1]),.dout(n1306),.clk(gclk));
	jxor g1243(.dina(w_n1306_0[1]),.dinb(w_n1291_0[1]),.dout(n1307),.clk(gclk));
	jxor g1244(.dina(w_n1307_0[1]),.dinb(w_n1288_0[1]),.dout(n1308),.clk(gclk));
	jxor g1245(.dina(w_n1308_0[1]),.dinb(w_n1286_0[1]),.dout(n1309),.clk(gclk));
	jxor g1246(.dina(w_n1309_0[1]),.dinb(w_n1283_0[1]),.dout(n1310),.clk(gclk));
	jxor g1247(.dina(w_n1310_0[1]),.dinb(w_n1281_0[1]),.dout(n1311),.clk(gclk));
	jxor g1248(.dina(w_n1311_0[1]),.dinb(w_n1278_0[1]),.dout(n1312),.clk(gclk));
	jxor g1249(.dina(w_n1312_0[1]),.dinb(w_n1276_0[1]),.dout(n1313),.clk(gclk));
	jxor g1250(.dina(w_n1313_0[1]),.dinb(w_n1273_0[1]),.dout(n1314),.clk(gclk));
	jxor g1251(.dina(w_n1314_0[1]),.dinb(w_n1271_0[1]),.dout(n1315),.clk(gclk));
	jxor g1252(.dina(w_n1315_0[1]),.dinb(w_n1268_0[1]),.dout(n1316),.clk(gclk));
	jxor g1253(.dina(w_n1316_0[1]),.dinb(w_n1266_0[1]),.dout(n1317),.clk(gclk));
	jxor g1254(.dina(w_n1317_0[1]),.dinb(w_n1263_0[1]),.dout(n1318),.clk(gclk));
	jxor g1255(.dina(w_n1318_0[1]),.dinb(w_n1261_0[1]),.dout(n1319),.clk(gclk));
	jxor g1256(.dina(w_n1319_0[1]),.dinb(w_n1258_0[1]),.dout(n1320),.clk(gclk));
	jxor g1257(.dina(w_n1320_0[1]),.dinb(w_n1256_0[1]),.dout(n1321),.clk(gclk));
	jxor g1258(.dina(w_n1321_0[1]),.dinb(w_n1253_0[1]),.dout(n1322),.clk(gclk));
	jxor g1259(.dina(w_n1322_0[1]),.dinb(w_n1251_0[1]),.dout(n1323),.clk(gclk));
	jnot g1260(.din(n1323),.dout(n1324),.clk(gclk));
	jxor g1261(.dina(w_n1324_0[1]),.dinb(w_n1248_0[1]),.dout(n1325),.clk(gclk));
	jxor g1262(.dina(w_n1325_0[1]),.dinb(w_n1247_0[1]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(w_n1326_0[1]),.dout(n1327),.clk(gclk));
	jxor g1264(.dina(w_dff_B_u11I65Fp8_0),.dinb(w_n1244_0[1]),.dout(w_dff_A_Mg1X7kYi3_2),.clk(gclk));
	jnot g1265(.din(w_n1325_0[0]),.dout(n1329),.clk(gclk));
	jor g1266(.dina(w_dff_B_urI1xCRA6_0),.dinb(w_n1247_0[0]),.dout(n1330),.clk(gclk));
	jor g1267(.dina(w_n1326_0[0]),.dinb(w_n1244_0[0]),.dout(n1331),.clk(gclk));
	jand g1268(.dina(n1331),.dinb(w_dff_B_GlvTNpIt5_1),.dout(n1332),.clk(gclk));
	jnot g1269(.din(w_n1251_0[0]),.dout(n1333),.clk(gclk));
	jnot g1270(.din(w_n1322_0[0]),.dout(n1334),.clk(gclk));
	jor g1271(.dina(w_dff_B_Ee5XMWLf9_0),.dinb(n1333),.dout(n1335),.clk(gclk));
	jor g1272(.dina(w_n1324_0[0]),.dinb(w_n1248_0[0]),.dout(n1336),.clk(gclk));
	jand g1273(.dina(n1336),.dinb(w_dff_B_2M717mWW2_1),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1320_0[0]),.dinb(w_n1256_0[0]),.dout(n1339),.clk(gclk));
	jand g1276(.dina(w_n1321_0[0]),.dinb(w_n1253_0[0]),.dout(n1340),.clk(gclk));
	jor g1277(.dina(n1340),.dinb(w_dff_B_j079FCM32_1),.dout(n1341),.clk(gclk));
	jand g1278(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1342),.clk(gclk));
	jnot g1279(.din(n1342),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1318_0[0]),.dinb(w_n1261_0[0]),.dout(n1344),.clk(gclk));
	jand g1281(.dina(w_n1319_0[0]),.dinb(w_n1258_0[0]),.dout(n1345),.clk(gclk));
	jor g1282(.dina(n1345),.dinb(w_dff_B_RZ68iGV39_1),.dout(n1346),.clk(gclk));
	jand g1283(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1347),.clk(gclk));
	jnot g1284(.din(n1347),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1316_0[0]),.dinb(w_n1266_0[0]),.dout(n1349),.clk(gclk));
	jand g1286(.dina(w_n1317_0[0]),.dinb(w_n1263_0[0]),.dout(n1350),.clk(gclk));
	jor g1287(.dina(n1350),.dinb(w_dff_B_HdN6e2QS5_1),.dout(n1351),.clk(gclk));
	jand g1288(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1352),.clk(gclk));
	jnot g1289(.din(n1352),.dout(n1353),.clk(gclk));
	jand g1290(.dina(w_n1314_0[0]),.dinb(w_n1271_0[0]),.dout(n1354),.clk(gclk));
	jand g1291(.dina(w_n1315_0[0]),.dinb(w_n1268_0[0]),.dout(n1355),.clk(gclk));
	jor g1292(.dina(n1355),.dinb(w_dff_B_ckoJgik34_1),.dout(n1356),.clk(gclk));
	jand g1293(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1357),.clk(gclk));
	jnot g1294(.din(n1357),.dout(n1358),.clk(gclk));
	jand g1295(.dina(w_n1312_0[0]),.dinb(w_n1276_0[0]),.dout(n1359),.clk(gclk));
	jand g1296(.dina(w_n1313_0[0]),.dinb(w_n1273_0[0]),.dout(n1360),.clk(gclk));
	jor g1297(.dina(n1360),.dinb(w_dff_B_r1QgCYWE8_1),.dout(n1361),.clk(gclk));
	jand g1298(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1362),.clk(gclk));
	jnot g1299(.din(n1362),.dout(n1363),.clk(gclk));
	jand g1300(.dina(w_n1310_0[0]),.dinb(w_n1281_0[0]),.dout(n1364),.clk(gclk));
	jand g1301(.dina(w_n1311_0[0]),.dinb(w_n1278_0[0]),.dout(n1365),.clk(gclk));
	jor g1302(.dina(n1365),.dinb(w_dff_B_bemMx2d96_1),.dout(n1366),.clk(gclk));
	jand g1303(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1367),.clk(gclk));
	jnot g1304(.din(n1367),.dout(n1368),.clk(gclk));
	jand g1305(.dina(w_n1308_0[0]),.dinb(w_n1286_0[0]),.dout(n1369),.clk(gclk));
	jand g1306(.dina(w_n1309_0[0]),.dinb(w_n1283_0[0]),.dout(n1370),.clk(gclk));
	jor g1307(.dina(n1370),.dinb(w_dff_B_lW6ZkaRh0_1),.dout(n1371),.clk(gclk));
	jand g1308(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1372),.clk(gclk));
	jnot g1309(.din(n1372),.dout(n1373),.clk(gclk));
	jand g1310(.dina(w_n1306_0[0]),.dinb(w_n1291_0[0]),.dout(n1374),.clk(gclk));
	jand g1311(.dina(w_n1307_0[0]),.dinb(w_n1288_0[0]),.dout(n1375),.clk(gclk));
	jor g1312(.dina(n1375),.dinb(w_dff_B_GJ7x2nk19_1),.dout(n1376),.clk(gclk));
	jand g1313(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jand g1315(.dina(w_n1304_0[0]),.dinb(w_n1296_0[0]),.dout(n1379),.clk(gclk));
	jand g1316(.dina(w_n1305_0[0]),.dinb(w_n1293_0[0]),.dout(n1380),.clk(gclk));
	jor g1317(.dina(n1380),.dinb(w_dff_B_qudcE3uE2_1),.dout(n1381),.clk(gclk));
	jand g1318(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1382),.clk(gclk));
	jand g1319(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1383),.clk(gclk));
	jor g1320(.dina(w_n1301_0[0]),.dinb(w_n1298_0[0]),.dout(n1384),.clk(gclk));
	jor g1321(.dina(w_n1303_0[0]),.dinb(w_n1297_0[0]),.dout(n1385),.clk(gclk));
	jand g1322(.dina(n1385),.dinb(w_dff_B_yvVQoDbq7_1),.dout(n1386),.clk(gclk));
	jxor g1323(.dina(w_n1386_0[1]),.dinb(w_n1383_0[1]),.dout(n1387),.clk(gclk));
	jnot g1324(.din(n1387),.dout(n1388),.clk(gclk));
	jxor g1325(.dina(w_n1388_0[1]),.dinb(w_n1382_0[1]),.dout(n1389),.clk(gclk));
	jxor g1326(.dina(w_n1389_0[1]),.dinb(w_n1381_0[1]),.dout(n1390),.clk(gclk));
	jxor g1327(.dina(w_n1390_0[1]),.dinb(w_n1378_0[1]),.dout(n1391),.clk(gclk));
	jxor g1328(.dina(w_n1391_0[1]),.dinb(w_n1376_0[1]),.dout(n1392),.clk(gclk));
	jxor g1329(.dina(w_n1392_0[1]),.dinb(w_n1373_0[1]),.dout(n1393),.clk(gclk));
	jxor g1330(.dina(w_n1393_0[1]),.dinb(w_n1371_0[1]),.dout(n1394),.clk(gclk));
	jxor g1331(.dina(w_n1394_0[1]),.dinb(w_n1368_0[1]),.dout(n1395),.clk(gclk));
	jxor g1332(.dina(w_n1395_0[1]),.dinb(w_n1366_0[1]),.dout(n1396),.clk(gclk));
	jxor g1333(.dina(w_n1396_0[1]),.dinb(w_n1363_0[1]),.dout(n1397),.clk(gclk));
	jxor g1334(.dina(w_n1397_0[1]),.dinb(w_n1361_0[1]),.dout(n1398),.clk(gclk));
	jxor g1335(.dina(w_n1398_0[1]),.dinb(w_n1358_0[1]),.dout(n1399),.clk(gclk));
	jxor g1336(.dina(w_n1399_0[1]),.dinb(w_n1356_0[1]),.dout(n1400),.clk(gclk));
	jxor g1337(.dina(w_n1400_0[1]),.dinb(w_n1353_0[1]),.dout(n1401),.clk(gclk));
	jxor g1338(.dina(w_n1401_0[1]),.dinb(w_n1351_0[1]),.dout(n1402),.clk(gclk));
	jxor g1339(.dina(w_n1402_0[1]),.dinb(w_n1348_0[1]),.dout(n1403),.clk(gclk));
	jxor g1340(.dina(w_n1403_0[1]),.dinb(w_n1346_0[1]),.dout(n1404),.clk(gclk));
	jxor g1341(.dina(w_n1404_0[1]),.dinb(w_n1343_0[1]),.dout(n1405),.clk(gclk));
	jxor g1342(.dina(w_n1405_0[1]),.dinb(w_n1341_0[1]),.dout(n1406),.clk(gclk));
	jnot g1343(.din(n1406),.dout(n1407),.clk(gclk));
	jxor g1344(.dina(w_n1407_0[1]),.dinb(w_n1338_0[1]),.dout(n1408),.clk(gclk));
	jnot g1345(.din(n1408),.dout(n1409),.clk(gclk));
	jxor g1346(.dina(w_n1409_0[1]),.dinb(w_n1337_0[1]),.dout(n1410),.clk(gclk));
	jxor g1347(.dina(w_n1410_0[1]),.dinb(w_n1332_0[1]),.dout(w_dff_A_CwhZzTZn9_2),.clk(gclk));
	jor g1348(.dina(w_n1409_0[0]),.dinb(w_n1337_0[0]),.dout(n1412),.clk(gclk));
	jnot g1349(.din(w_n1410_0[0]),.dout(n1413),.clk(gclk));
	jor g1350(.dina(w_dff_B_SJt7GV7E3_0),.dinb(w_n1332_0[0]),.dout(n1414),.clk(gclk));
	jand g1351(.dina(n1414),.dinb(w_dff_B_G3MHIb661_1),.dout(n1415),.clk(gclk));
	jnot g1352(.din(w_n1341_0[0]),.dout(n1416),.clk(gclk));
	jnot g1353(.din(w_n1405_0[0]),.dout(n1417),.clk(gclk));
	jor g1354(.dina(n1417),.dinb(n1416),.dout(n1418),.clk(gclk));
	jor g1355(.dina(w_n1407_0[0]),.dinb(w_n1338_0[0]),.dout(n1419),.clk(gclk));
	jand g1356(.dina(n1419),.dinb(w_dff_B_3bupPnHd6_1),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1403_0[0]),.dinb(w_n1346_0[0]),.dout(n1422),.clk(gclk));
	jand g1359(.dina(w_n1404_0[0]),.dinb(w_n1343_0[0]),.dout(n1423),.clk(gclk));
	jor g1360(.dina(n1423),.dinb(w_dff_B_gMOD04LK8_1),.dout(n1424),.clk(gclk));
	jand g1361(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1425),.clk(gclk));
	jnot g1362(.din(n1425),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1401_0[0]),.dinb(w_n1351_0[0]),.dout(n1427),.clk(gclk));
	jand g1364(.dina(w_n1402_0[0]),.dinb(w_n1348_0[0]),.dout(n1428),.clk(gclk));
	jor g1365(.dina(n1428),.dinb(w_dff_B_9e3ArnSM4_1),.dout(n1429),.clk(gclk));
	jand g1366(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1430),.clk(gclk));
	jnot g1367(.din(n1430),.dout(n1431),.clk(gclk));
	jand g1368(.dina(w_n1399_0[0]),.dinb(w_n1356_0[0]),.dout(n1432),.clk(gclk));
	jand g1369(.dina(w_n1400_0[0]),.dinb(w_n1353_0[0]),.dout(n1433),.clk(gclk));
	jor g1370(.dina(n1433),.dinb(w_dff_B_1JFEX1qQ4_1),.dout(n1434),.clk(gclk));
	jand g1371(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1435),.clk(gclk));
	jnot g1372(.din(n1435),.dout(n1436),.clk(gclk));
	jand g1373(.dina(w_n1397_0[0]),.dinb(w_n1361_0[0]),.dout(n1437),.clk(gclk));
	jand g1374(.dina(w_n1398_0[0]),.dinb(w_n1358_0[0]),.dout(n1438),.clk(gclk));
	jor g1375(.dina(n1438),.dinb(w_dff_B_3ivT3rTn6_1),.dout(n1439),.clk(gclk));
	jand g1376(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1440),.clk(gclk));
	jnot g1377(.din(n1440),.dout(n1441),.clk(gclk));
	jand g1378(.dina(w_n1395_0[0]),.dinb(w_n1366_0[0]),.dout(n1442),.clk(gclk));
	jand g1379(.dina(w_n1396_0[0]),.dinb(w_n1363_0[0]),.dout(n1443),.clk(gclk));
	jor g1380(.dina(n1443),.dinb(w_dff_B_6TwkF4Yo1_1),.dout(n1444),.clk(gclk));
	jand g1381(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1445),.clk(gclk));
	jnot g1382(.din(n1445),.dout(n1446),.clk(gclk));
	jand g1383(.dina(w_n1393_0[0]),.dinb(w_n1371_0[0]),.dout(n1447),.clk(gclk));
	jand g1384(.dina(w_n1394_0[0]),.dinb(w_n1368_0[0]),.dout(n1448),.clk(gclk));
	jor g1385(.dina(n1448),.dinb(w_dff_B_t0a1Cb0x2_1),.dout(n1449),.clk(gclk));
	jand g1386(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1450),.clk(gclk));
	jnot g1387(.din(n1450),.dout(n1451),.clk(gclk));
	jand g1388(.dina(w_n1391_0[0]),.dinb(w_n1376_0[0]),.dout(n1452),.clk(gclk));
	jand g1389(.dina(w_n1392_0[0]),.dinb(w_n1373_0[0]),.dout(n1453),.clk(gclk));
	jor g1390(.dina(n1453),.dinb(w_dff_B_oNsStTFp5_1),.dout(n1454),.clk(gclk));
	jand g1391(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1455),.clk(gclk));
	jnot g1392(.din(n1455),.dout(n1456),.clk(gclk));
	jand g1393(.dina(w_n1389_0[0]),.dinb(w_n1381_0[0]),.dout(n1457),.clk(gclk));
	jand g1394(.dina(w_n1390_0[0]),.dinb(w_n1378_0[0]),.dout(n1458),.clk(gclk));
	jor g1395(.dina(n1458),.dinb(w_dff_B_0k0xiUEN0_1),.dout(n1459),.clk(gclk));
	jand g1396(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1460),.clk(gclk));
	jand g1397(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1461),.clk(gclk));
	jor g1398(.dina(w_n1386_0[0]),.dinb(w_n1383_0[0]),.dout(n1462),.clk(gclk));
	jor g1399(.dina(w_n1388_0[0]),.dinb(w_n1382_0[0]),.dout(n1463),.clk(gclk));
	jand g1400(.dina(n1463),.dinb(w_dff_B_CzlX2EJb3_1),.dout(n1464),.clk(gclk));
	jxor g1401(.dina(w_n1464_0[1]),.dinb(w_n1461_0[1]),.dout(n1465),.clk(gclk));
	jnot g1402(.din(n1465),.dout(n1466),.clk(gclk));
	jxor g1403(.dina(w_n1466_0[1]),.dinb(w_n1460_0[1]),.dout(n1467),.clk(gclk));
	jxor g1404(.dina(w_n1467_0[1]),.dinb(w_n1459_0[1]),.dout(n1468),.clk(gclk));
	jxor g1405(.dina(w_n1468_0[1]),.dinb(w_n1456_0[1]),.dout(n1469),.clk(gclk));
	jxor g1406(.dina(w_n1469_0[1]),.dinb(w_n1454_0[1]),.dout(n1470),.clk(gclk));
	jxor g1407(.dina(w_n1470_0[1]),.dinb(w_n1451_0[1]),.dout(n1471),.clk(gclk));
	jxor g1408(.dina(w_n1471_0[1]),.dinb(w_n1449_0[1]),.dout(n1472),.clk(gclk));
	jxor g1409(.dina(w_n1472_0[1]),.dinb(w_n1446_0[1]),.dout(n1473),.clk(gclk));
	jxor g1410(.dina(w_n1473_0[1]),.dinb(w_n1444_0[1]),.dout(n1474),.clk(gclk));
	jxor g1411(.dina(w_n1474_0[1]),.dinb(w_n1441_0[1]),.dout(n1475),.clk(gclk));
	jxor g1412(.dina(w_n1475_0[1]),.dinb(w_n1439_0[1]),.dout(n1476),.clk(gclk));
	jxor g1413(.dina(w_n1476_0[1]),.dinb(w_n1436_0[1]),.dout(n1477),.clk(gclk));
	jxor g1414(.dina(w_n1477_0[1]),.dinb(w_n1434_0[1]),.dout(n1478),.clk(gclk));
	jxor g1415(.dina(w_n1478_0[1]),.dinb(w_n1431_0[1]),.dout(n1479),.clk(gclk));
	jxor g1416(.dina(w_n1479_0[1]),.dinb(w_n1429_0[1]),.dout(n1480),.clk(gclk));
	jxor g1417(.dina(w_n1480_0[1]),.dinb(w_n1426_0[1]),.dout(n1481),.clk(gclk));
	jxor g1418(.dina(w_n1481_0[1]),.dinb(w_n1424_0[1]),.dout(n1482),.clk(gclk));
	jnot g1419(.din(n1482),.dout(n1483),.clk(gclk));
	jxor g1420(.dina(w_n1483_0[1]),.dinb(w_n1421_0[1]),.dout(n1484),.clk(gclk));
	jnot g1421(.din(n1484),.dout(n1485),.clk(gclk));
	jxor g1422(.dina(w_n1485_0[1]),.dinb(w_n1420_0[1]),.dout(n1486),.clk(gclk));
	jxor g1423(.dina(w_n1486_0[1]),.dinb(w_n1415_0[1]),.dout(w_dff_A_6Ai86vBq2_2),.clk(gclk));
	jor g1424(.dina(w_n1485_0[0]),.dinb(w_n1420_0[0]),.dout(n1488),.clk(gclk));
	jnot g1425(.din(w_n1486_0[0]),.dout(n1489),.clk(gclk));
	jor g1426(.dina(w_dff_B_l8h2kqKv1_0),.dinb(w_n1415_0[0]),.dout(n1490),.clk(gclk));
	jand g1427(.dina(n1490),.dinb(w_dff_B_PspZc4QJ1_1),.dout(n1491),.clk(gclk));
	jnot g1428(.din(w_n1424_0[0]),.dout(n1492),.clk(gclk));
	jnot g1429(.din(w_n1481_0[0]),.dout(n1493),.clk(gclk));
	jor g1430(.dina(n1493),.dinb(n1492),.dout(n1494),.clk(gclk));
	jor g1431(.dina(w_n1483_0[0]),.dinb(w_n1421_0[0]),.dout(n1495),.clk(gclk));
	jand g1432(.dina(n1495),.dinb(w_dff_B_ldfrfag78_1),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1479_0[0]),.dinb(w_n1429_0[0]),.dout(n1498),.clk(gclk));
	jand g1435(.dina(w_n1480_0[0]),.dinb(w_n1426_0[0]),.dout(n1499),.clk(gclk));
	jor g1436(.dina(n1499),.dinb(w_dff_B_pVRMKH112_1),.dout(n1500),.clk(gclk));
	jand g1437(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1501),.clk(gclk));
	jnot g1438(.din(n1501),.dout(n1502),.clk(gclk));
	jand g1439(.dina(w_n1477_0[0]),.dinb(w_n1434_0[0]),.dout(n1503),.clk(gclk));
	jand g1440(.dina(w_n1478_0[0]),.dinb(w_n1431_0[0]),.dout(n1504),.clk(gclk));
	jor g1441(.dina(n1504),.dinb(w_dff_B_XiSKkmLA7_1),.dout(n1505),.clk(gclk));
	jand g1442(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1506),.clk(gclk));
	jnot g1443(.din(n1506),.dout(n1507),.clk(gclk));
	jand g1444(.dina(w_n1475_0[0]),.dinb(w_n1439_0[0]),.dout(n1508),.clk(gclk));
	jand g1445(.dina(w_n1476_0[0]),.dinb(w_n1436_0[0]),.dout(n1509),.clk(gclk));
	jor g1446(.dina(n1509),.dinb(w_dff_B_K41MyTbU4_1),.dout(n1510),.clk(gclk));
	jand g1447(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1511),.clk(gclk));
	jnot g1448(.din(n1511),.dout(n1512),.clk(gclk));
	jand g1449(.dina(w_n1473_0[0]),.dinb(w_n1444_0[0]),.dout(n1513),.clk(gclk));
	jand g1450(.dina(w_n1474_0[0]),.dinb(w_n1441_0[0]),.dout(n1514),.clk(gclk));
	jor g1451(.dina(n1514),.dinb(w_dff_B_dEwrKoGB5_1),.dout(n1515),.clk(gclk));
	jand g1452(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1516),.clk(gclk));
	jnot g1453(.din(n1516),.dout(n1517),.clk(gclk));
	jand g1454(.dina(w_n1471_0[0]),.dinb(w_n1449_0[0]),.dout(n1518),.clk(gclk));
	jand g1455(.dina(w_n1472_0[0]),.dinb(w_n1446_0[0]),.dout(n1519),.clk(gclk));
	jor g1456(.dina(n1519),.dinb(w_dff_B_ojVnhXCC2_1),.dout(n1520),.clk(gclk));
	jand g1457(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1521),.clk(gclk));
	jnot g1458(.din(n1521),.dout(n1522),.clk(gclk));
	jand g1459(.dina(w_n1469_0[0]),.dinb(w_n1454_0[0]),.dout(n1523),.clk(gclk));
	jand g1460(.dina(w_n1470_0[0]),.dinb(w_n1451_0[0]),.dout(n1524),.clk(gclk));
	jor g1461(.dina(n1524),.dinb(w_dff_B_9L9nGFxd7_1),.dout(n1525),.clk(gclk));
	jand g1462(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1526),.clk(gclk));
	jnot g1463(.din(n1526),.dout(n1527),.clk(gclk));
	jand g1464(.dina(w_n1467_0[0]),.dinb(w_n1459_0[0]),.dout(n1528),.clk(gclk));
	jand g1465(.dina(w_n1468_0[0]),.dinb(w_n1456_0[0]),.dout(n1529),.clk(gclk));
	jor g1466(.dina(n1529),.dinb(w_dff_B_LWNVmBBi8_1),.dout(n1530),.clk(gclk));
	jand g1467(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1531),.clk(gclk));
	jand g1468(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1532),.clk(gclk));
	jor g1469(.dina(w_n1464_0[0]),.dinb(w_n1461_0[0]),.dout(n1533),.clk(gclk));
	jor g1470(.dina(w_n1466_0[0]),.dinb(w_n1460_0[0]),.dout(n1534),.clk(gclk));
	jand g1471(.dina(n1534),.dinb(w_dff_B_4Q00MYR71_1),.dout(n1535),.clk(gclk));
	jxor g1472(.dina(w_n1535_0[1]),.dinb(w_n1532_0[1]),.dout(n1536),.clk(gclk));
	jnot g1473(.din(n1536),.dout(n1537),.clk(gclk));
	jxor g1474(.dina(w_n1537_0[1]),.dinb(w_n1531_0[1]),.dout(n1538),.clk(gclk));
	jxor g1475(.dina(w_n1538_0[1]),.dinb(w_n1530_0[1]),.dout(n1539),.clk(gclk));
	jxor g1476(.dina(w_n1539_0[1]),.dinb(w_n1527_0[1]),.dout(n1540),.clk(gclk));
	jxor g1477(.dina(w_n1540_0[1]),.dinb(w_n1525_0[1]),.dout(n1541),.clk(gclk));
	jxor g1478(.dina(w_n1541_0[1]),.dinb(w_n1522_0[1]),.dout(n1542),.clk(gclk));
	jxor g1479(.dina(w_n1542_0[1]),.dinb(w_n1520_0[1]),.dout(n1543),.clk(gclk));
	jxor g1480(.dina(w_n1543_0[1]),.dinb(w_n1517_0[1]),.dout(n1544),.clk(gclk));
	jxor g1481(.dina(w_n1544_0[1]),.dinb(w_n1515_0[1]),.dout(n1545),.clk(gclk));
	jxor g1482(.dina(w_n1545_0[1]),.dinb(w_n1512_0[1]),.dout(n1546),.clk(gclk));
	jxor g1483(.dina(w_n1546_0[1]),.dinb(w_n1510_0[1]),.dout(n1547),.clk(gclk));
	jxor g1484(.dina(w_n1547_0[1]),.dinb(w_n1507_0[1]),.dout(n1548),.clk(gclk));
	jxor g1485(.dina(w_n1548_0[1]),.dinb(w_n1505_0[1]),.dout(n1549),.clk(gclk));
	jxor g1486(.dina(w_n1549_0[1]),.dinb(w_n1502_0[1]),.dout(n1550),.clk(gclk));
	jxor g1487(.dina(w_n1550_0[1]),.dinb(w_n1500_0[1]),.dout(n1551),.clk(gclk));
	jnot g1488(.din(n1551),.dout(n1552),.clk(gclk));
	jxor g1489(.dina(w_n1552_0[1]),.dinb(w_n1497_0[1]),.dout(n1553),.clk(gclk));
	jnot g1490(.din(n1553),.dout(n1554),.clk(gclk));
	jxor g1491(.dina(w_n1554_0[1]),.dinb(w_n1496_0[1]),.dout(n1555),.clk(gclk));
	jxor g1492(.dina(w_n1555_0[1]),.dinb(w_n1491_0[1]),.dout(w_dff_A_L32hW2LS1_2),.clk(gclk));
	jor g1493(.dina(w_n1554_0[0]),.dinb(w_n1496_0[0]),.dout(n1557),.clk(gclk));
	jnot g1494(.din(w_n1555_0[0]),.dout(n1558),.clk(gclk));
	jor g1495(.dina(w_dff_B_vDfTjoF11_0),.dinb(w_n1491_0[0]),.dout(n1559),.clk(gclk));
	jand g1496(.dina(n1559),.dinb(w_dff_B_a8uOOsQh7_1),.dout(n1560),.clk(gclk));
	jnot g1497(.din(w_n1500_0[0]),.dout(n1561),.clk(gclk));
	jnot g1498(.din(w_n1550_0[0]),.dout(n1562),.clk(gclk));
	jor g1499(.dina(w_dff_B_rSxV2MYi3_0),.dinb(n1561),.dout(n1563),.clk(gclk));
	jor g1500(.dina(w_n1552_0[0]),.dinb(w_n1497_0[0]),.dout(n1564),.clk(gclk));
	jand g1501(.dina(n1564),.dinb(w_dff_B_dNZdGybo7_1),.dout(n1565),.clk(gclk));
	jand g1502(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1566),.clk(gclk));
	jand g1503(.dina(w_n1548_0[0]),.dinb(w_n1505_0[0]),.dout(n1567),.clk(gclk));
	jand g1504(.dina(w_n1549_0[0]),.dinb(w_n1502_0[0]),.dout(n1568),.clk(gclk));
	jor g1505(.dina(n1568),.dinb(w_dff_B_rwbfXufI7_1),.dout(n1569),.clk(gclk));
	jand g1506(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1570),.clk(gclk));
	jnot g1507(.din(n1570),.dout(n1571),.clk(gclk));
	jand g1508(.dina(w_n1546_0[0]),.dinb(w_n1510_0[0]),.dout(n1572),.clk(gclk));
	jand g1509(.dina(w_n1547_0[0]),.dinb(w_n1507_0[0]),.dout(n1573),.clk(gclk));
	jor g1510(.dina(n1573),.dinb(w_dff_B_pagIvr6A9_1),.dout(n1574),.clk(gclk));
	jand g1511(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1575),.clk(gclk));
	jnot g1512(.din(n1575),.dout(n1576),.clk(gclk));
	jand g1513(.dina(w_n1544_0[0]),.dinb(w_n1515_0[0]),.dout(n1577),.clk(gclk));
	jand g1514(.dina(w_n1545_0[0]),.dinb(w_n1512_0[0]),.dout(n1578),.clk(gclk));
	jor g1515(.dina(n1578),.dinb(w_dff_B_WXGUjXj40_1),.dout(n1579),.clk(gclk));
	jand g1516(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1580),.clk(gclk));
	jnot g1517(.din(n1580),.dout(n1581),.clk(gclk));
	jand g1518(.dina(w_n1542_0[0]),.dinb(w_n1520_0[0]),.dout(n1582),.clk(gclk));
	jand g1519(.dina(w_n1543_0[0]),.dinb(w_n1517_0[0]),.dout(n1583),.clk(gclk));
	jor g1520(.dina(n1583),.dinb(w_dff_B_OAaZjvPj1_1),.dout(n1584),.clk(gclk));
	jand g1521(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1585),.clk(gclk));
	jnot g1522(.din(n1585),.dout(n1586),.clk(gclk));
	jand g1523(.dina(w_n1540_0[0]),.dinb(w_n1525_0[0]),.dout(n1587),.clk(gclk));
	jand g1524(.dina(w_n1541_0[0]),.dinb(w_n1522_0[0]),.dout(n1588),.clk(gclk));
	jor g1525(.dina(n1588),.dinb(w_dff_B_h6vcaayM6_1),.dout(n1589),.clk(gclk));
	jand g1526(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1590),.clk(gclk));
	jnot g1527(.din(n1590),.dout(n1591),.clk(gclk));
	jand g1528(.dina(w_n1538_0[0]),.dinb(w_n1530_0[0]),.dout(n1592),.clk(gclk));
	jand g1529(.dina(w_n1539_0[0]),.dinb(w_n1527_0[0]),.dout(n1593),.clk(gclk));
	jor g1530(.dina(n1593),.dinb(w_dff_B_bBKY3IsN3_1),.dout(n1594),.clk(gclk));
	jand g1531(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1595),.clk(gclk));
	jand g1532(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1596),.clk(gclk));
	jor g1533(.dina(w_n1535_0[0]),.dinb(w_n1532_0[0]),.dout(n1597),.clk(gclk));
	jor g1534(.dina(w_n1537_0[0]),.dinb(w_n1531_0[0]),.dout(n1598),.clk(gclk));
	jand g1535(.dina(n1598),.dinb(w_dff_B_p0m5Rv4t8_1),.dout(n1599),.clk(gclk));
	jxor g1536(.dina(w_n1599_0[1]),.dinb(w_n1596_0[1]),.dout(n1600),.clk(gclk));
	jnot g1537(.din(n1600),.dout(n1601),.clk(gclk));
	jxor g1538(.dina(w_n1601_0[1]),.dinb(w_n1595_0[1]),.dout(n1602),.clk(gclk));
	jxor g1539(.dina(w_n1602_0[1]),.dinb(w_n1594_0[1]),.dout(n1603),.clk(gclk));
	jxor g1540(.dina(w_n1603_0[1]),.dinb(w_n1591_0[1]),.dout(n1604),.clk(gclk));
	jxor g1541(.dina(w_n1604_0[1]),.dinb(w_n1589_0[1]),.dout(n1605),.clk(gclk));
	jxor g1542(.dina(w_n1605_0[1]),.dinb(w_n1586_0[1]),.dout(n1606),.clk(gclk));
	jxor g1543(.dina(w_n1606_0[1]),.dinb(w_n1584_0[1]),.dout(n1607),.clk(gclk));
	jxor g1544(.dina(w_n1607_0[1]),.dinb(w_n1581_0[1]),.dout(n1608),.clk(gclk));
	jxor g1545(.dina(w_n1608_0[1]),.dinb(w_n1579_0[1]),.dout(n1609),.clk(gclk));
	jxor g1546(.dina(w_n1609_0[1]),.dinb(w_n1576_0[1]),.dout(n1610),.clk(gclk));
	jxor g1547(.dina(w_n1610_0[1]),.dinb(w_n1574_0[1]),.dout(n1611),.clk(gclk));
	jxor g1548(.dina(w_n1611_0[1]),.dinb(w_n1571_0[1]),.dout(n1612),.clk(gclk));
	jxor g1549(.dina(w_n1612_0[1]),.dinb(w_n1569_0[1]),.dout(n1613),.clk(gclk));
	jnot g1550(.din(n1613),.dout(n1614),.clk(gclk));
	jxor g1551(.dina(w_n1614_0[1]),.dinb(w_n1566_0[1]),.dout(n1615),.clk(gclk));
	jnot g1552(.din(n1615),.dout(n1616),.clk(gclk));
	jxor g1553(.dina(w_n1616_0[1]),.dinb(w_n1565_0[1]),.dout(n1617),.clk(gclk));
	jxor g1554(.dina(w_n1617_0[1]),.dinb(w_n1560_0[1]),.dout(w_dff_A_U4vuyFKf9_2),.clk(gclk));
	jor g1555(.dina(w_n1616_0[0]),.dinb(w_n1565_0[0]),.dout(n1619),.clk(gclk));
	jnot g1556(.din(w_n1617_0[0]),.dout(n1620),.clk(gclk));
	jor g1557(.dina(w_dff_B_JCTp6ct86_0),.dinb(w_n1560_0[0]),.dout(n1621),.clk(gclk));
	jand g1558(.dina(n1621),.dinb(w_dff_B_9hYt5XTP8_1),.dout(n1622),.clk(gclk));
	jnot g1559(.din(w_n1569_0[0]),.dout(n1623),.clk(gclk));
	jnot g1560(.din(w_n1612_0[0]),.dout(n1624),.clk(gclk));
	jor g1561(.dina(n1624),.dinb(n1623),.dout(n1625),.clk(gclk));
	jor g1562(.dina(w_n1614_0[0]),.dinb(w_n1566_0[0]),.dout(n1626),.clk(gclk));
	jand g1563(.dina(n1626),.dinb(w_dff_B_sOht3dtF1_1),.dout(n1627),.clk(gclk));
	jand g1564(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1628),.clk(gclk));
	jand g1565(.dina(w_n1610_0[0]),.dinb(w_n1574_0[0]),.dout(n1629),.clk(gclk));
	jand g1566(.dina(w_n1611_0[0]),.dinb(w_n1571_0[0]),.dout(n1630),.clk(gclk));
	jor g1567(.dina(n1630),.dinb(w_dff_B_5Zokezc54_1),.dout(n1631),.clk(gclk));
	jand g1568(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1632),.clk(gclk));
	jnot g1569(.din(n1632),.dout(n1633),.clk(gclk));
	jand g1570(.dina(w_n1608_0[0]),.dinb(w_n1579_0[0]),.dout(n1634),.clk(gclk));
	jand g1571(.dina(w_n1609_0[0]),.dinb(w_n1576_0[0]),.dout(n1635),.clk(gclk));
	jor g1572(.dina(n1635),.dinb(w_dff_B_UDKKrrrV9_1),.dout(n1636),.clk(gclk));
	jand g1573(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jand g1575(.dina(w_n1606_0[0]),.dinb(w_n1584_0[0]),.dout(n1639),.clk(gclk));
	jand g1576(.dina(w_n1607_0[0]),.dinb(w_n1581_0[0]),.dout(n1640),.clk(gclk));
	jor g1577(.dina(n1640),.dinb(w_dff_B_PuxHg3Gn7_1),.dout(n1641),.clk(gclk));
	jand g1578(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1642),.clk(gclk));
	jnot g1579(.din(n1642),.dout(n1643),.clk(gclk));
	jand g1580(.dina(w_n1604_0[0]),.dinb(w_n1589_0[0]),.dout(n1644),.clk(gclk));
	jand g1581(.dina(w_n1605_0[0]),.dinb(w_n1586_0[0]),.dout(n1645),.clk(gclk));
	jor g1582(.dina(n1645),.dinb(w_dff_B_xk3vPnoh0_1),.dout(n1646),.clk(gclk));
	jand g1583(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(n1647),.dout(n1648),.clk(gclk));
	jand g1585(.dina(w_n1602_0[0]),.dinb(w_n1594_0[0]),.dout(n1649),.clk(gclk));
	jand g1586(.dina(w_n1603_0[0]),.dinb(w_n1591_0[0]),.dout(n1650),.clk(gclk));
	jor g1587(.dina(n1650),.dinb(w_dff_B_WSfU75pS8_1),.dout(n1651),.clk(gclk));
	jand g1588(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1652),.clk(gclk));
	jand g1589(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1653),.clk(gclk));
	jor g1590(.dina(w_n1599_0[0]),.dinb(w_n1596_0[0]),.dout(n1654),.clk(gclk));
	jor g1591(.dina(w_n1601_0[0]),.dinb(w_n1595_0[0]),.dout(n1655),.clk(gclk));
	jand g1592(.dina(n1655),.dinb(w_dff_B_Hrnhfkl04_1),.dout(n1656),.clk(gclk));
	jxor g1593(.dina(w_n1656_0[1]),.dinb(w_n1653_0[1]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jxor g1595(.dina(w_n1658_0[1]),.dinb(w_n1652_0[1]),.dout(n1659),.clk(gclk));
	jxor g1596(.dina(w_n1659_0[1]),.dinb(w_n1651_0[1]),.dout(n1660),.clk(gclk));
	jxor g1597(.dina(w_n1660_0[1]),.dinb(w_n1648_0[1]),.dout(n1661),.clk(gclk));
	jxor g1598(.dina(w_n1661_0[1]),.dinb(w_n1646_0[1]),.dout(n1662),.clk(gclk));
	jxor g1599(.dina(w_n1662_0[1]),.dinb(w_n1643_0[1]),.dout(n1663),.clk(gclk));
	jxor g1600(.dina(w_n1663_0[1]),.dinb(w_n1641_0[1]),.dout(n1664),.clk(gclk));
	jxor g1601(.dina(w_n1664_0[1]),.dinb(w_n1638_0[1]),.dout(n1665),.clk(gclk));
	jxor g1602(.dina(w_n1665_0[1]),.dinb(w_n1636_0[1]),.dout(n1666),.clk(gclk));
	jxor g1603(.dina(w_n1666_0[1]),.dinb(w_n1633_0[1]),.dout(n1667),.clk(gclk));
	jxor g1604(.dina(w_n1667_0[1]),.dinb(w_n1631_0[1]),.dout(n1668),.clk(gclk));
	jnot g1605(.din(n1668),.dout(n1669),.clk(gclk));
	jxor g1606(.dina(w_n1669_0[1]),.dinb(w_n1628_0[1]),.dout(n1670),.clk(gclk));
	jnot g1607(.din(n1670),.dout(n1671),.clk(gclk));
	jxor g1608(.dina(w_n1671_0[1]),.dinb(w_n1627_0[1]),.dout(n1672),.clk(gclk));
	jxor g1609(.dina(w_n1672_0[1]),.dinb(w_n1622_0[1]),.dout(w_dff_A_nROzBrc79_2),.clk(gclk));
	jor g1610(.dina(w_n1671_0[0]),.dinb(w_n1627_0[0]),.dout(n1674),.clk(gclk));
	jnot g1611(.din(w_n1672_0[0]),.dout(n1675),.clk(gclk));
	jor g1612(.dina(w_dff_B_a4Snyv5j7_0),.dinb(w_n1622_0[0]),.dout(n1676),.clk(gclk));
	jand g1613(.dina(n1676),.dinb(w_dff_B_Hczv6KUZ7_1),.dout(n1677),.clk(gclk));
	jnot g1614(.din(w_n1631_0[0]),.dout(n1678),.clk(gclk));
	jnot g1615(.din(w_n1667_0[0]),.dout(n1679),.clk(gclk));
	jor g1616(.dina(n1679),.dinb(w_dff_B_BpAGy5bV6_1),.dout(n1680),.clk(gclk));
	jor g1617(.dina(w_n1669_0[0]),.dinb(w_n1628_0[0]),.dout(n1681),.clk(gclk));
	jand g1618(.dina(n1681),.dinb(w_dff_B_YpIpUHEK4_1),.dout(n1682),.clk(gclk));
	jand g1619(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1683),.clk(gclk));
	jnot g1620(.din(n1683),.dout(n1684),.clk(gclk));
	jand g1621(.dina(w_n1665_0[0]),.dinb(w_n1636_0[0]),.dout(n1685),.clk(gclk));
	jand g1622(.dina(w_n1666_0[0]),.dinb(w_n1633_0[0]),.dout(n1686),.clk(gclk));
	jor g1623(.dina(n1686),.dinb(w_dff_B_rH54O8kr0_1),.dout(n1687),.clk(gclk));
	jand g1624(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1688),.clk(gclk));
	jnot g1625(.din(n1688),.dout(n1689),.clk(gclk));
	jand g1626(.dina(w_n1663_0[0]),.dinb(w_n1641_0[0]),.dout(n1690),.clk(gclk));
	jand g1627(.dina(w_n1664_0[0]),.dinb(w_n1638_0[0]),.dout(n1691),.clk(gclk));
	jor g1628(.dina(n1691),.dinb(w_dff_B_JljeUlJQ0_1),.dout(n1692),.clk(gclk));
	jand g1629(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1693),.clk(gclk));
	jnot g1630(.din(n1693),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1661_0[0]),.dinb(w_n1646_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1662_0[0]),.dinb(w_n1643_0[0]),.dout(n1696),.clk(gclk));
	jor g1633(.dina(n1696),.dinb(w_dff_B_lFIuXwu42_1),.dout(n1697),.clk(gclk));
	jand g1634(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1659_0[0]),.dinb(w_n1651_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1660_0[0]),.dinb(w_n1648_0[0]),.dout(n1701),.clk(gclk));
	jor g1638(.dina(n1701),.dinb(w_dff_B_FYAmhI927_1),.dout(n1702),.clk(gclk));
	jand g1639(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1703),.clk(gclk));
	jand g1640(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1704),.clk(gclk));
	jor g1641(.dina(w_n1656_0[0]),.dinb(w_n1653_0[0]),.dout(n1705),.clk(gclk));
	jor g1642(.dina(w_n1658_0[0]),.dinb(w_n1652_0[0]),.dout(n1706),.clk(gclk));
	jand g1643(.dina(n1706),.dinb(w_dff_B_6xgTCNBr0_1),.dout(n1707),.clk(gclk));
	jxor g1644(.dina(w_n1707_0[1]),.dinb(w_n1704_0[1]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jxor g1646(.dina(w_n1709_0[1]),.dinb(w_n1703_0[1]),.dout(n1710),.clk(gclk));
	jxor g1647(.dina(w_n1710_0[1]),.dinb(w_n1702_0[1]),.dout(n1711),.clk(gclk));
	jxor g1648(.dina(w_n1711_0[1]),.dinb(w_n1699_0[1]),.dout(n1712),.clk(gclk));
	jxor g1649(.dina(w_n1712_0[1]),.dinb(w_n1697_0[1]),.dout(n1713),.clk(gclk));
	jxor g1650(.dina(w_n1713_0[1]),.dinb(w_n1694_0[1]),.dout(n1714),.clk(gclk));
	jxor g1651(.dina(w_n1714_0[1]),.dinb(w_n1692_0[1]),.dout(n1715),.clk(gclk));
	jxor g1652(.dina(w_n1715_0[1]),.dinb(w_n1689_0[1]),.dout(n1716),.clk(gclk));
	jxor g1653(.dina(w_n1716_0[1]),.dinb(w_n1687_0[1]),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1684_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1682_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1677_0[1]),.dout(w_dff_A_Hct20z8J2_2),.clk(gclk));
	jor g1658(.dina(w_n1719_0[0]),.dinb(w_n1682_0[0]),.dout(n1722),.clk(gclk));
	jnot g1659(.din(w_n1720_0[0]),.dout(n1723),.clk(gclk));
	jor g1660(.dina(w_dff_B_apjOOWYS0_0),.dinb(w_n1677_0[0]),.dout(n1724),.clk(gclk));
	jand g1661(.dina(n1724),.dinb(w_dff_B_Wq2Kv3s35_1),.dout(n1725),.clk(gclk));
	jand g1662(.dina(w_n1716_0[0]),.dinb(w_n1687_0[0]),.dout(n1726),.clk(gclk));
	jand g1663(.dina(w_n1717_0[0]),.dinb(w_n1684_0[0]),.dout(n1727),.clk(gclk));
	jor g1664(.dina(n1727),.dinb(w_dff_B_apJ5POHG4_1),.dout(n1728),.clk(gclk));
	jand g1665(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(n1729),.dout(n1730),.clk(gclk));
	jand g1667(.dina(w_n1714_0[0]),.dinb(w_n1692_0[0]),.dout(n1731),.clk(gclk));
	jand g1668(.dina(w_n1715_0[0]),.dinb(w_n1689_0[0]),.dout(n1732),.clk(gclk));
	jor g1669(.dina(n1732),.dinb(w_dff_B_tYvUEpmN3_1),.dout(n1733),.clk(gclk));
	jand g1670(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1734),.clk(gclk));
	jnot g1671(.din(n1734),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1712_0[0]),.dinb(w_n1697_0[0]),.dout(n1736),.clk(gclk));
	jand g1673(.dina(w_n1713_0[0]),.dinb(w_n1694_0[0]),.dout(n1737),.clk(gclk));
	jor g1674(.dina(n1737),.dinb(w_dff_B_th8nxmQb1_1),.dout(n1738),.clk(gclk));
	jand g1675(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1739),.clk(gclk));
	jnot g1676(.din(n1739),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1710_0[0]),.dinb(w_n1702_0[0]),.dout(n1741),.clk(gclk));
	jand g1678(.dina(w_n1711_0[0]),.dinb(w_n1699_0[0]),.dout(n1742),.clk(gclk));
	jor g1679(.dina(n1742),.dinb(w_dff_B_4Bt6y4zt0_1),.dout(n1743),.clk(gclk));
	jand g1680(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1745),.clk(gclk));
	jor g1682(.dina(w_n1707_0[0]),.dinb(w_n1704_0[0]),.dout(n1746),.clk(gclk));
	jor g1683(.dina(w_n1709_0[0]),.dinb(w_n1703_0[0]),.dout(n1747),.clk(gclk));
	jand g1684(.dina(n1747),.dinb(w_dff_B_UoYNGMjq0_1),.dout(n1748),.clk(gclk));
	jxor g1685(.dina(w_n1748_0[1]),.dinb(w_n1745_0[1]),.dout(n1749),.clk(gclk));
	jnot g1686(.din(n1749),.dout(n1750),.clk(gclk));
	jxor g1687(.dina(w_n1750_0[1]),.dinb(w_n1744_0[1]),.dout(n1751),.clk(gclk));
	jxor g1688(.dina(w_n1751_0[1]),.dinb(w_n1743_0[1]),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1740_0[1]),.dout(n1753),.clk(gclk));
	jxor g1690(.dina(w_n1753_0[1]),.dinb(w_n1738_0[1]),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1735_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1733_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1730_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1728_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1725_0[1]),.dout(w_dff_A_48KSIqDl5_2),.clk(gclk));
	jnot g1696(.din(w_n1728_0[0]),.dout(n1760),.clk(gclk));
	jnot g1697(.din(w_n1757_0[0]),.dout(n1761),.clk(gclk));
	jor g1698(.dina(n1761),.dinb(w_dff_B_ujHNKIta2_1),.dout(n1762),.clk(gclk));
	jnot g1699(.din(w_n1758_0[0]),.dout(n1763),.clk(gclk));
	jor g1700(.dina(w_dff_B_3nD9Myey6_0),.dinb(w_n1725_0[0]),.dout(n1764),.clk(gclk));
	jand g1701(.dina(n1764),.dinb(w_dff_B_yegT27uo2_1),.dout(n1765),.clk(gclk));
	jand g1702(.dina(w_n1755_0[0]),.dinb(w_n1733_0[0]),.dout(n1766),.clk(gclk));
	jand g1703(.dina(w_n1756_0[0]),.dinb(w_n1730_0[0]),.dout(n1767),.clk(gclk));
	jor g1704(.dina(n1767),.dinb(w_dff_B_K1E8wuCf6_1),.dout(n1768),.clk(gclk));
	jand g1705(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1769),.clk(gclk));
	jnot g1706(.din(n1769),.dout(n1770),.clk(gclk));
	jand g1707(.dina(w_n1753_0[0]),.dinb(w_n1738_0[0]),.dout(n1771),.clk(gclk));
	jand g1708(.dina(w_n1754_0[0]),.dinb(w_n1735_0[0]),.dout(n1772),.clk(gclk));
	jor g1709(.dina(n1772),.dinb(w_dff_B_DfFTOkR05_1),.dout(n1773),.clk(gclk));
	jand g1710(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1774),.clk(gclk));
	jnot g1711(.din(n1774),.dout(n1775),.clk(gclk));
	jand g1712(.dina(w_n1751_0[0]),.dinb(w_n1743_0[0]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_n1752_0[0]),.dinb(w_n1740_0[0]),.dout(n1777),.clk(gclk));
	jor g1714(.dina(n1777),.dinb(w_dff_B_L2SDGRk72_1),.dout(n1778),.clk(gclk));
	jand g1715(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1779),.clk(gclk));
	jand g1716(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1780),.clk(gclk));
	jor g1717(.dina(w_n1748_0[0]),.dinb(w_n1745_0[0]),.dout(n1781),.clk(gclk));
	jor g1718(.dina(w_n1750_0[0]),.dinb(w_n1744_0[0]),.dout(n1782),.clk(gclk));
	jand g1719(.dina(n1782),.dinb(w_dff_B_Zw6pdW2B7_1),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1780_0[1]),.dout(n1784),.clk(gclk));
	jnot g1721(.din(n1784),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1779_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1778_0[1]),.dout(n1787),.clk(gclk));
	jxor g1724(.dina(w_n1787_0[1]),.dinb(w_n1775_0[1]),.dout(n1788),.clk(gclk));
	jxor g1725(.dina(w_n1788_0[1]),.dinb(w_n1773_0[1]),.dout(n1789),.clk(gclk));
	jxor g1726(.dina(w_n1789_0[1]),.dinb(w_n1770_0[1]),.dout(n1790),.clk(gclk));
	jxor g1727(.dina(w_n1790_0[1]),.dinb(w_n1768_0[1]),.dout(n1791),.clk(gclk));
	jxor g1728(.dina(w_n1791_0[1]),.dinb(w_n1765_0[1]),.dout(w_dff_A_uIbrthHL5_2),.clk(gclk));
	jnot g1729(.din(w_n1768_0[0]),.dout(n1793),.clk(gclk));
	jnot g1730(.din(w_n1790_0[0]),.dout(n1794),.clk(gclk));
	jor g1731(.dina(n1794),.dinb(w_dff_B_zTqoFgxU7_1),.dout(n1795),.clk(gclk));
	jnot g1732(.din(w_n1791_0[0]),.dout(n1796),.clk(gclk));
	jor g1733(.dina(w_dff_B_tvgH6RWW3_0),.dinb(w_n1765_0[0]),.dout(n1797),.clk(gclk));
	jand g1734(.dina(n1797),.dinb(w_dff_B_fdbJkxX72_1),.dout(n1798),.clk(gclk));
	jand g1735(.dina(w_n1788_0[0]),.dinb(w_n1773_0[0]),.dout(n1799),.clk(gclk));
	jand g1736(.dina(w_n1789_0[0]),.dinb(w_n1770_0[0]),.dout(n1800),.clk(gclk));
	jor g1737(.dina(n1800),.dinb(w_dff_B_M3dpZsFI7_1),.dout(n1801),.clk(gclk));
	jand g1738(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jand g1740(.dina(w_n1786_0[0]),.dinb(w_n1778_0[0]),.dout(n1804),.clk(gclk));
	jand g1741(.dina(w_n1787_0[0]),.dinb(w_n1775_0[0]),.dout(n1805),.clk(gclk));
	jor g1742(.dina(n1805),.dinb(w_dff_B_F4FHKNsW0_1),.dout(n1806),.clk(gclk));
	jand g1743(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1807),.clk(gclk));
	jand g1744(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1808),.clk(gclk));
	jor g1745(.dina(w_n1783_0[0]),.dinb(w_n1780_0[0]),.dout(n1809),.clk(gclk));
	jor g1746(.dina(w_n1785_0[0]),.dinb(w_n1779_0[0]),.dout(n1810),.clk(gclk));
	jand g1747(.dina(n1810),.dinb(w_dff_B_4SA924Xj6_1),.dout(n1811),.clk(gclk));
	jxor g1748(.dina(w_n1811_0[1]),.dinb(w_n1808_0[1]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(n1812),.dout(n1813),.clk(gclk));
	jxor g1750(.dina(w_n1813_0[1]),.dinb(w_n1807_0[1]),.dout(n1814),.clk(gclk));
	jxor g1751(.dina(w_n1814_0[1]),.dinb(w_n1806_0[1]),.dout(n1815),.clk(gclk));
	jxor g1752(.dina(w_n1815_0[1]),.dinb(w_n1803_0[1]),.dout(n1816),.clk(gclk));
	jxor g1753(.dina(w_n1816_0[1]),.dinb(w_n1801_0[1]),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1817_0[1]),.dinb(w_n1798_0[1]),.dout(w_dff_A_UUSXDR6i6_2),.clk(gclk));
	jnot g1755(.din(w_n1801_0[0]),.dout(n1819),.clk(gclk));
	jnot g1756(.din(w_n1816_0[0]),.dout(n1820),.clk(gclk));
	jor g1757(.dina(n1820),.dinb(w_dff_B_YhTOozlg0_1),.dout(n1821),.clk(gclk));
	jnot g1758(.din(w_n1817_0[0]),.dout(n1822),.clk(gclk));
	jor g1759(.dina(w_dff_B_EHataNLT3_0),.dinb(w_n1798_0[0]),.dout(n1823),.clk(gclk));
	jand g1760(.dina(n1823),.dinb(w_dff_B_NQTZLS0q4_1),.dout(n1824),.clk(gclk));
	jand g1761(.dina(w_n1814_0[0]),.dinb(w_n1806_0[0]),.dout(n1825),.clk(gclk));
	jand g1762(.dina(w_n1815_0[0]),.dinb(w_n1803_0[0]),.dout(n1826),.clk(gclk));
	jor g1763(.dina(n1826),.dinb(w_dff_B_tNkfSlSJ7_1),.dout(n1827),.clk(gclk));
	jand g1764(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1828),.clk(gclk));
	jand g1765(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1829),.clk(gclk));
	jor g1766(.dina(w_n1811_0[0]),.dinb(w_n1808_0[0]),.dout(n1830),.clk(gclk));
	jor g1767(.dina(w_n1813_0[0]),.dinb(w_n1807_0[0]),.dout(n1831),.clk(gclk));
	jand g1768(.dina(n1831),.dinb(w_dff_B_SykyZ5wE9_1),.dout(n1832),.clk(gclk));
	jxor g1769(.dina(w_n1832_0[1]),.dinb(w_n1829_0[1]),.dout(n1833),.clk(gclk));
	jnot g1770(.din(n1833),.dout(n1834),.clk(gclk));
	jxor g1771(.dina(w_n1834_0[1]),.dinb(w_n1828_0[1]),.dout(n1835),.clk(gclk));
	jxor g1772(.dina(w_n1835_0[1]),.dinb(w_n1827_0[1]),.dout(n1836),.clk(gclk));
	jxor g1773(.dina(w_n1836_0[1]),.dinb(w_n1824_0[1]),.dout(w_dff_A_zwUMdALK2_2),.clk(gclk));
	jand g1774(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1838),.clk(gclk));
	jor g1775(.dina(w_n1832_0[0]),.dinb(w_n1829_0[0]),.dout(n1839),.clk(gclk));
	jor g1776(.dina(w_n1834_0[0]),.dinb(w_n1828_0[0]),.dout(n1840),.clk(gclk));
	jand g1777(.dina(n1840),.dinb(w_dff_B_WOnb8SOF2_1),.dout(n1841),.clk(gclk));
	jor g1778(.dina(w_n1841_0[1]),.dinb(w_n1838_0[1]),.dout(n1842),.clk(gclk));
	jnot g1779(.din(w_n1827_0[0]),.dout(n1843),.clk(gclk));
	jnot g1780(.din(w_n1835_0[0]),.dout(n1844),.clk(gclk));
	jor g1781(.dina(n1844),.dinb(w_dff_B_jCAK1uKJ6_1),.dout(n1845),.clk(gclk));
	jnot g1782(.din(w_n1836_0[0]),.dout(n1846),.clk(gclk));
	jor g1783(.dina(w_dff_B_qFQVdwG56_0),.dinb(w_n1824_0[0]),.dout(n1847),.clk(gclk));
	jand g1784(.dina(n1847),.dinb(w_dff_B_9BjyQurF6_1),.dout(n1848),.clk(gclk));
	jxor g1785(.dina(w_n1841_0[0]),.dinb(w_n1838_0[0]),.dout(n1849),.clk(gclk));
	jnot g1786(.din(w_n1849_0[1]),.dout(n1850),.clk(gclk));
	jor g1787(.dina(w_dff_B_3PRkUcnj7_0),.dinb(w_n1848_0[1]),.dout(n1851),.clk(gclk));
	jand g1788(.dina(n1851),.dinb(w_dff_B_CRQgdMGd2_1),.dout(G6287gat),.clk(gclk));
	jxor g1789(.dina(w_n1849_0[0]),.dinb(w_n1848_0[0]),.dout(w_dff_A_KQCoHiXA8_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl3 jspl3_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.doutc(w_G18gat_7[2]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl3 jspl3_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.doutc(w_G273gat_7[2]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_dff_A_x4eBRqMp2_1),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl3 jspl3_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.doutc(w_G307gat_7[2]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(w_dff_A_qLYUvskc7_1),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n69_0(.douta(w_dff_A_qNtSau7H0_0),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_dff_A_jVSOrltG9_0),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n72_0(.douta(w_dff_A_yQlDCY0r9_0),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.din(n81));
	jspl3 jspl3_w_n82_0(.douta(w_n82_0[0]),.doutb(w_dff_A_2wtDOQkA6_1),.doutc(w_dff_A_isb7tLK02_2),.din(n82));
	jspl jspl_w_n82_1(.douta(w_n82_1[0]),.doutb(w_dff_A_wzFeeiny6_1),.din(w_n82_0[0]));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n85_0(.douta(w_dff_A_zA7efneb1_0),.doutb(w_n85_0[1]),.din(n85));
	jspl jspl_w_n87_0(.douta(w_n87_0[0]),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_dff_A_3bc51pMd5_0),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n94_0(.douta(w_dff_A_o96JgnLg3_0),.doutb(w_n94_0[1]),.din(n94));
	jspl jspl_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n100_0(.douta(w_n100_0[0]),.doutb(w_dff_A_IqkzQ5Xs0_1),.doutc(w_dff_A_Z0PxXlJi4_2),.din(n100));
	jspl jspl_w_n100_1(.douta(w_dff_A_wRGR6vxt7_0),.doutb(w_n100_1[1]),.din(w_n100_0[0]));
	jspl3 jspl3_w_n101_0(.douta(w_dff_A_jIE5RpNV8_0),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_dff_A_ULikrVqh5_0),.doutb(w_n103_0[1]),.din(n103));
	jspl jspl_w_n104_0(.douta(w_dff_A_IGVxKSBU0_0),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_dff_A_CTRaqL9B3_1),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n110_0(.douta(w_dff_A_1tP4Ojsj6_0),.doutb(w_n110_0[1]),.din(n110));
	jspl jspl_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.din(n115));
	jspl jspl_w_n116_0(.douta(w_dff_A_t8goGsCr9_0),.doutb(w_n116_0[1]),.din(n116));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(w_dff_B_LmbkEhOm2_2));
	jspl jspl_w_n129_0(.douta(w_n129_0[0]),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_dff_A_kaDeBZSS5_1),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_dff_A_dBh5L1BT2_0),.doutb(w_dff_A_nybzF4DU4_1),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.doutc(w_n133_0[2]),.din(n133));
	jspl jspl_w_n138_0(.douta(w_n138_0[0]),.doutb(w_n138_0[1]),.din(n138));
	jspl jspl_w_n139_0(.douta(w_dff_A_1LCq0UX68_0),.doutb(w_n139_0[1]),.din(n139));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_dff_A_16lnEayP7_1),.din(n142));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl jspl_w_n145_0(.douta(w_dff_A_zXoueFPQ6_0),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n150_0(.douta(w_n150_0[0]),.doutb(w_n150_0[1]),.din(n150));
	jspl jspl_w_n151_0(.douta(w_dff_A_Npyp55tc1_0),.doutb(w_n151_0[1]),.din(n151));
	jspl3 jspl3_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.doutc(w_n156_0[2]),.din(n156));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(w_dff_B_6WHuhTtx4_2));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(w_dff_B_kzWq9imN9_2));
	jspl jspl_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.din(n166));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n169_0(.douta(w_dff_A_a8R000an1_0),.doutb(w_dff_A_gZCz23As0_1),.doutc(w_n169_0[2]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(w_dff_B_CZmZ4Z1s3_2));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl jspl_w_n177_0(.douta(w_dff_A_JG8iwnZG5_0),.doutb(w_n177_0[1]),.din(n177));
	jspl jspl_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.din(n178));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_dff_A_t5eeBDnN5_1),.din(n180));
	jspl jspl_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.din(n181));
	jspl jspl_w_n183_0(.douta(w_dff_A_VZPaFjUV4_0),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_dff_A_ashIQI344_0),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.doutc(w_n194_0[2]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.din(w_dff_B_SL8ZdoEa6_2));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(w_dff_B_mfADympr8_2));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(w_dff_B_eL30RuV68_2));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.din(n209));
	jspl3 jspl3_w_n210_0(.douta(w_n210_0[0]),.doutb(w_dff_A_ihGef0np8_1),.doutc(w_dff_A_ME7jCby71_2),.din(n210));
	jspl jspl_w_n210_1(.douta(w_dff_A_ab6agvHO7_0),.doutb(w_n210_1[1]),.din(w_n210_0[0]));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl jspl_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.din(n215));
	jspl jspl_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.din(w_dff_B_my4An37E2_2));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(w_dff_B_BwpPDbDd4_2));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_dff_A_DPpMOZQn6_0),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.din(n221));
	jspl jspl_w_n223_0(.douta(w_n223_0[0]),.doutb(w_dff_A_jlM84O8q0_1),.din(n223));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n226_0(.douta(w_dff_A_r7OMeDpp7_0),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.din(n231));
	jspl jspl_w_n232_0(.douta(w_dff_A_jgurZwdt9_0),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n237_0(.douta(w_n237_0[0]),.doutb(w_n237_0[1]),.doutc(w_n237_0[2]),.din(n237));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(w_dff_B_z2IB3KoP5_2));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.din(w_dff_B_oKHH0kyI4_2));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_60eohaZi9_2));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(w_dff_B_NxmFnLMh2_2));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_n257_0[1]),.din(n257));
	jspl3 jspl3_w_n258_0(.douta(w_dff_A_aBDBlh6d9_0),.doutb(w_dff_A_eBdNRukX7_1),.doutc(w_n258_0[2]),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(w_dff_B_2ccDlXr84_2));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(w_dff_B_1ynuhIjH3_2));
	jspl jspl_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.din(n268));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.din(w_dff_B_lNc23o2r7_2));
	jspl jspl_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.din(n270));
	jspl jspl_w_n271_0(.douta(w_dff_A_6MqYMjVg1_0),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_uk6LQE8m1_1),.din(n274));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl jspl_w_n277_0(.douta(w_dff_A_WJYgSSeq1_0),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n283_0(.douta(w_dff_A_OPdTFdsX8_0),.doutb(w_n283_0[1]),.din(n283));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(w_dff_B_KvgfoixZ0_2));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(w_dff_B_OiP437gK3_2));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_n300_0[1]),.din(w_dff_B_gwbk1L7D7_2));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(w_dff_B_qiqaGBdF2_2));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(w_dff_B_CpkB4cPl0_2));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n314_0(.douta(w_dff_A_BCYGFEtJ4_0),.doutb(w_dff_A_TShp7RaZ3_1),.doutc(w_n314_0[2]),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.din(n317));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.din(w_dff_B_GQJav8ev3_2));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(w_dff_B_in7sRfZw5_2));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(w_dff_B_XBXvx0H27_2));
	jspl jspl_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.din(n326));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(w_dff_B_otGOyUp50_2));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n329_0(.douta(w_dff_A_iWTcsfKo0_0),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(n330));
	jspl jspl_w_n332_0(.douta(w_n332_0[0]),.doutb(w_dff_A_VidqzFNW6_1),.din(n332));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_dff_A_PEKduRXH7_0),.doutb(w_n335_0[1]),.din(n335));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl jspl_w_n341_0(.douta(w_dff_A_wwsr9i9c7_0),.doutb(w_n341_0[1]),.din(n341));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(w_dff_B_InpKIDaf8_2));
	jspl jspl_w_n351_0(.douta(w_n351_0[0]),.doutb(w_n351_0[1]),.din(n351));
	jspl jspl_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.din(w_dff_B_N8WbGEM79_2));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(n356));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(w_dff_B_d7k18fMk7_2));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(w_dff_B_VkUFP3RP6_2));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(n366));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(w_dff_B_9r95EjvW0_2));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_Fn4KLys41_1),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl3 jspl3_w_n376_0(.douta(w_dff_A_vbg071tF9_0),.doutb(w_dff_A_zMPDIusV4_1),.doutc(w_n376_0[2]),.din(n376));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.din(n377));
	jspl jspl_w_n380_0(.douta(w_dff_A_FNgLIZwm6_0),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.din(n382));
	jspl jspl_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.din(n383));
	jspl jspl_w_n384_0(.douta(w_n384_0[0]),.doutb(w_n384_0[1]),.din(n384));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(w_dff_B_io9CbdDf0_2));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl jspl_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.din(w_dff_B_OSIDnEiA1_2));
	jspl jspl_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.din(n388));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.din(w_dff_B_6D1veawk7_2));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(n390));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(w_dff_B_Cv00onWb5_2));
	jspl jspl_w_n392_0(.douta(w_n392_0[0]),.doutb(w_n392_0[1]),.din(n392));
	jspl jspl_w_n393_0(.douta(w_dff_A_kU40C3S38_0),.doutb(w_n393_0[1]),.din(n393));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_dff_A_3CJq4Na68_1),.din(n396));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n399_0(.douta(w_dff_A_pnmCap4I7_0),.doutb(w_n399_0[1]),.din(n399));
	jspl jspl_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_dff_A_QtvxpQdK0_0),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_n410_0[2]),.din(n410));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(w_dff_B_vJ5JRxYC2_2));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl jspl_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.din(w_dff_B_YprPyH070_2));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.din(n420));
	jspl jspl_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.din(w_dff_B_bCkENo171_2));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(w_dff_B_ip1OYZXP2_2));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(w_dff_B_wz3dzYdM9_2));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(w_dff_B_j6F4Nlxt6_2));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(w_dff_B_mJYNJxgE9_2));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_dff_A_tRz3lwnQ9_1),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n446_0(.douta(w_dff_A_TrtfMKBO0_0),.doutb(w_dff_A_hDjMxZIc3_1),.doutc(w_n446_0[2]),.din(n446));
	jspl jspl_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.din(n447));
	jspl jspl_w_n450_0(.douta(w_dff_A_1dQUkF5l2_0),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.din(w_dff_B_pOhTzdCH3_2));
	jspl jspl_w_n454_0(.douta(w_n454_0[0]),.doutb(w_n454_0[1]),.din(n454));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.din(n455));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl jspl_w_n458_0(.douta(w_n458_0[0]),.doutb(w_n458_0[1]),.din(n458));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(w_dff_B_joj2jMnZ3_2));
	jspl jspl_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.din(n460));
	jspl jspl_w_n461_0(.douta(w_n461_0[0]),.doutb(w_n461_0[1]),.din(w_dff_B_g1o7SUW86_2));
	jspl jspl_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.din(n462));
	jspl jspl_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.din(w_dff_B_Moc7km7x7_2));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(n464));
	jspl jspl_w_n465_0(.douta(w_dff_A_pvQlB12I5_0),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(n466));
	jspl jspl_w_n468_0(.douta(w_n468_0[0]),.doutb(w_dff_A_JKTgIqrw1_1),.din(n468));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(n469));
	jspl jspl_w_n471_0(.douta(w_dff_A_3ewd5nH07_0),.doutb(w_n471_0[1]),.din(n471));
	jspl jspl_w_n476_0(.douta(w_n476_0[0]),.doutb(w_n476_0[1]),.din(n476));
	jspl jspl_w_n477_0(.douta(w_dff_A_CoUUaYe63_0),.doutb(w_n477_0[1]),.din(n477));
	jspl3 jspl3_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.doutc(w_n482_0[2]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(w_dff_B_ukBH0eR21_2));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(w_dff_B_vtYozoDN3_2));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(w_dff_B_P90XYJTQ4_2));
	jspl jspl_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.din(n497));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(w_dff_B_2oiaiKTi4_2));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(w_dff_B_UOTUdhWY3_2));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_c848xsSQ9_2));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(w_dff_B_ldFlnqha2_2));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_dff_A_rAkL1biL0_1),.din(n519));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_dff_A_okRv4hTg5_0),.doutb(w_dff_A_w7exM3Ua5_1),.doutc(w_n523_0[2]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n527_0(.douta(w_dff_A_ORLsOMXy6_0),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_n529_0[0]),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(w_dff_B_AaPrnNlc1_2));
	jspl jspl_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.din(n531));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(w_dff_B_upS3G5Yz1_2));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.din(n535));
	jspl jspl_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.din(n536));
	jspl jspl_w_n537_0(.douta(w_n537_0[0]),.doutb(w_n537_0[1]),.din(n537));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(w_dff_B_dPQiGyWm2_2));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(w_dff_B_Jjsyq7Hc5_2));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(w_dff_B_PlMEJB0o9_2));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n544_0(.douta(w_dff_A_OzxLbf6k9_0),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_dff_A_iE7a1jkd8_1),.din(n547));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_dff_A_B7YqcfYP3_0),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n556_0(.douta(w_dff_A_V61aGOcA3_0),.doutb(w_n556_0[1]),.din(n556));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(w_dff_B_OO7HPbty9_2));
	jspl jspl_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.din(n566));
	jspl jspl_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.din(w_dff_B_DAT7my1X3_2));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.din(n571));
	jspl jspl_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.din(w_dff_B_X1JJlNGf9_2));
	jspl jspl_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.din(n576));
	jspl jspl_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.din(w_dff_B_UEsYEI8b8_2));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl jspl_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.din(w_dff_B_fFbzYEDd7_2));
	jspl jspl_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(w_dff_B_KZqUSP9O5_2));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(w_dff_B_NZTP6NYu9_2));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(n596));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(w_dff_B_9ozcuxUk2_2));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_dff_A_uAiNKDt00_1),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(n606));
	jspl3 jspl3_w_n607_0(.douta(w_dff_A_NXNylrvi2_0),.doutb(w_dff_A_M9IiwrW08_1),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n611_0(.douta(w_dff_A_p1ExIVA06_0),.doutb(w_n611_0[1]),.din(n611));
	jspl jspl_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.din(n613));
	jspl jspl_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.din(w_dff_B_pV3RM8kO6_2));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(w_dff_B_fZAO0HLr4_2));
	jspl jspl_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.din(n617));
	jspl jspl_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.din(w_dff_B_Y2egNx893_2));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.din(n620));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.din(n621));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(w_dff_B_TuOrFy6A8_2));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.din(n625));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(w_dff_B_YdHV0KgQ8_2));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(w_dff_B_WD6Ur2R19_2));
	jspl jspl_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.din(n629));
	jspl jspl_w_n630_0(.douta(w_dff_A_8nZPzhWn0_0),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n633_0(.douta(w_n633_0[0]),.doutb(w_dff_A_VEujq0b56_1),.din(n633));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl jspl_w_n636_0(.douta(w_dff_A_iTXaZvbS8_0),.doutb(w_n636_0[1]),.din(n636));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_dff_A_ovFp6XYL3_0),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.doutc(w_n647_0[2]),.din(n647));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(w_dff_B_69glCq6x7_2));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(w_dff_B_YybAkBW14_2));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(w_dff_B_1yZeRs0z3_2));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(n662));
	jspl jspl_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.din(w_dff_B_jReiZpSs1_2));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(n667));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(w_dff_B_Ef4mkVVx3_2));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(w_dff_B_hsU6ID7L5_2));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.din(w_dff_B_k2iDG3JR1_2));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(w_dff_B_bFjrIidG9_2));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(w_dff_B_3vDR8Cz34_2));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_dff_A_pFIzj7hA7_1),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_dff_A_WbOULxLr1_0),.doutb(w_n695_0[1]),.doutc(w_n695_0[2]),.din(n695));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl3 jspl3_w_n698_0(.douta(w_dff_A_T2OwA3n83_0),.doutb(w_dff_A_45MFTm1j1_1),.doutc(w_n698_0[2]),.din(n698));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n702_0(.douta(w_dff_A_PuqeexTg5_0),.doutb(w_n702_0[1]),.din(n702));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(w_dff_B_zqjynpTp0_2));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.din(w_dff_B_4IdKWKoN1_2));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.din(n708));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(w_dff_B_rnu65OlP0_2));
	jspl jspl_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(w_dff_B_wuzspgXl2_2));
	jspl jspl_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl jspl_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.din(n714));
	jspl jspl_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.din(n715));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(w_dff_B_wQdkmXAX3_2));
	jspl jspl_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.din(n718));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(w_dff_B_5HHz45KX0_2));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(w_dff_B_G3QqpJfF0_2));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n723_0(.douta(w_dff_A_hp903XOU7_0),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(n724));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_dff_A_9NszZZ8G3_1),.din(n726));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_dff_A_rg9oEtRT9_0),.doutb(w_n729_0[1]),.din(n729));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(n734));
	jspl jspl_w_n735_0(.douta(w_dff_A_Bb9hNL731_0),.doutb(w_n735_0[1]),.din(n735));
	jspl3 jspl3_w_n740_0(.douta(w_n740_0[0]),.doutb(w_n740_0[1]),.doutc(w_n740_0[2]),.din(n740));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(w_dff_B_X2BvY5948_2));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(w_dff_B_98cUKTy00_2));
	jspl jspl_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(w_dff_B_s1oEiOdU9_2));
	jspl jspl_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.din(n755));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(w_dff_B_3UUv34cF6_2));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(w_dff_B_jXm3dBaj8_2));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(w_dff_B_Z8L1CnUT9_2));
	jspl jspl_w_n770_0(.douta(w_n770_0[0]),.doutb(w_n770_0[1]),.din(n770));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(w_dff_B_ikKPjnGQ6_2));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(w_dff_B_zmwDxNgR1_2));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(w_dff_B_AxSNxK3Y9_2));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_khvspGQO6_2));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_dff_A_kO1gTAnV0_1),.din(n792));
	jspl jspl_w_n793_0(.douta(w_dff_A_t44wiNYu7_0),.doutb(w_n793_0[1]),.din(n793));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl jspl_w_n800_0(.douta(w_dff_A_CxS8Eef66_0),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(w_dff_B_z0LSDmXY5_2));
	jspl jspl_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.din(n804));
	jspl jspl_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.din(w_dff_B_RFXlgBXa0_2));
	jspl jspl_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.din(n806));
	jspl jspl_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.din(w_dff_B_ybKDPPf21_2));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.din(n808));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(w_dff_B_szXqKr1U5_2));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(w_dff_B_WSBkRGqV8_2));
	jspl jspl_w_n812_0(.douta(w_n812_0[0]),.doutb(w_n812_0[1]),.din(n812));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl jspl_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.din(n814));
	jspl jspl_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(w_dff_B_sJWUG6142_2));
	jspl jspl_w_n818_0(.douta(w_n818_0[0]),.doutb(w_n818_0[1]),.din(n818));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(w_dff_B_WcmNniVo7_2));
	jspl jspl_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.din(n820));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(w_dff_B_0o7XpGAz9_2));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(n822));
	jspl jspl_w_n823_0(.douta(w_dff_A_ykRVGLmZ7_0),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n826_0(.douta(w_n826_0[0]),.doutb(w_dff_A_HUmEwnRZ3_1),.din(n826));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n829_0(.douta(w_dff_A_kyZTZRFM8_0),.doutb(w_n829_0[1]),.din(n829));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(w_dff_B_wO10LduC0_2));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl jspl_w_n840_0(.douta(w_dff_A_8g1bLN284_0),.doutb(w_n840_0[1]),.din(n840));
	jspl3 jspl3_w_n844_0(.douta(w_n844_0[0]),.doutb(w_n844_0[1]),.doutc(w_n844_0[2]),.din(n844));
	jspl jspl_w_n846_0(.douta(w_n846_0[0]),.doutb(w_n846_0[1]),.din(w_dff_B_jU74dILT4_2));
	jspl jspl_w_n849_0(.douta(w_n849_0[0]),.doutb(w_n849_0[1]),.din(n849));
	jspl jspl_w_n851_0(.douta(w_n851_0[0]),.doutb(w_n851_0[1]),.din(w_dff_B_hS6AMZ2m3_2));
	jspl jspl_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.din(n854));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(w_dff_B_dJ60ay428_2));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(w_dff_B_bsFbhQmc0_2));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(w_dff_B_Iell99iK5_2));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(w_dff_B_22rxImAM4_2));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(n874));
	jspl jspl_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.din(w_dff_B_DFyjm9Ys5_2));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(w_dff_B_iSePcQlc6_2));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(w_dff_B_WSaq7kmt7_2));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(w_dff_B_3FIpdvcG0_2));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_dff_A_QgymNIau6_1),.din(n896));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(w_dff_B_Ycy7sUPW7_2));
	jspl jspl_w_n901_0(.douta(w_n901_0[0]),.doutb(w_n901_0[1]),.din(n901));
	jspl jspl_w_n903_0(.douta(w_dff_A_UYrp90wJ3_0),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n906_0(.douta(w_n906_0[0]),.doutb(w_n906_0[1]),.din(n906));
	jspl jspl_w_n907_0(.douta(w_n907_0[0]),.doutb(w_n907_0[1]),.din(w_dff_B_CF3fq3pc5_2));
	jspl jspl_w_n908_0(.douta(w_n908_0[0]),.doutb(w_n908_0[1]),.din(n908));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(w_dff_B_HJJXPDLJ1_2));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(n910));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(w_dff_B_r3cc26Gc8_2));
	jspl jspl_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.din(n912));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(w_dff_B_pK0UmoXy1_2));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.din(w_dff_B_znWFqW642_2));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(n916));
	jspl jspl_w_n917_0(.douta(w_n917_0[0]),.doutb(w_n917_0[1]),.din(w_dff_B_fIPyYPm37_2));
	jspl jspl_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.din(n918));
	jspl jspl_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.din(n919));
	jspl jspl_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.din(n920));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(w_dff_B_y0ItLKzh4_2));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(n924));
	jspl jspl_w_n925_0(.douta(w_n925_0[0]),.doutb(w_n925_0[1]),.din(w_dff_B_7XoFcijs1_2));
	jspl jspl_w_n926_0(.douta(w_n926_0[0]),.doutb(w_n926_0[1]),.din(n926));
	jspl3 jspl3_w_n927_0(.douta(w_n927_0[0]),.doutb(w_dff_A_3epEYrKA2_1),.doutc(w_dff_A_axzWNOhv0_2),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_dff_A_Oj2QZeXD0_1),.din(n929));
	jspl jspl_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.din(n930));
	jspl jspl_w_n931_0(.douta(w_n931_0[0]),.doutb(w_dff_A_rPD8mdkc9_1),.din(n931));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(w_dff_B_UgomcaYM9_2));
	jspl3 jspl3_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.doutc(w_n942_0[2]),.din(n942));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_n943_0[1]),.din(w_dff_B_OlErDkei0_2));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(n949));
	jspl jspl_w_n951_0(.douta(w_n951_0[0]),.doutb(w_n951_0[1]),.din(w_dff_B_AHIF6KrI3_2));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n956_0(.douta(w_n956_0[0]),.doutb(w_n956_0[1]),.din(w_dff_B_KSl44vcR5_2));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(n959));
	jspl jspl_w_n961_0(.douta(w_n961_0[0]),.doutb(w_n961_0[1]),.din(w_dff_B_vAKqYFTu3_2));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.din(w_dff_B_hSUeKmrL0_2));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_n971_0[1]),.din(w_dff_B_MjkJMhHw9_2));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n976_0(.douta(w_n976_0[0]),.doutb(w_n976_0[1]),.din(w_dff_B_g97xEijh0_2));
	jspl jspl_w_n979_0(.douta(w_n979_0[0]),.doutb(w_n979_0[1]),.din(n979));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(w_dff_B_thbvFUV31_2));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(w_dff_B_ZWgEyIQa3_2));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(w_dff_B_oOUT4ZHk3_2));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(w_dff_B_23rRmjYY1_2));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(w_dff_B_fFN9NgEZ6_2));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_dff_A_3cWmQLSM5_1),.din(n1006));
	jspl jspl_w_n1008_0(.douta(w_dff_A_N9UzwRK64_0),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1010_0(.douta(w_n1010_0[0]),.doutb(w_n1010_0[1]),.din(w_dff_B_WsuEKtQ94_2));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.din(w_dff_B_ok5zClye5_2));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl jspl_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.din(w_dff_B_BmViWpj58_2));
	jspl jspl_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.din(n1015));
	jspl jspl_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.din(w_dff_B_CvCblr1X9_2));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(w_dff_B_ao4BY8oo8_2));
	jspl jspl_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.din(n1019));
	jspl jspl_w_n1020_0(.douta(w_n1020_0[0]),.doutb(w_n1020_0[1]),.din(w_dff_B_FNpHUw6v3_2));
	jspl jspl_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.din(n1021));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.din(w_dff_B_BLi57DKT7_2));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(n1023));
	jspl jspl_w_n1024_0(.douta(w_n1024_0[0]),.doutb(w_n1024_0[1]),.din(n1024));
	jspl jspl_w_n1025_0(.douta(w_n1025_0[0]),.doutb(w_n1025_0[1]),.din(n1025));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1027_0(.douta(w_n1027_0[0]),.doutb(w_n1027_0[1]),.din(n1027));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(w_dff_B_n7NZzqfv9_2));
	jspl jspl_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.din(n1029));
	jspl jspl_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.din(w_dff_B_m3dEVGtb0_2));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_dff_A_rzHhCtPL6_1),.din(n1032));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1034_0(.douta(w_dff_A_IYu9QDqv2_0),.doutb(w_n1034_0[1]),.din(n1034));
	jspl jspl_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.din(n1035));
	jspl jspl_w_n1037_0(.douta(w_n1037_0[0]),.doutb(w_n1037_0[1]),.din(w_dff_B_sIVTiUs64_2));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_dff_A_8iyxgJFi0_1),.din(n1039));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(n1043));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(w_dff_B_aZrjLaUP2_2));
	jspl jspl_w_n1048_0(.douta(w_dff_A_kLeTUCqx2_0),.doutb(w_n1048_0[1]),.din(n1048));
	jspl jspl_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.din(w_dff_B_AbRIsUjF5_2));
	jspl jspl_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.din(w_dff_B_e94QfI5g5_2));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.din(n1057));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(w_dff_B_jgMd85UI9_2));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.din(n1062));
	jspl jspl_w_n1064_0(.douta(w_n1064_0[0]),.doutb(w_n1064_0[1]),.din(w_dff_B_K9MfCiiH9_2));
	jspl jspl_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.din(n1067));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(w_dff_B_QMuW436K2_2));
	jspl jspl_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.din(n1072));
	jspl jspl_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.din(w_dff_B_YDUtoW4R7_2));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(n1077));
	jspl jspl_w_n1079_0(.douta(w_n1079_0[0]),.doutb(w_n1079_0[1]),.din(w_dff_B_czjghiQe6_2));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(w_dff_B_E8f9MlnF1_2));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(n1087));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(w_dff_B_W4qd8b791_2));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(w_dff_B_ZfiCaKEH3_2));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(w_dff_B_ZwivAUV38_2));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(w_dff_B_hwGPVRFa1_2));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1110_0(.douta(w_dff_A_QejrMFgQ1_0),.doutb(w_n1110_0[1]),.din(w_dff_B_BWx1odqe4_2));
	jspl jspl_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.din(n1114));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.din(n1116));
	jspl jspl_w_n1117_0(.douta(w_n1117_0[0]),.doutb(w_n1117_0[1]),.din(w_dff_B_tsN5TVO52_2));
	jspl jspl_w_n1118_0(.douta(w_n1118_0[0]),.doutb(w_n1118_0[1]),.din(n1118));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(w_dff_B_6X1GQTtL4_2));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl jspl_w_n1121_0(.douta(w_n1121_0[0]),.doutb(w_n1121_0[1]),.din(w_dff_B_zGdvxZ9X5_2));
	jspl jspl_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.din(n1122));
	jspl jspl_w_n1123_0(.douta(w_n1123_0[0]),.doutb(w_n1123_0[1]),.din(w_dff_B_RuQq9Eub5_2));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.din(w_dff_B_EisvOOA97_2));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(n1126));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(w_dff_B_tK1POAiv8_2));
	jspl jspl_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.din(n1128));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(n1131));
	jspl jspl_w_n1132_0(.douta(w_n1132_0[0]),.doutb(w_n1132_0[1]),.din(n1132));
	jspl jspl_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.din(w_dff_B_5LD0MFNh0_2));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1135_0(.douta(w_n1135_0[0]),.doutb(w_n1135_0[1]),.din(w_dff_B_rdvUAVGU5_2));
	jspl jspl_w_n1137_0(.douta(w_n1137_0[0]),.doutb(w_n1137_0[1]),.din(n1137));
	jspl jspl_w_n1138_0(.douta(w_n1138_0[0]),.doutb(w_n1138_0[1]),.din(n1138));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1140_0(.douta(w_n1140_0[0]),.doutb(w_dff_A_Om9vCIER8_1),.din(n1140));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(n1141));
	jspl jspl_w_n1147_0(.douta(w_n1147_0[0]),.doutb(w_n1147_0[1]),.din(n1147));
	jspl jspl_w_n1151_0(.douta(w_dff_A_1qgBAHnM3_0),.doutb(w_n1151_0[1]),.din(w_dff_B_BmLhtFuJ1_2));
	jspl jspl_w_n1152_0(.douta(w_n1152_0[0]),.doutb(w_n1152_0[1]),.din(w_dff_B_OFFb5aQu2_2));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(n1156));
	jspl jspl_w_n1158_0(.douta(w_n1158_0[0]),.doutb(w_n1158_0[1]),.din(w_dff_B_2ErB38d85_2));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(n1161));
	jspl jspl_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.din(w_dff_B_7O8tEm8a3_2));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl jspl_w_n1168_0(.douta(w_n1168_0[0]),.doutb(w_n1168_0[1]),.din(w_dff_B_f2fXMfxO2_2));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(n1171));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(w_dff_B_Za3PwOC99_2));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(n1176));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.din(w_dff_B_xlGvVhf30_2));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(w_dff_B_IwuZxtfj9_2));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(n1186));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(w_dff_B_Qb35jaaX6_2));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(n1191));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(w_dff_B_3zLaC3ht5_2));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(w_dff_B_65EnfEbg5_2));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(w_dff_B_n8FDE26z7_2));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(w_dff_B_ZkUGvUdg8_2));
	jspl jspl_w_n1207_0(.douta(w_n1207_0[0]),.doutb(w_n1207_0[1]),.din(w_dff_B_Xn6nswdx1_2));
	jspl jspl_w_n1208_0(.douta(w_n1208_0[0]),.doutb(w_n1208_0[1]),.din(w_dff_B_TRYhdKbR3_2));
	jspl jspl_w_n1210_0(.douta(w_n1210_0[0]),.doutb(w_n1210_0[1]),.din(n1210));
	jspl jspl_w_n1212_0(.douta(w_n1212_0[0]),.doutb(w_n1212_0[1]),.din(n1212));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1214_0(.douta(w_n1214_0[0]),.doutb(w_n1214_0[1]),.din(n1214));
	jspl jspl_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.din(w_dff_B_OSqXrNmC5_2));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(w_dff_B_ajak31ho7_2));
	jspl jspl_w_n1218_0(.douta(w_n1218_0[0]),.doutb(w_n1218_0[1]),.din(n1218));
	jspl jspl_w_n1219_0(.douta(w_n1219_0[0]),.doutb(w_n1219_0[1]),.din(w_dff_B_26ORQgZm0_2));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1221_0(.douta(w_n1221_0[0]),.doutb(w_n1221_0[1]),.din(w_dff_B_rFjJMvLB6_2));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(n1222));
	jspl jspl_w_n1223_0(.douta(w_n1223_0[0]),.doutb(w_n1223_0[1]),.din(w_dff_B_dW6wxl6L3_2));
	jspl jspl_w_n1224_0(.douta(w_n1224_0[0]),.doutb(w_n1224_0[1]),.din(n1224));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(w_dff_B_AvICfoV98_2));
	jspl jspl_w_n1226_0(.douta(w_n1226_0[0]),.doutb(w_n1226_0[1]),.din(n1226));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(n1227));
	jspl jspl_w_n1228_0(.douta(w_n1228_0[0]),.doutb(w_n1228_0[1]),.din(n1228));
	jspl jspl_w_n1229_0(.douta(w_n1229_0[0]),.doutb(w_n1229_0[1]),.din(n1229));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1231_0(.douta(w_n1231_0[0]),.doutb(w_n1231_0[1]),.din(w_dff_B_mr1nHZhz7_2));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(n1232));
	jspl jspl_w_n1234_0(.douta(w_n1234_0[0]),.doutb(w_n1234_0[1]),.din(w_dff_B_QyiOm4660_2));
	jspl jspl_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(n1237));
	jspl jspl_w_n1238_0(.douta(w_dff_A_YtIxMlso6_0),.doutb(w_n1238_0[1]),.din(n1238));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(n1247));
	jspl jspl_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.din(w_dff_B_0xiW4LK49_2));
	jspl jspl_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.din(n1251));
	jspl jspl_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.din(w_dff_B_cOfaW6Mn8_2));
	jspl jspl_w_n1256_0(.douta(w_n1256_0[0]),.doutb(w_n1256_0[1]),.din(n1256));
	jspl jspl_w_n1258_0(.douta(w_n1258_0[0]),.doutb(w_n1258_0[1]),.din(w_dff_B_WDf10k9W8_2));
	jspl jspl_w_n1261_0(.douta(w_n1261_0[0]),.doutb(w_n1261_0[1]),.din(n1261));
	jspl jspl_w_n1263_0(.douta(w_n1263_0[0]),.doutb(w_n1263_0[1]),.din(w_dff_B_LczfR24N0_2));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(n1266));
	jspl jspl_w_n1268_0(.douta(w_n1268_0[0]),.doutb(w_n1268_0[1]),.din(w_dff_B_eC9RpPVU6_2));
	jspl jspl_w_n1271_0(.douta(w_n1271_0[0]),.doutb(w_n1271_0[1]),.din(n1271));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(w_dff_B_kFyMKoK27_2));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(n1276));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(w_dff_B_MuvFa1BM3_2));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(n1281));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(w_dff_B_LPIVmATe5_2));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(n1286));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(w_dff_B_sEnDKUqv7_2));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_n1291_0[1]),.din(n1291));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(w_dff_B_zz2U9j7y4_2));
	jspl jspl_w_n1296_0(.douta(w_n1296_0[0]),.doutb(w_n1296_0[1]),.din(w_dff_B_gXAYdozV7_2));
	jspl jspl_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.din(w_dff_B_l7vSSOB04_2));
	jspl jspl_w_n1298_0(.douta(w_n1298_0[0]),.doutb(w_n1298_0[1]),.din(w_dff_B_q0E3ocqJ8_2));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1303_0(.douta(w_n1303_0[0]),.doutb(w_n1303_0[1]),.din(n1303));
	jspl jspl_w_n1304_0(.douta(w_n1304_0[0]),.doutb(w_n1304_0[1]),.din(n1304));
	jspl jspl_w_n1305_0(.douta(w_n1305_0[0]),.doutb(w_n1305_0[1]),.din(n1305));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(n1307));
	jspl jspl_w_n1308_0(.douta(w_n1308_0[0]),.doutb(w_n1308_0[1]),.din(w_dff_B_sajY995T2_2));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(w_dff_B_KrtcCkho1_2));
	jspl jspl_w_n1311_0(.douta(w_n1311_0[0]),.doutb(w_n1311_0[1]),.din(n1311));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(w_dff_B_bBFQ8uv53_2));
	jspl jspl_w_n1313_0(.douta(w_n1313_0[0]),.doutb(w_n1313_0[1]),.din(n1313));
	jspl jspl_w_n1314_0(.douta(w_n1314_0[0]),.doutb(w_n1314_0[1]),.din(w_dff_B_2UwdX7bc2_2));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.din(w_dff_B_iqP04Ira2_2));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1318_0(.douta(w_n1318_0[0]),.doutb(w_n1318_0[1]),.din(n1318));
	jspl jspl_w_n1319_0(.douta(w_n1319_0[0]),.doutb(w_n1319_0[1]),.din(n1319));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.din(n1321));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_dff_A_w51f6fKg9_1),.din(n1322));
	jspl jspl_w_n1324_0(.douta(w_n1324_0[0]),.doutb(w_n1324_0[1]),.din(n1324));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_dff_A_YmfkltVR9_1),.din(n1325));
	jspl jspl_w_n1326_0(.douta(w_dff_A_Fc4YPKTA5_0),.doutb(w_n1326_0[1]),.din(n1326));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(n1332));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(n1337));
	jspl jspl_w_n1338_0(.douta(w_n1338_0[0]),.doutb(w_n1338_0[1]),.din(w_dff_B_1eQL6QIs8_2));
	jspl jspl_w_n1341_0(.douta(w_n1341_0[0]),.doutb(w_n1341_0[1]),.din(n1341));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(w_dff_B_48lD1CKl9_2));
	jspl jspl_w_n1346_0(.douta(w_n1346_0[0]),.doutb(w_n1346_0[1]),.din(n1346));
	jspl jspl_w_n1348_0(.douta(w_n1348_0[0]),.doutb(w_n1348_0[1]),.din(w_dff_B_mTGVb2Y87_2));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(n1351));
	jspl jspl_w_n1353_0(.douta(w_n1353_0[0]),.doutb(w_n1353_0[1]),.din(w_dff_B_4jwkYf7z2_2));
	jspl jspl_w_n1356_0(.douta(w_n1356_0[0]),.doutb(w_n1356_0[1]),.din(n1356));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(w_dff_B_5S7Cx1Wo0_2));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(w_dff_B_vCLHSOEX6_2));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(n1366));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(w_dff_B_dOjXQLHZ1_2));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(w_dff_B_Dq6CTl2L9_2));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(w_dff_B_IYIt1woL4_2));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(w_dff_B_1jCtZI1E6_2));
	jspl jspl_w_n1381_0(.douta(w_n1381_0[0]),.doutb(w_n1381_0[1]),.din(w_dff_B_Dh6JNuk36_2));
	jspl jspl_w_n1382_0(.douta(w_n1382_0[0]),.doutb(w_n1382_0[1]),.din(w_dff_B_k8Ala0aO3_2));
	jspl jspl_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.din(w_dff_B_1Mlva9xD5_2));
	jspl jspl_w_n1386_0(.douta(w_n1386_0[0]),.doutb(w_n1386_0[1]),.din(n1386));
	jspl jspl_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_n1388_0[1]),.din(n1388));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(n1389));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(n1390));
	jspl jspl_w_n1391_0(.douta(w_n1391_0[0]),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1392_0(.douta(w_n1392_0[0]),.doutb(w_n1392_0[1]),.din(n1392));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(w_dff_B_sSCut7rS2_2));
	jspl jspl_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.din(n1396));
	jspl jspl_w_n1397_0(.douta(w_n1397_0[0]),.doutb(w_n1397_0[1]),.din(w_dff_B_eRYndxZQ9_2));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(w_dff_B_Fjw6Mauc8_2));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(n1400));
	jspl jspl_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_n1401_0[1]),.din(w_dff_B_wRhOut4q0_2));
	jspl jspl_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_n1402_0[1]),.din(n1402));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_n1404_0[1]),.din(n1404));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl jspl_w_n1407_0(.douta(w_n1407_0[0]),.doutb(w_n1407_0[1]),.din(n1407));
	jspl jspl_w_n1409_0(.douta(w_n1409_0[0]),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_dff_A_lgICghwQ9_1),.din(n1410));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(n1415));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(w_dff_B_Cngn24uH1_2));
	jspl jspl_w_n1421_0(.douta(w_n1421_0[0]),.doutb(w_n1421_0[1]),.din(w_dff_B_Vzsvtm4e3_2));
	jspl jspl_w_n1424_0(.douta(w_n1424_0[0]),.doutb(w_n1424_0[1]),.din(n1424));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(w_dff_B_Z9LoOTDA7_2));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(w_dff_B_dZq68j420_2));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(w_dff_B_itcEa49g7_2));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(w_dff_B_Lm7RFGGj8_2));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(n1444));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(w_dff_B_StFokFFU0_2));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(w_dff_B_iLfpviWR0_2));
	jspl jspl_w_n1451_0(.douta(w_n1451_0[0]),.doutb(w_n1451_0[1]),.din(w_dff_B_1Nd5QAbS8_2));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(w_dff_B_hg36VsNB6_2));
	jspl jspl_w_n1456_0(.douta(w_n1456_0[0]),.doutb(w_n1456_0[1]),.din(w_dff_B_jxzYtriR6_2));
	jspl jspl_w_n1459_0(.douta(w_n1459_0[0]),.doutb(w_n1459_0[1]),.din(w_dff_B_eCwWw4tB1_2));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(w_dff_B_hYRIFJQP7_2));
	jspl jspl_w_n1461_0(.douta(w_n1461_0[0]),.doutb(w_n1461_0[1]),.din(w_dff_B_20Kyx2j61_2));
	jspl jspl_w_n1464_0(.douta(w_n1464_0[0]),.doutb(w_n1464_0[1]),.din(n1464));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(n1466));
	jspl jspl_w_n1467_0(.douta(w_n1467_0[0]),.doutb(w_n1467_0[1]),.din(n1467));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_n1468_0[1]),.din(n1468));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1470_0(.douta(w_n1470_0[0]),.doutb(w_n1470_0[1]),.din(n1470));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(n1471));
	jspl jspl_w_n1472_0(.douta(w_n1472_0[0]),.doutb(w_n1472_0[1]),.din(n1472));
	jspl jspl_w_n1473_0(.douta(w_n1473_0[0]),.doutb(w_n1473_0[1]),.din(n1473));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(n1474));
	jspl jspl_w_n1475_0(.douta(w_n1475_0[0]),.doutb(w_n1475_0[1]),.din(w_dff_B_bYfsVfi42_2));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(n1476));
	jspl jspl_w_n1477_0(.douta(w_n1477_0[0]),.doutb(w_n1477_0[1]),.din(w_dff_B_HDcp3aG34_2));
	jspl jspl_w_n1478_0(.douta(w_n1478_0[0]),.doutb(w_n1478_0[1]),.din(n1478));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(w_dff_B_8w6Vab4P0_2));
	jspl jspl_w_n1480_0(.douta(w_n1480_0[0]),.doutb(w_n1480_0[1]),.din(n1480));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(n1481));
	jspl jspl_w_n1483_0(.douta(w_n1483_0[0]),.doutb(w_n1483_0[1]),.din(n1483));
	jspl jspl_w_n1485_0(.douta(w_n1485_0[0]),.doutb(w_n1485_0[1]),.din(n1485));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_dff_A_6OXjizs55_1),.din(n1486));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(n1491));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(w_dff_B_a33fP2nu5_2));
	jspl jspl_w_n1497_0(.douta(w_n1497_0[0]),.doutb(w_n1497_0[1]),.din(w_dff_B_f5hCBJZx7_2));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(n1500));
	jspl jspl_w_n1502_0(.douta(w_n1502_0[0]),.doutb(w_n1502_0[1]),.din(w_dff_B_TV43XzgL1_2));
	jspl jspl_w_n1505_0(.douta(w_n1505_0[0]),.doutb(w_n1505_0[1]),.din(n1505));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(w_dff_B_4CzgkvPs3_2));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(w_dff_B_vWEqRT4V1_2));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(w_dff_B_IcO8rX5a7_2));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(w_dff_B_y9GIDU0I4_2));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.din(w_dff_B_uIocQ37G6_2));
	jspl jspl_w_n1522_0(.douta(w_n1522_0[0]),.doutb(w_n1522_0[1]),.din(w_dff_B_1Wmbdlxi2_2));
	jspl jspl_w_n1525_0(.douta(w_n1525_0[0]),.doutb(w_n1525_0[1]),.din(w_dff_B_JFgwEwTC7_2));
	jspl jspl_w_n1527_0(.douta(w_n1527_0[0]),.doutb(w_n1527_0[1]),.din(w_dff_B_e01CU9l05_2));
	jspl jspl_w_n1530_0(.douta(w_n1530_0[0]),.doutb(w_n1530_0[1]),.din(w_dff_B_J0E8nPgL3_2));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(w_dff_B_BLj5OV3O9_2));
	jspl jspl_w_n1532_0(.douta(w_n1532_0[0]),.doutb(w_n1532_0[1]),.din(w_dff_B_HTirBmXv6_2));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(n1535));
	jspl jspl_w_n1537_0(.douta(w_n1537_0[0]),.doutb(w_n1537_0[1]),.din(n1537));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.din(n1539));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(n1540));
	jspl jspl_w_n1541_0(.douta(w_n1541_0[0]),.doutb(w_n1541_0[1]),.din(n1541));
	jspl jspl_w_n1542_0(.douta(w_n1542_0[0]),.doutb(w_n1542_0[1]),.din(n1542));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1544_0(.douta(w_n1544_0[0]),.doutb(w_n1544_0[1]),.din(n1544));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1546_0(.douta(w_n1546_0[0]),.doutb(w_n1546_0[1]),.din(n1546));
	jspl jspl_w_n1547_0(.douta(w_n1547_0[0]),.doutb(w_n1547_0[1]),.din(n1547));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(w_dff_B_BwMT4r4s5_2));
	jspl jspl_w_n1549_0(.douta(w_n1549_0[0]),.doutb(w_n1549_0[1]),.din(n1549));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_dff_A_fK9qtCNH5_1),.din(n1550));
	jspl jspl_w_n1552_0(.douta(w_n1552_0[0]),.doutb(w_n1552_0[1]),.din(n1552));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_dff_A_GWaUef9G5_1),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(n1565));
	jspl jspl_w_n1566_0(.douta(w_n1566_0[0]),.doutb(w_n1566_0[1]),.din(w_dff_B_NFOVWNVB8_2));
	jspl jspl_w_n1569_0(.douta(w_n1569_0[0]),.doutb(w_n1569_0[1]),.din(n1569));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(w_dff_B_SsRb6lpj6_2));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(w_dff_B_2R8NMV0v3_2));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(w_dff_B_ZP7WsaNU0_2));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(w_dff_B_diTzV2yZ9_2));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_n1581_0[1]),.din(w_dff_B_Sddow3bz4_2));
	jspl jspl_w_n1584_0(.douta(w_n1584_0[0]),.doutb(w_n1584_0[1]),.din(w_dff_B_LAskapZm5_2));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.din(w_dff_B_OncjjOTl6_2));
	jspl jspl_w_n1589_0(.douta(w_n1589_0[0]),.doutb(w_n1589_0[1]),.din(w_dff_B_nlDQTvOA9_2));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(w_dff_B_8WbYio3T6_2));
	jspl jspl_w_n1594_0(.douta(w_n1594_0[0]),.doutb(w_n1594_0[1]),.din(w_dff_B_DoJLaGXc5_2));
	jspl jspl_w_n1595_0(.douta(w_n1595_0[0]),.doutb(w_n1595_0[1]),.din(w_dff_B_fpEPPbdR3_2));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(w_dff_B_b1k1UvD19_2));
	jspl jspl_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_n1603_0[1]),.din(n1603));
	jspl jspl_w_n1604_0(.douta(w_n1604_0[0]),.doutb(w_n1604_0[1]),.din(n1604));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1606_0(.douta(w_n1606_0[0]),.doutb(w_n1606_0[1]),.din(n1606));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1608_0(.douta(w_n1608_0[0]),.doutb(w_n1608_0[1]),.din(n1608));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.din(n1611));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(n1612));
	jspl jspl_w_n1614_0(.douta(w_n1614_0[0]),.doutb(w_n1614_0[1]),.din(n1614));
	jspl jspl_w_n1616_0(.douta(w_n1616_0[0]),.doutb(w_n1616_0[1]),.din(n1616));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_dff_A_IMnnVenA9_1),.din(n1617));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(n1622));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(w_dff_B_eA7aoaMJ9_2));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(w_dff_B_okOZllCj2_2));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_dff_A_Wswiurrn4_1),.din(n1631));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(w_dff_B_vDxlcce85_2));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(w_dff_B_uIBjKJe90_2));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(w_dff_B_dz0k26vB2_2));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_n1641_0[1]),.din(w_dff_B_tEmEHAdO5_2));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(w_dff_B_pLG9O1LA0_2));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(w_dff_B_sWdREgKP8_2));
	jspl jspl_w_n1648_0(.douta(w_n1648_0[0]),.doutb(w_n1648_0[1]),.din(w_dff_B_rQO4g00b5_2));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(w_dff_B_NRAchYUb4_2));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_n1652_0[1]),.din(w_dff_B_2q3rfz6I1_2));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(w_dff_B_4fxGLIjY0_2));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(n1656));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(n1658));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1660_0(.douta(w_n1660_0[0]),.doutb(w_n1660_0[1]),.din(n1660));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(n1661));
	jspl jspl_w_n1662_0(.douta(w_n1662_0[0]),.doutb(w_n1662_0[1]),.din(n1662));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(n1663));
	jspl jspl_w_n1664_0(.douta(w_n1664_0[0]),.doutb(w_n1664_0[1]),.din(n1664));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(n1666));
	jspl jspl_w_n1667_0(.douta(w_n1667_0[0]),.doutb(w_n1667_0[1]),.din(n1667));
	jspl jspl_w_n1669_0(.douta(w_n1669_0[0]),.doutb(w_n1669_0[1]),.din(n1669));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(n1671));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_dff_A_7o8BL2rh8_1),.din(n1672));
	jspl jspl_w_n1677_0(.douta(w_n1677_0[0]),.doutb(w_n1677_0[1]),.din(n1677));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(w_dff_B_AsdTUFM99_2));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(w_dff_B_Md1qSbaj1_2));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_n1687_0[1]),.din(w_dff_B_GZgJyiDF4_2));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(w_dff_B_wWyQm1T04_2));
	jspl jspl_w_n1692_0(.douta(w_n1692_0[0]),.doutb(w_n1692_0[1]),.din(w_dff_B_EzRe3tCe8_2));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(w_dff_B_Eg9FkntX4_2));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_n1697_0[1]),.din(w_dff_B_j8LajU4o8_2));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(w_dff_B_0DfkFQY61_2));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(w_dff_B_jmMqyqcm9_2));
	jspl jspl_w_n1703_0(.douta(w_n1703_0[0]),.doutb(w_n1703_0[1]),.din(w_dff_B_Yf9oaDTh0_2));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(w_dff_B_GMBo0y002_2));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(n1707));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(n1709));
	jspl jspl_w_n1710_0(.douta(w_n1710_0[0]),.doutb(w_n1710_0[1]),.din(n1710));
	jspl jspl_w_n1711_0(.douta(w_n1711_0[0]),.doutb(w_n1711_0[1]),.din(n1711));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(n1712));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(n1713));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(n1714));
	jspl jspl_w_n1715_0(.douta(w_n1715_0[0]),.doutb(w_n1715_0[1]),.din(n1715));
	jspl jspl_w_n1716_0(.douta(w_n1716_0[0]),.doutb(w_n1716_0[1]),.din(n1716));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_dff_A_HV3sCXwW3_1),.din(n1720));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1728_0(.douta(w_n1728_0[0]),.doutb(w_dff_A_KO0EuAWu9_1),.din(n1728));
	jspl jspl_w_n1730_0(.douta(w_n1730_0[0]),.doutb(w_n1730_0[1]),.din(w_dff_B_YqZFdzjd8_2));
	jspl jspl_w_n1733_0(.douta(w_n1733_0[0]),.doutb(w_n1733_0[1]),.din(w_dff_B_eWqtMJtR2_2));
	jspl jspl_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.din(w_dff_B_jlXX2w2d4_2));
	jspl jspl_w_n1738_0(.douta(w_n1738_0[0]),.doutb(w_n1738_0[1]),.din(w_dff_B_4bnrSVb15_2));
	jspl jspl_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.din(w_dff_B_3kFUTehD8_2));
	jspl jspl_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.din(w_dff_B_2E4qR4cc6_2));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(w_dff_B_ziA82jg42_2));
	jspl jspl_w_n1745_0(.douta(w_n1745_0[0]),.doutb(w_n1745_0[1]),.din(w_dff_B_kT7sBeMi1_2));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(n1748));
	jspl jspl_w_n1750_0(.douta(w_n1750_0[0]),.doutb(w_n1750_0[1]),.din(n1750));
	jspl jspl_w_n1751_0(.douta(w_n1751_0[0]),.doutb(w_n1751_0[1]),.din(n1751));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1753_0(.douta(w_n1753_0[0]),.doutb(w_n1753_0[1]),.din(n1753));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_dff_A_E6PWdTsO3_1),.din(n1758));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl jspl_w_n1768_0(.douta(w_n1768_0[0]),.doutb(w_dff_A_9n7XV7sv6_1),.din(n1768));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(w_dff_B_ZmKqx6aG2_2));
	jspl jspl_w_n1773_0(.douta(w_n1773_0[0]),.doutb(w_n1773_0[1]),.din(w_dff_B_LyBfnB659_2));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(w_dff_B_D4NOgbEQ5_2));
	jspl jspl_w_n1778_0(.douta(w_n1778_0[0]),.doutb(w_n1778_0[1]),.din(w_dff_B_nodTVjh30_2));
	jspl jspl_w_n1779_0(.douta(w_n1779_0[0]),.doutb(w_n1779_0[1]),.din(w_dff_B_BBmT6JTF2_2));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(w_dff_B_Pk8E9oz23_2));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_n1786_0[1]),.din(n1786));
	jspl jspl_w_n1787_0(.douta(w_n1787_0[0]),.doutb(w_n1787_0[1]),.din(n1787));
	jspl jspl_w_n1788_0(.douta(w_n1788_0[0]),.doutb(w_n1788_0[1]),.din(n1788));
	jspl jspl_w_n1789_0(.douta(w_n1789_0[0]),.doutb(w_n1789_0[1]),.din(n1789));
	jspl jspl_w_n1790_0(.douta(w_n1790_0[0]),.doutb(w_n1790_0[1]),.din(n1790));
	jspl jspl_w_n1791_0(.douta(w_n1791_0[0]),.doutb(w_dff_A_xi9bByvv3_1),.din(n1791));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(n1798));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_dff_A_forErhb54_1),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(w_dff_B_BDl4KhBR6_2));
	jspl jspl_w_n1806_0(.douta(w_n1806_0[0]),.doutb(w_n1806_0[1]),.din(w_dff_B_MHVvfctY5_2));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(w_dff_B_cMF3AuPD1_2));
	jspl jspl_w_n1808_0(.douta(w_n1808_0[0]),.doutb(w_n1808_0[1]),.din(w_dff_B_liKzinUN3_2));
	jspl jspl_w_n1811_0(.douta(w_n1811_0[0]),.doutb(w_n1811_0[1]),.din(n1811));
	jspl jspl_w_n1813_0(.douta(w_n1813_0[0]),.doutb(w_n1813_0[1]),.din(n1813));
	jspl jspl_w_n1814_0(.douta(w_n1814_0[0]),.doutb(w_n1814_0[1]),.din(n1814));
	jspl jspl_w_n1815_0(.douta(w_n1815_0[0]),.doutb(w_n1815_0[1]),.din(n1815));
	jspl jspl_w_n1816_0(.douta(w_n1816_0[0]),.doutb(w_n1816_0[1]),.din(n1816));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_dff_A_2B9FjQxb3_1),.din(n1817));
	jspl jspl_w_n1824_0(.douta(w_n1824_0[0]),.doutb(w_n1824_0[1]),.din(n1824));
	jspl jspl_w_n1827_0(.douta(w_n1827_0[0]),.doutb(w_dff_A_PxkUvdjD5_1),.din(n1827));
	jspl jspl_w_n1828_0(.douta(w_n1828_0[0]),.doutb(w_n1828_0[1]),.din(w_dff_B_LrVQ6VMx0_2));
	jspl jspl_w_n1829_0(.douta(w_n1829_0[0]),.doutb(w_n1829_0[1]),.din(w_dff_B_JpaPDBvt5_2));
	jspl jspl_w_n1832_0(.douta(w_n1832_0[0]),.doutb(w_n1832_0[1]),.din(n1832));
	jspl jspl_w_n1834_0(.douta(w_n1834_0[0]),.doutb(w_n1834_0[1]),.din(n1834));
	jspl jspl_w_n1835_0(.douta(w_n1835_0[0]),.doutb(w_n1835_0[1]),.din(n1835));
	jspl jspl_w_n1836_0(.douta(w_n1836_0[0]),.doutb(w_dff_A_zIOHEaBV8_1),.din(n1836));
	jspl jspl_w_n1838_0(.douta(w_n1838_0[0]),.doutb(w_n1838_0[1]),.din(w_dff_B_ePcqAiRz6_2));
	jspl jspl_w_n1841_0(.douta(w_n1841_0[0]),.doutb(w_n1841_0[1]),.din(n1841));
	jspl jspl_w_n1848_0(.douta(w_n1848_0[0]),.doutb(w_n1848_0[1]),.din(n1848));
	jspl jspl_w_n1849_0(.douta(w_dff_A_S3oaBWKP4_0),.doutb(w_n1849_0[1]),.din(n1849));
	jdff dff_B_FlnRawTX7_1(.din(n67),.dout(w_dff_B_FlnRawTX7_1),.clk(gclk));
	jdff dff_B_wCMHpDOi5_1(.din(n73),.dout(w_dff_B_wCMHpDOi5_1),.clk(gclk));
	jdff dff_B_sdJfy7uL5_1(.din(w_dff_B_wCMHpDOi5_1),.dout(w_dff_B_sdJfy7uL5_1),.clk(gclk));
	jdff dff_B_STxbppBs3_1(.din(w_dff_B_sdJfy7uL5_1),.dout(w_dff_B_STxbppBs3_1),.clk(gclk));
	jdff dff_B_HbMs7I9A8_1(.din(w_dff_B_STxbppBs3_1),.dout(w_dff_B_HbMs7I9A8_1),.clk(gclk));
	jdff dff_B_60O3SjDB7_1(.din(n90),.dout(w_dff_B_60O3SjDB7_1),.clk(gclk));
	jdff dff_B_ERxjwXja7_1(.din(w_dff_B_60O3SjDB7_1),.dout(w_dff_B_ERxjwXja7_1),.clk(gclk));
	jdff dff_B_0F0VZf8u2_1(.din(w_dff_B_ERxjwXja7_1),.dout(w_dff_B_0F0VZf8u2_1),.clk(gclk));
	jdff dff_B_Lr8oXvTq9_1(.din(w_dff_B_0F0VZf8u2_1),.dout(w_dff_B_Lr8oXvTq9_1),.clk(gclk));
	jdff dff_B_ilYyFsgQ3_1(.din(w_dff_B_Lr8oXvTq9_1),.dout(w_dff_B_ilYyFsgQ3_1),.clk(gclk));
	jdff dff_B_4iotCQpn5_1(.din(w_dff_B_ilYyFsgQ3_1),.dout(w_dff_B_4iotCQpn5_1),.clk(gclk));
	jdff dff_B_Zp5c4yA99_1(.din(w_dff_B_4iotCQpn5_1),.dout(w_dff_B_Zp5c4yA99_1),.clk(gclk));
	jdff dff_B_rRivL0kd8_1(.din(n111),.dout(w_dff_B_rRivL0kd8_1),.clk(gclk));
	jdff dff_B_SJSr3X7k5_1(.din(w_dff_B_rRivL0kd8_1),.dout(w_dff_B_SJSr3X7k5_1),.clk(gclk));
	jdff dff_B_VvhWuhwe8_1(.din(w_dff_B_SJSr3X7k5_1),.dout(w_dff_B_VvhWuhwe8_1),.clk(gclk));
	jdff dff_B_aSgInQzn5_1(.din(w_dff_B_VvhWuhwe8_1),.dout(w_dff_B_aSgInQzn5_1),.clk(gclk));
	jdff dff_B_IIVETUCY5_1(.din(w_dff_B_aSgInQzn5_1),.dout(w_dff_B_IIVETUCY5_1),.clk(gclk));
	jdff dff_B_O86EOvnT3_1(.din(w_dff_B_IIVETUCY5_1),.dout(w_dff_B_O86EOvnT3_1),.clk(gclk));
	jdff dff_B_Gufbg2BB4_1(.din(w_dff_B_O86EOvnT3_1),.dout(w_dff_B_Gufbg2BB4_1),.clk(gclk));
	jdff dff_B_zjxJOgeN3_1(.din(w_dff_B_Gufbg2BB4_1),.dout(w_dff_B_zjxJOgeN3_1),.clk(gclk));
	jdff dff_B_gl7VcSe70_1(.din(w_dff_B_zjxJOgeN3_1),.dout(w_dff_B_gl7VcSe70_1),.clk(gclk));
	jdff dff_B_oWExCNQ75_1(.din(w_dff_B_gl7VcSe70_1),.dout(w_dff_B_oWExCNQ75_1),.clk(gclk));
	jdff dff_B_vtS2lXxj3_1(.din(n146),.dout(w_dff_B_vtS2lXxj3_1),.clk(gclk));
	jdff dff_B_UbgYM5jy7_1(.din(w_dff_B_vtS2lXxj3_1),.dout(w_dff_B_UbgYM5jy7_1),.clk(gclk));
	jdff dff_B_T2EdSbCF4_1(.din(w_dff_B_UbgYM5jy7_1),.dout(w_dff_B_T2EdSbCF4_1),.clk(gclk));
	jdff dff_B_G9KAKXTI4_1(.din(w_dff_B_T2EdSbCF4_1),.dout(w_dff_B_G9KAKXTI4_1),.clk(gclk));
	jdff dff_B_BCjl6DfE9_1(.din(w_dff_B_G9KAKXTI4_1),.dout(w_dff_B_BCjl6DfE9_1),.clk(gclk));
	jdff dff_B_shKcgyAq3_1(.din(w_dff_B_BCjl6DfE9_1),.dout(w_dff_B_shKcgyAq3_1),.clk(gclk));
	jdff dff_B_1fo167qq5_1(.din(w_dff_B_shKcgyAq3_1),.dout(w_dff_B_1fo167qq5_1),.clk(gclk));
	jdff dff_B_DsEquqky4_1(.din(w_dff_B_1fo167qq5_1),.dout(w_dff_B_DsEquqky4_1),.clk(gclk));
	jdff dff_B_Iw9Bbdmu3_1(.din(w_dff_B_DsEquqky4_1),.dout(w_dff_B_Iw9Bbdmu3_1),.clk(gclk));
	jdff dff_B_4593GmyZ5_1(.din(w_dff_B_Iw9Bbdmu3_1),.dout(w_dff_B_4593GmyZ5_1),.clk(gclk));
	jdff dff_B_8BOnlKVH7_1(.din(w_dff_B_4593GmyZ5_1),.dout(w_dff_B_8BOnlKVH7_1),.clk(gclk));
	jdff dff_B_9sJ4FH923_1(.din(w_dff_B_8BOnlKVH7_1),.dout(w_dff_B_9sJ4FH923_1),.clk(gclk));
	jdff dff_B_nEJzxkY00_1(.din(w_dff_B_9sJ4FH923_1),.dout(w_dff_B_nEJzxkY00_1),.clk(gclk));
	jdff dff_B_6Q1zjGBA2_1(.din(n184),.dout(w_dff_B_6Q1zjGBA2_1),.clk(gclk));
	jdff dff_B_sLWALcqO7_1(.din(w_dff_B_6Q1zjGBA2_1),.dout(w_dff_B_sLWALcqO7_1),.clk(gclk));
	jdff dff_B_VGKpUuhp3_1(.din(w_dff_B_sLWALcqO7_1),.dout(w_dff_B_VGKpUuhp3_1),.clk(gclk));
	jdff dff_B_SXvicOZ97_1(.din(w_dff_B_VGKpUuhp3_1),.dout(w_dff_B_SXvicOZ97_1),.clk(gclk));
	jdff dff_B_8nFYkbrA6_1(.din(w_dff_B_SXvicOZ97_1),.dout(w_dff_B_8nFYkbrA6_1),.clk(gclk));
	jdff dff_B_brptCj5c0_1(.din(w_dff_B_8nFYkbrA6_1),.dout(w_dff_B_brptCj5c0_1),.clk(gclk));
	jdff dff_B_R31P1xF99_1(.din(w_dff_B_brptCj5c0_1),.dout(w_dff_B_R31P1xF99_1),.clk(gclk));
	jdff dff_B_5oPOPCIv2_1(.din(w_dff_B_R31P1xF99_1),.dout(w_dff_B_5oPOPCIv2_1),.clk(gclk));
	jdff dff_B_MKZEa4wR8_1(.din(w_dff_B_5oPOPCIv2_1),.dout(w_dff_B_MKZEa4wR8_1),.clk(gclk));
	jdff dff_B_DBHOqC0l8_1(.din(w_dff_B_MKZEa4wR8_1),.dout(w_dff_B_DBHOqC0l8_1),.clk(gclk));
	jdff dff_B_B3Z3reUi3_1(.din(w_dff_B_DBHOqC0l8_1),.dout(w_dff_B_B3Z3reUi3_1),.clk(gclk));
	jdff dff_B_Ak2Bm4ee3_1(.din(w_dff_B_B3Z3reUi3_1),.dout(w_dff_B_Ak2Bm4ee3_1),.clk(gclk));
	jdff dff_B_3F6TGqKX7_1(.din(w_dff_B_Ak2Bm4ee3_1),.dout(w_dff_B_3F6TGqKX7_1),.clk(gclk));
	jdff dff_B_9fUtzQSP0_1(.din(w_dff_B_3F6TGqKX7_1),.dout(w_dff_B_9fUtzQSP0_1),.clk(gclk));
	jdff dff_B_wDHTkjfr6_1(.din(w_dff_B_9fUtzQSP0_1),.dout(w_dff_B_wDHTkjfr6_1),.clk(gclk));
	jdff dff_B_YCIsNlDY6_1(.din(w_dff_B_wDHTkjfr6_1),.dout(w_dff_B_YCIsNlDY6_1),.clk(gclk));
	jdff dff_B_whqYXsbT0_1(.din(n227),.dout(w_dff_B_whqYXsbT0_1),.clk(gclk));
	jdff dff_B_S96bL5oT8_1(.din(w_dff_B_whqYXsbT0_1),.dout(w_dff_B_S96bL5oT8_1),.clk(gclk));
	jdff dff_B_EaGbqYTL1_1(.din(w_dff_B_S96bL5oT8_1),.dout(w_dff_B_EaGbqYTL1_1),.clk(gclk));
	jdff dff_B_PI3bVm1B4_1(.din(w_dff_B_EaGbqYTL1_1),.dout(w_dff_B_PI3bVm1B4_1),.clk(gclk));
	jdff dff_B_qqi9RPW07_1(.din(w_dff_B_PI3bVm1B4_1),.dout(w_dff_B_qqi9RPW07_1),.clk(gclk));
	jdff dff_B_dzhTTeFT2_1(.din(w_dff_B_qqi9RPW07_1),.dout(w_dff_B_dzhTTeFT2_1),.clk(gclk));
	jdff dff_B_CuLD6BCu9_1(.din(w_dff_B_dzhTTeFT2_1),.dout(w_dff_B_CuLD6BCu9_1),.clk(gclk));
	jdff dff_B_cLVzMxuz2_1(.din(w_dff_B_CuLD6BCu9_1),.dout(w_dff_B_cLVzMxuz2_1),.clk(gclk));
	jdff dff_B_B2XPbEAQ1_1(.din(w_dff_B_cLVzMxuz2_1),.dout(w_dff_B_B2XPbEAQ1_1),.clk(gclk));
	jdff dff_B_uO8pLFjw1_1(.din(w_dff_B_B2XPbEAQ1_1),.dout(w_dff_B_uO8pLFjw1_1),.clk(gclk));
	jdff dff_B_m5IUpABs2_1(.din(w_dff_B_uO8pLFjw1_1),.dout(w_dff_B_m5IUpABs2_1),.clk(gclk));
	jdff dff_B_dmF44GG68_1(.din(w_dff_B_m5IUpABs2_1),.dout(w_dff_B_dmF44GG68_1),.clk(gclk));
	jdff dff_B_5gBjBoyz1_1(.din(w_dff_B_dmF44GG68_1),.dout(w_dff_B_5gBjBoyz1_1),.clk(gclk));
	jdff dff_B_u41Sj2Aq7_1(.din(w_dff_B_5gBjBoyz1_1),.dout(w_dff_B_u41Sj2Aq7_1),.clk(gclk));
	jdff dff_B_wYKy2GAs8_1(.din(w_dff_B_u41Sj2Aq7_1),.dout(w_dff_B_wYKy2GAs8_1),.clk(gclk));
	jdff dff_B_05xGj70w6_1(.din(w_dff_B_wYKy2GAs8_1),.dout(w_dff_B_05xGj70w6_1),.clk(gclk));
	jdff dff_B_ykSk5iGP3_1(.din(w_dff_B_05xGj70w6_1),.dout(w_dff_B_ykSk5iGP3_1),.clk(gclk));
	jdff dff_B_6aNrz2ZU6_1(.din(w_dff_B_ykSk5iGP3_1),.dout(w_dff_B_6aNrz2ZU6_1),.clk(gclk));
	jdff dff_B_rVL77JfP0_1(.din(w_dff_B_6aNrz2ZU6_1),.dout(w_dff_B_rVL77JfP0_1),.clk(gclk));
	jdff dff_B_a2zzzpxG1_1(.din(n278),.dout(w_dff_B_a2zzzpxG1_1),.clk(gclk));
	jdff dff_B_0lqUBRAk6_1(.din(w_dff_B_a2zzzpxG1_1),.dout(w_dff_B_0lqUBRAk6_1),.clk(gclk));
	jdff dff_B_q0MGXqm38_1(.din(w_dff_B_0lqUBRAk6_1),.dout(w_dff_B_q0MGXqm38_1),.clk(gclk));
	jdff dff_B_dsNivNOQ9_1(.din(w_dff_B_q0MGXqm38_1),.dout(w_dff_B_dsNivNOQ9_1),.clk(gclk));
	jdff dff_B_Iwv3UNpM2_1(.din(w_dff_B_dsNivNOQ9_1),.dout(w_dff_B_Iwv3UNpM2_1),.clk(gclk));
	jdff dff_B_2gRP9Kha2_1(.din(w_dff_B_Iwv3UNpM2_1),.dout(w_dff_B_2gRP9Kha2_1),.clk(gclk));
	jdff dff_B_SbEy35GQ2_1(.din(w_dff_B_2gRP9Kha2_1),.dout(w_dff_B_SbEy35GQ2_1),.clk(gclk));
	jdff dff_B_MHas7a3Z4_1(.din(w_dff_B_SbEy35GQ2_1),.dout(w_dff_B_MHas7a3Z4_1),.clk(gclk));
	jdff dff_B_SsfSV83S3_1(.din(w_dff_B_MHas7a3Z4_1),.dout(w_dff_B_SsfSV83S3_1),.clk(gclk));
	jdff dff_B_VJ4NDuJq5_1(.din(w_dff_B_SsfSV83S3_1),.dout(w_dff_B_VJ4NDuJq5_1),.clk(gclk));
	jdff dff_B_3xCvqsgU0_1(.din(w_dff_B_VJ4NDuJq5_1),.dout(w_dff_B_3xCvqsgU0_1),.clk(gclk));
	jdff dff_B_Hvnz8wtV3_1(.din(w_dff_B_3xCvqsgU0_1),.dout(w_dff_B_Hvnz8wtV3_1),.clk(gclk));
	jdff dff_B_GRHxvnvb1_1(.din(w_dff_B_Hvnz8wtV3_1),.dout(w_dff_B_GRHxvnvb1_1),.clk(gclk));
	jdff dff_B_copsStCz9_1(.din(w_dff_B_GRHxvnvb1_1),.dout(w_dff_B_copsStCz9_1),.clk(gclk));
	jdff dff_B_g54p5iyo6_1(.din(w_dff_B_copsStCz9_1),.dout(w_dff_B_g54p5iyo6_1),.clk(gclk));
	jdff dff_B_IaJhPYqY2_1(.din(w_dff_B_g54p5iyo6_1),.dout(w_dff_B_IaJhPYqY2_1),.clk(gclk));
	jdff dff_B_kyPMqsYh0_1(.din(w_dff_B_IaJhPYqY2_1),.dout(w_dff_B_kyPMqsYh0_1),.clk(gclk));
	jdff dff_B_W6V02sKH1_1(.din(w_dff_B_kyPMqsYh0_1),.dout(w_dff_B_W6V02sKH1_1),.clk(gclk));
	jdff dff_B_gzhWT1iK0_1(.din(w_dff_B_W6V02sKH1_1),.dout(w_dff_B_gzhWT1iK0_1),.clk(gclk));
	jdff dff_B_AmtNKtQH0_1(.din(w_dff_B_gzhWT1iK0_1),.dout(w_dff_B_AmtNKtQH0_1),.clk(gclk));
	jdff dff_B_TNbf3rd33_1(.din(w_dff_B_AmtNKtQH0_1),.dout(w_dff_B_TNbf3rd33_1),.clk(gclk));
	jdff dff_B_oH3KqGwB4_1(.din(w_dff_B_TNbf3rd33_1),.dout(w_dff_B_oH3KqGwB4_1),.clk(gclk));
	jdff dff_B_wEIEdFzp5_1(.din(n336),.dout(w_dff_B_wEIEdFzp5_1),.clk(gclk));
	jdff dff_B_7QXIm5Yn0_1(.din(w_dff_B_wEIEdFzp5_1),.dout(w_dff_B_7QXIm5Yn0_1),.clk(gclk));
	jdff dff_B_oYSEhs1h1_1(.din(w_dff_B_7QXIm5Yn0_1),.dout(w_dff_B_oYSEhs1h1_1),.clk(gclk));
	jdff dff_B_NxNILxUd8_1(.din(w_dff_B_oYSEhs1h1_1),.dout(w_dff_B_NxNILxUd8_1),.clk(gclk));
	jdff dff_B_cWchFx2B2_1(.din(w_dff_B_NxNILxUd8_1),.dout(w_dff_B_cWchFx2B2_1),.clk(gclk));
	jdff dff_B_Saglca3F8_1(.din(w_dff_B_cWchFx2B2_1),.dout(w_dff_B_Saglca3F8_1),.clk(gclk));
	jdff dff_B_dyXn8XrA1_1(.din(w_dff_B_Saglca3F8_1),.dout(w_dff_B_dyXn8XrA1_1),.clk(gclk));
	jdff dff_B_ZbQhgMU97_1(.din(w_dff_B_dyXn8XrA1_1),.dout(w_dff_B_ZbQhgMU97_1),.clk(gclk));
	jdff dff_B_Aax07fdp0_1(.din(w_dff_B_ZbQhgMU97_1),.dout(w_dff_B_Aax07fdp0_1),.clk(gclk));
	jdff dff_B_1vQ5ORq25_1(.din(w_dff_B_Aax07fdp0_1),.dout(w_dff_B_1vQ5ORq25_1),.clk(gclk));
	jdff dff_B_CjQAJZ9z5_1(.din(w_dff_B_1vQ5ORq25_1),.dout(w_dff_B_CjQAJZ9z5_1),.clk(gclk));
	jdff dff_B_ZE1xVrXg4_1(.din(w_dff_B_CjQAJZ9z5_1),.dout(w_dff_B_ZE1xVrXg4_1),.clk(gclk));
	jdff dff_B_Fa4hIdED2_1(.din(w_dff_B_ZE1xVrXg4_1),.dout(w_dff_B_Fa4hIdED2_1),.clk(gclk));
	jdff dff_B_WUvc9dgb7_1(.din(w_dff_B_Fa4hIdED2_1),.dout(w_dff_B_WUvc9dgb7_1),.clk(gclk));
	jdff dff_B_h1ZqDlFJ3_1(.din(w_dff_B_WUvc9dgb7_1),.dout(w_dff_B_h1ZqDlFJ3_1),.clk(gclk));
	jdff dff_B_KFiCfCiN7_1(.din(w_dff_B_h1ZqDlFJ3_1),.dout(w_dff_B_KFiCfCiN7_1),.clk(gclk));
	jdff dff_B_c2Igsh980_1(.din(w_dff_B_KFiCfCiN7_1),.dout(w_dff_B_c2Igsh980_1),.clk(gclk));
	jdff dff_B_OXCMwMYx9_1(.din(w_dff_B_c2Igsh980_1),.dout(w_dff_B_OXCMwMYx9_1),.clk(gclk));
	jdff dff_B_Xs4uT3ic5_1(.din(w_dff_B_OXCMwMYx9_1),.dout(w_dff_B_Xs4uT3ic5_1),.clk(gclk));
	jdff dff_B_UxQEuFzx7_1(.din(w_dff_B_Xs4uT3ic5_1),.dout(w_dff_B_UxQEuFzx7_1),.clk(gclk));
	jdff dff_B_V23efQt70_1(.din(w_dff_B_UxQEuFzx7_1),.dout(w_dff_B_V23efQt70_1),.clk(gclk));
	jdff dff_B_a2Q06y577_1(.din(w_dff_B_V23efQt70_1),.dout(w_dff_B_a2Q06y577_1),.clk(gclk));
	jdff dff_B_p4C8DXdO9_1(.din(w_dff_B_a2Q06y577_1),.dout(w_dff_B_p4C8DXdO9_1),.clk(gclk));
	jdff dff_B_AlgJPJUD7_1(.din(w_dff_B_p4C8DXdO9_1),.dout(w_dff_B_AlgJPJUD7_1),.clk(gclk));
	jdff dff_B_piHzdoiB6_1(.din(w_dff_B_AlgJPJUD7_1),.dout(w_dff_B_piHzdoiB6_1),.clk(gclk));
	jdff dff_B_twgeBedW1_1(.din(n400),.dout(w_dff_B_twgeBedW1_1),.clk(gclk));
	jdff dff_B_wxuHUL808_1(.din(w_dff_B_twgeBedW1_1),.dout(w_dff_B_wxuHUL808_1),.clk(gclk));
	jdff dff_B_EiKE7WDD1_1(.din(w_dff_B_wxuHUL808_1),.dout(w_dff_B_EiKE7WDD1_1),.clk(gclk));
	jdff dff_B_mcgllPVV0_1(.din(w_dff_B_EiKE7WDD1_1),.dout(w_dff_B_mcgllPVV0_1),.clk(gclk));
	jdff dff_B_mi42vg061_1(.din(w_dff_B_mcgllPVV0_1),.dout(w_dff_B_mi42vg061_1),.clk(gclk));
	jdff dff_B_sylcrNYg0_1(.din(w_dff_B_mi42vg061_1),.dout(w_dff_B_sylcrNYg0_1),.clk(gclk));
	jdff dff_B_s9HluGJc9_1(.din(w_dff_B_sylcrNYg0_1),.dout(w_dff_B_s9HluGJc9_1),.clk(gclk));
	jdff dff_B_9oAPPFJD4_1(.din(w_dff_B_s9HluGJc9_1),.dout(w_dff_B_9oAPPFJD4_1),.clk(gclk));
	jdff dff_B_r1BgwDeh7_1(.din(w_dff_B_9oAPPFJD4_1),.dout(w_dff_B_r1BgwDeh7_1),.clk(gclk));
	jdff dff_B_keb4xBe01_1(.din(w_dff_B_r1BgwDeh7_1),.dout(w_dff_B_keb4xBe01_1),.clk(gclk));
	jdff dff_B_PmQBQZJ82_1(.din(w_dff_B_keb4xBe01_1),.dout(w_dff_B_PmQBQZJ82_1),.clk(gclk));
	jdff dff_B_EXJ4tpse4_1(.din(w_dff_B_PmQBQZJ82_1),.dout(w_dff_B_EXJ4tpse4_1),.clk(gclk));
	jdff dff_B_XXn03XVt7_1(.din(w_dff_B_EXJ4tpse4_1),.dout(w_dff_B_XXn03XVt7_1),.clk(gclk));
	jdff dff_B_L2Do306Q9_1(.din(w_dff_B_XXn03XVt7_1),.dout(w_dff_B_L2Do306Q9_1),.clk(gclk));
	jdff dff_B_bWAoU4x65_1(.din(w_dff_B_L2Do306Q9_1),.dout(w_dff_B_bWAoU4x65_1),.clk(gclk));
	jdff dff_B_ak3ovxsm3_1(.din(w_dff_B_bWAoU4x65_1),.dout(w_dff_B_ak3ovxsm3_1),.clk(gclk));
	jdff dff_B_fK0Zv3Bt1_1(.din(w_dff_B_ak3ovxsm3_1),.dout(w_dff_B_fK0Zv3Bt1_1),.clk(gclk));
	jdff dff_B_zR2l0qQX4_1(.din(w_dff_B_fK0Zv3Bt1_1),.dout(w_dff_B_zR2l0qQX4_1),.clk(gclk));
	jdff dff_B_7vS8L6GY2_1(.din(w_dff_B_zR2l0qQX4_1),.dout(w_dff_B_7vS8L6GY2_1),.clk(gclk));
	jdff dff_B_gRLERNxY0_1(.din(w_dff_B_7vS8L6GY2_1),.dout(w_dff_B_gRLERNxY0_1),.clk(gclk));
	jdff dff_B_qkHWLBlB4_1(.din(w_dff_B_gRLERNxY0_1),.dout(w_dff_B_qkHWLBlB4_1),.clk(gclk));
	jdff dff_B_PybMpjAB1_1(.din(w_dff_B_qkHWLBlB4_1),.dout(w_dff_B_PybMpjAB1_1),.clk(gclk));
	jdff dff_B_HFhK5X3L2_1(.din(w_dff_B_PybMpjAB1_1),.dout(w_dff_B_HFhK5X3L2_1),.clk(gclk));
	jdff dff_B_kOkW5tSF7_1(.din(w_dff_B_HFhK5X3L2_1),.dout(w_dff_B_kOkW5tSF7_1),.clk(gclk));
	jdff dff_B_mkB5CaAJ5_1(.din(w_dff_B_kOkW5tSF7_1),.dout(w_dff_B_mkB5CaAJ5_1),.clk(gclk));
	jdff dff_B_1HiSq3Lm1_1(.din(w_dff_B_mkB5CaAJ5_1),.dout(w_dff_B_1HiSq3Lm1_1),.clk(gclk));
	jdff dff_B_NBLTAN7Q0_1(.din(w_dff_B_1HiSq3Lm1_1),.dout(w_dff_B_NBLTAN7Q0_1),.clk(gclk));
	jdff dff_B_erQVcywS2_1(.din(w_dff_B_NBLTAN7Q0_1),.dout(w_dff_B_erQVcywS2_1),.clk(gclk));
	jdff dff_B_NYGj0Y1o1_1(.din(n472),.dout(w_dff_B_NYGj0Y1o1_1),.clk(gclk));
	jdff dff_B_IldXXGwX6_1(.din(w_dff_B_NYGj0Y1o1_1),.dout(w_dff_B_IldXXGwX6_1),.clk(gclk));
	jdff dff_B_QYrHQz6Q2_1(.din(w_dff_B_IldXXGwX6_1),.dout(w_dff_B_QYrHQz6Q2_1),.clk(gclk));
	jdff dff_B_ILTw8DYX2_1(.din(w_dff_B_QYrHQz6Q2_1),.dout(w_dff_B_ILTw8DYX2_1),.clk(gclk));
	jdff dff_B_hjRQWfnk3_1(.din(w_dff_B_ILTw8DYX2_1),.dout(w_dff_B_hjRQWfnk3_1),.clk(gclk));
	jdff dff_B_A2p1NaP77_1(.din(w_dff_B_hjRQWfnk3_1),.dout(w_dff_B_A2p1NaP77_1),.clk(gclk));
	jdff dff_B_sCTWq8G43_1(.din(w_dff_B_A2p1NaP77_1),.dout(w_dff_B_sCTWq8G43_1),.clk(gclk));
	jdff dff_B_yA6YbsKe0_1(.din(w_dff_B_sCTWq8G43_1),.dout(w_dff_B_yA6YbsKe0_1),.clk(gclk));
	jdff dff_B_yT2TeJI65_1(.din(w_dff_B_yA6YbsKe0_1),.dout(w_dff_B_yT2TeJI65_1),.clk(gclk));
	jdff dff_B_gZqqw59y5_1(.din(w_dff_B_yT2TeJI65_1),.dout(w_dff_B_gZqqw59y5_1),.clk(gclk));
	jdff dff_B_qcdJzEly7_1(.din(w_dff_B_gZqqw59y5_1),.dout(w_dff_B_qcdJzEly7_1),.clk(gclk));
	jdff dff_B_GSQHUgRC2_1(.din(w_dff_B_qcdJzEly7_1),.dout(w_dff_B_GSQHUgRC2_1),.clk(gclk));
	jdff dff_B_OkR3p2hZ6_1(.din(w_dff_B_GSQHUgRC2_1),.dout(w_dff_B_OkR3p2hZ6_1),.clk(gclk));
	jdff dff_B_fhJQTi3w3_1(.din(w_dff_B_OkR3p2hZ6_1),.dout(w_dff_B_fhJQTi3w3_1),.clk(gclk));
	jdff dff_B_vdgutqrR8_1(.din(w_dff_B_fhJQTi3w3_1),.dout(w_dff_B_vdgutqrR8_1),.clk(gclk));
	jdff dff_B_yHJfLbJI9_1(.din(w_dff_B_vdgutqrR8_1),.dout(w_dff_B_yHJfLbJI9_1),.clk(gclk));
	jdff dff_B_SljHnOOY0_1(.din(w_dff_B_yHJfLbJI9_1),.dout(w_dff_B_SljHnOOY0_1),.clk(gclk));
	jdff dff_B_lJKQxDEb3_1(.din(w_dff_B_SljHnOOY0_1),.dout(w_dff_B_lJKQxDEb3_1),.clk(gclk));
	jdff dff_B_Wl3a5Hia0_1(.din(w_dff_B_lJKQxDEb3_1),.dout(w_dff_B_Wl3a5Hia0_1),.clk(gclk));
	jdff dff_B_3Ry4I1MU7_1(.din(w_dff_B_Wl3a5Hia0_1),.dout(w_dff_B_3Ry4I1MU7_1),.clk(gclk));
	jdff dff_B_I7q5oAJW0_1(.din(w_dff_B_3Ry4I1MU7_1),.dout(w_dff_B_I7q5oAJW0_1),.clk(gclk));
	jdff dff_B_ryj4xiuG5_1(.din(w_dff_B_I7q5oAJW0_1),.dout(w_dff_B_ryj4xiuG5_1),.clk(gclk));
	jdff dff_B_FkILoM930_1(.din(w_dff_B_ryj4xiuG5_1),.dout(w_dff_B_FkILoM930_1),.clk(gclk));
	jdff dff_B_4OpwQnyS8_1(.din(w_dff_B_FkILoM930_1),.dout(w_dff_B_4OpwQnyS8_1),.clk(gclk));
	jdff dff_B_BtFzJvlK8_1(.din(w_dff_B_4OpwQnyS8_1),.dout(w_dff_B_BtFzJvlK8_1),.clk(gclk));
	jdff dff_B_xevlMDq26_1(.din(w_dff_B_BtFzJvlK8_1),.dout(w_dff_B_xevlMDq26_1),.clk(gclk));
	jdff dff_B_DCzy1yr71_1(.din(w_dff_B_xevlMDq26_1),.dout(w_dff_B_DCzy1yr71_1),.clk(gclk));
	jdff dff_B_ttirPb0p5_1(.din(w_dff_B_DCzy1yr71_1),.dout(w_dff_B_ttirPb0p5_1),.clk(gclk));
	jdff dff_B_V6OycExF9_1(.din(w_dff_B_ttirPb0p5_1),.dout(w_dff_B_V6OycExF9_1),.clk(gclk));
	jdff dff_B_d4Dqqnfg6_1(.din(w_dff_B_V6OycExF9_1),.dout(w_dff_B_d4Dqqnfg6_1),.clk(gclk));
	jdff dff_B_OwwZINRB0_1(.din(w_dff_B_d4Dqqnfg6_1),.dout(w_dff_B_OwwZINRB0_1),.clk(gclk));
	jdff dff_B_ktBhtVTz7_1(.din(n551),.dout(w_dff_B_ktBhtVTz7_1),.clk(gclk));
	jdff dff_B_RzNlVu1r1_1(.din(w_dff_B_ktBhtVTz7_1),.dout(w_dff_B_RzNlVu1r1_1),.clk(gclk));
	jdff dff_B_HLDLkxPu9_1(.din(w_dff_B_RzNlVu1r1_1),.dout(w_dff_B_HLDLkxPu9_1),.clk(gclk));
	jdff dff_B_gtQXxrHa1_1(.din(w_dff_B_HLDLkxPu9_1),.dout(w_dff_B_gtQXxrHa1_1),.clk(gclk));
	jdff dff_B_8aA5e3yu7_1(.din(w_dff_B_gtQXxrHa1_1),.dout(w_dff_B_8aA5e3yu7_1),.clk(gclk));
	jdff dff_B_6rM5mEZx0_1(.din(w_dff_B_8aA5e3yu7_1),.dout(w_dff_B_6rM5mEZx0_1),.clk(gclk));
	jdff dff_B_N1FIAjYu3_1(.din(w_dff_B_6rM5mEZx0_1),.dout(w_dff_B_N1FIAjYu3_1),.clk(gclk));
	jdff dff_B_uuZLULmc9_1(.din(w_dff_B_N1FIAjYu3_1),.dout(w_dff_B_uuZLULmc9_1),.clk(gclk));
	jdff dff_B_y39mqIOx5_1(.din(w_dff_B_uuZLULmc9_1),.dout(w_dff_B_y39mqIOx5_1),.clk(gclk));
	jdff dff_B_N66UojaU8_1(.din(w_dff_B_y39mqIOx5_1),.dout(w_dff_B_N66UojaU8_1),.clk(gclk));
	jdff dff_B_kzgJ6SHl0_1(.din(w_dff_B_N66UojaU8_1),.dout(w_dff_B_kzgJ6SHl0_1),.clk(gclk));
	jdff dff_B_aW1bQlwx5_1(.din(w_dff_B_kzgJ6SHl0_1),.dout(w_dff_B_aW1bQlwx5_1),.clk(gclk));
	jdff dff_B_DCsPMNPK1_1(.din(w_dff_B_aW1bQlwx5_1),.dout(w_dff_B_DCsPMNPK1_1),.clk(gclk));
	jdff dff_B_VPO3duGm6_1(.din(w_dff_B_DCsPMNPK1_1),.dout(w_dff_B_VPO3duGm6_1),.clk(gclk));
	jdff dff_B_ObMTLEoV8_1(.din(w_dff_B_VPO3duGm6_1),.dout(w_dff_B_ObMTLEoV8_1),.clk(gclk));
	jdff dff_B_yqQPOCkE4_1(.din(w_dff_B_ObMTLEoV8_1),.dout(w_dff_B_yqQPOCkE4_1),.clk(gclk));
	jdff dff_B_etbc91OF2_1(.din(w_dff_B_yqQPOCkE4_1),.dout(w_dff_B_etbc91OF2_1),.clk(gclk));
	jdff dff_B_BPzNYXxU8_1(.din(w_dff_B_etbc91OF2_1),.dout(w_dff_B_BPzNYXxU8_1),.clk(gclk));
	jdff dff_B_YRzLklgY1_1(.din(w_dff_B_BPzNYXxU8_1),.dout(w_dff_B_YRzLklgY1_1),.clk(gclk));
	jdff dff_B_THBOFXCS7_1(.din(w_dff_B_YRzLklgY1_1),.dout(w_dff_B_THBOFXCS7_1),.clk(gclk));
	jdff dff_B_LwRIqg1o0_1(.din(w_dff_B_THBOFXCS7_1),.dout(w_dff_B_LwRIqg1o0_1),.clk(gclk));
	jdff dff_B_wfSShkjz8_1(.din(w_dff_B_LwRIqg1o0_1),.dout(w_dff_B_wfSShkjz8_1),.clk(gclk));
	jdff dff_B_ongBu5qs5_1(.din(w_dff_B_wfSShkjz8_1),.dout(w_dff_B_ongBu5qs5_1),.clk(gclk));
	jdff dff_B_sYEdVRJL3_1(.din(w_dff_B_ongBu5qs5_1),.dout(w_dff_B_sYEdVRJL3_1),.clk(gclk));
	jdff dff_B_ZAAZaKp33_1(.din(w_dff_B_sYEdVRJL3_1),.dout(w_dff_B_ZAAZaKp33_1),.clk(gclk));
	jdff dff_B_WV6TQTm70_1(.din(w_dff_B_ZAAZaKp33_1),.dout(w_dff_B_WV6TQTm70_1),.clk(gclk));
	jdff dff_B_IdOjdoJ26_1(.din(w_dff_B_WV6TQTm70_1),.dout(w_dff_B_IdOjdoJ26_1),.clk(gclk));
	jdff dff_B_qw3yPsm44_1(.din(w_dff_B_IdOjdoJ26_1),.dout(w_dff_B_qw3yPsm44_1),.clk(gclk));
	jdff dff_B_ZDiVBwSW1_1(.din(w_dff_B_qw3yPsm44_1),.dout(w_dff_B_ZDiVBwSW1_1),.clk(gclk));
	jdff dff_B_OYW74MFD7_1(.din(w_dff_B_ZDiVBwSW1_1),.dout(w_dff_B_OYW74MFD7_1),.clk(gclk));
	jdff dff_B_82QcN2bB2_1(.din(w_dff_B_OYW74MFD7_1),.dout(w_dff_B_82QcN2bB2_1),.clk(gclk));
	jdff dff_B_F9V7fWIk4_1(.din(w_dff_B_82QcN2bB2_1),.dout(w_dff_B_F9V7fWIk4_1),.clk(gclk));
	jdff dff_B_y9UtJkD21_1(.din(w_dff_B_F9V7fWIk4_1),.dout(w_dff_B_y9UtJkD21_1),.clk(gclk));
	jdff dff_B_kK36N8uP3_1(.din(w_dff_B_y9UtJkD21_1),.dout(w_dff_B_kK36N8uP3_1),.clk(gclk));
	jdff dff_B_ZEYgtjty0_1(.din(n637),.dout(w_dff_B_ZEYgtjty0_1),.clk(gclk));
	jdff dff_B_oqDz8hAC1_1(.din(w_dff_B_ZEYgtjty0_1),.dout(w_dff_B_oqDz8hAC1_1),.clk(gclk));
	jdff dff_B_unukIL8g8_1(.din(w_dff_B_oqDz8hAC1_1),.dout(w_dff_B_unukIL8g8_1),.clk(gclk));
	jdff dff_B_LNj8l2Mm3_1(.din(w_dff_B_unukIL8g8_1),.dout(w_dff_B_LNj8l2Mm3_1),.clk(gclk));
	jdff dff_B_rpPXZwUs2_1(.din(w_dff_B_LNj8l2Mm3_1),.dout(w_dff_B_rpPXZwUs2_1),.clk(gclk));
	jdff dff_B_sSMNNu0M6_1(.din(w_dff_B_rpPXZwUs2_1),.dout(w_dff_B_sSMNNu0M6_1),.clk(gclk));
	jdff dff_B_VbDqiQwg3_1(.din(w_dff_B_sSMNNu0M6_1),.dout(w_dff_B_VbDqiQwg3_1),.clk(gclk));
	jdff dff_B_ozUNbSNK1_1(.din(w_dff_B_VbDqiQwg3_1),.dout(w_dff_B_ozUNbSNK1_1),.clk(gclk));
	jdff dff_B_98Shzfw17_1(.din(w_dff_B_ozUNbSNK1_1),.dout(w_dff_B_98Shzfw17_1),.clk(gclk));
	jdff dff_B_2IY5qGhI4_1(.din(w_dff_B_98Shzfw17_1),.dout(w_dff_B_2IY5qGhI4_1),.clk(gclk));
	jdff dff_B_SLvFabNq4_1(.din(w_dff_B_2IY5qGhI4_1),.dout(w_dff_B_SLvFabNq4_1),.clk(gclk));
	jdff dff_B_qxZSQcba9_1(.din(w_dff_B_SLvFabNq4_1),.dout(w_dff_B_qxZSQcba9_1),.clk(gclk));
	jdff dff_B_KJsQRmJY9_1(.din(w_dff_B_qxZSQcba9_1),.dout(w_dff_B_KJsQRmJY9_1),.clk(gclk));
	jdff dff_B_Xn7QxX964_1(.din(w_dff_B_KJsQRmJY9_1),.dout(w_dff_B_Xn7QxX964_1),.clk(gclk));
	jdff dff_B_mXNgArBm6_1(.din(w_dff_B_Xn7QxX964_1),.dout(w_dff_B_mXNgArBm6_1),.clk(gclk));
	jdff dff_B_x0SIfecO0_1(.din(w_dff_B_mXNgArBm6_1),.dout(w_dff_B_x0SIfecO0_1),.clk(gclk));
	jdff dff_B_3Pfl5ZEQ4_1(.din(w_dff_B_x0SIfecO0_1),.dout(w_dff_B_3Pfl5ZEQ4_1),.clk(gclk));
	jdff dff_B_m51UgDzc6_1(.din(w_dff_B_3Pfl5ZEQ4_1),.dout(w_dff_B_m51UgDzc6_1),.clk(gclk));
	jdff dff_B_XIa552yP9_1(.din(w_dff_B_m51UgDzc6_1),.dout(w_dff_B_XIa552yP9_1),.clk(gclk));
	jdff dff_B_tzj67nvd6_1(.din(w_dff_B_XIa552yP9_1),.dout(w_dff_B_tzj67nvd6_1),.clk(gclk));
	jdff dff_B_Nanzewwn2_1(.din(w_dff_B_tzj67nvd6_1),.dout(w_dff_B_Nanzewwn2_1),.clk(gclk));
	jdff dff_B_3yRAxRhV6_1(.din(w_dff_B_Nanzewwn2_1),.dout(w_dff_B_3yRAxRhV6_1),.clk(gclk));
	jdff dff_B_DZXN19Ym3_1(.din(w_dff_B_3yRAxRhV6_1),.dout(w_dff_B_DZXN19Ym3_1),.clk(gclk));
	jdff dff_B_6XQ7hKEd0_1(.din(w_dff_B_DZXN19Ym3_1),.dout(w_dff_B_6XQ7hKEd0_1),.clk(gclk));
	jdff dff_B_ckUrSzjC9_1(.din(w_dff_B_6XQ7hKEd0_1),.dout(w_dff_B_ckUrSzjC9_1),.clk(gclk));
	jdff dff_B_gS1NIQse5_1(.din(w_dff_B_ckUrSzjC9_1),.dout(w_dff_B_gS1NIQse5_1),.clk(gclk));
	jdff dff_B_X5qHLXuE6_1(.din(w_dff_B_gS1NIQse5_1),.dout(w_dff_B_X5qHLXuE6_1),.clk(gclk));
	jdff dff_B_TsvRSnEh7_1(.din(w_dff_B_X5qHLXuE6_1),.dout(w_dff_B_TsvRSnEh7_1),.clk(gclk));
	jdff dff_B_FcIdlVHP6_1(.din(w_dff_B_TsvRSnEh7_1),.dout(w_dff_B_FcIdlVHP6_1),.clk(gclk));
	jdff dff_B_y53I3yOU9_1(.din(w_dff_B_FcIdlVHP6_1),.dout(w_dff_B_y53I3yOU9_1),.clk(gclk));
	jdff dff_B_EY0OYSmp4_1(.din(w_dff_B_y53I3yOU9_1),.dout(w_dff_B_EY0OYSmp4_1),.clk(gclk));
	jdff dff_B_gvARfhkR2_1(.din(w_dff_B_EY0OYSmp4_1),.dout(w_dff_B_gvARfhkR2_1),.clk(gclk));
	jdff dff_B_NpKctRtW2_1(.din(w_dff_B_gvARfhkR2_1),.dout(w_dff_B_NpKctRtW2_1),.clk(gclk));
	jdff dff_B_0E9cUlez9_1(.din(w_dff_B_NpKctRtW2_1),.dout(w_dff_B_0E9cUlez9_1),.clk(gclk));
	jdff dff_B_ibRxwUPP8_1(.din(w_dff_B_0E9cUlez9_1),.dout(w_dff_B_ibRxwUPP8_1),.clk(gclk));
	jdff dff_B_xs3BxYij3_1(.din(w_dff_B_ibRxwUPP8_1),.dout(w_dff_B_xs3BxYij3_1),.clk(gclk));
	jdff dff_B_r8jvjtir1_1(.din(w_dff_B_xs3BxYij3_1),.dout(w_dff_B_r8jvjtir1_1),.clk(gclk));
	jdff dff_B_kaDOa3CU8_1(.din(n730),.dout(w_dff_B_kaDOa3CU8_1),.clk(gclk));
	jdff dff_B_BPW3frcf6_1(.din(w_dff_B_kaDOa3CU8_1),.dout(w_dff_B_BPW3frcf6_1),.clk(gclk));
	jdff dff_B_7kNDhn4b4_1(.din(w_dff_B_BPW3frcf6_1),.dout(w_dff_B_7kNDhn4b4_1),.clk(gclk));
	jdff dff_B_8ScdTIkO8_1(.din(w_dff_B_7kNDhn4b4_1),.dout(w_dff_B_8ScdTIkO8_1),.clk(gclk));
	jdff dff_B_zHPOdMG66_1(.din(w_dff_B_8ScdTIkO8_1),.dout(w_dff_B_zHPOdMG66_1),.clk(gclk));
	jdff dff_B_nZJqR1a20_1(.din(w_dff_B_zHPOdMG66_1),.dout(w_dff_B_nZJqR1a20_1),.clk(gclk));
	jdff dff_B_XnphZwK74_1(.din(w_dff_B_nZJqR1a20_1),.dout(w_dff_B_XnphZwK74_1),.clk(gclk));
	jdff dff_B_3voclOSs7_1(.din(w_dff_B_XnphZwK74_1),.dout(w_dff_B_3voclOSs7_1),.clk(gclk));
	jdff dff_B_O2kuxKOs0_1(.din(w_dff_B_3voclOSs7_1),.dout(w_dff_B_O2kuxKOs0_1),.clk(gclk));
	jdff dff_B_xpL578oA7_1(.din(w_dff_B_O2kuxKOs0_1),.dout(w_dff_B_xpL578oA7_1),.clk(gclk));
	jdff dff_B_USkmvQ2t4_1(.din(w_dff_B_xpL578oA7_1),.dout(w_dff_B_USkmvQ2t4_1),.clk(gclk));
	jdff dff_B_zIZtKdkO8_1(.din(w_dff_B_USkmvQ2t4_1),.dout(w_dff_B_zIZtKdkO8_1),.clk(gclk));
	jdff dff_B_REkL5Tur8_1(.din(w_dff_B_zIZtKdkO8_1),.dout(w_dff_B_REkL5Tur8_1),.clk(gclk));
	jdff dff_B_XcsPeYpc6_1(.din(w_dff_B_REkL5Tur8_1),.dout(w_dff_B_XcsPeYpc6_1),.clk(gclk));
	jdff dff_B_0xOEg74p3_1(.din(w_dff_B_XcsPeYpc6_1),.dout(w_dff_B_0xOEg74p3_1),.clk(gclk));
	jdff dff_B_ONtpKoir0_1(.din(w_dff_B_0xOEg74p3_1),.dout(w_dff_B_ONtpKoir0_1),.clk(gclk));
	jdff dff_B_8OQ14b2L7_1(.din(w_dff_B_ONtpKoir0_1),.dout(w_dff_B_8OQ14b2L7_1),.clk(gclk));
	jdff dff_B_G9KYFOPh5_1(.din(w_dff_B_8OQ14b2L7_1),.dout(w_dff_B_G9KYFOPh5_1),.clk(gclk));
	jdff dff_B_uQRYcA7X6_1(.din(w_dff_B_G9KYFOPh5_1),.dout(w_dff_B_uQRYcA7X6_1),.clk(gclk));
	jdff dff_B_kbomD1TL5_1(.din(w_dff_B_uQRYcA7X6_1),.dout(w_dff_B_kbomD1TL5_1),.clk(gclk));
	jdff dff_B_ArfNz0o08_1(.din(w_dff_B_kbomD1TL5_1),.dout(w_dff_B_ArfNz0o08_1),.clk(gclk));
	jdff dff_B_T7YQxieu8_1(.din(w_dff_B_ArfNz0o08_1),.dout(w_dff_B_T7YQxieu8_1),.clk(gclk));
	jdff dff_B_3kBdBnNv0_1(.din(w_dff_B_T7YQxieu8_1),.dout(w_dff_B_3kBdBnNv0_1),.clk(gclk));
	jdff dff_B_dCiJrYpe1_1(.din(w_dff_B_3kBdBnNv0_1),.dout(w_dff_B_dCiJrYpe1_1),.clk(gclk));
	jdff dff_B_dAEAkRyB1_1(.din(w_dff_B_dCiJrYpe1_1),.dout(w_dff_B_dAEAkRyB1_1),.clk(gclk));
	jdff dff_B_6MefftY48_1(.din(w_dff_B_dAEAkRyB1_1),.dout(w_dff_B_6MefftY48_1),.clk(gclk));
	jdff dff_B_JKi06wMq4_1(.din(w_dff_B_6MefftY48_1),.dout(w_dff_B_JKi06wMq4_1),.clk(gclk));
	jdff dff_B_JezrVyNm5_1(.din(w_dff_B_JKi06wMq4_1),.dout(w_dff_B_JezrVyNm5_1),.clk(gclk));
	jdff dff_B_ebkeY8eE6_1(.din(w_dff_B_JezrVyNm5_1),.dout(w_dff_B_ebkeY8eE6_1),.clk(gclk));
	jdff dff_B_1KXdIPwK7_1(.din(w_dff_B_ebkeY8eE6_1),.dout(w_dff_B_1KXdIPwK7_1),.clk(gclk));
	jdff dff_B_wG01vPSr8_1(.din(w_dff_B_1KXdIPwK7_1),.dout(w_dff_B_wG01vPSr8_1),.clk(gclk));
	jdff dff_B_2qgeSkaM3_1(.din(w_dff_B_wG01vPSr8_1),.dout(w_dff_B_2qgeSkaM3_1),.clk(gclk));
	jdff dff_B_3JBG7tbr1_1(.din(w_dff_B_2qgeSkaM3_1),.dout(w_dff_B_3JBG7tbr1_1),.clk(gclk));
	jdff dff_B_nImkeq1M7_1(.din(w_dff_B_3JBG7tbr1_1),.dout(w_dff_B_nImkeq1M7_1),.clk(gclk));
	jdff dff_B_TkuOc68t9_1(.din(w_dff_B_nImkeq1M7_1),.dout(w_dff_B_TkuOc68t9_1),.clk(gclk));
	jdff dff_B_ZwTUEMLH1_1(.din(w_dff_B_TkuOc68t9_1),.dout(w_dff_B_ZwTUEMLH1_1),.clk(gclk));
	jdff dff_B_m7MKIcwi0_1(.din(w_dff_B_ZwTUEMLH1_1),.dout(w_dff_B_m7MKIcwi0_1),.clk(gclk));
	jdff dff_B_DxUyB6ww3_1(.din(w_dff_B_m7MKIcwi0_1),.dout(w_dff_B_DxUyB6ww3_1),.clk(gclk));
	jdff dff_B_OfJVT3ax0_1(.din(w_dff_B_DxUyB6ww3_1),.dout(w_dff_B_OfJVT3ax0_1),.clk(gclk));
	jdff dff_B_eVLHXhof4_1(.din(w_dff_B_OfJVT3ax0_1),.dout(w_dff_B_eVLHXhof4_1),.clk(gclk));
	jdff dff_B_0HGfBFmk8_1(.din(n830),.dout(w_dff_B_0HGfBFmk8_1),.clk(gclk));
	jdff dff_B_B7Ah3vti3_1(.din(w_dff_B_0HGfBFmk8_1),.dout(w_dff_B_B7Ah3vti3_1),.clk(gclk));
	jdff dff_B_tolJagxi0_1(.din(w_dff_B_B7Ah3vti3_1),.dout(w_dff_B_tolJagxi0_1),.clk(gclk));
	jdff dff_B_yfR3WOZH0_1(.din(w_dff_B_tolJagxi0_1),.dout(w_dff_B_yfR3WOZH0_1),.clk(gclk));
	jdff dff_B_ZD3T5Btk8_1(.din(w_dff_B_yfR3WOZH0_1),.dout(w_dff_B_ZD3T5Btk8_1),.clk(gclk));
	jdff dff_B_eHHOcdQg9_1(.din(w_dff_B_ZD3T5Btk8_1),.dout(w_dff_B_eHHOcdQg9_1),.clk(gclk));
	jdff dff_B_MzMZgsoR4_1(.din(w_dff_B_eHHOcdQg9_1),.dout(w_dff_B_MzMZgsoR4_1),.clk(gclk));
	jdff dff_B_zPTnjEN10_1(.din(w_dff_B_MzMZgsoR4_1),.dout(w_dff_B_zPTnjEN10_1),.clk(gclk));
	jdff dff_B_9IgSwGIK9_1(.din(w_dff_B_zPTnjEN10_1),.dout(w_dff_B_9IgSwGIK9_1),.clk(gclk));
	jdff dff_B_lBw163TE5_1(.din(w_dff_B_9IgSwGIK9_1),.dout(w_dff_B_lBw163TE5_1),.clk(gclk));
	jdff dff_B_bNjQ7o7w2_1(.din(w_dff_B_lBw163TE5_1),.dout(w_dff_B_bNjQ7o7w2_1),.clk(gclk));
	jdff dff_B_7LdLhKzY1_1(.din(w_dff_B_bNjQ7o7w2_1),.dout(w_dff_B_7LdLhKzY1_1),.clk(gclk));
	jdff dff_B_bKqTumec4_1(.din(w_dff_B_7LdLhKzY1_1),.dout(w_dff_B_bKqTumec4_1),.clk(gclk));
	jdff dff_B_FFdO61uq1_1(.din(w_dff_B_bKqTumec4_1),.dout(w_dff_B_FFdO61uq1_1),.clk(gclk));
	jdff dff_B_HHMDA5zG7_1(.din(w_dff_B_FFdO61uq1_1),.dout(w_dff_B_HHMDA5zG7_1),.clk(gclk));
	jdff dff_B_gyYYBCfy4_1(.din(w_dff_B_HHMDA5zG7_1),.dout(w_dff_B_gyYYBCfy4_1),.clk(gclk));
	jdff dff_B_wi7HRvc36_1(.din(w_dff_B_gyYYBCfy4_1),.dout(w_dff_B_wi7HRvc36_1),.clk(gclk));
	jdff dff_B_el9pkpPi1_1(.din(w_dff_B_wi7HRvc36_1),.dout(w_dff_B_el9pkpPi1_1),.clk(gclk));
	jdff dff_B_llOe2NHT7_1(.din(w_dff_B_el9pkpPi1_1),.dout(w_dff_B_llOe2NHT7_1),.clk(gclk));
	jdff dff_B_cR8OxUy66_1(.din(w_dff_B_llOe2NHT7_1),.dout(w_dff_B_cR8OxUy66_1),.clk(gclk));
	jdff dff_B_ML6Af0WK5_1(.din(w_dff_B_cR8OxUy66_1),.dout(w_dff_B_ML6Af0WK5_1),.clk(gclk));
	jdff dff_B_n7lek9Bk3_1(.din(w_dff_B_ML6Af0WK5_1),.dout(w_dff_B_n7lek9Bk3_1),.clk(gclk));
	jdff dff_B_6kHImbUL5_1(.din(w_dff_B_n7lek9Bk3_1),.dout(w_dff_B_6kHImbUL5_1),.clk(gclk));
	jdff dff_B_1fYz7J8g3_1(.din(w_dff_B_6kHImbUL5_1),.dout(w_dff_B_1fYz7J8g3_1),.clk(gclk));
	jdff dff_B_P2PIbB795_1(.din(w_dff_B_1fYz7J8g3_1),.dout(w_dff_B_P2PIbB795_1),.clk(gclk));
	jdff dff_B_BUerrUPW6_1(.din(w_dff_B_P2PIbB795_1),.dout(w_dff_B_BUerrUPW6_1),.clk(gclk));
	jdff dff_B_IEBvoBpi7_1(.din(w_dff_B_BUerrUPW6_1),.dout(w_dff_B_IEBvoBpi7_1),.clk(gclk));
	jdff dff_B_wqUt48lV2_1(.din(w_dff_B_IEBvoBpi7_1),.dout(w_dff_B_wqUt48lV2_1),.clk(gclk));
	jdff dff_B_vHtlslYq7_1(.din(w_dff_B_wqUt48lV2_1),.dout(w_dff_B_vHtlslYq7_1),.clk(gclk));
	jdff dff_B_6qiNbwWT0_1(.din(w_dff_B_vHtlslYq7_1),.dout(w_dff_B_6qiNbwWT0_1),.clk(gclk));
	jdff dff_B_dro4N5VE5_1(.din(w_dff_B_6qiNbwWT0_1),.dout(w_dff_B_dro4N5VE5_1),.clk(gclk));
	jdff dff_B_4VsBXKE91_1(.din(w_dff_B_dro4N5VE5_1),.dout(w_dff_B_4VsBXKE91_1),.clk(gclk));
	jdff dff_B_Q0I7I8ae0_1(.din(w_dff_B_4VsBXKE91_1),.dout(w_dff_B_Q0I7I8ae0_1),.clk(gclk));
	jdff dff_B_xv0YMTVj1_1(.din(w_dff_B_Q0I7I8ae0_1),.dout(w_dff_B_xv0YMTVj1_1),.clk(gclk));
	jdff dff_B_a1QxwmEr6_1(.din(w_dff_B_xv0YMTVj1_1),.dout(w_dff_B_a1QxwmEr6_1),.clk(gclk));
	jdff dff_B_PrYNMY7t2_1(.din(w_dff_B_a1QxwmEr6_1),.dout(w_dff_B_PrYNMY7t2_1),.clk(gclk));
	jdff dff_B_X7aRTx155_1(.din(w_dff_B_PrYNMY7t2_1),.dout(w_dff_B_X7aRTx155_1),.clk(gclk));
	jdff dff_B_2DeyiiQs4_1(.din(w_dff_B_X7aRTx155_1),.dout(w_dff_B_2DeyiiQs4_1),.clk(gclk));
	jdff dff_B_dYDUkzgO3_1(.din(w_dff_B_2DeyiiQs4_1),.dout(w_dff_B_dYDUkzgO3_1),.clk(gclk));
	jdff dff_B_VQNox5Wu7_1(.din(w_dff_B_dYDUkzgO3_1),.dout(w_dff_B_VQNox5Wu7_1),.clk(gclk));
	jdff dff_B_kik3iT5f1_1(.din(w_dff_B_VQNox5Wu7_1),.dout(w_dff_B_kik3iT5f1_1),.clk(gclk));
	jdff dff_B_qG0HeMm17_1(.din(w_dff_B_kik3iT5f1_1),.dout(w_dff_B_qG0HeMm17_1),.clk(gclk));
	jdff dff_B_0R1rp4Wc2_1(.din(w_dff_B_qG0HeMm17_1),.dout(w_dff_B_0R1rp4Wc2_1),.clk(gclk));
	jdff dff_B_u11I65Fp8_0(.din(n1327),.dout(w_dff_B_u11I65Fp8_0),.clk(gclk));
	jdff dff_B_n0LX8HK47_1(.din(n1842),.dout(w_dff_B_n0LX8HK47_1),.clk(gclk));
	jdff dff_B_6ns2AneW4_1(.din(w_dff_B_n0LX8HK47_1),.dout(w_dff_B_6ns2AneW4_1),.clk(gclk));
	jdff dff_B_1koqxMBQ5_1(.din(w_dff_B_6ns2AneW4_1),.dout(w_dff_B_1koqxMBQ5_1),.clk(gclk));
	jdff dff_B_dFS5DP7C6_1(.din(w_dff_B_1koqxMBQ5_1),.dout(w_dff_B_dFS5DP7C6_1),.clk(gclk));
	jdff dff_B_Z9aypmpx9_1(.din(w_dff_B_dFS5DP7C6_1),.dout(w_dff_B_Z9aypmpx9_1),.clk(gclk));
	jdff dff_B_eH4ngXJK0_1(.din(w_dff_B_Z9aypmpx9_1),.dout(w_dff_B_eH4ngXJK0_1),.clk(gclk));
	jdff dff_B_mk1sOs1A8_1(.din(w_dff_B_eH4ngXJK0_1),.dout(w_dff_B_mk1sOs1A8_1),.clk(gclk));
	jdff dff_B_9Cy1jNDN7_1(.din(w_dff_B_mk1sOs1A8_1),.dout(w_dff_B_9Cy1jNDN7_1),.clk(gclk));
	jdff dff_B_LrXHFHu72_1(.din(w_dff_B_9Cy1jNDN7_1),.dout(w_dff_B_LrXHFHu72_1),.clk(gclk));
	jdff dff_B_iPdCQyZc7_1(.din(w_dff_B_LrXHFHu72_1),.dout(w_dff_B_iPdCQyZc7_1),.clk(gclk));
	jdff dff_B_AOIVlaK13_1(.din(w_dff_B_iPdCQyZc7_1),.dout(w_dff_B_AOIVlaK13_1),.clk(gclk));
	jdff dff_B_fjcqt6UR5_1(.din(w_dff_B_AOIVlaK13_1),.dout(w_dff_B_fjcqt6UR5_1),.clk(gclk));
	jdff dff_B_CRQgdMGd2_1(.din(w_dff_B_fjcqt6UR5_1),.dout(w_dff_B_CRQgdMGd2_1),.clk(gclk));
	jdff dff_B_Bp1dfDng5_0(.din(n1850),.dout(w_dff_B_Bp1dfDng5_0),.clk(gclk));
	jdff dff_B_z1qPUNpM0_0(.din(w_dff_B_Bp1dfDng5_0),.dout(w_dff_B_z1qPUNpM0_0),.clk(gclk));
	jdff dff_B_XCngyXQD0_0(.din(w_dff_B_z1qPUNpM0_0),.dout(w_dff_B_XCngyXQD0_0),.clk(gclk));
	jdff dff_B_fZWO75Y52_0(.din(w_dff_B_XCngyXQD0_0),.dout(w_dff_B_fZWO75Y52_0),.clk(gclk));
	jdff dff_B_ZEjg1Ehh8_0(.din(w_dff_B_fZWO75Y52_0),.dout(w_dff_B_ZEjg1Ehh8_0),.clk(gclk));
	jdff dff_B_JBwtRBqg2_0(.din(w_dff_B_ZEjg1Ehh8_0),.dout(w_dff_B_JBwtRBqg2_0),.clk(gclk));
	jdff dff_B_HrtTerQR4_0(.din(w_dff_B_JBwtRBqg2_0),.dout(w_dff_B_HrtTerQR4_0),.clk(gclk));
	jdff dff_B_dJbWj8eF4_0(.din(w_dff_B_HrtTerQR4_0),.dout(w_dff_B_dJbWj8eF4_0),.clk(gclk));
	jdff dff_B_SbVYbqqq7_0(.din(w_dff_B_dJbWj8eF4_0),.dout(w_dff_B_SbVYbqqq7_0),.clk(gclk));
	jdff dff_B_5mEyW3ZQ4_0(.din(w_dff_B_SbVYbqqq7_0),.dout(w_dff_B_5mEyW3ZQ4_0),.clk(gclk));
	jdff dff_B_3PRkUcnj7_0(.din(w_dff_B_5mEyW3ZQ4_0),.dout(w_dff_B_3PRkUcnj7_0),.clk(gclk));
	jdff dff_A_BJ4y7Wle8_0(.dout(w_n1849_0[0]),.din(w_dff_A_BJ4y7Wle8_0),.clk(gclk));
	jdff dff_A_wh3y0wNg4_0(.dout(w_dff_A_BJ4y7Wle8_0),.din(w_dff_A_wh3y0wNg4_0),.clk(gclk));
	jdff dff_A_rDD0R9Uk3_0(.dout(w_dff_A_wh3y0wNg4_0),.din(w_dff_A_rDD0R9Uk3_0),.clk(gclk));
	jdff dff_A_y2g2Omgw0_0(.dout(w_dff_A_rDD0R9Uk3_0),.din(w_dff_A_y2g2Omgw0_0),.clk(gclk));
	jdff dff_A_dIvK8EgK9_0(.dout(w_dff_A_y2g2Omgw0_0),.din(w_dff_A_dIvK8EgK9_0),.clk(gclk));
	jdff dff_A_OSycrRUc6_0(.dout(w_dff_A_dIvK8EgK9_0),.din(w_dff_A_OSycrRUc6_0),.clk(gclk));
	jdff dff_A_GPXpLpwF7_0(.dout(w_dff_A_OSycrRUc6_0),.din(w_dff_A_GPXpLpwF7_0),.clk(gclk));
	jdff dff_A_d5Ti3UEX0_0(.dout(w_dff_A_GPXpLpwF7_0),.din(w_dff_A_d5Ti3UEX0_0),.clk(gclk));
	jdff dff_A_vhdZGHMM4_0(.dout(w_dff_A_d5Ti3UEX0_0),.din(w_dff_A_vhdZGHMM4_0),.clk(gclk));
	jdff dff_A_vlFk7etE4_0(.dout(w_dff_A_vhdZGHMM4_0),.din(w_dff_A_vlFk7etE4_0),.clk(gclk));
	jdff dff_A_eTZknVkp3_0(.dout(w_dff_A_vlFk7etE4_0),.din(w_dff_A_eTZknVkp3_0),.clk(gclk));
	jdff dff_A_S3oaBWKP4_0(.dout(w_dff_A_eTZknVkp3_0),.din(w_dff_A_S3oaBWKP4_0),.clk(gclk));
	jdff dff_B_koBkdfDe4_1(.din(n1839),.dout(w_dff_B_koBkdfDe4_1),.clk(gclk));
	jdff dff_B_WOnb8SOF2_1(.din(w_dff_B_koBkdfDe4_1),.dout(w_dff_B_WOnb8SOF2_1),.clk(gclk));
	jdff dff_B_nEuXBt0h1_2(.din(n1838),.dout(w_dff_B_nEuXBt0h1_2),.clk(gclk));
	jdff dff_B_JOzWbBhU9_2(.din(w_dff_B_nEuXBt0h1_2),.dout(w_dff_B_JOzWbBhU9_2),.clk(gclk));
	jdff dff_B_fUgv6U4v4_2(.din(w_dff_B_JOzWbBhU9_2),.dout(w_dff_B_fUgv6U4v4_2),.clk(gclk));
	jdff dff_B_tHlkeFko2_2(.din(w_dff_B_fUgv6U4v4_2),.dout(w_dff_B_tHlkeFko2_2),.clk(gclk));
	jdff dff_B_dqBnVESn8_2(.din(w_dff_B_tHlkeFko2_2),.dout(w_dff_B_dqBnVESn8_2),.clk(gclk));
	jdff dff_B_jgzWMh1h8_2(.din(w_dff_B_dqBnVESn8_2),.dout(w_dff_B_jgzWMh1h8_2),.clk(gclk));
	jdff dff_B_9IqJ6khm4_2(.din(w_dff_B_jgzWMh1h8_2),.dout(w_dff_B_9IqJ6khm4_2),.clk(gclk));
	jdff dff_B_JMbEtx3p4_2(.din(w_dff_B_9IqJ6khm4_2),.dout(w_dff_B_JMbEtx3p4_2),.clk(gclk));
	jdff dff_B_F8Kl8dPW8_2(.din(w_dff_B_JMbEtx3p4_2),.dout(w_dff_B_F8Kl8dPW8_2),.clk(gclk));
	jdff dff_B_CVcCcHL35_2(.din(w_dff_B_F8Kl8dPW8_2),.dout(w_dff_B_CVcCcHL35_2),.clk(gclk));
	jdff dff_B_bZEdkymb4_2(.din(w_dff_B_CVcCcHL35_2),.dout(w_dff_B_bZEdkymb4_2),.clk(gclk));
	jdff dff_B_IRnNEqf71_2(.din(w_dff_B_bZEdkymb4_2),.dout(w_dff_B_IRnNEqf71_2),.clk(gclk));
	jdff dff_B_YM5kcdg20_2(.din(w_dff_B_IRnNEqf71_2),.dout(w_dff_B_YM5kcdg20_2),.clk(gclk));
	jdff dff_B_8CZW2qvp4_2(.din(w_dff_B_YM5kcdg20_2),.dout(w_dff_B_8CZW2qvp4_2),.clk(gclk));
	jdff dff_B_sNv1zJeD5_2(.din(w_dff_B_8CZW2qvp4_2),.dout(w_dff_B_sNv1zJeD5_2),.clk(gclk));
	jdff dff_B_k0K2nnHz3_2(.din(w_dff_B_sNv1zJeD5_2),.dout(w_dff_B_k0K2nnHz3_2),.clk(gclk));
	jdff dff_B_rb1w8U7q5_2(.din(w_dff_B_k0K2nnHz3_2),.dout(w_dff_B_rb1w8U7q5_2),.clk(gclk));
	jdff dff_B_sCXdE0Tt4_2(.din(w_dff_B_rb1w8U7q5_2),.dout(w_dff_B_sCXdE0Tt4_2),.clk(gclk));
	jdff dff_B_HBTy6h9n8_2(.din(w_dff_B_sCXdE0Tt4_2),.dout(w_dff_B_HBTy6h9n8_2),.clk(gclk));
	jdff dff_B_jBWqYXq38_2(.din(w_dff_B_HBTy6h9n8_2),.dout(w_dff_B_jBWqYXq38_2),.clk(gclk));
	jdff dff_B_jujs5ISR1_2(.din(w_dff_B_jBWqYXq38_2),.dout(w_dff_B_jujs5ISR1_2),.clk(gclk));
	jdff dff_B_AT4jU38D8_2(.din(w_dff_B_jujs5ISR1_2),.dout(w_dff_B_AT4jU38D8_2),.clk(gclk));
	jdff dff_B_IqqRYEiy4_2(.din(w_dff_B_AT4jU38D8_2),.dout(w_dff_B_IqqRYEiy4_2),.clk(gclk));
	jdff dff_B_2IVRv3ae7_2(.din(w_dff_B_IqqRYEiy4_2),.dout(w_dff_B_2IVRv3ae7_2),.clk(gclk));
	jdff dff_B_JdbAeKTF4_2(.din(w_dff_B_2IVRv3ae7_2),.dout(w_dff_B_JdbAeKTF4_2),.clk(gclk));
	jdff dff_B_NIdbV4B44_2(.din(w_dff_B_JdbAeKTF4_2),.dout(w_dff_B_NIdbV4B44_2),.clk(gclk));
	jdff dff_B_yjSWPEpy6_2(.din(w_dff_B_NIdbV4B44_2),.dout(w_dff_B_yjSWPEpy6_2),.clk(gclk));
	jdff dff_B_N3XxefAG9_2(.din(w_dff_B_yjSWPEpy6_2),.dout(w_dff_B_N3XxefAG9_2),.clk(gclk));
	jdff dff_B_cepbRAYc7_2(.din(w_dff_B_N3XxefAG9_2),.dout(w_dff_B_cepbRAYc7_2),.clk(gclk));
	jdff dff_B_XCfK2yRO3_2(.din(w_dff_B_cepbRAYc7_2),.dout(w_dff_B_XCfK2yRO3_2),.clk(gclk));
	jdff dff_B_8dlMRbOE5_2(.din(w_dff_B_XCfK2yRO3_2),.dout(w_dff_B_8dlMRbOE5_2),.clk(gclk));
	jdff dff_B_hyXwfLLg6_2(.din(w_dff_B_8dlMRbOE5_2),.dout(w_dff_B_hyXwfLLg6_2),.clk(gclk));
	jdff dff_B_hdxH3QjP6_2(.din(w_dff_B_hyXwfLLg6_2),.dout(w_dff_B_hdxH3QjP6_2),.clk(gclk));
	jdff dff_B_xAcshE6C9_2(.din(w_dff_B_hdxH3QjP6_2),.dout(w_dff_B_xAcshE6C9_2),.clk(gclk));
	jdff dff_B_wZIRk25T4_2(.din(w_dff_B_xAcshE6C9_2),.dout(w_dff_B_wZIRk25T4_2),.clk(gclk));
	jdff dff_B_d9ARTDuk8_2(.din(w_dff_B_wZIRk25T4_2),.dout(w_dff_B_d9ARTDuk8_2),.clk(gclk));
	jdff dff_B_tg4T8bQB5_2(.din(w_dff_B_d9ARTDuk8_2),.dout(w_dff_B_tg4T8bQB5_2),.clk(gclk));
	jdff dff_B_MsXe6ssV0_2(.din(w_dff_B_tg4T8bQB5_2),.dout(w_dff_B_MsXe6ssV0_2),.clk(gclk));
	jdff dff_B_z7R67VBi6_2(.din(w_dff_B_MsXe6ssV0_2),.dout(w_dff_B_z7R67VBi6_2),.clk(gclk));
	jdff dff_B_I48V4YaI3_2(.din(w_dff_B_z7R67VBi6_2),.dout(w_dff_B_I48V4YaI3_2),.clk(gclk));
	jdff dff_B_nhlUiY0X9_2(.din(w_dff_B_I48V4YaI3_2),.dout(w_dff_B_nhlUiY0X9_2),.clk(gclk));
	jdff dff_B_UCUluUy38_2(.din(w_dff_B_nhlUiY0X9_2),.dout(w_dff_B_UCUluUy38_2),.clk(gclk));
	jdff dff_B_6tHIm0Zj1_2(.din(w_dff_B_UCUluUy38_2),.dout(w_dff_B_6tHIm0Zj1_2),.clk(gclk));
	jdff dff_B_fDrxW39B4_2(.din(w_dff_B_6tHIm0Zj1_2),.dout(w_dff_B_fDrxW39B4_2),.clk(gclk));
	jdff dff_B_zUhDUf382_2(.din(w_dff_B_fDrxW39B4_2),.dout(w_dff_B_zUhDUf382_2),.clk(gclk));
	jdff dff_B_hdtmYOMd1_2(.din(w_dff_B_zUhDUf382_2),.dout(w_dff_B_hdtmYOMd1_2),.clk(gclk));
	jdff dff_B_HHIV3MQM1_2(.din(w_dff_B_hdtmYOMd1_2),.dout(w_dff_B_HHIV3MQM1_2),.clk(gclk));
	jdff dff_B_LRdvF6EQ6_2(.din(w_dff_B_HHIV3MQM1_2),.dout(w_dff_B_LRdvF6EQ6_2),.clk(gclk));
	jdff dff_B_CVZWGe6c4_2(.din(w_dff_B_LRdvF6EQ6_2),.dout(w_dff_B_CVZWGe6c4_2),.clk(gclk));
	jdff dff_B_x8EtMWeH1_2(.din(w_dff_B_CVZWGe6c4_2),.dout(w_dff_B_x8EtMWeH1_2),.clk(gclk));
	jdff dff_B_oaMw4zbH6_2(.din(w_dff_B_x8EtMWeH1_2),.dout(w_dff_B_oaMw4zbH6_2),.clk(gclk));
	jdff dff_B_hWBi9QTS3_2(.din(w_dff_B_oaMw4zbH6_2),.dout(w_dff_B_hWBi9QTS3_2),.clk(gclk));
	jdff dff_B_MsJNs49r5_2(.din(w_dff_B_hWBi9QTS3_2),.dout(w_dff_B_MsJNs49r5_2),.clk(gclk));
	jdff dff_B_tB4TPbVH7_2(.din(w_dff_B_MsJNs49r5_2),.dout(w_dff_B_tB4TPbVH7_2),.clk(gclk));
	jdff dff_B_rZzduNnC5_2(.din(w_dff_B_tB4TPbVH7_2),.dout(w_dff_B_rZzduNnC5_2),.clk(gclk));
	jdff dff_B_lv8uBgJO8_2(.din(w_dff_B_rZzduNnC5_2),.dout(w_dff_B_lv8uBgJO8_2),.clk(gclk));
	jdff dff_B_VapzC66b9_2(.din(w_dff_B_lv8uBgJO8_2),.dout(w_dff_B_VapzC66b9_2),.clk(gclk));
	jdff dff_B_JoxeLlV34_2(.din(w_dff_B_VapzC66b9_2),.dout(w_dff_B_JoxeLlV34_2),.clk(gclk));
	jdff dff_B_Z8eS5z1F6_2(.din(w_dff_B_JoxeLlV34_2),.dout(w_dff_B_Z8eS5z1F6_2),.clk(gclk));
	jdff dff_B_ePcqAiRz6_2(.din(w_dff_B_Z8eS5z1F6_2),.dout(w_dff_B_ePcqAiRz6_2),.clk(gclk));
	jdff dff_B_JnwV1ZWt8_1(.din(n1845),.dout(w_dff_B_JnwV1ZWt8_1),.clk(gclk));
	jdff dff_B_qXSxj49q2_1(.din(w_dff_B_JnwV1ZWt8_1),.dout(w_dff_B_qXSxj49q2_1),.clk(gclk));
	jdff dff_B_5CsEPWPS6_1(.din(w_dff_B_qXSxj49q2_1),.dout(w_dff_B_5CsEPWPS6_1),.clk(gclk));
	jdff dff_B_GW4GZKY47_1(.din(w_dff_B_5CsEPWPS6_1),.dout(w_dff_B_GW4GZKY47_1),.clk(gclk));
	jdff dff_B_xEw3p8Zd7_1(.din(w_dff_B_GW4GZKY47_1),.dout(w_dff_B_xEw3p8Zd7_1),.clk(gclk));
	jdff dff_B_qOxhTNHt7_1(.din(w_dff_B_xEw3p8Zd7_1),.dout(w_dff_B_qOxhTNHt7_1),.clk(gclk));
	jdff dff_B_0JORbhdS1_1(.din(w_dff_B_qOxhTNHt7_1),.dout(w_dff_B_0JORbhdS1_1),.clk(gclk));
	jdff dff_B_LM8C4jpA7_1(.din(w_dff_B_0JORbhdS1_1),.dout(w_dff_B_LM8C4jpA7_1),.clk(gclk));
	jdff dff_B_Ehttn7093_1(.din(w_dff_B_LM8C4jpA7_1),.dout(w_dff_B_Ehttn7093_1),.clk(gclk));
	jdff dff_B_H66ywrZl3_1(.din(w_dff_B_Ehttn7093_1),.dout(w_dff_B_H66ywrZl3_1),.clk(gclk));
	jdff dff_B_9BjyQurF6_1(.din(w_dff_B_H66ywrZl3_1),.dout(w_dff_B_9BjyQurF6_1),.clk(gclk));
	jdff dff_B_PYOtlqJO2_0(.din(n1846),.dout(w_dff_B_PYOtlqJO2_0),.clk(gclk));
	jdff dff_B_vWoNWi672_0(.din(w_dff_B_PYOtlqJO2_0),.dout(w_dff_B_vWoNWi672_0),.clk(gclk));
	jdff dff_B_Yp3G70995_0(.din(w_dff_B_vWoNWi672_0),.dout(w_dff_B_Yp3G70995_0),.clk(gclk));
	jdff dff_B_aYeKkPR34_0(.din(w_dff_B_Yp3G70995_0),.dout(w_dff_B_aYeKkPR34_0),.clk(gclk));
	jdff dff_B_8amJfuLy1_0(.din(w_dff_B_aYeKkPR34_0),.dout(w_dff_B_8amJfuLy1_0),.clk(gclk));
	jdff dff_B_Pk2uFOrX4_0(.din(w_dff_B_8amJfuLy1_0),.dout(w_dff_B_Pk2uFOrX4_0),.clk(gclk));
	jdff dff_B_OLgVuWOW8_0(.din(w_dff_B_Pk2uFOrX4_0),.dout(w_dff_B_OLgVuWOW8_0),.clk(gclk));
	jdff dff_B_WYbEhz6C4_0(.din(w_dff_B_OLgVuWOW8_0),.dout(w_dff_B_WYbEhz6C4_0),.clk(gclk));
	jdff dff_B_fxyJUvnQ9_0(.din(w_dff_B_WYbEhz6C4_0),.dout(w_dff_B_fxyJUvnQ9_0),.clk(gclk));
	jdff dff_B_qFQVdwG56_0(.din(w_dff_B_fxyJUvnQ9_0),.dout(w_dff_B_qFQVdwG56_0),.clk(gclk));
	jdff dff_A_nk87A8Dq2_1(.dout(w_n1836_0[1]),.din(w_dff_A_nk87A8Dq2_1),.clk(gclk));
	jdff dff_A_Mcdi5QNK0_1(.dout(w_dff_A_nk87A8Dq2_1),.din(w_dff_A_Mcdi5QNK0_1),.clk(gclk));
	jdff dff_A_ghVWx5al9_1(.dout(w_dff_A_Mcdi5QNK0_1),.din(w_dff_A_ghVWx5al9_1),.clk(gclk));
	jdff dff_A_f6FrMDOM6_1(.dout(w_dff_A_ghVWx5al9_1),.din(w_dff_A_f6FrMDOM6_1),.clk(gclk));
	jdff dff_A_akaDuShF5_1(.dout(w_dff_A_f6FrMDOM6_1),.din(w_dff_A_akaDuShF5_1),.clk(gclk));
	jdff dff_A_cFeDyn1d0_1(.dout(w_dff_A_akaDuShF5_1),.din(w_dff_A_cFeDyn1d0_1),.clk(gclk));
	jdff dff_A_WoOF1ovi5_1(.dout(w_dff_A_cFeDyn1d0_1),.din(w_dff_A_WoOF1ovi5_1),.clk(gclk));
	jdff dff_A_A7m0i16D3_1(.dout(w_dff_A_WoOF1ovi5_1),.din(w_dff_A_A7m0i16D3_1),.clk(gclk));
	jdff dff_A_X8l1TA9i6_1(.dout(w_dff_A_A7m0i16D3_1),.din(w_dff_A_X8l1TA9i6_1),.clk(gclk));
	jdff dff_A_75M4gMx63_1(.dout(w_dff_A_X8l1TA9i6_1),.din(w_dff_A_75M4gMx63_1),.clk(gclk));
	jdff dff_A_zIOHEaBV8_1(.dout(w_dff_A_75M4gMx63_1),.din(w_dff_A_zIOHEaBV8_1),.clk(gclk));
	jdff dff_B_YpfZXQss1_1(.din(n1821),.dout(w_dff_B_YpfZXQss1_1),.clk(gclk));
	jdff dff_B_ax82Dsdr0_1(.din(w_dff_B_YpfZXQss1_1),.dout(w_dff_B_ax82Dsdr0_1),.clk(gclk));
	jdff dff_B_cm0kPttC7_1(.din(w_dff_B_ax82Dsdr0_1),.dout(w_dff_B_cm0kPttC7_1),.clk(gclk));
	jdff dff_B_XE2IO5qy3_1(.din(w_dff_B_cm0kPttC7_1),.dout(w_dff_B_XE2IO5qy3_1),.clk(gclk));
	jdff dff_B_OuOoZMZN4_1(.din(w_dff_B_XE2IO5qy3_1),.dout(w_dff_B_OuOoZMZN4_1),.clk(gclk));
	jdff dff_B_nnBCEnVs7_1(.din(w_dff_B_OuOoZMZN4_1),.dout(w_dff_B_nnBCEnVs7_1),.clk(gclk));
	jdff dff_B_6pROSCHP8_1(.din(w_dff_B_nnBCEnVs7_1),.dout(w_dff_B_6pROSCHP8_1),.clk(gclk));
	jdff dff_B_2SBE1Oq47_1(.din(w_dff_B_6pROSCHP8_1),.dout(w_dff_B_2SBE1Oq47_1),.clk(gclk));
	jdff dff_B_ehtuY3Tn8_1(.din(w_dff_B_2SBE1Oq47_1),.dout(w_dff_B_ehtuY3Tn8_1),.clk(gclk));
	jdff dff_B_Gp4NQj3s2_1(.din(w_dff_B_ehtuY3Tn8_1),.dout(w_dff_B_Gp4NQj3s2_1),.clk(gclk));
	jdff dff_B_NQTZLS0q4_1(.din(w_dff_B_Gp4NQj3s2_1),.dout(w_dff_B_NQTZLS0q4_1),.clk(gclk));
	jdff dff_B_4jBcN43r6_0(.din(n1822),.dout(w_dff_B_4jBcN43r6_0),.clk(gclk));
	jdff dff_B_CGkeXy6N7_0(.din(w_dff_B_4jBcN43r6_0),.dout(w_dff_B_CGkeXy6N7_0),.clk(gclk));
	jdff dff_B_o3HO7RTu9_0(.din(w_dff_B_CGkeXy6N7_0),.dout(w_dff_B_o3HO7RTu9_0),.clk(gclk));
	jdff dff_B_Y1CNqHxN0_0(.din(w_dff_B_o3HO7RTu9_0),.dout(w_dff_B_Y1CNqHxN0_0),.clk(gclk));
	jdff dff_B_C4VeJW8r2_0(.din(w_dff_B_Y1CNqHxN0_0),.dout(w_dff_B_C4VeJW8r2_0),.clk(gclk));
	jdff dff_B_1CAcnE9l7_0(.din(w_dff_B_C4VeJW8r2_0),.dout(w_dff_B_1CAcnE9l7_0),.clk(gclk));
	jdff dff_B_vqAhaM5b6_0(.din(w_dff_B_1CAcnE9l7_0),.dout(w_dff_B_vqAhaM5b6_0),.clk(gclk));
	jdff dff_B_nGS1uDC61_0(.din(w_dff_B_vqAhaM5b6_0),.dout(w_dff_B_nGS1uDC61_0),.clk(gclk));
	jdff dff_B_5sbpvJjw0_0(.din(w_dff_B_nGS1uDC61_0),.dout(w_dff_B_5sbpvJjw0_0),.clk(gclk));
	jdff dff_B_EHataNLT3_0(.din(w_dff_B_5sbpvJjw0_0),.dout(w_dff_B_EHataNLT3_0),.clk(gclk));
	jdff dff_A_QE8AgDb75_1(.dout(w_n1817_0[1]),.din(w_dff_A_QE8AgDb75_1),.clk(gclk));
	jdff dff_A_0mUsjU6w3_1(.dout(w_dff_A_QE8AgDb75_1),.din(w_dff_A_0mUsjU6w3_1),.clk(gclk));
	jdff dff_A_aF4XfnDL2_1(.dout(w_dff_A_0mUsjU6w3_1),.din(w_dff_A_aF4XfnDL2_1),.clk(gclk));
	jdff dff_A_gbt5IOib1_1(.dout(w_dff_A_aF4XfnDL2_1),.din(w_dff_A_gbt5IOib1_1),.clk(gclk));
	jdff dff_A_1oH8ZtIp1_1(.dout(w_dff_A_gbt5IOib1_1),.din(w_dff_A_1oH8ZtIp1_1),.clk(gclk));
	jdff dff_A_TBAGzUVs1_1(.dout(w_dff_A_1oH8ZtIp1_1),.din(w_dff_A_TBAGzUVs1_1),.clk(gclk));
	jdff dff_A_FuYVuRKB3_1(.dout(w_dff_A_TBAGzUVs1_1),.din(w_dff_A_FuYVuRKB3_1),.clk(gclk));
	jdff dff_A_ncEp9u7e5_1(.dout(w_dff_A_FuYVuRKB3_1),.din(w_dff_A_ncEp9u7e5_1),.clk(gclk));
	jdff dff_A_XSva6HVo6_1(.dout(w_dff_A_ncEp9u7e5_1),.din(w_dff_A_XSva6HVo6_1),.clk(gclk));
	jdff dff_A_lOHNcVEa5_1(.dout(w_dff_A_XSva6HVo6_1),.din(w_dff_A_lOHNcVEa5_1),.clk(gclk));
	jdff dff_A_2B9FjQxb3_1(.dout(w_dff_A_lOHNcVEa5_1),.din(w_dff_A_2B9FjQxb3_1),.clk(gclk));
	jdff dff_B_i52lIxVR4_1(.din(n1795),.dout(w_dff_B_i52lIxVR4_1),.clk(gclk));
	jdff dff_B_Dr5ldv727_1(.din(w_dff_B_i52lIxVR4_1),.dout(w_dff_B_Dr5ldv727_1),.clk(gclk));
	jdff dff_B_lhzLMJYF4_1(.din(w_dff_B_Dr5ldv727_1),.dout(w_dff_B_lhzLMJYF4_1),.clk(gclk));
	jdff dff_B_xbZ3ChDl6_1(.din(w_dff_B_lhzLMJYF4_1),.dout(w_dff_B_xbZ3ChDl6_1),.clk(gclk));
	jdff dff_B_FhL4hDBK2_1(.din(w_dff_B_xbZ3ChDl6_1),.dout(w_dff_B_FhL4hDBK2_1),.clk(gclk));
	jdff dff_B_48HKwAtk5_1(.din(w_dff_B_FhL4hDBK2_1),.dout(w_dff_B_48HKwAtk5_1),.clk(gclk));
	jdff dff_B_jSK22BhL5_1(.din(w_dff_B_48HKwAtk5_1),.dout(w_dff_B_jSK22BhL5_1),.clk(gclk));
	jdff dff_B_P5IiImCZ2_1(.din(w_dff_B_jSK22BhL5_1),.dout(w_dff_B_P5IiImCZ2_1),.clk(gclk));
	jdff dff_B_zAkpJhzv9_1(.din(w_dff_B_P5IiImCZ2_1),.dout(w_dff_B_zAkpJhzv9_1),.clk(gclk));
	jdff dff_B_An3zfZ9k7_1(.din(w_dff_B_zAkpJhzv9_1),.dout(w_dff_B_An3zfZ9k7_1),.clk(gclk));
	jdff dff_B_fdbJkxX72_1(.din(w_dff_B_An3zfZ9k7_1),.dout(w_dff_B_fdbJkxX72_1),.clk(gclk));
	jdff dff_B_EiUK8CGZ9_0(.din(n1796),.dout(w_dff_B_EiUK8CGZ9_0),.clk(gclk));
	jdff dff_B_AytBTrla6_0(.din(w_dff_B_EiUK8CGZ9_0),.dout(w_dff_B_AytBTrla6_0),.clk(gclk));
	jdff dff_B_HU5yLeRN6_0(.din(w_dff_B_AytBTrla6_0),.dout(w_dff_B_HU5yLeRN6_0),.clk(gclk));
	jdff dff_B_lFt0TUh56_0(.din(w_dff_B_HU5yLeRN6_0),.dout(w_dff_B_lFt0TUh56_0),.clk(gclk));
	jdff dff_B_VhFZKmrQ3_0(.din(w_dff_B_lFt0TUh56_0),.dout(w_dff_B_VhFZKmrQ3_0),.clk(gclk));
	jdff dff_B_8uuVBiwE2_0(.din(w_dff_B_VhFZKmrQ3_0),.dout(w_dff_B_8uuVBiwE2_0),.clk(gclk));
	jdff dff_B_PWajHzqd0_0(.din(w_dff_B_8uuVBiwE2_0),.dout(w_dff_B_PWajHzqd0_0),.clk(gclk));
	jdff dff_B_Lcsf8UQD7_0(.din(w_dff_B_PWajHzqd0_0),.dout(w_dff_B_Lcsf8UQD7_0),.clk(gclk));
	jdff dff_B_U0J3qJw59_0(.din(w_dff_B_Lcsf8UQD7_0),.dout(w_dff_B_U0J3qJw59_0),.clk(gclk));
	jdff dff_B_tvgH6RWW3_0(.din(w_dff_B_U0J3qJw59_0),.dout(w_dff_B_tvgH6RWW3_0),.clk(gclk));
	jdff dff_A_G0CghVSE2_1(.dout(w_n1791_0[1]),.din(w_dff_A_G0CghVSE2_1),.clk(gclk));
	jdff dff_A_mXmWR6iq6_1(.dout(w_dff_A_G0CghVSE2_1),.din(w_dff_A_mXmWR6iq6_1),.clk(gclk));
	jdff dff_A_eATnJKXS0_1(.dout(w_dff_A_mXmWR6iq6_1),.din(w_dff_A_eATnJKXS0_1),.clk(gclk));
	jdff dff_A_5amLb5yT3_1(.dout(w_dff_A_eATnJKXS0_1),.din(w_dff_A_5amLb5yT3_1),.clk(gclk));
	jdff dff_A_geN1YJdJ8_1(.dout(w_dff_A_5amLb5yT3_1),.din(w_dff_A_geN1YJdJ8_1),.clk(gclk));
	jdff dff_A_NcAAZBOy2_1(.dout(w_dff_A_geN1YJdJ8_1),.din(w_dff_A_NcAAZBOy2_1),.clk(gclk));
	jdff dff_A_zCvsgT2n8_1(.dout(w_dff_A_NcAAZBOy2_1),.din(w_dff_A_zCvsgT2n8_1),.clk(gclk));
	jdff dff_A_xaus8U144_1(.dout(w_dff_A_zCvsgT2n8_1),.din(w_dff_A_xaus8U144_1),.clk(gclk));
	jdff dff_A_Fs5VNS545_1(.dout(w_dff_A_xaus8U144_1),.din(w_dff_A_Fs5VNS545_1),.clk(gclk));
	jdff dff_A_5J14Okyl9_1(.dout(w_dff_A_Fs5VNS545_1),.din(w_dff_A_5J14Okyl9_1),.clk(gclk));
	jdff dff_A_xi9bByvv3_1(.dout(w_dff_A_5J14Okyl9_1),.din(w_dff_A_xi9bByvv3_1),.clk(gclk));
	jdff dff_B_apthHD0e7_1(.din(n1762),.dout(w_dff_B_apthHD0e7_1),.clk(gclk));
	jdff dff_B_3CNzG3aN4_1(.din(w_dff_B_apthHD0e7_1),.dout(w_dff_B_3CNzG3aN4_1),.clk(gclk));
	jdff dff_B_PzWddbZx0_1(.din(w_dff_B_3CNzG3aN4_1),.dout(w_dff_B_PzWddbZx0_1),.clk(gclk));
	jdff dff_B_CITiLbRG3_1(.din(w_dff_B_PzWddbZx0_1),.dout(w_dff_B_CITiLbRG3_1),.clk(gclk));
	jdff dff_B_NmzAodJC2_1(.din(w_dff_B_CITiLbRG3_1),.dout(w_dff_B_NmzAodJC2_1),.clk(gclk));
	jdff dff_B_XNOh7ZWf3_1(.din(w_dff_B_NmzAodJC2_1),.dout(w_dff_B_XNOh7ZWf3_1),.clk(gclk));
	jdff dff_B_1LpawFoo9_1(.din(w_dff_B_XNOh7ZWf3_1),.dout(w_dff_B_1LpawFoo9_1),.clk(gclk));
	jdff dff_B_6YCGpQLP2_1(.din(w_dff_B_1LpawFoo9_1),.dout(w_dff_B_6YCGpQLP2_1),.clk(gclk));
	jdff dff_B_Ohoibt1s9_1(.din(w_dff_B_6YCGpQLP2_1),.dout(w_dff_B_Ohoibt1s9_1),.clk(gclk));
	jdff dff_B_MvQb0VFd2_1(.din(w_dff_B_Ohoibt1s9_1),.dout(w_dff_B_MvQb0VFd2_1),.clk(gclk));
	jdff dff_B_yegT27uo2_1(.din(w_dff_B_MvQb0VFd2_1),.dout(w_dff_B_yegT27uo2_1),.clk(gclk));
	jdff dff_B_64NhoyK05_0(.din(n1763),.dout(w_dff_B_64NhoyK05_0),.clk(gclk));
	jdff dff_B_d3hNrJBK0_0(.din(w_dff_B_64NhoyK05_0),.dout(w_dff_B_d3hNrJBK0_0),.clk(gclk));
	jdff dff_B_DrIMhhQN8_0(.din(w_dff_B_d3hNrJBK0_0),.dout(w_dff_B_DrIMhhQN8_0),.clk(gclk));
	jdff dff_B_vfYykq8t3_0(.din(w_dff_B_DrIMhhQN8_0),.dout(w_dff_B_vfYykq8t3_0),.clk(gclk));
	jdff dff_B_mj6D7phu8_0(.din(w_dff_B_vfYykq8t3_0),.dout(w_dff_B_mj6D7phu8_0),.clk(gclk));
	jdff dff_B_2eSu4Mxe3_0(.din(w_dff_B_mj6D7phu8_0),.dout(w_dff_B_2eSu4Mxe3_0),.clk(gclk));
	jdff dff_B_tfxb9vAU6_0(.din(w_dff_B_2eSu4Mxe3_0),.dout(w_dff_B_tfxb9vAU6_0),.clk(gclk));
	jdff dff_B_2tc02Oid4_0(.din(w_dff_B_tfxb9vAU6_0),.dout(w_dff_B_2tc02Oid4_0),.clk(gclk));
	jdff dff_B_1UsXatsV3_0(.din(w_dff_B_2tc02Oid4_0),.dout(w_dff_B_1UsXatsV3_0),.clk(gclk));
	jdff dff_B_3nD9Myey6_0(.din(w_dff_B_1UsXatsV3_0),.dout(w_dff_B_3nD9Myey6_0),.clk(gclk));
	jdff dff_A_9mQsSc2g5_1(.dout(w_n1758_0[1]),.din(w_dff_A_9mQsSc2g5_1),.clk(gclk));
	jdff dff_A_Sjtr7ByO3_1(.dout(w_dff_A_9mQsSc2g5_1),.din(w_dff_A_Sjtr7ByO3_1),.clk(gclk));
	jdff dff_A_IcP6V3Gg1_1(.dout(w_dff_A_Sjtr7ByO3_1),.din(w_dff_A_IcP6V3Gg1_1),.clk(gclk));
	jdff dff_A_6pYpxFGI2_1(.dout(w_dff_A_IcP6V3Gg1_1),.din(w_dff_A_6pYpxFGI2_1),.clk(gclk));
	jdff dff_A_qTjsp5wm9_1(.dout(w_dff_A_6pYpxFGI2_1),.din(w_dff_A_qTjsp5wm9_1),.clk(gclk));
	jdff dff_A_vjUs6s9b9_1(.dout(w_dff_A_qTjsp5wm9_1),.din(w_dff_A_vjUs6s9b9_1),.clk(gclk));
	jdff dff_A_C7Mk18sD1_1(.dout(w_dff_A_vjUs6s9b9_1),.din(w_dff_A_C7Mk18sD1_1),.clk(gclk));
	jdff dff_A_fAbhAN8Z0_1(.dout(w_dff_A_C7Mk18sD1_1),.din(w_dff_A_fAbhAN8Z0_1),.clk(gclk));
	jdff dff_A_oP21dmZr9_1(.dout(w_dff_A_fAbhAN8Z0_1),.din(w_dff_A_oP21dmZr9_1),.clk(gclk));
	jdff dff_A_KjjI57cC0_1(.dout(w_dff_A_oP21dmZr9_1),.din(w_dff_A_KjjI57cC0_1),.clk(gclk));
	jdff dff_A_E6PWdTsO3_1(.dout(w_dff_A_KjjI57cC0_1),.din(w_dff_A_E6PWdTsO3_1),.clk(gclk));
	jdff dff_B_lH4AGOPK9_1(.din(n1722),.dout(w_dff_B_lH4AGOPK9_1),.clk(gclk));
	jdff dff_B_pZCIYfz65_1(.din(w_dff_B_lH4AGOPK9_1),.dout(w_dff_B_pZCIYfz65_1),.clk(gclk));
	jdff dff_B_aN1T8Bvq5_1(.din(w_dff_B_pZCIYfz65_1),.dout(w_dff_B_aN1T8Bvq5_1),.clk(gclk));
	jdff dff_B_drALFYzw0_1(.din(w_dff_B_aN1T8Bvq5_1),.dout(w_dff_B_drALFYzw0_1),.clk(gclk));
	jdff dff_B_mqANwPTm8_1(.din(w_dff_B_drALFYzw0_1),.dout(w_dff_B_mqANwPTm8_1),.clk(gclk));
	jdff dff_B_bzga3F7h5_1(.din(w_dff_B_mqANwPTm8_1),.dout(w_dff_B_bzga3F7h5_1),.clk(gclk));
	jdff dff_B_tmtsrMiO3_1(.din(w_dff_B_bzga3F7h5_1),.dout(w_dff_B_tmtsrMiO3_1),.clk(gclk));
	jdff dff_B_JrbHG7JQ6_1(.din(w_dff_B_tmtsrMiO3_1),.dout(w_dff_B_JrbHG7JQ6_1),.clk(gclk));
	jdff dff_B_D8UuVnSp3_1(.din(w_dff_B_JrbHG7JQ6_1),.dout(w_dff_B_D8UuVnSp3_1),.clk(gclk));
	jdff dff_B_BIWYyO460_1(.din(w_dff_B_D8UuVnSp3_1),.dout(w_dff_B_BIWYyO460_1),.clk(gclk));
	jdff dff_B_Wq2Kv3s35_1(.din(w_dff_B_BIWYyO460_1),.dout(w_dff_B_Wq2Kv3s35_1),.clk(gclk));
	jdff dff_B_rScQOwiB1_0(.din(n1723),.dout(w_dff_B_rScQOwiB1_0),.clk(gclk));
	jdff dff_B_wggJHljV9_0(.din(w_dff_B_rScQOwiB1_0),.dout(w_dff_B_wggJHljV9_0),.clk(gclk));
	jdff dff_B_a9eyFLI59_0(.din(w_dff_B_wggJHljV9_0),.dout(w_dff_B_a9eyFLI59_0),.clk(gclk));
	jdff dff_B_6mFfBnNw7_0(.din(w_dff_B_a9eyFLI59_0),.dout(w_dff_B_6mFfBnNw7_0),.clk(gclk));
	jdff dff_B_ZNYORSge3_0(.din(w_dff_B_6mFfBnNw7_0),.dout(w_dff_B_ZNYORSge3_0),.clk(gclk));
	jdff dff_B_50Jg3p789_0(.din(w_dff_B_ZNYORSge3_0),.dout(w_dff_B_50Jg3p789_0),.clk(gclk));
	jdff dff_B_JD6PozWB6_0(.din(w_dff_B_50Jg3p789_0),.dout(w_dff_B_JD6PozWB6_0),.clk(gclk));
	jdff dff_B_yb3ddDnU1_0(.din(w_dff_B_JD6PozWB6_0),.dout(w_dff_B_yb3ddDnU1_0),.clk(gclk));
	jdff dff_B_apjOOWYS0_0(.din(w_dff_B_yb3ddDnU1_0),.dout(w_dff_B_apjOOWYS0_0),.clk(gclk));
	jdff dff_A_ZBUv3hRO5_1(.dout(w_n1720_0[1]),.din(w_dff_A_ZBUv3hRO5_1),.clk(gclk));
	jdff dff_A_fnYVZVd12_1(.dout(w_dff_A_ZBUv3hRO5_1),.din(w_dff_A_fnYVZVd12_1),.clk(gclk));
	jdff dff_A_CMyBLQ227_1(.dout(w_dff_A_fnYVZVd12_1),.din(w_dff_A_CMyBLQ227_1),.clk(gclk));
	jdff dff_A_3qhdM4hb1_1(.dout(w_dff_A_CMyBLQ227_1),.din(w_dff_A_3qhdM4hb1_1),.clk(gclk));
	jdff dff_A_fKZfkly18_1(.dout(w_dff_A_3qhdM4hb1_1),.din(w_dff_A_fKZfkly18_1),.clk(gclk));
	jdff dff_A_sUQCH0aM0_1(.dout(w_dff_A_fKZfkly18_1),.din(w_dff_A_sUQCH0aM0_1),.clk(gclk));
	jdff dff_A_jWvFyAXy9_1(.dout(w_dff_A_sUQCH0aM0_1),.din(w_dff_A_jWvFyAXy9_1),.clk(gclk));
	jdff dff_A_9fOCJ18c2_1(.dout(w_dff_A_jWvFyAXy9_1),.din(w_dff_A_9fOCJ18c2_1),.clk(gclk));
	jdff dff_A_qbZioxW05_1(.dout(w_dff_A_9fOCJ18c2_1),.din(w_dff_A_qbZioxW05_1),.clk(gclk));
	jdff dff_A_HV3sCXwW3_1(.dout(w_dff_A_qbZioxW05_1),.din(w_dff_A_HV3sCXwW3_1),.clk(gclk));
	jdff dff_B_QrDZuXk75_1(.din(n1674),.dout(w_dff_B_QrDZuXk75_1),.clk(gclk));
	jdff dff_B_8U7dz88v0_1(.din(w_dff_B_QrDZuXk75_1),.dout(w_dff_B_8U7dz88v0_1),.clk(gclk));
	jdff dff_B_4eQubw3Y2_1(.din(w_dff_B_8U7dz88v0_1),.dout(w_dff_B_4eQubw3Y2_1),.clk(gclk));
	jdff dff_B_EyYA1Y8n3_1(.din(w_dff_B_4eQubw3Y2_1),.dout(w_dff_B_EyYA1Y8n3_1),.clk(gclk));
	jdff dff_B_vpjXqzBJ5_1(.din(w_dff_B_EyYA1Y8n3_1),.dout(w_dff_B_vpjXqzBJ5_1),.clk(gclk));
	jdff dff_B_v4zOHPYL9_1(.din(w_dff_B_vpjXqzBJ5_1),.dout(w_dff_B_v4zOHPYL9_1),.clk(gclk));
	jdff dff_B_tGZy8yPl4_1(.din(w_dff_B_v4zOHPYL9_1),.dout(w_dff_B_tGZy8yPl4_1),.clk(gclk));
	jdff dff_B_ih7J4Yym1_1(.din(w_dff_B_tGZy8yPl4_1),.dout(w_dff_B_ih7J4Yym1_1),.clk(gclk));
	jdff dff_B_iHJZqq0E4_1(.din(w_dff_B_ih7J4Yym1_1),.dout(w_dff_B_iHJZqq0E4_1),.clk(gclk));
	jdff dff_B_Hczv6KUZ7_1(.din(w_dff_B_iHJZqq0E4_1),.dout(w_dff_B_Hczv6KUZ7_1),.clk(gclk));
	jdff dff_B_60htQl7F3_0(.din(n1675),.dout(w_dff_B_60htQl7F3_0),.clk(gclk));
	jdff dff_B_44xPq9ta6_0(.din(w_dff_B_60htQl7F3_0),.dout(w_dff_B_44xPq9ta6_0),.clk(gclk));
	jdff dff_B_BZYUnd6j5_0(.din(w_dff_B_44xPq9ta6_0),.dout(w_dff_B_BZYUnd6j5_0),.clk(gclk));
	jdff dff_B_ymnNBS8V3_0(.din(w_dff_B_BZYUnd6j5_0),.dout(w_dff_B_ymnNBS8V3_0),.clk(gclk));
	jdff dff_B_aCjEXt151_0(.din(w_dff_B_ymnNBS8V3_0),.dout(w_dff_B_aCjEXt151_0),.clk(gclk));
	jdff dff_B_vCJ1xMxt7_0(.din(w_dff_B_aCjEXt151_0),.dout(w_dff_B_vCJ1xMxt7_0),.clk(gclk));
	jdff dff_B_pkYusNoI1_0(.din(w_dff_B_vCJ1xMxt7_0),.dout(w_dff_B_pkYusNoI1_0),.clk(gclk));
	jdff dff_B_a4Snyv5j7_0(.din(w_dff_B_pkYusNoI1_0),.dout(w_dff_B_a4Snyv5j7_0),.clk(gclk));
	jdff dff_A_kte2a3xO4_1(.dout(w_n1672_0[1]),.din(w_dff_A_kte2a3xO4_1),.clk(gclk));
	jdff dff_A_sJigHy9A3_1(.dout(w_dff_A_kte2a3xO4_1),.din(w_dff_A_sJigHy9A3_1),.clk(gclk));
	jdff dff_A_c8gRWP3l6_1(.dout(w_dff_A_sJigHy9A3_1),.din(w_dff_A_c8gRWP3l6_1),.clk(gclk));
	jdff dff_A_WtoWpsNH6_1(.dout(w_dff_A_c8gRWP3l6_1),.din(w_dff_A_WtoWpsNH6_1),.clk(gclk));
	jdff dff_A_W4V3Bqox1_1(.dout(w_dff_A_WtoWpsNH6_1),.din(w_dff_A_W4V3Bqox1_1),.clk(gclk));
	jdff dff_A_4qbFL7Py8_1(.dout(w_dff_A_W4V3Bqox1_1),.din(w_dff_A_4qbFL7Py8_1),.clk(gclk));
	jdff dff_A_8jqlQjjl5_1(.dout(w_dff_A_4qbFL7Py8_1),.din(w_dff_A_8jqlQjjl5_1),.clk(gclk));
	jdff dff_A_rwhWemd01_1(.dout(w_dff_A_8jqlQjjl5_1),.din(w_dff_A_rwhWemd01_1),.clk(gclk));
	jdff dff_A_7o8BL2rh8_1(.dout(w_dff_A_rwhWemd01_1),.din(w_dff_A_7o8BL2rh8_1),.clk(gclk));
	jdff dff_B_WyKDqC1u0_1(.din(n1619),.dout(w_dff_B_WyKDqC1u0_1),.clk(gclk));
	jdff dff_B_DSabBSQw0_1(.din(w_dff_B_WyKDqC1u0_1),.dout(w_dff_B_DSabBSQw0_1),.clk(gclk));
	jdff dff_B_wYbgBOcU3_1(.din(w_dff_B_DSabBSQw0_1),.dout(w_dff_B_wYbgBOcU3_1),.clk(gclk));
	jdff dff_B_7BPj9n451_1(.din(w_dff_B_wYbgBOcU3_1),.dout(w_dff_B_7BPj9n451_1),.clk(gclk));
	jdff dff_B_nQ2cNvO85_1(.din(w_dff_B_7BPj9n451_1),.dout(w_dff_B_nQ2cNvO85_1),.clk(gclk));
	jdff dff_B_OjKeyUXM1_1(.din(w_dff_B_nQ2cNvO85_1),.dout(w_dff_B_OjKeyUXM1_1),.clk(gclk));
	jdff dff_B_ctM5bRNX0_1(.din(w_dff_B_OjKeyUXM1_1),.dout(w_dff_B_ctM5bRNX0_1),.clk(gclk));
	jdff dff_B_j1GPd84g8_1(.din(w_dff_B_ctM5bRNX0_1),.dout(w_dff_B_j1GPd84g8_1),.clk(gclk));
	jdff dff_B_qDT9jkU24_1(.din(w_dff_B_j1GPd84g8_1),.dout(w_dff_B_qDT9jkU24_1),.clk(gclk));
	jdff dff_B_9hYt5XTP8_1(.din(w_dff_B_qDT9jkU24_1),.dout(w_dff_B_9hYt5XTP8_1),.clk(gclk));
	jdff dff_B_nxXT2Woi2_0(.din(n1620),.dout(w_dff_B_nxXT2Woi2_0),.clk(gclk));
	jdff dff_B_5fQYakNd8_0(.din(w_dff_B_nxXT2Woi2_0),.dout(w_dff_B_5fQYakNd8_0),.clk(gclk));
	jdff dff_B_IqNuwjlM2_0(.din(w_dff_B_5fQYakNd8_0),.dout(w_dff_B_IqNuwjlM2_0),.clk(gclk));
	jdff dff_B_cWKUjQgH9_0(.din(w_dff_B_IqNuwjlM2_0),.dout(w_dff_B_cWKUjQgH9_0),.clk(gclk));
	jdff dff_B_7mwu9n2e0_0(.din(w_dff_B_cWKUjQgH9_0),.dout(w_dff_B_7mwu9n2e0_0),.clk(gclk));
	jdff dff_B_zY4VCRG69_0(.din(w_dff_B_7mwu9n2e0_0),.dout(w_dff_B_zY4VCRG69_0),.clk(gclk));
	jdff dff_B_Nie2abV93_0(.din(w_dff_B_zY4VCRG69_0),.dout(w_dff_B_Nie2abV93_0),.clk(gclk));
	jdff dff_B_JCTp6ct86_0(.din(w_dff_B_Nie2abV93_0),.dout(w_dff_B_JCTp6ct86_0),.clk(gclk));
	jdff dff_A_Vm8e3S9c9_1(.dout(w_n1617_0[1]),.din(w_dff_A_Vm8e3S9c9_1),.clk(gclk));
	jdff dff_A_LTLZkO4D4_1(.dout(w_dff_A_Vm8e3S9c9_1),.din(w_dff_A_LTLZkO4D4_1),.clk(gclk));
	jdff dff_A_YNaUGyI08_1(.dout(w_dff_A_LTLZkO4D4_1),.din(w_dff_A_YNaUGyI08_1),.clk(gclk));
	jdff dff_A_YdmhWq4o0_1(.dout(w_dff_A_YNaUGyI08_1),.din(w_dff_A_YdmhWq4o0_1),.clk(gclk));
	jdff dff_A_aH0kG7nK6_1(.dout(w_dff_A_YdmhWq4o0_1),.din(w_dff_A_aH0kG7nK6_1),.clk(gclk));
	jdff dff_A_nkz9XtE07_1(.dout(w_dff_A_aH0kG7nK6_1),.din(w_dff_A_nkz9XtE07_1),.clk(gclk));
	jdff dff_A_H7g02P1A2_1(.dout(w_dff_A_nkz9XtE07_1),.din(w_dff_A_H7g02P1A2_1),.clk(gclk));
	jdff dff_A_eDaLSKlu8_1(.dout(w_dff_A_H7g02P1A2_1),.din(w_dff_A_eDaLSKlu8_1),.clk(gclk));
	jdff dff_A_IMnnVenA9_1(.dout(w_dff_A_eDaLSKlu8_1),.din(w_dff_A_IMnnVenA9_1),.clk(gclk));
	jdff dff_B_n4RELTC35_1(.din(n1557),.dout(w_dff_B_n4RELTC35_1),.clk(gclk));
	jdff dff_B_XgKRyzh94_1(.din(w_dff_B_n4RELTC35_1),.dout(w_dff_B_XgKRyzh94_1),.clk(gclk));
	jdff dff_B_RhTGLby80_1(.din(w_dff_B_XgKRyzh94_1),.dout(w_dff_B_RhTGLby80_1),.clk(gclk));
	jdff dff_B_ZRKTzA5T5_1(.din(w_dff_B_RhTGLby80_1),.dout(w_dff_B_ZRKTzA5T5_1),.clk(gclk));
	jdff dff_B_BGWNLnmi0_1(.din(w_dff_B_ZRKTzA5T5_1),.dout(w_dff_B_BGWNLnmi0_1),.clk(gclk));
	jdff dff_B_DP6C2C9o9_1(.din(w_dff_B_BGWNLnmi0_1),.dout(w_dff_B_DP6C2C9o9_1),.clk(gclk));
	jdff dff_B_LfiWfs5q6_1(.din(w_dff_B_DP6C2C9o9_1),.dout(w_dff_B_LfiWfs5q6_1),.clk(gclk));
	jdff dff_B_a8uOOsQh7_1(.din(w_dff_B_LfiWfs5q6_1),.dout(w_dff_B_a8uOOsQh7_1),.clk(gclk));
	jdff dff_B_kZXr2ywO9_0(.din(n1558),.dout(w_dff_B_kZXr2ywO9_0),.clk(gclk));
	jdff dff_B_tfKKtK025_0(.din(w_dff_B_kZXr2ywO9_0),.dout(w_dff_B_tfKKtK025_0),.clk(gclk));
	jdff dff_B_SSCxDJ4F7_0(.din(w_dff_B_tfKKtK025_0),.dout(w_dff_B_SSCxDJ4F7_0),.clk(gclk));
	jdff dff_B_nr4biGt38_0(.din(w_dff_B_SSCxDJ4F7_0),.dout(w_dff_B_nr4biGt38_0),.clk(gclk));
	jdff dff_B_CZlildiN7_0(.din(w_dff_B_nr4biGt38_0),.dout(w_dff_B_CZlildiN7_0),.clk(gclk));
	jdff dff_B_vDfTjoF11_0(.din(w_dff_B_CZlildiN7_0),.dout(w_dff_B_vDfTjoF11_0),.clk(gclk));
	jdff dff_A_b56HJCUi8_1(.dout(w_n1555_0[1]),.din(w_dff_A_b56HJCUi8_1),.clk(gclk));
	jdff dff_A_qSmd7q688_1(.dout(w_dff_A_b56HJCUi8_1),.din(w_dff_A_qSmd7q688_1),.clk(gclk));
	jdff dff_A_ZTURvvJv4_1(.dout(w_dff_A_qSmd7q688_1),.din(w_dff_A_ZTURvvJv4_1),.clk(gclk));
	jdff dff_A_qir4WC4H3_1(.dout(w_dff_A_ZTURvvJv4_1),.din(w_dff_A_qir4WC4H3_1),.clk(gclk));
	jdff dff_A_qTk1zyAX2_1(.dout(w_dff_A_qir4WC4H3_1),.din(w_dff_A_qTk1zyAX2_1),.clk(gclk));
	jdff dff_A_YdbMfr8e5_1(.dout(w_dff_A_qTk1zyAX2_1),.din(w_dff_A_YdbMfr8e5_1),.clk(gclk));
	jdff dff_A_GWaUef9G5_1(.dout(w_dff_A_YdbMfr8e5_1),.din(w_dff_A_GWaUef9G5_1),.clk(gclk));
	jdff dff_B_USfsmGXm0_1(.din(n1488),.dout(w_dff_B_USfsmGXm0_1),.clk(gclk));
	jdff dff_B_lWRSwoYc0_1(.din(w_dff_B_USfsmGXm0_1),.dout(w_dff_B_lWRSwoYc0_1),.clk(gclk));
	jdff dff_B_sdsv42lk8_1(.din(w_dff_B_lWRSwoYc0_1),.dout(w_dff_B_sdsv42lk8_1),.clk(gclk));
	jdff dff_B_XQRFyYYN7_1(.din(w_dff_B_sdsv42lk8_1),.dout(w_dff_B_XQRFyYYN7_1),.clk(gclk));
	jdff dff_B_HeOI2PSo2_1(.din(w_dff_B_XQRFyYYN7_1),.dout(w_dff_B_HeOI2PSo2_1),.clk(gclk));
	jdff dff_B_Ry5I1mhL5_1(.din(w_dff_B_HeOI2PSo2_1),.dout(w_dff_B_Ry5I1mhL5_1),.clk(gclk));
	jdff dff_B_PspZc4QJ1_1(.din(w_dff_B_Ry5I1mhL5_1),.dout(w_dff_B_PspZc4QJ1_1),.clk(gclk));
	jdff dff_B_mpPu7rD83_0(.din(n1489),.dout(w_dff_B_mpPu7rD83_0),.clk(gclk));
	jdff dff_B_i3HfL7z81_0(.din(w_dff_B_mpPu7rD83_0),.dout(w_dff_B_i3HfL7z81_0),.clk(gclk));
	jdff dff_B_NvseCO2M7_0(.din(w_dff_B_i3HfL7z81_0),.dout(w_dff_B_NvseCO2M7_0),.clk(gclk));
	jdff dff_B_veZRmBQf5_0(.din(w_dff_B_NvseCO2M7_0),.dout(w_dff_B_veZRmBQf5_0),.clk(gclk));
	jdff dff_B_l8h2kqKv1_0(.din(w_dff_B_veZRmBQf5_0),.dout(w_dff_B_l8h2kqKv1_0),.clk(gclk));
	jdff dff_A_Tz4EQcmS4_1(.dout(w_n1486_0[1]),.din(w_dff_A_Tz4EQcmS4_1),.clk(gclk));
	jdff dff_A_pLs5YupV5_1(.dout(w_dff_A_Tz4EQcmS4_1),.din(w_dff_A_pLs5YupV5_1),.clk(gclk));
	jdff dff_A_W3HsODiu8_1(.dout(w_dff_A_pLs5YupV5_1),.din(w_dff_A_W3HsODiu8_1),.clk(gclk));
	jdff dff_A_gtlsd8vm0_1(.dout(w_dff_A_W3HsODiu8_1),.din(w_dff_A_gtlsd8vm0_1),.clk(gclk));
	jdff dff_A_ac1VM2QA6_1(.dout(w_dff_A_gtlsd8vm0_1),.din(w_dff_A_ac1VM2QA6_1),.clk(gclk));
	jdff dff_A_6OXjizs55_1(.dout(w_dff_A_ac1VM2QA6_1),.din(w_dff_A_6OXjizs55_1),.clk(gclk));
	jdff dff_B_tjKHlDfa3_1(.din(n1412),.dout(w_dff_B_tjKHlDfa3_1),.clk(gclk));
	jdff dff_B_FKK0XW893_1(.din(w_dff_B_tjKHlDfa3_1),.dout(w_dff_B_FKK0XW893_1),.clk(gclk));
	jdff dff_B_9NEI6zxU5_1(.din(w_dff_B_FKK0XW893_1),.dout(w_dff_B_9NEI6zxU5_1),.clk(gclk));
	jdff dff_B_GTSAcAkx5_1(.din(w_dff_B_9NEI6zxU5_1),.dout(w_dff_B_GTSAcAkx5_1),.clk(gclk));
	jdff dff_B_J2ojcNg75_1(.din(w_dff_B_GTSAcAkx5_1),.dout(w_dff_B_J2ojcNg75_1),.clk(gclk));
	jdff dff_B_G3MHIb661_1(.din(w_dff_B_J2ojcNg75_1),.dout(w_dff_B_G3MHIb661_1),.clk(gclk));
	jdff dff_B_rgvWZtm54_0(.din(n1413),.dout(w_dff_B_rgvWZtm54_0),.clk(gclk));
	jdff dff_B_jazBqxMe8_0(.din(w_dff_B_rgvWZtm54_0),.dout(w_dff_B_jazBqxMe8_0),.clk(gclk));
	jdff dff_B_saUc9m3L0_0(.din(w_dff_B_jazBqxMe8_0),.dout(w_dff_B_saUc9m3L0_0),.clk(gclk));
	jdff dff_B_SJt7GV7E3_0(.din(w_dff_B_saUc9m3L0_0),.dout(w_dff_B_SJt7GV7E3_0),.clk(gclk));
	jdff dff_A_teWPpJ3x2_1(.dout(w_n1410_0[1]),.din(w_dff_A_teWPpJ3x2_1),.clk(gclk));
	jdff dff_A_f3GD0nUL2_1(.dout(w_dff_A_teWPpJ3x2_1),.din(w_dff_A_f3GD0nUL2_1),.clk(gclk));
	jdff dff_A_BTauswms8_1(.dout(w_dff_A_f3GD0nUL2_1),.din(w_dff_A_BTauswms8_1),.clk(gclk));
	jdff dff_A_IBuaDJlC0_1(.dout(w_dff_A_BTauswms8_1),.din(w_dff_A_IBuaDJlC0_1),.clk(gclk));
	jdff dff_A_lgICghwQ9_1(.dout(w_dff_A_IBuaDJlC0_1),.din(w_dff_A_lgICghwQ9_1),.clk(gclk));
	jdff dff_B_frxD2xVz1_1(.din(n1330),.dout(w_dff_B_frxD2xVz1_1),.clk(gclk));
	jdff dff_B_g5XiQJX29_1(.din(w_dff_B_frxD2xVz1_1),.dout(w_dff_B_g5XiQJX29_1),.clk(gclk));
	jdff dff_B_GlvTNpIt5_1(.din(w_dff_B_g5XiQJX29_1),.dout(w_dff_B_GlvTNpIt5_1),.clk(gclk));
	jdff dff_A_mSqC7HeX1_0(.dout(w_n1326_0[0]),.din(w_dff_A_mSqC7HeX1_0),.clk(gclk));
	jdff dff_A_Fc4YPKTA5_0(.dout(w_dff_A_mSqC7HeX1_0),.din(w_dff_A_Fc4YPKTA5_0),.clk(gclk));
	jdff dff_B_2vRuOUkq5_1(.din(n1242),.dout(w_dff_B_2vRuOUkq5_1),.clk(gclk));
	jdff dff_A_YtIxMlso6_0(.dout(w_n1238_0[0]),.din(w_dff_A_YtIxMlso6_0),.clk(gclk));
	jdff dff_B_jo2C4wSM4_1(.din(n1145),.dout(w_dff_B_jo2C4wSM4_1),.clk(gclk));
	jdff dff_A_8iyxgJFi0_1(.dout(w_n1039_0[1]),.din(w_dff_A_8iyxgJFi0_1),.clk(gclk));
	jdff dff_B_sIVTiUs64_2(.din(n1037),.dout(w_dff_B_sIVTiUs64_2),.clk(gclk));
	jdff dff_B_byKfvmww9_1(.din(n935),.dout(w_dff_B_byKfvmww9_1),.clk(gclk));
	jdff dff_A_qNRg8aGX1_0(.dout(w_n829_0[0]),.din(w_dff_A_qNRg8aGX1_0),.clk(gclk));
	jdff dff_A_JgXN2zTt1_0(.dout(w_dff_A_qNRg8aGX1_0),.din(w_dff_A_JgXN2zTt1_0),.clk(gclk));
	jdff dff_A_DfQ8exKU5_0(.dout(w_dff_A_JgXN2zTt1_0),.din(w_dff_A_DfQ8exKU5_0),.clk(gclk));
	jdff dff_A_XtxeZWxf2_0(.dout(w_dff_A_DfQ8exKU5_0),.din(w_dff_A_XtxeZWxf2_0),.clk(gclk));
	jdff dff_A_HCtayFC97_0(.dout(w_dff_A_XtxeZWxf2_0),.din(w_dff_A_HCtayFC97_0),.clk(gclk));
	jdff dff_A_80Tal6Wq3_0(.dout(w_dff_A_HCtayFC97_0),.din(w_dff_A_80Tal6Wq3_0),.clk(gclk));
	jdff dff_A_17tMaAR57_0(.dout(w_dff_A_80Tal6Wq3_0),.din(w_dff_A_17tMaAR57_0),.clk(gclk));
	jdff dff_A_UBTuDwGq1_0(.dout(w_dff_A_17tMaAR57_0),.din(w_dff_A_UBTuDwGq1_0),.clk(gclk));
	jdff dff_A_oUoOvbm24_0(.dout(w_dff_A_UBTuDwGq1_0),.din(w_dff_A_oUoOvbm24_0),.clk(gclk));
	jdff dff_A_hBNQuMGh6_0(.dout(w_dff_A_oUoOvbm24_0),.din(w_dff_A_hBNQuMGh6_0),.clk(gclk));
	jdff dff_A_ZYSSPDsR3_0(.dout(w_dff_A_hBNQuMGh6_0),.din(w_dff_A_ZYSSPDsR3_0),.clk(gclk));
	jdff dff_A_lvVskOPa4_0(.dout(w_dff_A_ZYSSPDsR3_0),.din(w_dff_A_lvVskOPa4_0),.clk(gclk));
	jdff dff_A_sifpBE7k8_0(.dout(w_dff_A_lvVskOPa4_0),.din(w_dff_A_sifpBE7k8_0),.clk(gclk));
	jdff dff_A_RmpMzXNi0_0(.dout(w_dff_A_sifpBE7k8_0),.din(w_dff_A_RmpMzXNi0_0),.clk(gclk));
	jdff dff_A_VO2i2IdE4_0(.dout(w_dff_A_RmpMzXNi0_0),.din(w_dff_A_VO2i2IdE4_0),.clk(gclk));
	jdff dff_A_GYSUPLGE8_0(.dout(w_dff_A_VO2i2IdE4_0),.din(w_dff_A_GYSUPLGE8_0),.clk(gclk));
	jdff dff_A_k1Zd2eOK2_0(.dout(w_dff_A_GYSUPLGE8_0),.din(w_dff_A_k1Zd2eOK2_0),.clk(gclk));
	jdff dff_A_alQEwqyh8_0(.dout(w_dff_A_k1Zd2eOK2_0),.din(w_dff_A_alQEwqyh8_0),.clk(gclk));
	jdff dff_A_Lby3IRmd5_0(.dout(w_dff_A_alQEwqyh8_0),.din(w_dff_A_Lby3IRmd5_0),.clk(gclk));
	jdff dff_A_STlUFQBE4_0(.dout(w_dff_A_Lby3IRmd5_0),.din(w_dff_A_STlUFQBE4_0),.clk(gclk));
	jdff dff_A_CburmB6r4_0(.dout(w_dff_A_STlUFQBE4_0),.din(w_dff_A_CburmB6r4_0),.clk(gclk));
	jdff dff_A_TwfLiWdX0_0(.dout(w_dff_A_CburmB6r4_0),.din(w_dff_A_TwfLiWdX0_0),.clk(gclk));
	jdff dff_A_phh4mHJV9_0(.dout(w_dff_A_TwfLiWdX0_0),.din(w_dff_A_phh4mHJV9_0),.clk(gclk));
	jdff dff_A_5kSOOloa8_0(.dout(w_dff_A_phh4mHJV9_0),.din(w_dff_A_5kSOOloa8_0),.clk(gclk));
	jdff dff_A_nRGcuvUV7_0(.dout(w_dff_A_5kSOOloa8_0),.din(w_dff_A_nRGcuvUV7_0),.clk(gclk));
	jdff dff_A_wMLIcOJV0_0(.dout(w_dff_A_nRGcuvUV7_0),.din(w_dff_A_wMLIcOJV0_0),.clk(gclk));
	jdff dff_A_AW3zlEQG8_0(.dout(w_dff_A_wMLIcOJV0_0),.din(w_dff_A_AW3zlEQG8_0),.clk(gclk));
	jdff dff_A_IHV4G6Sb8_0(.dout(w_dff_A_AW3zlEQG8_0),.din(w_dff_A_IHV4G6Sb8_0),.clk(gclk));
	jdff dff_A_5b8AV0XN8_0(.dout(w_dff_A_IHV4G6Sb8_0),.din(w_dff_A_5b8AV0XN8_0),.clk(gclk));
	jdff dff_A_DGqxklfv6_0(.dout(w_dff_A_5b8AV0XN8_0),.din(w_dff_A_DGqxklfv6_0),.clk(gclk));
	jdff dff_A_MjMeCmeQ8_0(.dout(w_dff_A_DGqxklfv6_0),.din(w_dff_A_MjMeCmeQ8_0),.clk(gclk));
	jdff dff_A_KDIwBGNi1_0(.dout(w_dff_A_MjMeCmeQ8_0),.din(w_dff_A_KDIwBGNi1_0),.clk(gclk));
	jdff dff_A_864cxI9s6_0(.dout(w_dff_A_KDIwBGNi1_0),.din(w_dff_A_864cxI9s6_0),.clk(gclk));
	jdff dff_A_PaXeYqjV7_0(.dout(w_dff_A_864cxI9s6_0),.din(w_dff_A_PaXeYqjV7_0),.clk(gclk));
	jdff dff_A_3xPJlGV88_0(.dout(w_dff_A_PaXeYqjV7_0),.din(w_dff_A_3xPJlGV88_0),.clk(gclk));
	jdff dff_A_R6u16fb98_0(.dout(w_dff_A_3xPJlGV88_0),.din(w_dff_A_R6u16fb98_0),.clk(gclk));
	jdff dff_A_tf8mc7TZ5_0(.dout(w_dff_A_R6u16fb98_0),.din(w_dff_A_tf8mc7TZ5_0),.clk(gclk));
	jdff dff_A_vDJPMjFE9_0(.dout(w_dff_A_tf8mc7TZ5_0),.din(w_dff_A_vDJPMjFE9_0),.clk(gclk));
	jdff dff_A_BvGu7WyE3_0(.dout(w_dff_A_vDJPMjFE9_0),.din(w_dff_A_BvGu7WyE3_0),.clk(gclk));
	jdff dff_A_h5l2llis0_0(.dout(w_dff_A_BvGu7WyE3_0),.din(w_dff_A_h5l2llis0_0),.clk(gclk));
	jdff dff_A_TvAQHO4q6_0(.dout(w_dff_A_h5l2llis0_0),.din(w_dff_A_TvAQHO4q6_0),.clk(gclk));
	jdff dff_A_xyr3zLB41_0(.dout(w_dff_A_TvAQHO4q6_0),.din(w_dff_A_xyr3zLB41_0),.clk(gclk));
	jdff dff_A_lMon71Tu2_0(.dout(w_dff_A_xyr3zLB41_0),.din(w_dff_A_lMon71Tu2_0),.clk(gclk));
	jdff dff_A_kyZTZRFM8_0(.dout(w_dff_A_lMon71Tu2_0),.din(w_dff_A_kyZTZRFM8_0),.clk(gclk));
	jdff dff_A_rPD8mdkc9_1(.dout(w_n931_0[1]),.din(w_dff_A_rPD8mdkc9_1),.clk(gclk));
	jdff dff_B_WUFQEIHg0_1(.din(n832),.dout(w_dff_B_WUFQEIHg0_1),.clk(gclk));
	jdff dff_A_t3yutd8v3_0(.dout(w_n729_0[0]),.din(w_dff_A_t3yutd8v3_0),.clk(gclk));
	jdff dff_A_2IW4mItI8_0(.dout(w_dff_A_t3yutd8v3_0),.din(w_dff_A_2IW4mItI8_0),.clk(gclk));
	jdff dff_A_vlMTcgpY1_0(.dout(w_dff_A_2IW4mItI8_0),.din(w_dff_A_vlMTcgpY1_0),.clk(gclk));
	jdff dff_A_fbo78wwa9_0(.dout(w_dff_A_vlMTcgpY1_0),.din(w_dff_A_fbo78wwa9_0),.clk(gclk));
	jdff dff_A_4R9mg1Gv7_0(.dout(w_dff_A_fbo78wwa9_0),.din(w_dff_A_4R9mg1Gv7_0),.clk(gclk));
	jdff dff_A_vTHGO2To3_0(.dout(w_dff_A_4R9mg1Gv7_0),.din(w_dff_A_vTHGO2To3_0),.clk(gclk));
	jdff dff_A_jQ28pvgX0_0(.dout(w_dff_A_vTHGO2To3_0),.din(w_dff_A_jQ28pvgX0_0),.clk(gclk));
	jdff dff_A_9q6bxR0N9_0(.dout(w_dff_A_jQ28pvgX0_0),.din(w_dff_A_9q6bxR0N9_0),.clk(gclk));
	jdff dff_A_Yahpox9g3_0(.dout(w_dff_A_9q6bxR0N9_0),.din(w_dff_A_Yahpox9g3_0),.clk(gclk));
	jdff dff_A_RKyrTVUw0_0(.dout(w_dff_A_Yahpox9g3_0),.din(w_dff_A_RKyrTVUw0_0),.clk(gclk));
	jdff dff_A_DrxZLU1J7_0(.dout(w_dff_A_RKyrTVUw0_0),.din(w_dff_A_DrxZLU1J7_0),.clk(gclk));
	jdff dff_A_drsOUfEZ3_0(.dout(w_dff_A_DrxZLU1J7_0),.din(w_dff_A_drsOUfEZ3_0),.clk(gclk));
	jdff dff_A_HuVd3Y6V7_0(.dout(w_dff_A_drsOUfEZ3_0),.din(w_dff_A_HuVd3Y6V7_0),.clk(gclk));
	jdff dff_A_e74l0oWE2_0(.dout(w_dff_A_HuVd3Y6V7_0),.din(w_dff_A_e74l0oWE2_0),.clk(gclk));
	jdff dff_A_I04age3X6_0(.dout(w_dff_A_e74l0oWE2_0),.din(w_dff_A_I04age3X6_0),.clk(gclk));
	jdff dff_A_cnvKZSoj3_0(.dout(w_dff_A_I04age3X6_0),.din(w_dff_A_cnvKZSoj3_0),.clk(gclk));
	jdff dff_A_rFllEZ7S9_0(.dout(w_dff_A_cnvKZSoj3_0),.din(w_dff_A_rFllEZ7S9_0),.clk(gclk));
	jdff dff_A_ArdhJ4v70_0(.dout(w_dff_A_rFllEZ7S9_0),.din(w_dff_A_ArdhJ4v70_0),.clk(gclk));
	jdff dff_A_t8FkTvUv5_0(.dout(w_dff_A_ArdhJ4v70_0),.din(w_dff_A_t8FkTvUv5_0),.clk(gclk));
	jdff dff_A_TIzXt2Qc1_0(.dout(w_dff_A_t8FkTvUv5_0),.din(w_dff_A_TIzXt2Qc1_0),.clk(gclk));
	jdff dff_A_wcACY4Mm1_0(.dout(w_dff_A_TIzXt2Qc1_0),.din(w_dff_A_wcACY4Mm1_0),.clk(gclk));
	jdff dff_A_9s1Sia4g4_0(.dout(w_dff_A_wcACY4Mm1_0),.din(w_dff_A_9s1Sia4g4_0),.clk(gclk));
	jdff dff_A_VMbvWN9B1_0(.dout(w_dff_A_9s1Sia4g4_0),.din(w_dff_A_VMbvWN9B1_0),.clk(gclk));
	jdff dff_A_es8PT67q7_0(.dout(w_dff_A_VMbvWN9B1_0),.din(w_dff_A_es8PT67q7_0),.clk(gclk));
	jdff dff_A_3tZjujnG8_0(.dout(w_dff_A_es8PT67q7_0),.din(w_dff_A_3tZjujnG8_0),.clk(gclk));
	jdff dff_A_nKUHsgCu2_0(.dout(w_dff_A_3tZjujnG8_0),.din(w_dff_A_nKUHsgCu2_0),.clk(gclk));
	jdff dff_A_XHaYsywL2_0(.dout(w_dff_A_nKUHsgCu2_0),.din(w_dff_A_XHaYsywL2_0),.clk(gclk));
	jdff dff_A_mqhKkZ8E0_0(.dout(w_dff_A_XHaYsywL2_0),.din(w_dff_A_mqhKkZ8E0_0),.clk(gclk));
	jdff dff_A_4cySiSeH1_0(.dout(w_dff_A_mqhKkZ8E0_0),.din(w_dff_A_4cySiSeH1_0),.clk(gclk));
	jdff dff_A_HB7cFgzJ3_0(.dout(w_dff_A_4cySiSeH1_0),.din(w_dff_A_HB7cFgzJ3_0),.clk(gclk));
	jdff dff_A_hwbYGpQC2_0(.dout(w_dff_A_HB7cFgzJ3_0),.din(w_dff_A_hwbYGpQC2_0),.clk(gclk));
	jdff dff_A_dCYxRYtA2_0(.dout(w_dff_A_hwbYGpQC2_0),.din(w_dff_A_dCYxRYtA2_0),.clk(gclk));
	jdff dff_A_rVwR51FL1_0(.dout(w_dff_A_dCYxRYtA2_0),.din(w_dff_A_rVwR51FL1_0),.clk(gclk));
	jdff dff_A_5tASqAVF5_0(.dout(w_dff_A_rVwR51FL1_0),.din(w_dff_A_5tASqAVF5_0),.clk(gclk));
	jdff dff_A_UGPkjZmw0_0(.dout(w_dff_A_5tASqAVF5_0),.din(w_dff_A_UGPkjZmw0_0),.clk(gclk));
	jdff dff_A_EvEAvwR46_0(.dout(w_dff_A_UGPkjZmw0_0),.din(w_dff_A_EvEAvwR46_0),.clk(gclk));
	jdff dff_A_WMyZgvck7_0(.dout(w_dff_A_EvEAvwR46_0),.din(w_dff_A_WMyZgvck7_0),.clk(gclk));
	jdff dff_A_N6AoFGDw4_0(.dout(w_dff_A_WMyZgvck7_0),.din(w_dff_A_N6AoFGDw4_0),.clk(gclk));
	jdff dff_A_ApnZFqMo9_0(.dout(w_dff_A_N6AoFGDw4_0),.din(w_dff_A_ApnZFqMo9_0),.clk(gclk));
	jdff dff_A_8Taggs821_0(.dout(w_dff_A_ApnZFqMo9_0),.din(w_dff_A_8Taggs821_0),.clk(gclk));
	jdff dff_A_rg9oEtRT9_0(.dout(w_dff_A_8Taggs821_0),.din(w_dff_A_rg9oEtRT9_0),.clk(gclk));
	jdff dff_A_HUmEwnRZ3_1(.dout(w_n826_0[1]),.din(w_dff_A_HUmEwnRZ3_1),.clk(gclk));
	jdff dff_B_3t9gZx5K6_1(.din(n736),.dout(w_dff_B_3t9gZx5K6_1),.clk(gclk));
	jdff dff_B_L7VvIAtI3_1(.din(w_dff_B_3t9gZx5K6_1),.dout(w_dff_B_L7VvIAtI3_1),.clk(gclk));
	jdff dff_B_okdm2yDn5_1(.din(w_dff_B_L7VvIAtI3_1),.dout(w_dff_B_okdm2yDn5_1),.clk(gclk));
	jdff dff_B_vlaR4Psj6_1(.din(w_dff_B_okdm2yDn5_1),.dout(w_dff_B_vlaR4Psj6_1),.clk(gclk));
	jdff dff_B_TsRoWXeD1_1(.din(w_dff_B_vlaR4Psj6_1),.dout(w_dff_B_TsRoWXeD1_1),.clk(gclk));
	jdff dff_B_L6p6CLBb1_1(.din(w_dff_B_TsRoWXeD1_1),.dout(w_dff_B_L6p6CLBb1_1),.clk(gclk));
	jdff dff_B_YiE75Lzf9_1(.din(w_dff_B_L6p6CLBb1_1),.dout(w_dff_B_YiE75Lzf9_1),.clk(gclk));
	jdff dff_B_2zV4ajEy0_1(.din(w_dff_B_YiE75Lzf9_1),.dout(w_dff_B_2zV4ajEy0_1),.clk(gclk));
	jdff dff_B_D5roRV2S7_1(.din(w_dff_B_2zV4ajEy0_1),.dout(w_dff_B_D5roRV2S7_1),.clk(gclk));
	jdff dff_B_VLSOsmEX6_1(.din(w_dff_B_D5roRV2S7_1),.dout(w_dff_B_VLSOsmEX6_1),.clk(gclk));
	jdff dff_B_8SXLJU0a1_1(.din(w_dff_B_VLSOsmEX6_1),.dout(w_dff_B_8SXLJU0a1_1),.clk(gclk));
	jdff dff_B_0hnHS7hT4_1(.din(w_dff_B_8SXLJU0a1_1),.dout(w_dff_B_0hnHS7hT4_1),.clk(gclk));
	jdff dff_B_MzaqPRWa0_1(.din(w_dff_B_0hnHS7hT4_1),.dout(w_dff_B_MzaqPRWa0_1),.clk(gclk));
	jdff dff_B_5dBb4DJN7_1(.din(w_dff_B_MzaqPRWa0_1),.dout(w_dff_B_5dBb4DJN7_1),.clk(gclk));
	jdff dff_B_bL39RRKl0_1(.din(w_dff_B_5dBb4DJN7_1),.dout(w_dff_B_bL39RRKl0_1),.clk(gclk));
	jdff dff_B_SqYK75VZ2_1(.din(w_dff_B_bL39RRKl0_1),.dout(w_dff_B_SqYK75VZ2_1),.clk(gclk));
	jdff dff_B_31AAucs20_1(.din(w_dff_B_SqYK75VZ2_1),.dout(w_dff_B_31AAucs20_1),.clk(gclk));
	jdff dff_B_otlpwXtr3_1(.din(w_dff_B_31AAucs20_1),.dout(w_dff_B_otlpwXtr3_1),.clk(gclk));
	jdff dff_B_v6pmgBCp7_1(.din(w_dff_B_otlpwXtr3_1),.dout(w_dff_B_v6pmgBCp7_1),.clk(gclk));
	jdff dff_B_B8LIxpM91_1(.din(w_dff_B_v6pmgBCp7_1),.dout(w_dff_B_B8LIxpM91_1),.clk(gclk));
	jdff dff_B_JPKN5Tqy6_1(.din(w_dff_B_B8LIxpM91_1),.dout(w_dff_B_JPKN5Tqy6_1),.clk(gclk));
	jdff dff_B_HxKgMiqD4_1(.din(w_dff_B_JPKN5Tqy6_1),.dout(w_dff_B_HxKgMiqD4_1),.clk(gclk));
	jdff dff_B_Scn7qKiP2_1(.din(w_dff_B_HxKgMiqD4_1),.dout(w_dff_B_Scn7qKiP2_1),.clk(gclk));
	jdff dff_B_HFWmZ27m9_1(.din(w_dff_B_Scn7qKiP2_1),.dout(w_dff_B_HFWmZ27m9_1),.clk(gclk));
	jdff dff_B_K3Nt58Zx1_1(.din(w_dff_B_HFWmZ27m9_1),.dout(w_dff_B_K3Nt58Zx1_1),.clk(gclk));
	jdff dff_B_NTV7a2sP9_1(.din(w_dff_B_K3Nt58Zx1_1),.dout(w_dff_B_NTV7a2sP9_1),.clk(gclk));
	jdff dff_B_sMCjv46i2_1(.din(w_dff_B_NTV7a2sP9_1),.dout(w_dff_B_sMCjv46i2_1),.clk(gclk));
	jdff dff_B_VHZkwYA20_1(.din(w_dff_B_sMCjv46i2_1),.dout(w_dff_B_VHZkwYA20_1),.clk(gclk));
	jdff dff_B_sfJyiSy11_1(.din(w_dff_B_VHZkwYA20_1),.dout(w_dff_B_sfJyiSy11_1),.clk(gclk));
	jdff dff_B_G652oqZV7_1(.din(w_dff_B_sfJyiSy11_1),.dout(w_dff_B_G652oqZV7_1),.clk(gclk));
	jdff dff_B_Kw3aQ7mJ5_1(.din(w_dff_B_G652oqZV7_1),.dout(w_dff_B_Kw3aQ7mJ5_1),.clk(gclk));
	jdff dff_B_7HOgLgjF9_1(.din(w_dff_B_Kw3aQ7mJ5_1),.dout(w_dff_B_7HOgLgjF9_1),.clk(gclk));
	jdff dff_B_2rB4suMf6_1(.din(w_dff_B_7HOgLgjF9_1),.dout(w_dff_B_2rB4suMf6_1),.clk(gclk));
	jdff dff_B_Tt7ssnoQ1_1(.din(w_dff_B_2rB4suMf6_1),.dout(w_dff_B_Tt7ssnoQ1_1),.clk(gclk));
	jdff dff_B_BAK52qaT6_1(.din(w_dff_B_Tt7ssnoQ1_1),.dout(w_dff_B_BAK52qaT6_1),.clk(gclk));
	jdff dff_B_08Y2FHn92_1(.din(w_dff_B_BAK52qaT6_1),.dout(w_dff_B_08Y2FHn92_1),.clk(gclk));
	jdff dff_B_APixYkF69_1(.din(w_dff_B_08Y2FHn92_1),.dout(w_dff_B_APixYkF69_1),.clk(gclk));
	jdff dff_B_jxu3HVWu3_1(.din(n732),.dout(w_dff_B_jxu3HVWu3_1),.clk(gclk));
	jdff dff_A_3Se68il30_0(.dout(w_n636_0[0]),.din(w_dff_A_3Se68il30_0),.clk(gclk));
	jdff dff_A_qegC0KNM3_0(.dout(w_dff_A_3Se68il30_0),.din(w_dff_A_qegC0KNM3_0),.clk(gclk));
	jdff dff_A_T7PijzyN8_0(.dout(w_dff_A_qegC0KNM3_0),.din(w_dff_A_T7PijzyN8_0),.clk(gclk));
	jdff dff_A_U99S566E9_0(.dout(w_dff_A_T7PijzyN8_0),.din(w_dff_A_U99S566E9_0),.clk(gclk));
	jdff dff_A_a5F5TQay5_0(.dout(w_dff_A_U99S566E9_0),.din(w_dff_A_a5F5TQay5_0),.clk(gclk));
	jdff dff_A_gYHFqeoV4_0(.dout(w_dff_A_a5F5TQay5_0),.din(w_dff_A_gYHFqeoV4_0),.clk(gclk));
	jdff dff_A_Ixnpqw4C1_0(.dout(w_dff_A_gYHFqeoV4_0),.din(w_dff_A_Ixnpqw4C1_0),.clk(gclk));
	jdff dff_A_H5hEAAHK7_0(.dout(w_dff_A_Ixnpqw4C1_0),.din(w_dff_A_H5hEAAHK7_0),.clk(gclk));
	jdff dff_A_tzzZlqe55_0(.dout(w_dff_A_H5hEAAHK7_0),.din(w_dff_A_tzzZlqe55_0),.clk(gclk));
	jdff dff_A_gsbXq6Qo4_0(.dout(w_dff_A_tzzZlqe55_0),.din(w_dff_A_gsbXq6Qo4_0),.clk(gclk));
	jdff dff_A_Eiy7Uz6W0_0(.dout(w_dff_A_gsbXq6Qo4_0),.din(w_dff_A_Eiy7Uz6W0_0),.clk(gclk));
	jdff dff_A_KtEIAcWO1_0(.dout(w_dff_A_Eiy7Uz6W0_0),.din(w_dff_A_KtEIAcWO1_0),.clk(gclk));
	jdff dff_A_CZOV7ISu0_0(.dout(w_dff_A_KtEIAcWO1_0),.din(w_dff_A_CZOV7ISu0_0),.clk(gclk));
	jdff dff_A_hom3Zi0f2_0(.dout(w_dff_A_CZOV7ISu0_0),.din(w_dff_A_hom3Zi0f2_0),.clk(gclk));
	jdff dff_A_I8A3ZDls4_0(.dout(w_dff_A_hom3Zi0f2_0),.din(w_dff_A_I8A3ZDls4_0),.clk(gclk));
	jdff dff_A_EAJPG4996_0(.dout(w_dff_A_I8A3ZDls4_0),.din(w_dff_A_EAJPG4996_0),.clk(gclk));
	jdff dff_A_O4TzIQaN9_0(.dout(w_dff_A_EAJPG4996_0),.din(w_dff_A_O4TzIQaN9_0),.clk(gclk));
	jdff dff_A_o6ONkrSf6_0(.dout(w_dff_A_O4TzIQaN9_0),.din(w_dff_A_o6ONkrSf6_0),.clk(gclk));
	jdff dff_A_3eR9Xw4o1_0(.dout(w_dff_A_o6ONkrSf6_0),.din(w_dff_A_3eR9Xw4o1_0),.clk(gclk));
	jdff dff_A_7NH5S5IB5_0(.dout(w_dff_A_3eR9Xw4o1_0),.din(w_dff_A_7NH5S5IB5_0),.clk(gclk));
	jdff dff_A_R7hFAMTz8_0(.dout(w_dff_A_7NH5S5IB5_0),.din(w_dff_A_R7hFAMTz8_0),.clk(gclk));
	jdff dff_A_Kish0dB56_0(.dout(w_dff_A_R7hFAMTz8_0),.din(w_dff_A_Kish0dB56_0),.clk(gclk));
	jdff dff_A_tsK7WZvd3_0(.dout(w_dff_A_Kish0dB56_0),.din(w_dff_A_tsK7WZvd3_0),.clk(gclk));
	jdff dff_A_xG60JkBl0_0(.dout(w_dff_A_tsK7WZvd3_0),.din(w_dff_A_xG60JkBl0_0),.clk(gclk));
	jdff dff_A_mlHfyNgV3_0(.dout(w_dff_A_xG60JkBl0_0),.din(w_dff_A_mlHfyNgV3_0),.clk(gclk));
	jdff dff_A_Rci0Molr9_0(.dout(w_dff_A_mlHfyNgV3_0),.din(w_dff_A_Rci0Molr9_0),.clk(gclk));
	jdff dff_A_PVZvRimo4_0(.dout(w_dff_A_Rci0Molr9_0),.din(w_dff_A_PVZvRimo4_0),.clk(gclk));
	jdff dff_A_cag03PwF6_0(.dout(w_dff_A_PVZvRimo4_0),.din(w_dff_A_cag03PwF6_0),.clk(gclk));
	jdff dff_A_j1DM6ePW0_0(.dout(w_dff_A_cag03PwF6_0),.din(w_dff_A_j1DM6ePW0_0),.clk(gclk));
	jdff dff_A_BQnAje3Q7_0(.dout(w_dff_A_j1DM6ePW0_0),.din(w_dff_A_BQnAje3Q7_0),.clk(gclk));
	jdff dff_A_NhyM3Bc79_0(.dout(w_dff_A_BQnAje3Q7_0),.din(w_dff_A_NhyM3Bc79_0),.clk(gclk));
	jdff dff_A_Unu0pAN28_0(.dout(w_dff_A_NhyM3Bc79_0),.din(w_dff_A_Unu0pAN28_0),.clk(gclk));
	jdff dff_A_0kKlBQdF0_0(.dout(w_dff_A_Unu0pAN28_0),.din(w_dff_A_0kKlBQdF0_0),.clk(gclk));
	jdff dff_A_BgfZlWBi2_0(.dout(w_dff_A_0kKlBQdF0_0),.din(w_dff_A_BgfZlWBi2_0),.clk(gclk));
	jdff dff_A_PDnNGCep8_0(.dout(w_dff_A_BgfZlWBi2_0),.din(w_dff_A_PDnNGCep8_0),.clk(gclk));
	jdff dff_A_BRoNz3jn2_0(.dout(w_dff_A_PDnNGCep8_0),.din(w_dff_A_BRoNz3jn2_0),.clk(gclk));
	jdff dff_A_14cqpYVj0_0(.dout(w_dff_A_BRoNz3jn2_0),.din(w_dff_A_14cqpYVj0_0),.clk(gclk));
	jdff dff_A_iTXaZvbS8_0(.dout(w_dff_A_14cqpYVj0_0),.din(w_dff_A_iTXaZvbS8_0),.clk(gclk));
	jdff dff_A_9NszZZ8G3_1(.dout(w_n726_0[1]),.din(w_dff_A_9NszZZ8G3_1),.clk(gclk));
	jdff dff_B_lU9l0C5p5_1(.din(n643),.dout(w_dff_B_lU9l0C5p5_1),.clk(gclk));
	jdff dff_B_xrLqgSAx0_1(.din(w_dff_B_lU9l0C5p5_1),.dout(w_dff_B_xrLqgSAx0_1),.clk(gclk));
	jdff dff_B_monT6oy97_1(.din(w_dff_B_xrLqgSAx0_1),.dout(w_dff_B_monT6oy97_1),.clk(gclk));
	jdff dff_B_Tyc6hKCI3_1(.din(w_dff_B_monT6oy97_1),.dout(w_dff_B_Tyc6hKCI3_1),.clk(gclk));
	jdff dff_B_vi922Aph6_1(.din(w_dff_B_Tyc6hKCI3_1),.dout(w_dff_B_vi922Aph6_1),.clk(gclk));
	jdff dff_B_qvDo52W75_1(.din(w_dff_B_vi922Aph6_1),.dout(w_dff_B_qvDo52W75_1),.clk(gclk));
	jdff dff_B_noQNMYPZ2_1(.din(w_dff_B_qvDo52W75_1),.dout(w_dff_B_noQNMYPZ2_1),.clk(gclk));
	jdff dff_B_t80WDKL63_1(.din(w_dff_B_noQNMYPZ2_1),.dout(w_dff_B_t80WDKL63_1),.clk(gclk));
	jdff dff_B_OFx7J3Sg9_1(.din(w_dff_B_t80WDKL63_1),.dout(w_dff_B_OFx7J3Sg9_1),.clk(gclk));
	jdff dff_B_oW5DSX7p3_1(.din(w_dff_B_OFx7J3Sg9_1),.dout(w_dff_B_oW5DSX7p3_1),.clk(gclk));
	jdff dff_B_ueSlggYk1_1(.din(w_dff_B_oW5DSX7p3_1),.dout(w_dff_B_ueSlggYk1_1),.clk(gclk));
	jdff dff_B_AqGEbTsd4_1(.din(w_dff_B_ueSlggYk1_1),.dout(w_dff_B_AqGEbTsd4_1),.clk(gclk));
	jdff dff_B_ggtqc0Wz1_1(.din(w_dff_B_AqGEbTsd4_1),.dout(w_dff_B_ggtqc0Wz1_1),.clk(gclk));
	jdff dff_B_6P39f6xr3_1(.din(w_dff_B_ggtqc0Wz1_1),.dout(w_dff_B_6P39f6xr3_1),.clk(gclk));
	jdff dff_B_3GqyIPiY7_1(.din(w_dff_B_6P39f6xr3_1),.dout(w_dff_B_3GqyIPiY7_1),.clk(gclk));
	jdff dff_B_2bK0TQyd9_1(.din(w_dff_B_3GqyIPiY7_1),.dout(w_dff_B_2bK0TQyd9_1),.clk(gclk));
	jdff dff_B_eGtVeBXP3_1(.din(w_dff_B_2bK0TQyd9_1),.dout(w_dff_B_eGtVeBXP3_1),.clk(gclk));
	jdff dff_B_oR4LQKt69_1(.din(w_dff_B_eGtVeBXP3_1),.dout(w_dff_B_oR4LQKt69_1),.clk(gclk));
	jdff dff_B_hB3YcFAy3_1(.din(w_dff_B_oR4LQKt69_1),.dout(w_dff_B_hB3YcFAy3_1),.clk(gclk));
	jdff dff_B_VysaI1qI3_1(.din(w_dff_B_hB3YcFAy3_1),.dout(w_dff_B_VysaI1qI3_1),.clk(gclk));
	jdff dff_B_eK0D9hSg1_1(.din(w_dff_B_VysaI1qI3_1),.dout(w_dff_B_eK0D9hSg1_1),.clk(gclk));
	jdff dff_B_v5yPIENZ2_1(.din(w_dff_B_eK0D9hSg1_1),.dout(w_dff_B_v5yPIENZ2_1),.clk(gclk));
	jdff dff_B_WlQVzxEd2_1(.din(w_dff_B_v5yPIENZ2_1),.dout(w_dff_B_WlQVzxEd2_1),.clk(gclk));
	jdff dff_B_2puEdKtI9_1(.din(w_dff_B_WlQVzxEd2_1),.dout(w_dff_B_2puEdKtI9_1),.clk(gclk));
	jdff dff_B_w4bNLSnL4_1(.din(w_dff_B_2puEdKtI9_1),.dout(w_dff_B_w4bNLSnL4_1),.clk(gclk));
	jdff dff_B_05lzDWlB2_1(.din(w_dff_B_w4bNLSnL4_1),.dout(w_dff_B_05lzDWlB2_1),.clk(gclk));
	jdff dff_B_OeihB6SH1_1(.din(w_dff_B_05lzDWlB2_1),.dout(w_dff_B_OeihB6SH1_1),.clk(gclk));
	jdff dff_B_BbmTrQTR7_1(.din(w_dff_B_OeihB6SH1_1),.dout(w_dff_B_BbmTrQTR7_1),.clk(gclk));
	jdff dff_B_FqDt8CYB4_1(.din(w_dff_B_BbmTrQTR7_1),.dout(w_dff_B_FqDt8CYB4_1),.clk(gclk));
	jdff dff_B_LysVxLLV6_1(.din(w_dff_B_FqDt8CYB4_1),.dout(w_dff_B_LysVxLLV6_1),.clk(gclk));
	jdff dff_B_Gh9WNbTS0_1(.din(w_dff_B_LysVxLLV6_1),.dout(w_dff_B_Gh9WNbTS0_1),.clk(gclk));
	jdff dff_B_oly3NsYK1_1(.din(w_dff_B_Gh9WNbTS0_1),.dout(w_dff_B_oly3NsYK1_1),.clk(gclk));
	jdff dff_B_VPvJsWGj0_1(.din(w_dff_B_oly3NsYK1_1),.dout(w_dff_B_VPvJsWGj0_1),.clk(gclk));
	jdff dff_B_XsTpae6H8_1(.din(w_dff_B_VPvJsWGj0_1),.dout(w_dff_B_XsTpae6H8_1),.clk(gclk));
	jdff dff_B_5vRFOpjz6_1(.din(n639),.dout(w_dff_B_5vRFOpjz6_1),.clk(gclk));
	jdff dff_A_28fmAf4M3_0(.dout(w_n550_0[0]),.din(w_dff_A_28fmAf4M3_0),.clk(gclk));
	jdff dff_A_gv55jvDa9_0(.dout(w_dff_A_28fmAf4M3_0),.din(w_dff_A_gv55jvDa9_0),.clk(gclk));
	jdff dff_A_mUVL712O0_0(.dout(w_dff_A_gv55jvDa9_0),.din(w_dff_A_mUVL712O0_0),.clk(gclk));
	jdff dff_A_EVGLiU8n8_0(.dout(w_dff_A_mUVL712O0_0),.din(w_dff_A_EVGLiU8n8_0),.clk(gclk));
	jdff dff_A_lLe2K2uN4_0(.dout(w_dff_A_EVGLiU8n8_0),.din(w_dff_A_lLe2K2uN4_0),.clk(gclk));
	jdff dff_A_Q83hYziu9_0(.dout(w_dff_A_lLe2K2uN4_0),.din(w_dff_A_Q83hYziu9_0),.clk(gclk));
	jdff dff_A_JhB8Y5r74_0(.dout(w_dff_A_Q83hYziu9_0),.din(w_dff_A_JhB8Y5r74_0),.clk(gclk));
	jdff dff_A_YcPnmJBb5_0(.dout(w_dff_A_JhB8Y5r74_0),.din(w_dff_A_YcPnmJBb5_0),.clk(gclk));
	jdff dff_A_wwubtDUj4_0(.dout(w_dff_A_YcPnmJBb5_0),.din(w_dff_A_wwubtDUj4_0),.clk(gclk));
	jdff dff_A_D94wLc9M4_0(.dout(w_dff_A_wwubtDUj4_0),.din(w_dff_A_D94wLc9M4_0),.clk(gclk));
	jdff dff_A_uwkHHHXP5_0(.dout(w_dff_A_D94wLc9M4_0),.din(w_dff_A_uwkHHHXP5_0),.clk(gclk));
	jdff dff_A_ev3T4ELG1_0(.dout(w_dff_A_uwkHHHXP5_0),.din(w_dff_A_ev3T4ELG1_0),.clk(gclk));
	jdff dff_A_YbTiujcb2_0(.dout(w_dff_A_ev3T4ELG1_0),.din(w_dff_A_YbTiujcb2_0),.clk(gclk));
	jdff dff_A_WsLhl5zJ4_0(.dout(w_dff_A_YbTiujcb2_0),.din(w_dff_A_WsLhl5zJ4_0),.clk(gclk));
	jdff dff_A_qeBLLR2w4_0(.dout(w_dff_A_WsLhl5zJ4_0),.din(w_dff_A_qeBLLR2w4_0),.clk(gclk));
	jdff dff_A_2Fgg3fG85_0(.dout(w_dff_A_qeBLLR2w4_0),.din(w_dff_A_2Fgg3fG85_0),.clk(gclk));
	jdff dff_A_JDd2GKi55_0(.dout(w_dff_A_2Fgg3fG85_0),.din(w_dff_A_JDd2GKi55_0),.clk(gclk));
	jdff dff_A_64SMlF383_0(.dout(w_dff_A_JDd2GKi55_0),.din(w_dff_A_64SMlF383_0),.clk(gclk));
	jdff dff_A_su2s0Tvr5_0(.dout(w_dff_A_64SMlF383_0),.din(w_dff_A_su2s0Tvr5_0),.clk(gclk));
	jdff dff_A_aRAuyn407_0(.dout(w_dff_A_su2s0Tvr5_0),.din(w_dff_A_aRAuyn407_0),.clk(gclk));
	jdff dff_A_xA13lmIc0_0(.dout(w_dff_A_aRAuyn407_0),.din(w_dff_A_xA13lmIc0_0),.clk(gclk));
	jdff dff_A_DTTdvm9I0_0(.dout(w_dff_A_xA13lmIc0_0),.din(w_dff_A_DTTdvm9I0_0),.clk(gclk));
	jdff dff_A_PTgevmWC4_0(.dout(w_dff_A_DTTdvm9I0_0),.din(w_dff_A_PTgevmWC4_0),.clk(gclk));
	jdff dff_A_NcbltGHV6_0(.dout(w_dff_A_PTgevmWC4_0),.din(w_dff_A_NcbltGHV6_0),.clk(gclk));
	jdff dff_A_kprWxV2v2_0(.dout(w_dff_A_NcbltGHV6_0),.din(w_dff_A_kprWxV2v2_0),.clk(gclk));
	jdff dff_A_sxDBOWrp1_0(.dout(w_dff_A_kprWxV2v2_0),.din(w_dff_A_sxDBOWrp1_0),.clk(gclk));
	jdff dff_A_RSMlVI9d3_0(.dout(w_dff_A_sxDBOWrp1_0),.din(w_dff_A_RSMlVI9d3_0),.clk(gclk));
	jdff dff_A_HrUUWE7i2_0(.dout(w_dff_A_RSMlVI9d3_0),.din(w_dff_A_HrUUWE7i2_0),.clk(gclk));
	jdff dff_A_XE4UNfHk2_0(.dout(w_dff_A_HrUUWE7i2_0),.din(w_dff_A_XE4UNfHk2_0),.clk(gclk));
	jdff dff_A_Thmjh4gW0_0(.dout(w_dff_A_XE4UNfHk2_0),.din(w_dff_A_Thmjh4gW0_0),.clk(gclk));
	jdff dff_A_2rnCKYeo7_0(.dout(w_dff_A_Thmjh4gW0_0),.din(w_dff_A_2rnCKYeo7_0),.clk(gclk));
	jdff dff_A_juz2ebfG8_0(.dout(w_dff_A_2rnCKYeo7_0),.din(w_dff_A_juz2ebfG8_0),.clk(gclk));
	jdff dff_A_WHW0Pjbg7_0(.dout(w_dff_A_juz2ebfG8_0),.din(w_dff_A_WHW0Pjbg7_0),.clk(gclk));
	jdff dff_A_qV0J2Adw5_0(.dout(w_dff_A_WHW0Pjbg7_0),.din(w_dff_A_qV0J2Adw5_0),.clk(gclk));
	jdff dff_A_B7YqcfYP3_0(.dout(w_dff_A_qV0J2Adw5_0),.din(w_dff_A_B7YqcfYP3_0),.clk(gclk));
	jdff dff_A_VEujq0b56_1(.dout(w_n633_0[1]),.din(w_dff_A_VEujq0b56_1),.clk(gclk));
	jdff dff_B_OJfJScoz0_1(.din(n557),.dout(w_dff_B_OJfJScoz0_1),.clk(gclk));
	jdff dff_B_joy5pEiW6_1(.din(w_dff_B_OJfJScoz0_1),.dout(w_dff_B_joy5pEiW6_1),.clk(gclk));
	jdff dff_B_3DAOgqIv0_1(.din(w_dff_B_joy5pEiW6_1),.dout(w_dff_B_3DAOgqIv0_1),.clk(gclk));
	jdff dff_B_YBPywL6Y7_1(.din(w_dff_B_3DAOgqIv0_1),.dout(w_dff_B_YBPywL6Y7_1),.clk(gclk));
	jdff dff_B_EnBhvp3R5_1(.din(w_dff_B_YBPywL6Y7_1),.dout(w_dff_B_EnBhvp3R5_1),.clk(gclk));
	jdff dff_B_C964AZh05_1(.din(w_dff_B_EnBhvp3R5_1),.dout(w_dff_B_C964AZh05_1),.clk(gclk));
	jdff dff_B_hL3MVVJ48_1(.din(w_dff_B_C964AZh05_1),.dout(w_dff_B_hL3MVVJ48_1),.clk(gclk));
	jdff dff_B_UVMXs8U84_1(.din(w_dff_B_hL3MVVJ48_1),.dout(w_dff_B_UVMXs8U84_1),.clk(gclk));
	jdff dff_B_NilN6uRf9_1(.din(w_dff_B_UVMXs8U84_1),.dout(w_dff_B_NilN6uRf9_1),.clk(gclk));
	jdff dff_B_lrcE3rTO2_1(.din(w_dff_B_NilN6uRf9_1),.dout(w_dff_B_lrcE3rTO2_1),.clk(gclk));
	jdff dff_B_OcEBqq0a0_1(.din(w_dff_B_lrcE3rTO2_1),.dout(w_dff_B_OcEBqq0a0_1),.clk(gclk));
	jdff dff_B_rGFg2lv54_1(.din(w_dff_B_OcEBqq0a0_1),.dout(w_dff_B_rGFg2lv54_1),.clk(gclk));
	jdff dff_B_C98GHJac1_1(.din(w_dff_B_rGFg2lv54_1),.dout(w_dff_B_C98GHJac1_1),.clk(gclk));
	jdff dff_B_SRazcrER0_1(.din(w_dff_B_C98GHJac1_1),.dout(w_dff_B_SRazcrER0_1),.clk(gclk));
	jdff dff_B_B5Mhl2501_1(.din(w_dff_B_SRazcrER0_1),.dout(w_dff_B_B5Mhl2501_1),.clk(gclk));
	jdff dff_B_XCivvqJI1_1(.din(w_dff_B_B5Mhl2501_1),.dout(w_dff_B_XCivvqJI1_1),.clk(gclk));
	jdff dff_B_yzdRFT6X2_1(.din(w_dff_B_XCivvqJI1_1),.dout(w_dff_B_yzdRFT6X2_1),.clk(gclk));
	jdff dff_B_8XdL0IZy2_1(.din(w_dff_B_yzdRFT6X2_1),.dout(w_dff_B_8XdL0IZy2_1),.clk(gclk));
	jdff dff_B_rd4GnHpT2_1(.din(w_dff_B_8XdL0IZy2_1),.dout(w_dff_B_rd4GnHpT2_1),.clk(gclk));
	jdff dff_B_GAred9fU3_1(.din(w_dff_B_rd4GnHpT2_1),.dout(w_dff_B_GAred9fU3_1),.clk(gclk));
	jdff dff_B_ScXbBoIh5_1(.din(w_dff_B_GAred9fU3_1),.dout(w_dff_B_ScXbBoIh5_1),.clk(gclk));
	jdff dff_B_CEfqVYqh2_1(.din(w_dff_B_ScXbBoIh5_1),.dout(w_dff_B_CEfqVYqh2_1),.clk(gclk));
	jdff dff_B_u2mvNLNg6_1(.din(w_dff_B_CEfqVYqh2_1),.dout(w_dff_B_u2mvNLNg6_1),.clk(gclk));
	jdff dff_B_rdiRkRYn2_1(.din(w_dff_B_u2mvNLNg6_1),.dout(w_dff_B_rdiRkRYn2_1),.clk(gclk));
	jdff dff_B_LFjcMIIR9_1(.din(w_dff_B_rdiRkRYn2_1),.dout(w_dff_B_LFjcMIIR9_1),.clk(gclk));
	jdff dff_B_qrdrG9vH9_1(.din(w_dff_B_LFjcMIIR9_1),.dout(w_dff_B_qrdrG9vH9_1),.clk(gclk));
	jdff dff_B_hA2MNSKg1_1(.din(w_dff_B_qrdrG9vH9_1),.dout(w_dff_B_hA2MNSKg1_1),.clk(gclk));
	jdff dff_B_paERo2nw3_1(.din(w_dff_B_hA2MNSKg1_1),.dout(w_dff_B_paERo2nw3_1),.clk(gclk));
	jdff dff_B_50uwYBqb8_1(.din(w_dff_B_paERo2nw3_1),.dout(w_dff_B_50uwYBqb8_1),.clk(gclk));
	jdff dff_B_5bCHPLMj2_1(.din(w_dff_B_50uwYBqb8_1),.dout(w_dff_B_5bCHPLMj2_1),.clk(gclk));
	jdff dff_B_roJGW98C6_1(.din(w_dff_B_5bCHPLMj2_1),.dout(w_dff_B_roJGW98C6_1),.clk(gclk));
	jdff dff_B_SiMRqYSP0_1(.din(n553),.dout(w_dff_B_SiMRqYSP0_1),.clk(gclk));
	jdff dff_A_TfVGntJz7_0(.dout(w_n471_0[0]),.din(w_dff_A_TfVGntJz7_0),.clk(gclk));
	jdff dff_A_cb660BSI2_0(.dout(w_dff_A_TfVGntJz7_0),.din(w_dff_A_cb660BSI2_0),.clk(gclk));
	jdff dff_A_wsJKOmr06_0(.dout(w_dff_A_cb660BSI2_0),.din(w_dff_A_wsJKOmr06_0),.clk(gclk));
	jdff dff_A_OarxkGwb9_0(.dout(w_dff_A_wsJKOmr06_0),.din(w_dff_A_OarxkGwb9_0),.clk(gclk));
	jdff dff_A_MJEZPcC65_0(.dout(w_dff_A_OarxkGwb9_0),.din(w_dff_A_MJEZPcC65_0),.clk(gclk));
	jdff dff_A_jE0oqnOV1_0(.dout(w_dff_A_MJEZPcC65_0),.din(w_dff_A_jE0oqnOV1_0),.clk(gclk));
	jdff dff_A_NgTIrXBe0_0(.dout(w_dff_A_jE0oqnOV1_0),.din(w_dff_A_NgTIrXBe0_0),.clk(gclk));
	jdff dff_A_WOEk7TDI7_0(.dout(w_dff_A_NgTIrXBe0_0),.din(w_dff_A_WOEk7TDI7_0),.clk(gclk));
	jdff dff_A_ZwcKZ1oD1_0(.dout(w_dff_A_WOEk7TDI7_0),.din(w_dff_A_ZwcKZ1oD1_0),.clk(gclk));
	jdff dff_A_1KYVI5oj1_0(.dout(w_dff_A_ZwcKZ1oD1_0),.din(w_dff_A_1KYVI5oj1_0),.clk(gclk));
	jdff dff_A_q3sEG3wu9_0(.dout(w_dff_A_1KYVI5oj1_0),.din(w_dff_A_q3sEG3wu9_0),.clk(gclk));
	jdff dff_A_FECjCLY76_0(.dout(w_dff_A_q3sEG3wu9_0),.din(w_dff_A_FECjCLY76_0),.clk(gclk));
	jdff dff_A_VVB6rwfg3_0(.dout(w_dff_A_FECjCLY76_0),.din(w_dff_A_VVB6rwfg3_0),.clk(gclk));
	jdff dff_A_RgaFQV2E3_0(.dout(w_dff_A_VVB6rwfg3_0),.din(w_dff_A_RgaFQV2E3_0),.clk(gclk));
	jdff dff_A_V0BsDLNf3_0(.dout(w_dff_A_RgaFQV2E3_0),.din(w_dff_A_V0BsDLNf3_0),.clk(gclk));
	jdff dff_A_PHckNOMP3_0(.dout(w_dff_A_V0BsDLNf3_0),.din(w_dff_A_PHckNOMP3_0),.clk(gclk));
	jdff dff_A_796bviRN4_0(.dout(w_dff_A_PHckNOMP3_0),.din(w_dff_A_796bviRN4_0),.clk(gclk));
	jdff dff_A_ha7oxkKw9_0(.dout(w_dff_A_796bviRN4_0),.din(w_dff_A_ha7oxkKw9_0),.clk(gclk));
	jdff dff_A_fJfDg6ol7_0(.dout(w_dff_A_ha7oxkKw9_0),.din(w_dff_A_fJfDg6ol7_0),.clk(gclk));
	jdff dff_A_m6oYLtBJ3_0(.dout(w_dff_A_fJfDg6ol7_0),.din(w_dff_A_m6oYLtBJ3_0),.clk(gclk));
	jdff dff_A_atYdfedi5_0(.dout(w_dff_A_m6oYLtBJ3_0),.din(w_dff_A_atYdfedi5_0),.clk(gclk));
	jdff dff_A_iQ4PABgr5_0(.dout(w_dff_A_atYdfedi5_0),.din(w_dff_A_iQ4PABgr5_0),.clk(gclk));
	jdff dff_A_jrbihYW94_0(.dout(w_dff_A_iQ4PABgr5_0),.din(w_dff_A_jrbihYW94_0),.clk(gclk));
	jdff dff_A_VNghTjrV4_0(.dout(w_dff_A_jrbihYW94_0),.din(w_dff_A_VNghTjrV4_0),.clk(gclk));
	jdff dff_A_uMVnOkCX0_0(.dout(w_dff_A_VNghTjrV4_0),.din(w_dff_A_uMVnOkCX0_0),.clk(gclk));
	jdff dff_A_T6f6kl7h9_0(.dout(w_dff_A_uMVnOkCX0_0),.din(w_dff_A_T6f6kl7h9_0),.clk(gclk));
	jdff dff_A_G7SOcXHi1_0(.dout(w_dff_A_T6f6kl7h9_0),.din(w_dff_A_G7SOcXHi1_0),.clk(gclk));
	jdff dff_A_Wpkx4X1d1_0(.dout(w_dff_A_G7SOcXHi1_0),.din(w_dff_A_Wpkx4X1d1_0),.clk(gclk));
	jdff dff_A_wON9vDc00_0(.dout(w_dff_A_Wpkx4X1d1_0),.din(w_dff_A_wON9vDc00_0),.clk(gclk));
	jdff dff_A_pKmVraOf9_0(.dout(w_dff_A_wON9vDc00_0),.din(w_dff_A_pKmVraOf9_0),.clk(gclk));
	jdff dff_A_ecIxD9CN5_0(.dout(w_dff_A_pKmVraOf9_0),.din(w_dff_A_ecIxD9CN5_0),.clk(gclk));
	jdff dff_A_3ewd5nH07_0(.dout(w_dff_A_ecIxD9CN5_0),.din(w_dff_A_3ewd5nH07_0),.clk(gclk));
	jdff dff_A_iE7a1jkd8_1(.dout(w_n547_0[1]),.din(w_dff_A_iE7a1jkd8_1),.clk(gclk));
	jdff dff_B_SHXBKMV59_1(.din(n478),.dout(w_dff_B_SHXBKMV59_1),.clk(gclk));
	jdff dff_B_KUkdH2Ek2_1(.din(w_dff_B_SHXBKMV59_1),.dout(w_dff_B_KUkdH2Ek2_1),.clk(gclk));
	jdff dff_B_jSczWzAw1_1(.din(w_dff_B_KUkdH2Ek2_1),.dout(w_dff_B_jSczWzAw1_1),.clk(gclk));
	jdff dff_B_e7XHIZua4_1(.din(w_dff_B_jSczWzAw1_1),.dout(w_dff_B_e7XHIZua4_1),.clk(gclk));
	jdff dff_B_oeIymY4S7_1(.din(w_dff_B_e7XHIZua4_1),.dout(w_dff_B_oeIymY4S7_1),.clk(gclk));
	jdff dff_B_qvpSU4mg0_1(.din(w_dff_B_oeIymY4S7_1),.dout(w_dff_B_qvpSU4mg0_1),.clk(gclk));
	jdff dff_B_YCHuXqUO9_1(.din(w_dff_B_qvpSU4mg0_1),.dout(w_dff_B_YCHuXqUO9_1),.clk(gclk));
	jdff dff_B_Dlg3pveE8_1(.din(w_dff_B_YCHuXqUO9_1),.dout(w_dff_B_Dlg3pveE8_1),.clk(gclk));
	jdff dff_B_Y6Ph1RZp8_1(.din(w_dff_B_Dlg3pveE8_1),.dout(w_dff_B_Y6Ph1RZp8_1),.clk(gclk));
	jdff dff_B_7bbmL7kk0_1(.din(w_dff_B_Y6Ph1RZp8_1),.dout(w_dff_B_7bbmL7kk0_1),.clk(gclk));
	jdff dff_B_82q5e7au1_1(.din(w_dff_B_7bbmL7kk0_1),.dout(w_dff_B_82q5e7au1_1),.clk(gclk));
	jdff dff_B_0NGNH7rw5_1(.din(w_dff_B_82q5e7au1_1),.dout(w_dff_B_0NGNH7rw5_1),.clk(gclk));
	jdff dff_B_sb2qU9gS3_1(.din(w_dff_B_0NGNH7rw5_1),.dout(w_dff_B_sb2qU9gS3_1),.clk(gclk));
	jdff dff_B_ca2ebekT1_1(.din(w_dff_B_sb2qU9gS3_1),.dout(w_dff_B_ca2ebekT1_1),.clk(gclk));
	jdff dff_B_WtQrNsz83_1(.din(w_dff_B_ca2ebekT1_1),.dout(w_dff_B_WtQrNsz83_1),.clk(gclk));
	jdff dff_B_DXAwpNOh7_1(.din(w_dff_B_WtQrNsz83_1),.dout(w_dff_B_DXAwpNOh7_1),.clk(gclk));
	jdff dff_B_LYqCxyIv1_1(.din(w_dff_B_DXAwpNOh7_1),.dout(w_dff_B_LYqCxyIv1_1),.clk(gclk));
	jdff dff_B_0xslFham9_1(.din(w_dff_B_LYqCxyIv1_1),.dout(w_dff_B_0xslFham9_1),.clk(gclk));
	jdff dff_B_BPA1vyTb9_1(.din(w_dff_B_0xslFham9_1),.dout(w_dff_B_BPA1vyTb9_1),.clk(gclk));
	jdff dff_B_SKAL9PmQ0_1(.din(w_dff_B_BPA1vyTb9_1),.dout(w_dff_B_SKAL9PmQ0_1),.clk(gclk));
	jdff dff_B_2CZqNCrI2_1(.din(w_dff_B_SKAL9PmQ0_1),.dout(w_dff_B_2CZqNCrI2_1),.clk(gclk));
	jdff dff_B_12IyrgCF9_1(.din(w_dff_B_2CZqNCrI2_1),.dout(w_dff_B_12IyrgCF9_1),.clk(gclk));
	jdff dff_B_cs4ZLtuU8_1(.din(w_dff_B_12IyrgCF9_1),.dout(w_dff_B_cs4ZLtuU8_1),.clk(gclk));
	jdff dff_B_ZgCJ9OWN6_1(.din(w_dff_B_cs4ZLtuU8_1),.dout(w_dff_B_ZgCJ9OWN6_1),.clk(gclk));
	jdff dff_B_oXIPgjlU4_1(.din(w_dff_B_ZgCJ9OWN6_1),.dout(w_dff_B_oXIPgjlU4_1),.clk(gclk));
	jdff dff_B_rRGPNQS83_1(.din(w_dff_B_oXIPgjlU4_1),.dout(w_dff_B_rRGPNQS83_1),.clk(gclk));
	jdff dff_B_SGNPYJPA7_1(.din(w_dff_B_rRGPNQS83_1),.dout(w_dff_B_SGNPYJPA7_1),.clk(gclk));
	jdff dff_B_KRdIAUVx8_1(.din(w_dff_B_SGNPYJPA7_1),.dout(w_dff_B_KRdIAUVx8_1),.clk(gclk));
	jdff dff_B_AYmBTs4D8_1(.din(n474),.dout(w_dff_B_AYmBTs4D8_1),.clk(gclk));
	jdff dff_A_MsZw9eL00_0(.dout(w_n399_0[0]),.din(w_dff_A_MsZw9eL00_0),.clk(gclk));
	jdff dff_A_S9aX8mER4_0(.dout(w_dff_A_MsZw9eL00_0),.din(w_dff_A_S9aX8mER4_0),.clk(gclk));
	jdff dff_A_mhz7RFrQ9_0(.dout(w_dff_A_S9aX8mER4_0),.din(w_dff_A_mhz7RFrQ9_0),.clk(gclk));
	jdff dff_A_eOpELvlj0_0(.dout(w_dff_A_mhz7RFrQ9_0),.din(w_dff_A_eOpELvlj0_0),.clk(gclk));
	jdff dff_A_fncPAUtS0_0(.dout(w_dff_A_eOpELvlj0_0),.din(w_dff_A_fncPAUtS0_0),.clk(gclk));
	jdff dff_A_7CsSnZhN1_0(.dout(w_dff_A_fncPAUtS0_0),.din(w_dff_A_7CsSnZhN1_0),.clk(gclk));
	jdff dff_A_nWL8wY5z6_0(.dout(w_dff_A_7CsSnZhN1_0),.din(w_dff_A_nWL8wY5z6_0),.clk(gclk));
	jdff dff_A_XvWY4woz7_0(.dout(w_dff_A_nWL8wY5z6_0),.din(w_dff_A_XvWY4woz7_0),.clk(gclk));
	jdff dff_A_V5Yvs6a06_0(.dout(w_dff_A_XvWY4woz7_0),.din(w_dff_A_V5Yvs6a06_0),.clk(gclk));
	jdff dff_A_aJmCCQqP3_0(.dout(w_dff_A_V5Yvs6a06_0),.din(w_dff_A_aJmCCQqP3_0),.clk(gclk));
	jdff dff_A_AF8J90EB8_0(.dout(w_dff_A_aJmCCQqP3_0),.din(w_dff_A_AF8J90EB8_0),.clk(gclk));
	jdff dff_A_DrVyjojO3_0(.dout(w_dff_A_AF8J90EB8_0),.din(w_dff_A_DrVyjojO3_0),.clk(gclk));
	jdff dff_A_SZnW5jyC4_0(.dout(w_dff_A_DrVyjojO3_0),.din(w_dff_A_SZnW5jyC4_0),.clk(gclk));
	jdff dff_A_Hput9qZ54_0(.dout(w_dff_A_SZnW5jyC4_0),.din(w_dff_A_Hput9qZ54_0),.clk(gclk));
	jdff dff_A_DCA00LGs1_0(.dout(w_dff_A_Hput9qZ54_0),.din(w_dff_A_DCA00LGs1_0),.clk(gclk));
	jdff dff_A_ifkn9wne2_0(.dout(w_dff_A_DCA00LGs1_0),.din(w_dff_A_ifkn9wne2_0),.clk(gclk));
	jdff dff_A_rnapPzg55_0(.dout(w_dff_A_ifkn9wne2_0),.din(w_dff_A_rnapPzg55_0),.clk(gclk));
	jdff dff_A_mbKfXsXN0_0(.dout(w_dff_A_rnapPzg55_0),.din(w_dff_A_mbKfXsXN0_0),.clk(gclk));
	jdff dff_A_LDsKEhHh2_0(.dout(w_dff_A_mbKfXsXN0_0),.din(w_dff_A_LDsKEhHh2_0),.clk(gclk));
	jdff dff_A_zzaQnLjh7_0(.dout(w_dff_A_LDsKEhHh2_0),.din(w_dff_A_zzaQnLjh7_0),.clk(gclk));
	jdff dff_A_ZYQKrtTy8_0(.dout(w_dff_A_zzaQnLjh7_0),.din(w_dff_A_ZYQKrtTy8_0),.clk(gclk));
	jdff dff_A_XRk1wtlT0_0(.dout(w_dff_A_ZYQKrtTy8_0),.din(w_dff_A_XRk1wtlT0_0),.clk(gclk));
	jdff dff_A_RXDF3Jaj7_0(.dout(w_dff_A_XRk1wtlT0_0),.din(w_dff_A_RXDF3Jaj7_0),.clk(gclk));
	jdff dff_A_KkKty4pY6_0(.dout(w_dff_A_RXDF3Jaj7_0),.din(w_dff_A_KkKty4pY6_0),.clk(gclk));
	jdff dff_A_PW1IC8L31_0(.dout(w_dff_A_KkKty4pY6_0),.din(w_dff_A_PW1IC8L31_0),.clk(gclk));
	jdff dff_A_Pi5vtkFv3_0(.dout(w_dff_A_PW1IC8L31_0),.din(w_dff_A_Pi5vtkFv3_0),.clk(gclk));
	jdff dff_A_Cq33Vq0E9_0(.dout(w_dff_A_Pi5vtkFv3_0),.din(w_dff_A_Cq33Vq0E9_0),.clk(gclk));
	jdff dff_A_PPh594NK9_0(.dout(w_dff_A_Cq33Vq0E9_0),.din(w_dff_A_PPh594NK9_0),.clk(gclk));
	jdff dff_A_pnmCap4I7_0(.dout(w_dff_A_PPh594NK9_0),.din(w_dff_A_pnmCap4I7_0),.clk(gclk));
	jdff dff_A_JKTgIqrw1_1(.dout(w_n468_0[1]),.din(w_dff_A_JKTgIqrw1_1),.clk(gclk));
	jdff dff_B_8tM1nnR65_1(.din(n406),.dout(w_dff_B_8tM1nnR65_1),.clk(gclk));
	jdff dff_B_expECOPx3_1(.din(w_dff_B_8tM1nnR65_1),.dout(w_dff_B_expECOPx3_1),.clk(gclk));
	jdff dff_B_dGtnS4Ig9_1(.din(w_dff_B_expECOPx3_1),.dout(w_dff_B_dGtnS4Ig9_1),.clk(gclk));
	jdff dff_B_WZX3xJTF5_1(.din(w_dff_B_dGtnS4Ig9_1),.dout(w_dff_B_WZX3xJTF5_1),.clk(gclk));
	jdff dff_B_AKeJy0H19_1(.din(w_dff_B_WZX3xJTF5_1),.dout(w_dff_B_AKeJy0H19_1),.clk(gclk));
	jdff dff_B_0L4ounem3_1(.din(w_dff_B_AKeJy0H19_1),.dout(w_dff_B_0L4ounem3_1),.clk(gclk));
	jdff dff_B_qNH2hI4z3_1(.din(w_dff_B_0L4ounem3_1),.dout(w_dff_B_qNH2hI4z3_1),.clk(gclk));
	jdff dff_B_qBuVi36n1_1(.din(w_dff_B_qNH2hI4z3_1),.dout(w_dff_B_qBuVi36n1_1),.clk(gclk));
	jdff dff_B_mWMq3leq7_1(.din(w_dff_B_qBuVi36n1_1),.dout(w_dff_B_mWMq3leq7_1),.clk(gclk));
	jdff dff_B_JVaVW0bZ0_1(.din(w_dff_B_mWMq3leq7_1),.dout(w_dff_B_JVaVW0bZ0_1),.clk(gclk));
	jdff dff_B_wTJPMqFx7_1(.din(w_dff_B_JVaVW0bZ0_1),.dout(w_dff_B_wTJPMqFx7_1),.clk(gclk));
	jdff dff_B_7NRFgcrF2_1(.din(w_dff_B_wTJPMqFx7_1),.dout(w_dff_B_7NRFgcrF2_1),.clk(gclk));
	jdff dff_B_ZrTlRkxe0_1(.din(w_dff_B_7NRFgcrF2_1),.dout(w_dff_B_ZrTlRkxe0_1),.clk(gclk));
	jdff dff_B_fE8E5YMv9_1(.din(w_dff_B_ZrTlRkxe0_1),.dout(w_dff_B_fE8E5YMv9_1),.clk(gclk));
	jdff dff_B_jxd1XQPV9_1(.din(w_dff_B_fE8E5YMv9_1),.dout(w_dff_B_jxd1XQPV9_1),.clk(gclk));
	jdff dff_B_xdaXtQ4L7_1(.din(w_dff_B_jxd1XQPV9_1),.dout(w_dff_B_xdaXtQ4L7_1),.clk(gclk));
	jdff dff_B_BSxM0G4N5_1(.din(w_dff_B_xdaXtQ4L7_1),.dout(w_dff_B_BSxM0G4N5_1),.clk(gclk));
	jdff dff_B_vos2f6LB7_1(.din(w_dff_B_BSxM0G4N5_1),.dout(w_dff_B_vos2f6LB7_1),.clk(gclk));
	jdff dff_B_OpBSgC7a5_1(.din(w_dff_B_vos2f6LB7_1),.dout(w_dff_B_OpBSgC7a5_1),.clk(gclk));
	jdff dff_B_gZP13rbP1_1(.din(w_dff_B_OpBSgC7a5_1),.dout(w_dff_B_gZP13rbP1_1),.clk(gclk));
	jdff dff_B_UNG6iTBt4_1(.din(w_dff_B_gZP13rbP1_1),.dout(w_dff_B_UNG6iTBt4_1),.clk(gclk));
	jdff dff_B_Ct6SxtCE4_1(.din(w_dff_B_UNG6iTBt4_1),.dout(w_dff_B_Ct6SxtCE4_1),.clk(gclk));
	jdff dff_B_v9jalWxg6_1(.din(w_dff_B_Ct6SxtCE4_1),.dout(w_dff_B_v9jalWxg6_1),.clk(gclk));
	jdff dff_B_qUdHmnrM6_1(.din(w_dff_B_v9jalWxg6_1),.dout(w_dff_B_qUdHmnrM6_1),.clk(gclk));
	jdff dff_B_5LHCkCEA4_1(.din(w_dff_B_qUdHmnrM6_1),.dout(w_dff_B_5LHCkCEA4_1),.clk(gclk));
	jdff dff_B_G8Fc5G387_1(.din(n402),.dout(w_dff_B_G8Fc5G387_1),.clk(gclk));
	jdff dff_A_o0IdYv1X2_0(.dout(w_n335_0[0]),.din(w_dff_A_o0IdYv1X2_0),.clk(gclk));
	jdff dff_A_41d7oRsv5_0(.dout(w_dff_A_o0IdYv1X2_0),.din(w_dff_A_41d7oRsv5_0),.clk(gclk));
	jdff dff_A_YlLJb8ht6_0(.dout(w_dff_A_41d7oRsv5_0),.din(w_dff_A_YlLJb8ht6_0),.clk(gclk));
	jdff dff_A_fFEXxIo36_0(.dout(w_dff_A_YlLJb8ht6_0),.din(w_dff_A_fFEXxIo36_0),.clk(gclk));
	jdff dff_A_f37HOTUI0_0(.dout(w_dff_A_fFEXxIo36_0),.din(w_dff_A_f37HOTUI0_0),.clk(gclk));
	jdff dff_A_hB5TfpfO7_0(.dout(w_dff_A_f37HOTUI0_0),.din(w_dff_A_hB5TfpfO7_0),.clk(gclk));
	jdff dff_A_U0MRCOKw7_0(.dout(w_dff_A_hB5TfpfO7_0),.din(w_dff_A_U0MRCOKw7_0),.clk(gclk));
	jdff dff_A_a49wjfty6_0(.dout(w_dff_A_U0MRCOKw7_0),.din(w_dff_A_a49wjfty6_0),.clk(gclk));
	jdff dff_A_ZDdbKGXc0_0(.dout(w_dff_A_a49wjfty6_0),.din(w_dff_A_ZDdbKGXc0_0),.clk(gclk));
	jdff dff_A_pJp30FFi1_0(.dout(w_dff_A_ZDdbKGXc0_0),.din(w_dff_A_pJp30FFi1_0),.clk(gclk));
	jdff dff_A_tfuJ1Uo45_0(.dout(w_dff_A_pJp30FFi1_0),.din(w_dff_A_tfuJ1Uo45_0),.clk(gclk));
	jdff dff_A_l6USH4Oj8_0(.dout(w_dff_A_tfuJ1Uo45_0),.din(w_dff_A_l6USH4Oj8_0),.clk(gclk));
	jdff dff_A_ic76lS2t2_0(.dout(w_dff_A_l6USH4Oj8_0),.din(w_dff_A_ic76lS2t2_0),.clk(gclk));
	jdff dff_A_PLur7qtH0_0(.dout(w_dff_A_ic76lS2t2_0),.din(w_dff_A_PLur7qtH0_0),.clk(gclk));
	jdff dff_A_gN9wrMQX9_0(.dout(w_dff_A_PLur7qtH0_0),.din(w_dff_A_gN9wrMQX9_0),.clk(gclk));
	jdff dff_A_dnwwuee63_0(.dout(w_dff_A_gN9wrMQX9_0),.din(w_dff_A_dnwwuee63_0),.clk(gclk));
	jdff dff_A_cpotRyDG6_0(.dout(w_dff_A_dnwwuee63_0),.din(w_dff_A_cpotRyDG6_0),.clk(gclk));
	jdff dff_A_zRKrqAC58_0(.dout(w_dff_A_cpotRyDG6_0),.din(w_dff_A_zRKrqAC58_0),.clk(gclk));
	jdff dff_A_0tUIz5fG9_0(.dout(w_dff_A_zRKrqAC58_0),.din(w_dff_A_0tUIz5fG9_0),.clk(gclk));
	jdff dff_A_Mtw9PDXq7_0(.dout(w_dff_A_0tUIz5fG9_0),.din(w_dff_A_Mtw9PDXq7_0),.clk(gclk));
	jdff dff_A_9KWDlbn13_0(.dout(w_dff_A_Mtw9PDXq7_0),.din(w_dff_A_9KWDlbn13_0),.clk(gclk));
	jdff dff_A_A5AhjcCE6_0(.dout(w_dff_A_9KWDlbn13_0),.din(w_dff_A_A5AhjcCE6_0),.clk(gclk));
	jdff dff_A_diIkPePp5_0(.dout(w_dff_A_A5AhjcCE6_0),.din(w_dff_A_diIkPePp5_0),.clk(gclk));
	jdff dff_A_Wb3qlsaT2_0(.dout(w_dff_A_diIkPePp5_0),.din(w_dff_A_Wb3qlsaT2_0),.clk(gclk));
	jdff dff_A_RNesFzje9_0(.dout(w_dff_A_Wb3qlsaT2_0),.din(w_dff_A_RNesFzje9_0),.clk(gclk));
	jdff dff_A_PEKduRXH7_0(.dout(w_dff_A_RNesFzje9_0),.din(w_dff_A_PEKduRXH7_0),.clk(gclk));
	jdff dff_A_3CJq4Na68_1(.dout(w_n396_0[1]),.din(w_dff_A_3CJq4Na68_1),.clk(gclk));
	jdff dff_B_VrrZgCmV6_1(.din(n342),.dout(w_dff_B_VrrZgCmV6_1),.clk(gclk));
	jdff dff_B_mDYnHiFa7_1(.din(w_dff_B_VrrZgCmV6_1),.dout(w_dff_B_mDYnHiFa7_1),.clk(gclk));
	jdff dff_B_xohbVPTK9_1(.din(w_dff_B_mDYnHiFa7_1),.dout(w_dff_B_xohbVPTK9_1),.clk(gclk));
	jdff dff_B_o7QfjYe32_1(.din(w_dff_B_xohbVPTK9_1),.dout(w_dff_B_o7QfjYe32_1),.clk(gclk));
	jdff dff_B_VbRvaQ872_1(.din(w_dff_B_o7QfjYe32_1),.dout(w_dff_B_VbRvaQ872_1),.clk(gclk));
	jdff dff_B_MjjmvXDn0_1(.din(w_dff_B_VbRvaQ872_1),.dout(w_dff_B_MjjmvXDn0_1),.clk(gclk));
	jdff dff_B_e3iHZ4Zg2_1(.din(w_dff_B_MjjmvXDn0_1),.dout(w_dff_B_e3iHZ4Zg2_1),.clk(gclk));
	jdff dff_B_USundpJN9_1(.din(w_dff_B_e3iHZ4Zg2_1),.dout(w_dff_B_USundpJN9_1),.clk(gclk));
	jdff dff_B_2WSZ42HF4_1(.din(w_dff_B_USundpJN9_1),.dout(w_dff_B_2WSZ42HF4_1),.clk(gclk));
	jdff dff_B_GaVuTz163_1(.din(w_dff_B_2WSZ42HF4_1),.dout(w_dff_B_GaVuTz163_1),.clk(gclk));
	jdff dff_B_llBApBEW4_1(.din(w_dff_B_GaVuTz163_1),.dout(w_dff_B_llBApBEW4_1),.clk(gclk));
	jdff dff_B_BNOntGvT6_1(.din(w_dff_B_llBApBEW4_1),.dout(w_dff_B_BNOntGvT6_1),.clk(gclk));
	jdff dff_B_aExB5qGr1_1(.din(w_dff_B_BNOntGvT6_1),.dout(w_dff_B_aExB5qGr1_1),.clk(gclk));
	jdff dff_B_Lwq3ozrN1_1(.din(w_dff_B_aExB5qGr1_1),.dout(w_dff_B_Lwq3ozrN1_1),.clk(gclk));
	jdff dff_B_diMeUvQl1_1(.din(w_dff_B_Lwq3ozrN1_1),.dout(w_dff_B_diMeUvQl1_1),.clk(gclk));
	jdff dff_B_CJGC58Sf0_1(.din(w_dff_B_diMeUvQl1_1),.dout(w_dff_B_CJGC58Sf0_1),.clk(gclk));
	jdff dff_B_feXLolQg1_1(.din(w_dff_B_CJGC58Sf0_1),.dout(w_dff_B_feXLolQg1_1),.clk(gclk));
	jdff dff_B_Cy9ppjHU9_1(.din(w_dff_B_feXLolQg1_1),.dout(w_dff_B_Cy9ppjHU9_1),.clk(gclk));
	jdff dff_B_Boy1qROf5_1(.din(w_dff_B_Cy9ppjHU9_1),.dout(w_dff_B_Boy1qROf5_1),.clk(gclk));
	jdff dff_B_aerMXmxU8_1(.din(w_dff_B_Boy1qROf5_1),.dout(w_dff_B_aerMXmxU8_1),.clk(gclk));
	jdff dff_B_zDDQiLEs8_1(.din(w_dff_B_aerMXmxU8_1),.dout(w_dff_B_zDDQiLEs8_1),.clk(gclk));
	jdff dff_B_qyHnPJs31_1(.din(w_dff_B_zDDQiLEs8_1),.dout(w_dff_B_qyHnPJs31_1),.clk(gclk));
	jdff dff_B_ibo5FJdy2_1(.din(n338),.dout(w_dff_B_ibo5FJdy2_1),.clk(gclk));
	jdff dff_A_MTGAcOxS8_0(.dout(w_n277_0[0]),.din(w_dff_A_MTGAcOxS8_0),.clk(gclk));
	jdff dff_A_Dqlxau3C9_0(.dout(w_dff_A_MTGAcOxS8_0),.din(w_dff_A_Dqlxau3C9_0),.clk(gclk));
	jdff dff_A_ZyvMiqwv7_0(.dout(w_dff_A_Dqlxau3C9_0),.din(w_dff_A_ZyvMiqwv7_0),.clk(gclk));
	jdff dff_A_AF5Godks4_0(.dout(w_dff_A_ZyvMiqwv7_0),.din(w_dff_A_AF5Godks4_0),.clk(gclk));
	jdff dff_A_t49iNQX13_0(.dout(w_dff_A_AF5Godks4_0),.din(w_dff_A_t49iNQX13_0),.clk(gclk));
	jdff dff_A_Vou0topv5_0(.dout(w_dff_A_t49iNQX13_0),.din(w_dff_A_Vou0topv5_0),.clk(gclk));
	jdff dff_A_8V5MMddR3_0(.dout(w_dff_A_Vou0topv5_0),.din(w_dff_A_8V5MMddR3_0),.clk(gclk));
	jdff dff_A_NDxk09Lm9_0(.dout(w_dff_A_8V5MMddR3_0),.din(w_dff_A_NDxk09Lm9_0),.clk(gclk));
	jdff dff_A_3bqzTno87_0(.dout(w_dff_A_NDxk09Lm9_0),.din(w_dff_A_3bqzTno87_0),.clk(gclk));
	jdff dff_A_u740gv2z5_0(.dout(w_dff_A_3bqzTno87_0),.din(w_dff_A_u740gv2z5_0),.clk(gclk));
	jdff dff_A_JUX6K2h81_0(.dout(w_dff_A_u740gv2z5_0),.din(w_dff_A_JUX6K2h81_0),.clk(gclk));
	jdff dff_A_qiFtbCbr5_0(.dout(w_dff_A_JUX6K2h81_0),.din(w_dff_A_qiFtbCbr5_0),.clk(gclk));
	jdff dff_A_MPJ39nPw9_0(.dout(w_dff_A_qiFtbCbr5_0),.din(w_dff_A_MPJ39nPw9_0),.clk(gclk));
	jdff dff_A_1uLbwkqc1_0(.dout(w_dff_A_MPJ39nPw9_0),.din(w_dff_A_1uLbwkqc1_0),.clk(gclk));
	jdff dff_A_cnvrGUbq3_0(.dout(w_dff_A_1uLbwkqc1_0),.din(w_dff_A_cnvrGUbq3_0),.clk(gclk));
	jdff dff_A_66IuD3qm1_0(.dout(w_dff_A_cnvrGUbq3_0),.din(w_dff_A_66IuD3qm1_0),.clk(gclk));
	jdff dff_A_vcHSnjrt3_0(.dout(w_dff_A_66IuD3qm1_0),.din(w_dff_A_vcHSnjrt3_0),.clk(gclk));
	jdff dff_A_Xol5qGsh0_0(.dout(w_dff_A_vcHSnjrt3_0),.din(w_dff_A_Xol5qGsh0_0),.clk(gclk));
	jdff dff_A_Rs6q3HyB2_0(.dout(w_dff_A_Xol5qGsh0_0),.din(w_dff_A_Rs6q3HyB2_0),.clk(gclk));
	jdff dff_A_7h3mI36C1_0(.dout(w_dff_A_Rs6q3HyB2_0),.din(w_dff_A_7h3mI36C1_0),.clk(gclk));
	jdff dff_A_GJNayBME6_0(.dout(w_dff_A_7h3mI36C1_0),.din(w_dff_A_GJNayBME6_0),.clk(gclk));
	jdff dff_A_vIIkb0HD7_0(.dout(w_dff_A_GJNayBME6_0),.din(w_dff_A_vIIkb0HD7_0),.clk(gclk));
	jdff dff_A_WJYgSSeq1_0(.dout(w_dff_A_vIIkb0HD7_0),.din(w_dff_A_WJYgSSeq1_0),.clk(gclk));
	jdff dff_A_VidqzFNW6_1(.dout(w_n332_0[1]),.din(w_dff_A_VidqzFNW6_1),.clk(gclk));
	jdff dff_B_f0vyNdGs6_1(.din(n284),.dout(w_dff_B_f0vyNdGs6_1),.clk(gclk));
	jdff dff_B_JFgCKWVc8_1(.din(w_dff_B_f0vyNdGs6_1),.dout(w_dff_B_JFgCKWVc8_1),.clk(gclk));
	jdff dff_B_MvkArjkZ4_1(.din(w_dff_B_JFgCKWVc8_1),.dout(w_dff_B_MvkArjkZ4_1),.clk(gclk));
	jdff dff_B_QfVfJSCB6_1(.din(w_dff_B_MvkArjkZ4_1),.dout(w_dff_B_QfVfJSCB6_1),.clk(gclk));
	jdff dff_B_aWIF8es22_1(.din(w_dff_B_QfVfJSCB6_1),.dout(w_dff_B_aWIF8es22_1),.clk(gclk));
	jdff dff_B_ay02jxqo6_1(.din(w_dff_B_aWIF8es22_1),.dout(w_dff_B_ay02jxqo6_1),.clk(gclk));
	jdff dff_B_dLsXYE3Z5_1(.din(w_dff_B_ay02jxqo6_1),.dout(w_dff_B_dLsXYE3Z5_1),.clk(gclk));
	jdff dff_B_zgHnO0sP7_1(.din(w_dff_B_dLsXYE3Z5_1),.dout(w_dff_B_zgHnO0sP7_1),.clk(gclk));
	jdff dff_B_n4NTiLWU4_1(.din(w_dff_B_zgHnO0sP7_1),.dout(w_dff_B_n4NTiLWU4_1),.clk(gclk));
	jdff dff_B_9DF1XkZM9_1(.din(w_dff_B_n4NTiLWU4_1),.dout(w_dff_B_9DF1XkZM9_1),.clk(gclk));
	jdff dff_B_6VFewGtb1_1(.din(w_dff_B_9DF1XkZM9_1),.dout(w_dff_B_6VFewGtb1_1),.clk(gclk));
	jdff dff_B_XspO4uMb3_1(.din(w_dff_B_6VFewGtb1_1),.dout(w_dff_B_XspO4uMb3_1),.clk(gclk));
	jdff dff_B_qyoP1Ca73_1(.din(w_dff_B_XspO4uMb3_1),.dout(w_dff_B_qyoP1Ca73_1),.clk(gclk));
	jdff dff_B_6tf9Yp4V8_1(.din(w_dff_B_qyoP1Ca73_1),.dout(w_dff_B_6tf9Yp4V8_1),.clk(gclk));
	jdff dff_B_qeR3ms464_1(.din(w_dff_B_6tf9Yp4V8_1),.dout(w_dff_B_qeR3ms464_1),.clk(gclk));
	jdff dff_B_Z2TokshB1_1(.din(w_dff_B_qeR3ms464_1),.dout(w_dff_B_Z2TokshB1_1),.clk(gclk));
	jdff dff_B_k3rcn5xi0_1(.din(w_dff_B_Z2TokshB1_1),.dout(w_dff_B_k3rcn5xi0_1),.clk(gclk));
	jdff dff_B_YQ8XFpW90_1(.din(w_dff_B_k3rcn5xi0_1),.dout(w_dff_B_YQ8XFpW90_1),.clk(gclk));
	jdff dff_B_qwvf0gmh5_1(.din(w_dff_B_YQ8XFpW90_1),.dout(w_dff_B_qwvf0gmh5_1),.clk(gclk));
	jdff dff_B_zvFQplgs5_1(.din(n280),.dout(w_dff_B_zvFQplgs5_1),.clk(gclk));
	jdff dff_A_DxyQf3yv1_0(.dout(w_n226_0[0]),.din(w_dff_A_DxyQf3yv1_0),.clk(gclk));
	jdff dff_A_WGEYsVGX8_0(.dout(w_dff_A_DxyQf3yv1_0),.din(w_dff_A_WGEYsVGX8_0),.clk(gclk));
	jdff dff_A_McTraJS24_0(.dout(w_dff_A_WGEYsVGX8_0),.din(w_dff_A_McTraJS24_0),.clk(gclk));
	jdff dff_A_sBNH4PME7_0(.dout(w_dff_A_McTraJS24_0),.din(w_dff_A_sBNH4PME7_0),.clk(gclk));
	jdff dff_A_sLsyXSrp2_0(.dout(w_dff_A_sBNH4PME7_0),.din(w_dff_A_sLsyXSrp2_0),.clk(gclk));
	jdff dff_A_a2o728ux5_0(.dout(w_dff_A_sLsyXSrp2_0),.din(w_dff_A_a2o728ux5_0),.clk(gclk));
	jdff dff_A_uf9mn53k1_0(.dout(w_dff_A_a2o728ux5_0),.din(w_dff_A_uf9mn53k1_0),.clk(gclk));
	jdff dff_A_mRaioLGc7_0(.dout(w_dff_A_uf9mn53k1_0),.din(w_dff_A_mRaioLGc7_0),.clk(gclk));
	jdff dff_A_YpSBvYFC1_0(.dout(w_dff_A_mRaioLGc7_0),.din(w_dff_A_YpSBvYFC1_0),.clk(gclk));
	jdff dff_A_aAAURnAq8_0(.dout(w_dff_A_YpSBvYFC1_0),.din(w_dff_A_aAAURnAq8_0),.clk(gclk));
	jdff dff_A_XCPjNbdl0_0(.dout(w_dff_A_aAAURnAq8_0),.din(w_dff_A_XCPjNbdl0_0),.clk(gclk));
	jdff dff_A_gOyCnO5A1_0(.dout(w_dff_A_XCPjNbdl0_0),.din(w_dff_A_gOyCnO5A1_0),.clk(gclk));
	jdff dff_A_4L6LIz1d6_0(.dout(w_dff_A_gOyCnO5A1_0),.din(w_dff_A_4L6LIz1d6_0),.clk(gclk));
	jdff dff_A_PoUpHa9o8_0(.dout(w_dff_A_4L6LIz1d6_0),.din(w_dff_A_PoUpHa9o8_0),.clk(gclk));
	jdff dff_A_MtB7Ibou8_0(.dout(w_dff_A_PoUpHa9o8_0),.din(w_dff_A_MtB7Ibou8_0),.clk(gclk));
	jdff dff_A_slhcY3sp1_0(.dout(w_dff_A_MtB7Ibou8_0),.din(w_dff_A_slhcY3sp1_0),.clk(gclk));
	jdff dff_A_8hqnuJXv0_0(.dout(w_dff_A_slhcY3sp1_0),.din(w_dff_A_8hqnuJXv0_0),.clk(gclk));
	jdff dff_A_teltklyC2_0(.dout(w_dff_A_8hqnuJXv0_0),.din(w_dff_A_teltklyC2_0),.clk(gclk));
	jdff dff_A_Nzpx970u6_0(.dout(w_dff_A_teltklyC2_0),.din(w_dff_A_Nzpx970u6_0),.clk(gclk));
	jdff dff_A_r7OMeDpp7_0(.dout(w_dff_A_Nzpx970u6_0),.din(w_dff_A_r7OMeDpp7_0),.clk(gclk));
	jdff dff_A_uk6LQE8m1_1(.dout(w_n274_0[1]),.din(w_dff_A_uk6LQE8m1_1),.clk(gclk));
	jdff dff_B_GXZScAZ97_1(.din(n233),.dout(w_dff_B_GXZScAZ97_1),.clk(gclk));
	jdff dff_B_sNXOD5Te5_1(.din(w_dff_B_GXZScAZ97_1),.dout(w_dff_B_sNXOD5Te5_1),.clk(gclk));
	jdff dff_B_mosPq6Iw7_1(.din(w_dff_B_sNXOD5Te5_1),.dout(w_dff_B_mosPq6Iw7_1),.clk(gclk));
	jdff dff_B_DmqVEt9h3_1(.din(w_dff_B_mosPq6Iw7_1),.dout(w_dff_B_DmqVEt9h3_1),.clk(gclk));
	jdff dff_B_WqQ9P0BI9_1(.din(w_dff_B_DmqVEt9h3_1),.dout(w_dff_B_WqQ9P0BI9_1),.clk(gclk));
	jdff dff_B_tYMvDHjF9_1(.din(w_dff_B_WqQ9P0BI9_1),.dout(w_dff_B_tYMvDHjF9_1),.clk(gclk));
	jdff dff_B_mYvwLHIE3_1(.din(w_dff_B_tYMvDHjF9_1),.dout(w_dff_B_mYvwLHIE3_1),.clk(gclk));
	jdff dff_B_jy7V7kH94_1(.din(w_dff_B_mYvwLHIE3_1),.dout(w_dff_B_jy7V7kH94_1),.clk(gclk));
	jdff dff_B_nYSoaTrs1_1(.din(w_dff_B_jy7V7kH94_1),.dout(w_dff_B_nYSoaTrs1_1),.clk(gclk));
	jdff dff_B_I7oXqdZX9_1(.din(w_dff_B_nYSoaTrs1_1),.dout(w_dff_B_I7oXqdZX9_1),.clk(gclk));
	jdff dff_B_xjCOxvEJ8_1(.din(w_dff_B_I7oXqdZX9_1),.dout(w_dff_B_xjCOxvEJ8_1),.clk(gclk));
	jdff dff_B_A0SwQJBz2_1(.din(w_dff_B_xjCOxvEJ8_1),.dout(w_dff_B_A0SwQJBz2_1),.clk(gclk));
	jdff dff_B_9neIFpWk8_1(.din(w_dff_B_A0SwQJBz2_1),.dout(w_dff_B_9neIFpWk8_1),.clk(gclk));
	jdff dff_B_9kGByPrb8_1(.din(w_dff_B_9neIFpWk8_1),.dout(w_dff_B_9kGByPrb8_1),.clk(gclk));
	jdff dff_B_KNAIm56a4_1(.din(w_dff_B_9kGByPrb8_1),.dout(w_dff_B_KNAIm56a4_1),.clk(gclk));
	jdff dff_B_zlTyNM2h9_1(.din(w_dff_B_KNAIm56a4_1),.dout(w_dff_B_zlTyNM2h9_1),.clk(gclk));
	jdff dff_B_0vmM2Dpk6_1(.din(n229),.dout(w_dff_B_0vmM2Dpk6_1),.clk(gclk));
	jdff dff_A_RQoc8dDu3_0(.dout(w_n183_0[0]),.din(w_dff_A_RQoc8dDu3_0),.clk(gclk));
	jdff dff_A_3UYvoCjL7_0(.dout(w_dff_A_RQoc8dDu3_0),.din(w_dff_A_3UYvoCjL7_0),.clk(gclk));
	jdff dff_A_JYJIqle31_0(.dout(w_dff_A_3UYvoCjL7_0),.din(w_dff_A_JYJIqle31_0),.clk(gclk));
	jdff dff_A_Zam404ga7_0(.dout(w_dff_A_JYJIqle31_0),.din(w_dff_A_Zam404ga7_0),.clk(gclk));
	jdff dff_A_xpaw3GIc3_0(.dout(w_dff_A_Zam404ga7_0),.din(w_dff_A_xpaw3GIc3_0),.clk(gclk));
	jdff dff_A_qtTvdTNd6_0(.dout(w_dff_A_xpaw3GIc3_0),.din(w_dff_A_qtTvdTNd6_0),.clk(gclk));
	jdff dff_A_b0WoWlA55_0(.dout(w_dff_A_qtTvdTNd6_0),.din(w_dff_A_b0WoWlA55_0),.clk(gclk));
	jdff dff_A_ipcMJtvZ3_0(.dout(w_dff_A_b0WoWlA55_0),.din(w_dff_A_ipcMJtvZ3_0),.clk(gclk));
	jdff dff_A_lllFJPyA9_0(.dout(w_dff_A_ipcMJtvZ3_0),.din(w_dff_A_lllFJPyA9_0),.clk(gclk));
	jdff dff_A_NIXy8Lja8_0(.dout(w_dff_A_lllFJPyA9_0),.din(w_dff_A_NIXy8Lja8_0),.clk(gclk));
	jdff dff_A_XuSvxjEP4_0(.dout(w_dff_A_NIXy8Lja8_0),.din(w_dff_A_XuSvxjEP4_0),.clk(gclk));
	jdff dff_A_evmWHlwv5_0(.dout(w_dff_A_XuSvxjEP4_0),.din(w_dff_A_evmWHlwv5_0),.clk(gclk));
	jdff dff_A_sRkSva2B6_0(.dout(w_dff_A_evmWHlwv5_0),.din(w_dff_A_sRkSva2B6_0),.clk(gclk));
	jdff dff_A_s7YYj71d7_0(.dout(w_dff_A_sRkSva2B6_0),.din(w_dff_A_s7YYj71d7_0),.clk(gclk));
	jdff dff_A_eI7iRPhF5_0(.dout(w_dff_A_s7YYj71d7_0),.din(w_dff_A_eI7iRPhF5_0),.clk(gclk));
	jdff dff_A_CKC3Yn8f7_0(.dout(w_dff_A_eI7iRPhF5_0),.din(w_dff_A_CKC3Yn8f7_0),.clk(gclk));
	jdff dff_A_VZPaFjUV4_0(.dout(w_dff_A_CKC3Yn8f7_0),.din(w_dff_A_VZPaFjUV4_0),.clk(gclk));
	jdff dff_A_jlM84O8q0_1(.dout(w_n223_0[1]),.din(w_dff_A_jlM84O8q0_1),.clk(gclk));
	jdff dff_B_zfuvNCQQ3_1(.din(n190),.dout(w_dff_B_zfuvNCQQ3_1),.clk(gclk));
	jdff dff_B_bpvSJBRK9_1(.din(w_dff_B_zfuvNCQQ3_1),.dout(w_dff_B_bpvSJBRK9_1),.clk(gclk));
	jdff dff_B_7oNspLiC5_1(.din(w_dff_B_bpvSJBRK9_1),.dout(w_dff_B_7oNspLiC5_1),.clk(gclk));
	jdff dff_B_EEACuwh76_1(.din(w_dff_B_7oNspLiC5_1),.dout(w_dff_B_EEACuwh76_1),.clk(gclk));
	jdff dff_B_Eu5engjA1_1(.din(w_dff_B_EEACuwh76_1),.dout(w_dff_B_Eu5engjA1_1),.clk(gclk));
	jdff dff_B_vQnexihB6_1(.din(w_dff_B_Eu5engjA1_1),.dout(w_dff_B_vQnexihB6_1),.clk(gclk));
	jdff dff_B_ILKNcXJf1_1(.din(w_dff_B_vQnexihB6_1),.dout(w_dff_B_ILKNcXJf1_1),.clk(gclk));
	jdff dff_B_nQtXH1jO1_1(.din(w_dff_B_ILKNcXJf1_1),.dout(w_dff_B_nQtXH1jO1_1),.clk(gclk));
	jdff dff_B_8ZTVRIvv5_1(.din(w_dff_B_nQtXH1jO1_1),.dout(w_dff_B_8ZTVRIvv5_1),.clk(gclk));
	jdff dff_B_xxPN8qXu7_1(.din(w_dff_B_8ZTVRIvv5_1),.dout(w_dff_B_xxPN8qXu7_1),.clk(gclk));
	jdff dff_B_MfqZ7y0c9_1(.din(w_dff_B_xxPN8qXu7_1),.dout(w_dff_B_MfqZ7y0c9_1),.clk(gclk));
	jdff dff_B_u1ziF5763_1(.din(w_dff_B_MfqZ7y0c9_1),.dout(w_dff_B_u1ziF5763_1),.clk(gclk));
	jdff dff_B_EHlu3dn94_1(.din(w_dff_B_u1ziF5763_1),.dout(w_dff_B_EHlu3dn94_1),.clk(gclk));
	jdff dff_B_NiuiUYAR7_1(.din(n186),.dout(w_dff_B_NiuiUYAR7_1),.clk(gclk));
	jdff dff_A_3morTeKC0_0(.dout(w_n145_0[0]),.din(w_dff_A_3morTeKC0_0),.clk(gclk));
	jdff dff_A_xHNVvKMT8_0(.dout(w_dff_A_3morTeKC0_0),.din(w_dff_A_xHNVvKMT8_0),.clk(gclk));
	jdff dff_A_nlkU3F5a8_0(.dout(w_dff_A_xHNVvKMT8_0),.din(w_dff_A_nlkU3F5a8_0),.clk(gclk));
	jdff dff_A_YRrVLZFO9_0(.dout(w_dff_A_nlkU3F5a8_0),.din(w_dff_A_YRrVLZFO9_0),.clk(gclk));
	jdff dff_A_aTQPuo2u3_0(.dout(w_dff_A_YRrVLZFO9_0),.din(w_dff_A_aTQPuo2u3_0),.clk(gclk));
	jdff dff_A_NBLHVlz99_0(.dout(w_dff_A_aTQPuo2u3_0),.din(w_dff_A_NBLHVlz99_0),.clk(gclk));
	jdff dff_A_svvjYLuG6_0(.dout(w_dff_A_NBLHVlz99_0),.din(w_dff_A_svvjYLuG6_0),.clk(gclk));
	jdff dff_A_8VOR3zpj2_0(.dout(w_dff_A_svvjYLuG6_0),.din(w_dff_A_8VOR3zpj2_0),.clk(gclk));
	jdff dff_A_ev0RHqGZ3_0(.dout(w_dff_A_8VOR3zpj2_0),.din(w_dff_A_ev0RHqGZ3_0),.clk(gclk));
	jdff dff_A_wHYSETMK7_0(.dout(w_dff_A_ev0RHqGZ3_0),.din(w_dff_A_wHYSETMK7_0),.clk(gclk));
	jdff dff_A_VCuonMYy9_0(.dout(w_dff_A_wHYSETMK7_0),.din(w_dff_A_VCuonMYy9_0),.clk(gclk));
	jdff dff_A_mvCLfD9x0_0(.dout(w_dff_A_VCuonMYy9_0),.din(w_dff_A_mvCLfD9x0_0),.clk(gclk));
	jdff dff_A_syDCTWfq5_0(.dout(w_dff_A_mvCLfD9x0_0),.din(w_dff_A_syDCTWfq5_0),.clk(gclk));
	jdff dff_A_zXoueFPQ6_0(.dout(w_dff_A_syDCTWfq5_0),.din(w_dff_A_zXoueFPQ6_0),.clk(gclk));
	jdff dff_A_t5eeBDnN5_1(.dout(w_n180_0[1]),.din(w_dff_A_t5eeBDnN5_1),.clk(gclk));
	jdff dff_B_9xiLlT4y2_1(.din(n152),.dout(w_dff_B_9xiLlT4y2_1),.clk(gclk));
	jdff dff_B_9KRAEmbh7_1(.din(w_dff_B_9xiLlT4y2_1),.dout(w_dff_B_9KRAEmbh7_1),.clk(gclk));
	jdff dff_B_ggZTS0gd1_1(.din(w_dff_B_9KRAEmbh7_1),.dout(w_dff_B_ggZTS0gd1_1),.clk(gclk));
	jdff dff_B_4LKlCLrA7_1(.din(w_dff_B_ggZTS0gd1_1),.dout(w_dff_B_4LKlCLrA7_1),.clk(gclk));
	jdff dff_B_2R25WAQK8_1(.din(w_dff_B_4LKlCLrA7_1),.dout(w_dff_B_2R25WAQK8_1),.clk(gclk));
	jdff dff_B_TppLyg4v4_1(.din(w_dff_B_2R25WAQK8_1),.dout(w_dff_B_TppLyg4v4_1),.clk(gclk));
	jdff dff_B_9nLxrKgD3_1(.din(w_dff_B_TppLyg4v4_1),.dout(w_dff_B_9nLxrKgD3_1),.clk(gclk));
	jdff dff_B_sNuIyDiq9_1(.din(w_dff_B_9nLxrKgD3_1),.dout(w_dff_B_sNuIyDiq9_1),.clk(gclk));
	jdff dff_B_M5kAxx6I7_1(.din(w_dff_B_sNuIyDiq9_1),.dout(w_dff_B_M5kAxx6I7_1),.clk(gclk));
	jdff dff_B_owl5xRXF4_1(.din(w_dff_B_M5kAxx6I7_1),.dout(w_dff_B_owl5xRXF4_1),.clk(gclk));
	jdff dff_B_2rxQ8rZv0_1(.din(n148),.dout(w_dff_B_2rxQ8rZv0_1),.clk(gclk));
	jdff dff_A_OpndN7z58_0(.dout(w_n110_0[0]),.din(w_dff_A_OpndN7z58_0),.clk(gclk));
	jdff dff_A_keAsB39M8_0(.dout(w_dff_A_OpndN7z58_0),.din(w_dff_A_keAsB39M8_0),.clk(gclk));
	jdff dff_A_gKgPIvD13_0(.dout(w_dff_A_keAsB39M8_0),.din(w_dff_A_gKgPIvD13_0),.clk(gclk));
	jdff dff_A_4cydyGjc7_0(.dout(w_dff_A_gKgPIvD13_0),.din(w_dff_A_4cydyGjc7_0),.clk(gclk));
	jdff dff_A_udABFOUe6_0(.dout(w_dff_A_4cydyGjc7_0),.din(w_dff_A_udABFOUe6_0),.clk(gclk));
	jdff dff_A_CCdgCSaS5_0(.dout(w_dff_A_udABFOUe6_0),.din(w_dff_A_CCdgCSaS5_0),.clk(gclk));
	jdff dff_A_YRpxcmXh3_0(.dout(w_dff_A_CCdgCSaS5_0),.din(w_dff_A_YRpxcmXh3_0),.clk(gclk));
	jdff dff_A_9KFj6Kic7_0(.dout(w_dff_A_YRpxcmXh3_0),.din(w_dff_A_9KFj6Kic7_0),.clk(gclk));
	jdff dff_A_fghwch2a5_0(.dout(w_dff_A_9KFj6Kic7_0),.din(w_dff_A_fghwch2a5_0),.clk(gclk));
	jdff dff_A_fswP8Brl5_0(.dout(w_dff_A_fghwch2a5_0),.din(w_dff_A_fswP8Brl5_0),.clk(gclk));
	jdff dff_A_1tP4Ojsj6_0(.dout(w_dff_A_fswP8Brl5_0),.din(w_dff_A_1tP4Ojsj6_0),.clk(gclk));
	jdff dff_A_16lnEayP7_1(.dout(w_n142_0[1]),.din(w_dff_A_16lnEayP7_1),.clk(gclk));
	jdff dff_B_ql0xxNOV8_1(.din(n117),.dout(w_dff_B_ql0xxNOV8_1),.clk(gclk));
	jdff dff_B_yEyi6Bcm2_1(.din(w_dff_B_ql0xxNOV8_1),.dout(w_dff_B_yEyi6Bcm2_1),.clk(gclk));
	jdff dff_B_dByFWDg89_1(.din(w_dff_B_yEyi6Bcm2_1),.dout(w_dff_B_dByFWDg89_1),.clk(gclk));
	jdff dff_B_3mjKI0g11_1(.din(w_dff_B_dByFWDg89_1),.dout(w_dff_B_3mjKI0g11_1),.clk(gclk));
	jdff dff_B_bu9REvml5_1(.din(w_dff_B_3mjKI0g11_1),.dout(w_dff_B_bu9REvml5_1),.clk(gclk));
	jdff dff_B_tmlWrp378_1(.din(w_dff_B_bu9REvml5_1),.dout(w_dff_B_tmlWrp378_1),.clk(gclk));
	jdff dff_B_WOKIVqPd1_1(.din(w_dff_B_tmlWrp378_1),.dout(w_dff_B_WOKIVqPd1_1),.clk(gclk));
	jdff dff_B_uBqySN0o4_1(.din(n113),.dout(w_dff_B_uBqySN0o4_1),.clk(gclk));
	jdff dff_A_6Iqt84Uz8_0(.dout(w_n89_0[0]),.din(w_dff_A_6Iqt84Uz8_0),.clk(gclk));
	jdff dff_A_lkj7oKoR0_0(.dout(w_dff_A_6Iqt84Uz8_0),.din(w_dff_A_lkj7oKoR0_0),.clk(gclk));
	jdff dff_A_RxECoBzC0_0(.dout(w_dff_A_lkj7oKoR0_0),.din(w_dff_A_RxECoBzC0_0),.clk(gclk));
	jdff dff_A_RJrAcvEy5_0(.dout(w_dff_A_RxECoBzC0_0),.din(w_dff_A_RJrAcvEy5_0),.clk(gclk));
	jdff dff_A_sMiz8vT45_0(.dout(w_dff_A_RJrAcvEy5_0),.din(w_dff_A_sMiz8vT45_0),.clk(gclk));
	jdff dff_A_zR5A5U2s7_0(.dout(w_dff_A_sMiz8vT45_0),.din(w_dff_A_zR5A5U2s7_0),.clk(gclk));
	jdff dff_A_ld20n9FH2_0(.dout(w_dff_A_zR5A5U2s7_0),.din(w_dff_A_ld20n9FH2_0),.clk(gclk));
	jdff dff_A_3bc51pMd5_0(.dout(w_dff_A_ld20n9FH2_0),.din(w_dff_A_3bc51pMd5_0),.clk(gclk));
	jdff dff_A_CTRaqL9B3_1(.dout(w_n107_0[1]),.din(w_dff_A_CTRaqL9B3_1),.clk(gclk));
	jdff dff_B_somNRr3K8_1(.din(n95),.dout(w_dff_B_somNRr3K8_1),.clk(gclk));
	jdff dff_B_3z8o40fg2_1(.din(w_dff_B_somNRr3K8_1),.dout(w_dff_B_3z8o40fg2_1),.clk(gclk));
	jdff dff_B_pGbrx3Wv3_1(.din(w_dff_B_3z8o40fg2_1),.dout(w_dff_B_pGbrx3Wv3_1),.clk(gclk));
	jdff dff_B_5uOOUoA52_1(.din(w_dff_B_pGbrx3Wv3_1),.dout(w_dff_B_5uOOUoA52_1),.clk(gclk));
	jdff dff_B_3MngmSLX7_1(.din(n91),.dout(w_dff_B_3MngmSLX7_1),.clk(gclk));
	jdff dff_B_8fabrxSB4_0(.din(n86),.dout(w_dff_B_8fabrxSB4_0),.clk(gclk));
	jdff dff_A_DuRvFlYK3_0(.dout(w_n72_0[0]),.din(w_dff_A_DuRvFlYK3_0),.clk(gclk));
	jdff dff_A_dzP8WDLp8_0(.dout(w_dff_A_DuRvFlYK3_0),.din(w_dff_A_dzP8WDLp8_0),.clk(gclk));
	jdff dff_A_XjuzOzbT6_0(.dout(w_dff_A_dzP8WDLp8_0),.din(w_dff_A_XjuzOzbT6_0),.clk(gclk));
	jdff dff_A_OePys8Kz6_0(.dout(w_dff_A_XjuzOzbT6_0),.din(w_dff_A_OePys8Kz6_0),.clk(gclk));
	jdff dff_A_yQlDCY0r9_0(.dout(w_dff_A_OePys8Kz6_0),.din(w_dff_A_yQlDCY0r9_0),.clk(gclk));
	jdff dff_A_jVSOrltG9_0(.dout(w_n70_0[0]),.din(w_dff_A_jVSOrltG9_0),.clk(gclk));
	jdff dff_A_qNtSau7H0_0(.dout(w_n69_0[0]),.din(w_dff_A_qNtSau7H0_0),.clk(gclk));
	jdff dff_A_Om9vCIER8_1(.dout(w_n1140_0[1]),.din(w_dff_A_Om9vCIER8_1),.clk(gclk));
	jdff dff_B_rxFTLE6m4_1(.din(n1040),.dout(w_dff_B_rxFTLE6m4_1),.clk(gclk));
	jdff dff_B_JeJeGQdS0_2(.din(n938),.dout(w_dff_B_JeJeGQdS0_2),.clk(gclk));
	jdff dff_B_eeC0TOx72_2(.din(w_dff_B_JeJeGQdS0_2),.dout(w_dff_B_eeC0TOx72_2),.clk(gclk));
	jdff dff_B_EqNcRvMn0_2(.din(w_dff_B_eeC0TOx72_2),.dout(w_dff_B_EqNcRvMn0_2),.clk(gclk));
	jdff dff_B_sd4iDbTu4_2(.din(w_dff_B_EqNcRvMn0_2),.dout(w_dff_B_sd4iDbTu4_2),.clk(gclk));
	jdff dff_B_4JqgDNrV1_2(.din(w_dff_B_sd4iDbTu4_2),.dout(w_dff_B_4JqgDNrV1_2),.clk(gclk));
	jdff dff_B_NhZ0ttCJ2_2(.din(w_dff_B_4JqgDNrV1_2),.dout(w_dff_B_NhZ0ttCJ2_2),.clk(gclk));
	jdff dff_B_u1Un5rHB2_2(.din(w_dff_B_NhZ0ttCJ2_2),.dout(w_dff_B_u1Un5rHB2_2),.clk(gclk));
	jdff dff_B_nI3qGxFd2_2(.din(w_dff_B_u1Un5rHB2_2),.dout(w_dff_B_nI3qGxFd2_2),.clk(gclk));
	jdff dff_B_HK9IvcZv5_2(.din(w_dff_B_nI3qGxFd2_2),.dout(w_dff_B_HK9IvcZv5_2),.clk(gclk));
	jdff dff_B_TY5MJ6X65_2(.din(w_dff_B_HK9IvcZv5_2),.dout(w_dff_B_TY5MJ6X65_2),.clk(gclk));
	jdff dff_B_KR9ir9qC3_2(.din(w_dff_B_TY5MJ6X65_2),.dout(w_dff_B_KR9ir9qC3_2),.clk(gclk));
	jdff dff_B_hwQDgPLZ3_2(.din(w_dff_B_KR9ir9qC3_2),.dout(w_dff_B_hwQDgPLZ3_2),.clk(gclk));
	jdff dff_B_KBRszzhj2_2(.din(w_dff_B_hwQDgPLZ3_2),.dout(w_dff_B_KBRszzhj2_2),.clk(gclk));
	jdff dff_B_4yDbemdy3_2(.din(w_dff_B_KBRszzhj2_2),.dout(w_dff_B_4yDbemdy3_2),.clk(gclk));
	jdff dff_B_dU7Dbcac8_2(.din(w_dff_B_4yDbemdy3_2),.dout(w_dff_B_dU7Dbcac8_2),.clk(gclk));
	jdff dff_B_aLJbCdnY1_2(.din(w_dff_B_dU7Dbcac8_2),.dout(w_dff_B_aLJbCdnY1_2),.clk(gclk));
	jdff dff_B_pZzzmzNk9_2(.din(w_dff_B_aLJbCdnY1_2),.dout(w_dff_B_pZzzmzNk9_2),.clk(gclk));
	jdff dff_B_jFmfJljb9_2(.din(w_dff_B_pZzzmzNk9_2),.dout(w_dff_B_jFmfJljb9_2),.clk(gclk));
	jdff dff_B_y0ggQzps5_2(.din(w_dff_B_jFmfJljb9_2),.dout(w_dff_B_y0ggQzps5_2),.clk(gclk));
	jdff dff_B_WLtX5I5J0_2(.din(w_dff_B_y0ggQzps5_2),.dout(w_dff_B_WLtX5I5J0_2),.clk(gclk));
	jdff dff_B_Px9ysO1c9_2(.din(w_dff_B_WLtX5I5J0_2),.dout(w_dff_B_Px9ysO1c9_2),.clk(gclk));
	jdff dff_B_2NAuces67_2(.din(w_dff_B_Px9ysO1c9_2),.dout(w_dff_B_2NAuces67_2),.clk(gclk));
	jdff dff_B_oUs2DGfX2_2(.din(w_dff_B_2NAuces67_2),.dout(w_dff_B_oUs2DGfX2_2),.clk(gclk));
	jdff dff_B_B2ynoS7N8_2(.din(w_dff_B_oUs2DGfX2_2),.dout(w_dff_B_B2ynoS7N8_2),.clk(gclk));
	jdff dff_B_Gv73NBPG9_2(.din(w_dff_B_B2ynoS7N8_2),.dout(w_dff_B_Gv73NBPG9_2),.clk(gclk));
	jdff dff_B_cGbWw0kq6_2(.din(w_dff_B_Gv73NBPG9_2),.dout(w_dff_B_cGbWw0kq6_2),.clk(gclk));
	jdff dff_B_hwS2Wrzm3_2(.din(w_dff_B_cGbWw0kq6_2),.dout(w_dff_B_hwS2Wrzm3_2),.clk(gclk));
	jdff dff_B_T0DtvykX4_2(.din(w_dff_B_hwS2Wrzm3_2),.dout(w_dff_B_T0DtvykX4_2),.clk(gclk));
	jdff dff_B_BLzPcQXz2_2(.din(w_dff_B_T0DtvykX4_2),.dout(w_dff_B_BLzPcQXz2_2),.clk(gclk));
	jdff dff_B_lCFiarFR4_2(.din(w_dff_B_BLzPcQXz2_2),.dout(w_dff_B_lCFiarFR4_2),.clk(gclk));
	jdff dff_B_EtTf68cC0_2(.din(w_dff_B_lCFiarFR4_2),.dout(w_dff_B_EtTf68cC0_2),.clk(gclk));
	jdff dff_B_O675cwWI4_2(.din(w_dff_B_EtTf68cC0_2),.dout(w_dff_B_O675cwWI4_2),.clk(gclk));
	jdff dff_B_w3paKbUS7_2(.din(w_dff_B_O675cwWI4_2),.dout(w_dff_B_w3paKbUS7_2),.clk(gclk));
	jdff dff_B_4e2zvKBd8_2(.din(w_dff_B_w3paKbUS7_2),.dout(w_dff_B_4e2zvKBd8_2),.clk(gclk));
	jdff dff_B_OsatqXEn2_2(.din(w_dff_B_4e2zvKBd8_2),.dout(w_dff_B_OsatqXEn2_2),.clk(gclk));
	jdff dff_B_6gcFq2qZ4_2(.din(w_dff_B_OsatqXEn2_2),.dout(w_dff_B_6gcFq2qZ4_2),.clk(gclk));
	jdff dff_B_43cWqXcJ9_2(.din(w_dff_B_6gcFq2qZ4_2),.dout(w_dff_B_43cWqXcJ9_2),.clk(gclk));
	jdff dff_B_XmiBbv9O8_2(.din(w_dff_B_43cWqXcJ9_2),.dout(w_dff_B_XmiBbv9O8_2),.clk(gclk));
	jdff dff_B_dbi9DG9r0_2(.din(w_dff_B_XmiBbv9O8_2),.dout(w_dff_B_dbi9DG9r0_2),.clk(gclk));
	jdff dff_B_cSCjdipF3_2(.din(w_dff_B_dbi9DG9r0_2),.dout(w_dff_B_cSCjdipF3_2),.clk(gclk));
	jdff dff_B_iQbbHtVj4_2(.din(w_dff_B_cSCjdipF3_2),.dout(w_dff_B_iQbbHtVj4_2),.clk(gclk));
	jdff dff_B_3iPC0LYk7_2(.din(w_dff_B_iQbbHtVj4_2),.dout(w_dff_B_3iPC0LYk7_2),.clk(gclk));
	jdff dff_B_xWKZTo7M7_2(.din(w_dff_B_3iPC0LYk7_2),.dout(w_dff_B_xWKZTo7M7_2),.clk(gclk));
	jdff dff_B_UgomcaYM9_2(.din(w_dff_B_xWKZTo7M7_2),.dout(w_dff_B_UgomcaYM9_2),.clk(gclk));
	jdff dff_A_IYu9QDqv2_0(.dout(w_n1034_0[0]),.din(w_dff_A_IYu9QDqv2_0),.clk(gclk));
	jdff dff_B_9J9G5dhP3_1(.din(n940),.dout(w_dff_B_9J9G5dhP3_1),.clk(gclk));
	jdff dff_B_TA4DWdGV8_2(.din(n835),.dout(w_dff_B_TA4DWdGV8_2),.clk(gclk));
	jdff dff_B_CLklGeY05_2(.din(w_dff_B_TA4DWdGV8_2),.dout(w_dff_B_CLklGeY05_2),.clk(gclk));
	jdff dff_B_QyBjJ8Vn9_2(.din(w_dff_B_CLklGeY05_2),.dout(w_dff_B_QyBjJ8Vn9_2),.clk(gclk));
	jdff dff_B_wTBYR0hu4_2(.din(w_dff_B_QyBjJ8Vn9_2),.dout(w_dff_B_wTBYR0hu4_2),.clk(gclk));
	jdff dff_B_TfGXVdAR0_2(.din(w_dff_B_wTBYR0hu4_2),.dout(w_dff_B_TfGXVdAR0_2),.clk(gclk));
	jdff dff_B_YJqXvrmm9_2(.din(w_dff_B_TfGXVdAR0_2),.dout(w_dff_B_YJqXvrmm9_2),.clk(gclk));
	jdff dff_B_k0IZG2Hc4_2(.din(w_dff_B_YJqXvrmm9_2),.dout(w_dff_B_k0IZG2Hc4_2),.clk(gclk));
	jdff dff_B_LMwbwHTU1_2(.din(w_dff_B_k0IZG2Hc4_2),.dout(w_dff_B_LMwbwHTU1_2),.clk(gclk));
	jdff dff_B_UGMUiXF57_2(.din(w_dff_B_LMwbwHTU1_2),.dout(w_dff_B_UGMUiXF57_2),.clk(gclk));
	jdff dff_B_AAgdIXzo4_2(.din(w_dff_B_UGMUiXF57_2),.dout(w_dff_B_AAgdIXzo4_2),.clk(gclk));
	jdff dff_B_wKENF1XL0_2(.din(w_dff_B_AAgdIXzo4_2),.dout(w_dff_B_wKENF1XL0_2),.clk(gclk));
	jdff dff_B_ZSJlHGs64_2(.din(w_dff_B_wKENF1XL0_2),.dout(w_dff_B_ZSJlHGs64_2),.clk(gclk));
	jdff dff_B_j4xQdnXq2_2(.din(w_dff_B_ZSJlHGs64_2),.dout(w_dff_B_j4xQdnXq2_2),.clk(gclk));
	jdff dff_B_kmFz5Dci2_2(.din(w_dff_B_j4xQdnXq2_2),.dout(w_dff_B_kmFz5Dci2_2),.clk(gclk));
	jdff dff_B_sucw9Ygt1_2(.din(w_dff_B_kmFz5Dci2_2),.dout(w_dff_B_sucw9Ygt1_2),.clk(gclk));
	jdff dff_B_IfUz4ndu2_2(.din(w_dff_B_sucw9Ygt1_2),.dout(w_dff_B_IfUz4ndu2_2),.clk(gclk));
	jdff dff_B_qVy19lph5_2(.din(w_dff_B_IfUz4ndu2_2),.dout(w_dff_B_qVy19lph5_2),.clk(gclk));
	jdff dff_B_zly0R7qp5_2(.din(w_dff_B_qVy19lph5_2),.dout(w_dff_B_zly0R7qp5_2),.clk(gclk));
	jdff dff_B_m7VVN3qx0_2(.din(w_dff_B_zly0R7qp5_2),.dout(w_dff_B_m7VVN3qx0_2),.clk(gclk));
	jdff dff_B_lywSVzBg9_2(.din(w_dff_B_m7VVN3qx0_2),.dout(w_dff_B_lywSVzBg9_2),.clk(gclk));
	jdff dff_B_SqR5ieOD9_2(.din(w_dff_B_lywSVzBg9_2),.dout(w_dff_B_SqR5ieOD9_2),.clk(gclk));
	jdff dff_B_qCfP3pXC0_2(.din(w_dff_B_SqR5ieOD9_2),.dout(w_dff_B_qCfP3pXC0_2),.clk(gclk));
	jdff dff_B_Ge9IynTe0_2(.din(w_dff_B_qCfP3pXC0_2),.dout(w_dff_B_Ge9IynTe0_2),.clk(gclk));
	jdff dff_B_pHsg5nmV1_2(.din(w_dff_B_Ge9IynTe0_2),.dout(w_dff_B_pHsg5nmV1_2),.clk(gclk));
	jdff dff_B_PouuHYAR1_2(.din(w_dff_B_pHsg5nmV1_2),.dout(w_dff_B_PouuHYAR1_2),.clk(gclk));
	jdff dff_B_2BO1y4Tc3_2(.din(w_dff_B_PouuHYAR1_2),.dout(w_dff_B_2BO1y4Tc3_2),.clk(gclk));
	jdff dff_B_hqLbpPmL6_2(.din(w_dff_B_2BO1y4Tc3_2),.dout(w_dff_B_hqLbpPmL6_2),.clk(gclk));
	jdff dff_B_hMjNrgmF9_2(.din(w_dff_B_hqLbpPmL6_2),.dout(w_dff_B_hMjNrgmF9_2),.clk(gclk));
	jdff dff_B_A23ukn8M6_2(.din(w_dff_B_hMjNrgmF9_2),.dout(w_dff_B_A23ukn8M6_2),.clk(gclk));
	jdff dff_B_NJyS9AiW9_2(.din(w_dff_B_A23ukn8M6_2),.dout(w_dff_B_NJyS9AiW9_2),.clk(gclk));
	jdff dff_B_QYCS95NF0_2(.din(w_dff_B_NJyS9AiW9_2),.dout(w_dff_B_QYCS95NF0_2),.clk(gclk));
	jdff dff_B_NdiLhKAS4_2(.din(w_dff_B_QYCS95NF0_2),.dout(w_dff_B_NdiLhKAS4_2),.clk(gclk));
	jdff dff_B_E70GJp9W9_2(.din(w_dff_B_NdiLhKAS4_2),.dout(w_dff_B_E70GJp9W9_2),.clk(gclk));
	jdff dff_B_rpYQZu1i4_2(.din(w_dff_B_E70GJp9W9_2),.dout(w_dff_B_rpYQZu1i4_2),.clk(gclk));
	jdff dff_B_ffCQGSql1_2(.din(w_dff_B_rpYQZu1i4_2),.dout(w_dff_B_ffCQGSql1_2),.clk(gclk));
	jdff dff_B_zNG8Nvgp8_2(.din(w_dff_B_ffCQGSql1_2),.dout(w_dff_B_zNG8Nvgp8_2),.clk(gclk));
	jdff dff_B_7pssP60b0_2(.din(w_dff_B_zNG8Nvgp8_2),.dout(w_dff_B_7pssP60b0_2),.clk(gclk));
	jdff dff_B_m2SC6Q7j9_2(.din(w_dff_B_7pssP60b0_2),.dout(w_dff_B_m2SC6Q7j9_2),.clk(gclk));
	jdff dff_B_yrfeAPaT5_2(.din(w_dff_B_m2SC6Q7j9_2),.dout(w_dff_B_yrfeAPaT5_2),.clk(gclk));
	jdff dff_B_JqAG9UCb9_2(.din(w_dff_B_yrfeAPaT5_2),.dout(w_dff_B_JqAG9UCb9_2),.clk(gclk));
	jdff dff_B_wO10LduC0_2(.din(w_dff_B_JqAG9UCb9_2),.dout(w_dff_B_wO10LduC0_2),.clk(gclk));
	jdff dff_A_Oj2QZeXD0_1(.dout(w_n929_0[1]),.din(w_dff_A_Oj2QZeXD0_1),.clk(gclk));
	jdff dff_B_V0dPnTPX0_1(.din(n841),.dout(w_dff_B_V0dPnTPX0_1),.clk(gclk));
	jdff dff_B_Ji9pX2ES4_1(.din(w_dff_B_V0dPnTPX0_1),.dout(w_dff_B_Ji9pX2ES4_1),.clk(gclk));
	jdff dff_B_0LUshjrx3_1(.din(w_dff_B_Ji9pX2ES4_1),.dout(w_dff_B_0LUshjrx3_1),.clk(gclk));
	jdff dff_B_T8rBcWFe3_1(.din(w_dff_B_0LUshjrx3_1),.dout(w_dff_B_T8rBcWFe3_1),.clk(gclk));
	jdff dff_B_HRWhvgFq4_1(.din(w_dff_B_T8rBcWFe3_1),.dout(w_dff_B_HRWhvgFq4_1),.clk(gclk));
	jdff dff_B_fd6niYRp1_1(.din(w_dff_B_HRWhvgFq4_1),.dout(w_dff_B_fd6niYRp1_1),.clk(gclk));
	jdff dff_B_xOW05q3B3_1(.din(w_dff_B_fd6niYRp1_1),.dout(w_dff_B_xOW05q3B3_1),.clk(gclk));
	jdff dff_B_DfFrf3BO6_1(.din(w_dff_B_xOW05q3B3_1),.dout(w_dff_B_DfFrf3BO6_1),.clk(gclk));
	jdff dff_B_FzFgK3iN0_1(.din(w_dff_B_DfFrf3BO6_1),.dout(w_dff_B_FzFgK3iN0_1),.clk(gclk));
	jdff dff_B_UbiBswyu7_1(.din(w_dff_B_FzFgK3iN0_1),.dout(w_dff_B_UbiBswyu7_1),.clk(gclk));
	jdff dff_B_DonOGi5j8_1(.din(w_dff_B_UbiBswyu7_1),.dout(w_dff_B_DonOGi5j8_1),.clk(gclk));
	jdff dff_B_DVlO2hi82_1(.din(w_dff_B_DonOGi5j8_1),.dout(w_dff_B_DVlO2hi82_1),.clk(gclk));
	jdff dff_B_sXy64Lbe9_1(.din(w_dff_B_DVlO2hi82_1),.dout(w_dff_B_sXy64Lbe9_1),.clk(gclk));
	jdff dff_B_yA48ylDb6_1(.din(w_dff_B_sXy64Lbe9_1),.dout(w_dff_B_yA48ylDb6_1),.clk(gclk));
	jdff dff_B_WqyKBDO63_1(.din(w_dff_B_yA48ylDb6_1),.dout(w_dff_B_WqyKBDO63_1),.clk(gclk));
	jdff dff_B_GEvAHh4Q7_1(.din(w_dff_B_WqyKBDO63_1),.dout(w_dff_B_GEvAHh4Q7_1),.clk(gclk));
	jdff dff_B_szhGWO7G2_1(.din(w_dff_B_GEvAHh4Q7_1),.dout(w_dff_B_szhGWO7G2_1),.clk(gclk));
	jdff dff_B_InNh9hGR3_1(.din(w_dff_B_szhGWO7G2_1),.dout(w_dff_B_InNh9hGR3_1),.clk(gclk));
	jdff dff_B_deOhBe0D3_1(.din(w_dff_B_InNh9hGR3_1),.dout(w_dff_B_deOhBe0D3_1),.clk(gclk));
	jdff dff_B_65BZeBJU7_1(.din(w_dff_B_deOhBe0D3_1),.dout(w_dff_B_65BZeBJU7_1),.clk(gclk));
	jdff dff_B_UTvbge8z0_1(.din(w_dff_B_65BZeBJU7_1),.dout(w_dff_B_UTvbge8z0_1),.clk(gclk));
	jdff dff_B_E2CMcfpL2_1(.din(w_dff_B_UTvbge8z0_1),.dout(w_dff_B_E2CMcfpL2_1),.clk(gclk));
	jdff dff_B_HoBcODdq0_1(.din(w_dff_B_E2CMcfpL2_1),.dout(w_dff_B_HoBcODdq0_1),.clk(gclk));
	jdff dff_B_xNpdHfJl8_1(.din(w_dff_B_HoBcODdq0_1),.dout(w_dff_B_xNpdHfJl8_1),.clk(gclk));
	jdff dff_B_SJcwfZQ30_1(.din(w_dff_B_xNpdHfJl8_1),.dout(w_dff_B_SJcwfZQ30_1),.clk(gclk));
	jdff dff_B_p86gTzkp7_1(.din(w_dff_B_SJcwfZQ30_1),.dout(w_dff_B_p86gTzkp7_1),.clk(gclk));
	jdff dff_B_wCHZHEGk1_1(.din(w_dff_B_p86gTzkp7_1),.dout(w_dff_B_wCHZHEGk1_1),.clk(gclk));
	jdff dff_B_TwMEC49E3_1(.din(w_dff_B_wCHZHEGk1_1),.dout(w_dff_B_TwMEC49E3_1),.clk(gclk));
	jdff dff_B_x1jdbZhI2_1(.din(w_dff_B_TwMEC49E3_1),.dout(w_dff_B_x1jdbZhI2_1),.clk(gclk));
	jdff dff_B_4wxA6eZn4_1(.din(w_dff_B_x1jdbZhI2_1),.dout(w_dff_B_4wxA6eZn4_1),.clk(gclk));
	jdff dff_B_pxfrCFT81_1(.din(w_dff_B_4wxA6eZn4_1),.dout(w_dff_B_pxfrCFT81_1),.clk(gclk));
	jdff dff_B_2zceQQ1i8_1(.din(w_dff_B_pxfrCFT81_1),.dout(w_dff_B_2zceQQ1i8_1),.clk(gclk));
	jdff dff_B_9Lah1VMm0_1(.din(w_dff_B_2zceQQ1i8_1),.dout(w_dff_B_9Lah1VMm0_1),.clk(gclk));
	jdff dff_B_ASKlD0uT5_1(.din(w_dff_B_9Lah1VMm0_1),.dout(w_dff_B_ASKlD0uT5_1),.clk(gclk));
	jdff dff_B_Cb7Bv95w9_1(.din(w_dff_B_ASKlD0uT5_1),.dout(w_dff_B_Cb7Bv95w9_1),.clk(gclk));
	jdff dff_B_xYDsoEwY9_1(.din(w_dff_B_Cb7Bv95w9_1),.dout(w_dff_B_xYDsoEwY9_1),.clk(gclk));
	jdff dff_B_sNHx9GFp7_1(.din(w_dff_B_xYDsoEwY9_1),.dout(w_dff_B_sNHx9GFp7_1),.clk(gclk));
	jdff dff_B_HWRDEJIq8_1(.din(n836),.dout(w_dff_B_HWRDEJIq8_1),.clk(gclk));
	jdff dff_A_8Ls6SQMY1_0(.dout(w_n735_0[0]),.din(w_dff_A_8Ls6SQMY1_0),.clk(gclk));
	jdff dff_A_jOD8LKnJ0_0(.dout(w_dff_A_8Ls6SQMY1_0),.din(w_dff_A_jOD8LKnJ0_0),.clk(gclk));
	jdff dff_A_xBUhKTzQ8_0(.dout(w_dff_A_jOD8LKnJ0_0),.din(w_dff_A_xBUhKTzQ8_0),.clk(gclk));
	jdff dff_A_ibTJclNI9_0(.dout(w_dff_A_xBUhKTzQ8_0),.din(w_dff_A_ibTJclNI9_0),.clk(gclk));
	jdff dff_A_CQtyuUFf5_0(.dout(w_dff_A_ibTJclNI9_0),.din(w_dff_A_CQtyuUFf5_0),.clk(gclk));
	jdff dff_A_k9P9u1CZ4_0(.dout(w_dff_A_CQtyuUFf5_0),.din(w_dff_A_k9P9u1CZ4_0),.clk(gclk));
	jdff dff_A_hnt2NgWO6_0(.dout(w_dff_A_k9P9u1CZ4_0),.din(w_dff_A_hnt2NgWO6_0),.clk(gclk));
	jdff dff_A_Sc62zVqh8_0(.dout(w_dff_A_hnt2NgWO6_0),.din(w_dff_A_Sc62zVqh8_0),.clk(gclk));
	jdff dff_A_3RBACpkU1_0(.dout(w_dff_A_Sc62zVqh8_0),.din(w_dff_A_3RBACpkU1_0),.clk(gclk));
	jdff dff_A_zP82B3G82_0(.dout(w_dff_A_3RBACpkU1_0),.din(w_dff_A_zP82B3G82_0),.clk(gclk));
	jdff dff_A_nIQTdYas5_0(.dout(w_dff_A_zP82B3G82_0),.din(w_dff_A_nIQTdYas5_0),.clk(gclk));
	jdff dff_A_kHK3pD0g0_0(.dout(w_dff_A_nIQTdYas5_0),.din(w_dff_A_kHK3pD0g0_0),.clk(gclk));
	jdff dff_A_LUAWhf7J4_0(.dout(w_dff_A_kHK3pD0g0_0),.din(w_dff_A_LUAWhf7J4_0),.clk(gclk));
	jdff dff_A_BTA1JJRI6_0(.dout(w_dff_A_LUAWhf7J4_0),.din(w_dff_A_BTA1JJRI6_0),.clk(gclk));
	jdff dff_A_NcKBC49r1_0(.dout(w_dff_A_BTA1JJRI6_0),.din(w_dff_A_NcKBC49r1_0),.clk(gclk));
	jdff dff_A_U36aJKzV6_0(.dout(w_dff_A_NcKBC49r1_0),.din(w_dff_A_U36aJKzV6_0),.clk(gclk));
	jdff dff_A_LGM7CuMA1_0(.dout(w_dff_A_U36aJKzV6_0),.din(w_dff_A_LGM7CuMA1_0),.clk(gclk));
	jdff dff_A_kX1Zn2fm0_0(.dout(w_dff_A_LGM7CuMA1_0),.din(w_dff_A_kX1Zn2fm0_0),.clk(gclk));
	jdff dff_A_z5RbAXbL2_0(.dout(w_dff_A_kX1Zn2fm0_0),.din(w_dff_A_z5RbAXbL2_0),.clk(gclk));
	jdff dff_A_9bIR5dQA7_0(.dout(w_dff_A_z5RbAXbL2_0),.din(w_dff_A_9bIR5dQA7_0),.clk(gclk));
	jdff dff_A_c3TXFA8I1_0(.dout(w_dff_A_9bIR5dQA7_0),.din(w_dff_A_c3TXFA8I1_0),.clk(gclk));
	jdff dff_A_fhBQCqvb4_0(.dout(w_dff_A_c3TXFA8I1_0),.din(w_dff_A_fhBQCqvb4_0),.clk(gclk));
	jdff dff_A_Gwt5aC6M9_0(.dout(w_dff_A_fhBQCqvb4_0),.din(w_dff_A_Gwt5aC6M9_0),.clk(gclk));
	jdff dff_A_un2q7DOg9_0(.dout(w_dff_A_Gwt5aC6M9_0),.din(w_dff_A_un2q7DOg9_0),.clk(gclk));
	jdff dff_A_Fw41wDSs7_0(.dout(w_dff_A_un2q7DOg9_0),.din(w_dff_A_Fw41wDSs7_0),.clk(gclk));
	jdff dff_A_gFL68rjQ3_0(.dout(w_dff_A_Fw41wDSs7_0),.din(w_dff_A_gFL68rjQ3_0),.clk(gclk));
	jdff dff_A_lJLprpNW4_0(.dout(w_dff_A_gFL68rjQ3_0),.din(w_dff_A_lJLprpNW4_0),.clk(gclk));
	jdff dff_A_9muuIYZa4_0(.dout(w_dff_A_lJLprpNW4_0),.din(w_dff_A_9muuIYZa4_0),.clk(gclk));
	jdff dff_A_XDBXbmDU9_0(.dout(w_dff_A_9muuIYZa4_0),.din(w_dff_A_XDBXbmDU9_0),.clk(gclk));
	jdff dff_A_zDsM3TAb9_0(.dout(w_dff_A_XDBXbmDU9_0),.din(w_dff_A_zDsM3TAb9_0),.clk(gclk));
	jdff dff_A_BtDzUKUL9_0(.dout(w_dff_A_zDsM3TAb9_0),.din(w_dff_A_BtDzUKUL9_0),.clk(gclk));
	jdff dff_A_W2ao1JDL2_0(.dout(w_dff_A_BtDzUKUL9_0),.din(w_dff_A_W2ao1JDL2_0),.clk(gclk));
	jdff dff_A_rZmwKjpC6_0(.dout(w_dff_A_W2ao1JDL2_0),.din(w_dff_A_rZmwKjpC6_0),.clk(gclk));
	jdff dff_A_FHz3OLs28_0(.dout(w_dff_A_rZmwKjpC6_0),.din(w_dff_A_FHz3OLs28_0),.clk(gclk));
	jdff dff_A_P6mwVooE5_0(.dout(w_dff_A_FHz3OLs28_0),.din(w_dff_A_P6mwVooE5_0),.clk(gclk));
	jdff dff_A_udAcokyh0_0(.dout(w_dff_A_P6mwVooE5_0),.din(w_dff_A_udAcokyh0_0),.clk(gclk));
	jdff dff_A_I6WCFdXQ7_0(.dout(w_dff_A_udAcokyh0_0),.din(w_dff_A_I6WCFdXQ7_0),.clk(gclk));
	jdff dff_A_Bb9hNL731_0(.dout(w_dff_A_I6WCFdXQ7_0),.din(w_dff_A_Bb9hNL731_0),.clk(gclk));
	jdff dff_A_ykRVGLmZ7_0(.dout(w_n823_0[0]),.din(w_dff_A_ykRVGLmZ7_0),.clk(gclk));
	jdff dff_B_3XNwPl930_1(.din(n737),.dout(w_dff_B_3XNwPl930_1),.clk(gclk));
	jdff dff_A_V0al9raf3_0(.dout(w_n642_0[0]),.din(w_dff_A_V0al9raf3_0),.clk(gclk));
	jdff dff_A_p7IMXphc6_0(.dout(w_dff_A_V0al9raf3_0),.din(w_dff_A_p7IMXphc6_0),.clk(gclk));
	jdff dff_A_b2PrGeK75_0(.dout(w_dff_A_p7IMXphc6_0),.din(w_dff_A_b2PrGeK75_0),.clk(gclk));
	jdff dff_A_ok5d407S7_0(.dout(w_dff_A_b2PrGeK75_0),.din(w_dff_A_ok5d407S7_0),.clk(gclk));
	jdff dff_A_5Zjy2mMT3_0(.dout(w_dff_A_ok5d407S7_0),.din(w_dff_A_5Zjy2mMT3_0),.clk(gclk));
	jdff dff_A_zHP9eEiN3_0(.dout(w_dff_A_5Zjy2mMT3_0),.din(w_dff_A_zHP9eEiN3_0),.clk(gclk));
	jdff dff_A_rUsxgoGb9_0(.dout(w_dff_A_zHP9eEiN3_0),.din(w_dff_A_rUsxgoGb9_0),.clk(gclk));
	jdff dff_A_UkVNKsnp5_0(.dout(w_dff_A_rUsxgoGb9_0),.din(w_dff_A_UkVNKsnp5_0),.clk(gclk));
	jdff dff_A_hzDffdzX1_0(.dout(w_dff_A_UkVNKsnp5_0),.din(w_dff_A_hzDffdzX1_0),.clk(gclk));
	jdff dff_A_WcQP0GVk7_0(.dout(w_dff_A_hzDffdzX1_0),.din(w_dff_A_WcQP0GVk7_0),.clk(gclk));
	jdff dff_A_kJPQVcKW1_0(.dout(w_dff_A_WcQP0GVk7_0),.din(w_dff_A_kJPQVcKW1_0),.clk(gclk));
	jdff dff_A_qhnUAuHw9_0(.dout(w_dff_A_kJPQVcKW1_0),.din(w_dff_A_qhnUAuHw9_0),.clk(gclk));
	jdff dff_A_oVsqIYz31_0(.dout(w_dff_A_qhnUAuHw9_0),.din(w_dff_A_oVsqIYz31_0),.clk(gclk));
	jdff dff_A_5tCBRLI28_0(.dout(w_dff_A_oVsqIYz31_0),.din(w_dff_A_5tCBRLI28_0),.clk(gclk));
	jdff dff_A_LNjcHkWh6_0(.dout(w_dff_A_5tCBRLI28_0),.din(w_dff_A_LNjcHkWh6_0),.clk(gclk));
	jdff dff_A_IM2OIQZE5_0(.dout(w_dff_A_LNjcHkWh6_0),.din(w_dff_A_IM2OIQZE5_0),.clk(gclk));
	jdff dff_A_F87PH2eY3_0(.dout(w_dff_A_IM2OIQZE5_0),.din(w_dff_A_F87PH2eY3_0),.clk(gclk));
	jdff dff_A_3WGIdDBq0_0(.dout(w_dff_A_F87PH2eY3_0),.din(w_dff_A_3WGIdDBq0_0),.clk(gclk));
	jdff dff_A_GXxg27Sd2_0(.dout(w_dff_A_3WGIdDBq0_0),.din(w_dff_A_GXxg27Sd2_0),.clk(gclk));
	jdff dff_A_swUgQyJJ3_0(.dout(w_dff_A_GXxg27Sd2_0),.din(w_dff_A_swUgQyJJ3_0),.clk(gclk));
	jdff dff_A_PP0Q3MYf6_0(.dout(w_dff_A_swUgQyJJ3_0),.din(w_dff_A_PP0Q3MYf6_0),.clk(gclk));
	jdff dff_A_lWUYQwJa5_0(.dout(w_dff_A_PP0Q3MYf6_0),.din(w_dff_A_lWUYQwJa5_0),.clk(gclk));
	jdff dff_A_XLGvzO3m2_0(.dout(w_dff_A_lWUYQwJa5_0),.din(w_dff_A_XLGvzO3m2_0),.clk(gclk));
	jdff dff_A_RCDgZQ4G3_0(.dout(w_dff_A_XLGvzO3m2_0),.din(w_dff_A_RCDgZQ4G3_0),.clk(gclk));
	jdff dff_A_T5knTiQt4_0(.dout(w_dff_A_RCDgZQ4G3_0),.din(w_dff_A_T5knTiQt4_0),.clk(gclk));
	jdff dff_A_2I5mb8x68_0(.dout(w_dff_A_T5knTiQt4_0),.din(w_dff_A_2I5mb8x68_0),.clk(gclk));
	jdff dff_A_x7BSejfI0_0(.dout(w_dff_A_2I5mb8x68_0),.din(w_dff_A_x7BSejfI0_0),.clk(gclk));
	jdff dff_A_6fOqBFAZ8_0(.dout(w_dff_A_x7BSejfI0_0),.din(w_dff_A_6fOqBFAZ8_0),.clk(gclk));
	jdff dff_A_SueV4pZG8_0(.dout(w_dff_A_6fOqBFAZ8_0),.din(w_dff_A_SueV4pZG8_0),.clk(gclk));
	jdff dff_A_a24faCMM5_0(.dout(w_dff_A_SueV4pZG8_0),.din(w_dff_A_a24faCMM5_0),.clk(gclk));
	jdff dff_A_oM5fdqOE2_0(.dout(w_dff_A_a24faCMM5_0),.din(w_dff_A_oM5fdqOE2_0),.clk(gclk));
	jdff dff_A_8D5ntETR4_0(.dout(w_dff_A_oM5fdqOE2_0),.din(w_dff_A_8D5ntETR4_0),.clk(gclk));
	jdff dff_A_MBWUmYwd6_0(.dout(w_dff_A_8D5ntETR4_0),.din(w_dff_A_MBWUmYwd6_0),.clk(gclk));
	jdff dff_A_s3ndbN176_0(.dout(w_dff_A_MBWUmYwd6_0),.din(w_dff_A_s3ndbN176_0),.clk(gclk));
	jdff dff_A_ovFp6XYL3_0(.dout(w_dff_A_s3ndbN176_0),.din(w_dff_A_ovFp6XYL3_0),.clk(gclk));
	jdff dff_A_hp903XOU7_0(.dout(w_n723_0[0]),.din(w_dff_A_hp903XOU7_0),.clk(gclk));
	jdff dff_B_wsW7Faqe1_1(.din(n644),.dout(w_dff_B_wsW7Faqe1_1),.clk(gclk));
	jdff dff_A_dd4K6fuO5_0(.dout(w_n556_0[0]),.din(w_dff_A_dd4K6fuO5_0),.clk(gclk));
	jdff dff_A_XpPiGr3x1_0(.dout(w_dff_A_dd4K6fuO5_0),.din(w_dff_A_XpPiGr3x1_0),.clk(gclk));
	jdff dff_A_yC0MeDY08_0(.dout(w_dff_A_XpPiGr3x1_0),.din(w_dff_A_yC0MeDY08_0),.clk(gclk));
	jdff dff_A_cGGgTJYQ8_0(.dout(w_dff_A_yC0MeDY08_0),.din(w_dff_A_cGGgTJYQ8_0),.clk(gclk));
	jdff dff_A_ukmfKaNG1_0(.dout(w_dff_A_cGGgTJYQ8_0),.din(w_dff_A_ukmfKaNG1_0),.clk(gclk));
	jdff dff_A_kV8hlzAE2_0(.dout(w_dff_A_ukmfKaNG1_0),.din(w_dff_A_kV8hlzAE2_0),.clk(gclk));
	jdff dff_A_8E0wrzOd7_0(.dout(w_dff_A_kV8hlzAE2_0),.din(w_dff_A_8E0wrzOd7_0),.clk(gclk));
	jdff dff_A_FGnF1Twi8_0(.dout(w_dff_A_8E0wrzOd7_0),.din(w_dff_A_FGnF1Twi8_0),.clk(gclk));
	jdff dff_A_8FWgaAg45_0(.dout(w_dff_A_FGnF1Twi8_0),.din(w_dff_A_8FWgaAg45_0),.clk(gclk));
	jdff dff_A_3IbXwgMp1_0(.dout(w_dff_A_8FWgaAg45_0),.din(w_dff_A_3IbXwgMp1_0),.clk(gclk));
	jdff dff_A_ZLevxzaJ1_0(.dout(w_dff_A_3IbXwgMp1_0),.din(w_dff_A_ZLevxzaJ1_0),.clk(gclk));
	jdff dff_A_BgRLUtul7_0(.dout(w_dff_A_ZLevxzaJ1_0),.din(w_dff_A_BgRLUtul7_0),.clk(gclk));
	jdff dff_A_sg8rqorY3_0(.dout(w_dff_A_BgRLUtul7_0),.din(w_dff_A_sg8rqorY3_0),.clk(gclk));
	jdff dff_A_fa6nMazo9_0(.dout(w_dff_A_sg8rqorY3_0),.din(w_dff_A_fa6nMazo9_0),.clk(gclk));
	jdff dff_A_p5UHkiEQ0_0(.dout(w_dff_A_fa6nMazo9_0),.din(w_dff_A_p5UHkiEQ0_0),.clk(gclk));
	jdff dff_A_Ye9ch74A0_0(.dout(w_dff_A_p5UHkiEQ0_0),.din(w_dff_A_Ye9ch74A0_0),.clk(gclk));
	jdff dff_A_spBK6mPB3_0(.dout(w_dff_A_Ye9ch74A0_0),.din(w_dff_A_spBK6mPB3_0),.clk(gclk));
	jdff dff_A_oFRqVpEZ1_0(.dout(w_dff_A_spBK6mPB3_0),.din(w_dff_A_oFRqVpEZ1_0),.clk(gclk));
	jdff dff_A_FYQN9leY6_0(.dout(w_dff_A_oFRqVpEZ1_0),.din(w_dff_A_FYQN9leY6_0),.clk(gclk));
	jdff dff_A_OeR9mgBf7_0(.dout(w_dff_A_FYQN9leY6_0),.din(w_dff_A_OeR9mgBf7_0),.clk(gclk));
	jdff dff_A_6IydYeZ35_0(.dout(w_dff_A_OeR9mgBf7_0),.din(w_dff_A_6IydYeZ35_0),.clk(gclk));
	jdff dff_A_fpoXmepm6_0(.dout(w_dff_A_6IydYeZ35_0),.din(w_dff_A_fpoXmepm6_0),.clk(gclk));
	jdff dff_A_QailJnZE4_0(.dout(w_dff_A_fpoXmepm6_0),.din(w_dff_A_QailJnZE4_0),.clk(gclk));
	jdff dff_A_PxFHXmx40_0(.dout(w_dff_A_QailJnZE4_0),.din(w_dff_A_PxFHXmx40_0),.clk(gclk));
	jdff dff_A_CaQIVJYX8_0(.dout(w_dff_A_PxFHXmx40_0),.din(w_dff_A_CaQIVJYX8_0),.clk(gclk));
	jdff dff_A_qSSv5qNJ3_0(.dout(w_dff_A_CaQIVJYX8_0),.din(w_dff_A_qSSv5qNJ3_0),.clk(gclk));
	jdff dff_A_lztAnQVH3_0(.dout(w_dff_A_qSSv5qNJ3_0),.din(w_dff_A_lztAnQVH3_0),.clk(gclk));
	jdff dff_A_wLoomBFP2_0(.dout(w_dff_A_lztAnQVH3_0),.din(w_dff_A_wLoomBFP2_0),.clk(gclk));
	jdff dff_A_MoHgFzyH7_0(.dout(w_dff_A_wLoomBFP2_0),.din(w_dff_A_MoHgFzyH7_0),.clk(gclk));
	jdff dff_A_m1KXgRUx1_0(.dout(w_dff_A_MoHgFzyH7_0),.din(w_dff_A_m1KXgRUx1_0),.clk(gclk));
	jdff dff_A_TP7SxmJx9_0(.dout(w_dff_A_m1KXgRUx1_0),.din(w_dff_A_TP7SxmJx9_0),.clk(gclk));
	jdff dff_A_V61aGOcA3_0(.dout(w_dff_A_TP7SxmJx9_0),.din(w_dff_A_V61aGOcA3_0),.clk(gclk));
	jdff dff_A_8nZPzhWn0_0(.dout(w_n630_0[0]),.din(w_dff_A_8nZPzhWn0_0),.clk(gclk));
	jdff dff_B_ceJJ1TqA2_1(.din(n558),.dout(w_dff_B_ceJJ1TqA2_1),.clk(gclk));
	jdff dff_A_P6dJldKc0_0(.dout(w_n477_0[0]),.din(w_dff_A_P6dJldKc0_0),.clk(gclk));
	jdff dff_A_x6mkCbD29_0(.dout(w_dff_A_P6dJldKc0_0),.din(w_dff_A_x6mkCbD29_0),.clk(gclk));
	jdff dff_A_hvsux0TA0_0(.dout(w_dff_A_x6mkCbD29_0),.din(w_dff_A_hvsux0TA0_0),.clk(gclk));
	jdff dff_A_U6oKz77h8_0(.dout(w_dff_A_hvsux0TA0_0),.din(w_dff_A_U6oKz77h8_0),.clk(gclk));
	jdff dff_A_2qflyQ9V8_0(.dout(w_dff_A_U6oKz77h8_0),.din(w_dff_A_2qflyQ9V8_0),.clk(gclk));
	jdff dff_A_r3vTuDxT8_0(.dout(w_dff_A_2qflyQ9V8_0),.din(w_dff_A_r3vTuDxT8_0),.clk(gclk));
	jdff dff_A_QKav6WDD9_0(.dout(w_dff_A_r3vTuDxT8_0),.din(w_dff_A_QKav6WDD9_0),.clk(gclk));
	jdff dff_A_wotP33kW4_0(.dout(w_dff_A_QKav6WDD9_0),.din(w_dff_A_wotP33kW4_0),.clk(gclk));
	jdff dff_A_FYhn0K6s0_0(.dout(w_dff_A_wotP33kW4_0),.din(w_dff_A_FYhn0K6s0_0),.clk(gclk));
	jdff dff_A_NEr2QcCr4_0(.dout(w_dff_A_FYhn0K6s0_0),.din(w_dff_A_NEr2QcCr4_0),.clk(gclk));
	jdff dff_A_fVHvH0Nz1_0(.dout(w_dff_A_NEr2QcCr4_0),.din(w_dff_A_fVHvH0Nz1_0),.clk(gclk));
	jdff dff_A_W4O9bCZS5_0(.dout(w_dff_A_fVHvH0Nz1_0),.din(w_dff_A_W4O9bCZS5_0),.clk(gclk));
	jdff dff_A_U8nw2nkM6_0(.dout(w_dff_A_W4O9bCZS5_0),.din(w_dff_A_U8nw2nkM6_0),.clk(gclk));
	jdff dff_A_oSDvXZGQ8_0(.dout(w_dff_A_U8nw2nkM6_0),.din(w_dff_A_oSDvXZGQ8_0),.clk(gclk));
	jdff dff_A_QTqKNitV0_0(.dout(w_dff_A_oSDvXZGQ8_0),.din(w_dff_A_QTqKNitV0_0),.clk(gclk));
	jdff dff_A_nzcDwDXq8_0(.dout(w_dff_A_QTqKNitV0_0),.din(w_dff_A_nzcDwDXq8_0),.clk(gclk));
	jdff dff_A_UDeiaAs46_0(.dout(w_dff_A_nzcDwDXq8_0),.din(w_dff_A_UDeiaAs46_0),.clk(gclk));
	jdff dff_A_2y9Kiczx8_0(.dout(w_dff_A_UDeiaAs46_0),.din(w_dff_A_2y9Kiczx8_0),.clk(gclk));
	jdff dff_A_rOYROLLh6_0(.dout(w_dff_A_2y9Kiczx8_0),.din(w_dff_A_rOYROLLh6_0),.clk(gclk));
	jdff dff_A_Aoo1p9QS5_0(.dout(w_dff_A_rOYROLLh6_0),.din(w_dff_A_Aoo1p9QS5_0),.clk(gclk));
	jdff dff_A_5CtkRo1O9_0(.dout(w_dff_A_Aoo1p9QS5_0),.din(w_dff_A_5CtkRo1O9_0),.clk(gclk));
	jdff dff_A_5KCFZhqS6_0(.dout(w_dff_A_5CtkRo1O9_0),.din(w_dff_A_5KCFZhqS6_0),.clk(gclk));
	jdff dff_A_XVNGvzzC1_0(.dout(w_dff_A_5KCFZhqS6_0),.din(w_dff_A_XVNGvzzC1_0),.clk(gclk));
	jdff dff_A_wyWBpMfD2_0(.dout(w_dff_A_XVNGvzzC1_0),.din(w_dff_A_wyWBpMfD2_0),.clk(gclk));
	jdff dff_A_2LZFltMa0_0(.dout(w_dff_A_wyWBpMfD2_0),.din(w_dff_A_2LZFltMa0_0),.clk(gclk));
	jdff dff_A_YI0jEpQn0_0(.dout(w_dff_A_2LZFltMa0_0),.din(w_dff_A_YI0jEpQn0_0),.clk(gclk));
	jdff dff_A_IyPEsJ6c7_0(.dout(w_dff_A_YI0jEpQn0_0),.din(w_dff_A_IyPEsJ6c7_0),.clk(gclk));
	jdff dff_A_dFHcTdGH8_0(.dout(w_dff_A_IyPEsJ6c7_0),.din(w_dff_A_dFHcTdGH8_0),.clk(gclk));
	jdff dff_A_CoUUaYe63_0(.dout(w_dff_A_dFHcTdGH8_0),.din(w_dff_A_CoUUaYe63_0),.clk(gclk));
	jdff dff_A_OzxLbf6k9_0(.dout(w_n544_0[0]),.din(w_dff_A_OzxLbf6k9_0),.clk(gclk));
	jdff dff_B_gogWROKv2_1(.din(n479),.dout(w_dff_B_gogWROKv2_1),.clk(gclk));
	jdff dff_A_v21n0fTZ4_0(.dout(w_n405_0[0]),.din(w_dff_A_v21n0fTZ4_0),.clk(gclk));
	jdff dff_A_VILfCfRD9_0(.dout(w_dff_A_v21n0fTZ4_0),.din(w_dff_A_VILfCfRD9_0),.clk(gclk));
	jdff dff_A_XKmlLdVR4_0(.dout(w_dff_A_VILfCfRD9_0),.din(w_dff_A_XKmlLdVR4_0),.clk(gclk));
	jdff dff_A_x92JFB3l0_0(.dout(w_dff_A_XKmlLdVR4_0),.din(w_dff_A_x92JFB3l0_0),.clk(gclk));
	jdff dff_A_pRdAAAwT4_0(.dout(w_dff_A_x92JFB3l0_0),.din(w_dff_A_pRdAAAwT4_0),.clk(gclk));
	jdff dff_A_vKtNUfFu8_0(.dout(w_dff_A_pRdAAAwT4_0),.din(w_dff_A_vKtNUfFu8_0),.clk(gclk));
	jdff dff_A_lbrnj7yG3_0(.dout(w_dff_A_vKtNUfFu8_0),.din(w_dff_A_lbrnj7yG3_0),.clk(gclk));
	jdff dff_A_7y4nNyga7_0(.dout(w_dff_A_lbrnj7yG3_0),.din(w_dff_A_7y4nNyga7_0),.clk(gclk));
	jdff dff_A_GbCvOvxI3_0(.dout(w_dff_A_7y4nNyga7_0),.din(w_dff_A_GbCvOvxI3_0),.clk(gclk));
	jdff dff_A_sm1ugC7Q9_0(.dout(w_dff_A_GbCvOvxI3_0),.din(w_dff_A_sm1ugC7Q9_0),.clk(gclk));
	jdff dff_A_BIg1jQKh9_0(.dout(w_dff_A_sm1ugC7Q9_0),.din(w_dff_A_BIg1jQKh9_0),.clk(gclk));
	jdff dff_A_aK53XAkd9_0(.dout(w_dff_A_BIg1jQKh9_0),.din(w_dff_A_aK53XAkd9_0),.clk(gclk));
	jdff dff_A_kUkYfGiZ6_0(.dout(w_dff_A_aK53XAkd9_0),.din(w_dff_A_kUkYfGiZ6_0),.clk(gclk));
	jdff dff_A_uHWkqcUh3_0(.dout(w_dff_A_kUkYfGiZ6_0),.din(w_dff_A_uHWkqcUh3_0),.clk(gclk));
	jdff dff_A_C9NYpTyg8_0(.dout(w_dff_A_uHWkqcUh3_0),.din(w_dff_A_C9NYpTyg8_0),.clk(gclk));
	jdff dff_A_1ZSlr2KI2_0(.dout(w_dff_A_C9NYpTyg8_0),.din(w_dff_A_1ZSlr2KI2_0),.clk(gclk));
	jdff dff_A_S7ZC8g7x1_0(.dout(w_dff_A_1ZSlr2KI2_0),.din(w_dff_A_S7ZC8g7x1_0),.clk(gclk));
	jdff dff_A_Qgvyx5An0_0(.dout(w_dff_A_S7ZC8g7x1_0),.din(w_dff_A_Qgvyx5An0_0),.clk(gclk));
	jdff dff_A_2vqSeVJR0_0(.dout(w_dff_A_Qgvyx5An0_0),.din(w_dff_A_2vqSeVJR0_0),.clk(gclk));
	jdff dff_A_viXzDErQ3_0(.dout(w_dff_A_2vqSeVJR0_0),.din(w_dff_A_viXzDErQ3_0),.clk(gclk));
	jdff dff_A_kpOJqIyM6_0(.dout(w_dff_A_viXzDErQ3_0),.din(w_dff_A_kpOJqIyM6_0),.clk(gclk));
	jdff dff_A_oEz2Eta81_0(.dout(w_dff_A_kpOJqIyM6_0),.din(w_dff_A_oEz2Eta81_0),.clk(gclk));
	jdff dff_A_bva2DfvG1_0(.dout(w_dff_A_oEz2Eta81_0),.din(w_dff_A_bva2DfvG1_0),.clk(gclk));
	jdff dff_A_DNk0Tqry6_0(.dout(w_dff_A_bva2DfvG1_0),.din(w_dff_A_DNk0Tqry6_0),.clk(gclk));
	jdff dff_A_VuyPjDBI5_0(.dout(w_dff_A_DNk0Tqry6_0),.din(w_dff_A_VuyPjDBI5_0),.clk(gclk));
	jdff dff_A_QtvxpQdK0_0(.dout(w_dff_A_VuyPjDBI5_0),.din(w_dff_A_QtvxpQdK0_0),.clk(gclk));
	jdff dff_A_pvQlB12I5_0(.dout(w_n465_0[0]),.din(w_dff_A_pvQlB12I5_0),.clk(gclk));
	jdff dff_B_NRDAfc2w1_1(.din(n407),.dout(w_dff_B_NRDAfc2w1_1),.clk(gclk));
	jdff dff_A_EFaKOvSU7_0(.dout(w_n341_0[0]),.din(w_dff_A_EFaKOvSU7_0),.clk(gclk));
	jdff dff_A_F9W2pI9J0_0(.dout(w_dff_A_EFaKOvSU7_0),.din(w_dff_A_F9W2pI9J0_0),.clk(gclk));
	jdff dff_A_MKkkEXvY5_0(.dout(w_dff_A_F9W2pI9J0_0),.din(w_dff_A_MKkkEXvY5_0),.clk(gclk));
	jdff dff_A_9wQh1g897_0(.dout(w_dff_A_MKkkEXvY5_0),.din(w_dff_A_9wQh1g897_0),.clk(gclk));
	jdff dff_A_pP0MZyNU7_0(.dout(w_dff_A_9wQh1g897_0),.din(w_dff_A_pP0MZyNU7_0),.clk(gclk));
	jdff dff_A_dafSOxb04_0(.dout(w_dff_A_pP0MZyNU7_0),.din(w_dff_A_dafSOxb04_0),.clk(gclk));
	jdff dff_A_SEhsINf50_0(.dout(w_dff_A_dafSOxb04_0),.din(w_dff_A_SEhsINf50_0),.clk(gclk));
	jdff dff_A_x5GVXpIL1_0(.dout(w_dff_A_SEhsINf50_0),.din(w_dff_A_x5GVXpIL1_0),.clk(gclk));
	jdff dff_A_SMUWz6sn9_0(.dout(w_dff_A_x5GVXpIL1_0),.din(w_dff_A_SMUWz6sn9_0),.clk(gclk));
	jdff dff_A_0MaEnKQ37_0(.dout(w_dff_A_SMUWz6sn9_0),.din(w_dff_A_0MaEnKQ37_0),.clk(gclk));
	jdff dff_A_uYojGnKC8_0(.dout(w_dff_A_0MaEnKQ37_0),.din(w_dff_A_uYojGnKC8_0),.clk(gclk));
	jdff dff_A_7b83H1by4_0(.dout(w_dff_A_uYojGnKC8_0),.din(w_dff_A_7b83H1by4_0),.clk(gclk));
	jdff dff_A_Ub93Ysst8_0(.dout(w_dff_A_7b83H1by4_0),.din(w_dff_A_Ub93Ysst8_0),.clk(gclk));
	jdff dff_A_yIPqrXrz2_0(.dout(w_dff_A_Ub93Ysst8_0),.din(w_dff_A_yIPqrXrz2_0),.clk(gclk));
	jdff dff_A_s33j0M6c0_0(.dout(w_dff_A_yIPqrXrz2_0),.din(w_dff_A_s33j0M6c0_0),.clk(gclk));
	jdff dff_A_u8e92U088_0(.dout(w_dff_A_s33j0M6c0_0),.din(w_dff_A_u8e92U088_0),.clk(gclk));
	jdff dff_A_KjTGQSAi7_0(.dout(w_dff_A_u8e92U088_0),.din(w_dff_A_KjTGQSAi7_0),.clk(gclk));
	jdff dff_A_Ohaj9CmS3_0(.dout(w_dff_A_KjTGQSAi7_0),.din(w_dff_A_Ohaj9CmS3_0),.clk(gclk));
	jdff dff_A_wCqiOfDk2_0(.dout(w_dff_A_Ohaj9CmS3_0),.din(w_dff_A_wCqiOfDk2_0),.clk(gclk));
	jdff dff_A_nek62cl68_0(.dout(w_dff_A_wCqiOfDk2_0),.din(w_dff_A_nek62cl68_0),.clk(gclk));
	jdff dff_A_9rEGXyCu4_0(.dout(w_dff_A_nek62cl68_0),.din(w_dff_A_9rEGXyCu4_0),.clk(gclk));
	jdff dff_A_M2X7AVgt9_0(.dout(w_dff_A_9rEGXyCu4_0),.din(w_dff_A_M2X7AVgt9_0),.clk(gclk));
	jdff dff_A_wwsr9i9c7_0(.dout(w_dff_A_M2X7AVgt9_0),.din(w_dff_A_wwsr9i9c7_0),.clk(gclk));
	jdff dff_A_kU40C3S38_0(.dout(w_n393_0[0]),.din(w_dff_A_kU40C3S38_0),.clk(gclk));
	jdff dff_B_MxR0tMp03_1(.din(n343),.dout(w_dff_B_MxR0tMp03_1),.clk(gclk));
	jdff dff_A_FLit4rH82_0(.dout(w_n283_0[0]),.din(w_dff_A_FLit4rH82_0),.clk(gclk));
	jdff dff_A_mP77Y0bP5_0(.dout(w_dff_A_FLit4rH82_0),.din(w_dff_A_mP77Y0bP5_0),.clk(gclk));
	jdff dff_A_uxR7mQh25_0(.dout(w_dff_A_mP77Y0bP5_0),.din(w_dff_A_uxR7mQh25_0),.clk(gclk));
	jdff dff_A_XD2yMGAe1_0(.dout(w_dff_A_uxR7mQh25_0),.din(w_dff_A_XD2yMGAe1_0),.clk(gclk));
	jdff dff_A_92gyhUh10_0(.dout(w_dff_A_XD2yMGAe1_0),.din(w_dff_A_92gyhUh10_0),.clk(gclk));
	jdff dff_A_TmepH2FY5_0(.dout(w_dff_A_92gyhUh10_0),.din(w_dff_A_TmepH2FY5_0),.clk(gclk));
	jdff dff_A_Pb1Ua0MB8_0(.dout(w_dff_A_TmepH2FY5_0),.din(w_dff_A_Pb1Ua0MB8_0),.clk(gclk));
	jdff dff_A_8dbla37a9_0(.dout(w_dff_A_Pb1Ua0MB8_0),.din(w_dff_A_8dbla37a9_0),.clk(gclk));
	jdff dff_A_XYdVrmuR4_0(.dout(w_dff_A_8dbla37a9_0),.din(w_dff_A_XYdVrmuR4_0),.clk(gclk));
	jdff dff_A_430wvDOS2_0(.dout(w_dff_A_XYdVrmuR4_0),.din(w_dff_A_430wvDOS2_0),.clk(gclk));
	jdff dff_A_AxfoHPAD1_0(.dout(w_dff_A_430wvDOS2_0),.din(w_dff_A_AxfoHPAD1_0),.clk(gclk));
	jdff dff_A_bCANLyk59_0(.dout(w_dff_A_AxfoHPAD1_0),.din(w_dff_A_bCANLyk59_0),.clk(gclk));
	jdff dff_A_IQiOv7Kf8_0(.dout(w_dff_A_bCANLyk59_0),.din(w_dff_A_IQiOv7Kf8_0),.clk(gclk));
	jdff dff_A_wHQKoMmj4_0(.dout(w_dff_A_IQiOv7Kf8_0),.din(w_dff_A_wHQKoMmj4_0),.clk(gclk));
	jdff dff_A_TFEjcWnh6_0(.dout(w_dff_A_wHQKoMmj4_0),.din(w_dff_A_TFEjcWnh6_0),.clk(gclk));
	jdff dff_A_OBycHW4B6_0(.dout(w_dff_A_TFEjcWnh6_0),.din(w_dff_A_OBycHW4B6_0),.clk(gclk));
	jdff dff_A_Tdsyh3pk5_0(.dout(w_dff_A_OBycHW4B6_0),.din(w_dff_A_Tdsyh3pk5_0),.clk(gclk));
	jdff dff_A_uUK32Z9q1_0(.dout(w_dff_A_Tdsyh3pk5_0),.din(w_dff_A_uUK32Z9q1_0),.clk(gclk));
	jdff dff_A_DUFK8B177_0(.dout(w_dff_A_uUK32Z9q1_0),.din(w_dff_A_DUFK8B177_0),.clk(gclk));
	jdff dff_A_OPdTFdsX8_0(.dout(w_dff_A_DUFK8B177_0),.din(w_dff_A_OPdTFdsX8_0),.clk(gclk));
	jdff dff_A_iWTcsfKo0_0(.dout(w_n329_0[0]),.din(w_dff_A_iWTcsfKo0_0),.clk(gclk));
	jdff dff_B_9jqgJuYA5_1(.din(n285),.dout(w_dff_B_9jqgJuYA5_1),.clk(gclk));
	jdff dff_A_gbicxs0O4_0(.dout(w_n232_0[0]),.din(w_dff_A_gbicxs0O4_0),.clk(gclk));
	jdff dff_A_cHAz5HE42_0(.dout(w_dff_A_gbicxs0O4_0),.din(w_dff_A_cHAz5HE42_0),.clk(gclk));
	jdff dff_A_RrNwHRsJ0_0(.dout(w_dff_A_cHAz5HE42_0),.din(w_dff_A_RrNwHRsJ0_0),.clk(gclk));
	jdff dff_A_SWr58CsJ3_0(.dout(w_dff_A_RrNwHRsJ0_0),.din(w_dff_A_SWr58CsJ3_0),.clk(gclk));
	jdff dff_A_rl4DFSnm6_0(.dout(w_dff_A_SWr58CsJ3_0),.din(w_dff_A_rl4DFSnm6_0),.clk(gclk));
	jdff dff_A_vj842KFM7_0(.dout(w_dff_A_rl4DFSnm6_0),.din(w_dff_A_vj842KFM7_0),.clk(gclk));
	jdff dff_A_vs0t15Ym1_0(.dout(w_dff_A_vj842KFM7_0),.din(w_dff_A_vs0t15Ym1_0),.clk(gclk));
	jdff dff_A_9njqBmUc0_0(.dout(w_dff_A_vs0t15Ym1_0),.din(w_dff_A_9njqBmUc0_0),.clk(gclk));
	jdff dff_A_fhxewFaJ4_0(.dout(w_dff_A_9njqBmUc0_0),.din(w_dff_A_fhxewFaJ4_0),.clk(gclk));
	jdff dff_A_vtSVeODc7_0(.dout(w_dff_A_fhxewFaJ4_0),.din(w_dff_A_vtSVeODc7_0),.clk(gclk));
	jdff dff_A_GNnBl4sc3_0(.dout(w_dff_A_vtSVeODc7_0),.din(w_dff_A_GNnBl4sc3_0),.clk(gclk));
	jdff dff_A_g5m0mqt44_0(.dout(w_dff_A_GNnBl4sc3_0),.din(w_dff_A_g5m0mqt44_0),.clk(gclk));
	jdff dff_A_pVJcJDce9_0(.dout(w_dff_A_g5m0mqt44_0),.din(w_dff_A_pVJcJDce9_0),.clk(gclk));
	jdff dff_A_Xe22HY7d1_0(.dout(w_dff_A_pVJcJDce9_0),.din(w_dff_A_Xe22HY7d1_0),.clk(gclk));
	jdff dff_A_DIlmSFjG2_0(.dout(w_dff_A_Xe22HY7d1_0),.din(w_dff_A_DIlmSFjG2_0),.clk(gclk));
	jdff dff_A_Mbt6qhLF3_0(.dout(w_dff_A_DIlmSFjG2_0),.din(w_dff_A_Mbt6qhLF3_0),.clk(gclk));
	jdff dff_A_jgurZwdt9_0(.dout(w_dff_A_Mbt6qhLF3_0),.din(w_dff_A_jgurZwdt9_0),.clk(gclk));
	jdff dff_A_6MqYMjVg1_0(.dout(w_n271_0[0]),.din(w_dff_A_6MqYMjVg1_0),.clk(gclk));
	jdff dff_B_dAuOBgIL1_1(.din(n234),.dout(w_dff_B_dAuOBgIL1_1),.clk(gclk));
	jdff dff_A_xR1gWTJD2_0(.dout(w_n189_0[0]),.din(w_dff_A_xR1gWTJD2_0),.clk(gclk));
	jdff dff_A_F0WIojUQ1_0(.dout(w_dff_A_xR1gWTJD2_0),.din(w_dff_A_F0WIojUQ1_0),.clk(gclk));
	jdff dff_A_640Skq8P8_0(.dout(w_dff_A_F0WIojUQ1_0),.din(w_dff_A_640Skq8P8_0),.clk(gclk));
	jdff dff_A_Nhn8XYwv4_0(.dout(w_dff_A_640Skq8P8_0),.din(w_dff_A_Nhn8XYwv4_0),.clk(gclk));
	jdff dff_A_RFyH1kny0_0(.dout(w_dff_A_Nhn8XYwv4_0),.din(w_dff_A_RFyH1kny0_0),.clk(gclk));
	jdff dff_A_LrCsXBUG6_0(.dout(w_dff_A_RFyH1kny0_0),.din(w_dff_A_LrCsXBUG6_0),.clk(gclk));
	jdff dff_A_DBQeq0Fo2_0(.dout(w_dff_A_LrCsXBUG6_0),.din(w_dff_A_DBQeq0Fo2_0),.clk(gclk));
	jdff dff_A_9mbuu8nP3_0(.dout(w_dff_A_DBQeq0Fo2_0),.din(w_dff_A_9mbuu8nP3_0),.clk(gclk));
	jdff dff_A_uy2i3tGS0_0(.dout(w_dff_A_9mbuu8nP3_0),.din(w_dff_A_uy2i3tGS0_0),.clk(gclk));
	jdff dff_A_eRscqzXf0_0(.dout(w_dff_A_uy2i3tGS0_0),.din(w_dff_A_eRscqzXf0_0),.clk(gclk));
	jdff dff_A_7XGsQS204_0(.dout(w_dff_A_eRscqzXf0_0),.din(w_dff_A_7XGsQS204_0),.clk(gclk));
	jdff dff_A_81lRWZBC6_0(.dout(w_dff_A_7XGsQS204_0),.din(w_dff_A_81lRWZBC6_0),.clk(gclk));
	jdff dff_A_jTQmQ8Kn5_0(.dout(w_dff_A_81lRWZBC6_0),.din(w_dff_A_jTQmQ8Kn5_0),.clk(gclk));
	jdff dff_A_ashIQI344_0(.dout(w_dff_A_jTQmQ8Kn5_0),.din(w_dff_A_ashIQI344_0),.clk(gclk));
	jdff dff_A_DPpMOZQn6_0(.dout(w_n220_0[0]),.din(w_dff_A_DPpMOZQn6_0),.clk(gclk));
	jdff dff_B_ScOtqCUR0_1(.din(n191),.dout(w_dff_B_ScOtqCUR0_1),.clk(gclk));
	jdff dff_A_pVE7kE5D0_0(.dout(w_n151_0[0]),.din(w_dff_A_pVE7kE5D0_0),.clk(gclk));
	jdff dff_A_nXxWpgoZ6_0(.dout(w_dff_A_pVE7kE5D0_0),.din(w_dff_A_nXxWpgoZ6_0),.clk(gclk));
	jdff dff_A_MbDdXnqq0_0(.dout(w_dff_A_nXxWpgoZ6_0),.din(w_dff_A_MbDdXnqq0_0),.clk(gclk));
	jdff dff_A_4Vysn0yB1_0(.dout(w_dff_A_MbDdXnqq0_0),.din(w_dff_A_4Vysn0yB1_0),.clk(gclk));
	jdff dff_A_AaMmI03z0_0(.dout(w_dff_A_4Vysn0yB1_0),.din(w_dff_A_AaMmI03z0_0),.clk(gclk));
	jdff dff_A_0wW5U7509_0(.dout(w_dff_A_AaMmI03z0_0),.din(w_dff_A_0wW5U7509_0),.clk(gclk));
	jdff dff_A_lnPhx0Ix4_0(.dout(w_dff_A_0wW5U7509_0),.din(w_dff_A_lnPhx0Ix4_0),.clk(gclk));
	jdff dff_A_Hmj2pzsU1_0(.dout(w_dff_A_lnPhx0Ix4_0),.din(w_dff_A_Hmj2pzsU1_0),.clk(gclk));
	jdff dff_A_VfvNn8Ru3_0(.dout(w_dff_A_Hmj2pzsU1_0),.din(w_dff_A_VfvNn8Ru3_0),.clk(gclk));
	jdff dff_A_lVMWhBhW4_0(.dout(w_dff_A_VfvNn8Ru3_0),.din(w_dff_A_lVMWhBhW4_0),.clk(gclk));
	jdff dff_A_Npyp55tc1_0(.dout(w_dff_A_lVMWhBhW4_0),.din(w_dff_A_Npyp55tc1_0),.clk(gclk));
	jdff dff_A_JG8iwnZG5_0(.dout(w_n177_0[0]),.din(w_dff_A_JG8iwnZG5_0),.clk(gclk));
	jdff dff_B_6qB0mknv3_1(.din(n153),.dout(w_dff_B_6qB0mknv3_1),.clk(gclk));
	jdff dff_A_JbFnYCS59_0(.dout(w_n116_0[0]),.din(w_dff_A_JbFnYCS59_0),.clk(gclk));
	jdff dff_A_i1TlMSzT1_0(.dout(w_dff_A_JbFnYCS59_0),.din(w_dff_A_i1TlMSzT1_0),.clk(gclk));
	jdff dff_A_55wZ5YOo2_0(.dout(w_dff_A_i1TlMSzT1_0),.din(w_dff_A_55wZ5YOo2_0),.clk(gclk));
	jdff dff_A_LYe7BlVf2_0(.dout(w_dff_A_55wZ5YOo2_0),.din(w_dff_A_LYe7BlVf2_0),.clk(gclk));
	jdff dff_A_e6xyxHaw5_0(.dout(w_dff_A_LYe7BlVf2_0),.din(w_dff_A_e6xyxHaw5_0),.clk(gclk));
	jdff dff_A_RryRbKAU6_0(.dout(w_dff_A_e6xyxHaw5_0),.din(w_dff_A_RryRbKAU6_0),.clk(gclk));
	jdff dff_A_zBfqEmkV3_0(.dout(w_dff_A_RryRbKAU6_0),.din(w_dff_A_zBfqEmkV3_0),.clk(gclk));
	jdff dff_A_t8goGsCr9_0(.dout(w_dff_A_zBfqEmkV3_0),.din(w_dff_A_t8goGsCr9_0),.clk(gclk));
	jdff dff_A_1LCq0UX68_0(.dout(w_n139_0[0]),.din(w_dff_A_1LCq0UX68_0),.clk(gclk));
	jdff dff_A_IGVxKSBU0_0(.dout(w_n104_0[0]),.din(w_dff_A_IGVxKSBU0_0),.clk(gclk));
	jdff dff_A_zA7efneb1_0(.dout(w_n85_0[0]),.din(w_dff_A_zA7efneb1_0),.clk(gclk));
	jdff dff_A_wzFeeiny6_1(.dout(w_n82_1[1]),.din(w_dff_A_wzFeeiny6_1),.clk(gclk));
	jdff dff_A_8wOEl3lt9_0(.dout(w_n94_0[0]),.din(w_dff_A_8wOEl3lt9_0),.clk(gclk));
	jdff dff_A_gxb0Kmdb6_0(.dout(w_dff_A_8wOEl3lt9_0),.din(w_dff_A_gxb0Kmdb6_0),.clk(gclk));
	jdff dff_A_LRuQbPIa4_0(.dout(w_dff_A_gxb0Kmdb6_0),.din(w_dff_A_LRuQbPIa4_0),.clk(gclk));
	jdff dff_A_BmzAGfJI1_0(.dout(w_dff_A_LRuQbPIa4_0),.din(w_dff_A_BmzAGfJI1_0),.clk(gclk));
	jdff dff_A_o96JgnLg3_0(.dout(w_dff_A_BmzAGfJI1_0),.din(w_dff_A_o96JgnLg3_0),.clk(gclk));
	jdff dff_A_GRJDodBM4_0(.dout(w_n103_0[0]),.din(w_dff_A_GRJDodBM4_0),.clk(gclk));
	jdff dff_A_ULikrVqh5_0(.dout(w_dff_A_GRJDodBM4_0),.din(w_dff_A_ULikrVqh5_0),.clk(gclk));
	jdff dff_B_GllUaxUV7_1(.din(n97),.dout(w_dff_B_GllUaxUV7_1),.clk(gclk));
	jdff dff_A_2wtDOQkA6_1(.dout(w_n82_0[1]),.din(w_dff_A_2wtDOQkA6_1),.clk(gclk));
	jdff dff_A_X3OPPVNu9_2(.dout(w_n82_0[2]),.din(w_dff_A_X3OPPVNu9_2),.clk(gclk));
	jdff dff_A_isb7tLK02_2(.dout(w_dff_A_X3OPPVNu9_2),.din(w_dff_A_isb7tLK02_2),.clk(gclk));
	jdff dff_A_1qgBAHnM3_0(.dout(w_n1151_0[0]),.din(w_dff_A_1qgBAHnM3_0),.clk(gclk));
	jdff dff_B_BmLhtFuJ1_2(.din(n1151),.dout(w_dff_B_BmLhtFuJ1_2),.clk(gclk));
	jdff dff_B_ocyQzzZ21_2(.din(n1044),.dout(w_dff_B_ocyQzzZ21_2),.clk(gclk));
	jdff dff_B_rlT6IMnw4_2(.din(w_dff_B_ocyQzzZ21_2),.dout(w_dff_B_rlT6IMnw4_2),.clk(gclk));
	jdff dff_B_S06AnL1I2_2(.din(w_dff_B_rlT6IMnw4_2),.dout(w_dff_B_S06AnL1I2_2),.clk(gclk));
	jdff dff_B_GVqKwmtX8_2(.din(w_dff_B_S06AnL1I2_2),.dout(w_dff_B_GVqKwmtX8_2),.clk(gclk));
	jdff dff_B_a2AGywqX0_2(.din(w_dff_B_GVqKwmtX8_2),.dout(w_dff_B_a2AGywqX0_2),.clk(gclk));
	jdff dff_B_wPdW3wBw0_2(.din(w_dff_B_a2AGywqX0_2),.dout(w_dff_B_wPdW3wBw0_2),.clk(gclk));
	jdff dff_B_FOn5djG20_2(.din(w_dff_B_wPdW3wBw0_2),.dout(w_dff_B_FOn5djG20_2),.clk(gclk));
	jdff dff_B_MuIMJzik6_2(.din(w_dff_B_FOn5djG20_2),.dout(w_dff_B_MuIMJzik6_2),.clk(gclk));
	jdff dff_B_t4louVvR6_2(.din(w_dff_B_MuIMJzik6_2),.dout(w_dff_B_t4louVvR6_2),.clk(gclk));
	jdff dff_B_8M1DNNVT9_2(.din(w_dff_B_t4louVvR6_2),.dout(w_dff_B_8M1DNNVT9_2),.clk(gclk));
	jdff dff_B_WMtLWxSR4_2(.din(w_dff_B_8M1DNNVT9_2),.dout(w_dff_B_WMtLWxSR4_2),.clk(gclk));
	jdff dff_B_D2hovTJA7_2(.din(w_dff_B_WMtLWxSR4_2),.dout(w_dff_B_D2hovTJA7_2),.clk(gclk));
	jdff dff_B_AiX9Q5Fi9_2(.din(w_dff_B_D2hovTJA7_2),.dout(w_dff_B_AiX9Q5Fi9_2),.clk(gclk));
	jdff dff_B_fxczt5X34_2(.din(w_dff_B_AiX9Q5Fi9_2),.dout(w_dff_B_fxczt5X34_2),.clk(gclk));
	jdff dff_B_HikhZ2YX1_2(.din(w_dff_B_fxczt5X34_2),.dout(w_dff_B_HikhZ2YX1_2),.clk(gclk));
	jdff dff_B_eaS9SxWf4_2(.din(w_dff_B_HikhZ2YX1_2),.dout(w_dff_B_eaS9SxWf4_2),.clk(gclk));
	jdff dff_B_ToWGlZ6L7_2(.din(w_dff_B_eaS9SxWf4_2),.dout(w_dff_B_ToWGlZ6L7_2),.clk(gclk));
	jdff dff_B_XqaD1iUu4_2(.din(w_dff_B_ToWGlZ6L7_2),.dout(w_dff_B_XqaD1iUu4_2),.clk(gclk));
	jdff dff_B_iMY4XgAd2_2(.din(w_dff_B_XqaD1iUu4_2),.dout(w_dff_B_iMY4XgAd2_2),.clk(gclk));
	jdff dff_B_ccy3aQBn2_2(.din(w_dff_B_iMY4XgAd2_2),.dout(w_dff_B_ccy3aQBn2_2),.clk(gclk));
	jdff dff_B_8mRcifVg1_2(.din(w_dff_B_ccy3aQBn2_2),.dout(w_dff_B_8mRcifVg1_2),.clk(gclk));
	jdff dff_B_Vtzj9JXw7_2(.din(w_dff_B_8mRcifVg1_2),.dout(w_dff_B_Vtzj9JXw7_2),.clk(gclk));
	jdff dff_B_NgY4FC6y5_2(.din(w_dff_B_Vtzj9JXw7_2),.dout(w_dff_B_NgY4FC6y5_2),.clk(gclk));
	jdff dff_B_jPjNxvub3_2(.din(w_dff_B_NgY4FC6y5_2),.dout(w_dff_B_jPjNxvub3_2),.clk(gclk));
	jdff dff_B_jW6skY2Y9_2(.din(w_dff_B_jPjNxvub3_2),.dout(w_dff_B_jW6skY2Y9_2),.clk(gclk));
	jdff dff_B_Mlb2ZzGS0_2(.din(w_dff_B_jW6skY2Y9_2),.dout(w_dff_B_Mlb2ZzGS0_2),.clk(gclk));
	jdff dff_B_0qcN5Jcl8_2(.din(w_dff_B_Mlb2ZzGS0_2),.dout(w_dff_B_0qcN5Jcl8_2),.clk(gclk));
	jdff dff_B_02whfXKO2_2(.din(w_dff_B_0qcN5Jcl8_2),.dout(w_dff_B_02whfXKO2_2),.clk(gclk));
	jdff dff_B_yii16jwC2_2(.din(w_dff_B_02whfXKO2_2),.dout(w_dff_B_yii16jwC2_2),.clk(gclk));
	jdff dff_B_hlyFtVtZ3_2(.din(w_dff_B_yii16jwC2_2),.dout(w_dff_B_hlyFtVtZ3_2),.clk(gclk));
	jdff dff_B_Yx4TN7v45_2(.din(w_dff_B_hlyFtVtZ3_2),.dout(w_dff_B_Yx4TN7v45_2),.clk(gclk));
	jdff dff_B_Sj6uyHAj9_2(.din(w_dff_B_Yx4TN7v45_2),.dout(w_dff_B_Sj6uyHAj9_2),.clk(gclk));
	jdff dff_B_ODy9GZzg9_2(.din(w_dff_B_Sj6uyHAj9_2),.dout(w_dff_B_ODy9GZzg9_2),.clk(gclk));
	jdff dff_B_N1ACvKMH5_2(.din(w_dff_B_ODy9GZzg9_2),.dout(w_dff_B_N1ACvKMH5_2),.clk(gclk));
	jdff dff_B_fl60HsEZ2_2(.din(w_dff_B_N1ACvKMH5_2),.dout(w_dff_B_fl60HsEZ2_2),.clk(gclk));
	jdff dff_B_pAuD7G3b6_2(.din(w_dff_B_fl60HsEZ2_2),.dout(w_dff_B_pAuD7G3b6_2),.clk(gclk));
	jdff dff_B_ErWk5laX0_2(.din(w_dff_B_pAuD7G3b6_2),.dout(w_dff_B_ErWk5laX0_2),.clk(gclk));
	jdff dff_B_XZjISiha4_2(.din(w_dff_B_ErWk5laX0_2),.dout(w_dff_B_XZjISiha4_2),.clk(gclk));
	jdff dff_B_UUXTOPCD8_2(.din(w_dff_B_XZjISiha4_2),.dout(w_dff_B_UUXTOPCD8_2),.clk(gclk));
	jdff dff_B_dHfnf7lJ6_2(.din(w_dff_B_UUXTOPCD8_2),.dout(w_dff_B_dHfnf7lJ6_2),.clk(gclk));
	jdff dff_B_fFjd9uOZ2_2(.din(w_dff_B_dHfnf7lJ6_2),.dout(w_dff_B_fFjd9uOZ2_2),.clk(gclk));
	jdff dff_B_ttZn8Y1j7_2(.din(w_dff_B_fFjd9uOZ2_2),.dout(w_dff_B_ttZn8Y1j7_2),.clk(gclk));
	jdff dff_B_q4ru4Yif6_2(.din(w_dff_B_ttZn8Y1j7_2),.dout(w_dff_B_q4ru4Yif6_2),.clk(gclk));
	jdff dff_B_aZrjLaUP2_2(.din(w_dff_B_q4ru4Yif6_2),.dout(w_dff_B_aZrjLaUP2_2),.clk(gclk));
	jdff dff_A_kLeTUCqx2_0(.dout(w_n1048_0[0]),.din(w_dff_A_kLeTUCqx2_0),.clk(gclk));
	jdff dff_B_UWPl9sBx1_1(.din(n1046),.dout(w_dff_B_UWPl9sBx1_1),.clk(gclk));
	jdff dff_B_6VcU4rsP4_2(.din(n943),.dout(w_dff_B_6VcU4rsP4_2),.clk(gclk));
	jdff dff_B_xXkI68eK1_2(.din(w_dff_B_6VcU4rsP4_2),.dout(w_dff_B_xXkI68eK1_2),.clk(gclk));
	jdff dff_B_j32ADvOg1_2(.din(w_dff_B_xXkI68eK1_2),.dout(w_dff_B_j32ADvOg1_2),.clk(gclk));
	jdff dff_B_apGrgngt8_2(.din(w_dff_B_j32ADvOg1_2),.dout(w_dff_B_apGrgngt8_2),.clk(gclk));
	jdff dff_B_SbNGzs4J6_2(.din(w_dff_B_apGrgngt8_2),.dout(w_dff_B_SbNGzs4J6_2),.clk(gclk));
	jdff dff_B_03NIjkI52_2(.din(w_dff_B_SbNGzs4J6_2),.dout(w_dff_B_03NIjkI52_2),.clk(gclk));
	jdff dff_B_bCRIOj3k1_2(.din(w_dff_B_03NIjkI52_2),.dout(w_dff_B_bCRIOj3k1_2),.clk(gclk));
	jdff dff_B_C8OKsyJY5_2(.din(w_dff_B_bCRIOj3k1_2),.dout(w_dff_B_C8OKsyJY5_2),.clk(gclk));
	jdff dff_B_yFH92Y7X3_2(.din(w_dff_B_C8OKsyJY5_2),.dout(w_dff_B_yFH92Y7X3_2),.clk(gclk));
	jdff dff_B_LRDRYvPu5_2(.din(w_dff_B_yFH92Y7X3_2),.dout(w_dff_B_LRDRYvPu5_2),.clk(gclk));
	jdff dff_B_EROViqrh7_2(.din(w_dff_B_LRDRYvPu5_2),.dout(w_dff_B_EROViqrh7_2),.clk(gclk));
	jdff dff_B_TPUpIvki3_2(.din(w_dff_B_EROViqrh7_2),.dout(w_dff_B_TPUpIvki3_2),.clk(gclk));
	jdff dff_B_DEg7uwmr2_2(.din(w_dff_B_TPUpIvki3_2),.dout(w_dff_B_DEg7uwmr2_2),.clk(gclk));
	jdff dff_B_is3IUrvB0_2(.din(w_dff_B_DEg7uwmr2_2),.dout(w_dff_B_is3IUrvB0_2),.clk(gclk));
	jdff dff_B_vWBpL7ha8_2(.din(w_dff_B_is3IUrvB0_2),.dout(w_dff_B_vWBpL7ha8_2),.clk(gclk));
	jdff dff_B_jvzpxm137_2(.din(w_dff_B_vWBpL7ha8_2),.dout(w_dff_B_jvzpxm137_2),.clk(gclk));
	jdff dff_B_HSCV1UZj3_2(.din(w_dff_B_jvzpxm137_2),.dout(w_dff_B_HSCV1UZj3_2),.clk(gclk));
	jdff dff_B_kbidfiAl4_2(.din(w_dff_B_HSCV1UZj3_2),.dout(w_dff_B_kbidfiAl4_2),.clk(gclk));
	jdff dff_B_FmCeQ5XW9_2(.din(w_dff_B_kbidfiAl4_2),.dout(w_dff_B_FmCeQ5XW9_2),.clk(gclk));
	jdff dff_B_hGAzrKfH0_2(.din(w_dff_B_FmCeQ5XW9_2),.dout(w_dff_B_hGAzrKfH0_2),.clk(gclk));
	jdff dff_B_sRsis2oF1_2(.din(w_dff_B_hGAzrKfH0_2),.dout(w_dff_B_sRsis2oF1_2),.clk(gclk));
	jdff dff_B_RrRBUQwa0_2(.din(w_dff_B_sRsis2oF1_2),.dout(w_dff_B_RrRBUQwa0_2),.clk(gclk));
	jdff dff_B_JECTympL4_2(.din(w_dff_B_RrRBUQwa0_2),.dout(w_dff_B_JECTympL4_2),.clk(gclk));
	jdff dff_B_UH5Pltlm0_2(.din(w_dff_B_JECTympL4_2),.dout(w_dff_B_UH5Pltlm0_2),.clk(gclk));
	jdff dff_B_RsuIk8EJ6_2(.din(w_dff_B_UH5Pltlm0_2),.dout(w_dff_B_RsuIk8EJ6_2),.clk(gclk));
	jdff dff_B_VBB7XORv4_2(.din(w_dff_B_RsuIk8EJ6_2),.dout(w_dff_B_VBB7XORv4_2),.clk(gclk));
	jdff dff_B_Mh2uFYUk4_2(.din(w_dff_B_VBB7XORv4_2),.dout(w_dff_B_Mh2uFYUk4_2),.clk(gclk));
	jdff dff_B_e2dKciYF1_2(.din(w_dff_B_Mh2uFYUk4_2),.dout(w_dff_B_e2dKciYF1_2),.clk(gclk));
	jdff dff_B_HW40Zgwk5_2(.din(w_dff_B_e2dKciYF1_2),.dout(w_dff_B_HW40Zgwk5_2),.clk(gclk));
	jdff dff_B_hlq2KFZ66_2(.din(w_dff_B_HW40Zgwk5_2),.dout(w_dff_B_hlq2KFZ66_2),.clk(gclk));
	jdff dff_B_d1iyb83h8_2(.din(w_dff_B_hlq2KFZ66_2),.dout(w_dff_B_d1iyb83h8_2),.clk(gclk));
	jdff dff_B_o4lWT9hn1_2(.din(w_dff_B_d1iyb83h8_2),.dout(w_dff_B_o4lWT9hn1_2),.clk(gclk));
	jdff dff_B_jYBENLzS3_2(.din(w_dff_B_o4lWT9hn1_2),.dout(w_dff_B_jYBENLzS3_2),.clk(gclk));
	jdff dff_B_L7mBxDtg2_2(.din(w_dff_B_jYBENLzS3_2),.dout(w_dff_B_L7mBxDtg2_2),.clk(gclk));
	jdff dff_B_AcX11O4H3_2(.din(w_dff_B_L7mBxDtg2_2),.dout(w_dff_B_AcX11O4H3_2),.clk(gclk));
	jdff dff_B_BtUbDKoU7_2(.din(w_dff_B_AcX11O4H3_2),.dout(w_dff_B_BtUbDKoU7_2),.clk(gclk));
	jdff dff_B_wEF0KkXg4_2(.din(w_dff_B_BtUbDKoU7_2),.dout(w_dff_B_wEF0KkXg4_2),.clk(gclk));
	jdff dff_B_u2KJDh9v3_2(.din(w_dff_B_wEF0KkXg4_2),.dout(w_dff_B_u2KJDh9v3_2),.clk(gclk));
	jdff dff_B_wG1EELJS9_2(.din(w_dff_B_u2KJDh9v3_2),.dout(w_dff_B_wG1EELJS9_2),.clk(gclk));
	jdff dff_B_C6GIKeOi4_2(.din(w_dff_B_wG1EELJS9_2),.dout(w_dff_B_C6GIKeOi4_2),.clk(gclk));
	jdff dff_B_OlErDkei0_2(.din(w_dff_B_C6GIKeOi4_2),.dout(w_dff_B_OlErDkei0_2),.clk(gclk));
	jdff dff_A_rzHhCtPL6_1(.dout(w_n1032_0[1]),.din(w_dff_A_rzHhCtPL6_1),.clk(gclk));
	jdff dff_A_sfvkaepl4_0(.dout(w_n840_0[0]),.din(w_dff_A_sfvkaepl4_0),.clk(gclk));
	jdff dff_A_j09C3lLo8_0(.dout(w_dff_A_sfvkaepl4_0),.din(w_dff_A_j09C3lLo8_0),.clk(gclk));
	jdff dff_A_tHCBWyJb3_0(.dout(w_dff_A_j09C3lLo8_0),.din(w_dff_A_tHCBWyJb3_0),.clk(gclk));
	jdff dff_A_55kyTyUN6_0(.dout(w_dff_A_tHCBWyJb3_0),.din(w_dff_A_55kyTyUN6_0),.clk(gclk));
	jdff dff_A_NkHF0lWc3_0(.dout(w_dff_A_55kyTyUN6_0),.din(w_dff_A_NkHF0lWc3_0),.clk(gclk));
	jdff dff_A_GL9lb41z9_0(.dout(w_dff_A_NkHF0lWc3_0),.din(w_dff_A_GL9lb41z9_0),.clk(gclk));
	jdff dff_A_u5qBhXCf2_0(.dout(w_dff_A_GL9lb41z9_0),.din(w_dff_A_u5qBhXCf2_0),.clk(gclk));
	jdff dff_A_Xurl298G2_0(.dout(w_dff_A_u5qBhXCf2_0),.din(w_dff_A_Xurl298G2_0),.clk(gclk));
	jdff dff_A_0r240fVN2_0(.dout(w_dff_A_Xurl298G2_0),.din(w_dff_A_0r240fVN2_0),.clk(gclk));
	jdff dff_A_iHrnoSBO6_0(.dout(w_dff_A_0r240fVN2_0),.din(w_dff_A_iHrnoSBO6_0),.clk(gclk));
	jdff dff_A_gRMC4qa37_0(.dout(w_dff_A_iHrnoSBO6_0),.din(w_dff_A_gRMC4qa37_0),.clk(gclk));
	jdff dff_A_NiK3pdK10_0(.dout(w_dff_A_gRMC4qa37_0),.din(w_dff_A_NiK3pdK10_0),.clk(gclk));
	jdff dff_A_POaw8Ohg6_0(.dout(w_dff_A_NiK3pdK10_0),.din(w_dff_A_POaw8Ohg6_0),.clk(gclk));
	jdff dff_A_ziWenKew8_0(.dout(w_dff_A_POaw8Ohg6_0),.din(w_dff_A_ziWenKew8_0),.clk(gclk));
	jdff dff_A_Z54ryrHP1_0(.dout(w_dff_A_ziWenKew8_0),.din(w_dff_A_Z54ryrHP1_0),.clk(gclk));
	jdff dff_A_DdlyYtEd5_0(.dout(w_dff_A_Z54ryrHP1_0),.din(w_dff_A_DdlyYtEd5_0),.clk(gclk));
	jdff dff_A_xmNPZfBT7_0(.dout(w_dff_A_DdlyYtEd5_0),.din(w_dff_A_xmNPZfBT7_0),.clk(gclk));
	jdff dff_A_axi8cN4E5_0(.dout(w_dff_A_xmNPZfBT7_0),.din(w_dff_A_axi8cN4E5_0),.clk(gclk));
	jdff dff_A_neikj1IE3_0(.dout(w_dff_A_axi8cN4E5_0),.din(w_dff_A_neikj1IE3_0),.clk(gclk));
	jdff dff_A_csYina3v8_0(.dout(w_dff_A_neikj1IE3_0),.din(w_dff_A_csYina3v8_0),.clk(gclk));
	jdff dff_A_oW39yD0f9_0(.dout(w_dff_A_csYina3v8_0),.din(w_dff_A_oW39yD0f9_0),.clk(gclk));
	jdff dff_A_QbXBvsLp1_0(.dout(w_dff_A_oW39yD0f9_0),.din(w_dff_A_QbXBvsLp1_0),.clk(gclk));
	jdff dff_A_ghnwqKhI1_0(.dout(w_dff_A_QbXBvsLp1_0),.din(w_dff_A_ghnwqKhI1_0),.clk(gclk));
	jdff dff_A_2LDLtKfd4_0(.dout(w_dff_A_ghnwqKhI1_0),.din(w_dff_A_2LDLtKfd4_0),.clk(gclk));
	jdff dff_A_I4C6SkdQ7_0(.dout(w_dff_A_2LDLtKfd4_0),.din(w_dff_A_I4C6SkdQ7_0),.clk(gclk));
	jdff dff_A_ThYMcMxK0_0(.dout(w_dff_A_I4C6SkdQ7_0),.din(w_dff_A_ThYMcMxK0_0),.clk(gclk));
	jdff dff_A_yfPUh4IJ2_0(.dout(w_dff_A_ThYMcMxK0_0),.din(w_dff_A_yfPUh4IJ2_0),.clk(gclk));
	jdff dff_A_WCTDRuKu5_0(.dout(w_dff_A_yfPUh4IJ2_0),.din(w_dff_A_WCTDRuKu5_0),.clk(gclk));
	jdff dff_A_XcFEmsJT1_0(.dout(w_dff_A_WCTDRuKu5_0),.din(w_dff_A_XcFEmsJT1_0),.clk(gclk));
	jdff dff_A_vNu79JpS6_0(.dout(w_dff_A_XcFEmsJT1_0),.din(w_dff_A_vNu79JpS6_0),.clk(gclk));
	jdff dff_A_ImD6d5LR1_0(.dout(w_dff_A_vNu79JpS6_0),.din(w_dff_A_ImD6d5LR1_0),.clk(gclk));
	jdff dff_A_OOiy5AA68_0(.dout(w_dff_A_ImD6d5LR1_0),.din(w_dff_A_OOiy5AA68_0),.clk(gclk));
	jdff dff_A_E9MTsjz49_0(.dout(w_dff_A_OOiy5AA68_0),.din(w_dff_A_E9MTsjz49_0),.clk(gclk));
	jdff dff_A_nbq3ehR25_0(.dout(w_dff_A_E9MTsjz49_0),.din(w_dff_A_nbq3ehR25_0),.clk(gclk));
	jdff dff_A_NWSDKE085_0(.dout(w_dff_A_nbq3ehR25_0),.din(w_dff_A_NWSDKE085_0),.clk(gclk));
	jdff dff_A_uKNqnDtx9_0(.dout(w_dff_A_NWSDKE085_0),.din(w_dff_A_uKNqnDtx9_0),.clk(gclk));
	jdff dff_A_8X035g628_0(.dout(w_dff_A_uKNqnDtx9_0),.din(w_dff_A_8X035g628_0),.clk(gclk));
	jdff dff_A_8g1bLN284_0(.dout(w_dff_A_8X035g628_0),.din(w_dff_A_8g1bLN284_0),.clk(gclk));
	jdff dff_A_3epEYrKA2_1(.dout(w_n927_0[1]),.din(w_dff_A_3epEYrKA2_1),.clk(gclk));
	jdff dff_A_axzWNOhv0_2(.dout(w_n927_0[2]),.din(w_dff_A_axzWNOhv0_2),.clk(gclk));
	jdff dff_B_KML9lAql1_1(.din(n842),.dout(w_dff_B_KML9lAql1_1),.clk(gclk));
	jdff dff_B_HMGSGBSP1_2(.din(n742),.dout(w_dff_B_HMGSGBSP1_2),.clk(gclk));
	jdff dff_B_viWuZVKu5_2(.din(w_dff_B_HMGSGBSP1_2),.dout(w_dff_B_viWuZVKu5_2),.clk(gclk));
	jdff dff_B_2Ip3rDe58_2(.din(w_dff_B_viWuZVKu5_2),.dout(w_dff_B_2Ip3rDe58_2),.clk(gclk));
	jdff dff_B_3f3pOnVF1_2(.din(w_dff_B_2Ip3rDe58_2),.dout(w_dff_B_3f3pOnVF1_2),.clk(gclk));
	jdff dff_B_E1cjXEZG9_2(.din(w_dff_B_3f3pOnVF1_2),.dout(w_dff_B_E1cjXEZG9_2),.clk(gclk));
	jdff dff_B_CgVBLYsv9_2(.din(w_dff_B_E1cjXEZG9_2),.dout(w_dff_B_CgVBLYsv9_2),.clk(gclk));
	jdff dff_B_ef0mOmRk2_2(.din(w_dff_B_CgVBLYsv9_2),.dout(w_dff_B_ef0mOmRk2_2),.clk(gclk));
	jdff dff_B_VPO8kEh80_2(.din(w_dff_B_ef0mOmRk2_2),.dout(w_dff_B_VPO8kEh80_2),.clk(gclk));
	jdff dff_B_tnCHmtY43_2(.din(w_dff_B_VPO8kEh80_2),.dout(w_dff_B_tnCHmtY43_2),.clk(gclk));
	jdff dff_B_NFqTWkbm1_2(.din(w_dff_B_tnCHmtY43_2),.dout(w_dff_B_NFqTWkbm1_2),.clk(gclk));
	jdff dff_B_4vm3ZSHt4_2(.din(w_dff_B_NFqTWkbm1_2),.dout(w_dff_B_4vm3ZSHt4_2),.clk(gclk));
	jdff dff_B_jCJebprb0_2(.din(w_dff_B_4vm3ZSHt4_2),.dout(w_dff_B_jCJebprb0_2),.clk(gclk));
	jdff dff_B_5g4GjFHb2_2(.din(w_dff_B_jCJebprb0_2),.dout(w_dff_B_5g4GjFHb2_2),.clk(gclk));
	jdff dff_B_GmQejb4D7_2(.din(w_dff_B_5g4GjFHb2_2),.dout(w_dff_B_GmQejb4D7_2),.clk(gclk));
	jdff dff_B_tmAxVij19_2(.din(w_dff_B_GmQejb4D7_2),.dout(w_dff_B_tmAxVij19_2),.clk(gclk));
	jdff dff_B_Eo0JXkHB4_2(.din(w_dff_B_tmAxVij19_2),.dout(w_dff_B_Eo0JXkHB4_2),.clk(gclk));
	jdff dff_B_hnZ2YC053_2(.din(w_dff_B_Eo0JXkHB4_2),.dout(w_dff_B_hnZ2YC053_2),.clk(gclk));
	jdff dff_B_v4KJ7nUd5_2(.din(w_dff_B_hnZ2YC053_2),.dout(w_dff_B_v4KJ7nUd5_2),.clk(gclk));
	jdff dff_B_1fYsJQyi3_2(.din(w_dff_B_v4KJ7nUd5_2),.dout(w_dff_B_1fYsJQyi3_2),.clk(gclk));
	jdff dff_B_Zo9Rq65i6_2(.din(w_dff_B_1fYsJQyi3_2),.dout(w_dff_B_Zo9Rq65i6_2),.clk(gclk));
	jdff dff_B_DawQzYpX3_2(.din(w_dff_B_Zo9Rq65i6_2),.dout(w_dff_B_DawQzYpX3_2),.clk(gclk));
	jdff dff_B_ckZuosHW4_2(.din(w_dff_B_DawQzYpX3_2),.dout(w_dff_B_ckZuosHW4_2),.clk(gclk));
	jdff dff_B_HEYw3L3e2_2(.din(w_dff_B_ckZuosHW4_2),.dout(w_dff_B_HEYw3L3e2_2),.clk(gclk));
	jdff dff_B_vwTgl1Pe5_2(.din(w_dff_B_HEYw3L3e2_2),.dout(w_dff_B_vwTgl1Pe5_2),.clk(gclk));
	jdff dff_B_S3tY8KDi6_2(.din(w_dff_B_vwTgl1Pe5_2),.dout(w_dff_B_S3tY8KDi6_2),.clk(gclk));
	jdff dff_B_orX2KXrt7_2(.din(w_dff_B_S3tY8KDi6_2),.dout(w_dff_B_orX2KXrt7_2),.clk(gclk));
	jdff dff_B_m7CL91jd0_2(.din(w_dff_B_orX2KXrt7_2),.dout(w_dff_B_m7CL91jd0_2),.clk(gclk));
	jdff dff_B_exGLuhs23_2(.din(w_dff_B_m7CL91jd0_2),.dout(w_dff_B_exGLuhs23_2),.clk(gclk));
	jdff dff_B_GVhOx6UT8_2(.din(w_dff_B_exGLuhs23_2),.dout(w_dff_B_GVhOx6UT8_2),.clk(gclk));
	jdff dff_B_thoognot0_2(.din(w_dff_B_GVhOx6UT8_2),.dout(w_dff_B_thoognot0_2),.clk(gclk));
	jdff dff_B_76CJ4OMI8_2(.din(w_dff_B_thoognot0_2),.dout(w_dff_B_76CJ4OMI8_2),.clk(gclk));
	jdff dff_B_vPIU9umq5_2(.din(w_dff_B_76CJ4OMI8_2),.dout(w_dff_B_vPIU9umq5_2),.clk(gclk));
	jdff dff_B_t2YhdeBC0_2(.din(w_dff_B_vPIU9umq5_2),.dout(w_dff_B_t2YhdeBC0_2),.clk(gclk));
	jdff dff_B_X2BvY5948_2(.din(w_dff_B_t2YhdeBC0_2),.dout(w_dff_B_X2BvY5948_2),.clk(gclk));
	jdff dff_B_0o7XpGAz9_2(.din(n821),.dout(w_dff_B_0o7XpGAz9_2),.clk(gclk));
	jdff dff_B_f52rD6cQ1_1(.din(n743),.dout(w_dff_B_f52rD6cQ1_1),.clk(gclk));
	jdff dff_B_Ez3ezwi98_2(.din(n649),.dout(w_dff_B_Ez3ezwi98_2),.clk(gclk));
	jdff dff_B_DsaySTek7_2(.din(w_dff_B_Ez3ezwi98_2),.dout(w_dff_B_DsaySTek7_2),.clk(gclk));
	jdff dff_B_pASD9vDS0_2(.din(w_dff_B_DsaySTek7_2),.dout(w_dff_B_pASD9vDS0_2),.clk(gclk));
	jdff dff_B_i545mfNE5_2(.din(w_dff_B_pASD9vDS0_2),.dout(w_dff_B_i545mfNE5_2),.clk(gclk));
	jdff dff_B_TEQPCNfb2_2(.din(w_dff_B_i545mfNE5_2),.dout(w_dff_B_TEQPCNfb2_2),.clk(gclk));
	jdff dff_B_QLoZTlQL2_2(.din(w_dff_B_TEQPCNfb2_2),.dout(w_dff_B_QLoZTlQL2_2),.clk(gclk));
	jdff dff_B_gXzPuCI46_2(.din(w_dff_B_QLoZTlQL2_2),.dout(w_dff_B_gXzPuCI46_2),.clk(gclk));
	jdff dff_B_MZSskENs3_2(.din(w_dff_B_gXzPuCI46_2),.dout(w_dff_B_MZSskENs3_2),.clk(gclk));
	jdff dff_B_EbkmuCLV9_2(.din(w_dff_B_MZSskENs3_2),.dout(w_dff_B_EbkmuCLV9_2),.clk(gclk));
	jdff dff_B_uRNj2x3J9_2(.din(w_dff_B_EbkmuCLV9_2),.dout(w_dff_B_uRNj2x3J9_2),.clk(gclk));
	jdff dff_B_GYlkhpAa9_2(.din(w_dff_B_uRNj2x3J9_2),.dout(w_dff_B_GYlkhpAa9_2),.clk(gclk));
	jdff dff_B_wQbd0lRN8_2(.din(w_dff_B_GYlkhpAa9_2),.dout(w_dff_B_wQbd0lRN8_2),.clk(gclk));
	jdff dff_B_5iSkpzgT3_2(.din(w_dff_B_wQbd0lRN8_2),.dout(w_dff_B_5iSkpzgT3_2),.clk(gclk));
	jdff dff_B_85IqjXRi8_2(.din(w_dff_B_5iSkpzgT3_2),.dout(w_dff_B_85IqjXRi8_2),.clk(gclk));
	jdff dff_B_D8MWlv167_2(.din(w_dff_B_85IqjXRi8_2),.dout(w_dff_B_D8MWlv167_2),.clk(gclk));
	jdff dff_B_qcfRUw7a2_2(.din(w_dff_B_D8MWlv167_2),.dout(w_dff_B_qcfRUw7a2_2),.clk(gclk));
	jdff dff_B_KnYwV7Ie8_2(.din(w_dff_B_qcfRUw7a2_2),.dout(w_dff_B_KnYwV7Ie8_2),.clk(gclk));
	jdff dff_B_nY1BbMpL2_2(.din(w_dff_B_KnYwV7Ie8_2),.dout(w_dff_B_nY1BbMpL2_2),.clk(gclk));
	jdff dff_B_xUBq8LUz9_2(.din(w_dff_B_nY1BbMpL2_2),.dout(w_dff_B_xUBq8LUz9_2),.clk(gclk));
	jdff dff_B_2L2fDyKB8_2(.din(w_dff_B_xUBq8LUz9_2),.dout(w_dff_B_2L2fDyKB8_2),.clk(gclk));
	jdff dff_B_mpkc6BD26_2(.din(w_dff_B_2L2fDyKB8_2),.dout(w_dff_B_mpkc6BD26_2),.clk(gclk));
	jdff dff_B_fJUf09Y04_2(.din(w_dff_B_mpkc6BD26_2),.dout(w_dff_B_fJUf09Y04_2),.clk(gclk));
	jdff dff_B_aCiqBmLW9_2(.din(w_dff_B_fJUf09Y04_2),.dout(w_dff_B_aCiqBmLW9_2),.clk(gclk));
	jdff dff_B_EhWBx6Cq5_2(.din(w_dff_B_aCiqBmLW9_2),.dout(w_dff_B_EhWBx6Cq5_2),.clk(gclk));
	jdff dff_B_bwI9yltF0_2(.din(w_dff_B_EhWBx6Cq5_2),.dout(w_dff_B_bwI9yltF0_2),.clk(gclk));
	jdff dff_B_Cp9nh4yP6_2(.din(w_dff_B_bwI9yltF0_2),.dout(w_dff_B_Cp9nh4yP6_2),.clk(gclk));
	jdff dff_B_6KF8uVbC1_2(.din(w_dff_B_Cp9nh4yP6_2),.dout(w_dff_B_6KF8uVbC1_2),.clk(gclk));
	jdff dff_B_Inpf2ij73_2(.din(w_dff_B_6KF8uVbC1_2),.dout(w_dff_B_Inpf2ij73_2),.clk(gclk));
	jdff dff_B_asRicJ5x4_2(.din(w_dff_B_Inpf2ij73_2),.dout(w_dff_B_asRicJ5x4_2),.clk(gclk));
	jdff dff_B_KWMNtjam0_2(.din(w_dff_B_asRicJ5x4_2),.dout(w_dff_B_KWMNtjam0_2),.clk(gclk));
	jdff dff_B_69glCq6x7_2(.din(w_dff_B_KWMNtjam0_2),.dout(w_dff_B_69glCq6x7_2),.clk(gclk));
	jdff dff_B_G3QqpJfF0_2(.din(n721),.dout(w_dff_B_G3QqpJfF0_2),.clk(gclk));
	jdff dff_B_X9AQeE1F8_1(.din(n650),.dout(w_dff_B_X9AQeE1F8_1),.clk(gclk));
	jdff dff_B_Srme0Lsp1_2(.din(n563),.dout(w_dff_B_Srme0Lsp1_2),.clk(gclk));
	jdff dff_B_MCA5sysm1_2(.din(w_dff_B_Srme0Lsp1_2),.dout(w_dff_B_MCA5sysm1_2),.clk(gclk));
	jdff dff_B_JC33sl7w7_2(.din(w_dff_B_MCA5sysm1_2),.dout(w_dff_B_JC33sl7w7_2),.clk(gclk));
	jdff dff_B_MESuZzuJ8_2(.din(w_dff_B_JC33sl7w7_2),.dout(w_dff_B_MESuZzuJ8_2),.clk(gclk));
	jdff dff_B_UYbyn5cS6_2(.din(w_dff_B_MESuZzuJ8_2),.dout(w_dff_B_UYbyn5cS6_2),.clk(gclk));
	jdff dff_B_0bZi3Wt47_2(.din(w_dff_B_UYbyn5cS6_2),.dout(w_dff_B_0bZi3Wt47_2),.clk(gclk));
	jdff dff_B_MV0H9icV7_2(.din(w_dff_B_0bZi3Wt47_2),.dout(w_dff_B_MV0H9icV7_2),.clk(gclk));
	jdff dff_B_c9VWh5OX0_2(.din(w_dff_B_MV0H9icV7_2),.dout(w_dff_B_c9VWh5OX0_2),.clk(gclk));
	jdff dff_B_rXITN77F3_2(.din(w_dff_B_c9VWh5OX0_2),.dout(w_dff_B_rXITN77F3_2),.clk(gclk));
	jdff dff_B_wUOv5E3n4_2(.din(w_dff_B_rXITN77F3_2),.dout(w_dff_B_wUOv5E3n4_2),.clk(gclk));
	jdff dff_B_wlul32NE4_2(.din(w_dff_B_wUOv5E3n4_2),.dout(w_dff_B_wlul32NE4_2),.clk(gclk));
	jdff dff_B_l6YuJYHl6_2(.din(w_dff_B_wlul32NE4_2),.dout(w_dff_B_l6YuJYHl6_2),.clk(gclk));
	jdff dff_B_MISHKE7b1_2(.din(w_dff_B_l6YuJYHl6_2),.dout(w_dff_B_MISHKE7b1_2),.clk(gclk));
	jdff dff_B_tbDNQlhJ1_2(.din(w_dff_B_MISHKE7b1_2),.dout(w_dff_B_tbDNQlhJ1_2),.clk(gclk));
	jdff dff_B_6DlFXdW13_2(.din(w_dff_B_tbDNQlhJ1_2),.dout(w_dff_B_6DlFXdW13_2),.clk(gclk));
	jdff dff_B_jrn2BW7N3_2(.din(w_dff_B_6DlFXdW13_2),.dout(w_dff_B_jrn2BW7N3_2),.clk(gclk));
	jdff dff_B_opw29W1Y4_2(.din(w_dff_B_jrn2BW7N3_2),.dout(w_dff_B_opw29W1Y4_2),.clk(gclk));
	jdff dff_B_sKks8iMG7_2(.din(w_dff_B_opw29W1Y4_2),.dout(w_dff_B_sKks8iMG7_2),.clk(gclk));
	jdff dff_B_EAIjP8xk8_2(.din(w_dff_B_sKks8iMG7_2),.dout(w_dff_B_EAIjP8xk8_2),.clk(gclk));
	jdff dff_B_ksWvyQwx3_2(.din(w_dff_B_EAIjP8xk8_2),.dout(w_dff_B_ksWvyQwx3_2),.clk(gclk));
	jdff dff_B_QcLFNgqx4_2(.din(w_dff_B_ksWvyQwx3_2),.dout(w_dff_B_QcLFNgqx4_2),.clk(gclk));
	jdff dff_B_A2PWGXGY4_2(.din(w_dff_B_QcLFNgqx4_2),.dout(w_dff_B_A2PWGXGY4_2),.clk(gclk));
	jdff dff_B_SKACZcwk2_2(.din(w_dff_B_A2PWGXGY4_2),.dout(w_dff_B_SKACZcwk2_2),.clk(gclk));
	jdff dff_B_8Ade8wf23_2(.din(w_dff_B_SKACZcwk2_2),.dout(w_dff_B_8Ade8wf23_2),.clk(gclk));
	jdff dff_B_AiBGui6H6_2(.din(w_dff_B_8Ade8wf23_2),.dout(w_dff_B_AiBGui6H6_2),.clk(gclk));
	jdff dff_B_xZoxIi9v4_2(.din(w_dff_B_AiBGui6H6_2),.dout(w_dff_B_xZoxIi9v4_2),.clk(gclk));
	jdff dff_B_bx3pvt1y4_2(.din(w_dff_B_xZoxIi9v4_2),.dout(w_dff_B_bx3pvt1y4_2),.clk(gclk));
	jdff dff_B_OO7HPbty9_2(.din(w_dff_B_bx3pvt1y4_2),.dout(w_dff_B_OO7HPbty9_2),.clk(gclk));
	jdff dff_B_WD6Ur2R19_2(.din(n628),.dout(w_dff_B_WD6Ur2R19_2),.clk(gclk));
	jdff dff_B_zFuVlLZs2_1(.din(n564),.dout(w_dff_B_zFuVlLZs2_1),.clk(gclk));
	jdff dff_B_fWL7QoAV2_2(.din(n484),.dout(w_dff_B_fWL7QoAV2_2),.clk(gclk));
	jdff dff_B_NrMuFbNg8_2(.din(w_dff_B_fWL7QoAV2_2),.dout(w_dff_B_NrMuFbNg8_2),.clk(gclk));
	jdff dff_B_614uzick1_2(.din(w_dff_B_NrMuFbNg8_2),.dout(w_dff_B_614uzick1_2),.clk(gclk));
	jdff dff_B_1TKcZNRU7_2(.din(w_dff_B_614uzick1_2),.dout(w_dff_B_1TKcZNRU7_2),.clk(gclk));
	jdff dff_B_Ak6k3QKo9_2(.din(w_dff_B_1TKcZNRU7_2),.dout(w_dff_B_Ak6k3QKo9_2),.clk(gclk));
	jdff dff_B_9s2dY15T7_2(.din(w_dff_B_Ak6k3QKo9_2),.dout(w_dff_B_9s2dY15T7_2),.clk(gclk));
	jdff dff_B_49VkbSUp9_2(.din(w_dff_B_9s2dY15T7_2),.dout(w_dff_B_49VkbSUp9_2),.clk(gclk));
	jdff dff_B_d6MHqYF23_2(.din(w_dff_B_49VkbSUp9_2),.dout(w_dff_B_d6MHqYF23_2),.clk(gclk));
	jdff dff_B_JeWNfWkH0_2(.din(w_dff_B_d6MHqYF23_2),.dout(w_dff_B_JeWNfWkH0_2),.clk(gclk));
	jdff dff_B_srGNjmG24_2(.din(w_dff_B_JeWNfWkH0_2),.dout(w_dff_B_srGNjmG24_2),.clk(gclk));
	jdff dff_B_x9Ddx2Xm5_2(.din(w_dff_B_srGNjmG24_2),.dout(w_dff_B_x9Ddx2Xm5_2),.clk(gclk));
	jdff dff_B_3TTVyZJ61_2(.din(w_dff_B_x9Ddx2Xm5_2),.dout(w_dff_B_3TTVyZJ61_2),.clk(gclk));
	jdff dff_B_id4z2nxo8_2(.din(w_dff_B_3TTVyZJ61_2),.dout(w_dff_B_id4z2nxo8_2),.clk(gclk));
	jdff dff_B_hOGl5MEE6_2(.din(w_dff_B_id4z2nxo8_2),.dout(w_dff_B_hOGl5MEE6_2),.clk(gclk));
	jdff dff_B_dx61HIkF0_2(.din(w_dff_B_hOGl5MEE6_2),.dout(w_dff_B_dx61HIkF0_2),.clk(gclk));
	jdff dff_B_EdzsSPAA7_2(.din(w_dff_B_dx61HIkF0_2),.dout(w_dff_B_EdzsSPAA7_2),.clk(gclk));
	jdff dff_B_zarxGLFy5_2(.din(w_dff_B_EdzsSPAA7_2),.dout(w_dff_B_zarxGLFy5_2),.clk(gclk));
	jdff dff_B_GnEUns0H7_2(.din(w_dff_B_zarxGLFy5_2),.dout(w_dff_B_GnEUns0H7_2),.clk(gclk));
	jdff dff_B_HvH16jII8_2(.din(w_dff_B_GnEUns0H7_2),.dout(w_dff_B_HvH16jII8_2),.clk(gclk));
	jdff dff_B_VwjtGjNL9_2(.din(w_dff_B_HvH16jII8_2),.dout(w_dff_B_VwjtGjNL9_2),.clk(gclk));
	jdff dff_B_HUK9nZOo4_2(.din(w_dff_B_VwjtGjNL9_2),.dout(w_dff_B_HUK9nZOo4_2),.clk(gclk));
	jdff dff_B_RUlh8mkv9_2(.din(w_dff_B_HUK9nZOo4_2),.dout(w_dff_B_RUlh8mkv9_2),.clk(gclk));
	jdff dff_B_y449ZoZd7_2(.din(w_dff_B_RUlh8mkv9_2),.dout(w_dff_B_y449ZoZd7_2),.clk(gclk));
	jdff dff_B_qTjIi8T84_2(.din(w_dff_B_y449ZoZd7_2),.dout(w_dff_B_qTjIi8T84_2),.clk(gclk));
	jdff dff_B_ukBH0eR21_2(.din(w_dff_B_qTjIi8T84_2),.dout(w_dff_B_ukBH0eR21_2),.clk(gclk));
	jdff dff_B_PlMEJB0o9_2(.din(n542),.dout(w_dff_B_PlMEJB0o9_2),.clk(gclk));
	jdff dff_B_cQqrFy9q4_1(.din(n485),.dout(w_dff_B_cQqrFy9q4_1),.clk(gclk));
	jdff dff_B_oGXZN2S17_2(.din(n412),.dout(w_dff_B_oGXZN2S17_2),.clk(gclk));
	jdff dff_B_dcmPLmwV5_2(.din(w_dff_B_oGXZN2S17_2),.dout(w_dff_B_dcmPLmwV5_2),.clk(gclk));
	jdff dff_B_OY363PeA3_2(.din(w_dff_B_dcmPLmwV5_2),.dout(w_dff_B_OY363PeA3_2),.clk(gclk));
	jdff dff_B_84f9GGzJ0_2(.din(w_dff_B_OY363PeA3_2),.dout(w_dff_B_84f9GGzJ0_2),.clk(gclk));
	jdff dff_B_wTdFwfpJ7_2(.din(w_dff_B_84f9GGzJ0_2),.dout(w_dff_B_wTdFwfpJ7_2),.clk(gclk));
	jdff dff_B_afeorywH9_2(.din(w_dff_B_wTdFwfpJ7_2),.dout(w_dff_B_afeorywH9_2),.clk(gclk));
	jdff dff_B_qEeyTEU21_2(.din(w_dff_B_afeorywH9_2),.dout(w_dff_B_qEeyTEU21_2),.clk(gclk));
	jdff dff_B_hmjmKlc68_2(.din(w_dff_B_qEeyTEU21_2),.dout(w_dff_B_hmjmKlc68_2),.clk(gclk));
	jdff dff_B_hfJE7aeS1_2(.din(w_dff_B_hmjmKlc68_2),.dout(w_dff_B_hfJE7aeS1_2),.clk(gclk));
	jdff dff_B_SEGgKQXj4_2(.din(w_dff_B_hfJE7aeS1_2),.dout(w_dff_B_SEGgKQXj4_2),.clk(gclk));
	jdff dff_B_YSbcQQLq3_2(.din(w_dff_B_SEGgKQXj4_2),.dout(w_dff_B_YSbcQQLq3_2),.clk(gclk));
	jdff dff_B_Z1dCurid3_2(.din(w_dff_B_YSbcQQLq3_2),.dout(w_dff_B_Z1dCurid3_2),.clk(gclk));
	jdff dff_B_8nG992SQ6_2(.din(w_dff_B_Z1dCurid3_2),.dout(w_dff_B_8nG992SQ6_2),.clk(gclk));
	jdff dff_B_DupaHDwX9_2(.din(w_dff_B_8nG992SQ6_2),.dout(w_dff_B_DupaHDwX9_2),.clk(gclk));
	jdff dff_B_MrsWqR4A0_2(.din(w_dff_B_DupaHDwX9_2),.dout(w_dff_B_MrsWqR4A0_2),.clk(gclk));
	jdff dff_B_DTPpgtrK7_2(.din(w_dff_B_MrsWqR4A0_2),.dout(w_dff_B_DTPpgtrK7_2),.clk(gclk));
	jdff dff_B_AqPc4pSF0_2(.din(w_dff_B_DTPpgtrK7_2),.dout(w_dff_B_AqPc4pSF0_2),.clk(gclk));
	jdff dff_B_AN0G1K7T0_2(.din(w_dff_B_AqPc4pSF0_2),.dout(w_dff_B_AN0G1K7T0_2),.clk(gclk));
	jdff dff_B_PPoL0E3m5_2(.din(w_dff_B_AN0G1K7T0_2),.dout(w_dff_B_PPoL0E3m5_2),.clk(gclk));
	jdff dff_B_bnRtv1O20_2(.din(w_dff_B_PPoL0E3m5_2),.dout(w_dff_B_bnRtv1O20_2),.clk(gclk));
	jdff dff_B_5oHCXnj42_2(.din(w_dff_B_bnRtv1O20_2),.dout(w_dff_B_5oHCXnj42_2),.clk(gclk));
	jdff dff_B_vJ5JRxYC2_2(.din(w_dff_B_5oHCXnj42_2),.dout(w_dff_B_vJ5JRxYC2_2),.clk(gclk));
	jdff dff_B_Moc7km7x7_2(.din(n463),.dout(w_dff_B_Moc7km7x7_2),.clk(gclk));
	jdff dff_B_vkyvK0Dy8_1(.din(n413),.dout(w_dff_B_vkyvK0Dy8_1),.clk(gclk));
	jdff dff_B_YDiGq3YV8_2(.din(n348),.dout(w_dff_B_YDiGq3YV8_2),.clk(gclk));
	jdff dff_B_1fbf1D4U9_2(.din(w_dff_B_YDiGq3YV8_2),.dout(w_dff_B_1fbf1D4U9_2),.clk(gclk));
	jdff dff_B_OGMxSz1Z2_2(.din(w_dff_B_1fbf1D4U9_2),.dout(w_dff_B_OGMxSz1Z2_2),.clk(gclk));
	jdff dff_B_1NxLQ00i4_2(.din(w_dff_B_OGMxSz1Z2_2),.dout(w_dff_B_1NxLQ00i4_2),.clk(gclk));
	jdff dff_B_5onlD2pa3_2(.din(w_dff_B_1NxLQ00i4_2),.dout(w_dff_B_5onlD2pa3_2),.clk(gclk));
	jdff dff_B_PQcHEGID9_2(.din(w_dff_B_5onlD2pa3_2),.dout(w_dff_B_PQcHEGID9_2),.clk(gclk));
	jdff dff_B_9CQLLmy53_2(.din(w_dff_B_PQcHEGID9_2),.dout(w_dff_B_9CQLLmy53_2),.clk(gclk));
	jdff dff_B_WSfaPRf54_2(.din(w_dff_B_9CQLLmy53_2),.dout(w_dff_B_WSfaPRf54_2),.clk(gclk));
	jdff dff_B_8IVexXC99_2(.din(w_dff_B_WSfaPRf54_2),.dout(w_dff_B_8IVexXC99_2),.clk(gclk));
	jdff dff_B_CwI58KiC7_2(.din(w_dff_B_8IVexXC99_2),.dout(w_dff_B_CwI58KiC7_2),.clk(gclk));
	jdff dff_B_1alBs9ag3_2(.din(w_dff_B_CwI58KiC7_2),.dout(w_dff_B_1alBs9ag3_2),.clk(gclk));
	jdff dff_B_sRYweDbj3_2(.din(w_dff_B_1alBs9ag3_2),.dout(w_dff_B_sRYweDbj3_2),.clk(gclk));
	jdff dff_B_gwIHCuXq4_2(.din(w_dff_B_sRYweDbj3_2),.dout(w_dff_B_gwIHCuXq4_2),.clk(gclk));
	jdff dff_B_O8NHjyGe1_2(.din(w_dff_B_gwIHCuXq4_2),.dout(w_dff_B_O8NHjyGe1_2),.clk(gclk));
	jdff dff_B_tn5qo77Q2_2(.din(w_dff_B_O8NHjyGe1_2),.dout(w_dff_B_tn5qo77Q2_2),.clk(gclk));
	jdff dff_B_2qljnYKr5_2(.din(w_dff_B_tn5qo77Q2_2),.dout(w_dff_B_2qljnYKr5_2),.clk(gclk));
	jdff dff_B_6lOs4cgo8_2(.din(w_dff_B_2qljnYKr5_2),.dout(w_dff_B_6lOs4cgo8_2),.clk(gclk));
	jdff dff_B_ei6UQS5s0_2(.din(w_dff_B_6lOs4cgo8_2),.dout(w_dff_B_ei6UQS5s0_2),.clk(gclk));
	jdff dff_B_InpKIDaf8_2(.din(w_dff_B_ei6UQS5s0_2),.dout(w_dff_B_InpKIDaf8_2),.clk(gclk));
	jdff dff_B_Cv00onWb5_2(.din(n391),.dout(w_dff_B_Cv00onWb5_2),.clk(gclk));
	jdff dff_B_KohjZSWe6_1(.din(n349),.dout(w_dff_B_KohjZSWe6_1),.clk(gclk));
	jdff dff_B_9RCnqk8y0_2(.din(n290),.dout(w_dff_B_9RCnqk8y0_2),.clk(gclk));
	jdff dff_B_kkfzAReT7_2(.din(w_dff_B_9RCnqk8y0_2),.dout(w_dff_B_kkfzAReT7_2),.clk(gclk));
	jdff dff_B_8dxjvqVf7_2(.din(w_dff_B_kkfzAReT7_2),.dout(w_dff_B_8dxjvqVf7_2),.clk(gclk));
	jdff dff_B_Ktm2YA779_2(.din(w_dff_B_8dxjvqVf7_2),.dout(w_dff_B_Ktm2YA779_2),.clk(gclk));
	jdff dff_B_f58Lg4jI1_2(.din(w_dff_B_Ktm2YA779_2),.dout(w_dff_B_f58Lg4jI1_2),.clk(gclk));
	jdff dff_B_3xP7YiDt0_2(.din(w_dff_B_f58Lg4jI1_2),.dout(w_dff_B_3xP7YiDt0_2),.clk(gclk));
	jdff dff_B_MjApJ2Ef2_2(.din(w_dff_B_3xP7YiDt0_2),.dout(w_dff_B_MjApJ2Ef2_2),.clk(gclk));
	jdff dff_B_RYj4j7GR7_2(.din(w_dff_B_MjApJ2Ef2_2),.dout(w_dff_B_RYj4j7GR7_2),.clk(gclk));
	jdff dff_B_JN8Rmjbu0_2(.din(w_dff_B_RYj4j7GR7_2),.dout(w_dff_B_JN8Rmjbu0_2),.clk(gclk));
	jdff dff_B_Zwgq2YQn4_2(.din(w_dff_B_JN8Rmjbu0_2),.dout(w_dff_B_Zwgq2YQn4_2),.clk(gclk));
	jdff dff_B_Qvv4S3gL1_2(.din(w_dff_B_Zwgq2YQn4_2),.dout(w_dff_B_Qvv4S3gL1_2),.clk(gclk));
	jdff dff_B_tXkMbQqq4_2(.din(w_dff_B_Qvv4S3gL1_2),.dout(w_dff_B_tXkMbQqq4_2),.clk(gclk));
	jdff dff_B_ItELkwND8_2(.din(w_dff_B_tXkMbQqq4_2),.dout(w_dff_B_ItELkwND8_2),.clk(gclk));
	jdff dff_B_7emjLOGz8_2(.din(w_dff_B_ItELkwND8_2),.dout(w_dff_B_7emjLOGz8_2),.clk(gclk));
	jdff dff_B_San30miK3_2(.din(w_dff_B_7emjLOGz8_2),.dout(w_dff_B_San30miK3_2),.clk(gclk));
	jdff dff_B_KvgfoixZ0_2(.din(w_dff_B_San30miK3_2),.dout(w_dff_B_KvgfoixZ0_2),.clk(gclk));
	jdff dff_B_otGOyUp50_2(.din(n327),.dout(w_dff_B_otGOyUp50_2),.clk(gclk));
	jdff dff_B_93cARDKC8_1(.din(n291),.dout(w_dff_B_93cARDKC8_1),.clk(gclk));
	jdff dff_B_0zxOQWab8_2(.din(n239),.dout(w_dff_B_0zxOQWab8_2),.clk(gclk));
	jdff dff_B_NB1dVVAN1_2(.din(w_dff_B_0zxOQWab8_2),.dout(w_dff_B_NB1dVVAN1_2),.clk(gclk));
	jdff dff_B_TY4KntTa0_2(.din(w_dff_B_NB1dVVAN1_2),.dout(w_dff_B_TY4KntTa0_2),.clk(gclk));
	jdff dff_B_1uek05gj7_2(.din(w_dff_B_TY4KntTa0_2),.dout(w_dff_B_1uek05gj7_2),.clk(gclk));
	jdff dff_B_nB2cmqc60_2(.din(w_dff_B_1uek05gj7_2),.dout(w_dff_B_nB2cmqc60_2),.clk(gclk));
	jdff dff_B_BFGcQ4OJ9_2(.din(w_dff_B_nB2cmqc60_2),.dout(w_dff_B_BFGcQ4OJ9_2),.clk(gclk));
	jdff dff_B_9pq8nSal8_2(.din(w_dff_B_BFGcQ4OJ9_2),.dout(w_dff_B_9pq8nSal8_2),.clk(gclk));
	jdff dff_B_i2pGKpnn3_2(.din(w_dff_B_9pq8nSal8_2),.dout(w_dff_B_i2pGKpnn3_2),.clk(gclk));
	jdff dff_B_XQCe5YRT3_2(.din(w_dff_B_i2pGKpnn3_2),.dout(w_dff_B_XQCe5YRT3_2),.clk(gclk));
	jdff dff_B_OlLvvtdM3_2(.din(w_dff_B_XQCe5YRT3_2),.dout(w_dff_B_OlLvvtdM3_2),.clk(gclk));
	jdff dff_B_ddhbREas5_2(.din(w_dff_B_OlLvvtdM3_2),.dout(w_dff_B_ddhbREas5_2),.clk(gclk));
	jdff dff_B_lDmu6JHi8_2(.din(w_dff_B_ddhbREas5_2),.dout(w_dff_B_lDmu6JHi8_2),.clk(gclk));
	jdff dff_B_z2IB3KoP5_2(.din(w_dff_B_lDmu6JHi8_2),.dout(w_dff_B_z2IB3KoP5_2),.clk(gclk));
	jdff dff_B_lNc23o2r7_2(.din(n269),.dout(w_dff_B_lNc23o2r7_2),.clk(gclk));
	jdff dff_B_Q7T7t4QA3_1(.din(n240),.dout(w_dff_B_Q7T7t4QA3_1),.clk(gclk));
	jdff dff_B_d10n6hdY6_2(.din(n196),.dout(w_dff_B_d10n6hdY6_2),.clk(gclk));
	jdff dff_B_vwJ3UIP02_2(.din(w_dff_B_d10n6hdY6_2),.dout(w_dff_B_vwJ3UIP02_2),.clk(gclk));
	jdff dff_B_kCJ6zncB5_2(.din(w_dff_B_vwJ3UIP02_2),.dout(w_dff_B_kCJ6zncB5_2),.clk(gclk));
	jdff dff_B_sQywHaUr9_2(.din(w_dff_B_kCJ6zncB5_2),.dout(w_dff_B_sQywHaUr9_2),.clk(gclk));
	jdff dff_B_pbbOhqe95_2(.din(w_dff_B_sQywHaUr9_2),.dout(w_dff_B_pbbOhqe95_2),.clk(gclk));
	jdff dff_B_TdgP8NmY8_2(.din(w_dff_B_pbbOhqe95_2),.dout(w_dff_B_TdgP8NmY8_2),.clk(gclk));
	jdff dff_B_fZMRQ7B03_2(.din(w_dff_B_TdgP8NmY8_2),.dout(w_dff_B_fZMRQ7B03_2),.clk(gclk));
	jdff dff_B_8WR5SiN83_2(.din(w_dff_B_fZMRQ7B03_2),.dout(w_dff_B_8WR5SiN83_2),.clk(gclk));
	jdff dff_B_SWtnxoTH5_2(.din(w_dff_B_8WR5SiN83_2),.dout(w_dff_B_SWtnxoTH5_2),.clk(gclk));
	jdff dff_B_SL8ZdoEa6_2(.din(w_dff_B_SWtnxoTH5_2),.dout(w_dff_B_SL8ZdoEa6_2),.clk(gclk));
	jdff dff_B_BwpPDbDd4_2(.din(n218),.dout(w_dff_B_BwpPDbDd4_2),.clk(gclk));
	jdff dff_B_rb5e9BaE9_1(.din(n197),.dout(w_dff_B_rb5e9BaE9_1),.clk(gclk));
	jdff dff_B_93yd9Np29_2(.din(n158),.dout(w_dff_B_93yd9Np29_2),.clk(gclk));
	jdff dff_B_KNPyR0fw0_2(.din(w_dff_B_93yd9Np29_2),.dout(w_dff_B_KNPyR0fw0_2),.clk(gclk));
	jdff dff_B_VUCyno7I9_2(.din(w_dff_B_KNPyR0fw0_2),.dout(w_dff_B_VUCyno7I9_2),.clk(gclk));
	jdff dff_B_ByoylkFx9_2(.din(w_dff_B_VUCyno7I9_2),.dout(w_dff_B_ByoylkFx9_2),.clk(gclk));
	jdff dff_B_FKoK8ueI5_2(.din(w_dff_B_ByoylkFx9_2),.dout(w_dff_B_FKoK8ueI5_2),.clk(gclk));
	jdff dff_B_wHPEqHOf6_2(.din(w_dff_B_FKoK8ueI5_2),.dout(w_dff_B_wHPEqHOf6_2),.clk(gclk));
	jdff dff_B_6WHuhTtx4_2(.din(w_dff_B_wHPEqHOf6_2),.dout(w_dff_B_6WHuhTtx4_2),.clk(gclk));
	jdff dff_B_CZmZ4Z1s3_2(.din(n175),.dout(w_dff_B_CZmZ4Z1s3_2),.clk(gclk));
	jdff dff_B_C0xixdSd6_1(.din(n161),.dout(w_dff_B_C0xixdSd6_1),.clk(gclk));
	jdff dff_B_CJuuASMf2_1(.din(w_dff_B_C0xixdSd6_1),.dout(w_dff_B_CJuuASMf2_1),.clk(gclk));
	jdff dff_B_TFIA9FbN7_2(.din(n128),.dout(w_dff_B_TFIA9FbN7_2),.clk(gclk));
	jdff dff_B_nx8LWBXN6_2(.din(w_dff_B_TFIA9FbN7_2),.dout(w_dff_B_nx8LWBXN6_2),.clk(gclk));
	jdff dff_B_7FwG0O9p1_2(.din(w_dff_B_nx8LWBXN6_2),.dout(w_dff_B_7FwG0O9p1_2),.clk(gclk));
	jdff dff_B_LmbkEhOm2_2(.din(w_dff_B_7FwG0O9p1_2),.dout(w_dff_B_LmbkEhOm2_2),.clk(gclk));
	jdff dff_A_kaDeBZSS5_1(.dout(w_n130_0[1]),.din(w_dff_A_kaDeBZSS5_1),.clk(gclk));
	jdff dff_A_jIE5RpNV8_0(.dout(w_n101_0[0]),.din(w_dff_A_jIE5RpNV8_0),.clk(gclk));
	jdff dff_A_wRGR6vxt7_0(.dout(w_n100_1[0]),.din(w_dff_A_wRGR6vxt7_0),.clk(gclk));
	jdff dff_A_IqkzQ5Xs0_1(.dout(w_n100_0[1]),.din(w_dff_A_IqkzQ5Xs0_1),.clk(gclk));
	jdff dff_A_iZRBN08a4_2(.dout(w_n100_0[2]),.din(w_dff_A_iZRBN08a4_2),.clk(gclk));
	jdff dff_A_Z0PxXlJi4_2(.dout(w_dff_A_iZRBN08a4_2),.din(w_dff_A_Z0PxXlJi4_2),.clk(gclk));
	jdff dff_B_urI1xCRA6_0(.din(n1329),.dout(w_dff_B_urI1xCRA6_0),.clk(gclk));
	jdff dff_A_9iBBkNyV8_1(.dout(w_n1325_0[1]),.din(w_dff_A_9iBBkNyV8_1),.clk(gclk));
	jdff dff_A_YmfkltVR9_1(.dout(w_dff_A_9iBBkNyV8_1),.din(w_dff_A_YmfkltVR9_1),.clk(gclk));
	jdff dff_B_X81WlWxz2_1(.din(n1245),.dout(w_dff_B_X81WlWxz2_1),.clk(gclk));
	jdff dff_B_RMb7G1lh3_1(.din(w_dff_B_X81WlWxz2_1),.dout(w_dff_B_RMb7G1lh3_1),.clk(gclk));
	jdff dff_B_jhpcgWXj2_2(.din(n1152),.dout(w_dff_B_jhpcgWXj2_2),.clk(gclk));
	jdff dff_B_EcjBM6v66_2(.din(w_dff_B_jhpcgWXj2_2),.dout(w_dff_B_EcjBM6v66_2),.clk(gclk));
	jdff dff_B_MzH7DKhg3_2(.din(w_dff_B_EcjBM6v66_2),.dout(w_dff_B_MzH7DKhg3_2),.clk(gclk));
	jdff dff_B_uzJEh9QK8_2(.din(w_dff_B_MzH7DKhg3_2),.dout(w_dff_B_uzJEh9QK8_2),.clk(gclk));
	jdff dff_B_fwHIOZsQ5_2(.din(w_dff_B_uzJEh9QK8_2),.dout(w_dff_B_fwHIOZsQ5_2),.clk(gclk));
	jdff dff_B_TzEie9ks1_2(.din(w_dff_B_fwHIOZsQ5_2),.dout(w_dff_B_TzEie9ks1_2),.clk(gclk));
	jdff dff_B_I9yRw00K5_2(.din(w_dff_B_TzEie9ks1_2),.dout(w_dff_B_I9yRw00K5_2),.clk(gclk));
	jdff dff_B_feK24Jrs0_2(.din(w_dff_B_I9yRw00K5_2),.dout(w_dff_B_feK24Jrs0_2),.clk(gclk));
	jdff dff_B_55uPTe7i2_2(.din(w_dff_B_feK24Jrs0_2),.dout(w_dff_B_55uPTe7i2_2),.clk(gclk));
	jdff dff_B_R1CqWste0_2(.din(w_dff_B_55uPTe7i2_2),.dout(w_dff_B_R1CqWste0_2),.clk(gclk));
	jdff dff_B_09BZpA1C9_2(.din(w_dff_B_R1CqWste0_2),.dout(w_dff_B_09BZpA1C9_2),.clk(gclk));
	jdff dff_B_s6E45NDp1_2(.din(w_dff_B_09BZpA1C9_2),.dout(w_dff_B_s6E45NDp1_2),.clk(gclk));
	jdff dff_B_UcicT4r90_2(.din(w_dff_B_s6E45NDp1_2),.dout(w_dff_B_UcicT4r90_2),.clk(gclk));
	jdff dff_B_0oW87VPB8_2(.din(w_dff_B_UcicT4r90_2),.dout(w_dff_B_0oW87VPB8_2),.clk(gclk));
	jdff dff_B_D2OBaIQS0_2(.din(w_dff_B_0oW87VPB8_2),.dout(w_dff_B_D2OBaIQS0_2),.clk(gclk));
	jdff dff_B_wm7YZmGz4_2(.din(w_dff_B_D2OBaIQS0_2),.dout(w_dff_B_wm7YZmGz4_2),.clk(gclk));
	jdff dff_B_SqgLxptV8_2(.din(w_dff_B_wm7YZmGz4_2),.dout(w_dff_B_SqgLxptV8_2),.clk(gclk));
	jdff dff_B_M49xPGwf2_2(.din(w_dff_B_SqgLxptV8_2),.dout(w_dff_B_M49xPGwf2_2),.clk(gclk));
	jdff dff_B_f6DXcH6h7_2(.din(w_dff_B_M49xPGwf2_2),.dout(w_dff_B_f6DXcH6h7_2),.clk(gclk));
	jdff dff_B_0OHa1wGY5_2(.din(w_dff_B_f6DXcH6h7_2),.dout(w_dff_B_0OHa1wGY5_2),.clk(gclk));
	jdff dff_B_Hygmnn8X4_2(.din(w_dff_B_0OHa1wGY5_2),.dout(w_dff_B_Hygmnn8X4_2),.clk(gclk));
	jdff dff_B_5BfroobQ8_2(.din(w_dff_B_Hygmnn8X4_2),.dout(w_dff_B_5BfroobQ8_2),.clk(gclk));
	jdff dff_B_gac5Wmuo4_2(.din(w_dff_B_5BfroobQ8_2),.dout(w_dff_B_gac5Wmuo4_2),.clk(gclk));
	jdff dff_B_M0PEp5102_2(.din(w_dff_B_gac5Wmuo4_2),.dout(w_dff_B_M0PEp5102_2),.clk(gclk));
	jdff dff_B_3gsk11nK3_2(.din(w_dff_B_M0PEp5102_2),.dout(w_dff_B_3gsk11nK3_2),.clk(gclk));
	jdff dff_B_rY1cNEMX2_2(.din(w_dff_B_3gsk11nK3_2),.dout(w_dff_B_rY1cNEMX2_2),.clk(gclk));
	jdff dff_B_1vGEAePT3_2(.din(w_dff_B_rY1cNEMX2_2),.dout(w_dff_B_1vGEAePT3_2),.clk(gclk));
	jdff dff_B_f3np73zH5_2(.din(w_dff_B_1vGEAePT3_2),.dout(w_dff_B_f3np73zH5_2),.clk(gclk));
	jdff dff_B_iDjT3xKg4_2(.din(w_dff_B_f3np73zH5_2),.dout(w_dff_B_iDjT3xKg4_2),.clk(gclk));
	jdff dff_B_eNsimHCv9_2(.din(w_dff_B_iDjT3xKg4_2),.dout(w_dff_B_eNsimHCv9_2),.clk(gclk));
	jdff dff_B_LQ0INL6c9_2(.din(w_dff_B_eNsimHCv9_2),.dout(w_dff_B_LQ0INL6c9_2),.clk(gclk));
	jdff dff_B_x27H9P4l9_2(.din(w_dff_B_LQ0INL6c9_2),.dout(w_dff_B_x27H9P4l9_2),.clk(gclk));
	jdff dff_B_oXeVwatv8_2(.din(w_dff_B_x27H9P4l9_2),.dout(w_dff_B_oXeVwatv8_2),.clk(gclk));
	jdff dff_B_qlOvGnHU8_2(.din(w_dff_B_oXeVwatv8_2),.dout(w_dff_B_qlOvGnHU8_2),.clk(gclk));
	jdff dff_B_d7us3JCG8_2(.din(w_dff_B_qlOvGnHU8_2),.dout(w_dff_B_d7us3JCG8_2),.clk(gclk));
	jdff dff_B_tZXwgX9O2_2(.din(w_dff_B_d7us3JCG8_2),.dout(w_dff_B_tZXwgX9O2_2),.clk(gclk));
	jdff dff_B_ecgv8P0H5_2(.din(w_dff_B_tZXwgX9O2_2),.dout(w_dff_B_ecgv8P0H5_2),.clk(gclk));
	jdff dff_B_7SBnluyj4_2(.din(w_dff_B_ecgv8P0H5_2),.dout(w_dff_B_7SBnluyj4_2),.clk(gclk));
	jdff dff_B_jCILsPOp8_2(.din(w_dff_B_7SBnluyj4_2),.dout(w_dff_B_jCILsPOp8_2),.clk(gclk));
	jdff dff_B_4UOyRuZP9_2(.din(w_dff_B_jCILsPOp8_2),.dout(w_dff_B_4UOyRuZP9_2),.clk(gclk));
	jdff dff_B_dkaREQ6B8_2(.din(w_dff_B_4UOyRuZP9_2),.dout(w_dff_B_dkaREQ6B8_2),.clk(gclk));
	jdff dff_B_xiS8vVXY8_2(.din(w_dff_B_dkaREQ6B8_2),.dout(w_dff_B_xiS8vVXY8_2),.clk(gclk));
	jdff dff_B_mfTSQzP12_2(.din(w_dff_B_xiS8vVXY8_2),.dout(w_dff_B_mfTSQzP12_2),.clk(gclk));
	jdff dff_B_6M2XYg5C5_2(.din(w_dff_B_mfTSQzP12_2),.dout(w_dff_B_6M2XYg5C5_2),.clk(gclk));
	jdff dff_B_HyFIu3p40_2(.din(w_dff_B_6M2XYg5C5_2),.dout(w_dff_B_HyFIu3p40_2),.clk(gclk));
	jdff dff_B_OFFb5aQu2_2(.din(w_dff_B_HyFIu3p40_2),.dout(w_dff_B_OFFb5aQu2_2),.clk(gclk));
	jdff dff_B_QyiOm4660_2(.din(n1234),.dout(w_dff_B_QyiOm4660_2),.clk(gclk));
	jdff dff_B_SnrhP7B65_1(.din(n1154),.dout(w_dff_B_SnrhP7B65_1),.clk(gclk));
	jdff dff_B_iNMnHjWV0_2(.din(n1049),.dout(w_dff_B_iNMnHjWV0_2),.clk(gclk));
	jdff dff_B_5HjPxClh0_2(.din(w_dff_B_iNMnHjWV0_2),.dout(w_dff_B_5HjPxClh0_2),.clk(gclk));
	jdff dff_B_OMV4n6lG3_2(.din(w_dff_B_5HjPxClh0_2),.dout(w_dff_B_OMV4n6lG3_2),.clk(gclk));
	jdff dff_B_hXRvGQNO1_2(.din(w_dff_B_OMV4n6lG3_2),.dout(w_dff_B_hXRvGQNO1_2),.clk(gclk));
	jdff dff_B_0kH68DPw6_2(.din(w_dff_B_hXRvGQNO1_2),.dout(w_dff_B_0kH68DPw6_2),.clk(gclk));
	jdff dff_B_15w2wBG63_2(.din(w_dff_B_0kH68DPw6_2),.dout(w_dff_B_15w2wBG63_2),.clk(gclk));
	jdff dff_B_scZFHE220_2(.din(w_dff_B_15w2wBG63_2),.dout(w_dff_B_scZFHE220_2),.clk(gclk));
	jdff dff_B_bmzkcFqB3_2(.din(w_dff_B_scZFHE220_2),.dout(w_dff_B_bmzkcFqB3_2),.clk(gclk));
	jdff dff_B_FcHGVivP9_2(.din(w_dff_B_bmzkcFqB3_2),.dout(w_dff_B_FcHGVivP9_2),.clk(gclk));
	jdff dff_B_T5T2sVXp3_2(.din(w_dff_B_FcHGVivP9_2),.dout(w_dff_B_T5T2sVXp3_2),.clk(gclk));
	jdff dff_B_zuMkanZg0_2(.din(w_dff_B_T5T2sVXp3_2),.dout(w_dff_B_zuMkanZg0_2),.clk(gclk));
	jdff dff_B_waRBfHkp0_2(.din(w_dff_B_zuMkanZg0_2),.dout(w_dff_B_waRBfHkp0_2),.clk(gclk));
	jdff dff_B_O2HnyURc9_2(.din(w_dff_B_waRBfHkp0_2),.dout(w_dff_B_O2HnyURc9_2),.clk(gclk));
	jdff dff_B_r8YJhsfO0_2(.din(w_dff_B_O2HnyURc9_2),.dout(w_dff_B_r8YJhsfO0_2),.clk(gclk));
	jdff dff_B_0yELmqbw9_2(.din(w_dff_B_r8YJhsfO0_2),.dout(w_dff_B_0yELmqbw9_2),.clk(gclk));
	jdff dff_B_uq6Sipvg6_2(.din(w_dff_B_0yELmqbw9_2),.dout(w_dff_B_uq6Sipvg6_2),.clk(gclk));
	jdff dff_B_n2ALeWO01_2(.din(w_dff_B_uq6Sipvg6_2),.dout(w_dff_B_n2ALeWO01_2),.clk(gclk));
	jdff dff_B_LUnbG5p03_2(.din(w_dff_B_n2ALeWO01_2),.dout(w_dff_B_LUnbG5p03_2),.clk(gclk));
	jdff dff_B_W1xe0KwH4_2(.din(w_dff_B_LUnbG5p03_2),.dout(w_dff_B_W1xe0KwH4_2),.clk(gclk));
	jdff dff_B_6kZjZzGb6_2(.din(w_dff_B_W1xe0KwH4_2),.dout(w_dff_B_6kZjZzGb6_2),.clk(gclk));
	jdff dff_B_SNG295vV5_2(.din(w_dff_B_6kZjZzGb6_2),.dout(w_dff_B_SNG295vV5_2),.clk(gclk));
	jdff dff_B_gRNLXhAW7_2(.din(w_dff_B_SNG295vV5_2),.dout(w_dff_B_gRNLXhAW7_2),.clk(gclk));
	jdff dff_B_Rsmzu8z67_2(.din(w_dff_B_gRNLXhAW7_2),.dout(w_dff_B_Rsmzu8z67_2),.clk(gclk));
	jdff dff_B_wHxO7Paz8_2(.din(w_dff_B_Rsmzu8z67_2),.dout(w_dff_B_wHxO7Paz8_2),.clk(gclk));
	jdff dff_B_gRYISlmU2_2(.din(w_dff_B_wHxO7Paz8_2),.dout(w_dff_B_gRYISlmU2_2),.clk(gclk));
	jdff dff_B_lLJ5ZAtj5_2(.din(w_dff_B_gRYISlmU2_2),.dout(w_dff_B_lLJ5ZAtj5_2),.clk(gclk));
	jdff dff_B_3JQvdVkT6_2(.din(w_dff_B_lLJ5ZAtj5_2),.dout(w_dff_B_3JQvdVkT6_2),.clk(gclk));
	jdff dff_B_uWdZWg122_2(.din(w_dff_B_3JQvdVkT6_2),.dout(w_dff_B_uWdZWg122_2),.clk(gclk));
	jdff dff_B_6wqui3nG3_2(.din(w_dff_B_uWdZWg122_2),.dout(w_dff_B_6wqui3nG3_2),.clk(gclk));
	jdff dff_B_FmUM072u5_2(.din(w_dff_B_6wqui3nG3_2),.dout(w_dff_B_FmUM072u5_2),.clk(gclk));
	jdff dff_B_WbZHUZFl1_2(.din(w_dff_B_FmUM072u5_2),.dout(w_dff_B_WbZHUZFl1_2),.clk(gclk));
	jdff dff_B_Yf8cyQ189_2(.din(w_dff_B_WbZHUZFl1_2),.dout(w_dff_B_Yf8cyQ189_2),.clk(gclk));
	jdff dff_B_vJf8brBr6_2(.din(w_dff_B_Yf8cyQ189_2),.dout(w_dff_B_vJf8brBr6_2),.clk(gclk));
	jdff dff_B_3xVWWNr32_2(.din(w_dff_B_vJf8brBr6_2),.dout(w_dff_B_3xVWWNr32_2),.clk(gclk));
	jdff dff_B_HXsqowzj6_2(.din(w_dff_B_3xVWWNr32_2),.dout(w_dff_B_HXsqowzj6_2),.clk(gclk));
	jdff dff_B_b2t2bj9c2_2(.din(w_dff_B_HXsqowzj6_2),.dout(w_dff_B_b2t2bj9c2_2),.clk(gclk));
	jdff dff_B_xkpS3onQ1_2(.din(w_dff_B_b2t2bj9c2_2),.dout(w_dff_B_xkpS3onQ1_2),.clk(gclk));
	jdff dff_B_8F4401XA9_2(.din(w_dff_B_xkpS3onQ1_2),.dout(w_dff_B_8F4401XA9_2),.clk(gclk));
	jdff dff_B_3ys7jXIa3_2(.din(w_dff_B_8F4401XA9_2),.dout(w_dff_B_3ys7jXIa3_2),.clk(gclk));
	jdff dff_B_1D5F9tCx2_2(.din(w_dff_B_3ys7jXIa3_2),.dout(w_dff_B_1D5F9tCx2_2),.clk(gclk));
	jdff dff_B_1ePHcbk11_2(.din(w_dff_B_1D5F9tCx2_2),.dout(w_dff_B_1ePHcbk11_2),.clk(gclk));
	jdff dff_B_AbRIsUjF5_2(.din(w_dff_B_1ePHcbk11_2),.dout(w_dff_B_AbRIsUjF5_2),.clk(gclk));
	jdff dff_B_rdvUAVGU5_2(.din(n1135),.dout(w_dff_B_rdvUAVGU5_2),.clk(gclk));
	jdff dff_B_meIcJku66_1(.din(n1050),.dout(w_dff_B_meIcJku66_1),.clk(gclk));
	jdff dff_B_eqQbwuD19_2(.din(n951),.dout(w_dff_B_eqQbwuD19_2),.clk(gclk));
	jdff dff_B_7ZEhjk2q5_2(.din(w_dff_B_eqQbwuD19_2),.dout(w_dff_B_7ZEhjk2q5_2),.clk(gclk));
	jdff dff_B_Mhh4rQ9h0_2(.din(w_dff_B_7ZEhjk2q5_2),.dout(w_dff_B_Mhh4rQ9h0_2),.clk(gclk));
	jdff dff_B_Ky6pV3WL6_2(.din(w_dff_B_Mhh4rQ9h0_2),.dout(w_dff_B_Ky6pV3WL6_2),.clk(gclk));
	jdff dff_B_T0ZUg2d78_2(.din(w_dff_B_Ky6pV3WL6_2),.dout(w_dff_B_T0ZUg2d78_2),.clk(gclk));
	jdff dff_B_DZX70JOu0_2(.din(w_dff_B_T0ZUg2d78_2),.dout(w_dff_B_DZX70JOu0_2),.clk(gclk));
	jdff dff_B_iRPohZZU0_2(.din(w_dff_B_DZX70JOu0_2),.dout(w_dff_B_iRPohZZU0_2),.clk(gclk));
	jdff dff_B_k8TgaVrf1_2(.din(w_dff_B_iRPohZZU0_2),.dout(w_dff_B_k8TgaVrf1_2),.clk(gclk));
	jdff dff_B_TRonZ1RH1_2(.din(w_dff_B_k8TgaVrf1_2),.dout(w_dff_B_TRonZ1RH1_2),.clk(gclk));
	jdff dff_B_nmb0H0LR2_2(.din(w_dff_B_TRonZ1RH1_2),.dout(w_dff_B_nmb0H0LR2_2),.clk(gclk));
	jdff dff_B_6PKRvAUd2_2(.din(w_dff_B_nmb0H0LR2_2),.dout(w_dff_B_6PKRvAUd2_2),.clk(gclk));
	jdff dff_B_NkxEajnw3_2(.din(w_dff_B_6PKRvAUd2_2),.dout(w_dff_B_NkxEajnw3_2),.clk(gclk));
	jdff dff_B_02xyN4cw8_2(.din(w_dff_B_NkxEajnw3_2),.dout(w_dff_B_02xyN4cw8_2),.clk(gclk));
	jdff dff_B_ViQZTLPK3_2(.din(w_dff_B_02xyN4cw8_2),.dout(w_dff_B_ViQZTLPK3_2),.clk(gclk));
	jdff dff_B_SUAiV7wt4_2(.din(w_dff_B_ViQZTLPK3_2),.dout(w_dff_B_SUAiV7wt4_2),.clk(gclk));
	jdff dff_B_QvBLEJa96_2(.din(w_dff_B_SUAiV7wt4_2),.dout(w_dff_B_QvBLEJa96_2),.clk(gclk));
	jdff dff_B_sOd6C8IF1_2(.din(w_dff_B_QvBLEJa96_2),.dout(w_dff_B_sOd6C8IF1_2),.clk(gclk));
	jdff dff_B_HmjaLFUn7_2(.din(w_dff_B_sOd6C8IF1_2),.dout(w_dff_B_HmjaLFUn7_2),.clk(gclk));
	jdff dff_B_9iBz9BZr0_2(.din(w_dff_B_HmjaLFUn7_2),.dout(w_dff_B_9iBz9BZr0_2),.clk(gclk));
	jdff dff_B_Br0IU2by3_2(.din(w_dff_B_9iBz9BZr0_2),.dout(w_dff_B_Br0IU2by3_2),.clk(gclk));
	jdff dff_B_SLRbH0SZ3_2(.din(w_dff_B_Br0IU2by3_2),.dout(w_dff_B_SLRbH0SZ3_2),.clk(gclk));
	jdff dff_B_akP5Pr0z6_2(.din(w_dff_B_SLRbH0SZ3_2),.dout(w_dff_B_akP5Pr0z6_2),.clk(gclk));
	jdff dff_B_i98bKQRl3_2(.din(w_dff_B_akP5Pr0z6_2),.dout(w_dff_B_i98bKQRl3_2),.clk(gclk));
	jdff dff_B_sLw84q5N1_2(.din(w_dff_B_i98bKQRl3_2),.dout(w_dff_B_sLw84q5N1_2),.clk(gclk));
	jdff dff_B_oGgnWCGX6_2(.din(w_dff_B_sLw84q5N1_2),.dout(w_dff_B_oGgnWCGX6_2),.clk(gclk));
	jdff dff_B_2hc1pEix2_2(.din(w_dff_B_oGgnWCGX6_2),.dout(w_dff_B_2hc1pEix2_2),.clk(gclk));
	jdff dff_B_RizyaOpd5_2(.din(w_dff_B_2hc1pEix2_2),.dout(w_dff_B_RizyaOpd5_2),.clk(gclk));
	jdff dff_B_UmSXSHi78_2(.din(w_dff_B_RizyaOpd5_2),.dout(w_dff_B_UmSXSHi78_2),.clk(gclk));
	jdff dff_B_oSXyEGlP8_2(.din(w_dff_B_UmSXSHi78_2),.dout(w_dff_B_oSXyEGlP8_2),.clk(gclk));
	jdff dff_B_PiAyqK7i8_2(.din(w_dff_B_oSXyEGlP8_2),.dout(w_dff_B_PiAyqK7i8_2),.clk(gclk));
	jdff dff_B_FGcdhoVp0_2(.din(w_dff_B_PiAyqK7i8_2),.dout(w_dff_B_FGcdhoVp0_2),.clk(gclk));
	jdff dff_B_QrRRimLK3_2(.din(w_dff_B_FGcdhoVp0_2),.dout(w_dff_B_QrRRimLK3_2),.clk(gclk));
	jdff dff_B_o7DzriGY2_2(.din(w_dff_B_QrRRimLK3_2),.dout(w_dff_B_o7DzriGY2_2),.clk(gclk));
	jdff dff_B_pcx0bA3k5_2(.din(w_dff_B_o7DzriGY2_2),.dout(w_dff_B_pcx0bA3k5_2),.clk(gclk));
	jdff dff_B_CmIl0sOT2_2(.din(w_dff_B_pcx0bA3k5_2),.dout(w_dff_B_CmIl0sOT2_2),.clk(gclk));
	jdff dff_B_D6a944kG4_2(.din(w_dff_B_CmIl0sOT2_2),.dout(w_dff_B_D6a944kG4_2),.clk(gclk));
	jdff dff_B_AHIF6KrI3_2(.din(w_dff_B_D6a944kG4_2),.dout(w_dff_B_AHIF6KrI3_2),.clk(gclk));
	jdff dff_B_m3dEVGtb0_2(.din(n1030),.dout(w_dff_B_m3dEVGtb0_2),.clk(gclk));
	jdff dff_B_mILTqqt04_1(.din(n952),.dout(w_dff_B_mILTqqt04_1),.clk(gclk));
	jdff dff_B_stFAc2Bj6_2(.din(n846),.dout(w_dff_B_stFAc2Bj6_2),.clk(gclk));
	jdff dff_B_AJ5NI2ek9_2(.din(w_dff_B_stFAc2Bj6_2),.dout(w_dff_B_AJ5NI2ek9_2),.clk(gclk));
	jdff dff_B_zgHu8R7O3_2(.din(w_dff_B_AJ5NI2ek9_2),.dout(w_dff_B_zgHu8R7O3_2),.clk(gclk));
	jdff dff_B_V5qaQwey2_2(.din(w_dff_B_zgHu8R7O3_2),.dout(w_dff_B_V5qaQwey2_2),.clk(gclk));
	jdff dff_B_ab4FaQyv0_2(.din(w_dff_B_V5qaQwey2_2),.dout(w_dff_B_ab4FaQyv0_2),.clk(gclk));
	jdff dff_B_uJUWv9AP1_2(.din(w_dff_B_ab4FaQyv0_2),.dout(w_dff_B_uJUWv9AP1_2),.clk(gclk));
	jdff dff_B_bWnqCw5C6_2(.din(w_dff_B_uJUWv9AP1_2),.dout(w_dff_B_bWnqCw5C6_2),.clk(gclk));
	jdff dff_B_PaWFGgsD9_2(.din(w_dff_B_bWnqCw5C6_2),.dout(w_dff_B_PaWFGgsD9_2),.clk(gclk));
	jdff dff_B_8Rvi8o8v8_2(.din(w_dff_B_PaWFGgsD9_2),.dout(w_dff_B_8Rvi8o8v8_2),.clk(gclk));
	jdff dff_B_8xmQrgpQ3_2(.din(w_dff_B_8Rvi8o8v8_2),.dout(w_dff_B_8xmQrgpQ3_2),.clk(gclk));
	jdff dff_B_NjSlqKvw5_2(.din(w_dff_B_8xmQrgpQ3_2),.dout(w_dff_B_NjSlqKvw5_2),.clk(gclk));
	jdff dff_B_zKfxGX9u6_2(.din(w_dff_B_NjSlqKvw5_2),.dout(w_dff_B_zKfxGX9u6_2),.clk(gclk));
	jdff dff_B_uyj7bbH26_2(.din(w_dff_B_zKfxGX9u6_2),.dout(w_dff_B_uyj7bbH26_2),.clk(gclk));
	jdff dff_B_Ix0kHojs9_2(.din(w_dff_B_uyj7bbH26_2),.dout(w_dff_B_Ix0kHojs9_2),.clk(gclk));
	jdff dff_B_HiZ5F0NJ0_2(.din(w_dff_B_Ix0kHojs9_2),.dout(w_dff_B_HiZ5F0NJ0_2),.clk(gclk));
	jdff dff_B_qQjwxNPs8_2(.din(w_dff_B_HiZ5F0NJ0_2),.dout(w_dff_B_qQjwxNPs8_2),.clk(gclk));
	jdff dff_B_9mPjWmwy7_2(.din(w_dff_B_qQjwxNPs8_2),.dout(w_dff_B_9mPjWmwy7_2),.clk(gclk));
	jdff dff_B_PzFpS3aL9_2(.din(w_dff_B_9mPjWmwy7_2),.dout(w_dff_B_PzFpS3aL9_2),.clk(gclk));
	jdff dff_B_IW8xLLZV9_2(.din(w_dff_B_PzFpS3aL9_2),.dout(w_dff_B_IW8xLLZV9_2),.clk(gclk));
	jdff dff_B_tWWScgaR0_2(.din(w_dff_B_IW8xLLZV9_2),.dout(w_dff_B_tWWScgaR0_2),.clk(gclk));
	jdff dff_B_QjwAqWEO9_2(.din(w_dff_B_tWWScgaR0_2),.dout(w_dff_B_QjwAqWEO9_2),.clk(gclk));
	jdff dff_B_lztXbDZL0_2(.din(w_dff_B_QjwAqWEO9_2),.dout(w_dff_B_lztXbDZL0_2),.clk(gclk));
	jdff dff_B_lO9uSmIZ2_2(.din(w_dff_B_lztXbDZL0_2),.dout(w_dff_B_lO9uSmIZ2_2),.clk(gclk));
	jdff dff_B_gM7O6HhC5_2(.din(w_dff_B_lO9uSmIZ2_2),.dout(w_dff_B_gM7O6HhC5_2),.clk(gclk));
	jdff dff_B_YeQYBF960_2(.din(w_dff_B_gM7O6HhC5_2),.dout(w_dff_B_YeQYBF960_2),.clk(gclk));
	jdff dff_B_A404kjfF5_2(.din(w_dff_B_YeQYBF960_2),.dout(w_dff_B_A404kjfF5_2),.clk(gclk));
	jdff dff_B_WgbQywpY3_2(.din(w_dff_B_A404kjfF5_2),.dout(w_dff_B_WgbQywpY3_2),.clk(gclk));
	jdff dff_B_SElweEU06_2(.din(w_dff_B_WgbQywpY3_2),.dout(w_dff_B_SElweEU06_2),.clk(gclk));
	jdff dff_B_6DmLUu9r0_2(.din(w_dff_B_SElweEU06_2),.dout(w_dff_B_6DmLUu9r0_2),.clk(gclk));
	jdff dff_B_hEL1jvx86_2(.din(w_dff_B_6DmLUu9r0_2),.dout(w_dff_B_hEL1jvx86_2),.clk(gclk));
	jdff dff_B_nn9nDP6E8_2(.din(w_dff_B_hEL1jvx86_2),.dout(w_dff_B_nn9nDP6E8_2),.clk(gclk));
	jdff dff_B_FEd5SPu67_2(.din(w_dff_B_nn9nDP6E8_2),.dout(w_dff_B_FEd5SPu67_2),.clk(gclk));
	jdff dff_B_QULM0WWm1_2(.din(w_dff_B_FEd5SPu67_2),.dout(w_dff_B_QULM0WWm1_2),.clk(gclk));
	jdff dff_B_jU74dILT4_2(.din(w_dff_B_QULM0WWm1_2),.dout(w_dff_B_jU74dILT4_2),.clk(gclk));
	jdff dff_B_7XoFcijs1_2(.din(n925),.dout(w_dff_B_7XoFcijs1_2),.clk(gclk));
	jdff dff_B_zyKCsiWb0_1(.din(n847),.dout(w_dff_B_zyKCsiWb0_1),.clk(gclk));
	jdff dff_B_We9Z8XBh8_2(.din(n747),.dout(w_dff_B_We9Z8XBh8_2),.clk(gclk));
	jdff dff_B_mdNiJjxS3_2(.din(w_dff_B_We9Z8XBh8_2),.dout(w_dff_B_mdNiJjxS3_2),.clk(gclk));
	jdff dff_B_p9xagXVH9_2(.din(w_dff_B_mdNiJjxS3_2),.dout(w_dff_B_p9xagXVH9_2),.clk(gclk));
	jdff dff_B_9YjJxp4u5_2(.din(w_dff_B_p9xagXVH9_2),.dout(w_dff_B_9YjJxp4u5_2),.clk(gclk));
	jdff dff_B_KYKnToLb7_2(.din(w_dff_B_9YjJxp4u5_2),.dout(w_dff_B_KYKnToLb7_2),.clk(gclk));
	jdff dff_B_J254yehR8_2(.din(w_dff_B_KYKnToLb7_2),.dout(w_dff_B_J254yehR8_2),.clk(gclk));
	jdff dff_B_1XtR4fN54_2(.din(w_dff_B_J254yehR8_2),.dout(w_dff_B_1XtR4fN54_2),.clk(gclk));
	jdff dff_B_v1FinV3Y0_2(.din(w_dff_B_1XtR4fN54_2),.dout(w_dff_B_v1FinV3Y0_2),.clk(gclk));
	jdff dff_B_vOF6JRXL2_2(.din(w_dff_B_v1FinV3Y0_2),.dout(w_dff_B_vOF6JRXL2_2),.clk(gclk));
	jdff dff_B_LsNQSsFU8_2(.din(w_dff_B_vOF6JRXL2_2),.dout(w_dff_B_LsNQSsFU8_2),.clk(gclk));
	jdff dff_B_mky0OAFw7_2(.din(w_dff_B_LsNQSsFU8_2),.dout(w_dff_B_mky0OAFw7_2),.clk(gclk));
	jdff dff_B_qIioBpRo0_2(.din(w_dff_B_mky0OAFw7_2),.dout(w_dff_B_qIioBpRo0_2),.clk(gclk));
	jdff dff_B_1aYFacmk1_2(.din(w_dff_B_qIioBpRo0_2),.dout(w_dff_B_1aYFacmk1_2),.clk(gclk));
	jdff dff_B_JDyPD08J4_2(.din(w_dff_B_1aYFacmk1_2),.dout(w_dff_B_JDyPD08J4_2),.clk(gclk));
	jdff dff_B_RlB8V2kd5_2(.din(w_dff_B_JDyPD08J4_2),.dout(w_dff_B_RlB8V2kd5_2),.clk(gclk));
	jdff dff_B_aqMNWGO69_2(.din(w_dff_B_RlB8V2kd5_2),.dout(w_dff_B_aqMNWGO69_2),.clk(gclk));
	jdff dff_B_pUn6F2fF2_2(.din(w_dff_B_aqMNWGO69_2),.dout(w_dff_B_pUn6F2fF2_2),.clk(gclk));
	jdff dff_B_2WaI5Fi15_2(.din(w_dff_B_pUn6F2fF2_2),.dout(w_dff_B_2WaI5Fi15_2),.clk(gclk));
	jdff dff_B_kKOUUeLy4_2(.din(w_dff_B_2WaI5Fi15_2),.dout(w_dff_B_kKOUUeLy4_2),.clk(gclk));
	jdff dff_B_xUUM9IQG0_2(.din(w_dff_B_kKOUUeLy4_2),.dout(w_dff_B_xUUM9IQG0_2),.clk(gclk));
	jdff dff_B_l4cFAL2j9_2(.din(w_dff_B_xUUM9IQG0_2),.dout(w_dff_B_l4cFAL2j9_2),.clk(gclk));
	jdff dff_B_OBvKMMPj5_2(.din(w_dff_B_l4cFAL2j9_2),.dout(w_dff_B_OBvKMMPj5_2),.clk(gclk));
	jdff dff_B_aAv4rUYN1_2(.din(w_dff_B_OBvKMMPj5_2),.dout(w_dff_B_aAv4rUYN1_2),.clk(gclk));
	jdff dff_B_xDnmvA5n8_2(.din(w_dff_B_aAv4rUYN1_2),.dout(w_dff_B_xDnmvA5n8_2),.clk(gclk));
	jdff dff_B_P0N2xsry4_2(.din(w_dff_B_xDnmvA5n8_2),.dout(w_dff_B_P0N2xsry4_2),.clk(gclk));
	jdff dff_B_ejzxZOMW8_2(.din(w_dff_B_P0N2xsry4_2),.dout(w_dff_B_ejzxZOMW8_2),.clk(gclk));
	jdff dff_B_lJscurRa6_2(.din(w_dff_B_ejzxZOMW8_2),.dout(w_dff_B_lJscurRa6_2),.clk(gclk));
	jdff dff_B_kBwr3cgl3_2(.din(w_dff_B_lJscurRa6_2),.dout(w_dff_B_kBwr3cgl3_2),.clk(gclk));
	jdff dff_B_8ASJgFOC1_2(.din(w_dff_B_kBwr3cgl3_2),.dout(w_dff_B_8ASJgFOC1_2),.clk(gclk));
	jdff dff_B_keIzBWij9_2(.din(w_dff_B_8ASJgFOC1_2),.dout(w_dff_B_keIzBWij9_2),.clk(gclk));
	jdff dff_B_98cUKTy00_2(.din(w_dff_B_keIzBWij9_2),.dout(w_dff_B_98cUKTy00_2),.clk(gclk));
	jdff dff_B_WcmNniVo7_2(.din(n819),.dout(w_dff_B_WcmNniVo7_2),.clk(gclk));
	jdff dff_B_Jrwnh8Ov3_1(.din(n748),.dout(w_dff_B_Jrwnh8Ov3_1),.clk(gclk));
	jdff dff_B_f00ZAlqR5_2(.din(n654),.dout(w_dff_B_f00ZAlqR5_2),.clk(gclk));
	jdff dff_B_yqK1LtDd4_2(.din(w_dff_B_f00ZAlqR5_2),.dout(w_dff_B_yqK1LtDd4_2),.clk(gclk));
	jdff dff_B_nP5fgjlh6_2(.din(w_dff_B_yqK1LtDd4_2),.dout(w_dff_B_nP5fgjlh6_2),.clk(gclk));
	jdff dff_B_AX33OKgJ0_2(.din(w_dff_B_nP5fgjlh6_2),.dout(w_dff_B_AX33OKgJ0_2),.clk(gclk));
	jdff dff_B_oBrERymj0_2(.din(w_dff_B_AX33OKgJ0_2),.dout(w_dff_B_oBrERymj0_2),.clk(gclk));
	jdff dff_B_tp3C8vCo8_2(.din(w_dff_B_oBrERymj0_2),.dout(w_dff_B_tp3C8vCo8_2),.clk(gclk));
	jdff dff_B_XEShJlEV0_2(.din(w_dff_B_tp3C8vCo8_2),.dout(w_dff_B_XEShJlEV0_2),.clk(gclk));
	jdff dff_B_uDKTL3zM7_2(.din(w_dff_B_XEShJlEV0_2),.dout(w_dff_B_uDKTL3zM7_2),.clk(gclk));
	jdff dff_B_CGADboC25_2(.din(w_dff_B_uDKTL3zM7_2),.dout(w_dff_B_CGADboC25_2),.clk(gclk));
	jdff dff_B_ji3YnJRP1_2(.din(w_dff_B_CGADboC25_2),.dout(w_dff_B_ji3YnJRP1_2),.clk(gclk));
	jdff dff_B_Fk6tUKYK7_2(.din(w_dff_B_ji3YnJRP1_2),.dout(w_dff_B_Fk6tUKYK7_2),.clk(gclk));
	jdff dff_B_gzq3zFZ36_2(.din(w_dff_B_Fk6tUKYK7_2),.dout(w_dff_B_gzq3zFZ36_2),.clk(gclk));
	jdff dff_B_0pJMLwpF8_2(.din(w_dff_B_gzq3zFZ36_2),.dout(w_dff_B_0pJMLwpF8_2),.clk(gclk));
	jdff dff_B_1HH0YJwX0_2(.din(w_dff_B_0pJMLwpF8_2),.dout(w_dff_B_1HH0YJwX0_2),.clk(gclk));
	jdff dff_B_AdOsjWVc7_2(.din(w_dff_B_1HH0YJwX0_2),.dout(w_dff_B_AdOsjWVc7_2),.clk(gclk));
	jdff dff_B_n8hsLvsJ5_2(.din(w_dff_B_AdOsjWVc7_2),.dout(w_dff_B_n8hsLvsJ5_2),.clk(gclk));
	jdff dff_B_bw8R6iq72_2(.din(w_dff_B_n8hsLvsJ5_2),.dout(w_dff_B_bw8R6iq72_2),.clk(gclk));
	jdff dff_B_8rQg8CkI4_2(.din(w_dff_B_bw8R6iq72_2),.dout(w_dff_B_8rQg8CkI4_2),.clk(gclk));
	jdff dff_B_npgGVab36_2(.din(w_dff_B_8rQg8CkI4_2),.dout(w_dff_B_npgGVab36_2),.clk(gclk));
	jdff dff_B_DHoi7CfD6_2(.din(w_dff_B_npgGVab36_2),.dout(w_dff_B_DHoi7CfD6_2),.clk(gclk));
	jdff dff_B_Wlbn5PPV2_2(.din(w_dff_B_DHoi7CfD6_2),.dout(w_dff_B_Wlbn5PPV2_2),.clk(gclk));
	jdff dff_B_ZtaRnt5t4_2(.din(w_dff_B_Wlbn5PPV2_2),.dout(w_dff_B_ZtaRnt5t4_2),.clk(gclk));
	jdff dff_B_PVi658TA6_2(.din(w_dff_B_ZtaRnt5t4_2),.dout(w_dff_B_PVi658TA6_2),.clk(gclk));
	jdff dff_B_OX7rEuTv8_2(.din(w_dff_B_PVi658TA6_2),.dout(w_dff_B_OX7rEuTv8_2),.clk(gclk));
	jdff dff_B_wlGdNU8N8_2(.din(w_dff_B_OX7rEuTv8_2),.dout(w_dff_B_wlGdNU8N8_2),.clk(gclk));
	jdff dff_B_DwIRPnk66_2(.din(w_dff_B_wlGdNU8N8_2),.dout(w_dff_B_DwIRPnk66_2),.clk(gclk));
	jdff dff_B_gRlJwIzp3_2(.din(w_dff_B_DwIRPnk66_2),.dout(w_dff_B_gRlJwIzp3_2),.clk(gclk));
	jdff dff_B_YybAkBW14_2(.din(w_dff_B_gRlJwIzp3_2),.dout(w_dff_B_YybAkBW14_2),.clk(gclk));
	jdff dff_B_5HHz45KX0_2(.din(n719),.dout(w_dff_B_5HHz45KX0_2),.clk(gclk));
	jdff dff_B_k3h97Z802_1(.din(n655),.dout(w_dff_B_k3h97Z802_1),.clk(gclk));
	jdff dff_B_Zhfs6oPJ0_2(.din(n568),.dout(w_dff_B_Zhfs6oPJ0_2),.clk(gclk));
	jdff dff_B_r4oaUgYX9_2(.din(w_dff_B_Zhfs6oPJ0_2),.dout(w_dff_B_r4oaUgYX9_2),.clk(gclk));
	jdff dff_B_pPeQXJGT4_2(.din(w_dff_B_r4oaUgYX9_2),.dout(w_dff_B_pPeQXJGT4_2),.clk(gclk));
	jdff dff_B_QulQVZjg9_2(.din(w_dff_B_pPeQXJGT4_2),.dout(w_dff_B_QulQVZjg9_2),.clk(gclk));
	jdff dff_B_KOPuALy08_2(.din(w_dff_B_QulQVZjg9_2),.dout(w_dff_B_KOPuALy08_2),.clk(gclk));
	jdff dff_B_adQbcNVJ6_2(.din(w_dff_B_KOPuALy08_2),.dout(w_dff_B_adQbcNVJ6_2),.clk(gclk));
	jdff dff_B_X32gJhcy3_2(.din(w_dff_B_adQbcNVJ6_2),.dout(w_dff_B_X32gJhcy3_2),.clk(gclk));
	jdff dff_B_GiLNzKdD2_2(.din(w_dff_B_X32gJhcy3_2),.dout(w_dff_B_GiLNzKdD2_2),.clk(gclk));
	jdff dff_B_KADIC0AV0_2(.din(w_dff_B_GiLNzKdD2_2),.dout(w_dff_B_KADIC0AV0_2),.clk(gclk));
	jdff dff_B_VJ0LrDsJ5_2(.din(w_dff_B_KADIC0AV0_2),.dout(w_dff_B_VJ0LrDsJ5_2),.clk(gclk));
	jdff dff_B_pbBzgsqh9_2(.din(w_dff_B_VJ0LrDsJ5_2),.dout(w_dff_B_pbBzgsqh9_2),.clk(gclk));
	jdff dff_B_ilkwgL9p6_2(.din(w_dff_B_pbBzgsqh9_2),.dout(w_dff_B_ilkwgL9p6_2),.clk(gclk));
	jdff dff_B_zpPXU2Yq2_2(.din(w_dff_B_ilkwgL9p6_2),.dout(w_dff_B_zpPXU2Yq2_2),.clk(gclk));
	jdff dff_B_9Hw1d2E67_2(.din(w_dff_B_zpPXU2Yq2_2),.dout(w_dff_B_9Hw1d2E67_2),.clk(gclk));
	jdff dff_B_ci6Xkj838_2(.din(w_dff_B_9Hw1d2E67_2),.dout(w_dff_B_ci6Xkj838_2),.clk(gclk));
	jdff dff_B_T6ThZ1VN7_2(.din(w_dff_B_ci6Xkj838_2),.dout(w_dff_B_T6ThZ1VN7_2),.clk(gclk));
	jdff dff_B_efEoOrsF5_2(.din(w_dff_B_T6ThZ1VN7_2),.dout(w_dff_B_efEoOrsF5_2),.clk(gclk));
	jdff dff_B_1xQnkExC8_2(.din(w_dff_B_efEoOrsF5_2),.dout(w_dff_B_1xQnkExC8_2),.clk(gclk));
	jdff dff_B_4UzZik378_2(.din(w_dff_B_1xQnkExC8_2),.dout(w_dff_B_4UzZik378_2),.clk(gclk));
	jdff dff_B_LKVDHP0r2_2(.din(w_dff_B_4UzZik378_2),.dout(w_dff_B_LKVDHP0r2_2),.clk(gclk));
	jdff dff_B_VtqfVqPy5_2(.din(w_dff_B_LKVDHP0r2_2),.dout(w_dff_B_VtqfVqPy5_2),.clk(gclk));
	jdff dff_B_ytQFanFC4_2(.din(w_dff_B_VtqfVqPy5_2),.dout(w_dff_B_ytQFanFC4_2),.clk(gclk));
	jdff dff_B_oHZMPEqB3_2(.din(w_dff_B_ytQFanFC4_2),.dout(w_dff_B_oHZMPEqB3_2),.clk(gclk));
	jdff dff_B_xayU2yD50_2(.din(w_dff_B_oHZMPEqB3_2),.dout(w_dff_B_xayU2yD50_2),.clk(gclk));
	jdff dff_B_DAT7my1X3_2(.din(w_dff_B_xayU2yD50_2),.dout(w_dff_B_DAT7my1X3_2),.clk(gclk));
	jdff dff_B_YdHV0KgQ8_2(.din(n626),.dout(w_dff_B_YdHV0KgQ8_2),.clk(gclk));
	jdff dff_B_1RE9BRv90_1(.din(n569),.dout(w_dff_B_1RE9BRv90_1),.clk(gclk));
	jdff dff_B_1xrU55Ru8_2(.din(n489),.dout(w_dff_B_1xrU55Ru8_2),.clk(gclk));
	jdff dff_B_YaV28dQQ3_2(.din(w_dff_B_1xrU55Ru8_2),.dout(w_dff_B_YaV28dQQ3_2),.clk(gclk));
	jdff dff_B_Yjrc6gJ42_2(.din(w_dff_B_YaV28dQQ3_2),.dout(w_dff_B_Yjrc6gJ42_2),.clk(gclk));
	jdff dff_B_Ukr3cB5x0_2(.din(w_dff_B_Yjrc6gJ42_2),.dout(w_dff_B_Ukr3cB5x0_2),.clk(gclk));
	jdff dff_B_ERwYQfkc0_2(.din(w_dff_B_Ukr3cB5x0_2),.dout(w_dff_B_ERwYQfkc0_2),.clk(gclk));
	jdff dff_B_oQal8ZrF4_2(.din(w_dff_B_ERwYQfkc0_2),.dout(w_dff_B_oQal8ZrF4_2),.clk(gclk));
	jdff dff_B_usZwKi3J4_2(.din(w_dff_B_oQal8ZrF4_2),.dout(w_dff_B_usZwKi3J4_2),.clk(gclk));
	jdff dff_B_bCqitPJ50_2(.din(w_dff_B_usZwKi3J4_2),.dout(w_dff_B_bCqitPJ50_2),.clk(gclk));
	jdff dff_B_2ZyK4bWL7_2(.din(w_dff_B_bCqitPJ50_2),.dout(w_dff_B_2ZyK4bWL7_2),.clk(gclk));
	jdff dff_B_7gN6gaJ66_2(.din(w_dff_B_2ZyK4bWL7_2),.dout(w_dff_B_7gN6gaJ66_2),.clk(gclk));
	jdff dff_B_w8L7IhV79_2(.din(w_dff_B_7gN6gaJ66_2),.dout(w_dff_B_w8L7IhV79_2),.clk(gclk));
	jdff dff_B_7KutKp0b0_2(.din(w_dff_B_w8L7IhV79_2),.dout(w_dff_B_7KutKp0b0_2),.clk(gclk));
	jdff dff_B_yT8tjpoK7_2(.din(w_dff_B_7KutKp0b0_2),.dout(w_dff_B_yT8tjpoK7_2),.clk(gclk));
	jdff dff_B_uMs7yRyT9_2(.din(w_dff_B_yT8tjpoK7_2),.dout(w_dff_B_uMs7yRyT9_2),.clk(gclk));
	jdff dff_B_i2f7Y6Yv4_2(.din(w_dff_B_uMs7yRyT9_2),.dout(w_dff_B_i2f7Y6Yv4_2),.clk(gclk));
	jdff dff_B_AZdkpHa16_2(.din(w_dff_B_i2f7Y6Yv4_2),.dout(w_dff_B_AZdkpHa16_2),.clk(gclk));
	jdff dff_B_QmRVezwg1_2(.din(w_dff_B_AZdkpHa16_2),.dout(w_dff_B_QmRVezwg1_2),.clk(gclk));
	jdff dff_B_kjwPxhGc7_2(.din(w_dff_B_QmRVezwg1_2),.dout(w_dff_B_kjwPxhGc7_2),.clk(gclk));
	jdff dff_B_m4TgB3lK0_2(.din(w_dff_B_kjwPxhGc7_2),.dout(w_dff_B_m4TgB3lK0_2),.clk(gclk));
	jdff dff_B_gYPxl9zq4_2(.din(w_dff_B_m4TgB3lK0_2),.dout(w_dff_B_gYPxl9zq4_2),.clk(gclk));
	jdff dff_B_VWWjJVTc9_2(.din(w_dff_B_gYPxl9zq4_2),.dout(w_dff_B_VWWjJVTc9_2),.clk(gclk));
	jdff dff_B_vtYozoDN3_2(.din(w_dff_B_VWWjJVTc9_2),.dout(w_dff_B_vtYozoDN3_2),.clk(gclk));
	jdff dff_B_Jjsyq7Hc5_2(.din(n540),.dout(w_dff_B_Jjsyq7Hc5_2),.clk(gclk));
	jdff dff_B_nNxqHRh25_1(.din(n490),.dout(w_dff_B_nNxqHRh25_1),.clk(gclk));
	jdff dff_B_6FVp7wfK9_2(.din(n417),.dout(w_dff_B_6FVp7wfK9_2),.clk(gclk));
	jdff dff_B_uSVM9zp24_2(.din(w_dff_B_6FVp7wfK9_2),.dout(w_dff_B_uSVM9zp24_2),.clk(gclk));
	jdff dff_B_ZbwXR7sd0_2(.din(w_dff_B_uSVM9zp24_2),.dout(w_dff_B_ZbwXR7sd0_2),.clk(gclk));
	jdff dff_B_GR5cHUbp3_2(.din(w_dff_B_ZbwXR7sd0_2),.dout(w_dff_B_GR5cHUbp3_2),.clk(gclk));
	jdff dff_B_xBPaiVfs0_2(.din(w_dff_B_GR5cHUbp3_2),.dout(w_dff_B_xBPaiVfs0_2),.clk(gclk));
	jdff dff_B_wf3B6y9T1_2(.din(w_dff_B_xBPaiVfs0_2),.dout(w_dff_B_wf3B6y9T1_2),.clk(gclk));
	jdff dff_B_7yUhBR1v1_2(.din(w_dff_B_wf3B6y9T1_2),.dout(w_dff_B_7yUhBR1v1_2),.clk(gclk));
	jdff dff_B_u7qckrIH4_2(.din(w_dff_B_7yUhBR1v1_2),.dout(w_dff_B_u7qckrIH4_2),.clk(gclk));
	jdff dff_B_GZEZDqxD6_2(.din(w_dff_B_u7qckrIH4_2),.dout(w_dff_B_GZEZDqxD6_2),.clk(gclk));
	jdff dff_B_uTWclKZB0_2(.din(w_dff_B_GZEZDqxD6_2),.dout(w_dff_B_uTWclKZB0_2),.clk(gclk));
	jdff dff_B_kuWK8RGY5_2(.din(w_dff_B_uTWclKZB0_2),.dout(w_dff_B_kuWK8RGY5_2),.clk(gclk));
	jdff dff_B_y3VFfP5Q0_2(.din(w_dff_B_kuWK8RGY5_2),.dout(w_dff_B_y3VFfP5Q0_2),.clk(gclk));
	jdff dff_B_gqIGHKLq7_2(.din(w_dff_B_y3VFfP5Q0_2),.dout(w_dff_B_gqIGHKLq7_2),.clk(gclk));
	jdff dff_B_BJbuCKz14_2(.din(w_dff_B_gqIGHKLq7_2),.dout(w_dff_B_BJbuCKz14_2),.clk(gclk));
	jdff dff_B_hEekkcA76_2(.din(w_dff_B_BJbuCKz14_2),.dout(w_dff_B_hEekkcA76_2),.clk(gclk));
	jdff dff_B_3Yq3fpC63_2(.din(w_dff_B_hEekkcA76_2),.dout(w_dff_B_3Yq3fpC63_2),.clk(gclk));
	jdff dff_B_EQFCMH9U8_2(.din(w_dff_B_3Yq3fpC63_2),.dout(w_dff_B_EQFCMH9U8_2),.clk(gclk));
	jdff dff_B_Bpc4qT336_2(.din(w_dff_B_EQFCMH9U8_2),.dout(w_dff_B_Bpc4qT336_2),.clk(gclk));
	jdff dff_B_YprPyH070_2(.din(w_dff_B_Bpc4qT336_2),.dout(w_dff_B_YprPyH070_2),.clk(gclk));
	jdff dff_B_g1o7SUW86_2(.din(n461),.dout(w_dff_B_g1o7SUW86_2),.clk(gclk));
	jdff dff_B_Wnsct9yN9_1(.din(n418),.dout(w_dff_B_Wnsct9yN9_1),.clk(gclk));
	jdff dff_B_WLEthIES4_2(.din(n353),.dout(w_dff_B_WLEthIES4_2),.clk(gclk));
	jdff dff_B_JPVB1Lln7_2(.din(w_dff_B_WLEthIES4_2),.dout(w_dff_B_JPVB1Lln7_2),.clk(gclk));
	jdff dff_B_zoNuClxX2_2(.din(w_dff_B_JPVB1Lln7_2),.dout(w_dff_B_zoNuClxX2_2),.clk(gclk));
	jdff dff_B_MCAlPrUI6_2(.din(w_dff_B_zoNuClxX2_2),.dout(w_dff_B_MCAlPrUI6_2),.clk(gclk));
	jdff dff_B_MveQxUIh7_2(.din(w_dff_B_MCAlPrUI6_2),.dout(w_dff_B_MveQxUIh7_2),.clk(gclk));
	jdff dff_B_0yqxMRmq8_2(.din(w_dff_B_MveQxUIh7_2),.dout(w_dff_B_0yqxMRmq8_2),.clk(gclk));
	jdff dff_B_1uR6By4x2_2(.din(w_dff_B_0yqxMRmq8_2),.dout(w_dff_B_1uR6By4x2_2),.clk(gclk));
	jdff dff_B_G9FjQpuX6_2(.din(w_dff_B_1uR6By4x2_2),.dout(w_dff_B_G9FjQpuX6_2),.clk(gclk));
	jdff dff_B_pTXcbLj86_2(.din(w_dff_B_G9FjQpuX6_2),.dout(w_dff_B_pTXcbLj86_2),.clk(gclk));
	jdff dff_B_13aWHWaf9_2(.din(w_dff_B_pTXcbLj86_2),.dout(w_dff_B_13aWHWaf9_2),.clk(gclk));
	jdff dff_B_5omikSVf3_2(.din(w_dff_B_13aWHWaf9_2),.dout(w_dff_B_5omikSVf3_2),.clk(gclk));
	jdff dff_B_4TOZWLV17_2(.din(w_dff_B_5omikSVf3_2),.dout(w_dff_B_4TOZWLV17_2),.clk(gclk));
	jdff dff_B_nZPCvxHK3_2(.din(w_dff_B_4TOZWLV17_2),.dout(w_dff_B_nZPCvxHK3_2),.clk(gclk));
	jdff dff_B_rMH96HVO0_2(.din(w_dff_B_nZPCvxHK3_2),.dout(w_dff_B_rMH96HVO0_2),.clk(gclk));
	jdff dff_B_Z3Zdxp6i2_2(.din(w_dff_B_rMH96HVO0_2),.dout(w_dff_B_Z3Zdxp6i2_2),.clk(gclk));
	jdff dff_B_N8WbGEM79_2(.din(w_dff_B_Z3Zdxp6i2_2),.dout(w_dff_B_N8WbGEM79_2),.clk(gclk));
	jdff dff_B_6D1veawk7_2(.din(n389),.dout(w_dff_B_6D1veawk7_2),.clk(gclk));
	jdff dff_B_ySOKwf7v3_1(.din(n354),.dout(w_dff_B_ySOKwf7v3_1),.clk(gclk));
	jdff dff_B_Bu5kDFb36_2(.din(n295),.dout(w_dff_B_Bu5kDFb36_2),.clk(gclk));
	jdff dff_B_1gvMluSc3_2(.din(w_dff_B_Bu5kDFb36_2),.dout(w_dff_B_1gvMluSc3_2),.clk(gclk));
	jdff dff_B_pBCjjGPm9_2(.din(w_dff_B_1gvMluSc3_2),.dout(w_dff_B_pBCjjGPm9_2),.clk(gclk));
	jdff dff_B_Dk3u8Pgi5_2(.din(w_dff_B_pBCjjGPm9_2),.dout(w_dff_B_Dk3u8Pgi5_2),.clk(gclk));
	jdff dff_B_IshrJwqg4_2(.din(w_dff_B_Dk3u8Pgi5_2),.dout(w_dff_B_IshrJwqg4_2),.clk(gclk));
	jdff dff_B_PMtM9BMi8_2(.din(w_dff_B_IshrJwqg4_2),.dout(w_dff_B_PMtM9BMi8_2),.clk(gclk));
	jdff dff_B_yRbYU5eQ1_2(.din(w_dff_B_PMtM9BMi8_2),.dout(w_dff_B_yRbYU5eQ1_2),.clk(gclk));
	jdff dff_B_kpwSXUlE6_2(.din(w_dff_B_yRbYU5eQ1_2),.dout(w_dff_B_kpwSXUlE6_2),.clk(gclk));
	jdff dff_B_O39suy319_2(.din(w_dff_B_kpwSXUlE6_2),.dout(w_dff_B_O39suy319_2),.clk(gclk));
	jdff dff_B_WArw8JPJ4_2(.din(w_dff_B_O39suy319_2),.dout(w_dff_B_WArw8JPJ4_2),.clk(gclk));
	jdff dff_B_uyBdwhtL5_2(.din(w_dff_B_WArw8JPJ4_2),.dout(w_dff_B_uyBdwhtL5_2),.clk(gclk));
	jdff dff_B_11zFcYfw0_2(.din(w_dff_B_uyBdwhtL5_2),.dout(w_dff_B_11zFcYfw0_2),.clk(gclk));
	jdff dff_B_OiP437gK3_2(.din(w_dff_B_11zFcYfw0_2),.dout(w_dff_B_OiP437gK3_2),.clk(gclk));
	jdff dff_B_XBXvx0H27_2(.din(n325),.dout(w_dff_B_XBXvx0H27_2),.clk(gclk));
	jdff dff_B_iRswQ0ey1_1(.din(n296),.dout(w_dff_B_iRswQ0ey1_1),.clk(gclk));
	jdff dff_B_jcTjOypa2_2(.din(n244),.dout(w_dff_B_jcTjOypa2_2),.clk(gclk));
	jdff dff_B_9JznZKBa8_2(.din(w_dff_B_jcTjOypa2_2),.dout(w_dff_B_9JznZKBa8_2),.clk(gclk));
	jdff dff_B_6dmY5Vls7_2(.din(w_dff_B_9JznZKBa8_2),.dout(w_dff_B_6dmY5Vls7_2),.clk(gclk));
	jdff dff_B_4tL5MAtu1_2(.din(w_dff_B_6dmY5Vls7_2),.dout(w_dff_B_4tL5MAtu1_2),.clk(gclk));
	jdff dff_B_BF3tYk9g0_2(.din(w_dff_B_4tL5MAtu1_2),.dout(w_dff_B_BF3tYk9g0_2),.clk(gclk));
	jdff dff_B_bZvf2xlb5_2(.din(w_dff_B_BF3tYk9g0_2),.dout(w_dff_B_bZvf2xlb5_2),.clk(gclk));
	jdff dff_B_pZgW24Ge1_2(.din(w_dff_B_bZvf2xlb5_2),.dout(w_dff_B_pZgW24Ge1_2),.clk(gclk));
	jdff dff_B_NG9iA7hD7_2(.din(w_dff_B_pZgW24Ge1_2),.dout(w_dff_B_NG9iA7hD7_2),.clk(gclk));
	jdff dff_B_GD7v6uAu6_2(.din(w_dff_B_NG9iA7hD7_2),.dout(w_dff_B_GD7v6uAu6_2),.clk(gclk));
	jdff dff_B_oKHH0kyI4_2(.din(w_dff_B_GD7v6uAu6_2),.dout(w_dff_B_oKHH0kyI4_2),.clk(gclk));
	jdff dff_B_1ynuhIjH3_2(.din(n267),.dout(w_dff_B_1ynuhIjH3_2),.clk(gclk));
	jdff dff_B_15bCaxtq3_1(.din(n245),.dout(w_dff_B_15bCaxtq3_1),.clk(gclk));
	jdff dff_B_PwWkD2i26_2(.din(n201),.dout(w_dff_B_PwWkD2i26_2),.clk(gclk));
	jdff dff_B_QuL2VtNh3_2(.din(w_dff_B_PwWkD2i26_2),.dout(w_dff_B_QuL2VtNh3_2),.clk(gclk));
	jdff dff_B_64nu832F7_2(.din(w_dff_B_QuL2VtNh3_2),.dout(w_dff_B_64nu832F7_2),.clk(gclk));
	jdff dff_B_JFjJ9UwW9_2(.din(w_dff_B_64nu832F7_2),.dout(w_dff_B_JFjJ9UwW9_2),.clk(gclk));
	jdff dff_B_cktnGQw64_2(.din(w_dff_B_JFjJ9UwW9_2),.dout(w_dff_B_cktnGQw64_2),.clk(gclk));
	jdff dff_B_3hfS6LpD7_2(.din(w_dff_B_cktnGQw64_2),.dout(w_dff_B_3hfS6LpD7_2),.clk(gclk));
	jdff dff_B_mfADympr8_2(.din(w_dff_B_3hfS6LpD7_2),.dout(w_dff_B_mfADympr8_2),.clk(gclk));
	jdff dff_B_my4An37E2_2(.din(n216),.dout(w_dff_B_my4An37E2_2),.clk(gclk));
	jdff dff_B_CnGC1LJ43_1(.din(n202),.dout(w_dff_B_CnGC1LJ43_1),.clk(gclk));
	jdff dff_B_WDlZjkOk6_0(.din(n173),.dout(w_dff_B_WDlZjkOk6_0),.clk(gclk));
	jdff dff_B_SzUfRClK4_2(.din(n165),.dout(w_dff_B_SzUfRClK4_2),.clk(gclk));
	jdff dff_B_OIrHpVDL6_2(.din(w_dff_B_SzUfRClK4_2),.dout(w_dff_B_OIrHpVDL6_2),.clk(gclk));
	jdff dff_B_BOnTrUgh6_2(.din(w_dff_B_OIrHpVDL6_2),.dout(w_dff_B_BOnTrUgh6_2),.clk(gclk));
	jdff dff_B_kzWq9imN9_2(.din(w_dff_B_BOnTrUgh6_2),.dout(w_dff_B_kzWq9imN9_2),.clk(gclk));
	jdff dff_B_pFdws3C57_1(.din(n167),.dout(w_dff_B_pFdws3C57_1),.clk(gclk));
	jdff dff_A_WuclRIoY1_0(.dout(w_n132_0[0]),.din(w_dff_A_WuclRIoY1_0),.clk(gclk));
	jdff dff_A_dBh5L1BT2_0(.dout(w_dff_A_WuclRIoY1_0),.din(w_dff_A_dBh5L1BT2_0),.clk(gclk));
	jdff dff_A_nybzF4DU4_1(.dout(w_n132_0[1]),.din(w_dff_A_nybzF4DU4_1),.clk(gclk));
	jdff dff_B_2M717mWW2_1(.din(n1335),.dout(w_dff_B_2M717mWW2_1),.clk(gclk));
	jdff dff_B_LSlQbbUc4_2(.din(n1248),.dout(w_dff_B_LSlQbbUc4_2),.clk(gclk));
	jdff dff_B_L7JheQjM9_2(.din(w_dff_B_LSlQbbUc4_2),.dout(w_dff_B_L7JheQjM9_2),.clk(gclk));
	jdff dff_B_OooR60JJ8_2(.din(w_dff_B_L7JheQjM9_2),.dout(w_dff_B_OooR60JJ8_2),.clk(gclk));
	jdff dff_B_eh7Up9Fu0_2(.din(w_dff_B_OooR60JJ8_2),.dout(w_dff_B_eh7Up9Fu0_2),.clk(gclk));
	jdff dff_B_NV1Z95S91_2(.din(w_dff_B_eh7Up9Fu0_2),.dout(w_dff_B_NV1Z95S91_2),.clk(gclk));
	jdff dff_B_CHB7EotM9_2(.din(w_dff_B_NV1Z95S91_2),.dout(w_dff_B_CHB7EotM9_2),.clk(gclk));
	jdff dff_B_IxPt0z7L4_2(.din(w_dff_B_CHB7EotM9_2),.dout(w_dff_B_IxPt0z7L4_2),.clk(gclk));
	jdff dff_B_knxtopdp1_2(.din(w_dff_B_IxPt0z7L4_2),.dout(w_dff_B_knxtopdp1_2),.clk(gclk));
	jdff dff_B_5hYVt8dC3_2(.din(w_dff_B_knxtopdp1_2),.dout(w_dff_B_5hYVt8dC3_2),.clk(gclk));
	jdff dff_B_CNUex1ct3_2(.din(w_dff_B_5hYVt8dC3_2),.dout(w_dff_B_CNUex1ct3_2),.clk(gclk));
	jdff dff_B_LCopGGo09_2(.din(w_dff_B_CNUex1ct3_2),.dout(w_dff_B_LCopGGo09_2),.clk(gclk));
	jdff dff_B_A6UB1nQT5_2(.din(w_dff_B_LCopGGo09_2),.dout(w_dff_B_A6UB1nQT5_2),.clk(gclk));
	jdff dff_B_7D7BeYab0_2(.din(w_dff_B_A6UB1nQT5_2),.dout(w_dff_B_7D7BeYab0_2),.clk(gclk));
	jdff dff_B_AmGCKWCi0_2(.din(w_dff_B_7D7BeYab0_2),.dout(w_dff_B_AmGCKWCi0_2),.clk(gclk));
	jdff dff_B_0w51Zm1m6_2(.din(w_dff_B_AmGCKWCi0_2),.dout(w_dff_B_0w51Zm1m6_2),.clk(gclk));
	jdff dff_B_U7wlVsm69_2(.din(w_dff_B_0w51Zm1m6_2),.dout(w_dff_B_U7wlVsm69_2),.clk(gclk));
	jdff dff_B_M7oa6wst3_2(.din(w_dff_B_U7wlVsm69_2),.dout(w_dff_B_M7oa6wst3_2),.clk(gclk));
	jdff dff_B_LtiZDGRA0_2(.din(w_dff_B_M7oa6wst3_2),.dout(w_dff_B_LtiZDGRA0_2),.clk(gclk));
	jdff dff_B_uMYL27yz2_2(.din(w_dff_B_LtiZDGRA0_2),.dout(w_dff_B_uMYL27yz2_2),.clk(gclk));
	jdff dff_B_Us7xfdiy0_2(.din(w_dff_B_uMYL27yz2_2),.dout(w_dff_B_Us7xfdiy0_2),.clk(gclk));
	jdff dff_B_CyVHJF063_2(.din(w_dff_B_Us7xfdiy0_2),.dout(w_dff_B_CyVHJF063_2),.clk(gclk));
	jdff dff_B_Prtpxoy29_2(.din(w_dff_B_CyVHJF063_2),.dout(w_dff_B_Prtpxoy29_2),.clk(gclk));
	jdff dff_B_hesYcBQ25_2(.din(w_dff_B_Prtpxoy29_2),.dout(w_dff_B_hesYcBQ25_2),.clk(gclk));
	jdff dff_B_MSFfHjxj9_2(.din(w_dff_B_hesYcBQ25_2),.dout(w_dff_B_MSFfHjxj9_2),.clk(gclk));
	jdff dff_B_ovwrTjgN8_2(.din(w_dff_B_MSFfHjxj9_2),.dout(w_dff_B_ovwrTjgN8_2),.clk(gclk));
	jdff dff_B_NIEcuV0g4_2(.din(w_dff_B_ovwrTjgN8_2),.dout(w_dff_B_NIEcuV0g4_2),.clk(gclk));
	jdff dff_B_6Q6vAWed1_2(.din(w_dff_B_NIEcuV0g4_2),.dout(w_dff_B_6Q6vAWed1_2),.clk(gclk));
	jdff dff_B_NVTlvgY32_2(.din(w_dff_B_6Q6vAWed1_2),.dout(w_dff_B_NVTlvgY32_2),.clk(gclk));
	jdff dff_B_KoJIRmpW9_2(.din(w_dff_B_NVTlvgY32_2),.dout(w_dff_B_KoJIRmpW9_2),.clk(gclk));
	jdff dff_B_Szg31fkN9_2(.din(w_dff_B_KoJIRmpW9_2),.dout(w_dff_B_Szg31fkN9_2),.clk(gclk));
	jdff dff_B_mioyXxj12_2(.din(w_dff_B_Szg31fkN9_2),.dout(w_dff_B_mioyXxj12_2),.clk(gclk));
	jdff dff_B_kf9bFCNS9_2(.din(w_dff_B_mioyXxj12_2),.dout(w_dff_B_kf9bFCNS9_2),.clk(gclk));
	jdff dff_B_eqosYD2w2_2(.din(w_dff_B_kf9bFCNS9_2),.dout(w_dff_B_eqosYD2w2_2),.clk(gclk));
	jdff dff_B_Dmf6m8BR0_2(.din(w_dff_B_eqosYD2w2_2),.dout(w_dff_B_Dmf6m8BR0_2),.clk(gclk));
	jdff dff_B_N9Qi9z0Q9_2(.din(w_dff_B_Dmf6m8BR0_2),.dout(w_dff_B_N9Qi9z0Q9_2),.clk(gclk));
	jdff dff_B_HpP7aRbU9_2(.din(w_dff_B_N9Qi9z0Q9_2),.dout(w_dff_B_HpP7aRbU9_2),.clk(gclk));
	jdff dff_B_b8e2FE217_2(.din(w_dff_B_HpP7aRbU9_2),.dout(w_dff_B_b8e2FE217_2),.clk(gclk));
	jdff dff_B_YexX2FXP8_2(.din(w_dff_B_b8e2FE217_2),.dout(w_dff_B_YexX2FXP8_2),.clk(gclk));
	jdff dff_B_v1u9n2wh9_2(.din(w_dff_B_YexX2FXP8_2),.dout(w_dff_B_v1u9n2wh9_2),.clk(gclk));
	jdff dff_B_IqiPKs9H6_2(.din(w_dff_B_v1u9n2wh9_2),.dout(w_dff_B_IqiPKs9H6_2),.clk(gclk));
	jdff dff_B_vkPk90SI4_2(.din(w_dff_B_IqiPKs9H6_2),.dout(w_dff_B_vkPk90SI4_2),.clk(gclk));
	jdff dff_B_dRHV32lw6_2(.din(w_dff_B_vkPk90SI4_2),.dout(w_dff_B_dRHV32lw6_2),.clk(gclk));
	jdff dff_B_w4YMeVRn7_2(.din(w_dff_B_dRHV32lw6_2),.dout(w_dff_B_w4YMeVRn7_2),.clk(gclk));
	jdff dff_B_gJ4jzwkt7_2(.din(w_dff_B_w4YMeVRn7_2),.dout(w_dff_B_gJ4jzwkt7_2),.clk(gclk));
	jdff dff_B_0xiW4LK49_2(.din(w_dff_B_gJ4jzwkt7_2),.dout(w_dff_B_0xiW4LK49_2),.clk(gclk));
	jdff dff_B_Ee5XMWLf9_0(.din(n1334),.dout(w_dff_B_Ee5XMWLf9_0),.clk(gclk));
	jdff dff_A_w51f6fKg9_1(.dout(w_n1322_0[1]),.din(w_dff_A_w51f6fKg9_1),.clk(gclk));
	jdff dff_B_xnCG75dL2_1(.din(n1249),.dout(w_dff_B_xnCG75dL2_1),.clk(gclk));
	jdff dff_B_53MaQN4X4_2(.din(n1158),.dout(w_dff_B_53MaQN4X4_2),.clk(gclk));
	jdff dff_B_KGanxDDu1_2(.din(w_dff_B_53MaQN4X4_2),.dout(w_dff_B_KGanxDDu1_2),.clk(gclk));
	jdff dff_B_Bs6gDwtV9_2(.din(w_dff_B_KGanxDDu1_2),.dout(w_dff_B_Bs6gDwtV9_2),.clk(gclk));
	jdff dff_B_ISeXTPpf9_2(.din(w_dff_B_Bs6gDwtV9_2),.dout(w_dff_B_ISeXTPpf9_2),.clk(gclk));
	jdff dff_B_lWNKAr9w4_2(.din(w_dff_B_ISeXTPpf9_2),.dout(w_dff_B_lWNKAr9w4_2),.clk(gclk));
	jdff dff_B_GmAjXuqL2_2(.din(w_dff_B_lWNKAr9w4_2),.dout(w_dff_B_GmAjXuqL2_2),.clk(gclk));
	jdff dff_B_Mnrrvqfb6_2(.din(w_dff_B_GmAjXuqL2_2),.dout(w_dff_B_Mnrrvqfb6_2),.clk(gclk));
	jdff dff_B_JUEOp0jP2_2(.din(w_dff_B_Mnrrvqfb6_2),.dout(w_dff_B_JUEOp0jP2_2),.clk(gclk));
	jdff dff_B_d1KfKdJO8_2(.din(w_dff_B_JUEOp0jP2_2),.dout(w_dff_B_d1KfKdJO8_2),.clk(gclk));
	jdff dff_B_43ejrfAY0_2(.din(w_dff_B_d1KfKdJO8_2),.dout(w_dff_B_43ejrfAY0_2),.clk(gclk));
	jdff dff_B_BjvUevhY5_2(.din(w_dff_B_43ejrfAY0_2),.dout(w_dff_B_BjvUevhY5_2),.clk(gclk));
	jdff dff_B_cnJSCd992_2(.din(w_dff_B_BjvUevhY5_2),.dout(w_dff_B_cnJSCd992_2),.clk(gclk));
	jdff dff_B_jUgNDZPm7_2(.din(w_dff_B_cnJSCd992_2),.dout(w_dff_B_jUgNDZPm7_2),.clk(gclk));
	jdff dff_B_xcCmmGRM3_2(.din(w_dff_B_jUgNDZPm7_2),.dout(w_dff_B_xcCmmGRM3_2),.clk(gclk));
	jdff dff_B_Hmhlsa1h3_2(.din(w_dff_B_xcCmmGRM3_2),.dout(w_dff_B_Hmhlsa1h3_2),.clk(gclk));
	jdff dff_B_QIkXkwcQ2_2(.din(w_dff_B_Hmhlsa1h3_2),.dout(w_dff_B_QIkXkwcQ2_2),.clk(gclk));
	jdff dff_B_jI0iw5Yv2_2(.din(w_dff_B_QIkXkwcQ2_2),.dout(w_dff_B_jI0iw5Yv2_2),.clk(gclk));
	jdff dff_B_93vMeepE7_2(.din(w_dff_B_jI0iw5Yv2_2),.dout(w_dff_B_93vMeepE7_2),.clk(gclk));
	jdff dff_B_NskGbCXo3_2(.din(w_dff_B_93vMeepE7_2),.dout(w_dff_B_NskGbCXo3_2),.clk(gclk));
	jdff dff_B_Q01G0jzX9_2(.din(w_dff_B_NskGbCXo3_2),.dout(w_dff_B_Q01G0jzX9_2),.clk(gclk));
	jdff dff_B_zHH4s5XG7_2(.din(w_dff_B_Q01G0jzX9_2),.dout(w_dff_B_zHH4s5XG7_2),.clk(gclk));
	jdff dff_B_qKiqwGLP5_2(.din(w_dff_B_zHH4s5XG7_2),.dout(w_dff_B_qKiqwGLP5_2),.clk(gclk));
	jdff dff_B_NfEjddmh5_2(.din(w_dff_B_qKiqwGLP5_2),.dout(w_dff_B_NfEjddmh5_2),.clk(gclk));
	jdff dff_B_9th4BbCO1_2(.din(w_dff_B_NfEjddmh5_2),.dout(w_dff_B_9th4BbCO1_2),.clk(gclk));
	jdff dff_B_DWX6gro16_2(.din(w_dff_B_9th4BbCO1_2),.dout(w_dff_B_DWX6gro16_2),.clk(gclk));
	jdff dff_B_jvwO0Dk37_2(.din(w_dff_B_DWX6gro16_2),.dout(w_dff_B_jvwO0Dk37_2),.clk(gclk));
	jdff dff_B_yyvrSAqx6_2(.din(w_dff_B_jvwO0Dk37_2),.dout(w_dff_B_yyvrSAqx6_2),.clk(gclk));
	jdff dff_B_kJII4sUl3_2(.din(w_dff_B_yyvrSAqx6_2),.dout(w_dff_B_kJII4sUl3_2),.clk(gclk));
	jdff dff_B_DCXxTNcP3_2(.din(w_dff_B_kJII4sUl3_2),.dout(w_dff_B_DCXxTNcP3_2),.clk(gclk));
	jdff dff_B_FhfigvyI6_2(.din(w_dff_B_DCXxTNcP3_2),.dout(w_dff_B_FhfigvyI6_2),.clk(gclk));
	jdff dff_B_gxHPoZ764_2(.din(w_dff_B_FhfigvyI6_2),.dout(w_dff_B_gxHPoZ764_2),.clk(gclk));
	jdff dff_B_uiGsonpX5_2(.din(w_dff_B_gxHPoZ764_2),.dout(w_dff_B_uiGsonpX5_2),.clk(gclk));
	jdff dff_B_jmigQF8R8_2(.din(w_dff_B_uiGsonpX5_2),.dout(w_dff_B_jmigQF8R8_2),.clk(gclk));
	jdff dff_B_1BkoRZqD4_2(.din(w_dff_B_jmigQF8R8_2),.dout(w_dff_B_1BkoRZqD4_2),.clk(gclk));
	jdff dff_B_xJJ4MQxu6_2(.din(w_dff_B_1BkoRZqD4_2),.dout(w_dff_B_xJJ4MQxu6_2),.clk(gclk));
	jdff dff_B_Af9XluMH3_2(.din(w_dff_B_xJJ4MQxu6_2),.dout(w_dff_B_Af9XluMH3_2),.clk(gclk));
	jdff dff_B_d0u4lOUS5_2(.din(w_dff_B_Af9XluMH3_2),.dout(w_dff_B_d0u4lOUS5_2),.clk(gclk));
	jdff dff_B_eSchcl8v1_2(.din(w_dff_B_d0u4lOUS5_2),.dout(w_dff_B_eSchcl8v1_2),.clk(gclk));
	jdff dff_B_Qs3PfOV91_2(.din(w_dff_B_eSchcl8v1_2),.dout(w_dff_B_Qs3PfOV91_2),.clk(gclk));
	jdff dff_B_2ErB38d85_2(.din(w_dff_B_Qs3PfOV91_2),.dout(w_dff_B_2ErB38d85_2),.clk(gclk));
	jdff dff_B_mr1nHZhz7_2(.din(n1231),.dout(w_dff_B_mr1nHZhz7_2),.clk(gclk));
	jdff dff_B_pNGp6yFR8_1(.din(n1159),.dout(w_dff_B_pNGp6yFR8_1),.clk(gclk));
	jdff dff_B_T1ijMHX20_2(.din(n1054),.dout(w_dff_B_T1ijMHX20_2),.clk(gclk));
	jdff dff_B_wFZKOjKB2_2(.din(w_dff_B_T1ijMHX20_2),.dout(w_dff_B_wFZKOjKB2_2),.clk(gclk));
	jdff dff_B_BbMdPf1Y1_2(.din(w_dff_B_wFZKOjKB2_2),.dout(w_dff_B_BbMdPf1Y1_2),.clk(gclk));
	jdff dff_B_FpTDjBFC9_2(.din(w_dff_B_BbMdPf1Y1_2),.dout(w_dff_B_FpTDjBFC9_2),.clk(gclk));
	jdff dff_B_BLBZhFu03_2(.din(w_dff_B_FpTDjBFC9_2),.dout(w_dff_B_BLBZhFu03_2),.clk(gclk));
	jdff dff_B_4gbJmk3O4_2(.din(w_dff_B_BLBZhFu03_2),.dout(w_dff_B_4gbJmk3O4_2),.clk(gclk));
	jdff dff_B_soxMN8Ja5_2(.din(w_dff_B_4gbJmk3O4_2),.dout(w_dff_B_soxMN8Ja5_2),.clk(gclk));
	jdff dff_B_oIvImuyX3_2(.din(w_dff_B_soxMN8Ja5_2),.dout(w_dff_B_oIvImuyX3_2),.clk(gclk));
	jdff dff_B_Shfkdzxj6_2(.din(w_dff_B_oIvImuyX3_2),.dout(w_dff_B_Shfkdzxj6_2),.clk(gclk));
	jdff dff_B_Fv119xlz5_2(.din(w_dff_B_Shfkdzxj6_2),.dout(w_dff_B_Fv119xlz5_2),.clk(gclk));
	jdff dff_B_LIRzKSoi3_2(.din(w_dff_B_Fv119xlz5_2),.dout(w_dff_B_LIRzKSoi3_2),.clk(gclk));
	jdff dff_B_ckSUSvKi3_2(.din(w_dff_B_LIRzKSoi3_2),.dout(w_dff_B_ckSUSvKi3_2),.clk(gclk));
	jdff dff_B_QX8ZCOEV9_2(.din(w_dff_B_ckSUSvKi3_2),.dout(w_dff_B_QX8ZCOEV9_2),.clk(gclk));
	jdff dff_B_biCmIdwW5_2(.din(w_dff_B_QX8ZCOEV9_2),.dout(w_dff_B_biCmIdwW5_2),.clk(gclk));
	jdff dff_B_In7ss3oz2_2(.din(w_dff_B_biCmIdwW5_2),.dout(w_dff_B_In7ss3oz2_2),.clk(gclk));
	jdff dff_B_m9R1ue6B1_2(.din(w_dff_B_In7ss3oz2_2),.dout(w_dff_B_m9R1ue6B1_2),.clk(gclk));
	jdff dff_B_jD5TeEdK8_2(.din(w_dff_B_m9R1ue6B1_2),.dout(w_dff_B_jD5TeEdK8_2),.clk(gclk));
	jdff dff_B_1tAT5HYP9_2(.din(w_dff_B_jD5TeEdK8_2),.dout(w_dff_B_1tAT5HYP9_2),.clk(gclk));
	jdff dff_B_w0lhWW4L0_2(.din(w_dff_B_1tAT5HYP9_2),.dout(w_dff_B_w0lhWW4L0_2),.clk(gclk));
	jdff dff_B_KaG9cDgs9_2(.din(w_dff_B_w0lhWW4L0_2),.dout(w_dff_B_KaG9cDgs9_2),.clk(gclk));
	jdff dff_B_t41gk4817_2(.din(w_dff_B_KaG9cDgs9_2),.dout(w_dff_B_t41gk4817_2),.clk(gclk));
	jdff dff_B_RRKOLcpu0_2(.din(w_dff_B_t41gk4817_2),.dout(w_dff_B_RRKOLcpu0_2),.clk(gclk));
	jdff dff_B_VPu0juO67_2(.din(w_dff_B_RRKOLcpu0_2),.dout(w_dff_B_VPu0juO67_2),.clk(gclk));
	jdff dff_B_sNgMEBVH1_2(.din(w_dff_B_VPu0juO67_2),.dout(w_dff_B_sNgMEBVH1_2),.clk(gclk));
	jdff dff_B_31fMGXW38_2(.din(w_dff_B_sNgMEBVH1_2),.dout(w_dff_B_31fMGXW38_2),.clk(gclk));
	jdff dff_B_ijDPh3q34_2(.din(w_dff_B_31fMGXW38_2),.dout(w_dff_B_ijDPh3q34_2),.clk(gclk));
	jdff dff_B_5BWcjAtN8_2(.din(w_dff_B_ijDPh3q34_2),.dout(w_dff_B_5BWcjAtN8_2),.clk(gclk));
	jdff dff_B_9gQurTIf8_2(.din(w_dff_B_5BWcjAtN8_2),.dout(w_dff_B_9gQurTIf8_2),.clk(gclk));
	jdff dff_B_vHMpXA5p1_2(.din(w_dff_B_9gQurTIf8_2),.dout(w_dff_B_vHMpXA5p1_2),.clk(gclk));
	jdff dff_B_C4hSN5h07_2(.din(w_dff_B_vHMpXA5p1_2),.dout(w_dff_B_C4hSN5h07_2),.clk(gclk));
	jdff dff_B_i6Kh2RHd0_2(.din(w_dff_B_C4hSN5h07_2),.dout(w_dff_B_i6Kh2RHd0_2),.clk(gclk));
	jdff dff_B_6ZXrghi65_2(.din(w_dff_B_i6Kh2RHd0_2),.dout(w_dff_B_6ZXrghi65_2),.clk(gclk));
	jdff dff_B_a94EnyxS3_2(.din(w_dff_B_6ZXrghi65_2),.dout(w_dff_B_a94EnyxS3_2),.clk(gclk));
	jdff dff_B_1sUde2R02_2(.din(w_dff_B_a94EnyxS3_2),.dout(w_dff_B_1sUde2R02_2),.clk(gclk));
	jdff dff_B_EMJpRulh7_2(.din(w_dff_B_1sUde2R02_2),.dout(w_dff_B_EMJpRulh7_2),.clk(gclk));
	jdff dff_B_UPNvuDtc2_2(.din(w_dff_B_EMJpRulh7_2),.dout(w_dff_B_UPNvuDtc2_2),.clk(gclk));
	jdff dff_B_e94QfI5g5_2(.din(w_dff_B_UPNvuDtc2_2),.dout(w_dff_B_e94QfI5g5_2),.clk(gclk));
	jdff dff_B_5LD0MFNh0_2(.din(n1133),.dout(w_dff_B_5LD0MFNh0_2),.clk(gclk));
	jdff dff_B_ECAasbK75_1(.din(n1055),.dout(w_dff_B_ECAasbK75_1),.clk(gclk));
	jdff dff_B_Ke20WAPe4_2(.din(n956),.dout(w_dff_B_Ke20WAPe4_2),.clk(gclk));
	jdff dff_B_1XjXP9l55_2(.din(w_dff_B_Ke20WAPe4_2),.dout(w_dff_B_1XjXP9l55_2),.clk(gclk));
	jdff dff_B_MMPIrmgd5_2(.din(w_dff_B_1XjXP9l55_2),.dout(w_dff_B_MMPIrmgd5_2),.clk(gclk));
	jdff dff_B_uAyCDodE7_2(.din(w_dff_B_MMPIrmgd5_2),.dout(w_dff_B_uAyCDodE7_2),.clk(gclk));
	jdff dff_B_c6lRLEDj9_2(.din(w_dff_B_uAyCDodE7_2),.dout(w_dff_B_c6lRLEDj9_2),.clk(gclk));
	jdff dff_B_o0bpbOf17_2(.din(w_dff_B_c6lRLEDj9_2),.dout(w_dff_B_o0bpbOf17_2),.clk(gclk));
	jdff dff_B_igfgnHTu4_2(.din(w_dff_B_o0bpbOf17_2),.dout(w_dff_B_igfgnHTu4_2),.clk(gclk));
	jdff dff_B_kNvsuaeZ6_2(.din(w_dff_B_igfgnHTu4_2),.dout(w_dff_B_kNvsuaeZ6_2),.clk(gclk));
	jdff dff_B_xy4bWwsH0_2(.din(w_dff_B_kNvsuaeZ6_2),.dout(w_dff_B_xy4bWwsH0_2),.clk(gclk));
	jdff dff_B_EbQJL6L00_2(.din(w_dff_B_xy4bWwsH0_2),.dout(w_dff_B_EbQJL6L00_2),.clk(gclk));
	jdff dff_B_cXD23sEV0_2(.din(w_dff_B_EbQJL6L00_2),.dout(w_dff_B_cXD23sEV0_2),.clk(gclk));
	jdff dff_B_lDxFzLCk0_2(.din(w_dff_B_cXD23sEV0_2),.dout(w_dff_B_lDxFzLCk0_2),.clk(gclk));
	jdff dff_B_whBou9vE4_2(.din(w_dff_B_lDxFzLCk0_2),.dout(w_dff_B_whBou9vE4_2),.clk(gclk));
	jdff dff_B_QksqPF8d0_2(.din(w_dff_B_whBou9vE4_2),.dout(w_dff_B_QksqPF8d0_2),.clk(gclk));
	jdff dff_B_u9vO1Nvb6_2(.din(w_dff_B_QksqPF8d0_2),.dout(w_dff_B_u9vO1Nvb6_2),.clk(gclk));
	jdff dff_B_J6XSEByu4_2(.din(w_dff_B_u9vO1Nvb6_2),.dout(w_dff_B_J6XSEByu4_2),.clk(gclk));
	jdff dff_B_oDqUxfck0_2(.din(w_dff_B_J6XSEByu4_2),.dout(w_dff_B_oDqUxfck0_2),.clk(gclk));
	jdff dff_B_tJIPaCUI7_2(.din(w_dff_B_oDqUxfck0_2),.dout(w_dff_B_tJIPaCUI7_2),.clk(gclk));
	jdff dff_B_j86xvJXf7_2(.din(w_dff_B_tJIPaCUI7_2),.dout(w_dff_B_j86xvJXf7_2),.clk(gclk));
	jdff dff_B_4N91gOOs5_2(.din(w_dff_B_j86xvJXf7_2),.dout(w_dff_B_4N91gOOs5_2),.clk(gclk));
	jdff dff_B_wVyFThKK2_2(.din(w_dff_B_4N91gOOs5_2),.dout(w_dff_B_wVyFThKK2_2),.clk(gclk));
	jdff dff_B_B1s2MeMh6_2(.din(w_dff_B_wVyFThKK2_2),.dout(w_dff_B_B1s2MeMh6_2),.clk(gclk));
	jdff dff_B_rb2LQZfP5_2(.din(w_dff_B_B1s2MeMh6_2),.dout(w_dff_B_rb2LQZfP5_2),.clk(gclk));
	jdff dff_B_RqShlrS31_2(.din(w_dff_B_rb2LQZfP5_2),.dout(w_dff_B_RqShlrS31_2),.clk(gclk));
	jdff dff_B_1GESWonR3_2(.din(w_dff_B_RqShlrS31_2),.dout(w_dff_B_1GESWonR3_2),.clk(gclk));
	jdff dff_B_2Ar4nirw1_2(.din(w_dff_B_1GESWonR3_2),.dout(w_dff_B_2Ar4nirw1_2),.clk(gclk));
	jdff dff_B_6yqp78Sn4_2(.din(w_dff_B_2Ar4nirw1_2),.dout(w_dff_B_6yqp78Sn4_2),.clk(gclk));
	jdff dff_B_q1ZkHdQL5_2(.din(w_dff_B_6yqp78Sn4_2),.dout(w_dff_B_q1ZkHdQL5_2),.clk(gclk));
	jdff dff_B_A9k3sJDT7_2(.din(w_dff_B_q1ZkHdQL5_2),.dout(w_dff_B_A9k3sJDT7_2),.clk(gclk));
	jdff dff_B_0fyOtX0z4_2(.din(w_dff_B_A9k3sJDT7_2),.dout(w_dff_B_0fyOtX0z4_2),.clk(gclk));
	jdff dff_B_EkfVU8YA2_2(.din(w_dff_B_0fyOtX0z4_2),.dout(w_dff_B_EkfVU8YA2_2),.clk(gclk));
	jdff dff_B_ropKusnn7_2(.din(w_dff_B_EkfVU8YA2_2),.dout(w_dff_B_ropKusnn7_2),.clk(gclk));
	jdff dff_B_nEgpEXPa6_2(.din(w_dff_B_ropKusnn7_2),.dout(w_dff_B_nEgpEXPa6_2),.clk(gclk));
	jdff dff_B_KSl44vcR5_2(.din(w_dff_B_nEgpEXPa6_2),.dout(w_dff_B_KSl44vcR5_2),.clk(gclk));
	jdff dff_B_n7NZzqfv9_2(.din(n1028),.dout(w_dff_B_n7NZzqfv9_2),.clk(gclk));
	jdff dff_B_uw7NCiMR7_1(.din(n957),.dout(w_dff_B_uw7NCiMR7_1),.clk(gclk));
	jdff dff_B_KvSqF5Xf6_2(.din(n851),.dout(w_dff_B_KvSqF5Xf6_2),.clk(gclk));
	jdff dff_B_zt9nszF87_2(.din(w_dff_B_KvSqF5Xf6_2),.dout(w_dff_B_zt9nszF87_2),.clk(gclk));
	jdff dff_B_vrcl4GP45_2(.din(w_dff_B_zt9nszF87_2),.dout(w_dff_B_vrcl4GP45_2),.clk(gclk));
	jdff dff_B_9IiAZcp32_2(.din(w_dff_B_vrcl4GP45_2),.dout(w_dff_B_9IiAZcp32_2),.clk(gclk));
	jdff dff_B_QYnN5lha2_2(.din(w_dff_B_9IiAZcp32_2),.dout(w_dff_B_QYnN5lha2_2),.clk(gclk));
	jdff dff_B_KrHSFf0N1_2(.din(w_dff_B_QYnN5lha2_2),.dout(w_dff_B_KrHSFf0N1_2),.clk(gclk));
	jdff dff_B_o4bt0WnC5_2(.din(w_dff_B_KrHSFf0N1_2),.dout(w_dff_B_o4bt0WnC5_2),.clk(gclk));
	jdff dff_B_nJnovh7Y1_2(.din(w_dff_B_o4bt0WnC5_2),.dout(w_dff_B_nJnovh7Y1_2),.clk(gclk));
	jdff dff_B_iFBffaZp4_2(.din(w_dff_B_nJnovh7Y1_2),.dout(w_dff_B_iFBffaZp4_2),.clk(gclk));
	jdff dff_B_FMGVtxxm0_2(.din(w_dff_B_iFBffaZp4_2),.dout(w_dff_B_FMGVtxxm0_2),.clk(gclk));
	jdff dff_B_ZDhITpnG4_2(.din(w_dff_B_FMGVtxxm0_2),.dout(w_dff_B_ZDhITpnG4_2),.clk(gclk));
	jdff dff_B_fG6TlCOR6_2(.din(w_dff_B_ZDhITpnG4_2),.dout(w_dff_B_fG6TlCOR6_2),.clk(gclk));
	jdff dff_B_1DB1riyM5_2(.din(w_dff_B_fG6TlCOR6_2),.dout(w_dff_B_1DB1riyM5_2),.clk(gclk));
	jdff dff_B_HBVtvih01_2(.din(w_dff_B_1DB1riyM5_2),.dout(w_dff_B_HBVtvih01_2),.clk(gclk));
	jdff dff_B_SBkTADVc5_2(.din(w_dff_B_HBVtvih01_2),.dout(w_dff_B_SBkTADVc5_2),.clk(gclk));
	jdff dff_B_gsO7nT6D4_2(.din(w_dff_B_SBkTADVc5_2),.dout(w_dff_B_gsO7nT6D4_2),.clk(gclk));
	jdff dff_B_AKbNUzs42_2(.din(w_dff_B_gsO7nT6D4_2),.dout(w_dff_B_AKbNUzs42_2),.clk(gclk));
	jdff dff_B_JPix2ID42_2(.din(w_dff_B_AKbNUzs42_2),.dout(w_dff_B_JPix2ID42_2),.clk(gclk));
	jdff dff_B_NF7cbl9P3_2(.din(w_dff_B_JPix2ID42_2),.dout(w_dff_B_NF7cbl9P3_2),.clk(gclk));
	jdff dff_B_tIBo4Md27_2(.din(w_dff_B_NF7cbl9P3_2),.dout(w_dff_B_tIBo4Md27_2),.clk(gclk));
	jdff dff_B_k7wjO0wN6_2(.din(w_dff_B_tIBo4Md27_2),.dout(w_dff_B_k7wjO0wN6_2),.clk(gclk));
	jdff dff_B_ovyvEWee1_2(.din(w_dff_B_k7wjO0wN6_2),.dout(w_dff_B_ovyvEWee1_2),.clk(gclk));
	jdff dff_B_X9jQoiQo6_2(.din(w_dff_B_ovyvEWee1_2),.dout(w_dff_B_X9jQoiQo6_2),.clk(gclk));
	jdff dff_B_7BOU26IH7_2(.din(w_dff_B_X9jQoiQo6_2),.dout(w_dff_B_7BOU26IH7_2),.clk(gclk));
	jdff dff_B_6yiJD5CE7_2(.din(w_dff_B_7BOU26IH7_2),.dout(w_dff_B_6yiJD5CE7_2),.clk(gclk));
	jdff dff_B_Dyf31tXD6_2(.din(w_dff_B_6yiJD5CE7_2),.dout(w_dff_B_Dyf31tXD6_2),.clk(gclk));
	jdff dff_B_cGnUEqZN1_2(.din(w_dff_B_Dyf31tXD6_2),.dout(w_dff_B_cGnUEqZN1_2),.clk(gclk));
	jdff dff_B_TULUFHFB5_2(.din(w_dff_B_cGnUEqZN1_2),.dout(w_dff_B_TULUFHFB5_2),.clk(gclk));
	jdff dff_B_mAr4DQtM5_2(.din(w_dff_B_TULUFHFB5_2),.dout(w_dff_B_mAr4DQtM5_2),.clk(gclk));
	jdff dff_B_IzK4a4Es8_2(.din(w_dff_B_mAr4DQtM5_2),.dout(w_dff_B_IzK4a4Es8_2),.clk(gclk));
	jdff dff_B_hS6AMZ2m3_2(.din(w_dff_B_IzK4a4Es8_2),.dout(w_dff_B_hS6AMZ2m3_2),.clk(gclk));
	jdff dff_B_y0ItLKzh4_2(.din(n923),.dout(w_dff_B_y0ItLKzh4_2),.clk(gclk));
	jdff dff_B_Dwps49C11_1(.din(n852),.dout(w_dff_B_Dwps49C11_1),.clk(gclk));
	jdff dff_B_LnBYv4ut4_2(.din(n752),.dout(w_dff_B_LnBYv4ut4_2),.clk(gclk));
	jdff dff_B_MRdZLkga7_2(.din(w_dff_B_LnBYv4ut4_2),.dout(w_dff_B_MRdZLkga7_2),.clk(gclk));
	jdff dff_B_Qv2GJThw2_2(.din(w_dff_B_MRdZLkga7_2),.dout(w_dff_B_Qv2GJThw2_2),.clk(gclk));
	jdff dff_B_AUs6zmqn3_2(.din(w_dff_B_Qv2GJThw2_2),.dout(w_dff_B_AUs6zmqn3_2),.clk(gclk));
	jdff dff_B_BgdQMJFT1_2(.din(w_dff_B_AUs6zmqn3_2),.dout(w_dff_B_BgdQMJFT1_2),.clk(gclk));
	jdff dff_B_4ATcdP1I6_2(.din(w_dff_B_BgdQMJFT1_2),.dout(w_dff_B_4ATcdP1I6_2),.clk(gclk));
	jdff dff_B_EPcGaCRJ9_2(.din(w_dff_B_4ATcdP1I6_2),.dout(w_dff_B_EPcGaCRJ9_2),.clk(gclk));
	jdff dff_B_b9YLYGBa5_2(.din(w_dff_B_EPcGaCRJ9_2),.dout(w_dff_B_b9YLYGBa5_2),.clk(gclk));
	jdff dff_B_VXtbv3575_2(.din(w_dff_B_b9YLYGBa5_2),.dout(w_dff_B_VXtbv3575_2),.clk(gclk));
	jdff dff_B_5riRUXIX6_2(.din(w_dff_B_VXtbv3575_2),.dout(w_dff_B_5riRUXIX6_2),.clk(gclk));
	jdff dff_B_GYAY10FO0_2(.din(w_dff_B_5riRUXIX6_2),.dout(w_dff_B_GYAY10FO0_2),.clk(gclk));
	jdff dff_B_quLp7gEl4_2(.din(w_dff_B_GYAY10FO0_2),.dout(w_dff_B_quLp7gEl4_2),.clk(gclk));
	jdff dff_B_ygIfWRUg1_2(.din(w_dff_B_quLp7gEl4_2),.dout(w_dff_B_ygIfWRUg1_2),.clk(gclk));
	jdff dff_B_M1W2GrJw3_2(.din(w_dff_B_ygIfWRUg1_2),.dout(w_dff_B_M1W2GrJw3_2),.clk(gclk));
	jdff dff_B_cXqLT28b1_2(.din(w_dff_B_M1W2GrJw3_2),.dout(w_dff_B_cXqLT28b1_2),.clk(gclk));
	jdff dff_B_ZaJZXSuO1_2(.din(w_dff_B_cXqLT28b1_2),.dout(w_dff_B_ZaJZXSuO1_2),.clk(gclk));
	jdff dff_B_1cObaf4I7_2(.din(w_dff_B_ZaJZXSuO1_2),.dout(w_dff_B_1cObaf4I7_2),.clk(gclk));
	jdff dff_B_P6bPwYBd5_2(.din(w_dff_B_1cObaf4I7_2),.dout(w_dff_B_P6bPwYBd5_2),.clk(gclk));
	jdff dff_B_k67Jsa5P8_2(.din(w_dff_B_P6bPwYBd5_2),.dout(w_dff_B_k67Jsa5P8_2),.clk(gclk));
	jdff dff_B_u9uXpZsG0_2(.din(w_dff_B_k67Jsa5P8_2),.dout(w_dff_B_u9uXpZsG0_2),.clk(gclk));
	jdff dff_B_WbeRbB8t3_2(.din(w_dff_B_u9uXpZsG0_2),.dout(w_dff_B_WbeRbB8t3_2),.clk(gclk));
	jdff dff_B_RDibWo8g7_2(.din(w_dff_B_WbeRbB8t3_2),.dout(w_dff_B_RDibWo8g7_2),.clk(gclk));
	jdff dff_B_Ttu6j5n41_2(.din(w_dff_B_RDibWo8g7_2),.dout(w_dff_B_Ttu6j5n41_2),.clk(gclk));
	jdff dff_B_mBkjRJXv2_2(.din(w_dff_B_Ttu6j5n41_2),.dout(w_dff_B_mBkjRJXv2_2),.clk(gclk));
	jdff dff_B_I9S76K1N0_2(.din(w_dff_B_mBkjRJXv2_2),.dout(w_dff_B_I9S76K1N0_2),.clk(gclk));
	jdff dff_B_DtafXJMb0_2(.din(w_dff_B_I9S76K1N0_2),.dout(w_dff_B_DtafXJMb0_2),.clk(gclk));
	jdff dff_B_u96r5TEf0_2(.din(w_dff_B_DtafXJMb0_2),.dout(w_dff_B_u96r5TEf0_2),.clk(gclk));
	jdff dff_B_s1oEiOdU9_2(.din(w_dff_B_u96r5TEf0_2),.dout(w_dff_B_s1oEiOdU9_2),.clk(gclk));
	jdff dff_B_sJWUG6142_2(.din(n817),.dout(w_dff_B_sJWUG6142_2),.clk(gclk));
	jdff dff_B_ZjSS2dJ77_1(.din(n753),.dout(w_dff_B_ZjSS2dJ77_1),.clk(gclk));
	jdff dff_B_OovdVmMD9_2(.din(n659),.dout(w_dff_B_OovdVmMD9_2),.clk(gclk));
	jdff dff_B_mbrfkRjZ6_2(.din(w_dff_B_OovdVmMD9_2),.dout(w_dff_B_mbrfkRjZ6_2),.clk(gclk));
	jdff dff_B_ph9WnQB71_2(.din(w_dff_B_mbrfkRjZ6_2),.dout(w_dff_B_ph9WnQB71_2),.clk(gclk));
	jdff dff_B_2hCHuFoX9_2(.din(w_dff_B_ph9WnQB71_2),.dout(w_dff_B_2hCHuFoX9_2),.clk(gclk));
	jdff dff_B_jyrAqK5y4_2(.din(w_dff_B_2hCHuFoX9_2),.dout(w_dff_B_jyrAqK5y4_2),.clk(gclk));
	jdff dff_B_kFs4xjBA9_2(.din(w_dff_B_jyrAqK5y4_2),.dout(w_dff_B_kFs4xjBA9_2),.clk(gclk));
	jdff dff_B_P6mMWZoB0_2(.din(w_dff_B_kFs4xjBA9_2),.dout(w_dff_B_P6mMWZoB0_2),.clk(gclk));
	jdff dff_B_cIFSHJkA6_2(.din(w_dff_B_P6mMWZoB0_2),.dout(w_dff_B_cIFSHJkA6_2),.clk(gclk));
	jdff dff_B_5h9pYmoR2_2(.din(w_dff_B_cIFSHJkA6_2),.dout(w_dff_B_5h9pYmoR2_2),.clk(gclk));
	jdff dff_B_LWGaaqau1_2(.din(w_dff_B_5h9pYmoR2_2),.dout(w_dff_B_LWGaaqau1_2),.clk(gclk));
	jdff dff_B_sTiLKptz2_2(.din(w_dff_B_LWGaaqau1_2),.dout(w_dff_B_sTiLKptz2_2),.clk(gclk));
	jdff dff_B_4QxDY0h17_2(.din(w_dff_B_sTiLKptz2_2),.dout(w_dff_B_4QxDY0h17_2),.clk(gclk));
	jdff dff_B_fs4NH9nC7_2(.din(w_dff_B_4QxDY0h17_2),.dout(w_dff_B_fs4NH9nC7_2),.clk(gclk));
	jdff dff_B_gLHlhhrj7_2(.din(w_dff_B_fs4NH9nC7_2),.dout(w_dff_B_gLHlhhrj7_2),.clk(gclk));
	jdff dff_B_CzNupRbp4_2(.din(w_dff_B_gLHlhhrj7_2),.dout(w_dff_B_CzNupRbp4_2),.clk(gclk));
	jdff dff_B_MdoKOw5Z7_2(.din(w_dff_B_CzNupRbp4_2),.dout(w_dff_B_MdoKOw5Z7_2),.clk(gclk));
	jdff dff_B_uM6XrG4b9_2(.din(w_dff_B_MdoKOw5Z7_2),.dout(w_dff_B_uM6XrG4b9_2),.clk(gclk));
	jdff dff_B_1aPqaaPW2_2(.din(w_dff_B_uM6XrG4b9_2),.dout(w_dff_B_1aPqaaPW2_2),.clk(gclk));
	jdff dff_B_j7IJ6u3j3_2(.din(w_dff_B_1aPqaaPW2_2),.dout(w_dff_B_j7IJ6u3j3_2),.clk(gclk));
	jdff dff_B_oaqFlQSI1_2(.din(w_dff_B_j7IJ6u3j3_2),.dout(w_dff_B_oaqFlQSI1_2),.clk(gclk));
	jdff dff_B_oFe5B9XV2_2(.din(w_dff_B_oaqFlQSI1_2),.dout(w_dff_B_oFe5B9XV2_2),.clk(gclk));
	jdff dff_B_BwPWjQ027_2(.din(w_dff_B_oFe5B9XV2_2),.dout(w_dff_B_BwPWjQ027_2),.clk(gclk));
	jdff dff_B_XFwmC7VM9_2(.din(w_dff_B_BwPWjQ027_2),.dout(w_dff_B_XFwmC7VM9_2),.clk(gclk));
	jdff dff_B_5z3krZC54_2(.din(w_dff_B_XFwmC7VM9_2),.dout(w_dff_B_5z3krZC54_2),.clk(gclk));
	jdff dff_B_1yZeRs0z3_2(.din(w_dff_B_5z3krZC54_2),.dout(w_dff_B_1yZeRs0z3_2),.clk(gclk));
	jdff dff_B_wQdkmXAX3_2(.din(n717),.dout(w_dff_B_wQdkmXAX3_2),.clk(gclk));
	jdff dff_B_PxDcOGDe3_1(.din(n660),.dout(w_dff_B_PxDcOGDe3_1),.clk(gclk));
	jdff dff_B_JZ8SG1Fu1_2(.din(n573),.dout(w_dff_B_JZ8SG1Fu1_2),.clk(gclk));
	jdff dff_B_p8YDnsjB4_2(.din(w_dff_B_JZ8SG1Fu1_2),.dout(w_dff_B_p8YDnsjB4_2),.clk(gclk));
	jdff dff_B_zd57863Y5_2(.din(w_dff_B_p8YDnsjB4_2),.dout(w_dff_B_zd57863Y5_2),.clk(gclk));
	jdff dff_B_Ir1YAI7m4_2(.din(w_dff_B_zd57863Y5_2),.dout(w_dff_B_Ir1YAI7m4_2),.clk(gclk));
	jdff dff_B_03C02Cah2_2(.din(w_dff_B_Ir1YAI7m4_2),.dout(w_dff_B_03C02Cah2_2),.clk(gclk));
	jdff dff_B_yvtZqhmy4_2(.din(w_dff_B_03C02Cah2_2),.dout(w_dff_B_yvtZqhmy4_2),.clk(gclk));
	jdff dff_B_p8HTkv9f6_2(.din(w_dff_B_yvtZqhmy4_2),.dout(w_dff_B_p8HTkv9f6_2),.clk(gclk));
	jdff dff_B_dt2I0D6d6_2(.din(w_dff_B_p8HTkv9f6_2),.dout(w_dff_B_dt2I0D6d6_2),.clk(gclk));
	jdff dff_B_umRCVLAJ1_2(.din(w_dff_B_dt2I0D6d6_2),.dout(w_dff_B_umRCVLAJ1_2),.clk(gclk));
	jdff dff_B_7qArkClW9_2(.din(w_dff_B_umRCVLAJ1_2),.dout(w_dff_B_7qArkClW9_2),.clk(gclk));
	jdff dff_B_myxRQu1h0_2(.din(w_dff_B_7qArkClW9_2),.dout(w_dff_B_myxRQu1h0_2),.clk(gclk));
	jdff dff_B_aurLMFSO6_2(.din(w_dff_B_myxRQu1h0_2),.dout(w_dff_B_aurLMFSO6_2),.clk(gclk));
	jdff dff_B_w5XKOL2x8_2(.din(w_dff_B_aurLMFSO6_2),.dout(w_dff_B_w5XKOL2x8_2),.clk(gclk));
	jdff dff_B_t0ytvEDT6_2(.din(w_dff_B_w5XKOL2x8_2),.dout(w_dff_B_t0ytvEDT6_2),.clk(gclk));
	jdff dff_B_IiC9sOro1_2(.din(w_dff_B_t0ytvEDT6_2),.dout(w_dff_B_IiC9sOro1_2),.clk(gclk));
	jdff dff_B_Z95Fs6UR2_2(.din(w_dff_B_IiC9sOro1_2),.dout(w_dff_B_Z95Fs6UR2_2),.clk(gclk));
	jdff dff_B_M4r6nRbe2_2(.din(w_dff_B_Z95Fs6UR2_2),.dout(w_dff_B_M4r6nRbe2_2),.clk(gclk));
	jdff dff_B_vCcrBO4m3_2(.din(w_dff_B_M4r6nRbe2_2),.dout(w_dff_B_vCcrBO4m3_2),.clk(gclk));
	jdff dff_B_MoG9zz6F2_2(.din(w_dff_B_vCcrBO4m3_2),.dout(w_dff_B_MoG9zz6F2_2),.clk(gclk));
	jdff dff_B_bJtg3bdA2_2(.din(w_dff_B_MoG9zz6F2_2),.dout(w_dff_B_bJtg3bdA2_2),.clk(gclk));
	jdff dff_B_YnVZirDT9_2(.din(w_dff_B_bJtg3bdA2_2),.dout(w_dff_B_YnVZirDT9_2),.clk(gclk));
	jdff dff_B_X1JJlNGf9_2(.din(w_dff_B_YnVZirDT9_2),.dout(w_dff_B_X1JJlNGf9_2),.clk(gclk));
	jdff dff_B_TuOrFy6A8_2(.din(n624),.dout(w_dff_B_TuOrFy6A8_2),.clk(gclk));
	jdff dff_B_8DXc4VHP2_1(.din(n574),.dout(w_dff_B_8DXc4VHP2_1),.clk(gclk));
	jdff dff_B_oIsN6uep7_2(.din(n494),.dout(w_dff_B_oIsN6uep7_2),.clk(gclk));
	jdff dff_B_Ih5CN3Tj0_2(.din(w_dff_B_oIsN6uep7_2),.dout(w_dff_B_Ih5CN3Tj0_2),.clk(gclk));
	jdff dff_B_4kcX0mzb1_2(.din(w_dff_B_Ih5CN3Tj0_2),.dout(w_dff_B_4kcX0mzb1_2),.clk(gclk));
	jdff dff_B_ZvltgaRF3_2(.din(w_dff_B_4kcX0mzb1_2),.dout(w_dff_B_ZvltgaRF3_2),.clk(gclk));
	jdff dff_B_koZp7SGU2_2(.din(w_dff_B_ZvltgaRF3_2),.dout(w_dff_B_koZp7SGU2_2),.clk(gclk));
	jdff dff_B_7kP5wfc11_2(.din(w_dff_B_koZp7SGU2_2),.dout(w_dff_B_7kP5wfc11_2),.clk(gclk));
	jdff dff_B_wR9LdgtU5_2(.din(w_dff_B_7kP5wfc11_2),.dout(w_dff_B_wR9LdgtU5_2),.clk(gclk));
	jdff dff_B_1GTjPDU11_2(.din(w_dff_B_wR9LdgtU5_2),.dout(w_dff_B_1GTjPDU11_2),.clk(gclk));
	jdff dff_B_AeK5lfvI7_2(.din(w_dff_B_1GTjPDU11_2),.dout(w_dff_B_AeK5lfvI7_2),.clk(gclk));
	jdff dff_B_q0iyvY4j2_2(.din(w_dff_B_AeK5lfvI7_2),.dout(w_dff_B_q0iyvY4j2_2),.clk(gclk));
	jdff dff_B_zRi0fW0q7_2(.din(w_dff_B_q0iyvY4j2_2),.dout(w_dff_B_zRi0fW0q7_2),.clk(gclk));
	jdff dff_B_J2u2ttDO0_2(.din(w_dff_B_zRi0fW0q7_2),.dout(w_dff_B_J2u2ttDO0_2),.clk(gclk));
	jdff dff_B_bEtRwI3i2_2(.din(w_dff_B_J2u2ttDO0_2),.dout(w_dff_B_bEtRwI3i2_2),.clk(gclk));
	jdff dff_B_5LR6fvlK2_2(.din(w_dff_B_bEtRwI3i2_2),.dout(w_dff_B_5LR6fvlK2_2),.clk(gclk));
	jdff dff_B_pAFZ88CO8_2(.din(w_dff_B_5LR6fvlK2_2),.dout(w_dff_B_pAFZ88CO8_2),.clk(gclk));
	jdff dff_B_3rWeH4hL8_2(.din(w_dff_B_pAFZ88CO8_2),.dout(w_dff_B_3rWeH4hL8_2),.clk(gclk));
	jdff dff_B_J2hirTEo0_2(.din(w_dff_B_3rWeH4hL8_2),.dout(w_dff_B_J2hirTEo0_2),.clk(gclk));
	jdff dff_B_vJKj6JTm9_2(.din(w_dff_B_J2hirTEo0_2),.dout(w_dff_B_vJKj6JTm9_2),.clk(gclk));
	jdff dff_B_P90XYJTQ4_2(.din(w_dff_B_vJKj6JTm9_2),.dout(w_dff_B_P90XYJTQ4_2),.clk(gclk));
	jdff dff_B_dPQiGyWm2_2(.din(n538),.dout(w_dff_B_dPQiGyWm2_2),.clk(gclk));
	jdff dff_B_UeXsh9uZ9_1(.din(n495),.dout(w_dff_B_UeXsh9uZ9_1),.clk(gclk));
	jdff dff_B_F82px3E89_2(.din(n422),.dout(w_dff_B_F82px3E89_2),.clk(gclk));
	jdff dff_B_Br0cfbnG1_2(.din(w_dff_B_F82px3E89_2),.dout(w_dff_B_Br0cfbnG1_2),.clk(gclk));
	jdff dff_B_pZrQ5QnB7_2(.din(w_dff_B_Br0cfbnG1_2),.dout(w_dff_B_pZrQ5QnB7_2),.clk(gclk));
	jdff dff_B_q9BiA5k03_2(.din(w_dff_B_pZrQ5QnB7_2),.dout(w_dff_B_q9BiA5k03_2),.clk(gclk));
	jdff dff_B_LiQDsVnC5_2(.din(w_dff_B_q9BiA5k03_2),.dout(w_dff_B_LiQDsVnC5_2),.clk(gclk));
	jdff dff_B_G0BU64Od8_2(.din(w_dff_B_LiQDsVnC5_2),.dout(w_dff_B_G0BU64Od8_2),.clk(gclk));
	jdff dff_B_6rtVPpiT1_2(.din(w_dff_B_G0BU64Od8_2),.dout(w_dff_B_6rtVPpiT1_2),.clk(gclk));
	jdff dff_B_2lvusSrS3_2(.din(w_dff_B_6rtVPpiT1_2),.dout(w_dff_B_2lvusSrS3_2),.clk(gclk));
	jdff dff_B_gfQtg04x3_2(.din(w_dff_B_2lvusSrS3_2),.dout(w_dff_B_gfQtg04x3_2),.clk(gclk));
	jdff dff_B_wq79QjT70_2(.din(w_dff_B_gfQtg04x3_2),.dout(w_dff_B_wq79QjT70_2),.clk(gclk));
	jdff dff_B_KViurxnT3_2(.din(w_dff_B_wq79QjT70_2),.dout(w_dff_B_KViurxnT3_2),.clk(gclk));
	jdff dff_B_lRr41Z7I0_2(.din(w_dff_B_KViurxnT3_2),.dout(w_dff_B_lRr41Z7I0_2),.clk(gclk));
	jdff dff_B_Q93eLLWX4_2(.din(w_dff_B_lRr41Z7I0_2),.dout(w_dff_B_Q93eLLWX4_2),.clk(gclk));
	jdff dff_B_IVnHvEPA5_2(.din(w_dff_B_Q93eLLWX4_2),.dout(w_dff_B_IVnHvEPA5_2),.clk(gclk));
	jdff dff_B_9IdZrWbO3_2(.din(w_dff_B_IVnHvEPA5_2),.dout(w_dff_B_9IdZrWbO3_2),.clk(gclk));
	jdff dff_B_bCkENo171_2(.din(w_dff_B_9IdZrWbO3_2),.dout(w_dff_B_bCkENo171_2),.clk(gclk));
	jdff dff_B_joj2jMnZ3_2(.din(n459),.dout(w_dff_B_joj2jMnZ3_2),.clk(gclk));
	jdff dff_B_S3LDvzAM3_1(.din(n423),.dout(w_dff_B_S3LDvzAM3_1),.clk(gclk));
	jdff dff_B_GKexaLQJ6_2(.din(n358),.dout(w_dff_B_GKexaLQJ6_2),.clk(gclk));
	jdff dff_B_Z677QtdV3_2(.din(w_dff_B_GKexaLQJ6_2),.dout(w_dff_B_Z677QtdV3_2),.clk(gclk));
	jdff dff_B_uVB1NLlq7_2(.din(w_dff_B_Z677QtdV3_2),.dout(w_dff_B_uVB1NLlq7_2),.clk(gclk));
	jdff dff_B_Xk1LeGoS3_2(.din(w_dff_B_uVB1NLlq7_2),.dout(w_dff_B_Xk1LeGoS3_2),.clk(gclk));
	jdff dff_B_wPG9Mjms5_2(.din(w_dff_B_Xk1LeGoS3_2),.dout(w_dff_B_wPG9Mjms5_2),.clk(gclk));
	jdff dff_B_uIo3Bg5t1_2(.din(w_dff_B_wPG9Mjms5_2),.dout(w_dff_B_uIo3Bg5t1_2),.clk(gclk));
	jdff dff_B_unD14ByA0_2(.din(w_dff_B_uIo3Bg5t1_2),.dout(w_dff_B_unD14ByA0_2),.clk(gclk));
	jdff dff_B_P4FCEVZp9_2(.din(w_dff_B_unD14ByA0_2),.dout(w_dff_B_P4FCEVZp9_2),.clk(gclk));
	jdff dff_B_bPnAOKI30_2(.din(w_dff_B_P4FCEVZp9_2),.dout(w_dff_B_bPnAOKI30_2),.clk(gclk));
	jdff dff_B_l01mquOU9_2(.din(w_dff_B_bPnAOKI30_2),.dout(w_dff_B_l01mquOU9_2),.clk(gclk));
	jdff dff_B_7tYK5xUI4_2(.din(w_dff_B_l01mquOU9_2),.dout(w_dff_B_7tYK5xUI4_2),.clk(gclk));
	jdff dff_B_PA96h7SR8_2(.din(w_dff_B_7tYK5xUI4_2),.dout(w_dff_B_PA96h7SR8_2),.clk(gclk));
	jdff dff_B_d7k18fMk7_2(.din(w_dff_B_PA96h7SR8_2),.dout(w_dff_B_d7k18fMk7_2),.clk(gclk));
	jdff dff_B_OSIDnEiA1_2(.din(n387),.dout(w_dff_B_OSIDnEiA1_2),.clk(gclk));
	jdff dff_B_OnsABkWv7_1(.din(n359),.dout(w_dff_B_OnsABkWv7_1),.clk(gclk));
	jdff dff_B_1vjrn6XB0_2(.din(n300),.dout(w_dff_B_1vjrn6XB0_2),.clk(gclk));
	jdff dff_B_RVQJDNk02_2(.din(w_dff_B_1vjrn6XB0_2),.dout(w_dff_B_RVQJDNk02_2),.clk(gclk));
	jdff dff_B_U01tVpCE9_2(.din(w_dff_B_RVQJDNk02_2),.dout(w_dff_B_U01tVpCE9_2),.clk(gclk));
	jdff dff_B_AZjQPbyp1_2(.din(w_dff_B_U01tVpCE9_2),.dout(w_dff_B_AZjQPbyp1_2),.clk(gclk));
	jdff dff_B_pQJyU4jZ5_2(.din(w_dff_B_AZjQPbyp1_2),.dout(w_dff_B_pQJyU4jZ5_2),.clk(gclk));
	jdff dff_B_alz9Qaub2_2(.din(w_dff_B_pQJyU4jZ5_2),.dout(w_dff_B_alz9Qaub2_2),.clk(gclk));
	jdff dff_B_qcvaPbNc8_2(.din(w_dff_B_alz9Qaub2_2),.dout(w_dff_B_qcvaPbNc8_2),.clk(gclk));
	jdff dff_B_de23805L4_2(.din(w_dff_B_qcvaPbNc8_2),.dout(w_dff_B_de23805L4_2),.clk(gclk));
	jdff dff_B_G6F0HEmv0_2(.din(w_dff_B_de23805L4_2),.dout(w_dff_B_G6F0HEmv0_2),.clk(gclk));
	jdff dff_B_gwbk1L7D7_2(.din(w_dff_B_G6F0HEmv0_2),.dout(w_dff_B_gwbk1L7D7_2),.clk(gclk));
	jdff dff_B_in7sRfZw5_2(.din(n323),.dout(w_dff_B_in7sRfZw5_2),.clk(gclk));
	jdff dff_B_OkUzAfi64_1(.din(n301),.dout(w_dff_B_OkUzAfi64_1),.clk(gclk));
	jdff dff_B_uO7Gtbni9_2(.din(n249),.dout(w_dff_B_uO7Gtbni9_2),.clk(gclk));
	jdff dff_B_2YxeOzGf2_2(.din(w_dff_B_uO7Gtbni9_2),.dout(w_dff_B_2YxeOzGf2_2),.clk(gclk));
	jdff dff_B_iQHxFL9o1_2(.din(w_dff_B_2YxeOzGf2_2),.dout(w_dff_B_iQHxFL9o1_2),.clk(gclk));
	jdff dff_B_ObLDN0uT1_2(.din(w_dff_B_iQHxFL9o1_2),.dout(w_dff_B_ObLDN0uT1_2),.clk(gclk));
	jdff dff_B_GvXDFjLQ8_2(.din(w_dff_B_ObLDN0uT1_2),.dout(w_dff_B_GvXDFjLQ8_2),.clk(gclk));
	jdff dff_B_cFWyPtRn7_2(.din(w_dff_B_GvXDFjLQ8_2),.dout(w_dff_B_cFWyPtRn7_2),.clk(gclk));
	jdff dff_B_60eohaZi9_2(.din(w_dff_B_cFWyPtRn7_2),.dout(w_dff_B_60eohaZi9_2),.clk(gclk));
	jdff dff_B_2ccDlXr84_2(.din(n265),.dout(w_dff_B_2ccDlXr84_2),.clk(gclk));
	jdff dff_B_f4uAbTBS5_1(.din(n250),.dout(w_dff_B_f4uAbTBS5_1),.clk(gclk));
	jdff dff_B_KeyIPZfW7_0(.din(n214),.dout(w_dff_B_KeyIPZfW7_0),.clk(gclk));
	jdff dff_B_ipChMsk04_2(.din(n206),.dout(w_dff_B_ipChMsk04_2),.clk(gclk));
	jdff dff_B_AIGDCwhD8_2(.din(w_dff_B_ipChMsk04_2),.dout(w_dff_B_AIGDCwhD8_2),.clk(gclk));
	jdff dff_B_zmvDwT8o8_2(.din(w_dff_B_AIGDCwhD8_2),.dout(w_dff_B_zmvDwT8o8_2),.clk(gclk));
	jdff dff_B_eL30RuV68_2(.din(w_dff_B_zmvDwT8o8_2),.dout(w_dff_B_eL30RuV68_2),.clk(gclk));
	jdff dff_B_x3G1lenS0_1(.din(n208),.dout(w_dff_B_x3G1lenS0_1),.clk(gclk));
	jdff dff_A_ab6agvHO7_0(.dout(w_n210_1[0]),.din(w_dff_A_ab6agvHO7_0),.clk(gclk));
	jdff dff_A_SLtjRVKq4_0(.dout(w_n169_0[0]),.din(w_dff_A_SLtjRVKq4_0),.clk(gclk));
	jdff dff_A_a8R000an1_0(.dout(w_dff_A_SLtjRVKq4_0),.din(w_dff_A_a8R000an1_0),.clk(gclk));
	jdff dff_A_gZCz23As0_1(.dout(w_n169_0[1]),.din(w_dff_A_gZCz23As0_1),.clk(gclk));
	jdff dff_B_Cngn24uH1_2(.din(n1420),.dout(w_dff_B_Cngn24uH1_2),.clk(gclk));
	jdff dff_B_3bupPnHd6_1(.din(n1418),.dout(w_dff_B_3bupPnHd6_1),.clk(gclk));
	jdff dff_B_aZ3jnh142_2(.din(n1338),.dout(w_dff_B_aZ3jnh142_2),.clk(gclk));
	jdff dff_B_vtqBcY7A7_2(.din(w_dff_B_aZ3jnh142_2),.dout(w_dff_B_vtqBcY7A7_2),.clk(gclk));
	jdff dff_B_bmTkb4Q08_2(.din(w_dff_B_vtqBcY7A7_2),.dout(w_dff_B_bmTkb4Q08_2),.clk(gclk));
	jdff dff_B_8HMpiAWT9_2(.din(w_dff_B_bmTkb4Q08_2),.dout(w_dff_B_8HMpiAWT9_2),.clk(gclk));
	jdff dff_B_oxlVLBY17_2(.din(w_dff_B_8HMpiAWT9_2),.dout(w_dff_B_oxlVLBY17_2),.clk(gclk));
	jdff dff_B_oJ57Udyv6_2(.din(w_dff_B_oxlVLBY17_2),.dout(w_dff_B_oJ57Udyv6_2),.clk(gclk));
	jdff dff_B_tB2jw37h8_2(.din(w_dff_B_oJ57Udyv6_2),.dout(w_dff_B_tB2jw37h8_2),.clk(gclk));
	jdff dff_B_dXUyMAfa5_2(.din(w_dff_B_tB2jw37h8_2),.dout(w_dff_B_dXUyMAfa5_2),.clk(gclk));
	jdff dff_B_7U5BNE2h3_2(.din(w_dff_B_dXUyMAfa5_2),.dout(w_dff_B_7U5BNE2h3_2),.clk(gclk));
	jdff dff_B_vT7X76Rv3_2(.din(w_dff_B_7U5BNE2h3_2),.dout(w_dff_B_vT7X76Rv3_2),.clk(gclk));
	jdff dff_B_zny6G3B55_2(.din(w_dff_B_vT7X76Rv3_2),.dout(w_dff_B_zny6G3B55_2),.clk(gclk));
	jdff dff_B_mR0cDyN53_2(.din(w_dff_B_zny6G3B55_2),.dout(w_dff_B_mR0cDyN53_2),.clk(gclk));
	jdff dff_B_2TyaRKCI0_2(.din(w_dff_B_mR0cDyN53_2),.dout(w_dff_B_2TyaRKCI0_2),.clk(gclk));
	jdff dff_B_NJOjni0j8_2(.din(w_dff_B_2TyaRKCI0_2),.dout(w_dff_B_NJOjni0j8_2),.clk(gclk));
	jdff dff_B_DRfNpyRh3_2(.din(w_dff_B_NJOjni0j8_2),.dout(w_dff_B_DRfNpyRh3_2),.clk(gclk));
	jdff dff_B_GmYBuXMx6_2(.din(w_dff_B_DRfNpyRh3_2),.dout(w_dff_B_GmYBuXMx6_2),.clk(gclk));
	jdff dff_B_ob7u66dA5_2(.din(w_dff_B_GmYBuXMx6_2),.dout(w_dff_B_ob7u66dA5_2),.clk(gclk));
	jdff dff_B_g1bXdf332_2(.din(w_dff_B_ob7u66dA5_2),.dout(w_dff_B_g1bXdf332_2),.clk(gclk));
	jdff dff_B_xcT8Hw5A6_2(.din(w_dff_B_g1bXdf332_2),.dout(w_dff_B_xcT8Hw5A6_2),.clk(gclk));
	jdff dff_B_JNoD57bK9_2(.din(w_dff_B_xcT8Hw5A6_2),.dout(w_dff_B_JNoD57bK9_2),.clk(gclk));
	jdff dff_B_P4IWm8Lw4_2(.din(w_dff_B_JNoD57bK9_2),.dout(w_dff_B_P4IWm8Lw4_2),.clk(gclk));
	jdff dff_B_t7xLGml19_2(.din(w_dff_B_P4IWm8Lw4_2),.dout(w_dff_B_t7xLGml19_2),.clk(gclk));
	jdff dff_B_u2nNLLRN7_2(.din(w_dff_B_t7xLGml19_2),.dout(w_dff_B_u2nNLLRN7_2),.clk(gclk));
	jdff dff_B_h90Ymaf81_2(.din(w_dff_B_u2nNLLRN7_2),.dout(w_dff_B_h90Ymaf81_2),.clk(gclk));
	jdff dff_B_RmhpkNBi2_2(.din(w_dff_B_h90Ymaf81_2),.dout(w_dff_B_RmhpkNBi2_2),.clk(gclk));
	jdff dff_B_Cb2JB3eH4_2(.din(w_dff_B_RmhpkNBi2_2),.dout(w_dff_B_Cb2JB3eH4_2),.clk(gclk));
	jdff dff_B_DlERetDA5_2(.din(w_dff_B_Cb2JB3eH4_2),.dout(w_dff_B_DlERetDA5_2),.clk(gclk));
	jdff dff_B_AtO0RiFG2_2(.din(w_dff_B_DlERetDA5_2),.dout(w_dff_B_AtO0RiFG2_2),.clk(gclk));
	jdff dff_B_cPKFPiaE4_2(.din(w_dff_B_AtO0RiFG2_2),.dout(w_dff_B_cPKFPiaE4_2),.clk(gclk));
	jdff dff_B_5bqZ0WpY3_2(.din(w_dff_B_cPKFPiaE4_2),.dout(w_dff_B_5bqZ0WpY3_2),.clk(gclk));
	jdff dff_B_p8vXaVt50_2(.din(w_dff_B_5bqZ0WpY3_2),.dout(w_dff_B_p8vXaVt50_2),.clk(gclk));
	jdff dff_B_kX8bOGQ94_2(.din(w_dff_B_p8vXaVt50_2),.dout(w_dff_B_kX8bOGQ94_2),.clk(gclk));
	jdff dff_B_8lO6u5X73_2(.din(w_dff_B_kX8bOGQ94_2),.dout(w_dff_B_8lO6u5X73_2),.clk(gclk));
	jdff dff_B_NvdEGkyk9_2(.din(w_dff_B_8lO6u5X73_2),.dout(w_dff_B_NvdEGkyk9_2),.clk(gclk));
	jdff dff_B_xto9W2mR5_2(.din(w_dff_B_NvdEGkyk9_2),.dout(w_dff_B_xto9W2mR5_2),.clk(gclk));
	jdff dff_B_vRuAq3F79_2(.din(w_dff_B_xto9W2mR5_2),.dout(w_dff_B_vRuAq3F79_2),.clk(gclk));
	jdff dff_B_OQkdBmkH5_2(.din(w_dff_B_vRuAq3F79_2),.dout(w_dff_B_OQkdBmkH5_2),.clk(gclk));
	jdff dff_B_gBTA61rt3_2(.din(w_dff_B_OQkdBmkH5_2),.dout(w_dff_B_gBTA61rt3_2),.clk(gclk));
	jdff dff_B_GYWVTZGF9_2(.din(w_dff_B_gBTA61rt3_2),.dout(w_dff_B_GYWVTZGF9_2),.clk(gclk));
	jdff dff_B_fPrVdaRI2_2(.din(w_dff_B_GYWVTZGF9_2),.dout(w_dff_B_fPrVdaRI2_2),.clk(gclk));
	jdff dff_B_d3KbCPHj1_2(.din(w_dff_B_fPrVdaRI2_2),.dout(w_dff_B_d3KbCPHj1_2),.clk(gclk));
	jdff dff_B_0LAtOIli8_2(.din(w_dff_B_d3KbCPHj1_2),.dout(w_dff_B_0LAtOIli8_2),.clk(gclk));
	jdff dff_B_Fn2HwZ4t2_2(.din(w_dff_B_0LAtOIli8_2),.dout(w_dff_B_Fn2HwZ4t2_2),.clk(gclk));
	jdff dff_B_wfVjBIIC1_2(.din(w_dff_B_Fn2HwZ4t2_2),.dout(w_dff_B_wfVjBIIC1_2),.clk(gclk));
	jdff dff_B_1eQL6QIs8_2(.din(w_dff_B_wfVjBIIC1_2),.dout(w_dff_B_1eQL6QIs8_2),.clk(gclk));
	jdff dff_B_j079FCM32_1(.din(n1339),.dout(w_dff_B_j079FCM32_1),.clk(gclk));
	jdff dff_B_PI422c360_2(.din(n1253),.dout(w_dff_B_PI422c360_2),.clk(gclk));
	jdff dff_B_0k1qYqts8_2(.din(w_dff_B_PI422c360_2),.dout(w_dff_B_0k1qYqts8_2),.clk(gclk));
	jdff dff_B_n4X64WQn4_2(.din(w_dff_B_0k1qYqts8_2),.dout(w_dff_B_n4X64WQn4_2),.clk(gclk));
	jdff dff_B_fkPcQl4o1_2(.din(w_dff_B_n4X64WQn4_2),.dout(w_dff_B_fkPcQl4o1_2),.clk(gclk));
	jdff dff_B_PpdQCT3Z0_2(.din(w_dff_B_fkPcQl4o1_2),.dout(w_dff_B_PpdQCT3Z0_2),.clk(gclk));
	jdff dff_B_8hCRoQ5t5_2(.din(w_dff_B_PpdQCT3Z0_2),.dout(w_dff_B_8hCRoQ5t5_2),.clk(gclk));
	jdff dff_B_APuEXC5e9_2(.din(w_dff_B_8hCRoQ5t5_2),.dout(w_dff_B_APuEXC5e9_2),.clk(gclk));
	jdff dff_B_GbCPCTYz1_2(.din(w_dff_B_APuEXC5e9_2),.dout(w_dff_B_GbCPCTYz1_2),.clk(gclk));
	jdff dff_B_K7jJE0Jy3_2(.din(w_dff_B_GbCPCTYz1_2),.dout(w_dff_B_K7jJE0Jy3_2),.clk(gclk));
	jdff dff_B_3TK67x301_2(.din(w_dff_B_K7jJE0Jy3_2),.dout(w_dff_B_3TK67x301_2),.clk(gclk));
	jdff dff_B_v5NBp9iH1_2(.din(w_dff_B_3TK67x301_2),.dout(w_dff_B_v5NBp9iH1_2),.clk(gclk));
	jdff dff_B_Y7fFNuvr6_2(.din(w_dff_B_v5NBp9iH1_2),.dout(w_dff_B_Y7fFNuvr6_2),.clk(gclk));
	jdff dff_B_Eu5KtEvZ1_2(.din(w_dff_B_Y7fFNuvr6_2),.dout(w_dff_B_Eu5KtEvZ1_2),.clk(gclk));
	jdff dff_B_aueFfBGV6_2(.din(w_dff_B_Eu5KtEvZ1_2),.dout(w_dff_B_aueFfBGV6_2),.clk(gclk));
	jdff dff_B_tQZZZIRE0_2(.din(w_dff_B_aueFfBGV6_2),.dout(w_dff_B_tQZZZIRE0_2),.clk(gclk));
	jdff dff_B_HQV4qQML0_2(.din(w_dff_B_tQZZZIRE0_2),.dout(w_dff_B_HQV4qQML0_2),.clk(gclk));
	jdff dff_B_0fbb3tXx2_2(.din(w_dff_B_HQV4qQML0_2),.dout(w_dff_B_0fbb3tXx2_2),.clk(gclk));
	jdff dff_B_1FHJatrq9_2(.din(w_dff_B_0fbb3tXx2_2),.dout(w_dff_B_1FHJatrq9_2),.clk(gclk));
	jdff dff_B_vi3PR3DX7_2(.din(w_dff_B_1FHJatrq9_2),.dout(w_dff_B_vi3PR3DX7_2),.clk(gclk));
	jdff dff_B_XuLUhRgw8_2(.din(w_dff_B_vi3PR3DX7_2),.dout(w_dff_B_XuLUhRgw8_2),.clk(gclk));
	jdff dff_B_Mvz7x8wc9_2(.din(w_dff_B_XuLUhRgw8_2),.dout(w_dff_B_Mvz7x8wc9_2),.clk(gclk));
	jdff dff_B_zAgSOMbJ1_2(.din(w_dff_B_Mvz7x8wc9_2),.dout(w_dff_B_zAgSOMbJ1_2),.clk(gclk));
	jdff dff_B_LEZ89wzN3_2(.din(w_dff_B_zAgSOMbJ1_2),.dout(w_dff_B_LEZ89wzN3_2),.clk(gclk));
	jdff dff_B_NOF0MlVd2_2(.din(w_dff_B_LEZ89wzN3_2),.dout(w_dff_B_NOF0MlVd2_2),.clk(gclk));
	jdff dff_B_gnkp2g2F3_2(.din(w_dff_B_NOF0MlVd2_2),.dout(w_dff_B_gnkp2g2F3_2),.clk(gclk));
	jdff dff_B_WhNPmtF40_2(.din(w_dff_B_gnkp2g2F3_2),.dout(w_dff_B_WhNPmtF40_2),.clk(gclk));
	jdff dff_B_J0cWdLFq7_2(.din(w_dff_B_WhNPmtF40_2),.dout(w_dff_B_J0cWdLFq7_2),.clk(gclk));
	jdff dff_B_cqEnRLDh7_2(.din(w_dff_B_J0cWdLFq7_2),.dout(w_dff_B_cqEnRLDh7_2),.clk(gclk));
	jdff dff_B_7MYw9aY48_2(.din(w_dff_B_cqEnRLDh7_2),.dout(w_dff_B_7MYw9aY48_2),.clk(gclk));
	jdff dff_B_tb6suika7_2(.din(w_dff_B_7MYw9aY48_2),.dout(w_dff_B_tb6suika7_2),.clk(gclk));
	jdff dff_B_xXZRh6PY2_2(.din(w_dff_B_tb6suika7_2),.dout(w_dff_B_xXZRh6PY2_2),.clk(gclk));
	jdff dff_B_TYtpAtfY6_2(.din(w_dff_B_xXZRh6PY2_2),.dout(w_dff_B_TYtpAtfY6_2),.clk(gclk));
	jdff dff_B_aN8JocuM8_2(.din(w_dff_B_TYtpAtfY6_2),.dout(w_dff_B_aN8JocuM8_2),.clk(gclk));
	jdff dff_B_Vq5kSKGY4_2(.din(w_dff_B_aN8JocuM8_2),.dout(w_dff_B_Vq5kSKGY4_2),.clk(gclk));
	jdff dff_B_4gq6v1Mr3_2(.din(w_dff_B_Vq5kSKGY4_2),.dout(w_dff_B_4gq6v1Mr3_2),.clk(gclk));
	jdff dff_B_9AkKwsAe4_2(.din(w_dff_B_4gq6v1Mr3_2),.dout(w_dff_B_9AkKwsAe4_2),.clk(gclk));
	jdff dff_B_POJg5BVq9_2(.din(w_dff_B_9AkKwsAe4_2),.dout(w_dff_B_POJg5BVq9_2),.clk(gclk));
	jdff dff_B_uqq4h8726_2(.din(w_dff_B_POJg5BVq9_2),.dout(w_dff_B_uqq4h8726_2),.clk(gclk));
	jdff dff_B_YfD2Hzhk8_2(.din(w_dff_B_uqq4h8726_2),.dout(w_dff_B_YfD2Hzhk8_2),.clk(gclk));
	jdff dff_B_cOfaW6Mn8_2(.din(w_dff_B_YfD2Hzhk8_2),.dout(w_dff_B_cOfaW6Mn8_2),.clk(gclk));
	jdff dff_B_Ve6XuVT70_1(.din(n1254),.dout(w_dff_B_Ve6XuVT70_1),.clk(gclk));
	jdff dff_B_nfOcNSbU3_2(.din(n1163),.dout(w_dff_B_nfOcNSbU3_2),.clk(gclk));
	jdff dff_B_NTvImXe40_2(.din(w_dff_B_nfOcNSbU3_2),.dout(w_dff_B_NTvImXe40_2),.clk(gclk));
	jdff dff_B_QcKZOX7W0_2(.din(w_dff_B_NTvImXe40_2),.dout(w_dff_B_QcKZOX7W0_2),.clk(gclk));
	jdff dff_B_wmjLikGs7_2(.din(w_dff_B_QcKZOX7W0_2),.dout(w_dff_B_wmjLikGs7_2),.clk(gclk));
	jdff dff_B_Pf16pe8T2_2(.din(w_dff_B_wmjLikGs7_2),.dout(w_dff_B_Pf16pe8T2_2),.clk(gclk));
	jdff dff_B_UvhsvRMM4_2(.din(w_dff_B_Pf16pe8T2_2),.dout(w_dff_B_UvhsvRMM4_2),.clk(gclk));
	jdff dff_B_ojG4mz3I3_2(.din(w_dff_B_UvhsvRMM4_2),.dout(w_dff_B_ojG4mz3I3_2),.clk(gclk));
	jdff dff_B_SkndRomy4_2(.din(w_dff_B_ojG4mz3I3_2),.dout(w_dff_B_SkndRomy4_2),.clk(gclk));
	jdff dff_B_dVZpe6im1_2(.din(w_dff_B_SkndRomy4_2),.dout(w_dff_B_dVZpe6im1_2),.clk(gclk));
	jdff dff_B_yT33qTN85_2(.din(w_dff_B_dVZpe6im1_2),.dout(w_dff_B_yT33qTN85_2),.clk(gclk));
	jdff dff_B_uNT2z6zX7_2(.din(w_dff_B_yT33qTN85_2),.dout(w_dff_B_uNT2z6zX7_2),.clk(gclk));
	jdff dff_B_YL1NPOqU4_2(.din(w_dff_B_uNT2z6zX7_2),.dout(w_dff_B_YL1NPOqU4_2),.clk(gclk));
	jdff dff_B_uBnxwzTY1_2(.din(w_dff_B_YL1NPOqU4_2),.dout(w_dff_B_uBnxwzTY1_2),.clk(gclk));
	jdff dff_B_xGQWlKlm2_2(.din(w_dff_B_uBnxwzTY1_2),.dout(w_dff_B_xGQWlKlm2_2),.clk(gclk));
	jdff dff_B_z5IbGw5I9_2(.din(w_dff_B_xGQWlKlm2_2),.dout(w_dff_B_z5IbGw5I9_2),.clk(gclk));
	jdff dff_B_9YUShBSr9_2(.din(w_dff_B_z5IbGw5I9_2),.dout(w_dff_B_9YUShBSr9_2),.clk(gclk));
	jdff dff_B_B6jRnsGT6_2(.din(w_dff_B_9YUShBSr9_2),.dout(w_dff_B_B6jRnsGT6_2),.clk(gclk));
	jdff dff_B_X6eKo2i10_2(.din(w_dff_B_B6jRnsGT6_2),.dout(w_dff_B_X6eKo2i10_2),.clk(gclk));
	jdff dff_B_lRAPt5F47_2(.din(w_dff_B_X6eKo2i10_2),.dout(w_dff_B_lRAPt5F47_2),.clk(gclk));
	jdff dff_B_4NuHBtki4_2(.din(w_dff_B_lRAPt5F47_2),.dout(w_dff_B_4NuHBtki4_2),.clk(gclk));
	jdff dff_B_Hstqz02F4_2(.din(w_dff_B_4NuHBtki4_2),.dout(w_dff_B_Hstqz02F4_2),.clk(gclk));
	jdff dff_B_7nDGbcRP0_2(.din(w_dff_B_Hstqz02F4_2),.dout(w_dff_B_7nDGbcRP0_2),.clk(gclk));
	jdff dff_B_FxvLFpN11_2(.din(w_dff_B_7nDGbcRP0_2),.dout(w_dff_B_FxvLFpN11_2),.clk(gclk));
	jdff dff_B_o8poyn7j6_2(.din(w_dff_B_FxvLFpN11_2),.dout(w_dff_B_o8poyn7j6_2),.clk(gclk));
	jdff dff_B_sm4MqfOX2_2(.din(w_dff_B_o8poyn7j6_2),.dout(w_dff_B_sm4MqfOX2_2),.clk(gclk));
	jdff dff_B_Xl17A2n18_2(.din(w_dff_B_sm4MqfOX2_2),.dout(w_dff_B_Xl17A2n18_2),.clk(gclk));
	jdff dff_B_9f07JttR6_2(.din(w_dff_B_Xl17A2n18_2),.dout(w_dff_B_9f07JttR6_2),.clk(gclk));
	jdff dff_B_b9V4tXMK4_2(.din(w_dff_B_9f07JttR6_2),.dout(w_dff_B_b9V4tXMK4_2),.clk(gclk));
	jdff dff_B_HUBpYrcV2_2(.din(w_dff_B_b9V4tXMK4_2),.dout(w_dff_B_HUBpYrcV2_2),.clk(gclk));
	jdff dff_B_Ps0V7Caa8_2(.din(w_dff_B_HUBpYrcV2_2),.dout(w_dff_B_Ps0V7Caa8_2),.clk(gclk));
	jdff dff_B_V2RoNlDE6_2(.din(w_dff_B_Ps0V7Caa8_2),.dout(w_dff_B_V2RoNlDE6_2),.clk(gclk));
	jdff dff_B_sVCQM1Ir8_2(.din(w_dff_B_V2RoNlDE6_2),.dout(w_dff_B_sVCQM1Ir8_2),.clk(gclk));
	jdff dff_B_mROPoYsL2_2(.din(w_dff_B_sVCQM1Ir8_2),.dout(w_dff_B_mROPoYsL2_2),.clk(gclk));
	jdff dff_B_h4CYYHiG5_2(.din(w_dff_B_mROPoYsL2_2),.dout(w_dff_B_h4CYYHiG5_2),.clk(gclk));
	jdff dff_B_1PGqQiA23_2(.din(w_dff_B_h4CYYHiG5_2),.dout(w_dff_B_1PGqQiA23_2),.clk(gclk));
	jdff dff_B_YpX0O3M52_2(.din(w_dff_B_1PGqQiA23_2),.dout(w_dff_B_YpX0O3M52_2),.clk(gclk));
	jdff dff_B_7O8tEm8a3_2(.din(w_dff_B_YpX0O3M52_2),.dout(w_dff_B_7O8tEm8a3_2),.clk(gclk));
	jdff dff_B_tzPycaO79_1(.din(n1164),.dout(w_dff_B_tzPycaO79_1),.clk(gclk));
	jdff dff_B_o2go5oBQ2_2(.din(n1059),.dout(w_dff_B_o2go5oBQ2_2),.clk(gclk));
	jdff dff_B_7oH5w5b32_2(.din(w_dff_B_o2go5oBQ2_2),.dout(w_dff_B_7oH5w5b32_2),.clk(gclk));
	jdff dff_B_7vc7kcyo9_2(.din(w_dff_B_7oH5w5b32_2),.dout(w_dff_B_7vc7kcyo9_2),.clk(gclk));
	jdff dff_B_FX0QTQVc8_2(.din(w_dff_B_7vc7kcyo9_2),.dout(w_dff_B_FX0QTQVc8_2),.clk(gclk));
	jdff dff_B_3yEABLAK2_2(.din(w_dff_B_FX0QTQVc8_2),.dout(w_dff_B_3yEABLAK2_2),.clk(gclk));
	jdff dff_B_EzfpCxNI3_2(.din(w_dff_B_3yEABLAK2_2),.dout(w_dff_B_EzfpCxNI3_2),.clk(gclk));
	jdff dff_B_jeQIlDFF1_2(.din(w_dff_B_EzfpCxNI3_2),.dout(w_dff_B_jeQIlDFF1_2),.clk(gclk));
	jdff dff_B_FpXZ0RLg1_2(.din(w_dff_B_jeQIlDFF1_2),.dout(w_dff_B_FpXZ0RLg1_2),.clk(gclk));
	jdff dff_B_mG9kDgzC6_2(.din(w_dff_B_FpXZ0RLg1_2),.dout(w_dff_B_mG9kDgzC6_2),.clk(gclk));
	jdff dff_B_lZg8j7oV9_2(.din(w_dff_B_mG9kDgzC6_2),.dout(w_dff_B_lZg8j7oV9_2),.clk(gclk));
	jdff dff_B_gvRoVTrJ8_2(.din(w_dff_B_lZg8j7oV9_2),.dout(w_dff_B_gvRoVTrJ8_2),.clk(gclk));
	jdff dff_B_Gn0TFo9s3_2(.din(w_dff_B_gvRoVTrJ8_2),.dout(w_dff_B_Gn0TFo9s3_2),.clk(gclk));
	jdff dff_B_LiQhnnfs6_2(.din(w_dff_B_Gn0TFo9s3_2),.dout(w_dff_B_LiQhnnfs6_2),.clk(gclk));
	jdff dff_B_SLIBLd9q1_2(.din(w_dff_B_LiQhnnfs6_2),.dout(w_dff_B_SLIBLd9q1_2),.clk(gclk));
	jdff dff_B_2NbuIvYu0_2(.din(w_dff_B_SLIBLd9q1_2),.dout(w_dff_B_2NbuIvYu0_2),.clk(gclk));
	jdff dff_B_sAiHmYUk3_2(.din(w_dff_B_2NbuIvYu0_2),.dout(w_dff_B_sAiHmYUk3_2),.clk(gclk));
	jdff dff_B_3FM4j2vm9_2(.din(w_dff_B_sAiHmYUk3_2),.dout(w_dff_B_3FM4j2vm9_2),.clk(gclk));
	jdff dff_B_ItvwI4py1_2(.din(w_dff_B_3FM4j2vm9_2),.dout(w_dff_B_ItvwI4py1_2),.clk(gclk));
	jdff dff_B_mDSpuFgx6_2(.din(w_dff_B_ItvwI4py1_2),.dout(w_dff_B_mDSpuFgx6_2),.clk(gclk));
	jdff dff_B_FwMBvBaX3_2(.din(w_dff_B_mDSpuFgx6_2),.dout(w_dff_B_FwMBvBaX3_2),.clk(gclk));
	jdff dff_B_3yNBNeIM2_2(.din(w_dff_B_FwMBvBaX3_2),.dout(w_dff_B_3yNBNeIM2_2),.clk(gclk));
	jdff dff_B_HVNi8iDy8_2(.din(w_dff_B_3yNBNeIM2_2),.dout(w_dff_B_HVNi8iDy8_2),.clk(gclk));
	jdff dff_B_TFLqg0jh5_2(.din(w_dff_B_HVNi8iDy8_2),.dout(w_dff_B_TFLqg0jh5_2),.clk(gclk));
	jdff dff_B_0SAOxi2C2_2(.din(w_dff_B_TFLqg0jh5_2),.dout(w_dff_B_0SAOxi2C2_2),.clk(gclk));
	jdff dff_B_plDDwwII2_2(.din(w_dff_B_0SAOxi2C2_2),.dout(w_dff_B_plDDwwII2_2),.clk(gclk));
	jdff dff_B_ZxBJxJsb5_2(.din(w_dff_B_plDDwwII2_2),.dout(w_dff_B_ZxBJxJsb5_2),.clk(gclk));
	jdff dff_B_5xG3zZT59_2(.din(w_dff_B_ZxBJxJsb5_2),.dout(w_dff_B_5xG3zZT59_2),.clk(gclk));
	jdff dff_B_ednsvzuj3_2(.din(w_dff_B_5xG3zZT59_2),.dout(w_dff_B_ednsvzuj3_2),.clk(gclk));
	jdff dff_B_bqNnc41A2_2(.din(w_dff_B_ednsvzuj3_2),.dout(w_dff_B_bqNnc41A2_2),.clk(gclk));
	jdff dff_B_NUxBqaob5_2(.din(w_dff_B_bqNnc41A2_2),.dout(w_dff_B_NUxBqaob5_2),.clk(gclk));
	jdff dff_B_WYutRZFW9_2(.din(w_dff_B_NUxBqaob5_2),.dout(w_dff_B_WYutRZFW9_2),.clk(gclk));
	jdff dff_B_4955CFnq5_2(.din(w_dff_B_WYutRZFW9_2),.dout(w_dff_B_4955CFnq5_2),.clk(gclk));
	jdff dff_B_3jmo5Plu7_2(.din(w_dff_B_4955CFnq5_2),.dout(w_dff_B_3jmo5Plu7_2),.clk(gclk));
	jdff dff_B_jgMd85UI9_2(.din(w_dff_B_3jmo5Plu7_2),.dout(w_dff_B_jgMd85UI9_2),.clk(gclk));
	jdff dff_B_5zfOOgKH1_1(.din(n1060),.dout(w_dff_B_5zfOOgKH1_1),.clk(gclk));
	jdff dff_B_QIxohLxn2_2(.din(n961),.dout(w_dff_B_QIxohLxn2_2),.clk(gclk));
	jdff dff_B_6hxwt7Fy4_2(.din(w_dff_B_QIxohLxn2_2),.dout(w_dff_B_6hxwt7Fy4_2),.clk(gclk));
	jdff dff_B_3XGwUPQP5_2(.din(w_dff_B_6hxwt7Fy4_2),.dout(w_dff_B_3XGwUPQP5_2),.clk(gclk));
	jdff dff_B_G7giD9hq9_2(.din(w_dff_B_3XGwUPQP5_2),.dout(w_dff_B_G7giD9hq9_2),.clk(gclk));
	jdff dff_B_xToTssDQ7_2(.din(w_dff_B_G7giD9hq9_2),.dout(w_dff_B_xToTssDQ7_2),.clk(gclk));
	jdff dff_B_e5iwbTld5_2(.din(w_dff_B_xToTssDQ7_2),.dout(w_dff_B_e5iwbTld5_2),.clk(gclk));
	jdff dff_B_Gph20BZe6_2(.din(w_dff_B_e5iwbTld5_2),.dout(w_dff_B_Gph20BZe6_2),.clk(gclk));
	jdff dff_B_hyqFPLER3_2(.din(w_dff_B_Gph20BZe6_2),.dout(w_dff_B_hyqFPLER3_2),.clk(gclk));
	jdff dff_B_lA07zuv24_2(.din(w_dff_B_hyqFPLER3_2),.dout(w_dff_B_lA07zuv24_2),.clk(gclk));
	jdff dff_B_wxoAQ9ZA1_2(.din(w_dff_B_lA07zuv24_2),.dout(w_dff_B_wxoAQ9ZA1_2),.clk(gclk));
	jdff dff_B_ujlAmiKJ0_2(.din(w_dff_B_wxoAQ9ZA1_2),.dout(w_dff_B_ujlAmiKJ0_2),.clk(gclk));
	jdff dff_B_sKJQqRI01_2(.din(w_dff_B_ujlAmiKJ0_2),.dout(w_dff_B_sKJQqRI01_2),.clk(gclk));
	jdff dff_B_PUwZJS0q9_2(.din(w_dff_B_sKJQqRI01_2),.dout(w_dff_B_PUwZJS0q9_2),.clk(gclk));
	jdff dff_B_EvvaHqgi8_2(.din(w_dff_B_PUwZJS0q9_2),.dout(w_dff_B_EvvaHqgi8_2),.clk(gclk));
	jdff dff_B_XYBGXCFu3_2(.din(w_dff_B_EvvaHqgi8_2),.dout(w_dff_B_XYBGXCFu3_2),.clk(gclk));
	jdff dff_B_JNYZAVaS6_2(.din(w_dff_B_XYBGXCFu3_2),.dout(w_dff_B_JNYZAVaS6_2),.clk(gclk));
	jdff dff_B_tXoteiTe4_2(.din(w_dff_B_JNYZAVaS6_2),.dout(w_dff_B_tXoteiTe4_2),.clk(gclk));
	jdff dff_B_9Dq2HxPU6_2(.din(w_dff_B_tXoteiTe4_2),.dout(w_dff_B_9Dq2HxPU6_2),.clk(gclk));
	jdff dff_B_jE9CHGHA6_2(.din(w_dff_B_9Dq2HxPU6_2),.dout(w_dff_B_jE9CHGHA6_2),.clk(gclk));
	jdff dff_B_9eHXxFAx0_2(.din(w_dff_B_jE9CHGHA6_2),.dout(w_dff_B_9eHXxFAx0_2),.clk(gclk));
	jdff dff_B_o0Co45uI2_2(.din(w_dff_B_9eHXxFAx0_2),.dout(w_dff_B_o0Co45uI2_2),.clk(gclk));
	jdff dff_B_84v3fYGE8_2(.din(w_dff_B_o0Co45uI2_2),.dout(w_dff_B_84v3fYGE8_2),.clk(gclk));
	jdff dff_B_VwQvWoxP5_2(.din(w_dff_B_84v3fYGE8_2),.dout(w_dff_B_VwQvWoxP5_2),.clk(gclk));
	jdff dff_B_HMMxcNY57_2(.din(w_dff_B_VwQvWoxP5_2),.dout(w_dff_B_HMMxcNY57_2),.clk(gclk));
	jdff dff_B_gE0BVxXE6_2(.din(w_dff_B_HMMxcNY57_2),.dout(w_dff_B_gE0BVxXE6_2),.clk(gclk));
	jdff dff_B_Pf201PmX5_2(.din(w_dff_B_gE0BVxXE6_2),.dout(w_dff_B_Pf201PmX5_2),.clk(gclk));
	jdff dff_B_CRxlwRcg9_2(.din(w_dff_B_Pf201PmX5_2),.dout(w_dff_B_CRxlwRcg9_2),.clk(gclk));
	jdff dff_B_sSNVoSWM0_2(.din(w_dff_B_CRxlwRcg9_2),.dout(w_dff_B_sSNVoSWM0_2),.clk(gclk));
	jdff dff_B_5HPx6JnY1_2(.din(w_dff_B_sSNVoSWM0_2),.dout(w_dff_B_5HPx6JnY1_2),.clk(gclk));
	jdff dff_B_B1c5aMwc9_2(.din(w_dff_B_5HPx6JnY1_2),.dout(w_dff_B_B1c5aMwc9_2),.clk(gclk));
	jdff dff_B_vAKqYFTu3_2(.din(w_dff_B_B1c5aMwc9_2),.dout(w_dff_B_vAKqYFTu3_2),.clk(gclk));
	jdff dff_B_P0j1A7UR7_1(.din(n962),.dout(w_dff_B_P0j1A7UR7_1),.clk(gclk));
	jdff dff_B_OXIUOoLh4_2(.din(n856),.dout(w_dff_B_OXIUOoLh4_2),.clk(gclk));
	jdff dff_B_CmZbFzZh6_2(.din(w_dff_B_OXIUOoLh4_2),.dout(w_dff_B_CmZbFzZh6_2),.clk(gclk));
	jdff dff_B_z1UvYoPe3_2(.din(w_dff_B_CmZbFzZh6_2),.dout(w_dff_B_z1UvYoPe3_2),.clk(gclk));
	jdff dff_B_8zS91aOP5_2(.din(w_dff_B_z1UvYoPe3_2),.dout(w_dff_B_8zS91aOP5_2),.clk(gclk));
	jdff dff_B_HaCrWVrX1_2(.din(w_dff_B_8zS91aOP5_2),.dout(w_dff_B_HaCrWVrX1_2),.clk(gclk));
	jdff dff_B_uon66A4t7_2(.din(w_dff_B_HaCrWVrX1_2),.dout(w_dff_B_uon66A4t7_2),.clk(gclk));
	jdff dff_B_CAVtoGyb2_2(.din(w_dff_B_uon66A4t7_2),.dout(w_dff_B_CAVtoGyb2_2),.clk(gclk));
	jdff dff_B_d38Y6Adh0_2(.din(w_dff_B_CAVtoGyb2_2),.dout(w_dff_B_d38Y6Adh0_2),.clk(gclk));
	jdff dff_B_qRpnyxTx7_2(.din(w_dff_B_d38Y6Adh0_2),.dout(w_dff_B_qRpnyxTx7_2),.clk(gclk));
	jdff dff_B_0KhrJO591_2(.din(w_dff_B_qRpnyxTx7_2),.dout(w_dff_B_0KhrJO591_2),.clk(gclk));
	jdff dff_B_fYYc96mb7_2(.din(w_dff_B_0KhrJO591_2),.dout(w_dff_B_fYYc96mb7_2),.clk(gclk));
	jdff dff_B_UAMoE8dV9_2(.din(w_dff_B_fYYc96mb7_2),.dout(w_dff_B_UAMoE8dV9_2),.clk(gclk));
	jdff dff_B_fKhjjdYX9_2(.din(w_dff_B_UAMoE8dV9_2),.dout(w_dff_B_fKhjjdYX9_2),.clk(gclk));
	jdff dff_B_KrdBSDVd2_2(.din(w_dff_B_fKhjjdYX9_2),.dout(w_dff_B_KrdBSDVd2_2),.clk(gclk));
	jdff dff_B_7zN15ypl5_2(.din(w_dff_B_KrdBSDVd2_2),.dout(w_dff_B_7zN15ypl5_2),.clk(gclk));
	jdff dff_B_QRhlHi2y5_2(.din(w_dff_B_7zN15ypl5_2),.dout(w_dff_B_QRhlHi2y5_2),.clk(gclk));
	jdff dff_B_OZcXcJNC6_2(.din(w_dff_B_QRhlHi2y5_2),.dout(w_dff_B_OZcXcJNC6_2),.clk(gclk));
	jdff dff_B_xsb35Enf5_2(.din(w_dff_B_OZcXcJNC6_2),.dout(w_dff_B_xsb35Enf5_2),.clk(gclk));
	jdff dff_B_iyTO8Kl67_2(.din(w_dff_B_xsb35Enf5_2),.dout(w_dff_B_iyTO8Kl67_2),.clk(gclk));
	jdff dff_B_ManyWFd04_2(.din(w_dff_B_iyTO8Kl67_2),.dout(w_dff_B_ManyWFd04_2),.clk(gclk));
	jdff dff_B_o9S6mCbt4_2(.din(w_dff_B_ManyWFd04_2),.dout(w_dff_B_o9S6mCbt4_2),.clk(gclk));
	jdff dff_B_hMoX1NjO8_2(.din(w_dff_B_o9S6mCbt4_2),.dout(w_dff_B_hMoX1NjO8_2),.clk(gclk));
	jdff dff_B_M6S4EStO2_2(.din(w_dff_B_hMoX1NjO8_2),.dout(w_dff_B_M6S4EStO2_2),.clk(gclk));
	jdff dff_B_hI21th195_2(.din(w_dff_B_M6S4EStO2_2),.dout(w_dff_B_hI21th195_2),.clk(gclk));
	jdff dff_B_NjjlAV5p3_2(.din(w_dff_B_hI21th195_2),.dout(w_dff_B_NjjlAV5p3_2),.clk(gclk));
	jdff dff_B_wliBZn6i9_2(.din(w_dff_B_NjjlAV5p3_2),.dout(w_dff_B_wliBZn6i9_2),.clk(gclk));
	jdff dff_B_Nhrj8v1l1_2(.din(w_dff_B_wliBZn6i9_2),.dout(w_dff_B_Nhrj8v1l1_2),.clk(gclk));
	jdff dff_B_dJ60ay428_2(.din(w_dff_B_Nhrj8v1l1_2),.dout(w_dff_B_dJ60ay428_2),.clk(gclk));
	jdff dff_B_UDL5hThD3_1(.din(n857),.dout(w_dff_B_UDL5hThD3_1),.clk(gclk));
	jdff dff_B_WYR6X4fS7_2(.din(n757),.dout(w_dff_B_WYR6X4fS7_2),.clk(gclk));
	jdff dff_B_1EiUASCF3_2(.din(w_dff_B_WYR6X4fS7_2),.dout(w_dff_B_1EiUASCF3_2),.clk(gclk));
	jdff dff_B_wNJco7zY9_2(.din(w_dff_B_1EiUASCF3_2),.dout(w_dff_B_wNJco7zY9_2),.clk(gclk));
	jdff dff_B_5Cj3yCW42_2(.din(w_dff_B_wNJco7zY9_2),.dout(w_dff_B_5Cj3yCW42_2),.clk(gclk));
	jdff dff_B_hT4hPMCR3_2(.din(w_dff_B_5Cj3yCW42_2),.dout(w_dff_B_hT4hPMCR3_2),.clk(gclk));
	jdff dff_B_vA6MhM9C2_2(.din(w_dff_B_hT4hPMCR3_2),.dout(w_dff_B_vA6MhM9C2_2),.clk(gclk));
	jdff dff_B_FIpGf8mP1_2(.din(w_dff_B_vA6MhM9C2_2),.dout(w_dff_B_FIpGf8mP1_2),.clk(gclk));
	jdff dff_B_MVsv0wPv0_2(.din(w_dff_B_FIpGf8mP1_2),.dout(w_dff_B_MVsv0wPv0_2),.clk(gclk));
	jdff dff_B_mg0O518l1_2(.din(w_dff_B_MVsv0wPv0_2),.dout(w_dff_B_mg0O518l1_2),.clk(gclk));
	jdff dff_B_kMt8oLOT1_2(.din(w_dff_B_mg0O518l1_2),.dout(w_dff_B_kMt8oLOT1_2),.clk(gclk));
	jdff dff_B_wSNUgtch3_2(.din(w_dff_B_kMt8oLOT1_2),.dout(w_dff_B_wSNUgtch3_2),.clk(gclk));
	jdff dff_B_8y9ykXg09_2(.din(w_dff_B_wSNUgtch3_2),.dout(w_dff_B_8y9ykXg09_2),.clk(gclk));
	jdff dff_B_uKuqM9kx5_2(.din(w_dff_B_8y9ykXg09_2),.dout(w_dff_B_uKuqM9kx5_2),.clk(gclk));
	jdff dff_B_XyAt3mok3_2(.din(w_dff_B_uKuqM9kx5_2),.dout(w_dff_B_XyAt3mok3_2),.clk(gclk));
	jdff dff_B_dnhHSFST4_2(.din(w_dff_B_XyAt3mok3_2),.dout(w_dff_B_dnhHSFST4_2),.clk(gclk));
	jdff dff_B_5cpiIYba4_2(.din(w_dff_B_dnhHSFST4_2),.dout(w_dff_B_5cpiIYba4_2),.clk(gclk));
	jdff dff_B_NGJkUk2B5_2(.din(w_dff_B_5cpiIYba4_2),.dout(w_dff_B_NGJkUk2B5_2),.clk(gclk));
	jdff dff_B_DWgZfIhi8_2(.din(w_dff_B_NGJkUk2B5_2),.dout(w_dff_B_DWgZfIhi8_2),.clk(gclk));
	jdff dff_B_qqAHShGX3_2(.din(w_dff_B_DWgZfIhi8_2),.dout(w_dff_B_qqAHShGX3_2),.clk(gclk));
	jdff dff_B_DAyPCTnv6_2(.din(w_dff_B_qqAHShGX3_2),.dout(w_dff_B_DAyPCTnv6_2),.clk(gclk));
	jdff dff_B_FfYx2GC76_2(.din(w_dff_B_DAyPCTnv6_2),.dout(w_dff_B_FfYx2GC76_2),.clk(gclk));
	jdff dff_B_NpaD1rYU5_2(.din(w_dff_B_FfYx2GC76_2),.dout(w_dff_B_NpaD1rYU5_2),.clk(gclk));
	jdff dff_B_9B3sKFAV5_2(.din(w_dff_B_NpaD1rYU5_2),.dout(w_dff_B_9B3sKFAV5_2),.clk(gclk));
	jdff dff_B_dn1IyzkQ2_2(.din(w_dff_B_9B3sKFAV5_2),.dout(w_dff_B_dn1IyzkQ2_2),.clk(gclk));
	jdff dff_B_3UUv34cF6_2(.din(w_dff_B_dn1IyzkQ2_2),.dout(w_dff_B_3UUv34cF6_2),.clk(gclk));
	jdff dff_B_TCeNeTdF2_1(.din(n758),.dout(w_dff_B_TCeNeTdF2_1),.clk(gclk));
	jdff dff_B_QcUiI7CH3_2(.din(n664),.dout(w_dff_B_QcUiI7CH3_2),.clk(gclk));
	jdff dff_B_p0mKxhVA7_2(.din(w_dff_B_QcUiI7CH3_2),.dout(w_dff_B_p0mKxhVA7_2),.clk(gclk));
	jdff dff_B_Gzj7WSl15_2(.din(w_dff_B_p0mKxhVA7_2),.dout(w_dff_B_Gzj7WSl15_2),.clk(gclk));
	jdff dff_B_Sj4h1qfx0_2(.din(w_dff_B_Gzj7WSl15_2),.dout(w_dff_B_Sj4h1qfx0_2),.clk(gclk));
	jdff dff_B_pkvnDbSG7_2(.din(w_dff_B_Sj4h1qfx0_2),.dout(w_dff_B_pkvnDbSG7_2),.clk(gclk));
	jdff dff_B_PenXEBXB5_2(.din(w_dff_B_pkvnDbSG7_2),.dout(w_dff_B_PenXEBXB5_2),.clk(gclk));
	jdff dff_B_GQXZorl61_2(.din(w_dff_B_PenXEBXB5_2),.dout(w_dff_B_GQXZorl61_2),.clk(gclk));
	jdff dff_B_ifYq9zLr9_2(.din(w_dff_B_GQXZorl61_2),.dout(w_dff_B_ifYq9zLr9_2),.clk(gclk));
	jdff dff_B_6w5OLoTf3_2(.din(w_dff_B_ifYq9zLr9_2),.dout(w_dff_B_6w5OLoTf3_2),.clk(gclk));
	jdff dff_B_glB7C4ag2_2(.din(w_dff_B_6w5OLoTf3_2),.dout(w_dff_B_glB7C4ag2_2),.clk(gclk));
	jdff dff_B_NV1kw4X71_2(.din(w_dff_B_glB7C4ag2_2),.dout(w_dff_B_NV1kw4X71_2),.clk(gclk));
	jdff dff_B_Yxm4oLyq7_2(.din(w_dff_B_NV1kw4X71_2),.dout(w_dff_B_Yxm4oLyq7_2),.clk(gclk));
	jdff dff_B_YqoqONaq2_2(.din(w_dff_B_Yxm4oLyq7_2),.dout(w_dff_B_YqoqONaq2_2),.clk(gclk));
	jdff dff_B_HYyigz4y9_2(.din(w_dff_B_YqoqONaq2_2),.dout(w_dff_B_HYyigz4y9_2),.clk(gclk));
	jdff dff_B_WMOHkmnw6_2(.din(w_dff_B_HYyigz4y9_2),.dout(w_dff_B_WMOHkmnw6_2),.clk(gclk));
	jdff dff_B_30Lm1NbZ3_2(.din(w_dff_B_WMOHkmnw6_2),.dout(w_dff_B_30Lm1NbZ3_2),.clk(gclk));
	jdff dff_B_ribJBYlS7_2(.din(w_dff_B_30Lm1NbZ3_2),.dout(w_dff_B_ribJBYlS7_2),.clk(gclk));
	jdff dff_B_z8FhWHer3_2(.din(w_dff_B_ribJBYlS7_2),.dout(w_dff_B_z8FhWHer3_2),.clk(gclk));
	jdff dff_B_67wGB1fs5_2(.din(w_dff_B_z8FhWHer3_2),.dout(w_dff_B_67wGB1fs5_2),.clk(gclk));
	jdff dff_B_oejDmRnQ4_2(.din(w_dff_B_67wGB1fs5_2),.dout(w_dff_B_oejDmRnQ4_2),.clk(gclk));
	jdff dff_B_qWIwacVh8_2(.din(w_dff_B_oejDmRnQ4_2),.dout(w_dff_B_qWIwacVh8_2),.clk(gclk));
	jdff dff_B_jReiZpSs1_2(.din(w_dff_B_qWIwacVh8_2),.dout(w_dff_B_jReiZpSs1_2),.clk(gclk));
	jdff dff_B_YElVKpLK0_1(.din(n665),.dout(w_dff_B_YElVKpLK0_1),.clk(gclk));
	jdff dff_B_xlbZDUBi6_2(.din(n578),.dout(w_dff_B_xlbZDUBi6_2),.clk(gclk));
	jdff dff_B_kLXiJHaK5_2(.din(w_dff_B_xlbZDUBi6_2),.dout(w_dff_B_kLXiJHaK5_2),.clk(gclk));
	jdff dff_B_3MZieGVZ5_2(.din(w_dff_B_kLXiJHaK5_2),.dout(w_dff_B_3MZieGVZ5_2),.clk(gclk));
	jdff dff_B_nvGxiWNk0_2(.din(w_dff_B_3MZieGVZ5_2),.dout(w_dff_B_nvGxiWNk0_2),.clk(gclk));
	jdff dff_B_7SBpEuGF3_2(.din(w_dff_B_nvGxiWNk0_2),.dout(w_dff_B_7SBpEuGF3_2),.clk(gclk));
	jdff dff_B_WoGYCLPa6_2(.din(w_dff_B_7SBpEuGF3_2),.dout(w_dff_B_WoGYCLPa6_2),.clk(gclk));
	jdff dff_B_hfEpRZxv5_2(.din(w_dff_B_WoGYCLPa6_2),.dout(w_dff_B_hfEpRZxv5_2),.clk(gclk));
	jdff dff_B_04pQeXka8_2(.din(w_dff_B_hfEpRZxv5_2),.dout(w_dff_B_04pQeXka8_2),.clk(gclk));
	jdff dff_B_LTIjk67s1_2(.din(w_dff_B_04pQeXka8_2),.dout(w_dff_B_LTIjk67s1_2),.clk(gclk));
	jdff dff_B_ZppctRjs8_2(.din(w_dff_B_LTIjk67s1_2),.dout(w_dff_B_ZppctRjs8_2),.clk(gclk));
	jdff dff_B_xCudkfpS0_2(.din(w_dff_B_ZppctRjs8_2),.dout(w_dff_B_xCudkfpS0_2),.clk(gclk));
	jdff dff_B_FAMxKb3Q8_2(.din(w_dff_B_xCudkfpS0_2),.dout(w_dff_B_FAMxKb3Q8_2),.clk(gclk));
	jdff dff_B_WbTqpJMO0_2(.din(w_dff_B_FAMxKb3Q8_2),.dout(w_dff_B_WbTqpJMO0_2),.clk(gclk));
	jdff dff_B_gZhJ61136_2(.din(w_dff_B_WbTqpJMO0_2),.dout(w_dff_B_gZhJ61136_2),.clk(gclk));
	jdff dff_B_LbLHEl9s2_2(.din(w_dff_B_gZhJ61136_2),.dout(w_dff_B_LbLHEl9s2_2),.clk(gclk));
	jdff dff_B_WplqsmkK7_2(.din(w_dff_B_LbLHEl9s2_2),.dout(w_dff_B_WplqsmkK7_2),.clk(gclk));
	jdff dff_B_cPkiZ6ip5_2(.din(w_dff_B_WplqsmkK7_2),.dout(w_dff_B_cPkiZ6ip5_2),.clk(gclk));
	jdff dff_B_KezsfKsU0_2(.din(w_dff_B_cPkiZ6ip5_2),.dout(w_dff_B_KezsfKsU0_2),.clk(gclk));
	jdff dff_B_UEsYEI8b8_2(.din(w_dff_B_KezsfKsU0_2),.dout(w_dff_B_UEsYEI8b8_2),.clk(gclk));
	jdff dff_B_o79ldpKl3_1(.din(n579),.dout(w_dff_B_o79ldpKl3_1),.clk(gclk));
	jdff dff_B_KLDDFsu83_2(.din(n499),.dout(w_dff_B_KLDDFsu83_2),.clk(gclk));
	jdff dff_B_FpqF9WsI6_2(.din(w_dff_B_KLDDFsu83_2),.dout(w_dff_B_FpqF9WsI6_2),.clk(gclk));
	jdff dff_B_jmIzYgfK4_2(.din(w_dff_B_FpqF9WsI6_2),.dout(w_dff_B_jmIzYgfK4_2),.clk(gclk));
	jdff dff_B_wtpiBXXw0_2(.din(w_dff_B_jmIzYgfK4_2),.dout(w_dff_B_wtpiBXXw0_2),.clk(gclk));
	jdff dff_B_u5QYdera1_2(.din(w_dff_B_wtpiBXXw0_2),.dout(w_dff_B_u5QYdera1_2),.clk(gclk));
	jdff dff_B_FQ9oS25q2_2(.din(w_dff_B_u5QYdera1_2),.dout(w_dff_B_FQ9oS25q2_2),.clk(gclk));
	jdff dff_B_PXb4sKmT7_2(.din(w_dff_B_FQ9oS25q2_2),.dout(w_dff_B_PXb4sKmT7_2),.clk(gclk));
	jdff dff_B_ctwbJgRX1_2(.din(w_dff_B_PXb4sKmT7_2),.dout(w_dff_B_ctwbJgRX1_2),.clk(gclk));
	jdff dff_B_HSQXpIsl9_2(.din(w_dff_B_ctwbJgRX1_2),.dout(w_dff_B_HSQXpIsl9_2),.clk(gclk));
	jdff dff_B_dlzBw1uu6_2(.din(w_dff_B_HSQXpIsl9_2),.dout(w_dff_B_dlzBw1uu6_2),.clk(gclk));
	jdff dff_B_8YaGXYWq7_2(.din(w_dff_B_dlzBw1uu6_2),.dout(w_dff_B_8YaGXYWq7_2),.clk(gclk));
	jdff dff_B_O5Pov7Hy9_2(.din(w_dff_B_8YaGXYWq7_2),.dout(w_dff_B_O5Pov7Hy9_2),.clk(gclk));
	jdff dff_B_K0kHUNdJ1_2(.din(w_dff_B_O5Pov7Hy9_2),.dout(w_dff_B_K0kHUNdJ1_2),.clk(gclk));
	jdff dff_B_T5OkNbqd0_2(.din(w_dff_B_K0kHUNdJ1_2),.dout(w_dff_B_T5OkNbqd0_2),.clk(gclk));
	jdff dff_B_ZlqvOwWy0_2(.din(w_dff_B_T5OkNbqd0_2),.dout(w_dff_B_ZlqvOwWy0_2),.clk(gclk));
	jdff dff_B_2oiaiKTi4_2(.din(w_dff_B_ZlqvOwWy0_2),.dout(w_dff_B_2oiaiKTi4_2),.clk(gclk));
	jdff dff_B_6jsqFIrz7_1(.din(n500),.dout(w_dff_B_6jsqFIrz7_1),.clk(gclk));
	jdff dff_B_u7E9BCYc3_2(.din(n427),.dout(w_dff_B_u7E9BCYc3_2),.clk(gclk));
	jdff dff_B_A3UpByrr6_2(.din(w_dff_B_u7E9BCYc3_2),.dout(w_dff_B_A3UpByrr6_2),.clk(gclk));
	jdff dff_B_ECMFJSbV7_2(.din(w_dff_B_A3UpByrr6_2),.dout(w_dff_B_ECMFJSbV7_2),.clk(gclk));
	jdff dff_B_97I8f5Tv9_2(.din(w_dff_B_ECMFJSbV7_2),.dout(w_dff_B_97I8f5Tv9_2),.clk(gclk));
	jdff dff_B_cbLYQat23_2(.din(w_dff_B_97I8f5Tv9_2),.dout(w_dff_B_cbLYQat23_2),.clk(gclk));
	jdff dff_B_VZbOWOIH8_2(.din(w_dff_B_cbLYQat23_2),.dout(w_dff_B_VZbOWOIH8_2),.clk(gclk));
	jdff dff_B_jCLVR2lx4_2(.din(w_dff_B_VZbOWOIH8_2),.dout(w_dff_B_jCLVR2lx4_2),.clk(gclk));
	jdff dff_B_HRevj4JV1_2(.din(w_dff_B_jCLVR2lx4_2),.dout(w_dff_B_HRevj4JV1_2),.clk(gclk));
	jdff dff_B_B6d6QJdc7_2(.din(w_dff_B_HRevj4JV1_2),.dout(w_dff_B_B6d6QJdc7_2),.clk(gclk));
	jdff dff_B_Q5eu5QZV0_2(.din(w_dff_B_B6d6QJdc7_2),.dout(w_dff_B_Q5eu5QZV0_2),.clk(gclk));
	jdff dff_B_dNJb3Yeb1_2(.din(w_dff_B_Q5eu5QZV0_2),.dout(w_dff_B_dNJb3Yeb1_2),.clk(gclk));
	jdff dff_B_zIQaBel87_2(.din(w_dff_B_dNJb3Yeb1_2),.dout(w_dff_B_zIQaBel87_2),.clk(gclk));
	jdff dff_B_ip1OYZXP2_2(.din(w_dff_B_zIQaBel87_2),.dout(w_dff_B_ip1OYZXP2_2),.clk(gclk));
	jdff dff_B_OxFG7zEq4_1(.din(n428),.dout(w_dff_B_OxFG7zEq4_1),.clk(gclk));
	jdff dff_B_IaqEn6cD0_2(.din(n363),.dout(w_dff_B_IaqEn6cD0_2),.clk(gclk));
	jdff dff_B_95LMWnMg1_2(.din(w_dff_B_IaqEn6cD0_2),.dout(w_dff_B_95LMWnMg1_2),.clk(gclk));
	jdff dff_B_wScDON8r5_2(.din(w_dff_B_95LMWnMg1_2),.dout(w_dff_B_wScDON8r5_2),.clk(gclk));
	jdff dff_B_gUmVQuXm4_2(.din(w_dff_B_wScDON8r5_2),.dout(w_dff_B_gUmVQuXm4_2),.clk(gclk));
	jdff dff_B_rqajqbQu9_2(.din(w_dff_B_gUmVQuXm4_2),.dout(w_dff_B_rqajqbQu9_2),.clk(gclk));
	jdff dff_B_ksSQGzqn5_2(.din(w_dff_B_rqajqbQu9_2),.dout(w_dff_B_ksSQGzqn5_2),.clk(gclk));
	jdff dff_B_r85wganR1_2(.din(w_dff_B_ksSQGzqn5_2),.dout(w_dff_B_r85wganR1_2),.clk(gclk));
	jdff dff_B_TXbdvrH06_2(.din(w_dff_B_r85wganR1_2),.dout(w_dff_B_TXbdvrH06_2),.clk(gclk));
	jdff dff_B_QPOFtPMW1_2(.din(w_dff_B_TXbdvrH06_2),.dout(w_dff_B_QPOFtPMW1_2),.clk(gclk));
	jdff dff_B_VkUFP3RP6_2(.din(w_dff_B_QPOFtPMW1_2),.dout(w_dff_B_VkUFP3RP6_2),.clk(gclk));
	jdff dff_B_io9CbdDf0_2(.din(n385),.dout(w_dff_B_io9CbdDf0_2),.clk(gclk));
	jdff dff_B_FqnL9AwD9_1(.din(n364),.dout(w_dff_B_FqnL9AwD9_1),.clk(gclk));
	jdff dff_B_DYZfqvEo8_2(.din(n305),.dout(w_dff_B_DYZfqvEo8_2),.clk(gclk));
	jdff dff_B_HGKg3pE81_2(.din(w_dff_B_DYZfqvEo8_2),.dout(w_dff_B_HGKg3pE81_2),.clk(gclk));
	jdff dff_B_X03eZoHQ5_2(.din(w_dff_B_HGKg3pE81_2),.dout(w_dff_B_X03eZoHQ5_2),.clk(gclk));
	jdff dff_B_UPMDiGPW9_2(.din(w_dff_B_X03eZoHQ5_2),.dout(w_dff_B_UPMDiGPW9_2),.clk(gclk));
	jdff dff_B_cxJ5nufr4_2(.din(w_dff_B_UPMDiGPW9_2),.dout(w_dff_B_cxJ5nufr4_2),.clk(gclk));
	jdff dff_B_VSZnugCs8_2(.din(w_dff_B_cxJ5nufr4_2),.dout(w_dff_B_VSZnugCs8_2),.clk(gclk));
	jdff dff_B_qiqaGBdF2_2(.din(w_dff_B_VSZnugCs8_2),.dout(w_dff_B_qiqaGBdF2_2),.clk(gclk));
	jdff dff_B_GQJav8ev3_2(.din(n321),.dout(w_dff_B_GQJav8ev3_2),.clk(gclk));
	jdff dff_B_Us5gRVrN8_1(.din(n306),.dout(w_dff_B_Us5gRVrN8_1),.clk(gclk));
	jdff dff_B_reSi97mk6_2(.din(n254),.dout(w_dff_B_reSi97mk6_2),.clk(gclk));
	jdff dff_B_plJwiYGs8_2(.din(w_dff_B_reSi97mk6_2),.dout(w_dff_B_plJwiYGs8_2),.clk(gclk));
	jdff dff_B_kqNS9IRA6_2(.din(w_dff_B_plJwiYGs8_2),.dout(w_dff_B_kqNS9IRA6_2),.clk(gclk));
	jdff dff_B_NxmFnLMh2_2(.din(w_dff_B_kqNS9IRA6_2),.dout(w_dff_B_NxmFnLMh2_2),.clk(gclk));
	jdff dff_B_ld0GMe2J5_1(.din(n256),.dout(w_dff_B_ld0GMe2J5_1),.clk(gclk));
	jdff dff_A_ihGef0np8_1(.dout(w_n210_0[1]),.din(w_dff_A_ihGef0np8_1),.clk(gclk));
	jdff dff_A_UFdfwBAu8_2(.dout(w_n210_0[2]),.din(w_dff_A_UFdfwBAu8_2),.clk(gclk));
	jdff dff_A_ME7jCby71_2(.dout(w_dff_A_UFdfwBAu8_2),.din(w_dff_A_ME7jCby71_2),.clk(gclk));
	jdff dff_B_a33fP2nu5_2(.din(n1496),.dout(w_dff_B_a33fP2nu5_2),.clk(gclk));
	jdff dff_B_ldfrfag78_1(.din(n1494),.dout(w_dff_B_ldfrfag78_1),.clk(gclk));
	jdff dff_B_YopbOVgc0_2(.din(n1421),.dout(w_dff_B_YopbOVgc0_2),.clk(gclk));
	jdff dff_B_eWIuPVRh6_2(.din(w_dff_B_YopbOVgc0_2),.dout(w_dff_B_eWIuPVRh6_2),.clk(gclk));
	jdff dff_B_GRDWU3Zx6_2(.din(w_dff_B_eWIuPVRh6_2),.dout(w_dff_B_GRDWU3Zx6_2),.clk(gclk));
	jdff dff_B_0fyB5x247_2(.din(w_dff_B_GRDWU3Zx6_2),.dout(w_dff_B_0fyB5x247_2),.clk(gclk));
	jdff dff_B_VLvMbGr95_2(.din(w_dff_B_0fyB5x247_2),.dout(w_dff_B_VLvMbGr95_2),.clk(gclk));
	jdff dff_B_kDS3O4KO7_2(.din(w_dff_B_VLvMbGr95_2),.dout(w_dff_B_kDS3O4KO7_2),.clk(gclk));
	jdff dff_B_06gyuQDf8_2(.din(w_dff_B_kDS3O4KO7_2),.dout(w_dff_B_06gyuQDf8_2),.clk(gclk));
	jdff dff_B_31MFiyW06_2(.din(w_dff_B_06gyuQDf8_2),.dout(w_dff_B_31MFiyW06_2),.clk(gclk));
	jdff dff_B_v2kQEH1V3_2(.din(w_dff_B_31MFiyW06_2),.dout(w_dff_B_v2kQEH1V3_2),.clk(gclk));
	jdff dff_B_hxE3nZQB8_2(.din(w_dff_B_v2kQEH1V3_2),.dout(w_dff_B_hxE3nZQB8_2),.clk(gclk));
	jdff dff_B_HBifSMOO0_2(.din(w_dff_B_hxE3nZQB8_2),.dout(w_dff_B_HBifSMOO0_2),.clk(gclk));
	jdff dff_B_4C4RFaPW2_2(.din(w_dff_B_HBifSMOO0_2),.dout(w_dff_B_4C4RFaPW2_2),.clk(gclk));
	jdff dff_B_wLYE6GuJ5_2(.din(w_dff_B_4C4RFaPW2_2),.dout(w_dff_B_wLYE6GuJ5_2),.clk(gclk));
	jdff dff_B_9m9kf7zg4_2(.din(w_dff_B_wLYE6GuJ5_2),.dout(w_dff_B_9m9kf7zg4_2),.clk(gclk));
	jdff dff_B_znXQe2J80_2(.din(w_dff_B_9m9kf7zg4_2),.dout(w_dff_B_znXQe2J80_2),.clk(gclk));
	jdff dff_B_teBCpntl9_2(.din(w_dff_B_znXQe2J80_2),.dout(w_dff_B_teBCpntl9_2),.clk(gclk));
	jdff dff_B_wicxiOmA5_2(.din(w_dff_B_teBCpntl9_2),.dout(w_dff_B_wicxiOmA5_2),.clk(gclk));
	jdff dff_B_Zy60lVAV2_2(.din(w_dff_B_wicxiOmA5_2),.dout(w_dff_B_Zy60lVAV2_2),.clk(gclk));
	jdff dff_B_lE6DP6rJ8_2(.din(w_dff_B_Zy60lVAV2_2),.dout(w_dff_B_lE6DP6rJ8_2),.clk(gclk));
	jdff dff_B_aKSAEdNP7_2(.din(w_dff_B_lE6DP6rJ8_2),.dout(w_dff_B_aKSAEdNP7_2),.clk(gclk));
	jdff dff_B_fSk7J3782_2(.din(w_dff_B_aKSAEdNP7_2),.dout(w_dff_B_fSk7J3782_2),.clk(gclk));
	jdff dff_B_pfO65SxL1_2(.din(w_dff_B_fSk7J3782_2),.dout(w_dff_B_pfO65SxL1_2),.clk(gclk));
	jdff dff_B_8b1SmzKf6_2(.din(w_dff_B_pfO65SxL1_2),.dout(w_dff_B_8b1SmzKf6_2),.clk(gclk));
	jdff dff_B_mJ85caAD8_2(.din(w_dff_B_8b1SmzKf6_2),.dout(w_dff_B_mJ85caAD8_2),.clk(gclk));
	jdff dff_B_miI1PorH1_2(.din(w_dff_B_mJ85caAD8_2),.dout(w_dff_B_miI1PorH1_2),.clk(gclk));
	jdff dff_B_HD7tQvOF1_2(.din(w_dff_B_miI1PorH1_2),.dout(w_dff_B_HD7tQvOF1_2),.clk(gclk));
	jdff dff_B_KbYHEZsq2_2(.din(w_dff_B_HD7tQvOF1_2),.dout(w_dff_B_KbYHEZsq2_2),.clk(gclk));
	jdff dff_B_WUSUN2y83_2(.din(w_dff_B_KbYHEZsq2_2),.dout(w_dff_B_WUSUN2y83_2),.clk(gclk));
	jdff dff_B_zM5xh3Ux3_2(.din(w_dff_B_WUSUN2y83_2),.dout(w_dff_B_zM5xh3Ux3_2),.clk(gclk));
	jdff dff_B_gYXFpMN14_2(.din(w_dff_B_zM5xh3Ux3_2),.dout(w_dff_B_gYXFpMN14_2),.clk(gclk));
	jdff dff_B_2vbDUsx77_2(.din(w_dff_B_gYXFpMN14_2),.dout(w_dff_B_2vbDUsx77_2),.clk(gclk));
	jdff dff_B_yGgFNGF35_2(.din(w_dff_B_2vbDUsx77_2),.dout(w_dff_B_yGgFNGF35_2),.clk(gclk));
	jdff dff_B_Ae60r8WL9_2(.din(w_dff_B_yGgFNGF35_2),.dout(w_dff_B_Ae60r8WL9_2),.clk(gclk));
	jdff dff_B_xHv7a9Jw2_2(.din(w_dff_B_Ae60r8WL9_2),.dout(w_dff_B_xHv7a9Jw2_2),.clk(gclk));
	jdff dff_B_NtRzrdJq3_2(.din(w_dff_B_xHv7a9Jw2_2),.dout(w_dff_B_NtRzrdJq3_2),.clk(gclk));
	jdff dff_B_8vEXte5I0_2(.din(w_dff_B_NtRzrdJq3_2),.dout(w_dff_B_8vEXte5I0_2),.clk(gclk));
	jdff dff_B_P19jcpSz5_2(.din(w_dff_B_8vEXte5I0_2),.dout(w_dff_B_P19jcpSz5_2),.clk(gclk));
	jdff dff_B_6udUZmPU9_2(.din(w_dff_B_P19jcpSz5_2),.dout(w_dff_B_6udUZmPU9_2),.clk(gclk));
	jdff dff_B_D3CIDLky0_2(.din(w_dff_B_6udUZmPU9_2),.dout(w_dff_B_D3CIDLky0_2),.clk(gclk));
	jdff dff_B_xByME6L32_2(.din(w_dff_B_D3CIDLky0_2),.dout(w_dff_B_xByME6L32_2),.clk(gclk));
	jdff dff_B_VPP5cuBQ8_2(.din(w_dff_B_xByME6L32_2),.dout(w_dff_B_VPP5cuBQ8_2),.clk(gclk));
	jdff dff_B_gUpcipTp4_2(.din(w_dff_B_VPP5cuBQ8_2),.dout(w_dff_B_gUpcipTp4_2),.clk(gclk));
	jdff dff_B_vlb96aLX1_2(.din(w_dff_B_gUpcipTp4_2),.dout(w_dff_B_vlb96aLX1_2),.clk(gclk));
	jdff dff_B_FsrhkoL98_2(.din(w_dff_B_vlb96aLX1_2),.dout(w_dff_B_FsrhkoL98_2),.clk(gclk));
	jdff dff_B_hFQBophy3_2(.din(w_dff_B_FsrhkoL98_2),.dout(w_dff_B_hFQBophy3_2),.clk(gclk));
	jdff dff_B_Vzsvtm4e3_2(.din(w_dff_B_hFQBophy3_2),.dout(w_dff_B_Vzsvtm4e3_2),.clk(gclk));
	jdff dff_B_gMOD04LK8_1(.din(n1422),.dout(w_dff_B_gMOD04LK8_1),.clk(gclk));
	jdff dff_B_JPKKkgyZ2_2(.din(n1343),.dout(w_dff_B_JPKKkgyZ2_2),.clk(gclk));
	jdff dff_B_XI1hN6LU8_2(.din(w_dff_B_JPKKkgyZ2_2),.dout(w_dff_B_XI1hN6LU8_2),.clk(gclk));
	jdff dff_B_OEp2csFP1_2(.din(w_dff_B_XI1hN6LU8_2),.dout(w_dff_B_OEp2csFP1_2),.clk(gclk));
	jdff dff_B_zSLDlSjR2_2(.din(w_dff_B_OEp2csFP1_2),.dout(w_dff_B_zSLDlSjR2_2),.clk(gclk));
	jdff dff_B_qroJzE191_2(.din(w_dff_B_zSLDlSjR2_2),.dout(w_dff_B_qroJzE191_2),.clk(gclk));
	jdff dff_B_HPeq6HI29_2(.din(w_dff_B_qroJzE191_2),.dout(w_dff_B_HPeq6HI29_2),.clk(gclk));
	jdff dff_B_IHE6y6hl2_2(.din(w_dff_B_HPeq6HI29_2),.dout(w_dff_B_IHE6y6hl2_2),.clk(gclk));
	jdff dff_B_TL7fwjhG1_2(.din(w_dff_B_IHE6y6hl2_2),.dout(w_dff_B_TL7fwjhG1_2),.clk(gclk));
	jdff dff_B_gnjlbvzi4_2(.din(w_dff_B_TL7fwjhG1_2),.dout(w_dff_B_gnjlbvzi4_2),.clk(gclk));
	jdff dff_B_wWluNzAv1_2(.din(w_dff_B_gnjlbvzi4_2),.dout(w_dff_B_wWluNzAv1_2),.clk(gclk));
	jdff dff_B_G8Ao3u3H9_2(.din(w_dff_B_wWluNzAv1_2),.dout(w_dff_B_G8Ao3u3H9_2),.clk(gclk));
	jdff dff_B_fUqjQJOO1_2(.din(w_dff_B_G8Ao3u3H9_2),.dout(w_dff_B_fUqjQJOO1_2),.clk(gclk));
	jdff dff_B_hbdkR3oi6_2(.din(w_dff_B_fUqjQJOO1_2),.dout(w_dff_B_hbdkR3oi6_2),.clk(gclk));
	jdff dff_B_iisJzLOF6_2(.din(w_dff_B_hbdkR3oi6_2),.dout(w_dff_B_iisJzLOF6_2),.clk(gclk));
	jdff dff_B_rlV2Adwh7_2(.din(w_dff_B_iisJzLOF6_2),.dout(w_dff_B_rlV2Adwh7_2),.clk(gclk));
	jdff dff_B_voFJmxMS9_2(.din(w_dff_B_rlV2Adwh7_2),.dout(w_dff_B_voFJmxMS9_2),.clk(gclk));
	jdff dff_B_QBGxZDqj4_2(.din(w_dff_B_voFJmxMS9_2),.dout(w_dff_B_QBGxZDqj4_2),.clk(gclk));
	jdff dff_B_GVEgjdkh0_2(.din(w_dff_B_QBGxZDqj4_2),.dout(w_dff_B_GVEgjdkh0_2),.clk(gclk));
	jdff dff_B_fiMewi637_2(.din(w_dff_B_GVEgjdkh0_2),.dout(w_dff_B_fiMewi637_2),.clk(gclk));
	jdff dff_B_TnyTLXOj3_2(.din(w_dff_B_fiMewi637_2),.dout(w_dff_B_TnyTLXOj3_2),.clk(gclk));
	jdff dff_B_tIBRf3oc1_2(.din(w_dff_B_TnyTLXOj3_2),.dout(w_dff_B_tIBRf3oc1_2),.clk(gclk));
	jdff dff_B_jeO4sf1y5_2(.din(w_dff_B_tIBRf3oc1_2),.dout(w_dff_B_jeO4sf1y5_2),.clk(gclk));
	jdff dff_B_9aiGenyJ0_2(.din(w_dff_B_jeO4sf1y5_2),.dout(w_dff_B_9aiGenyJ0_2),.clk(gclk));
	jdff dff_B_KgMIuiRv3_2(.din(w_dff_B_9aiGenyJ0_2),.dout(w_dff_B_KgMIuiRv3_2),.clk(gclk));
	jdff dff_B_maD6bYUp0_2(.din(w_dff_B_KgMIuiRv3_2),.dout(w_dff_B_maD6bYUp0_2),.clk(gclk));
	jdff dff_B_E3hVxtbw5_2(.din(w_dff_B_maD6bYUp0_2),.dout(w_dff_B_E3hVxtbw5_2),.clk(gclk));
	jdff dff_B_jnNrYOPt7_2(.din(w_dff_B_E3hVxtbw5_2),.dout(w_dff_B_jnNrYOPt7_2),.clk(gclk));
	jdff dff_B_mJSkHJbU7_2(.din(w_dff_B_jnNrYOPt7_2),.dout(w_dff_B_mJSkHJbU7_2),.clk(gclk));
	jdff dff_B_m3eRQ6ht4_2(.din(w_dff_B_mJSkHJbU7_2),.dout(w_dff_B_m3eRQ6ht4_2),.clk(gclk));
	jdff dff_B_NkWAB6qo9_2(.din(w_dff_B_m3eRQ6ht4_2),.dout(w_dff_B_NkWAB6qo9_2),.clk(gclk));
	jdff dff_B_6iqaITqX3_2(.din(w_dff_B_NkWAB6qo9_2),.dout(w_dff_B_6iqaITqX3_2),.clk(gclk));
	jdff dff_B_Q6cPTMuz3_2(.din(w_dff_B_6iqaITqX3_2),.dout(w_dff_B_Q6cPTMuz3_2),.clk(gclk));
	jdff dff_B_Q72KRGlz9_2(.din(w_dff_B_Q6cPTMuz3_2),.dout(w_dff_B_Q72KRGlz9_2),.clk(gclk));
	jdff dff_B_j9AdApCh5_2(.din(w_dff_B_Q72KRGlz9_2),.dout(w_dff_B_j9AdApCh5_2),.clk(gclk));
	jdff dff_B_GEDCO0BG4_2(.din(w_dff_B_j9AdApCh5_2),.dout(w_dff_B_GEDCO0BG4_2),.clk(gclk));
	jdff dff_B_MN5QEbox8_2(.din(w_dff_B_GEDCO0BG4_2),.dout(w_dff_B_MN5QEbox8_2),.clk(gclk));
	jdff dff_B_faP0WOb70_2(.din(w_dff_B_MN5QEbox8_2),.dout(w_dff_B_faP0WOb70_2),.clk(gclk));
	jdff dff_B_iNdENpZB7_2(.din(w_dff_B_faP0WOb70_2),.dout(w_dff_B_iNdENpZB7_2),.clk(gclk));
	jdff dff_B_TcqLODSQ1_2(.din(w_dff_B_iNdENpZB7_2),.dout(w_dff_B_TcqLODSQ1_2),.clk(gclk));
	jdff dff_B_uRxpRYjz2_2(.din(w_dff_B_TcqLODSQ1_2),.dout(w_dff_B_uRxpRYjz2_2),.clk(gclk));
	jdff dff_B_48lD1CKl9_2(.din(w_dff_B_uRxpRYjz2_2),.dout(w_dff_B_48lD1CKl9_2),.clk(gclk));
	jdff dff_B_RZ68iGV39_1(.din(n1344),.dout(w_dff_B_RZ68iGV39_1),.clk(gclk));
	jdff dff_B_KFJiuq5N9_2(.din(n1258),.dout(w_dff_B_KFJiuq5N9_2),.clk(gclk));
	jdff dff_B_0YKe3tCR5_2(.din(w_dff_B_KFJiuq5N9_2),.dout(w_dff_B_0YKe3tCR5_2),.clk(gclk));
	jdff dff_B_3rbb7qLk6_2(.din(w_dff_B_0YKe3tCR5_2),.dout(w_dff_B_3rbb7qLk6_2),.clk(gclk));
	jdff dff_B_sJUeJWGk0_2(.din(w_dff_B_3rbb7qLk6_2),.dout(w_dff_B_sJUeJWGk0_2),.clk(gclk));
	jdff dff_B_75jZM8Ny8_2(.din(w_dff_B_sJUeJWGk0_2),.dout(w_dff_B_75jZM8Ny8_2),.clk(gclk));
	jdff dff_B_djLFzpT95_2(.din(w_dff_B_75jZM8Ny8_2),.dout(w_dff_B_djLFzpT95_2),.clk(gclk));
	jdff dff_B_reFHK3Yc4_2(.din(w_dff_B_djLFzpT95_2),.dout(w_dff_B_reFHK3Yc4_2),.clk(gclk));
	jdff dff_B_BHvNkurK6_2(.din(w_dff_B_reFHK3Yc4_2),.dout(w_dff_B_BHvNkurK6_2),.clk(gclk));
	jdff dff_B_kAeCw6A77_2(.din(w_dff_B_BHvNkurK6_2),.dout(w_dff_B_kAeCw6A77_2),.clk(gclk));
	jdff dff_B_pqociOfC7_2(.din(w_dff_B_kAeCw6A77_2),.dout(w_dff_B_pqociOfC7_2),.clk(gclk));
	jdff dff_B_89rbMWGo2_2(.din(w_dff_B_pqociOfC7_2),.dout(w_dff_B_89rbMWGo2_2),.clk(gclk));
	jdff dff_B_g7c2nQDA0_2(.din(w_dff_B_89rbMWGo2_2),.dout(w_dff_B_g7c2nQDA0_2),.clk(gclk));
	jdff dff_B_rG3yH1Hq7_2(.din(w_dff_B_g7c2nQDA0_2),.dout(w_dff_B_rG3yH1Hq7_2),.clk(gclk));
	jdff dff_B_liKv9Xwc3_2(.din(w_dff_B_rG3yH1Hq7_2),.dout(w_dff_B_liKv9Xwc3_2),.clk(gclk));
	jdff dff_B_rY5h51Sy4_2(.din(w_dff_B_liKv9Xwc3_2),.dout(w_dff_B_rY5h51Sy4_2),.clk(gclk));
	jdff dff_B_L5JkQPZ33_2(.din(w_dff_B_rY5h51Sy4_2),.dout(w_dff_B_L5JkQPZ33_2),.clk(gclk));
	jdff dff_B_yU6BNIox6_2(.din(w_dff_B_L5JkQPZ33_2),.dout(w_dff_B_yU6BNIox6_2),.clk(gclk));
	jdff dff_B_ko1uQX8q9_2(.din(w_dff_B_yU6BNIox6_2),.dout(w_dff_B_ko1uQX8q9_2),.clk(gclk));
	jdff dff_B_94YFYyOb3_2(.din(w_dff_B_ko1uQX8q9_2),.dout(w_dff_B_94YFYyOb3_2),.clk(gclk));
	jdff dff_B_cLWsJTfx5_2(.din(w_dff_B_94YFYyOb3_2),.dout(w_dff_B_cLWsJTfx5_2),.clk(gclk));
	jdff dff_B_Nc7jlJOn1_2(.din(w_dff_B_cLWsJTfx5_2),.dout(w_dff_B_Nc7jlJOn1_2),.clk(gclk));
	jdff dff_B_bpA98IQ31_2(.din(w_dff_B_Nc7jlJOn1_2),.dout(w_dff_B_bpA98IQ31_2),.clk(gclk));
	jdff dff_B_crlLbWCT1_2(.din(w_dff_B_bpA98IQ31_2),.dout(w_dff_B_crlLbWCT1_2),.clk(gclk));
	jdff dff_B_FbxaMjPy3_2(.din(w_dff_B_crlLbWCT1_2),.dout(w_dff_B_FbxaMjPy3_2),.clk(gclk));
	jdff dff_B_2fl6Fxwo8_2(.din(w_dff_B_FbxaMjPy3_2),.dout(w_dff_B_2fl6Fxwo8_2),.clk(gclk));
	jdff dff_B_TPbtqJO76_2(.din(w_dff_B_2fl6Fxwo8_2),.dout(w_dff_B_TPbtqJO76_2),.clk(gclk));
	jdff dff_B_V1Yo2WOt2_2(.din(w_dff_B_TPbtqJO76_2),.dout(w_dff_B_V1Yo2WOt2_2),.clk(gclk));
	jdff dff_B_6PHdLnga7_2(.din(w_dff_B_V1Yo2WOt2_2),.dout(w_dff_B_6PHdLnga7_2),.clk(gclk));
	jdff dff_B_cnaKGKw74_2(.din(w_dff_B_6PHdLnga7_2),.dout(w_dff_B_cnaKGKw74_2),.clk(gclk));
	jdff dff_B_236yhGDc5_2(.din(w_dff_B_cnaKGKw74_2),.dout(w_dff_B_236yhGDc5_2),.clk(gclk));
	jdff dff_B_git90gTn4_2(.din(w_dff_B_236yhGDc5_2),.dout(w_dff_B_git90gTn4_2),.clk(gclk));
	jdff dff_B_YFZr2Nw31_2(.din(w_dff_B_git90gTn4_2),.dout(w_dff_B_YFZr2Nw31_2),.clk(gclk));
	jdff dff_B_npnLzxhn2_2(.din(w_dff_B_YFZr2Nw31_2),.dout(w_dff_B_npnLzxhn2_2),.clk(gclk));
	jdff dff_B_AAQ7mzk81_2(.din(w_dff_B_npnLzxhn2_2),.dout(w_dff_B_AAQ7mzk81_2),.clk(gclk));
	jdff dff_B_KMmU36vm5_2(.din(w_dff_B_AAQ7mzk81_2),.dout(w_dff_B_KMmU36vm5_2),.clk(gclk));
	jdff dff_B_6zEDXQG32_2(.din(w_dff_B_KMmU36vm5_2),.dout(w_dff_B_6zEDXQG32_2),.clk(gclk));
	jdff dff_B_ftoLNtMu0_2(.din(w_dff_B_6zEDXQG32_2),.dout(w_dff_B_ftoLNtMu0_2),.clk(gclk));
	jdff dff_B_WDf10k9W8_2(.din(w_dff_B_ftoLNtMu0_2),.dout(w_dff_B_WDf10k9W8_2),.clk(gclk));
	jdff dff_B_ZI9ttziG9_1(.din(n1259),.dout(w_dff_B_ZI9ttziG9_1),.clk(gclk));
	jdff dff_B_5H3rShpr7_2(.din(n1168),.dout(w_dff_B_5H3rShpr7_2),.clk(gclk));
	jdff dff_B_8VVajlqj1_2(.din(w_dff_B_5H3rShpr7_2),.dout(w_dff_B_8VVajlqj1_2),.clk(gclk));
	jdff dff_B_bAVnja4l2_2(.din(w_dff_B_8VVajlqj1_2),.dout(w_dff_B_bAVnja4l2_2),.clk(gclk));
	jdff dff_B_Uc6xRWYa9_2(.din(w_dff_B_bAVnja4l2_2),.dout(w_dff_B_Uc6xRWYa9_2),.clk(gclk));
	jdff dff_B_LRvRgw2j0_2(.din(w_dff_B_Uc6xRWYa9_2),.dout(w_dff_B_LRvRgw2j0_2),.clk(gclk));
	jdff dff_B_xcJPdG8w2_2(.din(w_dff_B_LRvRgw2j0_2),.dout(w_dff_B_xcJPdG8w2_2),.clk(gclk));
	jdff dff_B_1bvD3nxm7_2(.din(w_dff_B_xcJPdG8w2_2),.dout(w_dff_B_1bvD3nxm7_2),.clk(gclk));
	jdff dff_B_ASBkdjsz7_2(.din(w_dff_B_1bvD3nxm7_2),.dout(w_dff_B_ASBkdjsz7_2),.clk(gclk));
	jdff dff_B_8I2C815e1_2(.din(w_dff_B_ASBkdjsz7_2),.dout(w_dff_B_8I2C815e1_2),.clk(gclk));
	jdff dff_B_z1QCF9jJ6_2(.din(w_dff_B_8I2C815e1_2),.dout(w_dff_B_z1QCF9jJ6_2),.clk(gclk));
	jdff dff_B_nxCQ0w4O1_2(.din(w_dff_B_z1QCF9jJ6_2),.dout(w_dff_B_nxCQ0w4O1_2),.clk(gclk));
	jdff dff_B_JDDM5JJs7_2(.din(w_dff_B_nxCQ0w4O1_2),.dout(w_dff_B_JDDM5JJs7_2),.clk(gclk));
	jdff dff_B_jGGTOKtQ5_2(.din(w_dff_B_JDDM5JJs7_2),.dout(w_dff_B_jGGTOKtQ5_2),.clk(gclk));
	jdff dff_B_tsV8RmVd3_2(.din(w_dff_B_jGGTOKtQ5_2),.dout(w_dff_B_tsV8RmVd3_2),.clk(gclk));
	jdff dff_B_lQjfcswZ6_2(.din(w_dff_B_tsV8RmVd3_2),.dout(w_dff_B_lQjfcswZ6_2),.clk(gclk));
	jdff dff_B_cO59nhhm8_2(.din(w_dff_B_lQjfcswZ6_2),.dout(w_dff_B_cO59nhhm8_2),.clk(gclk));
	jdff dff_B_pyoOHU246_2(.din(w_dff_B_cO59nhhm8_2),.dout(w_dff_B_pyoOHU246_2),.clk(gclk));
	jdff dff_B_mJlORRbv0_2(.din(w_dff_B_pyoOHU246_2),.dout(w_dff_B_mJlORRbv0_2),.clk(gclk));
	jdff dff_B_SUStyfXp9_2(.din(w_dff_B_mJlORRbv0_2),.dout(w_dff_B_SUStyfXp9_2),.clk(gclk));
	jdff dff_B_bHfjIWcU9_2(.din(w_dff_B_SUStyfXp9_2),.dout(w_dff_B_bHfjIWcU9_2),.clk(gclk));
	jdff dff_B_3NuufQ5J1_2(.din(w_dff_B_bHfjIWcU9_2),.dout(w_dff_B_3NuufQ5J1_2),.clk(gclk));
	jdff dff_B_u2X4psDd6_2(.din(w_dff_B_3NuufQ5J1_2),.dout(w_dff_B_u2X4psDd6_2),.clk(gclk));
	jdff dff_B_2pH2f6uW9_2(.din(w_dff_B_u2X4psDd6_2),.dout(w_dff_B_2pH2f6uW9_2),.clk(gclk));
	jdff dff_B_lwC2gSPs2_2(.din(w_dff_B_2pH2f6uW9_2),.dout(w_dff_B_lwC2gSPs2_2),.clk(gclk));
	jdff dff_B_fSBAsAr70_2(.din(w_dff_B_lwC2gSPs2_2),.dout(w_dff_B_fSBAsAr70_2),.clk(gclk));
	jdff dff_B_3CeHHTiH2_2(.din(w_dff_B_fSBAsAr70_2),.dout(w_dff_B_3CeHHTiH2_2),.clk(gclk));
	jdff dff_B_twBWysc17_2(.din(w_dff_B_3CeHHTiH2_2),.dout(w_dff_B_twBWysc17_2),.clk(gclk));
	jdff dff_B_iZWSx8Ib7_2(.din(w_dff_B_twBWysc17_2),.dout(w_dff_B_iZWSx8Ib7_2),.clk(gclk));
	jdff dff_B_xu8kWeZT1_2(.din(w_dff_B_iZWSx8Ib7_2),.dout(w_dff_B_xu8kWeZT1_2),.clk(gclk));
	jdff dff_B_YoSLBF7D6_2(.din(w_dff_B_xu8kWeZT1_2),.dout(w_dff_B_YoSLBF7D6_2),.clk(gclk));
	jdff dff_B_4X8NU8Ze6_2(.din(w_dff_B_YoSLBF7D6_2),.dout(w_dff_B_4X8NU8Ze6_2),.clk(gclk));
	jdff dff_B_MrRiON2f2_2(.din(w_dff_B_4X8NU8Ze6_2),.dout(w_dff_B_MrRiON2f2_2),.clk(gclk));
	jdff dff_B_M13MTssq1_2(.din(w_dff_B_MrRiON2f2_2),.dout(w_dff_B_M13MTssq1_2),.clk(gclk));
	jdff dff_B_iZoOIOJk2_2(.din(w_dff_B_M13MTssq1_2),.dout(w_dff_B_iZoOIOJk2_2),.clk(gclk));
	jdff dff_B_f2fXMfxO2_2(.din(w_dff_B_iZoOIOJk2_2),.dout(w_dff_B_f2fXMfxO2_2),.clk(gclk));
	jdff dff_B_h96iplJp8_1(.din(n1169),.dout(w_dff_B_h96iplJp8_1),.clk(gclk));
	jdff dff_B_qf1KbyvZ9_2(.din(n1064),.dout(w_dff_B_qf1KbyvZ9_2),.clk(gclk));
	jdff dff_B_GiRXq2pD7_2(.din(w_dff_B_qf1KbyvZ9_2),.dout(w_dff_B_GiRXq2pD7_2),.clk(gclk));
	jdff dff_B_sFXmxg8H3_2(.din(w_dff_B_GiRXq2pD7_2),.dout(w_dff_B_sFXmxg8H3_2),.clk(gclk));
	jdff dff_B_0yoVnBMw0_2(.din(w_dff_B_sFXmxg8H3_2),.dout(w_dff_B_0yoVnBMw0_2),.clk(gclk));
	jdff dff_B_RwYS4Orm3_2(.din(w_dff_B_0yoVnBMw0_2),.dout(w_dff_B_RwYS4Orm3_2),.clk(gclk));
	jdff dff_B_oIzowEBO4_2(.din(w_dff_B_RwYS4Orm3_2),.dout(w_dff_B_oIzowEBO4_2),.clk(gclk));
	jdff dff_B_1m30Jtb47_2(.din(w_dff_B_oIzowEBO4_2),.dout(w_dff_B_1m30Jtb47_2),.clk(gclk));
	jdff dff_B_G3DM9bid2_2(.din(w_dff_B_1m30Jtb47_2),.dout(w_dff_B_G3DM9bid2_2),.clk(gclk));
	jdff dff_B_ko52E0RT1_2(.din(w_dff_B_G3DM9bid2_2),.dout(w_dff_B_ko52E0RT1_2),.clk(gclk));
	jdff dff_B_16dFWnR53_2(.din(w_dff_B_ko52E0RT1_2),.dout(w_dff_B_16dFWnR53_2),.clk(gclk));
	jdff dff_B_wSzjwccF5_2(.din(w_dff_B_16dFWnR53_2),.dout(w_dff_B_wSzjwccF5_2),.clk(gclk));
	jdff dff_B_YvuMUbEI9_2(.din(w_dff_B_wSzjwccF5_2),.dout(w_dff_B_YvuMUbEI9_2),.clk(gclk));
	jdff dff_B_JFGP2rfe0_2(.din(w_dff_B_YvuMUbEI9_2),.dout(w_dff_B_JFGP2rfe0_2),.clk(gclk));
	jdff dff_B_17Hop5s74_2(.din(w_dff_B_JFGP2rfe0_2),.dout(w_dff_B_17Hop5s74_2),.clk(gclk));
	jdff dff_B_6ZYgppYs0_2(.din(w_dff_B_17Hop5s74_2),.dout(w_dff_B_6ZYgppYs0_2),.clk(gclk));
	jdff dff_B_w5Qj2VkR7_2(.din(w_dff_B_6ZYgppYs0_2),.dout(w_dff_B_w5Qj2VkR7_2),.clk(gclk));
	jdff dff_B_p80WPCGv9_2(.din(w_dff_B_w5Qj2VkR7_2),.dout(w_dff_B_p80WPCGv9_2),.clk(gclk));
	jdff dff_B_IvxFYclK9_2(.din(w_dff_B_p80WPCGv9_2),.dout(w_dff_B_IvxFYclK9_2),.clk(gclk));
	jdff dff_B_83514W5S9_2(.din(w_dff_B_IvxFYclK9_2),.dout(w_dff_B_83514W5S9_2),.clk(gclk));
	jdff dff_B_gagttwTN8_2(.din(w_dff_B_83514W5S9_2),.dout(w_dff_B_gagttwTN8_2),.clk(gclk));
	jdff dff_B_fagEDV9h5_2(.din(w_dff_B_gagttwTN8_2),.dout(w_dff_B_fagEDV9h5_2),.clk(gclk));
	jdff dff_B_Wf05x0wK6_2(.din(w_dff_B_fagEDV9h5_2),.dout(w_dff_B_Wf05x0wK6_2),.clk(gclk));
	jdff dff_B_AHPGsVDo8_2(.din(w_dff_B_Wf05x0wK6_2),.dout(w_dff_B_AHPGsVDo8_2),.clk(gclk));
	jdff dff_B_eImlIFJa4_2(.din(w_dff_B_AHPGsVDo8_2),.dout(w_dff_B_eImlIFJa4_2),.clk(gclk));
	jdff dff_B_EQlOIpa20_2(.din(w_dff_B_eImlIFJa4_2),.dout(w_dff_B_EQlOIpa20_2),.clk(gclk));
	jdff dff_B_bTKE2vxA3_2(.din(w_dff_B_EQlOIpa20_2),.dout(w_dff_B_bTKE2vxA3_2),.clk(gclk));
	jdff dff_B_dMcF30JL8_2(.din(w_dff_B_bTKE2vxA3_2),.dout(w_dff_B_dMcF30JL8_2),.clk(gclk));
	jdff dff_B_XDxMHo5Z4_2(.din(w_dff_B_dMcF30JL8_2),.dout(w_dff_B_XDxMHo5Z4_2),.clk(gclk));
	jdff dff_B_rdtuf9CZ9_2(.din(w_dff_B_XDxMHo5Z4_2),.dout(w_dff_B_rdtuf9CZ9_2),.clk(gclk));
	jdff dff_B_UQtSHOaW8_2(.din(w_dff_B_rdtuf9CZ9_2),.dout(w_dff_B_UQtSHOaW8_2),.clk(gclk));
	jdff dff_B_Ymx0eTka8_2(.din(w_dff_B_UQtSHOaW8_2),.dout(w_dff_B_Ymx0eTka8_2),.clk(gclk));
	jdff dff_B_K9MfCiiH9_2(.din(w_dff_B_Ymx0eTka8_2),.dout(w_dff_B_K9MfCiiH9_2),.clk(gclk));
	jdff dff_B_gKd82W6n2_1(.din(n1065),.dout(w_dff_B_gKd82W6n2_1),.clk(gclk));
	jdff dff_B_k0xdLmBg4_2(.din(n966),.dout(w_dff_B_k0xdLmBg4_2),.clk(gclk));
	jdff dff_B_VRLMVOOx8_2(.din(w_dff_B_k0xdLmBg4_2),.dout(w_dff_B_VRLMVOOx8_2),.clk(gclk));
	jdff dff_B_BRIZJtgZ4_2(.din(w_dff_B_VRLMVOOx8_2),.dout(w_dff_B_BRIZJtgZ4_2),.clk(gclk));
	jdff dff_B_IkzqHC132_2(.din(w_dff_B_BRIZJtgZ4_2),.dout(w_dff_B_IkzqHC132_2),.clk(gclk));
	jdff dff_B_tNdueXcE1_2(.din(w_dff_B_IkzqHC132_2),.dout(w_dff_B_tNdueXcE1_2),.clk(gclk));
	jdff dff_B_ffOYEBMO4_2(.din(w_dff_B_tNdueXcE1_2),.dout(w_dff_B_ffOYEBMO4_2),.clk(gclk));
	jdff dff_B_ESnLHkbH0_2(.din(w_dff_B_ffOYEBMO4_2),.dout(w_dff_B_ESnLHkbH0_2),.clk(gclk));
	jdff dff_B_FUYTKE2j4_2(.din(w_dff_B_ESnLHkbH0_2),.dout(w_dff_B_FUYTKE2j4_2),.clk(gclk));
	jdff dff_B_G8btJlP34_2(.din(w_dff_B_FUYTKE2j4_2),.dout(w_dff_B_G8btJlP34_2),.clk(gclk));
	jdff dff_B_k4qDj2Ga0_2(.din(w_dff_B_G8btJlP34_2),.dout(w_dff_B_k4qDj2Ga0_2),.clk(gclk));
	jdff dff_B_BXDDCU8X4_2(.din(w_dff_B_k4qDj2Ga0_2),.dout(w_dff_B_BXDDCU8X4_2),.clk(gclk));
	jdff dff_B_0rgr56EP8_2(.din(w_dff_B_BXDDCU8X4_2),.dout(w_dff_B_0rgr56EP8_2),.clk(gclk));
	jdff dff_B_NgqsGmwE2_2(.din(w_dff_B_0rgr56EP8_2),.dout(w_dff_B_NgqsGmwE2_2),.clk(gclk));
	jdff dff_B_lpKppnX52_2(.din(w_dff_B_NgqsGmwE2_2),.dout(w_dff_B_lpKppnX52_2),.clk(gclk));
	jdff dff_B_NiP8qZpS5_2(.din(w_dff_B_lpKppnX52_2),.dout(w_dff_B_NiP8qZpS5_2),.clk(gclk));
	jdff dff_B_uzvUZMxA4_2(.din(w_dff_B_NiP8qZpS5_2),.dout(w_dff_B_uzvUZMxA4_2),.clk(gclk));
	jdff dff_B_ZlbwXcYs5_2(.din(w_dff_B_uzvUZMxA4_2),.dout(w_dff_B_ZlbwXcYs5_2),.clk(gclk));
	jdff dff_B_N01fWury7_2(.din(w_dff_B_ZlbwXcYs5_2),.dout(w_dff_B_N01fWury7_2),.clk(gclk));
	jdff dff_B_izJRony38_2(.din(w_dff_B_N01fWury7_2),.dout(w_dff_B_izJRony38_2),.clk(gclk));
	jdff dff_B_tEBojRND8_2(.din(w_dff_B_izJRony38_2),.dout(w_dff_B_tEBojRND8_2),.clk(gclk));
	jdff dff_B_0hkuzV6i5_2(.din(w_dff_B_tEBojRND8_2),.dout(w_dff_B_0hkuzV6i5_2),.clk(gclk));
	jdff dff_B_dgR86CNW8_2(.din(w_dff_B_0hkuzV6i5_2),.dout(w_dff_B_dgR86CNW8_2),.clk(gclk));
	jdff dff_B_zYhZMvND2_2(.din(w_dff_B_dgR86CNW8_2),.dout(w_dff_B_zYhZMvND2_2),.clk(gclk));
	jdff dff_B_FLVCCj0G8_2(.din(w_dff_B_zYhZMvND2_2),.dout(w_dff_B_FLVCCj0G8_2),.clk(gclk));
	jdff dff_B_hAwQIO8k7_2(.din(w_dff_B_FLVCCj0G8_2),.dout(w_dff_B_hAwQIO8k7_2),.clk(gclk));
	jdff dff_B_cmJXqYMn6_2(.din(w_dff_B_hAwQIO8k7_2),.dout(w_dff_B_cmJXqYMn6_2),.clk(gclk));
	jdff dff_B_qeQMGMeM3_2(.din(w_dff_B_cmJXqYMn6_2),.dout(w_dff_B_qeQMGMeM3_2),.clk(gclk));
	jdff dff_B_U38vW7tC1_2(.din(w_dff_B_qeQMGMeM3_2),.dout(w_dff_B_U38vW7tC1_2),.clk(gclk));
	jdff dff_B_hSUeKmrL0_2(.din(w_dff_B_U38vW7tC1_2),.dout(w_dff_B_hSUeKmrL0_2),.clk(gclk));
	jdff dff_B_kCfO6Aus2_1(.din(n967),.dout(w_dff_B_kCfO6Aus2_1),.clk(gclk));
	jdff dff_B_PbN4Eizn7_2(.din(n861),.dout(w_dff_B_PbN4Eizn7_2),.clk(gclk));
	jdff dff_B_dwGTMwxF7_2(.din(w_dff_B_PbN4Eizn7_2),.dout(w_dff_B_dwGTMwxF7_2),.clk(gclk));
	jdff dff_B_cog3cDJ09_2(.din(w_dff_B_dwGTMwxF7_2),.dout(w_dff_B_cog3cDJ09_2),.clk(gclk));
	jdff dff_B_PO7USqUY7_2(.din(w_dff_B_cog3cDJ09_2),.dout(w_dff_B_PO7USqUY7_2),.clk(gclk));
	jdff dff_B_4DxmM4Yi2_2(.din(w_dff_B_PO7USqUY7_2),.dout(w_dff_B_4DxmM4Yi2_2),.clk(gclk));
	jdff dff_B_fpKF7vWF4_2(.din(w_dff_B_4DxmM4Yi2_2),.dout(w_dff_B_fpKF7vWF4_2),.clk(gclk));
	jdff dff_B_E6J55IHH9_2(.din(w_dff_B_fpKF7vWF4_2),.dout(w_dff_B_E6J55IHH9_2),.clk(gclk));
	jdff dff_B_ptzncvBY9_2(.din(w_dff_B_E6J55IHH9_2),.dout(w_dff_B_ptzncvBY9_2),.clk(gclk));
	jdff dff_B_cyAbCoaC9_2(.din(w_dff_B_ptzncvBY9_2),.dout(w_dff_B_cyAbCoaC9_2),.clk(gclk));
	jdff dff_B_bWapu2ob4_2(.din(w_dff_B_cyAbCoaC9_2),.dout(w_dff_B_bWapu2ob4_2),.clk(gclk));
	jdff dff_B_7ry2q6NH6_2(.din(w_dff_B_bWapu2ob4_2),.dout(w_dff_B_7ry2q6NH6_2),.clk(gclk));
	jdff dff_B_eP9fNeyA4_2(.din(w_dff_B_7ry2q6NH6_2),.dout(w_dff_B_eP9fNeyA4_2),.clk(gclk));
	jdff dff_B_eGQr13TS4_2(.din(w_dff_B_eP9fNeyA4_2),.dout(w_dff_B_eGQr13TS4_2),.clk(gclk));
	jdff dff_B_OxZD4LAk5_2(.din(w_dff_B_eGQr13TS4_2),.dout(w_dff_B_OxZD4LAk5_2),.clk(gclk));
	jdff dff_B_UBY4ksMm9_2(.din(w_dff_B_OxZD4LAk5_2),.dout(w_dff_B_UBY4ksMm9_2),.clk(gclk));
	jdff dff_B_tTd7OPdb0_2(.din(w_dff_B_UBY4ksMm9_2),.dout(w_dff_B_tTd7OPdb0_2),.clk(gclk));
	jdff dff_B_SHeUR4Sv5_2(.din(w_dff_B_tTd7OPdb0_2),.dout(w_dff_B_SHeUR4Sv5_2),.clk(gclk));
	jdff dff_B_8eaMojvU9_2(.din(w_dff_B_SHeUR4Sv5_2),.dout(w_dff_B_8eaMojvU9_2),.clk(gclk));
	jdff dff_B_OUWETMbk1_2(.din(w_dff_B_8eaMojvU9_2),.dout(w_dff_B_OUWETMbk1_2),.clk(gclk));
	jdff dff_B_90v5L3Bz6_2(.din(w_dff_B_OUWETMbk1_2),.dout(w_dff_B_90v5L3Bz6_2),.clk(gclk));
	jdff dff_B_xO9qI2a85_2(.din(w_dff_B_90v5L3Bz6_2),.dout(w_dff_B_xO9qI2a85_2),.clk(gclk));
	jdff dff_B_EfJ9Vx9R3_2(.din(w_dff_B_xO9qI2a85_2),.dout(w_dff_B_EfJ9Vx9R3_2),.clk(gclk));
	jdff dff_B_Rvcy1IOO3_2(.din(w_dff_B_EfJ9Vx9R3_2),.dout(w_dff_B_Rvcy1IOO3_2),.clk(gclk));
	jdff dff_B_vIhzUtvF0_2(.din(w_dff_B_Rvcy1IOO3_2),.dout(w_dff_B_vIhzUtvF0_2),.clk(gclk));
	jdff dff_B_ldwTfSl73_2(.din(w_dff_B_vIhzUtvF0_2),.dout(w_dff_B_ldwTfSl73_2),.clk(gclk));
	jdff dff_B_bsFbhQmc0_2(.din(w_dff_B_ldwTfSl73_2),.dout(w_dff_B_bsFbhQmc0_2),.clk(gclk));
	jdff dff_B_Nv9sc4k00_1(.din(n862),.dout(w_dff_B_Nv9sc4k00_1),.clk(gclk));
	jdff dff_B_J9T8q5a18_2(.din(n762),.dout(w_dff_B_J9T8q5a18_2),.clk(gclk));
	jdff dff_B_ZbyGjajf2_2(.din(w_dff_B_J9T8q5a18_2),.dout(w_dff_B_ZbyGjajf2_2),.clk(gclk));
	jdff dff_B_NUel66ar8_2(.din(w_dff_B_ZbyGjajf2_2),.dout(w_dff_B_NUel66ar8_2),.clk(gclk));
	jdff dff_B_TNfSqxTJ1_2(.din(w_dff_B_NUel66ar8_2),.dout(w_dff_B_TNfSqxTJ1_2),.clk(gclk));
	jdff dff_B_OYSSLdlg7_2(.din(w_dff_B_TNfSqxTJ1_2),.dout(w_dff_B_OYSSLdlg7_2),.clk(gclk));
	jdff dff_B_OeFb2pvZ6_2(.din(w_dff_B_OYSSLdlg7_2),.dout(w_dff_B_OeFb2pvZ6_2),.clk(gclk));
	jdff dff_B_xiEhIQEO9_2(.din(w_dff_B_OeFb2pvZ6_2),.dout(w_dff_B_xiEhIQEO9_2),.clk(gclk));
	jdff dff_B_GxzQNKvI3_2(.din(w_dff_B_xiEhIQEO9_2),.dout(w_dff_B_GxzQNKvI3_2),.clk(gclk));
	jdff dff_B_2rAVyXYa2_2(.din(w_dff_B_GxzQNKvI3_2),.dout(w_dff_B_2rAVyXYa2_2),.clk(gclk));
	jdff dff_B_9XTBTupQ8_2(.din(w_dff_B_2rAVyXYa2_2),.dout(w_dff_B_9XTBTupQ8_2),.clk(gclk));
	jdff dff_B_28YkXFdP4_2(.din(w_dff_B_9XTBTupQ8_2),.dout(w_dff_B_28YkXFdP4_2),.clk(gclk));
	jdff dff_B_PPAgc3366_2(.din(w_dff_B_28YkXFdP4_2),.dout(w_dff_B_PPAgc3366_2),.clk(gclk));
	jdff dff_B_NP0XiZvg9_2(.din(w_dff_B_PPAgc3366_2),.dout(w_dff_B_NP0XiZvg9_2),.clk(gclk));
	jdff dff_B_yDuHGVi34_2(.din(w_dff_B_NP0XiZvg9_2),.dout(w_dff_B_yDuHGVi34_2),.clk(gclk));
	jdff dff_B_wj3lF2p25_2(.din(w_dff_B_yDuHGVi34_2),.dout(w_dff_B_wj3lF2p25_2),.clk(gclk));
	jdff dff_B_yJ5YPjel7_2(.din(w_dff_B_wj3lF2p25_2),.dout(w_dff_B_yJ5YPjel7_2),.clk(gclk));
	jdff dff_B_rqKP1Z425_2(.din(w_dff_B_yJ5YPjel7_2),.dout(w_dff_B_rqKP1Z425_2),.clk(gclk));
	jdff dff_B_h2d35uWt7_2(.din(w_dff_B_rqKP1Z425_2),.dout(w_dff_B_h2d35uWt7_2),.clk(gclk));
	jdff dff_B_5SmefWIh7_2(.din(w_dff_B_h2d35uWt7_2),.dout(w_dff_B_5SmefWIh7_2),.clk(gclk));
	jdff dff_B_8qpIUJ1q2_2(.din(w_dff_B_5SmefWIh7_2),.dout(w_dff_B_8qpIUJ1q2_2),.clk(gclk));
	jdff dff_B_WV1L8tsl5_2(.din(w_dff_B_8qpIUJ1q2_2),.dout(w_dff_B_WV1L8tsl5_2),.clk(gclk));
	jdff dff_B_bB0kAjRn7_2(.din(w_dff_B_WV1L8tsl5_2),.dout(w_dff_B_bB0kAjRn7_2),.clk(gclk));
	jdff dff_B_jXm3dBaj8_2(.din(w_dff_B_bB0kAjRn7_2),.dout(w_dff_B_jXm3dBaj8_2),.clk(gclk));
	jdff dff_B_NfzOU8uG7_1(.din(n763),.dout(w_dff_B_NfzOU8uG7_1),.clk(gclk));
	jdff dff_B_UddFAk9F3_2(.din(n669),.dout(w_dff_B_UddFAk9F3_2),.clk(gclk));
	jdff dff_B_aF20CRb32_2(.din(w_dff_B_UddFAk9F3_2),.dout(w_dff_B_aF20CRb32_2),.clk(gclk));
	jdff dff_B_Mm38oxW87_2(.din(w_dff_B_aF20CRb32_2),.dout(w_dff_B_Mm38oxW87_2),.clk(gclk));
	jdff dff_B_0AWD1DAx1_2(.din(w_dff_B_Mm38oxW87_2),.dout(w_dff_B_0AWD1DAx1_2),.clk(gclk));
	jdff dff_B_j55uUv796_2(.din(w_dff_B_0AWD1DAx1_2),.dout(w_dff_B_j55uUv796_2),.clk(gclk));
	jdff dff_B_zcBHRLik0_2(.din(w_dff_B_j55uUv796_2),.dout(w_dff_B_zcBHRLik0_2),.clk(gclk));
	jdff dff_B_a2gGLxfn6_2(.din(w_dff_B_zcBHRLik0_2),.dout(w_dff_B_a2gGLxfn6_2),.clk(gclk));
	jdff dff_B_CODX0LgQ2_2(.din(w_dff_B_a2gGLxfn6_2),.dout(w_dff_B_CODX0LgQ2_2),.clk(gclk));
	jdff dff_B_KJRbJor27_2(.din(w_dff_B_CODX0LgQ2_2),.dout(w_dff_B_KJRbJor27_2),.clk(gclk));
	jdff dff_B_Zn7slPYZ7_2(.din(w_dff_B_KJRbJor27_2),.dout(w_dff_B_Zn7slPYZ7_2),.clk(gclk));
	jdff dff_B_EGJCjpjA7_2(.din(w_dff_B_Zn7slPYZ7_2),.dout(w_dff_B_EGJCjpjA7_2),.clk(gclk));
	jdff dff_B_alIpKFw52_2(.din(w_dff_B_EGJCjpjA7_2),.dout(w_dff_B_alIpKFw52_2),.clk(gclk));
	jdff dff_B_w5LNbcyV9_2(.din(w_dff_B_alIpKFw52_2),.dout(w_dff_B_w5LNbcyV9_2),.clk(gclk));
	jdff dff_B_983xOmMV2_2(.din(w_dff_B_w5LNbcyV9_2),.dout(w_dff_B_983xOmMV2_2),.clk(gclk));
	jdff dff_B_h8Q7jCOb0_2(.din(w_dff_B_983xOmMV2_2),.dout(w_dff_B_h8Q7jCOb0_2),.clk(gclk));
	jdff dff_B_wGWHjVzP5_2(.din(w_dff_B_h8Q7jCOb0_2),.dout(w_dff_B_wGWHjVzP5_2),.clk(gclk));
	jdff dff_B_eQ816E361_2(.din(w_dff_B_wGWHjVzP5_2),.dout(w_dff_B_eQ816E361_2),.clk(gclk));
	jdff dff_B_C7wYALGK1_2(.din(w_dff_B_eQ816E361_2),.dout(w_dff_B_C7wYALGK1_2),.clk(gclk));
	jdff dff_B_aI2f7H149_2(.din(w_dff_B_C7wYALGK1_2),.dout(w_dff_B_aI2f7H149_2),.clk(gclk));
	jdff dff_B_Ef4mkVVx3_2(.din(w_dff_B_aI2f7H149_2),.dout(w_dff_B_Ef4mkVVx3_2),.clk(gclk));
	jdff dff_B_aS9WQCEK1_1(.din(n670),.dout(w_dff_B_aS9WQCEK1_1),.clk(gclk));
	jdff dff_B_XvBRwcpl7_2(.din(n583),.dout(w_dff_B_XvBRwcpl7_2),.clk(gclk));
	jdff dff_B_EHf0HZtO6_2(.din(w_dff_B_XvBRwcpl7_2),.dout(w_dff_B_EHf0HZtO6_2),.clk(gclk));
	jdff dff_B_FFe7cNla8_2(.din(w_dff_B_EHf0HZtO6_2),.dout(w_dff_B_FFe7cNla8_2),.clk(gclk));
	jdff dff_B_5RicMekn8_2(.din(w_dff_B_FFe7cNla8_2),.dout(w_dff_B_5RicMekn8_2),.clk(gclk));
	jdff dff_B_o3ALsuSM7_2(.din(w_dff_B_5RicMekn8_2),.dout(w_dff_B_o3ALsuSM7_2),.clk(gclk));
	jdff dff_B_Ctyu6zb89_2(.din(w_dff_B_o3ALsuSM7_2),.dout(w_dff_B_Ctyu6zb89_2),.clk(gclk));
	jdff dff_B_ccLgiHjv4_2(.din(w_dff_B_Ctyu6zb89_2),.dout(w_dff_B_ccLgiHjv4_2),.clk(gclk));
	jdff dff_B_CN69VyeF0_2(.din(w_dff_B_ccLgiHjv4_2),.dout(w_dff_B_CN69VyeF0_2),.clk(gclk));
	jdff dff_B_jHP4GolN1_2(.din(w_dff_B_CN69VyeF0_2),.dout(w_dff_B_jHP4GolN1_2),.clk(gclk));
	jdff dff_B_7VzO5X2y9_2(.din(w_dff_B_jHP4GolN1_2),.dout(w_dff_B_7VzO5X2y9_2),.clk(gclk));
	jdff dff_B_1zwhxOMR1_2(.din(w_dff_B_7VzO5X2y9_2),.dout(w_dff_B_1zwhxOMR1_2),.clk(gclk));
	jdff dff_B_dcc151WO0_2(.din(w_dff_B_1zwhxOMR1_2),.dout(w_dff_B_dcc151WO0_2),.clk(gclk));
	jdff dff_B_VGhdKhtI2_2(.din(w_dff_B_dcc151WO0_2),.dout(w_dff_B_VGhdKhtI2_2),.clk(gclk));
	jdff dff_B_YnkYjL2D3_2(.din(w_dff_B_VGhdKhtI2_2),.dout(w_dff_B_YnkYjL2D3_2),.clk(gclk));
	jdff dff_B_cs1K0E3V8_2(.din(w_dff_B_YnkYjL2D3_2),.dout(w_dff_B_cs1K0E3V8_2),.clk(gclk));
	jdff dff_B_lwA8I24v7_2(.din(w_dff_B_cs1K0E3V8_2),.dout(w_dff_B_lwA8I24v7_2),.clk(gclk));
	jdff dff_B_fFbzYEDd7_2(.din(w_dff_B_lwA8I24v7_2),.dout(w_dff_B_fFbzYEDd7_2),.clk(gclk));
	jdff dff_B_OlGt9Uuj4_1(.din(n584),.dout(w_dff_B_OlGt9Uuj4_1),.clk(gclk));
	jdff dff_B_ukYQadji0_2(.din(n504),.dout(w_dff_B_ukYQadji0_2),.clk(gclk));
	jdff dff_B_W4KVTdUj5_2(.din(w_dff_B_ukYQadji0_2),.dout(w_dff_B_W4KVTdUj5_2),.clk(gclk));
	jdff dff_B_hxCJIC1i1_2(.din(w_dff_B_W4KVTdUj5_2),.dout(w_dff_B_hxCJIC1i1_2),.clk(gclk));
	jdff dff_B_YkFgylAc6_2(.din(w_dff_B_hxCJIC1i1_2),.dout(w_dff_B_YkFgylAc6_2),.clk(gclk));
	jdff dff_B_azSjNYVm9_2(.din(w_dff_B_YkFgylAc6_2),.dout(w_dff_B_azSjNYVm9_2),.clk(gclk));
	jdff dff_B_nhe4O2Va9_2(.din(w_dff_B_azSjNYVm9_2),.dout(w_dff_B_nhe4O2Va9_2),.clk(gclk));
	jdff dff_B_RpVEfoGQ7_2(.din(w_dff_B_nhe4O2Va9_2),.dout(w_dff_B_RpVEfoGQ7_2),.clk(gclk));
	jdff dff_B_zH4DftIt4_2(.din(w_dff_B_RpVEfoGQ7_2),.dout(w_dff_B_zH4DftIt4_2),.clk(gclk));
	jdff dff_B_eCttojSS2_2(.din(w_dff_B_zH4DftIt4_2),.dout(w_dff_B_eCttojSS2_2),.clk(gclk));
	jdff dff_B_dVKWTuVr6_2(.din(w_dff_B_eCttojSS2_2),.dout(w_dff_B_dVKWTuVr6_2),.clk(gclk));
	jdff dff_B_tAecjG1c2_2(.din(w_dff_B_dVKWTuVr6_2),.dout(w_dff_B_tAecjG1c2_2),.clk(gclk));
	jdff dff_B_MQ9nJEQ77_2(.din(w_dff_B_tAecjG1c2_2),.dout(w_dff_B_MQ9nJEQ77_2),.clk(gclk));
	jdff dff_B_H8BgJNg37_2(.din(w_dff_B_MQ9nJEQ77_2),.dout(w_dff_B_H8BgJNg37_2),.clk(gclk));
	jdff dff_B_UOTUdhWY3_2(.din(w_dff_B_H8BgJNg37_2),.dout(w_dff_B_UOTUdhWY3_2),.clk(gclk));
	jdff dff_B_g62wjsut6_1(.din(n505),.dout(w_dff_B_g62wjsut6_1),.clk(gclk));
	jdff dff_B_mofUbUYw9_2(.din(n432),.dout(w_dff_B_mofUbUYw9_2),.clk(gclk));
	jdff dff_B_niybe1Iv7_2(.din(w_dff_B_mofUbUYw9_2),.dout(w_dff_B_niybe1Iv7_2),.clk(gclk));
	jdff dff_B_ZyESmRrZ5_2(.din(w_dff_B_niybe1Iv7_2),.dout(w_dff_B_ZyESmRrZ5_2),.clk(gclk));
	jdff dff_B_EPUifdh25_2(.din(w_dff_B_ZyESmRrZ5_2),.dout(w_dff_B_EPUifdh25_2),.clk(gclk));
	jdff dff_B_rja1QFI06_2(.din(w_dff_B_EPUifdh25_2),.dout(w_dff_B_rja1QFI06_2),.clk(gclk));
	jdff dff_B_R8tjpMQq4_2(.din(w_dff_B_rja1QFI06_2),.dout(w_dff_B_R8tjpMQq4_2),.clk(gclk));
	jdff dff_B_vCFwQKYd9_2(.din(w_dff_B_R8tjpMQq4_2),.dout(w_dff_B_vCFwQKYd9_2),.clk(gclk));
	jdff dff_B_nzeE4d2Q3_2(.din(w_dff_B_vCFwQKYd9_2),.dout(w_dff_B_nzeE4d2Q3_2),.clk(gclk));
	jdff dff_B_wzXhIDkY3_2(.din(w_dff_B_nzeE4d2Q3_2),.dout(w_dff_B_wzXhIDkY3_2),.clk(gclk));
	jdff dff_B_YYVXrBV72_2(.din(w_dff_B_wzXhIDkY3_2),.dout(w_dff_B_YYVXrBV72_2),.clk(gclk));
	jdff dff_B_wz3dzYdM9_2(.din(w_dff_B_YYVXrBV72_2),.dout(w_dff_B_wz3dzYdM9_2),.clk(gclk));
	jdff dff_B_j6F4Nlxt6_2(.din(n435),.dout(w_dff_B_j6F4Nlxt6_2),.clk(gclk));
	jdff dff_B_qL2BFsb78_1(.din(n433),.dout(w_dff_B_qL2BFsb78_1),.clk(gclk));
	jdff dff_B_3Se7Sk4K0_2(.din(n368),.dout(w_dff_B_3Se7Sk4K0_2),.clk(gclk));
	jdff dff_B_2osNilFo9_2(.din(w_dff_B_3Se7Sk4K0_2),.dout(w_dff_B_2osNilFo9_2),.clk(gclk));
	jdff dff_B_xnS6lx2i0_2(.din(w_dff_B_2osNilFo9_2),.dout(w_dff_B_xnS6lx2i0_2),.clk(gclk));
	jdff dff_B_ehvJyKEo2_2(.din(w_dff_B_xnS6lx2i0_2),.dout(w_dff_B_ehvJyKEo2_2),.clk(gclk));
	jdff dff_B_AdIRERwX0_2(.din(w_dff_B_ehvJyKEo2_2),.dout(w_dff_B_AdIRERwX0_2),.clk(gclk));
	jdff dff_B_OkaMSu4h5_2(.din(w_dff_B_AdIRERwX0_2),.dout(w_dff_B_OkaMSu4h5_2),.clk(gclk));
	jdff dff_B_9r95EjvW0_2(.din(w_dff_B_OkaMSu4h5_2),.dout(w_dff_B_9r95EjvW0_2),.clk(gclk));
	jdff dff_B_8bw6Fr9D8_1(.din(n369),.dout(w_dff_B_8bw6Fr9D8_1),.clk(gclk));
	jdff dff_B_F4LgOeMa1_2(.din(n310),.dout(w_dff_B_F4LgOeMa1_2),.clk(gclk));
	jdff dff_B_Uly7U9a64_2(.din(w_dff_B_F4LgOeMa1_2),.dout(w_dff_B_Uly7U9a64_2),.clk(gclk));
	jdff dff_B_Ytmx2Tpe3_2(.din(w_dff_B_Uly7U9a64_2),.dout(w_dff_B_Ytmx2Tpe3_2),.clk(gclk));
	jdff dff_B_CpkB4cPl0_2(.din(w_dff_B_Ytmx2Tpe3_2),.dout(w_dff_B_CpkB4cPl0_2),.clk(gclk));
	jdff dff_B_COEn0i7q4_1(.din(n312),.dout(w_dff_B_COEn0i7q4_1),.clk(gclk));
	jdff dff_A_aBDBlh6d9_0(.dout(w_n258_0[0]),.din(w_dff_A_aBDBlh6d9_0),.clk(gclk));
	jdff dff_A_OWBOdTT50_1(.dout(w_n258_0[1]),.din(w_dff_A_OWBOdTT50_1),.clk(gclk));
	jdff dff_A_eBdNRukX7_1(.dout(w_dff_A_OWBOdTT50_1),.din(w_dff_A_eBdNRukX7_1),.clk(gclk));
	jdff dff_B_dNZdGybo7_1(.din(n1563),.dout(w_dff_B_dNZdGybo7_1),.clk(gclk));
	jdff dff_B_OaC6pXkf2_2(.din(n1497),.dout(w_dff_B_OaC6pXkf2_2),.clk(gclk));
	jdff dff_B_bzQZHME51_2(.din(w_dff_B_OaC6pXkf2_2),.dout(w_dff_B_bzQZHME51_2),.clk(gclk));
	jdff dff_B_qjo4ML0j0_2(.din(w_dff_B_bzQZHME51_2),.dout(w_dff_B_qjo4ML0j0_2),.clk(gclk));
	jdff dff_B_lW6ummAk4_2(.din(w_dff_B_qjo4ML0j0_2),.dout(w_dff_B_lW6ummAk4_2),.clk(gclk));
	jdff dff_B_HAMdJXqj4_2(.din(w_dff_B_lW6ummAk4_2),.dout(w_dff_B_HAMdJXqj4_2),.clk(gclk));
	jdff dff_B_SP7WhHL67_2(.din(w_dff_B_HAMdJXqj4_2),.dout(w_dff_B_SP7WhHL67_2),.clk(gclk));
	jdff dff_B_LaQCwOWy0_2(.din(w_dff_B_SP7WhHL67_2),.dout(w_dff_B_LaQCwOWy0_2),.clk(gclk));
	jdff dff_B_14Xlus2t8_2(.din(w_dff_B_LaQCwOWy0_2),.dout(w_dff_B_14Xlus2t8_2),.clk(gclk));
	jdff dff_B_xOSKmMFo8_2(.din(w_dff_B_14Xlus2t8_2),.dout(w_dff_B_xOSKmMFo8_2),.clk(gclk));
	jdff dff_B_V5YreD3D5_2(.din(w_dff_B_xOSKmMFo8_2),.dout(w_dff_B_V5YreD3D5_2),.clk(gclk));
	jdff dff_B_uvhoH1SS8_2(.din(w_dff_B_V5YreD3D5_2),.dout(w_dff_B_uvhoH1SS8_2),.clk(gclk));
	jdff dff_B_f8BKMykT4_2(.din(w_dff_B_uvhoH1SS8_2),.dout(w_dff_B_f8BKMykT4_2),.clk(gclk));
	jdff dff_B_zSr0kpJE8_2(.din(w_dff_B_f8BKMykT4_2),.dout(w_dff_B_zSr0kpJE8_2),.clk(gclk));
	jdff dff_B_xZbkgrvL4_2(.din(w_dff_B_zSr0kpJE8_2),.dout(w_dff_B_xZbkgrvL4_2),.clk(gclk));
	jdff dff_B_dXkBzECY6_2(.din(w_dff_B_xZbkgrvL4_2),.dout(w_dff_B_dXkBzECY6_2),.clk(gclk));
	jdff dff_B_yjUKA5dm2_2(.din(w_dff_B_dXkBzECY6_2),.dout(w_dff_B_yjUKA5dm2_2),.clk(gclk));
	jdff dff_B_vZeAWra68_2(.din(w_dff_B_yjUKA5dm2_2),.dout(w_dff_B_vZeAWra68_2),.clk(gclk));
	jdff dff_B_eB5GVjmy3_2(.din(w_dff_B_vZeAWra68_2),.dout(w_dff_B_eB5GVjmy3_2),.clk(gclk));
	jdff dff_B_ZwGW23gW1_2(.din(w_dff_B_eB5GVjmy3_2),.dout(w_dff_B_ZwGW23gW1_2),.clk(gclk));
	jdff dff_B_0gVfbluu6_2(.din(w_dff_B_ZwGW23gW1_2),.dout(w_dff_B_0gVfbluu6_2),.clk(gclk));
	jdff dff_B_eFVkGurk6_2(.din(w_dff_B_0gVfbluu6_2),.dout(w_dff_B_eFVkGurk6_2),.clk(gclk));
	jdff dff_B_XJM0d1OB9_2(.din(w_dff_B_eFVkGurk6_2),.dout(w_dff_B_XJM0d1OB9_2),.clk(gclk));
	jdff dff_B_ouWZbJ9b9_2(.din(w_dff_B_XJM0d1OB9_2),.dout(w_dff_B_ouWZbJ9b9_2),.clk(gclk));
	jdff dff_B_19cuWiUj1_2(.din(w_dff_B_ouWZbJ9b9_2),.dout(w_dff_B_19cuWiUj1_2),.clk(gclk));
	jdff dff_B_IvR2Vxpf3_2(.din(w_dff_B_19cuWiUj1_2),.dout(w_dff_B_IvR2Vxpf3_2),.clk(gclk));
	jdff dff_B_sAfgoOGC1_2(.din(w_dff_B_IvR2Vxpf3_2),.dout(w_dff_B_sAfgoOGC1_2),.clk(gclk));
	jdff dff_B_oI9oCBLJ8_2(.din(w_dff_B_sAfgoOGC1_2),.dout(w_dff_B_oI9oCBLJ8_2),.clk(gclk));
	jdff dff_B_GAGxHBL25_2(.din(w_dff_B_oI9oCBLJ8_2),.dout(w_dff_B_GAGxHBL25_2),.clk(gclk));
	jdff dff_B_57mQVH8X6_2(.din(w_dff_B_GAGxHBL25_2),.dout(w_dff_B_57mQVH8X6_2),.clk(gclk));
	jdff dff_B_Ahei8Xw10_2(.din(w_dff_B_57mQVH8X6_2),.dout(w_dff_B_Ahei8Xw10_2),.clk(gclk));
	jdff dff_B_zNAtCrG97_2(.din(w_dff_B_Ahei8Xw10_2),.dout(w_dff_B_zNAtCrG97_2),.clk(gclk));
	jdff dff_B_zG7eIA2k6_2(.din(w_dff_B_zNAtCrG97_2),.dout(w_dff_B_zG7eIA2k6_2),.clk(gclk));
	jdff dff_B_WLeD4J7R0_2(.din(w_dff_B_zG7eIA2k6_2),.dout(w_dff_B_WLeD4J7R0_2),.clk(gclk));
	jdff dff_B_x1VE0BXf2_2(.din(w_dff_B_WLeD4J7R0_2),.dout(w_dff_B_x1VE0BXf2_2),.clk(gclk));
	jdff dff_B_3UDgbXl85_2(.din(w_dff_B_x1VE0BXf2_2),.dout(w_dff_B_3UDgbXl85_2),.clk(gclk));
	jdff dff_B_w7r14DpS8_2(.din(w_dff_B_3UDgbXl85_2),.dout(w_dff_B_w7r14DpS8_2),.clk(gclk));
	jdff dff_B_TLOdqBCR5_2(.din(w_dff_B_w7r14DpS8_2),.dout(w_dff_B_TLOdqBCR5_2),.clk(gclk));
	jdff dff_B_oqcAXjZY4_2(.din(w_dff_B_TLOdqBCR5_2),.dout(w_dff_B_oqcAXjZY4_2),.clk(gclk));
	jdff dff_B_WCVgGZJd3_2(.din(w_dff_B_oqcAXjZY4_2),.dout(w_dff_B_WCVgGZJd3_2),.clk(gclk));
	jdff dff_B_gxzjjlWO1_2(.din(w_dff_B_WCVgGZJd3_2),.dout(w_dff_B_gxzjjlWO1_2),.clk(gclk));
	jdff dff_B_JQKp7SRZ4_2(.din(w_dff_B_gxzjjlWO1_2),.dout(w_dff_B_JQKp7SRZ4_2),.clk(gclk));
	jdff dff_B_dqZnbUCp3_2(.din(w_dff_B_JQKp7SRZ4_2),.dout(w_dff_B_dqZnbUCp3_2),.clk(gclk));
	jdff dff_B_p47rBmF72_2(.din(w_dff_B_dqZnbUCp3_2),.dout(w_dff_B_p47rBmF72_2),.clk(gclk));
	jdff dff_B_rFbxQWOV3_2(.din(w_dff_B_p47rBmF72_2),.dout(w_dff_B_rFbxQWOV3_2),.clk(gclk));
	jdff dff_B_syuyrcj01_2(.din(w_dff_B_rFbxQWOV3_2),.dout(w_dff_B_syuyrcj01_2),.clk(gclk));
	jdff dff_B_p6FGVhTh7_2(.din(w_dff_B_syuyrcj01_2),.dout(w_dff_B_p6FGVhTh7_2),.clk(gclk));
	jdff dff_B_f5hCBJZx7_2(.din(w_dff_B_p6FGVhTh7_2),.dout(w_dff_B_f5hCBJZx7_2),.clk(gclk));
	jdff dff_B_rSxV2MYi3_0(.din(n1562),.dout(w_dff_B_rSxV2MYi3_0),.clk(gclk));
	jdff dff_A_fK9qtCNH5_1(.dout(w_n1550_0[1]),.din(w_dff_A_fK9qtCNH5_1),.clk(gclk));
	jdff dff_B_pVRMKH112_1(.din(n1498),.dout(w_dff_B_pVRMKH112_1),.clk(gclk));
	jdff dff_B_2s4yTaNW8_2(.din(n1426),.dout(w_dff_B_2s4yTaNW8_2),.clk(gclk));
	jdff dff_B_339u2ylJ9_2(.din(w_dff_B_2s4yTaNW8_2),.dout(w_dff_B_339u2ylJ9_2),.clk(gclk));
	jdff dff_B_pqbFETGt8_2(.din(w_dff_B_339u2ylJ9_2),.dout(w_dff_B_pqbFETGt8_2),.clk(gclk));
	jdff dff_B_NG2Kevfy5_2(.din(w_dff_B_pqbFETGt8_2),.dout(w_dff_B_NG2Kevfy5_2),.clk(gclk));
	jdff dff_B_nlJtgKHu2_2(.din(w_dff_B_NG2Kevfy5_2),.dout(w_dff_B_nlJtgKHu2_2),.clk(gclk));
	jdff dff_B_LE3cqdHL7_2(.din(w_dff_B_nlJtgKHu2_2),.dout(w_dff_B_LE3cqdHL7_2),.clk(gclk));
	jdff dff_B_WfpD5SbF6_2(.din(w_dff_B_LE3cqdHL7_2),.dout(w_dff_B_WfpD5SbF6_2),.clk(gclk));
	jdff dff_B_LKhtnuhk3_2(.din(w_dff_B_WfpD5SbF6_2),.dout(w_dff_B_LKhtnuhk3_2),.clk(gclk));
	jdff dff_B_j0c0Kj3Y1_2(.din(w_dff_B_LKhtnuhk3_2),.dout(w_dff_B_j0c0Kj3Y1_2),.clk(gclk));
	jdff dff_B_njHtBhzj3_2(.din(w_dff_B_j0c0Kj3Y1_2),.dout(w_dff_B_njHtBhzj3_2),.clk(gclk));
	jdff dff_B_kAtIHfPU9_2(.din(w_dff_B_njHtBhzj3_2),.dout(w_dff_B_kAtIHfPU9_2),.clk(gclk));
	jdff dff_B_LHFPeuCu5_2(.din(w_dff_B_kAtIHfPU9_2),.dout(w_dff_B_LHFPeuCu5_2),.clk(gclk));
	jdff dff_B_5UO3cQxI7_2(.din(w_dff_B_LHFPeuCu5_2),.dout(w_dff_B_5UO3cQxI7_2),.clk(gclk));
	jdff dff_B_MspLqAmI8_2(.din(w_dff_B_5UO3cQxI7_2),.dout(w_dff_B_MspLqAmI8_2),.clk(gclk));
	jdff dff_B_16qeeGLi6_2(.din(w_dff_B_MspLqAmI8_2),.dout(w_dff_B_16qeeGLi6_2),.clk(gclk));
	jdff dff_B_77yuZhVP2_2(.din(w_dff_B_16qeeGLi6_2),.dout(w_dff_B_77yuZhVP2_2),.clk(gclk));
	jdff dff_B_p5eHDbOQ4_2(.din(w_dff_B_77yuZhVP2_2),.dout(w_dff_B_p5eHDbOQ4_2),.clk(gclk));
	jdff dff_B_iPzakK8z5_2(.din(w_dff_B_p5eHDbOQ4_2),.dout(w_dff_B_iPzakK8z5_2),.clk(gclk));
	jdff dff_B_PcNY3Rs13_2(.din(w_dff_B_iPzakK8z5_2),.dout(w_dff_B_PcNY3Rs13_2),.clk(gclk));
	jdff dff_B_a0ifAPls6_2(.din(w_dff_B_PcNY3Rs13_2),.dout(w_dff_B_a0ifAPls6_2),.clk(gclk));
	jdff dff_B_IzEMmRMk8_2(.din(w_dff_B_a0ifAPls6_2),.dout(w_dff_B_IzEMmRMk8_2),.clk(gclk));
	jdff dff_B_uDY1FGLF6_2(.din(w_dff_B_IzEMmRMk8_2),.dout(w_dff_B_uDY1FGLF6_2),.clk(gclk));
	jdff dff_B_YWYEcBk66_2(.din(w_dff_B_uDY1FGLF6_2),.dout(w_dff_B_YWYEcBk66_2),.clk(gclk));
	jdff dff_B_Jzjomdso8_2(.din(w_dff_B_YWYEcBk66_2),.dout(w_dff_B_Jzjomdso8_2),.clk(gclk));
	jdff dff_B_BOFqJPvP0_2(.din(w_dff_B_Jzjomdso8_2),.dout(w_dff_B_BOFqJPvP0_2),.clk(gclk));
	jdff dff_B_tBXtUiTt4_2(.din(w_dff_B_BOFqJPvP0_2),.dout(w_dff_B_tBXtUiTt4_2),.clk(gclk));
	jdff dff_B_U3lGBHK96_2(.din(w_dff_B_tBXtUiTt4_2),.dout(w_dff_B_U3lGBHK96_2),.clk(gclk));
	jdff dff_B_oqA7mvpU6_2(.din(w_dff_B_U3lGBHK96_2),.dout(w_dff_B_oqA7mvpU6_2),.clk(gclk));
	jdff dff_B_Wge6w4UP6_2(.din(w_dff_B_oqA7mvpU6_2),.dout(w_dff_B_Wge6w4UP6_2),.clk(gclk));
	jdff dff_B_TZBI3ML91_2(.din(w_dff_B_Wge6w4UP6_2),.dout(w_dff_B_TZBI3ML91_2),.clk(gclk));
	jdff dff_B_e3m7vQf03_2(.din(w_dff_B_TZBI3ML91_2),.dout(w_dff_B_e3m7vQf03_2),.clk(gclk));
	jdff dff_B_l9h8n5uz4_2(.din(w_dff_B_e3m7vQf03_2),.dout(w_dff_B_l9h8n5uz4_2),.clk(gclk));
	jdff dff_B_2smcDJBn8_2(.din(w_dff_B_l9h8n5uz4_2),.dout(w_dff_B_2smcDJBn8_2),.clk(gclk));
	jdff dff_B_l5yMxhnj3_2(.din(w_dff_B_2smcDJBn8_2),.dout(w_dff_B_l5yMxhnj3_2),.clk(gclk));
	jdff dff_B_S1eIQdOD7_2(.din(w_dff_B_l5yMxhnj3_2),.dout(w_dff_B_S1eIQdOD7_2),.clk(gclk));
	jdff dff_B_FWzn2Zgp8_2(.din(w_dff_B_S1eIQdOD7_2),.dout(w_dff_B_FWzn2Zgp8_2),.clk(gclk));
	jdff dff_B_Gr5JGbmA5_2(.din(w_dff_B_FWzn2Zgp8_2),.dout(w_dff_B_Gr5JGbmA5_2),.clk(gclk));
	jdff dff_B_cMdYXuJ37_2(.din(w_dff_B_Gr5JGbmA5_2),.dout(w_dff_B_cMdYXuJ37_2),.clk(gclk));
	jdff dff_B_HguAhdNx3_2(.din(w_dff_B_cMdYXuJ37_2),.dout(w_dff_B_HguAhdNx3_2),.clk(gclk));
	jdff dff_B_6Sa4aOd89_2(.din(w_dff_B_HguAhdNx3_2),.dout(w_dff_B_6Sa4aOd89_2),.clk(gclk));
	jdff dff_B_nEVlyori2_2(.din(w_dff_B_6Sa4aOd89_2),.dout(w_dff_B_nEVlyori2_2),.clk(gclk));
	jdff dff_B_Z9LoOTDA7_2(.din(w_dff_B_nEVlyori2_2),.dout(w_dff_B_Z9LoOTDA7_2),.clk(gclk));
	jdff dff_B_8w6Vab4P0_2(.din(n1479),.dout(w_dff_B_8w6Vab4P0_2),.clk(gclk));
	jdff dff_B_9e3ArnSM4_1(.din(n1427),.dout(w_dff_B_9e3ArnSM4_1),.clk(gclk));
	jdff dff_B_XfwUtztd4_2(.din(n1348),.dout(w_dff_B_XfwUtztd4_2),.clk(gclk));
	jdff dff_B_ZYpPyd7D8_2(.din(w_dff_B_XfwUtztd4_2),.dout(w_dff_B_ZYpPyd7D8_2),.clk(gclk));
	jdff dff_B_o8JqlCPX7_2(.din(w_dff_B_ZYpPyd7D8_2),.dout(w_dff_B_o8JqlCPX7_2),.clk(gclk));
	jdff dff_B_5PIcEdNX7_2(.din(w_dff_B_o8JqlCPX7_2),.dout(w_dff_B_5PIcEdNX7_2),.clk(gclk));
	jdff dff_B_omAJYMEv7_2(.din(w_dff_B_5PIcEdNX7_2),.dout(w_dff_B_omAJYMEv7_2),.clk(gclk));
	jdff dff_B_Wasq2FvN5_2(.din(w_dff_B_omAJYMEv7_2),.dout(w_dff_B_Wasq2FvN5_2),.clk(gclk));
	jdff dff_B_WscfOdyS2_2(.din(w_dff_B_Wasq2FvN5_2),.dout(w_dff_B_WscfOdyS2_2),.clk(gclk));
	jdff dff_B_5KsJoTbB1_2(.din(w_dff_B_WscfOdyS2_2),.dout(w_dff_B_5KsJoTbB1_2),.clk(gclk));
	jdff dff_B_Gu6FDvBM0_2(.din(w_dff_B_5KsJoTbB1_2),.dout(w_dff_B_Gu6FDvBM0_2),.clk(gclk));
	jdff dff_B_AMrgHlco9_2(.din(w_dff_B_Gu6FDvBM0_2),.dout(w_dff_B_AMrgHlco9_2),.clk(gclk));
	jdff dff_B_jTrfBuMJ3_2(.din(w_dff_B_AMrgHlco9_2),.dout(w_dff_B_jTrfBuMJ3_2),.clk(gclk));
	jdff dff_B_s60lqEXF6_2(.din(w_dff_B_jTrfBuMJ3_2),.dout(w_dff_B_s60lqEXF6_2),.clk(gclk));
	jdff dff_B_tqwzxJFg1_2(.din(w_dff_B_s60lqEXF6_2),.dout(w_dff_B_tqwzxJFg1_2),.clk(gclk));
	jdff dff_B_fBToE5Ig5_2(.din(w_dff_B_tqwzxJFg1_2),.dout(w_dff_B_fBToE5Ig5_2),.clk(gclk));
	jdff dff_B_KlosOtsY3_2(.din(w_dff_B_fBToE5Ig5_2),.dout(w_dff_B_KlosOtsY3_2),.clk(gclk));
	jdff dff_B_EtYeH5jM2_2(.din(w_dff_B_KlosOtsY3_2),.dout(w_dff_B_EtYeH5jM2_2),.clk(gclk));
	jdff dff_B_RDhSc2Hj0_2(.din(w_dff_B_EtYeH5jM2_2),.dout(w_dff_B_RDhSc2Hj0_2),.clk(gclk));
	jdff dff_B_9CaG2y445_2(.din(w_dff_B_RDhSc2Hj0_2),.dout(w_dff_B_9CaG2y445_2),.clk(gclk));
	jdff dff_B_zD1M4WBq9_2(.din(w_dff_B_9CaG2y445_2),.dout(w_dff_B_zD1M4WBq9_2),.clk(gclk));
	jdff dff_B_VCoDaFvr7_2(.din(w_dff_B_zD1M4WBq9_2),.dout(w_dff_B_VCoDaFvr7_2),.clk(gclk));
	jdff dff_B_qpvjGOiZ6_2(.din(w_dff_B_VCoDaFvr7_2),.dout(w_dff_B_qpvjGOiZ6_2),.clk(gclk));
	jdff dff_B_p176txV42_2(.din(w_dff_B_qpvjGOiZ6_2),.dout(w_dff_B_p176txV42_2),.clk(gclk));
	jdff dff_B_yH86lC9q1_2(.din(w_dff_B_p176txV42_2),.dout(w_dff_B_yH86lC9q1_2),.clk(gclk));
	jdff dff_B_VxUcgy9p7_2(.din(w_dff_B_yH86lC9q1_2),.dout(w_dff_B_VxUcgy9p7_2),.clk(gclk));
	jdff dff_B_e1u9NH2T7_2(.din(w_dff_B_VxUcgy9p7_2),.dout(w_dff_B_e1u9NH2T7_2),.clk(gclk));
	jdff dff_B_8ZXWSOco2_2(.din(w_dff_B_e1u9NH2T7_2),.dout(w_dff_B_8ZXWSOco2_2),.clk(gclk));
	jdff dff_B_Yslkd1rH1_2(.din(w_dff_B_8ZXWSOco2_2),.dout(w_dff_B_Yslkd1rH1_2),.clk(gclk));
	jdff dff_B_viwLNiED5_2(.din(w_dff_B_Yslkd1rH1_2),.dout(w_dff_B_viwLNiED5_2),.clk(gclk));
	jdff dff_B_oRVTyjUm3_2(.din(w_dff_B_viwLNiED5_2),.dout(w_dff_B_oRVTyjUm3_2),.clk(gclk));
	jdff dff_B_sOmRu7fn8_2(.din(w_dff_B_oRVTyjUm3_2),.dout(w_dff_B_sOmRu7fn8_2),.clk(gclk));
	jdff dff_B_ImAHvpZZ1_2(.din(w_dff_B_sOmRu7fn8_2),.dout(w_dff_B_ImAHvpZZ1_2),.clk(gclk));
	jdff dff_B_dLpTrMyX5_2(.din(w_dff_B_ImAHvpZZ1_2),.dout(w_dff_B_dLpTrMyX5_2),.clk(gclk));
	jdff dff_B_JtrT2PDz5_2(.din(w_dff_B_dLpTrMyX5_2),.dout(w_dff_B_JtrT2PDz5_2),.clk(gclk));
	jdff dff_B_2lOJk4B49_2(.din(w_dff_B_JtrT2PDz5_2),.dout(w_dff_B_2lOJk4B49_2),.clk(gclk));
	jdff dff_B_nc1ovFbM5_2(.din(w_dff_B_2lOJk4B49_2),.dout(w_dff_B_nc1ovFbM5_2),.clk(gclk));
	jdff dff_B_b28KNNQc0_2(.din(w_dff_B_nc1ovFbM5_2),.dout(w_dff_B_b28KNNQc0_2),.clk(gclk));
	jdff dff_B_JBxP3dqb3_2(.din(w_dff_B_b28KNNQc0_2),.dout(w_dff_B_JBxP3dqb3_2),.clk(gclk));
	jdff dff_B_e12GkItb2_2(.din(w_dff_B_JBxP3dqb3_2),.dout(w_dff_B_e12GkItb2_2),.clk(gclk));
	jdff dff_B_mTGVb2Y87_2(.din(w_dff_B_e12GkItb2_2),.dout(w_dff_B_mTGVb2Y87_2),.clk(gclk));
	jdff dff_B_wRhOut4q0_2(.din(n1401),.dout(w_dff_B_wRhOut4q0_2),.clk(gclk));
	jdff dff_B_HdN6e2QS5_1(.din(n1349),.dout(w_dff_B_HdN6e2QS5_1),.clk(gclk));
	jdff dff_B_cfbh6X9D7_2(.din(n1263),.dout(w_dff_B_cfbh6X9D7_2),.clk(gclk));
	jdff dff_B_pOT4qoYE9_2(.din(w_dff_B_cfbh6X9D7_2),.dout(w_dff_B_pOT4qoYE9_2),.clk(gclk));
	jdff dff_B_rjq7m8fe5_2(.din(w_dff_B_pOT4qoYE9_2),.dout(w_dff_B_rjq7m8fe5_2),.clk(gclk));
	jdff dff_B_MTuFUmnU5_2(.din(w_dff_B_rjq7m8fe5_2),.dout(w_dff_B_MTuFUmnU5_2),.clk(gclk));
	jdff dff_B_wvJP5jEF0_2(.din(w_dff_B_MTuFUmnU5_2),.dout(w_dff_B_wvJP5jEF0_2),.clk(gclk));
	jdff dff_B_Nk7tMNV87_2(.din(w_dff_B_wvJP5jEF0_2),.dout(w_dff_B_Nk7tMNV87_2),.clk(gclk));
	jdff dff_B_F9uI3vXr8_2(.din(w_dff_B_Nk7tMNV87_2),.dout(w_dff_B_F9uI3vXr8_2),.clk(gclk));
	jdff dff_B_9ESwFd571_2(.din(w_dff_B_F9uI3vXr8_2),.dout(w_dff_B_9ESwFd571_2),.clk(gclk));
	jdff dff_B_CTQr98h62_2(.din(w_dff_B_9ESwFd571_2),.dout(w_dff_B_CTQr98h62_2),.clk(gclk));
	jdff dff_B_O6Cj7JoH4_2(.din(w_dff_B_CTQr98h62_2),.dout(w_dff_B_O6Cj7JoH4_2),.clk(gclk));
	jdff dff_B_ynsDrXfz9_2(.din(w_dff_B_O6Cj7JoH4_2),.dout(w_dff_B_ynsDrXfz9_2),.clk(gclk));
	jdff dff_B_Uf3367ra5_2(.din(w_dff_B_ynsDrXfz9_2),.dout(w_dff_B_Uf3367ra5_2),.clk(gclk));
	jdff dff_B_0af13xxu5_2(.din(w_dff_B_Uf3367ra5_2),.dout(w_dff_B_0af13xxu5_2),.clk(gclk));
	jdff dff_B_Kw7vO2ZE4_2(.din(w_dff_B_0af13xxu5_2),.dout(w_dff_B_Kw7vO2ZE4_2),.clk(gclk));
	jdff dff_B_A50lyDmP1_2(.din(w_dff_B_Kw7vO2ZE4_2),.dout(w_dff_B_A50lyDmP1_2),.clk(gclk));
	jdff dff_B_B12yDqG91_2(.din(w_dff_B_A50lyDmP1_2),.dout(w_dff_B_B12yDqG91_2),.clk(gclk));
	jdff dff_B_5uO59pTn4_2(.din(w_dff_B_B12yDqG91_2),.dout(w_dff_B_5uO59pTn4_2),.clk(gclk));
	jdff dff_B_gtldhGR49_2(.din(w_dff_B_5uO59pTn4_2),.dout(w_dff_B_gtldhGR49_2),.clk(gclk));
	jdff dff_B_btLbHQG55_2(.din(w_dff_B_gtldhGR49_2),.dout(w_dff_B_btLbHQG55_2),.clk(gclk));
	jdff dff_B_jdCCI9yg0_2(.din(w_dff_B_btLbHQG55_2),.dout(w_dff_B_jdCCI9yg0_2),.clk(gclk));
	jdff dff_B_b3oEeMNT3_2(.din(w_dff_B_jdCCI9yg0_2),.dout(w_dff_B_b3oEeMNT3_2),.clk(gclk));
	jdff dff_B_rpLcmaKz7_2(.din(w_dff_B_b3oEeMNT3_2),.dout(w_dff_B_rpLcmaKz7_2),.clk(gclk));
	jdff dff_B_GIpjYGQf5_2(.din(w_dff_B_rpLcmaKz7_2),.dout(w_dff_B_GIpjYGQf5_2),.clk(gclk));
	jdff dff_B_4XeTKFQn7_2(.din(w_dff_B_GIpjYGQf5_2),.dout(w_dff_B_4XeTKFQn7_2),.clk(gclk));
	jdff dff_B_v6ceRsv35_2(.din(w_dff_B_4XeTKFQn7_2),.dout(w_dff_B_v6ceRsv35_2),.clk(gclk));
	jdff dff_B_i8lKL3H85_2(.din(w_dff_B_v6ceRsv35_2),.dout(w_dff_B_i8lKL3H85_2),.clk(gclk));
	jdff dff_B_6EyYZzVG6_2(.din(w_dff_B_i8lKL3H85_2),.dout(w_dff_B_6EyYZzVG6_2),.clk(gclk));
	jdff dff_B_zKpleKsM8_2(.din(w_dff_B_6EyYZzVG6_2),.dout(w_dff_B_zKpleKsM8_2),.clk(gclk));
	jdff dff_B_X3hfhygc5_2(.din(w_dff_B_zKpleKsM8_2),.dout(w_dff_B_X3hfhygc5_2),.clk(gclk));
	jdff dff_B_9yGH2G2T3_2(.din(w_dff_B_X3hfhygc5_2),.dout(w_dff_B_9yGH2G2T3_2),.clk(gclk));
	jdff dff_B_rqUVYrVU9_2(.din(w_dff_B_9yGH2G2T3_2),.dout(w_dff_B_rqUVYrVU9_2),.clk(gclk));
	jdff dff_B_HFkZRdSW2_2(.din(w_dff_B_rqUVYrVU9_2),.dout(w_dff_B_HFkZRdSW2_2),.clk(gclk));
	jdff dff_B_hv2AnX7z3_2(.din(w_dff_B_HFkZRdSW2_2),.dout(w_dff_B_hv2AnX7z3_2),.clk(gclk));
	jdff dff_B_djjgwTXb7_2(.din(w_dff_B_hv2AnX7z3_2),.dout(w_dff_B_djjgwTXb7_2),.clk(gclk));
	jdff dff_B_Wx6OaocS6_2(.din(w_dff_B_djjgwTXb7_2),.dout(w_dff_B_Wx6OaocS6_2),.clk(gclk));
	jdff dff_B_LczfR24N0_2(.din(w_dff_B_Wx6OaocS6_2),.dout(w_dff_B_LczfR24N0_2),.clk(gclk));
	jdff dff_B_iqP04Ira2_2(.din(n1316),.dout(w_dff_B_iqP04Ira2_2),.clk(gclk));
	jdff dff_B_z5RhBe3P9_1(.din(n1264),.dout(w_dff_B_z5RhBe3P9_1),.clk(gclk));
	jdff dff_B_ahExX52R0_2(.din(n1173),.dout(w_dff_B_ahExX52R0_2),.clk(gclk));
	jdff dff_B_v1RNsA6J9_2(.din(w_dff_B_ahExX52R0_2),.dout(w_dff_B_v1RNsA6J9_2),.clk(gclk));
	jdff dff_B_cJL8jU797_2(.din(w_dff_B_v1RNsA6J9_2),.dout(w_dff_B_cJL8jU797_2),.clk(gclk));
	jdff dff_B_eA16Gydg5_2(.din(w_dff_B_cJL8jU797_2),.dout(w_dff_B_eA16Gydg5_2),.clk(gclk));
	jdff dff_B_HzZ6NIKZ0_2(.din(w_dff_B_eA16Gydg5_2),.dout(w_dff_B_HzZ6NIKZ0_2),.clk(gclk));
	jdff dff_B_lIS2M8i35_2(.din(w_dff_B_HzZ6NIKZ0_2),.dout(w_dff_B_lIS2M8i35_2),.clk(gclk));
	jdff dff_B_BlvSV2fL8_2(.din(w_dff_B_lIS2M8i35_2),.dout(w_dff_B_BlvSV2fL8_2),.clk(gclk));
	jdff dff_B_IYhS2iSa6_2(.din(w_dff_B_BlvSV2fL8_2),.dout(w_dff_B_IYhS2iSa6_2),.clk(gclk));
	jdff dff_B_amg2TSHd5_2(.din(w_dff_B_IYhS2iSa6_2),.dout(w_dff_B_amg2TSHd5_2),.clk(gclk));
	jdff dff_B_CBRTIi9H5_2(.din(w_dff_B_amg2TSHd5_2),.dout(w_dff_B_CBRTIi9H5_2),.clk(gclk));
	jdff dff_B_9RfQCK361_2(.din(w_dff_B_CBRTIi9H5_2),.dout(w_dff_B_9RfQCK361_2),.clk(gclk));
	jdff dff_B_Y3ycp56H7_2(.din(w_dff_B_9RfQCK361_2),.dout(w_dff_B_Y3ycp56H7_2),.clk(gclk));
	jdff dff_B_UqpjfU9K1_2(.din(w_dff_B_Y3ycp56H7_2),.dout(w_dff_B_UqpjfU9K1_2),.clk(gclk));
	jdff dff_B_WerwZNX65_2(.din(w_dff_B_UqpjfU9K1_2),.dout(w_dff_B_WerwZNX65_2),.clk(gclk));
	jdff dff_B_XIXe867m6_2(.din(w_dff_B_WerwZNX65_2),.dout(w_dff_B_XIXe867m6_2),.clk(gclk));
	jdff dff_B_UiRo5sdd1_2(.din(w_dff_B_XIXe867m6_2),.dout(w_dff_B_UiRo5sdd1_2),.clk(gclk));
	jdff dff_B_NwydGrbz1_2(.din(w_dff_B_UiRo5sdd1_2),.dout(w_dff_B_NwydGrbz1_2),.clk(gclk));
	jdff dff_B_YLDc6gkU2_2(.din(w_dff_B_NwydGrbz1_2),.dout(w_dff_B_YLDc6gkU2_2),.clk(gclk));
	jdff dff_B_2N1Yr9ex1_2(.din(w_dff_B_YLDc6gkU2_2),.dout(w_dff_B_2N1Yr9ex1_2),.clk(gclk));
	jdff dff_B_QXlBy0AW5_2(.din(w_dff_B_2N1Yr9ex1_2),.dout(w_dff_B_QXlBy0AW5_2),.clk(gclk));
	jdff dff_B_P4ZlhUqU8_2(.din(w_dff_B_QXlBy0AW5_2),.dout(w_dff_B_P4ZlhUqU8_2),.clk(gclk));
	jdff dff_B_leDsltOd6_2(.din(w_dff_B_P4ZlhUqU8_2),.dout(w_dff_B_leDsltOd6_2),.clk(gclk));
	jdff dff_B_4oJiMfPy2_2(.din(w_dff_B_leDsltOd6_2),.dout(w_dff_B_4oJiMfPy2_2),.clk(gclk));
	jdff dff_B_SVfCfHwD8_2(.din(w_dff_B_4oJiMfPy2_2),.dout(w_dff_B_SVfCfHwD8_2),.clk(gclk));
	jdff dff_B_q3wKuDe99_2(.din(w_dff_B_SVfCfHwD8_2),.dout(w_dff_B_q3wKuDe99_2),.clk(gclk));
	jdff dff_B_650xjR7n2_2(.din(w_dff_B_q3wKuDe99_2),.dout(w_dff_B_650xjR7n2_2),.clk(gclk));
	jdff dff_B_Slrvo9Ty9_2(.din(w_dff_B_650xjR7n2_2),.dout(w_dff_B_Slrvo9Ty9_2),.clk(gclk));
	jdff dff_B_89vM4sNl6_2(.din(w_dff_B_Slrvo9Ty9_2),.dout(w_dff_B_89vM4sNl6_2),.clk(gclk));
	jdff dff_B_pfgS2cDN7_2(.din(w_dff_B_89vM4sNl6_2),.dout(w_dff_B_pfgS2cDN7_2),.clk(gclk));
	jdff dff_B_7mbIxNWX3_2(.din(w_dff_B_pfgS2cDN7_2),.dout(w_dff_B_7mbIxNWX3_2),.clk(gclk));
	jdff dff_B_xJj2QTNd3_2(.din(w_dff_B_7mbIxNWX3_2),.dout(w_dff_B_xJj2QTNd3_2),.clk(gclk));
	jdff dff_B_V0XZExdl1_2(.din(w_dff_B_xJj2QTNd3_2),.dout(w_dff_B_V0XZExdl1_2),.clk(gclk));
	jdff dff_B_Za3PwOC99_2(.din(w_dff_B_V0XZExdl1_2),.dout(w_dff_B_Za3PwOC99_2),.clk(gclk));
	jdff dff_B_AvICfoV98_2(.din(n1225),.dout(w_dff_B_AvICfoV98_2),.clk(gclk));
	jdff dff_B_gkznpBEf4_1(.din(n1174),.dout(w_dff_B_gkznpBEf4_1),.clk(gclk));
	jdff dff_B_Um5dOghd3_2(.din(n1069),.dout(w_dff_B_Um5dOghd3_2),.clk(gclk));
	jdff dff_B_H9E6PndJ4_2(.din(w_dff_B_Um5dOghd3_2),.dout(w_dff_B_H9E6PndJ4_2),.clk(gclk));
	jdff dff_B_mLYq6oUH3_2(.din(w_dff_B_H9E6PndJ4_2),.dout(w_dff_B_mLYq6oUH3_2),.clk(gclk));
	jdff dff_B_qOMWTWBP5_2(.din(w_dff_B_mLYq6oUH3_2),.dout(w_dff_B_qOMWTWBP5_2),.clk(gclk));
	jdff dff_B_1whUBTFv3_2(.din(w_dff_B_qOMWTWBP5_2),.dout(w_dff_B_1whUBTFv3_2),.clk(gclk));
	jdff dff_B_Mwfq03dg8_2(.din(w_dff_B_1whUBTFv3_2),.dout(w_dff_B_Mwfq03dg8_2),.clk(gclk));
	jdff dff_B_srBU42iG0_2(.din(w_dff_B_Mwfq03dg8_2),.dout(w_dff_B_srBU42iG0_2),.clk(gclk));
	jdff dff_B_AKkFTaAY9_2(.din(w_dff_B_srBU42iG0_2),.dout(w_dff_B_AKkFTaAY9_2),.clk(gclk));
	jdff dff_B_hEVWqqtR3_2(.din(w_dff_B_AKkFTaAY9_2),.dout(w_dff_B_hEVWqqtR3_2),.clk(gclk));
	jdff dff_B_JmZnRLM25_2(.din(w_dff_B_hEVWqqtR3_2),.dout(w_dff_B_JmZnRLM25_2),.clk(gclk));
	jdff dff_B_7jVS0mXv5_2(.din(w_dff_B_JmZnRLM25_2),.dout(w_dff_B_7jVS0mXv5_2),.clk(gclk));
	jdff dff_B_UHmDUxO57_2(.din(w_dff_B_7jVS0mXv5_2),.dout(w_dff_B_UHmDUxO57_2),.clk(gclk));
	jdff dff_B_CjtcbXPy7_2(.din(w_dff_B_UHmDUxO57_2),.dout(w_dff_B_CjtcbXPy7_2),.clk(gclk));
	jdff dff_B_7lY1tv9g5_2(.din(w_dff_B_CjtcbXPy7_2),.dout(w_dff_B_7lY1tv9g5_2),.clk(gclk));
	jdff dff_B_WwvHEjaQ0_2(.din(w_dff_B_7lY1tv9g5_2),.dout(w_dff_B_WwvHEjaQ0_2),.clk(gclk));
	jdff dff_B_snmFQfGG1_2(.din(w_dff_B_WwvHEjaQ0_2),.dout(w_dff_B_snmFQfGG1_2),.clk(gclk));
	jdff dff_B_qyeUTYx37_2(.din(w_dff_B_snmFQfGG1_2),.dout(w_dff_B_qyeUTYx37_2),.clk(gclk));
	jdff dff_B_uW37g5LN3_2(.din(w_dff_B_qyeUTYx37_2),.dout(w_dff_B_uW37g5LN3_2),.clk(gclk));
	jdff dff_B_equ5fY3g1_2(.din(w_dff_B_uW37g5LN3_2),.dout(w_dff_B_equ5fY3g1_2),.clk(gclk));
	jdff dff_B_cdQk5QfP5_2(.din(w_dff_B_equ5fY3g1_2),.dout(w_dff_B_cdQk5QfP5_2),.clk(gclk));
	jdff dff_B_AviJSpvS3_2(.din(w_dff_B_cdQk5QfP5_2),.dout(w_dff_B_AviJSpvS3_2),.clk(gclk));
	jdff dff_B_owY0euqi6_2(.din(w_dff_B_AviJSpvS3_2),.dout(w_dff_B_owY0euqi6_2),.clk(gclk));
	jdff dff_B_yvbmzEOI3_2(.din(w_dff_B_owY0euqi6_2),.dout(w_dff_B_yvbmzEOI3_2),.clk(gclk));
	jdff dff_B_7E72KJj92_2(.din(w_dff_B_yvbmzEOI3_2),.dout(w_dff_B_7E72KJj92_2),.clk(gclk));
	jdff dff_B_vXbupGDE7_2(.din(w_dff_B_7E72KJj92_2),.dout(w_dff_B_vXbupGDE7_2),.clk(gclk));
	jdff dff_B_LiKea8F97_2(.din(w_dff_B_vXbupGDE7_2),.dout(w_dff_B_LiKea8F97_2),.clk(gclk));
	jdff dff_B_X3kIljoC4_2(.din(w_dff_B_LiKea8F97_2),.dout(w_dff_B_X3kIljoC4_2),.clk(gclk));
	jdff dff_B_vRZtnJ3b7_2(.din(w_dff_B_X3kIljoC4_2),.dout(w_dff_B_vRZtnJ3b7_2),.clk(gclk));
	jdff dff_B_dlF8wpcl4_2(.din(w_dff_B_vRZtnJ3b7_2),.dout(w_dff_B_dlF8wpcl4_2),.clk(gclk));
	jdff dff_B_QMuW436K2_2(.din(w_dff_B_dlF8wpcl4_2),.dout(w_dff_B_QMuW436K2_2),.clk(gclk));
	jdff dff_B_tK1POAiv8_2(.din(n1127),.dout(w_dff_B_tK1POAiv8_2),.clk(gclk));
	jdff dff_B_AWEkbpKd1_1(.din(n1070),.dout(w_dff_B_AWEkbpKd1_1),.clk(gclk));
	jdff dff_B_5vBfRpeh4_2(.din(n971),.dout(w_dff_B_5vBfRpeh4_2),.clk(gclk));
	jdff dff_B_M2ILRsz14_2(.din(w_dff_B_5vBfRpeh4_2),.dout(w_dff_B_M2ILRsz14_2),.clk(gclk));
	jdff dff_B_QjrNtuYS3_2(.din(w_dff_B_M2ILRsz14_2),.dout(w_dff_B_QjrNtuYS3_2),.clk(gclk));
	jdff dff_B_kb4jkFpI7_2(.din(w_dff_B_QjrNtuYS3_2),.dout(w_dff_B_kb4jkFpI7_2),.clk(gclk));
	jdff dff_B_1RBGOdJH1_2(.din(w_dff_B_kb4jkFpI7_2),.dout(w_dff_B_1RBGOdJH1_2),.clk(gclk));
	jdff dff_B_enG3Nk1C4_2(.din(w_dff_B_1RBGOdJH1_2),.dout(w_dff_B_enG3Nk1C4_2),.clk(gclk));
	jdff dff_B_9gFfoXFU0_2(.din(w_dff_B_enG3Nk1C4_2),.dout(w_dff_B_9gFfoXFU0_2),.clk(gclk));
	jdff dff_B_ZFHIbfop4_2(.din(w_dff_B_9gFfoXFU0_2),.dout(w_dff_B_ZFHIbfop4_2),.clk(gclk));
	jdff dff_B_8SNUpDdJ0_2(.din(w_dff_B_ZFHIbfop4_2),.dout(w_dff_B_8SNUpDdJ0_2),.clk(gclk));
	jdff dff_B_8EDZHkR78_2(.din(w_dff_B_8SNUpDdJ0_2),.dout(w_dff_B_8EDZHkR78_2),.clk(gclk));
	jdff dff_B_H52xUj512_2(.din(w_dff_B_8EDZHkR78_2),.dout(w_dff_B_H52xUj512_2),.clk(gclk));
	jdff dff_B_Hcx913mr2_2(.din(w_dff_B_H52xUj512_2),.dout(w_dff_B_Hcx913mr2_2),.clk(gclk));
	jdff dff_B_GJBaQ3Y26_2(.din(w_dff_B_Hcx913mr2_2),.dout(w_dff_B_GJBaQ3Y26_2),.clk(gclk));
	jdff dff_B_AXk6Rmex0_2(.din(w_dff_B_GJBaQ3Y26_2),.dout(w_dff_B_AXk6Rmex0_2),.clk(gclk));
	jdff dff_B_tBAQOmxm2_2(.din(w_dff_B_AXk6Rmex0_2),.dout(w_dff_B_tBAQOmxm2_2),.clk(gclk));
	jdff dff_B_JwLdyZUt0_2(.din(w_dff_B_tBAQOmxm2_2),.dout(w_dff_B_JwLdyZUt0_2),.clk(gclk));
	jdff dff_B_2Uys5daT8_2(.din(w_dff_B_JwLdyZUt0_2),.dout(w_dff_B_2Uys5daT8_2),.clk(gclk));
	jdff dff_B_VvDPI0nO7_2(.din(w_dff_B_2Uys5daT8_2),.dout(w_dff_B_VvDPI0nO7_2),.clk(gclk));
	jdff dff_B_QAnNtVyB4_2(.din(w_dff_B_VvDPI0nO7_2),.dout(w_dff_B_QAnNtVyB4_2),.clk(gclk));
	jdff dff_B_fImbjnfv7_2(.din(w_dff_B_QAnNtVyB4_2),.dout(w_dff_B_fImbjnfv7_2),.clk(gclk));
	jdff dff_B_193FPRAe6_2(.din(w_dff_B_fImbjnfv7_2),.dout(w_dff_B_193FPRAe6_2),.clk(gclk));
	jdff dff_B_0XLaWxPT5_2(.din(w_dff_B_193FPRAe6_2),.dout(w_dff_B_0XLaWxPT5_2),.clk(gclk));
	jdff dff_B_gNZp66ua7_2(.din(w_dff_B_0XLaWxPT5_2),.dout(w_dff_B_gNZp66ua7_2),.clk(gclk));
	jdff dff_B_uURC9QOx5_2(.din(w_dff_B_gNZp66ua7_2),.dout(w_dff_B_uURC9QOx5_2),.clk(gclk));
	jdff dff_B_Hywtq1Vt1_2(.din(w_dff_B_uURC9QOx5_2),.dout(w_dff_B_Hywtq1Vt1_2),.clk(gclk));
	jdff dff_B_VUUqCtZM2_2(.din(w_dff_B_Hywtq1Vt1_2),.dout(w_dff_B_VUUqCtZM2_2),.clk(gclk));
	jdff dff_B_MjkJMhHw9_2(.din(w_dff_B_VUUqCtZM2_2),.dout(w_dff_B_MjkJMhHw9_2),.clk(gclk));
	jdff dff_B_BLi57DKT7_2(.din(n1022),.dout(w_dff_B_BLi57DKT7_2),.clk(gclk));
	jdff dff_B_qwmlGLoC7_1(.din(n972),.dout(w_dff_B_qwmlGLoC7_1),.clk(gclk));
	jdff dff_B_euHYX45B4_2(.din(n866),.dout(w_dff_B_euHYX45B4_2),.clk(gclk));
	jdff dff_B_A1z9AQnR1_2(.din(w_dff_B_euHYX45B4_2),.dout(w_dff_B_A1z9AQnR1_2),.clk(gclk));
	jdff dff_B_UejawuOu4_2(.din(w_dff_B_A1z9AQnR1_2),.dout(w_dff_B_UejawuOu4_2),.clk(gclk));
	jdff dff_B_qrnNWu0h4_2(.din(w_dff_B_UejawuOu4_2),.dout(w_dff_B_qrnNWu0h4_2),.clk(gclk));
	jdff dff_B_UN6E8hBU2_2(.din(w_dff_B_qrnNWu0h4_2),.dout(w_dff_B_UN6E8hBU2_2),.clk(gclk));
	jdff dff_B_GZc0UFjg3_2(.din(w_dff_B_UN6E8hBU2_2),.dout(w_dff_B_GZc0UFjg3_2),.clk(gclk));
	jdff dff_B_Sziofqbt8_2(.din(w_dff_B_GZc0UFjg3_2),.dout(w_dff_B_Sziofqbt8_2),.clk(gclk));
	jdff dff_B_wP0DZBgY8_2(.din(w_dff_B_Sziofqbt8_2),.dout(w_dff_B_wP0DZBgY8_2),.clk(gclk));
	jdff dff_B_yLXbKVKd0_2(.din(w_dff_B_wP0DZBgY8_2),.dout(w_dff_B_yLXbKVKd0_2),.clk(gclk));
	jdff dff_B_b3WXyUQe3_2(.din(w_dff_B_yLXbKVKd0_2),.dout(w_dff_B_b3WXyUQe3_2),.clk(gclk));
	jdff dff_B_sK9bpa6M6_2(.din(w_dff_B_b3WXyUQe3_2),.dout(w_dff_B_sK9bpa6M6_2),.clk(gclk));
	jdff dff_B_eQWzRKi33_2(.din(w_dff_B_sK9bpa6M6_2),.dout(w_dff_B_eQWzRKi33_2),.clk(gclk));
	jdff dff_B_P6aWvTaA8_2(.din(w_dff_B_eQWzRKi33_2),.dout(w_dff_B_P6aWvTaA8_2),.clk(gclk));
	jdff dff_B_qZmgXeD04_2(.din(w_dff_B_P6aWvTaA8_2),.dout(w_dff_B_qZmgXeD04_2),.clk(gclk));
	jdff dff_B_rPhT8Vtk6_2(.din(w_dff_B_qZmgXeD04_2),.dout(w_dff_B_rPhT8Vtk6_2),.clk(gclk));
	jdff dff_B_LNrPLZp47_2(.din(w_dff_B_rPhT8Vtk6_2),.dout(w_dff_B_LNrPLZp47_2),.clk(gclk));
	jdff dff_B_tgrg1QM66_2(.din(w_dff_B_LNrPLZp47_2),.dout(w_dff_B_tgrg1QM66_2),.clk(gclk));
	jdff dff_B_PokZ6lb99_2(.din(w_dff_B_tgrg1QM66_2),.dout(w_dff_B_PokZ6lb99_2),.clk(gclk));
	jdff dff_B_1EwewgJP1_2(.din(w_dff_B_PokZ6lb99_2),.dout(w_dff_B_1EwewgJP1_2),.clk(gclk));
	jdff dff_B_rrtrXJzX3_2(.din(w_dff_B_1EwewgJP1_2),.dout(w_dff_B_rrtrXJzX3_2),.clk(gclk));
	jdff dff_B_pzAnSdtX1_2(.din(w_dff_B_rrtrXJzX3_2),.dout(w_dff_B_pzAnSdtX1_2),.clk(gclk));
	jdff dff_B_UABLJ9ch4_2(.din(w_dff_B_pzAnSdtX1_2),.dout(w_dff_B_UABLJ9ch4_2),.clk(gclk));
	jdff dff_B_hWnCGiGP0_2(.din(w_dff_B_UABLJ9ch4_2),.dout(w_dff_B_hWnCGiGP0_2),.clk(gclk));
	jdff dff_B_Iell99iK5_2(.din(w_dff_B_hWnCGiGP0_2),.dout(w_dff_B_Iell99iK5_2),.clk(gclk));
	jdff dff_B_fIPyYPm37_2(.din(n917),.dout(w_dff_B_fIPyYPm37_2),.clk(gclk));
	jdff dff_B_5qkz8cg51_1(.din(n867),.dout(w_dff_B_5qkz8cg51_1),.clk(gclk));
	jdff dff_B_BoEwLXE98_2(.din(n767),.dout(w_dff_B_BoEwLXE98_2),.clk(gclk));
	jdff dff_B_s3DLjG1M5_2(.din(w_dff_B_BoEwLXE98_2),.dout(w_dff_B_s3DLjG1M5_2),.clk(gclk));
	jdff dff_B_72R1pmrG2_2(.din(w_dff_B_s3DLjG1M5_2),.dout(w_dff_B_72R1pmrG2_2),.clk(gclk));
	jdff dff_B_N8CUq8oI7_2(.din(w_dff_B_72R1pmrG2_2),.dout(w_dff_B_N8CUq8oI7_2),.clk(gclk));
	jdff dff_B_ZrPzR4LO1_2(.din(w_dff_B_N8CUq8oI7_2),.dout(w_dff_B_ZrPzR4LO1_2),.clk(gclk));
	jdff dff_B_zOVgel6M8_2(.din(w_dff_B_ZrPzR4LO1_2),.dout(w_dff_B_zOVgel6M8_2),.clk(gclk));
	jdff dff_B_ooH9eEDJ8_2(.din(w_dff_B_zOVgel6M8_2),.dout(w_dff_B_ooH9eEDJ8_2),.clk(gclk));
	jdff dff_B_prHYvDcF8_2(.din(w_dff_B_ooH9eEDJ8_2),.dout(w_dff_B_prHYvDcF8_2),.clk(gclk));
	jdff dff_B_LoJzzz282_2(.din(w_dff_B_prHYvDcF8_2),.dout(w_dff_B_LoJzzz282_2),.clk(gclk));
	jdff dff_B_KG9YTMnp0_2(.din(w_dff_B_LoJzzz282_2),.dout(w_dff_B_KG9YTMnp0_2),.clk(gclk));
	jdff dff_B_NPG4eW0u9_2(.din(w_dff_B_KG9YTMnp0_2),.dout(w_dff_B_NPG4eW0u9_2),.clk(gclk));
	jdff dff_B_sr5SH9mf4_2(.din(w_dff_B_NPG4eW0u9_2),.dout(w_dff_B_sr5SH9mf4_2),.clk(gclk));
	jdff dff_B_PYtNlISA0_2(.din(w_dff_B_sr5SH9mf4_2),.dout(w_dff_B_PYtNlISA0_2),.clk(gclk));
	jdff dff_B_2noJLMqk7_2(.din(w_dff_B_PYtNlISA0_2),.dout(w_dff_B_2noJLMqk7_2),.clk(gclk));
	jdff dff_B_9NFdoTIe5_2(.din(w_dff_B_2noJLMqk7_2),.dout(w_dff_B_9NFdoTIe5_2),.clk(gclk));
	jdff dff_B_Y3j9pDfy8_2(.din(w_dff_B_9NFdoTIe5_2),.dout(w_dff_B_Y3j9pDfy8_2),.clk(gclk));
	jdff dff_B_kPVOvwrw1_2(.din(w_dff_B_Y3j9pDfy8_2),.dout(w_dff_B_kPVOvwrw1_2),.clk(gclk));
	jdff dff_B_D2eo2n0s1_2(.din(w_dff_B_kPVOvwrw1_2),.dout(w_dff_B_D2eo2n0s1_2),.clk(gclk));
	jdff dff_B_jpcMik465_2(.din(w_dff_B_D2eo2n0s1_2),.dout(w_dff_B_jpcMik465_2),.clk(gclk));
	jdff dff_B_Paijxd6A3_2(.din(w_dff_B_jpcMik465_2),.dout(w_dff_B_Paijxd6A3_2),.clk(gclk));
	jdff dff_B_Z8L1CnUT9_2(.din(w_dff_B_Paijxd6A3_2),.dout(w_dff_B_Z8L1CnUT9_2),.clk(gclk));
	jdff dff_B_WSBkRGqV8_2(.din(n811),.dout(w_dff_B_WSBkRGqV8_2),.clk(gclk));
	jdff dff_B_at4LAabB1_1(.din(n768),.dout(w_dff_B_at4LAabB1_1),.clk(gclk));
	jdff dff_B_xm9sL97L3_2(.din(n674),.dout(w_dff_B_xm9sL97L3_2),.clk(gclk));
	jdff dff_B_IJM3OSEj6_2(.din(w_dff_B_xm9sL97L3_2),.dout(w_dff_B_IJM3OSEj6_2),.clk(gclk));
	jdff dff_B_UaIeGqz83_2(.din(w_dff_B_IJM3OSEj6_2),.dout(w_dff_B_UaIeGqz83_2),.clk(gclk));
	jdff dff_B_2PDd1dUx3_2(.din(w_dff_B_UaIeGqz83_2),.dout(w_dff_B_2PDd1dUx3_2),.clk(gclk));
	jdff dff_B_diK9KQf09_2(.din(w_dff_B_2PDd1dUx3_2),.dout(w_dff_B_diK9KQf09_2),.clk(gclk));
	jdff dff_B_CgqCN6Ob6_2(.din(w_dff_B_diK9KQf09_2),.dout(w_dff_B_CgqCN6Ob6_2),.clk(gclk));
	jdff dff_B_yrbs7l8d4_2(.din(w_dff_B_CgqCN6Ob6_2),.dout(w_dff_B_yrbs7l8d4_2),.clk(gclk));
	jdff dff_B_apjji1UT0_2(.din(w_dff_B_yrbs7l8d4_2),.dout(w_dff_B_apjji1UT0_2),.clk(gclk));
	jdff dff_B_ek5MbE8t4_2(.din(w_dff_B_apjji1UT0_2),.dout(w_dff_B_ek5MbE8t4_2),.clk(gclk));
	jdff dff_B_A8GwERoR6_2(.din(w_dff_B_ek5MbE8t4_2),.dout(w_dff_B_A8GwERoR6_2),.clk(gclk));
	jdff dff_B_llqUQRuw1_2(.din(w_dff_B_A8GwERoR6_2),.dout(w_dff_B_llqUQRuw1_2),.clk(gclk));
	jdff dff_B_RoFBmCux9_2(.din(w_dff_B_llqUQRuw1_2),.dout(w_dff_B_RoFBmCux9_2),.clk(gclk));
	jdff dff_B_B8SSFgt11_2(.din(w_dff_B_RoFBmCux9_2),.dout(w_dff_B_B8SSFgt11_2),.clk(gclk));
	jdff dff_B_h79TveDr7_2(.din(w_dff_B_B8SSFgt11_2),.dout(w_dff_B_h79TveDr7_2),.clk(gclk));
	jdff dff_B_XsGsk21n0_2(.din(w_dff_B_h79TveDr7_2),.dout(w_dff_B_XsGsk21n0_2),.clk(gclk));
	jdff dff_B_Hi2RD2N60_2(.din(w_dff_B_XsGsk21n0_2),.dout(w_dff_B_Hi2RD2N60_2),.clk(gclk));
	jdff dff_B_wFOIOPRv5_2(.din(w_dff_B_Hi2RD2N60_2),.dout(w_dff_B_wFOIOPRv5_2),.clk(gclk));
	jdff dff_B_hsU6ID7L5_2(.din(w_dff_B_wFOIOPRv5_2),.dout(w_dff_B_hsU6ID7L5_2),.clk(gclk));
	jdff dff_B_wuzspgXl2_2(.din(n711),.dout(w_dff_B_wuzspgXl2_2),.clk(gclk));
	jdff dff_B_7p28RDIn2_1(.din(n675),.dout(w_dff_B_7p28RDIn2_1),.clk(gclk));
	jdff dff_B_IvhAtpny5_2(.din(n588),.dout(w_dff_B_IvhAtpny5_2),.clk(gclk));
	jdff dff_B_ntUjpUV23_2(.din(w_dff_B_IvhAtpny5_2),.dout(w_dff_B_ntUjpUV23_2),.clk(gclk));
	jdff dff_B_aXQJ4Nol2_2(.din(w_dff_B_ntUjpUV23_2),.dout(w_dff_B_aXQJ4Nol2_2),.clk(gclk));
	jdff dff_B_F6eAuYKZ0_2(.din(w_dff_B_aXQJ4Nol2_2),.dout(w_dff_B_F6eAuYKZ0_2),.clk(gclk));
	jdff dff_B_Udhy0t6J0_2(.din(w_dff_B_F6eAuYKZ0_2),.dout(w_dff_B_Udhy0t6J0_2),.clk(gclk));
	jdff dff_B_lmWiHY131_2(.din(w_dff_B_Udhy0t6J0_2),.dout(w_dff_B_lmWiHY131_2),.clk(gclk));
	jdff dff_B_OvqtrIH24_2(.din(w_dff_B_lmWiHY131_2),.dout(w_dff_B_OvqtrIH24_2),.clk(gclk));
	jdff dff_B_Ai7eka4U2_2(.din(w_dff_B_OvqtrIH24_2),.dout(w_dff_B_Ai7eka4U2_2),.clk(gclk));
	jdff dff_B_iLaE0e8Z1_2(.din(w_dff_B_Ai7eka4U2_2),.dout(w_dff_B_iLaE0e8Z1_2),.clk(gclk));
	jdff dff_B_Inh5uVQS7_2(.din(w_dff_B_iLaE0e8Z1_2),.dout(w_dff_B_Inh5uVQS7_2),.clk(gclk));
	jdff dff_B_EMq02nqV4_2(.din(w_dff_B_Inh5uVQS7_2),.dout(w_dff_B_EMq02nqV4_2),.clk(gclk));
	jdff dff_B_KFImtiDl6_2(.din(w_dff_B_EMq02nqV4_2),.dout(w_dff_B_KFImtiDl6_2),.clk(gclk));
	jdff dff_B_tSfP3CgY5_2(.din(w_dff_B_KFImtiDl6_2),.dout(w_dff_B_tSfP3CgY5_2),.clk(gclk));
	jdff dff_B_UlTiNIbn1_2(.din(w_dff_B_tSfP3CgY5_2),.dout(w_dff_B_UlTiNIbn1_2),.clk(gclk));
	jdff dff_B_KZqUSP9O5_2(.din(w_dff_B_UlTiNIbn1_2),.dout(w_dff_B_KZqUSP9O5_2),.clk(gclk));
	jdff dff_B_Y2egNx893_2(.din(n618),.dout(w_dff_B_Y2egNx893_2),.clk(gclk));
	jdff dff_B_31QFqtey6_1(.din(n589),.dout(w_dff_B_31QFqtey6_1),.clk(gclk));
	jdff dff_B_vP52Pb2a6_2(.din(n509),.dout(w_dff_B_vP52Pb2a6_2),.clk(gclk));
	jdff dff_B_1t8bvtjs3_2(.din(w_dff_B_vP52Pb2a6_2),.dout(w_dff_B_1t8bvtjs3_2),.clk(gclk));
	jdff dff_B_NrlT1bAy1_2(.din(w_dff_B_1t8bvtjs3_2),.dout(w_dff_B_NrlT1bAy1_2),.clk(gclk));
	jdff dff_B_Z9SNXE2q4_2(.din(w_dff_B_NrlT1bAy1_2),.dout(w_dff_B_Z9SNXE2q4_2),.clk(gclk));
	jdff dff_B_WKUyCBj38_2(.din(w_dff_B_Z9SNXE2q4_2),.dout(w_dff_B_WKUyCBj38_2),.clk(gclk));
	jdff dff_B_LB8L9Yvo7_2(.din(w_dff_B_WKUyCBj38_2),.dout(w_dff_B_LB8L9Yvo7_2),.clk(gclk));
	jdff dff_B_p2RIrWX56_2(.din(w_dff_B_LB8L9Yvo7_2),.dout(w_dff_B_p2RIrWX56_2),.clk(gclk));
	jdff dff_B_pNC0CmEc3_2(.din(w_dff_B_p2RIrWX56_2),.dout(w_dff_B_pNC0CmEc3_2),.clk(gclk));
	jdff dff_B_RyrqkUYe9_2(.din(w_dff_B_pNC0CmEc3_2),.dout(w_dff_B_RyrqkUYe9_2),.clk(gclk));
	jdff dff_B_zCXSiF3q7_2(.din(w_dff_B_RyrqkUYe9_2),.dout(w_dff_B_zCXSiF3q7_2),.clk(gclk));
	jdff dff_B_kAILsstx7_2(.din(w_dff_B_zCXSiF3q7_2),.dout(w_dff_B_kAILsstx7_2),.clk(gclk));
	jdff dff_B_c848xsSQ9_2(.din(w_dff_B_kAILsstx7_2),.dout(w_dff_B_c848xsSQ9_2),.clk(gclk));
	jdff dff_B_upS3G5Yz1_2(.din(n532),.dout(w_dff_B_upS3G5Yz1_2),.clk(gclk));
	jdff dff_B_d1adPsZB7_1(.din(n510),.dout(w_dff_B_d1adPsZB7_1),.clk(gclk));
	jdff dff_B_fw470LLj2_2(.din(n437),.dout(w_dff_B_fw470LLj2_2),.clk(gclk));
	jdff dff_B_6EfH1EH60_2(.din(w_dff_B_fw470LLj2_2),.dout(w_dff_B_6EfH1EH60_2),.clk(gclk));
	jdff dff_B_9WPp3wtB4_2(.din(w_dff_B_6EfH1EH60_2),.dout(w_dff_B_9WPp3wtB4_2),.clk(gclk));
	jdff dff_B_g4yDPvSI4_2(.din(w_dff_B_9WPp3wtB4_2),.dout(w_dff_B_g4yDPvSI4_2),.clk(gclk));
	jdff dff_B_6ZYf0Wku2_2(.din(w_dff_B_g4yDPvSI4_2),.dout(w_dff_B_6ZYf0Wku2_2),.clk(gclk));
	jdff dff_B_nTiI5cAn6_2(.din(w_dff_B_6ZYf0Wku2_2),.dout(w_dff_B_nTiI5cAn6_2),.clk(gclk));
	jdff dff_B_RKafCkak1_2(.din(w_dff_B_nTiI5cAn6_2),.dout(w_dff_B_RKafCkak1_2),.clk(gclk));
	jdff dff_B_qYiD3Cj93_2(.din(w_dff_B_RKafCkak1_2),.dout(w_dff_B_qYiD3Cj93_2),.clk(gclk));
	jdff dff_B_mJYNJxgE9_2(.din(w_dff_B_qYiD3Cj93_2),.dout(w_dff_B_mJYNJxgE9_2),.clk(gclk));
	jdff dff_B_hguGGLuJ8_2(.din(n453),.dout(w_dff_B_hguGGLuJ8_2),.clk(gclk));
	jdff dff_B_pOhTzdCH3_2(.din(w_dff_B_hguGGLuJ8_2),.dout(w_dff_B_pOhTzdCH3_2),.clk(gclk));
	jdff dff_B_oo7D6KYu1_1(.din(n438),.dout(w_dff_B_oo7D6KYu1_1),.clk(gclk));
	jdff dff_B_sjyUoo7r6_1(.din(w_dff_B_oo7D6KYu1_1),.dout(w_dff_B_sjyUoo7r6_1),.clk(gclk));
	jdff dff_B_miAtFRV98_1(.din(w_dff_B_sjyUoo7r6_1),.dout(w_dff_B_miAtFRV98_1),.clk(gclk));
	jdff dff_B_8EBzYBeb4_1(.din(w_dff_B_miAtFRV98_1),.dout(w_dff_B_8EBzYBeb4_1),.clk(gclk));
	jdff dff_B_NQ3EdVAi2_1(.din(w_dff_B_8EBzYBeb4_1),.dout(w_dff_B_NQ3EdVAi2_1),.clk(gclk));
	jdff dff_B_Un0ukGf28_1(.din(w_dff_B_NQ3EdVAi2_1),.dout(w_dff_B_Un0ukGf28_1),.clk(gclk));
	jdff dff_B_WX9qKg549_0(.din(n381),.dout(w_dff_B_WX9qKg549_0),.clk(gclk));
	jdff dff_B_4BpUftWB8_0(.din(w_dff_B_WX9qKg549_0),.dout(w_dff_B_4BpUftWB8_0),.clk(gclk));
	jdff dff_A_l59cnuZg1_0(.dout(w_n380_0[0]),.din(w_dff_A_l59cnuZg1_0),.clk(gclk));
	jdff dff_A_kSDZ4KsA5_0(.dout(w_dff_A_l59cnuZg1_0),.din(w_dff_A_kSDZ4KsA5_0),.clk(gclk));
	jdff dff_A_FNgLIZwm6_0(.dout(w_dff_A_kSDZ4KsA5_0),.din(w_dff_A_FNgLIZwm6_0),.clk(gclk));
	jdff dff_B_qmu8Bjy34_1(.din(n374),.dout(w_dff_B_qmu8Bjy34_1),.clk(gclk));
	jdff dff_A_BCYGFEtJ4_0(.dout(w_n314_0[0]),.din(w_dff_A_BCYGFEtJ4_0),.clk(gclk));
	jdff dff_A_XTS216BY7_1(.dout(w_n314_0[1]),.din(w_dff_A_XTS216BY7_1),.clk(gclk));
	jdff dff_A_TShp7RaZ3_1(.dout(w_dff_A_XTS216BY7_1),.din(w_dff_A_TShp7RaZ3_1),.clk(gclk));
	jdff dff_A_xGyqHUB36_1(.dout(w_n372_0[1]),.din(w_dff_A_xGyqHUB36_1),.clk(gclk));
	jdff dff_A_gzqnjVnz3_1(.dout(w_dff_A_xGyqHUB36_1),.din(w_dff_A_gzqnjVnz3_1),.clk(gclk));
	jdff dff_A_vBbfU2UW7_1(.dout(w_dff_A_gzqnjVnz3_1),.din(w_dff_A_vBbfU2UW7_1),.clk(gclk));
	jdff dff_A_Fin152cb7_1(.dout(w_dff_A_vBbfU2UW7_1),.din(w_dff_A_Fin152cb7_1),.clk(gclk));
	jdff dff_A_AIO1wok05_1(.dout(w_dff_A_Fin152cb7_1),.din(w_dff_A_AIO1wok05_1),.clk(gclk));
	jdff dff_A_Fn4KLys41_1(.dout(w_dff_A_AIO1wok05_1),.din(w_dff_A_Fn4KLys41_1),.clk(gclk));
	jdff dff_B_SRfgufy24_2(.din(n1627),.dout(w_dff_B_SRfgufy24_2),.clk(gclk));
	jdff dff_B_eA7aoaMJ9_2(.din(w_dff_B_SRfgufy24_2),.dout(w_dff_B_eA7aoaMJ9_2),.clk(gclk));
	jdff dff_B_sOht3dtF1_1(.din(n1625),.dout(w_dff_B_sOht3dtF1_1),.clk(gclk));
	jdff dff_B_7UQ2vDpt1_2(.din(n1566),.dout(w_dff_B_7UQ2vDpt1_2),.clk(gclk));
	jdff dff_B_huhSvj3r8_2(.din(w_dff_B_7UQ2vDpt1_2),.dout(w_dff_B_huhSvj3r8_2),.clk(gclk));
	jdff dff_B_871pwHoW0_2(.din(w_dff_B_huhSvj3r8_2),.dout(w_dff_B_871pwHoW0_2),.clk(gclk));
	jdff dff_B_S5GWN62B7_2(.din(w_dff_B_871pwHoW0_2),.dout(w_dff_B_S5GWN62B7_2),.clk(gclk));
	jdff dff_B_r78LakDc8_2(.din(w_dff_B_S5GWN62B7_2),.dout(w_dff_B_r78LakDc8_2),.clk(gclk));
	jdff dff_B_tBkInLPj6_2(.din(w_dff_B_r78LakDc8_2),.dout(w_dff_B_tBkInLPj6_2),.clk(gclk));
	jdff dff_B_XONPbD7x5_2(.din(w_dff_B_tBkInLPj6_2),.dout(w_dff_B_XONPbD7x5_2),.clk(gclk));
	jdff dff_B_xk9jNLee5_2(.din(w_dff_B_XONPbD7x5_2),.dout(w_dff_B_xk9jNLee5_2),.clk(gclk));
	jdff dff_B_h78Cr5E01_2(.din(w_dff_B_xk9jNLee5_2),.dout(w_dff_B_h78Cr5E01_2),.clk(gclk));
	jdff dff_B_qwMZolfl7_2(.din(w_dff_B_h78Cr5E01_2),.dout(w_dff_B_qwMZolfl7_2),.clk(gclk));
	jdff dff_B_jB0rlgym9_2(.din(w_dff_B_qwMZolfl7_2),.dout(w_dff_B_jB0rlgym9_2),.clk(gclk));
	jdff dff_B_PDPXy9p86_2(.din(w_dff_B_jB0rlgym9_2),.dout(w_dff_B_PDPXy9p86_2),.clk(gclk));
	jdff dff_B_IMQ55Fku5_2(.din(w_dff_B_PDPXy9p86_2),.dout(w_dff_B_IMQ55Fku5_2),.clk(gclk));
	jdff dff_B_FqKH4nCt2_2(.din(w_dff_B_IMQ55Fku5_2),.dout(w_dff_B_FqKH4nCt2_2),.clk(gclk));
	jdff dff_B_LSj3fhoK4_2(.din(w_dff_B_FqKH4nCt2_2),.dout(w_dff_B_LSj3fhoK4_2),.clk(gclk));
	jdff dff_B_oLxYCPow6_2(.din(w_dff_B_LSj3fhoK4_2),.dout(w_dff_B_oLxYCPow6_2),.clk(gclk));
	jdff dff_B_LRzd3Ust8_2(.din(w_dff_B_oLxYCPow6_2),.dout(w_dff_B_LRzd3Ust8_2),.clk(gclk));
	jdff dff_B_38XKmR9x9_2(.din(w_dff_B_LRzd3Ust8_2),.dout(w_dff_B_38XKmR9x9_2),.clk(gclk));
	jdff dff_B_7aqk4jRV4_2(.din(w_dff_B_38XKmR9x9_2),.dout(w_dff_B_7aqk4jRV4_2),.clk(gclk));
	jdff dff_B_zkkDv3E37_2(.din(w_dff_B_7aqk4jRV4_2),.dout(w_dff_B_zkkDv3E37_2),.clk(gclk));
	jdff dff_B_MdZXwrO87_2(.din(w_dff_B_zkkDv3E37_2),.dout(w_dff_B_MdZXwrO87_2),.clk(gclk));
	jdff dff_B_RWiWCDx43_2(.din(w_dff_B_MdZXwrO87_2),.dout(w_dff_B_RWiWCDx43_2),.clk(gclk));
	jdff dff_B_pfZ4jjN22_2(.din(w_dff_B_RWiWCDx43_2),.dout(w_dff_B_pfZ4jjN22_2),.clk(gclk));
	jdff dff_B_5yxv7tkq0_2(.din(w_dff_B_pfZ4jjN22_2),.dout(w_dff_B_5yxv7tkq0_2),.clk(gclk));
	jdff dff_B_iI5Wie4t2_2(.din(w_dff_B_5yxv7tkq0_2),.dout(w_dff_B_iI5Wie4t2_2),.clk(gclk));
	jdff dff_B_W5IwKxo92_2(.din(w_dff_B_iI5Wie4t2_2),.dout(w_dff_B_W5IwKxo92_2),.clk(gclk));
	jdff dff_B_xhY1LQaj5_2(.din(w_dff_B_W5IwKxo92_2),.dout(w_dff_B_xhY1LQaj5_2),.clk(gclk));
	jdff dff_B_lCgs9Int7_2(.din(w_dff_B_xhY1LQaj5_2),.dout(w_dff_B_lCgs9Int7_2),.clk(gclk));
	jdff dff_B_jUamT2Mz3_2(.din(w_dff_B_lCgs9Int7_2),.dout(w_dff_B_jUamT2Mz3_2),.clk(gclk));
	jdff dff_B_UQbfboNu6_2(.din(w_dff_B_jUamT2Mz3_2),.dout(w_dff_B_UQbfboNu6_2),.clk(gclk));
	jdff dff_B_hPou34aI7_2(.din(w_dff_B_UQbfboNu6_2),.dout(w_dff_B_hPou34aI7_2),.clk(gclk));
	jdff dff_B_hwJ0obT02_2(.din(w_dff_B_hPou34aI7_2),.dout(w_dff_B_hwJ0obT02_2),.clk(gclk));
	jdff dff_B_2AQTaIZL4_2(.din(w_dff_B_hwJ0obT02_2),.dout(w_dff_B_2AQTaIZL4_2),.clk(gclk));
	jdff dff_B_0kuy7kFZ9_2(.din(w_dff_B_2AQTaIZL4_2),.dout(w_dff_B_0kuy7kFZ9_2),.clk(gclk));
	jdff dff_B_Z6HkTEQZ8_2(.din(w_dff_B_0kuy7kFZ9_2),.dout(w_dff_B_Z6HkTEQZ8_2),.clk(gclk));
	jdff dff_B_8aMgngwz9_2(.din(w_dff_B_Z6HkTEQZ8_2),.dout(w_dff_B_8aMgngwz9_2),.clk(gclk));
	jdff dff_B_rvc7jwsb6_2(.din(w_dff_B_8aMgngwz9_2),.dout(w_dff_B_rvc7jwsb6_2),.clk(gclk));
	jdff dff_B_oGK8bSH33_2(.din(w_dff_B_rvc7jwsb6_2),.dout(w_dff_B_oGK8bSH33_2),.clk(gclk));
	jdff dff_B_InQRtAr46_2(.din(w_dff_B_oGK8bSH33_2),.dout(w_dff_B_InQRtAr46_2),.clk(gclk));
	jdff dff_B_QnJnjJhi7_2(.din(w_dff_B_InQRtAr46_2),.dout(w_dff_B_QnJnjJhi7_2),.clk(gclk));
	jdff dff_B_QuMjzmJb6_2(.din(w_dff_B_QnJnjJhi7_2),.dout(w_dff_B_QuMjzmJb6_2),.clk(gclk));
	jdff dff_B_HpTYzOoU6_2(.din(w_dff_B_QuMjzmJb6_2),.dout(w_dff_B_HpTYzOoU6_2),.clk(gclk));
	jdff dff_B_tnFkS6LD3_2(.din(w_dff_B_HpTYzOoU6_2),.dout(w_dff_B_tnFkS6LD3_2),.clk(gclk));
	jdff dff_B_7nSIKhlr0_2(.din(w_dff_B_tnFkS6LD3_2),.dout(w_dff_B_7nSIKhlr0_2),.clk(gclk));
	jdff dff_B_H5P1Ru7E9_2(.din(w_dff_B_7nSIKhlr0_2),.dout(w_dff_B_H5P1Ru7E9_2),.clk(gclk));
	jdff dff_B_x57F2QSf8_2(.din(w_dff_B_H5P1Ru7E9_2),.dout(w_dff_B_x57F2QSf8_2),.clk(gclk));
	jdff dff_B_NFOVWNVB8_2(.din(w_dff_B_x57F2QSf8_2),.dout(w_dff_B_NFOVWNVB8_2),.clk(gclk));
	jdff dff_B_rwbfXufI7_1(.din(n1567),.dout(w_dff_B_rwbfXufI7_1),.clk(gclk));
	jdff dff_B_Mvf2yZgD3_2(.din(n1502),.dout(w_dff_B_Mvf2yZgD3_2),.clk(gclk));
	jdff dff_B_pQvDS6CJ8_2(.din(w_dff_B_Mvf2yZgD3_2),.dout(w_dff_B_pQvDS6CJ8_2),.clk(gclk));
	jdff dff_B_9isAehT03_2(.din(w_dff_B_pQvDS6CJ8_2),.dout(w_dff_B_9isAehT03_2),.clk(gclk));
	jdff dff_B_NPzyMXyw8_2(.din(w_dff_B_9isAehT03_2),.dout(w_dff_B_NPzyMXyw8_2),.clk(gclk));
	jdff dff_B_JDaUb3UT0_2(.din(w_dff_B_NPzyMXyw8_2),.dout(w_dff_B_JDaUb3UT0_2),.clk(gclk));
	jdff dff_B_4HkQPYwG4_2(.din(w_dff_B_JDaUb3UT0_2),.dout(w_dff_B_4HkQPYwG4_2),.clk(gclk));
	jdff dff_B_wUAZFx8i3_2(.din(w_dff_B_4HkQPYwG4_2),.dout(w_dff_B_wUAZFx8i3_2),.clk(gclk));
	jdff dff_B_kqgyDSbB7_2(.din(w_dff_B_wUAZFx8i3_2),.dout(w_dff_B_kqgyDSbB7_2),.clk(gclk));
	jdff dff_B_WBU4xJDb6_2(.din(w_dff_B_kqgyDSbB7_2),.dout(w_dff_B_WBU4xJDb6_2),.clk(gclk));
	jdff dff_B_Txeyitlz0_2(.din(w_dff_B_WBU4xJDb6_2),.dout(w_dff_B_Txeyitlz0_2),.clk(gclk));
	jdff dff_B_3gEGxFem4_2(.din(w_dff_B_Txeyitlz0_2),.dout(w_dff_B_3gEGxFem4_2),.clk(gclk));
	jdff dff_B_GagQk1B23_2(.din(w_dff_B_3gEGxFem4_2),.dout(w_dff_B_GagQk1B23_2),.clk(gclk));
	jdff dff_B_K9MDhRgH9_2(.din(w_dff_B_GagQk1B23_2),.dout(w_dff_B_K9MDhRgH9_2),.clk(gclk));
	jdff dff_B_bVpb0vZx3_2(.din(w_dff_B_K9MDhRgH9_2),.dout(w_dff_B_bVpb0vZx3_2),.clk(gclk));
	jdff dff_B_ysoCoTuV6_2(.din(w_dff_B_bVpb0vZx3_2),.dout(w_dff_B_ysoCoTuV6_2),.clk(gclk));
	jdff dff_B_CjHb5NVu2_2(.din(w_dff_B_ysoCoTuV6_2),.dout(w_dff_B_CjHb5NVu2_2),.clk(gclk));
	jdff dff_B_zbeL8hEc1_2(.din(w_dff_B_CjHb5NVu2_2),.dout(w_dff_B_zbeL8hEc1_2),.clk(gclk));
	jdff dff_B_FqnPh0Ac3_2(.din(w_dff_B_zbeL8hEc1_2),.dout(w_dff_B_FqnPh0Ac3_2),.clk(gclk));
	jdff dff_B_mEzzAhU84_2(.din(w_dff_B_FqnPh0Ac3_2),.dout(w_dff_B_mEzzAhU84_2),.clk(gclk));
	jdff dff_B_DHNhYu8h6_2(.din(w_dff_B_mEzzAhU84_2),.dout(w_dff_B_DHNhYu8h6_2),.clk(gclk));
	jdff dff_B_jIlodVVD3_2(.din(w_dff_B_DHNhYu8h6_2),.dout(w_dff_B_jIlodVVD3_2),.clk(gclk));
	jdff dff_B_NQEFVnjF8_2(.din(w_dff_B_jIlodVVD3_2),.dout(w_dff_B_NQEFVnjF8_2),.clk(gclk));
	jdff dff_B_vXDTy26G7_2(.din(w_dff_B_NQEFVnjF8_2),.dout(w_dff_B_vXDTy26G7_2),.clk(gclk));
	jdff dff_B_f3ccBAjS1_2(.din(w_dff_B_vXDTy26G7_2),.dout(w_dff_B_f3ccBAjS1_2),.clk(gclk));
	jdff dff_B_DWNrcmau4_2(.din(w_dff_B_f3ccBAjS1_2),.dout(w_dff_B_DWNrcmau4_2),.clk(gclk));
	jdff dff_B_GNGYj2926_2(.din(w_dff_B_DWNrcmau4_2),.dout(w_dff_B_GNGYj2926_2),.clk(gclk));
	jdff dff_B_MhkjpI8u8_2(.din(w_dff_B_GNGYj2926_2),.dout(w_dff_B_MhkjpI8u8_2),.clk(gclk));
	jdff dff_B_m3iwztcT4_2(.din(w_dff_B_MhkjpI8u8_2),.dout(w_dff_B_m3iwztcT4_2),.clk(gclk));
	jdff dff_B_yzcaKUmW1_2(.din(w_dff_B_m3iwztcT4_2),.dout(w_dff_B_yzcaKUmW1_2),.clk(gclk));
	jdff dff_B_4o77uoY66_2(.din(w_dff_B_yzcaKUmW1_2),.dout(w_dff_B_4o77uoY66_2),.clk(gclk));
	jdff dff_B_JskkLIcq3_2(.din(w_dff_B_4o77uoY66_2),.dout(w_dff_B_JskkLIcq3_2),.clk(gclk));
	jdff dff_B_ObfWJ0v77_2(.din(w_dff_B_JskkLIcq3_2),.dout(w_dff_B_ObfWJ0v77_2),.clk(gclk));
	jdff dff_B_Z5x83MkA7_2(.din(w_dff_B_ObfWJ0v77_2),.dout(w_dff_B_Z5x83MkA7_2),.clk(gclk));
	jdff dff_B_0o0WE9rC9_2(.din(w_dff_B_Z5x83MkA7_2),.dout(w_dff_B_0o0WE9rC9_2),.clk(gclk));
	jdff dff_B_0eA6watc4_2(.din(w_dff_B_0o0WE9rC9_2),.dout(w_dff_B_0eA6watc4_2),.clk(gclk));
	jdff dff_B_dHiVH9Qm0_2(.din(w_dff_B_0eA6watc4_2),.dout(w_dff_B_dHiVH9Qm0_2),.clk(gclk));
	jdff dff_B_18vL9vgB9_2(.din(w_dff_B_dHiVH9Qm0_2),.dout(w_dff_B_18vL9vgB9_2),.clk(gclk));
	jdff dff_B_oBmBB0qd8_2(.din(w_dff_B_18vL9vgB9_2),.dout(w_dff_B_oBmBB0qd8_2),.clk(gclk));
	jdff dff_B_smj5HRXp3_2(.din(w_dff_B_oBmBB0qd8_2),.dout(w_dff_B_smj5HRXp3_2),.clk(gclk));
	jdff dff_B_iAHRBxRd4_2(.din(w_dff_B_smj5HRXp3_2),.dout(w_dff_B_iAHRBxRd4_2),.clk(gclk));
	jdff dff_B_9VX2uy3g5_2(.din(w_dff_B_iAHRBxRd4_2),.dout(w_dff_B_9VX2uy3g5_2),.clk(gclk));
	jdff dff_B_TV43XzgL1_2(.din(w_dff_B_9VX2uy3g5_2),.dout(w_dff_B_TV43XzgL1_2),.clk(gclk));
	jdff dff_B_BwMT4r4s5_2(.din(n1548),.dout(w_dff_B_BwMT4r4s5_2),.clk(gclk));
	jdff dff_B_XiSKkmLA7_1(.din(n1503),.dout(w_dff_B_XiSKkmLA7_1),.clk(gclk));
	jdff dff_B_UFZsLjkw2_2(.din(n1431),.dout(w_dff_B_UFZsLjkw2_2),.clk(gclk));
	jdff dff_B_OxU07TAa7_2(.din(w_dff_B_UFZsLjkw2_2),.dout(w_dff_B_OxU07TAa7_2),.clk(gclk));
	jdff dff_B_b3kbwmDA4_2(.din(w_dff_B_OxU07TAa7_2),.dout(w_dff_B_b3kbwmDA4_2),.clk(gclk));
	jdff dff_B_uzCmvRUr1_2(.din(w_dff_B_b3kbwmDA4_2),.dout(w_dff_B_uzCmvRUr1_2),.clk(gclk));
	jdff dff_B_Q3yPZTjQ0_2(.din(w_dff_B_uzCmvRUr1_2),.dout(w_dff_B_Q3yPZTjQ0_2),.clk(gclk));
	jdff dff_B_JtNrimHy7_2(.din(w_dff_B_Q3yPZTjQ0_2),.dout(w_dff_B_JtNrimHy7_2),.clk(gclk));
	jdff dff_B_vHKvY9xx8_2(.din(w_dff_B_JtNrimHy7_2),.dout(w_dff_B_vHKvY9xx8_2),.clk(gclk));
	jdff dff_B_LYmqUexy1_2(.din(w_dff_B_vHKvY9xx8_2),.dout(w_dff_B_LYmqUexy1_2),.clk(gclk));
	jdff dff_B_nzXB5Axe0_2(.din(w_dff_B_LYmqUexy1_2),.dout(w_dff_B_nzXB5Axe0_2),.clk(gclk));
	jdff dff_B_o0KuoGH45_2(.din(w_dff_B_nzXB5Axe0_2),.dout(w_dff_B_o0KuoGH45_2),.clk(gclk));
	jdff dff_B_HrqJFEGP7_2(.din(w_dff_B_o0KuoGH45_2),.dout(w_dff_B_HrqJFEGP7_2),.clk(gclk));
	jdff dff_B_vwEbBfa66_2(.din(w_dff_B_HrqJFEGP7_2),.dout(w_dff_B_vwEbBfa66_2),.clk(gclk));
	jdff dff_B_j4FjnTbs3_2(.din(w_dff_B_vwEbBfa66_2),.dout(w_dff_B_j4FjnTbs3_2),.clk(gclk));
	jdff dff_B_XTStYCP62_2(.din(w_dff_B_j4FjnTbs3_2),.dout(w_dff_B_XTStYCP62_2),.clk(gclk));
	jdff dff_B_lXXVWJKZ8_2(.din(w_dff_B_XTStYCP62_2),.dout(w_dff_B_lXXVWJKZ8_2),.clk(gclk));
	jdff dff_B_d9bnuhPI1_2(.din(w_dff_B_lXXVWJKZ8_2),.dout(w_dff_B_d9bnuhPI1_2),.clk(gclk));
	jdff dff_B_O00mVJWo6_2(.din(w_dff_B_d9bnuhPI1_2),.dout(w_dff_B_O00mVJWo6_2),.clk(gclk));
	jdff dff_B_OmdAFn3f6_2(.din(w_dff_B_O00mVJWo6_2),.dout(w_dff_B_OmdAFn3f6_2),.clk(gclk));
	jdff dff_B_QrG3MQFZ8_2(.din(w_dff_B_OmdAFn3f6_2),.dout(w_dff_B_QrG3MQFZ8_2),.clk(gclk));
	jdff dff_B_PBiylGLt6_2(.din(w_dff_B_QrG3MQFZ8_2),.dout(w_dff_B_PBiylGLt6_2),.clk(gclk));
	jdff dff_B_UKFjPI116_2(.din(w_dff_B_PBiylGLt6_2),.dout(w_dff_B_UKFjPI116_2),.clk(gclk));
	jdff dff_B_WuS5Uz2n7_2(.din(w_dff_B_UKFjPI116_2),.dout(w_dff_B_WuS5Uz2n7_2),.clk(gclk));
	jdff dff_B_niOnAxFJ5_2(.din(w_dff_B_WuS5Uz2n7_2),.dout(w_dff_B_niOnAxFJ5_2),.clk(gclk));
	jdff dff_B_v9QocWb95_2(.din(w_dff_B_niOnAxFJ5_2),.dout(w_dff_B_v9QocWb95_2),.clk(gclk));
	jdff dff_B_buf3OLjB7_2(.din(w_dff_B_v9QocWb95_2),.dout(w_dff_B_buf3OLjB7_2),.clk(gclk));
	jdff dff_B_yRftY1Vk2_2(.din(w_dff_B_buf3OLjB7_2),.dout(w_dff_B_yRftY1Vk2_2),.clk(gclk));
	jdff dff_B_onEH6jfg7_2(.din(w_dff_B_yRftY1Vk2_2),.dout(w_dff_B_onEH6jfg7_2),.clk(gclk));
	jdff dff_B_tcI9A7fe1_2(.din(w_dff_B_onEH6jfg7_2),.dout(w_dff_B_tcI9A7fe1_2),.clk(gclk));
	jdff dff_B_9mt8ZGc07_2(.din(w_dff_B_tcI9A7fe1_2),.dout(w_dff_B_9mt8ZGc07_2),.clk(gclk));
	jdff dff_B_Tslrz7OR0_2(.din(w_dff_B_9mt8ZGc07_2),.dout(w_dff_B_Tslrz7OR0_2),.clk(gclk));
	jdff dff_B_1OcW82H66_2(.din(w_dff_B_Tslrz7OR0_2),.dout(w_dff_B_1OcW82H66_2),.clk(gclk));
	jdff dff_B_1lC2vAhN2_2(.din(w_dff_B_1OcW82H66_2),.dout(w_dff_B_1lC2vAhN2_2),.clk(gclk));
	jdff dff_B_8Ds5zo293_2(.din(w_dff_B_1lC2vAhN2_2),.dout(w_dff_B_8Ds5zo293_2),.clk(gclk));
	jdff dff_B_6eiamWys7_2(.din(w_dff_B_8Ds5zo293_2),.dout(w_dff_B_6eiamWys7_2),.clk(gclk));
	jdff dff_B_C4rtvTfn2_2(.din(w_dff_B_6eiamWys7_2),.dout(w_dff_B_C4rtvTfn2_2),.clk(gclk));
	jdff dff_B_SjAAH8dP5_2(.din(w_dff_B_C4rtvTfn2_2),.dout(w_dff_B_SjAAH8dP5_2),.clk(gclk));
	jdff dff_B_cXN8GZMR2_2(.din(w_dff_B_SjAAH8dP5_2),.dout(w_dff_B_cXN8GZMR2_2),.clk(gclk));
	jdff dff_B_RFzc39rY8_2(.din(w_dff_B_cXN8GZMR2_2),.dout(w_dff_B_RFzc39rY8_2),.clk(gclk));
	jdff dff_B_dZq68j420_2(.din(w_dff_B_RFzc39rY8_2),.dout(w_dff_B_dZq68j420_2),.clk(gclk));
	jdff dff_B_HDcp3aG34_2(.din(n1477),.dout(w_dff_B_HDcp3aG34_2),.clk(gclk));
	jdff dff_B_1JFEX1qQ4_1(.din(n1432),.dout(w_dff_B_1JFEX1qQ4_1),.clk(gclk));
	jdff dff_B_HZGu3cma2_2(.din(n1353),.dout(w_dff_B_HZGu3cma2_2),.clk(gclk));
	jdff dff_B_XNIyxbBy3_2(.din(w_dff_B_HZGu3cma2_2),.dout(w_dff_B_XNIyxbBy3_2),.clk(gclk));
	jdff dff_B_I98fVVhP9_2(.din(w_dff_B_XNIyxbBy3_2),.dout(w_dff_B_I98fVVhP9_2),.clk(gclk));
	jdff dff_B_ZSGFVfg87_2(.din(w_dff_B_I98fVVhP9_2),.dout(w_dff_B_ZSGFVfg87_2),.clk(gclk));
	jdff dff_B_Q11PkA5z9_2(.din(w_dff_B_ZSGFVfg87_2),.dout(w_dff_B_Q11PkA5z9_2),.clk(gclk));
	jdff dff_B_oIDAby5q5_2(.din(w_dff_B_Q11PkA5z9_2),.dout(w_dff_B_oIDAby5q5_2),.clk(gclk));
	jdff dff_B_qgDDOgEK5_2(.din(w_dff_B_oIDAby5q5_2),.dout(w_dff_B_qgDDOgEK5_2),.clk(gclk));
	jdff dff_B_CmEJZYRf7_2(.din(w_dff_B_qgDDOgEK5_2),.dout(w_dff_B_CmEJZYRf7_2),.clk(gclk));
	jdff dff_B_AZQy3XSX2_2(.din(w_dff_B_CmEJZYRf7_2),.dout(w_dff_B_AZQy3XSX2_2),.clk(gclk));
	jdff dff_B_YHB9kQED6_2(.din(w_dff_B_AZQy3XSX2_2),.dout(w_dff_B_YHB9kQED6_2),.clk(gclk));
	jdff dff_B_s7wvoDhq8_2(.din(w_dff_B_YHB9kQED6_2),.dout(w_dff_B_s7wvoDhq8_2),.clk(gclk));
	jdff dff_B_vY3Anbyk1_2(.din(w_dff_B_s7wvoDhq8_2),.dout(w_dff_B_vY3Anbyk1_2),.clk(gclk));
	jdff dff_B_odDdmaQV4_2(.din(w_dff_B_vY3Anbyk1_2),.dout(w_dff_B_odDdmaQV4_2),.clk(gclk));
	jdff dff_B_Wzpp64Y94_2(.din(w_dff_B_odDdmaQV4_2),.dout(w_dff_B_Wzpp64Y94_2),.clk(gclk));
	jdff dff_B_L8OC3DjU9_2(.din(w_dff_B_Wzpp64Y94_2),.dout(w_dff_B_L8OC3DjU9_2),.clk(gclk));
	jdff dff_B_jIfNha519_2(.din(w_dff_B_L8OC3DjU9_2),.dout(w_dff_B_jIfNha519_2),.clk(gclk));
	jdff dff_B_92Bf2roA2_2(.din(w_dff_B_jIfNha519_2),.dout(w_dff_B_92Bf2roA2_2),.clk(gclk));
	jdff dff_B_Sblvx5pt6_2(.din(w_dff_B_92Bf2roA2_2),.dout(w_dff_B_Sblvx5pt6_2),.clk(gclk));
	jdff dff_B_dR5qpD550_2(.din(w_dff_B_Sblvx5pt6_2),.dout(w_dff_B_dR5qpD550_2),.clk(gclk));
	jdff dff_B_T8zy2mK06_2(.din(w_dff_B_dR5qpD550_2),.dout(w_dff_B_T8zy2mK06_2),.clk(gclk));
	jdff dff_B_4wktHXKN7_2(.din(w_dff_B_T8zy2mK06_2),.dout(w_dff_B_4wktHXKN7_2),.clk(gclk));
	jdff dff_B_PXdDBign1_2(.din(w_dff_B_4wktHXKN7_2),.dout(w_dff_B_PXdDBign1_2),.clk(gclk));
	jdff dff_B_ltelvjfZ1_2(.din(w_dff_B_PXdDBign1_2),.dout(w_dff_B_ltelvjfZ1_2),.clk(gclk));
	jdff dff_B_rdjL7JGq1_2(.din(w_dff_B_ltelvjfZ1_2),.dout(w_dff_B_rdjL7JGq1_2),.clk(gclk));
	jdff dff_B_bx2Zq2VQ7_2(.din(w_dff_B_rdjL7JGq1_2),.dout(w_dff_B_bx2Zq2VQ7_2),.clk(gclk));
	jdff dff_B_rSmeVuHS9_2(.din(w_dff_B_bx2Zq2VQ7_2),.dout(w_dff_B_rSmeVuHS9_2),.clk(gclk));
	jdff dff_B_FDqiVCnI7_2(.din(w_dff_B_rSmeVuHS9_2),.dout(w_dff_B_FDqiVCnI7_2),.clk(gclk));
	jdff dff_B_pq9IWWZu5_2(.din(w_dff_B_FDqiVCnI7_2),.dout(w_dff_B_pq9IWWZu5_2),.clk(gclk));
	jdff dff_B_33Z4DPbN0_2(.din(w_dff_B_pq9IWWZu5_2),.dout(w_dff_B_33Z4DPbN0_2),.clk(gclk));
	jdff dff_B_OjK0KNgq1_2(.din(w_dff_B_33Z4DPbN0_2),.dout(w_dff_B_OjK0KNgq1_2),.clk(gclk));
	jdff dff_B_L3eFov7W4_2(.din(w_dff_B_OjK0KNgq1_2),.dout(w_dff_B_L3eFov7W4_2),.clk(gclk));
	jdff dff_B_b87Rd3sz6_2(.din(w_dff_B_L3eFov7W4_2),.dout(w_dff_B_b87Rd3sz6_2),.clk(gclk));
	jdff dff_B_cSb3M2FH2_2(.din(w_dff_B_b87Rd3sz6_2),.dout(w_dff_B_cSb3M2FH2_2),.clk(gclk));
	jdff dff_B_ixZfKWQW1_2(.din(w_dff_B_cSb3M2FH2_2),.dout(w_dff_B_ixZfKWQW1_2),.clk(gclk));
	jdff dff_B_h44IoPU77_2(.din(w_dff_B_ixZfKWQW1_2),.dout(w_dff_B_h44IoPU77_2),.clk(gclk));
	jdff dff_B_4jwkYf7z2_2(.din(w_dff_B_h44IoPU77_2),.dout(w_dff_B_4jwkYf7z2_2),.clk(gclk));
	jdff dff_B_Fjw6Mauc8_2(.din(n1399),.dout(w_dff_B_Fjw6Mauc8_2),.clk(gclk));
	jdff dff_B_ckoJgik34_1(.din(n1354),.dout(w_dff_B_ckoJgik34_1),.clk(gclk));
	jdff dff_B_BUzwAzmW1_2(.din(n1268),.dout(w_dff_B_BUzwAzmW1_2),.clk(gclk));
	jdff dff_B_nhGAj5Hc6_2(.din(w_dff_B_BUzwAzmW1_2),.dout(w_dff_B_nhGAj5Hc6_2),.clk(gclk));
	jdff dff_B_goePkZZT3_2(.din(w_dff_B_nhGAj5Hc6_2),.dout(w_dff_B_goePkZZT3_2),.clk(gclk));
	jdff dff_B_LQsgcfT99_2(.din(w_dff_B_goePkZZT3_2),.dout(w_dff_B_LQsgcfT99_2),.clk(gclk));
	jdff dff_B_xkuW47bO8_2(.din(w_dff_B_LQsgcfT99_2),.dout(w_dff_B_xkuW47bO8_2),.clk(gclk));
	jdff dff_B_ZXGmVv0z9_2(.din(w_dff_B_xkuW47bO8_2),.dout(w_dff_B_ZXGmVv0z9_2),.clk(gclk));
	jdff dff_B_L6EvGvoJ5_2(.din(w_dff_B_ZXGmVv0z9_2),.dout(w_dff_B_L6EvGvoJ5_2),.clk(gclk));
	jdff dff_B_TS6mNVD46_2(.din(w_dff_B_L6EvGvoJ5_2),.dout(w_dff_B_TS6mNVD46_2),.clk(gclk));
	jdff dff_B_jfFICcWr8_2(.din(w_dff_B_TS6mNVD46_2),.dout(w_dff_B_jfFICcWr8_2),.clk(gclk));
	jdff dff_B_R1sKQJhC0_2(.din(w_dff_B_jfFICcWr8_2),.dout(w_dff_B_R1sKQJhC0_2),.clk(gclk));
	jdff dff_B_Ze2Ww4tU6_2(.din(w_dff_B_R1sKQJhC0_2),.dout(w_dff_B_Ze2Ww4tU6_2),.clk(gclk));
	jdff dff_B_BTBcaIhU8_2(.din(w_dff_B_Ze2Ww4tU6_2),.dout(w_dff_B_BTBcaIhU8_2),.clk(gclk));
	jdff dff_B_pt1L801d0_2(.din(w_dff_B_BTBcaIhU8_2),.dout(w_dff_B_pt1L801d0_2),.clk(gclk));
	jdff dff_B_OwH5Bnl94_2(.din(w_dff_B_pt1L801d0_2),.dout(w_dff_B_OwH5Bnl94_2),.clk(gclk));
	jdff dff_B_kUUqCF2v9_2(.din(w_dff_B_OwH5Bnl94_2),.dout(w_dff_B_kUUqCF2v9_2),.clk(gclk));
	jdff dff_B_1ezRevFb5_2(.din(w_dff_B_kUUqCF2v9_2),.dout(w_dff_B_1ezRevFb5_2),.clk(gclk));
	jdff dff_B_7EaYkE927_2(.din(w_dff_B_1ezRevFb5_2),.dout(w_dff_B_7EaYkE927_2),.clk(gclk));
	jdff dff_B_FkC94jJG1_2(.din(w_dff_B_7EaYkE927_2),.dout(w_dff_B_FkC94jJG1_2),.clk(gclk));
	jdff dff_B_MRv00Cms0_2(.din(w_dff_B_FkC94jJG1_2),.dout(w_dff_B_MRv00Cms0_2),.clk(gclk));
	jdff dff_B_bRLP17tr7_2(.din(w_dff_B_MRv00Cms0_2),.dout(w_dff_B_bRLP17tr7_2),.clk(gclk));
	jdff dff_B_GVDXnYiT3_2(.din(w_dff_B_bRLP17tr7_2),.dout(w_dff_B_GVDXnYiT3_2),.clk(gclk));
	jdff dff_B_tmmyJO6H8_2(.din(w_dff_B_GVDXnYiT3_2),.dout(w_dff_B_tmmyJO6H8_2),.clk(gclk));
	jdff dff_B_KCuZ7vS78_2(.din(w_dff_B_tmmyJO6H8_2),.dout(w_dff_B_KCuZ7vS78_2),.clk(gclk));
	jdff dff_B_8jOKard33_2(.din(w_dff_B_KCuZ7vS78_2),.dout(w_dff_B_8jOKard33_2),.clk(gclk));
	jdff dff_B_I1ZoLuMB0_2(.din(w_dff_B_8jOKard33_2),.dout(w_dff_B_I1ZoLuMB0_2),.clk(gclk));
	jdff dff_B_CjplzZ6j5_2(.din(w_dff_B_I1ZoLuMB0_2),.dout(w_dff_B_CjplzZ6j5_2),.clk(gclk));
	jdff dff_B_W94DCY7N9_2(.din(w_dff_B_CjplzZ6j5_2),.dout(w_dff_B_W94DCY7N9_2),.clk(gclk));
	jdff dff_B_8IRTFaGX9_2(.din(w_dff_B_W94DCY7N9_2),.dout(w_dff_B_8IRTFaGX9_2),.clk(gclk));
	jdff dff_B_T9Hi2CWP2_2(.din(w_dff_B_8IRTFaGX9_2),.dout(w_dff_B_T9Hi2CWP2_2),.clk(gclk));
	jdff dff_B_vGJjGu0s8_2(.din(w_dff_B_T9Hi2CWP2_2),.dout(w_dff_B_vGJjGu0s8_2),.clk(gclk));
	jdff dff_B_TRXvdSrD5_2(.din(w_dff_B_vGJjGu0s8_2),.dout(w_dff_B_TRXvdSrD5_2),.clk(gclk));
	jdff dff_B_rB5tgRum1_2(.din(w_dff_B_TRXvdSrD5_2),.dout(w_dff_B_rB5tgRum1_2),.clk(gclk));
	jdff dff_B_eC9RpPVU6_2(.din(w_dff_B_rB5tgRum1_2),.dout(w_dff_B_eC9RpPVU6_2),.clk(gclk));
	jdff dff_B_2UwdX7bc2_2(.din(n1314),.dout(w_dff_B_2UwdX7bc2_2),.clk(gclk));
	jdff dff_B_q3cqk8wI7_1(.din(n1269),.dout(w_dff_B_q3cqk8wI7_1),.clk(gclk));
	jdff dff_B_auwTIVFR1_2(.din(n1178),.dout(w_dff_B_auwTIVFR1_2),.clk(gclk));
	jdff dff_B_0DsliCtt0_2(.din(w_dff_B_auwTIVFR1_2),.dout(w_dff_B_0DsliCtt0_2),.clk(gclk));
	jdff dff_B_bkOpRP0e6_2(.din(w_dff_B_0DsliCtt0_2),.dout(w_dff_B_bkOpRP0e6_2),.clk(gclk));
	jdff dff_B_LaTCcrM55_2(.din(w_dff_B_bkOpRP0e6_2),.dout(w_dff_B_LaTCcrM55_2),.clk(gclk));
	jdff dff_B_8T85ZtNL2_2(.din(w_dff_B_LaTCcrM55_2),.dout(w_dff_B_8T85ZtNL2_2),.clk(gclk));
	jdff dff_B_oJSSqais1_2(.din(w_dff_B_8T85ZtNL2_2),.dout(w_dff_B_oJSSqais1_2),.clk(gclk));
	jdff dff_B_nJvTM4YU0_2(.din(w_dff_B_oJSSqais1_2),.dout(w_dff_B_nJvTM4YU0_2),.clk(gclk));
	jdff dff_B_tYsAHgzx2_2(.din(w_dff_B_nJvTM4YU0_2),.dout(w_dff_B_tYsAHgzx2_2),.clk(gclk));
	jdff dff_B_DSTjxvUO3_2(.din(w_dff_B_tYsAHgzx2_2),.dout(w_dff_B_DSTjxvUO3_2),.clk(gclk));
	jdff dff_B_FGLdiDzD1_2(.din(w_dff_B_DSTjxvUO3_2),.dout(w_dff_B_FGLdiDzD1_2),.clk(gclk));
	jdff dff_B_5syXlhcn3_2(.din(w_dff_B_FGLdiDzD1_2),.dout(w_dff_B_5syXlhcn3_2),.clk(gclk));
	jdff dff_B_PoHsGxcf9_2(.din(w_dff_B_5syXlhcn3_2),.dout(w_dff_B_PoHsGxcf9_2),.clk(gclk));
	jdff dff_B_pdl2veQ49_2(.din(w_dff_B_PoHsGxcf9_2),.dout(w_dff_B_pdl2veQ49_2),.clk(gclk));
	jdff dff_B_EgZqF5cf8_2(.din(w_dff_B_pdl2veQ49_2),.dout(w_dff_B_EgZqF5cf8_2),.clk(gclk));
	jdff dff_B_PLN4BaHI4_2(.din(w_dff_B_EgZqF5cf8_2),.dout(w_dff_B_PLN4BaHI4_2),.clk(gclk));
	jdff dff_B_TcNQNQQ27_2(.din(w_dff_B_PLN4BaHI4_2),.dout(w_dff_B_TcNQNQQ27_2),.clk(gclk));
	jdff dff_B_ndL5Mfm68_2(.din(w_dff_B_TcNQNQQ27_2),.dout(w_dff_B_ndL5Mfm68_2),.clk(gclk));
	jdff dff_B_JDGjRaL27_2(.din(w_dff_B_ndL5Mfm68_2),.dout(w_dff_B_JDGjRaL27_2),.clk(gclk));
	jdff dff_B_FUppF7bS9_2(.din(w_dff_B_JDGjRaL27_2),.dout(w_dff_B_FUppF7bS9_2),.clk(gclk));
	jdff dff_B_3IPEXlJ09_2(.din(w_dff_B_FUppF7bS9_2),.dout(w_dff_B_3IPEXlJ09_2),.clk(gclk));
	jdff dff_B_URgeEkML7_2(.din(w_dff_B_3IPEXlJ09_2),.dout(w_dff_B_URgeEkML7_2),.clk(gclk));
	jdff dff_B_3AKeL1FL9_2(.din(w_dff_B_URgeEkML7_2),.dout(w_dff_B_3AKeL1FL9_2),.clk(gclk));
	jdff dff_B_SFaYoCVH2_2(.din(w_dff_B_3AKeL1FL9_2),.dout(w_dff_B_SFaYoCVH2_2),.clk(gclk));
	jdff dff_B_S4C5hUq79_2(.din(w_dff_B_SFaYoCVH2_2),.dout(w_dff_B_S4C5hUq79_2),.clk(gclk));
	jdff dff_B_JqsryJaH7_2(.din(w_dff_B_S4C5hUq79_2),.dout(w_dff_B_JqsryJaH7_2),.clk(gclk));
	jdff dff_B_tlftLW2g3_2(.din(w_dff_B_JqsryJaH7_2),.dout(w_dff_B_tlftLW2g3_2),.clk(gclk));
	jdff dff_B_3tMK8PX95_2(.din(w_dff_B_tlftLW2g3_2),.dout(w_dff_B_3tMK8PX95_2),.clk(gclk));
	jdff dff_B_c44AnU8s7_2(.din(w_dff_B_3tMK8PX95_2),.dout(w_dff_B_c44AnU8s7_2),.clk(gclk));
	jdff dff_B_JVPyZeaB5_2(.din(w_dff_B_c44AnU8s7_2),.dout(w_dff_B_JVPyZeaB5_2),.clk(gclk));
	jdff dff_B_xlGvVhf30_2(.din(w_dff_B_JVPyZeaB5_2),.dout(w_dff_B_xlGvVhf30_2),.clk(gclk));
	jdff dff_B_dW6wxl6L3_2(.din(n1223),.dout(w_dff_B_dW6wxl6L3_2),.clk(gclk));
	jdff dff_B_XgFFSGbv9_1(.din(n1179),.dout(w_dff_B_XgFFSGbv9_1),.clk(gclk));
	jdff dff_B_2o09OKuV8_2(.din(n1074),.dout(w_dff_B_2o09OKuV8_2),.clk(gclk));
	jdff dff_B_zgYJ0pHr6_2(.din(w_dff_B_2o09OKuV8_2),.dout(w_dff_B_zgYJ0pHr6_2),.clk(gclk));
	jdff dff_B_nLOEvRYt2_2(.din(w_dff_B_zgYJ0pHr6_2),.dout(w_dff_B_nLOEvRYt2_2),.clk(gclk));
	jdff dff_B_NCjfJO1t4_2(.din(w_dff_B_nLOEvRYt2_2),.dout(w_dff_B_NCjfJO1t4_2),.clk(gclk));
	jdff dff_B_4PD5ByvA2_2(.din(w_dff_B_NCjfJO1t4_2),.dout(w_dff_B_4PD5ByvA2_2),.clk(gclk));
	jdff dff_B_n8SZAGFl6_2(.din(w_dff_B_4PD5ByvA2_2),.dout(w_dff_B_n8SZAGFl6_2),.clk(gclk));
	jdff dff_B_rllWA5NL2_2(.din(w_dff_B_n8SZAGFl6_2),.dout(w_dff_B_rllWA5NL2_2),.clk(gclk));
	jdff dff_B_1TlrS8Wi4_2(.din(w_dff_B_rllWA5NL2_2),.dout(w_dff_B_1TlrS8Wi4_2),.clk(gclk));
	jdff dff_B_4mXHrKEz8_2(.din(w_dff_B_1TlrS8Wi4_2),.dout(w_dff_B_4mXHrKEz8_2),.clk(gclk));
	jdff dff_B_RiGlJB8F7_2(.din(w_dff_B_4mXHrKEz8_2),.dout(w_dff_B_RiGlJB8F7_2),.clk(gclk));
	jdff dff_B_7ErlvpRI7_2(.din(w_dff_B_RiGlJB8F7_2),.dout(w_dff_B_7ErlvpRI7_2),.clk(gclk));
	jdff dff_B_VGQaozw35_2(.din(w_dff_B_7ErlvpRI7_2),.dout(w_dff_B_VGQaozw35_2),.clk(gclk));
	jdff dff_B_iDcCYbTy9_2(.din(w_dff_B_VGQaozw35_2),.dout(w_dff_B_iDcCYbTy9_2),.clk(gclk));
	jdff dff_B_hFnnzyKg9_2(.din(w_dff_B_iDcCYbTy9_2),.dout(w_dff_B_hFnnzyKg9_2),.clk(gclk));
	jdff dff_B_36aCdQqs1_2(.din(w_dff_B_hFnnzyKg9_2),.dout(w_dff_B_36aCdQqs1_2),.clk(gclk));
	jdff dff_B_zJWHwpmw2_2(.din(w_dff_B_36aCdQqs1_2),.dout(w_dff_B_zJWHwpmw2_2),.clk(gclk));
	jdff dff_B_xu99mW7m6_2(.din(w_dff_B_zJWHwpmw2_2),.dout(w_dff_B_xu99mW7m6_2),.clk(gclk));
	jdff dff_B_L9WJ1Hq10_2(.din(w_dff_B_xu99mW7m6_2),.dout(w_dff_B_L9WJ1Hq10_2),.clk(gclk));
	jdff dff_B_OzzuWtfr4_2(.din(w_dff_B_L9WJ1Hq10_2),.dout(w_dff_B_OzzuWtfr4_2),.clk(gclk));
	jdff dff_B_eSSNZ9hf2_2(.din(w_dff_B_OzzuWtfr4_2),.dout(w_dff_B_eSSNZ9hf2_2),.clk(gclk));
	jdff dff_B_0cSgwv064_2(.din(w_dff_B_eSSNZ9hf2_2),.dout(w_dff_B_0cSgwv064_2),.clk(gclk));
	jdff dff_B_Yk2TGZCQ6_2(.din(w_dff_B_0cSgwv064_2),.dout(w_dff_B_Yk2TGZCQ6_2),.clk(gclk));
	jdff dff_B_MeEXKSJ12_2(.din(w_dff_B_Yk2TGZCQ6_2),.dout(w_dff_B_MeEXKSJ12_2),.clk(gclk));
	jdff dff_B_w7HHdtyQ2_2(.din(w_dff_B_MeEXKSJ12_2),.dout(w_dff_B_w7HHdtyQ2_2),.clk(gclk));
	jdff dff_B_RWcd2X5d0_2(.din(w_dff_B_w7HHdtyQ2_2),.dout(w_dff_B_RWcd2X5d0_2),.clk(gclk));
	jdff dff_B_Me1QunXb1_2(.din(w_dff_B_RWcd2X5d0_2),.dout(w_dff_B_Me1QunXb1_2),.clk(gclk));
	jdff dff_B_YDUtoW4R7_2(.din(w_dff_B_Me1QunXb1_2),.dout(w_dff_B_YDUtoW4R7_2),.clk(gclk));
	jdff dff_B_EisvOOA97_2(.din(n1125),.dout(w_dff_B_EisvOOA97_2),.clk(gclk));
	jdff dff_B_UXKY7mn06_1(.din(n1075),.dout(w_dff_B_UXKY7mn06_1),.clk(gclk));
	jdff dff_B_8sgDm9NF2_2(.din(n976),.dout(w_dff_B_8sgDm9NF2_2),.clk(gclk));
	jdff dff_B_TBDdfDyR2_2(.din(w_dff_B_8sgDm9NF2_2),.dout(w_dff_B_TBDdfDyR2_2),.clk(gclk));
	jdff dff_B_r6JjjiU71_2(.din(w_dff_B_TBDdfDyR2_2),.dout(w_dff_B_r6JjjiU71_2),.clk(gclk));
	jdff dff_B_XGovgof19_2(.din(w_dff_B_r6JjjiU71_2),.dout(w_dff_B_XGovgof19_2),.clk(gclk));
	jdff dff_B_Fo1XGixH7_2(.din(w_dff_B_XGovgof19_2),.dout(w_dff_B_Fo1XGixH7_2),.clk(gclk));
	jdff dff_B_C9pKSjZ53_2(.din(w_dff_B_Fo1XGixH7_2),.dout(w_dff_B_C9pKSjZ53_2),.clk(gclk));
	jdff dff_B_BZ0JSpxN5_2(.din(w_dff_B_C9pKSjZ53_2),.dout(w_dff_B_BZ0JSpxN5_2),.clk(gclk));
	jdff dff_B_JOaHNq4c1_2(.din(w_dff_B_BZ0JSpxN5_2),.dout(w_dff_B_JOaHNq4c1_2),.clk(gclk));
	jdff dff_B_HfweC5BM9_2(.din(w_dff_B_JOaHNq4c1_2),.dout(w_dff_B_HfweC5BM9_2),.clk(gclk));
	jdff dff_B_girXWb537_2(.din(w_dff_B_HfweC5BM9_2),.dout(w_dff_B_girXWb537_2),.clk(gclk));
	jdff dff_B_wVH4Xcqz8_2(.din(w_dff_B_girXWb537_2),.dout(w_dff_B_wVH4Xcqz8_2),.clk(gclk));
	jdff dff_B_3ZZ3Zrdy8_2(.din(w_dff_B_wVH4Xcqz8_2),.dout(w_dff_B_3ZZ3Zrdy8_2),.clk(gclk));
	jdff dff_B_MZzN1EZd7_2(.din(w_dff_B_3ZZ3Zrdy8_2),.dout(w_dff_B_MZzN1EZd7_2),.clk(gclk));
	jdff dff_B_qwGsE8z64_2(.din(w_dff_B_MZzN1EZd7_2),.dout(w_dff_B_qwGsE8z64_2),.clk(gclk));
	jdff dff_B_5DkLULiV4_2(.din(w_dff_B_qwGsE8z64_2),.dout(w_dff_B_5DkLULiV4_2),.clk(gclk));
	jdff dff_B_hNzpbAAV5_2(.din(w_dff_B_5DkLULiV4_2),.dout(w_dff_B_hNzpbAAV5_2),.clk(gclk));
	jdff dff_B_hXs4bfJi6_2(.din(w_dff_B_hNzpbAAV5_2),.dout(w_dff_B_hXs4bfJi6_2),.clk(gclk));
	jdff dff_B_F1VjSATd5_2(.din(w_dff_B_hXs4bfJi6_2),.dout(w_dff_B_F1VjSATd5_2),.clk(gclk));
	jdff dff_B_TwQghdDz1_2(.din(w_dff_B_F1VjSATd5_2),.dout(w_dff_B_TwQghdDz1_2),.clk(gclk));
	jdff dff_B_EtLqrdVo4_2(.din(w_dff_B_TwQghdDz1_2),.dout(w_dff_B_EtLqrdVo4_2),.clk(gclk));
	jdff dff_B_xKke7LSc0_2(.din(w_dff_B_EtLqrdVo4_2),.dout(w_dff_B_xKke7LSc0_2),.clk(gclk));
	jdff dff_B_IAYLx7mw7_2(.din(w_dff_B_xKke7LSc0_2),.dout(w_dff_B_IAYLx7mw7_2),.clk(gclk));
	jdff dff_B_6dGQuVQ40_2(.din(w_dff_B_IAYLx7mw7_2),.dout(w_dff_B_6dGQuVQ40_2),.clk(gclk));
	jdff dff_B_g97xEijh0_2(.din(w_dff_B_6dGQuVQ40_2),.dout(w_dff_B_g97xEijh0_2),.clk(gclk));
	jdff dff_B_FNpHUw6v3_2(.din(n1020),.dout(w_dff_B_FNpHUw6v3_2),.clk(gclk));
	jdff dff_B_hxo8JQPg8_1(.din(n977),.dout(w_dff_B_hxo8JQPg8_1),.clk(gclk));
	jdff dff_B_mYCkYm2d2_2(.din(n871),.dout(w_dff_B_mYCkYm2d2_2),.clk(gclk));
	jdff dff_B_VYQj7Cxz5_2(.din(w_dff_B_mYCkYm2d2_2),.dout(w_dff_B_VYQj7Cxz5_2),.clk(gclk));
	jdff dff_B_fB3zviGM0_2(.din(w_dff_B_VYQj7Cxz5_2),.dout(w_dff_B_fB3zviGM0_2),.clk(gclk));
	jdff dff_B_5iPVPvLl8_2(.din(w_dff_B_fB3zviGM0_2),.dout(w_dff_B_5iPVPvLl8_2),.clk(gclk));
	jdff dff_B_MveOTinn4_2(.din(w_dff_B_5iPVPvLl8_2),.dout(w_dff_B_MveOTinn4_2),.clk(gclk));
	jdff dff_B_Jz4oOYo95_2(.din(w_dff_B_MveOTinn4_2),.dout(w_dff_B_Jz4oOYo95_2),.clk(gclk));
	jdff dff_B_wHK2ikOq9_2(.din(w_dff_B_Jz4oOYo95_2),.dout(w_dff_B_wHK2ikOq9_2),.clk(gclk));
	jdff dff_B_I8Epqzad1_2(.din(w_dff_B_wHK2ikOq9_2),.dout(w_dff_B_I8Epqzad1_2),.clk(gclk));
	jdff dff_B_qQDpREwL1_2(.din(w_dff_B_I8Epqzad1_2),.dout(w_dff_B_qQDpREwL1_2),.clk(gclk));
	jdff dff_B_FnVBqF0B2_2(.din(w_dff_B_qQDpREwL1_2),.dout(w_dff_B_FnVBqF0B2_2),.clk(gclk));
	jdff dff_B_6G4OdG8v9_2(.din(w_dff_B_FnVBqF0B2_2),.dout(w_dff_B_6G4OdG8v9_2),.clk(gclk));
	jdff dff_B_RpOu18NR3_2(.din(w_dff_B_6G4OdG8v9_2),.dout(w_dff_B_RpOu18NR3_2),.clk(gclk));
	jdff dff_B_AnvPfdSS4_2(.din(w_dff_B_RpOu18NR3_2),.dout(w_dff_B_AnvPfdSS4_2),.clk(gclk));
	jdff dff_B_heKggPzN9_2(.din(w_dff_B_AnvPfdSS4_2),.dout(w_dff_B_heKggPzN9_2),.clk(gclk));
	jdff dff_B_YnvwImeh3_2(.din(w_dff_B_heKggPzN9_2),.dout(w_dff_B_YnvwImeh3_2),.clk(gclk));
	jdff dff_B_hdgmBAZ34_2(.din(w_dff_B_YnvwImeh3_2),.dout(w_dff_B_hdgmBAZ34_2),.clk(gclk));
	jdff dff_B_diaAH8yP6_2(.din(w_dff_B_hdgmBAZ34_2),.dout(w_dff_B_diaAH8yP6_2),.clk(gclk));
	jdff dff_B_3LujCoJV6_2(.din(w_dff_B_diaAH8yP6_2),.dout(w_dff_B_3LujCoJV6_2),.clk(gclk));
	jdff dff_B_a4iW99d93_2(.din(w_dff_B_3LujCoJV6_2),.dout(w_dff_B_a4iW99d93_2),.clk(gclk));
	jdff dff_B_CjApRlu04_2(.din(w_dff_B_a4iW99d93_2),.dout(w_dff_B_CjApRlu04_2),.clk(gclk));
	jdff dff_B_22rxImAM4_2(.din(w_dff_B_CjApRlu04_2),.dout(w_dff_B_22rxImAM4_2),.clk(gclk));
	jdff dff_B_znWFqW642_2(.din(n915),.dout(w_dff_B_znWFqW642_2),.clk(gclk));
	jdff dff_B_7ThjlGih2_1(.din(n872),.dout(w_dff_B_7ThjlGih2_1),.clk(gclk));
	jdff dff_B_XaOk3fSX7_2(.din(n772),.dout(w_dff_B_XaOk3fSX7_2),.clk(gclk));
	jdff dff_B_JO6KkWhK4_2(.din(w_dff_B_XaOk3fSX7_2),.dout(w_dff_B_JO6KkWhK4_2),.clk(gclk));
	jdff dff_B_lfY27dJP3_2(.din(w_dff_B_JO6KkWhK4_2),.dout(w_dff_B_lfY27dJP3_2),.clk(gclk));
	jdff dff_B_jneRnVpk7_2(.din(w_dff_B_lfY27dJP3_2),.dout(w_dff_B_jneRnVpk7_2),.clk(gclk));
	jdff dff_B_yB8FO8Wb0_2(.din(w_dff_B_jneRnVpk7_2),.dout(w_dff_B_yB8FO8Wb0_2),.clk(gclk));
	jdff dff_B_fr8RiATb0_2(.din(w_dff_B_yB8FO8Wb0_2),.dout(w_dff_B_fr8RiATb0_2),.clk(gclk));
	jdff dff_B_droAkZxZ3_2(.din(w_dff_B_fr8RiATb0_2),.dout(w_dff_B_droAkZxZ3_2),.clk(gclk));
	jdff dff_B_CGHNnbgz0_2(.din(w_dff_B_droAkZxZ3_2),.dout(w_dff_B_CGHNnbgz0_2),.clk(gclk));
	jdff dff_B_XRuruMet1_2(.din(w_dff_B_CGHNnbgz0_2),.dout(w_dff_B_XRuruMet1_2),.clk(gclk));
	jdff dff_B_UrkMKO8C4_2(.din(w_dff_B_XRuruMet1_2),.dout(w_dff_B_UrkMKO8C4_2),.clk(gclk));
	jdff dff_B_uZXURiRo4_2(.din(w_dff_B_UrkMKO8C4_2),.dout(w_dff_B_uZXURiRo4_2),.clk(gclk));
	jdff dff_B_vK2tTix46_2(.din(w_dff_B_uZXURiRo4_2),.dout(w_dff_B_vK2tTix46_2),.clk(gclk));
	jdff dff_B_JELBREoE1_2(.din(w_dff_B_vK2tTix46_2),.dout(w_dff_B_JELBREoE1_2),.clk(gclk));
	jdff dff_B_hi6wsLRV7_2(.din(w_dff_B_JELBREoE1_2),.dout(w_dff_B_hi6wsLRV7_2),.clk(gclk));
	jdff dff_B_EUHJQGSs1_2(.din(w_dff_B_hi6wsLRV7_2),.dout(w_dff_B_EUHJQGSs1_2),.clk(gclk));
	jdff dff_B_QlcaS6xt6_2(.din(w_dff_B_EUHJQGSs1_2),.dout(w_dff_B_QlcaS6xt6_2),.clk(gclk));
	jdff dff_B_CpTTwEOK3_2(.din(w_dff_B_QlcaS6xt6_2),.dout(w_dff_B_CpTTwEOK3_2),.clk(gclk));
	jdff dff_B_ikKPjnGQ6_2(.din(w_dff_B_CpTTwEOK3_2),.dout(w_dff_B_ikKPjnGQ6_2),.clk(gclk));
	jdff dff_B_szXqKr1U5_2(.din(n809),.dout(w_dff_B_szXqKr1U5_2),.clk(gclk));
	jdff dff_B_EHm0L3KP9_1(.din(n773),.dout(w_dff_B_EHm0L3KP9_1),.clk(gclk));
	jdff dff_B_HyrPJHJQ3_2(.din(n679),.dout(w_dff_B_HyrPJHJQ3_2),.clk(gclk));
	jdff dff_B_GDAsc6sk7_2(.din(w_dff_B_HyrPJHJQ3_2),.dout(w_dff_B_GDAsc6sk7_2),.clk(gclk));
	jdff dff_B_NDxrJoVg9_2(.din(w_dff_B_GDAsc6sk7_2),.dout(w_dff_B_NDxrJoVg9_2),.clk(gclk));
	jdff dff_B_SEvZthWw3_2(.din(w_dff_B_NDxrJoVg9_2),.dout(w_dff_B_SEvZthWw3_2),.clk(gclk));
	jdff dff_B_EdB1Pe199_2(.din(w_dff_B_SEvZthWw3_2),.dout(w_dff_B_EdB1Pe199_2),.clk(gclk));
	jdff dff_B_GguUIXlm3_2(.din(w_dff_B_EdB1Pe199_2),.dout(w_dff_B_GguUIXlm3_2),.clk(gclk));
	jdff dff_B_U4KAo54S1_2(.din(w_dff_B_GguUIXlm3_2),.dout(w_dff_B_U4KAo54S1_2),.clk(gclk));
	jdff dff_B_K1waBADP9_2(.din(w_dff_B_U4KAo54S1_2),.dout(w_dff_B_K1waBADP9_2),.clk(gclk));
	jdff dff_B_SWPEdXiK2_2(.din(w_dff_B_K1waBADP9_2),.dout(w_dff_B_SWPEdXiK2_2),.clk(gclk));
	jdff dff_B_9byeOhXv5_2(.din(w_dff_B_SWPEdXiK2_2),.dout(w_dff_B_9byeOhXv5_2),.clk(gclk));
	jdff dff_B_Shz1Aqw69_2(.din(w_dff_B_9byeOhXv5_2),.dout(w_dff_B_Shz1Aqw69_2),.clk(gclk));
	jdff dff_B_4e2VIIbb2_2(.din(w_dff_B_Shz1Aqw69_2),.dout(w_dff_B_4e2VIIbb2_2),.clk(gclk));
	jdff dff_B_oKTa9Z6e8_2(.din(w_dff_B_4e2VIIbb2_2),.dout(w_dff_B_oKTa9Z6e8_2),.clk(gclk));
	jdff dff_B_PnGStDAv7_2(.din(w_dff_B_oKTa9Z6e8_2),.dout(w_dff_B_PnGStDAv7_2),.clk(gclk));
	jdff dff_B_k2iDG3JR1_2(.din(w_dff_B_PnGStDAv7_2),.dout(w_dff_B_k2iDG3JR1_2),.clk(gclk));
	jdff dff_B_rnu65OlP0_2(.din(n709),.dout(w_dff_B_rnu65OlP0_2),.clk(gclk));
	jdff dff_B_Y9MhPSzk2_1(.din(n680),.dout(w_dff_B_Y9MhPSzk2_1),.clk(gclk));
	jdff dff_B_LIXcAc2O5_2(.din(n593),.dout(w_dff_B_LIXcAc2O5_2),.clk(gclk));
	jdff dff_B_mvFRcGWT2_2(.din(w_dff_B_LIXcAc2O5_2),.dout(w_dff_B_mvFRcGWT2_2),.clk(gclk));
	jdff dff_B_onSIMLQJ6_2(.din(w_dff_B_mvFRcGWT2_2),.dout(w_dff_B_onSIMLQJ6_2),.clk(gclk));
	jdff dff_B_z7hSY4bY5_2(.din(w_dff_B_onSIMLQJ6_2),.dout(w_dff_B_z7hSY4bY5_2),.clk(gclk));
	jdff dff_B_4T76rDuK2_2(.din(w_dff_B_z7hSY4bY5_2),.dout(w_dff_B_4T76rDuK2_2),.clk(gclk));
	jdff dff_B_DlqGR35S1_2(.din(w_dff_B_4T76rDuK2_2),.dout(w_dff_B_DlqGR35S1_2),.clk(gclk));
	jdff dff_B_IYdwAWZH0_2(.din(w_dff_B_DlqGR35S1_2),.dout(w_dff_B_IYdwAWZH0_2),.clk(gclk));
	jdff dff_B_ypl0N8wR2_2(.din(w_dff_B_IYdwAWZH0_2),.dout(w_dff_B_ypl0N8wR2_2),.clk(gclk));
	jdff dff_B_ZHpkIu0s7_2(.din(w_dff_B_ypl0N8wR2_2),.dout(w_dff_B_ZHpkIu0s7_2),.clk(gclk));
	jdff dff_B_XLpWBxtc2_2(.din(w_dff_B_ZHpkIu0s7_2),.dout(w_dff_B_XLpWBxtc2_2),.clk(gclk));
	jdff dff_B_hepGxWQP0_2(.din(w_dff_B_XLpWBxtc2_2),.dout(w_dff_B_hepGxWQP0_2),.clk(gclk));
	jdff dff_B_NZTP6NYu9_2(.din(w_dff_B_hepGxWQP0_2),.dout(w_dff_B_NZTP6NYu9_2),.clk(gclk));
	jdff dff_B_fZAO0HLr4_2(.din(n616),.dout(w_dff_B_fZAO0HLr4_2),.clk(gclk));
	jdff dff_B_9ghebZGk8_1(.din(n594),.dout(w_dff_B_9ghebZGk8_1),.clk(gclk));
	jdff dff_B_lQCrSu5l7_2(.din(n514),.dout(w_dff_B_lQCrSu5l7_2),.clk(gclk));
	jdff dff_B_oIP1yoqL8_2(.din(w_dff_B_lQCrSu5l7_2),.dout(w_dff_B_oIP1yoqL8_2),.clk(gclk));
	jdff dff_B_IcS8Xf7q7_2(.din(w_dff_B_oIP1yoqL8_2),.dout(w_dff_B_IcS8Xf7q7_2),.clk(gclk));
	jdff dff_B_VIutb0F06_2(.din(w_dff_B_IcS8Xf7q7_2),.dout(w_dff_B_VIutb0F06_2),.clk(gclk));
	jdff dff_B_9QkdcicG0_2(.din(w_dff_B_VIutb0F06_2),.dout(w_dff_B_9QkdcicG0_2),.clk(gclk));
	jdff dff_B_P5mEoDRL9_2(.din(w_dff_B_9QkdcicG0_2),.dout(w_dff_B_P5mEoDRL9_2),.clk(gclk));
	jdff dff_B_IwPzVIZl5_2(.din(w_dff_B_P5mEoDRL9_2),.dout(w_dff_B_IwPzVIZl5_2),.clk(gclk));
	jdff dff_B_a0lQqF4h6_2(.din(w_dff_B_IwPzVIZl5_2),.dout(w_dff_B_a0lQqF4h6_2),.clk(gclk));
	jdff dff_B_ldFlnqha2_2(.din(w_dff_B_a0lQqF4h6_2),.dout(w_dff_B_ldFlnqha2_2),.clk(gclk));
	jdff dff_B_2i1IVh7i6_2(.din(n530),.dout(w_dff_B_2i1IVh7i6_2),.clk(gclk));
	jdff dff_B_AaPrnNlc1_2(.din(w_dff_B_2i1IVh7i6_2),.dout(w_dff_B_AaPrnNlc1_2),.clk(gclk));
	jdff dff_B_8EbeydnL5_1(.din(n515),.dout(w_dff_B_8EbeydnL5_1),.clk(gclk));
	jdff dff_B_ttxOODxp4_1(.din(w_dff_B_8EbeydnL5_1),.dout(w_dff_B_ttxOODxp4_1),.clk(gclk));
	jdff dff_B_SNA3vDRz5_1(.din(w_dff_B_ttxOODxp4_1),.dout(w_dff_B_SNA3vDRz5_1),.clk(gclk));
	jdff dff_B_isjKHTxj5_1(.din(w_dff_B_SNA3vDRz5_1),.dout(w_dff_B_isjKHTxj5_1),.clk(gclk));
	jdff dff_B_3ZRXdkm85_1(.din(w_dff_B_isjKHTxj5_1),.dout(w_dff_B_3ZRXdkm85_1),.clk(gclk));
	jdff dff_B_qyNN8air7_1(.din(w_dff_B_3ZRXdkm85_1),.dout(w_dff_B_qyNN8air7_1),.clk(gclk));
	jdff dff_B_tFPh4Pe25_0(.din(n451),.dout(w_dff_B_tFPh4Pe25_0),.clk(gclk));
	jdff dff_B_RAreoxw01_0(.din(w_dff_B_tFPh4Pe25_0),.dout(w_dff_B_RAreoxw01_0),.clk(gclk));
	jdff dff_A_tAE24NYn6_0(.dout(w_n450_0[0]),.din(w_dff_A_tAE24NYn6_0),.clk(gclk));
	jdff dff_A_SiIxT2xb8_0(.dout(w_dff_A_tAE24NYn6_0),.din(w_dff_A_SiIxT2xb8_0),.clk(gclk));
	jdff dff_A_1dQUkF5l2_0(.dout(w_dff_A_SiIxT2xb8_0),.din(w_dff_A_1dQUkF5l2_0),.clk(gclk));
	jdff dff_B_N7i4VHMt8_1(.din(n444),.dout(w_dff_B_N7i4VHMt8_1),.clk(gclk));
	jdff dff_A_vbg071tF9_0(.dout(w_n376_0[0]),.din(w_dff_A_vbg071tF9_0),.clk(gclk));
	jdff dff_A_Wwcu4ipG4_1(.dout(w_n376_0[1]),.din(w_dff_A_Wwcu4ipG4_1),.clk(gclk));
	jdff dff_A_zMPDIusV4_1(.dout(w_dff_A_Wwcu4ipG4_1),.din(w_dff_A_zMPDIusV4_1),.clk(gclk));
	jdff dff_A_W4w189eW0_1(.dout(w_n442_0[1]),.din(w_dff_A_W4w189eW0_1),.clk(gclk));
	jdff dff_A_a2mVrLoC1_1(.dout(w_dff_A_W4w189eW0_1),.din(w_dff_A_a2mVrLoC1_1),.clk(gclk));
	jdff dff_A_SrNpZSN95_1(.dout(w_dff_A_a2mVrLoC1_1),.din(w_dff_A_SrNpZSN95_1),.clk(gclk));
	jdff dff_A_Dm8KbRbH0_1(.dout(w_dff_A_SrNpZSN95_1),.din(w_dff_A_Dm8KbRbH0_1),.clk(gclk));
	jdff dff_A_smyor4li1_1(.dout(w_dff_A_Dm8KbRbH0_1),.din(w_dff_A_smyor4li1_1),.clk(gclk));
	jdff dff_A_tRz3lwnQ9_1(.dout(w_dff_A_smyor4li1_1),.din(w_dff_A_tRz3lwnQ9_1),.clk(gclk));
	jdff dff_B_AsdTUFM99_2(.din(n1682),.dout(w_dff_B_AsdTUFM99_2),.clk(gclk));
	jdff dff_B_YpIpUHEK4_1(.din(n1680),.dout(w_dff_B_YpIpUHEK4_1),.clk(gclk));
	jdff dff_B_PArHlcTp7_2(.din(n1628),.dout(w_dff_B_PArHlcTp7_2),.clk(gclk));
	jdff dff_B_qiwI0KSH8_2(.din(w_dff_B_PArHlcTp7_2),.dout(w_dff_B_qiwI0KSH8_2),.clk(gclk));
	jdff dff_B_cKtvtclL9_2(.din(w_dff_B_qiwI0KSH8_2),.dout(w_dff_B_cKtvtclL9_2),.clk(gclk));
	jdff dff_B_0LNSKlF92_2(.din(w_dff_B_cKtvtclL9_2),.dout(w_dff_B_0LNSKlF92_2),.clk(gclk));
	jdff dff_B_J4sxSRGO4_2(.din(w_dff_B_0LNSKlF92_2),.dout(w_dff_B_J4sxSRGO4_2),.clk(gclk));
	jdff dff_B_z8U5FOiJ5_2(.din(w_dff_B_J4sxSRGO4_2),.dout(w_dff_B_z8U5FOiJ5_2),.clk(gclk));
	jdff dff_B_dLOTGVoM0_2(.din(w_dff_B_z8U5FOiJ5_2),.dout(w_dff_B_dLOTGVoM0_2),.clk(gclk));
	jdff dff_B_YlSTYzZj9_2(.din(w_dff_B_dLOTGVoM0_2),.dout(w_dff_B_YlSTYzZj9_2),.clk(gclk));
	jdff dff_B_JyIuXjHS8_2(.din(w_dff_B_YlSTYzZj9_2),.dout(w_dff_B_JyIuXjHS8_2),.clk(gclk));
	jdff dff_B_YgBJPPjW0_2(.din(w_dff_B_JyIuXjHS8_2),.dout(w_dff_B_YgBJPPjW0_2),.clk(gclk));
	jdff dff_B_Szt3aTFi8_2(.din(w_dff_B_YgBJPPjW0_2),.dout(w_dff_B_Szt3aTFi8_2),.clk(gclk));
	jdff dff_B_snRKwoe24_2(.din(w_dff_B_Szt3aTFi8_2),.dout(w_dff_B_snRKwoe24_2),.clk(gclk));
	jdff dff_B_MpW5awIF6_2(.din(w_dff_B_snRKwoe24_2),.dout(w_dff_B_MpW5awIF6_2),.clk(gclk));
	jdff dff_B_FxxATGpD3_2(.din(w_dff_B_MpW5awIF6_2),.dout(w_dff_B_FxxATGpD3_2),.clk(gclk));
	jdff dff_B_amgqkloe2_2(.din(w_dff_B_FxxATGpD3_2),.dout(w_dff_B_amgqkloe2_2),.clk(gclk));
	jdff dff_B_WsOKPWoK0_2(.din(w_dff_B_amgqkloe2_2),.dout(w_dff_B_WsOKPWoK0_2),.clk(gclk));
	jdff dff_B_PEQ2wayV7_2(.din(w_dff_B_WsOKPWoK0_2),.dout(w_dff_B_PEQ2wayV7_2),.clk(gclk));
	jdff dff_B_GVk2yZF33_2(.din(w_dff_B_PEQ2wayV7_2),.dout(w_dff_B_GVk2yZF33_2),.clk(gclk));
	jdff dff_B_xDf3TU6n5_2(.din(w_dff_B_GVk2yZF33_2),.dout(w_dff_B_xDf3TU6n5_2),.clk(gclk));
	jdff dff_B_GBlKSAWE9_2(.din(w_dff_B_xDf3TU6n5_2),.dout(w_dff_B_GBlKSAWE9_2),.clk(gclk));
	jdff dff_B_V03I3ieu8_2(.din(w_dff_B_GBlKSAWE9_2),.dout(w_dff_B_V03I3ieu8_2),.clk(gclk));
	jdff dff_B_Sd3JDFYY6_2(.din(w_dff_B_V03I3ieu8_2),.dout(w_dff_B_Sd3JDFYY6_2),.clk(gclk));
	jdff dff_B_bZJ2N5px0_2(.din(w_dff_B_Sd3JDFYY6_2),.dout(w_dff_B_bZJ2N5px0_2),.clk(gclk));
	jdff dff_B_AowOnzXc9_2(.din(w_dff_B_bZJ2N5px0_2),.dout(w_dff_B_AowOnzXc9_2),.clk(gclk));
	jdff dff_B_dpQU4WUr3_2(.din(w_dff_B_AowOnzXc9_2),.dout(w_dff_B_dpQU4WUr3_2),.clk(gclk));
	jdff dff_B_s3U6reL44_2(.din(w_dff_B_dpQU4WUr3_2),.dout(w_dff_B_s3U6reL44_2),.clk(gclk));
	jdff dff_B_P58tzSC07_2(.din(w_dff_B_s3U6reL44_2),.dout(w_dff_B_P58tzSC07_2),.clk(gclk));
	jdff dff_B_5lApa9jI1_2(.din(w_dff_B_P58tzSC07_2),.dout(w_dff_B_5lApa9jI1_2),.clk(gclk));
	jdff dff_B_GKWVAdBZ3_2(.din(w_dff_B_5lApa9jI1_2),.dout(w_dff_B_GKWVAdBZ3_2),.clk(gclk));
	jdff dff_B_C6jXFXyJ4_2(.din(w_dff_B_GKWVAdBZ3_2),.dout(w_dff_B_C6jXFXyJ4_2),.clk(gclk));
	jdff dff_B_a83QJQJW7_2(.din(w_dff_B_C6jXFXyJ4_2),.dout(w_dff_B_a83QJQJW7_2),.clk(gclk));
	jdff dff_B_ImdX8alE0_2(.din(w_dff_B_a83QJQJW7_2),.dout(w_dff_B_ImdX8alE0_2),.clk(gclk));
	jdff dff_B_N5mzrMAR5_2(.din(w_dff_B_ImdX8alE0_2),.dout(w_dff_B_N5mzrMAR5_2),.clk(gclk));
	jdff dff_B_SC5LjA8y3_2(.din(w_dff_B_N5mzrMAR5_2),.dout(w_dff_B_SC5LjA8y3_2),.clk(gclk));
	jdff dff_B_UaAiIiiB6_2(.din(w_dff_B_SC5LjA8y3_2),.dout(w_dff_B_UaAiIiiB6_2),.clk(gclk));
	jdff dff_B_ZEMXU4sU1_2(.din(w_dff_B_UaAiIiiB6_2),.dout(w_dff_B_ZEMXU4sU1_2),.clk(gclk));
	jdff dff_B_r8ryJgr71_2(.din(w_dff_B_ZEMXU4sU1_2),.dout(w_dff_B_r8ryJgr71_2),.clk(gclk));
	jdff dff_B_ij2djt9q8_2(.din(w_dff_B_r8ryJgr71_2),.dout(w_dff_B_ij2djt9q8_2),.clk(gclk));
	jdff dff_B_If8Kb8MC5_2(.din(w_dff_B_ij2djt9q8_2),.dout(w_dff_B_If8Kb8MC5_2),.clk(gclk));
	jdff dff_B_r4cU4sKg0_2(.din(w_dff_B_If8Kb8MC5_2),.dout(w_dff_B_r4cU4sKg0_2),.clk(gclk));
	jdff dff_B_i3zVcTM01_2(.din(w_dff_B_r4cU4sKg0_2),.dout(w_dff_B_i3zVcTM01_2),.clk(gclk));
	jdff dff_B_4k1mpOB02_2(.din(w_dff_B_i3zVcTM01_2),.dout(w_dff_B_4k1mpOB02_2),.clk(gclk));
	jdff dff_B_wykz0jUS4_2(.din(w_dff_B_4k1mpOB02_2),.dout(w_dff_B_wykz0jUS4_2),.clk(gclk));
	jdff dff_B_4sxKzeg92_2(.din(w_dff_B_wykz0jUS4_2),.dout(w_dff_B_4sxKzeg92_2),.clk(gclk));
	jdff dff_B_VzGOJpHZ2_2(.din(w_dff_B_4sxKzeg92_2),.dout(w_dff_B_VzGOJpHZ2_2),.clk(gclk));
	jdff dff_B_ppU07i4X5_2(.din(w_dff_B_VzGOJpHZ2_2),.dout(w_dff_B_ppU07i4X5_2),.clk(gclk));
	jdff dff_B_SOd0D7wR4_2(.din(w_dff_B_ppU07i4X5_2),.dout(w_dff_B_SOd0D7wR4_2),.clk(gclk));
	jdff dff_B_WUkWgVNA1_2(.din(w_dff_B_SOd0D7wR4_2),.dout(w_dff_B_WUkWgVNA1_2),.clk(gclk));
	jdff dff_B_okOZllCj2_2(.din(w_dff_B_WUkWgVNA1_2),.dout(w_dff_B_okOZllCj2_2),.clk(gclk));
	jdff dff_B_BpAGy5bV6_1(.din(n1678),.dout(w_dff_B_BpAGy5bV6_1),.clk(gclk));
	jdff dff_A_Wswiurrn4_1(.dout(w_n1631_0[1]),.din(w_dff_A_Wswiurrn4_1),.clk(gclk));
	jdff dff_B_5Zokezc54_1(.din(n1629),.dout(w_dff_B_5Zokezc54_1),.clk(gclk));
	jdff dff_B_EII6tz7c4_2(.din(n1571),.dout(w_dff_B_EII6tz7c4_2),.clk(gclk));
	jdff dff_B_5iBeThyd4_2(.din(w_dff_B_EII6tz7c4_2),.dout(w_dff_B_5iBeThyd4_2),.clk(gclk));
	jdff dff_B_X06eB6e28_2(.din(w_dff_B_5iBeThyd4_2),.dout(w_dff_B_X06eB6e28_2),.clk(gclk));
	jdff dff_B_0Q2tU6qi6_2(.din(w_dff_B_X06eB6e28_2),.dout(w_dff_B_0Q2tU6qi6_2),.clk(gclk));
	jdff dff_B_rCvZpAjm5_2(.din(w_dff_B_0Q2tU6qi6_2),.dout(w_dff_B_rCvZpAjm5_2),.clk(gclk));
	jdff dff_B_dXyaVulQ1_2(.din(w_dff_B_rCvZpAjm5_2),.dout(w_dff_B_dXyaVulQ1_2),.clk(gclk));
	jdff dff_B_FYtV1i0B1_2(.din(w_dff_B_dXyaVulQ1_2),.dout(w_dff_B_FYtV1i0B1_2),.clk(gclk));
	jdff dff_B_XEC6lTLt3_2(.din(w_dff_B_FYtV1i0B1_2),.dout(w_dff_B_XEC6lTLt3_2),.clk(gclk));
	jdff dff_B_ZMzzyrzm2_2(.din(w_dff_B_XEC6lTLt3_2),.dout(w_dff_B_ZMzzyrzm2_2),.clk(gclk));
	jdff dff_B_kyp6GfXr6_2(.din(w_dff_B_ZMzzyrzm2_2),.dout(w_dff_B_kyp6GfXr6_2),.clk(gclk));
	jdff dff_B_4vyHJ6G09_2(.din(w_dff_B_kyp6GfXr6_2),.dout(w_dff_B_4vyHJ6G09_2),.clk(gclk));
	jdff dff_B_5SOLiOdu3_2(.din(w_dff_B_4vyHJ6G09_2),.dout(w_dff_B_5SOLiOdu3_2),.clk(gclk));
	jdff dff_B_o1GIZ1Sd5_2(.din(w_dff_B_5SOLiOdu3_2),.dout(w_dff_B_o1GIZ1Sd5_2),.clk(gclk));
	jdff dff_B_3la8R4sz0_2(.din(w_dff_B_o1GIZ1Sd5_2),.dout(w_dff_B_3la8R4sz0_2),.clk(gclk));
	jdff dff_B_hu7kdU4w6_2(.din(w_dff_B_3la8R4sz0_2),.dout(w_dff_B_hu7kdU4w6_2),.clk(gclk));
	jdff dff_B_h07Pw2yX7_2(.din(w_dff_B_hu7kdU4w6_2),.dout(w_dff_B_h07Pw2yX7_2),.clk(gclk));
	jdff dff_B_9V2VZvxe5_2(.din(w_dff_B_h07Pw2yX7_2),.dout(w_dff_B_9V2VZvxe5_2),.clk(gclk));
	jdff dff_B_ASsZyJm94_2(.din(w_dff_B_9V2VZvxe5_2),.dout(w_dff_B_ASsZyJm94_2),.clk(gclk));
	jdff dff_B_A9yI4gMT4_2(.din(w_dff_B_ASsZyJm94_2),.dout(w_dff_B_A9yI4gMT4_2),.clk(gclk));
	jdff dff_B_u5Omsozp9_2(.din(w_dff_B_A9yI4gMT4_2),.dout(w_dff_B_u5Omsozp9_2),.clk(gclk));
	jdff dff_B_yprUHcKH6_2(.din(w_dff_B_u5Omsozp9_2),.dout(w_dff_B_yprUHcKH6_2),.clk(gclk));
	jdff dff_B_s3PM9E6V0_2(.din(w_dff_B_yprUHcKH6_2),.dout(w_dff_B_s3PM9E6V0_2),.clk(gclk));
	jdff dff_B_mBAHCuQW4_2(.din(w_dff_B_s3PM9E6V0_2),.dout(w_dff_B_mBAHCuQW4_2),.clk(gclk));
	jdff dff_B_wa7If9a09_2(.din(w_dff_B_mBAHCuQW4_2),.dout(w_dff_B_wa7If9a09_2),.clk(gclk));
	jdff dff_B_ZPzbgEgX5_2(.din(w_dff_B_wa7If9a09_2),.dout(w_dff_B_ZPzbgEgX5_2),.clk(gclk));
	jdff dff_B_GGYKYHp36_2(.din(w_dff_B_ZPzbgEgX5_2),.dout(w_dff_B_GGYKYHp36_2),.clk(gclk));
	jdff dff_B_hki1wbsE5_2(.din(w_dff_B_GGYKYHp36_2),.dout(w_dff_B_hki1wbsE5_2),.clk(gclk));
	jdff dff_B_vSXcGfHH8_2(.din(w_dff_B_hki1wbsE5_2),.dout(w_dff_B_vSXcGfHH8_2),.clk(gclk));
	jdff dff_B_gRcf7Shg7_2(.din(w_dff_B_vSXcGfHH8_2),.dout(w_dff_B_gRcf7Shg7_2),.clk(gclk));
	jdff dff_B_YUEU3PB34_2(.din(w_dff_B_gRcf7Shg7_2),.dout(w_dff_B_YUEU3PB34_2),.clk(gclk));
	jdff dff_B_v7IBVsMS7_2(.din(w_dff_B_YUEU3PB34_2),.dout(w_dff_B_v7IBVsMS7_2),.clk(gclk));
	jdff dff_B_jXEB89iI1_2(.din(w_dff_B_v7IBVsMS7_2),.dout(w_dff_B_jXEB89iI1_2),.clk(gclk));
	jdff dff_B_4cQLnrIp3_2(.din(w_dff_B_jXEB89iI1_2),.dout(w_dff_B_4cQLnrIp3_2),.clk(gclk));
	jdff dff_B_k2y5Llhv9_2(.din(w_dff_B_4cQLnrIp3_2),.dout(w_dff_B_k2y5Llhv9_2),.clk(gclk));
	jdff dff_B_jzle25lS0_2(.din(w_dff_B_k2y5Llhv9_2),.dout(w_dff_B_jzle25lS0_2),.clk(gclk));
	jdff dff_B_7j9wF6AW7_2(.din(w_dff_B_jzle25lS0_2),.dout(w_dff_B_7j9wF6AW7_2),.clk(gclk));
	jdff dff_B_rSElkkp40_2(.din(w_dff_B_7j9wF6AW7_2),.dout(w_dff_B_rSElkkp40_2),.clk(gclk));
	jdff dff_B_oMDpZC6N7_2(.din(w_dff_B_rSElkkp40_2),.dout(w_dff_B_oMDpZC6N7_2),.clk(gclk));
	jdff dff_B_nlzTKguN6_2(.din(w_dff_B_oMDpZC6N7_2),.dout(w_dff_B_nlzTKguN6_2),.clk(gclk));
	jdff dff_B_tAEciqjq9_2(.din(w_dff_B_nlzTKguN6_2),.dout(w_dff_B_tAEciqjq9_2),.clk(gclk));
	jdff dff_B_yrwraxs34_2(.din(w_dff_B_tAEciqjq9_2),.dout(w_dff_B_yrwraxs34_2),.clk(gclk));
	jdff dff_B_gOCfkhlM7_2(.din(w_dff_B_yrwraxs34_2),.dout(w_dff_B_gOCfkhlM7_2),.clk(gclk));
	jdff dff_B_SsRb6lpj6_2(.din(w_dff_B_gOCfkhlM7_2),.dout(w_dff_B_SsRb6lpj6_2),.clk(gclk));
	jdff dff_B_2R8NMV0v3_2(.din(n1574),.dout(w_dff_B_2R8NMV0v3_2),.clk(gclk));
	jdff dff_B_pagIvr6A9_1(.din(n1572),.dout(w_dff_B_pagIvr6A9_1),.clk(gclk));
	jdff dff_B_TLuVNcfx0_2(.din(n1507),.dout(w_dff_B_TLuVNcfx0_2),.clk(gclk));
	jdff dff_B_WRy6xeMn3_2(.din(w_dff_B_TLuVNcfx0_2),.dout(w_dff_B_WRy6xeMn3_2),.clk(gclk));
	jdff dff_B_91c7I6DH5_2(.din(w_dff_B_WRy6xeMn3_2),.dout(w_dff_B_91c7I6DH5_2),.clk(gclk));
	jdff dff_B_aBp54Wtv4_2(.din(w_dff_B_91c7I6DH5_2),.dout(w_dff_B_aBp54Wtv4_2),.clk(gclk));
	jdff dff_B_CODpvkFf0_2(.din(w_dff_B_aBp54Wtv4_2),.dout(w_dff_B_CODpvkFf0_2),.clk(gclk));
	jdff dff_B_1iRxiGVT0_2(.din(w_dff_B_CODpvkFf0_2),.dout(w_dff_B_1iRxiGVT0_2),.clk(gclk));
	jdff dff_B_vdQYW4Hw1_2(.din(w_dff_B_1iRxiGVT0_2),.dout(w_dff_B_vdQYW4Hw1_2),.clk(gclk));
	jdff dff_B_reTqCqZp4_2(.din(w_dff_B_vdQYW4Hw1_2),.dout(w_dff_B_reTqCqZp4_2),.clk(gclk));
	jdff dff_B_voqJWS125_2(.din(w_dff_B_reTqCqZp4_2),.dout(w_dff_B_voqJWS125_2),.clk(gclk));
	jdff dff_B_yl3ejYsE6_2(.din(w_dff_B_voqJWS125_2),.dout(w_dff_B_yl3ejYsE6_2),.clk(gclk));
	jdff dff_B_kjCn1hoO6_2(.din(w_dff_B_yl3ejYsE6_2),.dout(w_dff_B_kjCn1hoO6_2),.clk(gclk));
	jdff dff_B_yuqiEWKI0_2(.din(w_dff_B_kjCn1hoO6_2),.dout(w_dff_B_yuqiEWKI0_2),.clk(gclk));
	jdff dff_B_0HFGYiWl6_2(.din(w_dff_B_yuqiEWKI0_2),.dout(w_dff_B_0HFGYiWl6_2),.clk(gclk));
	jdff dff_B_oP3nAfxX5_2(.din(w_dff_B_0HFGYiWl6_2),.dout(w_dff_B_oP3nAfxX5_2),.clk(gclk));
	jdff dff_B_08jXME4B6_2(.din(w_dff_B_oP3nAfxX5_2),.dout(w_dff_B_08jXME4B6_2),.clk(gclk));
	jdff dff_B_GMloJzhW1_2(.din(w_dff_B_08jXME4B6_2),.dout(w_dff_B_GMloJzhW1_2),.clk(gclk));
	jdff dff_B_pa8eGOHw3_2(.din(w_dff_B_GMloJzhW1_2),.dout(w_dff_B_pa8eGOHw3_2),.clk(gclk));
	jdff dff_B_aGfszCib8_2(.din(w_dff_B_pa8eGOHw3_2),.dout(w_dff_B_aGfszCib8_2),.clk(gclk));
	jdff dff_B_B2uFpXqJ9_2(.din(w_dff_B_aGfszCib8_2),.dout(w_dff_B_B2uFpXqJ9_2),.clk(gclk));
	jdff dff_B_h0qAKFFr9_2(.din(w_dff_B_B2uFpXqJ9_2),.dout(w_dff_B_h0qAKFFr9_2),.clk(gclk));
	jdff dff_B_m71BTlAj1_2(.din(w_dff_B_h0qAKFFr9_2),.dout(w_dff_B_m71BTlAj1_2),.clk(gclk));
	jdff dff_B_jamaZ3bo1_2(.din(w_dff_B_m71BTlAj1_2),.dout(w_dff_B_jamaZ3bo1_2),.clk(gclk));
	jdff dff_B_Tc0hrw154_2(.din(w_dff_B_jamaZ3bo1_2),.dout(w_dff_B_Tc0hrw154_2),.clk(gclk));
	jdff dff_B_WsdiyoMh8_2(.din(w_dff_B_Tc0hrw154_2),.dout(w_dff_B_WsdiyoMh8_2),.clk(gclk));
	jdff dff_B_dJOOY7kP7_2(.din(w_dff_B_WsdiyoMh8_2),.dout(w_dff_B_dJOOY7kP7_2),.clk(gclk));
	jdff dff_B_tpVz6Gsm7_2(.din(w_dff_B_dJOOY7kP7_2),.dout(w_dff_B_tpVz6Gsm7_2),.clk(gclk));
	jdff dff_B_55SGtvPf6_2(.din(w_dff_B_tpVz6Gsm7_2),.dout(w_dff_B_55SGtvPf6_2),.clk(gclk));
	jdff dff_B_AXwMpPAh1_2(.din(w_dff_B_55SGtvPf6_2),.dout(w_dff_B_AXwMpPAh1_2),.clk(gclk));
	jdff dff_B_0zhgQm5e9_2(.din(w_dff_B_AXwMpPAh1_2),.dout(w_dff_B_0zhgQm5e9_2),.clk(gclk));
	jdff dff_B_3qGD6MkH2_2(.din(w_dff_B_0zhgQm5e9_2),.dout(w_dff_B_3qGD6MkH2_2),.clk(gclk));
	jdff dff_B_IUUhIEmi9_2(.din(w_dff_B_3qGD6MkH2_2),.dout(w_dff_B_IUUhIEmi9_2),.clk(gclk));
	jdff dff_B_jQqc8zqU4_2(.din(w_dff_B_IUUhIEmi9_2),.dout(w_dff_B_jQqc8zqU4_2),.clk(gclk));
	jdff dff_B_829tdbsk5_2(.din(w_dff_B_jQqc8zqU4_2),.dout(w_dff_B_829tdbsk5_2),.clk(gclk));
	jdff dff_B_DTEQhiTy4_2(.din(w_dff_B_829tdbsk5_2),.dout(w_dff_B_DTEQhiTy4_2),.clk(gclk));
	jdff dff_B_lzgvobre2_2(.din(w_dff_B_DTEQhiTy4_2),.dout(w_dff_B_lzgvobre2_2),.clk(gclk));
	jdff dff_B_JUoSF68r3_2(.din(w_dff_B_lzgvobre2_2),.dout(w_dff_B_JUoSF68r3_2),.clk(gclk));
	jdff dff_B_XK4FhS402_2(.din(w_dff_B_JUoSF68r3_2),.dout(w_dff_B_XK4FhS402_2),.clk(gclk));
	jdff dff_B_6mmEAo6i4_2(.din(w_dff_B_XK4FhS402_2),.dout(w_dff_B_6mmEAo6i4_2),.clk(gclk));
	jdff dff_B_4CzgkvPs3_2(.din(w_dff_B_6mmEAo6i4_2),.dout(w_dff_B_4CzgkvPs3_2),.clk(gclk));
	jdff dff_B_K41MyTbU4_1(.din(n1508),.dout(w_dff_B_K41MyTbU4_1),.clk(gclk));
	jdff dff_B_TyK5dQqj5_2(.din(n1436),.dout(w_dff_B_TyK5dQqj5_2),.clk(gclk));
	jdff dff_B_arrXisRy6_2(.din(w_dff_B_TyK5dQqj5_2),.dout(w_dff_B_arrXisRy6_2),.clk(gclk));
	jdff dff_B_Zk13VLht1_2(.din(w_dff_B_arrXisRy6_2),.dout(w_dff_B_Zk13VLht1_2),.clk(gclk));
	jdff dff_B_TW86E0Zv5_2(.din(w_dff_B_Zk13VLht1_2),.dout(w_dff_B_TW86E0Zv5_2),.clk(gclk));
	jdff dff_B_9pVyEPLW4_2(.din(w_dff_B_TW86E0Zv5_2),.dout(w_dff_B_9pVyEPLW4_2),.clk(gclk));
	jdff dff_B_7s6xVT6I4_2(.din(w_dff_B_9pVyEPLW4_2),.dout(w_dff_B_7s6xVT6I4_2),.clk(gclk));
	jdff dff_B_0uIMJlZc9_2(.din(w_dff_B_7s6xVT6I4_2),.dout(w_dff_B_0uIMJlZc9_2),.clk(gclk));
	jdff dff_B_AEQteULq6_2(.din(w_dff_B_0uIMJlZc9_2),.dout(w_dff_B_AEQteULq6_2),.clk(gclk));
	jdff dff_B_mQgpQWQO8_2(.din(w_dff_B_AEQteULq6_2),.dout(w_dff_B_mQgpQWQO8_2),.clk(gclk));
	jdff dff_B_Du1S8MxW8_2(.din(w_dff_B_mQgpQWQO8_2),.dout(w_dff_B_Du1S8MxW8_2),.clk(gclk));
	jdff dff_B_snbtd5uG4_2(.din(w_dff_B_Du1S8MxW8_2),.dout(w_dff_B_snbtd5uG4_2),.clk(gclk));
	jdff dff_B_R7HZpIr20_2(.din(w_dff_B_snbtd5uG4_2),.dout(w_dff_B_R7HZpIr20_2),.clk(gclk));
	jdff dff_B_QGdQG0sN8_2(.din(w_dff_B_R7HZpIr20_2),.dout(w_dff_B_QGdQG0sN8_2),.clk(gclk));
	jdff dff_B_1JuYYxyY3_2(.din(w_dff_B_QGdQG0sN8_2),.dout(w_dff_B_1JuYYxyY3_2),.clk(gclk));
	jdff dff_B_69TUTZL13_2(.din(w_dff_B_1JuYYxyY3_2),.dout(w_dff_B_69TUTZL13_2),.clk(gclk));
	jdff dff_B_eWu280fD2_2(.din(w_dff_B_69TUTZL13_2),.dout(w_dff_B_eWu280fD2_2),.clk(gclk));
	jdff dff_B_OqfR5k8g6_2(.din(w_dff_B_eWu280fD2_2),.dout(w_dff_B_OqfR5k8g6_2),.clk(gclk));
	jdff dff_B_Sesxpo9h3_2(.din(w_dff_B_OqfR5k8g6_2),.dout(w_dff_B_Sesxpo9h3_2),.clk(gclk));
	jdff dff_B_ozzNEXzh1_2(.din(w_dff_B_Sesxpo9h3_2),.dout(w_dff_B_ozzNEXzh1_2),.clk(gclk));
	jdff dff_B_uDazpirA8_2(.din(w_dff_B_ozzNEXzh1_2),.dout(w_dff_B_uDazpirA8_2),.clk(gclk));
	jdff dff_B_L6QxvCDs1_2(.din(w_dff_B_uDazpirA8_2),.dout(w_dff_B_L6QxvCDs1_2),.clk(gclk));
	jdff dff_B_ThLEIJR14_2(.din(w_dff_B_L6QxvCDs1_2),.dout(w_dff_B_ThLEIJR14_2),.clk(gclk));
	jdff dff_B_oo2V7gSP7_2(.din(w_dff_B_ThLEIJR14_2),.dout(w_dff_B_oo2V7gSP7_2),.clk(gclk));
	jdff dff_B_eJ8H1CBG3_2(.din(w_dff_B_oo2V7gSP7_2),.dout(w_dff_B_eJ8H1CBG3_2),.clk(gclk));
	jdff dff_B_SvzLXKei0_2(.din(w_dff_B_eJ8H1CBG3_2),.dout(w_dff_B_SvzLXKei0_2),.clk(gclk));
	jdff dff_B_kntGFaS84_2(.din(w_dff_B_SvzLXKei0_2),.dout(w_dff_B_kntGFaS84_2),.clk(gclk));
	jdff dff_B_KCi92yq28_2(.din(w_dff_B_kntGFaS84_2),.dout(w_dff_B_KCi92yq28_2),.clk(gclk));
	jdff dff_B_mYEcX1I12_2(.din(w_dff_B_KCi92yq28_2),.dout(w_dff_B_mYEcX1I12_2),.clk(gclk));
	jdff dff_B_LZNvlh2l6_2(.din(w_dff_B_mYEcX1I12_2),.dout(w_dff_B_LZNvlh2l6_2),.clk(gclk));
	jdff dff_B_AmcbLqlN5_2(.din(w_dff_B_LZNvlh2l6_2),.dout(w_dff_B_AmcbLqlN5_2),.clk(gclk));
	jdff dff_B_avgG7PRt1_2(.din(w_dff_B_AmcbLqlN5_2),.dout(w_dff_B_avgG7PRt1_2),.clk(gclk));
	jdff dff_B_cGP2vjTw7_2(.din(w_dff_B_avgG7PRt1_2),.dout(w_dff_B_cGP2vjTw7_2),.clk(gclk));
	jdff dff_B_Qc3ocyp11_2(.din(w_dff_B_cGP2vjTw7_2),.dout(w_dff_B_Qc3ocyp11_2),.clk(gclk));
	jdff dff_B_6Xsy4sUD5_2(.din(w_dff_B_Qc3ocyp11_2),.dout(w_dff_B_6Xsy4sUD5_2),.clk(gclk));
	jdff dff_B_O80VdUpm7_2(.din(w_dff_B_6Xsy4sUD5_2),.dout(w_dff_B_O80VdUpm7_2),.clk(gclk));
	jdff dff_B_itcEa49g7_2(.din(w_dff_B_O80VdUpm7_2),.dout(w_dff_B_itcEa49g7_2),.clk(gclk));
	jdff dff_B_bYfsVfi42_2(.din(n1475),.dout(w_dff_B_bYfsVfi42_2),.clk(gclk));
	jdff dff_B_3ivT3rTn6_1(.din(n1437),.dout(w_dff_B_3ivT3rTn6_1),.clk(gclk));
	jdff dff_B_flQf7tPn4_2(.din(n1358),.dout(w_dff_B_flQf7tPn4_2),.clk(gclk));
	jdff dff_B_56Pqgc8c1_2(.din(w_dff_B_flQf7tPn4_2),.dout(w_dff_B_56Pqgc8c1_2),.clk(gclk));
	jdff dff_B_7dtkclOw9_2(.din(w_dff_B_56Pqgc8c1_2),.dout(w_dff_B_7dtkclOw9_2),.clk(gclk));
	jdff dff_B_KlDK33Mf7_2(.din(w_dff_B_7dtkclOw9_2),.dout(w_dff_B_KlDK33Mf7_2),.clk(gclk));
	jdff dff_B_eHFgj4Ve3_2(.din(w_dff_B_KlDK33Mf7_2),.dout(w_dff_B_eHFgj4Ve3_2),.clk(gclk));
	jdff dff_B_d7Wy6wTi6_2(.din(w_dff_B_eHFgj4Ve3_2),.dout(w_dff_B_d7Wy6wTi6_2),.clk(gclk));
	jdff dff_B_D0d9A9qJ6_2(.din(w_dff_B_d7Wy6wTi6_2),.dout(w_dff_B_D0d9A9qJ6_2),.clk(gclk));
	jdff dff_B_P6mjiWLb0_2(.din(w_dff_B_D0d9A9qJ6_2),.dout(w_dff_B_P6mjiWLb0_2),.clk(gclk));
	jdff dff_B_tBCFtUkA8_2(.din(w_dff_B_P6mjiWLb0_2),.dout(w_dff_B_tBCFtUkA8_2),.clk(gclk));
	jdff dff_B_FBTOGR5y4_2(.din(w_dff_B_tBCFtUkA8_2),.dout(w_dff_B_FBTOGR5y4_2),.clk(gclk));
	jdff dff_B_V34flryK0_2(.din(w_dff_B_FBTOGR5y4_2),.dout(w_dff_B_V34flryK0_2),.clk(gclk));
	jdff dff_B_wdQgBuBB6_2(.din(w_dff_B_V34flryK0_2),.dout(w_dff_B_wdQgBuBB6_2),.clk(gclk));
	jdff dff_B_Hgs3QckX9_2(.din(w_dff_B_wdQgBuBB6_2),.dout(w_dff_B_Hgs3QckX9_2),.clk(gclk));
	jdff dff_B_sc8IGDxq3_2(.din(w_dff_B_Hgs3QckX9_2),.dout(w_dff_B_sc8IGDxq3_2),.clk(gclk));
	jdff dff_B_MwTtwYIr2_2(.din(w_dff_B_sc8IGDxq3_2),.dout(w_dff_B_MwTtwYIr2_2),.clk(gclk));
	jdff dff_B_EyFblM9y6_2(.din(w_dff_B_MwTtwYIr2_2),.dout(w_dff_B_EyFblM9y6_2),.clk(gclk));
	jdff dff_B_6MxbI05r8_2(.din(w_dff_B_EyFblM9y6_2),.dout(w_dff_B_6MxbI05r8_2),.clk(gclk));
	jdff dff_B_VVAKi3DV0_2(.din(w_dff_B_6MxbI05r8_2),.dout(w_dff_B_VVAKi3DV0_2),.clk(gclk));
	jdff dff_B_hk35RDvd0_2(.din(w_dff_B_VVAKi3DV0_2),.dout(w_dff_B_hk35RDvd0_2),.clk(gclk));
	jdff dff_B_PSrJARcw7_2(.din(w_dff_B_hk35RDvd0_2),.dout(w_dff_B_PSrJARcw7_2),.clk(gclk));
	jdff dff_B_owJ0xV6P1_2(.din(w_dff_B_PSrJARcw7_2),.dout(w_dff_B_owJ0xV6P1_2),.clk(gclk));
	jdff dff_B_376C6p1S1_2(.din(w_dff_B_owJ0xV6P1_2),.dout(w_dff_B_376C6p1S1_2),.clk(gclk));
	jdff dff_B_tQNyFucx4_2(.din(w_dff_B_376C6p1S1_2),.dout(w_dff_B_tQNyFucx4_2),.clk(gclk));
	jdff dff_B_Q4xVar3X0_2(.din(w_dff_B_tQNyFucx4_2),.dout(w_dff_B_Q4xVar3X0_2),.clk(gclk));
	jdff dff_B_a2AdSJ5e5_2(.din(w_dff_B_Q4xVar3X0_2),.dout(w_dff_B_a2AdSJ5e5_2),.clk(gclk));
	jdff dff_B_rJHnmdi38_2(.din(w_dff_B_a2AdSJ5e5_2),.dout(w_dff_B_rJHnmdi38_2),.clk(gclk));
	jdff dff_B_ZgWZNZGs6_2(.din(w_dff_B_rJHnmdi38_2),.dout(w_dff_B_ZgWZNZGs6_2),.clk(gclk));
	jdff dff_B_VkjFSMyx0_2(.din(w_dff_B_ZgWZNZGs6_2),.dout(w_dff_B_VkjFSMyx0_2),.clk(gclk));
	jdff dff_B_mMgjSKlN0_2(.din(w_dff_B_VkjFSMyx0_2),.dout(w_dff_B_mMgjSKlN0_2),.clk(gclk));
	jdff dff_B_2cmTMOFd7_2(.din(w_dff_B_mMgjSKlN0_2),.dout(w_dff_B_2cmTMOFd7_2),.clk(gclk));
	jdff dff_B_ckOJNAx06_2(.din(w_dff_B_2cmTMOFd7_2),.dout(w_dff_B_ckOJNAx06_2),.clk(gclk));
	jdff dff_B_Zvq4qjqE0_2(.din(w_dff_B_ckOJNAx06_2),.dout(w_dff_B_Zvq4qjqE0_2),.clk(gclk));
	jdff dff_B_5S7Cx1Wo0_2(.din(w_dff_B_Zvq4qjqE0_2),.dout(w_dff_B_5S7Cx1Wo0_2),.clk(gclk));
	jdff dff_B_eRYndxZQ9_2(.din(n1397),.dout(w_dff_B_eRYndxZQ9_2),.clk(gclk));
	jdff dff_B_r1QgCYWE8_1(.din(n1359),.dout(w_dff_B_r1QgCYWE8_1),.clk(gclk));
	jdff dff_B_mAp5Wr2U3_2(.din(n1273),.dout(w_dff_B_mAp5Wr2U3_2),.clk(gclk));
	jdff dff_B_jZRyMvmh3_2(.din(w_dff_B_mAp5Wr2U3_2),.dout(w_dff_B_jZRyMvmh3_2),.clk(gclk));
	jdff dff_B_xAe6ydeR9_2(.din(w_dff_B_jZRyMvmh3_2),.dout(w_dff_B_xAe6ydeR9_2),.clk(gclk));
	jdff dff_B_9EdJwgCh9_2(.din(w_dff_B_xAe6ydeR9_2),.dout(w_dff_B_9EdJwgCh9_2),.clk(gclk));
	jdff dff_B_vdzOl8vN5_2(.din(w_dff_B_9EdJwgCh9_2),.dout(w_dff_B_vdzOl8vN5_2),.clk(gclk));
	jdff dff_B_eqZXP6sM3_2(.din(w_dff_B_vdzOl8vN5_2),.dout(w_dff_B_eqZXP6sM3_2),.clk(gclk));
	jdff dff_B_4D0HCNlm1_2(.din(w_dff_B_eqZXP6sM3_2),.dout(w_dff_B_4D0HCNlm1_2),.clk(gclk));
	jdff dff_B_6UWdwD3b1_2(.din(w_dff_B_4D0HCNlm1_2),.dout(w_dff_B_6UWdwD3b1_2),.clk(gclk));
	jdff dff_B_JAXKTocg6_2(.din(w_dff_B_6UWdwD3b1_2),.dout(w_dff_B_JAXKTocg6_2),.clk(gclk));
	jdff dff_B_38PoEDjK5_2(.din(w_dff_B_JAXKTocg6_2),.dout(w_dff_B_38PoEDjK5_2),.clk(gclk));
	jdff dff_B_FDHm8uDc8_2(.din(w_dff_B_38PoEDjK5_2),.dout(w_dff_B_FDHm8uDc8_2),.clk(gclk));
	jdff dff_B_DER76iIo3_2(.din(w_dff_B_FDHm8uDc8_2),.dout(w_dff_B_DER76iIo3_2),.clk(gclk));
	jdff dff_B_8lS6xrSr4_2(.din(w_dff_B_DER76iIo3_2),.dout(w_dff_B_8lS6xrSr4_2),.clk(gclk));
	jdff dff_B_4XGQjpMt0_2(.din(w_dff_B_8lS6xrSr4_2),.dout(w_dff_B_4XGQjpMt0_2),.clk(gclk));
	jdff dff_B_tOyO4qrW9_2(.din(w_dff_B_4XGQjpMt0_2),.dout(w_dff_B_tOyO4qrW9_2),.clk(gclk));
	jdff dff_B_R1BRX1oa3_2(.din(w_dff_B_tOyO4qrW9_2),.dout(w_dff_B_R1BRX1oa3_2),.clk(gclk));
	jdff dff_B_l9io95j56_2(.din(w_dff_B_R1BRX1oa3_2),.dout(w_dff_B_l9io95j56_2),.clk(gclk));
	jdff dff_B_U2nah3FP2_2(.din(w_dff_B_l9io95j56_2),.dout(w_dff_B_U2nah3FP2_2),.clk(gclk));
	jdff dff_B_ICOJaBic1_2(.din(w_dff_B_U2nah3FP2_2),.dout(w_dff_B_ICOJaBic1_2),.clk(gclk));
	jdff dff_B_u6t4UeYS9_2(.din(w_dff_B_ICOJaBic1_2),.dout(w_dff_B_u6t4UeYS9_2),.clk(gclk));
	jdff dff_B_iyr9dA2w2_2(.din(w_dff_B_u6t4UeYS9_2),.dout(w_dff_B_iyr9dA2w2_2),.clk(gclk));
	jdff dff_B_Gc4LD6193_2(.din(w_dff_B_iyr9dA2w2_2),.dout(w_dff_B_Gc4LD6193_2),.clk(gclk));
	jdff dff_B_PJB8swyl7_2(.din(w_dff_B_Gc4LD6193_2),.dout(w_dff_B_PJB8swyl7_2),.clk(gclk));
	jdff dff_B_W3BSKrt41_2(.din(w_dff_B_PJB8swyl7_2),.dout(w_dff_B_W3BSKrt41_2),.clk(gclk));
	jdff dff_B_nnKpUWXO7_2(.din(w_dff_B_W3BSKrt41_2),.dout(w_dff_B_nnKpUWXO7_2),.clk(gclk));
	jdff dff_B_44aVBxuU2_2(.din(w_dff_B_nnKpUWXO7_2),.dout(w_dff_B_44aVBxuU2_2),.clk(gclk));
	jdff dff_B_gllUJLha2_2(.din(w_dff_B_44aVBxuU2_2),.dout(w_dff_B_gllUJLha2_2),.clk(gclk));
	jdff dff_B_JofmrGE47_2(.din(w_dff_B_gllUJLha2_2),.dout(w_dff_B_JofmrGE47_2),.clk(gclk));
	jdff dff_B_k60LU9g95_2(.din(w_dff_B_JofmrGE47_2),.dout(w_dff_B_k60LU9g95_2),.clk(gclk));
	jdff dff_B_kFyMKoK27_2(.din(w_dff_B_k60LU9g95_2),.dout(w_dff_B_kFyMKoK27_2),.clk(gclk));
	jdff dff_B_bBFQ8uv53_2(.din(n1312),.dout(w_dff_B_bBFQ8uv53_2),.clk(gclk));
	jdff dff_B_wagfIO683_1(.din(n1274),.dout(w_dff_B_wagfIO683_1),.clk(gclk));
	jdff dff_B_PdHUiMdJ8_2(.din(n1183),.dout(w_dff_B_PdHUiMdJ8_2),.clk(gclk));
	jdff dff_B_UpRxfvD89_2(.din(w_dff_B_PdHUiMdJ8_2),.dout(w_dff_B_UpRxfvD89_2),.clk(gclk));
	jdff dff_B_tkGe4RU20_2(.din(w_dff_B_UpRxfvD89_2),.dout(w_dff_B_tkGe4RU20_2),.clk(gclk));
	jdff dff_B_wczrDmUN1_2(.din(w_dff_B_tkGe4RU20_2),.dout(w_dff_B_wczrDmUN1_2),.clk(gclk));
	jdff dff_B_oBmvKOG43_2(.din(w_dff_B_wczrDmUN1_2),.dout(w_dff_B_oBmvKOG43_2),.clk(gclk));
	jdff dff_B_IEimpLLb4_2(.din(w_dff_B_oBmvKOG43_2),.dout(w_dff_B_IEimpLLb4_2),.clk(gclk));
	jdff dff_B_RiZfGMyU6_2(.din(w_dff_B_IEimpLLb4_2),.dout(w_dff_B_RiZfGMyU6_2),.clk(gclk));
	jdff dff_B_dJafIPej1_2(.din(w_dff_B_RiZfGMyU6_2),.dout(w_dff_B_dJafIPej1_2),.clk(gclk));
	jdff dff_B_PA2s1AEB4_2(.din(w_dff_B_dJafIPej1_2),.dout(w_dff_B_PA2s1AEB4_2),.clk(gclk));
	jdff dff_B_3vqY1THw9_2(.din(w_dff_B_PA2s1AEB4_2),.dout(w_dff_B_3vqY1THw9_2),.clk(gclk));
	jdff dff_B_1dOSfdRo8_2(.din(w_dff_B_3vqY1THw9_2),.dout(w_dff_B_1dOSfdRo8_2),.clk(gclk));
	jdff dff_B_hWh6G7eG3_2(.din(w_dff_B_1dOSfdRo8_2),.dout(w_dff_B_hWh6G7eG3_2),.clk(gclk));
	jdff dff_B_LuGowNgP7_2(.din(w_dff_B_hWh6G7eG3_2),.dout(w_dff_B_LuGowNgP7_2),.clk(gclk));
	jdff dff_B_hMAT3ppX4_2(.din(w_dff_B_LuGowNgP7_2),.dout(w_dff_B_hMAT3ppX4_2),.clk(gclk));
	jdff dff_B_hN2Og05J4_2(.din(w_dff_B_hMAT3ppX4_2),.dout(w_dff_B_hN2Og05J4_2),.clk(gclk));
	jdff dff_B_GFGmnGVU7_2(.din(w_dff_B_hN2Og05J4_2),.dout(w_dff_B_GFGmnGVU7_2),.clk(gclk));
	jdff dff_B_D5IPn25S0_2(.din(w_dff_B_GFGmnGVU7_2),.dout(w_dff_B_D5IPn25S0_2),.clk(gclk));
	jdff dff_B_vYPnYFYf5_2(.din(w_dff_B_D5IPn25S0_2),.dout(w_dff_B_vYPnYFYf5_2),.clk(gclk));
	jdff dff_B_eN7zp82a4_2(.din(w_dff_B_vYPnYFYf5_2),.dout(w_dff_B_eN7zp82a4_2),.clk(gclk));
	jdff dff_B_vb6Wdhxy4_2(.din(w_dff_B_eN7zp82a4_2),.dout(w_dff_B_vb6Wdhxy4_2),.clk(gclk));
	jdff dff_B_a0kRmkz70_2(.din(w_dff_B_vb6Wdhxy4_2),.dout(w_dff_B_a0kRmkz70_2),.clk(gclk));
	jdff dff_B_kQM9N60a5_2(.din(w_dff_B_a0kRmkz70_2),.dout(w_dff_B_kQM9N60a5_2),.clk(gclk));
	jdff dff_B_U7kB5AXn3_2(.din(w_dff_B_kQM9N60a5_2),.dout(w_dff_B_U7kB5AXn3_2),.clk(gclk));
	jdff dff_B_PKA8kakU5_2(.din(w_dff_B_U7kB5AXn3_2),.dout(w_dff_B_PKA8kakU5_2),.clk(gclk));
	jdff dff_B_1o7Vschu5_2(.din(w_dff_B_PKA8kakU5_2),.dout(w_dff_B_1o7Vschu5_2),.clk(gclk));
	jdff dff_B_BWgj89hY8_2(.din(w_dff_B_1o7Vschu5_2),.dout(w_dff_B_BWgj89hY8_2),.clk(gclk));
	jdff dff_B_IwuZxtfj9_2(.din(w_dff_B_BWgj89hY8_2),.dout(w_dff_B_IwuZxtfj9_2),.clk(gclk));
	jdff dff_B_rFjJMvLB6_2(.din(n1221),.dout(w_dff_B_rFjJMvLB6_2),.clk(gclk));
	jdff dff_B_xYPBzUfi5_1(.din(n1184),.dout(w_dff_B_xYPBzUfi5_1),.clk(gclk));
	jdff dff_B_ZlQXV9LP0_2(.din(n1079),.dout(w_dff_B_ZlQXV9LP0_2),.clk(gclk));
	jdff dff_B_Oor7oGdn0_2(.din(w_dff_B_ZlQXV9LP0_2),.dout(w_dff_B_Oor7oGdn0_2),.clk(gclk));
	jdff dff_B_Bh1fsua58_2(.din(w_dff_B_Oor7oGdn0_2),.dout(w_dff_B_Bh1fsua58_2),.clk(gclk));
	jdff dff_B_Jf3z8ZEo1_2(.din(w_dff_B_Bh1fsua58_2),.dout(w_dff_B_Jf3z8ZEo1_2),.clk(gclk));
	jdff dff_B_n9kziAFO6_2(.din(w_dff_B_Jf3z8ZEo1_2),.dout(w_dff_B_n9kziAFO6_2),.clk(gclk));
	jdff dff_B_D5EpSTut7_2(.din(w_dff_B_n9kziAFO6_2),.dout(w_dff_B_D5EpSTut7_2),.clk(gclk));
	jdff dff_B_rsGyHwG74_2(.din(w_dff_B_D5EpSTut7_2),.dout(w_dff_B_rsGyHwG74_2),.clk(gclk));
	jdff dff_B_rvyRnOh60_2(.din(w_dff_B_rsGyHwG74_2),.dout(w_dff_B_rvyRnOh60_2),.clk(gclk));
	jdff dff_B_fuDwmqRr1_2(.din(w_dff_B_rvyRnOh60_2),.dout(w_dff_B_fuDwmqRr1_2),.clk(gclk));
	jdff dff_B_Eq7Pr4C17_2(.din(w_dff_B_fuDwmqRr1_2),.dout(w_dff_B_Eq7Pr4C17_2),.clk(gclk));
	jdff dff_B_IJ0O3Nk72_2(.din(w_dff_B_Eq7Pr4C17_2),.dout(w_dff_B_IJ0O3Nk72_2),.clk(gclk));
	jdff dff_B_KRvi5V9U8_2(.din(w_dff_B_IJ0O3Nk72_2),.dout(w_dff_B_KRvi5V9U8_2),.clk(gclk));
	jdff dff_B_cukbiTFI2_2(.din(w_dff_B_KRvi5V9U8_2),.dout(w_dff_B_cukbiTFI2_2),.clk(gclk));
	jdff dff_B_pHA1L4m16_2(.din(w_dff_B_cukbiTFI2_2),.dout(w_dff_B_pHA1L4m16_2),.clk(gclk));
	jdff dff_B_jWlWgwqZ9_2(.din(w_dff_B_pHA1L4m16_2),.dout(w_dff_B_jWlWgwqZ9_2),.clk(gclk));
	jdff dff_B_onhZauR79_2(.din(w_dff_B_jWlWgwqZ9_2),.dout(w_dff_B_onhZauR79_2),.clk(gclk));
	jdff dff_B_U8cur0Jw2_2(.din(w_dff_B_onhZauR79_2),.dout(w_dff_B_U8cur0Jw2_2),.clk(gclk));
	jdff dff_B_jnn794fg4_2(.din(w_dff_B_U8cur0Jw2_2),.dout(w_dff_B_jnn794fg4_2),.clk(gclk));
	jdff dff_B_hxT1HbQd3_2(.din(w_dff_B_jnn794fg4_2),.dout(w_dff_B_hxT1HbQd3_2),.clk(gclk));
	jdff dff_B_Rv0JryFq4_2(.din(w_dff_B_hxT1HbQd3_2),.dout(w_dff_B_Rv0JryFq4_2),.clk(gclk));
	jdff dff_B_k4bGixr26_2(.din(w_dff_B_Rv0JryFq4_2),.dout(w_dff_B_k4bGixr26_2),.clk(gclk));
	jdff dff_B_7CKXMnQ41_2(.din(w_dff_B_k4bGixr26_2),.dout(w_dff_B_7CKXMnQ41_2),.clk(gclk));
	jdff dff_B_TsgmmHrT5_2(.din(w_dff_B_7CKXMnQ41_2),.dout(w_dff_B_TsgmmHrT5_2),.clk(gclk));
	jdff dff_B_czjghiQe6_2(.din(w_dff_B_TsgmmHrT5_2),.dout(w_dff_B_czjghiQe6_2),.clk(gclk));
	jdff dff_B_RuQq9Eub5_2(.din(n1123),.dout(w_dff_B_RuQq9Eub5_2),.clk(gclk));
	jdff dff_B_pcewXHOL5_1(.din(n1080),.dout(w_dff_B_pcewXHOL5_1),.clk(gclk));
	jdff dff_B_V8XIUyyD9_2(.din(n981),.dout(w_dff_B_V8XIUyyD9_2),.clk(gclk));
	jdff dff_B_mnaP1wgb4_2(.din(w_dff_B_V8XIUyyD9_2),.dout(w_dff_B_mnaP1wgb4_2),.clk(gclk));
	jdff dff_B_Zedg13GE5_2(.din(w_dff_B_mnaP1wgb4_2),.dout(w_dff_B_Zedg13GE5_2),.clk(gclk));
	jdff dff_B_D4JC1RTp0_2(.din(w_dff_B_Zedg13GE5_2),.dout(w_dff_B_D4JC1RTp0_2),.clk(gclk));
	jdff dff_B_Xx2gwmqm1_2(.din(w_dff_B_D4JC1RTp0_2),.dout(w_dff_B_Xx2gwmqm1_2),.clk(gclk));
	jdff dff_B_ZgY6m3Il0_2(.din(w_dff_B_Xx2gwmqm1_2),.dout(w_dff_B_ZgY6m3Il0_2),.clk(gclk));
	jdff dff_B_sgwBHFZn2_2(.din(w_dff_B_ZgY6m3Il0_2),.dout(w_dff_B_sgwBHFZn2_2),.clk(gclk));
	jdff dff_B_gINrAaA18_2(.din(w_dff_B_sgwBHFZn2_2),.dout(w_dff_B_gINrAaA18_2),.clk(gclk));
	jdff dff_B_0GOtKah77_2(.din(w_dff_B_gINrAaA18_2),.dout(w_dff_B_0GOtKah77_2),.clk(gclk));
	jdff dff_B_XuSJ6VgI9_2(.din(w_dff_B_0GOtKah77_2),.dout(w_dff_B_XuSJ6VgI9_2),.clk(gclk));
	jdff dff_B_gNIDXnNk7_2(.din(w_dff_B_XuSJ6VgI9_2),.dout(w_dff_B_gNIDXnNk7_2),.clk(gclk));
	jdff dff_B_VPNAr3yf0_2(.din(w_dff_B_gNIDXnNk7_2),.dout(w_dff_B_VPNAr3yf0_2),.clk(gclk));
	jdff dff_B_zyNYa4Zf0_2(.din(w_dff_B_VPNAr3yf0_2),.dout(w_dff_B_zyNYa4Zf0_2),.clk(gclk));
	jdff dff_B_lZ58jvSi3_2(.din(w_dff_B_zyNYa4Zf0_2),.dout(w_dff_B_lZ58jvSi3_2),.clk(gclk));
	jdff dff_B_JvaKCZre8_2(.din(w_dff_B_lZ58jvSi3_2),.dout(w_dff_B_JvaKCZre8_2),.clk(gclk));
	jdff dff_B_3vXwOkX01_2(.din(w_dff_B_JvaKCZre8_2),.dout(w_dff_B_3vXwOkX01_2),.clk(gclk));
	jdff dff_B_ixZqhkfJ8_2(.din(w_dff_B_3vXwOkX01_2),.dout(w_dff_B_ixZqhkfJ8_2),.clk(gclk));
	jdff dff_B_TaXcv2j70_2(.din(w_dff_B_ixZqhkfJ8_2),.dout(w_dff_B_TaXcv2j70_2),.clk(gclk));
	jdff dff_B_T7MIpknU2_2(.din(w_dff_B_TaXcv2j70_2),.dout(w_dff_B_T7MIpknU2_2),.clk(gclk));
	jdff dff_B_Dm1VWGbe4_2(.din(w_dff_B_T7MIpknU2_2),.dout(w_dff_B_Dm1VWGbe4_2),.clk(gclk));
	jdff dff_B_thbvFUV31_2(.din(w_dff_B_Dm1VWGbe4_2),.dout(w_dff_B_thbvFUV31_2),.clk(gclk));
	jdff dff_B_ao4BY8oo8_2(.din(n1018),.dout(w_dff_B_ao4BY8oo8_2),.clk(gclk));
	jdff dff_B_DZRvO2GV2_1(.din(n982),.dout(w_dff_B_DZRvO2GV2_1),.clk(gclk));
	jdff dff_B_tSSnxbXa8_2(.din(n876),.dout(w_dff_B_tSSnxbXa8_2),.clk(gclk));
	jdff dff_B_76t1DMNq6_2(.din(w_dff_B_tSSnxbXa8_2),.dout(w_dff_B_76t1DMNq6_2),.clk(gclk));
	jdff dff_B_6zSNXt7N2_2(.din(w_dff_B_76t1DMNq6_2),.dout(w_dff_B_6zSNXt7N2_2),.clk(gclk));
	jdff dff_B_fteipKbY6_2(.din(w_dff_B_6zSNXt7N2_2),.dout(w_dff_B_fteipKbY6_2),.clk(gclk));
	jdff dff_B_JfjY3Nog7_2(.din(w_dff_B_fteipKbY6_2),.dout(w_dff_B_JfjY3Nog7_2),.clk(gclk));
	jdff dff_B_KcNaJbXd4_2(.din(w_dff_B_JfjY3Nog7_2),.dout(w_dff_B_KcNaJbXd4_2),.clk(gclk));
	jdff dff_B_MDSMfXng6_2(.din(w_dff_B_KcNaJbXd4_2),.dout(w_dff_B_MDSMfXng6_2),.clk(gclk));
	jdff dff_B_f6n8BLPv9_2(.din(w_dff_B_MDSMfXng6_2),.dout(w_dff_B_f6n8BLPv9_2),.clk(gclk));
	jdff dff_B_3Wyhvwui8_2(.din(w_dff_B_f6n8BLPv9_2),.dout(w_dff_B_3Wyhvwui8_2),.clk(gclk));
	jdff dff_B_vvbHeEAI8_2(.din(w_dff_B_3Wyhvwui8_2),.dout(w_dff_B_vvbHeEAI8_2),.clk(gclk));
	jdff dff_B_SbSxcFOS3_2(.din(w_dff_B_vvbHeEAI8_2),.dout(w_dff_B_SbSxcFOS3_2),.clk(gclk));
	jdff dff_B_kZzSmu0J0_2(.din(w_dff_B_SbSxcFOS3_2),.dout(w_dff_B_kZzSmu0J0_2),.clk(gclk));
	jdff dff_B_vlvc2Jgj6_2(.din(w_dff_B_kZzSmu0J0_2),.dout(w_dff_B_vlvc2Jgj6_2),.clk(gclk));
	jdff dff_B_konWLJGr2_2(.din(w_dff_B_vlvc2Jgj6_2),.dout(w_dff_B_konWLJGr2_2),.clk(gclk));
	jdff dff_B_C7HhDz9u0_2(.din(w_dff_B_konWLJGr2_2),.dout(w_dff_B_C7HhDz9u0_2),.clk(gclk));
	jdff dff_B_izwclW5u7_2(.din(w_dff_B_C7HhDz9u0_2),.dout(w_dff_B_izwclW5u7_2),.clk(gclk));
	jdff dff_B_3BVpdZpE4_2(.din(w_dff_B_izwclW5u7_2),.dout(w_dff_B_3BVpdZpE4_2),.clk(gclk));
	jdff dff_B_DFyjm9Ys5_2(.din(w_dff_B_3BVpdZpE4_2),.dout(w_dff_B_DFyjm9Ys5_2),.clk(gclk));
	jdff dff_B_pK0UmoXy1_2(.din(n913),.dout(w_dff_B_pK0UmoXy1_2),.clk(gclk));
	jdff dff_B_FCxt0qPm9_1(.din(n877),.dout(w_dff_B_FCxt0qPm9_1),.clk(gclk));
	jdff dff_B_b34qV6ic3_2(.din(n777),.dout(w_dff_B_b34qV6ic3_2),.clk(gclk));
	jdff dff_B_4YiGYZGb6_2(.din(w_dff_B_b34qV6ic3_2),.dout(w_dff_B_4YiGYZGb6_2),.clk(gclk));
	jdff dff_B_B8NqnJWJ9_2(.din(w_dff_B_4YiGYZGb6_2),.dout(w_dff_B_B8NqnJWJ9_2),.clk(gclk));
	jdff dff_B_7HJiycvM3_2(.din(w_dff_B_B8NqnJWJ9_2),.dout(w_dff_B_7HJiycvM3_2),.clk(gclk));
	jdff dff_B_SzadATYM5_2(.din(w_dff_B_7HJiycvM3_2),.dout(w_dff_B_SzadATYM5_2),.clk(gclk));
	jdff dff_B_it1ksGdT6_2(.din(w_dff_B_SzadATYM5_2),.dout(w_dff_B_it1ksGdT6_2),.clk(gclk));
	jdff dff_B_RkngrY8w2_2(.din(w_dff_B_it1ksGdT6_2),.dout(w_dff_B_RkngrY8w2_2),.clk(gclk));
	jdff dff_B_iim0fEk80_2(.din(w_dff_B_RkngrY8w2_2),.dout(w_dff_B_iim0fEk80_2),.clk(gclk));
	jdff dff_B_NEwVDMBL5_2(.din(w_dff_B_iim0fEk80_2),.dout(w_dff_B_NEwVDMBL5_2),.clk(gclk));
	jdff dff_B_UVljeYQg8_2(.din(w_dff_B_NEwVDMBL5_2),.dout(w_dff_B_UVljeYQg8_2),.clk(gclk));
	jdff dff_B_vFP3rCBv2_2(.din(w_dff_B_UVljeYQg8_2),.dout(w_dff_B_vFP3rCBv2_2),.clk(gclk));
	jdff dff_B_Quv42M9X6_2(.din(w_dff_B_vFP3rCBv2_2),.dout(w_dff_B_Quv42M9X6_2),.clk(gclk));
	jdff dff_B_FYcs07zF6_2(.din(w_dff_B_Quv42M9X6_2),.dout(w_dff_B_FYcs07zF6_2),.clk(gclk));
	jdff dff_B_hh67WdTi6_2(.din(w_dff_B_FYcs07zF6_2),.dout(w_dff_B_hh67WdTi6_2),.clk(gclk));
	jdff dff_B_zmwDxNgR1_2(.din(w_dff_B_hh67WdTi6_2),.dout(w_dff_B_zmwDxNgR1_2),.clk(gclk));
	jdff dff_B_ybKDPPf21_2(.din(n807),.dout(w_dff_B_ybKDPPf21_2),.clk(gclk));
	jdff dff_B_GEBf26LN1_1(.din(n778),.dout(w_dff_B_GEBf26LN1_1),.clk(gclk));
	jdff dff_B_tquyCFwV4_2(.din(n684),.dout(w_dff_B_tquyCFwV4_2),.clk(gclk));
	jdff dff_B_eQMVtQdk8_2(.din(w_dff_B_tquyCFwV4_2),.dout(w_dff_B_eQMVtQdk8_2),.clk(gclk));
	jdff dff_B_lE8BO4Ak8_2(.din(w_dff_B_eQMVtQdk8_2),.dout(w_dff_B_lE8BO4Ak8_2),.clk(gclk));
	jdff dff_B_Z4DX1izX5_2(.din(w_dff_B_lE8BO4Ak8_2),.dout(w_dff_B_Z4DX1izX5_2),.clk(gclk));
	jdff dff_B_tu2IuUGn9_2(.din(w_dff_B_Z4DX1izX5_2),.dout(w_dff_B_tu2IuUGn9_2),.clk(gclk));
	jdff dff_B_hmkxXFmX5_2(.din(w_dff_B_tu2IuUGn9_2),.dout(w_dff_B_hmkxXFmX5_2),.clk(gclk));
	jdff dff_B_N7Rujm9g6_2(.din(w_dff_B_hmkxXFmX5_2),.dout(w_dff_B_N7Rujm9g6_2),.clk(gclk));
	jdff dff_B_PMYZG2Gs1_2(.din(w_dff_B_N7Rujm9g6_2),.dout(w_dff_B_PMYZG2Gs1_2),.clk(gclk));
	jdff dff_B_H6Hjpk5R6_2(.din(w_dff_B_PMYZG2Gs1_2),.dout(w_dff_B_H6Hjpk5R6_2),.clk(gclk));
	jdff dff_B_neCTmOi35_2(.din(w_dff_B_H6Hjpk5R6_2),.dout(w_dff_B_neCTmOi35_2),.clk(gclk));
	jdff dff_B_6IlgLLGe7_2(.din(w_dff_B_neCTmOi35_2),.dout(w_dff_B_6IlgLLGe7_2),.clk(gclk));
	jdff dff_B_bFjrIidG9_2(.din(w_dff_B_6IlgLLGe7_2),.dout(w_dff_B_bFjrIidG9_2),.clk(gclk));
	jdff dff_B_4IdKWKoN1_2(.din(n707),.dout(w_dff_B_4IdKWKoN1_2),.clk(gclk));
	jdff dff_B_cAHDlMdl3_1(.din(n685),.dout(w_dff_B_cAHDlMdl3_1),.clk(gclk));
	jdff dff_B_Tmwl9KId3_2(.din(n598),.dout(w_dff_B_Tmwl9KId3_2),.clk(gclk));
	jdff dff_B_kgt4KW890_2(.din(w_dff_B_Tmwl9KId3_2),.dout(w_dff_B_kgt4KW890_2),.clk(gclk));
	jdff dff_B_BH4dHiRb6_2(.din(w_dff_B_kgt4KW890_2),.dout(w_dff_B_BH4dHiRb6_2),.clk(gclk));
	jdff dff_B_2OqAu5By9_2(.din(w_dff_B_BH4dHiRb6_2),.dout(w_dff_B_2OqAu5By9_2),.clk(gclk));
	jdff dff_B_tTRWVKnj0_2(.din(w_dff_B_2OqAu5By9_2),.dout(w_dff_B_tTRWVKnj0_2),.clk(gclk));
	jdff dff_B_G2VAy9Qs4_2(.din(w_dff_B_tTRWVKnj0_2),.dout(w_dff_B_G2VAy9Qs4_2),.clk(gclk));
	jdff dff_B_yZ9mZk8C6_2(.din(w_dff_B_G2VAy9Qs4_2),.dout(w_dff_B_yZ9mZk8C6_2),.clk(gclk));
	jdff dff_B_B6uDATif7_2(.din(w_dff_B_yZ9mZk8C6_2),.dout(w_dff_B_B6uDATif7_2),.clk(gclk));
	jdff dff_B_9ozcuxUk2_2(.din(w_dff_B_B6uDATif7_2),.dout(w_dff_B_9ozcuxUk2_2),.clk(gclk));
	jdff dff_B_cHkEKdtp7_2(.din(n614),.dout(w_dff_B_cHkEKdtp7_2),.clk(gclk));
	jdff dff_B_pV3RM8kO6_2(.din(w_dff_B_cHkEKdtp7_2),.dout(w_dff_B_pV3RM8kO6_2),.clk(gclk));
	jdff dff_B_SSi1Nx618_1(.din(n599),.dout(w_dff_B_SSi1Nx618_1),.clk(gclk));
	jdff dff_B_PWgDQNB48_1(.din(w_dff_B_SSi1Nx618_1),.dout(w_dff_B_PWgDQNB48_1),.clk(gclk));
	jdff dff_B_eEqzv1yO6_1(.din(w_dff_B_PWgDQNB48_1),.dout(w_dff_B_eEqzv1yO6_1),.clk(gclk));
	jdff dff_B_NBSVDX3K8_1(.din(w_dff_B_eEqzv1yO6_1),.dout(w_dff_B_NBSVDX3K8_1),.clk(gclk));
	jdff dff_B_uawajdVm2_1(.din(w_dff_B_NBSVDX3K8_1),.dout(w_dff_B_uawajdVm2_1),.clk(gclk));
	jdff dff_B_nDYSgVV54_1(.din(w_dff_B_uawajdVm2_1),.dout(w_dff_B_nDYSgVV54_1),.clk(gclk));
	jdff dff_B_1ZmkyheE0_0(.din(n528),.dout(w_dff_B_1ZmkyheE0_0),.clk(gclk));
	jdff dff_B_n7fgtk1y8_0(.din(w_dff_B_1ZmkyheE0_0),.dout(w_dff_B_n7fgtk1y8_0),.clk(gclk));
	jdff dff_A_OlbhUUiF2_0(.dout(w_n527_0[0]),.din(w_dff_A_OlbhUUiF2_0),.clk(gclk));
	jdff dff_A_bUW1CBpB1_0(.dout(w_dff_A_OlbhUUiF2_0),.din(w_dff_A_bUW1CBpB1_0),.clk(gclk));
	jdff dff_A_ORLsOMXy6_0(.dout(w_dff_A_bUW1CBpB1_0),.din(w_dff_A_ORLsOMXy6_0),.clk(gclk));
	jdff dff_B_oQXcnDpm6_1(.din(n521),.dout(w_dff_B_oQXcnDpm6_1),.clk(gclk));
	jdff dff_A_TrtfMKBO0_0(.dout(w_n446_0[0]),.din(w_dff_A_TrtfMKBO0_0),.clk(gclk));
	jdff dff_A_TiCADdSY4_1(.dout(w_n446_0[1]),.din(w_dff_A_TiCADdSY4_1),.clk(gclk));
	jdff dff_A_hDjMxZIc3_1(.dout(w_dff_A_TiCADdSY4_1),.din(w_dff_A_hDjMxZIc3_1),.clk(gclk));
	jdff dff_A_TAdN2pcZ7_1(.dout(w_n519_0[1]),.din(w_dff_A_TAdN2pcZ7_1),.clk(gclk));
	jdff dff_A_TpDKr2Pl4_1(.dout(w_dff_A_TAdN2pcZ7_1),.din(w_dff_A_TpDKr2Pl4_1),.clk(gclk));
	jdff dff_A_q3D9U0OS2_1(.dout(w_dff_A_TpDKr2Pl4_1),.din(w_dff_A_q3D9U0OS2_1),.clk(gclk));
	jdff dff_A_tlK2ukNF8_1(.dout(w_dff_A_q3D9U0OS2_1),.din(w_dff_A_tlK2ukNF8_1),.clk(gclk));
	jdff dff_A_fmims8R39_1(.dout(w_dff_A_tlK2ukNF8_1),.din(w_dff_A_fmims8R39_1),.clk(gclk));
	jdff dff_A_rAkL1biL0_1(.dout(w_dff_A_fmims8R39_1),.din(w_dff_A_rAkL1biL0_1),.clk(gclk));
	jdff dff_B_ujHNKIta2_1(.din(n1760),.dout(w_dff_B_ujHNKIta2_1),.clk(gclk));
	jdff dff_A_KO0EuAWu9_1(.dout(w_n1728_0[1]),.din(w_dff_A_KO0EuAWu9_1),.clk(gclk));
	jdff dff_B_apJ5POHG4_1(.din(n1726),.dout(w_dff_B_apJ5POHG4_1),.clk(gclk));
	jdff dff_B_9xz2TAaz5_2(.din(n1684),.dout(w_dff_B_9xz2TAaz5_2),.clk(gclk));
	jdff dff_B_osJnFlgF0_2(.din(w_dff_B_9xz2TAaz5_2),.dout(w_dff_B_osJnFlgF0_2),.clk(gclk));
	jdff dff_B_oLKqF3Bw1_2(.din(w_dff_B_osJnFlgF0_2),.dout(w_dff_B_oLKqF3Bw1_2),.clk(gclk));
	jdff dff_B_q9exviJh9_2(.din(w_dff_B_oLKqF3Bw1_2),.dout(w_dff_B_q9exviJh9_2),.clk(gclk));
	jdff dff_B_MbBfWPil6_2(.din(w_dff_B_q9exviJh9_2),.dout(w_dff_B_MbBfWPil6_2),.clk(gclk));
	jdff dff_B_3CSI38gN1_2(.din(w_dff_B_MbBfWPil6_2),.dout(w_dff_B_3CSI38gN1_2),.clk(gclk));
	jdff dff_B_LjxN97AI1_2(.din(w_dff_B_3CSI38gN1_2),.dout(w_dff_B_LjxN97AI1_2),.clk(gclk));
	jdff dff_B_sdzPZ9Sw3_2(.din(w_dff_B_LjxN97AI1_2),.dout(w_dff_B_sdzPZ9Sw3_2),.clk(gclk));
	jdff dff_B_CPsJ53rU2_2(.din(w_dff_B_sdzPZ9Sw3_2),.dout(w_dff_B_CPsJ53rU2_2),.clk(gclk));
	jdff dff_B_la46kmkC6_2(.din(w_dff_B_CPsJ53rU2_2),.dout(w_dff_B_la46kmkC6_2),.clk(gclk));
	jdff dff_B_Y1iJcdN41_2(.din(w_dff_B_la46kmkC6_2),.dout(w_dff_B_Y1iJcdN41_2),.clk(gclk));
	jdff dff_B_mtLx5q6a1_2(.din(w_dff_B_Y1iJcdN41_2),.dout(w_dff_B_mtLx5q6a1_2),.clk(gclk));
	jdff dff_B_QPk1gBoU5_2(.din(w_dff_B_mtLx5q6a1_2),.dout(w_dff_B_QPk1gBoU5_2),.clk(gclk));
	jdff dff_B_GUxVZLTq6_2(.din(w_dff_B_QPk1gBoU5_2),.dout(w_dff_B_GUxVZLTq6_2),.clk(gclk));
	jdff dff_B_HxGEV71P4_2(.din(w_dff_B_GUxVZLTq6_2),.dout(w_dff_B_HxGEV71P4_2),.clk(gclk));
	jdff dff_B_UUFraiRB4_2(.din(w_dff_B_HxGEV71P4_2),.dout(w_dff_B_UUFraiRB4_2),.clk(gclk));
	jdff dff_B_Muyuscta5_2(.din(w_dff_B_UUFraiRB4_2),.dout(w_dff_B_Muyuscta5_2),.clk(gclk));
	jdff dff_B_LZdvBhbe2_2(.din(w_dff_B_Muyuscta5_2),.dout(w_dff_B_LZdvBhbe2_2),.clk(gclk));
	jdff dff_B_l2uNAhBI8_2(.din(w_dff_B_LZdvBhbe2_2),.dout(w_dff_B_l2uNAhBI8_2),.clk(gclk));
	jdff dff_B_FcDlXBvW1_2(.din(w_dff_B_l2uNAhBI8_2),.dout(w_dff_B_FcDlXBvW1_2),.clk(gclk));
	jdff dff_B_3fxmqe3e9_2(.din(w_dff_B_FcDlXBvW1_2),.dout(w_dff_B_3fxmqe3e9_2),.clk(gclk));
	jdff dff_B_yho9OXWh9_2(.din(w_dff_B_3fxmqe3e9_2),.dout(w_dff_B_yho9OXWh9_2),.clk(gclk));
	jdff dff_B_CBHIiu7x3_2(.din(w_dff_B_yho9OXWh9_2),.dout(w_dff_B_CBHIiu7x3_2),.clk(gclk));
	jdff dff_B_F1Bx0yKk5_2(.din(w_dff_B_CBHIiu7x3_2),.dout(w_dff_B_F1Bx0yKk5_2),.clk(gclk));
	jdff dff_B_e92sGs230_2(.din(w_dff_B_F1Bx0yKk5_2),.dout(w_dff_B_e92sGs230_2),.clk(gclk));
	jdff dff_B_DAIOBDHK2_2(.din(w_dff_B_e92sGs230_2),.dout(w_dff_B_DAIOBDHK2_2),.clk(gclk));
	jdff dff_B_1ovJIxFL4_2(.din(w_dff_B_DAIOBDHK2_2),.dout(w_dff_B_1ovJIxFL4_2),.clk(gclk));
	jdff dff_B_SWDD36d69_2(.din(w_dff_B_1ovJIxFL4_2),.dout(w_dff_B_SWDD36d69_2),.clk(gclk));
	jdff dff_B_7LPw1nqW3_2(.din(w_dff_B_SWDD36d69_2),.dout(w_dff_B_7LPw1nqW3_2),.clk(gclk));
	jdff dff_B_HyHON5LR1_2(.din(w_dff_B_7LPw1nqW3_2),.dout(w_dff_B_HyHON5LR1_2),.clk(gclk));
	jdff dff_B_Bvfy7t9D9_2(.din(w_dff_B_HyHON5LR1_2),.dout(w_dff_B_Bvfy7t9D9_2),.clk(gclk));
	jdff dff_B_En6pPMKo1_2(.din(w_dff_B_Bvfy7t9D9_2),.dout(w_dff_B_En6pPMKo1_2),.clk(gclk));
	jdff dff_B_o50OStId1_2(.din(w_dff_B_En6pPMKo1_2),.dout(w_dff_B_o50OStId1_2),.clk(gclk));
	jdff dff_B_3DSU8NNU4_2(.din(w_dff_B_o50OStId1_2),.dout(w_dff_B_3DSU8NNU4_2),.clk(gclk));
	jdff dff_B_Bd7DnAjV1_2(.din(w_dff_B_3DSU8NNU4_2),.dout(w_dff_B_Bd7DnAjV1_2),.clk(gclk));
	jdff dff_B_0Xxlr55z2_2(.din(w_dff_B_Bd7DnAjV1_2),.dout(w_dff_B_0Xxlr55z2_2),.clk(gclk));
	jdff dff_B_mm9FWPiT4_2(.din(w_dff_B_0Xxlr55z2_2),.dout(w_dff_B_mm9FWPiT4_2),.clk(gclk));
	jdff dff_B_qFm6eFQb1_2(.din(w_dff_B_mm9FWPiT4_2),.dout(w_dff_B_qFm6eFQb1_2),.clk(gclk));
	jdff dff_B_w9Maiqfx9_2(.din(w_dff_B_qFm6eFQb1_2),.dout(w_dff_B_w9Maiqfx9_2),.clk(gclk));
	jdff dff_B_nHcQtLIw8_2(.din(w_dff_B_w9Maiqfx9_2),.dout(w_dff_B_nHcQtLIw8_2),.clk(gclk));
	jdff dff_B_N0VRdw9b2_2(.din(w_dff_B_nHcQtLIw8_2),.dout(w_dff_B_N0VRdw9b2_2),.clk(gclk));
	jdff dff_B_DSx5GGT06_2(.din(w_dff_B_N0VRdw9b2_2),.dout(w_dff_B_DSx5GGT06_2),.clk(gclk));
	jdff dff_B_Qa1UIgWT5_2(.din(w_dff_B_DSx5GGT06_2),.dout(w_dff_B_Qa1UIgWT5_2),.clk(gclk));
	jdff dff_B_a1ZSYa9u1_2(.din(w_dff_B_Qa1UIgWT5_2),.dout(w_dff_B_a1ZSYa9u1_2),.clk(gclk));
	jdff dff_B_qhsrqwUt1_2(.din(w_dff_B_a1ZSYa9u1_2),.dout(w_dff_B_qhsrqwUt1_2),.clk(gclk));
	jdff dff_B_XK2uILrM8_2(.din(w_dff_B_qhsrqwUt1_2),.dout(w_dff_B_XK2uILrM8_2),.clk(gclk));
	jdff dff_B_2XFUkYcT6_2(.din(w_dff_B_XK2uILrM8_2),.dout(w_dff_B_2XFUkYcT6_2),.clk(gclk));
	jdff dff_B_xiZ0u1Xr4_2(.din(w_dff_B_2XFUkYcT6_2),.dout(w_dff_B_xiZ0u1Xr4_2),.clk(gclk));
	jdff dff_B_Md1qSbaj1_2(.din(w_dff_B_xiZ0u1Xr4_2),.dout(w_dff_B_Md1qSbaj1_2),.clk(gclk));
	jdff dff_B_GZgJyiDF4_2(.din(n1687),.dout(w_dff_B_GZgJyiDF4_2),.clk(gclk));
	jdff dff_B_rH54O8kr0_1(.din(n1685),.dout(w_dff_B_rH54O8kr0_1),.clk(gclk));
	jdff dff_B_k66MwJLp8_2(.din(n1633),.dout(w_dff_B_k66MwJLp8_2),.clk(gclk));
	jdff dff_B_bkeVVpIO9_2(.din(w_dff_B_k66MwJLp8_2),.dout(w_dff_B_bkeVVpIO9_2),.clk(gclk));
	jdff dff_B_4pebG2L49_2(.din(w_dff_B_bkeVVpIO9_2),.dout(w_dff_B_4pebG2L49_2),.clk(gclk));
	jdff dff_B_J1VdQMTL7_2(.din(w_dff_B_4pebG2L49_2),.dout(w_dff_B_J1VdQMTL7_2),.clk(gclk));
	jdff dff_B_fb4IbUOw3_2(.din(w_dff_B_J1VdQMTL7_2),.dout(w_dff_B_fb4IbUOw3_2),.clk(gclk));
	jdff dff_B_FrA7bjqF2_2(.din(w_dff_B_fb4IbUOw3_2),.dout(w_dff_B_FrA7bjqF2_2),.clk(gclk));
	jdff dff_B_CovZDhnp4_2(.din(w_dff_B_FrA7bjqF2_2),.dout(w_dff_B_CovZDhnp4_2),.clk(gclk));
	jdff dff_B_lrlDqXVL1_2(.din(w_dff_B_CovZDhnp4_2),.dout(w_dff_B_lrlDqXVL1_2),.clk(gclk));
	jdff dff_B_psq5de8v6_2(.din(w_dff_B_lrlDqXVL1_2),.dout(w_dff_B_psq5de8v6_2),.clk(gclk));
	jdff dff_B_Vz4VUZNa6_2(.din(w_dff_B_psq5de8v6_2),.dout(w_dff_B_Vz4VUZNa6_2),.clk(gclk));
	jdff dff_B_zZi9vpUJ3_2(.din(w_dff_B_Vz4VUZNa6_2),.dout(w_dff_B_zZi9vpUJ3_2),.clk(gclk));
	jdff dff_B_bei4QNnw6_2(.din(w_dff_B_zZi9vpUJ3_2),.dout(w_dff_B_bei4QNnw6_2),.clk(gclk));
	jdff dff_B_9PYZaKk22_2(.din(w_dff_B_bei4QNnw6_2),.dout(w_dff_B_9PYZaKk22_2),.clk(gclk));
	jdff dff_B_MACv1VX81_2(.din(w_dff_B_9PYZaKk22_2),.dout(w_dff_B_MACv1VX81_2),.clk(gclk));
	jdff dff_B_bmuiqEK48_2(.din(w_dff_B_MACv1VX81_2),.dout(w_dff_B_bmuiqEK48_2),.clk(gclk));
	jdff dff_B_RXpBW1OE1_2(.din(w_dff_B_bmuiqEK48_2),.dout(w_dff_B_RXpBW1OE1_2),.clk(gclk));
	jdff dff_B_cMAqL4IR1_2(.din(w_dff_B_RXpBW1OE1_2),.dout(w_dff_B_cMAqL4IR1_2),.clk(gclk));
	jdff dff_B_UdPbB9rR5_2(.din(w_dff_B_cMAqL4IR1_2),.dout(w_dff_B_UdPbB9rR5_2),.clk(gclk));
	jdff dff_B_z6YKWQYh4_2(.din(w_dff_B_UdPbB9rR5_2),.dout(w_dff_B_z6YKWQYh4_2),.clk(gclk));
	jdff dff_B_B59K5Qmb4_2(.din(w_dff_B_z6YKWQYh4_2),.dout(w_dff_B_B59K5Qmb4_2),.clk(gclk));
	jdff dff_B_zl22vhKO1_2(.din(w_dff_B_B59K5Qmb4_2),.dout(w_dff_B_zl22vhKO1_2),.clk(gclk));
	jdff dff_B_MD0eqtep3_2(.din(w_dff_B_zl22vhKO1_2),.dout(w_dff_B_MD0eqtep3_2),.clk(gclk));
	jdff dff_B_wtVkrcJt5_2(.din(w_dff_B_MD0eqtep3_2),.dout(w_dff_B_wtVkrcJt5_2),.clk(gclk));
	jdff dff_B_K42KxeUG1_2(.din(w_dff_B_wtVkrcJt5_2),.dout(w_dff_B_K42KxeUG1_2),.clk(gclk));
	jdff dff_B_9UR64zlS8_2(.din(w_dff_B_K42KxeUG1_2),.dout(w_dff_B_9UR64zlS8_2),.clk(gclk));
	jdff dff_B_pAWjWLdN1_2(.din(w_dff_B_9UR64zlS8_2),.dout(w_dff_B_pAWjWLdN1_2),.clk(gclk));
	jdff dff_B_MRoQTFT48_2(.din(w_dff_B_pAWjWLdN1_2),.dout(w_dff_B_MRoQTFT48_2),.clk(gclk));
	jdff dff_B_mMoH7CHO8_2(.din(w_dff_B_MRoQTFT48_2),.dout(w_dff_B_mMoH7CHO8_2),.clk(gclk));
	jdff dff_B_xaz2qoEw2_2(.din(w_dff_B_mMoH7CHO8_2),.dout(w_dff_B_xaz2qoEw2_2),.clk(gclk));
	jdff dff_B_BwYFzB2s0_2(.din(w_dff_B_xaz2qoEw2_2),.dout(w_dff_B_BwYFzB2s0_2),.clk(gclk));
	jdff dff_B_1RZ1TZC06_2(.din(w_dff_B_BwYFzB2s0_2),.dout(w_dff_B_1RZ1TZC06_2),.clk(gclk));
	jdff dff_B_8vJGM7z75_2(.din(w_dff_B_1RZ1TZC06_2),.dout(w_dff_B_8vJGM7z75_2),.clk(gclk));
	jdff dff_B_t9uBPWse6_2(.din(w_dff_B_8vJGM7z75_2),.dout(w_dff_B_t9uBPWse6_2),.clk(gclk));
	jdff dff_B_Zoo3vDB21_2(.din(w_dff_B_t9uBPWse6_2),.dout(w_dff_B_Zoo3vDB21_2),.clk(gclk));
	jdff dff_B_Nge3wDfC4_2(.din(w_dff_B_Zoo3vDB21_2),.dout(w_dff_B_Nge3wDfC4_2),.clk(gclk));
	jdff dff_B_16v6yqL68_2(.din(w_dff_B_Nge3wDfC4_2),.dout(w_dff_B_16v6yqL68_2),.clk(gclk));
	jdff dff_B_qo7QaHEe8_2(.din(w_dff_B_16v6yqL68_2),.dout(w_dff_B_qo7QaHEe8_2),.clk(gclk));
	jdff dff_B_mJYvVkCf4_2(.din(w_dff_B_qo7QaHEe8_2),.dout(w_dff_B_mJYvVkCf4_2),.clk(gclk));
	jdff dff_B_0h7UaMMb7_2(.din(w_dff_B_mJYvVkCf4_2),.dout(w_dff_B_0h7UaMMb7_2),.clk(gclk));
	jdff dff_B_IAqsdOpI8_2(.din(w_dff_B_0h7UaMMb7_2),.dout(w_dff_B_IAqsdOpI8_2),.clk(gclk));
	jdff dff_B_CUFAMhhL3_2(.din(w_dff_B_IAqsdOpI8_2),.dout(w_dff_B_CUFAMhhL3_2),.clk(gclk));
	jdff dff_B_rxe1wSSc2_2(.din(w_dff_B_CUFAMhhL3_2),.dout(w_dff_B_rxe1wSSc2_2),.clk(gclk));
	jdff dff_B_YdhuBDJN6_2(.din(w_dff_B_rxe1wSSc2_2),.dout(w_dff_B_YdhuBDJN6_2),.clk(gclk));
	jdff dff_B_gLWcJpwC8_2(.din(w_dff_B_YdhuBDJN6_2),.dout(w_dff_B_gLWcJpwC8_2),.clk(gclk));
	jdff dff_B_vDxlcce85_2(.din(w_dff_B_gLWcJpwC8_2),.dout(w_dff_B_vDxlcce85_2),.clk(gclk));
	jdff dff_B_uIBjKJe90_2(.din(n1636),.dout(w_dff_B_uIBjKJe90_2),.clk(gclk));
	jdff dff_B_UDKKrrrV9_1(.din(n1634),.dout(w_dff_B_UDKKrrrV9_1),.clk(gclk));
	jdff dff_B_bO1HDDwj3_2(.din(n1576),.dout(w_dff_B_bO1HDDwj3_2),.clk(gclk));
	jdff dff_B_chIXy3lL2_2(.din(w_dff_B_bO1HDDwj3_2),.dout(w_dff_B_chIXy3lL2_2),.clk(gclk));
	jdff dff_B_r3Gu3hpD8_2(.din(w_dff_B_chIXy3lL2_2),.dout(w_dff_B_r3Gu3hpD8_2),.clk(gclk));
	jdff dff_B_qpJxfoZs3_2(.din(w_dff_B_r3Gu3hpD8_2),.dout(w_dff_B_qpJxfoZs3_2),.clk(gclk));
	jdff dff_B_NKy6GcsM3_2(.din(w_dff_B_qpJxfoZs3_2),.dout(w_dff_B_NKy6GcsM3_2),.clk(gclk));
	jdff dff_B_BxgWGTsK4_2(.din(w_dff_B_NKy6GcsM3_2),.dout(w_dff_B_BxgWGTsK4_2),.clk(gclk));
	jdff dff_B_BDbAN8D03_2(.din(w_dff_B_BxgWGTsK4_2),.dout(w_dff_B_BDbAN8D03_2),.clk(gclk));
	jdff dff_B_WyaPA5Ay1_2(.din(w_dff_B_BDbAN8D03_2),.dout(w_dff_B_WyaPA5Ay1_2),.clk(gclk));
	jdff dff_B_rumB24580_2(.din(w_dff_B_WyaPA5Ay1_2),.dout(w_dff_B_rumB24580_2),.clk(gclk));
	jdff dff_B_IoaFiZMh7_2(.din(w_dff_B_rumB24580_2),.dout(w_dff_B_IoaFiZMh7_2),.clk(gclk));
	jdff dff_B_3reBQm4S5_2(.din(w_dff_B_IoaFiZMh7_2),.dout(w_dff_B_3reBQm4S5_2),.clk(gclk));
	jdff dff_B_hKVPuUGl2_2(.din(w_dff_B_3reBQm4S5_2),.dout(w_dff_B_hKVPuUGl2_2),.clk(gclk));
	jdff dff_B_w2onzORz0_2(.din(w_dff_B_hKVPuUGl2_2),.dout(w_dff_B_w2onzORz0_2),.clk(gclk));
	jdff dff_B_Wu3zD1GT5_2(.din(w_dff_B_w2onzORz0_2),.dout(w_dff_B_Wu3zD1GT5_2),.clk(gclk));
	jdff dff_B_3oRQ7EPQ5_2(.din(w_dff_B_Wu3zD1GT5_2),.dout(w_dff_B_3oRQ7EPQ5_2),.clk(gclk));
	jdff dff_B_V2T2MCnd2_2(.din(w_dff_B_3oRQ7EPQ5_2),.dout(w_dff_B_V2T2MCnd2_2),.clk(gclk));
	jdff dff_B_D62z7zpH8_2(.din(w_dff_B_V2T2MCnd2_2),.dout(w_dff_B_D62z7zpH8_2),.clk(gclk));
	jdff dff_B_xO1lNm0a8_2(.din(w_dff_B_D62z7zpH8_2),.dout(w_dff_B_xO1lNm0a8_2),.clk(gclk));
	jdff dff_B_RcoLN56Y8_2(.din(w_dff_B_xO1lNm0a8_2),.dout(w_dff_B_RcoLN56Y8_2),.clk(gclk));
	jdff dff_B_9Sfyq3fq3_2(.din(w_dff_B_RcoLN56Y8_2),.dout(w_dff_B_9Sfyq3fq3_2),.clk(gclk));
	jdff dff_B_GCtRIySl5_2(.din(w_dff_B_9Sfyq3fq3_2),.dout(w_dff_B_GCtRIySl5_2),.clk(gclk));
	jdff dff_B_Rxzq6Hj58_2(.din(w_dff_B_GCtRIySl5_2),.dout(w_dff_B_Rxzq6Hj58_2),.clk(gclk));
	jdff dff_B_MVwDUCoH2_2(.din(w_dff_B_Rxzq6Hj58_2),.dout(w_dff_B_MVwDUCoH2_2),.clk(gclk));
	jdff dff_B_U4ZsiqT29_2(.din(w_dff_B_MVwDUCoH2_2),.dout(w_dff_B_U4ZsiqT29_2),.clk(gclk));
	jdff dff_B_21KJvFnr3_2(.din(w_dff_B_U4ZsiqT29_2),.dout(w_dff_B_21KJvFnr3_2),.clk(gclk));
	jdff dff_B_HWFBSknv5_2(.din(w_dff_B_21KJvFnr3_2),.dout(w_dff_B_HWFBSknv5_2),.clk(gclk));
	jdff dff_B_f0A0QqQH0_2(.din(w_dff_B_HWFBSknv5_2),.dout(w_dff_B_f0A0QqQH0_2),.clk(gclk));
	jdff dff_B_vjyf2qyx1_2(.din(w_dff_B_f0A0QqQH0_2),.dout(w_dff_B_vjyf2qyx1_2),.clk(gclk));
	jdff dff_B_QlaCx6Ry9_2(.din(w_dff_B_vjyf2qyx1_2),.dout(w_dff_B_QlaCx6Ry9_2),.clk(gclk));
	jdff dff_B_UH0OclH40_2(.din(w_dff_B_QlaCx6Ry9_2),.dout(w_dff_B_UH0OclH40_2),.clk(gclk));
	jdff dff_B_Q67uGzm68_2(.din(w_dff_B_UH0OclH40_2),.dout(w_dff_B_Q67uGzm68_2),.clk(gclk));
	jdff dff_B_EaeVlffx3_2(.din(w_dff_B_Q67uGzm68_2),.dout(w_dff_B_EaeVlffx3_2),.clk(gclk));
	jdff dff_B_Onr2JCiq4_2(.din(w_dff_B_EaeVlffx3_2),.dout(w_dff_B_Onr2JCiq4_2),.clk(gclk));
	jdff dff_B_waqcrjzC2_2(.din(w_dff_B_Onr2JCiq4_2),.dout(w_dff_B_waqcrjzC2_2),.clk(gclk));
	jdff dff_B_jPtQqvO00_2(.din(w_dff_B_waqcrjzC2_2),.dout(w_dff_B_jPtQqvO00_2),.clk(gclk));
	jdff dff_B_noyzE1Lq2_2(.din(w_dff_B_jPtQqvO00_2),.dout(w_dff_B_noyzE1Lq2_2),.clk(gclk));
	jdff dff_B_atTiopd40_2(.din(w_dff_B_noyzE1Lq2_2),.dout(w_dff_B_atTiopd40_2),.clk(gclk));
	jdff dff_B_czSDJJiW8_2(.din(w_dff_B_atTiopd40_2),.dout(w_dff_B_czSDJJiW8_2),.clk(gclk));
	jdff dff_B_bAjjmrUk2_2(.din(w_dff_B_czSDJJiW8_2),.dout(w_dff_B_bAjjmrUk2_2),.clk(gclk));
	jdff dff_B_HzXNkwGQ5_2(.din(w_dff_B_bAjjmrUk2_2),.dout(w_dff_B_HzXNkwGQ5_2),.clk(gclk));
	jdff dff_B_ZP7WsaNU0_2(.din(w_dff_B_HzXNkwGQ5_2),.dout(w_dff_B_ZP7WsaNU0_2),.clk(gclk));
	jdff dff_B_diTzV2yZ9_2(.din(n1579),.dout(w_dff_B_diTzV2yZ9_2),.clk(gclk));
	jdff dff_B_WXGUjXj40_1(.din(n1577),.dout(w_dff_B_WXGUjXj40_1),.clk(gclk));
	jdff dff_B_5ppg6Ajf3_2(.din(n1512),.dout(w_dff_B_5ppg6Ajf3_2),.clk(gclk));
	jdff dff_B_W7yAxnHD6_2(.din(w_dff_B_5ppg6Ajf3_2),.dout(w_dff_B_W7yAxnHD6_2),.clk(gclk));
	jdff dff_B_5NqwLzV36_2(.din(w_dff_B_W7yAxnHD6_2),.dout(w_dff_B_5NqwLzV36_2),.clk(gclk));
	jdff dff_B_CeGX5VUo4_2(.din(w_dff_B_5NqwLzV36_2),.dout(w_dff_B_CeGX5VUo4_2),.clk(gclk));
	jdff dff_B_GHlkrBiz1_2(.din(w_dff_B_CeGX5VUo4_2),.dout(w_dff_B_GHlkrBiz1_2),.clk(gclk));
	jdff dff_B_OR7FTlHf7_2(.din(w_dff_B_GHlkrBiz1_2),.dout(w_dff_B_OR7FTlHf7_2),.clk(gclk));
	jdff dff_B_kSwtPMCL1_2(.din(w_dff_B_OR7FTlHf7_2),.dout(w_dff_B_kSwtPMCL1_2),.clk(gclk));
	jdff dff_B_mlEsU0SL2_2(.din(w_dff_B_kSwtPMCL1_2),.dout(w_dff_B_mlEsU0SL2_2),.clk(gclk));
	jdff dff_B_RwDcWrAK2_2(.din(w_dff_B_mlEsU0SL2_2),.dout(w_dff_B_RwDcWrAK2_2),.clk(gclk));
	jdff dff_B_h1NsZ8C62_2(.din(w_dff_B_RwDcWrAK2_2),.dout(w_dff_B_h1NsZ8C62_2),.clk(gclk));
	jdff dff_B_stCasSyO9_2(.din(w_dff_B_h1NsZ8C62_2),.dout(w_dff_B_stCasSyO9_2),.clk(gclk));
	jdff dff_B_KvRttgXt2_2(.din(w_dff_B_stCasSyO9_2),.dout(w_dff_B_KvRttgXt2_2),.clk(gclk));
	jdff dff_B_FfBVZBr27_2(.din(w_dff_B_KvRttgXt2_2),.dout(w_dff_B_FfBVZBr27_2),.clk(gclk));
	jdff dff_B_0soXRjRa4_2(.din(w_dff_B_FfBVZBr27_2),.dout(w_dff_B_0soXRjRa4_2),.clk(gclk));
	jdff dff_B_z4tShkuq0_2(.din(w_dff_B_0soXRjRa4_2),.dout(w_dff_B_z4tShkuq0_2),.clk(gclk));
	jdff dff_B_Wmm1juw91_2(.din(w_dff_B_z4tShkuq0_2),.dout(w_dff_B_Wmm1juw91_2),.clk(gclk));
	jdff dff_B_4Uowic3k0_2(.din(w_dff_B_Wmm1juw91_2),.dout(w_dff_B_4Uowic3k0_2),.clk(gclk));
	jdff dff_B_S1lm61At7_2(.din(w_dff_B_4Uowic3k0_2),.dout(w_dff_B_S1lm61At7_2),.clk(gclk));
	jdff dff_B_pChfuww06_2(.din(w_dff_B_S1lm61At7_2),.dout(w_dff_B_pChfuww06_2),.clk(gclk));
	jdff dff_B_qgAKR1ne5_2(.din(w_dff_B_pChfuww06_2),.dout(w_dff_B_qgAKR1ne5_2),.clk(gclk));
	jdff dff_B_SYWtNSKa2_2(.din(w_dff_B_qgAKR1ne5_2),.dout(w_dff_B_SYWtNSKa2_2),.clk(gclk));
	jdff dff_B_xd8kkPwt5_2(.din(w_dff_B_SYWtNSKa2_2),.dout(w_dff_B_xd8kkPwt5_2),.clk(gclk));
	jdff dff_B_LQgl3NRM4_2(.din(w_dff_B_xd8kkPwt5_2),.dout(w_dff_B_LQgl3NRM4_2),.clk(gclk));
	jdff dff_B_oyWHq5wA9_2(.din(w_dff_B_LQgl3NRM4_2),.dout(w_dff_B_oyWHq5wA9_2),.clk(gclk));
	jdff dff_B_bnUwPA7f9_2(.din(w_dff_B_oyWHq5wA9_2),.dout(w_dff_B_bnUwPA7f9_2),.clk(gclk));
	jdff dff_B_2sJRKZjp7_2(.din(w_dff_B_bnUwPA7f9_2),.dout(w_dff_B_2sJRKZjp7_2),.clk(gclk));
	jdff dff_B_grEGwFDf6_2(.din(w_dff_B_2sJRKZjp7_2),.dout(w_dff_B_grEGwFDf6_2),.clk(gclk));
	jdff dff_B_L9PRyrWY3_2(.din(w_dff_B_grEGwFDf6_2),.dout(w_dff_B_L9PRyrWY3_2),.clk(gclk));
	jdff dff_B_M7FDF4N17_2(.din(w_dff_B_L9PRyrWY3_2),.dout(w_dff_B_M7FDF4N17_2),.clk(gclk));
	jdff dff_B_VI1Dtueh6_2(.din(w_dff_B_M7FDF4N17_2),.dout(w_dff_B_VI1Dtueh6_2),.clk(gclk));
	jdff dff_B_Gnz4gFRi6_2(.din(w_dff_B_VI1Dtueh6_2),.dout(w_dff_B_Gnz4gFRi6_2),.clk(gclk));
	jdff dff_B_seSrTjLh5_2(.din(w_dff_B_Gnz4gFRi6_2),.dout(w_dff_B_seSrTjLh5_2),.clk(gclk));
	jdff dff_B_aYfvuTza0_2(.din(w_dff_B_seSrTjLh5_2),.dout(w_dff_B_aYfvuTza0_2),.clk(gclk));
	jdff dff_B_LIo79Tfs1_2(.din(w_dff_B_aYfvuTza0_2),.dout(w_dff_B_LIo79Tfs1_2),.clk(gclk));
	jdff dff_B_zHXtUCGX5_2(.din(w_dff_B_LIo79Tfs1_2),.dout(w_dff_B_zHXtUCGX5_2),.clk(gclk));
	jdff dff_B_Luf9Nf274_2(.din(w_dff_B_zHXtUCGX5_2),.dout(w_dff_B_Luf9Nf274_2),.clk(gclk));
	jdff dff_B_vWEqRT4V1_2(.din(w_dff_B_Luf9Nf274_2),.dout(w_dff_B_vWEqRT4V1_2),.clk(gclk));
	jdff dff_B_IcO8rX5a7_2(.din(n1515),.dout(w_dff_B_IcO8rX5a7_2),.clk(gclk));
	jdff dff_B_dEwrKoGB5_1(.din(n1513),.dout(w_dff_B_dEwrKoGB5_1),.clk(gclk));
	jdff dff_B_j5H20azp7_2(.din(n1441),.dout(w_dff_B_j5H20azp7_2),.clk(gclk));
	jdff dff_B_F5wZsKrk6_2(.din(w_dff_B_j5H20azp7_2),.dout(w_dff_B_F5wZsKrk6_2),.clk(gclk));
	jdff dff_B_nw90zict1_2(.din(w_dff_B_F5wZsKrk6_2),.dout(w_dff_B_nw90zict1_2),.clk(gclk));
	jdff dff_B_7vDRSFeR0_2(.din(w_dff_B_nw90zict1_2),.dout(w_dff_B_7vDRSFeR0_2),.clk(gclk));
	jdff dff_B_wHzxIEBr5_2(.din(w_dff_B_7vDRSFeR0_2),.dout(w_dff_B_wHzxIEBr5_2),.clk(gclk));
	jdff dff_B_Mc71VNGq4_2(.din(w_dff_B_wHzxIEBr5_2),.dout(w_dff_B_Mc71VNGq4_2),.clk(gclk));
	jdff dff_B_oNbjh2yC5_2(.din(w_dff_B_Mc71VNGq4_2),.dout(w_dff_B_oNbjh2yC5_2),.clk(gclk));
	jdff dff_B_nGTDOzjN8_2(.din(w_dff_B_oNbjh2yC5_2),.dout(w_dff_B_nGTDOzjN8_2),.clk(gclk));
	jdff dff_B_taxqBUud3_2(.din(w_dff_B_nGTDOzjN8_2),.dout(w_dff_B_taxqBUud3_2),.clk(gclk));
	jdff dff_B_9yUfE9mN0_2(.din(w_dff_B_taxqBUud3_2),.dout(w_dff_B_9yUfE9mN0_2),.clk(gclk));
	jdff dff_B_elH7HKcZ1_2(.din(w_dff_B_9yUfE9mN0_2),.dout(w_dff_B_elH7HKcZ1_2),.clk(gclk));
	jdff dff_B_QeYhkzT07_2(.din(w_dff_B_elH7HKcZ1_2),.dout(w_dff_B_QeYhkzT07_2),.clk(gclk));
	jdff dff_B_XnRU8dS32_2(.din(w_dff_B_QeYhkzT07_2),.dout(w_dff_B_XnRU8dS32_2),.clk(gclk));
	jdff dff_B_kuokYYNo3_2(.din(w_dff_B_XnRU8dS32_2),.dout(w_dff_B_kuokYYNo3_2),.clk(gclk));
	jdff dff_B_YDfAOY1p7_2(.din(w_dff_B_kuokYYNo3_2),.dout(w_dff_B_YDfAOY1p7_2),.clk(gclk));
	jdff dff_B_veox868p9_2(.din(w_dff_B_YDfAOY1p7_2),.dout(w_dff_B_veox868p9_2),.clk(gclk));
	jdff dff_B_nvOSqB0B4_2(.din(w_dff_B_veox868p9_2),.dout(w_dff_B_nvOSqB0B4_2),.clk(gclk));
	jdff dff_B_7uh7XS7l9_2(.din(w_dff_B_nvOSqB0B4_2),.dout(w_dff_B_7uh7XS7l9_2),.clk(gclk));
	jdff dff_B_4BSMdsXu5_2(.din(w_dff_B_7uh7XS7l9_2),.dout(w_dff_B_4BSMdsXu5_2),.clk(gclk));
	jdff dff_B_LEs3JQ704_2(.din(w_dff_B_4BSMdsXu5_2),.dout(w_dff_B_LEs3JQ704_2),.clk(gclk));
	jdff dff_B_pnvOZK6z4_2(.din(w_dff_B_LEs3JQ704_2),.dout(w_dff_B_pnvOZK6z4_2),.clk(gclk));
	jdff dff_B_0ajzQRWW9_2(.din(w_dff_B_pnvOZK6z4_2),.dout(w_dff_B_0ajzQRWW9_2),.clk(gclk));
	jdff dff_B_6IVayNTO5_2(.din(w_dff_B_0ajzQRWW9_2),.dout(w_dff_B_6IVayNTO5_2),.clk(gclk));
	jdff dff_B_j4aMwnCJ3_2(.din(w_dff_B_6IVayNTO5_2),.dout(w_dff_B_j4aMwnCJ3_2),.clk(gclk));
	jdff dff_B_IrdULxle6_2(.din(w_dff_B_j4aMwnCJ3_2),.dout(w_dff_B_IrdULxle6_2),.clk(gclk));
	jdff dff_B_PlYmr6iJ2_2(.din(w_dff_B_IrdULxle6_2),.dout(w_dff_B_PlYmr6iJ2_2),.clk(gclk));
	jdff dff_B_h2itkcX45_2(.din(w_dff_B_PlYmr6iJ2_2),.dout(w_dff_B_h2itkcX45_2),.clk(gclk));
	jdff dff_B_kleeMFqW0_2(.din(w_dff_B_h2itkcX45_2),.dout(w_dff_B_kleeMFqW0_2),.clk(gclk));
	jdff dff_B_wcWwAPLW3_2(.din(w_dff_B_kleeMFqW0_2),.dout(w_dff_B_wcWwAPLW3_2),.clk(gclk));
	jdff dff_B_2AjHcWcm6_2(.din(w_dff_B_wcWwAPLW3_2),.dout(w_dff_B_2AjHcWcm6_2),.clk(gclk));
	jdff dff_B_9dZpEyNN0_2(.din(w_dff_B_2AjHcWcm6_2),.dout(w_dff_B_9dZpEyNN0_2),.clk(gclk));
	jdff dff_B_MiSq2gaE4_2(.din(w_dff_B_9dZpEyNN0_2),.dout(w_dff_B_MiSq2gaE4_2),.clk(gclk));
	jdff dff_B_Lm7RFGGj8_2(.din(w_dff_B_MiSq2gaE4_2),.dout(w_dff_B_Lm7RFGGj8_2),.clk(gclk));
	jdff dff_B_6TwkF4Yo1_1(.din(n1442),.dout(w_dff_B_6TwkF4Yo1_1),.clk(gclk));
	jdff dff_B_svmI7hRn1_2(.din(n1363),.dout(w_dff_B_svmI7hRn1_2),.clk(gclk));
	jdff dff_B_RlCsqdxM7_2(.din(w_dff_B_svmI7hRn1_2),.dout(w_dff_B_RlCsqdxM7_2),.clk(gclk));
	jdff dff_B_O6OPwk9x2_2(.din(w_dff_B_RlCsqdxM7_2),.dout(w_dff_B_O6OPwk9x2_2),.clk(gclk));
	jdff dff_B_ebBitJCz4_2(.din(w_dff_B_O6OPwk9x2_2),.dout(w_dff_B_ebBitJCz4_2),.clk(gclk));
	jdff dff_B_WmmHSPAr8_2(.din(w_dff_B_ebBitJCz4_2),.dout(w_dff_B_WmmHSPAr8_2),.clk(gclk));
	jdff dff_B_TIBZ03Xc2_2(.din(w_dff_B_WmmHSPAr8_2),.dout(w_dff_B_TIBZ03Xc2_2),.clk(gclk));
	jdff dff_B_zG5oYa8T0_2(.din(w_dff_B_TIBZ03Xc2_2),.dout(w_dff_B_zG5oYa8T0_2),.clk(gclk));
	jdff dff_B_N3keFv7v3_2(.din(w_dff_B_zG5oYa8T0_2),.dout(w_dff_B_N3keFv7v3_2),.clk(gclk));
	jdff dff_B_nzvJ5CoE7_2(.din(w_dff_B_N3keFv7v3_2),.dout(w_dff_B_nzvJ5CoE7_2),.clk(gclk));
	jdff dff_B_uBSzNkwD9_2(.din(w_dff_B_nzvJ5CoE7_2),.dout(w_dff_B_uBSzNkwD9_2),.clk(gclk));
	jdff dff_B_FFkodaBl1_2(.din(w_dff_B_uBSzNkwD9_2),.dout(w_dff_B_FFkodaBl1_2),.clk(gclk));
	jdff dff_B_MtD9L4fq2_2(.din(w_dff_B_FFkodaBl1_2),.dout(w_dff_B_MtD9L4fq2_2),.clk(gclk));
	jdff dff_B_wtNZsY9p5_2(.din(w_dff_B_MtD9L4fq2_2),.dout(w_dff_B_wtNZsY9p5_2),.clk(gclk));
	jdff dff_B_H4qA5dOq5_2(.din(w_dff_B_wtNZsY9p5_2),.dout(w_dff_B_H4qA5dOq5_2),.clk(gclk));
	jdff dff_B_imVBRHtE0_2(.din(w_dff_B_H4qA5dOq5_2),.dout(w_dff_B_imVBRHtE0_2),.clk(gclk));
	jdff dff_B_20nZ7xzd7_2(.din(w_dff_B_imVBRHtE0_2),.dout(w_dff_B_20nZ7xzd7_2),.clk(gclk));
	jdff dff_B_pIx08jGb9_2(.din(w_dff_B_20nZ7xzd7_2),.dout(w_dff_B_pIx08jGb9_2),.clk(gclk));
	jdff dff_B_SIWUZzmW4_2(.din(w_dff_B_pIx08jGb9_2),.dout(w_dff_B_SIWUZzmW4_2),.clk(gclk));
	jdff dff_B_Ub0zW7589_2(.din(w_dff_B_SIWUZzmW4_2),.dout(w_dff_B_Ub0zW7589_2),.clk(gclk));
	jdff dff_B_QXuqqmhL8_2(.din(w_dff_B_Ub0zW7589_2),.dout(w_dff_B_QXuqqmhL8_2),.clk(gclk));
	jdff dff_B_jzJVLdmV8_2(.din(w_dff_B_QXuqqmhL8_2),.dout(w_dff_B_jzJVLdmV8_2),.clk(gclk));
	jdff dff_B_2A2K6pco0_2(.din(w_dff_B_jzJVLdmV8_2),.dout(w_dff_B_2A2K6pco0_2),.clk(gclk));
	jdff dff_B_Q6e4xXjn6_2(.din(w_dff_B_2A2K6pco0_2),.dout(w_dff_B_Q6e4xXjn6_2),.clk(gclk));
	jdff dff_B_pJ6jJO6X4_2(.din(w_dff_B_Q6e4xXjn6_2),.dout(w_dff_B_pJ6jJO6X4_2),.clk(gclk));
	jdff dff_B_Giaq3oEH5_2(.din(w_dff_B_pJ6jJO6X4_2),.dout(w_dff_B_Giaq3oEH5_2),.clk(gclk));
	jdff dff_B_F1pyfHCD8_2(.din(w_dff_B_Giaq3oEH5_2),.dout(w_dff_B_F1pyfHCD8_2),.clk(gclk));
	jdff dff_B_LFCXrPL63_2(.din(w_dff_B_F1pyfHCD8_2),.dout(w_dff_B_LFCXrPL63_2),.clk(gclk));
	jdff dff_B_OG3yEUGn6_2(.din(w_dff_B_LFCXrPL63_2),.dout(w_dff_B_OG3yEUGn6_2),.clk(gclk));
	jdff dff_B_DeO4FRWO6_2(.din(w_dff_B_OG3yEUGn6_2),.dout(w_dff_B_DeO4FRWO6_2),.clk(gclk));
	jdff dff_B_vCLHSOEX6_2(.din(w_dff_B_DeO4FRWO6_2),.dout(w_dff_B_vCLHSOEX6_2),.clk(gclk));
	jdff dff_B_sSCut7rS2_2(.din(n1395),.dout(w_dff_B_sSCut7rS2_2),.clk(gclk));
	jdff dff_B_bemMx2d96_1(.din(n1364),.dout(w_dff_B_bemMx2d96_1),.clk(gclk));
	jdff dff_B_4AC5pT9Q8_2(.din(n1278),.dout(w_dff_B_4AC5pT9Q8_2),.clk(gclk));
	jdff dff_B_28tN70Jt4_2(.din(w_dff_B_4AC5pT9Q8_2),.dout(w_dff_B_28tN70Jt4_2),.clk(gclk));
	jdff dff_B_XigzSZeI8_2(.din(w_dff_B_28tN70Jt4_2),.dout(w_dff_B_XigzSZeI8_2),.clk(gclk));
	jdff dff_B_7087JP5Z0_2(.din(w_dff_B_XigzSZeI8_2),.dout(w_dff_B_7087JP5Z0_2),.clk(gclk));
	jdff dff_B_FZvQ8w9q8_2(.din(w_dff_B_7087JP5Z0_2),.dout(w_dff_B_FZvQ8w9q8_2),.clk(gclk));
	jdff dff_B_ljSEm1H61_2(.din(w_dff_B_FZvQ8w9q8_2),.dout(w_dff_B_ljSEm1H61_2),.clk(gclk));
	jdff dff_B_YW2hYdpE4_2(.din(w_dff_B_ljSEm1H61_2),.dout(w_dff_B_YW2hYdpE4_2),.clk(gclk));
	jdff dff_B_kMFhGTuv6_2(.din(w_dff_B_YW2hYdpE4_2),.dout(w_dff_B_kMFhGTuv6_2),.clk(gclk));
	jdff dff_B_aA8uHYOJ9_2(.din(w_dff_B_kMFhGTuv6_2),.dout(w_dff_B_aA8uHYOJ9_2),.clk(gclk));
	jdff dff_B_a09USQzg9_2(.din(w_dff_B_aA8uHYOJ9_2),.dout(w_dff_B_a09USQzg9_2),.clk(gclk));
	jdff dff_B_HlBs94x52_2(.din(w_dff_B_a09USQzg9_2),.dout(w_dff_B_HlBs94x52_2),.clk(gclk));
	jdff dff_B_RjlK8Ewe4_2(.din(w_dff_B_HlBs94x52_2),.dout(w_dff_B_RjlK8Ewe4_2),.clk(gclk));
	jdff dff_B_0gwwOZZh3_2(.din(w_dff_B_RjlK8Ewe4_2),.dout(w_dff_B_0gwwOZZh3_2),.clk(gclk));
	jdff dff_B_5b65wC8t8_2(.din(w_dff_B_0gwwOZZh3_2),.dout(w_dff_B_5b65wC8t8_2),.clk(gclk));
	jdff dff_B_Aqt3R2jC1_2(.din(w_dff_B_5b65wC8t8_2),.dout(w_dff_B_Aqt3R2jC1_2),.clk(gclk));
	jdff dff_B_6rSPOryw7_2(.din(w_dff_B_Aqt3R2jC1_2),.dout(w_dff_B_6rSPOryw7_2),.clk(gclk));
	jdff dff_B_4sbSCeOV9_2(.din(w_dff_B_6rSPOryw7_2),.dout(w_dff_B_4sbSCeOV9_2),.clk(gclk));
	jdff dff_B_Ucw76F171_2(.din(w_dff_B_4sbSCeOV9_2),.dout(w_dff_B_Ucw76F171_2),.clk(gclk));
	jdff dff_B_vfiwW1cI5_2(.din(w_dff_B_Ucw76F171_2),.dout(w_dff_B_vfiwW1cI5_2),.clk(gclk));
	jdff dff_B_BaPgsUkv8_2(.din(w_dff_B_vfiwW1cI5_2),.dout(w_dff_B_BaPgsUkv8_2),.clk(gclk));
	jdff dff_B_C0w1Xh9z6_2(.din(w_dff_B_BaPgsUkv8_2),.dout(w_dff_B_C0w1Xh9z6_2),.clk(gclk));
	jdff dff_B_ySMyQfaL6_2(.din(w_dff_B_C0w1Xh9z6_2),.dout(w_dff_B_ySMyQfaL6_2),.clk(gclk));
	jdff dff_B_xger0zA40_2(.din(w_dff_B_ySMyQfaL6_2),.dout(w_dff_B_xger0zA40_2),.clk(gclk));
	jdff dff_B_2qLdy5R17_2(.din(w_dff_B_xger0zA40_2),.dout(w_dff_B_2qLdy5R17_2),.clk(gclk));
	jdff dff_B_7UwSXrye8_2(.din(w_dff_B_2qLdy5R17_2),.dout(w_dff_B_7UwSXrye8_2),.clk(gclk));
	jdff dff_B_7ol1otzE3_2(.din(w_dff_B_7UwSXrye8_2),.dout(w_dff_B_7ol1otzE3_2),.clk(gclk));
	jdff dff_B_MuvFa1BM3_2(.din(w_dff_B_7ol1otzE3_2),.dout(w_dff_B_MuvFa1BM3_2),.clk(gclk));
	jdff dff_B_KrtcCkho1_2(.din(n1310),.dout(w_dff_B_KrtcCkho1_2),.clk(gclk));
	jdff dff_B_Mhl3G5ff3_1(.din(n1279),.dout(w_dff_B_Mhl3G5ff3_1),.clk(gclk));
	jdff dff_B_JF4915eS3_2(.din(n1188),.dout(w_dff_B_JF4915eS3_2),.clk(gclk));
	jdff dff_B_jpfrmX392_2(.din(w_dff_B_JF4915eS3_2),.dout(w_dff_B_jpfrmX392_2),.clk(gclk));
	jdff dff_B_WGARxPBc3_2(.din(w_dff_B_jpfrmX392_2),.dout(w_dff_B_WGARxPBc3_2),.clk(gclk));
	jdff dff_B_z25QBqam0_2(.din(w_dff_B_WGARxPBc3_2),.dout(w_dff_B_z25QBqam0_2),.clk(gclk));
	jdff dff_B_o9T6pYs51_2(.din(w_dff_B_z25QBqam0_2),.dout(w_dff_B_o9T6pYs51_2),.clk(gclk));
	jdff dff_B_90HNUajS3_2(.din(w_dff_B_o9T6pYs51_2),.dout(w_dff_B_90HNUajS3_2),.clk(gclk));
	jdff dff_B_AzmHqcUH8_2(.din(w_dff_B_90HNUajS3_2),.dout(w_dff_B_AzmHqcUH8_2),.clk(gclk));
	jdff dff_B_RKOPdOCw7_2(.din(w_dff_B_AzmHqcUH8_2),.dout(w_dff_B_RKOPdOCw7_2),.clk(gclk));
	jdff dff_B_dQdVIRSe7_2(.din(w_dff_B_RKOPdOCw7_2),.dout(w_dff_B_dQdVIRSe7_2),.clk(gclk));
	jdff dff_B_EIJQmjBq7_2(.din(w_dff_B_dQdVIRSe7_2),.dout(w_dff_B_EIJQmjBq7_2),.clk(gclk));
	jdff dff_B_mHWjMcIl5_2(.din(w_dff_B_EIJQmjBq7_2),.dout(w_dff_B_mHWjMcIl5_2),.clk(gclk));
	jdff dff_B_3706xz309_2(.din(w_dff_B_mHWjMcIl5_2),.dout(w_dff_B_3706xz309_2),.clk(gclk));
	jdff dff_B_aXZB5NRb8_2(.din(w_dff_B_3706xz309_2),.dout(w_dff_B_aXZB5NRb8_2),.clk(gclk));
	jdff dff_B_9k1Sy2v61_2(.din(w_dff_B_aXZB5NRb8_2),.dout(w_dff_B_9k1Sy2v61_2),.clk(gclk));
	jdff dff_B_8OYUEyyz1_2(.din(w_dff_B_9k1Sy2v61_2),.dout(w_dff_B_8OYUEyyz1_2),.clk(gclk));
	jdff dff_B_jmNlidCd0_2(.din(w_dff_B_8OYUEyyz1_2),.dout(w_dff_B_jmNlidCd0_2),.clk(gclk));
	jdff dff_B_0SJ0gnuq1_2(.din(w_dff_B_jmNlidCd0_2),.dout(w_dff_B_0SJ0gnuq1_2),.clk(gclk));
	jdff dff_B_yFFtZVHl8_2(.din(w_dff_B_0SJ0gnuq1_2),.dout(w_dff_B_yFFtZVHl8_2),.clk(gclk));
	jdff dff_B_I4HaKqUQ0_2(.din(w_dff_B_yFFtZVHl8_2),.dout(w_dff_B_I4HaKqUQ0_2),.clk(gclk));
	jdff dff_B_zZLvfhrD0_2(.din(w_dff_B_I4HaKqUQ0_2),.dout(w_dff_B_zZLvfhrD0_2),.clk(gclk));
	jdff dff_B_NmKAB2KR4_2(.din(w_dff_B_zZLvfhrD0_2),.dout(w_dff_B_NmKAB2KR4_2),.clk(gclk));
	jdff dff_B_q5mlOs9c6_2(.din(w_dff_B_NmKAB2KR4_2),.dout(w_dff_B_q5mlOs9c6_2),.clk(gclk));
	jdff dff_B_IgJPhkhL0_2(.din(w_dff_B_q5mlOs9c6_2),.dout(w_dff_B_IgJPhkhL0_2),.clk(gclk));
	jdff dff_B_Qb35jaaX6_2(.din(w_dff_B_IgJPhkhL0_2),.dout(w_dff_B_Qb35jaaX6_2),.clk(gclk));
	jdff dff_B_26ORQgZm0_2(.din(n1219),.dout(w_dff_B_26ORQgZm0_2),.clk(gclk));
	jdff dff_B_y1QTgYa17_1(.din(n1189),.dout(w_dff_B_y1QTgYa17_1),.clk(gclk));
	jdff dff_B_3I0pdiAz6_2(.din(n1084),.dout(w_dff_B_3I0pdiAz6_2),.clk(gclk));
	jdff dff_B_Qwey936N3_2(.din(w_dff_B_3I0pdiAz6_2),.dout(w_dff_B_Qwey936N3_2),.clk(gclk));
	jdff dff_B_BGGLXxHc5_2(.din(w_dff_B_Qwey936N3_2),.dout(w_dff_B_BGGLXxHc5_2),.clk(gclk));
	jdff dff_B_pdzRoFHZ1_2(.din(w_dff_B_BGGLXxHc5_2),.dout(w_dff_B_pdzRoFHZ1_2),.clk(gclk));
	jdff dff_B_D8daikzJ5_2(.din(w_dff_B_pdzRoFHZ1_2),.dout(w_dff_B_D8daikzJ5_2),.clk(gclk));
	jdff dff_B_Wduch9Zu9_2(.din(w_dff_B_D8daikzJ5_2),.dout(w_dff_B_Wduch9Zu9_2),.clk(gclk));
	jdff dff_B_92e2RsYI5_2(.din(w_dff_B_Wduch9Zu9_2),.dout(w_dff_B_92e2RsYI5_2),.clk(gclk));
	jdff dff_B_9tTjV6HB5_2(.din(w_dff_B_92e2RsYI5_2),.dout(w_dff_B_9tTjV6HB5_2),.clk(gclk));
	jdff dff_B_PhXhOdmP9_2(.din(w_dff_B_9tTjV6HB5_2),.dout(w_dff_B_PhXhOdmP9_2),.clk(gclk));
	jdff dff_B_gFxfOnAp5_2(.din(w_dff_B_PhXhOdmP9_2),.dout(w_dff_B_gFxfOnAp5_2),.clk(gclk));
	jdff dff_B_6VfZPh0A2_2(.din(w_dff_B_gFxfOnAp5_2),.dout(w_dff_B_6VfZPh0A2_2),.clk(gclk));
	jdff dff_B_DfHUZZgs5_2(.din(w_dff_B_6VfZPh0A2_2),.dout(w_dff_B_DfHUZZgs5_2),.clk(gclk));
	jdff dff_B_fRkCD2Mu6_2(.din(w_dff_B_DfHUZZgs5_2),.dout(w_dff_B_fRkCD2Mu6_2),.clk(gclk));
	jdff dff_B_GGbfKkwR8_2(.din(w_dff_B_fRkCD2Mu6_2),.dout(w_dff_B_GGbfKkwR8_2),.clk(gclk));
	jdff dff_B_yf7b5EYl3_2(.din(w_dff_B_GGbfKkwR8_2),.dout(w_dff_B_yf7b5EYl3_2),.clk(gclk));
	jdff dff_B_jGHlGI6w4_2(.din(w_dff_B_yf7b5EYl3_2),.dout(w_dff_B_jGHlGI6w4_2),.clk(gclk));
	jdff dff_B_47WLpT4Z0_2(.din(w_dff_B_jGHlGI6w4_2),.dout(w_dff_B_47WLpT4Z0_2),.clk(gclk));
	jdff dff_B_c259OeZs9_2(.din(w_dff_B_47WLpT4Z0_2),.dout(w_dff_B_c259OeZs9_2),.clk(gclk));
	jdff dff_B_9gvvRstr6_2(.din(w_dff_B_c259OeZs9_2),.dout(w_dff_B_9gvvRstr6_2),.clk(gclk));
	jdff dff_B_ctAfkzK51_2(.din(w_dff_B_9gvvRstr6_2),.dout(w_dff_B_ctAfkzK51_2),.clk(gclk));
	jdff dff_B_E8f9MlnF1_2(.din(w_dff_B_ctAfkzK51_2),.dout(w_dff_B_E8f9MlnF1_2),.clk(gclk));
	jdff dff_B_zGdvxZ9X5_2(.din(n1121),.dout(w_dff_B_zGdvxZ9X5_2),.clk(gclk));
	jdff dff_B_ITjObB5K9_1(.din(n1085),.dout(w_dff_B_ITjObB5K9_1),.clk(gclk));
	jdff dff_B_N7TCNxmV2_2(.din(n986),.dout(w_dff_B_N7TCNxmV2_2),.clk(gclk));
	jdff dff_B_6RLHAqst4_2(.din(w_dff_B_N7TCNxmV2_2),.dout(w_dff_B_6RLHAqst4_2),.clk(gclk));
	jdff dff_B_weu18uus0_2(.din(w_dff_B_6RLHAqst4_2),.dout(w_dff_B_weu18uus0_2),.clk(gclk));
	jdff dff_B_dMckLTxl9_2(.din(w_dff_B_weu18uus0_2),.dout(w_dff_B_dMckLTxl9_2),.clk(gclk));
	jdff dff_B_YYehwJwc0_2(.din(w_dff_B_dMckLTxl9_2),.dout(w_dff_B_YYehwJwc0_2),.clk(gclk));
	jdff dff_B_GE8Zn5Oz5_2(.din(w_dff_B_YYehwJwc0_2),.dout(w_dff_B_GE8Zn5Oz5_2),.clk(gclk));
	jdff dff_B_BhW9enfR8_2(.din(w_dff_B_GE8Zn5Oz5_2),.dout(w_dff_B_BhW9enfR8_2),.clk(gclk));
	jdff dff_B_FtgXLwPf4_2(.din(w_dff_B_BhW9enfR8_2),.dout(w_dff_B_FtgXLwPf4_2),.clk(gclk));
	jdff dff_B_2HUK1EPC7_2(.din(w_dff_B_FtgXLwPf4_2),.dout(w_dff_B_2HUK1EPC7_2),.clk(gclk));
	jdff dff_B_LIsFbDa67_2(.din(w_dff_B_2HUK1EPC7_2),.dout(w_dff_B_LIsFbDa67_2),.clk(gclk));
	jdff dff_B_x61XG7fo3_2(.din(w_dff_B_LIsFbDa67_2),.dout(w_dff_B_x61XG7fo3_2),.clk(gclk));
	jdff dff_B_YdDsdxE02_2(.din(w_dff_B_x61XG7fo3_2),.dout(w_dff_B_YdDsdxE02_2),.clk(gclk));
	jdff dff_B_jY7xnavw9_2(.din(w_dff_B_YdDsdxE02_2),.dout(w_dff_B_jY7xnavw9_2),.clk(gclk));
	jdff dff_B_82ANAqHI4_2(.din(w_dff_B_jY7xnavw9_2),.dout(w_dff_B_82ANAqHI4_2),.clk(gclk));
	jdff dff_B_JLQenPXC9_2(.din(w_dff_B_82ANAqHI4_2),.dout(w_dff_B_JLQenPXC9_2),.clk(gclk));
	jdff dff_B_DaNXQWe25_2(.din(w_dff_B_JLQenPXC9_2),.dout(w_dff_B_DaNXQWe25_2),.clk(gclk));
	jdff dff_B_868EQ2Rv7_2(.din(w_dff_B_DaNXQWe25_2),.dout(w_dff_B_868EQ2Rv7_2),.clk(gclk));
	jdff dff_B_ZWgEyIQa3_2(.din(w_dff_B_868EQ2Rv7_2),.dout(w_dff_B_ZWgEyIQa3_2),.clk(gclk));
	jdff dff_B_CvCblr1X9_2(.din(n1016),.dout(w_dff_B_CvCblr1X9_2),.clk(gclk));
	jdff dff_B_UnQj650K1_1(.din(n987),.dout(w_dff_B_UnQj650K1_1),.clk(gclk));
	jdff dff_B_lSW0Sf5z8_2(.din(n881),.dout(w_dff_B_lSW0Sf5z8_2),.clk(gclk));
	jdff dff_B_As7dHRBf6_2(.din(w_dff_B_lSW0Sf5z8_2),.dout(w_dff_B_As7dHRBf6_2),.clk(gclk));
	jdff dff_B_y7zUfQeL0_2(.din(w_dff_B_As7dHRBf6_2),.dout(w_dff_B_y7zUfQeL0_2),.clk(gclk));
	jdff dff_B_q9xohqDe9_2(.din(w_dff_B_y7zUfQeL0_2),.dout(w_dff_B_q9xohqDe9_2),.clk(gclk));
	jdff dff_B_7Ck9HBFN0_2(.din(w_dff_B_q9xohqDe9_2),.dout(w_dff_B_7Ck9HBFN0_2),.clk(gclk));
	jdff dff_B_5uZJCWtN4_2(.din(w_dff_B_7Ck9HBFN0_2),.dout(w_dff_B_5uZJCWtN4_2),.clk(gclk));
	jdff dff_B_KK6Lbwbz1_2(.din(w_dff_B_5uZJCWtN4_2),.dout(w_dff_B_KK6Lbwbz1_2),.clk(gclk));
	jdff dff_B_76jY0EUF1_2(.din(w_dff_B_KK6Lbwbz1_2),.dout(w_dff_B_76jY0EUF1_2),.clk(gclk));
	jdff dff_B_kM1yDmwx5_2(.din(w_dff_B_76jY0EUF1_2),.dout(w_dff_B_kM1yDmwx5_2),.clk(gclk));
	jdff dff_B_nUDDhB3m6_2(.din(w_dff_B_kM1yDmwx5_2),.dout(w_dff_B_nUDDhB3m6_2),.clk(gclk));
	jdff dff_B_6C7m0p0u1_2(.din(w_dff_B_nUDDhB3m6_2),.dout(w_dff_B_6C7m0p0u1_2),.clk(gclk));
	jdff dff_B_FAL7FRdG4_2(.din(w_dff_B_6C7m0p0u1_2),.dout(w_dff_B_FAL7FRdG4_2),.clk(gclk));
	jdff dff_B_kOQqsB679_2(.din(w_dff_B_FAL7FRdG4_2),.dout(w_dff_B_kOQqsB679_2),.clk(gclk));
	jdff dff_B_AB5qckfb4_2(.din(w_dff_B_kOQqsB679_2),.dout(w_dff_B_AB5qckfb4_2),.clk(gclk));
	jdff dff_B_iSePcQlc6_2(.din(w_dff_B_AB5qckfb4_2),.dout(w_dff_B_iSePcQlc6_2),.clk(gclk));
	jdff dff_B_r3cc26Gc8_2(.din(n911),.dout(w_dff_B_r3cc26Gc8_2),.clk(gclk));
	jdff dff_B_A83BQhCB9_1(.din(n882),.dout(w_dff_B_A83BQhCB9_1),.clk(gclk));
	jdff dff_B_BTA1Y7983_2(.din(n782),.dout(w_dff_B_BTA1Y7983_2),.clk(gclk));
	jdff dff_B_dod5aWcE3_2(.din(w_dff_B_BTA1Y7983_2),.dout(w_dff_B_dod5aWcE3_2),.clk(gclk));
	jdff dff_B_TEBdbmRm8_2(.din(w_dff_B_dod5aWcE3_2),.dout(w_dff_B_TEBdbmRm8_2),.clk(gclk));
	jdff dff_B_HJa9TXUS7_2(.din(w_dff_B_TEBdbmRm8_2),.dout(w_dff_B_HJa9TXUS7_2),.clk(gclk));
	jdff dff_B_KBNOUwhS6_2(.din(w_dff_B_HJa9TXUS7_2),.dout(w_dff_B_KBNOUwhS6_2),.clk(gclk));
	jdff dff_B_WXsuBGhM2_2(.din(w_dff_B_KBNOUwhS6_2),.dout(w_dff_B_WXsuBGhM2_2),.clk(gclk));
	jdff dff_B_hIgtUtU92_2(.din(w_dff_B_WXsuBGhM2_2),.dout(w_dff_B_hIgtUtU92_2),.clk(gclk));
	jdff dff_B_R8KQHlkm7_2(.din(w_dff_B_hIgtUtU92_2),.dout(w_dff_B_R8KQHlkm7_2),.clk(gclk));
	jdff dff_B_uCaSF1VP0_2(.din(w_dff_B_R8KQHlkm7_2),.dout(w_dff_B_uCaSF1VP0_2),.clk(gclk));
	jdff dff_B_sAONswcD3_2(.din(w_dff_B_uCaSF1VP0_2),.dout(w_dff_B_sAONswcD3_2),.clk(gclk));
	jdff dff_B_hPr8WnV05_2(.din(w_dff_B_sAONswcD3_2),.dout(w_dff_B_hPr8WnV05_2),.clk(gclk));
	jdff dff_B_AxSNxK3Y9_2(.din(w_dff_B_hPr8WnV05_2),.dout(w_dff_B_AxSNxK3Y9_2),.clk(gclk));
	jdff dff_B_RFXlgBXa0_2(.din(n805),.dout(w_dff_B_RFXlgBXa0_2),.clk(gclk));
	jdff dff_B_0sWTkjSX6_1(.din(n783),.dout(w_dff_B_0sWTkjSX6_1),.clk(gclk));
	jdff dff_B_Nw7rkneU4_2(.din(n689),.dout(w_dff_B_Nw7rkneU4_2),.clk(gclk));
	jdff dff_B_aX5oDOtj1_2(.din(w_dff_B_Nw7rkneU4_2),.dout(w_dff_B_aX5oDOtj1_2),.clk(gclk));
	jdff dff_B_gRw1XyA56_2(.din(w_dff_B_aX5oDOtj1_2),.dout(w_dff_B_gRw1XyA56_2),.clk(gclk));
	jdff dff_B_ri45ITj27_2(.din(w_dff_B_gRw1XyA56_2),.dout(w_dff_B_ri45ITj27_2),.clk(gclk));
	jdff dff_B_0SiDLvBJ1_2(.din(w_dff_B_ri45ITj27_2),.dout(w_dff_B_0SiDLvBJ1_2),.clk(gclk));
	jdff dff_B_0WmB5jlO3_2(.din(w_dff_B_0SiDLvBJ1_2),.dout(w_dff_B_0WmB5jlO3_2),.clk(gclk));
	jdff dff_B_q6eho9w43_2(.din(w_dff_B_0WmB5jlO3_2),.dout(w_dff_B_q6eho9w43_2),.clk(gclk));
	jdff dff_B_sMHNr9xq6_2(.din(w_dff_B_q6eho9w43_2),.dout(w_dff_B_sMHNr9xq6_2),.clk(gclk));
	jdff dff_B_3vDR8Cz34_2(.din(w_dff_B_sMHNr9xq6_2),.dout(w_dff_B_3vDR8Cz34_2),.clk(gclk));
	jdff dff_B_rAYZzfgx4_2(.din(n705),.dout(w_dff_B_rAYZzfgx4_2),.clk(gclk));
	jdff dff_B_zqjynpTp0_2(.din(w_dff_B_rAYZzfgx4_2),.dout(w_dff_B_zqjynpTp0_2),.clk(gclk));
	jdff dff_B_f5CxgFtA9_1(.din(n690),.dout(w_dff_B_f5CxgFtA9_1),.clk(gclk));
	jdff dff_B_PdCCOk0H0_1(.din(w_dff_B_f5CxgFtA9_1),.dout(w_dff_B_PdCCOk0H0_1),.clk(gclk));
	jdff dff_B_ZcJnCOHM2_1(.din(w_dff_B_PdCCOk0H0_1),.dout(w_dff_B_ZcJnCOHM2_1),.clk(gclk));
	jdff dff_B_3NgXzHpP7_1(.din(w_dff_B_ZcJnCOHM2_1),.dout(w_dff_B_3NgXzHpP7_1),.clk(gclk));
	jdff dff_B_kZNmdq1V6_1(.din(w_dff_B_3NgXzHpP7_1),.dout(w_dff_B_kZNmdq1V6_1),.clk(gclk));
	jdff dff_B_1BovEjzp0_1(.din(w_dff_B_kZNmdq1V6_1),.dout(w_dff_B_1BovEjzp0_1),.clk(gclk));
	jdff dff_B_PFpMQHd80_0(.din(n612),.dout(w_dff_B_PFpMQHd80_0),.clk(gclk));
	jdff dff_B_oqDe2AjM2_0(.din(w_dff_B_PFpMQHd80_0),.dout(w_dff_B_oqDe2AjM2_0),.clk(gclk));
	jdff dff_A_z98Y48qf6_0(.dout(w_n611_0[0]),.din(w_dff_A_z98Y48qf6_0),.clk(gclk));
	jdff dff_A_d6xTdqEj1_0(.dout(w_dff_A_z98Y48qf6_0),.din(w_dff_A_d6xTdqEj1_0),.clk(gclk));
	jdff dff_A_p1ExIVA06_0(.dout(w_dff_A_d6xTdqEj1_0),.din(w_dff_A_p1ExIVA06_0),.clk(gclk));
	jdff dff_B_TWlLduFk8_1(.din(n605),.dout(w_dff_B_TWlLduFk8_1),.clk(gclk));
	jdff dff_A_okRv4hTg5_0(.dout(w_n523_0[0]),.din(w_dff_A_okRv4hTg5_0),.clk(gclk));
	jdff dff_A_DVRWxS9i3_1(.dout(w_n523_0[1]),.din(w_dff_A_DVRWxS9i3_1),.clk(gclk));
	jdff dff_A_w7exM3Ua5_1(.dout(w_dff_A_DVRWxS9i3_1),.din(w_dff_A_w7exM3Ua5_1),.clk(gclk));
	jdff dff_A_LWJKdsaV1_1(.dout(w_n603_0[1]),.din(w_dff_A_LWJKdsaV1_1),.clk(gclk));
	jdff dff_A_uvCOXY9n2_1(.dout(w_dff_A_LWJKdsaV1_1),.din(w_dff_A_uvCOXY9n2_1),.clk(gclk));
	jdff dff_A_Eai8yYZ14_1(.dout(w_dff_A_uvCOXY9n2_1),.din(w_dff_A_Eai8yYZ14_1),.clk(gclk));
	jdff dff_A_9Ad9Y1rS2_1(.dout(w_dff_A_Eai8yYZ14_1),.din(w_dff_A_9Ad9Y1rS2_1),.clk(gclk));
	jdff dff_A_rB9uUE8L9_1(.dout(w_dff_A_9Ad9Y1rS2_1),.din(w_dff_A_rB9uUE8L9_1),.clk(gclk));
	jdff dff_A_uAiNKDt00_1(.dout(w_dff_A_rB9uUE8L9_1),.din(w_dff_A_uAiNKDt00_1),.clk(gclk));
	jdff dff_B_zTqoFgxU7_1(.din(n1793),.dout(w_dff_B_zTqoFgxU7_1),.clk(gclk));
	jdff dff_A_9n7XV7sv6_1(.dout(w_n1768_0[1]),.din(w_dff_A_9n7XV7sv6_1),.clk(gclk));
	jdff dff_B_K1E8wuCf6_1(.din(n1766),.dout(w_dff_B_K1E8wuCf6_1),.clk(gclk));
	jdff dff_B_SkQNsE0M6_2(.din(n1730),.dout(w_dff_B_SkQNsE0M6_2),.clk(gclk));
	jdff dff_B_w3i1aKTt9_2(.din(w_dff_B_SkQNsE0M6_2),.dout(w_dff_B_w3i1aKTt9_2),.clk(gclk));
	jdff dff_B_hCIO0l0H0_2(.din(w_dff_B_w3i1aKTt9_2),.dout(w_dff_B_hCIO0l0H0_2),.clk(gclk));
	jdff dff_B_HUsAG0Bc3_2(.din(w_dff_B_hCIO0l0H0_2),.dout(w_dff_B_HUsAG0Bc3_2),.clk(gclk));
	jdff dff_B_sDwQ91w46_2(.din(w_dff_B_HUsAG0Bc3_2),.dout(w_dff_B_sDwQ91w46_2),.clk(gclk));
	jdff dff_B_JuYwKgke5_2(.din(w_dff_B_sDwQ91w46_2),.dout(w_dff_B_JuYwKgke5_2),.clk(gclk));
	jdff dff_B_yZashIj38_2(.din(w_dff_B_JuYwKgke5_2),.dout(w_dff_B_yZashIj38_2),.clk(gclk));
	jdff dff_B_DWfgVCHX7_2(.din(w_dff_B_yZashIj38_2),.dout(w_dff_B_DWfgVCHX7_2),.clk(gclk));
	jdff dff_B_Yc5Rit5X9_2(.din(w_dff_B_DWfgVCHX7_2),.dout(w_dff_B_Yc5Rit5X9_2),.clk(gclk));
	jdff dff_B_aqevY56E3_2(.din(w_dff_B_Yc5Rit5X9_2),.dout(w_dff_B_aqevY56E3_2),.clk(gclk));
	jdff dff_B_1izovzXb4_2(.din(w_dff_B_aqevY56E3_2),.dout(w_dff_B_1izovzXb4_2),.clk(gclk));
	jdff dff_B_xk8K3NKn4_2(.din(w_dff_B_1izovzXb4_2),.dout(w_dff_B_xk8K3NKn4_2),.clk(gclk));
	jdff dff_B_NW2TZ1SI7_2(.din(w_dff_B_xk8K3NKn4_2),.dout(w_dff_B_NW2TZ1SI7_2),.clk(gclk));
	jdff dff_B_ow8MaT5U3_2(.din(w_dff_B_NW2TZ1SI7_2),.dout(w_dff_B_ow8MaT5U3_2),.clk(gclk));
	jdff dff_B_ok1lrZg16_2(.din(w_dff_B_ow8MaT5U3_2),.dout(w_dff_B_ok1lrZg16_2),.clk(gclk));
	jdff dff_B_YljKQU2P6_2(.din(w_dff_B_ok1lrZg16_2),.dout(w_dff_B_YljKQU2P6_2),.clk(gclk));
	jdff dff_B_YqoBb55R4_2(.din(w_dff_B_YljKQU2P6_2),.dout(w_dff_B_YqoBb55R4_2),.clk(gclk));
	jdff dff_B_ekYBECWE4_2(.din(w_dff_B_YqoBb55R4_2),.dout(w_dff_B_ekYBECWE4_2),.clk(gclk));
	jdff dff_B_vnu85MWu4_2(.din(w_dff_B_ekYBECWE4_2),.dout(w_dff_B_vnu85MWu4_2),.clk(gclk));
	jdff dff_B_KumHp6UV7_2(.din(w_dff_B_vnu85MWu4_2),.dout(w_dff_B_KumHp6UV7_2),.clk(gclk));
	jdff dff_B_G3nIlvgo2_2(.din(w_dff_B_KumHp6UV7_2),.dout(w_dff_B_G3nIlvgo2_2),.clk(gclk));
	jdff dff_B_MY3V3YK05_2(.din(w_dff_B_G3nIlvgo2_2),.dout(w_dff_B_MY3V3YK05_2),.clk(gclk));
	jdff dff_B_wgqfjphk6_2(.din(w_dff_B_MY3V3YK05_2),.dout(w_dff_B_wgqfjphk6_2),.clk(gclk));
	jdff dff_B_SQUwVAfB3_2(.din(w_dff_B_wgqfjphk6_2),.dout(w_dff_B_SQUwVAfB3_2),.clk(gclk));
	jdff dff_B_6A4tvn5k5_2(.din(w_dff_B_SQUwVAfB3_2),.dout(w_dff_B_6A4tvn5k5_2),.clk(gclk));
	jdff dff_B_6P8tyPpl9_2(.din(w_dff_B_6A4tvn5k5_2),.dout(w_dff_B_6P8tyPpl9_2),.clk(gclk));
	jdff dff_B_J8XDlvFm4_2(.din(w_dff_B_6P8tyPpl9_2),.dout(w_dff_B_J8XDlvFm4_2),.clk(gclk));
	jdff dff_B_c7t0rdZN5_2(.din(w_dff_B_J8XDlvFm4_2),.dout(w_dff_B_c7t0rdZN5_2),.clk(gclk));
	jdff dff_B_hBHlLwk92_2(.din(w_dff_B_c7t0rdZN5_2),.dout(w_dff_B_hBHlLwk92_2),.clk(gclk));
	jdff dff_B_1GkWyzn78_2(.din(w_dff_B_hBHlLwk92_2),.dout(w_dff_B_1GkWyzn78_2),.clk(gclk));
	jdff dff_B_JxF8Aspo5_2(.din(w_dff_B_1GkWyzn78_2),.dout(w_dff_B_JxF8Aspo5_2),.clk(gclk));
	jdff dff_B_UvdGenDh4_2(.din(w_dff_B_JxF8Aspo5_2),.dout(w_dff_B_UvdGenDh4_2),.clk(gclk));
	jdff dff_B_evC6RRMu9_2(.din(w_dff_B_UvdGenDh4_2),.dout(w_dff_B_evC6RRMu9_2),.clk(gclk));
	jdff dff_B_6FPuRBBm1_2(.din(w_dff_B_evC6RRMu9_2),.dout(w_dff_B_6FPuRBBm1_2),.clk(gclk));
	jdff dff_B_MzHYpbmN9_2(.din(w_dff_B_6FPuRBBm1_2),.dout(w_dff_B_MzHYpbmN9_2),.clk(gclk));
	jdff dff_B_691UAJeL7_2(.din(w_dff_B_MzHYpbmN9_2),.dout(w_dff_B_691UAJeL7_2),.clk(gclk));
	jdff dff_B_VPRZIXJZ7_2(.din(w_dff_B_691UAJeL7_2),.dout(w_dff_B_VPRZIXJZ7_2),.clk(gclk));
	jdff dff_B_DtWwtbae9_2(.din(w_dff_B_VPRZIXJZ7_2),.dout(w_dff_B_DtWwtbae9_2),.clk(gclk));
	jdff dff_B_flGWL8Yd0_2(.din(w_dff_B_DtWwtbae9_2),.dout(w_dff_B_flGWL8Yd0_2),.clk(gclk));
	jdff dff_B_0b1gWJAs8_2(.din(w_dff_B_flGWL8Yd0_2),.dout(w_dff_B_0b1gWJAs8_2),.clk(gclk));
	jdff dff_B_aMeCVaG10_2(.din(w_dff_B_0b1gWJAs8_2),.dout(w_dff_B_aMeCVaG10_2),.clk(gclk));
	jdff dff_B_AhiHYvNf7_2(.din(w_dff_B_aMeCVaG10_2),.dout(w_dff_B_AhiHYvNf7_2),.clk(gclk));
	jdff dff_B_5uCvNK794_2(.din(w_dff_B_AhiHYvNf7_2),.dout(w_dff_B_5uCvNK794_2),.clk(gclk));
	jdff dff_B_Ha2VZqoK3_2(.din(w_dff_B_5uCvNK794_2),.dout(w_dff_B_Ha2VZqoK3_2),.clk(gclk));
	jdff dff_B_usbleS4f2_2(.din(w_dff_B_Ha2VZqoK3_2),.dout(w_dff_B_usbleS4f2_2),.clk(gclk));
	jdff dff_B_omIE2QMI7_2(.din(w_dff_B_usbleS4f2_2),.dout(w_dff_B_omIE2QMI7_2),.clk(gclk));
	jdff dff_B_T22nB26N6_2(.din(w_dff_B_omIE2QMI7_2),.dout(w_dff_B_T22nB26N6_2),.clk(gclk));
	jdff dff_B_Jky6HVNF1_2(.din(w_dff_B_T22nB26N6_2),.dout(w_dff_B_Jky6HVNF1_2),.clk(gclk));
	jdff dff_B_8qzRylMw2_2(.din(w_dff_B_Jky6HVNF1_2),.dout(w_dff_B_8qzRylMw2_2),.clk(gclk));
	jdff dff_B_wLlSA1MN9_2(.din(w_dff_B_8qzRylMw2_2),.dout(w_dff_B_wLlSA1MN9_2),.clk(gclk));
	jdff dff_B_YqZFdzjd8_2(.din(w_dff_B_wLlSA1MN9_2),.dout(w_dff_B_YqZFdzjd8_2),.clk(gclk));
	jdff dff_B_eWqtMJtR2_2(.din(n1733),.dout(w_dff_B_eWqtMJtR2_2),.clk(gclk));
	jdff dff_B_tYvUEpmN3_1(.din(n1731),.dout(w_dff_B_tYvUEpmN3_1),.clk(gclk));
	jdff dff_B_xjz1kvxf4_2(.din(n1689),.dout(w_dff_B_xjz1kvxf4_2),.clk(gclk));
	jdff dff_B_UKazAOJP9_2(.din(w_dff_B_xjz1kvxf4_2),.dout(w_dff_B_UKazAOJP9_2),.clk(gclk));
	jdff dff_B_QZTb955o4_2(.din(w_dff_B_UKazAOJP9_2),.dout(w_dff_B_QZTb955o4_2),.clk(gclk));
	jdff dff_B_u8kKB4xi8_2(.din(w_dff_B_QZTb955o4_2),.dout(w_dff_B_u8kKB4xi8_2),.clk(gclk));
	jdff dff_B_WDQG8Xzs0_2(.din(w_dff_B_u8kKB4xi8_2),.dout(w_dff_B_WDQG8Xzs0_2),.clk(gclk));
	jdff dff_B_PNBdtUvD7_2(.din(w_dff_B_WDQG8Xzs0_2),.dout(w_dff_B_PNBdtUvD7_2),.clk(gclk));
	jdff dff_B_8RhFjxJJ7_2(.din(w_dff_B_PNBdtUvD7_2),.dout(w_dff_B_8RhFjxJJ7_2),.clk(gclk));
	jdff dff_B_IQTDBg2f4_2(.din(w_dff_B_8RhFjxJJ7_2),.dout(w_dff_B_IQTDBg2f4_2),.clk(gclk));
	jdff dff_B_ORLxoJ2g3_2(.din(w_dff_B_IQTDBg2f4_2),.dout(w_dff_B_ORLxoJ2g3_2),.clk(gclk));
	jdff dff_B_uLUTfVXl5_2(.din(w_dff_B_ORLxoJ2g3_2),.dout(w_dff_B_uLUTfVXl5_2),.clk(gclk));
	jdff dff_B_hcNAJMin2_2(.din(w_dff_B_uLUTfVXl5_2),.dout(w_dff_B_hcNAJMin2_2),.clk(gclk));
	jdff dff_B_iAY9FUAB4_2(.din(w_dff_B_hcNAJMin2_2),.dout(w_dff_B_iAY9FUAB4_2),.clk(gclk));
	jdff dff_B_bDhbvrd39_2(.din(w_dff_B_iAY9FUAB4_2),.dout(w_dff_B_bDhbvrd39_2),.clk(gclk));
	jdff dff_B_Pz7ULMi99_2(.din(w_dff_B_bDhbvrd39_2),.dout(w_dff_B_Pz7ULMi99_2),.clk(gclk));
	jdff dff_B_3duShExP0_2(.din(w_dff_B_Pz7ULMi99_2),.dout(w_dff_B_3duShExP0_2),.clk(gclk));
	jdff dff_B_0bIIEBpI1_2(.din(w_dff_B_3duShExP0_2),.dout(w_dff_B_0bIIEBpI1_2),.clk(gclk));
	jdff dff_B_nFbHJGNl0_2(.din(w_dff_B_0bIIEBpI1_2),.dout(w_dff_B_nFbHJGNl0_2),.clk(gclk));
	jdff dff_B_lwGAUJsl3_2(.din(w_dff_B_nFbHJGNl0_2),.dout(w_dff_B_lwGAUJsl3_2),.clk(gclk));
	jdff dff_B_BEXyloxr5_2(.din(w_dff_B_lwGAUJsl3_2),.dout(w_dff_B_BEXyloxr5_2),.clk(gclk));
	jdff dff_B_wEf2Nuqw1_2(.din(w_dff_B_BEXyloxr5_2),.dout(w_dff_B_wEf2Nuqw1_2),.clk(gclk));
	jdff dff_B_GlXLRHWq2_2(.din(w_dff_B_wEf2Nuqw1_2),.dout(w_dff_B_GlXLRHWq2_2),.clk(gclk));
	jdff dff_B_KRHJzMcj7_2(.din(w_dff_B_GlXLRHWq2_2),.dout(w_dff_B_KRHJzMcj7_2),.clk(gclk));
	jdff dff_B_gcwYpLyo3_2(.din(w_dff_B_KRHJzMcj7_2),.dout(w_dff_B_gcwYpLyo3_2),.clk(gclk));
	jdff dff_B_eQ0q6MuY7_2(.din(w_dff_B_gcwYpLyo3_2),.dout(w_dff_B_eQ0q6MuY7_2),.clk(gclk));
	jdff dff_B_dENTBUA79_2(.din(w_dff_B_eQ0q6MuY7_2),.dout(w_dff_B_dENTBUA79_2),.clk(gclk));
	jdff dff_B_3dOZS4Kg8_2(.din(w_dff_B_dENTBUA79_2),.dout(w_dff_B_3dOZS4Kg8_2),.clk(gclk));
	jdff dff_B_dsDenCKx9_2(.din(w_dff_B_3dOZS4Kg8_2),.dout(w_dff_B_dsDenCKx9_2),.clk(gclk));
	jdff dff_B_RKUxxegn4_2(.din(w_dff_B_dsDenCKx9_2),.dout(w_dff_B_RKUxxegn4_2),.clk(gclk));
	jdff dff_B_znAGUxhz9_2(.din(w_dff_B_RKUxxegn4_2),.dout(w_dff_B_znAGUxhz9_2),.clk(gclk));
	jdff dff_B_Cif6COd73_2(.din(w_dff_B_znAGUxhz9_2),.dout(w_dff_B_Cif6COd73_2),.clk(gclk));
	jdff dff_B_hJMqL0hB1_2(.din(w_dff_B_Cif6COd73_2),.dout(w_dff_B_hJMqL0hB1_2),.clk(gclk));
	jdff dff_B_4IzAYm0o3_2(.din(w_dff_B_hJMqL0hB1_2),.dout(w_dff_B_4IzAYm0o3_2),.clk(gclk));
	jdff dff_B_C2COPUGV2_2(.din(w_dff_B_4IzAYm0o3_2),.dout(w_dff_B_C2COPUGV2_2),.clk(gclk));
	jdff dff_B_xHxTZdoA7_2(.din(w_dff_B_C2COPUGV2_2),.dout(w_dff_B_xHxTZdoA7_2),.clk(gclk));
	jdff dff_B_FU12nnqy4_2(.din(w_dff_B_xHxTZdoA7_2),.dout(w_dff_B_FU12nnqy4_2),.clk(gclk));
	jdff dff_B_K6mIsrgp0_2(.din(w_dff_B_FU12nnqy4_2),.dout(w_dff_B_K6mIsrgp0_2),.clk(gclk));
	jdff dff_B_BRnou9A14_2(.din(w_dff_B_K6mIsrgp0_2),.dout(w_dff_B_BRnou9A14_2),.clk(gclk));
	jdff dff_B_Rq0sGR780_2(.din(w_dff_B_BRnou9A14_2),.dout(w_dff_B_Rq0sGR780_2),.clk(gclk));
	jdff dff_B_V0WEGXW86_2(.din(w_dff_B_Rq0sGR780_2),.dout(w_dff_B_V0WEGXW86_2),.clk(gclk));
	jdff dff_B_CCNeJ2CH6_2(.din(w_dff_B_V0WEGXW86_2),.dout(w_dff_B_CCNeJ2CH6_2),.clk(gclk));
	jdff dff_B_pXd4sEYr6_2(.din(w_dff_B_CCNeJ2CH6_2),.dout(w_dff_B_pXd4sEYr6_2),.clk(gclk));
	jdff dff_B_avZv5ACW8_2(.din(w_dff_B_pXd4sEYr6_2),.dout(w_dff_B_avZv5ACW8_2),.clk(gclk));
	jdff dff_B_bexQZ2CP0_2(.din(w_dff_B_avZv5ACW8_2),.dout(w_dff_B_bexQZ2CP0_2),.clk(gclk));
	jdff dff_B_X1U51X8C8_2(.din(w_dff_B_bexQZ2CP0_2),.dout(w_dff_B_X1U51X8C8_2),.clk(gclk));
	jdff dff_B_fxO94WAp4_2(.din(w_dff_B_X1U51X8C8_2),.dout(w_dff_B_fxO94WAp4_2),.clk(gclk));
	jdff dff_B_2nJbfz1l7_2(.din(w_dff_B_fxO94WAp4_2),.dout(w_dff_B_2nJbfz1l7_2),.clk(gclk));
	jdff dff_B_wWyQm1T04_2(.din(w_dff_B_2nJbfz1l7_2),.dout(w_dff_B_wWyQm1T04_2),.clk(gclk));
	jdff dff_B_EzRe3tCe8_2(.din(n1692),.dout(w_dff_B_EzRe3tCe8_2),.clk(gclk));
	jdff dff_B_JljeUlJQ0_1(.din(n1690),.dout(w_dff_B_JljeUlJQ0_1),.clk(gclk));
	jdff dff_B_DBqr7t5P3_2(.din(n1638),.dout(w_dff_B_DBqr7t5P3_2),.clk(gclk));
	jdff dff_B_M2vUMp7K1_2(.din(w_dff_B_DBqr7t5P3_2),.dout(w_dff_B_M2vUMp7K1_2),.clk(gclk));
	jdff dff_B_CpigqGl21_2(.din(w_dff_B_M2vUMp7K1_2),.dout(w_dff_B_CpigqGl21_2),.clk(gclk));
	jdff dff_B_WNmUCUVW1_2(.din(w_dff_B_CpigqGl21_2),.dout(w_dff_B_WNmUCUVW1_2),.clk(gclk));
	jdff dff_B_wAIm0fYC7_2(.din(w_dff_B_WNmUCUVW1_2),.dout(w_dff_B_wAIm0fYC7_2),.clk(gclk));
	jdff dff_B_bGz67cqn3_2(.din(w_dff_B_wAIm0fYC7_2),.dout(w_dff_B_bGz67cqn3_2),.clk(gclk));
	jdff dff_B_gpBi5Byj0_2(.din(w_dff_B_bGz67cqn3_2),.dout(w_dff_B_gpBi5Byj0_2),.clk(gclk));
	jdff dff_B_gzDQXrBx2_2(.din(w_dff_B_gpBi5Byj0_2),.dout(w_dff_B_gzDQXrBx2_2),.clk(gclk));
	jdff dff_B_BnwCrT4V8_2(.din(w_dff_B_gzDQXrBx2_2),.dout(w_dff_B_BnwCrT4V8_2),.clk(gclk));
	jdff dff_B_MZ78ol9p4_2(.din(w_dff_B_BnwCrT4V8_2),.dout(w_dff_B_MZ78ol9p4_2),.clk(gclk));
	jdff dff_B_64QAvVpK5_2(.din(w_dff_B_MZ78ol9p4_2),.dout(w_dff_B_64QAvVpK5_2),.clk(gclk));
	jdff dff_B_T2tIO3I22_2(.din(w_dff_B_64QAvVpK5_2),.dout(w_dff_B_T2tIO3I22_2),.clk(gclk));
	jdff dff_B_Xk6LG3D73_2(.din(w_dff_B_T2tIO3I22_2),.dout(w_dff_B_Xk6LG3D73_2),.clk(gclk));
	jdff dff_B_i1Z1PAty5_2(.din(w_dff_B_Xk6LG3D73_2),.dout(w_dff_B_i1Z1PAty5_2),.clk(gclk));
	jdff dff_B_6sv6gaOj2_2(.din(w_dff_B_i1Z1PAty5_2),.dout(w_dff_B_6sv6gaOj2_2),.clk(gclk));
	jdff dff_B_DAj1jKV31_2(.din(w_dff_B_6sv6gaOj2_2),.dout(w_dff_B_DAj1jKV31_2),.clk(gclk));
	jdff dff_B_ZxYpR0Ov1_2(.din(w_dff_B_DAj1jKV31_2),.dout(w_dff_B_ZxYpR0Ov1_2),.clk(gclk));
	jdff dff_B_yPsvRPbX9_2(.din(w_dff_B_ZxYpR0Ov1_2),.dout(w_dff_B_yPsvRPbX9_2),.clk(gclk));
	jdff dff_B_gcJvnEP77_2(.din(w_dff_B_yPsvRPbX9_2),.dout(w_dff_B_gcJvnEP77_2),.clk(gclk));
	jdff dff_B_6GfsG9kL5_2(.din(w_dff_B_gcJvnEP77_2),.dout(w_dff_B_6GfsG9kL5_2),.clk(gclk));
	jdff dff_B_07glfzRU9_2(.din(w_dff_B_6GfsG9kL5_2),.dout(w_dff_B_07glfzRU9_2),.clk(gclk));
	jdff dff_B_YDRyvsVQ5_2(.din(w_dff_B_07glfzRU9_2),.dout(w_dff_B_YDRyvsVQ5_2),.clk(gclk));
	jdff dff_B_VJRMPvHG5_2(.din(w_dff_B_YDRyvsVQ5_2),.dout(w_dff_B_VJRMPvHG5_2),.clk(gclk));
	jdff dff_B_Xk2AC1qs0_2(.din(w_dff_B_VJRMPvHG5_2),.dout(w_dff_B_Xk2AC1qs0_2),.clk(gclk));
	jdff dff_B_X5ev7AnE6_2(.din(w_dff_B_Xk2AC1qs0_2),.dout(w_dff_B_X5ev7AnE6_2),.clk(gclk));
	jdff dff_B_AKFIMH0n2_2(.din(w_dff_B_X5ev7AnE6_2),.dout(w_dff_B_AKFIMH0n2_2),.clk(gclk));
	jdff dff_B_RUUmnh4T6_2(.din(w_dff_B_AKFIMH0n2_2),.dout(w_dff_B_RUUmnh4T6_2),.clk(gclk));
	jdff dff_B_KEa06emA7_2(.din(w_dff_B_RUUmnh4T6_2),.dout(w_dff_B_KEa06emA7_2),.clk(gclk));
	jdff dff_B_xXSYyKvA2_2(.din(w_dff_B_KEa06emA7_2),.dout(w_dff_B_xXSYyKvA2_2),.clk(gclk));
	jdff dff_B_iI8u8BKe5_2(.din(w_dff_B_xXSYyKvA2_2),.dout(w_dff_B_iI8u8BKe5_2),.clk(gclk));
	jdff dff_B_UjUHYEMc3_2(.din(w_dff_B_iI8u8BKe5_2),.dout(w_dff_B_UjUHYEMc3_2),.clk(gclk));
	jdff dff_B_6bZtp23N2_2(.din(w_dff_B_UjUHYEMc3_2),.dout(w_dff_B_6bZtp23N2_2),.clk(gclk));
	jdff dff_B_C2SozrwU2_2(.din(w_dff_B_6bZtp23N2_2),.dout(w_dff_B_C2SozrwU2_2),.clk(gclk));
	jdff dff_B_NFZfAwyU8_2(.din(w_dff_B_C2SozrwU2_2),.dout(w_dff_B_NFZfAwyU8_2),.clk(gclk));
	jdff dff_B_WQKBUYiM7_2(.din(w_dff_B_NFZfAwyU8_2),.dout(w_dff_B_WQKBUYiM7_2),.clk(gclk));
	jdff dff_B_2Js7OGcF1_2(.din(w_dff_B_WQKBUYiM7_2),.dout(w_dff_B_2Js7OGcF1_2),.clk(gclk));
	jdff dff_B_2Q56mQTX6_2(.din(w_dff_B_2Js7OGcF1_2),.dout(w_dff_B_2Q56mQTX6_2),.clk(gclk));
	jdff dff_B_oirdcrNs4_2(.din(w_dff_B_2Q56mQTX6_2),.dout(w_dff_B_oirdcrNs4_2),.clk(gclk));
	jdff dff_B_6e6IMxZ20_2(.din(w_dff_B_oirdcrNs4_2),.dout(w_dff_B_6e6IMxZ20_2),.clk(gclk));
	jdff dff_B_NeaCHM014_2(.din(w_dff_B_6e6IMxZ20_2),.dout(w_dff_B_NeaCHM014_2),.clk(gclk));
	jdff dff_B_K1KHXBW88_2(.din(w_dff_B_NeaCHM014_2),.dout(w_dff_B_K1KHXBW88_2),.clk(gclk));
	jdff dff_B_ChUkjOSL6_2(.din(w_dff_B_K1KHXBW88_2),.dout(w_dff_B_ChUkjOSL6_2),.clk(gclk));
	jdff dff_B_dz0k26vB2_2(.din(w_dff_B_ChUkjOSL6_2),.dout(w_dff_B_dz0k26vB2_2),.clk(gclk));
	jdff dff_B_tEmEHAdO5_2(.din(n1641),.dout(w_dff_B_tEmEHAdO5_2),.clk(gclk));
	jdff dff_B_PuxHg3Gn7_1(.din(n1639),.dout(w_dff_B_PuxHg3Gn7_1),.clk(gclk));
	jdff dff_B_NiV5Ry3s4_2(.din(n1581),.dout(w_dff_B_NiV5Ry3s4_2),.clk(gclk));
	jdff dff_B_MbTDFteX9_2(.din(w_dff_B_NiV5Ry3s4_2),.dout(w_dff_B_MbTDFteX9_2),.clk(gclk));
	jdff dff_B_z9ZR1lCT3_2(.din(w_dff_B_MbTDFteX9_2),.dout(w_dff_B_z9ZR1lCT3_2),.clk(gclk));
	jdff dff_B_cBvxXdsU4_2(.din(w_dff_B_z9ZR1lCT3_2),.dout(w_dff_B_cBvxXdsU4_2),.clk(gclk));
	jdff dff_B_cLGkST2x8_2(.din(w_dff_B_cBvxXdsU4_2),.dout(w_dff_B_cLGkST2x8_2),.clk(gclk));
	jdff dff_B_Ut6etf7H3_2(.din(w_dff_B_cLGkST2x8_2),.dout(w_dff_B_Ut6etf7H3_2),.clk(gclk));
	jdff dff_B_KA75vRZH2_2(.din(w_dff_B_Ut6etf7H3_2),.dout(w_dff_B_KA75vRZH2_2),.clk(gclk));
	jdff dff_B_hhQWxWsW0_2(.din(w_dff_B_KA75vRZH2_2),.dout(w_dff_B_hhQWxWsW0_2),.clk(gclk));
	jdff dff_B_g9cGFbmd5_2(.din(w_dff_B_hhQWxWsW0_2),.dout(w_dff_B_g9cGFbmd5_2),.clk(gclk));
	jdff dff_B_n4Th0laP3_2(.din(w_dff_B_g9cGFbmd5_2),.dout(w_dff_B_n4Th0laP3_2),.clk(gclk));
	jdff dff_B_xuof9Mpq7_2(.din(w_dff_B_n4Th0laP3_2),.dout(w_dff_B_xuof9Mpq7_2),.clk(gclk));
	jdff dff_B_7XlAPCrD7_2(.din(w_dff_B_xuof9Mpq7_2),.dout(w_dff_B_7XlAPCrD7_2),.clk(gclk));
	jdff dff_B_OAyvb5cV0_2(.din(w_dff_B_7XlAPCrD7_2),.dout(w_dff_B_OAyvb5cV0_2),.clk(gclk));
	jdff dff_B_jazKxcXp4_2(.din(w_dff_B_OAyvb5cV0_2),.dout(w_dff_B_jazKxcXp4_2),.clk(gclk));
	jdff dff_B_Al86i8bD1_2(.din(w_dff_B_jazKxcXp4_2),.dout(w_dff_B_Al86i8bD1_2),.clk(gclk));
	jdff dff_B_AlLf2q5C1_2(.din(w_dff_B_Al86i8bD1_2),.dout(w_dff_B_AlLf2q5C1_2),.clk(gclk));
	jdff dff_B_ZItTtAfd6_2(.din(w_dff_B_AlLf2q5C1_2),.dout(w_dff_B_ZItTtAfd6_2),.clk(gclk));
	jdff dff_B_JMKddtrc4_2(.din(w_dff_B_ZItTtAfd6_2),.dout(w_dff_B_JMKddtrc4_2),.clk(gclk));
	jdff dff_B_ACa5mpu87_2(.din(w_dff_B_JMKddtrc4_2),.dout(w_dff_B_ACa5mpu87_2),.clk(gclk));
	jdff dff_B_SGuNUVAz9_2(.din(w_dff_B_ACa5mpu87_2),.dout(w_dff_B_SGuNUVAz9_2),.clk(gclk));
	jdff dff_B_nZCvjOUe4_2(.din(w_dff_B_SGuNUVAz9_2),.dout(w_dff_B_nZCvjOUe4_2),.clk(gclk));
	jdff dff_B_7AFXXhwe9_2(.din(w_dff_B_nZCvjOUe4_2),.dout(w_dff_B_7AFXXhwe9_2),.clk(gclk));
	jdff dff_B_FLGJ8WNf6_2(.din(w_dff_B_7AFXXhwe9_2),.dout(w_dff_B_FLGJ8WNf6_2),.clk(gclk));
	jdff dff_B_yLdseEDo5_2(.din(w_dff_B_FLGJ8WNf6_2),.dout(w_dff_B_yLdseEDo5_2),.clk(gclk));
	jdff dff_B_7057YDcd2_2(.din(w_dff_B_yLdseEDo5_2),.dout(w_dff_B_7057YDcd2_2),.clk(gclk));
	jdff dff_B_y4Yu8g8X3_2(.din(w_dff_B_7057YDcd2_2),.dout(w_dff_B_y4Yu8g8X3_2),.clk(gclk));
	jdff dff_B_Gl3NF1rb1_2(.din(w_dff_B_y4Yu8g8X3_2),.dout(w_dff_B_Gl3NF1rb1_2),.clk(gclk));
	jdff dff_B_e8DEKZqL1_2(.din(w_dff_B_Gl3NF1rb1_2),.dout(w_dff_B_e8DEKZqL1_2),.clk(gclk));
	jdff dff_B_xqymBRys9_2(.din(w_dff_B_e8DEKZqL1_2),.dout(w_dff_B_xqymBRys9_2),.clk(gclk));
	jdff dff_B_wxedBgbg0_2(.din(w_dff_B_xqymBRys9_2),.dout(w_dff_B_wxedBgbg0_2),.clk(gclk));
	jdff dff_B_2VWZ8N0X9_2(.din(w_dff_B_wxedBgbg0_2),.dout(w_dff_B_2VWZ8N0X9_2),.clk(gclk));
	jdff dff_B_LY4kAkbG8_2(.din(w_dff_B_2VWZ8N0X9_2),.dout(w_dff_B_LY4kAkbG8_2),.clk(gclk));
	jdff dff_B_o6OC3ZCQ1_2(.din(w_dff_B_LY4kAkbG8_2),.dout(w_dff_B_o6OC3ZCQ1_2),.clk(gclk));
	jdff dff_B_XdqYoZuF3_2(.din(w_dff_B_o6OC3ZCQ1_2),.dout(w_dff_B_XdqYoZuF3_2),.clk(gclk));
	jdff dff_B_jAHP4GMu9_2(.din(w_dff_B_XdqYoZuF3_2),.dout(w_dff_B_jAHP4GMu9_2),.clk(gclk));
	jdff dff_B_NVPOjIt99_2(.din(w_dff_B_jAHP4GMu9_2),.dout(w_dff_B_NVPOjIt99_2),.clk(gclk));
	jdff dff_B_iW66WLK87_2(.din(w_dff_B_NVPOjIt99_2),.dout(w_dff_B_iW66WLK87_2),.clk(gclk));
	jdff dff_B_VEHPxe3j2_2(.din(w_dff_B_iW66WLK87_2),.dout(w_dff_B_VEHPxe3j2_2),.clk(gclk));
	jdff dff_B_Sddow3bz4_2(.din(w_dff_B_VEHPxe3j2_2),.dout(w_dff_B_Sddow3bz4_2),.clk(gclk));
	jdff dff_B_LAskapZm5_2(.din(n1584),.dout(w_dff_B_LAskapZm5_2),.clk(gclk));
	jdff dff_B_OAaZjvPj1_1(.din(n1582),.dout(w_dff_B_OAaZjvPj1_1),.clk(gclk));
	jdff dff_B_YvArSvkU1_2(.din(n1517),.dout(w_dff_B_YvArSvkU1_2),.clk(gclk));
	jdff dff_B_9Amf4eFI1_2(.din(w_dff_B_YvArSvkU1_2),.dout(w_dff_B_9Amf4eFI1_2),.clk(gclk));
	jdff dff_B_b1Yq46iO8_2(.din(w_dff_B_9Amf4eFI1_2),.dout(w_dff_B_b1Yq46iO8_2),.clk(gclk));
	jdff dff_B_PBDpsqR14_2(.din(w_dff_B_b1Yq46iO8_2),.dout(w_dff_B_PBDpsqR14_2),.clk(gclk));
	jdff dff_B_dt0BS1H90_2(.din(w_dff_B_PBDpsqR14_2),.dout(w_dff_B_dt0BS1H90_2),.clk(gclk));
	jdff dff_B_tejImq9y6_2(.din(w_dff_B_dt0BS1H90_2),.dout(w_dff_B_tejImq9y6_2),.clk(gclk));
	jdff dff_B_5dEDRGNQ8_2(.din(w_dff_B_tejImq9y6_2),.dout(w_dff_B_5dEDRGNQ8_2),.clk(gclk));
	jdff dff_B_X2H6td5e5_2(.din(w_dff_B_5dEDRGNQ8_2),.dout(w_dff_B_X2H6td5e5_2),.clk(gclk));
	jdff dff_B_pTLxAzCZ9_2(.din(w_dff_B_X2H6td5e5_2),.dout(w_dff_B_pTLxAzCZ9_2),.clk(gclk));
	jdff dff_B_GDvjLGlX3_2(.din(w_dff_B_pTLxAzCZ9_2),.dout(w_dff_B_GDvjLGlX3_2),.clk(gclk));
	jdff dff_B_EN1qjhzT2_2(.din(w_dff_B_GDvjLGlX3_2),.dout(w_dff_B_EN1qjhzT2_2),.clk(gclk));
	jdff dff_B_VmMD9niZ8_2(.din(w_dff_B_EN1qjhzT2_2),.dout(w_dff_B_VmMD9niZ8_2),.clk(gclk));
	jdff dff_B_a7geb3ul0_2(.din(w_dff_B_VmMD9niZ8_2),.dout(w_dff_B_a7geb3ul0_2),.clk(gclk));
	jdff dff_B_6fKO13WA4_2(.din(w_dff_B_a7geb3ul0_2),.dout(w_dff_B_6fKO13WA4_2),.clk(gclk));
	jdff dff_B_ywRatiSP5_2(.din(w_dff_B_6fKO13WA4_2),.dout(w_dff_B_ywRatiSP5_2),.clk(gclk));
	jdff dff_B_HQ2tvnZ50_2(.din(w_dff_B_ywRatiSP5_2),.dout(w_dff_B_HQ2tvnZ50_2),.clk(gclk));
	jdff dff_B_QG5kuPBS3_2(.din(w_dff_B_HQ2tvnZ50_2),.dout(w_dff_B_QG5kuPBS3_2),.clk(gclk));
	jdff dff_B_CD3OADq45_2(.din(w_dff_B_QG5kuPBS3_2),.dout(w_dff_B_CD3OADq45_2),.clk(gclk));
	jdff dff_B_zYpnQ2Ig0_2(.din(w_dff_B_CD3OADq45_2),.dout(w_dff_B_zYpnQ2Ig0_2),.clk(gclk));
	jdff dff_B_cEGvPtLY2_2(.din(w_dff_B_zYpnQ2Ig0_2),.dout(w_dff_B_cEGvPtLY2_2),.clk(gclk));
	jdff dff_B_oirJ4AZ60_2(.din(w_dff_B_cEGvPtLY2_2),.dout(w_dff_B_oirJ4AZ60_2),.clk(gclk));
	jdff dff_B_hGizR7cq6_2(.din(w_dff_B_oirJ4AZ60_2),.dout(w_dff_B_hGizR7cq6_2),.clk(gclk));
	jdff dff_B_qJeZbiVS0_2(.din(w_dff_B_hGizR7cq6_2),.dout(w_dff_B_qJeZbiVS0_2),.clk(gclk));
	jdff dff_B_SV8i3JPX5_2(.din(w_dff_B_qJeZbiVS0_2),.dout(w_dff_B_SV8i3JPX5_2),.clk(gclk));
	jdff dff_B_cDQJ7fM50_2(.din(w_dff_B_SV8i3JPX5_2),.dout(w_dff_B_cDQJ7fM50_2),.clk(gclk));
	jdff dff_B_P5cb6zY73_2(.din(w_dff_B_cDQJ7fM50_2),.dout(w_dff_B_P5cb6zY73_2),.clk(gclk));
	jdff dff_B_vDXw7Xci5_2(.din(w_dff_B_P5cb6zY73_2),.dout(w_dff_B_vDXw7Xci5_2),.clk(gclk));
	jdff dff_B_HqQiNcsV3_2(.din(w_dff_B_vDXw7Xci5_2),.dout(w_dff_B_HqQiNcsV3_2),.clk(gclk));
	jdff dff_B_acsSjEvN0_2(.din(w_dff_B_HqQiNcsV3_2),.dout(w_dff_B_acsSjEvN0_2),.clk(gclk));
	jdff dff_B_hvPFtZkC6_2(.din(w_dff_B_acsSjEvN0_2),.dout(w_dff_B_hvPFtZkC6_2),.clk(gclk));
	jdff dff_B_HciZw9o28_2(.din(w_dff_B_hvPFtZkC6_2),.dout(w_dff_B_HciZw9o28_2),.clk(gclk));
	jdff dff_B_xbllgv9y5_2(.din(w_dff_B_HciZw9o28_2),.dout(w_dff_B_xbllgv9y5_2),.clk(gclk));
	jdff dff_B_hQ5NkmOB9_2(.din(w_dff_B_xbllgv9y5_2),.dout(w_dff_B_hQ5NkmOB9_2),.clk(gclk));
	jdff dff_B_jLRC9c199_2(.din(w_dff_B_hQ5NkmOB9_2),.dout(w_dff_B_jLRC9c199_2),.clk(gclk));
	jdff dff_B_y9GIDU0I4_2(.din(w_dff_B_jLRC9c199_2),.dout(w_dff_B_y9GIDU0I4_2),.clk(gclk));
	jdff dff_B_uIocQ37G6_2(.din(n1520),.dout(w_dff_B_uIocQ37G6_2),.clk(gclk));
	jdff dff_B_ojVnhXCC2_1(.din(n1518),.dout(w_dff_B_ojVnhXCC2_1),.clk(gclk));
	jdff dff_B_daI1jvuT4_2(.din(n1446),.dout(w_dff_B_daI1jvuT4_2),.clk(gclk));
	jdff dff_B_sAPYZK8Y7_2(.din(w_dff_B_daI1jvuT4_2),.dout(w_dff_B_sAPYZK8Y7_2),.clk(gclk));
	jdff dff_B_Gk4uQ0640_2(.din(w_dff_B_sAPYZK8Y7_2),.dout(w_dff_B_Gk4uQ0640_2),.clk(gclk));
	jdff dff_B_LmAKy6Eo2_2(.din(w_dff_B_Gk4uQ0640_2),.dout(w_dff_B_LmAKy6Eo2_2),.clk(gclk));
	jdff dff_B_QrPblEgJ0_2(.din(w_dff_B_LmAKy6Eo2_2),.dout(w_dff_B_QrPblEgJ0_2),.clk(gclk));
	jdff dff_B_207anArg1_2(.din(w_dff_B_QrPblEgJ0_2),.dout(w_dff_B_207anArg1_2),.clk(gclk));
	jdff dff_B_pAbdW2I46_2(.din(w_dff_B_207anArg1_2),.dout(w_dff_B_pAbdW2I46_2),.clk(gclk));
	jdff dff_B_zvHk8ibg3_2(.din(w_dff_B_pAbdW2I46_2),.dout(w_dff_B_zvHk8ibg3_2),.clk(gclk));
	jdff dff_B_lFKr3KxZ5_2(.din(w_dff_B_zvHk8ibg3_2),.dout(w_dff_B_lFKr3KxZ5_2),.clk(gclk));
	jdff dff_B_mlzJ81VE7_2(.din(w_dff_B_lFKr3KxZ5_2),.dout(w_dff_B_mlzJ81VE7_2),.clk(gclk));
	jdff dff_B_jJcPbM4i2_2(.din(w_dff_B_mlzJ81VE7_2),.dout(w_dff_B_jJcPbM4i2_2),.clk(gclk));
	jdff dff_B_LrcQsu8Z2_2(.din(w_dff_B_jJcPbM4i2_2),.dout(w_dff_B_LrcQsu8Z2_2),.clk(gclk));
	jdff dff_B_0GbhOBaB3_2(.din(w_dff_B_LrcQsu8Z2_2),.dout(w_dff_B_0GbhOBaB3_2),.clk(gclk));
	jdff dff_B_9zDx6fE76_2(.din(w_dff_B_0GbhOBaB3_2),.dout(w_dff_B_9zDx6fE76_2),.clk(gclk));
	jdff dff_B_ZaHYn9Kk4_2(.din(w_dff_B_9zDx6fE76_2),.dout(w_dff_B_ZaHYn9Kk4_2),.clk(gclk));
	jdff dff_B_9ggUCfBK7_2(.din(w_dff_B_ZaHYn9Kk4_2),.dout(w_dff_B_9ggUCfBK7_2),.clk(gclk));
	jdff dff_B_zoZRn6Nl4_2(.din(w_dff_B_9ggUCfBK7_2),.dout(w_dff_B_zoZRn6Nl4_2),.clk(gclk));
	jdff dff_B_469OYTAY2_2(.din(w_dff_B_zoZRn6Nl4_2),.dout(w_dff_B_469OYTAY2_2),.clk(gclk));
	jdff dff_B_5e8tB98s3_2(.din(w_dff_B_469OYTAY2_2),.dout(w_dff_B_5e8tB98s3_2),.clk(gclk));
	jdff dff_B_dBNHdffZ6_2(.din(w_dff_B_5e8tB98s3_2),.dout(w_dff_B_dBNHdffZ6_2),.clk(gclk));
	jdff dff_B_THr6khAD3_2(.din(w_dff_B_dBNHdffZ6_2),.dout(w_dff_B_THr6khAD3_2),.clk(gclk));
	jdff dff_B_ybIgZP7g0_2(.din(w_dff_B_THr6khAD3_2),.dout(w_dff_B_ybIgZP7g0_2),.clk(gclk));
	jdff dff_B_uT77OrPm8_2(.din(w_dff_B_ybIgZP7g0_2),.dout(w_dff_B_uT77OrPm8_2),.clk(gclk));
	jdff dff_B_smPQwfaU6_2(.din(w_dff_B_uT77OrPm8_2),.dout(w_dff_B_smPQwfaU6_2),.clk(gclk));
	jdff dff_B_bZB3Cq7N1_2(.din(w_dff_B_smPQwfaU6_2),.dout(w_dff_B_bZB3Cq7N1_2),.clk(gclk));
	jdff dff_B_BWDsVCAw7_2(.din(w_dff_B_bZB3Cq7N1_2),.dout(w_dff_B_BWDsVCAw7_2),.clk(gclk));
	jdff dff_B_b1bbbxGR2_2(.din(w_dff_B_BWDsVCAw7_2),.dout(w_dff_B_b1bbbxGR2_2),.clk(gclk));
	jdff dff_B_QnheOsAk7_2(.din(w_dff_B_b1bbbxGR2_2),.dout(w_dff_B_QnheOsAk7_2),.clk(gclk));
	jdff dff_B_EwS4Zgpp6_2(.din(w_dff_B_QnheOsAk7_2),.dout(w_dff_B_EwS4Zgpp6_2),.clk(gclk));
	jdff dff_B_bJddEd148_2(.din(w_dff_B_EwS4Zgpp6_2),.dout(w_dff_B_bJddEd148_2),.clk(gclk));
	jdff dff_B_StFokFFU0_2(.din(w_dff_B_bJddEd148_2),.dout(w_dff_B_StFokFFU0_2),.clk(gclk));
	jdff dff_B_iLfpviWR0_2(.din(n1449),.dout(w_dff_B_iLfpviWR0_2),.clk(gclk));
	jdff dff_B_t0a1Cb0x2_1(.din(n1447),.dout(w_dff_B_t0a1Cb0x2_1),.clk(gclk));
	jdff dff_B_gbLdcTBz1_2(.din(n1368),.dout(w_dff_B_gbLdcTBz1_2),.clk(gclk));
	jdff dff_B_3yPBi7Xl0_2(.din(w_dff_B_gbLdcTBz1_2),.dout(w_dff_B_3yPBi7Xl0_2),.clk(gclk));
	jdff dff_B_zPcgEp8b9_2(.din(w_dff_B_3yPBi7Xl0_2),.dout(w_dff_B_zPcgEp8b9_2),.clk(gclk));
	jdff dff_B_OCdsBj5S9_2(.din(w_dff_B_zPcgEp8b9_2),.dout(w_dff_B_OCdsBj5S9_2),.clk(gclk));
	jdff dff_B_J1YdYyb88_2(.din(w_dff_B_OCdsBj5S9_2),.dout(w_dff_B_J1YdYyb88_2),.clk(gclk));
	jdff dff_B_RrPFprv53_2(.din(w_dff_B_J1YdYyb88_2),.dout(w_dff_B_RrPFprv53_2),.clk(gclk));
	jdff dff_B_TWY3H4s41_2(.din(w_dff_B_RrPFprv53_2),.dout(w_dff_B_TWY3H4s41_2),.clk(gclk));
	jdff dff_B_8b7HdJju7_2(.din(w_dff_B_TWY3H4s41_2),.dout(w_dff_B_8b7HdJju7_2),.clk(gclk));
	jdff dff_B_5szc8Lyv9_2(.din(w_dff_B_8b7HdJju7_2),.dout(w_dff_B_5szc8Lyv9_2),.clk(gclk));
	jdff dff_B_5prMed0M1_2(.din(w_dff_B_5szc8Lyv9_2),.dout(w_dff_B_5prMed0M1_2),.clk(gclk));
	jdff dff_B_mSexEWmK2_2(.din(w_dff_B_5prMed0M1_2),.dout(w_dff_B_mSexEWmK2_2),.clk(gclk));
	jdff dff_B_Q4r0viye4_2(.din(w_dff_B_mSexEWmK2_2),.dout(w_dff_B_Q4r0viye4_2),.clk(gclk));
	jdff dff_B_J71A9wNR8_2(.din(w_dff_B_Q4r0viye4_2),.dout(w_dff_B_J71A9wNR8_2),.clk(gclk));
	jdff dff_B_RDohniPh7_2(.din(w_dff_B_J71A9wNR8_2),.dout(w_dff_B_RDohniPh7_2),.clk(gclk));
	jdff dff_B_lfFljG9L5_2(.din(w_dff_B_RDohniPh7_2),.dout(w_dff_B_lfFljG9L5_2),.clk(gclk));
	jdff dff_B_lNOsGHfN4_2(.din(w_dff_B_lfFljG9L5_2),.dout(w_dff_B_lNOsGHfN4_2),.clk(gclk));
	jdff dff_B_qH7mVeSB1_2(.din(w_dff_B_lNOsGHfN4_2),.dout(w_dff_B_qH7mVeSB1_2),.clk(gclk));
	jdff dff_B_k7UpXjk40_2(.din(w_dff_B_qH7mVeSB1_2),.dout(w_dff_B_k7UpXjk40_2),.clk(gclk));
	jdff dff_B_gxkE9eGk8_2(.din(w_dff_B_k7UpXjk40_2),.dout(w_dff_B_gxkE9eGk8_2),.clk(gclk));
	jdff dff_B_kTFSDjs02_2(.din(w_dff_B_gxkE9eGk8_2),.dout(w_dff_B_kTFSDjs02_2),.clk(gclk));
	jdff dff_B_KIFSxei32_2(.din(w_dff_B_kTFSDjs02_2),.dout(w_dff_B_KIFSxei32_2),.clk(gclk));
	jdff dff_B_lS8iLh7H7_2(.din(w_dff_B_KIFSxei32_2),.dout(w_dff_B_lS8iLh7H7_2),.clk(gclk));
	jdff dff_B_PQp5RMD44_2(.din(w_dff_B_lS8iLh7H7_2),.dout(w_dff_B_PQp5RMD44_2),.clk(gclk));
	jdff dff_B_0uNv9ZCo7_2(.din(w_dff_B_PQp5RMD44_2),.dout(w_dff_B_0uNv9ZCo7_2),.clk(gclk));
	jdff dff_B_b2HnPl0F6_2(.din(w_dff_B_0uNv9ZCo7_2),.dout(w_dff_B_b2HnPl0F6_2),.clk(gclk));
	jdff dff_B_aIE8N9OT4_2(.din(w_dff_B_b2HnPl0F6_2),.dout(w_dff_B_aIE8N9OT4_2),.clk(gclk));
	jdff dff_B_dOjXQLHZ1_2(.din(w_dff_B_aIE8N9OT4_2),.dout(w_dff_B_dOjXQLHZ1_2),.clk(gclk));
	jdff dff_B_lW6ZkaRh0_1(.din(n1369),.dout(w_dff_B_lW6ZkaRh0_1),.clk(gclk));
	jdff dff_B_G26W0DGU8_2(.din(n1283),.dout(w_dff_B_G26W0DGU8_2),.clk(gclk));
	jdff dff_B_HgZ7q5jk5_2(.din(w_dff_B_G26W0DGU8_2),.dout(w_dff_B_HgZ7q5jk5_2),.clk(gclk));
	jdff dff_B_a5yJQUzD8_2(.din(w_dff_B_HgZ7q5jk5_2),.dout(w_dff_B_a5yJQUzD8_2),.clk(gclk));
	jdff dff_B_o2BMIsvw4_2(.din(w_dff_B_a5yJQUzD8_2),.dout(w_dff_B_o2BMIsvw4_2),.clk(gclk));
	jdff dff_B_K93xpsFb6_2(.din(w_dff_B_o2BMIsvw4_2),.dout(w_dff_B_K93xpsFb6_2),.clk(gclk));
	jdff dff_B_mcofuDX07_2(.din(w_dff_B_K93xpsFb6_2),.dout(w_dff_B_mcofuDX07_2),.clk(gclk));
	jdff dff_B_dxjETRKv3_2(.din(w_dff_B_mcofuDX07_2),.dout(w_dff_B_dxjETRKv3_2),.clk(gclk));
	jdff dff_B_HTWBfWzI0_2(.din(w_dff_B_dxjETRKv3_2),.dout(w_dff_B_HTWBfWzI0_2),.clk(gclk));
	jdff dff_B_g9fWyUSA1_2(.din(w_dff_B_HTWBfWzI0_2),.dout(w_dff_B_g9fWyUSA1_2),.clk(gclk));
	jdff dff_B_uA1SB5e10_2(.din(w_dff_B_g9fWyUSA1_2),.dout(w_dff_B_uA1SB5e10_2),.clk(gclk));
	jdff dff_B_MQj0Ym9K7_2(.din(w_dff_B_uA1SB5e10_2),.dout(w_dff_B_MQj0Ym9K7_2),.clk(gclk));
	jdff dff_B_aSg1ez8S6_2(.din(w_dff_B_MQj0Ym9K7_2),.dout(w_dff_B_aSg1ez8S6_2),.clk(gclk));
	jdff dff_B_DvOTFCWY4_2(.din(w_dff_B_aSg1ez8S6_2),.dout(w_dff_B_DvOTFCWY4_2),.clk(gclk));
	jdff dff_B_e4OMPagk2_2(.din(w_dff_B_DvOTFCWY4_2),.dout(w_dff_B_e4OMPagk2_2),.clk(gclk));
	jdff dff_B_94PG2yZX9_2(.din(w_dff_B_e4OMPagk2_2),.dout(w_dff_B_94PG2yZX9_2),.clk(gclk));
	jdff dff_B_z25d29tI2_2(.din(w_dff_B_94PG2yZX9_2),.dout(w_dff_B_z25d29tI2_2),.clk(gclk));
	jdff dff_B_kxh2SXZf6_2(.din(w_dff_B_z25d29tI2_2),.dout(w_dff_B_kxh2SXZf6_2),.clk(gclk));
	jdff dff_B_bbKUNQuY0_2(.din(w_dff_B_kxh2SXZf6_2),.dout(w_dff_B_bbKUNQuY0_2),.clk(gclk));
	jdff dff_B_Hofe42hk7_2(.din(w_dff_B_bbKUNQuY0_2),.dout(w_dff_B_Hofe42hk7_2),.clk(gclk));
	jdff dff_B_32zujJz23_2(.din(w_dff_B_Hofe42hk7_2),.dout(w_dff_B_32zujJz23_2),.clk(gclk));
	jdff dff_B_14Iop9Gf0_2(.din(w_dff_B_32zujJz23_2),.dout(w_dff_B_14Iop9Gf0_2),.clk(gclk));
	jdff dff_B_VOZWeydZ5_2(.din(w_dff_B_14Iop9Gf0_2),.dout(w_dff_B_VOZWeydZ5_2),.clk(gclk));
	jdff dff_B_f1YkdpU64_2(.din(w_dff_B_VOZWeydZ5_2),.dout(w_dff_B_f1YkdpU64_2),.clk(gclk));
	jdff dff_B_LPIVmATe5_2(.din(w_dff_B_f1YkdpU64_2),.dout(w_dff_B_LPIVmATe5_2),.clk(gclk));
	jdff dff_B_sajY995T2_2(.din(n1308),.dout(w_dff_B_sajY995T2_2),.clk(gclk));
	jdff dff_B_Mq3GucuZ0_1(.din(n1284),.dout(w_dff_B_Mq3GucuZ0_1),.clk(gclk));
	jdff dff_B_FGkQiYP45_2(.din(n1193),.dout(w_dff_B_FGkQiYP45_2),.clk(gclk));
	jdff dff_B_jjTzbVSN0_2(.din(w_dff_B_FGkQiYP45_2),.dout(w_dff_B_jjTzbVSN0_2),.clk(gclk));
	jdff dff_B_GXxEVzKw7_2(.din(w_dff_B_jjTzbVSN0_2),.dout(w_dff_B_GXxEVzKw7_2),.clk(gclk));
	jdff dff_B_AGYJOGDB8_2(.din(w_dff_B_GXxEVzKw7_2),.dout(w_dff_B_AGYJOGDB8_2),.clk(gclk));
	jdff dff_B_FuCZzOor0_2(.din(w_dff_B_AGYJOGDB8_2),.dout(w_dff_B_FuCZzOor0_2),.clk(gclk));
	jdff dff_B_2X6svhfX3_2(.din(w_dff_B_FuCZzOor0_2),.dout(w_dff_B_2X6svhfX3_2),.clk(gclk));
	jdff dff_B_EWTXv7YF9_2(.din(w_dff_B_2X6svhfX3_2),.dout(w_dff_B_EWTXv7YF9_2),.clk(gclk));
	jdff dff_B_POKoi7GG1_2(.din(w_dff_B_EWTXv7YF9_2),.dout(w_dff_B_POKoi7GG1_2),.clk(gclk));
	jdff dff_B_pNkfxMLZ1_2(.din(w_dff_B_POKoi7GG1_2),.dout(w_dff_B_pNkfxMLZ1_2),.clk(gclk));
	jdff dff_B_soEM9Kco3_2(.din(w_dff_B_pNkfxMLZ1_2),.dout(w_dff_B_soEM9Kco3_2),.clk(gclk));
	jdff dff_B_GBbWMwcr4_2(.din(w_dff_B_soEM9Kco3_2),.dout(w_dff_B_GBbWMwcr4_2),.clk(gclk));
	jdff dff_B_f3q3hBLW0_2(.din(w_dff_B_GBbWMwcr4_2),.dout(w_dff_B_f3q3hBLW0_2),.clk(gclk));
	jdff dff_B_TOgBGkuo6_2(.din(w_dff_B_f3q3hBLW0_2),.dout(w_dff_B_TOgBGkuo6_2),.clk(gclk));
	jdff dff_B_xOL9zfQv9_2(.din(w_dff_B_TOgBGkuo6_2),.dout(w_dff_B_xOL9zfQv9_2),.clk(gclk));
	jdff dff_B_MbdUYURa1_2(.din(w_dff_B_xOL9zfQv9_2),.dout(w_dff_B_MbdUYURa1_2),.clk(gclk));
	jdff dff_B_rYVRGUli5_2(.din(w_dff_B_MbdUYURa1_2),.dout(w_dff_B_rYVRGUli5_2),.clk(gclk));
	jdff dff_B_855Ns1t19_2(.din(w_dff_B_rYVRGUli5_2),.dout(w_dff_B_855Ns1t19_2),.clk(gclk));
	jdff dff_B_bRXgNsFt9_2(.din(w_dff_B_855Ns1t19_2),.dout(w_dff_B_bRXgNsFt9_2),.clk(gclk));
	jdff dff_B_UeGESLzn7_2(.din(w_dff_B_bRXgNsFt9_2),.dout(w_dff_B_UeGESLzn7_2),.clk(gclk));
	jdff dff_B_hBlHuSKQ7_2(.din(w_dff_B_UeGESLzn7_2),.dout(w_dff_B_hBlHuSKQ7_2),.clk(gclk));
	jdff dff_B_3zLaC3ht5_2(.din(w_dff_B_hBlHuSKQ7_2),.dout(w_dff_B_3zLaC3ht5_2),.clk(gclk));
	jdff dff_B_ajak31ho7_2(.din(n1217),.dout(w_dff_B_ajak31ho7_2),.clk(gclk));
	jdff dff_B_Qjvy0QeU2_1(.din(n1194),.dout(w_dff_B_Qjvy0QeU2_1),.clk(gclk));
	jdff dff_B_mUoqfXpb6_2(.din(n1089),.dout(w_dff_B_mUoqfXpb6_2),.clk(gclk));
	jdff dff_B_I5ekQYDB4_2(.din(w_dff_B_mUoqfXpb6_2),.dout(w_dff_B_I5ekQYDB4_2),.clk(gclk));
	jdff dff_B_Vxpr2bKG5_2(.din(w_dff_B_I5ekQYDB4_2),.dout(w_dff_B_Vxpr2bKG5_2),.clk(gclk));
	jdff dff_B_AGojQlLr7_2(.din(w_dff_B_Vxpr2bKG5_2),.dout(w_dff_B_AGojQlLr7_2),.clk(gclk));
	jdff dff_B_6ZQeAD4R5_2(.din(w_dff_B_AGojQlLr7_2),.dout(w_dff_B_6ZQeAD4R5_2),.clk(gclk));
	jdff dff_B_svxZVkm66_2(.din(w_dff_B_6ZQeAD4R5_2),.dout(w_dff_B_svxZVkm66_2),.clk(gclk));
	jdff dff_B_MXek9y2s8_2(.din(w_dff_B_svxZVkm66_2),.dout(w_dff_B_MXek9y2s8_2),.clk(gclk));
	jdff dff_B_7iQWFiJG2_2(.din(w_dff_B_MXek9y2s8_2),.dout(w_dff_B_7iQWFiJG2_2),.clk(gclk));
	jdff dff_B_xRUPNnY77_2(.din(w_dff_B_7iQWFiJG2_2),.dout(w_dff_B_xRUPNnY77_2),.clk(gclk));
	jdff dff_B_RWVtGkIZ4_2(.din(w_dff_B_xRUPNnY77_2),.dout(w_dff_B_RWVtGkIZ4_2),.clk(gclk));
	jdff dff_B_xtJpvz2c0_2(.din(w_dff_B_RWVtGkIZ4_2),.dout(w_dff_B_xtJpvz2c0_2),.clk(gclk));
	jdff dff_B_VO0qJIZt6_2(.din(w_dff_B_xtJpvz2c0_2),.dout(w_dff_B_VO0qJIZt6_2),.clk(gclk));
	jdff dff_B_kv3EngaH2_2(.din(w_dff_B_VO0qJIZt6_2),.dout(w_dff_B_kv3EngaH2_2),.clk(gclk));
	jdff dff_B_47QfcKSa2_2(.din(w_dff_B_kv3EngaH2_2),.dout(w_dff_B_47QfcKSa2_2),.clk(gclk));
	jdff dff_B_Xp8eM6Dc5_2(.din(w_dff_B_47QfcKSa2_2),.dout(w_dff_B_Xp8eM6Dc5_2),.clk(gclk));
	jdff dff_B_vyo7kTGM4_2(.din(w_dff_B_Xp8eM6Dc5_2),.dout(w_dff_B_vyo7kTGM4_2),.clk(gclk));
	jdff dff_B_3YLVvh6J3_2(.din(w_dff_B_vyo7kTGM4_2),.dout(w_dff_B_3YLVvh6J3_2),.clk(gclk));
	jdff dff_B_W4qd8b791_2(.din(w_dff_B_3YLVvh6J3_2),.dout(w_dff_B_W4qd8b791_2),.clk(gclk));
	jdff dff_B_6X1GQTtL4_2(.din(n1119),.dout(w_dff_B_6X1GQTtL4_2),.clk(gclk));
	jdff dff_B_P3kYKh2x3_1(.din(n1090),.dout(w_dff_B_P3kYKh2x3_1),.clk(gclk));
	jdff dff_B_n9PjZANv1_2(.din(n991),.dout(w_dff_B_n9PjZANv1_2),.clk(gclk));
	jdff dff_B_BaxYGzmB6_2(.din(w_dff_B_n9PjZANv1_2),.dout(w_dff_B_BaxYGzmB6_2),.clk(gclk));
	jdff dff_B_Cltch9Dv1_2(.din(w_dff_B_BaxYGzmB6_2),.dout(w_dff_B_Cltch9Dv1_2),.clk(gclk));
	jdff dff_B_J7td25uE2_2(.din(w_dff_B_Cltch9Dv1_2),.dout(w_dff_B_J7td25uE2_2),.clk(gclk));
	jdff dff_B_W2wE3Ibc1_2(.din(w_dff_B_J7td25uE2_2),.dout(w_dff_B_W2wE3Ibc1_2),.clk(gclk));
	jdff dff_B_tS8MYGS40_2(.din(w_dff_B_W2wE3Ibc1_2),.dout(w_dff_B_tS8MYGS40_2),.clk(gclk));
	jdff dff_B_HrDbt5qB8_2(.din(w_dff_B_tS8MYGS40_2),.dout(w_dff_B_HrDbt5qB8_2),.clk(gclk));
	jdff dff_B_ICxvdQxH0_2(.din(w_dff_B_HrDbt5qB8_2),.dout(w_dff_B_ICxvdQxH0_2),.clk(gclk));
	jdff dff_B_W3Sw7jZn6_2(.din(w_dff_B_ICxvdQxH0_2),.dout(w_dff_B_W3Sw7jZn6_2),.clk(gclk));
	jdff dff_B_0GcYqEDU9_2(.din(w_dff_B_W3Sw7jZn6_2),.dout(w_dff_B_0GcYqEDU9_2),.clk(gclk));
	jdff dff_B_3IuKSbMU0_2(.din(w_dff_B_0GcYqEDU9_2),.dout(w_dff_B_3IuKSbMU0_2),.clk(gclk));
	jdff dff_B_Dqd4RCCR4_2(.din(w_dff_B_3IuKSbMU0_2),.dout(w_dff_B_Dqd4RCCR4_2),.clk(gclk));
	jdff dff_B_4dUU2XSZ9_2(.din(w_dff_B_Dqd4RCCR4_2),.dout(w_dff_B_4dUU2XSZ9_2),.clk(gclk));
	jdff dff_B_oeuxeKZW7_2(.din(w_dff_B_4dUU2XSZ9_2),.dout(w_dff_B_oeuxeKZW7_2),.clk(gclk));
	jdff dff_B_oOUT4ZHk3_2(.din(w_dff_B_oeuxeKZW7_2),.dout(w_dff_B_oOUT4ZHk3_2),.clk(gclk));
	jdff dff_B_BmViWpj58_2(.din(n1014),.dout(w_dff_B_BmViWpj58_2),.clk(gclk));
	jdff dff_B_SIoX6JBv3_1(.din(n992),.dout(w_dff_B_SIoX6JBv3_1),.clk(gclk));
	jdff dff_B_dzEnWlGx0_2(.din(n886),.dout(w_dff_B_dzEnWlGx0_2),.clk(gclk));
	jdff dff_B_Ry4equLn1_2(.din(w_dff_B_dzEnWlGx0_2),.dout(w_dff_B_Ry4equLn1_2),.clk(gclk));
	jdff dff_B_kt5DRlV32_2(.din(w_dff_B_Ry4equLn1_2),.dout(w_dff_B_kt5DRlV32_2),.clk(gclk));
	jdff dff_B_ZSQoWJbJ6_2(.din(w_dff_B_kt5DRlV32_2),.dout(w_dff_B_ZSQoWJbJ6_2),.clk(gclk));
	jdff dff_B_mVklfNNI6_2(.din(w_dff_B_ZSQoWJbJ6_2),.dout(w_dff_B_mVklfNNI6_2),.clk(gclk));
	jdff dff_B_XHI14um30_2(.din(w_dff_B_mVklfNNI6_2),.dout(w_dff_B_XHI14um30_2),.clk(gclk));
	jdff dff_B_qtgCMpEG1_2(.din(w_dff_B_XHI14um30_2),.dout(w_dff_B_qtgCMpEG1_2),.clk(gclk));
	jdff dff_B_3Ul1QpQD9_2(.din(w_dff_B_qtgCMpEG1_2),.dout(w_dff_B_3Ul1QpQD9_2),.clk(gclk));
	jdff dff_B_udoSRypK6_2(.din(w_dff_B_3Ul1QpQD9_2),.dout(w_dff_B_udoSRypK6_2),.clk(gclk));
	jdff dff_B_ufUGcuMS3_2(.din(w_dff_B_udoSRypK6_2),.dout(w_dff_B_ufUGcuMS3_2),.clk(gclk));
	jdff dff_B_d18ygHiN3_2(.din(w_dff_B_ufUGcuMS3_2),.dout(w_dff_B_d18ygHiN3_2),.clk(gclk));
	jdff dff_B_WSaq7kmt7_2(.din(w_dff_B_d18ygHiN3_2),.dout(w_dff_B_WSaq7kmt7_2),.clk(gclk));
	jdff dff_B_HJJXPDLJ1_2(.din(n909),.dout(w_dff_B_HJJXPDLJ1_2),.clk(gclk));
	jdff dff_B_EybfvUYZ7_1(.din(n887),.dout(w_dff_B_EybfvUYZ7_1),.clk(gclk));
	jdff dff_B_t2PhiEwp8_2(.din(n787),.dout(w_dff_B_t2PhiEwp8_2),.clk(gclk));
	jdff dff_B_HawM9VKV6_2(.din(w_dff_B_t2PhiEwp8_2),.dout(w_dff_B_HawM9VKV6_2),.clk(gclk));
	jdff dff_B_AcRAbhG65_2(.din(w_dff_B_HawM9VKV6_2),.dout(w_dff_B_AcRAbhG65_2),.clk(gclk));
	jdff dff_B_2vL1UFbj1_2(.din(w_dff_B_AcRAbhG65_2),.dout(w_dff_B_2vL1UFbj1_2),.clk(gclk));
	jdff dff_B_xB3fdIPI6_2(.din(w_dff_B_2vL1UFbj1_2),.dout(w_dff_B_xB3fdIPI6_2),.clk(gclk));
	jdff dff_B_ESApYGXA1_2(.din(w_dff_B_xB3fdIPI6_2),.dout(w_dff_B_ESApYGXA1_2),.clk(gclk));
	jdff dff_B_nSWEkW2E6_2(.din(w_dff_B_ESApYGXA1_2),.dout(w_dff_B_nSWEkW2E6_2),.clk(gclk));
	jdff dff_B_PgfyodEI6_2(.din(w_dff_B_nSWEkW2E6_2),.dout(w_dff_B_PgfyodEI6_2),.clk(gclk));
	jdff dff_B_khvspGQO6_2(.din(w_dff_B_PgfyodEI6_2),.dout(w_dff_B_khvspGQO6_2),.clk(gclk));
	jdff dff_B_9Ib3rFrG2_2(.din(n803),.dout(w_dff_B_9Ib3rFrG2_2),.clk(gclk));
	jdff dff_B_z0LSDmXY5_2(.din(w_dff_B_9Ib3rFrG2_2),.dout(w_dff_B_z0LSDmXY5_2),.clk(gclk));
	jdff dff_B_7ooSOI542_1(.din(n788),.dout(w_dff_B_7ooSOI542_1),.clk(gclk));
	jdff dff_B_p4ZKqOaR0_1(.din(w_dff_B_7ooSOI542_1),.dout(w_dff_B_p4ZKqOaR0_1),.clk(gclk));
	jdff dff_B_35davhdi4_1(.din(w_dff_B_p4ZKqOaR0_1),.dout(w_dff_B_35davhdi4_1),.clk(gclk));
	jdff dff_B_JTDIvzWL1_1(.din(w_dff_B_35davhdi4_1),.dout(w_dff_B_JTDIvzWL1_1),.clk(gclk));
	jdff dff_B_mhpKh3z56_1(.din(w_dff_B_JTDIvzWL1_1),.dout(w_dff_B_mhpKh3z56_1),.clk(gclk));
	jdff dff_B_AbMIWrjY2_1(.din(w_dff_B_mhpKh3z56_1),.dout(w_dff_B_AbMIWrjY2_1),.clk(gclk));
	jdff dff_B_lewCl6F46_0(.din(n703),.dout(w_dff_B_lewCl6F46_0),.clk(gclk));
	jdff dff_B_FN4EiElf2_0(.din(w_dff_B_lewCl6F46_0),.dout(w_dff_B_FN4EiElf2_0),.clk(gclk));
	jdff dff_A_LtKs6naQ4_0(.dout(w_n702_0[0]),.din(w_dff_A_LtKs6naQ4_0),.clk(gclk));
	jdff dff_A_QmNirHTN5_0(.dout(w_dff_A_LtKs6naQ4_0),.din(w_dff_A_QmNirHTN5_0),.clk(gclk));
	jdff dff_A_PuqeexTg5_0(.dout(w_dff_A_QmNirHTN5_0),.din(w_dff_A_PuqeexTg5_0),.clk(gclk));
	jdff dff_B_y9utSxa10_1(.din(n696),.dout(w_dff_B_y9utSxa10_1),.clk(gclk));
	jdff dff_A_NXNylrvi2_0(.dout(w_n607_0[0]),.din(w_dff_A_NXNylrvi2_0),.clk(gclk));
	jdff dff_A_L65x3gO94_1(.dout(w_n607_0[1]),.din(w_dff_A_L65x3gO94_1),.clk(gclk));
	jdff dff_A_M9IiwrW08_1(.dout(w_dff_A_L65x3gO94_1),.din(w_dff_A_M9IiwrW08_1),.clk(gclk));
	jdff dff_A_EGLeKxBN2_1(.dout(w_n694_0[1]),.din(w_dff_A_EGLeKxBN2_1),.clk(gclk));
	jdff dff_A_TJuwWHQb8_1(.dout(w_dff_A_EGLeKxBN2_1),.din(w_dff_A_TJuwWHQb8_1),.clk(gclk));
	jdff dff_A_1A2Pl0kz0_1(.dout(w_dff_A_TJuwWHQb8_1),.din(w_dff_A_1A2Pl0kz0_1),.clk(gclk));
	jdff dff_A_pp2KJSQw2_1(.dout(w_dff_A_1A2Pl0kz0_1),.din(w_dff_A_pp2KJSQw2_1),.clk(gclk));
	jdff dff_A_UVrgwKqi2_1(.dout(w_dff_A_pp2KJSQw2_1),.din(w_dff_A_UVrgwKqi2_1),.clk(gclk));
	jdff dff_A_pFIzj7hA7_1(.dout(w_dff_A_UVrgwKqi2_1),.din(w_dff_A_pFIzj7hA7_1),.clk(gclk));
	jdff dff_B_YhTOozlg0_1(.din(n1819),.dout(w_dff_B_YhTOozlg0_1),.clk(gclk));
	jdff dff_A_forErhb54_1(.dout(w_n1801_0[1]),.din(w_dff_A_forErhb54_1),.clk(gclk));
	jdff dff_B_M3dpZsFI7_1(.din(n1799),.dout(w_dff_B_M3dpZsFI7_1),.clk(gclk));
	jdff dff_B_0HaB0axa1_2(.din(n1770),.dout(w_dff_B_0HaB0axa1_2),.clk(gclk));
	jdff dff_B_7k4QvExD2_2(.din(w_dff_B_0HaB0axa1_2),.dout(w_dff_B_7k4QvExD2_2),.clk(gclk));
	jdff dff_B_ff95Fdir3_2(.din(w_dff_B_7k4QvExD2_2),.dout(w_dff_B_ff95Fdir3_2),.clk(gclk));
	jdff dff_B_TfongzZn7_2(.din(w_dff_B_ff95Fdir3_2),.dout(w_dff_B_TfongzZn7_2),.clk(gclk));
	jdff dff_B_wZEHvA7F2_2(.din(w_dff_B_TfongzZn7_2),.dout(w_dff_B_wZEHvA7F2_2),.clk(gclk));
	jdff dff_B_pXmYulmf2_2(.din(w_dff_B_wZEHvA7F2_2),.dout(w_dff_B_pXmYulmf2_2),.clk(gclk));
	jdff dff_B_hyAbOmRm7_2(.din(w_dff_B_pXmYulmf2_2),.dout(w_dff_B_hyAbOmRm7_2),.clk(gclk));
	jdff dff_B_NdWtZAad5_2(.din(w_dff_B_hyAbOmRm7_2),.dout(w_dff_B_NdWtZAad5_2),.clk(gclk));
	jdff dff_B_2EvYEiLO7_2(.din(w_dff_B_NdWtZAad5_2),.dout(w_dff_B_2EvYEiLO7_2),.clk(gclk));
	jdff dff_B_P6BeF5Ic8_2(.din(w_dff_B_2EvYEiLO7_2),.dout(w_dff_B_P6BeF5Ic8_2),.clk(gclk));
	jdff dff_B_3iyorYZv3_2(.din(w_dff_B_P6BeF5Ic8_2),.dout(w_dff_B_3iyorYZv3_2),.clk(gclk));
	jdff dff_B_ohECjMdP8_2(.din(w_dff_B_3iyorYZv3_2),.dout(w_dff_B_ohECjMdP8_2),.clk(gclk));
	jdff dff_B_vsmlhH618_2(.din(w_dff_B_ohECjMdP8_2),.dout(w_dff_B_vsmlhH618_2),.clk(gclk));
	jdff dff_B_mhVZrwmK5_2(.din(w_dff_B_vsmlhH618_2),.dout(w_dff_B_mhVZrwmK5_2),.clk(gclk));
	jdff dff_B_26FmZxsk4_2(.din(w_dff_B_mhVZrwmK5_2),.dout(w_dff_B_26FmZxsk4_2),.clk(gclk));
	jdff dff_B_FITgjqxD6_2(.din(w_dff_B_26FmZxsk4_2),.dout(w_dff_B_FITgjqxD6_2),.clk(gclk));
	jdff dff_B_SCjdpMpj2_2(.din(w_dff_B_FITgjqxD6_2),.dout(w_dff_B_SCjdpMpj2_2),.clk(gclk));
	jdff dff_B_saCfgQqm9_2(.din(w_dff_B_SCjdpMpj2_2),.dout(w_dff_B_saCfgQqm9_2),.clk(gclk));
	jdff dff_B_z8m9NxYF4_2(.din(w_dff_B_saCfgQqm9_2),.dout(w_dff_B_z8m9NxYF4_2),.clk(gclk));
	jdff dff_B_t7lFsx1r8_2(.din(w_dff_B_z8m9NxYF4_2),.dout(w_dff_B_t7lFsx1r8_2),.clk(gclk));
	jdff dff_B_WC7aDjPC7_2(.din(w_dff_B_t7lFsx1r8_2),.dout(w_dff_B_WC7aDjPC7_2),.clk(gclk));
	jdff dff_B_YDzMMs3k4_2(.din(w_dff_B_WC7aDjPC7_2),.dout(w_dff_B_YDzMMs3k4_2),.clk(gclk));
	jdff dff_B_snInNUvF6_2(.din(w_dff_B_YDzMMs3k4_2),.dout(w_dff_B_snInNUvF6_2),.clk(gclk));
	jdff dff_B_Eb2mfGpu2_2(.din(w_dff_B_snInNUvF6_2),.dout(w_dff_B_Eb2mfGpu2_2),.clk(gclk));
	jdff dff_B_C67XFGMj4_2(.din(w_dff_B_Eb2mfGpu2_2),.dout(w_dff_B_C67XFGMj4_2),.clk(gclk));
	jdff dff_B_Et0VyXD14_2(.din(w_dff_B_C67XFGMj4_2),.dout(w_dff_B_Et0VyXD14_2),.clk(gclk));
	jdff dff_B_ghyagT206_2(.din(w_dff_B_Et0VyXD14_2),.dout(w_dff_B_ghyagT206_2),.clk(gclk));
	jdff dff_B_1TcmJCxp3_2(.din(w_dff_B_ghyagT206_2),.dout(w_dff_B_1TcmJCxp3_2),.clk(gclk));
	jdff dff_B_2pibV6v52_2(.din(w_dff_B_1TcmJCxp3_2),.dout(w_dff_B_2pibV6v52_2),.clk(gclk));
	jdff dff_B_37YNWjfG8_2(.din(w_dff_B_2pibV6v52_2),.dout(w_dff_B_37YNWjfG8_2),.clk(gclk));
	jdff dff_B_P72XedN77_2(.din(w_dff_B_37YNWjfG8_2),.dout(w_dff_B_P72XedN77_2),.clk(gclk));
	jdff dff_B_xIP8GnzF5_2(.din(w_dff_B_P72XedN77_2),.dout(w_dff_B_xIP8GnzF5_2),.clk(gclk));
	jdff dff_B_U5rJyya81_2(.din(w_dff_B_xIP8GnzF5_2),.dout(w_dff_B_U5rJyya81_2),.clk(gclk));
	jdff dff_B_Cgri6rUs1_2(.din(w_dff_B_U5rJyya81_2),.dout(w_dff_B_Cgri6rUs1_2),.clk(gclk));
	jdff dff_B_V3iVCQRR9_2(.din(w_dff_B_Cgri6rUs1_2),.dout(w_dff_B_V3iVCQRR9_2),.clk(gclk));
	jdff dff_B_xWmgI4ER5_2(.din(w_dff_B_V3iVCQRR9_2),.dout(w_dff_B_xWmgI4ER5_2),.clk(gclk));
	jdff dff_B_PUcZxIoQ2_2(.din(w_dff_B_xWmgI4ER5_2),.dout(w_dff_B_PUcZxIoQ2_2),.clk(gclk));
	jdff dff_B_KtU4aUNN1_2(.din(w_dff_B_PUcZxIoQ2_2),.dout(w_dff_B_KtU4aUNN1_2),.clk(gclk));
	jdff dff_B_mZCFkYAs3_2(.din(w_dff_B_KtU4aUNN1_2),.dout(w_dff_B_mZCFkYAs3_2),.clk(gclk));
	jdff dff_B_YqQupxO30_2(.din(w_dff_B_mZCFkYAs3_2),.dout(w_dff_B_YqQupxO30_2),.clk(gclk));
	jdff dff_B_GgZharOd3_2(.din(w_dff_B_YqQupxO30_2),.dout(w_dff_B_GgZharOd3_2),.clk(gclk));
	jdff dff_B_Tl8NSNbd4_2(.din(w_dff_B_GgZharOd3_2),.dout(w_dff_B_Tl8NSNbd4_2),.clk(gclk));
	jdff dff_B_8l0m3WpH6_2(.din(w_dff_B_Tl8NSNbd4_2),.dout(w_dff_B_8l0m3WpH6_2),.clk(gclk));
	jdff dff_B_tSfQJftd3_2(.din(w_dff_B_8l0m3WpH6_2),.dout(w_dff_B_tSfQJftd3_2),.clk(gclk));
	jdff dff_B_X4Yd2b2h3_2(.din(w_dff_B_tSfQJftd3_2),.dout(w_dff_B_X4Yd2b2h3_2),.clk(gclk));
	jdff dff_B_JKWxCRqU5_2(.din(w_dff_B_X4Yd2b2h3_2),.dout(w_dff_B_JKWxCRqU5_2),.clk(gclk));
	jdff dff_B_weWzC20v2_2(.din(w_dff_B_JKWxCRqU5_2),.dout(w_dff_B_weWzC20v2_2),.clk(gclk));
	jdff dff_B_qpOnFZqU3_2(.din(w_dff_B_weWzC20v2_2),.dout(w_dff_B_qpOnFZqU3_2),.clk(gclk));
	jdff dff_B_zLPUFKln0_2(.din(w_dff_B_qpOnFZqU3_2),.dout(w_dff_B_zLPUFKln0_2),.clk(gclk));
	jdff dff_B_frcMyTb66_2(.din(w_dff_B_zLPUFKln0_2),.dout(w_dff_B_frcMyTb66_2),.clk(gclk));
	jdff dff_B_XZ7ZVWWB7_2(.din(w_dff_B_frcMyTb66_2),.dout(w_dff_B_XZ7ZVWWB7_2),.clk(gclk));
	jdff dff_B_8MOyUki03_2(.din(w_dff_B_XZ7ZVWWB7_2),.dout(w_dff_B_8MOyUki03_2),.clk(gclk));
	jdff dff_B_ZmKqx6aG2_2(.din(w_dff_B_8MOyUki03_2),.dout(w_dff_B_ZmKqx6aG2_2),.clk(gclk));
	jdff dff_B_LyBfnB659_2(.din(n1773),.dout(w_dff_B_LyBfnB659_2),.clk(gclk));
	jdff dff_B_DfFTOkR05_1(.din(n1771),.dout(w_dff_B_DfFTOkR05_1),.clk(gclk));
	jdff dff_B_YRZNjY0L5_2(.din(n1735),.dout(w_dff_B_YRZNjY0L5_2),.clk(gclk));
	jdff dff_B_gGnvlyNI1_2(.din(w_dff_B_YRZNjY0L5_2),.dout(w_dff_B_gGnvlyNI1_2),.clk(gclk));
	jdff dff_B_9RO4XDfu8_2(.din(w_dff_B_gGnvlyNI1_2),.dout(w_dff_B_9RO4XDfu8_2),.clk(gclk));
	jdff dff_B_XYGfNuor9_2(.din(w_dff_B_9RO4XDfu8_2),.dout(w_dff_B_XYGfNuor9_2),.clk(gclk));
	jdff dff_B_89Mem6RN5_2(.din(w_dff_B_XYGfNuor9_2),.dout(w_dff_B_89Mem6RN5_2),.clk(gclk));
	jdff dff_B_vi1Xy4W39_2(.din(w_dff_B_89Mem6RN5_2),.dout(w_dff_B_vi1Xy4W39_2),.clk(gclk));
	jdff dff_B_YgBCan3K2_2(.din(w_dff_B_vi1Xy4W39_2),.dout(w_dff_B_YgBCan3K2_2),.clk(gclk));
	jdff dff_B_9BusRFDI9_2(.din(w_dff_B_YgBCan3K2_2),.dout(w_dff_B_9BusRFDI9_2),.clk(gclk));
	jdff dff_B_0lHoUBJZ3_2(.din(w_dff_B_9BusRFDI9_2),.dout(w_dff_B_0lHoUBJZ3_2),.clk(gclk));
	jdff dff_B_JlD1X6Zy2_2(.din(w_dff_B_0lHoUBJZ3_2),.dout(w_dff_B_JlD1X6Zy2_2),.clk(gclk));
	jdff dff_B_MgqiZD7h9_2(.din(w_dff_B_JlD1X6Zy2_2),.dout(w_dff_B_MgqiZD7h9_2),.clk(gclk));
	jdff dff_B_CIluDLVX6_2(.din(w_dff_B_MgqiZD7h9_2),.dout(w_dff_B_CIluDLVX6_2),.clk(gclk));
	jdff dff_B_SFCQgHe50_2(.din(w_dff_B_CIluDLVX6_2),.dout(w_dff_B_SFCQgHe50_2),.clk(gclk));
	jdff dff_B_YJjqGf9e7_2(.din(w_dff_B_SFCQgHe50_2),.dout(w_dff_B_YJjqGf9e7_2),.clk(gclk));
	jdff dff_B_k43PoL7w5_2(.din(w_dff_B_YJjqGf9e7_2),.dout(w_dff_B_k43PoL7w5_2),.clk(gclk));
	jdff dff_B_3QikwAPS3_2(.din(w_dff_B_k43PoL7w5_2),.dout(w_dff_B_3QikwAPS3_2),.clk(gclk));
	jdff dff_B_Dxm82Scn5_2(.din(w_dff_B_3QikwAPS3_2),.dout(w_dff_B_Dxm82Scn5_2),.clk(gclk));
	jdff dff_B_Tne9fqnL2_2(.din(w_dff_B_Dxm82Scn5_2),.dout(w_dff_B_Tne9fqnL2_2),.clk(gclk));
	jdff dff_B_rZctT1pP5_2(.din(w_dff_B_Tne9fqnL2_2),.dout(w_dff_B_rZctT1pP5_2),.clk(gclk));
	jdff dff_B_40kpmGss3_2(.din(w_dff_B_rZctT1pP5_2),.dout(w_dff_B_40kpmGss3_2),.clk(gclk));
	jdff dff_B_Uer9rEWK1_2(.din(w_dff_B_40kpmGss3_2),.dout(w_dff_B_Uer9rEWK1_2),.clk(gclk));
	jdff dff_B_765oAwsF8_2(.din(w_dff_B_Uer9rEWK1_2),.dout(w_dff_B_765oAwsF8_2),.clk(gclk));
	jdff dff_B_1R5ZorMF6_2(.din(w_dff_B_765oAwsF8_2),.dout(w_dff_B_1R5ZorMF6_2),.clk(gclk));
	jdff dff_B_qkNxMDal8_2(.din(w_dff_B_1R5ZorMF6_2),.dout(w_dff_B_qkNxMDal8_2),.clk(gclk));
	jdff dff_B_HA4bT9nV5_2(.din(w_dff_B_qkNxMDal8_2),.dout(w_dff_B_HA4bT9nV5_2),.clk(gclk));
	jdff dff_B_oiooNBCM8_2(.din(w_dff_B_HA4bT9nV5_2),.dout(w_dff_B_oiooNBCM8_2),.clk(gclk));
	jdff dff_B_J8sTyzIM5_2(.din(w_dff_B_oiooNBCM8_2),.dout(w_dff_B_J8sTyzIM5_2),.clk(gclk));
	jdff dff_B_KMKTM12T8_2(.din(w_dff_B_J8sTyzIM5_2),.dout(w_dff_B_KMKTM12T8_2),.clk(gclk));
	jdff dff_B_zIA0RoIn2_2(.din(w_dff_B_KMKTM12T8_2),.dout(w_dff_B_zIA0RoIn2_2),.clk(gclk));
	jdff dff_B_C1AJAiKq3_2(.din(w_dff_B_zIA0RoIn2_2),.dout(w_dff_B_C1AJAiKq3_2),.clk(gclk));
	jdff dff_B_5fr6FxiB9_2(.din(w_dff_B_C1AJAiKq3_2),.dout(w_dff_B_5fr6FxiB9_2),.clk(gclk));
	jdff dff_B_U0TSpj3E9_2(.din(w_dff_B_5fr6FxiB9_2),.dout(w_dff_B_U0TSpj3E9_2),.clk(gclk));
	jdff dff_B_n5lHouWi7_2(.din(w_dff_B_U0TSpj3E9_2),.dout(w_dff_B_n5lHouWi7_2),.clk(gclk));
	jdff dff_B_p4jnIHe76_2(.din(w_dff_B_n5lHouWi7_2),.dout(w_dff_B_p4jnIHe76_2),.clk(gclk));
	jdff dff_B_1Jf62CBt7_2(.din(w_dff_B_p4jnIHe76_2),.dout(w_dff_B_1Jf62CBt7_2),.clk(gclk));
	jdff dff_B_Bq6k7Bc37_2(.din(w_dff_B_1Jf62CBt7_2),.dout(w_dff_B_Bq6k7Bc37_2),.clk(gclk));
	jdff dff_B_DiRQqmv01_2(.din(w_dff_B_Bq6k7Bc37_2),.dout(w_dff_B_DiRQqmv01_2),.clk(gclk));
	jdff dff_B_H2XFhAhq2_2(.din(w_dff_B_DiRQqmv01_2),.dout(w_dff_B_H2XFhAhq2_2),.clk(gclk));
	jdff dff_B_hKB2wtra9_2(.din(w_dff_B_H2XFhAhq2_2),.dout(w_dff_B_hKB2wtra9_2),.clk(gclk));
	jdff dff_B_mfFIpu5e7_2(.din(w_dff_B_hKB2wtra9_2),.dout(w_dff_B_mfFIpu5e7_2),.clk(gclk));
	jdff dff_B_Sd5nOAgD9_2(.din(w_dff_B_mfFIpu5e7_2),.dout(w_dff_B_Sd5nOAgD9_2),.clk(gclk));
	jdff dff_B_olUqor7E8_2(.din(w_dff_B_Sd5nOAgD9_2),.dout(w_dff_B_olUqor7E8_2),.clk(gclk));
	jdff dff_B_ESaHf6bM1_2(.din(w_dff_B_olUqor7E8_2),.dout(w_dff_B_ESaHf6bM1_2),.clk(gclk));
	jdff dff_B_EXBnntxx7_2(.din(w_dff_B_ESaHf6bM1_2),.dout(w_dff_B_EXBnntxx7_2),.clk(gclk));
	jdff dff_B_WcLJcDnf9_2(.din(w_dff_B_EXBnntxx7_2),.dout(w_dff_B_WcLJcDnf9_2),.clk(gclk));
	jdff dff_B_sfl1UaQe2_2(.din(w_dff_B_WcLJcDnf9_2),.dout(w_dff_B_sfl1UaQe2_2),.clk(gclk));
	jdff dff_B_N6P56TQY2_2(.din(w_dff_B_sfl1UaQe2_2),.dout(w_dff_B_N6P56TQY2_2),.clk(gclk));
	jdff dff_B_3c4LTtp89_2(.din(w_dff_B_N6P56TQY2_2),.dout(w_dff_B_3c4LTtp89_2),.clk(gclk));
	jdff dff_B_jlXX2w2d4_2(.din(w_dff_B_3c4LTtp89_2),.dout(w_dff_B_jlXX2w2d4_2),.clk(gclk));
	jdff dff_B_4bnrSVb15_2(.din(n1738),.dout(w_dff_B_4bnrSVb15_2),.clk(gclk));
	jdff dff_B_th8nxmQb1_1(.din(n1736),.dout(w_dff_B_th8nxmQb1_1),.clk(gclk));
	jdff dff_B_spksI4KI0_2(.din(n1694),.dout(w_dff_B_spksI4KI0_2),.clk(gclk));
	jdff dff_B_gHoaugaJ5_2(.din(w_dff_B_spksI4KI0_2),.dout(w_dff_B_gHoaugaJ5_2),.clk(gclk));
	jdff dff_B_viVHGa2t2_2(.din(w_dff_B_gHoaugaJ5_2),.dout(w_dff_B_viVHGa2t2_2),.clk(gclk));
	jdff dff_B_UdS3I12J1_2(.din(w_dff_B_viVHGa2t2_2),.dout(w_dff_B_UdS3I12J1_2),.clk(gclk));
	jdff dff_B_AOLr9xT47_2(.din(w_dff_B_UdS3I12J1_2),.dout(w_dff_B_AOLr9xT47_2),.clk(gclk));
	jdff dff_B_9NBuqUrL2_2(.din(w_dff_B_AOLr9xT47_2),.dout(w_dff_B_9NBuqUrL2_2),.clk(gclk));
	jdff dff_B_cnniJind8_2(.din(w_dff_B_9NBuqUrL2_2),.dout(w_dff_B_cnniJind8_2),.clk(gclk));
	jdff dff_B_Plx1KvFc4_2(.din(w_dff_B_cnniJind8_2),.dout(w_dff_B_Plx1KvFc4_2),.clk(gclk));
	jdff dff_B_yCEQ6V7U7_2(.din(w_dff_B_Plx1KvFc4_2),.dout(w_dff_B_yCEQ6V7U7_2),.clk(gclk));
	jdff dff_B_aKePuP7k2_2(.din(w_dff_B_yCEQ6V7U7_2),.dout(w_dff_B_aKePuP7k2_2),.clk(gclk));
	jdff dff_B_MkIVpLcQ4_2(.din(w_dff_B_aKePuP7k2_2),.dout(w_dff_B_MkIVpLcQ4_2),.clk(gclk));
	jdff dff_B_kDx8BLnU9_2(.din(w_dff_B_MkIVpLcQ4_2),.dout(w_dff_B_kDx8BLnU9_2),.clk(gclk));
	jdff dff_B_6UEBJIhl9_2(.din(w_dff_B_kDx8BLnU9_2),.dout(w_dff_B_6UEBJIhl9_2),.clk(gclk));
	jdff dff_B_UtZSgd8F0_2(.din(w_dff_B_6UEBJIhl9_2),.dout(w_dff_B_UtZSgd8F0_2),.clk(gclk));
	jdff dff_B_OQMvVDlt5_2(.din(w_dff_B_UtZSgd8F0_2),.dout(w_dff_B_OQMvVDlt5_2),.clk(gclk));
	jdff dff_B_8YfpEEqJ8_2(.din(w_dff_B_OQMvVDlt5_2),.dout(w_dff_B_8YfpEEqJ8_2),.clk(gclk));
	jdff dff_B_ga1HpFPy4_2(.din(w_dff_B_8YfpEEqJ8_2),.dout(w_dff_B_ga1HpFPy4_2),.clk(gclk));
	jdff dff_B_YsuQS3bt7_2(.din(w_dff_B_ga1HpFPy4_2),.dout(w_dff_B_YsuQS3bt7_2),.clk(gclk));
	jdff dff_B_Kgw5zafA2_2(.din(w_dff_B_YsuQS3bt7_2),.dout(w_dff_B_Kgw5zafA2_2),.clk(gclk));
	jdff dff_B_mxnlupeJ6_2(.din(w_dff_B_Kgw5zafA2_2),.dout(w_dff_B_mxnlupeJ6_2),.clk(gclk));
	jdff dff_B_XCeZ6X786_2(.din(w_dff_B_mxnlupeJ6_2),.dout(w_dff_B_XCeZ6X786_2),.clk(gclk));
	jdff dff_B_U7h8D77U3_2(.din(w_dff_B_XCeZ6X786_2),.dout(w_dff_B_U7h8D77U3_2),.clk(gclk));
	jdff dff_B_zGSSVDbV3_2(.din(w_dff_B_U7h8D77U3_2),.dout(w_dff_B_zGSSVDbV3_2),.clk(gclk));
	jdff dff_B_4dFxaZsZ6_2(.din(w_dff_B_zGSSVDbV3_2),.dout(w_dff_B_4dFxaZsZ6_2),.clk(gclk));
	jdff dff_B_dW2WJBGK4_2(.din(w_dff_B_4dFxaZsZ6_2),.dout(w_dff_B_dW2WJBGK4_2),.clk(gclk));
	jdff dff_B_eBkrm5Sx6_2(.din(w_dff_B_dW2WJBGK4_2),.dout(w_dff_B_eBkrm5Sx6_2),.clk(gclk));
	jdff dff_B_IbEw2Xca7_2(.din(w_dff_B_eBkrm5Sx6_2),.dout(w_dff_B_IbEw2Xca7_2),.clk(gclk));
	jdff dff_B_5MXoy1wm3_2(.din(w_dff_B_IbEw2Xca7_2),.dout(w_dff_B_5MXoy1wm3_2),.clk(gclk));
	jdff dff_B_UWiHhwvR6_2(.din(w_dff_B_5MXoy1wm3_2),.dout(w_dff_B_UWiHhwvR6_2),.clk(gclk));
	jdff dff_B_vN9s1hvP2_2(.din(w_dff_B_UWiHhwvR6_2),.dout(w_dff_B_vN9s1hvP2_2),.clk(gclk));
	jdff dff_B_Ah8tPILE5_2(.din(w_dff_B_vN9s1hvP2_2),.dout(w_dff_B_Ah8tPILE5_2),.clk(gclk));
	jdff dff_B_Sml7fttA9_2(.din(w_dff_B_Ah8tPILE5_2),.dout(w_dff_B_Sml7fttA9_2),.clk(gclk));
	jdff dff_B_3n7fR1TM1_2(.din(w_dff_B_Sml7fttA9_2),.dout(w_dff_B_3n7fR1TM1_2),.clk(gclk));
	jdff dff_B_tCttBEOm2_2(.din(w_dff_B_3n7fR1TM1_2),.dout(w_dff_B_tCttBEOm2_2),.clk(gclk));
	jdff dff_B_7lD3d9d15_2(.din(w_dff_B_tCttBEOm2_2),.dout(w_dff_B_7lD3d9d15_2),.clk(gclk));
	jdff dff_B_UAbuuPvg5_2(.din(w_dff_B_7lD3d9d15_2),.dout(w_dff_B_UAbuuPvg5_2),.clk(gclk));
	jdff dff_B_5ePkDAKo5_2(.din(w_dff_B_UAbuuPvg5_2),.dout(w_dff_B_5ePkDAKo5_2),.clk(gclk));
	jdff dff_B_7UIwb4sd0_2(.din(w_dff_B_5ePkDAKo5_2),.dout(w_dff_B_7UIwb4sd0_2),.clk(gclk));
	jdff dff_B_rZ6uSX1I1_2(.din(w_dff_B_7UIwb4sd0_2),.dout(w_dff_B_rZ6uSX1I1_2),.clk(gclk));
	jdff dff_B_bI1QfeL17_2(.din(w_dff_B_rZ6uSX1I1_2),.dout(w_dff_B_bI1QfeL17_2),.clk(gclk));
	jdff dff_B_QfTPBrKg4_2(.din(w_dff_B_bI1QfeL17_2),.dout(w_dff_B_QfTPBrKg4_2),.clk(gclk));
	jdff dff_B_lxgyNDby2_2(.din(w_dff_B_QfTPBrKg4_2),.dout(w_dff_B_lxgyNDby2_2),.clk(gclk));
	jdff dff_B_u1V6BJSX0_2(.din(w_dff_B_lxgyNDby2_2),.dout(w_dff_B_u1V6BJSX0_2),.clk(gclk));
	jdff dff_B_mldm1BE82_2(.din(w_dff_B_u1V6BJSX0_2),.dout(w_dff_B_mldm1BE82_2),.clk(gclk));
	jdff dff_B_Eg9FkntX4_2(.din(w_dff_B_mldm1BE82_2),.dout(w_dff_B_Eg9FkntX4_2),.clk(gclk));
	jdff dff_B_j8LajU4o8_2(.din(n1697),.dout(w_dff_B_j8LajU4o8_2),.clk(gclk));
	jdff dff_B_lFIuXwu42_1(.din(n1695),.dout(w_dff_B_lFIuXwu42_1),.clk(gclk));
	jdff dff_B_Qs3ojZcJ0_2(.din(n1643),.dout(w_dff_B_Qs3ojZcJ0_2),.clk(gclk));
	jdff dff_B_uIbXlQDa0_2(.din(w_dff_B_Qs3ojZcJ0_2),.dout(w_dff_B_uIbXlQDa0_2),.clk(gclk));
	jdff dff_B_dcBuCuRl6_2(.din(w_dff_B_uIbXlQDa0_2),.dout(w_dff_B_dcBuCuRl6_2),.clk(gclk));
	jdff dff_B_gsMoO4Be2_2(.din(w_dff_B_dcBuCuRl6_2),.dout(w_dff_B_gsMoO4Be2_2),.clk(gclk));
	jdff dff_B_PN9urS541_2(.din(w_dff_B_gsMoO4Be2_2),.dout(w_dff_B_PN9urS541_2),.clk(gclk));
	jdff dff_B_RXGdaVUM3_2(.din(w_dff_B_PN9urS541_2),.dout(w_dff_B_RXGdaVUM3_2),.clk(gclk));
	jdff dff_B_hFY1IdO71_2(.din(w_dff_B_RXGdaVUM3_2),.dout(w_dff_B_hFY1IdO71_2),.clk(gclk));
	jdff dff_B_RhxEi5HN8_2(.din(w_dff_B_hFY1IdO71_2),.dout(w_dff_B_RhxEi5HN8_2),.clk(gclk));
	jdff dff_B_Ml4x5f5j1_2(.din(w_dff_B_RhxEi5HN8_2),.dout(w_dff_B_Ml4x5f5j1_2),.clk(gclk));
	jdff dff_B_LV5TmCsu1_2(.din(w_dff_B_Ml4x5f5j1_2),.dout(w_dff_B_LV5TmCsu1_2),.clk(gclk));
	jdff dff_B_Zn7zUcSl6_2(.din(w_dff_B_LV5TmCsu1_2),.dout(w_dff_B_Zn7zUcSl6_2),.clk(gclk));
	jdff dff_B_Bw97XVjD4_2(.din(w_dff_B_Zn7zUcSl6_2),.dout(w_dff_B_Bw97XVjD4_2),.clk(gclk));
	jdff dff_B_PNa2N3v14_2(.din(w_dff_B_Bw97XVjD4_2),.dout(w_dff_B_PNa2N3v14_2),.clk(gclk));
	jdff dff_B_rPT91Zz68_2(.din(w_dff_B_PNa2N3v14_2),.dout(w_dff_B_rPT91Zz68_2),.clk(gclk));
	jdff dff_B_6ESbXcw15_2(.din(w_dff_B_rPT91Zz68_2),.dout(w_dff_B_6ESbXcw15_2),.clk(gclk));
	jdff dff_B_lM21z01S2_2(.din(w_dff_B_6ESbXcw15_2),.dout(w_dff_B_lM21z01S2_2),.clk(gclk));
	jdff dff_B_6VHY6elh1_2(.din(w_dff_B_lM21z01S2_2),.dout(w_dff_B_6VHY6elh1_2),.clk(gclk));
	jdff dff_B_5QK2eMPN4_2(.din(w_dff_B_6VHY6elh1_2),.dout(w_dff_B_5QK2eMPN4_2),.clk(gclk));
	jdff dff_B_AkX6FeFy1_2(.din(w_dff_B_5QK2eMPN4_2),.dout(w_dff_B_AkX6FeFy1_2),.clk(gclk));
	jdff dff_B_OmAPtIcb8_2(.din(w_dff_B_AkX6FeFy1_2),.dout(w_dff_B_OmAPtIcb8_2),.clk(gclk));
	jdff dff_B_3mOYujGQ7_2(.din(w_dff_B_OmAPtIcb8_2),.dout(w_dff_B_3mOYujGQ7_2),.clk(gclk));
	jdff dff_B_0oO0W1rO1_2(.din(w_dff_B_3mOYujGQ7_2),.dout(w_dff_B_0oO0W1rO1_2),.clk(gclk));
	jdff dff_B_4804Unir7_2(.din(w_dff_B_0oO0W1rO1_2),.dout(w_dff_B_4804Unir7_2),.clk(gclk));
	jdff dff_B_QWZeIdVw4_2(.din(w_dff_B_4804Unir7_2),.dout(w_dff_B_QWZeIdVw4_2),.clk(gclk));
	jdff dff_B_Zb6eP5zx5_2(.din(w_dff_B_QWZeIdVw4_2),.dout(w_dff_B_Zb6eP5zx5_2),.clk(gclk));
	jdff dff_B_Mbfv9tEX3_2(.din(w_dff_B_Zb6eP5zx5_2),.dout(w_dff_B_Mbfv9tEX3_2),.clk(gclk));
	jdff dff_B_y14YbYYC8_2(.din(w_dff_B_Mbfv9tEX3_2),.dout(w_dff_B_y14YbYYC8_2),.clk(gclk));
	jdff dff_B_MEB5eMOl8_2(.din(w_dff_B_y14YbYYC8_2),.dout(w_dff_B_MEB5eMOl8_2),.clk(gclk));
	jdff dff_B_UyIA1UxH8_2(.din(w_dff_B_MEB5eMOl8_2),.dout(w_dff_B_UyIA1UxH8_2),.clk(gclk));
	jdff dff_B_RlgI2S1y2_2(.din(w_dff_B_UyIA1UxH8_2),.dout(w_dff_B_RlgI2S1y2_2),.clk(gclk));
	jdff dff_B_gL60ooUd5_2(.din(w_dff_B_RlgI2S1y2_2),.dout(w_dff_B_gL60ooUd5_2),.clk(gclk));
	jdff dff_B_LYVrfjo41_2(.din(w_dff_B_gL60ooUd5_2),.dout(w_dff_B_LYVrfjo41_2),.clk(gclk));
	jdff dff_B_ZbhGg4gX2_2(.din(w_dff_B_LYVrfjo41_2),.dout(w_dff_B_ZbhGg4gX2_2),.clk(gclk));
	jdff dff_B_td786v915_2(.din(w_dff_B_ZbhGg4gX2_2),.dout(w_dff_B_td786v915_2),.clk(gclk));
	jdff dff_B_iMPfI7pk1_2(.din(w_dff_B_td786v915_2),.dout(w_dff_B_iMPfI7pk1_2),.clk(gclk));
	jdff dff_B_ZQWJoX5c6_2(.din(w_dff_B_iMPfI7pk1_2),.dout(w_dff_B_ZQWJoX5c6_2),.clk(gclk));
	jdff dff_B_VD1PKCFu3_2(.din(w_dff_B_ZQWJoX5c6_2),.dout(w_dff_B_VD1PKCFu3_2),.clk(gclk));
	jdff dff_B_WSo1ZvR09_2(.din(w_dff_B_VD1PKCFu3_2),.dout(w_dff_B_WSo1ZvR09_2),.clk(gclk));
	jdff dff_B_B3u1pvnC9_2(.din(w_dff_B_WSo1ZvR09_2),.dout(w_dff_B_B3u1pvnC9_2),.clk(gclk));
	jdff dff_B_oB3QjWB10_2(.din(w_dff_B_B3u1pvnC9_2),.dout(w_dff_B_oB3QjWB10_2),.clk(gclk));
	jdff dff_B_pLG9O1LA0_2(.din(w_dff_B_oB3QjWB10_2),.dout(w_dff_B_pLG9O1LA0_2),.clk(gclk));
	jdff dff_B_sWdREgKP8_2(.din(n1646),.dout(w_dff_B_sWdREgKP8_2),.clk(gclk));
	jdff dff_B_xk3vPnoh0_1(.din(n1644),.dout(w_dff_B_xk3vPnoh0_1),.clk(gclk));
	jdff dff_B_uxfWC7P78_2(.din(n1586),.dout(w_dff_B_uxfWC7P78_2),.clk(gclk));
	jdff dff_B_GJib9xOZ1_2(.din(w_dff_B_uxfWC7P78_2),.dout(w_dff_B_GJib9xOZ1_2),.clk(gclk));
	jdff dff_B_3ez7Cg612_2(.din(w_dff_B_GJib9xOZ1_2),.dout(w_dff_B_3ez7Cg612_2),.clk(gclk));
	jdff dff_B_LG7u3Kno1_2(.din(w_dff_B_3ez7Cg612_2),.dout(w_dff_B_LG7u3Kno1_2),.clk(gclk));
	jdff dff_B_v3wBOw1y6_2(.din(w_dff_B_LG7u3Kno1_2),.dout(w_dff_B_v3wBOw1y6_2),.clk(gclk));
	jdff dff_B_6e14Ipz25_2(.din(w_dff_B_v3wBOw1y6_2),.dout(w_dff_B_6e14Ipz25_2),.clk(gclk));
	jdff dff_B_tpddZU6i5_2(.din(w_dff_B_6e14Ipz25_2),.dout(w_dff_B_tpddZU6i5_2),.clk(gclk));
	jdff dff_B_3aX0VfXz2_2(.din(w_dff_B_tpddZU6i5_2),.dout(w_dff_B_3aX0VfXz2_2),.clk(gclk));
	jdff dff_B_kXJGuqJH4_2(.din(w_dff_B_3aX0VfXz2_2),.dout(w_dff_B_kXJGuqJH4_2),.clk(gclk));
	jdff dff_B_gHmvmxyR7_2(.din(w_dff_B_kXJGuqJH4_2),.dout(w_dff_B_gHmvmxyR7_2),.clk(gclk));
	jdff dff_B_7JAUW5HU3_2(.din(w_dff_B_gHmvmxyR7_2),.dout(w_dff_B_7JAUW5HU3_2),.clk(gclk));
	jdff dff_B_nlt359wa6_2(.din(w_dff_B_7JAUW5HU3_2),.dout(w_dff_B_nlt359wa6_2),.clk(gclk));
	jdff dff_B_Vrl86BMW7_2(.din(w_dff_B_nlt359wa6_2),.dout(w_dff_B_Vrl86BMW7_2),.clk(gclk));
	jdff dff_B_NKtHwobk8_2(.din(w_dff_B_Vrl86BMW7_2),.dout(w_dff_B_NKtHwobk8_2),.clk(gclk));
	jdff dff_B_bUSfSCpp7_2(.din(w_dff_B_NKtHwobk8_2),.dout(w_dff_B_bUSfSCpp7_2),.clk(gclk));
	jdff dff_B_97LlHUBV3_2(.din(w_dff_B_bUSfSCpp7_2),.dout(w_dff_B_97LlHUBV3_2),.clk(gclk));
	jdff dff_B_rcHDfZcH4_2(.din(w_dff_B_97LlHUBV3_2),.dout(w_dff_B_rcHDfZcH4_2),.clk(gclk));
	jdff dff_B_8hUEyB7o2_2(.din(w_dff_B_rcHDfZcH4_2),.dout(w_dff_B_8hUEyB7o2_2),.clk(gclk));
	jdff dff_B_0GY5Vt3I3_2(.din(w_dff_B_8hUEyB7o2_2),.dout(w_dff_B_0GY5Vt3I3_2),.clk(gclk));
	jdff dff_B_Zo7e0ClY7_2(.din(w_dff_B_0GY5Vt3I3_2),.dout(w_dff_B_Zo7e0ClY7_2),.clk(gclk));
	jdff dff_B_x4TZboyO8_2(.din(w_dff_B_Zo7e0ClY7_2),.dout(w_dff_B_x4TZboyO8_2),.clk(gclk));
	jdff dff_B_mEol29mC6_2(.din(w_dff_B_x4TZboyO8_2),.dout(w_dff_B_mEol29mC6_2),.clk(gclk));
	jdff dff_B_sP7jbFzi9_2(.din(w_dff_B_mEol29mC6_2),.dout(w_dff_B_sP7jbFzi9_2),.clk(gclk));
	jdff dff_B_jdlrES7f4_2(.din(w_dff_B_sP7jbFzi9_2),.dout(w_dff_B_jdlrES7f4_2),.clk(gclk));
	jdff dff_B_FVRPTocC9_2(.din(w_dff_B_jdlrES7f4_2),.dout(w_dff_B_FVRPTocC9_2),.clk(gclk));
	jdff dff_B_A7NlLIC69_2(.din(w_dff_B_FVRPTocC9_2),.dout(w_dff_B_A7NlLIC69_2),.clk(gclk));
	jdff dff_B_DlUjNFQq2_2(.din(w_dff_B_A7NlLIC69_2),.dout(w_dff_B_DlUjNFQq2_2),.clk(gclk));
	jdff dff_B_uTBzcYKo6_2(.din(w_dff_B_DlUjNFQq2_2),.dout(w_dff_B_uTBzcYKo6_2),.clk(gclk));
	jdff dff_B_7GTTzrjg5_2(.din(w_dff_B_uTBzcYKo6_2),.dout(w_dff_B_7GTTzrjg5_2),.clk(gclk));
	jdff dff_B_Hm5u2qJ15_2(.din(w_dff_B_7GTTzrjg5_2),.dout(w_dff_B_Hm5u2qJ15_2),.clk(gclk));
	jdff dff_B_RrjHD4372_2(.din(w_dff_B_Hm5u2qJ15_2),.dout(w_dff_B_RrjHD4372_2),.clk(gclk));
	jdff dff_B_f7wSfMtQ4_2(.din(w_dff_B_RrjHD4372_2),.dout(w_dff_B_f7wSfMtQ4_2),.clk(gclk));
	jdff dff_B_s6n4OxjG2_2(.din(w_dff_B_f7wSfMtQ4_2),.dout(w_dff_B_s6n4OxjG2_2),.clk(gclk));
	jdff dff_B_AG23YI9i6_2(.din(w_dff_B_s6n4OxjG2_2),.dout(w_dff_B_AG23YI9i6_2),.clk(gclk));
	jdff dff_B_HjmzoJX10_2(.din(w_dff_B_AG23YI9i6_2),.dout(w_dff_B_HjmzoJX10_2),.clk(gclk));
	jdff dff_B_0QPLeRFa5_2(.din(w_dff_B_HjmzoJX10_2),.dout(w_dff_B_0QPLeRFa5_2),.clk(gclk));
	jdff dff_B_OncjjOTl6_2(.din(w_dff_B_0QPLeRFa5_2),.dout(w_dff_B_OncjjOTl6_2),.clk(gclk));
	jdff dff_B_nlDQTvOA9_2(.din(n1589),.dout(w_dff_B_nlDQTvOA9_2),.clk(gclk));
	jdff dff_B_h6vcaayM6_1(.din(n1587),.dout(w_dff_B_h6vcaayM6_1),.clk(gclk));
	jdff dff_B_LN1KLsKG0_2(.din(n1522),.dout(w_dff_B_LN1KLsKG0_2),.clk(gclk));
	jdff dff_B_EKv3aaBO9_2(.din(w_dff_B_LN1KLsKG0_2),.dout(w_dff_B_EKv3aaBO9_2),.clk(gclk));
	jdff dff_B_ih1LFmet0_2(.din(w_dff_B_EKv3aaBO9_2),.dout(w_dff_B_ih1LFmet0_2),.clk(gclk));
	jdff dff_B_TE6bvH520_2(.din(w_dff_B_ih1LFmet0_2),.dout(w_dff_B_TE6bvH520_2),.clk(gclk));
	jdff dff_B_jbA2pDBE3_2(.din(w_dff_B_TE6bvH520_2),.dout(w_dff_B_jbA2pDBE3_2),.clk(gclk));
	jdff dff_B_6GS2D6WL2_2(.din(w_dff_B_jbA2pDBE3_2),.dout(w_dff_B_6GS2D6WL2_2),.clk(gclk));
	jdff dff_B_bahWkaCj8_2(.din(w_dff_B_6GS2D6WL2_2),.dout(w_dff_B_bahWkaCj8_2),.clk(gclk));
	jdff dff_B_P4I6i2BR0_2(.din(w_dff_B_bahWkaCj8_2),.dout(w_dff_B_P4I6i2BR0_2),.clk(gclk));
	jdff dff_B_wmB8RHgA4_2(.din(w_dff_B_P4I6i2BR0_2),.dout(w_dff_B_wmB8RHgA4_2),.clk(gclk));
	jdff dff_B_8MtvksDq9_2(.din(w_dff_B_wmB8RHgA4_2),.dout(w_dff_B_8MtvksDq9_2),.clk(gclk));
	jdff dff_B_9rkhLf1N1_2(.din(w_dff_B_8MtvksDq9_2),.dout(w_dff_B_9rkhLf1N1_2),.clk(gclk));
	jdff dff_B_20zguyvu0_2(.din(w_dff_B_9rkhLf1N1_2),.dout(w_dff_B_20zguyvu0_2),.clk(gclk));
	jdff dff_B_eem8j2Qn0_2(.din(w_dff_B_20zguyvu0_2),.dout(w_dff_B_eem8j2Qn0_2),.clk(gclk));
	jdff dff_B_ytUTXs197_2(.din(w_dff_B_eem8j2Qn0_2),.dout(w_dff_B_ytUTXs197_2),.clk(gclk));
	jdff dff_B_0KZ9AP1K8_2(.din(w_dff_B_ytUTXs197_2),.dout(w_dff_B_0KZ9AP1K8_2),.clk(gclk));
	jdff dff_B_0vm24MMq6_2(.din(w_dff_B_0KZ9AP1K8_2),.dout(w_dff_B_0vm24MMq6_2),.clk(gclk));
	jdff dff_B_XkyvqK3f5_2(.din(w_dff_B_0vm24MMq6_2),.dout(w_dff_B_XkyvqK3f5_2),.clk(gclk));
	jdff dff_B_1opj1cZ63_2(.din(w_dff_B_XkyvqK3f5_2),.dout(w_dff_B_1opj1cZ63_2),.clk(gclk));
	jdff dff_B_hpXRjjSe9_2(.din(w_dff_B_1opj1cZ63_2),.dout(w_dff_B_hpXRjjSe9_2),.clk(gclk));
	jdff dff_B_43zgnGut4_2(.din(w_dff_B_hpXRjjSe9_2),.dout(w_dff_B_43zgnGut4_2),.clk(gclk));
	jdff dff_B_A9Ks2ZsT2_2(.din(w_dff_B_43zgnGut4_2),.dout(w_dff_B_A9Ks2ZsT2_2),.clk(gclk));
	jdff dff_B_DsWwJvHK1_2(.din(w_dff_B_A9Ks2ZsT2_2),.dout(w_dff_B_DsWwJvHK1_2),.clk(gclk));
	jdff dff_B_uBt2GzZg2_2(.din(w_dff_B_DsWwJvHK1_2),.dout(w_dff_B_uBt2GzZg2_2),.clk(gclk));
	jdff dff_B_0fsiTw3x3_2(.din(w_dff_B_uBt2GzZg2_2),.dout(w_dff_B_0fsiTw3x3_2),.clk(gclk));
	jdff dff_B_jFZNP46H3_2(.din(w_dff_B_0fsiTw3x3_2),.dout(w_dff_B_jFZNP46H3_2),.clk(gclk));
	jdff dff_B_SWmWQhEh6_2(.din(w_dff_B_jFZNP46H3_2),.dout(w_dff_B_SWmWQhEh6_2),.clk(gclk));
	jdff dff_B_n6F17ieo9_2(.din(w_dff_B_SWmWQhEh6_2),.dout(w_dff_B_n6F17ieo9_2),.clk(gclk));
	jdff dff_B_bwYKO1Fa7_2(.din(w_dff_B_n6F17ieo9_2),.dout(w_dff_B_bwYKO1Fa7_2),.clk(gclk));
	jdff dff_B_vVJPDswb5_2(.din(w_dff_B_bwYKO1Fa7_2),.dout(w_dff_B_vVJPDswb5_2),.clk(gclk));
	jdff dff_B_nCC9fcAH6_2(.din(w_dff_B_vVJPDswb5_2),.dout(w_dff_B_nCC9fcAH6_2),.clk(gclk));
	jdff dff_B_Q9418DGX7_2(.din(w_dff_B_nCC9fcAH6_2),.dout(w_dff_B_Q9418DGX7_2),.clk(gclk));
	jdff dff_B_zHfX8UyQ3_2(.din(w_dff_B_Q9418DGX7_2),.dout(w_dff_B_zHfX8UyQ3_2),.clk(gclk));
	jdff dff_B_1Wmbdlxi2_2(.din(w_dff_B_zHfX8UyQ3_2),.dout(w_dff_B_1Wmbdlxi2_2),.clk(gclk));
	jdff dff_B_JFgwEwTC7_2(.din(n1525),.dout(w_dff_B_JFgwEwTC7_2),.clk(gclk));
	jdff dff_B_9L9nGFxd7_1(.din(n1523),.dout(w_dff_B_9L9nGFxd7_1),.clk(gclk));
	jdff dff_B_fav47N7a8_2(.din(n1451),.dout(w_dff_B_fav47N7a8_2),.clk(gclk));
	jdff dff_B_vUEzVpX84_2(.din(w_dff_B_fav47N7a8_2),.dout(w_dff_B_vUEzVpX84_2),.clk(gclk));
	jdff dff_B_mSeKqQ5c7_2(.din(w_dff_B_vUEzVpX84_2),.dout(w_dff_B_mSeKqQ5c7_2),.clk(gclk));
	jdff dff_B_yGvZgSGm0_2(.din(w_dff_B_mSeKqQ5c7_2),.dout(w_dff_B_yGvZgSGm0_2),.clk(gclk));
	jdff dff_B_tzXtrQJ47_2(.din(w_dff_B_yGvZgSGm0_2),.dout(w_dff_B_tzXtrQJ47_2),.clk(gclk));
	jdff dff_B_fsYCljgR8_2(.din(w_dff_B_tzXtrQJ47_2),.dout(w_dff_B_fsYCljgR8_2),.clk(gclk));
	jdff dff_B_zOUDat0H1_2(.din(w_dff_B_fsYCljgR8_2),.dout(w_dff_B_zOUDat0H1_2),.clk(gclk));
	jdff dff_B_XOJTIFOE6_2(.din(w_dff_B_zOUDat0H1_2),.dout(w_dff_B_XOJTIFOE6_2),.clk(gclk));
	jdff dff_B_7v3WGehJ8_2(.din(w_dff_B_XOJTIFOE6_2),.dout(w_dff_B_7v3WGehJ8_2),.clk(gclk));
	jdff dff_B_zwNYJRdG9_2(.din(w_dff_B_7v3WGehJ8_2),.dout(w_dff_B_zwNYJRdG9_2),.clk(gclk));
	jdff dff_B_zM3snEyE4_2(.din(w_dff_B_zwNYJRdG9_2),.dout(w_dff_B_zM3snEyE4_2),.clk(gclk));
	jdff dff_B_lL1Lr7pY7_2(.din(w_dff_B_zM3snEyE4_2),.dout(w_dff_B_lL1Lr7pY7_2),.clk(gclk));
	jdff dff_B_5C1maZMv7_2(.din(w_dff_B_lL1Lr7pY7_2),.dout(w_dff_B_5C1maZMv7_2),.clk(gclk));
	jdff dff_B_Hv9BOByu3_2(.din(w_dff_B_5C1maZMv7_2),.dout(w_dff_B_Hv9BOByu3_2),.clk(gclk));
	jdff dff_B_TXexaVhe4_2(.din(w_dff_B_Hv9BOByu3_2),.dout(w_dff_B_TXexaVhe4_2),.clk(gclk));
	jdff dff_B_8CUlMfc80_2(.din(w_dff_B_TXexaVhe4_2),.dout(w_dff_B_8CUlMfc80_2),.clk(gclk));
	jdff dff_B_ouH1gUc92_2(.din(w_dff_B_8CUlMfc80_2),.dout(w_dff_B_ouH1gUc92_2),.clk(gclk));
	jdff dff_B_h9PFo6nE5_2(.din(w_dff_B_ouH1gUc92_2),.dout(w_dff_B_h9PFo6nE5_2),.clk(gclk));
	jdff dff_B_xdJXjwU11_2(.din(w_dff_B_h9PFo6nE5_2),.dout(w_dff_B_xdJXjwU11_2),.clk(gclk));
	jdff dff_B_LKbqQDaE5_2(.din(w_dff_B_xdJXjwU11_2),.dout(w_dff_B_LKbqQDaE5_2),.clk(gclk));
	jdff dff_B_eoHwu7zi4_2(.din(w_dff_B_LKbqQDaE5_2),.dout(w_dff_B_eoHwu7zi4_2),.clk(gclk));
	jdff dff_B_ib0wdVZA5_2(.din(w_dff_B_eoHwu7zi4_2),.dout(w_dff_B_ib0wdVZA5_2),.clk(gclk));
	jdff dff_B_kHLkJIBB8_2(.din(w_dff_B_ib0wdVZA5_2),.dout(w_dff_B_kHLkJIBB8_2),.clk(gclk));
	jdff dff_B_nTmDnv9l4_2(.din(w_dff_B_kHLkJIBB8_2),.dout(w_dff_B_nTmDnv9l4_2),.clk(gclk));
	jdff dff_B_rjZuGj266_2(.din(w_dff_B_nTmDnv9l4_2),.dout(w_dff_B_rjZuGj266_2),.clk(gclk));
	jdff dff_B_LE2cHTDX0_2(.din(w_dff_B_rjZuGj266_2),.dout(w_dff_B_LE2cHTDX0_2),.clk(gclk));
	jdff dff_B_R7eja0Cs2_2(.din(w_dff_B_LE2cHTDX0_2),.dout(w_dff_B_R7eja0Cs2_2),.clk(gclk));
	jdff dff_B_4NG8Ychw2_2(.din(w_dff_B_R7eja0Cs2_2),.dout(w_dff_B_4NG8Ychw2_2),.clk(gclk));
	jdff dff_B_1Nd5QAbS8_2(.din(w_dff_B_4NG8Ychw2_2),.dout(w_dff_B_1Nd5QAbS8_2),.clk(gclk));
	jdff dff_B_hg36VsNB6_2(.din(n1454),.dout(w_dff_B_hg36VsNB6_2),.clk(gclk));
	jdff dff_B_oNsStTFp5_1(.din(n1452),.dout(w_dff_B_oNsStTFp5_1),.clk(gclk));
	jdff dff_B_oHmv5qXR6_2(.din(n1373),.dout(w_dff_B_oHmv5qXR6_2),.clk(gclk));
	jdff dff_B_NZgkpkxH2_2(.din(w_dff_B_oHmv5qXR6_2),.dout(w_dff_B_NZgkpkxH2_2),.clk(gclk));
	jdff dff_B_rDQfFCGb5_2(.din(w_dff_B_NZgkpkxH2_2),.dout(w_dff_B_rDQfFCGb5_2),.clk(gclk));
	jdff dff_B_aCA50iKr5_2(.din(w_dff_B_rDQfFCGb5_2),.dout(w_dff_B_aCA50iKr5_2),.clk(gclk));
	jdff dff_B_6k1sIwv72_2(.din(w_dff_B_aCA50iKr5_2),.dout(w_dff_B_6k1sIwv72_2),.clk(gclk));
	jdff dff_B_F22AP4UG6_2(.din(w_dff_B_6k1sIwv72_2),.dout(w_dff_B_F22AP4UG6_2),.clk(gclk));
	jdff dff_B_B0ucpamH0_2(.din(w_dff_B_F22AP4UG6_2),.dout(w_dff_B_B0ucpamH0_2),.clk(gclk));
	jdff dff_B_ZpIMM9nD3_2(.din(w_dff_B_B0ucpamH0_2),.dout(w_dff_B_ZpIMM9nD3_2),.clk(gclk));
	jdff dff_B_nrmH1mBP0_2(.din(w_dff_B_ZpIMM9nD3_2),.dout(w_dff_B_nrmH1mBP0_2),.clk(gclk));
	jdff dff_B_yxFTUBzI4_2(.din(w_dff_B_nrmH1mBP0_2),.dout(w_dff_B_yxFTUBzI4_2),.clk(gclk));
	jdff dff_B_p6vil0Wl2_2(.din(w_dff_B_yxFTUBzI4_2),.dout(w_dff_B_p6vil0Wl2_2),.clk(gclk));
	jdff dff_B_cHaKcw4M2_2(.din(w_dff_B_p6vil0Wl2_2),.dout(w_dff_B_cHaKcw4M2_2),.clk(gclk));
	jdff dff_B_aogjyaBg9_2(.din(w_dff_B_cHaKcw4M2_2),.dout(w_dff_B_aogjyaBg9_2),.clk(gclk));
	jdff dff_B_wtCTFTy29_2(.din(w_dff_B_aogjyaBg9_2),.dout(w_dff_B_wtCTFTy29_2),.clk(gclk));
	jdff dff_B_0i6o4roQ2_2(.din(w_dff_B_wtCTFTy29_2),.dout(w_dff_B_0i6o4roQ2_2),.clk(gclk));
	jdff dff_B_DFu1ENa23_2(.din(w_dff_B_0i6o4roQ2_2),.dout(w_dff_B_DFu1ENa23_2),.clk(gclk));
	jdff dff_B_kjPesmOp9_2(.din(w_dff_B_DFu1ENa23_2),.dout(w_dff_B_kjPesmOp9_2),.clk(gclk));
	jdff dff_B_Ytcb8UoX6_2(.din(w_dff_B_kjPesmOp9_2),.dout(w_dff_B_Ytcb8UoX6_2),.clk(gclk));
	jdff dff_B_OfeB5gDa3_2(.din(w_dff_B_Ytcb8UoX6_2),.dout(w_dff_B_OfeB5gDa3_2),.clk(gclk));
	jdff dff_B_GLibKxEC7_2(.din(w_dff_B_OfeB5gDa3_2),.dout(w_dff_B_GLibKxEC7_2),.clk(gclk));
	jdff dff_B_gYCGV48K5_2(.din(w_dff_B_GLibKxEC7_2),.dout(w_dff_B_gYCGV48K5_2),.clk(gclk));
	jdff dff_B_Ak3YZDbs5_2(.din(w_dff_B_gYCGV48K5_2),.dout(w_dff_B_Ak3YZDbs5_2),.clk(gclk));
	jdff dff_B_oMftZqqS6_2(.din(w_dff_B_Ak3YZDbs5_2),.dout(w_dff_B_oMftZqqS6_2),.clk(gclk));
	jdff dff_B_2PNucZHP1_2(.din(w_dff_B_oMftZqqS6_2),.dout(w_dff_B_2PNucZHP1_2),.clk(gclk));
	jdff dff_B_Dq6CTl2L9_2(.din(w_dff_B_2PNucZHP1_2),.dout(w_dff_B_Dq6CTl2L9_2),.clk(gclk));
	jdff dff_B_IYIt1woL4_2(.din(n1376),.dout(w_dff_B_IYIt1woL4_2),.clk(gclk));
	jdff dff_B_GJ7x2nk19_1(.din(n1374),.dout(w_dff_B_GJ7x2nk19_1),.clk(gclk));
	jdff dff_B_YrNXONms6_2(.din(n1288),.dout(w_dff_B_YrNXONms6_2),.clk(gclk));
	jdff dff_B_5ZG9u9ZI9_2(.din(w_dff_B_YrNXONms6_2),.dout(w_dff_B_5ZG9u9ZI9_2),.clk(gclk));
	jdff dff_B_1Ze3lasn0_2(.din(w_dff_B_5ZG9u9ZI9_2),.dout(w_dff_B_1Ze3lasn0_2),.clk(gclk));
	jdff dff_B_zSvF6KbM8_2(.din(w_dff_B_1Ze3lasn0_2),.dout(w_dff_B_zSvF6KbM8_2),.clk(gclk));
	jdff dff_B_YXlU9lrF2_2(.din(w_dff_B_zSvF6KbM8_2),.dout(w_dff_B_YXlU9lrF2_2),.clk(gclk));
	jdff dff_B_EPTjINBL6_2(.din(w_dff_B_YXlU9lrF2_2),.dout(w_dff_B_EPTjINBL6_2),.clk(gclk));
	jdff dff_B_qaMRMaTs9_2(.din(w_dff_B_EPTjINBL6_2),.dout(w_dff_B_qaMRMaTs9_2),.clk(gclk));
	jdff dff_B_OgC9dRfe4_2(.din(w_dff_B_qaMRMaTs9_2),.dout(w_dff_B_OgC9dRfe4_2),.clk(gclk));
	jdff dff_B_OcOJGZyC7_2(.din(w_dff_B_OgC9dRfe4_2),.dout(w_dff_B_OcOJGZyC7_2),.clk(gclk));
	jdff dff_B_BxtNQLdp8_2(.din(w_dff_B_OcOJGZyC7_2),.dout(w_dff_B_BxtNQLdp8_2),.clk(gclk));
	jdff dff_B_qgFBy6918_2(.din(w_dff_B_BxtNQLdp8_2),.dout(w_dff_B_qgFBy6918_2),.clk(gclk));
	jdff dff_B_n5GFp7w90_2(.din(w_dff_B_qgFBy6918_2),.dout(w_dff_B_n5GFp7w90_2),.clk(gclk));
	jdff dff_B_8MBLqyIJ4_2(.din(w_dff_B_n5GFp7w90_2),.dout(w_dff_B_8MBLqyIJ4_2),.clk(gclk));
	jdff dff_B_HDEZdqV55_2(.din(w_dff_B_8MBLqyIJ4_2),.dout(w_dff_B_HDEZdqV55_2),.clk(gclk));
	jdff dff_B_SDJSmfqO0_2(.din(w_dff_B_HDEZdqV55_2),.dout(w_dff_B_SDJSmfqO0_2),.clk(gclk));
	jdff dff_B_LXZwxnQa9_2(.din(w_dff_B_SDJSmfqO0_2),.dout(w_dff_B_LXZwxnQa9_2),.clk(gclk));
	jdff dff_B_3Q1D1rBf2_2(.din(w_dff_B_LXZwxnQa9_2),.dout(w_dff_B_3Q1D1rBf2_2),.clk(gclk));
	jdff dff_B_pVFPtswd1_2(.din(w_dff_B_3Q1D1rBf2_2),.dout(w_dff_B_pVFPtswd1_2),.clk(gclk));
	jdff dff_B_w0kiJNFI2_2(.din(w_dff_B_pVFPtswd1_2),.dout(w_dff_B_w0kiJNFI2_2),.clk(gclk));
	jdff dff_B_uVhiqHwO3_2(.din(w_dff_B_w0kiJNFI2_2),.dout(w_dff_B_uVhiqHwO3_2),.clk(gclk));
	jdff dff_B_sEnDKUqv7_2(.din(w_dff_B_uVhiqHwO3_2),.dout(w_dff_B_sEnDKUqv7_2),.clk(gclk));
	jdff dff_B_3ek4XcaU4_1(.din(n1289),.dout(w_dff_B_3ek4XcaU4_1),.clk(gclk));
	jdff dff_B_lJ7C1RDt4_2(.din(n1198),.dout(w_dff_B_lJ7C1RDt4_2),.clk(gclk));
	jdff dff_B_FO3yi2lv8_2(.din(w_dff_B_lJ7C1RDt4_2),.dout(w_dff_B_FO3yi2lv8_2),.clk(gclk));
	jdff dff_B_GUmy7p0p6_2(.din(w_dff_B_FO3yi2lv8_2),.dout(w_dff_B_GUmy7p0p6_2),.clk(gclk));
	jdff dff_B_DyutjSWN5_2(.din(w_dff_B_GUmy7p0p6_2),.dout(w_dff_B_DyutjSWN5_2),.clk(gclk));
	jdff dff_B_MXBeQyFu9_2(.din(w_dff_B_DyutjSWN5_2),.dout(w_dff_B_MXBeQyFu9_2),.clk(gclk));
	jdff dff_B_3A2UMLPS5_2(.din(w_dff_B_MXBeQyFu9_2),.dout(w_dff_B_3A2UMLPS5_2),.clk(gclk));
	jdff dff_B_EbZpbqqa4_2(.din(w_dff_B_3A2UMLPS5_2),.dout(w_dff_B_EbZpbqqa4_2),.clk(gclk));
	jdff dff_B_rL8qINCn0_2(.din(w_dff_B_EbZpbqqa4_2),.dout(w_dff_B_rL8qINCn0_2),.clk(gclk));
	jdff dff_B_cvGRX6as8_2(.din(w_dff_B_rL8qINCn0_2),.dout(w_dff_B_cvGRX6as8_2),.clk(gclk));
	jdff dff_B_kUGaiZG37_2(.din(w_dff_B_cvGRX6as8_2),.dout(w_dff_B_kUGaiZG37_2),.clk(gclk));
	jdff dff_B_6eYryBY42_2(.din(w_dff_B_kUGaiZG37_2),.dout(w_dff_B_6eYryBY42_2),.clk(gclk));
	jdff dff_B_0z6X96Rf4_2(.din(w_dff_B_6eYryBY42_2),.dout(w_dff_B_0z6X96Rf4_2),.clk(gclk));
	jdff dff_B_dpRxWuvB5_2(.din(w_dff_B_0z6X96Rf4_2),.dout(w_dff_B_dpRxWuvB5_2),.clk(gclk));
	jdff dff_B_CyniIOTJ5_2(.din(w_dff_B_dpRxWuvB5_2),.dout(w_dff_B_CyniIOTJ5_2),.clk(gclk));
	jdff dff_B_RyO1k4AJ4_2(.din(w_dff_B_CyniIOTJ5_2),.dout(w_dff_B_RyO1k4AJ4_2),.clk(gclk));
	jdff dff_B_Nsh1AuaP6_2(.din(w_dff_B_RyO1k4AJ4_2),.dout(w_dff_B_Nsh1AuaP6_2),.clk(gclk));
	jdff dff_B_n59VXHVa0_2(.din(w_dff_B_Nsh1AuaP6_2),.dout(w_dff_B_n59VXHVa0_2),.clk(gclk));
	jdff dff_B_65EnfEbg5_2(.din(w_dff_B_n59VXHVa0_2),.dout(w_dff_B_65EnfEbg5_2),.clk(gclk));
	jdff dff_B_OSqXrNmC5_2(.din(n1215),.dout(w_dff_B_OSqXrNmC5_2),.clk(gclk));
	jdff dff_B_AINmtyNJ6_1(.din(n1199),.dout(w_dff_B_AINmtyNJ6_1),.clk(gclk));
	jdff dff_B_iK2mAFDW3_2(.din(n1094),.dout(w_dff_B_iK2mAFDW3_2),.clk(gclk));
	jdff dff_B_PCD0TPj07_2(.din(w_dff_B_iK2mAFDW3_2),.dout(w_dff_B_PCD0TPj07_2),.clk(gclk));
	jdff dff_B_b6276lxL4_2(.din(w_dff_B_PCD0TPj07_2),.dout(w_dff_B_b6276lxL4_2),.clk(gclk));
	jdff dff_B_wTwB5vvR5_2(.din(w_dff_B_b6276lxL4_2),.dout(w_dff_B_wTwB5vvR5_2),.clk(gclk));
	jdff dff_B_eqJobM641_2(.din(w_dff_B_wTwB5vvR5_2),.dout(w_dff_B_eqJobM641_2),.clk(gclk));
	jdff dff_B_V5uOjYkI2_2(.din(w_dff_B_eqJobM641_2),.dout(w_dff_B_V5uOjYkI2_2),.clk(gclk));
	jdff dff_B_FWrQbHA09_2(.din(w_dff_B_V5uOjYkI2_2),.dout(w_dff_B_FWrQbHA09_2),.clk(gclk));
	jdff dff_B_QpfJ0azY9_2(.din(w_dff_B_FWrQbHA09_2),.dout(w_dff_B_QpfJ0azY9_2),.clk(gclk));
	jdff dff_B_2kAvn4pW1_2(.din(w_dff_B_QpfJ0azY9_2),.dout(w_dff_B_2kAvn4pW1_2),.clk(gclk));
	jdff dff_B_siEFPnIM9_2(.din(w_dff_B_2kAvn4pW1_2),.dout(w_dff_B_siEFPnIM9_2),.clk(gclk));
	jdff dff_B_IwFsrmHY7_2(.din(w_dff_B_siEFPnIM9_2),.dout(w_dff_B_IwFsrmHY7_2),.clk(gclk));
	jdff dff_B_4ZJQmA1u2_2(.din(w_dff_B_IwFsrmHY7_2),.dout(w_dff_B_4ZJQmA1u2_2),.clk(gclk));
	jdff dff_B_Jyg6YH0c9_2(.din(w_dff_B_4ZJQmA1u2_2),.dout(w_dff_B_Jyg6YH0c9_2),.clk(gclk));
	jdff dff_B_2MCgcwcC5_2(.din(w_dff_B_Jyg6YH0c9_2),.dout(w_dff_B_2MCgcwcC5_2),.clk(gclk));
	jdff dff_B_ZfiCaKEH3_2(.din(w_dff_B_2MCgcwcC5_2),.dout(w_dff_B_ZfiCaKEH3_2),.clk(gclk));
	jdff dff_B_hQnr7CKb1_2(.din(n1117),.dout(w_dff_B_hQnr7CKb1_2),.clk(gclk));
	jdff dff_B_tsN5TVO52_2(.din(w_dff_B_hQnr7CKb1_2),.dout(w_dff_B_tsN5TVO52_2),.clk(gclk));
	jdff dff_B_9lRe7hy55_1(.din(n1095),.dout(w_dff_B_9lRe7hy55_1),.clk(gclk));
	jdff dff_B_1lJKtMc85_2(.din(n996),.dout(w_dff_B_1lJKtMc85_2),.clk(gclk));
	jdff dff_B_jppu77Gt1_2(.din(w_dff_B_1lJKtMc85_2),.dout(w_dff_B_jppu77Gt1_2),.clk(gclk));
	jdff dff_B_LSv5OsKr9_2(.din(w_dff_B_jppu77Gt1_2),.dout(w_dff_B_LSv5OsKr9_2),.clk(gclk));
	jdff dff_B_UFnpmM8a5_2(.din(w_dff_B_LSv5OsKr9_2),.dout(w_dff_B_UFnpmM8a5_2),.clk(gclk));
	jdff dff_B_mmUVITa76_2(.din(w_dff_B_UFnpmM8a5_2),.dout(w_dff_B_mmUVITa76_2),.clk(gclk));
	jdff dff_B_WAzqaay31_2(.din(w_dff_B_mmUVITa76_2),.dout(w_dff_B_WAzqaay31_2),.clk(gclk));
	jdff dff_B_3BPAC2gE2_2(.din(w_dff_B_WAzqaay31_2),.dout(w_dff_B_3BPAC2gE2_2),.clk(gclk));
	jdff dff_B_OPDbgvjk9_2(.din(w_dff_B_3BPAC2gE2_2),.dout(w_dff_B_OPDbgvjk9_2),.clk(gclk));
	jdff dff_B_gRQjQGh94_2(.din(w_dff_B_OPDbgvjk9_2),.dout(w_dff_B_gRQjQGh94_2),.clk(gclk));
	jdff dff_B_pcqWMDNl5_2(.din(w_dff_B_gRQjQGh94_2),.dout(w_dff_B_pcqWMDNl5_2),.clk(gclk));
	jdff dff_B_nFu9CEJG0_2(.din(w_dff_B_pcqWMDNl5_2),.dout(w_dff_B_nFu9CEJG0_2),.clk(gclk));
	jdff dff_B_23rRmjYY1_2(.din(w_dff_B_nFu9CEJG0_2),.dout(w_dff_B_23rRmjYY1_2),.clk(gclk));
	jdff dff_B_FiJjNlFe1_2(.din(n1012),.dout(w_dff_B_FiJjNlFe1_2),.clk(gclk));
	jdff dff_B_ok5zClye5_2(.din(w_dff_B_FiJjNlFe1_2),.dout(w_dff_B_ok5zClye5_2),.clk(gclk));
	jdff dff_B_aSMKxdg69_1(.din(n997),.dout(w_dff_B_aSMKxdg69_1),.clk(gclk));
	jdff dff_B_mjik72bq7_2(.din(n891),.dout(w_dff_B_mjik72bq7_2),.clk(gclk));
	jdff dff_B_RY9mRFZd0_2(.din(w_dff_B_mjik72bq7_2),.dout(w_dff_B_RY9mRFZd0_2),.clk(gclk));
	jdff dff_B_xSHMoOkf1_2(.din(w_dff_B_RY9mRFZd0_2),.dout(w_dff_B_xSHMoOkf1_2),.clk(gclk));
	jdff dff_B_K0Lx7DLD7_2(.din(w_dff_B_xSHMoOkf1_2),.dout(w_dff_B_K0Lx7DLD7_2),.clk(gclk));
	jdff dff_B_AeZXW2289_2(.din(w_dff_B_K0Lx7DLD7_2),.dout(w_dff_B_AeZXW2289_2),.clk(gclk));
	jdff dff_B_QaVHFWPL4_2(.din(w_dff_B_AeZXW2289_2),.dout(w_dff_B_QaVHFWPL4_2),.clk(gclk));
	jdff dff_B_zaEV6AUQ7_2(.din(w_dff_B_QaVHFWPL4_2),.dout(w_dff_B_zaEV6AUQ7_2),.clk(gclk));
	jdff dff_B_OSsHow5H5_2(.din(w_dff_B_zaEV6AUQ7_2),.dout(w_dff_B_OSsHow5H5_2),.clk(gclk));
	jdff dff_B_3FIpdvcG0_2(.din(w_dff_B_OSsHow5H5_2),.dout(w_dff_B_3FIpdvcG0_2),.clk(gclk));
	jdff dff_B_tcFqXBI95_2(.din(n907),.dout(w_dff_B_tcFqXBI95_2),.clk(gclk));
	jdff dff_B_43zDDGAx6_2(.din(w_dff_B_tcFqXBI95_2),.dout(w_dff_B_43zDDGAx6_2),.clk(gclk));
	jdff dff_B_CF3fq3pc5_2(.din(w_dff_B_43zDDGAx6_2),.dout(w_dff_B_CF3fq3pc5_2),.clk(gclk));
	jdff dff_B_YfhrVjh72_1(.din(n892),.dout(w_dff_B_YfhrVjh72_1),.clk(gclk));
	jdff dff_B_6849uQSw6_1(.din(w_dff_B_YfhrVjh72_1),.dout(w_dff_B_6849uQSw6_1),.clk(gclk));
	jdff dff_B_wWYbSLJf7_1(.din(w_dff_B_6849uQSw6_1),.dout(w_dff_B_wWYbSLJf7_1),.clk(gclk));
	jdff dff_B_FFR5M8UT0_1(.din(w_dff_B_wWYbSLJf7_1),.dout(w_dff_B_FFR5M8UT0_1),.clk(gclk));
	jdff dff_B_xmythnXI6_1(.din(w_dff_B_FFR5M8UT0_1),.dout(w_dff_B_xmythnXI6_1),.clk(gclk));
	jdff dff_B_ewdCX36A1_1(.din(w_dff_B_xmythnXI6_1),.dout(w_dff_B_ewdCX36A1_1),.clk(gclk));
	jdff dff_B_8judfUTY8_0(.din(n801),.dout(w_dff_B_8judfUTY8_0),.clk(gclk));
	jdff dff_B_d7N1ZYqq2_0(.din(w_dff_B_8judfUTY8_0),.dout(w_dff_B_d7N1ZYqq2_0),.clk(gclk));
	jdff dff_A_l2pq6lHB9_0(.dout(w_n800_0[0]),.din(w_dff_A_l2pq6lHB9_0),.clk(gclk));
	jdff dff_A_7YwHJFsi2_0(.dout(w_dff_A_l2pq6lHB9_0),.din(w_dff_A_7YwHJFsi2_0),.clk(gclk));
	jdff dff_A_CxS8Eef66_0(.dout(w_dff_A_7YwHJFsi2_0),.din(w_dff_A_CxS8Eef66_0),.clk(gclk));
	jdff dff_B_zrpbKDpH7_1(.din(n794),.dout(w_dff_B_zrpbKDpH7_1),.clk(gclk));
	jdff dff_A_T2OwA3n83_0(.dout(w_n698_0[0]),.din(w_dff_A_T2OwA3n83_0),.clk(gclk));
	jdff dff_A_NGDQpmyY8_1(.dout(w_n698_0[1]),.din(w_dff_A_NGDQpmyY8_1),.clk(gclk));
	jdff dff_A_45MFTm1j1_1(.dout(w_dff_A_NGDQpmyY8_1),.din(w_dff_A_45MFTm1j1_1),.clk(gclk));
	jdff dff_A_d2Qncvh02_1(.dout(w_n792_0[1]),.din(w_dff_A_d2Qncvh02_1),.clk(gclk));
	jdff dff_A_U5mbdxMM8_1(.dout(w_dff_A_d2Qncvh02_1),.din(w_dff_A_U5mbdxMM8_1),.clk(gclk));
	jdff dff_A_4LbXaeqt2_1(.dout(w_dff_A_U5mbdxMM8_1),.din(w_dff_A_4LbXaeqt2_1),.clk(gclk));
	jdff dff_A_fFWhP3vZ1_1(.dout(w_dff_A_4LbXaeqt2_1),.din(w_dff_A_fFWhP3vZ1_1),.clk(gclk));
	jdff dff_A_evkcmivS0_1(.dout(w_dff_A_fFWhP3vZ1_1),.din(w_dff_A_evkcmivS0_1),.clk(gclk));
	jdff dff_A_kO1gTAnV0_1(.dout(w_dff_A_evkcmivS0_1),.din(w_dff_A_kO1gTAnV0_1),.clk(gclk));
	jdff dff_B_jCAK1uKJ6_1(.din(n1843),.dout(w_dff_B_jCAK1uKJ6_1),.clk(gclk));
	jdff dff_B_m74SQWxQ6_1(.din(n1830),.dout(w_dff_B_m74SQWxQ6_1),.clk(gclk));
	jdff dff_B_SykyZ5wE9_1(.din(w_dff_B_m74SQWxQ6_1),.dout(w_dff_B_SykyZ5wE9_1),.clk(gclk));
	jdff dff_B_CUxnaWaM1_2(.din(n1829),.dout(w_dff_B_CUxnaWaM1_2),.clk(gclk));
	jdff dff_B_b28AAknA0_2(.din(w_dff_B_CUxnaWaM1_2),.dout(w_dff_B_b28AAknA0_2),.clk(gclk));
	jdff dff_B_2F6PUUyV0_2(.din(w_dff_B_b28AAknA0_2),.dout(w_dff_B_2F6PUUyV0_2),.clk(gclk));
	jdff dff_B_skppOEvw0_2(.din(w_dff_B_2F6PUUyV0_2),.dout(w_dff_B_skppOEvw0_2),.clk(gclk));
	jdff dff_B_qCm9mVjM7_2(.din(w_dff_B_skppOEvw0_2),.dout(w_dff_B_qCm9mVjM7_2),.clk(gclk));
	jdff dff_B_3XdIOSMc7_2(.din(w_dff_B_qCm9mVjM7_2),.dout(w_dff_B_3XdIOSMc7_2),.clk(gclk));
	jdff dff_B_BK5kXT6W0_2(.din(w_dff_B_3XdIOSMc7_2),.dout(w_dff_B_BK5kXT6W0_2),.clk(gclk));
	jdff dff_B_9FxtHGkt3_2(.din(w_dff_B_BK5kXT6W0_2),.dout(w_dff_B_9FxtHGkt3_2),.clk(gclk));
	jdff dff_B_YrICbcdI5_2(.din(w_dff_B_9FxtHGkt3_2),.dout(w_dff_B_YrICbcdI5_2),.clk(gclk));
	jdff dff_B_8qfAlAIl3_2(.din(w_dff_B_YrICbcdI5_2),.dout(w_dff_B_8qfAlAIl3_2),.clk(gclk));
	jdff dff_B_NVIIEGVa5_2(.din(w_dff_B_8qfAlAIl3_2),.dout(w_dff_B_NVIIEGVa5_2),.clk(gclk));
	jdff dff_B_iSr6Q6Ml7_2(.din(w_dff_B_NVIIEGVa5_2),.dout(w_dff_B_iSr6Q6Ml7_2),.clk(gclk));
	jdff dff_B_iSNbBS7X0_2(.din(w_dff_B_iSr6Q6Ml7_2),.dout(w_dff_B_iSNbBS7X0_2),.clk(gclk));
	jdff dff_B_iXZyuVYv1_2(.din(w_dff_B_iSNbBS7X0_2),.dout(w_dff_B_iXZyuVYv1_2),.clk(gclk));
	jdff dff_B_3v1zFld53_2(.din(w_dff_B_iXZyuVYv1_2),.dout(w_dff_B_3v1zFld53_2),.clk(gclk));
	jdff dff_B_t6yA3jm96_2(.din(w_dff_B_3v1zFld53_2),.dout(w_dff_B_t6yA3jm96_2),.clk(gclk));
	jdff dff_B_eDKF1vgK6_2(.din(w_dff_B_t6yA3jm96_2),.dout(w_dff_B_eDKF1vgK6_2),.clk(gclk));
	jdff dff_B_g0hTqjNL0_2(.din(w_dff_B_eDKF1vgK6_2),.dout(w_dff_B_g0hTqjNL0_2),.clk(gclk));
	jdff dff_B_KkZANGyg3_2(.din(w_dff_B_g0hTqjNL0_2),.dout(w_dff_B_KkZANGyg3_2),.clk(gclk));
	jdff dff_B_S4c2Pgr29_2(.din(w_dff_B_KkZANGyg3_2),.dout(w_dff_B_S4c2Pgr29_2),.clk(gclk));
	jdff dff_B_4NnsSIQ28_2(.din(w_dff_B_S4c2Pgr29_2),.dout(w_dff_B_4NnsSIQ28_2),.clk(gclk));
	jdff dff_B_YsQ2ps2v5_2(.din(w_dff_B_4NnsSIQ28_2),.dout(w_dff_B_YsQ2ps2v5_2),.clk(gclk));
	jdff dff_B_OuqYkvnT0_2(.din(w_dff_B_YsQ2ps2v5_2),.dout(w_dff_B_OuqYkvnT0_2),.clk(gclk));
	jdff dff_B_Tcb3BKtD3_2(.din(w_dff_B_OuqYkvnT0_2),.dout(w_dff_B_Tcb3BKtD3_2),.clk(gclk));
	jdff dff_B_pqwEOZ3h2_2(.din(w_dff_B_Tcb3BKtD3_2),.dout(w_dff_B_pqwEOZ3h2_2),.clk(gclk));
	jdff dff_B_HOgzSMcM2_2(.din(w_dff_B_pqwEOZ3h2_2),.dout(w_dff_B_HOgzSMcM2_2),.clk(gclk));
	jdff dff_B_FQ59q70x2_2(.din(w_dff_B_HOgzSMcM2_2),.dout(w_dff_B_FQ59q70x2_2),.clk(gclk));
	jdff dff_B_yvBEuBC50_2(.din(w_dff_B_FQ59q70x2_2),.dout(w_dff_B_yvBEuBC50_2),.clk(gclk));
	jdff dff_B_oWrJkv4c0_2(.din(w_dff_B_yvBEuBC50_2),.dout(w_dff_B_oWrJkv4c0_2),.clk(gclk));
	jdff dff_B_O1VL38gO8_2(.din(w_dff_B_oWrJkv4c0_2),.dout(w_dff_B_O1VL38gO8_2),.clk(gclk));
	jdff dff_B_0b5JWE0C3_2(.din(w_dff_B_O1VL38gO8_2),.dout(w_dff_B_0b5JWE0C3_2),.clk(gclk));
	jdff dff_B_JIkDY88H5_2(.din(w_dff_B_0b5JWE0C3_2),.dout(w_dff_B_JIkDY88H5_2),.clk(gclk));
	jdff dff_B_PgwT66Ft0_2(.din(w_dff_B_JIkDY88H5_2),.dout(w_dff_B_PgwT66Ft0_2),.clk(gclk));
	jdff dff_B_x1E0QGhx9_2(.din(w_dff_B_PgwT66Ft0_2),.dout(w_dff_B_x1E0QGhx9_2),.clk(gclk));
	jdff dff_B_ca5zKw4h8_2(.din(w_dff_B_x1E0QGhx9_2),.dout(w_dff_B_ca5zKw4h8_2),.clk(gclk));
	jdff dff_B_uzznCBdC5_2(.din(w_dff_B_ca5zKw4h8_2),.dout(w_dff_B_uzznCBdC5_2),.clk(gclk));
	jdff dff_B_pBLwVpBR3_2(.din(w_dff_B_uzznCBdC5_2),.dout(w_dff_B_pBLwVpBR3_2),.clk(gclk));
	jdff dff_B_2vBVMB5V7_2(.din(w_dff_B_pBLwVpBR3_2),.dout(w_dff_B_2vBVMB5V7_2),.clk(gclk));
	jdff dff_B_PAPhILIy3_2(.din(w_dff_B_2vBVMB5V7_2),.dout(w_dff_B_PAPhILIy3_2),.clk(gclk));
	jdff dff_B_WRwiQj2L4_2(.din(w_dff_B_PAPhILIy3_2),.dout(w_dff_B_WRwiQj2L4_2),.clk(gclk));
	jdff dff_B_EHldMUyZ4_2(.din(w_dff_B_WRwiQj2L4_2),.dout(w_dff_B_EHldMUyZ4_2),.clk(gclk));
	jdff dff_B_6pIPIOnR0_2(.din(w_dff_B_EHldMUyZ4_2),.dout(w_dff_B_6pIPIOnR0_2),.clk(gclk));
	jdff dff_B_xGLIlCo35_2(.din(w_dff_B_6pIPIOnR0_2),.dout(w_dff_B_xGLIlCo35_2),.clk(gclk));
	jdff dff_B_6SDlchVF5_2(.din(w_dff_B_xGLIlCo35_2),.dout(w_dff_B_6SDlchVF5_2),.clk(gclk));
	jdff dff_B_QVJawq5M1_2(.din(w_dff_B_6SDlchVF5_2),.dout(w_dff_B_QVJawq5M1_2),.clk(gclk));
	jdff dff_B_33JjJkgE1_2(.din(w_dff_B_QVJawq5M1_2),.dout(w_dff_B_33JjJkgE1_2),.clk(gclk));
	jdff dff_B_xYrxdJeJ8_2(.din(w_dff_B_33JjJkgE1_2),.dout(w_dff_B_xYrxdJeJ8_2),.clk(gclk));
	jdff dff_B_zlYVAhuQ2_2(.din(w_dff_B_xYrxdJeJ8_2),.dout(w_dff_B_zlYVAhuQ2_2),.clk(gclk));
	jdff dff_B_UdVcBu1Y2_2(.din(w_dff_B_zlYVAhuQ2_2),.dout(w_dff_B_UdVcBu1Y2_2),.clk(gclk));
	jdff dff_B_GSay1yMy4_2(.din(w_dff_B_UdVcBu1Y2_2),.dout(w_dff_B_GSay1yMy4_2),.clk(gclk));
	jdff dff_B_uJDcT60q3_2(.din(w_dff_B_GSay1yMy4_2),.dout(w_dff_B_uJDcT60q3_2),.clk(gclk));
	jdff dff_B_Vl3RO6UD6_2(.din(w_dff_B_uJDcT60q3_2),.dout(w_dff_B_Vl3RO6UD6_2),.clk(gclk));
	jdff dff_B_ic6kJmWQ0_2(.din(w_dff_B_Vl3RO6UD6_2),.dout(w_dff_B_ic6kJmWQ0_2),.clk(gclk));
	jdff dff_B_o3w5aTvI6_2(.din(w_dff_B_ic6kJmWQ0_2),.dout(w_dff_B_o3w5aTvI6_2),.clk(gclk));
	jdff dff_B_tS3OpCkK8_2(.din(w_dff_B_o3w5aTvI6_2),.dout(w_dff_B_tS3OpCkK8_2),.clk(gclk));
	jdff dff_B_JpaPDBvt5_2(.din(w_dff_B_tS3OpCkK8_2),.dout(w_dff_B_JpaPDBvt5_2),.clk(gclk));
	jdff dff_B_Io0C18lm3_2(.din(n1828),.dout(w_dff_B_Io0C18lm3_2),.clk(gclk));
	jdff dff_B_0JpSH0Ks5_2(.din(w_dff_B_Io0C18lm3_2),.dout(w_dff_B_0JpSH0Ks5_2),.clk(gclk));
	jdff dff_B_JcwB5xj55_2(.din(w_dff_B_0JpSH0Ks5_2),.dout(w_dff_B_JcwB5xj55_2),.clk(gclk));
	jdff dff_B_3XafXdoa3_2(.din(w_dff_B_JcwB5xj55_2),.dout(w_dff_B_3XafXdoa3_2),.clk(gclk));
	jdff dff_B_6eWBLgkO9_2(.din(w_dff_B_3XafXdoa3_2),.dout(w_dff_B_6eWBLgkO9_2),.clk(gclk));
	jdff dff_B_zwOG9EMm1_2(.din(w_dff_B_6eWBLgkO9_2),.dout(w_dff_B_zwOG9EMm1_2),.clk(gclk));
	jdff dff_B_fAMpavzh5_2(.din(w_dff_B_zwOG9EMm1_2),.dout(w_dff_B_fAMpavzh5_2),.clk(gclk));
	jdff dff_B_43CkqX3Q6_2(.din(w_dff_B_fAMpavzh5_2),.dout(w_dff_B_43CkqX3Q6_2),.clk(gclk));
	jdff dff_B_Oajl5QBZ0_2(.din(w_dff_B_43CkqX3Q6_2),.dout(w_dff_B_Oajl5QBZ0_2),.clk(gclk));
	jdff dff_B_XbSfiRoT2_2(.din(w_dff_B_Oajl5QBZ0_2),.dout(w_dff_B_XbSfiRoT2_2),.clk(gclk));
	jdff dff_B_2JzFZOws9_2(.din(w_dff_B_XbSfiRoT2_2),.dout(w_dff_B_2JzFZOws9_2),.clk(gclk));
	jdff dff_B_JUogRO798_2(.din(w_dff_B_2JzFZOws9_2),.dout(w_dff_B_JUogRO798_2),.clk(gclk));
	jdff dff_B_6BTKIP6a1_2(.din(w_dff_B_JUogRO798_2),.dout(w_dff_B_6BTKIP6a1_2),.clk(gclk));
	jdff dff_B_9QV78O5O7_2(.din(w_dff_B_6BTKIP6a1_2),.dout(w_dff_B_9QV78O5O7_2),.clk(gclk));
	jdff dff_B_UbrfE7eD8_2(.din(w_dff_B_9QV78O5O7_2),.dout(w_dff_B_UbrfE7eD8_2),.clk(gclk));
	jdff dff_B_PxKKlXrO1_2(.din(w_dff_B_UbrfE7eD8_2),.dout(w_dff_B_PxKKlXrO1_2),.clk(gclk));
	jdff dff_B_OBCWGu427_2(.din(w_dff_B_PxKKlXrO1_2),.dout(w_dff_B_OBCWGu427_2),.clk(gclk));
	jdff dff_B_Ftt84J4K6_2(.din(w_dff_B_OBCWGu427_2),.dout(w_dff_B_Ftt84J4K6_2),.clk(gclk));
	jdff dff_B_kXcQg8lf6_2(.din(w_dff_B_Ftt84J4K6_2),.dout(w_dff_B_kXcQg8lf6_2),.clk(gclk));
	jdff dff_B_g5fyCOod0_2(.din(w_dff_B_kXcQg8lf6_2),.dout(w_dff_B_g5fyCOod0_2),.clk(gclk));
	jdff dff_B_WAIpNcRT3_2(.din(w_dff_B_g5fyCOod0_2),.dout(w_dff_B_WAIpNcRT3_2),.clk(gclk));
	jdff dff_B_yGZJ0dbg3_2(.din(w_dff_B_WAIpNcRT3_2),.dout(w_dff_B_yGZJ0dbg3_2),.clk(gclk));
	jdff dff_B_5aPNFg957_2(.din(w_dff_B_yGZJ0dbg3_2),.dout(w_dff_B_5aPNFg957_2),.clk(gclk));
	jdff dff_B_UWkzjN9W7_2(.din(w_dff_B_5aPNFg957_2),.dout(w_dff_B_UWkzjN9W7_2),.clk(gclk));
	jdff dff_B_P8ozYtQT3_2(.din(w_dff_B_UWkzjN9W7_2),.dout(w_dff_B_P8ozYtQT3_2),.clk(gclk));
	jdff dff_B_EGpFVIuC6_2(.din(w_dff_B_P8ozYtQT3_2),.dout(w_dff_B_EGpFVIuC6_2),.clk(gclk));
	jdff dff_B_8sVdXMeF4_2(.din(w_dff_B_EGpFVIuC6_2),.dout(w_dff_B_8sVdXMeF4_2),.clk(gclk));
	jdff dff_B_mLXGekro9_2(.din(w_dff_B_8sVdXMeF4_2),.dout(w_dff_B_mLXGekro9_2),.clk(gclk));
	jdff dff_B_e0aBAl9o2_2(.din(w_dff_B_mLXGekro9_2),.dout(w_dff_B_e0aBAl9o2_2),.clk(gclk));
	jdff dff_B_xbANQquN3_2(.din(w_dff_B_e0aBAl9o2_2),.dout(w_dff_B_xbANQquN3_2),.clk(gclk));
	jdff dff_B_YwtbcyEk0_2(.din(w_dff_B_xbANQquN3_2),.dout(w_dff_B_YwtbcyEk0_2),.clk(gclk));
	jdff dff_B_ezY8Qn7m3_2(.din(w_dff_B_YwtbcyEk0_2),.dout(w_dff_B_ezY8Qn7m3_2),.clk(gclk));
	jdff dff_B_4hHymzK85_2(.din(w_dff_B_ezY8Qn7m3_2),.dout(w_dff_B_4hHymzK85_2),.clk(gclk));
	jdff dff_B_0FiXl07T4_2(.din(w_dff_B_4hHymzK85_2),.dout(w_dff_B_0FiXl07T4_2),.clk(gclk));
	jdff dff_B_gRthv1q88_2(.din(w_dff_B_0FiXl07T4_2),.dout(w_dff_B_gRthv1q88_2),.clk(gclk));
	jdff dff_B_zw7zxnwg9_2(.din(w_dff_B_gRthv1q88_2),.dout(w_dff_B_zw7zxnwg9_2),.clk(gclk));
	jdff dff_B_jxC1T4AV6_2(.din(w_dff_B_zw7zxnwg9_2),.dout(w_dff_B_jxC1T4AV6_2),.clk(gclk));
	jdff dff_B_E2dozOxm0_2(.din(w_dff_B_jxC1T4AV6_2),.dout(w_dff_B_E2dozOxm0_2),.clk(gclk));
	jdff dff_B_BSDbIl0Z8_2(.din(w_dff_B_E2dozOxm0_2),.dout(w_dff_B_BSDbIl0Z8_2),.clk(gclk));
	jdff dff_B_i3i2BuvJ5_2(.din(w_dff_B_BSDbIl0Z8_2),.dout(w_dff_B_i3i2BuvJ5_2),.clk(gclk));
	jdff dff_B_lqrZSR975_2(.din(w_dff_B_i3i2BuvJ5_2),.dout(w_dff_B_lqrZSR975_2),.clk(gclk));
	jdff dff_B_LDhrNUaG9_2(.din(w_dff_B_lqrZSR975_2),.dout(w_dff_B_LDhrNUaG9_2),.clk(gclk));
	jdff dff_B_vblGXDUh3_2(.din(w_dff_B_LDhrNUaG9_2),.dout(w_dff_B_vblGXDUh3_2),.clk(gclk));
	jdff dff_B_Vh7J7k9B3_2(.din(w_dff_B_vblGXDUh3_2),.dout(w_dff_B_Vh7J7k9B3_2),.clk(gclk));
	jdff dff_B_uGbOiL3U2_2(.din(w_dff_B_Vh7J7k9B3_2),.dout(w_dff_B_uGbOiL3U2_2),.clk(gclk));
	jdff dff_B_nTSBBC977_2(.din(w_dff_B_uGbOiL3U2_2),.dout(w_dff_B_nTSBBC977_2),.clk(gclk));
	jdff dff_B_DxOxGhbg6_2(.din(w_dff_B_nTSBBC977_2),.dout(w_dff_B_DxOxGhbg6_2),.clk(gclk));
	jdff dff_B_A9ejUpU21_2(.din(w_dff_B_DxOxGhbg6_2),.dout(w_dff_B_A9ejUpU21_2),.clk(gclk));
	jdff dff_B_w5EglXWf4_2(.din(w_dff_B_A9ejUpU21_2),.dout(w_dff_B_w5EglXWf4_2),.clk(gclk));
	jdff dff_B_yx5ZLr0Q9_2(.din(w_dff_B_w5EglXWf4_2),.dout(w_dff_B_yx5ZLr0Q9_2),.clk(gclk));
	jdff dff_B_S3CfbWQj4_2(.din(w_dff_B_yx5ZLr0Q9_2),.dout(w_dff_B_S3CfbWQj4_2),.clk(gclk));
	jdff dff_B_3NNnZg2w2_2(.din(w_dff_B_S3CfbWQj4_2),.dout(w_dff_B_3NNnZg2w2_2),.clk(gclk));
	jdff dff_B_p8UVPiSB4_2(.din(w_dff_B_3NNnZg2w2_2),.dout(w_dff_B_p8UVPiSB4_2),.clk(gclk));
	jdff dff_B_eEHRC27B2_2(.din(w_dff_B_p8UVPiSB4_2),.dout(w_dff_B_eEHRC27B2_2),.clk(gclk));
	jdff dff_B_mcyc9t8e2_2(.din(w_dff_B_eEHRC27B2_2),.dout(w_dff_B_mcyc9t8e2_2),.clk(gclk));
	jdff dff_B_HAS1H0Vi8_2(.din(w_dff_B_mcyc9t8e2_2),.dout(w_dff_B_HAS1H0Vi8_2),.clk(gclk));
	jdff dff_B_xBEtQaQ09_2(.din(w_dff_B_HAS1H0Vi8_2),.dout(w_dff_B_xBEtQaQ09_2),.clk(gclk));
	jdff dff_B_LrVQ6VMx0_2(.din(w_dff_B_xBEtQaQ09_2),.dout(w_dff_B_LrVQ6VMx0_2),.clk(gclk));
	jdff dff_A_PxkUvdjD5_1(.dout(w_n1827_0[1]),.din(w_dff_A_PxkUvdjD5_1),.clk(gclk));
	jdff dff_B_tNkfSlSJ7_1(.din(n1825),.dout(w_dff_B_tNkfSlSJ7_1),.clk(gclk));
	jdff dff_B_4dLvkYWc8_2(.din(n1803),.dout(w_dff_B_4dLvkYWc8_2),.clk(gclk));
	jdff dff_B_sLQsfsQl0_2(.din(w_dff_B_4dLvkYWc8_2),.dout(w_dff_B_sLQsfsQl0_2),.clk(gclk));
	jdff dff_B_oTplcCrl8_2(.din(w_dff_B_sLQsfsQl0_2),.dout(w_dff_B_oTplcCrl8_2),.clk(gclk));
	jdff dff_B_a6odMmZx5_2(.din(w_dff_B_oTplcCrl8_2),.dout(w_dff_B_a6odMmZx5_2),.clk(gclk));
	jdff dff_B_YUE9JYIw7_2(.din(w_dff_B_a6odMmZx5_2),.dout(w_dff_B_YUE9JYIw7_2),.clk(gclk));
	jdff dff_B_scrNy5P06_2(.din(w_dff_B_YUE9JYIw7_2),.dout(w_dff_B_scrNy5P06_2),.clk(gclk));
	jdff dff_B_I1FQNfmj5_2(.din(w_dff_B_scrNy5P06_2),.dout(w_dff_B_I1FQNfmj5_2),.clk(gclk));
	jdff dff_B_VmxyKjzi0_2(.din(w_dff_B_I1FQNfmj5_2),.dout(w_dff_B_VmxyKjzi0_2),.clk(gclk));
	jdff dff_B_fsLTpXFY3_2(.din(w_dff_B_VmxyKjzi0_2),.dout(w_dff_B_fsLTpXFY3_2),.clk(gclk));
	jdff dff_B_7ZwsPFYy8_2(.din(w_dff_B_fsLTpXFY3_2),.dout(w_dff_B_7ZwsPFYy8_2),.clk(gclk));
	jdff dff_B_qOoOHsiR9_2(.din(w_dff_B_7ZwsPFYy8_2),.dout(w_dff_B_qOoOHsiR9_2),.clk(gclk));
	jdff dff_B_BbupKVlH9_2(.din(w_dff_B_qOoOHsiR9_2),.dout(w_dff_B_BbupKVlH9_2),.clk(gclk));
	jdff dff_B_P1Ih1j6K5_2(.din(w_dff_B_BbupKVlH9_2),.dout(w_dff_B_P1Ih1j6K5_2),.clk(gclk));
	jdff dff_B_DgXScoMA0_2(.din(w_dff_B_P1Ih1j6K5_2),.dout(w_dff_B_DgXScoMA0_2),.clk(gclk));
	jdff dff_B_NmBS3vZW2_2(.din(w_dff_B_DgXScoMA0_2),.dout(w_dff_B_NmBS3vZW2_2),.clk(gclk));
	jdff dff_B_Q77MKcYK8_2(.din(w_dff_B_NmBS3vZW2_2),.dout(w_dff_B_Q77MKcYK8_2),.clk(gclk));
	jdff dff_B_WuHLpyfd9_2(.din(w_dff_B_Q77MKcYK8_2),.dout(w_dff_B_WuHLpyfd9_2),.clk(gclk));
	jdff dff_B_lo6BSgHR0_2(.din(w_dff_B_WuHLpyfd9_2),.dout(w_dff_B_lo6BSgHR0_2),.clk(gclk));
	jdff dff_B_HqPjGSw55_2(.din(w_dff_B_lo6BSgHR0_2),.dout(w_dff_B_HqPjGSw55_2),.clk(gclk));
	jdff dff_B_IYTCDilo3_2(.din(w_dff_B_HqPjGSw55_2),.dout(w_dff_B_IYTCDilo3_2),.clk(gclk));
	jdff dff_B_LJCdHRll0_2(.din(w_dff_B_IYTCDilo3_2),.dout(w_dff_B_LJCdHRll0_2),.clk(gclk));
	jdff dff_B_fZnb51im9_2(.din(w_dff_B_LJCdHRll0_2),.dout(w_dff_B_fZnb51im9_2),.clk(gclk));
	jdff dff_B_cs7d5pUm3_2(.din(w_dff_B_fZnb51im9_2),.dout(w_dff_B_cs7d5pUm3_2),.clk(gclk));
	jdff dff_B_kNTNVw497_2(.din(w_dff_B_cs7d5pUm3_2),.dout(w_dff_B_kNTNVw497_2),.clk(gclk));
	jdff dff_B_uVOH9iV53_2(.din(w_dff_B_kNTNVw497_2),.dout(w_dff_B_uVOH9iV53_2),.clk(gclk));
	jdff dff_B_pd8cr83u1_2(.din(w_dff_B_uVOH9iV53_2),.dout(w_dff_B_pd8cr83u1_2),.clk(gclk));
	jdff dff_B_x0ZdlwOg4_2(.din(w_dff_B_pd8cr83u1_2),.dout(w_dff_B_x0ZdlwOg4_2),.clk(gclk));
	jdff dff_B_dxU6Rwjq1_2(.din(w_dff_B_x0ZdlwOg4_2),.dout(w_dff_B_dxU6Rwjq1_2),.clk(gclk));
	jdff dff_B_0HHP96Ct3_2(.din(w_dff_B_dxU6Rwjq1_2),.dout(w_dff_B_0HHP96Ct3_2),.clk(gclk));
	jdff dff_B_FnpccuzM3_2(.din(w_dff_B_0HHP96Ct3_2),.dout(w_dff_B_FnpccuzM3_2),.clk(gclk));
	jdff dff_B_JYGUfNFJ6_2(.din(w_dff_B_FnpccuzM3_2),.dout(w_dff_B_JYGUfNFJ6_2),.clk(gclk));
	jdff dff_B_KQVbYU6k0_2(.din(w_dff_B_JYGUfNFJ6_2),.dout(w_dff_B_KQVbYU6k0_2),.clk(gclk));
	jdff dff_B_0avmNBE58_2(.din(w_dff_B_KQVbYU6k0_2),.dout(w_dff_B_0avmNBE58_2),.clk(gclk));
	jdff dff_B_tQU9bh5X8_2(.din(w_dff_B_0avmNBE58_2),.dout(w_dff_B_tQU9bh5X8_2),.clk(gclk));
	jdff dff_B_td7Gawrf0_2(.din(w_dff_B_tQU9bh5X8_2),.dout(w_dff_B_td7Gawrf0_2),.clk(gclk));
	jdff dff_B_BifjfJIz2_2(.din(w_dff_B_td7Gawrf0_2),.dout(w_dff_B_BifjfJIz2_2),.clk(gclk));
	jdff dff_B_LNtVcsYs7_2(.din(w_dff_B_BifjfJIz2_2),.dout(w_dff_B_LNtVcsYs7_2),.clk(gclk));
	jdff dff_B_JATmf3Qr5_2(.din(w_dff_B_LNtVcsYs7_2),.dout(w_dff_B_JATmf3Qr5_2),.clk(gclk));
	jdff dff_B_909Y0NrD1_2(.din(w_dff_B_JATmf3Qr5_2),.dout(w_dff_B_909Y0NrD1_2),.clk(gclk));
	jdff dff_B_DCHDFsZj8_2(.din(w_dff_B_909Y0NrD1_2),.dout(w_dff_B_DCHDFsZj8_2),.clk(gclk));
	jdff dff_B_0XEov4yd9_2(.din(w_dff_B_DCHDFsZj8_2),.dout(w_dff_B_0XEov4yd9_2),.clk(gclk));
	jdff dff_B_A0hF8aBU9_2(.din(w_dff_B_0XEov4yd9_2),.dout(w_dff_B_A0hF8aBU9_2),.clk(gclk));
	jdff dff_B_ksdZnOE90_2(.din(w_dff_B_A0hF8aBU9_2),.dout(w_dff_B_ksdZnOE90_2),.clk(gclk));
	jdff dff_B_47ZBgnGh9_2(.din(w_dff_B_ksdZnOE90_2),.dout(w_dff_B_47ZBgnGh9_2),.clk(gclk));
	jdff dff_B_Orxy2JUP1_2(.din(w_dff_B_47ZBgnGh9_2),.dout(w_dff_B_Orxy2JUP1_2),.clk(gclk));
	jdff dff_B_tJgmbYCk6_2(.din(w_dff_B_Orxy2JUP1_2),.dout(w_dff_B_tJgmbYCk6_2),.clk(gclk));
	jdff dff_B_dHAPEObs9_2(.din(w_dff_B_tJgmbYCk6_2),.dout(w_dff_B_dHAPEObs9_2),.clk(gclk));
	jdff dff_B_FQuRCi891_2(.din(w_dff_B_dHAPEObs9_2),.dout(w_dff_B_FQuRCi891_2),.clk(gclk));
	jdff dff_B_Y3F4Ii1O1_2(.din(w_dff_B_FQuRCi891_2),.dout(w_dff_B_Y3F4Ii1O1_2),.clk(gclk));
	jdff dff_B_t2O9zU334_2(.din(w_dff_B_Y3F4Ii1O1_2),.dout(w_dff_B_t2O9zU334_2),.clk(gclk));
	jdff dff_B_IfzgHusX8_2(.din(w_dff_B_t2O9zU334_2),.dout(w_dff_B_IfzgHusX8_2),.clk(gclk));
	jdff dff_B_GOI5AjxA5_2(.din(w_dff_B_IfzgHusX8_2),.dout(w_dff_B_GOI5AjxA5_2),.clk(gclk));
	jdff dff_B_BqzcS7iz9_2(.din(w_dff_B_GOI5AjxA5_2),.dout(w_dff_B_BqzcS7iz9_2),.clk(gclk));
	jdff dff_B_B12W2YLo8_2(.din(w_dff_B_BqzcS7iz9_2),.dout(w_dff_B_B12W2YLo8_2),.clk(gclk));
	jdff dff_B_BDl4KhBR6_2(.din(w_dff_B_B12W2YLo8_2),.dout(w_dff_B_BDl4KhBR6_2),.clk(gclk));
	jdff dff_B_sZ0n4Hta5_1(.din(n1809),.dout(w_dff_B_sZ0n4Hta5_1),.clk(gclk));
	jdff dff_B_4SA924Xj6_1(.din(w_dff_B_sZ0n4Hta5_1),.dout(w_dff_B_4SA924Xj6_1),.clk(gclk));
	jdff dff_B_pYtGxsg74_2(.din(n1808),.dout(w_dff_B_pYtGxsg74_2),.clk(gclk));
	jdff dff_B_6wcyaKks7_2(.din(w_dff_B_pYtGxsg74_2),.dout(w_dff_B_6wcyaKks7_2),.clk(gclk));
	jdff dff_B_tYVFheJu1_2(.din(w_dff_B_6wcyaKks7_2),.dout(w_dff_B_tYVFheJu1_2),.clk(gclk));
	jdff dff_B_ZXdJCphm5_2(.din(w_dff_B_tYVFheJu1_2),.dout(w_dff_B_ZXdJCphm5_2),.clk(gclk));
	jdff dff_B_SgtXfrKJ1_2(.din(w_dff_B_ZXdJCphm5_2),.dout(w_dff_B_SgtXfrKJ1_2),.clk(gclk));
	jdff dff_B_JUgGGi8m3_2(.din(w_dff_B_SgtXfrKJ1_2),.dout(w_dff_B_JUgGGi8m3_2),.clk(gclk));
	jdff dff_B_BWMXU5Od6_2(.din(w_dff_B_JUgGGi8m3_2),.dout(w_dff_B_BWMXU5Od6_2),.clk(gclk));
	jdff dff_B_gXZI6gMM4_2(.din(w_dff_B_BWMXU5Od6_2),.dout(w_dff_B_gXZI6gMM4_2),.clk(gclk));
	jdff dff_B_sqKFri9O2_2(.din(w_dff_B_gXZI6gMM4_2),.dout(w_dff_B_sqKFri9O2_2),.clk(gclk));
	jdff dff_B_KHD8PpI99_2(.din(w_dff_B_sqKFri9O2_2),.dout(w_dff_B_KHD8PpI99_2),.clk(gclk));
	jdff dff_B_D5HvEX1H6_2(.din(w_dff_B_KHD8PpI99_2),.dout(w_dff_B_D5HvEX1H6_2),.clk(gclk));
	jdff dff_B_1MsBVYxW1_2(.din(w_dff_B_D5HvEX1H6_2),.dout(w_dff_B_1MsBVYxW1_2),.clk(gclk));
	jdff dff_B_HP6jWg9P9_2(.din(w_dff_B_1MsBVYxW1_2),.dout(w_dff_B_HP6jWg9P9_2),.clk(gclk));
	jdff dff_B_OgEhbXF22_2(.din(w_dff_B_HP6jWg9P9_2),.dout(w_dff_B_OgEhbXF22_2),.clk(gclk));
	jdff dff_B_HGZZxS0u1_2(.din(w_dff_B_OgEhbXF22_2),.dout(w_dff_B_HGZZxS0u1_2),.clk(gclk));
	jdff dff_B_skp5RAy89_2(.din(w_dff_B_HGZZxS0u1_2),.dout(w_dff_B_skp5RAy89_2),.clk(gclk));
	jdff dff_B_AKnNt36s7_2(.din(w_dff_B_skp5RAy89_2),.dout(w_dff_B_AKnNt36s7_2),.clk(gclk));
	jdff dff_B_0TDGUQG90_2(.din(w_dff_B_AKnNt36s7_2),.dout(w_dff_B_0TDGUQG90_2),.clk(gclk));
	jdff dff_B_FCnxYKVA8_2(.din(w_dff_B_0TDGUQG90_2),.dout(w_dff_B_FCnxYKVA8_2),.clk(gclk));
	jdff dff_B_1o47LyxD5_2(.din(w_dff_B_FCnxYKVA8_2),.dout(w_dff_B_1o47LyxD5_2),.clk(gclk));
	jdff dff_B_KbJkTd8h5_2(.din(w_dff_B_1o47LyxD5_2),.dout(w_dff_B_KbJkTd8h5_2),.clk(gclk));
	jdff dff_B_gkWCoAB23_2(.din(w_dff_B_KbJkTd8h5_2),.dout(w_dff_B_gkWCoAB23_2),.clk(gclk));
	jdff dff_B_UQmXc7to0_2(.din(w_dff_B_gkWCoAB23_2),.dout(w_dff_B_UQmXc7to0_2),.clk(gclk));
	jdff dff_B_4UTup3KZ6_2(.din(w_dff_B_UQmXc7to0_2),.dout(w_dff_B_4UTup3KZ6_2),.clk(gclk));
	jdff dff_B_LhTZJTzn6_2(.din(w_dff_B_4UTup3KZ6_2),.dout(w_dff_B_LhTZJTzn6_2),.clk(gclk));
	jdff dff_B_4cS2J8M68_2(.din(w_dff_B_LhTZJTzn6_2),.dout(w_dff_B_4cS2J8M68_2),.clk(gclk));
	jdff dff_B_M6rGNXHB9_2(.din(w_dff_B_4cS2J8M68_2),.dout(w_dff_B_M6rGNXHB9_2),.clk(gclk));
	jdff dff_B_MGhtXBaN5_2(.din(w_dff_B_M6rGNXHB9_2),.dout(w_dff_B_MGhtXBaN5_2),.clk(gclk));
	jdff dff_B_68U2CJkr2_2(.din(w_dff_B_MGhtXBaN5_2),.dout(w_dff_B_68U2CJkr2_2),.clk(gclk));
	jdff dff_B_ufurvf7s9_2(.din(w_dff_B_68U2CJkr2_2),.dout(w_dff_B_ufurvf7s9_2),.clk(gclk));
	jdff dff_B_XZPkNmnU2_2(.din(w_dff_B_ufurvf7s9_2),.dout(w_dff_B_XZPkNmnU2_2),.clk(gclk));
	jdff dff_B_VCQI0V6X0_2(.din(w_dff_B_XZPkNmnU2_2),.dout(w_dff_B_VCQI0V6X0_2),.clk(gclk));
	jdff dff_B_ZKBNlK0a0_2(.din(w_dff_B_VCQI0V6X0_2),.dout(w_dff_B_ZKBNlK0a0_2),.clk(gclk));
	jdff dff_B_UYT9ceN93_2(.din(w_dff_B_ZKBNlK0a0_2),.dout(w_dff_B_UYT9ceN93_2),.clk(gclk));
	jdff dff_B_FMCpWyC84_2(.din(w_dff_B_UYT9ceN93_2),.dout(w_dff_B_FMCpWyC84_2),.clk(gclk));
	jdff dff_B_5Z13YJdr9_2(.din(w_dff_B_FMCpWyC84_2),.dout(w_dff_B_5Z13YJdr9_2),.clk(gclk));
	jdff dff_B_S1UFURAg6_2(.din(w_dff_B_5Z13YJdr9_2),.dout(w_dff_B_S1UFURAg6_2),.clk(gclk));
	jdff dff_B_pVaxPmDY7_2(.din(w_dff_B_S1UFURAg6_2),.dout(w_dff_B_pVaxPmDY7_2),.clk(gclk));
	jdff dff_B_ezxlfzdC5_2(.din(w_dff_B_pVaxPmDY7_2),.dout(w_dff_B_ezxlfzdC5_2),.clk(gclk));
	jdff dff_B_Rm2GF1Gd0_2(.din(w_dff_B_ezxlfzdC5_2),.dout(w_dff_B_Rm2GF1Gd0_2),.clk(gclk));
	jdff dff_B_q2uh49Nx8_2(.din(w_dff_B_Rm2GF1Gd0_2),.dout(w_dff_B_q2uh49Nx8_2),.clk(gclk));
	jdff dff_B_e6DDI9pT2_2(.din(w_dff_B_q2uh49Nx8_2),.dout(w_dff_B_e6DDI9pT2_2),.clk(gclk));
	jdff dff_B_90gFSyaO2_2(.din(w_dff_B_e6DDI9pT2_2),.dout(w_dff_B_90gFSyaO2_2),.clk(gclk));
	jdff dff_B_L8DhqAQa1_2(.din(w_dff_B_90gFSyaO2_2),.dout(w_dff_B_L8DhqAQa1_2),.clk(gclk));
	jdff dff_B_0THf7X6Y9_2(.din(w_dff_B_L8DhqAQa1_2),.dout(w_dff_B_0THf7X6Y9_2),.clk(gclk));
	jdff dff_B_CFuopNKt8_2(.din(w_dff_B_0THf7X6Y9_2),.dout(w_dff_B_CFuopNKt8_2),.clk(gclk));
	jdff dff_B_eRw48RmR9_2(.din(w_dff_B_CFuopNKt8_2),.dout(w_dff_B_eRw48RmR9_2),.clk(gclk));
	jdff dff_B_gY0Fu8SE1_2(.din(w_dff_B_eRw48RmR9_2),.dout(w_dff_B_gY0Fu8SE1_2),.clk(gclk));
	jdff dff_B_dcPATMxg5_2(.din(w_dff_B_gY0Fu8SE1_2),.dout(w_dff_B_dcPATMxg5_2),.clk(gclk));
	jdff dff_B_daCfm07m0_2(.din(w_dff_B_dcPATMxg5_2),.dout(w_dff_B_daCfm07m0_2),.clk(gclk));
	jdff dff_B_rgODx5oW3_2(.din(w_dff_B_daCfm07m0_2),.dout(w_dff_B_rgODx5oW3_2),.clk(gclk));
	jdff dff_B_liKzinUN3_2(.din(w_dff_B_rgODx5oW3_2),.dout(w_dff_B_liKzinUN3_2),.clk(gclk));
	jdff dff_B_BsaTgHYw4_2(.din(n1807),.dout(w_dff_B_BsaTgHYw4_2),.clk(gclk));
	jdff dff_B_t1O6oKSq9_2(.din(w_dff_B_BsaTgHYw4_2),.dout(w_dff_B_t1O6oKSq9_2),.clk(gclk));
	jdff dff_B_ffSl9Cab9_2(.din(w_dff_B_t1O6oKSq9_2),.dout(w_dff_B_ffSl9Cab9_2),.clk(gclk));
	jdff dff_B_rGwecK6y3_2(.din(w_dff_B_ffSl9Cab9_2),.dout(w_dff_B_rGwecK6y3_2),.clk(gclk));
	jdff dff_B_iePs9Un07_2(.din(w_dff_B_rGwecK6y3_2),.dout(w_dff_B_iePs9Un07_2),.clk(gclk));
	jdff dff_B_P7LeVSks1_2(.din(w_dff_B_iePs9Un07_2),.dout(w_dff_B_P7LeVSks1_2),.clk(gclk));
	jdff dff_B_X9bENC9z3_2(.din(w_dff_B_P7LeVSks1_2),.dout(w_dff_B_X9bENC9z3_2),.clk(gclk));
	jdff dff_B_Kpkcmpxd9_2(.din(w_dff_B_X9bENC9z3_2),.dout(w_dff_B_Kpkcmpxd9_2),.clk(gclk));
	jdff dff_B_f7Ms2toJ7_2(.din(w_dff_B_Kpkcmpxd9_2),.dout(w_dff_B_f7Ms2toJ7_2),.clk(gclk));
	jdff dff_B_9UUunrXK7_2(.din(w_dff_B_f7Ms2toJ7_2),.dout(w_dff_B_9UUunrXK7_2),.clk(gclk));
	jdff dff_B_1D2L7WHF8_2(.din(w_dff_B_9UUunrXK7_2),.dout(w_dff_B_1D2L7WHF8_2),.clk(gclk));
	jdff dff_B_xflbiNQm5_2(.din(w_dff_B_1D2L7WHF8_2),.dout(w_dff_B_xflbiNQm5_2),.clk(gclk));
	jdff dff_B_O8R6TIUu0_2(.din(w_dff_B_xflbiNQm5_2),.dout(w_dff_B_O8R6TIUu0_2),.clk(gclk));
	jdff dff_B_YyY3S8tN5_2(.din(w_dff_B_O8R6TIUu0_2),.dout(w_dff_B_YyY3S8tN5_2),.clk(gclk));
	jdff dff_B_tac62QeS5_2(.din(w_dff_B_YyY3S8tN5_2),.dout(w_dff_B_tac62QeS5_2),.clk(gclk));
	jdff dff_B_1ZNPkkAa9_2(.din(w_dff_B_tac62QeS5_2),.dout(w_dff_B_1ZNPkkAa9_2),.clk(gclk));
	jdff dff_B_mvwwcEob5_2(.din(w_dff_B_1ZNPkkAa9_2),.dout(w_dff_B_mvwwcEob5_2),.clk(gclk));
	jdff dff_B_XsPAtI5j4_2(.din(w_dff_B_mvwwcEob5_2),.dout(w_dff_B_XsPAtI5j4_2),.clk(gclk));
	jdff dff_B_ym3FaRK93_2(.din(w_dff_B_XsPAtI5j4_2),.dout(w_dff_B_ym3FaRK93_2),.clk(gclk));
	jdff dff_B_9VbxueTl5_2(.din(w_dff_B_ym3FaRK93_2),.dout(w_dff_B_9VbxueTl5_2),.clk(gclk));
	jdff dff_B_nxuuSiIL1_2(.din(w_dff_B_9VbxueTl5_2),.dout(w_dff_B_nxuuSiIL1_2),.clk(gclk));
	jdff dff_B_FaGLtmmB8_2(.din(w_dff_B_nxuuSiIL1_2),.dout(w_dff_B_FaGLtmmB8_2),.clk(gclk));
	jdff dff_B_ziSHAdvN8_2(.din(w_dff_B_FaGLtmmB8_2),.dout(w_dff_B_ziSHAdvN8_2),.clk(gclk));
	jdff dff_B_bvhQ0Iwp7_2(.din(w_dff_B_ziSHAdvN8_2),.dout(w_dff_B_bvhQ0Iwp7_2),.clk(gclk));
	jdff dff_B_uSY1jnWt4_2(.din(w_dff_B_bvhQ0Iwp7_2),.dout(w_dff_B_uSY1jnWt4_2),.clk(gclk));
	jdff dff_B_VHF6EVyl6_2(.din(w_dff_B_uSY1jnWt4_2),.dout(w_dff_B_VHF6EVyl6_2),.clk(gclk));
	jdff dff_B_npCI8OJT0_2(.din(w_dff_B_VHF6EVyl6_2),.dout(w_dff_B_npCI8OJT0_2),.clk(gclk));
	jdff dff_B_ag9mSPOG2_2(.din(w_dff_B_npCI8OJT0_2),.dout(w_dff_B_ag9mSPOG2_2),.clk(gclk));
	jdff dff_B_IrtbiRLW6_2(.din(w_dff_B_ag9mSPOG2_2),.dout(w_dff_B_IrtbiRLW6_2),.clk(gclk));
	jdff dff_B_ddDhfMnS6_2(.din(w_dff_B_IrtbiRLW6_2),.dout(w_dff_B_ddDhfMnS6_2),.clk(gclk));
	jdff dff_B_J5JQUBGL5_2(.din(w_dff_B_ddDhfMnS6_2),.dout(w_dff_B_J5JQUBGL5_2),.clk(gclk));
	jdff dff_B_502FbmUk1_2(.din(w_dff_B_J5JQUBGL5_2),.dout(w_dff_B_502FbmUk1_2),.clk(gclk));
	jdff dff_B_x3i6euFo9_2(.din(w_dff_B_502FbmUk1_2),.dout(w_dff_B_x3i6euFo9_2),.clk(gclk));
	jdff dff_B_7LY5gOsh0_2(.din(w_dff_B_x3i6euFo9_2),.dout(w_dff_B_7LY5gOsh0_2),.clk(gclk));
	jdff dff_B_pfohpeQA2_2(.din(w_dff_B_7LY5gOsh0_2),.dout(w_dff_B_pfohpeQA2_2),.clk(gclk));
	jdff dff_B_S3xA4Bdw5_2(.din(w_dff_B_pfohpeQA2_2),.dout(w_dff_B_S3xA4Bdw5_2),.clk(gclk));
	jdff dff_B_hanA9ou25_2(.din(w_dff_B_S3xA4Bdw5_2),.dout(w_dff_B_hanA9ou25_2),.clk(gclk));
	jdff dff_B_zTIxwpjW0_2(.din(w_dff_B_hanA9ou25_2),.dout(w_dff_B_zTIxwpjW0_2),.clk(gclk));
	jdff dff_B_rQbUJ0ru3_2(.din(w_dff_B_zTIxwpjW0_2),.dout(w_dff_B_rQbUJ0ru3_2),.clk(gclk));
	jdff dff_B_fwqoqcxC6_2(.din(w_dff_B_rQbUJ0ru3_2),.dout(w_dff_B_fwqoqcxC6_2),.clk(gclk));
	jdff dff_B_2EmyCWth1_2(.din(w_dff_B_fwqoqcxC6_2),.dout(w_dff_B_2EmyCWth1_2),.clk(gclk));
	jdff dff_B_ioHhMvB60_2(.din(w_dff_B_2EmyCWth1_2),.dout(w_dff_B_ioHhMvB60_2),.clk(gclk));
	jdff dff_B_qUrc4GBi7_2(.din(w_dff_B_ioHhMvB60_2),.dout(w_dff_B_qUrc4GBi7_2),.clk(gclk));
	jdff dff_B_ktSeaH7l9_2(.din(w_dff_B_qUrc4GBi7_2),.dout(w_dff_B_ktSeaH7l9_2),.clk(gclk));
	jdff dff_B_hQUK7uvr6_2(.din(w_dff_B_ktSeaH7l9_2),.dout(w_dff_B_hQUK7uvr6_2),.clk(gclk));
	jdff dff_B_OU9X3bAu4_2(.din(w_dff_B_hQUK7uvr6_2),.dout(w_dff_B_OU9X3bAu4_2),.clk(gclk));
	jdff dff_B_HMeGfbQN8_2(.din(w_dff_B_OU9X3bAu4_2),.dout(w_dff_B_HMeGfbQN8_2),.clk(gclk));
	jdff dff_B_Cjs9p1UA5_2(.din(w_dff_B_HMeGfbQN8_2),.dout(w_dff_B_Cjs9p1UA5_2),.clk(gclk));
	jdff dff_B_ZXGHL8ZM3_2(.din(w_dff_B_Cjs9p1UA5_2),.dout(w_dff_B_ZXGHL8ZM3_2),.clk(gclk));
	jdff dff_B_zlajOHoB8_2(.din(w_dff_B_ZXGHL8ZM3_2),.dout(w_dff_B_zlajOHoB8_2),.clk(gclk));
	jdff dff_B_ikPHQRGp4_2(.din(w_dff_B_zlajOHoB8_2),.dout(w_dff_B_ikPHQRGp4_2),.clk(gclk));
	jdff dff_B_6EMyCyQB3_2(.din(w_dff_B_ikPHQRGp4_2),.dout(w_dff_B_6EMyCyQB3_2),.clk(gclk));
	jdff dff_B_MKqAvzv91_2(.din(w_dff_B_6EMyCyQB3_2),.dout(w_dff_B_MKqAvzv91_2),.clk(gclk));
	jdff dff_B_cMF3AuPD1_2(.din(w_dff_B_MKqAvzv91_2),.dout(w_dff_B_cMF3AuPD1_2),.clk(gclk));
	jdff dff_B_MHVvfctY5_2(.din(n1806),.dout(w_dff_B_MHVvfctY5_2),.clk(gclk));
	jdff dff_B_F4FHKNsW0_1(.din(n1804),.dout(w_dff_B_F4FHKNsW0_1),.clk(gclk));
	jdff dff_B_7th5Eu8k8_2(.din(n1775),.dout(w_dff_B_7th5Eu8k8_2),.clk(gclk));
	jdff dff_B_eNtQf8L76_2(.din(w_dff_B_7th5Eu8k8_2),.dout(w_dff_B_eNtQf8L76_2),.clk(gclk));
	jdff dff_B_ezqvSYVZ6_2(.din(w_dff_B_eNtQf8L76_2),.dout(w_dff_B_ezqvSYVZ6_2),.clk(gclk));
	jdff dff_B_9fcBDFs02_2(.din(w_dff_B_ezqvSYVZ6_2),.dout(w_dff_B_9fcBDFs02_2),.clk(gclk));
	jdff dff_B_qsmmEwuc5_2(.din(w_dff_B_9fcBDFs02_2),.dout(w_dff_B_qsmmEwuc5_2),.clk(gclk));
	jdff dff_B_tfyTaVAS2_2(.din(w_dff_B_qsmmEwuc5_2),.dout(w_dff_B_tfyTaVAS2_2),.clk(gclk));
	jdff dff_B_zOb538h45_2(.din(w_dff_B_tfyTaVAS2_2),.dout(w_dff_B_zOb538h45_2),.clk(gclk));
	jdff dff_B_RJjmI3QK1_2(.din(w_dff_B_zOb538h45_2),.dout(w_dff_B_RJjmI3QK1_2),.clk(gclk));
	jdff dff_B_EYDSJ1sE8_2(.din(w_dff_B_RJjmI3QK1_2),.dout(w_dff_B_EYDSJ1sE8_2),.clk(gclk));
	jdff dff_B_DO0oLwq75_2(.din(w_dff_B_EYDSJ1sE8_2),.dout(w_dff_B_DO0oLwq75_2),.clk(gclk));
	jdff dff_B_CuyjJIYD9_2(.din(w_dff_B_DO0oLwq75_2),.dout(w_dff_B_CuyjJIYD9_2),.clk(gclk));
	jdff dff_B_6ozzNfPh4_2(.din(w_dff_B_CuyjJIYD9_2),.dout(w_dff_B_6ozzNfPh4_2),.clk(gclk));
	jdff dff_B_7YzEt90d8_2(.din(w_dff_B_6ozzNfPh4_2),.dout(w_dff_B_7YzEt90d8_2),.clk(gclk));
	jdff dff_B_Dxn49qfq0_2(.din(w_dff_B_7YzEt90d8_2),.dout(w_dff_B_Dxn49qfq0_2),.clk(gclk));
	jdff dff_B_5GdsDPw96_2(.din(w_dff_B_Dxn49qfq0_2),.dout(w_dff_B_5GdsDPw96_2),.clk(gclk));
	jdff dff_B_22QqtQ808_2(.din(w_dff_B_5GdsDPw96_2),.dout(w_dff_B_22QqtQ808_2),.clk(gclk));
	jdff dff_B_RqYL07YI1_2(.din(w_dff_B_22QqtQ808_2),.dout(w_dff_B_RqYL07YI1_2),.clk(gclk));
	jdff dff_B_aNcYWcOO0_2(.din(w_dff_B_RqYL07YI1_2),.dout(w_dff_B_aNcYWcOO0_2),.clk(gclk));
	jdff dff_B_MXDMfUh82_2(.din(w_dff_B_aNcYWcOO0_2),.dout(w_dff_B_MXDMfUh82_2),.clk(gclk));
	jdff dff_B_dj062R2L6_2(.din(w_dff_B_MXDMfUh82_2),.dout(w_dff_B_dj062R2L6_2),.clk(gclk));
	jdff dff_B_FMniWWpY4_2(.din(w_dff_B_dj062R2L6_2),.dout(w_dff_B_FMniWWpY4_2),.clk(gclk));
	jdff dff_B_gwBjsHvd8_2(.din(w_dff_B_FMniWWpY4_2),.dout(w_dff_B_gwBjsHvd8_2),.clk(gclk));
	jdff dff_B_8Js46k7n8_2(.din(w_dff_B_gwBjsHvd8_2),.dout(w_dff_B_8Js46k7n8_2),.clk(gclk));
	jdff dff_B_GxZMVNUd0_2(.din(w_dff_B_8Js46k7n8_2),.dout(w_dff_B_GxZMVNUd0_2),.clk(gclk));
	jdff dff_B_Y1jUCgmY4_2(.din(w_dff_B_GxZMVNUd0_2),.dout(w_dff_B_Y1jUCgmY4_2),.clk(gclk));
	jdff dff_B_VHOplYd21_2(.din(w_dff_B_Y1jUCgmY4_2),.dout(w_dff_B_VHOplYd21_2),.clk(gclk));
	jdff dff_B_sqHp7r664_2(.din(w_dff_B_VHOplYd21_2),.dout(w_dff_B_sqHp7r664_2),.clk(gclk));
	jdff dff_B_FJfdvBIf9_2(.din(w_dff_B_sqHp7r664_2),.dout(w_dff_B_FJfdvBIf9_2),.clk(gclk));
	jdff dff_B_DoIa5PwG1_2(.din(w_dff_B_FJfdvBIf9_2),.dout(w_dff_B_DoIa5PwG1_2),.clk(gclk));
	jdff dff_B_zN4Rv6WV8_2(.din(w_dff_B_DoIa5PwG1_2),.dout(w_dff_B_zN4Rv6WV8_2),.clk(gclk));
	jdff dff_B_CuONGkfX1_2(.din(w_dff_B_zN4Rv6WV8_2),.dout(w_dff_B_CuONGkfX1_2),.clk(gclk));
	jdff dff_B_cPwlPMfn0_2(.din(w_dff_B_CuONGkfX1_2),.dout(w_dff_B_cPwlPMfn0_2),.clk(gclk));
	jdff dff_B_cDJhrIkx9_2(.din(w_dff_B_cPwlPMfn0_2),.dout(w_dff_B_cDJhrIkx9_2),.clk(gclk));
	jdff dff_B_Iw2lApEp2_2(.din(w_dff_B_cDJhrIkx9_2),.dout(w_dff_B_Iw2lApEp2_2),.clk(gclk));
	jdff dff_B_Jz6mZXIg2_2(.din(w_dff_B_Iw2lApEp2_2),.dout(w_dff_B_Jz6mZXIg2_2),.clk(gclk));
	jdff dff_B_dXfV98yg9_2(.din(w_dff_B_Jz6mZXIg2_2),.dout(w_dff_B_dXfV98yg9_2),.clk(gclk));
	jdff dff_B_9KmcZ8cl8_2(.din(w_dff_B_dXfV98yg9_2),.dout(w_dff_B_9KmcZ8cl8_2),.clk(gclk));
	jdff dff_B_zbFxFGgO2_2(.din(w_dff_B_9KmcZ8cl8_2),.dout(w_dff_B_zbFxFGgO2_2),.clk(gclk));
	jdff dff_B_vO8nQTRu6_2(.din(w_dff_B_zbFxFGgO2_2),.dout(w_dff_B_vO8nQTRu6_2),.clk(gclk));
	jdff dff_B_hsKuwM0e2_2(.din(w_dff_B_vO8nQTRu6_2),.dout(w_dff_B_hsKuwM0e2_2),.clk(gclk));
	jdff dff_B_O796C1Mu8_2(.din(w_dff_B_hsKuwM0e2_2),.dout(w_dff_B_O796C1Mu8_2),.clk(gclk));
	jdff dff_B_UClX28LH5_2(.din(w_dff_B_O796C1Mu8_2),.dout(w_dff_B_UClX28LH5_2),.clk(gclk));
	jdff dff_B_nldJQdoc6_2(.din(w_dff_B_UClX28LH5_2),.dout(w_dff_B_nldJQdoc6_2),.clk(gclk));
	jdff dff_B_6XfxOawj1_2(.din(w_dff_B_nldJQdoc6_2),.dout(w_dff_B_6XfxOawj1_2),.clk(gclk));
	jdff dff_B_BtpAo8wy3_2(.din(w_dff_B_6XfxOawj1_2),.dout(w_dff_B_BtpAo8wy3_2),.clk(gclk));
	jdff dff_B_8tKzbF3I9_2(.din(w_dff_B_BtpAo8wy3_2),.dout(w_dff_B_8tKzbF3I9_2),.clk(gclk));
	jdff dff_B_3KXoA0oy1_2(.din(w_dff_B_8tKzbF3I9_2),.dout(w_dff_B_3KXoA0oy1_2),.clk(gclk));
	jdff dff_B_6wMB7NcD8_2(.din(w_dff_B_3KXoA0oy1_2),.dout(w_dff_B_6wMB7NcD8_2),.clk(gclk));
	jdff dff_B_jmGBCNw90_2(.din(w_dff_B_6wMB7NcD8_2),.dout(w_dff_B_jmGBCNw90_2),.clk(gclk));
	jdff dff_B_PSwzMt0B0_2(.din(w_dff_B_jmGBCNw90_2),.dout(w_dff_B_PSwzMt0B0_2),.clk(gclk));
	jdff dff_B_D4NOgbEQ5_2(.din(w_dff_B_PSwzMt0B0_2),.dout(w_dff_B_D4NOgbEQ5_2),.clk(gclk));
	jdff dff_B_oYaDfUxp0_1(.din(n1781),.dout(w_dff_B_oYaDfUxp0_1),.clk(gclk));
	jdff dff_B_Zw6pdW2B7_1(.din(w_dff_B_oYaDfUxp0_1),.dout(w_dff_B_Zw6pdW2B7_1),.clk(gclk));
	jdff dff_B_OV4LUR9w6_2(.din(n1780),.dout(w_dff_B_OV4LUR9w6_2),.clk(gclk));
	jdff dff_B_7xVEc9Hf6_2(.din(w_dff_B_OV4LUR9w6_2),.dout(w_dff_B_7xVEc9Hf6_2),.clk(gclk));
	jdff dff_B_9zawBzxn9_2(.din(w_dff_B_7xVEc9Hf6_2),.dout(w_dff_B_9zawBzxn9_2),.clk(gclk));
	jdff dff_B_MieYUYhc0_2(.din(w_dff_B_9zawBzxn9_2),.dout(w_dff_B_MieYUYhc0_2),.clk(gclk));
	jdff dff_B_z5ZvKtdP1_2(.din(w_dff_B_MieYUYhc0_2),.dout(w_dff_B_z5ZvKtdP1_2),.clk(gclk));
	jdff dff_B_B1iToAsH0_2(.din(w_dff_B_z5ZvKtdP1_2),.dout(w_dff_B_B1iToAsH0_2),.clk(gclk));
	jdff dff_B_5gUBTiEV8_2(.din(w_dff_B_B1iToAsH0_2),.dout(w_dff_B_5gUBTiEV8_2),.clk(gclk));
	jdff dff_B_OuEIFy7O2_2(.din(w_dff_B_5gUBTiEV8_2),.dout(w_dff_B_OuEIFy7O2_2),.clk(gclk));
	jdff dff_B_Zm7Vb1ab6_2(.din(w_dff_B_OuEIFy7O2_2),.dout(w_dff_B_Zm7Vb1ab6_2),.clk(gclk));
	jdff dff_B_GOhfNCV89_2(.din(w_dff_B_Zm7Vb1ab6_2),.dout(w_dff_B_GOhfNCV89_2),.clk(gclk));
	jdff dff_B_IRBZdozG4_2(.din(w_dff_B_GOhfNCV89_2),.dout(w_dff_B_IRBZdozG4_2),.clk(gclk));
	jdff dff_B_yN02whnS4_2(.din(w_dff_B_IRBZdozG4_2),.dout(w_dff_B_yN02whnS4_2),.clk(gclk));
	jdff dff_B_RHotYsHB3_2(.din(w_dff_B_yN02whnS4_2),.dout(w_dff_B_RHotYsHB3_2),.clk(gclk));
	jdff dff_B_aiTtJlBd0_2(.din(w_dff_B_RHotYsHB3_2),.dout(w_dff_B_aiTtJlBd0_2),.clk(gclk));
	jdff dff_B_30NKNu9z1_2(.din(w_dff_B_aiTtJlBd0_2),.dout(w_dff_B_30NKNu9z1_2),.clk(gclk));
	jdff dff_B_J9XBmAWz3_2(.din(w_dff_B_30NKNu9z1_2),.dout(w_dff_B_J9XBmAWz3_2),.clk(gclk));
	jdff dff_B_KRdQabDh0_2(.din(w_dff_B_J9XBmAWz3_2),.dout(w_dff_B_KRdQabDh0_2),.clk(gclk));
	jdff dff_B_8xt4TcaS7_2(.din(w_dff_B_KRdQabDh0_2),.dout(w_dff_B_8xt4TcaS7_2),.clk(gclk));
	jdff dff_B_DdQebRkn8_2(.din(w_dff_B_8xt4TcaS7_2),.dout(w_dff_B_DdQebRkn8_2),.clk(gclk));
	jdff dff_B_5ndfVFLi2_2(.din(w_dff_B_DdQebRkn8_2),.dout(w_dff_B_5ndfVFLi2_2),.clk(gclk));
	jdff dff_B_EJRUeUsm9_2(.din(w_dff_B_5ndfVFLi2_2),.dout(w_dff_B_EJRUeUsm9_2),.clk(gclk));
	jdff dff_B_Rsr9SgWK7_2(.din(w_dff_B_EJRUeUsm9_2),.dout(w_dff_B_Rsr9SgWK7_2),.clk(gclk));
	jdff dff_B_UgIiy5Kt6_2(.din(w_dff_B_Rsr9SgWK7_2),.dout(w_dff_B_UgIiy5Kt6_2),.clk(gclk));
	jdff dff_B_CU6wx5aF5_2(.din(w_dff_B_UgIiy5Kt6_2),.dout(w_dff_B_CU6wx5aF5_2),.clk(gclk));
	jdff dff_B_bCX4Ajy76_2(.din(w_dff_B_CU6wx5aF5_2),.dout(w_dff_B_bCX4Ajy76_2),.clk(gclk));
	jdff dff_B_TMm5lXh39_2(.din(w_dff_B_bCX4Ajy76_2),.dout(w_dff_B_TMm5lXh39_2),.clk(gclk));
	jdff dff_B_hrHhPy0U8_2(.din(w_dff_B_TMm5lXh39_2),.dout(w_dff_B_hrHhPy0U8_2),.clk(gclk));
	jdff dff_B_VlUjF8JE3_2(.din(w_dff_B_hrHhPy0U8_2),.dout(w_dff_B_VlUjF8JE3_2),.clk(gclk));
	jdff dff_B_PG7edLz47_2(.din(w_dff_B_VlUjF8JE3_2),.dout(w_dff_B_PG7edLz47_2),.clk(gclk));
	jdff dff_B_YeZoBVpI3_2(.din(w_dff_B_PG7edLz47_2),.dout(w_dff_B_YeZoBVpI3_2),.clk(gclk));
	jdff dff_B_2vuAxxcz5_2(.din(w_dff_B_YeZoBVpI3_2),.dout(w_dff_B_2vuAxxcz5_2),.clk(gclk));
	jdff dff_B_Zo7pIShD4_2(.din(w_dff_B_2vuAxxcz5_2),.dout(w_dff_B_Zo7pIShD4_2),.clk(gclk));
	jdff dff_B_YM1UwXZe3_2(.din(w_dff_B_Zo7pIShD4_2),.dout(w_dff_B_YM1UwXZe3_2),.clk(gclk));
	jdff dff_B_XHW13VCe7_2(.din(w_dff_B_YM1UwXZe3_2),.dout(w_dff_B_XHW13VCe7_2),.clk(gclk));
	jdff dff_B_O3ViLOwi6_2(.din(w_dff_B_XHW13VCe7_2),.dout(w_dff_B_O3ViLOwi6_2),.clk(gclk));
	jdff dff_B_ZJrLVXEH9_2(.din(w_dff_B_O3ViLOwi6_2),.dout(w_dff_B_ZJrLVXEH9_2),.clk(gclk));
	jdff dff_B_dwrjPAOO5_2(.din(w_dff_B_ZJrLVXEH9_2),.dout(w_dff_B_dwrjPAOO5_2),.clk(gclk));
	jdff dff_B_KcxmlSch9_2(.din(w_dff_B_dwrjPAOO5_2),.dout(w_dff_B_KcxmlSch9_2),.clk(gclk));
	jdff dff_B_PnhtiqsM1_2(.din(w_dff_B_KcxmlSch9_2),.dout(w_dff_B_PnhtiqsM1_2),.clk(gclk));
	jdff dff_B_AXtIdQhT6_2(.din(w_dff_B_PnhtiqsM1_2),.dout(w_dff_B_AXtIdQhT6_2),.clk(gclk));
	jdff dff_B_xWAgze7w9_2(.din(w_dff_B_AXtIdQhT6_2),.dout(w_dff_B_xWAgze7w9_2),.clk(gclk));
	jdff dff_B_ZJAz3KHS8_2(.din(w_dff_B_xWAgze7w9_2),.dout(w_dff_B_ZJAz3KHS8_2),.clk(gclk));
	jdff dff_B_e0XZZnYI7_2(.din(w_dff_B_ZJAz3KHS8_2),.dout(w_dff_B_e0XZZnYI7_2),.clk(gclk));
	jdff dff_B_zLltfwQ73_2(.din(w_dff_B_e0XZZnYI7_2),.dout(w_dff_B_zLltfwQ73_2),.clk(gclk));
	jdff dff_B_BqDVFM0I9_2(.din(w_dff_B_zLltfwQ73_2),.dout(w_dff_B_BqDVFM0I9_2),.clk(gclk));
	jdff dff_B_YB20j6aj7_2(.din(w_dff_B_BqDVFM0I9_2),.dout(w_dff_B_YB20j6aj7_2),.clk(gclk));
	jdff dff_B_pAwqq2H84_2(.din(w_dff_B_YB20j6aj7_2),.dout(w_dff_B_pAwqq2H84_2),.clk(gclk));
	jdff dff_B_Pk8E9oz23_2(.din(w_dff_B_pAwqq2H84_2),.dout(w_dff_B_Pk8E9oz23_2),.clk(gclk));
	jdff dff_B_JbmMvYa28_2(.din(n1779),.dout(w_dff_B_JbmMvYa28_2),.clk(gclk));
	jdff dff_B_HLYmbXXu4_2(.din(w_dff_B_JbmMvYa28_2),.dout(w_dff_B_HLYmbXXu4_2),.clk(gclk));
	jdff dff_B_Bbe2et671_2(.din(w_dff_B_HLYmbXXu4_2),.dout(w_dff_B_Bbe2et671_2),.clk(gclk));
	jdff dff_B_MP2LU5qv2_2(.din(w_dff_B_Bbe2et671_2),.dout(w_dff_B_MP2LU5qv2_2),.clk(gclk));
	jdff dff_B_bPL2csOe3_2(.din(w_dff_B_MP2LU5qv2_2),.dout(w_dff_B_bPL2csOe3_2),.clk(gclk));
	jdff dff_B_KvEjsbWD6_2(.din(w_dff_B_bPL2csOe3_2),.dout(w_dff_B_KvEjsbWD6_2),.clk(gclk));
	jdff dff_B_YUhrlVBC6_2(.din(w_dff_B_KvEjsbWD6_2),.dout(w_dff_B_YUhrlVBC6_2),.clk(gclk));
	jdff dff_B_jOefrOrM7_2(.din(w_dff_B_YUhrlVBC6_2),.dout(w_dff_B_jOefrOrM7_2),.clk(gclk));
	jdff dff_B_9d3OhIBC0_2(.din(w_dff_B_jOefrOrM7_2),.dout(w_dff_B_9d3OhIBC0_2),.clk(gclk));
	jdff dff_B_eKpd4oYH6_2(.din(w_dff_B_9d3OhIBC0_2),.dout(w_dff_B_eKpd4oYH6_2),.clk(gclk));
	jdff dff_B_080ijP9M4_2(.din(w_dff_B_eKpd4oYH6_2),.dout(w_dff_B_080ijP9M4_2),.clk(gclk));
	jdff dff_B_yCaNAeC87_2(.din(w_dff_B_080ijP9M4_2),.dout(w_dff_B_yCaNAeC87_2),.clk(gclk));
	jdff dff_B_bKPjXg5E8_2(.din(w_dff_B_yCaNAeC87_2),.dout(w_dff_B_bKPjXg5E8_2),.clk(gclk));
	jdff dff_B_F7Cnun5r4_2(.din(w_dff_B_bKPjXg5E8_2),.dout(w_dff_B_F7Cnun5r4_2),.clk(gclk));
	jdff dff_B_yKzMgUDd6_2(.din(w_dff_B_F7Cnun5r4_2),.dout(w_dff_B_yKzMgUDd6_2),.clk(gclk));
	jdff dff_B_fkr5epSt1_2(.din(w_dff_B_yKzMgUDd6_2),.dout(w_dff_B_fkr5epSt1_2),.clk(gclk));
	jdff dff_B_pEXQ0zAK8_2(.din(w_dff_B_fkr5epSt1_2),.dout(w_dff_B_pEXQ0zAK8_2),.clk(gclk));
	jdff dff_B_DdwJof3h4_2(.din(w_dff_B_pEXQ0zAK8_2),.dout(w_dff_B_DdwJof3h4_2),.clk(gclk));
	jdff dff_B_Ry7Emped2_2(.din(w_dff_B_DdwJof3h4_2),.dout(w_dff_B_Ry7Emped2_2),.clk(gclk));
	jdff dff_B_ZvyBeOMc0_2(.din(w_dff_B_Ry7Emped2_2),.dout(w_dff_B_ZvyBeOMc0_2),.clk(gclk));
	jdff dff_B_er71KSAg2_2(.din(w_dff_B_ZvyBeOMc0_2),.dout(w_dff_B_er71KSAg2_2),.clk(gclk));
	jdff dff_B_TU1ZtA7S9_2(.din(w_dff_B_er71KSAg2_2),.dout(w_dff_B_TU1ZtA7S9_2),.clk(gclk));
	jdff dff_B_TTQ0rCYZ5_2(.din(w_dff_B_TU1ZtA7S9_2),.dout(w_dff_B_TTQ0rCYZ5_2),.clk(gclk));
	jdff dff_B_eq8TzAIK3_2(.din(w_dff_B_TTQ0rCYZ5_2),.dout(w_dff_B_eq8TzAIK3_2),.clk(gclk));
	jdff dff_B_wg6UR4za2_2(.din(w_dff_B_eq8TzAIK3_2),.dout(w_dff_B_wg6UR4za2_2),.clk(gclk));
	jdff dff_B_ovCrJYmZ1_2(.din(w_dff_B_wg6UR4za2_2),.dout(w_dff_B_ovCrJYmZ1_2),.clk(gclk));
	jdff dff_B_uXlVHjDb6_2(.din(w_dff_B_ovCrJYmZ1_2),.dout(w_dff_B_uXlVHjDb6_2),.clk(gclk));
	jdff dff_B_A8I7fDO20_2(.din(w_dff_B_uXlVHjDb6_2),.dout(w_dff_B_A8I7fDO20_2),.clk(gclk));
	jdff dff_B_iNxsZu442_2(.din(w_dff_B_A8I7fDO20_2),.dout(w_dff_B_iNxsZu442_2),.clk(gclk));
	jdff dff_B_U8TTNHZv1_2(.din(w_dff_B_iNxsZu442_2),.dout(w_dff_B_U8TTNHZv1_2),.clk(gclk));
	jdff dff_B_JjzevDjA3_2(.din(w_dff_B_U8TTNHZv1_2),.dout(w_dff_B_JjzevDjA3_2),.clk(gclk));
	jdff dff_B_LdtPjObD7_2(.din(w_dff_B_JjzevDjA3_2),.dout(w_dff_B_LdtPjObD7_2),.clk(gclk));
	jdff dff_B_aNEvkxOt6_2(.din(w_dff_B_LdtPjObD7_2),.dout(w_dff_B_aNEvkxOt6_2),.clk(gclk));
	jdff dff_B_cGjC7Z618_2(.din(w_dff_B_aNEvkxOt6_2),.dout(w_dff_B_cGjC7Z618_2),.clk(gclk));
	jdff dff_B_05Ha8Hq07_2(.din(w_dff_B_cGjC7Z618_2),.dout(w_dff_B_05Ha8Hq07_2),.clk(gclk));
	jdff dff_B_JBoKDsAG6_2(.din(w_dff_B_05Ha8Hq07_2),.dout(w_dff_B_JBoKDsAG6_2),.clk(gclk));
	jdff dff_B_5LjpxmwP3_2(.din(w_dff_B_JBoKDsAG6_2),.dout(w_dff_B_5LjpxmwP3_2),.clk(gclk));
	jdff dff_B_TeoLBedL4_2(.din(w_dff_B_5LjpxmwP3_2),.dout(w_dff_B_TeoLBedL4_2),.clk(gclk));
	jdff dff_B_owtTLooF9_2(.din(w_dff_B_TeoLBedL4_2),.dout(w_dff_B_owtTLooF9_2),.clk(gclk));
	jdff dff_B_m1RR29ev5_2(.din(w_dff_B_owtTLooF9_2),.dout(w_dff_B_m1RR29ev5_2),.clk(gclk));
	jdff dff_B_21nNhFmo1_2(.din(w_dff_B_m1RR29ev5_2),.dout(w_dff_B_21nNhFmo1_2),.clk(gclk));
	jdff dff_B_VCGXyKEd7_2(.din(w_dff_B_21nNhFmo1_2),.dout(w_dff_B_VCGXyKEd7_2),.clk(gclk));
	jdff dff_B_kljDPrGO5_2(.din(w_dff_B_VCGXyKEd7_2),.dout(w_dff_B_kljDPrGO5_2),.clk(gclk));
	jdff dff_B_Ug5oEP0f3_2(.din(w_dff_B_kljDPrGO5_2),.dout(w_dff_B_Ug5oEP0f3_2),.clk(gclk));
	jdff dff_B_RESDTSlx4_2(.din(w_dff_B_Ug5oEP0f3_2),.dout(w_dff_B_RESDTSlx4_2),.clk(gclk));
	jdff dff_B_I8mhd0fK9_2(.din(w_dff_B_RESDTSlx4_2),.dout(w_dff_B_I8mhd0fK9_2),.clk(gclk));
	jdff dff_B_IXvPLQhX8_2(.din(w_dff_B_I8mhd0fK9_2),.dout(w_dff_B_IXvPLQhX8_2),.clk(gclk));
	jdff dff_B_KvOeL6FU1_2(.din(w_dff_B_IXvPLQhX8_2),.dout(w_dff_B_KvOeL6FU1_2),.clk(gclk));
	jdff dff_B_BG45Licz8_2(.din(w_dff_B_KvOeL6FU1_2),.dout(w_dff_B_BG45Licz8_2),.clk(gclk));
	jdff dff_B_BBmT6JTF2_2(.din(w_dff_B_BG45Licz8_2),.dout(w_dff_B_BBmT6JTF2_2),.clk(gclk));
	jdff dff_B_nodTVjh30_2(.din(n1778),.dout(w_dff_B_nodTVjh30_2),.clk(gclk));
	jdff dff_B_L2SDGRk72_1(.din(n1776),.dout(w_dff_B_L2SDGRk72_1),.clk(gclk));
	jdff dff_B_ZWkI9xn98_2(.din(n1740),.dout(w_dff_B_ZWkI9xn98_2),.clk(gclk));
	jdff dff_B_RvkAJ08B5_2(.din(w_dff_B_ZWkI9xn98_2),.dout(w_dff_B_RvkAJ08B5_2),.clk(gclk));
	jdff dff_B_VeZ4sR612_2(.din(w_dff_B_RvkAJ08B5_2),.dout(w_dff_B_VeZ4sR612_2),.clk(gclk));
	jdff dff_B_T4b7XMC90_2(.din(w_dff_B_VeZ4sR612_2),.dout(w_dff_B_T4b7XMC90_2),.clk(gclk));
	jdff dff_B_ZTQaUEub6_2(.din(w_dff_B_T4b7XMC90_2),.dout(w_dff_B_ZTQaUEub6_2),.clk(gclk));
	jdff dff_B_0ujpAZ0z9_2(.din(w_dff_B_ZTQaUEub6_2),.dout(w_dff_B_0ujpAZ0z9_2),.clk(gclk));
	jdff dff_B_SL921Pt80_2(.din(w_dff_B_0ujpAZ0z9_2),.dout(w_dff_B_SL921Pt80_2),.clk(gclk));
	jdff dff_B_Bg7uuIgI8_2(.din(w_dff_B_SL921Pt80_2),.dout(w_dff_B_Bg7uuIgI8_2),.clk(gclk));
	jdff dff_B_Iv1CUzmx8_2(.din(w_dff_B_Bg7uuIgI8_2),.dout(w_dff_B_Iv1CUzmx8_2),.clk(gclk));
	jdff dff_B_yPcKFBWT3_2(.din(w_dff_B_Iv1CUzmx8_2),.dout(w_dff_B_yPcKFBWT3_2),.clk(gclk));
	jdff dff_B_kUBVjpyw2_2(.din(w_dff_B_yPcKFBWT3_2),.dout(w_dff_B_kUBVjpyw2_2),.clk(gclk));
	jdff dff_B_c5rXOnPh5_2(.din(w_dff_B_kUBVjpyw2_2),.dout(w_dff_B_c5rXOnPh5_2),.clk(gclk));
	jdff dff_B_y2X4KWtG6_2(.din(w_dff_B_c5rXOnPh5_2),.dout(w_dff_B_y2X4KWtG6_2),.clk(gclk));
	jdff dff_B_qap6YxH67_2(.din(w_dff_B_y2X4KWtG6_2),.dout(w_dff_B_qap6YxH67_2),.clk(gclk));
	jdff dff_B_dkeqJFbi4_2(.din(w_dff_B_qap6YxH67_2),.dout(w_dff_B_dkeqJFbi4_2),.clk(gclk));
	jdff dff_B_iCjWJ5809_2(.din(w_dff_B_dkeqJFbi4_2),.dout(w_dff_B_iCjWJ5809_2),.clk(gclk));
	jdff dff_B_0ahnppPY8_2(.din(w_dff_B_iCjWJ5809_2),.dout(w_dff_B_0ahnppPY8_2),.clk(gclk));
	jdff dff_B_mhG9EiKt7_2(.din(w_dff_B_0ahnppPY8_2),.dout(w_dff_B_mhG9EiKt7_2),.clk(gclk));
	jdff dff_B_ourMqqw07_2(.din(w_dff_B_mhG9EiKt7_2),.dout(w_dff_B_ourMqqw07_2),.clk(gclk));
	jdff dff_B_1jzBeIjY9_2(.din(w_dff_B_ourMqqw07_2),.dout(w_dff_B_1jzBeIjY9_2),.clk(gclk));
	jdff dff_B_BuZnoyKm4_2(.din(w_dff_B_1jzBeIjY9_2),.dout(w_dff_B_BuZnoyKm4_2),.clk(gclk));
	jdff dff_B_xR8vUvqk4_2(.din(w_dff_B_BuZnoyKm4_2),.dout(w_dff_B_xR8vUvqk4_2),.clk(gclk));
	jdff dff_B_ZxSQhSYP7_2(.din(w_dff_B_xR8vUvqk4_2),.dout(w_dff_B_ZxSQhSYP7_2),.clk(gclk));
	jdff dff_B_0b1WvJfR3_2(.din(w_dff_B_ZxSQhSYP7_2),.dout(w_dff_B_0b1WvJfR3_2),.clk(gclk));
	jdff dff_B_ogytpNaq0_2(.din(w_dff_B_0b1WvJfR3_2),.dout(w_dff_B_ogytpNaq0_2),.clk(gclk));
	jdff dff_B_Jv6k8U4S0_2(.din(w_dff_B_ogytpNaq0_2),.dout(w_dff_B_Jv6k8U4S0_2),.clk(gclk));
	jdff dff_B_iYbHOVF81_2(.din(w_dff_B_Jv6k8U4S0_2),.dout(w_dff_B_iYbHOVF81_2),.clk(gclk));
	jdff dff_B_mNivilHR3_2(.din(w_dff_B_iYbHOVF81_2),.dout(w_dff_B_mNivilHR3_2),.clk(gclk));
	jdff dff_B_3Bxzm1gu5_2(.din(w_dff_B_mNivilHR3_2),.dout(w_dff_B_3Bxzm1gu5_2),.clk(gclk));
	jdff dff_B_PNOtDNoa6_2(.din(w_dff_B_3Bxzm1gu5_2),.dout(w_dff_B_PNOtDNoa6_2),.clk(gclk));
	jdff dff_B_V2T9ES6U0_2(.din(w_dff_B_PNOtDNoa6_2),.dout(w_dff_B_V2T9ES6U0_2),.clk(gclk));
	jdff dff_B_DxUyRIN37_2(.din(w_dff_B_V2T9ES6U0_2),.dout(w_dff_B_DxUyRIN37_2),.clk(gclk));
	jdff dff_B_suJtMlCG3_2(.din(w_dff_B_DxUyRIN37_2),.dout(w_dff_B_suJtMlCG3_2),.clk(gclk));
	jdff dff_B_uvYZZWps6_2(.din(w_dff_B_suJtMlCG3_2),.dout(w_dff_B_uvYZZWps6_2),.clk(gclk));
	jdff dff_B_jOBpItFi5_2(.din(w_dff_B_uvYZZWps6_2),.dout(w_dff_B_jOBpItFi5_2),.clk(gclk));
	jdff dff_B_pFtKX6H66_2(.din(w_dff_B_jOBpItFi5_2),.dout(w_dff_B_pFtKX6H66_2),.clk(gclk));
	jdff dff_B_1cJgRuth6_2(.din(w_dff_B_pFtKX6H66_2),.dout(w_dff_B_1cJgRuth6_2),.clk(gclk));
	jdff dff_B_sGfhoS9A5_2(.din(w_dff_B_1cJgRuth6_2),.dout(w_dff_B_sGfhoS9A5_2),.clk(gclk));
	jdff dff_B_A4o8wSGS5_2(.din(w_dff_B_sGfhoS9A5_2),.dout(w_dff_B_A4o8wSGS5_2),.clk(gclk));
	jdff dff_B_z8ukxAKN1_2(.din(w_dff_B_A4o8wSGS5_2),.dout(w_dff_B_z8ukxAKN1_2),.clk(gclk));
	jdff dff_B_udZwhBoH5_2(.din(w_dff_B_z8ukxAKN1_2),.dout(w_dff_B_udZwhBoH5_2),.clk(gclk));
	jdff dff_B_Qx1bUMC01_2(.din(w_dff_B_udZwhBoH5_2),.dout(w_dff_B_Qx1bUMC01_2),.clk(gclk));
	jdff dff_B_3VzIIUf90_2(.din(w_dff_B_Qx1bUMC01_2),.dout(w_dff_B_3VzIIUf90_2),.clk(gclk));
	jdff dff_B_9Qkthlom1_2(.din(w_dff_B_3VzIIUf90_2),.dout(w_dff_B_9Qkthlom1_2),.clk(gclk));
	jdff dff_B_DQDjo2Hn4_2(.din(w_dff_B_9Qkthlom1_2),.dout(w_dff_B_DQDjo2Hn4_2),.clk(gclk));
	jdff dff_B_5NGm393O6_2(.din(w_dff_B_DQDjo2Hn4_2),.dout(w_dff_B_5NGm393O6_2),.clk(gclk));
	jdff dff_B_3kFUTehD8_2(.din(w_dff_B_5NGm393O6_2),.dout(w_dff_B_3kFUTehD8_2),.clk(gclk));
	jdff dff_B_QKVueGWt5_1(.din(n1746),.dout(w_dff_B_QKVueGWt5_1),.clk(gclk));
	jdff dff_B_UoYNGMjq0_1(.din(w_dff_B_QKVueGWt5_1),.dout(w_dff_B_UoYNGMjq0_1),.clk(gclk));
	jdff dff_B_t5MPMgJ02_2(.din(n1745),.dout(w_dff_B_t5MPMgJ02_2),.clk(gclk));
	jdff dff_B_lrW06qFI9_2(.din(w_dff_B_t5MPMgJ02_2),.dout(w_dff_B_lrW06qFI9_2),.clk(gclk));
	jdff dff_B_EoIaXoH00_2(.din(w_dff_B_lrW06qFI9_2),.dout(w_dff_B_EoIaXoH00_2),.clk(gclk));
	jdff dff_B_GDcqgL9b0_2(.din(w_dff_B_EoIaXoH00_2),.dout(w_dff_B_GDcqgL9b0_2),.clk(gclk));
	jdff dff_B_d1cknSAX0_2(.din(w_dff_B_GDcqgL9b0_2),.dout(w_dff_B_d1cknSAX0_2),.clk(gclk));
	jdff dff_B_iJOkd3Pb9_2(.din(w_dff_B_d1cknSAX0_2),.dout(w_dff_B_iJOkd3Pb9_2),.clk(gclk));
	jdff dff_B_g7jpPLsb0_2(.din(w_dff_B_iJOkd3Pb9_2),.dout(w_dff_B_g7jpPLsb0_2),.clk(gclk));
	jdff dff_B_LQOt9SSH5_2(.din(w_dff_B_g7jpPLsb0_2),.dout(w_dff_B_LQOt9SSH5_2),.clk(gclk));
	jdff dff_B_rIUQq1Mi8_2(.din(w_dff_B_LQOt9SSH5_2),.dout(w_dff_B_rIUQq1Mi8_2),.clk(gclk));
	jdff dff_B_WrZtnV7W3_2(.din(w_dff_B_rIUQq1Mi8_2),.dout(w_dff_B_WrZtnV7W3_2),.clk(gclk));
	jdff dff_B_1ckAXzvD5_2(.din(w_dff_B_WrZtnV7W3_2),.dout(w_dff_B_1ckAXzvD5_2),.clk(gclk));
	jdff dff_B_OiRVNyhP4_2(.din(w_dff_B_1ckAXzvD5_2),.dout(w_dff_B_OiRVNyhP4_2),.clk(gclk));
	jdff dff_B_FLveHS3u5_2(.din(w_dff_B_OiRVNyhP4_2),.dout(w_dff_B_FLveHS3u5_2),.clk(gclk));
	jdff dff_B_ppEP7JEA1_2(.din(w_dff_B_FLveHS3u5_2),.dout(w_dff_B_ppEP7JEA1_2),.clk(gclk));
	jdff dff_B_KiWTMxKC7_2(.din(w_dff_B_ppEP7JEA1_2),.dout(w_dff_B_KiWTMxKC7_2),.clk(gclk));
	jdff dff_B_dkqkfHcX3_2(.din(w_dff_B_KiWTMxKC7_2),.dout(w_dff_B_dkqkfHcX3_2),.clk(gclk));
	jdff dff_B_v0BD1dhP2_2(.din(w_dff_B_dkqkfHcX3_2),.dout(w_dff_B_v0BD1dhP2_2),.clk(gclk));
	jdff dff_B_vvUL2odx1_2(.din(w_dff_B_v0BD1dhP2_2),.dout(w_dff_B_vvUL2odx1_2),.clk(gclk));
	jdff dff_B_xDkxHkET9_2(.din(w_dff_B_vvUL2odx1_2),.dout(w_dff_B_xDkxHkET9_2),.clk(gclk));
	jdff dff_B_DDfNJLV50_2(.din(w_dff_B_xDkxHkET9_2),.dout(w_dff_B_DDfNJLV50_2),.clk(gclk));
	jdff dff_B_yMK4XQrG6_2(.din(w_dff_B_DDfNJLV50_2),.dout(w_dff_B_yMK4XQrG6_2),.clk(gclk));
	jdff dff_B_E7co62372_2(.din(w_dff_B_yMK4XQrG6_2),.dout(w_dff_B_E7co62372_2),.clk(gclk));
	jdff dff_B_Vs09CW373_2(.din(w_dff_B_E7co62372_2),.dout(w_dff_B_Vs09CW373_2),.clk(gclk));
	jdff dff_B_meUnrAjw7_2(.din(w_dff_B_Vs09CW373_2),.dout(w_dff_B_meUnrAjw7_2),.clk(gclk));
	jdff dff_B_lnKdbOrZ5_2(.din(w_dff_B_meUnrAjw7_2),.dout(w_dff_B_lnKdbOrZ5_2),.clk(gclk));
	jdff dff_B_jEPxsSch6_2(.din(w_dff_B_lnKdbOrZ5_2),.dout(w_dff_B_jEPxsSch6_2),.clk(gclk));
	jdff dff_B_1UbQTLs96_2(.din(w_dff_B_jEPxsSch6_2),.dout(w_dff_B_1UbQTLs96_2),.clk(gclk));
	jdff dff_B_ulXr90JH4_2(.din(w_dff_B_1UbQTLs96_2),.dout(w_dff_B_ulXr90JH4_2),.clk(gclk));
	jdff dff_B_qB7fgw5D7_2(.din(w_dff_B_ulXr90JH4_2),.dout(w_dff_B_qB7fgw5D7_2),.clk(gclk));
	jdff dff_B_Pey73YRh2_2(.din(w_dff_B_qB7fgw5D7_2),.dout(w_dff_B_Pey73YRh2_2),.clk(gclk));
	jdff dff_B_FZG5XH1I7_2(.din(w_dff_B_Pey73YRh2_2),.dout(w_dff_B_FZG5XH1I7_2),.clk(gclk));
	jdff dff_B_H98D4H0h5_2(.din(w_dff_B_FZG5XH1I7_2),.dout(w_dff_B_H98D4H0h5_2),.clk(gclk));
	jdff dff_B_Xq2bfW3m3_2(.din(w_dff_B_H98D4H0h5_2),.dout(w_dff_B_Xq2bfW3m3_2),.clk(gclk));
	jdff dff_B_4wh0O9dz1_2(.din(w_dff_B_Xq2bfW3m3_2),.dout(w_dff_B_4wh0O9dz1_2),.clk(gclk));
	jdff dff_B_SXKCb8oS9_2(.din(w_dff_B_4wh0O9dz1_2),.dout(w_dff_B_SXKCb8oS9_2),.clk(gclk));
	jdff dff_B_cwKLAzCP2_2(.din(w_dff_B_SXKCb8oS9_2),.dout(w_dff_B_cwKLAzCP2_2),.clk(gclk));
	jdff dff_B_4HbENNXZ3_2(.din(w_dff_B_cwKLAzCP2_2),.dout(w_dff_B_4HbENNXZ3_2),.clk(gclk));
	jdff dff_B_3BE3aLDE4_2(.din(w_dff_B_4HbENNXZ3_2),.dout(w_dff_B_3BE3aLDE4_2),.clk(gclk));
	jdff dff_B_Q4sWiyoZ0_2(.din(w_dff_B_3BE3aLDE4_2),.dout(w_dff_B_Q4sWiyoZ0_2),.clk(gclk));
	jdff dff_B_lVKF3b875_2(.din(w_dff_B_Q4sWiyoZ0_2),.dout(w_dff_B_lVKF3b875_2),.clk(gclk));
	jdff dff_B_38muVdk36_2(.din(w_dff_B_lVKF3b875_2),.dout(w_dff_B_38muVdk36_2),.clk(gclk));
	jdff dff_B_yopqtJGK1_2(.din(w_dff_B_38muVdk36_2),.dout(w_dff_B_yopqtJGK1_2),.clk(gclk));
	jdff dff_B_jArYjGoD7_2(.din(w_dff_B_yopqtJGK1_2),.dout(w_dff_B_jArYjGoD7_2),.clk(gclk));
	jdff dff_B_kT7sBeMi1_2(.din(w_dff_B_jArYjGoD7_2),.dout(w_dff_B_kT7sBeMi1_2),.clk(gclk));
	jdff dff_B_21mEbh8I0_2(.din(n1744),.dout(w_dff_B_21mEbh8I0_2),.clk(gclk));
	jdff dff_B_x71n1UtL6_2(.din(w_dff_B_21mEbh8I0_2),.dout(w_dff_B_x71n1UtL6_2),.clk(gclk));
	jdff dff_B_Xz6RaKpE9_2(.din(w_dff_B_x71n1UtL6_2),.dout(w_dff_B_Xz6RaKpE9_2),.clk(gclk));
	jdff dff_B_ZITUsOKo8_2(.din(w_dff_B_Xz6RaKpE9_2),.dout(w_dff_B_ZITUsOKo8_2),.clk(gclk));
	jdff dff_B_TF8YGS6n8_2(.din(w_dff_B_ZITUsOKo8_2),.dout(w_dff_B_TF8YGS6n8_2),.clk(gclk));
	jdff dff_B_y0gQJKMr9_2(.din(w_dff_B_TF8YGS6n8_2),.dout(w_dff_B_y0gQJKMr9_2),.clk(gclk));
	jdff dff_B_A5VmTtr62_2(.din(w_dff_B_y0gQJKMr9_2),.dout(w_dff_B_A5VmTtr62_2),.clk(gclk));
	jdff dff_B_srEb0CD73_2(.din(w_dff_B_A5VmTtr62_2),.dout(w_dff_B_srEb0CD73_2),.clk(gclk));
	jdff dff_B_yIM3PIHa5_2(.din(w_dff_B_srEb0CD73_2),.dout(w_dff_B_yIM3PIHa5_2),.clk(gclk));
	jdff dff_B_bbPAVANc9_2(.din(w_dff_B_yIM3PIHa5_2),.dout(w_dff_B_bbPAVANc9_2),.clk(gclk));
	jdff dff_B_NnziGxkV6_2(.din(w_dff_B_bbPAVANc9_2),.dout(w_dff_B_NnziGxkV6_2),.clk(gclk));
	jdff dff_B_Tu8GgzAT2_2(.din(w_dff_B_NnziGxkV6_2),.dout(w_dff_B_Tu8GgzAT2_2),.clk(gclk));
	jdff dff_B_pvbCDjg29_2(.din(w_dff_B_Tu8GgzAT2_2),.dout(w_dff_B_pvbCDjg29_2),.clk(gclk));
	jdff dff_B_jr9uTGXa7_2(.din(w_dff_B_pvbCDjg29_2),.dout(w_dff_B_jr9uTGXa7_2),.clk(gclk));
	jdff dff_B_vsfo1Fp33_2(.din(w_dff_B_jr9uTGXa7_2),.dout(w_dff_B_vsfo1Fp33_2),.clk(gclk));
	jdff dff_B_rInyRAr98_2(.din(w_dff_B_vsfo1Fp33_2),.dout(w_dff_B_rInyRAr98_2),.clk(gclk));
	jdff dff_B_q34B6lAI9_2(.din(w_dff_B_rInyRAr98_2),.dout(w_dff_B_q34B6lAI9_2),.clk(gclk));
	jdff dff_B_xXnwfbrR8_2(.din(w_dff_B_q34B6lAI9_2),.dout(w_dff_B_xXnwfbrR8_2),.clk(gclk));
	jdff dff_B_bXNbAUji5_2(.din(w_dff_B_xXnwfbrR8_2),.dout(w_dff_B_bXNbAUji5_2),.clk(gclk));
	jdff dff_B_Gh591ANM2_2(.din(w_dff_B_bXNbAUji5_2),.dout(w_dff_B_Gh591ANM2_2),.clk(gclk));
	jdff dff_B_3wibqupe7_2(.din(w_dff_B_Gh591ANM2_2),.dout(w_dff_B_3wibqupe7_2),.clk(gclk));
	jdff dff_B_QHEbQg640_2(.din(w_dff_B_3wibqupe7_2),.dout(w_dff_B_QHEbQg640_2),.clk(gclk));
	jdff dff_B_uNs538Jp8_2(.din(w_dff_B_QHEbQg640_2),.dout(w_dff_B_uNs538Jp8_2),.clk(gclk));
	jdff dff_B_pkx9ikNH4_2(.din(w_dff_B_uNs538Jp8_2),.dout(w_dff_B_pkx9ikNH4_2),.clk(gclk));
	jdff dff_B_yiDogyUX2_2(.din(w_dff_B_pkx9ikNH4_2),.dout(w_dff_B_yiDogyUX2_2),.clk(gclk));
	jdff dff_B_xYrUPg4e8_2(.din(w_dff_B_yiDogyUX2_2),.dout(w_dff_B_xYrUPg4e8_2),.clk(gclk));
	jdff dff_B_jhDuClEt7_2(.din(w_dff_B_xYrUPg4e8_2),.dout(w_dff_B_jhDuClEt7_2),.clk(gclk));
	jdff dff_B_ZAxmcxZr4_2(.din(w_dff_B_jhDuClEt7_2),.dout(w_dff_B_ZAxmcxZr4_2),.clk(gclk));
	jdff dff_B_KJJV1X3J4_2(.din(w_dff_B_ZAxmcxZr4_2),.dout(w_dff_B_KJJV1X3J4_2),.clk(gclk));
	jdff dff_B_VDMfBjA53_2(.din(w_dff_B_KJJV1X3J4_2),.dout(w_dff_B_VDMfBjA53_2),.clk(gclk));
	jdff dff_B_69J16IMU4_2(.din(w_dff_B_VDMfBjA53_2),.dout(w_dff_B_69J16IMU4_2),.clk(gclk));
	jdff dff_B_YhxIyYQG3_2(.din(w_dff_B_69J16IMU4_2),.dout(w_dff_B_YhxIyYQG3_2),.clk(gclk));
	jdff dff_B_2K4ObXET2_2(.din(w_dff_B_YhxIyYQG3_2),.dout(w_dff_B_2K4ObXET2_2),.clk(gclk));
	jdff dff_B_RqV1isF89_2(.din(w_dff_B_2K4ObXET2_2),.dout(w_dff_B_RqV1isF89_2),.clk(gclk));
	jdff dff_B_xuQuZlGa8_2(.din(w_dff_B_RqV1isF89_2),.dout(w_dff_B_xuQuZlGa8_2),.clk(gclk));
	jdff dff_B_R4bdEiuo9_2(.din(w_dff_B_xuQuZlGa8_2),.dout(w_dff_B_R4bdEiuo9_2),.clk(gclk));
	jdff dff_B_6MT5HUZl8_2(.din(w_dff_B_R4bdEiuo9_2),.dout(w_dff_B_6MT5HUZl8_2),.clk(gclk));
	jdff dff_B_7p8E9svd4_2(.din(w_dff_B_6MT5HUZl8_2),.dout(w_dff_B_7p8E9svd4_2),.clk(gclk));
	jdff dff_B_qOMa1gSn6_2(.din(w_dff_B_7p8E9svd4_2),.dout(w_dff_B_qOMa1gSn6_2),.clk(gclk));
	jdff dff_B_RcHkkidg7_2(.din(w_dff_B_qOMa1gSn6_2),.dout(w_dff_B_RcHkkidg7_2),.clk(gclk));
	jdff dff_B_g5tMIoOe7_2(.din(w_dff_B_RcHkkidg7_2),.dout(w_dff_B_g5tMIoOe7_2),.clk(gclk));
	jdff dff_B_E2sHLCiD5_2(.din(w_dff_B_g5tMIoOe7_2),.dout(w_dff_B_E2sHLCiD5_2),.clk(gclk));
	jdff dff_B_g7pGMShE4_2(.din(w_dff_B_E2sHLCiD5_2),.dout(w_dff_B_g7pGMShE4_2),.clk(gclk));
	jdff dff_B_IWFQQsI89_2(.din(w_dff_B_g7pGMShE4_2),.dout(w_dff_B_IWFQQsI89_2),.clk(gclk));
	jdff dff_B_N4xurE2H7_2(.din(w_dff_B_IWFQQsI89_2),.dout(w_dff_B_N4xurE2H7_2),.clk(gclk));
	jdff dff_B_ziA82jg42_2(.din(w_dff_B_N4xurE2H7_2),.dout(w_dff_B_ziA82jg42_2),.clk(gclk));
	jdff dff_B_2E4qR4cc6_2(.din(n1743),.dout(w_dff_B_2E4qR4cc6_2),.clk(gclk));
	jdff dff_B_4Bt6y4zt0_1(.din(n1741),.dout(w_dff_B_4Bt6y4zt0_1),.clk(gclk));
	jdff dff_B_99QiTFjo3_2(.din(n1699),.dout(w_dff_B_99QiTFjo3_2),.clk(gclk));
	jdff dff_B_puupNxe36_2(.din(w_dff_B_99QiTFjo3_2),.dout(w_dff_B_puupNxe36_2),.clk(gclk));
	jdff dff_B_gmfk8Z0c1_2(.din(w_dff_B_puupNxe36_2),.dout(w_dff_B_gmfk8Z0c1_2),.clk(gclk));
	jdff dff_B_55CQjVaE2_2(.din(w_dff_B_gmfk8Z0c1_2),.dout(w_dff_B_55CQjVaE2_2),.clk(gclk));
	jdff dff_B_YdQAmE2O8_2(.din(w_dff_B_55CQjVaE2_2),.dout(w_dff_B_YdQAmE2O8_2),.clk(gclk));
	jdff dff_B_50zTlLwx8_2(.din(w_dff_B_YdQAmE2O8_2),.dout(w_dff_B_50zTlLwx8_2),.clk(gclk));
	jdff dff_B_EbqiYn3y9_2(.din(w_dff_B_50zTlLwx8_2),.dout(w_dff_B_EbqiYn3y9_2),.clk(gclk));
	jdff dff_B_XKTlDXUp7_2(.din(w_dff_B_EbqiYn3y9_2),.dout(w_dff_B_XKTlDXUp7_2),.clk(gclk));
	jdff dff_B_J9eUGxIC7_2(.din(w_dff_B_XKTlDXUp7_2),.dout(w_dff_B_J9eUGxIC7_2),.clk(gclk));
	jdff dff_B_upil0NRb5_2(.din(w_dff_B_J9eUGxIC7_2),.dout(w_dff_B_upil0NRb5_2),.clk(gclk));
	jdff dff_B_XQ00n42s0_2(.din(w_dff_B_upil0NRb5_2),.dout(w_dff_B_XQ00n42s0_2),.clk(gclk));
	jdff dff_B_0N8rdUdi5_2(.din(w_dff_B_XQ00n42s0_2),.dout(w_dff_B_0N8rdUdi5_2),.clk(gclk));
	jdff dff_B_op4gHcy56_2(.din(w_dff_B_0N8rdUdi5_2),.dout(w_dff_B_op4gHcy56_2),.clk(gclk));
	jdff dff_B_zBgIB6pW4_2(.din(w_dff_B_op4gHcy56_2),.dout(w_dff_B_zBgIB6pW4_2),.clk(gclk));
	jdff dff_B_P18SjuOx9_2(.din(w_dff_B_zBgIB6pW4_2),.dout(w_dff_B_P18SjuOx9_2),.clk(gclk));
	jdff dff_B_8nVLgy2D1_2(.din(w_dff_B_P18SjuOx9_2),.dout(w_dff_B_8nVLgy2D1_2),.clk(gclk));
	jdff dff_B_4UjSdbpg6_2(.din(w_dff_B_8nVLgy2D1_2),.dout(w_dff_B_4UjSdbpg6_2),.clk(gclk));
	jdff dff_B_H63wemc78_2(.din(w_dff_B_4UjSdbpg6_2),.dout(w_dff_B_H63wemc78_2),.clk(gclk));
	jdff dff_B_TsuXj3H28_2(.din(w_dff_B_H63wemc78_2),.dout(w_dff_B_TsuXj3H28_2),.clk(gclk));
	jdff dff_B_6pSlz7uU4_2(.din(w_dff_B_TsuXj3H28_2),.dout(w_dff_B_6pSlz7uU4_2),.clk(gclk));
	jdff dff_B_1RDq1Ei12_2(.din(w_dff_B_6pSlz7uU4_2),.dout(w_dff_B_1RDq1Ei12_2),.clk(gclk));
	jdff dff_B_N5vehd0F0_2(.din(w_dff_B_1RDq1Ei12_2),.dout(w_dff_B_N5vehd0F0_2),.clk(gclk));
	jdff dff_B_smXfCofL7_2(.din(w_dff_B_N5vehd0F0_2),.dout(w_dff_B_smXfCofL7_2),.clk(gclk));
	jdff dff_B_fGhviDAs9_2(.din(w_dff_B_smXfCofL7_2),.dout(w_dff_B_fGhviDAs9_2),.clk(gclk));
	jdff dff_B_FkjDaoI48_2(.din(w_dff_B_fGhviDAs9_2),.dout(w_dff_B_FkjDaoI48_2),.clk(gclk));
	jdff dff_B_pTgCKzc72_2(.din(w_dff_B_FkjDaoI48_2),.dout(w_dff_B_pTgCKzc72_2),.clk(gclk));
	jdff dff_B_kFprMZUL1_2(.din(w_dff_B_pTgCKzc72_2),.dout(w_dff_B_kFprMZUL1_2),.clk(gclk));
	jdff dff_B_DylwgarZ7_2(.din(w_dff_B_kFprMZUL1_2),.dout(w_dff_B_DylwgarZ7_2),.clk(gclk));
	jdff dff_B_9Zoh5yMy3_2(.din(w_dff_B_DylwgarZ7_2),.dout(w_dff_B_9Zoh5yMy3_2),.clk(gclk));
	jdff dff_B_cQg39ptg1_2(.din(w_dff_B_9Zoh5yMy3_2),.dout(w_dff_B_cQg39ptg1_2),.clk(gclk));
	jdff dff_B_W8Se07348_2(.din(w_dff_B_cQg39ptg1_2),.dout(w_dff_B_W8Se07348_2),.clk(gclk));
	jdff dff_B_rTnB1yrs8_2(.din(w_dff_B_W8Se07348_2),.dout(w_dff_B_rTnB1yrs8_2),.clk(gclk));
	jdff dff_B_4Lvv8VEr4_2(.din(w_dff_B_rTnB1yrs8_2),.dout(w_dff_B_4Lvv8VEr4_2),.clk(gclk));
	jdff dff_B_2ELtoSym4_2(.din(w_dff_B_4Lvv8VEr4_2),.dout(w_dff_B_2ELtoSym4_2),.clk(gclk));
	jdff dff_B_2hmTYA1d8_2(.din(w_dff_B_2ELtoSym4_2),.dout(w_dff_B_2hmTYA1d8_2),.clk(gclk));
	jdff dff_B_1oIU5lsy4_2(.din(w_dff_B_2hmTYA1d8_2),.dout(w_dff_B_1oIU5lsy4_2),.clk(gclk));
	jdff dff_B_8tnOjYpD1_2(.din(w_dff_B_1oIU5lsy4_2),.dout(w_dff_B_8tnOjYpD1_2),.clk(gclk));
	jdff dff_B_JFD7i89n1_2(.din(w_dff_B_8tnOjYpD1_2),.dout(w_dff_B_JFD7i89n1_2),.clk(gclk));
	jdff dff_B_Zf8WhofN0_2(.din(w_dff_B_JFD7i89n1_2),.dout(w_dff_B_Zf8WhofN0_2),.clk(gclk));
	jdff dff_B_tHwOVsXV7_2(.din(w_dff_B_Zf8WhofN0_2),.dout(w_dff_B_tHwOVsXV7_2),.clk(gclk));
	jdff dff_B_Y9t54LXk6_2(.din(w_dff_B_tHwOVsXV7_2),.dout(w_dff_B_Y9t54LXk6_2),.clk(gclk));
	jdff dff_B_mUrMKwmt8_2(.din(w_dff_B_Y9t54LXk6_2),.dout(w_dff_B_mUrMKwmt8_2),.clk(gclk));
	jdff dff_B_0DfkFQY61_2(.din(w_dff_B_mUrMKwmt8_2),.dout(w_dff_B_0DfkFQY61_2),.clk(gclk));
	jdff dff_B_GFrhTRzC6_1(.din(n1705),.dout(w_dff_B_GFrhTRzC6_1),.clk(gclk));
	jdff dff_B_6xgTCNBr0_1(.din(w_dff_B_GFrhTRzC6_1),.dout(w_dff_B_6xgTCNBr0_1),.clk(gclk));
	jdff dff_B_HtI17TAk1_2(.din(n1704),.dout(w_dff_B_HtI17TAk1_2),.clk(gclk));
	jdff dff_B_gAMR6wl58_2(.din(w_dff_B_HtI17TAk1_2),.dout(w_dff_B_gAMR6wl58_2),.clk(gclk));
	jdff dff_B_KVN4DUkP1_2(.din(w_dff_B_gAMR6wl58_2),.dout(w_dff_B_KVN4DUkP1_2),.clk(gclk));
	jdff dff_B_XxjmFJb54_2(.din(w_dff_B_KVN4DUkP1_2),.dout(w_dff_B_XxjmFJb54_2),.clk(gclk));
	jdff dff_B_v0lSXM3x3_2(.din(w_dff_B_XxjmFJb54_2),.dout(w_dff_B_v0lSXM3x3_2),.clk(gclk));
	jdff dff_B_R7odIVcI1_2(.din(w_dff_B_v0lSXM3x3_2),.dout(w_dff_B_R7odIVcI1_2),.clk(gclk));
	jdff dff_B_ng9zFUrw5_2(.din(w_dff_B_R7odIVcI1_2),.dout(w_dff_B_ng9zFUrw5_2),.clk(gclk));
	jdff dff_B_RqejzdbV0_2(.din(w_dff_B_ng9zFUrw5_2),.dout(w_dff_B_RqejzdbV0_2),.clk(gclk));
	jdff dff_B_HlUJwcvE6_2(.din(w_dff_B_RqejzdbV0_2),.dout(w_dff_B_HlUJwcvE6_2),.clk(gclk));
	jdff dff_B_X7qDLgT79_2(.din(w_dff_B_HlUJwcvE6_2),.dout(w_dff_B_X7qDLgT79_2),.clk(gclk));
	jdff dff_B_bwROm8Dp8_2(.din(w_dff_B_X7qDLgT79_2),.dout(w_dff_B_bwROm8Dp8_2),.clk(gclk));
	jdff dff_B_jDmUArPP6_2(.din(w_dff_B_bwROm8Dp8_2),.dout(w_dff_B_jDmUArPP6_2),.clk(gclk));
	jdff dff_B_z3cttkUb5_2(.din(w_dff_B_jDmUArPP6_2),.dout(w_dff_B_z3cttkUb5_2),.clk(gclk));
	jdff dff_B_FSJYm9Vn8_2(.din(w_dff_B_z3cttkUb5_2),.dout(w_dff_B_FSJYm9Vn8_2),.clk(gclk));
	jdff dff_B_gBK1f5QN1_2(.din(w_dff_B_FSJYm9Vn8_2),.dout(w_dff_B_gBK1f5QN1_2),.clk(gclk));
	jdff dff_B_36taeYWU1_2(.din(w_dff_B_gBK1f5QN1_2),.dout(w_dff_B_36taeYWU1_2),.clk(gclk));
	jdff dff_B_NPRxi8OQ9_2(.din(w_dff_B_36taeYWU1_2),.dout(w_dff_B_NPRxi8OQ9_2),.clk(gclk));
	jdff dff_B_buj56fGq6_2(.din(w_dff_B_NPRxi8OQ9_2),.dout(w_dff_B_buj56fGq6_2),.clk(gclk));
	jdff dff_B_L0PTnb5n9_2(.din(w_dff_B_buj56fGq6_2),.dout(w_dff_B_L0PTnb5n9_2),.clk(gclk));
	jdff dff_B_VWSX9ZV76_2(.din(w_dff_B_L0PTnb5n9_2),.dout(w_dff_B_VWSX9ZV76_2),.clk(gclk));
	jdff dff_B_zQI3K1NZ0_2(.din(w_dff_B_VWSX9ZV76_2),.dout(w_dff_B_zQI3K1NZ0_2),.clk(gclk));
	jdff dff_B_s7afqwyq1_2(.din(w_dff_B_zQI3K1NZ0_2),.dout(w_dff_B_s7afqwyq1_2),.clk(gclk));
	jdff dff_B_55siENpu6_2(.din(w_dff_B_s7afqwyq1_2),.dout(w_dff_B_55siENpu6_2),.clk(gclk));
	jdff dff_B_5LFHCW8g7_2(.din(w_dff_B_55siENpu6_2),.dout(w_dff_B_5LFHCW8g7_2),.clk(gclk));
	jdff dff_B_Vl9j5ygu2_2(.din(w_dff_B_5LFHCW8g7_2),.dout(w_dff_B_Vl9j5ygu2_2),.clk(gclk));
	jdff dff_B_u8IcZ4Sm7_2(.din(w_dff_B_Vl9j5ygu2_2),.dout(w_dff_B_u8IcZ4Sm7_2),.clk(gclk));
	jdff dff_B_HgXMQ7ya9_2(.din(w_dff_B_u8IcZ4Sm7_2),.dout(w_dff_B_HgXMQ7ya9_2),.clk(gclk));
	jdff dff_B_YgMHxllh6_2(.din(w_dff_B_HgXMQ7ya9_2),.dout(w_dff_B_YgMHxllh6_2),.clk(gclk));
	jdff dff_B_unGaVVXG1_2(.din(w_dff_B_YgMHxllh6_2),.dout(w_dff_B_unGaVVXG1_2),.clk(gclk));
	jdff dff_B_Vc7kbnJk1_2(.din(w_dff_B_unGaVVXG1_2),.dout(w_dff_B_Vc7kbnJk1_2),.clk(gclk));
	jdff dff_B_1Vbt5vQf8_2(.din(w_dff_B_Vc7kbnJk1_2),.dout(w_dff_B_1Vbt5vQf8_2),.clk(gclk));
	jdff dff_B_6BBe5St64_2(.din(w_dff_B_1Vbt5vQf8_2),.dout(w_dff_B_6BBe5St64_2),.clk(gclk));
	jdff dff_B_3CEOJI8g6_2(.din(w_dff_B_6BBe5St64_2),.dout(w_dff_B_3CEOJI8g6_2),.clk(gclk));
	jdff dff_B_Cvpd7jbn4_2(.din(w_dff_B_3CEOJI8g6_2),.dout(w_dff_B_Cvpd7jbn4_2),.clk(gclk));
	jdff dff_B_62vw1PCN2_2(.din(w_dff_B_Cvpd7jbn4_2),.dout(w_dff_B_62vw1PCN2_2),.clk(gclk));
	jdff dff_B_g9EhUTMJ3_2(.din(w_dff_B_62vw1PCN2_2),.dout(w_dff_B_g9EhUTMJ3_2),.clk(gclk));
	jdff dff_B_PBlEnHlZ2_2(.din(w_dff_B_g9EhUTMJ3_2),.dout(w_dff_B_PBlEnHlZ2_2),.clk(gclk));
	jdff dff_B_Zby2zGPG7_2(.din(w_dff_B_PBlEnHlZ2_2),.dout(w_dff_B_Zby2zGPG7_2),.clk(gclk));
	jdff dff_B_uhgPa5op1_2(.din(w_dff_B_Zby2zGPG7_2),.dout(w_dff_B_uhgPa5op1_2),.clk(gclk));
	jdff dff_B_GMBo0y002_2(.din(w_dff_B_uhgPa5op1_2),.dout(w_dff_B_GMBo0y002_2),.clk(gclk));
	jdff dff_B_uKRD97Xl5_2(.din(n1703),.dout(w_dff_B_uKRD97Xl5_2),.clk(gclk));
	jdff dff_B_uJrXNTd85_2(.din(w_dff_B_uKRD97Xl5_2),.dout(w_dff_B_uJrXNTd85_2),.clk(gclk));
	jdff dff_B_pwbLZByw2_2(.din(w_dff_B_uJrXNTd85_2),.dout(w_dff_B_pwbLZByw2_2),.clk(gclk));
	jdff dff_B_NJqILe4L0_2(.din(w_dff_B_pwbLZByw2_2),.dout(w_dff_B_NJqILe4L0_2),.clk(gclk));
	jdff dff_B_Uwkfa8z69_2(.din(w_dff_B_NJqILe4L0_2),.dout(w_dff_B_Uwkfa8z69_2),.clk(gclk));
	jdff dff_B_XUthNvBx5_2(.din(w_dff_B_Uwkfa8z69_2),.dout(w_dff_B_XUthNvBx5_2),.clk(gclk));
	jdff dff_B_A0lD3kJz7_2(.din(w_dff_B_XUthNvBx5_2),.dout(w_dff_B_A0lD3kJz7_2),.clk(gclk));
	jdff dff_B_am6QIkWZ5_2(.din(w_dff_B_A0lD3kJz7_2),.dout(w_dff_B_am6QIkWZ5_2),.clk(gclk));
	jdff dff_B_vSN9umEr5_2(.din(w_dff_B_am6QIkWZ5_2),.dout(w_dff_B_vSN9umEr5_2),.clk(gclk));
	jdff dff_B_WuM1gtbH4_2(.din(w_dff_B_vSN9umEr5_2),.dout(w_dff_B_WuM1gtbH4_2),.clk(gclk));
	jdff dff_B_OU1O8fij0_2(.din(w_dff_B_WuM1gtbH4_2),.dout(w_dff_B_OU1O8fij0_2),.clk(gclk));
	jdff dff_B_ecMNIr6G1_2(.din(w_dff_B_OU1O8fij0_2),.dout(w_dff_B_ecMNIr6G1_2),.clk(gclk));
	jdff dff_B_BOPwxFL67_2(.din(w_dff_B_ecMNIr6G1_2),.dout(w_dff_B_BOPwxFL67_2),.clk(gclk));
	jdff dff_B_7HtFwwe50_2(.din(w_dff_B_BOPwxFL67_2),.dout(w_dff_B_7HtFwwe50_2),.clk(gclk));
	jdff dff_B_QEaLeHvU7_2(.din(w_dff_B_7HtFwwe50_2),.dout(w_dff_B_QEaLeHvU7_2),.clk(gclk));
	jdff dff_B_fDy71Ei10_2(.din(w_dff_B_QEaLeHvU7_2),.dout(w_dff_B_fDy71Ei10_2),.clk(gclk));
	jdff dff_B_PmBQaupu9_2(.din(w_dff_B_fDy71Ei10_2),.dout(w_dff_B_PmBQaupu9_2),.clk(gclk));
	jdff dff_B_srpOVKbr2_2(.din(w_dff_B_PmBQaupu9_2),.dout(w_dff_B_srpOVKbr2_2),.clk(gclk));
	jdff dff_B_fWM9lthE8_2(.din(w_dff_B_srpOVKbr2_2),.dout(w_dff_B_fWM9lthE8_2),.clk(gclk));
	jdff dff_B_3nJq1qak6_2(.din(w_dff_B_fWM9lthE8_2),.dout(w_dff_B_3nJq1qak6_2),.clk(gclk));
	jdff dff_B_JWO8f5rj0_2(.din(w_dff_B_3nJq1qak6_2),.dout(w_dff_B_JWO8f5rj0_2),.clk(gclk));
	jdff dff_B_HMkCkOnn1_2(.din(w_dff_B_JWO8f5rj0_2),.dout(w_dff_B_HMkCkOnn1_2),.clk(gclk));
	jdff dff_B_rmpInCQi9_2(.din(w_dff_B_HMkCkOnn1_2),.dout(w_dff_B_rmpInCQi9_2),.clk(gclk));
	jdff dff_B_5LcFkU4d1_2(.din(w_dff_B_rmpInCQi9_2),.dout(w_dff_B_5LcFkU4d1_2),.clk(gclk));
	jdff dff_B_fy6DyESh8_2(.din(w_dff_B_5LcFkU4d1_2),.dout(w_dff_B_fy6DyESh8_2),.clk(gclk));
	jdff dff_B_gGHflhEb5_2(.din(w_dff_B_fy6DyESh8_2),.dout(w_dff_B_gGHflhEb5_2),.clk(gclk));
	jdff dff_B_6pt5q2tr5_2(.din(w_dff_B_gGHflhEb5_2),.dout(w_dff_B_6pt5q2tr5_2),.clk(gclk));
	jdff dff_B_61jeyu9q3_2(.din(w_dff_B_6pt5q2tr5_2),.dout(w_dff_B_61jeyu9q3_2),.clk(gclk));
	jdff dff_B_GD17m7B46_2(.din(w_dff_B_61jeyu9q3_2),.dout(w_dff_B_GD17m7B46_2),.clk(gclk));
	jdff dff_B_8XUYucIN7_2(.din(w_dff_B_GD17m7B46_2),.dout(w_dff_B_8XUYucIN7_2),.clk(gclk));
	jdff dff_B_8BIw16mB0_2(.din(w_dff_B_8XUYucIN7_2),.dout(w_dff_B_8BIw16mB0_2),.clk(gclk));
	jdff dff_B_2Fduc4aY2_2(.din(w_dff_B_8BIw16mB0_2),.dout(w_dff_B_2Fduc4aY2_2),.clk(gclk));
	jdff dff_B_821GBm5b2_2(.din(w_dff_B_2Fduc4aY2_2),.dout(w_dff_B_821GBm5b2_2),.clk(gclk));
	jdff dff_B_nSgVZuvB2_2(.din(w_dff_B_821GBm5b2_2),.dout(w_dff_B_nSgVZuvB2_2),.clk(gclk));
	jdff dff_B_THRcDXML9_2(.din(w_dff_B_nSgVZuvB2_2),.dout(w_dff_B_THRcDXML9_2),.clk(gclk));
	jdff dff_B_DxNT2And2_2(.din(w_dff_B_THRcDXML9_2),.dout(w_dff_B_DxNT2And2_2),.clk(gclk));
	jdff dff_B_UIQV9kfH2_2(.din(w_dff_B_DxNT2And2_2),.dout(w_dff_B_UIQV9kfH2_2),.clk(gclk));
	jdff dff_B_hqHSZuvW4_2(.din(w_dff_B_UIQV9kfH2_2),.dout(w_dff_B_hqHSZuvW4_2),.clk(gclk));
	jdff dff_B_UsfujUSL3_2(.din(w_dff_B_hqHSZuvW4_2),.dout(w_dff_B_UsfujUSL3_2),.clk(gclk));
	jdff dff_B_QZeg2vO21_2(.din(w_dff_B_UsfujUSL3_2),.dout(w_dff_B_QZeg2vO21_2),.clk(gclk));
	jdff dff_B_RNw92S2o0_2(.din(w_dff_B_QZeg2vO21_2),.dout(w_dff_B_RNw92S2o0_2),.clk(gclk));
	jdff dff_B_Yf9oaDTh0_2(.din(w_dff_B_RNw92S2o0_2),.dout(w_dff_B_Yf9oaDTh0_2),.clk(gclk));
	jdff dff_B_jmMqyqcm9_2(.din(n1702),.dout(w_dff_B_jmMqyqcm9_2),.clk(gclk));
	jdff dff_B_FYAmhI927_1(.din(n1700),.dout(w_dff_B_FYAmhI927_1),.clk(gclk));
	jdff dff_B_hHjWGShV1_2(.din(n1648),.dout(w_dff_B_hHjWGShV1_2),.clk(gclk));
	jdff dff_B_UL9m2h943_2(.din(w_dff_B_hHjWGShV1_2),.dout(w_dff_B_UL9m2h943_2),.clk(gclk));
	jdff dff_B_uK8eEL0y1_2(.din(w_dff_B_UL9m2h943_2),.dout(w_dff_B_uK8eEL0y1_2),.clk(gclk));
	jdff dff_B_qaujD78D0_2(.din(w_dff_B_uK8eEL0y1_2),.dout(w_dff_B_qaujD78D0_2),.clk(gclk));
	jdff dff_B_e6BIrDic3_2(.din(w_dff_B_qaujD78D0_2),.dout(w_dff_B_e6BIrDic3_2),.clk(gclk));
	jdff dff_B_bz3w8n586_2(.din(w_dff_B_e6BIrDic3_2),.dout(w_dff_B_bz3w8n586_2),.clk(gclk));
	jdff dff_B_ABBDbDiQ0_2(.din(w_dff_B_bz3w8n586_2),.dout(w_dff_B_ABBDbDiQ0_2),.clk(gclk));
	jdff dff_B_g8wW0jOW5_2(.din(w_dff_B_ABBDbDiQ0_2),.dout(w_dff_B_g8wW0jOW5_2),.clk(gclk));
	jdff dff_B_veUdx0l33_2(.din(w_dff_B_g8wW0jOW5_2),.dout(w_dff_B_veUdx0l33_2),.clk(gclk));
	jdff dff_B_jO3H6MLN1_2(.din(w_dff_B_veUdx0l33_2),.dout(w_dff_B_jO3H6MLN1_2),.clk(gclk));
	jdff dff_B_LYmXvikb1_2(.din(w_dff_B_jO3H6MLN1_2),.dout(w_dff_B_LYmXvikb1_2),.clk(gclk));
	jdff dff_B_LOSSiULb0_2(.din(w_dff_B_LYmXvikb1_2),.dout(w_dff_B_LOSSiULb0_2),.clk(gclk));
	jdff dff_B_HERjnJit9_2(.din(w_dff_B_LOSSiULb0_2),.dout(w_dff_B_HERjnJit9_2),.clk(gclk));
	jdff dff_B_bWRSBSn73_2(.din(w_dff_B_HERjnJit9_2),.dout(w_dff_B_bWRSBSn73_2),.clk(gclk));
	jdff dff_B_GWqy7FtZ7_2(.din(w_dff_B_bWRSBSn73_2),.dout(w_dff_B_GWqy7FtZ7_2),.clk(gclk));
	jdff dff_B_C509QPgg1_2(.din(w_dff_B_GWqy7FtZ7_2),.dout(w_dff_B_C509QPgg1_2),.clk(gclk));
	jdff dff_B_Fxb7o3wR7_2(.din(w_dff_B_C509QPgg1_2),.dout(w_dff_B_Fxb7o3wR7_2),.clk(gclk));
	jdff dff_B_ruzmsfsF0_2(.din(w_dff_B_Fxb7o3wR7_2),.dout(w_dff_B_ruzmsfsF0_2),.clk(gclk));
	jdff dff_B_LtLCSeUH3_2(.din(w_dff_B_ruzmsfsF0_2),.dout(w_dff_B_LtLCSeUH3_2),.clk(gclk));
	jdff dff_B_Slm2Hbcx8_2(.din(w_dff_B_LtLCSeUH3_2),.dout(w_dff_B_Slm2Hbcx8_2),.clk(gclk));
	jdff dff_B_SbdBcWsb4_2(.din(w_dff_B_Slm2Hbcx8_2),.dout(w_dff_B_SbdBcWsb4_2),.clk(gclk));
	jdff dff_B_36GZfrMK8_2(.din(w_dff_B_SbdBcWsb4_2),.dout(w_dff_B_36GZfrMK8_2),.clk(gclk));
	jdff dff_B_3aPlP3zY3_2(.din(w_dff_B_36GZfrMK8_2),.dout(w_dff_B_3aPlP3zY3_2),.clk(gclk));
	jdff dff_B_sdF3dOd54_2(.din(w_dff_B_3aPlP3zY3_2),.dout(w_dff_B_sdF3dOd54_2),.clk(gclk));
	jdff dff_B_qByIQEVR2_2(.din(w_dff_B_sdF3dOd54_2),.dout(w_dff_B_qByIQEVR2_2),.clk(gclk));
	jdff dff_B_xdbSU1DA6_2(.din(w_dff_B_qByIQEVR2_2),.dout(w_dff_B_xdbSU1DA6_2),.clk(gclk));
	jdff dff_B_nssK0Cdd5_2(.din(w_dff_B_xdbSU1DA6_2),.dout(w_dff_B_nssK0Cdd5_2),.clk(gclk));
	jdff dff_B_dNQoKXOx3_2(.din(w_dff_B_nssK0Cdd5_2),.dout(w_dff_B_dNQoKXOx3_2),.clk(gclk));
	jdff dff_B_0XHagwRG1_2(.din(w_dff_B_dNQoKXOx3_2),.dout(w_dff_B_0XHagwRG1_2),.clk(gclk));
	jdff dff_B_erVG94Jm5_2(.din(w_dff_B_0XHagwRG1_2),.dout(w_dff_B_erVG94Jm5_2),.clk(gclk));
	jdff dff_B_O9iQwq537_2(.din(w_dff_B_erVG94Jm5_2),.dout(w_dff_B_O9iQwq537_2),.clk(gclk));
	jdff dff_B_zzUhDKMB8_2(.din(w_dff_B_O9iQwq537_2),.dout(w_dff_B_zzUhDKMB8_2),.clk(gclk));
	jdff dff_B_3vAkFII14_2(.din(w_dff_B_zzUhDKMB8_2),.dout(w_dff_B_3vAkFII14_2),.clk(gclk));
	jdff dff_B_iRkRLu2k1_2(.din(w_dff_B_3vAkFII14_2),.dout(w_dff_B_iRkRLu2k1_2),.clk(gclk));
	jdff dff_B_CpE1fB8t3_2(.din(w_dff_B_iRkRLu2k1_2),.dout(w_dff_B_CpE1fB8t3_2),.clk(gclk));
	jdff dff_B_OHmUMgqe9_2(.din(w_dff_B_CpE1fB8t3_2),.dout(w_dff_B_OHmUMgqe9_2),.clk(gclk));
	jdff dff_B_Big0HdWt4_2(.din(w_dff_B_OHmUMgqe9_2),.dout(w_dff_B_Big0HdWt4_2),.clk(gclk));
	jdff dff_B_nYaLSc6g8_2(.din(w_dff_B_Big0HdWt4_2),.dout(w_dff_B_nYaLSc6g8_2),.clk(gclk));
	jdff dff_B_rQO4g00b5_2(.din(w_dff_B_nYaLSc6g8_2),.dout(w_dff_B_rQO4g00b5_2),.clk(gclk));
	jdff dff_B_xNpPTo8O6_1(.din(n1654),.dout(w_dff_B_xNpPTo8O6_1),.clk(gclk));
	jdff dff_B_Hrnhfkl04_1(.din(w_dff_B_xNpPTo8O6_1),.dout(w_dff_B_Hrnhfkl04_1),.clk(gclk));
	jdff dff_B_aiAv9iMA3_2(.din(n1653),.dout(w_dff_B_aiAv9iMA3_2),.clk(gclk));
	jdff dff_B_4qQoKklD7_2(.din(w_dff_B_aiAv9iMA3_2),.dout(w_dff_B_4qQoKklD7_2),.clk(gclk));
	jdff dff_B_ky0nFzQR3_2(.din(w_dff_B_4qQoKklD7_2),.dout(w_dff_B_ky0nFzQR3_2),.clk(gclk));
	jdff dff_B_DXAkzDQ93_2(.din(w_dff_B_ky0nFzQR3_2),.dout(w_dff_B_DXAkzDQ93_2),.clk(gclk));
	jdff dff_B_DJToPCO48_2(.din(w_dff_B_DXAkzDQ93_2),.dout(w_dff_B_DJToPCO48_2),.clk(gclk));
	jdff dff_B_unAENyFN0_2(.din(w_dff_B_DJToPCO48_2),.dout(w_dff_B_unAENyFN0_2),.clk(gclk));
	jdff dff_B_33wbuzg13_2(.din(w_dff_B_unAENyFN0_2),.dout(w_dff_B_33wbuzg13_2),.clk(gclk));
	jdff dff_B_ZOilHMra3_2(.din(w_dff_B_33wbuzg13_2),.dout(w_dff_B_ZOilHMra3_2),.clk(gclk));
	jdff dff_B_xqC0jtwH6_2(.din(w_dff_B_ZOilHMra3_2),.dout(w_dff_B_xqC0jtwH6_2),.clk(gclk));
	jdff dff_B_cuglOGOZ2_2(.din(w_dff_B_xqC0jtwH6_2),.dout(w_dff_B_cuglOGOZ2_2),.clk(gclk));
	jdff dff_B_nK7loTJd2_2(.din(w_dff_B_cuglOGOZ2_2),.dout(w_dff_B_nK7loTJd2_2),.clk(gclk));
	jdff dff_B_qMskERQP1_2(.din(w_dff_B_nK7loTJd2_2),.dout(w_dff_B_qMskERQP1_2),.clk(gclk));
	jdff dff_B_NxqkiUSf0_2(.din(w_dff_B_qMskERQP1_2),.dout(w_dff_B_NxqkiUSf0_2),.clk(gclk));
	jdff dff_B_UqrGwyf40_2(.din(w_dff_B_NxqkiUSf0_2),.dout(w_dff_B_UqrGwyf40_2),.clk(gclk));
	jdff dff_B_Nzw9a53j2_2(.din(w_dff_B_UqrGwyf40_2),.dout(w_dff_B_Nzw9a53j2_2),.clk(gclk));
	jdff dff_B_hBXJ9mjI7_2(.din(w_dff_B_Nzw9a53j2_2),.dout(w_dff_B_hBXJ9mjI7_2),.clk(gclk));
	jdff dff_B_Lan52Tx93_2(.din(w_dff_B_hBXJ9mjI7_2),.dout(w_dff_B_Lan52Tx93_2),.clk(gclk));
	jdff dff_B_TgLl0Zq53_2(.din(w_dff_B_Lan52Tx93_2),.dout(w_dff_B_TgLl0Zq53_2),.clk(gclk));
	jdff dff_B_0VmyhUMs9_2(.din(w_dff_B_TgLl0Zq53_2),.dout(w_dff_B_0VmyhUMs9_2),.clk(gclk));
	jdff dff_B_yXudTNvo4_2(.din(w_dff_B_0VmyhUMs9_2),.dout(w_dff_B_yXudTNvo4_2),.clk(gclk));
	jdff dff_B_1G4XNrYe0_2(.din(w_dff_B_yXudTNvo4_2),.dout(w_dff_B_1G4XNrYe0_2),.clk(gclk));
	jdff dff_B_3kQhJqD36_2(.din(w_dff_B_1G4XNrYe0_2),.dout(w_dff_B_3kQhJqD36_2),.clk(gclk));
	jdff dff_B_X89BGa8y1_2(.din(w_dff_B_3kQhJqD36_2),.dout(w_dff_B_X89BGa8y1_2),.clk(gclk));
	jdff dff_B_NMO1wSXk8_2(.din(w_dff_B_X89BGa8y1_2),.dout(w_dff_B_NMO1wSXk8_2),.clk(gclk));
	jdff dff_B_ng0dt2gY4_2(.din(w_dff_B_NMO1wSXk8_2),.dout(w_dff_B_ng0dt2gY4_2),.clk(gclk));
	jdff dff_B_gGtKYGyA7_2(.din(w_dff_B_ng0dt2gY4_2),.dout(w_dff_B_gGtKYGyA7_2),.clk(gclk));
	jdff dff_B_xs93OViw3_2(.din(w_dff_B_gGtKYGyA7_2),.dout(w_dff_B_xs93OViw3_2),.clk(gclk));
	jdff dff_B_ckgbo0At9_2(.din(w_dff_B_xs93OViw3_2),.dout(w_dff_B_ckgbo0At9_2),.clk(gclk));
	jdff dff_B_xuEFvlmC0_2(.din(w_dff_B_ckgbo0At9_2),.dout(w_dff_B_xuEFvlmC0_2),.clk(gclk));
	jdff dff_B_ysxzvZzi7_2(.din(w_dff_B_xuEFvlmC0_2),.dout(w_dff_B_ysxzvZzi7_2),.clk(gclk));
	jdff dff_B_IN8DNn2W9_2(.din(w_dff_B_ysxzvZzi7_2),.dout(w_dff_B_IN8DNn2W9_2),.clk(gclk));
	jdff dff_B_uTHUNJco7_2(.din(w_dff_B_IN8DNn2W9_2),.dout(w_dff_B_uTHUNJco7_2),.clk(gclk));
	jdff dff_B_MlXZxz3L3_2(.din(w_dff_B_uTHUNJco7_2),.dout(w_dff_B_MlXZxz3L3_2),.clk(gclk));
	jdff dff_B_YR980bIB9_2(.din(w_dff_B_MlXZxz3L3_2),.dout(w_dff_B_YR980bIB9_2),.clk(gclk));
	jdff dff_B_7xWgjYg03_2(.din(w_dff_B_YR980bIB9_2),.dout(w_dff_B_7xWgjYg03_2),.clk(gclk));
	jdff dff_B_4fxGLIjY0_2(.din(w_dff_B_7xWgjYg03_2),.dout(w_dff_B_4fxGLIjY0_2),.clk(gclk));
	jdff dff_B_ahMLwZnv2_2(.din(n1652),.dout(w_dff_B_ahMLwZnv2_2),.clk(gclk));
	jdff dff_B_DoWjBlSB7_2(.din(w_dff_B_ahMLwZnv2_2),.dout(w_dff_B_DoWjBlSB7_2),.clk(gclk));
	jdff dff_B_P2XHzwit2_2(.din(w_dff_B_DoWjBlSB7_2),.dout(w_dff_B_P2XHzwit2_2),.clk(gclk));
	jdff dff_B_luz8iKn08_2(.din(w_dff_B_P2XHzwit2_2),.dout(w_dff_B_luz8iKn08_2),.clk(gclk));
	jdff dff_B_i1p9MT3M9_2(.din(w_dff_B_luz8iKn08_2),.dout(w_dff_B_i1p9MT3M9_2),.clk(gclk));
	jdff dff_B_EGjfu9GG1_2(.din(w_dff_B_i1p9MT3M9_2),.dout(w_dff_B_EGjfu9GG1_2),.clk(gclk));
	jdff dff_B_0ZJYfDSc2_2(.din(w_dff_B_EGjfu9GG1_2),.dout(w_dff_B_0ZJYfDSc2_2),.clk(gclk));
	jdff dff_B_zL4NKhxe8_2(.din(w_dff_B_0ZJYfDSc2_2),.dout(w_dff_B_zL4NKhxe8_2),.clk(gclk));
	jdff dff_B_Ydpl4CyJ9_2(.din(w_dff_B_zL4NKhxe8_2),.dout(w_dff_B_Ydpl4CyJ9_2),.clk(gclk));
	jdff dff_B_DnFdFUol0_2(.din(w_dff_B_Ydpl4CyJ9_2),.dout(w_dff_B_DnFdFUol0_2),.clk(gclk));
	jdff dff_B_MRjghXZe9_2(.din(w_dff_B_DnFdFUol0_2),.dout(w_dff_B_MRjghXZe9_2),.clk(gclk));
	jdff dff_B_IMoRia2E5_2(.din(w_dff_B_MRjghXZe9_2),.dout(w_dff_B_IMoRia2E5_2),.clk(gclk));
	jdff dff_B_O37zx7IJ9_2(.din(w_dff_B_IMoRia2E5_2),.dout(w_dff_B_O37zx7IJ9_2),.clk(gclk));
	jdff dff_B_mst2NUll6_2(.din(w_dff_B_O37zx7IJ9_2),.dout(w_dff_B_mst2NUll6_2),.clk(gclk));
	jdff dff_B_h9AEQIZW8_2(.din(w_dff_B_mst2NUll6_2),.dout(w_dff_B_h9AEQIZW8_2),.clk(gclk));
	jdff dff_B_6pY2AjZt4_2(.din(w_dff_B_h9AEQIZW8_2),.dout(w_dff_B_6pY2AjZt4_2),.clk(gclk));
	jdff dff_B_otJtoaek1_2(.din(w_dff_B_6pY2AjZt4_2),.dout(w_dff_B_otJtoaek1_2),.clk(gclk));
	jdff dff_B_NHdx7Krz7_2(.din(w_dff_B_otJtoaek1_2),.dout(w_dff_B_NHdx7Krz7_2),.clk(gclk));
	jdff dff_B_JOO2VYIq7_2(.din(w_dff_B_NHdx7Krz7_2),.dout(w_dff_B_JOO2VYIq7_2),.clk(gclk));
	jdff dff_B_3NExsbid3_2(.din(w_dff_B_JOO2VYIq7_2),.dout(w_dff_B_3NExsbid3_2),.clk(gclk));
	jdff dff_B_Ky1UEWae1_2(.din(w_dff_B_3NExsbid3_2),.dout(w_dff_B_Ky1UEWae1_2),.clk(gclk));
	jdff dff_B_r2HUpSFV1_2(.din(w_dff_B_Ky1UEWae1_2),.dout(w_dff_B_r2HUpSFV1_2),.clk(gclk));
	jdff dff_B_Yln5KWxh8_2(.din(w_dff_B_r2HUpSFV1_2),.dout(w_dff_B_Yln5KWxh8_2),.clk(gclk));
	jdff dff_B_3U6QBMYZ3_2(.din(w_dff_B_Yln5KWxh8_2),.dout(w_dff_B_3U6QBMYZ3_2),.clk(gclk));
	jdff dff_B_15MVkSzs4_2(.din(w_dff_B_3U6QBMYZ3_2),.dout(w_dff_B_15MVkSzs4_2),.clk(gclk));
	jdff dff_B_JYu6r52R4_2(.din(w_dff_B_15MVkSzs4_2),.dout(w_dff_B_JYu6r52R4_2),.clk(gclk));
	jdff dff_B_D5NHkI6b2_2(.din(w_dff_B_JYu6r52R4_2),.dout(w_dff_B_D5NHkI6b2_2),.clk(gclk));
	jdff dff_B_cpcDl0Io7_2(.din(w_dff_B_D5NHkI6b2_2),.dout(w_dff_B_cpcDl0Io7_2),.clk(gclk));
	jdff dff_B_T2QZDKY06_2(.din(w_dff_B_cpcDl0Io7_2),.dout(w_dff_B_T2QZDKY06_2),.clk(gclk));
	jdff dff_B_e9FP3Sq65_2(.din(w_dff_B_T2QZDKY06_2),.dout(w_dff_B_e9FP3Sq65_2),.clk(gclk));
	jdff dff_B_s9AsVBm07_2(.din(w_dff_B_e9FP3Sq65_2),.dout(w_dff_B_s9AsVBm07_2),.clk(gclk));
	jdff dff_B_auyUwOzI0_2(.din(w_dff_B_s9AsVBm07_2),.dout(w_dff_B_auyUwOzI0_2),.clk(gclk));
	jdff dff_B_TZbnHOKy5_2(.din(w_dff_B_auyUwOzI0_2),.dout(w_dff_B_TZbnHOKy5_2),.clk(gclk));
	jdff dff_B_D7GJBkBS3_2(.din(w_dff_B_TZbnHOKy5_2),.dout(w_dff_B_D7GJBkBS3_2),.clk(gclk));
	jdff dff_B_Pk1qeRbR0_2(.din(w_dff_B_D7GJBkBS3_2),.dout(w_dff_B_Pk1qeRbR0_2),.clk(gclk));
	jdff dff_B_iyL8tIMv1_2(.din(w_dff_B_Pk1qeRbR0_2),.dout(w_dff_B_iyL8tIMv1_2),.clk(gclk));
	jdff dff_B_4MBxpGec8_2(.din(w_dff_B_iyL8tIMv1_2),.dout(w_dff_B_4MBxpGec8_2),.clk(gclk));
	jdff dff_B_2q3rfz6I1_2(.din(w_dff_B_4MBxpGec8_2),.dout(w_dff_B_2q3rfz6I1_2),.clk(gclk));
	jdff dff_B_NRAchYUb4_2(.din(n1651),.dout(w_dff_B_NRAchYUb4_2),.clk(gclk));
	jdff dff_B_WSfU75pS8_1(.din(n1649),.dout(w_dff_B_WSfU75pS8_1),.clk(gclk));
	jdff dff_B_9YqY937n1_2(.din(n1591),.dout(w_dff_B_9YqY937n1_2),.clk(gclk));
	jdff dff_B_TW2XgW4e9_2(.din(w_dff_B_9YqY937n1_2),.dout(w_dff_B_TW2XgW4e9_2),.clk(gclk));
	jdff dff_B_YrWW2sWS9_2(.din(w_dff_B_TW2XgW4e9_2),.dout(w_dff_B_YrWW2sWS9_2),.clk(gclk));
	jdff dff_B_BZ5ZWk8T9_2(.din(w_dff_B_YrWW2sWS9_2),.dout(w_dff_B_BZ5ZWk8T9_2),.clk(gclk));
	jdff dff_B_dK7QjaNy4_2(.din(w_dff_B_BZ5ZWk8T9_2),.dout(w_dff_B_dK7QjaNy4_2),.clk(gclk));
	jdff dff_B_b49xwTzO0_2(.din(w_dff_B_dK7QjaNy4_2),.dout(w_dff_B_b49xwTzO0_2),.clk(gclk));
	jdff dff_B_27NgSyOQ6_2(.din(w_dff_B_b49xwTzO0_2),.dout(w_dff_B_27NgSyOQ6_2),.clk(gclk));
	jdff dff_B_TNSyfA4P2_2(.din(w_dff_B_27NgSyOQ6_2),.dout(w_dff_B_TNSyfA4P2_2),.clk(gclk));
	jdff dff_B_58Ra11ci7_2(.din(w_dff_B_TNSyfA4P2_2),.dout(w_dff_B_58Ra11ci7_2),.clk(gclk));
	jdff dff_B_yvvCVGsR9_2(.din(w_dff_B_58Ra11ci7_2),.dout(w_dff_B_yvvCVGsR9_2),.clk(gclk));
	jdff dff_B_IIAeljsp1_2(.din(w_dff_B_yvvCVGsR9_2),.dout(w_dff_B_IIAeljsp1_2),.clk(gclk));
	jdff dff_B_T2OsNlBx2_2(.din(w_dff_B_IIAeljsp1_2),.dout(w_dff_B_T2OsNlBx2_2),.clk(gclk));
	jdff dff_B_IIuxMkak0_2(.din(w_dff_B_T2OsNlBx2_2),.dout(w_dff_B_IIuxMkak0_2),.clk(gclk));
	jdff dff_B_S4hAwUkp0_2(.din(w_dff_B_IIuxMkak0_2),.dout(w_dff_B_S4hAwUkp0_2),.clk(gclk));
	jdff dff_B_Xx5hVm8c0_2(.din(w_dff_B_S4hAwUkp0_2),.dout(w_dff_B_Xx5hVm8c0_2),.clk(gclk));
	jdff dff_B_q6150sBa4_2(.din(w_dff_B_Xx5hVm8c0_2),.dout(w_dff_B_q6150sBa4_2),.clk(gclk));
	jdff dff_B_gGVaxCJh9_2(.din(w_dff_B_q6150sBa4_2),.dout(w_dff_B_gGVaxCJh9_2),.clk(gclk));
	jdff dff_B_7RVl3BZv2_2(.din(w_dff_B_gGVaxCJh9_2),.dout(w_dff_B_7RVl3BZv2_2),.clk(gclk));
	jdff dff_B_u3wzTDDL2_2(.din(w_dff_B_7RVl3BZv2_2),.dout(w_dff_B_u3wzTDDL2_2),.clk(gclk));
	jdff dff_B_qz7PjDcJ2_2(.din(w_dff_B_u3wzTDDL2_2),.dout(w_dff_B_qz7PjDcJ2_2),.clk(gclk));
	jdff dff_B_8CZyNRgL3_2(.din(w_dff_B_qz7PjDcJ2_2),.dout(w_dff_B_8CZyNRgL3_2),.clk(gclk));
	jdff dff_B_2mkUKDoB5_2(.din(w_dff_B_8CZyNRgL3_2),.dout(w_dff_B_2mkUKDoB5_2),.clk(gclk));
	jdff dff_B_Ej8lV7WY5_2(.din(w_dff_B_2mkUKDoB5_2),.dout(w_dff_B_Ej8lV7WY5_2),.clk(gclk));
	jdff dff_B_AtOxWHWd8_2(.din(w_dff_B_Ej8lV7WY5_2),.dout(w_dff_B_AtOxWHWd8_2),.clk(gclk));
	jdff dff_B_cADvcp5S9_2(.din(w_dff_B_AtOxWHWd8_2),.dout(w_dff_B_cADvcp5S9_2),.clk(gclk));
	jdff dff_B_I6kc8B7O6_2(.din(w_dff_B_cADvcp5S9_2),.dout(w_dff_B_I6kc8B7O6_2),.clk(gclk));
	jdff dff_B_el5nAwQ95_2(.din(w_dff_B_I6kc8B7O6_2),.dout(w_dff_B_el5nAwQ95_2),.clk(gclk));
	jdff dff_B_1bqxx8AJ0_2(.din(w_dff_B_el5nAwQ95_2),.dout(w_dff_B_1bqxx8AJ0_2),.clk(gclk));
	jdff dff_B_xhKGldnU6_2(.din(w_dff_B_1bqxx8AJ0_2),.dout(w_dff_B_xhKGldnU6_2),.clk(gclk));
	jdff dff_B_knhMGzkE6_2(.din(w_dff_B_xhKGldnU6_2),.dout(w_dff_B_knhMGzkE6_2),.clk(gclk));
	jdff dff_B_vWwshD5o0_2(.din(w_dff_B_knhMGzkE6_2),.dout(w_dff_B_vWwshD5o0_2),.clk(gclk));
	jdff dff_B_W1Z4epbj6_2(.din(w_dff_B_vWwshD5o0_2),.dout(w_dff_B_W1Z4epbj6_2),.clk(gclk));
	jdff dff_B_BNTCPf5U2_2(.din(w_dff_B_W1Z4epbj6_2),.dout(w_dff_B_BNTCPf5U2_2),.clk(gclk));
	jdff dff_B_RdvNckQa5_2(.din(w_dff_B_BNTCPf5U2_2),.dout(w_dff_B_RdvNckQa5_2),.clk(gclk));
	jdff dff_B_8WbYio3T6_2(.din(w_dff_B_RdvNckQa5_2),.dout(w_dff_B_8WbYio3T6_2),.clk(gclk));
	jdff dff_B_wVC0Od8X5_1(.din(n1597),.dout(w_dff_B_wVC0Od8X5_1),.clk(gclk));
	jdff dff_B_p0m5Rv4t8_1(.din(w_dff_B_wVC0Od8X5_1),.dout(w_dff_B_p0m5Rv4t8_1),.clk(gclk));
	jdff dff_B_hsVj3i1c3_2(.din(n1596),.dout(w_dff_B_hsVj3i1c3_2),.clk(gclk));
	jdff dff_B_ZT0dNhtU2_2(.din(w_dff_B_hsVj3i1c3_2),.dout(w_dff_B_ZT0dNhtU2_2),.clk(gclk));
	jdff dff_B_GPC05KQe3_2(.din(w_dff_B_ZT0dNhtU2_2),.dout(w_dff_B_GPC05KQe3_2),.clk(gclk));
	jdff dff_B_BC8DyLQX1_2(.din(w_dff_B_GPC05KQe3_2),.dout(w_dff_B_BC8DyLQX1_2),.clk(gclk));
	jdff dff_B_q7KhCkDr1_2(.din(w_dff_B_BC8DyLQX1_2),.dout(w_dff_B_q7KhCkDr1_2),.clk(gclk));
	jdff dff_B_fwS1yGYl4_2(.din(w_dff_B_q7KhCkDr1_2),.dout(w_dff_B_fwS1yGYl4_2),.clk(gclk));
	jdff dff_B_J07C6Oyn3_2(.din(w_dff_B_fwS1yGYl4_2),.dout(w_dff_B_J07C6Oyn3_2),.clk(gclk));
	jdff dff_B_6oAxxxwR9_2(.din(w_dff_B_J07C6Oyn3_2),.dout(w_dff_B_6oAxxxwR9_2),.clk(gclk));
	jdff dff_B_1Gq7FYcR8_2(.din(w_dff_B_6oAxxxwR9_2),.dout(w_dff_B_1Gq7FYcR8_2),.clk(gclk));
	jdff dff_B_TEmXnqMZ0_2(.din(w_dff_B_1Gq7FYcR8_2),.dout(w_dff_B_TEmXnqMZ0_2),.clk(gclk));
	jdff dff_B_6hKH2YtQ9_2(.din(w_dff_B_TEmXnqMZ0_2),.dout(w_dff_B_6hKH2YtQ9_2),.clk(gclk));
	jdff dff_B_Z8QBaZt10_2(.din(w_dff_B_6hKH2YtQ9_2),.dout(w_dff_B_Z8QBaZt10_2),.clk(gclk));
	jdff dff_B_KkWRe1nx5_2(.din(w_dff_B_Z8QBaZt10_2),.dout(w_dff_B_KkWRe1nx5_2),.clk(gclk));
	jdff dff_B_UfwHAyvR2_2(.din(w_dff_B_KkWRe1nx5_2),.dout(w_dff_B_UfwHAyvR2_2),.clk(gclk));
	jdff dff_B_9jJtGC1b4_2(.din(w_dff_B_UfwHAyvR2_2),.dout(w_dff_B_9jJtGC1b4_2),.clk(gclk));
	jdff dff_B_ml0YPfgJ6_2(.din(w_dff_B_9jJtGC1b4_2),.dout(w_dff_B_ml0YPfgJ6_2),.clk(gclk));
	jdff dff_B_jU4cg11p9_2(.din(w_dff_B_ml0YPfgJ6_2),.dout(w_dff_B_jU4cg11p9_2),.clk(gclk));
	jdff dff_B_YJnKEkYz6_2(.din(w_dff_B_jU4cg11p9_2),.dout(w_dff_B_YJnKEkYz6_2),.clk(gclk));
	jdff dff_B_mtI54M7h6_2(.din(w_dff_B_YJnKEkYz6_2),.dout(w_dff_B_mtI54M7h6_2),.clk(gclk));
	jdff dff_B_kngdEsDq6_2(.din(w_dff_B_mtI54M7h6_2),.dout(w_dff_B_kngdEsDq6_2),.clk(gclk));
	jdff dff_B_2sg2GHlP5_2(.din(w_dff_B_kngdEsDq6_2),.dout(w_dff_B_2sg2GHlP5_2),.clk(gclk));
	jdff dff_B_8WaSW2uw4_2(.din(w_dff_B_2sg2GHlP5_2),.dout(w_dff_B_8WaSW2uw4_2),.clk(gclk));
	jdff dff_B_qH1qv8SU0_2(.din(w_dff_B_8WaSW2uw4_2),.dout(w_dff_B_qH1qv8SU0_2),.clk(gclk));
	jdff dff_B_AMlJ2WeA6_2(.din(w_dff_B_qH1qv8SU0_2),.dout(w_dff_B_AMlJ2WeA6_2),.clk(gclk));
	jdff dff_B_JvsFduZG8_2(.din(w_dff_B_AMlJ2WeA6_2),.dout(w_dff_B_JvsFduZG8_2),.clk(gclk));
	jdff dff_B_lABYoHf46_2(.din(w_dff_B_JvsFduZG8_2),.dout(w_dff_B_lABYoHf46_2),.clk(gclk));
	jdff dff_B_AkWFt7wP1_2(.din(w_dff_B_lABYoHf46_2),.dout(w_dff_B_AkWFt7wP1_2),.clk(gclk));
	jdff dff_B_JUlQF8ek7_2(.din(w_dff_B_AkWFt7wP1_2),.dout(w_dff_B_JUlQF8ek7_2),.clk(gclk));
	jdff dff_B_uicXuqRs0_2(.din(w_dff_B_JUlQF8ek7_2),.dout(w_dff_B_uicXuqRs0_2),.clk(gclk));
	jdff dff_B_KAfbg7po1_2(.din(w_dff_B_uicXuqRs0_2),.dout(w_dff_B_KAfbg7po1_2),.clk(gclk));
	jdff dff_B_E7J8dNYc1_2(.din(w_dff_B_KAfbg7po1_2),.dout(w_dff_B_E7J8dNYc1_2),.clk(gclk));
	jdff dff_B_b1k1UvD19_2(.din(w_dff_B_E7J8dNYc1_2),.dout(w_dff_B_b1k1UvD19_2),.clk(gclk));
	jdff dff_B_qzyA06vm8_2(.din(n1595),.dout(w_dff_B_qzyA06vm8_2),.clk(gclk));
	jdff dff_B_2kB1rdeo4_2(.din(w_dff_B_qzyA06vm8_2),.dout(w_dff_B_2kB1rdeo4_2),.clk(gclk));
	jdff dff_B_i3kPQFn68_2(.din(w_dff_B_2kB1rdeo4_2),.dout(w_dff_B_i3kPQFn68_2),.clk(gclk));
	jdff dff_B_rBbVVXzk3_2(.din(w_dff_B_i3kPQFn68_2),.dout(w_dff_B_rBbVVXzk3_2),.clk(gclk));
	jdff dff_B_OLMdOwMG3_2(.din(w_dff_B_rBbVVXzk3_2),.dout(w_dff_B_OLMdOwMG3_2),.clk(gclk));
	jdff dff_B_b6NPsDK31_2(.din(w_dff_B_OLMdOwMG3_2),.dout(w_dff_B_b6NPsDK31_2),.clk(gclk));
	jdff dff_B_ybw575GR9_2(.din(w_dff_B_b6NPsDK31_2),.dout(w_dff_B_ybw575GR9_2),.clk(gclk));
	jdff dff_B_dy9kZaq41_2(.din(w_dff_B_ybw575GR9_2),.dout(w_dff_B_dy9kZaq41_2),.clk(gclk));
	jdff dff_B_uwIXpi7K9_2(.din(w_dff_B_dy9kZaq41_2),.dout(w_dff_B_uwIXpi7K9_2),.clk(gclk));
	jdff dff_B_cWXnl7XS5_2(.din(w_dff_B_uwIXpi7K9_2),.dout(w_dff_B_cWXnl7XS5_2),.clk(gclk));
	jdff dff_B_KTN1cKTp9_2(.din(w_dff_B_cWXnl7XS5_2),.dout(w_dff_B_KTN1cKTp9_2),.clk(gclk));
	jdff dff_B_x1cTF8kr4_2(.din(w_dff_B_KTN1cKTp9_2),.dout(w_dff_B_x1cTF8kr4_2),.clk(gclk));
	jdff dff_B_LeIqCTrk5_2(.din(w_dff_B_x1cTF8kr4_2),.dout(w_dff_B_LeIqCTrk5_2),.clk(gclk));
	jdff dff_B_vWCYQ6mF5_2(.din(w_dff_B_LeIqCTrk5_2),.dout(w_dff_B_vWCYQ6mF5_2),.clk(gclk));
	jdff dff_B_PBmy3mMv5_2(.din(w_dff_B_vWCYQ6mF5_2),.dout(w_dff_B_PBmy3mMv5_2),.clk(gclk));
	jdff dff_B_mQBbPX3g1_2(.din(w_dff_B_PBmy3mMv5_2),.dout(w_dff_B_mQBbPX3g1_2),.clk(gclk));
	jdff dff_B_f65ZQx3T4_2(.din(w_dff_B_mQBbPX3g1_2),.dout(w_dff_B_f65ZQx3T4_2),.clk(gclk));
	jdff dff_B_czRJXl6b0_2(.din(w_dff_B_f65ZQx3T4_2),.dout(w_dff_B_czRJXl6b0_2),.clk(gclk));
	jdff dff_B_YzHV5fm95_2(.din(w_dff_B_czRJXl6b0_2),.dout(w_dff_B_YzHV5fm95_2),.clk(gclk));
	jdff dff_B_Dg4U9h9C8_2(.din(w_dff_B_YzHV5fm95_2),.dout(w_dff_B_Dg4U9h9C8_2),.clk(gclk));
	jdff dff_B_0PjPSnM23_2(.din(w_dff_B_Dg4U9h9C8_2),.dout(w_dff_B_0PjPSnM23_2),.clk(gclk));
	jdff dff_B_xJNoHB8o2_2(.din(w_dff_B_0PjPSnM23_2),.dout(w_dff_B_xJNoHB8o2_2),.clk(gclk));
	jdff dff_B_Mr35CR9c0_2(.din(w_dff_B_xJNoHB8o2_2),.dout(w_dff_B_Mr35CR9c0_2),.clk(gclk));
	jdff dff_B_zV26xBQO9_2(.din(w_dff_B_Mr35CR9c0_2),.dout(w_dff_B_zV26xBQO9_2),.clk(gclk));
	jdff dff_B_UTC1WjZF3_2(.din(w_dff_B_zV26xBQO9_2),.dout(w_dff_B_UTC1WjZF3_2),.clk(gclk));
	jdff dff_B_LA4S2oE08_2(.din(w_dff_B_UTC1WjZF3_2),.dout(w_dff_B_LA4S2oE08_2),.clk(gclk));
	jdff dff_B_fRWjaOCM8_2(.din(w_dff_B_LA4S2oE08_2),.dout(w_dff_B_fRWjaOCM8_2),.clk(gclk));
	jdff dff_B_9kTK7JHq5_2(.din(w_dff_B_fRWjaOCM8_2),.dout(w_dff_B_9kTK7JHq5_2),.clk(gclk));
	jdff dff_B_O9MgvkTA0_2(.din(w_dff_B_9kTK7JHq5_2),.dout(w_dff_B_O9MgvkTA0_2),.clk(gclk));
	jdff dff_B_TKdnRh3l9_2(.din(w_dff_B_O9MgvkTA0_2),.dout(w_dff_B_TKdnRh3l9_2),.clk(gclk));
	jdff dff_B_E6ymctXg9_2(.din(w_dff_B_TKdnRh3l9_2),.dout(w_dff_B_E6ymctXg9_2),.clk(gclk));
	jdff dff_B_09sY0hXy6_2(.din(w_dff_B_E6ymctXg9_2),.dout(w_dff_B_09sY0hXy6_2),.clk(gclk));
	jdff dff_B_5ocwuLjD9_2(.din(w_dff_B_09sY0hXy6_2),.dout(w_dff_B_5ocwuLjD9_2),.clk(gclk));
	jdff dff_B_fpEPPbdR3_2(.din(w_dff_B_5ocwuLjD9_2),.dout(w_dff_B_fpEPPbdR3_2),.clk(gclk));
	jdff dff_B_DoJLaGXc5_2(.din(n1594),.dout(w_dff_B_DoJLaGXc5_2),.clk(gclk));
	jdff dff_B_bBKY3IsN3_1(.din(n1592),.dout(w_dff_B_bBKY3IsN3_1),.clk(gclk));
	jdff dff_B_S0E1Sgjj8_2(.din(n1527),.dout(w_dff_B_S0E1Sgjj8_2),.clk(gclk));
	jdff dff_B_ihIBvree0_2(.din(w_dff_B_S0E1Sgjj8_2),.dout(w_dff_B_ihIBvree0_2),.clk(gclk));
	jdff dff_B_2iquHi9D1_2(.din(w_dff_B_ihIBvree0_2),.dout(w_dff_B_2iquHi9D1_2),.clk(gclk));
	jdff dff_B_CzZ6HtAg6_2(.din(w_dff_B_2iquHi9D1_2),.dout(w_dff_B_CzZ6HtAg6_2),.clk(gclk));
	jdff dff_B_kKufEeyC7_2(.din(w_dff_B_CzZ6HtAg6_2),.dout(w_dff_B_kKufEeyC7_2),.clk(gclk));
	jdff dff_B_yTZrpuH99_2(.din(w_dff_B_kKufEeyC7_2),.dout(w_dff_B_yTZrpuH99_2),.clk(gclk));
	jdff dff_B_Bu3Tw3l13_2(.din(w_dff_B_yTZrpuH99_2),.dout(w_dff_B_Bu3Tw3l13_2),.clk(gclk));
	jdff dff_B_M18nt3R75_2(.din(w_dff_B_Bu3Tw3l13_2),.dout(w_dff_B_M18nt3R75_2),.clk(gclk));
	jdff dff_B_D1fpOwLX2_2(.din(w_dff_B_M18nt3R75_2),.dout(w_dff_B_D1fpOwLX2_2),.clk(gclk));
	jdff dff_B_zmWh65cA3_2(.din(w_dff_B_D1fpOwLX2_2),.dout(w_dff_B_zmWh65cA3_2),.clk(gclk));
	jdff dff_B_uxgOLdre9_2(.din(w_dff_B_zmWh65cA3_2),.dout(w_dff_B_uxgOLdre9_2),.clk(gclk));
	jdff dff_B_hWPQHs9E8_2(.din(w_dff_B_uxgOLdre9_2),.dout(w_dff_B_hWPQHs9E8_2),.clk(gclk));
	jdff dff_B_HTuYlEEF3_2(.din(w_dff_B_hWPQHs9E8_2),.dout(w_dff_B_HTuYlEEF3_2),.clk(gclk));
	jdff dff_B_jrhrHsHm6_2(.din(w_dff_B_HTuYlEEF3_2),.dout(w_dff_B_jrhrHsHm6_2),.clk(gclk));
	jdff dff_B_BH59cvnu4_2(.din(w_dff_B_jrhrHsHm6_2),.dout(w_dff_B_BH59cvnu4_2),.clk(gclk));
	jdff dff_B_omuUOhtQ2_2(.din(w_dff_B_BH59cvnu4_2),.dout(w_dff_B_omuUOhtQ2_2),.clk(gclk));
	jdff dff_B_ODdj48S42_2(.din(w_dff_B_omuUOhtQ2_2),.dout(w_dff_B_ODdj48S42_2),.clk(gclk));
	jdff dff_B_kHniHcMu6_2(.din(w_dff_B_ODdj48S42_2),.dout(w_dff_B_kHniHcMu6_2),.clk(gclk));
	jdff dff_B_WqFMNQPa6_2(.din(w_dff_B_kHniHcMu6_2),.dout(w_dff_B_WqFMNQPa6_2),.clk(gclk));
	jdff dff_B_IG64Vhwe4_2(.din(w_dff_B_WqFMNQPa6_2),.dout(w_dff_B_IG64Vhwe4_2),.clk(gclk));
	jdff dff_B_FUQTqP3s7_2(.din(w_dff_B_IG64Vhwe4_2),.dout(w_dff_B_FUQTqP3s7_2),.clk(gclk));
	jdff dff_B_ppIssLh38_2(.din(w_dff_B_FUQTqP3s7_2),.dout(w_dff_B_ppIssLh38_2),.clk(gclk));
	jdff dff_B_7ujWo1wp4_2(.din(w_dff_B_ppIssLh38_2),.dout(w_dff_B_7ujWo1wp4_2),.clk(gclk));
	jdff dff_B_xnWLW3Hf4_2(.din(w_dff_B_7ujWo1wp4_2),.dout(w_dff_B_xnWLW3Hf4_2),.clk(gclk));
	jdff dff_B_wAT6RGA13_2(.din(w_dff_B_xnWLW3Hf4_2),.dout(w_dff_B_wAT6RGA13_2),.clk(gclk));
	jdff dff_B_7AnPn6AK1_2(.din(w_dff_B_wAT6RGA13_2),.dout(w_dff_B_7AnPn6AK1_2),.clk(gclk));
	jdff dff_B_cuNydATm6_2(.din(w_dff_B_7AnPn6AK1_2),.dout(w_dff_B_cuNydATm6_2),.clk(gclk));
	jdff dff_B_mry06MKl3_2(.din(w_dff_B_cuNydATm6_2),.dout(w_dff_B_mry06MKl3_2),.clk(gclk));
	jdff dff_B_B9OZct8I1_2(.din(w_dff_B_mry06MKl3_2),.dout(w_dff_B_B9OZct8I1_2),.clk(gclk));
	jdff dff_B_EVsL6J9n5_2(.din(w_dff_B_B9OZct8I1_2),.dout(w_dff_B_EVsL6J9n5_2),.clk(gclk));
	jdff dff_B_e01CU9l05_2(.din(w_dff_B_EVsL6J9n5_2),.dout(w_dff_B_e01CU9l05_2),.clk(gclk));
	jdff dff_B_dmn7JpAz0_1(.din(n1533),.dout(w_dff_B_dmn7JpAz0_1),.clk(gclk));
	jdff dff_B_4Q00MYR71_1(.din(w_dff_B_dmn7JpAz0_1),.dout(w_dff_B_4Q00MYR71_1),.clk(gclk));
	jdff dff_B_scurrzbR6_2(.din(n1532),.dout(w_dff_B_scurrzbR6_2),.clk(gclk));
	jdff dff_B_fuhby7C86_2(.din(w_dff_B_scurrzbR6_2),.dout(w_dff_B_fuhby7C86_2),.clk(gclk));
	jdff dff_B_mDgyuTP89_2(.din(w_dff_B_fuhby7C86_2),.dout(w_dff_B_mDgyuTP89_2),.clk(gclk));
	jdff dff_B_da6GawuY7_2(.din(w_dff_B_mDgyuTP89_2),.dout(w_dff_B_da6GawuY7_2),.clk(gclk));
	jdff dff_B_QXIo7UYj7_2(.din(w_dff_B_da6GawuY7_2),.dout(w_dff_B_QXIo7UYj7_2),.clk(gclk));
	jdff dff_B_KQ1pBGtY2_2(.din(w_dff_B_QXIo7UYj7_2),.dout(w_dff_B_KQ1pBGtY2_2),.clk(gclk));
	jdff dff_B_uOkudGRp9_2(.din(w_dff_B_KQ1pBGtY2_2),.dout(w_dff_B_uOkudGRp9_2),.clk(gclk));
	jdff dff_B_CzTm0Stv3_2(.din(w_dff_B_uOkudGRp9_2),.dout(w_dff_B_CzTm0Stv3_2),.clk(gclk));
	jdff dff_B_cknq3JRn7_2(.din(w_dff_B_CzTm0Stv3_2),.dout(w_dff_B_cknq3JRn7_2),.clk(gclk));
	jdff dff_B_ws6DwHoa7_2(.din(w_dff_B_cknq3JRn7_2),.dout(w_dff_B_ws6DwHoa7_2),.clk(gclk));
	jdff dff_B_EQiyyne30_2(.din(w_dff_B_ws6DwHoa7_2),.dout(w_dff_B_EQiyyne30_2),.clk(gclk));
	jdff dff_B_4Vbre3vb8_2(.din(w_dff_B_EQiyyne30_2),.dout(w_dff_B_4Vbre3vb8_2),.clk(gclk));
	jdff dff_B_qy4THqZw2_2(.din(w_dff_B_4Vbre3vb8_2),.dout(w_dff_B_qy4THqZw2_2),.clk(gclk));
	jdff dff_B_w5pch2gz4_2(.din(w_dff_B_qy4THqZw2_2),.dout(w_dff_B_w5pch2gz4_2),.clk(gclk));
	jdff dff_B_nH2gAAy46_2(.din(w_dff_B_w5pch2gz4_2),.dout(w_dff_B_nH2gAAy46_2),.clk(gclk));
	jdff dff_B_XLGlIs8w1_2(.din(w_dff_B_nH2gAAy46_2),.dout(w_dff_B_XLGlIs8w1_2),.clk(gclk));
	jdff dff_B_7R8rTkqg7_2(.din(w_dff_B_XLGlIs8w1_2),.dout(w_dff_B_7R8rTkqg7_2),.clk(gclk));
	jdff dff_B_q1b0CAl68_2(.din(w_dff_B_7R8rTkqg7_2),.dout(w_dff_B_q1b0CAl68_2),.clk(gclk));
	jdff dff_B_zPg8FF8V3_2(.din(w_dff_B_q1b0CAl68_2),.dout(w_dff_B_zPg8FF8V3_2),.clk(gclk));
	jdff dff_B_6RPAaIEA7_2(.din(w_dff_B_zPg8FF8V3_2),.dout(w_dff_B_6RPAaIEA7_2),.clk(gclk));
	jdff dff_B_XmjSXXtT9_2(.din(w_dff_B_6RPAaIEA7_2),.dout(w_dff_B_XmjSXXtT9_2),.clk(gclk));
	jdff dff_B_SccjLZju5_2(.din(w_dff_B_XmjSXXtT9_2),.dout(w_dff_B_SccjLZju5_2),.clk(gclk));
	jdff dff_B_mmlEdfil5_2(.din(w_dff_B_SccjLZju5_2),.dout(w_dff_B_mmlEdfil5_2),.clk(gclk));
	jdff dff_B_WRsAhEQ13_2(.din(w_dff_B_mmlEdfil5_2),.dout(w_dff_B_WRsAhEQ13_2),.clk(gclk));
	jdff dff_B_ENUEjEXN2_2(.din(w_dff_B_WRsAhEQ13_2),.dout(w_dff_B_ENUEjEXN2_2),.clk(gclk));
	jdff dff_B_Zf4A8C0H6_2(.din(w_dff_B_ENUEjEXN2_2),.dout(w_dff_B_Zf4A8C0H6_2),.clk(gclk));
	jdff dff_B_6MRi33Rv2_2(.din(w_dff_B_Zf4A8C0H6_2),.dout(w_dff_B_6MRi33Rv2_2),.clk(gclk));
	jdff dff_B_HTirBmXv6_2(.din(w_dff_B_6MRi33Rv2_2),.dout(w_dff_B_HTirBmXv6_2),.clk(gclk));
	jdff dff_B_9Wk412pn0_2(.din(n1531),.dout(w_dff_B_9Wk412pn0_2),.clk(gclk));
	jdff dff_B_grQkBCCC6_2(.din(w_dff_B_9Wk412pn0_2),.dout(w_dff_B_grQkBCCC6_2),.clk(gclk));
	jdff dff_B_te9FeiMN5_2(.din(w_dff_B_grQkBCCC6_2),.dout(w_dff_B_te9FeiMN5_2),.clk(gclk));
	jdff dff_B_qCGkUKpX2_2(.din(w_dff_B_te9FeiMN5_2),.dout(w_dff_B_qCGkUKpX2_2),.clk(gclk));
	jdff dff_B_fYafNUsP7_2(.din(w_dff_B_qCGkUKpX2_2),.dout(w_dff_B_fYafNUsP7_2),.clk(gclk));
	jdff dff_B_5a2WX4Mw9_2(.din(w_dff_B_fYafNUsP7_2),.dout(w_dff_B_5a2WX4Mw9_2),.clk(gclk));
	jdff dff_B_E8VE4UNc9_2(.din(w_dff_B_5a2WX4Mw9_2),.dout(w_dff_B_E8VE4UNc9_2),.clk(gclk));
	jdff dff_B_MBIVnSCj8_2(.din(w_dff_B_E8VE4UNc9_2),.dout(w_dff_B_MBIVnSCj8_2),.clk(gclk));
	jdff dff_B_2vh6456A7_2(.din(w_dff_B_MBIVnSCj8_2),.dout(w_dff_B_2vh6456A7_2),.clk(gclk));
	jdff dff_B_xngfjrw92_2(.din(w_dff_B_2vh6456A7_2),.dout(w_dff_B_xngfjrw92_2),.clk(gclk));
	jdff dff_B_1GR3noE43_2(.din(w_dff_B_xngfjrw92_2),.dout(w_dff_B_1GR3noE43_2),.clk(gclk));
	jdff dff_B_bhIN0PzF4_2(.din(w_dff_B_1GR3noE43_2),.dout(w_dff_B_bhIN0PzF4_2),.clk(gclk));
	jdff dff_B_dDvhnWjM9_2(.din(w_dff_B_bhIN0PzF4_2),.dout(w_dff_B_dDvhnWjM9_2),.clk(gclk));
	jdff dff_B_U6fTCYAX7_2(.din(w_dff_B_dDvhnWjM9_2),.dout(w_dff_B_U6fTCYAX7_2),.clk(gclk));
	jdff dff_B_JT229aKv2_2(.din(w_dff_B_U6fTCYAX7_2),.dout(w_dff_B_JT229aKv2_2),.clk(gclk));
	jdff dff_B_XvQqza6q9_2(.din(w_dff_B_JT229aKv2_2),.dout(w_dff_B_XvQqza6q9_2),.clk(gclk));
	jdff dff_B_czJwQZmA5_2(.din(w_dff_B_XvQqza6q9_2),.dout(w_dff_B_czJwQZmA5_2),.clk(gclk));
	jdff dff_B_0qeOyR0j8_2(.din(w_dff_B_czJwQZmA5_2),.dout(w_dff_B_0qeOyR0j8_2),.clk(gclk));
	jdff dff_B_VY8LuFNI5_2(.din(w_dff_B_0qeOyR0j8_2),.dout(w_dff_B_VY8LuFNI5_2),.clk(gclk));
	jdff dff_B_x6QElvNv7_2(.din(w_dff_B_VY8LuFNI5_2),.dout(w_dff_B_x6QElvNv7_2),.clk(gclk));
	jdff dff_B_I9Kzl9jC0_2(.din(w_dff_B_x6QElvNv7_2),.dout(w_dff_B_I9Kzl9jC0_2),.clk(gclk));
	jdff dff_B_rlqbqyq75_2(.din(w_dff_B_I9Kzl9jC0_2),.dout(w_dff_B_rlqbqyq75_2),.clk(gclk));
	jdff dff_B_8q8zOGDW6_2(.din(w_dff_B_rlqbqyq75_2),.dout(w_dff_B_8q8zOGDW6_2),.clk(gclk));
	jdff dff_B_iRAklezC6_2(.din(w_dff_B_8q8zOGDW6_2),.dout(w_dff_B_iRAklezC6_2),.clk(gclk));
	jdff dff_B_YXSfQCqT9_2(.din(w_dff_B_iRAklezC6_2),.dout(w_dff_B_YXSfQCqT9_2),.clk(gclk));
	jdff dff_B_8uXW4JLO6_2(.din(w_dff_B_YXSfQCqT9_2),.dout(w_dff_B_8uXW4JLO6_2),.clk(gclk));
	jdff dff_B_9VziUF1K0_2(.din(w_dff_B_8uXW4JLO6_2),.dout(w_dff_B_9VziUF1K0_2),.clk(gclk));
	jdff dff_B_sGHKFza19_2(.din(w_dff_B_9VziUF1K0_2),.dout(w_dff_B_sGHKFza19_2),.clk(gclk));
	jdff dff_B_4tJZXsBh5_2(.din(w_dff_B_sGHKFza19_2),.dout(w_dff_B_4tJZXsBh5_2),.clk(gclk));
	jdff dff_B_BLj5OV3O9_2(.din(w_dff_B_4tJZXsBh5_2),.dout(w_dff_B_BLj5OV3O9_2),.clk(gclk));
	jdff dff_B_J0E8nPgL3_2(.din(n1530),.dout(w_dff_B_J0E8nPgL3_2),.clk(gclk));
	jdff dff_B_LWNVmBBi8_1(.din(n1528),.dout(w_dff_B_LWNVmBBi8_1),.clk(gclk));
	jdff dff_B_XIF0rP9a6_2(.din(n1456),.dout(w_dff_B_XIF0rP9a6_2),.clk(gclk));
	jdff dff_B_lo71QW9n0_2(.din(w_dff_B_XIF0rP9a6_2),.dout(w_dff_B_lo71QW9n0_2),.clk(gclk));
	jdff dff_B_aEbaNfxu6_2(.din(w_dff_B_lo71QW9n0_2),.dout(w_dff_B_aEbaNfxu6_2),.clk(gclk));
	jdff dff_B_auFmes176_2(.din(w_dff_B_aEbaNfxu6_2),.dout(w_dff_B_auFmes176_2),.clk(gclk));
	jdff dff_B_74P68oUx6_2(.din(w_dff_B_auFmes176_2),.dout(w_dff_B_74P68oUx6_2),.clk(gclk));
	jdff dff_B_QPTXPFBP8_2(.din(w_dff_B_74P68oUx6_2),.dout(w_dff_B_QPTXPFBP8_2),.clk(gclk));
	jdff dff_B_Cs6xXPxZ2_2(.din(w_dff_B_QPTXPFBP8_2),.dout(w_dff_B_Cs6xXPxZ2_2),.clk(gclk));
	jdff dff_B_mRKdPi8a7_2(.din(w_dff_B_Cs6xXPxZ2_2),.dout(w_dff_B_mRKdPi8a7_2),.clk(gclk));
	jdff dff_B_Unfnpv300_2(.din(w_dff_B_mRKdPi8a7_2),.dout(w_dff_B_Unfnpv300_2),.clk(gclk));
	jdff dff_B_Nsz6DUQ24_2(.din(w_dff_B_Unfnpv300_2),.dout(w_dff_B_Nsz6DUQ24_2),.clk(gclk));
	jdff dff_B_l39oDSQO8_2(.din(w_dff_B_Nsz6DUQ24_2),.dout(w_dff_B_l39oDSQO8_2),.clk(gclk));
	jdff dff_B_fJxi8moJ3_2(.din(w_dff_B_l39oDSQO8_2),.dout(w_dff_B_fJxi8moJ3_2),.clk(gclk));
	jdff dff_B_vCFdGXyA6_2(.din(w_dff_B_fJxi8moJ3_2),.dout(w_dff_B_vCFdGXyA6_2),.clk(gclk));
	jdff dff_B_7ku762rr3_2(.din(w_dff_B_vCFdGXyA6_2),.dout(w_dff_B_7ku762rr3_2),.clk(gclk));
	jdff dff_B_1TRYjNuL0_2(.din(w_dff_B_7ku762rr3_2),.dout(w_dff_B_1TRYjNuL0_2),.clk(gclk));
	jdff dff_B_LQ5cLO5H0_2(.din(w_dff_B_1TRYjNuL0_2),.dout(w_dff_B_LQ5cLO5H0_2),.clk(gclk));
	jdff dff_B_oj15eDZ95_2(.din(w_dff_B_LQ5cLO5H0_2),.dout(w_dff_B_oj15eDZ95_2),.clk(gclk));
	jdff dff_B_jwGDfejS6_2(.din(w_dff_B_oj15eDZ95_2),.dout(w_dff_B_jwGDfejS6_2),.clk(gclk));
	jdff dff_B_gfDtRAlj2_2(.din(w_dff_B_jwGDfejS6_2),.dout(w_dff_B_gfDtRAlj2_2),.clk(gclk));
	jdff dff_B_ZyHxGm152_2(.din(w_dff_B_gfDtRAlj2_2),.dout(w_dff_B_ZyHxGm152_2),.clk(gclk));
	jdff dff_B_WmQrnVJf4_2(.din(w_dff_B_ZyHxGm152_2),.dout(w_dff_B_WmQrnVJf4_2),.clk(gclk));
	jdff dff_B_zKUzstGZ3_2(.din(w_dff_B_WmQrnVJf4_2),.dout(w_dff_B_zKUzstGZ3_2),.clk(gclk));
	jdff dff_B_DfpeIN7G4_2(.din(w_dff_B_zKUzstGZ3_2),.dout(w_dff_B_DfpeIN7G4_2),.clk(gclk));
	jdff dff_B_SLJ8rhx79_2(.din(w_dff_B_DfpeIN7G4_2),.dout(w_dff_B_SLJ8rhx79_2),.clk(gclk));
	jdff dff_B_d3ki5epJ3_2(.din(w_dff_B_SLJ8rhx79_2),.dout(w_dff_B_d3ki5epJ3_2),.clk(gclk));
	jdff dff_B_tnVmR1Is8_2(.din(w_dff_B_d3ki5epJ3_2),.dout(w_dff_B_tnVmR1Is8_2),.clk(gclk));
	jdff dff_B_jxzYtriR6_2(.din(w_dff_B_tnVmR1Is8_2),.dout(w_dff_B_jxzYtriR6_2),.clk(gclk));
	jdff dff_B_MglutVNZ3_1(.din(n1462),.dout(w_dff_B_MglutVNZ3_1),.clk(gclk));
	jdff dff_B_CzlX2EJb3_1(.din(w_dff_B_MglutVNZ3_1),.dout(w_dff_B_CzlX2EJb3_1),.clk(gclk));
	jdff dff_B_24lQ92Uj5_2(.din(n1461),.dout(w_dff_B_24lQ92Uj5_2),.clk(gclk));
	jdff dff_B_VqePKXnN5_2(.din(w_dff_B_24lQ92Uj5_2),.dout(w_dff_B_VqePKXnN5_2),.clk(gclk));
	jdff dff_B_luNLzTs68_2(.din(w_dff_B_VqePKXnN5_2),.dout(w_dff_B_luNLzTs68_2),.clk(gclk));
	jdff dff_B_CfEQACIT1_2(.din(w_dff_B_luNLzTs68_2),.dout(w_dff_B_CfEQACIT1_2),.clk(gclk));
	jdff dff_B_oU9vCJA57_2(.din(w_dff_B_CfEQACIT1_2),.dout(w_dff_B_oU9vCJA57_2),.clk(gclk));
	jdff dff_B_I5s5Yn1E4_2(.din(w_dff_B_oU9vCJA57_2),.dout(w_dff_B_I5s5Yn1E4_2),.clk(gclk));
	jdff dff_B_8DoLXLE22_2(.din(w_dff_B_I5s5Yn1E4_2),.dout(w_dff_B_8DoLXLE22_2),.clk(gclk));
	jdff dff_B_pEmF8jXS9_2(.din(w_dff_B_8DoLXLE22_2),.dout(w_dff_B_pEmF8jXS9_2),.clk(gclk));
	jdff dff_B_bAkR8X8O4_2(.din(w_dff_B_pEmF8jXS9_2),.dout(w_dff_B_bAkR8X8O4_2),.clk(gclk));
	jdff dff_B_jn9Hd0rS2_2(.din(w_dff_B_bAkR8X8O4_2),.dout(w_dff_B_jn9Hd0rS2_2),.clk(gclk));
	jdff dff_B_liOd6g2o0_2(.din(w_dff_B_jn9Hd0rS2_2),.dout(w_dff_B_liOd6g2o0_2),.clk(gclk));
	jdff dff_B_iCqlXK5G2_2(.din(w_dff_B_liOd6g2o0_2),.dout(w_dff_B_iCqlXK5G2_2),.clk(gclk));
	jdff dff_B_KYStjnHp2_2(.din(w_dff_B_iCqlXK5G2_2),.dout(w_dff_B_KYStjnHp2_2),.clk(gclk));
	jdff dff_B_svIlcXZ58_2(.din(w_dff_B_KYStjnHp2_2),.dout(w_dff_B_svIlcXZ58_2),.clk(gclk));
	jdff dff_B_ZyP1ffpY5_2(.din(w_dff_B_svIlcXZ58_2),.dout(w_dff_B_ZyP1ffpY5_2),.clk(gclk));
	jdff dff_B_iqVRy71S2_2(.din(w_dff_B_ZyP1ffpY5_2),.dout(w_dff_B_iqVRy71S2_2),.clk(gclk));
	jdff dff_B_je1NiQkl5_2(.din(w_dff_B_iqVRy71S2_2),.dout(w_dff_B_je1NiQkl5_2),.clk(gclk));
	jdff dff_B_JP53Soyp6_2(.din(w_dff_B_je1NiQkl5_2),.dout(w_dff_B_JP53Soyp6_2),.clk(gclk));
	jdff dff_B_zxRBowWI9_2(.din(w_dff_B_JP53Soyp6_2),.dout(w_dff_B_zxRBowWI9_2),.clk(gclk));
	jdff dff_B_45ysJ7Du6_2(.din(w_dff_B_zxRBowWI9_2),.dout(w_dff_B_45ysJ7Du6_2),.clk(gclk));
	jdff dff_B_QHMbO7P43_2(.din(w_dff_B_45ysJ7Du6_2),.dout(w_dff_B_QHMbO7P43_2),.clk(gclk));
	jdff dff_B_LzDVF6rA3_2(.din(w_dff_B_QHMbO7P43_2),.dout(w_dff_B_LzDVF6rA3_2),.clk(gclk));
	jdff dff_B_cFXRF5md3_2(.din(w_dff_B_LzDVF6rA3_2),.dout(w_dff_B_cFXRF5md3_2),.clk(gclk));
	jdff dff_B_20Kyx2j61_2(.din(w_dff_B_cFXRF5md3_2),.dout(w_dff_B_20Kyx2j61_2),.clk(gclk));
	jdff dff_B_92FKZmHE8_2(.din(n1460),.dout(w_dff_B_92FKZmHE8_2),.clk(gclk));
	jdff dff_B_1icfifE90_2(.din(w_dff_B_92FKZmHE8_2),.dout(w_dff_B_1icfifE90_2),.clk(gclk));
	jdff dff_B_Aem7Old88_2(.din(w_dff_B_1icfifE90_2),.dout(w_dff_B_Aem7Old88_2),.clk(gclk));
	jdff dff_B_aw4v8y6v6_2(.din(w_dff_B_Aem7Old88_2),.dout(w_dff_B_aw4v8y6v6_2),.clk(gclk));
	jdff dff_B_cQGfxCNI5_2(.din(w_dff_B_aw4v8y6v6_2),.dout(w_dff_B_cQGfxCNI5_2),.clk(gclk));
	jdff dff_B_NiD73eUP4_2(.din(w_dff_B_cQGfxCNI5_2),.dout(w_dff_B_NiD73eUP4_2),.clk(gclk));
	jdff dff_B_wKV4GvXD7_2(.din(w_dff_B_NiD73eUP4_2),.dout(w_dff_B_wKV4GvXD7_2),.clk(gclk));
	jdff dff_B_WdkR7PEB2_2(.din(w_dff_B_wKV4GvXD7_2),.dout(w_dff_B_WdkR7PEB2_2),.clk(gclk));
	jdff dff_B_3lHCz7hc8_2(.din(w_dff_B_WdkR7PEB2_2),.dout(w_dff_B_3lHCz7hc8_2),.clk(gclk));
	jdff dff_B_MDjeQiY99_2(.din(w_dff_B_3lHCz7hc8_2),.dout(w_dff_B_MDjeQiY99_2),.clk(gclk));
	jdff dff_B_I2zqQL898_2(.din(w_dff_B_MDjeQiY99_2),.dout(w_dff_B_I2zqQL898_2),.clk(gclk));
	jdff dff_B_MI3Y3TUG8_2(.din(w_dff_B_I2zqQL898_2),.dout(w_dff_B_MI3Y3TUG8_2),.clk(gclk));
	jdff dff_B_DccHJvuu3_2(.din(w_dff_B_MI3Y3TUG8_2),.dout(w_dff_B_DccHJvuu3_2),.clk(gclk));
	jdff dff_B_2Ss5OX0X1_2(.din(w_dff_B_DccHJvuu3_2),.dout(w_dff_B_2Ss5OX0X1_2),.clk(gclk));
	jdff dff_B_FtBqalmJ7_2(.din(w_dff_B_2Ss5OX0X1_2),.dout(w_dff_B_FtBqalmJ7_2),.clk(gclk));
	jdff dff_B_XqVAPHix5_2(.din(w_dff_B_FtBqalmJ7_2),.dout(w_dff_B_XqVAPHix5_2),.clk(gclk));
	jdff dff_B_ihROzAI25_2(.din(w_dff_B_XqVAPHix5_2),.dout(w_dff_B_ihROzAI25_2),.clk(gclk));
	jdff dff_B_BGrJD9gu5_2(.din(w_dff_B_ihROzAI25_2),.dout(w_dff_B_BGrJD9gu5_2),.clk(gclk));
	jdff dff_B_mZxX5Rsn6_2(.din(w_dff_B_BGrJD9gu5_2),.dout(w_dff_B_mZxX5Rsn6_2),.clk(gclk));
	jdff dff_B_srjii0rw8_2(.din(w_dff_B_mZxX5Rsn6_2),.dout(w_dff_B_srjii0rw8_2),.clk(gclk));
	jdff dff_B_DuFglYDS0_2(.din(w_dff_B_srjii0rw8_2),.dout(w_dff_B_DuFglYDS0_2),.clk(gclk));
	jdff dff_B_nAVRZE284_2(.din(w_dff_B_DuFglYDS0_2),.dout(w_dff_B_nAVRZE284_2),.clk(gclk));
	jdff dff_B_CEhV7ef81_2(.din(w_dff_B_nAVRZE284_2),.dout(w_dff_B_CEhV7ef81_2),.clk(gclk));
	jdff dff_B_wRiG9jvG0_2(.din(w_dff_B_CEhV7ef81_2),.dout(w_dff_B_wRiG9jvG0_2),.clk(gclk));
	jdff dff_B_xncYHh4L1_2(.din(w_dff_B_wRiG9jvG0_2),.dout(w_dff_B_xncYHh4L1_2),.clk(gclk));
	jdff dff_B_hYRIFJQP7_2(.din(w_dff_B_xncYHh4L1_2),.dout(w_dff_B_hYRIFJQP7_2),.clk(gclk));
	jdff dff_B_eCwWw4tB1_2(.din(n1459),.dout(w_dff_B_eCwWw4tB1_2),.clk(gclk));
	jdff dff_B_0k0xiUEN0_1(.din(n1457),.dout(w_dff_B_0k0xiUEN0_1),.clk(gclk));
	jdff dff_B_dAFThpXq4_2(.din(n1378),.dout(w_dff_B_dAFThpXq4_2),.clk(gclk));
	jdff dff_B_aXsj5ag90_2(.din(w_dff_B_dAFThpXq4_2),.dout(w_dff_B_aXsj5ag90_2),.clk(gclk));
	jdff dff_B_UjqjOdZq3_2(.din(w_dff_B_aXsj5ag90_2),.dout(w_dff_B_UjqjOdZq3_2),.clk(gclk));
	jdff dff_B_Fd2Zhzq67_2(.din(w_dff_B_UjqjOdZq3_2),.dout(w_dff_B_Fd2Zhzq67_2),.clk(gclk));
	jdff dff_B_omlmCLLu2_2(.din(w_dff_B_Fd2Zhzq67_2),.dout(w_dff_B_omlmCLLu2_2),.clk(gclk));
	jdff dff_B_G5DPJV9X7_2(.din(w_dff_B_omlmCLLu2_2),.dout(w_dff_B_G5DPJV9X7_2),.clk(gclk));
	jdff dff_B_hIU0b7953_2(.din(w_dff_B_G5DPJV9X7_2),.dout(w_dff_B_hIU0b7953_2),.clk(gclk));
	jdff dff_B_IxtO8r7g2_2(.din(w_dff_B_hIU0b7953_2),.dout(w_dff_B_IxtO8r7g2_2),.clk(gclk));
	jdff dff_B_eQnNQWVM4_2(.din(w_dff_B_IxtO8r7g2_2),.dout(w_dff_B_eQnNQWVM4_2),.clk(gclk));
	jdff dff_B_cWaK1ZaQ8_2(.din(w_dff_B_eQnNQWVM4_2),.dout(w_dff_B_cWaK1ZaQ8_2),.clk(gclk));
	jdff dff_B_uHwp6gUm2_2(.din(w_dff_B_cWaK1ZaQ8_2),.dout(w_dff_B_uHwp6gUm2_2),.clk(gclk));
	jdff dff_B_HcDL6hYO4_2(.din(w_dff_B_uHwp6gUm2_2),.dout(w_dff_B_HcDL6hYO4_2),.clk(gclk));
	jdff dff_B_6sKYNW9V3_2(.din(w_dff_B_HcDL6hYO4_2),.dout(w_dff_B_6sKYNW9V3_2),.clk(gclk));
	jdff dff_B_bPYMBBJD3_2(.din(w_dff_B_6sKYNW9V3_2),.dout(w_dff_B_bPYMBBJD3_2),.clk(gclk));
	jdff dff_B_fRCMW0K32_2(.din(w_dff_B_bPYMBBJD3_2),.dout(w_dff_B_fRCMW0K32_2),.clk(gclk));
	jdff dff_B_04kN3zBI2_2(.din(w_dff_B_fRCMW0K32_2),.dout(w_dff_B_04kN3zBI2_2),.clk(gclk));
	jdff dff_B_aT2rmnRT5_2(.din(w_dff_B_04kN3zBI2_2),.dout(w_dff_B_aT2rmnRT5_2),.clk(gclk));
	jdff dff_B_9jdbiOqK4_2(.din(w_dff_B_aT2rmnRT5_2),.dout(w_dff_B_9jdbiOqK4_2),.clk(gclk));
	jdff dff_B_H6KYvTQw7_2(.din(w_dff_B_9jdbiOqK4_2),.dout(w_dff_B_H6KYvTQw7_2),.clk(gclk));
	jdff dff_B_qZKyA1Ne3_2(.din(w_dff_B_H6KYvTQw7_2),.dout(w_dff_B_qZKyA1Ne3_2),.clk(gclk));
	jdff dff_B_OJ5jeE0E4_2(.din(w_dff_B_qZKyA1Ne3_2),.dout(w_dff_B_OJ5jeE0E4_2),.clk(gclk));
	jdff dff_B_adR5r4CT0_2(.din(w_dff_B_OJ5jeE0E4_2),.dout(w_dff_B_adR5r4CT0_2),.clk(gclk));
	jdff dff_B_1jCtZI1E6_2(.din(w_dff_B_adR5r4CT0_2),.dout(w_dff_B_1jCtZI1E6_2),.clk(gclk));
	jdff dff_B_CnGbuHTM8_1(.din(n1384),.dout(w_dff_B_CnGbuHTM8_1),.clk(gclk));
	jdff dff_B_yvVQoDbq7_1(.din(w_dff_B_CnGbuHTM8_1),.dout(w_dff_B_yvVQoDbq7_1),.clk(gclk));
	jdff dff_B_WemccfOp4_2(.din(n1383),.dout(w_dff_B_WemccfOp4_2),.clk(gclk));
	jdff dff_B_aQG8d6OU9_2(.din(w_dff_B_WemccfOp4_2),.dout(w_dff_B_aQG8d6OU9_2),.clk(gclk));
	jdff dff_B_OdQAZ9Am7_2(.din(w_dff_B_aQG8d6OU9_2),.dout(w_dff_B_OdQAZ9Am7_2),.clk(gclk));
	jdff dff_B_MB6ov2St0_2(.din(w_dff_B_OdQAZ9Am7_2),.dout(w_dff_B_MB6ov2St0_2),.clk(gclk));
	jdff dff_B_d8dcbpx88_2(.din(w_dff_B_MB6ov2St0_2),.dout(w_dff_B_d8dcbpx88_2),.clk(gclk));
	jdff dff_B_ciU02CoR8_2(.din(w_dff_B_d8dcbpx88_2),.dout(w_dff_B_ciU02CoR8_2),.clk(gclk));
	jdff dff_B_ywrgHNzR9_2(.din(w_dff_B_ciU02CoR8_2),.dout(w_dff_B_ywrgHNzR9_2),.clk(gclk));
	jdff dff_B_nstDVpDs8_2(.din(w_dff_B_ywrgHNzR9_2),.dout(w_dff_B_nstDVpDs8_2),.clk(gclk));
	jdff dff_B_wlr0YWQL8_2(.din(w_dff_B_nstDVpDs8_2),.dout(w_dff_B_wlr0YWQL8_2),.clk(gclk));
	jdff dff_B_RsW0tuP66_2(.din(w_dff_B_wlr0YWQL8_2),.dout(w_dff_B_RsW0tuP66_2),.clk(gclk));
	jdff dff_B_3p1hX5M57_2(.din(w_dff_B_RsW0tuP66_2),.dout(w_dff_B_3p1hX5M57_2),.clk(gclk));
	jdff dff_B_XYhPx7PJ1_2(.din(w_dff_B_3p1hX5M57_2),.dout(w_dff_B_XYhPx7PJ1_2),.clk(gclk));
	jdff dff_B_KsAvWhQ68_2(.din(w_dff_B_XYhPx7PJ1_2),.dout(w_dff_B_KsAvWhQ68_2),.clk(gclk));
	jdff dff_B_ZCZzxZ5k2_2(.din(w_dff_B_KsAvWhQ68_2),.dout(w_dff_B_ZCZzxZ5k2_2),.clk(gclk));
	jdff dff_B_oSPh2pBG4_2(.din(w_dff_B_ZCZzxZ5k2_2),.dout(w_dff_B_oSPh2pBG4_2),.clk(gclk));
	jdff dff_B_l9nU6ptR2_2(.din(w_dff_B_oSPh2pBG4_2),.dout(w_dff_B_l9nU6ptR2_2),.clk(gclk));
	jdff dff_B_F15NscN18_2(.din(w_dff_B_l9nU6ptR2_2),.dout(w_dff_B_F15NscN18_2),.clk(gclk));
	jdff dff_B_Wo2KnIhZ1_2(.din(w_dff_B_F15NscN18_2),.dout(w_dff_B_Wo2KnIhZ1_2),.clk(gclk));
	jdff dff_B_D9ArtEgt2_2(.din(w_dff_B_Wo2KnIhZ1_2),.dout(w_dff_B_D9ArtEgt2_2),.clk(gclk));
	jdff dff_B_1Mlva9xD5_2(.din(w_dff_B_D9ArtEgt2_2),.dout(w_dff_B_1Mlva9xD5_2),.clk(gclk));
	jdff dff_B_IPzQLyDL4_2(.din(n1382),.dout(w_dff_B_IPzQLyDL4_2),.clk(gclk));
	jdff dff_B_7Zpip4VS2_2(.din(w_dff_B_IPzQLyDL4_2),.dout(w_dff_B_7Zpip4VS2_2),.clk(gclk));
	jdff dff_B_4Vnrbr6y4_2(.din(w_dff_B_7Zpip4VS2_2),.dout(w_dff_B_4Vnrbr6y4_2),.clk(gclk));
	jdff dff_B_089zXg7m1_2(.din(w_dff_B_4Vnrbr6y4_2),.dout(w_dff_B_089zXg7m1_2),.clk(gclk));
	jdff dff_B_DLpVpjLg4_2(.din(w_dff_B_089zXg7m1_2),.dout(w_dff_B_DLpVpjLg4_2),.clk(gclk));
	jdff dff_B_6Gjf5fC50_2(.din(w_dff_B_DLpVpjLg4_2),.dout(w_dff_B_6Gjf5fC50_2),.clk(gclk));
	jdff dff_B_7qitiaO06_2(.din(w_dff_B_6Gjf5fC50_2),.dout(w_dff_B_7qitiaO06_2),.clk(gclk));
	jdff dff_B_bS2gYdg69_2(.din(w_dff_B_7qitiaO06_2),.dout(w_dff_B_bS2gYdg69_2),.clk(gclk));
	jdff dff_B_KlAJC3fs6_2(.din(w_dff_B_bS2gYdg69_2),.dout(w_dff_B_KlAJC3fs6_2),.clk(gclk));
	jdff dff_B_xvjmtu9Y6_2(.din(w_dff_B_KlAJC3fs6_2),.dout(w_dff_B_xvjmtu9Y6_2),.clk(gclk));
	jdff dff_B_lp3dBn8P0_2(.din(w_dff_B_xvjmtu9Y6_2),.dout(w_dff_B_lp3dBn8P0_2),.clk(gclk));
	jdff dff_B_iahT1t9A2_2(.din(w_dff_B_lp3dBn8P0_2),.dout(w_dff_B_iahT1t9A2_2),.clk(gclk));
	jdff dff_B_bZDlMVdR8_2(.din(w_dff_B_iahT1t9A2_2),.dout(w_dff_B_bZDlMVdR8_2),.clk(gclk));
	jdff dff_B_IbroD1ny2_2(.din(w_dff_B_bZDlMVdR8_2),.dout(w_dff_B_IbroD1ny2_2),.clk(gclk));
	jdff dff_B_MQCCYPdm0_2(.din(w_dff_B_IbroD1ny2_2),.dout(w_dff_B_MQCCYPdm0_2),.clk(gclk));
	jdff dff_B_ruqNx9nc0_2(.din(w_dff_B_MQCCYPdm0_2),.dout(w_dff_B_ruqNx9nc0_2),.clk(gclk));
	jdff dff_B_vHUPRim29_2(.din(w_dff_B_ruqNx9nc0_2),.dout(w_dff_B_vHUPRim29_2),.clk(gclk));
	jdff dff_B_yffsoico2_2(.din(w_dff_B_vHUPRim29_2),.dout(w_dff_B_yffsoico2_2),.clk(gclk));
	jdff dff_B_LIoIJQCz5_2(.din(w_dff_B_yffsoico2_2),.dout(w_dff_B_LIoIJQCz5_2),.clk(gclk));
	jdff dff_B_ch5qPKIW8_2(.din(w_dff_B_LIoIJQCz5_2),.dout(w_dff_B_ch5qPKIW8_2),.clk(gclk));
	jdff dff_B_RlL0fRtE4_2(.din(w_dff_B_ch5qPKIW8_2),.dout(w_dff_B_RlL0fRtE4_2),.clk(gclk));
	jdff dff_B_k8Ala0aO3_2(.din(w_dff_B_RlL0fRtE4_2),.dout(w_dff_B_k8Ala0aO3_2),.clk(gclk));
	jdff dff_B_Dh6JNuk36_2(.din(n1381),.dout(w_dff_B_Dh6JNuk36_2),.clk(gclk));
	jdff dff_B_qudcE3uE2_1(.din(n1379),.dout(w_dff_B_qudcE3uE2_1),.clk(gclk));
	jdff dff_B_iiRm5VJO6_2(.din(n1293),.dout(w_dff_B_iiRm5VJO6_2),.clk(gclk));
	jdff dff_B_osfoBoGh4_2(.din(w_dff_B_iiRm5VJO6_2),.dout(w_dff_B_osfoBoGh4_2),.clk(gclk));
	jdff dff_B_RNAiMMtZ9_2(.din(w_dff_B_osfoBoGh4_2),.dout(w_dff_B_RNAiMMtZ9_2),.clk(gclk));
	jdff dff_B_xn9o05H20_2(.din(w_dff_B_RNAiMMtZ9_2),.dout(w_dff_B_xn9o05H20_2),.clk(gclk));
	jdff dff_B_Nz7ycwM99_2(.din(w_dff_B_xn9o05H20_2),.dout(w_dff_B_Nz7ycwM99_2),.clk(gclk));
	jdff dff_B_EXBJhQLh2_2(.din(w_dff_B_Nz7ycwM99_2),.dout(w_dff_B_EXBJhQLh2_2),.clk(gclk));
	jdff dff_B_uoYL7YAf0_2(.din(w_dff_B_EXBJhQLh2_2),.dout(w_dff_B_uoYL7YAf0_2),.clk(gclk));
	jdff dff_B_Kc9WJSp76_2(.din(w_dff_B_uoYL7YAf0_2),.dout(w_dff_B_Kc9WJSp76_2),.clk(gclk));
	jdff dff_B_Dvx2WFBE6_2(.din(w_dff_B_Kc9WJSp76_2),.dout(w_dff_B_Dvx2WFBE6_2),.clk(gclk));
	jdff dff_B_o2JZBoql4_2(.din(w_dff_B_Dvx2WFBE6_2),.dout(w_dff_B_o2JZBoql4_2),.clk(gclk));
	jdff dff_B_ElPwNQEa3_2(.din(w_dff_B_o2JZBoql4_2),.dout(w_dff_B_ElPwNQEa3_2),.clk(gclk));
	jdff dff_B_xuNH8mrY4_2(.din(w_dff_B_ElPwNQEa3_2),.dout(w_dff_B_xuNH8mrY4_2),.clk(gclk));
	jdff dff_B_GcsqxNbq7_2(.din(w_dff_B_xuNH8mrY4_2),.dout(w_dff_B_GcsqxNbq7_2),.clk(gclk));
	jdff dff_B_mYS8SCNT5_2(.din(w_dff_B_GcsqxNbq7_2),.dout(w_dff_B_mYS8SCNT5_2),.clk(gclk));
	jdff dff_B_X7AgxXXx9_2(.din(w_dff_B_mYS8SCNT5_2),.dout(w_dff_B_X7AgxXXx9_2),.clk(gclk));
	jdff dff_B_mUIbw0n03_2(.din(w_dff_B_X7AgxXXx9_2),.dout(w_dff_B_mUIbw0n03_2),.clk(gclk));
	jdff dff_B_kmn7GrF83_2(.din(w_dff_B_mUIbw0n03_2),.dout(w_dff_B_kmn7GrF83_2),.clk(gclk));
	jdff dff_B_dye1D9Xh4_2(.din(w_dff_B_kmn7GrF83_2),.dout(w_dff_B_dye1D9Xh4_2),.clk(gclk));
	jdff dff_B_zz2U9j7y4_2(.din(w_dff_B_dye1D9Xh4_2),.dout(w_dff_B_zz2U9j7y4_2),.clk(gclk));
	jdff dff_B_hzgYHQ3m3_1(.din(n1299),.dout(w_dff_B_hzgYHQ3m3_1),.clk(gclk));
	jdff dff_B_VUJ8kK6J4_1(.din(w_dff_B_hzgYHQ3m3_1),.dout(w_dff_B_VUJ8kK6J4_1),.clk(gclk));
	jdff dff_B_XUwPFccG1_2(.din(n1298),.dout(w_dff_B_XUwPFccG1_2),.clk(gclk));
	jdff dff_B_qDf8yzvU8_2(.din(w_dff_B_XUwPFccG1_2),.dout(w_dff_B_qDf8yzvU8_2),.clk(gclk));
	jdff dff_B_YfFESv7Y2_2(.din(w_dff_B_qDf8yzvU8_2),.dout(w_dff_B_YfFESv7Y2_2),.clk(gclk));
	jdff dff_B_6hGqH0oQ4_2(.din(w_dff_B_YfFESv7Y2_2),.dout(w_dff_B_6hGqH0oQ4_2),.clk(gclk));
	jdff dff_B_meMNprm84_2(.din(w_dff_B_6hGqH0oQ4_2),.dout(w_dff_B_meMNprm84_2),.clk(gclk));
	jdff dff_B_Eaa4tlWh8_2(.din(w_dff_B_meMNprm84_2),.dout(w_dff_B_Eaa4tlWh8_2),.clk(gclk));
	jdff dff_B_KMoxkrgq0_2(.din(w_dff_B_Eaa4tlWh8_2),.dout(w_dff_B_KMoxkrgq0_2),.clk(gclk));
	jdff dff_B_Ux04TXkM2_2(.din(w_dff_B_KMoxkrgq0_2),.dout(w_dff_B_Ux04TXkM2_2),.clk(gclk));
	jdff dff_B_tGhiMtQG1_2(.din(w_dff_B_Ux04TXkM2_2),.dout(w_dff_B_tGhiMtQG1_2),.clk(gclk));
	jdff dff_B_1rwjxNxj5_2(.din(w_dff_B_tGhiMtQG1_2),.dout(w_dff_B_1rwjxNxj5_2),.clk(gclk));
	jdff dff_B_sOGu36Ju5_2(.din(w_dff_B_1rwjxNxj5_2),.dout(w_dff_B_sOGu36Ju5_2),.clk(gclk));
	jdff dff_B_cxoNxekd9_2(.din(w_dff_B_sOGu36Ju5_2),.dout(w_dff_B_cxoNxekd9_2),.clk(gclk));
	jdff dff_B_euAX7Zcr6_2(.din(w_dff_B_cxoNxekd9_2),.dout(w_dff_B_euAX7Zcr6_2),.clk(gclk));
	jdff dff_B_tSq8EBt09_2(.din(w_dff_B_euAX7Zcr6_2),.dout(w_dff_B_tSq8EBt09_2),.clk(gclk));
	jdff dff_B_6O732Ypn7_2(.din(w_dff_B_tSq8EBt09_2),.dout(w_dff_B_6O732Ypn7_2),.clk(gclk));
	jdff dff_B_q0E3ocqJ8_2(.din(w_dff_B_6O732Ypn7_2),.dout(w_dff_B_q0E3ocqJ8_2),.clk(gclk));
	jdff dff_B_r6SG1ciY6_2(.din(n1297),.dout(w_dff_B_r6SG1ciY6_2),.clk(gclk));
	jdff dff_B_oHPu7e6b0_2(.din(w_dff_B_r6SG1ciY6_2),.dout(w_dff_B_oHPu7e6b0_2),.clk(gclk));
	jdff dff_B_CwIFVtBx7_2(.din(w_dff_B_oHPu7e6b0_2),.dout(w_dff_B_CwIFVtBx7_2),.clk(gclk));
	jdff dff_B_ncpZs0IK5_2(.din(w_dff_B_CwIFVtBx7_2),.dout(w_dff_B_ncpZs0IK5_2),.clk(gclk));
	jdff dff_B_c4XT9CKg9_2(.din(w_dff_B_ncpZs0IK5_2),.dout(w_dff_B_c4XT9CKg9_2),.clk(gclk));
	jdff dff_B_mZOzL4Oo1_2(.din(w_dff_B_c4XT9CKg9_2),.dout(w_dff_B_mZOzL4Oo1_2),.clk(gclk));
	jdff dff_B_q7o620Wi1_2(.din(w_dff_B_mZOzL4Oo1_2),.dout(w_dff_B_q7o620Wi1_2),.clk(gclk));
	jdff dff_B_wzOJCRbd9_2(.din(w_dff_B_q7o620Wi1_2),.dout(w_dff_B_wzOJCRbd9_2),.clk(gclk));
	jdff dff_B_OVmNq2RK6_2(.din(w_dff_B_wzOJCRbd9_2),.dout(w_dff_B_OVmNq2RK6_2),.clk(gclk));
	jdff dff_B_2jbcJW0z1_2(.din(w_dff_B_OVmNq2RK6_2),.dout(w_dff_B_2jbcJW0z1_2),.clk(gclk));
	jdff dff_B_B1T78iHV5_2(.din(w_dff_B_2jbcJW0z1_2),.dout(w_dff_B_B1T78iHV5_2),.clk(gclk));
	jdff dff_B_yBkBYxM09_2(.din(w_dff_B_B1T78iHV5_2),.dout(w_dff_B_yBkBYxM09_2),.clk(gclk));
	jdff dff_B_1zay1wks4_2(.din(w_dff_B_yBkBYxM09_2),.dout(w_dff_B_1zay1wks4_2),.clk(gclk));
	jdff dff_B_gYPRlT7H4_2(.din(w_dff_B_1zay1wks4_2),.dout(w_dff_B_gYPRlT7H4_2),.clk(gclk));
	jdff dff_B_yY6qZYRD5_2(.din(w_dff_B_gYPRlT7H4_2),.dout(w_dff_B_yY6qZYRD5_2),.clk(gclk));
	jdff dff_B_hUt2ukSY0_2(.din(w_dff_B_yY6qZYRD5_2),.dout(w_dff_B_hUt2ukSY0_2),.clk(gclk));
	jdff dff_B_P0PV6YsP7_2(.din(w_dff_B_hUt2ukSY0_2),.dout(w_dff_B_P0PV6YsP7_2),.clk(gclk));
	jdff dff_B_l7vSSOB04_2(.din(w_dff_B_P0PV6YsP7_2),.dout(w_dff_B_l7vSSOB04_2),.clk(gclk));
	jdff dff_B_gXAYdozV7_2(.din(n1296),.dout(w_dff_B_gXAYdozV7_2),.clk(gclk));
	jdff dff_B_3kYMEyRn3_1(.din(n1294),.dout(w_dff_B_3kYMEyRn3_1),.clk(gclk));
	jdff dff_B_MWdZUw5y2_2(.din(n1203),.dout(w_dff_B_MWdZUw5y2_2),.clk(gclk));
	jdff dff_B_LqlzNphT4_2(.din(w_dff_B_MWdZUw5y2_2),.dout(w_dff_B_LqlzNphT4_2),.clk(gclk));
	jdff dff_B_nj9zwWel5_2(.din(w_dff_B_LqlzNphT4_2),.dout(w_dff_B_nj9zwWel5_2),.clk(gclk));
	jdff dff_B_hYDwZY0m3_2(.din(w_dff_B_nj9zwWel5_2),.dout(w_dff_B_hYDwZY0m3_2),.clk(gclk));
	jdff dff_B_IDqj7peY7_2(.din(w_dff_B_hYDwZY0m3_2),.dout(w_dff_B_IDqj7peY7_2),.clk(gclk));
	jdff dff_B_HQYJAkKg8_2(.din(w_dff_B_IDqj7peY7_2),.dout(w_dff_B_HQYJAkKg8_2),.clk(gclk));
	jdff dff_B_qVhPU3vs7_2(.din(w_dff_B_HQYJAkKg8_2),.dout(w_dff_B_qVhPU3vs7_2),.clk(gclk));
	jdff dff_B_mBYEv04h1_2(.din(w_dff_B_qVhPU3vs7_2),.dout(w_dff_B_mBYEv04h1_2),.clk(gclk));
	jdff dff_B_Ql9u6AKD5_2(.din(w_dff_B_mBYEv04h1_2),.dout(w_dff_B_Ql9u6AKD5_2),.clk(gclk));
	jdff dff_B_yxJc6eEw4_2(.din(w_dff_B_Ql9u6AKD5_2),.dout(w_dff_B_yxJc6eEw4_2),.clk(gclk));
	jdff dff_B_SoV47NXv2_2(.din(w_dff_B_yxJc6eEw4_2),.dout(w_dff_B_SoV47NXv2_2),.clk(gclk));
	jdff dff_B_TakxGcfK5_2(.din(w_dff_B_SoV47NXv2_2),.dout(w_dff_B_TakxGcfK5_2),.clk(gclk));
	jdff dff_B_OJf8jh5j0_2(.din(w_dff_B_TakxGcfK5_2),.dout(w_dff_B_OJf8jh5j0_2),.clk(gclk));
	jdff dff_B_hAx1BpvH7_2(.din(w_dff_B_OJf8jh5j0_2),.dout(w_dff_B_hAx1BpvH7_2),.clk(gclk));
	jdff dff_B_n8FDE26z7_2(.din(w_dff_B_hAx1BpvH7_2),.dout(w_dff_B_n8FDE26z7_2),.clk(gclk));
	jdff dff_B_DXKOYRm12_2(.din(n1208),.dout(w_dff_B_DXKOYRm12_2),.clk(gclk));
	jdff dff_B_915OFzsM2_2(.din(w_dff_B_DXKOYRm12_2),.dout(w_dff_B_915OFzsM2_2),.clk(gclk));
	jdff dff_B_Qe6BCVrA4_2(.din(w_dff_B_915OFzsM2_2),.dout(w_dff_B_Qe6BCVrA4_2),.clk(gclk));
	jdff dff_B_OwqyJRuL6_2(.din(w_dff_B_Qe6BCVrA4_2),.dout(w_dff_B_OwqyJRuL6_2),.clk(gclk));
	jdff dff_B_UYvk1XaJ9_2(.din(w_dff_B_OwqyJRuL6_2),.dout(w_dff_B_UYvk1XaJ9_2),.clk(gclk));
	jdff dff_B_63czp9M95_2(.din(w_dff_B_UYvk1XaJ9_2),.dout(w_dff_B_63czp9M95_2),.clk(gclk));
	jdff dff_B_PoIkLgfo5_2(.din(w_dff_B_63czp9M95_2),.dout(w_dff_B_PoIkLgfo5_2),.clk(gclk));
	jdff dff_B_lJSoJzUj9_2(.din(w_dff_B_PoIkLgfo5_2),.dout(w_dff_B_lJSoJzUj9_2),.clk(gclk));
	jdff dff_B_jnyN9bbn6_2(.din(w_dff_B_lJSoJzUj9_2),.dout(w_dff_B_jnyN9bbn6_2),.clk(gclk));
	jdff dff_B_VyhTxvWP0_2(.din(w_dff_B_jnyN9bbn6_2),.dout(w_dff_B_VyhTxvWP0_2),.clk(gclk));
	jdff dff_B_fJPyw12V8_2(.din(w_dff_B_VyhTxvWP0_2),.dout(w_dff_B_fJPyw12V8_2),.clk(gclk));
	jdff dff_B_TRYhdKbR3_2(.din(w_dff_B_fJPyw12V8_2),.dout(w_dff_B_TRYhdKbR3_2),.clk(gclk));
	jdff dff_B_XgHBT7UW8_2(.din(n1207),.dout(w_dff_B_XgHBT7UW8_2),.clk(gclk));
	jdff dff_B_98jFRaQa7_2(.din(w_dff_B_XgHBT7UW8_2),.dout(w_dff_B_98jFRaQa7_2),.clk(gclk));
	jdff dff_B_nE0TC1Ml7_2(.din(w_dff_B_98jFRaQa7_2),.dout(w_dff_B_nE0TC1Ml7_2),.clk(gclk));
	jdff dff_B_FGJPNzIn4_2(.din(w_dff_B_nE0TC1Ml7_2),.dout(w_dff_B_FGJPNzIn4_2),.clk(gclk));
	jdff dff_B_3faphIZx1_2(.din(w_dff_B_FGJPNzIn4_2),.dout(w_dff_B_3faphIZx1_2),.clk(gclk));
	jdff dff_B_CegCFhZV5_2(.din(w_dff_B_3faphIZx1_2),.dout(w_dff_B_CegCFhZV5_2),.clk(gclk));
	jdff dff_B_XXuOwCFI6_2(.din(w_dff_B_CegCFhZV5_2),.dout(w_dff_B_XXuOwCFI6_2),.clk(gclk));
	jdff dff_B_X4cpIIKq4_2(.din(w_dff_B_XXuOwCFI6_2),.dout(w_dff_B_X4cpIIKq4_2),.clk(gclk));
	jdff dff_B_SkwsX9Kf0_2(.din(w_dff_B_X4cpIIKq4_2),.dout(w_dff_B_SkwsX9Kf0_2),.clk(gclk));
	jdff dff_B_ZALXm2qD7_2(.din(w_dff_B_SkwsX9Kf0_2),.dout(w_dff_B_ZALXm2qD7_2),.clk(gclk));
	jdff dff_B_wisMNCrq6_2(.din(w_dff_B_ZALXm2qD7_2),.dout(w_dff_B_wisMNCrq6_2),.clk(gclk));
	jdff dff_B_fmfsgtvM9_2(.din(w_dff_B_wisMNCrq6_2),.dout(w_dff_B_fmfsgtvM9_2),.clk(gclk));
	jdff dff_B_WtDL9gqU3_2(.din(w_dff_B_fmfsgtvM9_2),.dout(w_dff_B_WtDL9gqU3_2),.clk(gclk));
	jdff dff_B_Xn6nswdx1_2(.din(w_dff_B_WtDL9gqU3_2),.dout(w_dff_B_Xn6nswdx1_2),.clk(gclk));
	jdff dff_B_ZkUGvUdg8_2(.din(n1206),.dout(w_dff_B_ZkUGvUdg8_2),.clk(gclk));
	jdff dff_B_XdgiEJGx6_1(.din(n1204),.dout(w_dff_B_XdgiEJGx6_1),.clk(gclk));
	jdff dff_B_8ojOxZMk7_2(.din(n1099),.dout(w_dff_B_8ojOxZMk7_2),.clk(gclk));
	jdff dff_B_KHBwC0mO7_2(.din(w_dff_B_8ojOxZMk7_2),.dout(w_dff_B_KHBwC0mO7_2),.clk(gclk));
	jdff dff_B_L9tymt2o7_2(.din(w_dff_B_KHBwC0mO7_2),.dout(w_dff_B_L9tymt2o7_2),.clk(gclk));
	jdff dff_B_gCEoc0ok0_2(.din(w_dff_B_L9tymt2o7_2),.dout(w_dff_B_gCEoc0ok0_2),.clk(gclk));
	jdff dff_B_MPxCxC8F7_2(.din(w_dff_B_gCEoc0ok0_2),.dout(w_dff_B_MPxCxC8F7_2),.clk(gclk));
	jdff dff_B_GkVu1s132_2(.din(w_dff_B_MPxCxC8F7_2),.dout(w_dff_B_GkVu1s132_2),.clk(gclk));
	jdff dff_B_81nsxWVJ6_2(.din(w_dff_B_GkVu1s132_2),.dout(w_dff_B_81nsxWVJ6_2),.clk(gclk));
	jdff dff_B_xftHJnTj0_2(.din(w_dff_B_81nsxWVJ6_2),.dout(w_dff_B_xftHJnTj0_2),.clk(gclk));
	jdff dff_B_jdfI6LIz8_2(.din(w_dff_B_xftHJnTj0_2),.dout(w_dff_B_jdfI6LIz8_2),.clk(gclk));
	jdff dff_B_WuLqmkvo0_2(.din(w_dff_B_jdfI6LIz8_2),.dout(w_dff_B_WuLqmkvo0_2),.clk(gclk));
	jdff dff_B_ZwivAUV38_2(.din(w_dff_B_WuLqmkvo0_2),.dout(w_dff_B_ZwivAUV38_2),.clk(gclk));
	jdff dff_A_XIjrmA6j7_0(.dout(w_n1110_0[0]),.din(w_dff_A_XIjrmA6j7_0),.clk(gclk));
	jdff dff_A_RnJEbFAG9_0(.dout(w_dff_A_XIjrmA6j7_0),.din(w_dff_A_RnJEbFAG9_0),.clk(gclk));
	jdff dff_A_QejrMFgQ1_0(.dout(w_dff_A_RnJEbFAG9_0),.din(w_dff_A_QejrMFgQ1_0),.clk(gclk));
	jdff dff_B_BWx1odqe4_2(.din(n1110),.dout(w_dff_B_BWx1odqe4_2),.clk(gclk));
	jdff dff_B_hLKPFkcp0_1(.din(n1104),.dout(w_dff_B_hLKPFkcp0_1),.clk(gclk));
	jdff dff_B_WKbR0yNr9_1(.din(w_dff_B_hLKPFkcp0_1),.dout(w_dff_B_WKbR0yNr9_1),.clk(gclk));
	jdff dff_B_2L9qJ39V7_1(.din(w_dff_B_WKbR0yNr9_1),.dout(w_dff_B_2L9qJ39V7_1),.clk(gclk));
	jdff dff_B_QyGA5kwr6_1(.din(w_dff_B_2L9qJ39V7_1),.dout(w_dff_B_QyGA5kwr6_1),.clk(gclk));
	jdff dff_B_2ajsOZOZ6_1(.din(w_dff_B_QyGA5kwr6_1),.dout(w_dff_B_2ajsOZOZ6_1),.clk(gclk));
	jdff dff_B_Ey840Zsi9_1(.din(w_dff_B_2ajsOZOZ6_1),.dout(w_dff_B_Ey840Zsi9_1),.clk(gclk));
	jdff dff_B_lNYAzxww7_1(.din(n1105),.dout(w_dff_B_lNYAzxww7_1),.clk(gclk));
	jdff dff_B_bNAI5svb2_1(.din(w_dff_B_lNYAzxww7_1),.dout(w_dff_B_bNAI5svb2_1),.clk(gclk));
	jdff dff_A_mVit9xwJ2_1(.dout(w_G307gat_2[1]),.din(w_dff_A_mVit9xwJ2_1),.clk(gclk));
	jdff dff_A_AZd2pNcg9_1(.dout(w_dff_A_mVit9xwJ2_1),.din(w_dff_A_AZd2pNcg9_1),.clk(gclk));
	jdff dff_A_ZYScIdGK7_1(.dout(w_dff_A_AZd2pNcg9_1),.din(w_dff_A_ZYScIdGK7_1),.clk(gclk));
	jdff dff_A_RuE7Rnip8_1(.dout(w_dff_A_ZYScIdGK7_1),.din(w_dff_A_RuE7Rnip8_1),.clk(gclk));
	jdff dff_A_1rfP5BYn6_1(.dout(w_dff_A_RuE7Rnip8_1),.din(w_dff_A_1rfP5BYn6_1),.clk(gclk));
	jdff dff_A_j2WdFBsr8_1(.dout(w_dff_A_1rfP5BYn6_1),.din(w_dff_A_j2WdFBsr8_1),.clk(gclk));
	jdff dff_A_x4eBRqMp2_1(.dout(w_dff_A_j2WdFBsr8_1),.din(w_dff_A_x4eBRqMp2_1),.clk(gclk));
	jdff dff_B_OdCm1bZC7_2(.din(n1103),.dout(w_dff_B_OdCm1bZC7_2),.clk(gclk));
	jdff dff_B_yuwvpGbi1_2(.din(w_dff_B_OdCm1bZC7_2),.dout(w_dff_B_yuwvpGbi1_2),.clk(gclk));
	jdff dff_B_CrfCmex16_2(.din(w_dff_B_yuwvpGbi1_2),.dout(w_dff_B_CrfCmex16_2),.clk(gclk));
	jdff dff_B_SLp8eusp2_2(.din(w_dff_B_CrfCmex16_2),.dout(w_dff_B_SLp8eusp2_2),.clk(gclk));
	jdff dff_B_9k9VjoeR7_2(.din(w_dff_B_SLp8eusp2_2),.dout(w_dff_B_9k9VjoeR7_2),.clk(gclk));
	jdff dff_B_1LKT2Gyp5_2(.din(w_dff_B_9k9VjoeR7_2),.dout(w_dff_B_1LKT2Gyp5_2),.clk(gclk));
	jdff dff_B_70ZJ2Mv85_2(.din(w_dff_B_1LKT2Gyp5_2),.dout(w_dff_B_70ZJ2Mv85_2),.clk(gclk));
	jdff dff_B_B9mgERzy1_2(.din(w_dff_B_70ZJ2Mv85_2),.dout(w_dff_B_B9mgERzy1_2),.clk(gclk));
	jdff dff_B_HO2IAvlh3_2(.din(w_dff_B_B9mgERzy1_2),.dout(w_dff_B_HO2IAvlh3_2),.clk(gclk));
	jdff dff_B_hwGPVRFa1_2(.din(w_dff_B_HO2IAvlh3_2),.dout(w_dff_B_hwGPVRFa1_2),.clk(gclk));
	jdff dff_B_dGU27aM66_1(.din(n1100),.dout(w_dff_B_dGU27aM66_1),.clk(gclk));
	jdff dff_B_4bTIsIFD2_2(.din(n1001),.dout(w_dff_B_4bTIsIFD2_2),.clk(gclk));
	jdff dff_B_63rqYGLh9_2(.din(w_dff_B_4bTIsIFD2_2),.dout(w_dff_B_63rqYGLh9_2),.clk(gclk));
	jdff dff_B_TEqF3pxj1_2(.din(w_dff_B_63rqYGLh9_2),.dout(w_dff_B_TEqF3pxj1_2),.clk(gclk));
	jdff dff_B_6SuRuAjx5_2(.din(w_dff_B_TEqF3pxj1_2),.dout(w_dff_B_6SuRuAjx5_2),.clk(gclk));
	jdff dff_B_yEBdZkIb7_2(.din(w_dff_B_6SuRuAjx5_2),.dout(w_dff_B_yEBdZkIb7_2),.clk(gclk));
	jdff dff_B_XFdW4tmv0_2(.din(w_dff_B_yEBdZkIb7_2),.dout(w_dff_B_XFdW4tmv0_2),.clk(gclk));
	jdff dff_B_DOlnnmWH3_2(.din(w_dff_B_XFdW4tmv0_2),.dout(w_dff_B_DOlnnmWH3_2),.clk(gclk));
	jdff dff_B_fFN9NgEZ6_2(.din(w_dff_B_DOlnnmWH3_2),.dout(w_dff_B_fFN9NgEZ6_2),.clk(gclk));
	jdff dff_B_EqFFoG9E7_2(.din(n1010),.dout(w_dff_B_EqFFoG9E7_2),.clk(gclk));
	jdff dff_B_gh7giJJg6_2(.din(w_dff_B_EqFFoG9E7_2),.dout(w_dff_B_gh7giJJg6_2),.clk(gclk));
	jdff dff_B_CPHW86HD7_2(.din(w_dff_B_gh7giJJg6_2),.dout(w_dff_B_CPHW86HD7_2),.clk(gclk));
	jdff dff_B_dgeRzY9T7_2(.din(w_dff_B_CPHW86HD7_2),.dout(w_dff_B_dgeRzY9T7_2),.clk(gclk));
	jdff dff_B_WsuEKtQ94_2(.din(w_dff_B_dgeRzY9T7_2),.dout(w_dff_B_WsuEKtQ94_2),.clk(gclk));
	jdff dff_A_QAVTmnh25_0(.dout(w_n1008_0[0]),.din(w_dff_A_QAVTmnh25_0),.clk(gclk));
	jdff dff_A_uvHSWtwa2_0(.dout(w_dff_A_QAVTmnh25_0),.din(w_dff_A_uvHSWtwa2_0),.clk(gclk));
	jdff dff_A_N9UzwRK64_0(.dout(w_dff_A_uvHSWtwa2_0),.din(w_dff_A_N9UzwRK64_0),.clk(gclk));
	jdff dff_A_t44wiNYu7_0(.dout(w_n793_0[0]),.din(w_dff_A_t44wiNYu7_0),.clk(gclk));
	jdff dff_A_QHOwzUSP9_1(.dout(w_n1006_0[1]),.din(w_dff_A_QHOwzUSP9_1),.clk(gclk));
	jdff dff_A_3cWmQLSM5_1(.dout(w_dff_A_QHOwzUSP9_1),.din(w_dff_A_3cWmQLSM5_1),.clk(gclk));
	jdff dff_B_hDAG1rPw4_1(.din(n1002),.dout(w_dff_B_hDAG1rPw4_1),.clk(gclk));
	jdff dff_B_ivgsdJ9S8_1(.din(w_dff_B_hDAG1rPw4_1),.dout(w_dff_B_ivgsdJ9S8_1),.clk(gclk));
	jdff dff_B_Y0XRAVZb6_1(.din(w_dff_B_ivgsdJ9S8_1),.dout(w_dff_B_Y0XRAVZb6_1),.clk(gclk));
	jdff dff_B_debJB5Lr6_1(.din(w_dff_B_Y0XRAVZb6_1),.dout(w_dff_B_debJB5Lr6_1),.clk(gclk));
	jdff dff_B_EWZpWhAQ7_1(.din(w_dff_B_debJB5Lr6_1),.dout(w_dff_B_EWZpWhAQ7_1),.clk(gclk));
	jdff dff_A_l0fFdRyQ1_0(.dout(w_n903_0[0]),.din(w_dff_A_l0fFdRyQ1_0),.clk(gclk));
	jdff dff_A_EHBpv6gX8_0(.dout(w_dff_A_l0fFdRyQ1_0),.din(w_dff_A_EHBpv6gX8_0),.clk(gclk));
	jdff dff_A_UYrp90wJ3_0(.dout(w_dff_A_EHBpv6gX8_0),.din(w_dff_A_UYrp90wJ3_0),.clk(gclk));
	jdff dff_A_H5gxb2DF1_0(.dout(w_n695_0[0]),.din(w_dff_A_H5gxb2DF1_0),.clk(gclk));
	jdff dff_A_zqS5QNMI5_0(.dout(w_dff_A_H5gxb2DF1_0),.din(w_dff_A_zqS5QNMI5_0),.clk(gclk));
	jdff dff_A_WbOULxLr1_0(.dout(w_dff_A_zqS5QNMI5_0),.din(w_dff_A_WbOULxLr1_0),.clk(gclk));
	jdff dff_B_Ycy7sUPW7_2(.din(n898),.dout(w_dff_B_Ycy7sUPW7_2),.clk(gclk));
	jdff dff_A_3d3NyK4D6_1(.dout(w_n896_0[1]),.din(w_dff_A_3d3NyK4D6_1),.clk(gclk));
	jdff dff_A_GAtiqGUf0_1(.dout(w_dff_A_3d3NyK4D6_1),.din(w_dff_A_GAtiqGUf0_1),.clk(gclk));
	jdff dff_A_Rese1iCp1_1(.dout(w_dff_A_GAtiqGUf0_1),.din(w_dff_A_Rese1iCp1_1),.clk(gclk));
	jdff dff_A_L2EGjFho3_1(.dout(w_dff_A_Rese1iCp1_1),.din(w_dff_A_L2EGjFho3_1),.clk(gclk));
	jdff dff_A_QgymNIau6_1(.dout(w_dff_A_L2EGjFho3_1),.din(w_dff_A_QgymNIau6_1),.clk(gclk));
	jdff dff_A_qLYUvskc7_1(.dout(w_dff_A_sPfUjL1l8_0),.din(w_dff_A_qLYUvskc7_1),.clk(gclk));
	jdff dff_A_sPfUjL1l8_0(.dout(w_dff_A_NE2GPuAv3_0),.din(w_dff_A_sPfUjL1l8_0),.clk(gclk));
	jdff dff_A_NE2GPuAv3_0(.dout(w_dff_A_PShVza2c8_0),.din(w_dff_A_NE2GPuAv3_0),.clk(gclk));
	jdff dff_A_PShVza2c8_0(.dout(w_dff_A_0zm7ulG42_0),.din(w_dff_A_PShVza2c8_0),.clk(gclk));
	jdff dff_A_0zm7ulG42_0(.dout(w_dff_A_j5VviUPL2_0),.din(w_dff_A_0zm7ulG42_0),.clk(gclk));
	jdff dff_A_j5VviUPL2_0(.dout(w_dff_A_tTC9FYLk4_0),.din(w_dff_A_j5VviUPL2_0),.clk(gclk));
	jdff dff_A_tTC9FYLk4_0(.dout(w_dff_A_eAwVwr0k7_0),.din(w_dff_A_tTC9FYLk4_0),.clk(gclk));
	jdff dff_A_eAwVwr0k7_0(.dout(w_dff_A_74UJSTH11_0),.din(w_dff_A_eAwVwr0k7_0),.clk(gclk));
	jdff dff_A_74UJSTH11_0(.dout(w_dff_A_64C90BHz5_0),.din(w_dff_A_74UJSTH11_0),.clk(gclk));
	jdff dff_A_64C90BHz5_0(.dout(w_dff_A_mrCsYqBD2_0),.din(w_dff_A_64C90BHz5_0),.clk(gclk));
	jdff dff_A_mrCsYqBD2_0(.dout(w_dff_A_ol9UgZWG4_0),.din(w_dff_A_mrCsYqBD2_0),.clk(gclk));
	jdff dff_A_ol9UgZWG4_0(.dout(w_dff_A_9flp1qGQ0_0),.din(w_dff_A_ol9UgZWG4_0),.clk(gclk));
	jdff dff_A_9flp1qGQ0_0(.dout(w_dff_A_t283ZKbl5_0),.din(w_dff_A_9flp1qGQ0_0),.clk(gclk));
	jdff dff_A_t283ZKbl5_0(.dout(w_dff_A_Ha7xGOky4_0),.din(w_dff_A_t283ZKbl5_0),.clk(gclk));
	jdff dff_A_Ha7xGOky4_0(.dout(w_dff_A_6uhpB0TI7_0),.din(w_dff_A_Ha7xGOky4_0),.clk(gclk));
	jdff dff_A_6uhpB0TI7_0(.dout(w_dff_A_FvP308hJ6_0),.din(w_dff_A_6uhpB0TI7_0),.clk(gclk));
	jdff dff_A_FvP308hJ6_0(.dout(w_dff_A_1ibXjjTB8_0),.din(w_dff_A_FvP308hJ6_0),.clk(gclk));
	jdff dff_A_1ibXjjTB8_0(.dout(w_dff_A_C57Ap0IH4_0),.din(w_dff_A_1ibXjjTB8_0),.clk(gclk));
	jdff dff_A_C57Ap0IH4_0(.dout(w_dff_A_Q46xReL81_0),.din(w_dff_A_C57Ap0IH4_0),.clk(gclk));
	jdff dff_A_Q46xReL81_0(.dout(w_dff_A_GwArLYlx8_0),.din(w_dff_A_Q46xReL81_0),.clk(gclk));
	jdff dff_A_GwArLYlx8_0(.dout(w_dff_A_j4xyXNnf3_0),.din(w_dff_A_GwArLYlx8_0),.clk(gclk));
	jdff dff_A_j4xyXNnf3_0(.dout(w_dff_A_7ISzBbUm8_0),.din(w_dff_A_j4xyXNnf3_0),.clk(gclk));
	jdff dff_A_7ISzBbUm8_0(.dout(w_dff_A_NRZdd1iT2_0),.din(w_dff_A_7ISzBbUm8_0),.clk(gclk));
	jdff dff_A_NRZdd1iT2_0(.dout(w_dff_A_oxjuRczw8_0),.din(w_dff_A_NRZdd1iT2_0),.clk(gclk));
	jdff dff_A_oxjuRczw8_0(.dout(w_dff_A_HH0UcsaP7_0),.din(w_dff_A_oxjuRczw8_0),.clk(gclk));
	jdff dff_A_HH0UcsaP7_0(.dout(w_dff_A_Jy3zRvlp3_0),.din(w_dff_A_HH0UcsaP7_0),.clk(gclk));
	jdff dff_A_Jy3zRvlp3_0(.dout(w_dff_A_ja392aA08_0),.din(w_dff_A_Jy3zRvlp3_0),.clk(gclk));
	jdff dff_A_ja392aA08_0(.dout(w_dff_A_7QTZYZG49_0),.din(w_dff_A_ja392aA08_0),.clk(gclk));
	jdff dff_A_7QTZYZG49_0(.dout(w_dff_A_kjOKyZAa7_0),.din(w_dff_A_7QTZYZG49_0),.clk(gclk));
	jdff dff_A_kjOKyZAa7_0(.dout(w_dff_A_jb79drfl2_0),.din(w_dff_A_kjOKyZAa7_0),.clk(gclk));
	jdff dff_A_jb79drfl2_0(.dout(w_dff_A_dkvrzT458_0),.din(w_dff_A_jb79drfl2_0),.clk(gclk));
	jdff dff_A_dkvrzT458_0(.dout(w_dff_A_qkk441TT3_0),.din(w_dff_A_dkvrzT458_0),.clk(gclk));
	jdff dff_A_qkk441TT3_0(.dout(w_dff_A_yWZ5wtNx4_0),.din(w_dff_A_qkk441TT3_0),.clk(gclk));
	jdff dff_A_yWZ5wtNx4_0(.dout(w_dff_A_yUhV3XZu0_0),.din(w_dff_A_yWZ5wtNx4_0),.clk(gclk));
	jdff dff_A_yUhV3XZu0_0(.dout(w_dff_A_T8KygEKp3_0),.din(w_dff_A_yUhV3XZu0_0),.clk(gclk));
	jdff dff_A_T8KygEKp3_0(.dout(w_dff_A_QZHR3Mel1_0),.din(w_dff_A_T8KygEKp3_0),.clk(gclk));
	jdff dff_A_QZHR3Mel1_0(.dout(w_dff_A_5Xdqzr8V9_0),.din(w_dff_A_QZHR3Mel1_0),.clk(gclk));
	jdff dff_A_5Xdqzr8V9_0(.dout(w_dff_A_GcQnaqOF9_0),.din(w_dff_A_5Xdqzr8V9_0),.clk(gclk));
	jdff dff_A_GcQnaqOF9_0(.dout(w_dff_A_AW643vpz2_0),.din(w_dff_A_GcQnaqOF9_0),.clk(gclk));
	jdff dff_A_AW643vpz2_0(.dout(w_dff_A_BOEsfZn71_0),.din(w_dff_A_AW643vpz2_0),.clk(gclk));
	jdff dff_A_BOEsfZn71_0(.dout(w_dff_A_quydwrrO7_0),.din(w_dff_A_BOEsfZn71_0),.clk(gclk));
	jdff dff_A_quydwrrO7_0(.dout(w_dff_A_lXfelNFT5_0),.din(w_dff_A_quydwrrO7_0),.clk(gclk));
	jdff dff_A_lXfelNFT5_0(.dout(w_dff_A_Manmdn8F2_0),.din(w_dff_A_lXfelNFT5_0),.clk(gclk));
	jdff dff_A_Manmdn8F2_0(.dout(w_dff_A_Xuv4eNEh6_0),.din(w_dff_A_Manmdn8F2_0),.clk(gclk));
	jdff dff_A_Xuv4eNEh6_0(.dout(w_dff_A_mj5JHtcG4_0),.din(w_dff_A_Xuv4eNEh6_0),.clk(gclk));
	jdff dff_A_mj5JHtcG4_0(.dout(w_dff_A_lr5i5jJ84_0),.din(w_dff_A_mj5JHtcG4_0),.clk(gclk));
	jdff dff_A_lr5i5jJ84_0(.dout(w_dff_A_0g0SfOiE8_0),.din(w_dff_A_lr5i5jJ84_0),.clk(gclk));
	jdff dff_A_0g0SfOiE8_0(.dout(w_dff_A_nuRitZCD0_0),.din(w_dff_A_0g0SfOiE8_0),.clk(gclk));
	jdff dff_A_nuRitZCD0_0(.dout(w_dff_A_kAkSPkP93_0),.din(w_dff_A_nuRitZCD0_0),.clk(gclk));
	jdff dff_A_kAkSPkP93_0(.dout(w_dff_A_Up5xdlKm4_0),.din(w_dff_A_kAkSPkP93_0),.clk(gclk));
	jdff dff_A_Up5xdlKm4_0(.dout(w_dff_A_d5qXlybP4_0),.din(w_dff_A_Up5xdlKm4_0),.clk(gclk));
	jdff dff_A_d5qXlybP4_0(.dout(w_dff_A_mHEjEAwr8_0),.din(w_dff_A_d5qXlybP4_0),.clk(gclk));
	jdff dff_A_mHEjEAwr8_0(.dout(w_dff_A_wiBrkzwd7_0),.din(w_dff_A_mHEjEAwr8_0),.clk(gclk));
	jdff dff_A_wiBrkzwd7_0(.dout(w_dff_A_QiXHZho40_0),.din(w_dff_A_wiBrkzwd7_0),.clk(gclk));
	jdff dff_A_QiXHZho40_0(.dout(w_dff_A_twFiy3y93_0),.din(w_dff_A_QiXHZho40_0),.clk(gclk));
	jdff dff_A_twFiy3y93_0(.dout(w_dff_A_qcCVN0BH5_0),.din(w_dff_A_twFiy3y93_0),.clk(gclk));
	jdff dff_A_qcCVN0BH5_0(.dout(w_dff_A_SlszP6vW7_0),.din(w_dff_A_qcCVN0BH5_0),.clk(gclk));
	jdff dff_A_SlszP6vW7_0(.dout(w_dff_A_78x6wCWu6_0),.din(w_dff_A_SlszP6vW7_0),.clk(gclk));
	jdff dff_A_78x6wCWu6_0(.dout(w_dff_A_3lSMzqo55_0),.din(w_dff_A_78x6wCWu6_0),.clk(gclk));
	jdff dff_A_3lSMzqo55_0(.dout(w_dff_A_BLmCA7UH9_0),.din(w_dff_A_3lSMzqo55_0),.clk(gclk));
	jdff dff_A_BLmCA7UH9_0(.dout(w_dff_A_uZLHxEEa3_0),.din(w_dff_A_BLmCA7UH9_0),.clk(gclk));
	jdff dff_A_uZLHxEEa3_0(.dout(w_dff_A_FSmdya4s2_0),.din(w_dff_A_uZLHxEEa3_0),.clk(gclk));
	jdff dff_A_FSmdya4s2_0(.dout(w_dff_A_nyYDZOFl4_0),.din(w_dff_A_FSmdya4s2_0),.clk(gclk));
	jdff dff_A_nyYDZOFl4_0(.dout(w_dff_A_q6O22de35_0),.din(w_dff_A_nyYDZOFl4_0),.clk(gclk));
	jdff dff_A_q6O22de35_0(.dout(w_dff_A_hAS4SyhA4_0),.din(w_dff_A_q6O22de35_0),.clk(gclk));
	jdff dff_A_hAS4SyhA4_0(.dout(w_dff_A_eDbKs2iV5_0),.din(w_dff_A_hAS4SyhA4_0),.clk(gclk));
	jdff dff_A_eDbKs2iV5_0(.dout(w_dff_A_ozHjHBjO1_0),.din(w_dff_A_eDbKs2iV5_0),.clk(gclk));
	jdff dff_A_ozHjHBjO1_0(.dout(w_dff_A_aRO1PoMv3_0),.din(w_dff_A_ozHjHBjO1_0),.clk(gclk));
	jdff dff_A_aRO1PoMv3_0(.dout(w_dff_A_iSJBwK9L3_0),.din(w_dff_A_aRO1PoMv3_0),.clk(gclk));
	jdff dff_A_iSJBwK9L3_0(.dout(w_dff_A_c7m5qKbU6_0),.din(w_dff_A_iSJBwK9L3_0),.clk(gclk));
	jdff dff_A_c7m5qKbU6_0(.dout(w_dff_A_mWuGthc55_0),.din(w_dff_A_c7m5qKbU6_0),.clk(gclk));
	jdff dff_A_mWuGthc55_0(.dout(w_dff_A_OStBu9fY9_0),.din(w_dff_A_mWuGthc55_0),.clk(gclk));
	jdff dff_A_OStBu9fY9_0(.dout(w_dff_A_yTWRKoSS5_0),.din(w_dff_A_OStBu9fY9_0),.clk(gclk));
	jdff dff_A_yTWRKoSS5_0(.dout(w_dff_A_cGgknGSv6_0),.din(w_dff_A_yTWRKoSS5_0),.clk(gclk));
	jdff dff_A_cGgknGSv6_0(.dout(G545gat),.din(w_dff_A_cGgknGSv6_0),.clk(gclk));
	jdff dff_A_oHlkIbp78_2(.dout(w_dff_A_Ioca4err9_0),.din(w_dff_A_oHlkIbp78_2),.clk(gclk));
	jdff dff_A_Ioca4err9_0(.dout(w_dff_A_lpOZ5Fvf1_0),.din(w_dff_A_Ioca4err9_0),.clk(gclk));
	jdff dff_A_lpOZ5Fvf1_0(.dout(w_dff_A_LFXldfUV3_0),.din(w_dff_A_lpOZ5Fvf1_0),.clk(gclk));
	jdff dff_A_LFXldfUV3_0(.dout(w_dff_A_xOJhOIUo9_0),.din(w_dff_A_LFXldfUV3_0),.clk(gclk));
	jdff dff_A_xOJhOIUo9_0(.dout(w_dff_A_j22KwikW4_0),.din(w_dff_A_xOJhOIUo9_0),.clk(gclk));
	jdff dff_A_j22KwikW4_0(.dout(w_dff_A_pfopnZP06_0),.din(w_dff_A_j22KwikW4_0),.clk(gclk));
	jdff dff_A_pfopnZP06_0(.dout(w_dff_A_ICeAF8Rv5_0),.din(w_dff_A_pfopnZP06_0),.clk(gclk));
	jdff dff_A_ICeAF8Rv5_0(.dout(w_dff_A_ZQbp5s5K0_0),.din(w_dff_A_ICeAF8Rv5_0),.clk(gclk));
	jdff dff_A_ZQbp5s5K0_0(.dout(w_dff_A_YlHX0BwN2_0),.din(w_dff_A_ZQbp5s5K0_0),.clk(gclk));
	jdff dff_A_YlHX0BwN2_0(.dout(w_dff_A_ETy9gqGD1_0),.din(w_dff_A_YlHX0BwN2_0),.clk(gclk));
	jdff dff_A_ETy9gqGD1_0(.dout(w_dff_A_tezJ3UVG9_0),.din(w_dff_A_ETy9gqGD1_0),.clk(gclk));
	jdff dff_A_tezJ3UVG9_0(.dout(w_dff_A_nDsct10I7_0),.din(w_dff_A_tezJ3UVG9_0),.clk(gclk));
	jdff dff_A_nDsct10I7_0(.dout(w_dff_A_pkxGh6lD7_0),.din(w_dff_A_nDsct10I7_0),.clk(gclk));
	jdff dff_A_pkxGh6lD7_0(.dout(w_dff_A_IoOVz7to6_0),.din(w_dff_A_pkxGh6lD7_0),.clk(gclk));
	jdff dff_A_IoOVz7to6_0(.dout(w_dff_A_ffVc2a3L0_0),.din(w_dff_A_IoOVz7to6_0),.clk(gclk));
	jdff dff_A_ffVc2a3L0_0(.dout(w_dff_A_GpB6YlP24_0),.din(w_dff_A_ffVc2a3L0_0),.clk(gclk));
	jdff dff_A_GpB6YlP24_0(.dout(w_dff_A_jT9aZRKk7_0),.din(w_dff_A_GpB6YlP24_0),.clk(gclk));
	jdff dff_A_jT9aZRKk7_0(.dout(w_dff_A_5PaOZazT8_0),.din(w_dff_A_jT9aZRKk7_0),.clk(gclk));
	jdff dff_A_5PaOZazT8_0(.dout(w_dff_A_wseCQdZJ7_0),.din(w_dff_A_5PaOZazT8_0),.clk(gclk));
	jdff dff_A_wseCQdZJ7_0(.dout(w_dff_A_ViE1QtRD1_0),.din(w_dff_A_wseCQdZJ7_0),.clk(gclk));
	jdff dff_A_ViE1QtRD1_0(.dout(w_dff_A_aYFLuSr96_0),.din(w_dff_A_ViE1QtRD1_0),.clk(gclk));
	jdff dff_A_aYFLuSr96_0(.dout(w_dff_A_YoHzFePB3_0),.din(w_dff_A_aYFLuSr96_0),.clk(gclk));
	jdff dff_A_YoHzFePB3_0(.dout(w_dff_A_3YhlgYa31_0),.din(w_dff_A_YoHzFePB3_0),.clk(gclk));
	jdff dff_A_3YhlgYa31_0(.dout(w_dff_A_fQwfeTq67_0),.din(w_dff_A_3YhlgYa31_0),.clk(gclk));
	jdff dff_A_fQwfeTq67_0(.dout(w_dff_A_a55hHrgC9_0),.din(w_dff_A_fQwfeTq67_0),.clk(gclk));
	jdff dff_A_a55hHrgC9_0(.dout(w_dff_A_YmbmVZ1Y5_0),.din(w_dff_A_a55hHrgC9_0),.clk(gclk));
	jdff dff_A_YmbmVZ1Y5_0(.dout(w_dff_A_noCuUxlZ2_0),.din(w_dff_A_YmbmVZ1Y5_0),.clk(gclk));
	jdff dff_A_noCuUxlZ2_0(.dout(w_dff_A_6uwxm9735_0),.din(w_dff_A_noCuUxlZ2_0),.clk(gclk));
	jdff dff_A_6uwxm9735_0(.dout(w_dff_A_M1eDYs1t8_0),.din(w_dff_A_6uwxm9735_0),.clk(gclk));
	jdff dff_A_M1eDYs1t8_0(.dout(w_dff_A_ZLrn5UZR6_0),.din(w_dff_A_M1eDYs1t8_0),.clk(gclk));
	jdff dff_A_ZLrn5UZR6_0(.dout(w_dff_A_jlMQbcnx0_0),.din(w_dff_A_ZLrn5UZR6_0),.clk(gclk));
	jdff dff_A_jlMQbcnx0_0(.dout(w_dff_A_FI99FQIq5_0),.din(w_dff_A_jlMQbcnx0_0),.clk(gclk));
	jdff dff_A_FI99FQIq5_0(.dout(w_dff_A_PY7d6QfG4_0),.din(w_dff_A_FI99FQIq5_0),.clk(gclk));
	jdff dff_A_PY7d6QfG4_0(.dout(w_dff_A_MsWnJVJo1_0),.din(w_dff_A_PY7d6QfG4_0),.clk(gclk));
	jdff dff_A_MsWnJVJo1_0(.dout(w_dff_A_HlLZehqt3_0),.din(w_dff_A_MsWnJVJo1_0),.clk(gclk));
	jdff dff_A_HlLZehqt3_0(.dout(w_dff_A_lpba5pzq6_0),.din(w_dff_A_HlLZehqt3_0),.clk(gclk));
	jdff dff_A_lpba5pzq6_0(.dout(w_dff_A_swV9s9Hu1_0),.din(w_dff_A_lpba5pzq6_0),.clk(gclk));
	jdff dff_A_swV9s9Hu1_0(.dout(w_dff_A_isf6Pk4w8_0),.din(w_dff_A_swV9s9Hu1_0),.clk(gclk));
	jdff dff_A_isf6Pk4w8_0(.dout(w_dff_A_54BANchH9_0),.din(w_dff_A_isf6Pk4w8_0),.clk(gclk));
	jdff dff_A_54BANchH9_0(.dout(w_dff_A_uBzSb6rx4_0),.din(w_dff_A_54BANchH9_0),.clk(gclk));
	jdff dff_A_uBzSb6rx4_0(.dout(w_dff_A_gm0HgLDu1_0),.din(w_dff_A_uBzSb6rx4_0),.clk(gclk));
	jdff dff_A_gm0HgLDu1_0(.dout(w_dff_A_hcXpsd3A4_0),.din(w_dff_A_gm0HgLDu1_0),.clk(gclk));
	jdff dff_A_hcXpsd3A4_0(.dout(w_dff_A_JTFCEfen1_0),.din(w_dff_A_hcXpsd3A4_0),.clk(gclk));
	jdff dff_A_JTFCEfen1_0(.dout(w_dff_A_IjNHmEwA4_0),.din(w_dff_A_JTFCEfen1_0),.clk(gclk));
	jdff dff_A_IjNHmEwA4_0(.dout(w_dff_A_jtOqDm0C1_0),.din(w_dff_A_IjNHmEwA4_0),.clk(gclk));
	jdff dff_A_jtOqDm0C1_0(.dout(w_dff_A_QjAaaF7K9_0),.din(w_dff_A_jtOqDm0C1_0),.clk(gclk));
	jdff dff_A_QjAaaF7K9_0(.dout(w_dff_A_8GVQLnTP6_0),.din(w_dff_A_QjAaaF7K9_0),.clk(gclk));
	jdff dff_A_8GVQLnTP6_0(.dout(w_dff_A_Vjrix28J7_0),.din(w_dff_A_8GVQLnTP6_0),.clk(gclk));
	jdff dff_A_Vjrix28J7_0(.dout(w_dff_A_cuvBx6Za0_0),.din(w_dff_A_Vjrix28J7_0),.clk(gclk));
	jdff dff_A_cuvBx6Za0_0(.dout(w_dff_A_47q9H7HX8_0),.din(w_dff_A_cuvBx6Za0_0),.clk(gclk));
	jdff dff_A_47q9H7HX8_0(.dout(w_dff_A_H6AhyeRT7_0),.din(w_dff_A_47q9H7HX8_0),.clk(gclk));
	jdff dff_A_H6AhyeRT7_0(.dout(w_dff_A_PKpdpdsd9_0),.din(w_dff_A_H6AhyeRT7_0),.clk(gclk));
	jdff dff_A_PKpdpdsd9_0(.dout(w_dff_A_hD7rAjk38_0),.din(w_dff_A_PKpdpdsd9_0),.clk(gclk));
	jdff dff_A_hD7rAjk38_0(.dout(w_dff_A_KthuUe4o7_0),.din(w_dff_A_hD7rAjk38_0),.clk(gclk));
	jdff dff_A_KthuUe4o7_0(.dout(w_dff_A_1IAF9V465_0),.din(w_dff_A_KthuUe4o7_0),.clk(gclk));
	jdff dff_A_1IAF9V465_0(.dout(w_dff_A_rXU0VyyZ5_0),.din(w_dff_A_1IAF9V465_0),.clk(gclk));
	jdff dff_A_rXU0VyyZ5_0(.dout(w_dff_A_WUe1CLaf3_0),.din(w_dff_A_rXU0VyyZ5_0),.clk(gclk));
	jdff dff_A_WUe1CLaf3_0(.dout(w_dff_A_ngZ23UFr9_0),.din(w_dff_A_WUe1CLaf3_0),.clk(gclk));
	jdff dff_A_ngZ23UFr9_0(.dout(w_dff_A_Cc4exuqA1_0),.din(w_dff_A_ngZ23UFr9_0),.clk(gclk));
	jdff dff_A_Cc4exuqA1_0(.dout(w_dff_A_otkrwkU45_0),.din(w_dff_A_Cc4exuqA1_0),.clk(gclk));
	jdff dff_A_otkrwkU45_0(.dout(w_dff_A_dpU3uiMi9_0),.din(w_dff_A_otkrwkU45_0),.clk(gclk));
	jdff dff_A_dpU3uiMi9_0(.dout(w_dff_A_Lz5bU8Ya3_0),.din(w_dff_A_dpU3uiMi9_0),.clk(gclk));
	jdff dff_A_Lz5bU8Ya3_0(.dout(w_dff_A_KhCeDE7y0_0),.din(w_dff_A_Lz5bU8Ya3_0),.clk(gclk));
	jdff dff_A_KhCeDE7y0_0(.dout(w_dff_A_JE5APblT2_0),.din(w_dff_A_KhCeDE7y0_0),.clk(gclk));
	jdff dff_A_JE5APblT2_0(.dout(w_dff_A_3fHyx1Jv4_0),.din(w_dff_A_JE5APblT2_0),.clk(gclk));
	jdff dff_A_3fHyx1Jv4_0(.dout(w_dff_A_9WSXcsoI9_0),.din(w_dff_A_3fHyx1Jv4_0),.clk(gclk));
	jdff dff_A_9WSXcsoI9_0(.dout(w_dff_A_CrqKC3nq1_0),.din(w_dff_A_9WSXcsoI9_0),.clk(gclk));
	jdff dff_A_CrqKC3nq1_0(.dout(w_dff_A_CMHjCS0L6_0),.din(w_dff_A_CrqKC3nq1_0),.clk(gclk));
	jdff dff_A_CMHjCS0L6_0(.dout(w_dff_A_Ice4I31p7_0),.din(w_dff_A_CMHjCS0L6_0),.clk(gclk));
	jdff dff_A_Ice4I31p7_0(.dout(w_dff_A_fpu40RXS1_0),.din(w_dff_A_Ice4I31p7_0),.clk(gclk));
	jdff dff_A_fpu40RXS1_0(.dout(w_dff_A_2GRSyJqq1_0),.din(w_dff_A_fpu40RXS1_0),.clk(gclk));
	jdff dff_A_2GRSyJqq1_0(.dout(G1581gat),.din(w_dff_A_2GRSyJqq1_0),.clk(gclk));
	jdff dff_A_vs4kgBu57_2(.dout(w_dff_A_vt4Y2m9N4_0),.din(w_dff_A_vs4kgBu57_2),.clk(gclk));
	jdff dff_A_vt4Y2m9N4_0(.dout(w_dff_A_tdJLxAiP5_0),.din(w_dff_A_vt4Y2m9N4_0),.clk(gclk));
	jdff dff_A_tdJLxAiP5_0(.dout(w_dff_A_ysaXoF5z7_0),.din(w_dff_A_tdJLxAiP5_0),.clk(gclk));
	jdff dff_A_ysaXoF5z7_0(.dout(w_dff_A_yb9lUVjw4_0),.din(w_dff_A_ysaXoF5z7_0),.clk(gclk));
	jdff dff_A_yb9lUVjw4_0(.dout(w_dff_A_DZ3QFxdG1_0),.din(w_dff_A_yb9lUVjw4_0),.clk(gclk));
	jdff dff_A_DZ3QFxdG1_0(.dout(w_dff_A_IKsb1xaL8_0),.din(w_dff_A_DZ3QFxdG1_0),.clk(gclk));
	jdff dff_A_IKsb1xaL8_0(.dout(w_dff_A_X4Tjeb5v1_0),.din(w_dff_A_IKsb1xaL8_0),.clk(gclk));
	jdff dff_A_X4Tjeb5v1_0(.dout(w_dff_A_LdUcYung7_0),.din(w_dff_A_X4Tjeb5v1_0),.clk(gclk));
	jdff dff_A_LdUcYung7_0(.dout(w_dff_A_UcmHguER2_0),.din(w_dff_A_LdUcYung7_0),.clk(gclk));
	jdff dff_A_UcmHguER2_0(.dout(w_dff_A_72XggFCi2_0),.din(w_dff_A_UcmHguER2_0),.clk(gclk));
	jdff dff_A_72XggFCi2_0(.dout(w_dff_A_BDzujJga3_0),.din(w_dff_A_72XggFCi2_0),.clk(gclk));
	jdff dff_A_BDzujJga3_0(.dout(w_dff_A_Ws06adqW6_0),.din(w_dff_A_BDzujJga3_0),.clk(gclk));
	jdff dff_A_Ws06adqW6_0(.dout(w_dff_A_8aQeNKaS1_0),.din(w_dff_A_Ws06adqW6_0),.clk(gclk));
	jdff dff_A_8aQeNKaS1_0(.dout(w_dff_A_eej1nWK37_0),.din(w_dff_A_8aQeNKaS1_0),.clk(gclk));
	jdff dff_A_eej1nWK37_0(.dout(w_dff_A_3zS0AzMv2_0),.din(w_dff_A_eej1nWK37_0),.clk(gclk));
	jdff dff_A_3zS0AzMv2_0(.dout(w_dff_A_NpqL8I028_0),.din(w_dff_A_3zS0AzMv2_0),.clk(gclk));
	jdff dff_A_NpqL8I028_0(.dout(w_dff_A_wavaedhY7_0),.din(w_dff_A_NpqL8I028_0),.clk(gclk));
	jdff dff_A_wavaedhY7_0(.dout(w_dff_A_Rqw8Vh8i6_0),.din(w_dff_A_wavaedhY7_0),.clk(gclk));
	jdff dff_A_Rqw8Vh8i6_0(.dout(w_dff_A_WHQiO8fC0_0),.din(w_dff_A_Rqw8Vh8i6_0),.clk(gclk));
	jdff dff_A_WHQiO8fC0_0(.dout(w_dff_A_7uDrAlfu4_0),.din(w_dff_A_WHQiO8fC0_0),.clk(gclk));
	jdff dff_A_7uDrAlfu4_0(.dout(w_dff_A_qmfrpfF93_0),.din(w_dff_A_7uDrAlfu4_0),.clk(gclk));
	jdff dff_A_qmfrpfF93_0(.dout(w_dff_A_KH2RYoTc0_0),.din(w_dff_A_qmfrpfF93_0),.clk(gclk));
	jdff dff_A_KH2RYoTc0_0(.dout(w_dff_A_TyYzH7Uv2_0),.din(w_dff_A_KH2RYoTc0_0),.clk(gclk));
	jdff dff_A_TyYzH7Uv2_0(.dout(w_dff_A_KfMod0ct7_0),.din(w_dff_A_TyYzH7Uv2_0),.clk(gclk));
	jdff dff_A_KfMod0ct7_0(.dout(w_dff_A_BVjaDU2z8_0),.din(w_dff_A_KfMod0ct7_0),.clk(gclk));
	jdff dff_A_BVjaDU2z8_0(.dout(w_dff_A_umMVj3Sw2_0),.din(w_dff_A_BVjaDU2z8_0),.clk(gclk));
	jdff dff_A_umMVj3Sw2_0(.dout(w_dff_A_8XdyYXqr5_0),.din(w_dff_A_umMVj3Sw2_0),.clk(gclk));
	jdff dff_A_8XdyYXqr5_0(.dout(w_dff_A_FdIxDJKN6_0),.din(w_dff_A_8XdyYXqr5_0),.clk(gclk));
	jdff dff_A_FdIxDJKN6_0(.dout(w_dff_A_uAXBNBkM6_0),.din(w_dff_A_FdIxDJKN6_0),.clk(gclk));
	jdff dff_A_uAXBNBkM6_0(.dout(w_dff_A_XC0zWnLJ8_0),.din(w_dff_A_uAXBNBkM6_0),.clk(gclk));
	jdff dff_A_XC0zWnLJ8_0(.dout(w_dff_A_u5SMg9nV2_0),.din(w_dff_A_XC0zWnLJ8_0),.clk(gclk));
	jdff dff_A_u5SMg9nV2_0(.dout(w_dff_A_jKEUbQ1I1_0),.din(w_dff_A_u5SMg9nV2_0),.clk(gclk));
	jdff dff_A_jKEUbQ1I1_0(.dout(w_dff_A_CDJ35Hec5_0),.din(w_dff_A_jKEUbQ1I1_0),.clk(gclk));
	jdff dff_A_CDJ35Hec5_0(.dout(w_dff_A_lJ68NMyc3_0),.din(w_dff_A_CDJ35Hec5_0),.clk(gclk));
	jdff dff_A_lJ68NMyc3_0(.dout(w_dff_A_QVMWhmzb5_0),.din(w_dff_A_lJ68NMyc3_0),.clk(gclk));
	jdff dff_A_QVMWhmzb5_0(.dout(w_dff_A_oFYx4XUi9_0),.din(w_dff_A_QVMWhmzb5_0),.clk(gclk));
	jdff dff_A_oFYx4XUi9_0(.dout(w_dff_A_VzovCNYm7_0),.din(w_dff_A_oFYx4XUi9_0),.clk(gclk));
	jdff dff_A_VzovCNYm7_0(.dout(w_dff_A_kUCaB2we9_0),.din(w_dff_A_VzovCNYm7_0),.clk(gclk));
	jdff dff_A_kUCaB2we9_0(.dout(w_dff_A_K0Ilz7YP0_0),.din(w_dff_A_kUCaB2we9_0),.clk(gclk));
	jdff dff_A_K0Ilz7YP0_0(.dout(w_dff_A_AlwT8s9K8_0),.din(w_dff_A_K0Ilz7YP0_0),.clk(gclk));
	jdff dff_A_AlwT8s9K8_0(.dout(w_dff_A_8bn5XCZH8_0),.din(w_dff_A_AlwT8s9K8_0),.clk(gclk));
	jdff dff_A_8bn5XCZH8_0(.dout(w_dff_A_SJntTOgD2_0),.din(w_dff_A_8bn5XCZH8_0),.clk(gclk));
	jdff dff_A_SJntTOgD2_0(.dout(w_dff_A_N7hK5Ywo5_0),.din(w_dff_A_SJntTOgD2_0),.clk(gclk));
	jdff dff_A_N7hK5Ywo5_0(.dout(w_dff_A_V1IkvfIo0_0),.din(w_dff_A_N7hK5Ywo5_0),.clk(gclk));
	jdff dff_A_V1IkvfIo0_0(.dout(w_dff_A_C8vVumad3_0),.din(w_dff_A_V1IkvfIo0_0),.clk(gclk));
	jdff dff_A_C8vVumad3_0(.dout(w_dff_A_aB2V1atm8_0),.din(w_dff_A_C8vVumad3_0),.clk(gclk));
	jdff dff_A_aB2V1atm8_0(.dout(w_dff_A_pIu8zC9C4_0),.din(w_dff_A_aB2V1atm8_0),.clk(gclk));
	jdff dff_A_pIu8zC9C4_0(.dout(w_dff_A_1ItMPxZD5_0),.din(w_dff_A_pIu8zC9C4_0),.clk(gclk));
	jdff dff_A_1ItMPxZD5_0(.dout(w_dff_A_nFjwKY4e4_0),.din(w_dff_A_1ItMPxZD5_0),.clk(gclk));
	jdff dff_A_nFjwKY4e4_0(.dout(w_dff_A_7ylqROtw0_0),.din(w_dff_A_nFjwKY4e4_0),.clk(gclk));
	jdff dff_A_7ylqROtw0_0(.dout(w_dff_A_vReCnBqg2_0),.din(w_dff_A_7ylqROtw0_0),.clk(gclk));
	jdff dff_A_vReCnBqg2_0(.dout(w_dff_A_wRKgzkYP8_0),.din(w_dff_A_vReCnBqg2_0),.clk(gclk));
	jdff dff_A_wRKgzkYP8_0(.dout(w_dff_A_ykqs3oh58_0),.din(w_dff_A_wRKgzkYP8_0),.clk(gclk));
	jdff dff_A_ykqs3oh58_0(.dout(w_dff_A_UBa2lvoL8_0),.din(w_dff_A_ykqs3oh58_0),.clk(gclk));
	jdff dff_A_UBa2lvoL8_0(.dout(w_dff_A_f6GTBfjN3_0),.din(w_dff_A_UBa2lvoL8_0),.clk(gclk));
	jdff dff_A_f6GTBfjN3_0(.dout(w_dff_A_WpFZOaXU6_0),.din(w_dff_A_f6GTBfjN3_0),.clk(gclk));
	jdff dff_A_WpFZOaXU6_0(.dout(w_dff_A_R1PDDnD57_0),.din(w_dff_A_WpFZOaXU6_0),.clk(gclk));
	jdff dff_A_R1PDDnD57_0(.dout(w_dff_A_yuUlPWbi8_0),.din(w_dff_A_R1PDDnD57_0),.clk(gclk));
	jdff dff_A_yuUlPWbi8_0(.dout(w_dff_A_oPpAL3Eb8_0),.din(w_dff_A_yuUlPWbi8_0),.clk(gclk));
	jdff dff_A_oPpAL3Eb8_0(.dout(w_dff_A_YOEyE2Ft4_0),.din(w_dff_A_oPpAL3Eb8_0),.clk(gclk));
	jdff dff_A_YOEyE2Ft4_0(.dout(w_dff_A_ymDkE7QA9_0),.din(w_dff_A_YOEyE2Ft4_0),.clk(gclk));
	jdff dff_A_ymDkE7QA9_0(.dout(w_dff_A_PcpGoIOS7_0),.din(w_dff_A_ymDkE7QA9_0),.clk(gclk));
	jdff dff_A_PcpGoIOS7_0(.dout(w_dff_A_GVHM0wzS0_0),.din(w_dff_A_PcpGoIOS7_0),.clk(gclk));
	jdff dff_A_GVHM0wzS0_0(.dout(w_dff_A_DPLpEJdk3_0),.din(w_dff_A_GVHM0wzS0_0),.clk(gclk));
	jdff dff_A_DPLpEJdk3_0(.dout(w_dff_A_h4nhCUpe5_0),.din(w_dff_A_DPLpEJdk3_0),.clk(gclk));
	jdff dff_A_h4nhCUpe5_0(.dout(w_dff_A_jFUWWvbN5_0),.din(w_dff_A_h4nhCUpe5_0),.clk(gclk));
	jdff dff_A_jFUWWvbN5_0(.dout(w_dff_A_X2qNxCpV7_0),.din(w_dff_A_jFUWWvbN5_0),.clk(gclk));
	jdff dff_A_X2qNxCpV7_0(.dout(w_dff_A_ot49Qtx87_0),.din(w_dff_A_X2qNxCpV7_0),.clk(gclk));
	jdff dff_A_ot49Qtx87_0(.dout(G1901gat),.din(w_dff_A_ot49Qtx87_0),.clk(gclk));
	jdff dff_A_D1J7lZ8S1_2(.dout(w_dff_A_5VdlFGQX8_0),.din(w_dff_A_D1J7lZ8S1_2),.clk(gclk));
	jdff dff_A_5VdlFGQX8_0(.dout(w_dff_A_11uqXQUt4_0),.din(w_dff_A_5VdlFGQX8_0),.clk(gclk));
	jdff dff_A_11uqXQUt4_0(.dout(w_dff_A_z0hbwh0k0_0),.din(w_dff_A_11uqXQUt4_0),.clk(gclk));
	jdff dff_A_z0hbwh0k0_0(.dout(w_dff_A_5Ea3pvvn7_0),.din(w_dff_A_z0hbwh0k0_0),.clk(gclk));
	jdff dff_A_5Ea3pvvn7_0(.dout(w_dff_A_3MSpyuVM9_0),.din(w_dff_A_5Ea3pvvn7_0),.clk(gclk));
	jdff dff_A_3MSpyuVM9_0(.dout(w_dff_A_NPlD3U850_0),.din(w_dff_A_3MSpyuVM9_0),.clk(gclk));
	jdff dff_A_NPlD3U850_0(.dout(w_dff_A_aY6hHetZ2_0),.din(w_dff_A_NPlD3U850_0),.clk(gclk));
	jdff dff_A_aY6hHetZ2_0(.dout(w_dff_A_AYeoMJMa5_0),.din(w_dff_A_aY6hHetZ2_0),.clk(gclk));
	jdff dff_A_AYeoMJMa5_0(.dout(w_dff_A_DOvmNg326_0),.din(w_dff_A_AYeoMJMa5_0),.clk(gclk));
	jdff dff_A_DOvmNg326_0(.dout(w_dff_A_KIgKS7ex0_0),.din(w_dff_A_DOvmNg326_0),.clk(gclk));
	jdff dff_A_KIgKS7ex0_0(.dout(w_dff_A_dPOfIh3R4_0),.din(w_dff_A_KIgKS7ex0_0),.clk(gclk));
	jdff dff_A_dPOfIh3R4_0(.dout(w_dff_A_xxd3ghpm2_0),.din(w_dff_A_dPOfIh3R4_0),.clk(gclk));
	jdff dff_A_xxd3ghpm2_0(.dout(w_dff_A_4fX1ZjQL2_0),.din(w_dff_A_xxd3ghpm2_0),.clk(gclk));
	jdff dff_A_4fX1ZjQL2_0(.dout(w_dff_A_9pAvsRqz4_0),.din(w_dff_A_4fX1ZjQL2_0),.clk(gclk));
	jdff dff_A_9pAvsRqz4_0(.dout(w_dff_A_x6XmJUgp0_0),.din(w_dff_A_9pAvsRqz4_0),.clk(gclk));
	jdff dff_A_x6XmJUgp0_0(.dout(w_dff_A_gu6RG1KW0_0),.din(w_dff_A_x6XmJUgp0_0),.clk(gclk));
	jdff dff_A_gu6RG1KW0_0(.dout(w_dff_A_XcB9VRBe6_0),.din(w_dff_A_gu6RG1KW0_0),.clk(gclk));
	jdff dff_A_XcB9VRBe6_0(.dout(w_dff_A_SiOvmyOY5_0),.din(w_dff_A_XcB9VRBe6_0),.clk(gclk));
	jdff dff_A_SiOvmyOY5_0(.dout(w_dff_A_N8pYPSn50_0),.din(w_dff_A_SiOvmyOY5_0),.clk(gclk));
	jdff dff_A_N8pYPSn50_0(.dout(w_dff_A_yjZxB4u51_0),.din(w_dff_A_N8pYPSn50_0),.clk(gclk));
	jdff dff_A_yjZxB4u51_0(.dout(w_dff_A_7kkk1XYh7_0),.din(w_dff_A_yjZxB4u51_0),.clk(gclk));
	jdff dff_A_7kkk1XYh7_0(.dout(w_dff_A_IHH1p1JI5_0),.din(w_dff_A_7kkk1XYh7_0),.clk(gclk));
	jdff dff_A_IHH1p1JI5_0(.dout(w_dff_A_LziHCwwI2_0),.din(w_dff_A_IHH1p1JI5_0),.clk(gclk));
	jdff dff_A_LziHCwwI2_0(.dout(w_dff_A_VQMpyaCL4_0),.din(w_dff_A_LziHCwwI2_0),.clk(gclk));
	jdff dff_A_VQMpyaCL4_0(.dout(w_dff_A_qZ43ZVAg2_0),.din(w_dff_A_VQMpyaCL4_0),.clk(gclk));
	jdff dff_A_qZ43ZVAg2_0(.dout(w_dff_A_ia4uFhAI3_0),.din(w_dff_A_qZ43ZVAg2_0),.clk(gclk));
	jdff dff_A_ia4uFhAI3_0(.dout(w_dff_A_JBgWHlnm6_0),.din(w_dff_A_ia4uFhAI3_0),.clk(gclk));
	jdff dff_A_JBgWHlnm6_0(.dout(w_dff_A_jrHgQmEH5_0),.din(w_dff_A_JBgWHlnm6_0),.clk(gclk));
	jdff dff_A_jrHgQmEH5_0(.dout(w_dff_A_Ol8FOpdB8_0),.din(w_dff_A_jrHgQmEH5_0),.clk(gclk));
	jdff dff_A_Ol8FOpdB8_0(.dout(w_dff_A_Ipo92fHW3_0),.din(w_dff_A_Ol8FOpdB8_0),.clk(gclk));
	jdff dff_A_Ipo92fHW3_0(.dout(w_dff_A_XnBgPrZf6_0),.din(w_dff_A_Ipo92fHW3_0),.clk(gclk));
	jdff dff_A_XnBgPrZf6_0(.dout(w_dff_A_qGfGdB2L8_0),.din(w_dff_A_XnBgPrZf6_0),.clk(gclk));
	jdff dff_A_qGfGdB2L8_0(.dout(w_dff_A_MwnirlbD0_0),.din(w_dff_A_qGfGdB2L8_0),.clk(gclk));
	jdff dff_A_MwnirlbD0_0(.dout(w_dff_A_ZFFw6czc6_0),.din(w_dff_A_MwnirlbD0_0),.clk(gclk));
	jdff dff_A_ZFFw6czc6_0(.dout(w_dff_A_m4Ze4Ssf3_0),.din(w_dff_A_ZFFw6czc6_0),.clk(gclk));
	jdff dff_A_m4Ze4Ssf3_0(.dout(w_dff_A_ATdCIE9I0_0),.din(w_dff_A_m4Ze4Ssf3_0),.clk(gclk));
	jdff dff_A_ATdCIE9I0_0(.dout(w_dff_A_mTZKJUhg0_0),.din(w_dff_A_ATdCIE9I0_0),.clk(gclk));
	jdff dff_A_mTZKJUhg0_0(.dout(w_dff_A_1ylxeht97_0),.din(w_dff_A_mTZKJUhg0_0),.clk(gclk));
	jdff dff_A_1ylxeht97_0(.dout(w_dff_A_11aitGHD7_0),.din(w_dff_A_1ylxeht97_0),.clk(gclk));
	jdff dff_A_11aitGHD7_0(.dout(w_dff_A_NhXWoq7n7_0),.din(w_dff_A_11aitGHD7_0),.clk(gclk));
	jdff dff_A_NhXWoq7n7_0(.dout(w_dff_A_jGAapAjR2_0),.din(w_dff_A_NhXWoq7n7_0),.clk(gclk));
	jdff dff_A_jGAapAjR2_0(.dout(w_dff_A_R34ICqlN3_0),.din(w_dff_A_jGAapAjR2_0),.clk(gclk));
	jdff dff_A_R34ICqlN3_0(.dout(w_dff_A_56vmJzb38_0),.din(w_dff_A_R34ICqlN3_0),.clk(gclk));
	jdff dff_A_56vmJzb38_0(.dout(w_dff_A_floHRrHw9_0),.din(w_dff_A_56vmJzb38_0),.clk(gclk));
	jdff dff_A_floHRrHw9_0(.dout(w_dff_A_a6CXb8Ng1_0),.din(w_dff_A_floHRrHw9_0),.clk(gclk));
	jdff dff_A_a6CXb8Ng1_0(.dout(w_dff_A_UYKcMncX9_0),.din(w_dff_A_a6CXb8Ng1_0),.clk(gclk));
	jdff dff_A_UYKcMncX9_0(.dout(w_dff_A_WRmRh7vK6_0),.din(w_dff_A_UYKcMncX9_0),.clk(gclk));
	jdff dff_A_WRmRh7vK6_0(.dout(w_dff_A_ATRCgMXG2_0),.din(w_dff_A_WRmRh7vK6_0),.clk(gclk));
	jdff dff_A_ATRCgMXG2_0(.dout(w_dff_A_g6OSqU0P0_0),.din(w_dff_A_ATRCgMXG2_0),.clk(gclk));
	jdff dff_A_g6OSqU0P0_0(.dout(w_dff_A_4mTXAxGe0_0),.din(w_dff_A_g6OSqU0P0_0),.clk(gclk));
	jdff dff_A_4mTXAxGe0_0(.dout(w_dff_A_BvAqLBDM8_0),.din(w_dff_A_4mTXAxGe0_0),.clk(gclk));
	jdff dff_A_BvAqLBDM8_0(.dout(w_dff_A_vd4bv5001_0),.din(w_dff_A_BvAqLBDM8_0),.clk(gclk));
	jdff dff_A_vd4bv5001_0(.dout(w_dff_A_RDzJZCix4_0),.din(w_dff_A_vd4bv5001_0),.clk(gclk));
	jdff dff_A_RDzJZCix4_0(.dout(w_dff_A_sZKMNCFf6_0),.din(w_dff_A_RDzJZCix4_0),.clk(gclk));
	jdff dff_A_sZKMNCFf6_0(.dout(w_dff_A_rgER3r5x9_0),.din(w_dff_A_sZKMNCFf6_0),.clk(gclk));
	jdff dff_A_rgER3r5x9_0(.dout(w_dff_A_CQLc17Wd1_0),.din(w_dff_A_rgER3r5x9_0),.clk(gclk));
	jdff dff_A_CQLc17Wd1_0(.dout(w_dff_A_agLNOFAh4_0),.din(w_dff_A_CQLc17Wd1_0),.clk(gclk));
	jdff dff_A_agLNOFAh4_0(.dout(w_dff_A_auIuwebJ2_0),.din(w_dff_A_agLNOFAh4_0),.clk(gclk));
	jdff dff_A_auIuwebJ2_0(.dout(w_dff_A_NjVTGFQ62_0),.din(w_dff_A_auIuwebJ2_0),.clk(gclk));
	jdff dff_A_NjVTGFQ62_0(.dout(w_dff_A_Vzs7Oa837_0),.din(w_dff_A_NjVTGFQ62_0),.clk(gclk));
	jdff dff_A_Vzs7Oa837_0(.dout(w_dff_A_7D3sDAAy3_0),.din(w_dff_A_Vzs7Oa837_0),.clk(gclk));
	jdff dff_A_7D3sDAAy3_0(.dout(w_dff_A_9gn8rMLL5_0),.din(w_dff_A_7D3sDAAy3_0),.clk(gclk));
	jdff dff_A_9gn8rMLL5_0(.dout(w_dff_A_nWwozueN8_0),.din(w_dff_A_9gn8rMLL5_0),.clk(gclk));
	jdff dff_A_nWwozueN8_0(.dout(w_dff_A_TmBQdEiT0_0),.din(w_dff_A_nWwozueN8_0),.clk(gclk));
	jdff dff_A_TmBQdEiT0_0(.dout(w_dff_A_C7GbskCZ8_0),.din(w_dff_A_TmBQdEiT0_0),.clk(gclk));
	jdff dff_A_C7GbskCZ8_0(.dout(G2223gat),.din(w_dff_A_C7GbskCZ8_0),.clk(gclk));
	jdff dff_A_PldpzvGS2_2(.dout(w_dff_A_QaN4hjlH1_0),.din(w_dff_A_PldpzvGS2_2),.clk(gclk));
	jdff dff_A_QaN4hjlH1_0(.dout(w_dff_A_ux1XDO1D5_0),.din(w_dff_A_QaN4hjlH1_0),.clk(gclk));
	jdff dff_A_ux1XDO1D5_0(.dout(w_dff_A_VVd3iCVb6_0),.din(w_dff_A_ux1XDO1D5_0),.clk(gclk));
	jdff dff_A_VVd3iCVb6_0(.dout(w_dff_A_BiukFx9j7_0),.din(w_dff_A_VVd3iCVb6_0),.clk(gclk));
	jdff dff_A_BiukFx9j7_0(.dout(w_dff_A_PDAsfrc99_0),.din(w_dff_A_BiukFx9j7_0),.clk(gclk));
	jdff dff_A_PDAsfrc99_0(.dout(w_dff_A_GSIKqZTW5_0),.din(w_dff_A_PDAsfrc99_0),.clk(gclk));
	jdff dff_A_GSIKqZTW5_0(.dout(w_dff_A_dIJmV9rb3_0),.din(w_dff_A_GSIKqZTW5_0),.clk(gclk));
	jdff dff_A_dIJmV9rb3_0(.dout(w_dff_A_cwgYcYzE4_0),.din(w_dff_A_dIJmV9rb3_0),.clk(gclk));
	jdff dff_A_cwgYcYzE4_0(.dout(w_dff_A_hOtfK5E33_0),.din(w_dff_A_cwgYcYzE4_0),.clk(gclk));
	jdff dff_A_hOtfK5E33_0(.dout(w_dff_A_1pHepJP47_0),.din(w_dff_A_hOtfK5E33_0),.clk(gclk));
	jdff dff_A_1pHepJP47_0(.dout(w_dff_A_BpE9rstO0_0),.din(w_dff_A_1pHepJP47_0),.clk(gclk));
	jdff dff_A_BpE9rstO0_0(.dout(w_dff_A_QXxbKmvC7_0),.din(w_dff_A_BpE9rstO0_0),.clk(gclk));
	jdff dff_A_QXxbKmvC7_0(.dout(w_dff_A_U2ceAQvx6_0),.din(w_dff_A_QXxbKmvC7_0),.clk(gclk));
	jdff dff_A_U2ceAQvx6_0(.dout(w_dff_A_TK3rNgCK0_0),.din(w_dff_A_U2ceAQvx6_0),.clk(gclk));
	jdff dff_A_TK3rNgCK0_0(.dout(w_dff_A_EMGVVePw8_0),.din(w_dff_A_TK3rNgCK0_0),.clk(gclk));
	jdff dff_A_EMGVVePw8_0(.dout(w_dff_A_WTfNUG740_0),.din(w_dff_A_EMGVVePw8_0),.clk(gclk));
	jdff dff_A_WTfNUG740_0(.dout(w_dff_A_HHJvtuQG2_0),.din(w_dff_A_WTfNUG740_0),.clk(gclk));
	jdff dff_A_HHJvtuQG2_0(.dout(w_dff_A_1AZotT3V1_0),.din(w_dff_A_HHJvtuQG2_0),.clk(gclk));
	jdff dff_A_1AZotT3V1_0(.dout(w_dff_A_uZp04kMa4_0),.din(w_dff_A_1AZotT3V1_0),.clk(gclk));
	jdff dff_A_uZp04kMa4_0(.dout(w_dff_A_2Qd176o97_0),.din(w_dff_A_uZp04kMa4_0),.clk(gclk));
	jdff dff_A_2Qd176o97_0(.dout(w_dff_A_Pg0ws8P03_0),.din(w_dff_A_2Qd176o97_0),.clk(gclk));
	jdff dff_A_Pg0ws8P03_0(.dout(w_dff_A_98A75F9Z1_0),.din(w_dff_A_Pg0ws8P03_0),.clk(gclk));
	jdff dff_A_98A75F9Z1_0(.dout(w_dff_A_zKruO8ht1_0),.din(w_dff_A_98A75F9Z1_0),.clk(gclk));
	jdff dff_A_zKruO8ht1_0(.dout(w_dff_A_vvt1aiZm5_0),.din(w_dff_A_zKruO8ht1_0),.clk(gclk));
	jdff dff_A_vvt1aiZm5_0(.dout(w_dff_A_I1tgTuJy7_0),.din(w_dff_A_vvt1aiZm5_0),.clk(gclk));
	jdff dff_A_I1tgTuJy7_0(.dout(w_dff_A_y0RZYSPV7_0),.din(w_dff_A_I1tgTuJy7_0),.clk(gclk));
	jdff dff_A_y0RZYSPV7_0(.dout(w_dff_A_jxl0YOe47_0),.din(w_dff_A_y0RZYSPV7_0),.clk(gclk));
	jdff dff_A_jxl0YOe47_0(.dout(w_dff_A_4k0oDl9z6_0),.din(w_dff_A_jxl0YOe47_0),.clk(gclk));
	jdff dff_A_4k0oDl9z6_0(.dout(w_dff_A_tNSDqPDw4_0),.din(w_dff_A_4k0oDl9z6_0),.clk(gclk));
	jdff dff_A_tNSDqPDw4_0(.dout(w_dff_A_D1MbQm2I7_0),.din(w_dff_A_tNSDqPDw4_0),.clk(gclk));
	jdff dff_A_D1MbQm2I7_0(.dout(w_dff_A_PIlN1MBS3_0),.din(w_dff_A_D1MbQm2I7_0),.clk(gclk));
	jdff dff_A_PIlN1MBS3_0(.dout(w_dff_A_8CeeJWxV9_0),.din(w_dff_A_PIlN1MBS3_0),.clk(gclk));
	jdff dff_A_8CeeJWxV9_0(.dout(w_dff_A_9hxGB0Dr6_0),.din(w_dff_A_8CeeJWxV9_0),.clk(gclk));
	jdff dff_A_9hxGB0Dr6_0(.dout(w_dff_A_7j24TzSO2_0),.din(w_dff_A_9hxGB0Dr6_0),.clk(gclk));
	jdff dff_A_7j24TzSO2_0(.dout(w_dff_A_ZrqnpYrO6_0),.din(w_dff_A_7j24TzSO2_0),.clk(gclk));
	jdff dff_A_ZrqnpYrO6_0(.dout(w_dff_A_NUuKzZNk9_0),.din(w_dff_A_ZrqnpYrO6_0),.clk(gclk));
	jdff dff_A_NUuKzZNk9_0(.dout(w_dff_A_1osgNuPS4_0),.din(w_dff_A_NUuKzZNk9_0),.clk(gclk));
	jdff dff_A_1osgNuPS4_0(.dout(w_dff_A_XtUBurmn0_0),.din(w_dff_A_1osgNuPS4_0),.clk(gclk));
	jdff dff_A_XtUBurmn0_0(.dout(w_dff_A_nCOAkcvA3_0),.din(w_dff_A_XtUBurmn0_0),.clk(gclk));
	jdff dff_A_nCOAkcvA3_0(.dout(w_dff_A_OfAwnrYR2_0),.din(w_dff_A_nCOAkcvA3_0),.clk(gclk));
	jdff dff_A_OfAwnrYR2_0(.dout(w_dff_A_OfdBXbLF8_0),.din(w_dff_A_OfAwnrYR2_0),.clk(gclk));
	jdff dff_A_OfdBXbLF8_0(.dout(w_dff_A_eH0MGLK35_0),.din(w_dff_A_OfdBXbLF8_0),.clk(gclk));
	jdff dff_A_eH0MGLK35_0(.dout(w_dff_A_whbKx2wh6_0),.din(w_dff_A_eH0MGLK35_0),.clk(gclk));
	jdff dff_A_whbKx2wh6_0(.dout(w_dff_A_5RoUYWqt7_0),.din(w_dff_A_whbKx2wh6_0),.clk(gclk));
	jdff dff_A_5RoUYWqt7_0(.dout(w_dff_A_MfljODPt6_0),.din(w_dff_A_5RoUYWqt7_0),.clk(gclk));
	jdff dff_A_MfljODPt6_0(.dout(w_dff_A_Mv7MkqSf1_0),.din(w_dff_A_MfljODPt6_0),.clk(gclk));
	jdff dff_A_Mv7MkqSf1_0(.dout(w_dff_A_spk3HlPx2_0),.din(w_dff_A_Mv7MkqSf1_0),.clk(gclk));
	jdff dff_A_spk3HlPx2_0(.dout(w_dff_A_59u8j0E63_0),.din(w_dff_A_spk3HlPx2_0),.clk(gclk));
	jdff dff_A_59u8j0E63_0(.dout(w_dff_A_FsmbLvpH8_0),.din(w_dff_A_59u8j0E63_0),.clk(gclk));
	jdff dff_A_FsmbLvpH8_0(.dout(w_dff_A_T2n6wKPW0_0),.din(w_dff_A_FsmbLvpH8_0),.clk(gclk));
	jdff dff_A_T2n6wKPW0_0(.dout(w_dff_A_Jh2YMt7n6_0),.din(w_dff_A_T2n6wKPW0_0),.clk(gclk));
	jdff dff_A_Jh2YMt7n6_0(.dout(w_dff_A_w9IxogiP3_0),.din(w_dff_A_Jh2YMt7n6_0),.clk(gclk));
	jdff dff_A_w9IxogiP3_0(.dout(w_dff_A_x22pA9Dg2_0),.din(w_dff_A_w9IxogiP3_0),.clk(gclk));
	jdff dff_A_x22pA9Dg2_0(.dout(w_dff_A_Nn3xoHwg4_0),.din(w_dff_A_x22pA9Dg2_0),.clk(gclk));
	jdff dff_A_Nn3xoHwg4_0(.dout(w_dff_A_iOplehm90_0),.din(w_dff_A_Nn3xoHwg4_0),.clk(gclk));
	jdff dff_A_iOplehm90_0(.dout(w_dff_A_SzGz9iH07_0),.din(w_dff_A_iOplehm90_0),.clk(gclk));
	jdff dff_A_SzGz9iH07_0(.dout(w_dff_A_wjnyXDYZ8_0),.din(w_dff_A_SzGz9iH07_0),.clk(gclk));
	jdff dff_A_wjnyXDYZ8_0(.dout(w_dff_A_lgjC48jg0_0),.din(w_dff_A_wjnyXDYZ8_0),.clk(gclk));
	jdff dff_A_lgjC48jg0_0(.dout(w_dff_A_ivBOeMVc6_0),.din(w_dff_A_lgjC48jg0_0),.clk(gclk));
	jdff dff_A_ivBOeMVc6_0(.dout(w_dff_A_Su5wLHVe0_0),.din(w_dff_A_ivBOeMVc6_0),.clk(gclk));
	jdff dff_A_Su5wLHVe0_0(.dout(w_dff_A_B3yINSX60_0),.din(w_dff_A_Su5wLHVe0_0),.clk(gclk));
	jdff dff_A_B3yINSX60_0(.dout(w_dff_A_W3AJC9D04_0),.din(w_dff_A_B3yINSX60_0),.clk(gclk));
	jdff dff_A_W3AJC9D04_0(.dout(G2548gat),.din(w_dff_A_W3AJC9D04_0),.clk(gclk));
	jdff dff_A_YL90IabU6_2(.dout(w_dff_A_hSbn9xYI2_0),.din(w_dff_A_YL90IabU6_2),.clk(gclk));
	jdff dff_A_hSbn9xYI2_0(.dout(w_dff_A_CVqIS5yc9_0),.din(w_dff_A_hSbn9xYI2_0),.clk(gclk));
	jdff dff_A_CVqIS5yc9_0(.dout(w_dff_A_8s2g5Me99_0),.din(w_dff_A_CVqIS5yc9_0),.clk(gclk));
	jdff dff_A_8s2g5Me99_0(.dout(w_dff_A_TC7gfXnH7_0),.din(w_dff_A_8s2g5Me99_0),.clk(gclk));
	jdff dff_A_TC7gfXnH7_0(.dout(w_dff_A_JjI8d8YY3_0),.din(w_dff_A_TC7gfXnH7_0),.clk(gclk));
	jdff dff_A_JjI8d8YY3_0(.dout(w_dff_A_etQJDmiQ9_0),.din(w_dff_A_JjI8d8YY3_0),.clk(gclk));
	jdff dff_A_etQJDmiQ9_0(.dout(w_dff_A_NbObjnJx2_0),.din(w_dff_A_etQJDmiQ9_0),.clk(gclk));
	jdff dff_A_NbObjnJx2_0(.dout(w_dff_A_Up1xVSlF6_0),.din(w_dff_A_NbObjnJx2_0),.clk(gclk));
	jdff dff_A_Up1xVSlF6_0(.dout(w_dff_A_dbZUezcG7_0),.din(w_dff_A_Up1xVSlF6_0),.clk(gclk));
	jdff dff_A_dbZUezcG7_0(.dout(w_dff_A_EdVkP9cB3_0),.din(w_dff_A_dbZUezcG7_0),.clk(gclk));
	jdff dff_A_EdVkP9cB3_0(.dout(w_dff_A_uDtCIdfn4_0),.din(w_dff_A_EdVkP9cB3_0),.clk(gclk));
	jdff dff_A_uDtCIdfn4_0(.dout(w_dff_A_cjIiqBUC8_0),.din(w_dff_A_uDtCIdfn4_0),.clk(gclk));
	jdff dff_A_cjIiqBUC8_0(.dout(w_dff_A_rjrB2rRP7_0),.din(w_dff_A_cjIiqBUC8_0),.clk(gclk));
	jdff dff_A_rjrB2rRP7_0(.dout(w_dff_A_pPMhbB8H3_0),.din(w_dff_A_rjrB2rRP7_0),.clk(gclk));
	jdff dff_A_pPMhbB8H3_0(.dout(w_dff_A_yVEumW7h3_0),.din(w_dff_A_pPMhbB8H3_0),.clk(gclk));
	jdff dff_A_yVEumW7h3_0(.dout(w_dff_A_LYwKI1nT2_0),.din(w_dff_A_yVEumW7h3_0),.clk(gclk));
	jdff dff_A_LYwKI1nT2_0(.dout(w_dff_A_DFMR8NpH6_0),.din(w_dff_A_LYwKI1nT2_0),.clk(gclk));
	jdff dff_A_DFMR8NpH6_0(.dout(w_dff_A_n3H0GgbP7_0),.din(w_dff_A_DFMR8NpH6_0),.clk(gclk));
	jdff dff_A_n3H0GgbP7_0(.dout(w_dff_A_WEIjJbIZ9_0),.din(w_dff_A_n3H0GgbP7_0),.clk(gclk));
	jdff dff_A_WEIjJbIZ9_0(.dout(w_dff_A_bJL5Zpll8_0),.din(w_dff_A_WEIjJbIZ9_0),.clk(gclk));
	jdff dff_A_bJL5Zpll8_0(.dout(w_dff_A_QvRfJ2HN2_0),.din(w_dff_A_bJL5Zpll8_0),.clk(gclk));
	jdff dff_A_QvRfJ2HN2_0(.dout(w_dff_A_W6CIbonm3_0),.din(w_dff_A_QvRfJ2HN2_0),.clk(gclk));
	jdff dff_A_W6CIbonm3_0(.dout(w_dff_A_DoZteobw0_0),.din(w_dff_A_W6CIbonm3_0),.clk(gclk));
	jdff dff_A_DoZteobw0_0(.dout(w_dff_A_7B6PW1H97_0),.din(w_dff_A_DoZteobw0_0),.clk(gclk));
	jdff dff_A_7B6PW1H97_0(.dout(w_dff_A_Glb9PYKR3_0),.din(w_dff_A_7B6PW1H97_0),.clk(gclk));
	jdff dff_A_Glb9PYKR3_0(.dout(w_dff_A_SWu8MAQi4_0),.din(w_dff_A_Glb9PYKR3_0),.clk(gclk));
	jdff dff_A_SWu8MAQi4_0(.dout(w_dff_A_ik55kIAn4_0),.din(w_dff_A_SWu8MAQi4_0),.clk(gclk));
	jdff dff_A_ik55kIAn4_0(.dout(w_dff_A_OA7tcb1Q1_0),.din(w_dff_A_ik55kIAn4_0),.clk(gclk));
	jdff dff_A_OA7tcb1Q1_0(.dout(w_dff_A_Pp6EtWCg9_0),.din(w_dff_A_OA7tcb1Q1_0),.clk(gclk));
	jdff dff_A_Pp6EtWCg9_0(.dout(w_dff_A_JOacAFEL0_0),.din(w_dff_A_Pp6EtWCg9_0),.clk(gclk));
	jdff dff_A_JOacAFEL0_0(.dout(w_dff_A_taAlJBcR7_0),.din(w_dff_A_JOacAFEL0_0),.clk(gclk));
	jdff dff_A_taAlJBcR7_0(.dout(w_dff_A_FlVssQCe7_0),.din(w_dff_A_taAlJBcR7_0),.clk(gclk));
	jdff dff_A_FlVssQCe7_0(.dout(w_dff_A_okKLQTvm0_0),.din(w_dff_A_FlVssQCe7_0),.clk(gclk));
	jdff dff_A_okKLQTvm0_0(.dout(w_dff_A_8nvJZ0Vo1_0),.din(w_dff_A_okKLQTvm0_0),.clk(gclk));
	jdff dff_A_8nvJZ0Vo1_0(.dout(w_dff_A_XsgQDMbk5_0),.din(w_dff_A_8nvJZ0Vo1_0),.clk(gclk));
	jdff dff_A_XsgQDMbk5_0(.dout(w_dff_A_F6EzjnPa6_0),.din(w_dff_A_XsgQDMbk5_0),.clk(gclk));
	jdff dff_A_F6EzjnPa6_0(.dout(w_dff_A_nDBPpSMl6_0),.din(w_dff_A_F6EzjnPa6_0),.clk(gclk));
	jdff dff_A_nDBPpSMl6_0(.dout(w_dff_A_n6jdrTl05_0),.din(w_dff_A_nDBPpSMl6_0),.clk(gclk));
	jdff dff_A_n6jdrTl05_0(.dout(w_dff_A_2AYU47VH7_0),.din(w_dff_A_n6jdrTl05_0),.clk(gclk));
	jdff dff_A_2AYU47VH7_0(.dout(w_dff_A_lITkqGhi2_0),.din(w_dff_A_2AYU47VH7_0),.clk(gclk));
	jdff dff_A_lITkqGhi2_0(.dout(w_dff_A_mPJxec0m8_0),.din(w_dff_A_lITkqGhi2_0),.clk(gclk));
	jdff dff_A_mPJxec0m8_0(.dout(w_dff_A_PydP6ym81_0),.din(w_dff_A_mPJxec0m8_0),.clk(gclk));
	jdff dff_A_PydP6ym81_0(.dout(w_dff_A_7B3GncZN1_0),.din(w_dff_A_PydP6ym81_0),.clk(gclk));
	jdff dff_A_7B3GncZN1_0(.dout(w_dff_A_lUPKBMOB1_0),.din(w_dff_A_7B3GncZN1_0),.clk(gclk));
	jdff dff_A_lUPKBMOB1_0(.dout(w_dff_A_71TYRVaG3_0),.din(w_dff_A_lUPKBMOB1_0),.clk(gclk));
	jdff dff_A_71TYRVaG3_0(.dout(w_dff_A_Vr0tPljX2_0),.din(w_dff_A_71TYRVaG3_0),.clk(gclk));
	jdff dff_A_Vr0tPljX2_0(.dout(w_dff_A_D7G1jR538_0),.din(w_dff_A_Vr0tPljX2_0),.clk(gclk));
	jdff dff_A_D7G1jR538_0(.dout(w_dff_A_zcL5PmoR3_0),.din(w_dff_A_D7G1jR538_0),.clk(gclk));
	jdff dff_A_zcL5PmoR3_0(.dout(w_dff_A_KQUOWqSc1_0),.din(w_dff_A_zcL5PmoR3_0),.clk(gclk));
	jdff dff_A_KQUOWqSc1_0(.dout(w_dff_A_KMp0WJip0_0),.din(w_dff_A_KQUOWqSc1_0),.clk(gclk));
	jdff dff_A_KMp0WJip0_0(.dout(w_dff_A_3y1YA1Oa6_0),.din(w_dff_A_KMp0WJip0_0),.clk(gclk));
	jdff dff_A_3y1YA1Oa6_0(.dout(w_dff_A_ly3ySnyv7_0),.din(w_dff_A_3y1YA1Oa6_0),.clk(gclk));
	jdff dff_A_ly3ySnyv7_0(.dout(w_dff_A_WXDRqHZG4_0),.din(w_dff_A_ly3ySnyv7_0),.clk(gclk));
	jdff dff_A_WXDRqHZG4_0(.dout(w_dff_A_msLZBPmv9_0),.din(w_dff_A_WXDRqHZG4_0),.clk(gclk));
	jdff dff_A_msLZBPmv9_0(.dout(w_dff_A_P1l6Dv7z1_0),.din(w_dff_A_msLZBPmv9_0),.clk(gclk));
	jdff dff_A_P1l6Dv7z1_0(.dout(w_dff_A_gzUGqGrS0_0),.din(w_dff_A_P1l6Dv7z1_0),.clk(gclk));
	jdff dff_A_gzUGqGrS0_0(.dout(w_dff_A_kv8RO6a14_0),.din(w_dff_A_gzUGqGrS0_0),.clk(gclk));
	jdff dff_A_kv8RO6a14_0(.dout(w_dff_A_p1jXc0CU5_0),.din(w_dff_A_kv8RO6a14_0),.clk(gclk));
	jdff dff_A_p1jXc0CU5_0(.dout(w_dff_A_3pnN2caj1_0),.din(w_dff_A_p1jXc0CU5_0),.clk(gclk));
	jdff dff_A_3pnN2caj1_0(.dout(G2877gat),.din(w_dff_A_3pnN2caj1_0),.clk(gclk));
	jdff dff_A_ML3PYmGw6_2(.dout(w_dff_A_k3hbTgbw1_0),.din(w_dff_A_ML3PYmGw6_2),.clk(gclk));
	jdff dff_A_k3hbTgbw1_0(.dout(w_dff_A_7gMWKem29_0),.din(w_dff_A_k3hbTgbw1_0),.clk(gclk));
	jdff dff_A_7gMWKem29_0(.dout(w_dff_A_OVagVgzt8_0),.din(w_dff_A_7gMWKem29_0),.clk(gclk));
	jdff dff_A_OVagVgzt8_0(.dout(w_dff_A_EQk1N8XE8_0),.din(w_dff_A_OVagVgzt8_0),.clk(gclk));
	jdff dff_A_EQk1N8XE8_0(.dout(w_dff_A_o5UxAA9t6_0),.din(w_dff_A_EQk1N8XE8_0),.clk(gclk));
	jdff dff_A_o5UxAA9t6_0(.dout(w_dff_A_4owISbqM2_0),.din(w_dff_A_o5UxAA9t6_0),.clk(gclk));
	jdff dff_A_4owISbqM2_0(.dout(w_dff_A_ifry3w2J0_0),.din(w_dff_A_4owISbqM2_0),.clk(gclk));
	jdff dff_A_ifry3w2J0_0(.dout(w_dff_A_19QwWR2D4_0),.din(w_dff_A_ifry3w2J0_0),.clk(gclk));
	jdff dff_A_19QwWR2D4_0(.dout(w_dff_A_Sz3kEFaI4_0),.din(w_dff_A_19QwWR2D4_0),.clk(gclk));
	jdff dff_A_Sz3kEFaI4_0(.dout(w_dff_A_8sPxZoJ60_0),.din(w_dff_A_Sz3kEFaI4_0),.clk(gclk));
	jdff dff_A_8sPxZoJ60_0(.dout(w_dff_A_OCHEaoC98_0),.din(w_dff_A_8sPxZoJ60_0),.clk(gclk));
	jdff dff_A_OCHEaoC98_0(.dout(w_dff_A_H6QVTEWY3_0),.din(w_dff_A_OCHEaoC98_0),.clk(gclk));
	jdff dff_A_H6QVTEWY3_0(.dout(w_dff_A_zaog7Hqm6_0),.din(w_dff_A_H6QVTEWY3_0),.clk(gclk));
	jdff dff_A_zaog7Hqm6_0(.dout(w_dff_A_IJpfjMiy3_0),.din(w_dff_A_zaog7Hqm6_0),.clk(gclk));
	jdff dff_A_IJpfjMiy3_0(.dout(w_dff_A_DUwSHHoa4_0),.din(w_dff_A_IJpfjMiy3_0),.clk(gclk));
	jdff dff_A_DUwSHHoa4_0(.dout(w_dff_A_ry5I9gVV6_0),.din(w_dff_A_DUwSHHoa4_0),.clk(gclk));
	jdff dff_A_ry5I9gVV6_0(.dout(w_dff_A_COyi6Itd1_0),.din(w_dff_A_ry5I9gVV6_0),.clk(gclk));
	jdff dff_A_COyi6Itd1_0(.dout(w_dff_A_yiq7gymJ9_0),.din(w_dff_A_COyi6Itd1_0),.clk(gclk));
	jdff dff_A_yiq7gymJ9_0(.dout(w_dff_A_eZsxtNCc5_0),.din(w_dff_A_yiq7gymJ9_0),.clk(gclk));
	jdff dff_A_eZsxtNCc5_0(.dout(w_dff_A_ocRW2mOu0_0),.din(w_dff_A_eZsxtNCc5_0),.clk(gclk));
	jdff dff_A_ocRW2mOu0_0(.dout(w_dff_A_f0w3GwGQ1_0),.din(w_dff_A_ocRW2mOu0_0),.clk(gclk));
	jdff dff_A_f0w3GwGQ1_0(.dout(w_dff_A_NdPr0yb54_0),.din(w_dff_A_f0w3GwGQ1_0),.clk(gclk));
	jdff dff_A_NdPr0yb54_0(.dout(w_dff_A_wm2ibPjd5_0),.din(w_dff_A_NdPr0yb54_0),.clk(gclk));
	jdff dff_A_wm2ibPjd5_0(.dout(w_dff_A_h9W6Xg6G7_0),.din(w_dff_A_wm2ibPjd5_0),.clk(gclk));
	jdff dff_A_h9W6Xg6G7_0(.dout(w_dff_A_P5ZI6iMN3_0),.din(w_dff_A_h9W6Xg6G7_0),.clk(gclk));
	jdff dff_A_P5ZI6iMN3_0(.dout(w_dff_A_t2s8Yrtq2_0),.din(w_dff_A_P5ZI6iMN3_0),.clk(gclk));
	jdff dff_A_t2s8Yrtq2_0(.dout(w_dff_A_1nzIiqnE1_0),.din(w_dff_A_t2s8Yrtq2_0),.clk(gclk));
	jdff dff_A_1nzIiqnE1_0(.dout(w_dff_A_d4HTecqI3_0),.din(w_dff_A_1nzIiqnE1_0),.clk(gclk));
	jdff dff_A_d4HTecqI3_0(.dout(w_dff_A_fk4qrDBu0_0),.din(w_dff_A_d4HTecqI3_0),.clk(gclk));
	jdff dff_A_fk4qrDBu0_0(.dout(w_dff_A_ox2hGdUL6_0),.din(w_dff_A_fk4qrDBu0_0),.clk(gclk));
	jdff dff_A_ox2hGdUL6_0(.dout(w_dff_A_VnKYrr3r1_0),.din(w_dff_A_ox2hGdUL6_0),.clk(gclk));
	jdff dff_A_VnKYrr3r1_0(.dout(w_dff_A_v7AsgOaS8_0),.din(w_dff_A_VnKYrr3r1_0),.clk(gclk));
	jdff dff_A_v7AsgOaS8_0(.dout(w_dff_A_J0SWVODD8_0),.din(w_dff_A_v7AsgOaS8_0),.clk(gclk));
	jdff dff_A_J0SWVODD8_0(.dout(w_dff_A_VjGxIN4R5_0),.din(w_dff_A_J0SWVODD8_0),.clk(gclk));
	jdff dff_A_VjGxIN4R5_0(.dout(w_dff_A_8jbEMAUT0_0),.din(w_dff_A_VjGxIN4R5_0),.clk(gclk));
	jdff dff_A_8jbEMAUT0_0(.dout(w_dff_A_59W2UrYY3_0),.din(w_dff_A_8jbEMAUT0_0),.clk(gclk));
	jdff dff_A_59W2UrYY3_0(.dout(w_dff_A_bMnUCCrQ0_0),.din(w_dff_A_59W2UrYY3_0),.clk(gclk));
	jdff dff_A_bMnUCCrQ0_0(.dout(w_dff_A_kKZM6Pi90_0),.din(w_dff_A_bMnUCCrQ0_0),.clk(gclk));
	jdff dff_A_kKZM6Pi90_0(.dout(w_dff_A_CgrReBRv0_0),.din(w_dff_A_kKZM6Pi90_0),.clk(gclk));
	jdff dff_A_CgrReBRv0_0(.dout(w_dff_A_7Icgqo6H8_0),.din(w_dff_A_CgrReBRv0_0),.clk(gclk));
	jdff dff_A_7Icgqo6H8_0(.dout(w_dff_A_iNriN8iw9_0),.din(w_dff_A_7Icgqo6H8_0),.clk(gclk));
	jdff dff_A_iNriN8iw9_0(.dout(w_dff_A_9hdkHlNi4_0),.din(w_dff_A_iNriN8iw9_0),.clk(gclk));
	jdff dff_A_9hdkHlNi4_0(.dout(w_dff_A_Ok6iiI9m3_0),.din(w_dff_A_9hdkHlNi4_0),.clk(gclk));
	jdff dff_A_Ok6iiI9m3_0(.dout(w_dff_A_wI49MFMv7_0),.din(w_dff_A_Ok6iiI9m3_0),.clk(gclk));
	jdff dff_A_wI49MFMv7_0(.dout(w_dff_A_A47xoUlP6_0),.din(w_dff_A_wI49MFMv7_0),.clk(gclk));
	jdff dff_A_A47xoUlP6_0(.dout(w_dff_A_asAKRf9w1_0),.din(w_dff_A_A47xoUlP6_0),.clk(gclk));
	jdff dff_A_asAKRf9w1_0(.dout(w_dff_A_XtuG2nkg8_0),.din(w_dff_A_asAKRf9w1_0),.clk(gclk));
	jdff dff_A_XtuG2nkg8_0(.dout(w_dff_A_kTzuItIH0_0),.din(w_dff_A_XtuG2nkg8_0),.clk(gclk));
	jdff dff_A_kTzuItIH0_0(.dout(w_dff_A_kcLgxgPP7_0),.din(w_dff_A_kTzuItIH0_0),.clk(gclk));
	jdff dff_A_kcLgxgPP7_0(.dout(w_dff_A_4HfSNL7E7_0),.din(w_dff_A_kcLgxgPP7_0),.clk(gclk));
	jdff dff_A_4HfSNL7E7_0(.dout(w_dff_A_bhTdnMuf2_0),.din(w_dff_A_4HfSNL7E7_0),.clk(gclk));
	jdff dff_A_bhTdnMuf2_0(.dout(w_dff_A_mV8wK1155_0),.din(w_dff_A_bhTdnMuf2_0),.clk(gclk));
	jdff dff_A_mV8wK1155_0(.dout(w_dff_A_ePVaFnM57_0),.din(w_dff_A_mV8wK1155_0),.clk(gclk));
	jdff dff_A_ePVaFnM57_0(.dout(w_dff_A_SpgU20S39_0),.din(w_dff_A_ePVaFnM57_0),.clk(gclk));
	jdff dff_A_SpgU20S39_0(.dout(w_dff_A_GPpo5IbF2_0),.din(w_dff_A_SpgU20S39_0),.clk(gclk));
	jdff dff_A_GPpo5IbF2_0(.dout(w_dff_A_F81vDXYA9_0),.din(w_dff_A_GPpo5IbF2_0),.clk(gclk));
	jdff dff_A_F81vDXYA9_0(.dout(G3211gat),.din(w_dff_A_F81vDXYA9_0),.clk(gclk));
	jdff dff_A_p8CWdcT47_2(.dout(w_dff_A_vIN3fXLZ2_0),.din(w_dff_A_p8CWdcT47_2),.clk(gclk));
	jdff dff_A_vIN3fXLZ2_0(.dout(w_dff_A_murdQeTr3_0),.din(w_dff_A_vIN3fXLZ2_0),.clk(gclk));
	jdff dff_A_murdQeTr3_0(.dout(w_dff_A_qyRBVjgt4_0),.din(w_dff_A_murdQeTr3_0),.clk(gclk));
	jdff dff_A_qyRBVjgt4_0(.dout(w_dff_A_UWdhPYhA8_0),.din(w_dff_A_qyRBVjgt4_0),.clk(gclk));
	jdff dff_A_UWdhPYhA8_0(.dout(w_dff_A_Zc4eXUwU6_0),.din(w_dff_A_UWdhPYhA8_0),.clk(gclk));
	jdff dff_A_Zc4eXUwU6_0(.dout(w_dff_A_Mc8Wha1q2_0),.din(w_dff_A_Zc4eXUwU6_0),.clk(gclk));
	jdff dff_A_Mc8Wha1q2_0(.dout(w_dff_A_VsphuY9H5_0),.din(w_dff_A_Mc8Wha1q2_0),.clk(gclk));
	jdff dff_A_VsphuY9H5_0(.dout(w_dff_A_HX2q0STK3_0),.din(w_dff_A_VsphuY9H5_0),.clk(gclk));
	jdff dff_A_HX2q0STK3_0(.dout(w_dff_A_8mvjjQ8w0_0),.din(w_dff_A_HX2q0STK3_0),.clk(gclk));
	jdff dff_A_8mvjjQ8w0_0(.dout(w_dff_A_bqESm2l63_0),.din(w_dff_A_8mvjjQ8w0_0),.clk(gclk));
	jdff dff_A_bqESm2l63_0(.dout(w_dff_A_5Nl4WnvC9_0),.din(w_dff_A_bqESm2l63_0),.clk(gclk));
	jdff dff_A_5Nl4WnvC9_0(.dout(w_dff_A_ykxwu6cd3_0),.din(w_dff_A_5Nl4WnvC9_0),.clk(gclk));
	jdff dff_A_ykxwu6cd3_0(.dout(w_dff_A_lhpgddm69_0),.din(w_dff_A_ykxwu6cd3_0),.clk(gclk));
	jdff dff_A_lhpgddm69_0(.dout(w_dff_A_CWkLmZ9f6_0),.din(w_dff_A_lhpgddm69_0),.clk(gclk));
	jdff dff_A_CWkLmZ9f6_0(.dout(w_dff_A_a0rjBk531_0),.din(w_dff_A_CWkLmZ9f6_0),.clk(gclk));
	jdff dff_A_a0rjBk531_0(.dout(w_dff_A_2iedVuis6_0),.din(w_dff_A_a0rjBk531_0),.clk(gclk));
	jdff dff_A_2iedVuis6_0(.dout(w_dff_A_2GNJRJN49_0),.din(w_dff_A_2iedVuis6_0),.clk(gclk));
	jdff dff_A_2GNJRJN49_0(.dout(w_dff_A_ENcapxbA2_0),.din(w_dff_A_2GNJRJN49_0),.clk(gclk));
	jdff dff_A_ENcapxbA2_0(.dout(w_dff_A_E7uQrMF42_0),.din(w_dff_A_ENcapxbA2_0),.clk(gclk));
	jdff dff_A_E7uQrMF42_0(.dout(w_dff_A_3xiSwC5F9_0),.din(w_dff_A_E7uQrMF42_0),.clk(gclk));
	jdff dff_A_3xiSwC5F9_0(.dout(w_dff_A_svNWcnZz2_0),.din(w_dff_A_3xiSwC5F9_0),.clk(gclk));
	jdff dff_A_svNWcnZz2_0(.dout(w_dff_A_6rhR35bC2_0),.din(w_dff_A_svNWcnZz2_0),.clk(gclk));
	jdff dff_A_6rhR35bC2_0(.dout(w_dff_A_n736qRW58_0),.din(w_dff_A_6rhR35bC2_0),.clk(gclk));
	jdff dff_A_n736qRW58_0(.dout(w_dff_A_9ixB6Oj44_0),.din(w_dff_A_n736qRW58_0),.clk(gclk));
	jdff dff_A_9ixB6Oj44_0(.dout(w_dff_A_TSPdbDcl6_0),.din(w_dff_A_9ixB6Oj44_0),.clk(gclk));
	jdff dff_A_TSPdbDcl6_0(.dout(w_dff_A_EOI67Sd87_0),.din(w_dff_A_TSPdbDcl6_0),.clk(gclk));
	jdff dff_A_EOI67Sd87_0(.dout(w_dff_A_BSHQMDeF5_0),.din(w_dff_A_EOI67Sd87_0),.clk(gclk));
	jdff dff_A_BSHQMDeF5_0(.dout(w_dff_A_dku6XVqK9_0),.din(w_dff_A_BSHQMDeF5_0),.clk(gclk));
	jdff dff_A_dku6XVqK9_0(.dout(w_dff_A_4IISccVA9_0),.din(w_dff_A_dku6XVqK9_0),.clk(gclk));
	jdff dff_A_4IISccVA9_0(.dout(w_dff_A_vCWreVNQ1_0),.din(w_dff_A_4IISccVA9_0),.clk(gclk));
	jdff dff_A_vCWreVNQ1_0(.dout(w_dff_A_7blmHrjB1_0),.din(w_dff_A_vCWreVNQ1_0),.clk(gclk));
	jdff dff_A_7blmHrjB1_0(.dout(w_dff_A_a6ZhVuG86_0),.din(w_dff_A_7blmHrjB1_0),.clk(gclk));
	jdff dff_A_a6ZhVuG86_0(.dout(w_dff_A_WmshASpB0_0),.din(w_dff_A_a6ZhVuG86_0),.clk(gclk));
	jdff dff_A_WmshASpB0_0(.dout(w_dff_A_eviCvvc00_0),.din(w_dff_A_WmshASpB0_0),.clk(gclk));
	jdff dff_A_eviCvvc00_0(.dout(w_dff_A_vvNLWVY49_0),.din(w_dff_A_eviCvvc00_0),.clk(gclk));
	jdff dff_A_vvNLWVY49_0(.dout(w_dff_A_2uH30iFi9_0),.din(w_dff_A_vvNLWVY49_0),.clk(gclk));
	jdff dff_A_2uH30iFi9_0(.dout(w_dff_A_73Jy1lAO5_0),.din(w_dff_A_2uH30iFi9_0),.clk(gclk));
	jdff dff_A_73Jy1lAO5_0(.dout(w_dff_A_IWyQhmTp6_0),.din(w_dff_A_73Jy1lAO5_0),.clk(gclk));
	jdff dff_A_IWyQhmTp6_0(.dout(w_dff_A_QGZRqCOG2_0),.din(w_dff_A_IWyQhmTp6_0),.clk(gclk));
	jdff dff_A_QGZRqCOG2_0(.dout(w_dff_A_O2pv5VvY8_0),.din(w_dff_A_QGZRqCOG2_0),.clk(gclk));
	jdff dff_A_O2pv5VvY8_0(.dout(w_dff_A_5kDnpyuh7_0),.din(w_dff_A_O2pv5VvY8_0),.clk(gclk));
	jdff dff_A_5kDnpyuh7_0(.dout(w_dff_A_4bAvnC9u7_0),.din(w_dff_A_5kDnpyuh7_0),.clk(gclk));
	jdff dff_A_4bAvnC9u7_0(.dout(w_dff_A_CSfaVj1b3_0),.din(w_dff_A_4bAvnC9u7_0),.clk(gclk));
	jdff dff_A_CSfaVj1b3_0(.dout(w_dff_A_j2OmXIcK8_0),.din(w_dff_A_CSfaVj1b3_0),.clk(gclk));
	jdff dff_A_j2OmXIcK8_0(.dout(w_dff_A_nSO9w3xe7_0),.din(w_dff_A_j2OmXIcK8_0),.clk(gclk));
	jdff dff_A_nSO9w3xe7_0(.dout(w_dff_A_uzzkA84e1_0),.din(w_dff_A_nSO9w3xe7_0),.clk(gclk));
	jdff dff_A_uzzkA84e1_0(.dout(w_dff_A_1EyFcUot8_0),.din(w_dff_A_uzzkA84e1_0),.clk(gclk));
	jdff dff_A_1EyFcUot8_0(.dout(w_dff_A_wMQ1QNGZ9_0),.din(w_dff_A_1EyFcUot8_0),.clk(gclk));
	jdff dff_A_wMQ1QNGZ9_0(.dout(w_dff_A_BA22Zhw80_0),.din(w_dff_A_wMQ1QNGZ9_0),.clk(gclk));
	jdff dff_A_BA22Zhw80_0(.dout(w_dff_A_qM72JduN4_0),.din(w_dff_A_BA22Zhw80_0),.clk(gclk));
	jdff dff_A_qM72JduN4_0(.dout(w_dff_A_0iRaUxIe4_0),.din(w_dff_A_qM72JduN4_0),.clk(gclk));
	jdff dff_A_0iRaUxIe4_0(.dout(w_dff_A_c7RE4A0A9_0),.din(w_dff_A_0iRaUxIe4_0),.clk(gclk));
	jdff dff_A_c7RE4A0A9_0(.dout(w_dff_A_5JwUzXPA2_0),.din(w_dff_A_c7RE4A0A9_0),.clk(gclk));
	jdff dff_A_5JwUzXPA2_0(.dout(G3552gat),.din(w_dff_A_5JwUzXPA2_0),.clk(gclk));
	jdff dff_A_aV8fpFrx0_2(.dout(w_dff_A_0U1eS1Nh1_0),.din(w_dff_A_aV8fpFrx0_2),.clk(gclk));
	jdff dff_A_0U1eS1Nh1_0(.dout(w_dff_A_XciRZcPX6_0),.din(w_dff_A_0U1eS1Nh1_0),.clk(gclk));
	jdff dff_A_XciRZcPX6_0(.dout(w_dff_A_dNsXdzoD6_0),.din(w_dff_A_XciRZcPX6_0),.clk(gclk));
	jdff dff_A_dNsXdzoD6_0(.dout(w_dff_A_DF4r45PI4_0),.din(w_dff_A_dNsXdzoD6_0),.clk(gclk));
	jdff dff_A_DF4r45PI4_0(.dout(w_dff_A_6ib9vVbp3_0),.din(w_dff_A_DF4r45PI4_0),.clk(gclk));
	jdff dff_A_6ib9vVbp3_0(.dout(w_dff_A_QbC4MRD40_0),.din(w_dff_A_6ib9vVbp3_0),.clk(gclk));
	jdff dff_A_QbC4MRD40_0(.dout(w_dff_A_rllvemIL9_0),.din(w_dff_A_QbC4MRD40_0),.clk(gclk));
	jdff dff_A_rllvemIL9_0(.dout(w_dff_A_cmiqokas9_0),.din(w_dff_A_rllvemIL9_0),.clk(gclk));
	jdff dff_A_cmiqokas9_0(.dout(w_dff_A_0aT3jov38_0),.din(w_dff_A_cmiqokas9_0),.clk(gclk));
	jdff dff_A_0aT3jov38_0(.dout(w_dff_A_Xjz9riNF7_0),.din(w_dff_A_0aT3jov38_0),.clk(gclk));
	jdff dff_A_Xjz9riNF7_0(.dout(w_dff_A_wZ7XgEnk5_0),.din(w_dff_A_Xjz9riNF7_0),.clk(gclk));
	jdff dff_A_wZ7XgEnk5_0(.dout(w_dff_A_jvj58AaU0_0),.din(w_dff_A_wZ7XgEnk5_0),.clk(gclk));
	jdff dff_A_jvj58AaU0_0(.dout(w_dff_A_WGrBtmzJ3_0),.din(w_dff_A_jvj58AaU0_0),.clk(gclk));
	jdff dff_A_WGrBtmzJ3_0(.dout(w_dff_A_qrnMsTzN6_0),.din(w_dff_A_WGrBtmzJ3_0),.clk(gclk));
	jdff dff_A_qrnMsTzN6_0(.dout(w_dff_A_IXZ4RphD5_0),.din(w_dff_A_qrnMsTzN6_0),.clk(gclk));
	jdff dff_A_IXZ4RphD5_0(.dout(w_dff_A_nDQT0Bqm9_0),.din(w_dff_A_IXZ4RphD5_0),.clk(gclk));
	jdff dff_A_nDQT0Bqm9_0(.dout(w_dff_A_7DxEEq538_0),.din(w_dff_A_nDQT0Bqm9_0),.clk(gclk));
	jdff dff_A_7DxEEq538_0(.dout(w_dff_A_VMbF0QFq1_0),.din(w_dff_A_7DxEEq538_0),.clk(gclk));
	jdff dff_A_VMbF0QFq1_0(.dout(w_dff_A_0h7Rnq0j9_0),.din(w_dff_A_VMbF0QFq1_0),.clk(gclk));
	jdff dff_A_0h7Rnq0j9_0(.dout(w_dff_A_tObv25cz7_0),.din(w_dff_A_0h7Rnq0j9_0),.clk(gclk));
	jdff dff_A_tObv25cz7_0(.dout(w_dff_A_edY2CSKo7_0),.din(w_dff_A_tObv25cz7_0),.clk(gclk));
	jdff dff_A_edY2CSKo7_0(.dout(w_dff_A_rcOxops84_0),.din(w_dff_A_edY2CSKo7_0),.clk(gclk));
	jdff dff_A_rcOxops84_0(.dout(w_dff_A_1XIZFMrL2_0),.din(w_dff_A_rcOxops84_0),.clk(gclk));
	jdff dff_A_1XIZFMrL2_0(.dout(w_dff_A_DecREavl0_0),.din(w_dff_A_1XIZFMrL2_0),.clk(gclk));
	jdff dff_A_DecREavl0_0(.dout(w_dff_A_ZnuiK6Me8_0),.din(w_dff_A_DecREavl0_0),.clk(gclk));
	jdff dff_A_ZnuiK6Me8_0(.dout(w_dff_A_V9Z3Fxt27_0),.din(w_dff_A_ZnuiK6Me8_0),.clk(gclk));
	jdff dff_A_V9Z3Fxt27_0(.dout(w_dff_A_XGxsuKCA0_0),.din(w_dff_A_V9Z3Fxt27_0),.clk(gclk));
	jdff dff_A_XGxsuKCA0_0(.dout(w_dff_A_jSFjKJnA5_0),.din(w_dff_A_XGxsuKCA0_0),.clk(gclk));
	jdff dff_A_jSFjKJnA5_0(.dout(w_dff_A_OBHTPb8G3_0),.din(w_dff_A_jSFjKJnA5_0),.clk(gclk));
	jdff dff_A_OBHTPb8G3_0(.dout(w_dff_A_hrMPtjRC3_0),.din(w_dff_A_OBHTPb8G3_0),.clk(gclk));
	jdff dff_A_hrMPtjRC3_0(.dout(w_dff_A_BEbtPiKp7_0),.din(w_dff_A_hrMPtjRC3_0),.clk(gclk));
	jdff dff_A_BEbtPiKp7_0(.dout(w_dff_A_fuPxVhmE3_0),.din(w_dff_A_BEbtPiKp7_0),.clk(gclk));
	jdff dff_A_fuPxVhmE3_0(.dout(w_dff_A_sxaPDRBN3_0),.din(w_dff_A_fuPxVhmE3_0),.clk(gclk));
	jdff dff_A_sxaPDRBN3_0(.dout(w_dff_A_FIHiv3Lw1_0),.din(w_dff_A_sxaPDRBN3_0),.clk(gclk));
	jdff dff_A_FIHiv3Lw1_0(.dout(w_dff_A_nYZZPLxt4_0),.din(w_dff_A_FIHiv3Lw1_0),.clk(gclk));
	jdff dff_A_nYZZPLxt4_0(.dout(w_dff_A_HKSJ8cgS3_0),.din(w_dff_A_nYZZPLxt4_0),.clk(gclk));
	jdff dff_A_HKSJ8cgS3_0(.dout(w_dff_A_oefFO2oq7_0),.din(w_dff_A_HKSJ8cgS3_0),.clk(gclk));
	jdff dff_A_oefFO2oq7_0(.dout(w_dff_A_kywkKTac8_0),.din(w_dff_A_oefFO2oq7_0),.clk(gclk));
	jdff dff_A_kywkKTac8_0(.dout(w_dff_A_u6LAQU9n0_0),.din(w_dff_A_kywkKTac8_0),.clk(gclk));
	jdff dff_A_u6LAQU9n0_0(.dout(w_dff_A_qyUEWSpa9_0),.din(w_dff_A_u6LAQU9n0_0),.clk(gclk));
	jdff dff_A_qyUEWSpa9_0(.dout(w_dff_A_nVfuuVEZ5_0),.din(w_dff_A_qyUEWSpa9_0),.clk(gclk));
	jdff dff_A_nVfuuVEZ5_0(.dout(w_dff_A_y3Mg9dp28_0),.din(w_dff_A_nVfuuVEZ5_0),.clk(gclk));
	jdff dff_A_y3Mg9dp28_0(.dout(w_dff_A_EJNd4H0Z3_0),.din(w_dff_A_y3Mg9dp28_0),.clk(gclk));
	jdff dff_A_EJNd4H0Z3_0(.dout(w_dff_A_MvZc0U2H5_0),.din(w_dff_A_EJNd4H0Z3_0),.clk(gclk));
	jdff dff_A_MvZc0U2H5_0(.dout(w_dff_A_R8zNVeUO6_0),.din(w_dff_A_MvZc0U2H5_0),.clk(gclk));
	jdff dff_A_R8zNVeUO6_0(.dout(w_dff_A_S69efoHJ6_0),.din(w_dff_A_R8zNVeUO6_0),.clk(gclk));
	jdff dff_A_S69efoHJ6_0(.dout(w_dff_A_vYthnCn77_0),.din(w_dff_A_S69efoHJ6_0),.clk(gclk));
	jdff dff_A_vYthnCn77_0(.dout(w_dff_A_dRhvuoNw9_0),.din(w_dff_A_vYthnCn77_0),.clk(gclk));
	jdff dff_A_dRhvuoNw9_0(.dout(w_dff_A_nk5z5N5r8_0),.din(w_dff_A_dRhvuoNw9_0),.clk(gclk));
	jdff dff_A_nk5z5N5r8_0(.dout(w_dff_A_9vRoFg8j0_0),.din(w_dff_A_nk5z5N5r8_0),.clk(gclk));
	jdff dff_A_9vRoFg8j0_0(.dout(G3895gat),.din(w_dff_A_9vRoFg8j0_0),.clk(gclk));
	jdff dff_A_xLPUpw6m3_2(.dout(w_dff_A_QK12NJAC1_0),.din(w_dff_A_xLPUpw6m3_2),.clk(gclk));
	jdff dff_A_QK12NJAC1_0(.dout(w_dff_A_QcGeXnrj0_0),.din(w_dff_A_QK12NJAC1_0),.clk(gclk));
	jdff dff_A_QcGeXnrj0_0(.dout(w_dff_A_odvBaEmS8_0),.din(w_dff_A_QcGeXnrj0_0),.clk(gclk));
	jdff dff_A_odvBaEmS8_0(.dout(w_dff_A_78ghDAb57_0),.din(w_dff_A_odvBaEmS8_0),.clk(gclk));
	jdff dff_A_78ghDAb57_0(.dout(w_dff_A_OQNNHVWy1_0),.din(w_dff_A_78ghDAb57_0),.clk(gclk));
	jdff dff_A_OQNNHVWy1_0(.dout(w_dff_A_GMTVX1TR2_0),.din(w_dff_A_OQNNHVWy1_0),.clk(gclk));
	jdff dff_A_GMTVX1TR2_0(.dout(w_dff_A_f5UPQVK13_0),.din(w_dff_A_GMTVX1TR2_0),.clk(gclk));
	jdff dff_A_f5UPQVK13_0(.dout(w_dff_A_DcUF1SkU7_0),.din(w_dff_A_f5UPQVK13_0),.clk(gclk));
	jdff dff_A_DcUF1SkU7_0(.dout(w_dff_A_UtNgAUgX5_0),.din(w_dff_A_DcUF1SkU7_0),.clk(gclk));
	jdff dff_A_UtNgAUgX5_0(.dout(w_dff_A_khITjU2X8_0),.din(w_dff_A_UtNgAUgX5_0),.clk(gclk));
	jdff dff_A_khITjU2X8_0(.dout(w_dff_A_i0QThDGl5_0),.din(w_dff_A_khITjU2X8_0),.clk(gclk));
	jdff dff_A_i0QThDGl5_0(.dout(w_dff_A_Y6p5te3r2_0),.din(w_dff_A_i0QThDGl5_0),.clk(gclk));
	jdff dff_A_Y6p5te3r2_0(.dout(w_dff_A_dMnp0QqG2_0),.din(w_dff_A_Y6p5te3r2_0),.clk(gclk));
	jdff dff_A_dMnp0QqG2_0(.dout(w_dff_A_3em5remO9_0),.din(w_dff_A_dMnp0QqG2_0),.clk(gclk));
	jdff dff_A_3em5remO9_0(.dout(w_dff_A_7GrAzDZs5_0),.din(w_dff_A_3em5remO9_0),.clk(gclk));
	jdff dff_A_7GrAzDZs5_0(.dout(w_dff_A_Q0WNY1Xl4_0),.din(w_dff_A_7GrAzDZs5_0),.clk(gclk));
	jdff dff_A_Q0WNY1Xl4_0(.dout(w_dff_A_JL52Oqix5_0),.din(w_dff_A_Q0WNY1Xl4_0),.clk(gclk));
	jdff dff_A_JL52Oqix5_0(.dout(w_dff_A_nuzg1xGW4_0),.din(w_dff_A_JL52Oqix5_0),.clk(gclk));
	jdff dff_A_nuzg1xGW4_0(.dout(w_dff_A_RCarGdSy2_0),.din(w_dff_A_nuzg1xGW4_0),.clk(gclk));
	jdff dff_A_RCarGdSy2_0(.dout(w_dff_A_K5rHSPpA1_0),.din(w_dff_A_RCarGdSy2_0),.clk(gclk));
	jdff dff_A_K5rHSPpA1_0(.dout(w_dff_A_HHMFfhmR4_0),.din(w_dff_A_K5rHSPpA1_0),.clk(gclk));
	jdff dff_A_HHMFfhmR4_0(.dout(w_dff_A_S6AS7W723_0),.din(w_dff_A_HHMFfhmR4_0),.clk(gclk));
	jdff dff_A_S6AS7W723_0(.dout(w_dff_A_zZNXjYWQ1_0),.din(w_dff_A_S6AS7W723_0),.clk(gclk));
	jdff dff_A_zZNXjYWQ1_0(.dout(w_dff_A_0Pawiz2H8_0),.din(w_dff_A_zZNXjYWQ1_0),.clk(gclk));
	jdff dff_A_0Pawiz2H8_0(.dout(w_dff_A_ZOqTnZRI1_0),.din(w_dff_A_0Pawiz2H8_0),.clk(gclk));
	jdff dff_A_ZOqTnZRI1_0(.dout(w_dff_A_frzqTFQU7_0),.din(w_dff_A_ZOqTnZRI1_0),.clk(gclk));
	jdff dff_A_frzqTFQU7_0(.dout(w_dff_A_ztZV15So3_0),.din(w_dff_A_frzqTFQU7_0),.clk(gclk));
	jdff dff_A_ztZV15So3_0(.dout(w_dff_A_zRR3ME1v8_0),.din(w_dff_A_ztZV15So3_0),.clk(gclk));
	jdff dff_A_zRR3ME1v8_0(.dout(w_dff_A_YlS9cwIT6_0),.din(w_dff_A_zRR3ME1v8_0),.clk(gclk));
	jdff dff_A_YlS9cwIT6_0(.dout(w_dff_A_RtBY4bb97_0),.din(w_dff_A_YlS9cwIT6_0),.clk(gclk));
	jdff dff_A_RtBY4bb97_0(.dout(w_dff_A_CVak30a55_0),.din(w_dff_A_RtBY4bb97_0),.clk(gclk));
	jdff dff_A_CVak30a55_0(.dout(w_dff_A_AwjAA4Kz2_0),.din(w_dff_A_CVak30a55_0),.clk(gclk));
	jdff dff_A_AwjAA4Kz2_0(.dout(w_dff_A_q6EBBycg5_0),.din(w_dff_A_AwjAA4Kz2_0),.clk(gclk));
	jdff dff_A_q6EBBycg5_0(.dout(w_dff_A_YQ6ZgHCP2_0),.din(w_dff_A_q6EBBycg5_0),.clk(gclk));
	jdff dff_A_YQ6ZgHCP2_0(.dout(w_dff_A_l6TnnlmD7_0),.din(w_dff_A_YQ6ZgHCP2_0),.clk(gclk));
	jdff dff_A_l6TnnlmD7_0(.dout(w_dff_A_zLhYjaVg5_0),.din(w_dff_A_l6TnnlmD7_0),.clk(gclk));
	jdff dff_A_zLhYjaVg5_0(.dout(w_dff_A_r6EIwhAa1_0),.din(w_dff_A_zLhYjaVg5_0),.clk(gclk));
	jdff dff_A_r6EIwhAa1_0(.dout(w_dff_A_XYCROZpX6_0),.din(w_dff_A_r6EIwhAa1_0),.clk(gclk));
	jdff dff_A_XYCROZpX6_0(.dout(w_dff_A_3n2ABVn97_0),.din(w_dff_A_XYCROZpX6_0),.clk(gclk));
	jdff dff_A_3n2ABVn97_0(.dout(w_dff_A_N2Jlv2Hl5_0),.din(w_dff_A_3n2ABVn97_0),.clk(gclk));
	jdff dff_A_N2Jlv2Hl5_0(.dout(w_dff_A_1xRXt6jg0_0),.din(w_dff_A_N2Jlv2Hl5_0),.clk(gclk));
	jdff dff_A_1xRXt6jg0_0(.dout(w_dff_A_N3chEZbv8_0),.din(w_dff_A_1xRXt6jg0_0),.clk(gclk));
	jdff dff_A_N3chEZbv8_0(.dout(w_dff_A_5XDC8Sma9_0),.din(w_dff_A_N3chEZbv8_0),.clk(gclk));
	jdff dff_A_5XDC8Sma9_0(.dout(w_dff_A_9pOJfBB00_0),.din(w_dff_A_5XDC8Sma9_0),.clk(gclk));
	jdff dff_A_9pOJfBB00_0(.dout(w_dff_A_APiTgBJb5_0),.din(w_dff_A_9pOJfBB00_0),.clk(gclk));
	jdff dff_A_APiTgBJb5_0(.dout(w_dff_A_ZVkuoleY1_0),.din(w_dff_A_APiTgBJb5_0),.clk(gclk));
	jdff dff_A_ZVkuoleY1_0(.dout(w_dff_A_GgZyM2mP0_0),.din(w_dff_A_ZVkuoleY1_0),.clk(gclk));
	jdff dff_A_GgZyM2mP0_0(.dout(G4241gat),.din(w_dff_A_GgZyM2mP0_0),.clk(gclk));
	jdff dff_A_0FjbwSqr7_2(.dout(w_dff_A_v2NlOv3r7_0),.din(w_dff_A_0FjbwSqr7_2),.clk(gclk));
	jdff dff_A_v2NlOv3r7_0(.dout(w_dff_A_vXtYIMoI8_0),.din(w_dff_A_v2NlOv3r7_0),.clk(gclk));
	jdff dff_A_vXtYIMoI8_0(.dout(w_dff_A_fWjPS95U8_0),.din(w_dff_A_vXtYIMoI8_0),.clk(gclk));
	jdff dff_A_fWjPS95U8_0(.dout(w_dff_A_shWmwZ4i6_0),.din(w_dff_A_fWjPS95U8_0),.clk(gclk));
	jdff dff_A_shWmwZ4i6_0(.dout(w_dff_A_vAk4AwuO0_0),.din(w_dff_A_shWmwZ4i6_0),.clk(gclk));
	jdff dff_A_vAk4AwuO0_0(.dout(w_dff_A_j3ZrDR6t3_0),.din(w_dff_A_vAk4AwuO0_0),.clk(gclk));
	jdff dff_A_j3ZrDR6t3_0(.dout(w_dff_A_Ovwf8QUQ8_0),.din(w_dff_A_j3ZrDR6t3_0),.clk(gclk));
	jdff dff_A_Ovwf8QUQ8_0(.dout(w_dff_A_Nf3Q58to4_0),.din(w_dff_A_Ovwf8QUQ8_0),.clk(gclk));
	jdff dff_A_Nf3Q58to4_0(.dout(w_dff_A_UrFSKH9n3_0),.din(w_dff_A_Nf3Q58to4_0),.clk(gclk));
	jdff dff_A_UrFSKH9n3_0(.dout(w_dff_A_BURDr2196_0),.din(w_dff_A_UrFSKH9n3_0),.clk(gclk));
	jdff dff_A_BURDr2196_0(.dout(w_dff_A_ujZTwe5P2_0),.din(w_dff_A_BURDr2196_0),.clk(gclk));
	jdff dff_A_ujZTwe5P2_0(.dout(w_dff_A_ugvHRZPQ8_0),.din(w_dff_A_ujZTwe5P2_0),.clk(gclk));
	jdff dff_A_ugvHRZPQ8_0(.dout(w_dff_A_ptqPrW0t5_0),.din(w_dff_A_ugvHRZPQ8_0),.clk(gclk));
	jdff dff_A_ptqPrW0t5_0(.dout(w_dff_A_D3V15u9R0_0),.din(w_dff_A_ptqPrW0t5_0),.clk(gclk));
	jdff dff_A_D3V15u9R0_0(.dout(w_dff_A_10xftJvC4_0),.din(w_dff_A_D3V15u9R0_0),.clk(gclk));
	jdff dff_A_10xftJvC4_0(.dout(w_dff_A_3jvctEhx4_0),.din(w_dff_A_10xftJvC4_0),.clk(gclk));
	jdff dff_A_3jvctEhx4_0(.dout(w_dff_A_Sd4w4de37_0),.din(w_dff_A_3jvctEhx4_0),.clk(gclk));
	jdff dff_A_Sd4w4de37_0(.dout(w_dff_A_SUDhWvOt1_0),.din(w_dff_A_Sd4w4de37_0),.clk(gclk));
	jdff dff_A_SUDhWvOt1_0(.dout(w_dff_A_ACkv5MI83_0),.din(w_dff_A_SUDhWvOt1_0),.clk(gclk));
	jdff dff_A_ACkv5MI83_0(.dout(w_dff_A_AkXJFaCi0_0),.din(w_dff_A_ACkv5MI83_0),.clk(gclk));
	jdff dff_A_AkXJFaCi0_0(.dout(w_dff_A_DcwAzE9I1_0),.din(w_dff_A_AkXJFaCi0_0),.clk(gclk));
	jdff dff_A_DcwAzE9I1_0(.dout(w_dff_A_BjJMKzPh1_0),.din(w_dff_A_DcwAzE9I1_0),.clk(gclk));
	jdff dff_A_BjJMKzPh1_0(.dout(w_dff_A_Wri9CrDy5_0),.din(w_dff_A_BjJMKzPh1_0),.clk(gclk));
	jdff dff_A_Wri9CrDy5_0(.dout(w_dff_A_fPcFWY5b5_0),.din(w_dff_A_Wri9CrDy5_0),.clk(gclk));
	jdff dff_A_fPcFWY5b5_0(.dout(w_dff_A_xf7iYQEE1_0),.din(w_dff_A_fPcFWY5b5_0),.clk(gclk));
	jdff dff_A_xf7iYQEE1_0(.dout(w_dff_A_hJst8t655_0),.din(w_dff_A_xf7iYQEE1_0),.clk(gclk));
	jdff dff_A_hJst8t655_0(.dout(w_dff_A_66b8KN7Z9_0),.din(w_dff_A_hJst8t655_0),.clk(gclk));
	jdff dff_A_66b8KN7Z9_0(.dout(w_dff_A_pfcZH3Ke6_0),.din(w_dff_A_66b8KN7Z9_0),.clk(gclk));
	jdff dff_A_pfcZH3Ke6_0(.dout(w_dff_A_vdcsjvKF9_0),.din(w_dff_A_pfcZH3Ke6_0),.clk(gclk));
	jdff dff_A_vdcsjvKF9_0(.dout(w_dff_A_QBNhy4Oo8_0),.din(w_dff_A_vdcsjvKF9_0),.clk(gclk));
	jdff dff_A_QBNhy4Oo8_0(.dout(w_dff_A_i518BMWU1_0),.din(w_dff_A_QBNhy4Oo8_0),.clk(gclk));
	jdff dff_A_i518BMWU1_0(.dout(w_dff_A_eGRyYK2v9_0),.din(w_dff_A_i518BMWU1_0),.clk(gclk));
	jdff dff_A_eGRyYK2v9_0(.dout(w_dff_A_RBsEs5yg9_0),.din(w_dff_A_eGRyYK2v9_0),.clk(gclk));
	jdff dff_A_RBsEs5yg9_0(.dout(w_dff_A_gxPcKutd1_0),.din(w_dff_A_RBsEs5yg9_0),.clk(gclk));
	jdff dff_A_gxPcKutd1_0(.dout(w_dff_A_y5PqvIz20_0),.din(w_dff_A_gxPcKutd1_0),.clk(gclk));
	jdff dff_A_y5PqvIz20_0(.dout(w_dff_A_ZXblgs8T7_0),.din(w_dff_A_y5PqvIz20_0),.clk(gclk));
	jdff dff_A_ZXblgs8T7_0(.dout(w_dff_A_MA85Bv5N4_0),.din(w_dff_A_ZXblgs8T7_0),.clk(gclk));
	jdff dff_A_MA85Bv5N4_0(.dout(w_dff_A_2Bp2y0Eh2_0),.din(w_dff_A_MA85Bv5N4_0),.clk(gclk));
	jdff dff_A_2Bp2y0Eh2_0(.dout(w_dff_A_pNyLUNaN5_0),.din(w_dff_A_2Bp2y0Eh2_0),.clk(gclk));
	jdff dff_A_pNyLUNaN5_0(.dout(w_dff_A_ifPUox836_0),.din(w_dff_A_pNyLUNaN5_0),.clk(gclk));
	jdff dff_A_ifPUox836_0(.dout(w_dff_A_Vl8klQJT9_0),.din(w_dff_A_ifPUox836_0),.clk(gclk));
	jdff dff_A_Vl8klQJT9_0(.dout(w_dff_A_PjwROmtr7_0),.din(w_dff_A_Vl8klQJT9_0),.clk(gclk));
	jdff dff_A_PjwROmtr7_0(.dout(w_dff_A_5jvpmlY93_0),.din(w_dff_A_PjwROmtr7_0),.clk(gclk));
	jdff dff_A_5jvpmlY93_0(.dout(w_dff_A_2zTuU5tl4_0),.din(w_dff_A_5jvpmlY93_0),.clk(gclk));
	jdff dff_A_2zTuU5tl4_0(.dout(G4591gat),.din(w_dff_A_2zTuU5tl4_0),.clk(gclk));
	jdff dff_A_TjdGLRLw9_2(.dout(w_dff_A_a6dW4Wnh8_0),.din(w_dff_A_TjdGLRLw9_2),.clk(gclk));
	jdff dff_A_a6dW4Wnh8_0(.dout(w_dff_A_NpRxMuo52_0),.din(w_dff_A_a6dW4Wnh8_0),.clk(gclk));
	jdff dff_A_NpRxMuo52_0(.dout(w_dff_A_c6flYkow7_0),.din(w_dff_A_NpRxMuo52_0),.clk(gclk));
	jdff dff_A_c6flYkow7_0(.dout(w_dff_A_sCc4a96U6_0),.din(w_dff_A_c6flYkow7_0),.clk(gclk));
	jdff dff_A_sCc4a96U6_0(.dout(w_dff_A_AwwDDlC17_0),.din(w_dff_A_sCc4a96U6_0),.clk(gclk));
	jdff dff_A_AwwDDlC17_0(.dout(w_dff_A_CiHco9fX7_0),.din(w_dff_A_AwwDDlC17_0),.clk(gclk));
	jdff dff_A_CiHco9fX7_0(.dout(w_dff_A_NzwOd8pu2_0),.din(w_dff_A_CiHco9fX7_0),.clk(gclk));
	jdff dff_A_NzwOd8pu2_0(.dout(w_dff_A_Z41jJ2T81_0),.din(w_dff_A_NzwOd8pu2_0),.clk(gclk));
	jdff dff_A_Z41jJ2T81_0(.dout(w_dff_A_wWAq8bYL9_0),.din(w_dff_A_Z41jJ2T81_0),.clk(gclk));
	jdff dff_A_wWAq8bYL9_0(.dout(w_dff_A_1I6dMjJc0_0),.din(w_dff_A_wWAq8bYL9_0),.clk(gclk));
	jdff dff_A_1I6dMjJc0_0(.dout(w_dff_A_jGxsFTrn7_0),.din(w_dff_A_1I6dMjJc0_0),.clk(gclk));
	jdff dff_A_jGxsFTrn7_0(.dout(w_dff_A_y5wssT002_0),.din(w_dff_A_jGxsFTrn7_0),.clk(gclk));
	jdff dff_A_y5wssT002_0(.dout(w_dff_A_vphPzTZF8_0),.din(w_dff_A_y5wssT002_0),.clk(gclk));
	jdff dff_A_vphPzTZF8_0(.dout(w_dff_A_Dg5TWWQc3_0),.din(w_dff_A_vphPzTZF8_0),.clk(gclk));
	jdff dff_A_Dg5TWWQc3_0(.dout(w_dff_A_Hjs7E3516_0),.din(w_dff_A_Dg5TWWQc3_0),.clk(gclk));
	jdff dff_A_Hjs7E3516_0(.dout(w_dff_A_r2bio3nM9_0),.din(w_dff_A_Hjs7E3516_0),.clk(gclk));
	jdff dff_A_r2bio3nM9_0(.dout(w_dff_A_FL9yVWlF8_0),.din(w_dff_A_r2bio3nM9_0),.clk(gclk));
	jdff dff_A_FL9yVWlF8_0(.dout(w_dff_A_8R3uGzBw0_0),.din(w_dff_A_FL9yVWlF8_0),.clk(gclk));
	jdff dff_A_8R3uGzBw0_0(.dout(w_dff_A_tk7jAMRt0_0),.din(w_dff_A_8R3uGzBw0_0),.clk(gclk));
	jdff dff_A_tk7jAMRt0_0(.dout(w_dff_A_ADSz6GLN9_0),.din(w_dff_A_tk7jAMRt0_0),.clk(gclk));
	jdff dff_A_ADSz6GLN9_0(.dout(w_dff_A_e6UcSutJ9_0),.din(w_dff_A_ADSz6GLN9_0),.clk(gclk));
	jdff dff_A_e6UcSutJ9_0(.dout(w_dff_A_SQ0a9nQC3_0),.din(w_dff_A_e6UcSutJ9_0),.clk(gclk));
	jdff dff_A_SQ0a9nQC3_0(.dout(w_dff_A_9nhDXwj06_0),.din(w_dff_A_SQ0a9nQC3_0),.clk(gclk));
	jdff dff_A_9nhDXwj06_0(.dout(w_dff_A_Md4bjF6Z9_0),.din(w_dff_A_9nhDXwj06_0),.clk(gclk));
	jdff dff_A_Md4bjF6Z9_0(.dout(w_dff_A_yMqzClJm9_0),.din(w_dff_A_Md4bjF6Z9_0),.clk(gclk));
	jdff dff_A_yMqzClJm9_0(.dout(w_dff_A_P2YcLkYv7_0),.din(w_dff_A_yMqzClJm9_0),.clk(gclk));
	jdff dff_A_P2YcLkYv7_0(.dout(w_dff_A_wDcNvaE75_0),.din(w_dff_A_P2YcLkYv7_0),.clk(gclk));
	jdff dff_A_wDcNvaE75_0(.dout(w_dff_A_zEjC8w5T5_0),.din(w_dff_A_wDcNvaE75_0),.clk(gclk));
	jdff dff_A_zEjC8w5T5_0(.dout(w_dff_A_9NlEIUAy3_0),.din(w_dff_A_zEjC8w5T5_0),.clk(gclk));
	jdff dff_A_9NlEIUAy3_0(.dout(w_dff_A_SxsaFq6y8_0),.din(w_dff_A_9NlEIUAy3_0),.clk(gclk));
	jdff dff_A_SxsaFq6y8_0(.dout(w_dff_A_Bp11NYbI2_0),.din(w_dff_A_SxsaFq6y8_0),.clk(gclk));
	jdff dff_A_Bp11NYbI2_0(.dout(w_dff_A_1KgPX6CE6_0),.din(w_dff_A_Bp11NYbI2_0),.clk(gclk));
	jdff dff_A_1KgPX6CE6_0(.dout(w_dff_A_0ZrandTC4_0),.din(w_dff_A_1KgPX6CE6_0),.clk(gclk));
	jdff dff_A_0ZrandTC4_0(.dout(w_dff_A_7bRrsiQk5_0),.din(w_dff_A_0ZrandTC4_0),.clk(gclk));
	jdff dff_A_7bRrsiQk5_0(.dout(w_dff_A_SJq5fYCH5_0),.din(w_dff_A_7bRrsiQk5_0),.clk(gclk));
	jdff dff_A_SJq5fYCH5_0(.dout(w_dff_A_gvGWBQZQ6_0),.din(w_dff_A_SJq5fYCH5_0),.clk(gclk));
	jdff dff_A_gvGWBQZQ6_0(.dout(w_dff_A_e7Ks6Wl86_0),.din(w_dff_A_gvGWBQZQ6_0),.clk(gclk));
	jdff dff_A_e7Ks6Wl86_0(.dout(w_dff_A_BZDT2QZj6_0),.din(w_dff_A_e7Ks6Wl86_0),.clk(gclk));
	jdff dff_A_BZDT2QZj6_0(.dout(w_dff_A_0UNyN9CL2_0),.din(w_dff_A_BZDT2QZj6_0),.clk(gclk));
	jdff dff_A_0UNyN9CL2_0(.dout(w_dff_A_u4mEd3e62_0),.din(w_dff_A_0UNyN9CL2_0),.clk(gclk));
	jdff dff_A_u4mEd3e62_0(.dout(w_dff_A_p1R9qLD41_0),.din(w_dff_A_u4mEd3e62_0),.clk(gclk));
	jdff dff_A_p1R9qLD41_0(.dout(G4946gat),.din(w_dff_A_p1R9qLD41_0),.clk(gclk));
	jdff dff_A_n39HOqln6_2(.dout(w_dff_A_PXYOGhAB5_0),.din(w_dff_A_n39HOqln6_2),.clk(gclk));
	jdff dff_A_PXYOGhAB5_0(.dout(w_dff_A_ccvQQc4W1_0),.din(w_dff_A_PXYOGhAB5_0),.clk(gclk));
	jdff dff_A_ccvQQc4W1_0(.dout(w_dff_A_v3OSxPsP3_0),.din(w_dff_A_ccvQQc4W1_0),.clk(gclk));
	jdff dff_A_v3OSxPsP3_0(.dout(w_dff_A_KrXAkzbj4_0),.din(w_dff_A_v3OSxPsP3_0),.clk(gclk));
	jdff dff_A_KrXAkzbj4_0(.dout(w_dff_A_QnyWjelI2_0),.din(w_dff_A_KrXAkzbj4_0),.clk(gclk));
	jdff dff_A_QnyWjelI2_0(.dout(w_dff_A_cQwWQltv2_0),.din(w_dff_A_QnyWjelI2_0),.clk(gclk));
	jdff dff_A_cQwWQltv2_0(.dout(w_dff_A_JMQ0IoUh4_0),.din(w_dff_A_cQwWQltv2_0),.clk(gclk));
	jdff dff_A_JMQ0IoUh4_0(.dout(w_dff_A_DGbuDETQ3_0),.din(w_dff_A_JMQ0IoUh4_0),.clk(gclk));
	jdff dff_A_DGbuDETQ3_0(.dout(w_dff_A_MGG4IEfF1_0),.din(w_dff_A_DGbuDETQ3_0),.clk(gclk));
	jdff dff_A_MGG4IEfF1_0(.dout(w_dff_A_KeSUoF4c3_0),.din(w_dff_A_MGG4IEfF1_0),.clk(gclk));
	jdff dff_A_KeSUoF4c3_0(.dout(w_dff_A_XUReLZzE0_0),.din(w_dff_A_KeSUoF4c3_0),.clk(gclk));
	jdff dff_A_XUReLZzE0_0(.dout(w_dff_A_I3tK6U1N1_0),.din(w_dff_A_XUReLZzE0_0),.clk(gclk));
	jdff dff_A_I3tK6U1N1_0(.dout(w_dff_A_GuwBZFwr8_0),.din(w_dff_A_I3tK6U1N1_0),.clk(gclk));
	jdff dff_A_GuwBZFwr8_0(.dout(w_dff_A_9eXdsHEP1_0),.din(w_dff_A_GuwBZFwr8_0),.clk(gclk));
	jdff dff_A_9eXdsHEP1_0(.dout(w_dff_A_UMpSS8Q03_0),.din(w_dff_A_9eXdsHEP1_0),.clk(gclk));
	jdff dff_A_UMpSS8Q03_0(.dout(w_dff_A_Pp0sLBA62_0),.din(w_dff_A_UMpSS8Q03_0),.clk(gclk));
	jdff dff_A_Pp0sLBA62_0(.dout(w_dff_A_skNgviXu7_0),.din(w_dff_A_Pp0sLBA62_0),.clk(gclk));
	jdff dff_A_skNgviXu7_0(.dout(w_dff_A_xTBEM8Fr0_0),.din(w_dff_A_skNgviXu7_0),.clk(gclk));
	jdff dff_A_xTBEM8Fr0_0(.dout(w_dff_A_ysDfatWY2_0),.din(w_dff_A_xTBEM8Fr0_0),.clk(gclk));
	jdff dff_A_ysDfatWY2_0(.dout(w_dff_A_sIBXIBgh7_0),.din(w_dff_A_ysDfatWY2_0),.clk(gclk));
	jdff dff_A_sIBXIBgh7_0(.dout(w_dff_A_D0BStk2N7_0),.din(w_dff_A_sIBXIBgh7_0),.clk(gclk));
	jdff dff_A_D0BStk2N7_0(.dout(w_dff_A_O6fynBIh5_0),.din(w_dff_A_D0BStk2N7_0),.clk(gclk));
	jdff dff_A_O6fynBIh5_0(.dout(w_dff_A_ZrEvEVVm9_0),.din(w_dff_A_O6fynBIh5_0),.clk(gclk));
	jdff dff_A_ZrEvEVVm9_0(.dout(w_dff_A_KrVUD9wZ5_0),.din(w_dff_A_ZrEvEVVm9_0),.clk(gclk));
	jdff dff_A_KrVUD9wZ5_0(.dout(w_dff_A_3rmwHDer8_0),.din(w_dff_A_KrVUD9wZ5_0),.clk(gclk));
	jdff dff_A_3rmwHDer8_0(.dout(w_dff_A_ZM4Q09M85_0),.din(w_dff_A_3rmwHDer8_0),.clk(gclk));
	jdff dff_A_ZM4Q09M85_0(.dout(w_dff_A_RLjrw6mG7_0),.din(w_dff_A_ZM4Q09M85_0),.clk(gclk));
	jdff dff_A_RLjrw6mG7_0(.dout(w_dff_A_7viF9eR54_0),.din(w_dff_A_RLjrw6mG7_0),.clk(gclk));
	jdff dff_A_7viF9eR54_0(.dout(w_dff_A_dQrwwRV21_0),.din(w_dff_A_7viF9eR54_0),.clk(gclk));
	jdff dff_A_dQrwwRV21_0(.dout(w_dff_A_Oc7eU37c1_0),.din(w_dff_A_dQrwwRV21_0),.clk(gclk));
	jdff dff_A_Oc7eU37c1_0(.dout(w_dff_A_TjjslqyG7_0),.din(w_dff_A_Oc7eU37c1_0),.clk(gclk));
	jdff dff_A_TjjslqyG7_0(.dout(w_dff_A_s4eG32rq3_0),.din(w_dff_A_TjjslqyG7_0),.clk(gclk));
	jdff dff_A_s4eG32rq3_0(.dout(w_dff_A_tgEVvcUC2_0),.din(w_dff_A_s4eG32rq3_0),.clk(gclk));
	jdff dff_A_tgEVvcUC2_0(.dout(w_dff_A_TojyohDe3_0),.din(w_dff_A_tgEVvcUC2_0),.clk(gclk));
	jdff dff_A_TojyohDe3_0(.dout(w_dff_A_bjCIdwKR9_0),.din(w_dff_A_TojyohDe3_0),.clk(gclk));
	jdff dff_A_bjCIdwKR9_0(.dout(w_dff_A_XPmKIEMU6_0),.din(w_dff_A_bjCIdwKR9_0),.clk(gclk));
	jdff dff_A_XPmKIEMU6_0(.dout(w_dff_A_eEbg3W3c2_0),.din(w_dff_A_XPmKIEMU6_0),.clk(gclk));
	jdff dff_A_eEbg3W3c2_0(.dout(w_dff_A_UmDYDhTC6_0),.din(w_dff_A_eEbg3W3c2_0),.clk(gclk));
	jdff dff_A_UmDYDhTC6_0(.dout(G5308gat),.din(w_dff_A_UmDYDhTC6_0),.clk(gclk));
	jdff dff_A_WSl0EIyE8_2(.dout(w_dff_A_xitS8AkT0_0),.din(w_dff_A_WSl0EIyE8_2),.clk(gclk));
	jdff dff_A_xitS8AkT0_0(.dout(w_dff_A_BSxvz88n7_0),.din(w_dff_A_xitS8AkT0_0),.clk(gclk));
	jdff dff_A_BSxvz88n7_0(.dout(w_dff_A_LSoJSI6f1_0),.din(w_dff_A_BSxvz88n7_0),.clk(gclk));
	jdff dff_A_LSoJSI6f1_0(.dout(w_dff_A_DGL0CW8y4_0),.din(w_dff_A_LSoJSI6f1_0),.clk(gclk));
	jdff dff_A_DGL0CW8y4_0(.dout(w_dff_A_oTDyi2rv0_0),.din(w_dff_A_DGL0CW8y4_0),.clk(gclk));
	jdff dff_A_oTDyi2rv0_0(.dout(w_dff_A_Y4euN9vd1_0),.din(w_dff_A_oTDyi2rv0_0),.clk(gclk));
	jdff dff_A_Y4euN9vd1_0(.dout(w_dff_A_INVqkSpx5_0),.din(w_dff_A_Y4euN9vd1_0),.clk(gclk));
	jdff dff_A_INVqkSpx5_0(.dout(w_dff_A_f2eq9Zt65_0),.din(w_dff_A_INVqkSpx5_0),.clk(gclk));
	jdff dff_A_f2eq9Zt65_0(.dout(w_dff_A_lqJ6VHIA4_0),.din(w_dff_A_f2eq9Zt65_0),.clk(gclk));
	jdff dff_A_lqJ6VHIA4_0(.dout(w_dff_A_a7SqyRw98_0),.din(w_dff_A_lqJ6VHIA4_0),.clk(gclk));
	jdff dff_A_a7SqyRw98_0(.dout(w_dff_A_N0SmX26K4_0),.din(w_dff_A_a7SqyRw98_0),.clk(gclk));
	jdff dff_A_N0SmX26K4_0(.dout(w_dff_A_BVmziCF87_0),.din(w_dff_A_N0SmX26K4_0),.clk(gclk));
	jdff dff_A_BVmziCF87_0(.dout(w_dff_A_wRb2ybTo8_0),.din(w_dff_A_BVmziCF87_0),.clk(gclk));
	jdff dff_A_wRb2ybTo8_0(.dout(w_dff_A_HBEf2gIx4_0),.din(w_dff_A_wRb2ybTo8_0),.clk(gclk));
	jdff dff_A_HBEf2gIx4_0(.dout(w_dff_A_x3jQrAfc2_0),.din(w_dff_A_HBEf2gIx4_0),.clk(gclk));
	jdff dff_A_x3jQrAfc2_0(.dout(w_dff_A_RYrsZBUM6_0),.din(w_dff_A_x3jQrAfc2_0),.clk(gclk));
	jdff dff_A_RYrsZBUM6_0(.dout(w_dff_A_qKJwP7Kc2_0),.din(w_dff_A_RYrsZBUM6_0),.clk(gclk));
	jdff dff_A_qKJwP7Kc2_0(.dout(w_dff_A_OrKjtW3x1_0),.din(w_dff_A_qKJwP7Kc2_0),.clk(gclk));
	jdff dff_A_OrKjtW3x1_0(.dout(w_dff_A_A9mUCM720_0),.din(w_dff_A_OrKjtW3x1_0),.clk(gclk));
	jdff dff_A_A9mUCM720_0(.dout(w_dff_A_QmJ8Ul4Y6_0),.din(w_dff_A_A9mUCM720_0),.clk(gclk));
	jdff dff_A_QmJ8Ul4Y6_0(.dout(w_dff_A_T9F5kV4w5_0),.din(w_dff_A_QmJ8Ul4Y6_0),.clk(gclk));
	jdff dff_A_T9F5kV4w5_0(.dout(w_dff_A_4aa6IcZh6_0),.din(w_dff_A_T9F5kV4w5_0),.clk(gclk));
	jdff dff_A_4aa6IcZh6_0(.dout(w_dff_A_86YsFzoF3_0),.din(w_dff_A_4aa6IcZh6_0),.clk(gclk));
	jdff dff_A_86YsFzoF3_0(.dout(w_dff_A_RvU0rqpO0_0),.din(w_dff_A_86YsFzoF3_0),.clk(gclk));
	jdff dff_A_RvU0rqpO0_0(.dout(w_dff_A_zREhpBw31_0),.din(w_dff_A_RvU0rqpO0_0),.clk(gclk));
	jdff dff_A_zREhpBw31_0(.dout(w_dff_A_7yGCrpIi9_0),.din(w_dff_A_zREhpBw31_0),.clk(gclk));
	jdff dff_A_7yGCrpIi9_0(.dout(w_dff_A_L3I894qR8_0),.din(w_dff_A_7yGCrpIi9_0),.clk(gclk));
	jdff dff_A_L3I894qR8_0(.dout(w_dff_A_6FNDU8F08_0),.din(w_dff_A_L3I894qR8_0),.clk(gclk));
	jdff dff_A_6FNDU8F08_0(.dout(w_dff_A_JZbZCbVK2_0),.din(w_dff_A_6FNDU8F08_0),.clk(gclk));
	jdff dff_A_JZbZCbVK2_0(.dout(w_dff_A_lZbtv4Dn2_0),.din(w_dff_A_JZbZCbVK2_0),.clk(gclk));
	jdff dff_A_lZbtv4Dn2_0(.dout(w_dff_A_xjQqyAC48_0),.din(w_dff_A_lZbtv4Dn2_0),.clk(gclk));
	jdff dff_A_xjQqyAC48_0(.dout(w_dff_A_NXVTaOIn1_0),.din(w_dff_A_xjQqyAC48_0),.clk(gclk));
	jdff dff_A_NXVTaOIn1_0(.dout(w_dff_A_Arr6ZWbq3_0),.din(w_dff_A_NXVTaOIn1_0),.clk(gclk));
	jdff dff_A_Arr6ZWbq3_0(.dout(w_dff_A_UEa5lEg98_0),.din(w_dff_A_Arr6ZWbq3_0),.clk(gclk));
	jdff dff_A_UEa5lEg98_0(.dout(w_dff_A_AgN3q7uf2_0),.din(w_dff_A_UEa5lEg98_0),.clk(gclk));
	jdff dff_A_AgN3q7uf2_0(.dout(G5672gat),.din(w_dff_A_AgN3q7uf2_0),.clk(gclk));
	jdff dff_A_ZhxLR9C13_2(.dout(w_dff_A_9WX7sZQQ7_0),.din(w_dff_A_ZhxLR9C13_2),.clk(gclk));
	jdff dff_A_9WX7sZQQ7_0(.dout(w_dff_A_Ba3QuFnW3_0),.din(w_dff_A_9WX7sZQQ7_0),.clk(gclk));
	jdff dff_A_Ba3QuFnW3_0(.dout(w_dff_A_kWVBo9Cp2_0),.din(w_dff_A_Ba3QuFnW3_0),.clk(gclk));
	jdff dff_A_kWVBo9Cp2_0(.dout(w_dff_A_lqVv0DfJ7_0),.din(w_dff_A_kWVBo9Cp2_0),.clk(gclk));
	jdff dff_A_lqVv0DfJ7_0(.dout(w_dff_A_ZeDiL4Ar9_0),.din(w_dff_A_lqVv0DfJ7_0),.clk(gclk));
	jdff dff_A_ZeDiL4Ar9_0(.dout(w_dff_A_JMvNQLNs0_0),.din(w_dff_A_ZeDiL4Ar9_0),.clk(gclk));
	jdff dff_A_JMvNQLNs0_0(.dout(w_dff_A_MzjB351A9_0),.din(w_dff_A_JMvNQLNs0_0),.clk(gclk));
	jdff dff_A_MzjB351A9_0(.dout(w_dff_A_CpuYyrwR5_0),.din(w_dff_A_MzjB351A9_0),.clk(gclk));
	jdff dff_A_CpuYyrwR5_0(.dout(w_dff_A_v7UpYvVh4_0),.din(w_dff_A_CpuYyrwR5_0),.clk(gclk));
	jdff dff_A_v7UpYvVh4_0(.dout(w_dff_A_YOXKoh117_0),.din(w_dff_A_v7UpYvVh4_0),.clk(gclk));
	jdff dff_A_YOXKoh117_0(.dout(w_dff_A_C6uF63eD0_0),.din(w_dff_A_YOXKoh117_0),.clk(gclk));
	jdff dff_A_C6uF63eD0_0(.dout(w_dff_A_wvJpvDsk0_0),.din(w_dff_A_C6uF63eD0_0),.clk(gclk));
	jdff dff_A_wvJpvDsk0_0(.dout(w_dff_A_dwkQyt1l6_0),.din(w_dff_A_wvJpvDsk0_0),.clk(gclk));
	jdff dff_A_dwkQyt1l6_0(.dout(w_dff_A_StsFwRK94_0),.din(w_dff_A_dwkQyt1l6_0),.clk(gclk));
	jdff dff_A_StsFwRK94_0(.dout(w_dff_A_njdFfX3w3_0),.din(w_dff_A_StsFwRK94_0),.clk(gclk));
	jdff dff_A_njdFfX3w3_0(.dout(w_dff_A_Ozixgr5S6_0),.din(w_dff_A_njdFfX3w3_0),.clk(gclk));
	jdff dff_A_Ozixgr5S6_0(.dout(w_dff_A_nG3rHP5V2_0),.din(w_dff_A_Ozixgr5S6_0),.clk(gclk));
	jdff dff_A_nG3rHP5V2_0(.dout(w_dff_A_ZJdGLJYx9_0),.din(w_dff_A_nG3rHP5V2_0),.clk(gclk));
	jdff dff_A_ZJdGLJYx9_0(.dout(w_dff_A_clh1lQBc8_0),.din(w_dff_A_ZJdGLJYx9_0),.clk(gclk));
	jdff dff_A_clh1lQBc8_0(.dout(w_dff_A_B1DojI7m5_0),.din(w_dff_A_clh1lQBc8_0),.clk(gclk));
	jdff dff_A_B1DojI7m5_0(.dout(w_dff_A_zOwrnuid2_0),.din(w_dff_A_B1DojI7m5_0),.clk(gclk));
	jdff dff_A_zOwrnuid2_0(.dout(w_dff_A_TRer6PZN2_0),.din(w_dff_A_zOwrnuid2_0),.clk(gclk));
	jdff dff_A_TRer6PZN2_0(.dout(w_dff_A_F5ym6srX2_0),.din(w_dff_A_TRer6PZN2_0),.clk(gclk));
	jdff dff_A_F5ym6srX2_0(.dout(w_dff_A_SxJqZXzi3_0),.din(w_dff_A_F5ym6srX2_0),.clk(gclk));
	jdff dff_A_SxJqZXzi3_0(.dout(w_dff_A_hmBfOyWc5_0),.din(w_dff_A_SxJqZXzi3_0),.clk(gclk));
	jdff dff_A_hmBfOyWc5_0(.dout(w_dff_A_xIqKHLJc8_0),.din(w_dff_A_hmBfOyWc5_0),.clk(gclk));
	jdff dff_A_xIqKHLJc8_0(.dout(w_dff_A_EAKZ0q5X5_0),.din(w_dff_A_xIqKHLJc8_0),.clk(gclk));
	jdff dff_A_EAKZ0q5X5_0(.dout(w_dff_A_Rc7ncFnQ7_0),.din(w_dff_A_EAKZ0q5X5_0),.clk(gclk));
	jdff dff_A_Rc7ncFnQ7_0(.dout(w_dff_A_qJOfDy521_0),.din(w_dff_A_Rc7ncFnQ7_0),.clk(gclk));
	jdff dff_A_qJOfDy521_0(.dout(w_dff_A_pzyh0SBC4_0),.din(w_dff_A_qJOfDy521_0),.clk(gclk));
	jdff dff_A_pzyh0SBC4_0(.dout(w_dff_A_XtjlzGCk4_0),.din(w_dff_A_pzyh0SBC4_0),.clk(gclk));
	jdff dff_A_XtjlzGCk4_0(.dout(w_dff_A_32zRcKXp9_0),.din(w_dff_A_XtjlzGCk4_0),.clk(gclk));
	jdff dff_A_32zRcKXp9_0(.dout(G5971gat),.din(w_dff_A_32zRcKXp9_0),.clk(gclk));
	jdff dff_A_RiGNgq0v5_2(.dout(w_dff_A_BRaODm1z6_0),.din(w_dff_A_RiGNgq0v5_2),.clk(gclk));
	jdff dff_A_BRaODm1z6_0(.dout(w_dff_A_y6YdgwjN3_0),.din(w_dff_A_BRaODm1z6_0),.clk(gclk));
	jdff dff_A_y6YdgwjN3_0(.dout(w_dff_A_sA3CfVXX8_0),.din(w_dff_A_y6YdgwjN3_0),.clk(gclk));
	jdff dff_A_sA3CfVXX8_0(.dout(w_dff_A_nMnbmvvI1_0),.din(w_dff_A_sA3CfVXX8_0),.clk(gclk));
	jdff dff_A_nMnbmvvI1_0(.dout(w_dff_A_sQlvJgaY8_0),.din(w_dff_A_nMnbmvvI1_0),.clk(gclk));
	jdff dff_A_sQlvJgaY8_0(.dout(w_dff_A_uoPjVtxN1_0),.din(w_dff_A_sQlvJgaY8_0),.clk(gclk));
	jdff dff_A_uoPjVtxN1_0(.dout(w_dff_A_7yrMR0ab4_0),.din(w_dff_A_uoPjVtxN1_0),.clk(gclk));
	jdff dff_A_7yrMR0ab4_0(.dout(w_dff_A_VTEG6IL61_0),.din(w_dff_A_7yrMR0ab4_0),.clk(gclk));
	jdff dff_A_VTEG6IL61_0(.dout(w_dff_A_4Uxi5dxr4_0),.din(w_dff_A_VTEG6IL61_0),.clk(gclk));
	jdff dff_A_4Uxi5dxr4_0(.dout(w_dff_A_YeTiCmJM6_0),.din(w_dff_A_4Uxi5dxr4_0),.clk(gclk));
	jdff dff_A_YeTiCmJM6_0(.dout(w_dff_A_XEOHnWHI5_0),.din(w_dff_A_YeTiCmJM6_0),.clk(gclk));
	jdff dff_A_XEOHnWHI5_0(.dout(w_dff_A_mYFAKh8B8_0),.din(w_dff_A_XEOHnWHI5_0),.clk(gclk));
	jdff dff_A_mYFAKh8B8_0(.dout(w_dff_A_2Rl10XbI4_0),.din(w_dff_A_mYFAKh8B8_0),.clk(gclk));
	jdff dff_A_2Rl10XbI4_0(.dout(w_dff_A_8PSniu2M8_0),.din(w_dff_A_2Rl10XbI4_0),.clk(gclk));
	jdff dff_A_8PSniu2M8_0(.dout(w_dff_A_WvLuzetH5_0),.din(w_dff_A_8PSniu2M8_0),.clk(gclk));
	jdff dff_A_WvLuzetH5_0(.dout(w_dff_A_7rhpeM8U9_0),.din(w_dff_A_WvLuzetH5_0),.clk(gclk));
	jdff dff_A_7rhpeM8U9_0(.dout(w_dff_A_H6GXloK48_0),.din(w_dff_A_7rhpeM8U9_0),.clk(gclk));
	jdff dff_A_H6GXloK48_0(.dout(w_dff_A_m2SXRMYS6_0),.din(w_dff_A_H6GXloK48_0),.clk(gclk));
	jdff dff_A_m2SXRMYS6_0(.dout(w_dff_A_dP2cDpOZ9_0),.din(w_dff_A_m2SXRMYS6_0),.clk(gclk));
	jdff dff_A_dP2cDpOZ9_0(.dout(w_dff_A_Ziz6r9ml4_0),.din(w_dff_A_dP2cDpOZ9_0),.clk(gclk));
	jdff dff_A_Ziz6r9ml4_0(.dout(w_dff_A_f8EEHrxG9_0),.din(w_dff_A_Ziz6r9ml4_0),.clk(gclk));
	jdff dff_A_f8EEHrxG9_0(.dout(w_dff_A_IoTughCQ0_0),.din(w_dff_A_f8EEHrxG9_0),.clk(gclk));
	jdff dff_A_IoTughCQ0_0(.dout(w_dff_A_akKqVMdM8_0),.din(w_dff_A_IoTughCQ0_0),.clk(gclk));
	jdff dff_A_akKqVMdM8_0(.dout(w_dff_A_pMCnnbfu9_0),.din(w_dff_A_akKqVMdM8_0),.clk(gclk));
	jdff dff_A_pMCnnbfu9_0(.dout(w_dff_A_CWhxHb8s9_0),.din(w_dff_A_pMCnnbfu9_0),.clk(gclk));
	jdff dff_A_CWhxHb8s9_0(.dout(w_dff_A_i6BPHUvn5_0),.din(w_dff_A_CWhxHb8s9_0),.clk(gclk));
	jdff dff_A_i6BPHUvn5_0(.dout(w_dff_A_B2W53vBp3_0),.din(w_dff_A_i6BPHUvn5_0),.clk(gclk));
	jdff dff_A_B2W53vBp3_0(.dout(w_dff_A_AjyUEPaL0_0),.din(w_dff_A_B2W53vBp3_0),.clk(gclk));
	jdff dff_A_AjyUEPaL0_0(.dout(w_dff_A_4BgyMPAM4_0),.din(w_dff_A_AjyUEPaL0_0),.clk(gclk));
	jdff dff_A_4BgyMPAM4_0(.dout(G6123gat),.din(w_dff_A_4BgyMPAM4_0),.clk(gclk));
	jdff dff_A_YCRvBVIi5_2(.dout(w_dff_A_HhMXcIse2_0),.din(w_dff_A_YCRvBVIi5_2),.clk(gclk));
	jdff dff_A_HhMXcIse2_0(.dout(w_dff_A_k2PgIPBi0_0),.din(w_dff_A_HhMXcIse2_0),.clk(gclk));
	jdff dff_A_k2PgIPBi0_0(.dout(w_dff_A_wJHW178i5_0),.din(w_dff_A_k2PgIPBi0_0),.clk(gclk));
	jdff dff_A_wJHW178i5_0(.dout(w_dff_A_KtLN4ZB32_0),.din(w_dff_A_wJHW178i5_0),.clk(gclk));
	jdff dff_A_KtLN4ZB32_0(.dout(w_dff_A_3ikgKnXR2_0),.din(w_dff_A_KtLN4ZB32_0),.clk(gclk));
	jdff dff_A_3ikgKnXR2_0(.dout(w_dff_A_UyHNsjUb8_0),.din(w_dff_A_3ikgKnXR2_0),.clk(gclk));
	jdff dff_A_UyHNsjUb8_0(.dout(w_dff_A_7S8vQGny7_0),.din(w_dff_A_UyHNsjUb8_0),.clk(gclk));
	jdff dff_A_7S8vQGny7_0(.dout(w_dff_A_uqCEpxMI5_0),.din(w_dff_A_7S8vQGny7_0),.clk(gclk));
	jdff dff_A_uqCEpxMI5_0(.dout(w_dff_A_Tlcq6KGg6_0),.din(w_dff_A_uqCEpxMI5_0),.clk(gclk));
	jdff dff_A_Tlcq6KGg6_0(.dout(w_dff_A_vKU23z184_0),.din(w_dff_A_Tlcq6KGg6_0),.clk(gclk));
	jdff dff_A_vKU23z184_0(.dout(w_dff_A_IgztpfZa8_0),.din(w_dff_A_vKU23z184_0),.clk(gclk));
	jdff dff_A_IgztpfZa8_0(.dout(w_dff_A_uoBjILui7_0),.din(w_dff_A_IgztpfZa8_0),.clk(gclk));
	jdff dff_A_uoBjILui7_0(.dout(w_dff_A_Cb9Hg85J4_0),.din(w_dff_A_uoBjILui7_0),.clk(gclk));
	jdff dff_A_Cb9Hg85J4_0(.dout(w_dff_A_6akwj2CO0_0),.din(w_dff_A_Cb9Hg85J4_0),.clk(gclk));
	jdff dff_A_6akwj2CO0_0(.dout(w_dff_A_bS45ZKch5_0),.din(w_dff_A_6akwj2CO0_0),.clk(gclk));
	jdff dff_A_bS45ZKch5_0(.dout(w_dff_A_5dZKLWRO0_0),.din(w_dff_A_bS45ZKch5_0),.clk(gclk));
	jdff dff_A_5dZKLWRO0_0(.dout(w_dff_A_3e9fCXZc2_0),.din(w_dff_A_5dZKLWRO0_0),.clk(gclk));
	jdff dff_A_3e9fCXZc2_0(.dout(w_dff_A_EH0zUNSa3_0),.din(w_dff_A_3e9fCXZc2_0),.clk(gclk));
	jdff dff_A_EH0zUNSa3_0(.dout(w_dff_A_jsneHnAm8_0),.din(w_dff_A_EH0zUNSa3_0),.clk(gclk));
	jdff dff_A_jsneHnAm8_0(.dout(w_dff_A_sjZouKhD0_0),.din(w_dff_A_jsneHnAm8_0),.clk(gclk));
	jdff dff_A_sjZouKhD0_0(.dout(w_dff_A_4cBQzAk47_0),.din(w_dff_A_sjZouKhD0_0),.clk(gclk));
	jdff dff_A_4cBQzAk47_0(.dout(w_dff_A_9HaDc8zY5_0),.din(w_dff_A_4cBQzAk47_0),.clk(gclk));
	jdff dff_A_9HaDc8zY5_0(.dout(w_dff_A_EQhHENGU5_0),.din(w_dff_A_9HaDc8zY5_0),.clk(gclk));
	jdff dff_A_EQhHENGU5_0(.dout(w_dff_A_cHkLUQnw4_0),.din(w_dff_A_EQhHENGU5_0),.clk(gclk));
	jdff dff_A_cHkLUQnw4_0(.dout(w_dff_A_4hAR9USW3_0),.din(w_dff_A_cHkLUQnw4_0),.clk(gclk));
	jdff dff_A_4hAR9USW3_0(.dout(w_dff_A_ZJWPtwWd1_0),.din(w_dff_A_4hAR9USW3_0),.clk(gclk));
	jdff dff_A_ZJWPtwWd1_0(.dout(w_dff_A_cO1UaNWW3_0),.din(w_dff_A_ZJWPtwWd1_0),.clk(gclk));
	jdff dff_A_cO1UaNWW3_0(.dout(G6150gat),.din(w_dff_A_cO1UaNWW3_0),.clk(gclk));
	jdff dff_A_3j1PEYfK3_2(.dout(w_dff_A_sO9qh7Ax4_0),.din(w_dff_A_3j1PEYfK3_2),.clk(gclk));
	jdff dff_A_sO9qh7Ax4_0(.dout(w_dff_A_GhHGmgVn7_0),.din(w_dff_A_sO9qh7Ax4_0),.clk(gclk));
	jdff dff_A_GhHGmgVn7_0(.dout(w_dff_A_BrBtDBV98_0),.din(w_dff_A_GhHGmgVn7_0),.clk(gclk));
	jdff dff_A_BrBtDBV98_0(.dout(w_dff_A_j3J5GqAj0_0),.din(w_dff_A_BrBtDBV98_0),.clk(gclk));
	jdff dff_A_j3J5GqAj0_0(.dout(w_dff_A_av1uvVys2_0),.din(w_dff_A_j3J5GqAj0_0),.clk(gclk));
	jdff dff_A_av1uvVys2_0(.dout(w_dff_A_XaX95qps8_0),.din(w_dff_A_av1uvVys2_0),.clk(gclk));
	jdff dff_A_XaX95qps8_0(.dout(w_dff_A_mktdfFWU4_0),.din(w_dff_A_XaX95qps8_0),.clk(gclk));
	jdff dff_A_mktdfFWU4_0(.dout(w_dff_A_kr2eQAx83_0),.din(w_dff_A_mktdfFWU4_0),.clk(gclk));
	jdff dff_A_kr2eQAx83_0(.dout(w_dff_A_BLsqHu6k6_0),.din(w_dff_A_kr2eQAx83_0),.clk(gclk));
	jdff dff_A_BLsqHu6k6_0(.dout(w_dff_A_c6yqcFoO5_0),.din(w_dff_A_BLsqHu6k6_0),.clk(gclk));
	jdff dff_A_c6yqcFoO5_0(.dout(w_dff_A_khXknZXq3_0),.din(w_dff_A_c6yqcFoO5_0),.clk(gclk));
	jdff dff_A_khXknZXq3_0(.dout(w_dff_A_DEbtyCtf3_0),.din(w_dff_A_khXknZXq3_0),.clk(gclk));
	jdff dff_A_DEbtyCtf3_0(.dout(w_dff_A_h7t1cluU1_0),.din(w_dff_A_DEbtyCtf3_0),.clk(gclk));
	jdff dff_A_h7t1cluU1_0(.dout(w_dff_A_jPpR8efA0_0),.din(w_dff_A_h7t1cluU1_0),.clk(gclk));
	jdff dff_A_jPpR8efA0_0(.dout(w_dff_A_rFk65SJ82_0),.din(w_dff_A_jPpR8efA0_0),.clk(gclk));
	jdff dff_A_rFk65SJ82_0(.dout(w_dff_A_wjJBQDJX9_0),.din(w_dff_A_rFk65SJ82_0),.clk(gclk));
	jdff dff_A_wjJBQDJX9_0(.dout(w_dff_A_25khai6V3_0),.din(w_dff_A_wjJBQDJX9_0),.clk(gclk));
	jdff dff_A_25khai6V3_0(.dout(w_dff_A_kQdSDMHx2_0),.din(w_dff_A_25khai6V3_0),.clk(gclk));
	jdff dff_A_kQdSDMHx2_0(.dout(w_dff_A_TKnrswjf5_0),.din(w_dff_A_kQdSDMHx2_0),.clk(gclk));
	jdff dff_A_TKnrswjf5_0(.dout(w_dff_A_k0T0mM0J9_0),.din(w_dff_A_TKnrswjf5_0),.clk(gclk));
	jdff dff_A_k0T0mM0J9_0(.dout(w_dff_A_3ltsmNx67_0),.din(w_dff_A_k0T0mM0J9_0),.clk(gclk));
	jdff dff_A_3ltsmNx67_0(.dout(w_dff_A_Z9Ci4EUj9_0),.din(w_dff_A_3ltsmNx67_0),.clk(gclk));
	jdff dff_A_Z9Ci4EUj9_0(.dout(w_dff_A_SBKcqrin0_0),.din(w_dff_A_Z9Ci4EUj9_0),.clk(gclk));
	jdff dff_A_SBKcqrin0_0(.dout(w_dff_A_tfMGGzxj6_0),.din(w_dff_A_SBKcqrin0_0),.clk(gclk));
	jdff dff_A_tfMGGzxj6_0(.dout(w_dff_A_Se8Tumc06_0),.din(w_dff_A_tfMGGzxj6_0),.clk(gclk));
	jdff dff_A_Se8Tumc06_0(.dout(G6160gat),.din(w_dff_A_Se8Tumc06_0),.clk(gclk));
	jdff dff_A_qleo09kn4_2(.dout(w_dff_A_lCBBv9QO2_0),.din(w_dff_A_qleo09kn4_2),.clk(gclk));
	jdff dff_A_lCBBv9QO2_0(.dout(w_dff_A_TtyIYZh40_0),.din(w_dff_A_lCBBv9QO2_0),.clk(gclk));
	jdff dff_A_TtyIYZh40_0(.dout(w_dff_A_RfM33e8G2_0),.din(w_dff_A_TtyIYZh40_0),.clk(gclk));
	jdff dff_A_RfM33e8G2_0(.dout(w_dff_A_LWO1MQ7j5_0),.din(w_dff_A_RfM33e8G2_0),.clk(gclk));
	jdff dff_A_LWO1MQ7j5_0(.dout(w_dff_A_VlMxCanH3_0),.din(w_dff_A_LWO1MQ7j5_0),.clk(gclk));
	jdff dff_A_VlMxCanH3_0(.dout(w_dff_A_s1UldOVh1_0),.din(w_dff_A_VlMxCanH3_0),.clk(gclk));
	jdff dff_A_s1UldOVh1_0(.dout(w_dff_A_7EA0wUEj3_0),.din(w_dff_A_s1UldOVh1_0),.clk(gclk));
	jdff dff_A_7EA0wUEj3_0(.dout(w_dff_A_XRwueToC5_0),.din(w_dff_A_7EA0wUEj3_0),.clk(gclk));
	jdff dff_A_XRwueToC5_0(.dout(w_dff_A_87h3UxEH1_0),.din(w_dff_A_XRwueToC5_0),.clk(gclk));
	jdff dff_A_87h3UxEH1_0(.dout(w_dff_A_WtGHggMp3_0),.din(w_dff_A_87h3UxEH1_0),.clk(gclk));
	jdff dff_A_WtGHggMp3_0(.dout(w_dff_A_6GAAc6RP9_0),.din(w_dff_A_WtGHggMp3_0),.clk(gclk));
	jdff dff_A_6GAAc6RP9_0(.dout(w_dff_A_NlVlxsS29_0),.din(w_dff_A_6GAAc6RP9_0),.clk(gclk));
	jdff dff_A_NlVlxsS29_0(.dout(w_dff_A_qEFfAEZq2_0),.din(w_dff_A_NlVlxsS29_0),.clk(gclk));
	jdff dff_A_qEFfAEZq2_0(.dout(w_dff_A_KAjV3HxG2_0),.din(w_dff_A_qEFfAEZq2_0),.clk(gclk));
	jdff dff_A_KAjV3HxG2_0(.dout(w_dff_A_zhSAuQKB4_0),.din(w_dff_A_KAjV3HxG2_0),.clk(gclk));
	jdff dff_A_zhSAuQKB4_0(.dout(w_dff_A_4lAkaNN30_0),.din(w_dff_A_zhSAuQKB4_0),.clk(gclk));
	jdff dff_A_4lAkaNN30_0(.dout(w_dff_A_mHHFsiDr7_0),.din(w_dff_A_4lAkaNN30_0),.clk(gclk));
	jdff dff_A_mHHFsiDr7_0(.dout(w_dff_A_JCOnup5O1_0),.din(w_dff_A_mHHFsiDr7_0),.clk(gclk));
	jdff dff_A_JCOnup5O1_0(.dout(w_dff_A_EScLjh3c1_0),.din(w_dff_A_JCOnup5O1_0),.clk(gclk));
	jdff dff_A_EScLjh3c1_0(.dout(w_dff_A_KK68eYoc4_0),.din(w_dff_A_EScLjh3c1_0),.clk(gclk));
	jdff dff_A_KK68eYoc4_0(.dout(w_dff_A_A3dIK2xS6_0),.din(w_dff_A_KK68eYoc4_0),.clk(gclk));
	jdff dff_A_A3dIK2xS6_0(.dout(w_dff_A_Adjwx5WL4_0),.din(w_dff_A_A3dIK2xS6_0),.clk(gclk));
	jdff dff_A_Adjwx5WL4_0(.dout(w_dff_A_zdxO5D4b5_0),.din(w_dff_A_Adjwx5WL4_0),.clk(gclk));
	jdff dff_A_zdxO5D4b5_0(.dout(w_dff_A_hsHi8AYr0_0),.din(w_dff_A_zdxO5D4b5_0),.clk(gclk));
	jdff dff_A_hsHi8AYr0_0(.dout(G6170gat),.din(w_dff_A_hsHi8AYr0_0),.clk(gclk));
	jdff dff_A_Mg1X7kYi3_2(.dout(w_dff_A_2qyJRMkA9_0),.din(w_dff_A_Mg1X7kYi3_2),.clk(gclk));
	jdff dff_A_2qyJRMkA9_0(.dout(w_dff_A_BvZPiXOZ1_0),.din(w_dff_A_2qyJRMkA9_0),.clk(gclk));
	jdff dff_A_BvZPiXOZ1_0(.dout(w_dff_A_TvY2d2tY5_0),.din(w_dff_A_BvZPiXOZ1_0),.clk(gclk));
	jdff dff_A_TvY2d2tY5_0(.dout(w_dff_A_7R5GOZxK4_0),.din(w_dff_A_TvY2d2tY5_0),.clk(gclk));
	jdff dff_A_7R5GOZxK4_0(.dout(w_dff_A_ATA3UeNa2_0),.din(w_dff_A_7R5GOZxK4_0),.clk(gclk));
	jdff dff_A_ATA3UeNa2_0(.dout(w_dff_A_NLanNwY27_0),.din(w_dff_A_ATA3UeNa2_0),.clk(gclk));
	jdff dff_A_NLanNwY27_0(.dout(w_dff_A_RfXxmmml3_0),.din(w_dff_A_NLanNwY27_0),.clk(gclk));
	jdff dff_A_RfXxmmml3_0(.dout(w_dff_A_Y6LGIcFt5_0),.din(w_dff_A_RfXxmmml3_0),.clk(gclk));
	jdff dff_A_Y6LGIcFt5_0(.dout(w_dff_A_IHAPyJVP3_0),.din(w_dff_A_Y6LGIcFt5_0),.clk(gclk));
	jdff dff_A_IHAPyJVP3_0(.dout(w_dff_A_dJ6Fhpld1_0),.din(w_dff_A_IHAPyJVP3_0),.clk(gclk));
	jdff dff_A_dJ6Fhpld1_0(.dout(w_dff_A_JHshYPrD9_0),.din(w_dff_A_dJ6Fhpld1_0),.clk(gclk));
	jdff dff_A_JHshYPrD9_0(.dout(w_dff_A_seeCy2Kh2_0),.din(w_dff_A_JHshYPrD9_0),.clk(gclk));
	jdff dff_A_seeCy2Kh2_0(.dout(w_dff_A_nhVTJuWH6_0),.din(w_dff_A_seeCy2Kh2_0),.clk(gclk));
	jdff dff_A_nhVTJuWH6_0(.dout(w_dff_A_H0NHJC9x9_0),.din(w_dff_A_nhVTJuWH6_0),.clk(gclk));
	jdff dff_A_H0NHJC9x9_0(.dout(w_dff_A_A8G9NNRv7_0),.din(w_dff_A_H0NHJC9x9_0),.clk(gclk));
	jdff dff_A_A8G9NNRv7_0(.dout(w_dff_A_FY8nLnZF1_0),.din(w_dff_A_A8G9NNRv7_0),.clk(gclk));
	jdff dff_A_FY8nLnZF1_0(.dout(w_dff_A_WMQTWhBY1_0),.din(w_dff_A_FY8nLnZF1_0),.clk(gclk));
	jdff dff_A_WMQTWhBY1_0(.dout(w_dff_A_76rm7cOk5_0),.din(w_dff_A_WMQTWhBY1_0),.clk(gclk));
	jdff dff_A_76rm7cOk5_0(.dout(w_dff_A_OBMLu1gw6_0),.din(w_dff_A_76rm7cOk5_0),.clk(gclk));
	jdff dff_A_OBMLu1gw6_0(.dout(w_dff_A_botBkKyD1_0),.din(w_dff_A_OBMLu1gw6_0),.clk(gclk));
	jdff dff_A_botBkKyD1_0(.dout(w_dff_A_HxraTx742_0),.din(w_dff_A_botBkKyD1_0),.clk(gclk));
	jdff dff_A_HxraTx742_0(.dout(w_dff_A_iv5Ka1kQ3_0),.din(w_dff_A_HxraTx742_0),.clk(gclk));
	jdff dff_A_iv5Ka1kQ3_0(.dout(G6180gat),.din(w_dff_A_iv5Ka1kQ3_0),.clk(gclk));
	jdff dff_A_CwhZzTZn9_2(.dout(w_dff_A_tbPRJOkG3_0),.din(w_dff_A_CwhZzTZn9_2),.clk(gclk));
	jdff dff_A_tbPRJOkG3_0(.dout(w_dff_A_XslWL3Q60_0),.din(w_dff_A_tbPRJOkG3_0),.clk(gclk));
	jdff dff_A_XslWL3Q60_0(.dout(w_dff_A_p12QtY3W0_0),.din(w_dff_A_XslWL3Q60_0),.clk(gclk));
	jdff dff_A_p12QtY3W0_0(.dout(w_dff_A_GAJ89qqD4_0),.din(w_dff_A_p12QtY3W0_0),.clk(gclk));
	jdff dff_A_GAJ89qqD4_0(.dout(w_dff_A_tZIVaVvy3_0),.din(w_dff_A_GAJ89qqD4_0),.clk(gclk));
	jdff dff_A_tZIVaVvy3_0(.dout(w_dff_A_Rvp6YINZ0_0),.din(w_dff_A_tZIVaVvy3_0),.clk(gclk));
	jdff dff_A_Rvp6YINZ0_0(.dout(w_dff_A_eeohvE6f8_0),.din(w_dff_A_Rvp6YINZ0_0),.clk(gclk));
	jdff dff_A_eeohvE6f8_0(.dout(w_dff_A_pWRahA418_0),.din(w_dff_A_eeohvE6f8_0),.clk(gclk));
	jdff dff_A_pWRahA418_0(.dout(w_dff_A_l0gaW0P47_0),.din(w_dff_A_pWRahA418_0),.clk(gclk));
	jdff dff_A_l0gaW0P47_0(.dout(w_dff_A_GfyRGFpY7_0),.din(w_dff_A_l0gaW0P47_0),.clk(gclk));
	jdff dff_A_GfyRGFpY7_0(.dout(w_dff_A_ekRWmT9K0_0),.din(w_dff_A_GfyRGFpY7_0),.clk(gclk));
	jdff dff_A_ekRWmT9K0_0(.dout(w_dff_A_zo52ntwV2_0),.din(w_dff_A_ekRWmT9K0_0),.clk(gclk));
	jdff dff_A_zo52ntwV2_0(.dout(w_dff_A_jqpPCvAa8_0),.din(w_dff_A_zo52ntwV2_0),.clk(gclk));
	jdff dff_A_jqpPCvAa8_0(.dout(w_dff_A_LftrWyT60_0),.din(w_dff_A_jqpPCvAa8_0),.clk(gclk));
	jdff dff_A_LftrWyT60_0(.dout(w_dff_A_HbxrLCr01_0),.din(w_dff_A_LftrWyT60_0),.clk(gclk));
	jdff dff_A_HbxrLCr01_0(.dout(w_dff_A_LCDLV67j8_0),.din(w_dff_A_HbxrLCr01_0),.clk(gclk));
	jdff dff_A_LCDLV67j8_0(.dout(w_dff_A_SJ9EuBEv5_0),.din(w_dff_A_LCDLV67j8_0),.clk(gclk));
	jdff dff_A_SJ9EuBEv5_0(.dout(w_dff_A_h5UXlaAh7_0),.din(w_dff_A_SJ9EuBEv5_0),.clk(gclk));
	jdff dff_A_h5UXlaAh7_0(.dout(w_dff_A_1sC049pU4_0),.din(w_dff_A_h5UXlaAh7_0),.clk(gclk));
	jdff dff_A_1sC049pU4_0(.dout(w_dff_A_5mAlZ4cm9_0),.din(w_dff_A_1sC049pU4_0),.clk(gclk));
	jdff dff_A_5mAlZ4cm9_0(.dout(G6190gat),.din(w_dff_A_5mAlZ4cm9_0),.clk(gclk));
	jdff dff_A_6Ai86vBq2_2(.dout(w_dff_A_a1VLTSCQ7_0),.din(w_dff_A_6Ai86vBq2_2),.clk(gclk));
	jdff dff_A_a1VLTSCQ7_0(.dout(w_dff_A_IRgXpY0P6_0),.din(w_dff_A_a1VLTSCQ7_0),.clk(gclk));
	jdff dff_A_IRgXpY0P6_0(.dout(w_dff_A_qDronPmb3_0),.din(w_dff_A_IRgXpY0P6_0),.clk(gclk));
	jdff dff_A_qDronPmb3_0(.dout(w_dff_A_FZN0y7y06_0),.din(w_dff_A_qDronPmb3_0),.clk(gclk));
	jdff dff_A_FZN0y7y06_0(.dout(w_dff_A_O4Lpzdwo0_0),.din(w_dff_A_FZN0y7y06_0),.clk(gclk));
	jdff dff_A_O4Lpzdwo0_0(.dout(w_dff_A_XJFN3vim8_0),.din(w_dff_A_O4Lpzdwo0_0),.clk(gclk));
	jdff dff_A_XJFN3vim8_0(.dout(w_dff_A_Q4HwkHwE8_0),.din(w_dff_A_XJFN3vim8_0),.clk(gclk));
	jdff dff_A_Q4HwkHwE8_0(.dout(w_dff_A_w9looatv2_0),.din(w_dff_A_Q4HwkHwE8_0),.clk(gclk));
	jdff dff_A_w9looatv2_0(.dout(w_dff_A_dMMYrJ129_0),.din(w_dff_A_w9looatv2_0),.clk(gclk));
	jdff dff_A_dMMYrJ129_0(.dout(w_dff_A_xJTKLktf7_0),.din(w_dff_A_dMMYrJ129_0),.clk(gclk));
	jdff dff_A_xJTKLktf7_0(.dout(w_dff_A_6wb2kHls0_0),.din(w_dff_A_xJTKLktf7_0),.clk(gclk));
	jdff dff_A_6wb2kHls0_0(.dout(w_dff_A_EEPKoRtu3_0),.din(w_dff_A_6wb2kHls0_0),.clk(gclk));
	jdff dff_A_EEPKoRtu3_0(.dout(w_dff_A_SLmZPEzj6_0),.din(w_dff_A_EEPKoRtu3_0),.clk(gclk));
	jdff dff_A_SLmZPEzj6_0(.dout(w_dff_A_0wp4JsRD2_0),.din(w_dff_A_SLmZPEzj6_0),.clk(gclk));
	jdff dff_A_0wp4JsRD2_0(.dout(w_dff_A_NecOSmkM1_0),.din(w_dff_A_0wp4JsRD2_0),.clk(gclk));
	jdff dff_A_NecOSmkM1_0(.dout(w_dff_A_6a1JAple9_0),.din(w_dff_A_NecOSmkM1_0),.clk(gclk));
	jdff dff_A_6a1JAple9_0(.dout(w_dff_A_GHovIGQH4_0),.din(w_dff_A_6a1JAple9_0),.clk(gclk));
	jdff dff_A_GHovIGQH4_0(.dout(w_dff_A_gprhUM183_0),.din(w_dff_A_GHovIGQH4_0),.clk(gclk));
	jdff dff_A_gprhUM183_0(.dout(G6200gat),.din(w_dff_A_gprhUM183_0),.clk(gclk));
	jdff dff_A_L32hW2LS1_2(.dout(w_dff_A_iBoSeqZ20_0),.din(w_dff_A_L32hW2LS1_2),.clk(gclk));
	jdff dff_A_iBoSeqZ20_0(.dout(w_dff_A_R1ARCxDp7_0),.din(w_dff_A_iBoSeqZ20_0),.clk(gclk));
	jdff dff_A_R1ARCxDp7_0(.dout(w_dff_A_FXDStuyO8_0),.din(w_dff_A_R1ARCxDp7_0),.clk(gclk));
	jdff dff_A_FXDStuyO8_0(.dout(w_dff_A_cYNaAvBj0_0),.din(w_dff_A_FXDStuyO8_0),.clk(gclk));
	jdff dff_A_cYNaAvBj0_0(.dout(w_dff_A_jUExLUyv5_0),.din(w_dff_A_cYNaAvBj0_0),.clk(gclk));
	jdff dff_A_jUExLUyv5_0(.dout(w_dff_A_71jGEFgd5_0),.din(w_dff_A_jUExLUyv5_0),.clk(gclk));
	jdff dff_A_71jGEFgd5_0(.dout(w_dff_A_s4THd8ww1_0),.din(w_dff_A_71jGEFgd5_0),.clk(gclk));
	jdff dff_A_s4THd8ww1_0(.dout(w_dff_A_4PPJga7z6_0),.din(w_dff_A_s4THd8ww1_0),.clk(gclk));
	jdff dff_A_4PPJga7z6_0(.dout(w_dff_A_m6g3Z6dN4_0),.din(w_dff_A_4PPJga7z6_0),.clk(gclk));
	jdff dff_A_m6g3Z6dN4_0(.dout(w_dff_A_Fvialyc24_0),.din(w_dff_A_m6g3Z6dN4_0),.clk(gclk));
	jdff dff_A_Fvialyc24_0(.dout(w_dff_A_S9UxOVWJ3_0),.din(w_dff_A_Fvialyc24_0),.clk(gclk));
	jdff dff_A_S9UxOVWJ3_0(.dout(w_dff_A_XN0ANblW1_0),.din(w_dff_A_S9UxOVWJ3_0),.clk(gclk));
	jdff dff_A_XN0ANblW1_0(.dout(w_dff_A_Vf4sA6Ky9_0),.din(w_dff_A_XN0ANblW1_0),.clk(gclk));
	jdff dff_A_Vf4sA6Ky9_0(.dout(w_dff_A_UqpThG0K5_0),.din(w_dff_A_Vf4sA6Ky9_0),.clk(gclk));
	jdff dff_A_UqpThG0K5_0(.dout(w_dff_A_ID7eH4Lh0_0),.din(w_dff_A_UqpThG0K5_0),.clk(gclk));
	jdff dff_A_ID7eH4Lh0_0(.dout(w_dff_A_q9MdTBve0_0),.din(w_dff_A_ID7eH4Lh0_0),.clk(gclk));
	jdff dff_A_q9MdTBve0_0(.dout(G6210gat),.din(w_dff_A_q9MdTBve0_0),.clk(gclk));
	jdff dff_A_U4vuyFKf9_2(.dout(w_dff_A_1EfTJIz48_0),.din(w_dff_A_U4vuyFKf9_2),.clk(gclk));
	jdff dff_A_1EfTJIz48_0(.dout(w_dff_A_ZD3ppNsg2_0),.din(w_dff_A_1EfTJIz48_0),.clk(gclk));
	jdff dff_A_ZD3ppNsg2_0(.dout(w_dff_A_dqws9YBK7_0),.din(w_dff_A_ZD3ppNsg2_0),.clk(gclk));
	jdff dff_A_dqws9YBK7_0(.dout(w_dff_A_hUuoMGJp2_0),.din(w_dff_A_dqws9YBK7_0),.clk(gclk));
	jdff dff_A_hUuoMGJp2_0(.dout(w_dff_A_9fFbRT7h1_0),.din(w_dff_A_hUuoMGJp2_0),.clk(gclk));
	jdff dff_A_9fFbRT7h1_0(.dout(w_dff_A_3EUl0YvF1_0),.din(w_dff_A_9fFbRT7h1_0),.clk(gclk));
	jdff dff_A_3EUl0YvF1_0(.dout(w_dff_A_HoHzlm9f1_0),.din(w_dff_A_3EUl0YvF1_0),.clk(gclk));
	jdff dff_A_HoHzlm9f1_0(.dout(w_dff_A_8WCLFQ7O6_0),.din(w_dff_A_HoHzlm9f1_0),.clk(gclk));
	jdff dff_A_8WCLFQ7O6_0(.dout(w_dff_A_tdvirqIT9_0),.din(w_dff_A_8WCLFQ7O6_0),.clk(gclk));
	jdff dff_A_tdvirqIT9_0(.dout(w_dff_A_ll3i0FjZ5_0),.din(w_dff_A_tdvirqIT9_0),.clk(gclk));
	jdff dff_A_ll3i0FjZ5_0(.dout(w_dff_A_EE7XoC5N7_0),.din(w_dff_A_ll3i0FjZ5_0),.clk(gclk));
	jdff dff_A_EE7XoC5N7_0(.dout(w_dff_A_rsW6fxGB1_0),.din(w_dff_A_EE7XoC5N7_0),.clk(gclk));
	jdff dff_A_rsW6fxGB1_0(.dout(w_dff_A_gYBEpimB0_0),.din(w_dff_A_rsW6fxGB1_0),.clk(gclk));
	jdff dff_A_gYBEpimB0_0(.dout(w_dff_A_0f26mPQq5_0),.din(w_dff_A_gYBEpimB0_0),.clk(gclk));
	jdff dff_A_0f26mPQq5_0(.dout(G6220gat),.din(w_dff_A_0f26mPQq5_0),.clk(gclk));
	jdff dff_A_nROzBrc79_2(.dout(w_dff_A_1vMYkrXz2_0),.din(w_dff_A_nROzBrc79_2),.clk(gclk));
	jdff dff_A_1vMYkrXz2_0(.dout(w_dff_A_XcRWpCha5_0),.din(w_dff_A_1vMYkrXz2_0),.clk(gclk));
	jdff dff_A_XcRWpCha5_0(.dout(w_dff_A_y2jtvMmp1_0),.din(w_dff_A_XcRWpCha5_0),.clk(gclk));
	jdff dff_A_y2jtvMmp1_0(.dout(w_dff_A_D9PLMhrS7_0),.din(w_dff_A_y2jtvMmp1_0),.clk(gclk));
	jdff dff_A_D9PLMhrS7_0(.dout(w_dff_A_O7AZxJAF0_0),.din(w_dff_A_D9PLMhrS7_0),.clk(gclk));
	jdff dff_A_O7AZxJAF0_0(.dout(w_dff_A_JpOTPatm4_0),.din(w_dff_A_O7AZxJAF0_0),.clk(gclk));
	jdff dff_A_JpOTPatm4_0(.dout(w_dff_A_U3alkdkB6_0),.din(w_dff_A_JpOTPatm4_0),.clk(gclk));
	jdff dff_A_U3alkdkB6_0(.dout(w_dff_A_aBjB7jI41_0),.din(w_dff_A_U3alkdkB6_0),.clk(gclk));
	jdff dff_A_aBjB7jI41_0(.dout(w_dff_A_SaEu00Pt2_0),.din(w_dff_A_aBjB7jI41_0),.clk(gclk));
	jdff dff_A_SaEu00Pt2_0(.dout(w_dff_A_DZtfkPET7_0),.din(w_dff_A_SaEu00Pt2_0),.clk(gclk));
	jdff dff_A_DZtfkPET7_0(.dout(w_dff_A_Lj47b4v46_0),.din(w_dff_A_DZtfkPET7_0),.clk(gclk));
	jdff dff_A_Lj47b4v46_0(.dout(w_dff_A_rjdUdsfB2_0),.din(w_dff_A_Lj47b4v46_0),.clk(gclk));
	jdff dff_A_rjdUdsfB2_0(.dout(G6230gat),.din(w_dff_A_rjdUdsfB2_0),.clk(gclk));
	jdff dff_A_Hct20z8J2_2(.dout(w_dff_A_2UwWnLJQ9_0),.din(w_dff_A_Hct20z8J2_2),.clk(gclk));
	jdff dff_A_2UwWnLJQ9_0(.dout(w_dff_A_35PE9aVP0_0),.din(w_dff_A_2UwWnLJQ9_0),.clk(gclk));
	jdff dff_A_35PE9aVP0_0(.dout(w_dff_A_rlxzxRmH2_0),.din(w_dff_A_35PE9aVP0_0),.clk(gclk));
	jdff dff_A_rlxzxRmH2_0(.dout(w_dff_A_kRC3yNG81_0),.din(w_dff_A_rlxzxRmH2_0),.clk(gclk));
	jdff dff_A_kRC3yNG81_0(.dout(w_dff_A_ikuaTzLq8_0),.din(w_dff_A_kRC3yNG81_0),.clk(gclk));
	jdff dff_A_ikuaTzLq8_0(.dout(w_dff_A_Nu0umgT08_0),.din(w_dff_A_ikuaTzLq8_0),.clk(gclk));
	jdff dff_A_Nu0umgT08_0(.dout(w_dff_A_9Vrmr2321_0),.din(w_dff_A_Nu0umgT08_0),.clk(gclk));
	jdff dff_A_9Vrmr2321_0(.dout(w_dff_A_NjidA3oc1_0),.din(w_dff_A_9Vrmr2321_0),.clk(gclk));
	jdff dff_A_NjidA3oc1_0(.dout(w_dff_A_1mrt8IqO9_0),.din(w_dff_A_NjidA3oc1_0),.clk(gclk));
	jdff dff_A_1mrt8IqO9_0(.dout(w_dff_A_alY01VwI7_0),.din(w_dff_A_1mrt8IqO9_0),.clk(gclk));
	jdff dff_A_alY01VwI7_0(.dout(G6240gat),.din(w_dff_A_alY01VwI7_0),.clk(gclk));
	jdff dff_A_48KSIqDl5_2(.dout(w_dff_A_asVgSdPS4_0),.din(w_dff_A_48KSIqDl5_2),.clk(gclk));
	jdff dff_A_asVgSdPS4_0(.dout(w_dff_A_o8KvXOaC8_0),.din(w_dff_A_asVgSdPS4_0),.clk(gclk));
	jdff dff_A_o8KvXOaC8_0(.dout(w_dff_A_mVAHhzcV7_0),.din(w_dff_A_o8KvXOaC8_0),.clk(gclk));
	jdff dff_A_mVAHhzcV7_0(.dout(w_dff_A_0WIRGioh0_0),.din(w_dff_A_mVAHhzcV7_0),.clk(gclk));
	jdff dff_A_0WIRGioh0_0(.dout(w_dff_A_Xnt55Kve0_0),.din(w_dff_A_0WIRGioh0_0),.clk(gclk));
	jdff dff_A_Xnt55Kve0_0(.dout(w_dff_A_ig11lh6X4_0),.din(w_dff_A_Xnt55Kve0_0),.clk(gclk));
	jdff dff_A_ig11lh6X4_0(.dout(w_dff_A_YU1PYqp05_0),.din(w_dff_A_ig11lh6X4_0),.clk(gclk));
	jdff dff_A_YU1PYqp05_0(.dout(w_dff_A_pJpFmTC08_0),.din(w_dff_A_YU1PYqp05_0),.clk(gclk));
	jdff dff_A_pJpFmTC08_0(.dout(G6250gat),.din(w_dff_A_pJpFmTC08_0),.clk(gclk));
	jdff dff_A_uIbrthHL5_2(.dout(w_dff_A_nvLQ7oa05_0),.din(w_dff_A_uIbrthHL5_2),.clk(gclk));
	jdff dff_A_nvLQ7oa05_0(.dout(w_dff_A_qEEUoxZz6_0),.din(w_dff_A_nvLQ7oa05_0),.clk(gclk));
	jdff dff_A_qEEUoxZz6_0(.dout(w_dff_A_e706UnFA6_0),.din(w_dff_A_qEEUoxZz6_0),.clk(gclk));
	jdff dff_A_e706UnFA6_0(.dout(w_dff_A_Wcb4ODzY8_0),.din(w_dff_A_e706UnFA6_0),.clk(gclk));
	jdff dff_A_Wcb4ODzY8_0(.dout(w_dff_A_UOVXcXQh8_0),.din(w_dff_A_Wcb4ODzY8_0),.clk(gclk));
	jdff dff_A_UOVXcXQh8_0(.dout(w_dff_A_XgkLyMkz7_0),.din(w_dff_A_UOVXcXQh8_0),.clk(gclk));
	jdff dff_A_XgkLyMkz7_0(.dout(G6260gat),.din(w_dff_A_XgkLyMkz7_0),.clk(gclk));
	jdff dff_A_UUSXDR6i6_2(.dout(w_dff_A_uBwifqyv9_0),.din(w_dff_A_UUSXDR6i6_2),.clk(gclk));
	jdff dff_A_uBwifqyv9_0(.dout(w_dff_A_oQ1DY9T72_0),.din(w_dff_A_uBwifqyv9_0),.clk(gclk));
	jdff dff_A_oQ1DY9T72_0(.dout(w_dff_A_IQ7iIc6H0_0),.din(w_dff_A_oQ1DY9T72_0),.clk(gclk));
	jdff dff_A_IQ7iIc6H0_0(.dout(w_dff_A_BKciDslk4_0),.din(w_dff_A_IQ7iIc6H0_0),.clk(gclk));
	jdff dff_A_BKciDslk4_0(.dout(G6270gat),.din(w_dff_A_BKciDslk4_0),.clk(gclk));
	jdff dff_A_zwUMdALK2_2(.dout(w_dff_A_xozSZBXo9_0),.din(w_dff_A_zwUMdALK2_2),.clk(gclk));
	jdff dff_A_xozSZBXo9_0(.dout(w_dff_A_odSiYtK84_0),.din(w_dff_A_xozSZBXo9_0),.clk(gclk));
	jdff dff_A_odSiYtK84_0(.dout(G6280gat),.din(w_dff_A_odSiYtK84_0),.clk(gclk));
	jdff dff_A_KQCoHiXA8_2(.dout(G6288gat),.din(w_dff_A_KQCoHiXA8_2),.clk(gclk));
endmodule

