/*

c880:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jdff: 1127
	jand: 153
	jor: 119

Summary:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jdff: 1127
	jand: 153
	jor: 119
*/

module c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n101;
	wire n102;
	wire n103;
	wire n105;
	wire n106;
	wire n107;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n118;
	wire n119;
	wire n121;
	wire n122;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire [2:0] w_G1gat_0;
	wire [1:0] w_G1gat_1;
	wire [1:0] w_G8gat_0;
	wire [1:0] w_G13gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G17gat_1;
	wire [2:0] w_G17gat_2;
	wire [1:0] w_G26gat_0;
	wire [2:0] w_G29gat_0;
	wire [1:0] w_G36gat_0;
	wire [2:0] w_G42gat_0;
	wire [2:0] w_G42gat_1;
	wire [1:0] w_G42gat_2;
	wire [2:0] w_G51gat_0;
	wire [1:0] w_G51gat_1;
	wire [2:0] w_G55gat_0;
	wire [2:0] w_G59gat_0;
	wire [1:0] w_G59gat_1;
	wire [1:0] w_G68gat_0;
	wire [1:0] w_G75gat_0;
	wire [2:0] w_G80gat_0;
	wire [2:0] w_G91gat_0;
	wire [2:0] w_G96gat_0;
	wire [2:0] w_G101gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G111gat_0;
	wire [2:0] w_G116gat_0;
	wire [2:0] w_G121gat_0;
	wire [1:0] w_G126gat_0;
	wire [1:0] w_G130gat_0;
	wire [2:0] w_G138gat_0;
	wire [1:0] w_G138gat_1;
	wire [1:0] w_G143gat_0;
	wire [1:0] w_G146gat_0;
	wire [1:0] w_G149gat_0;
	wire [2:0] w_G153gat_0;
	wire [1:0] w_G156gat_0;
	wire [2:0] w_G159gat_0;
	wire [2:0] w_G159gat_1;
	wire [1:0] w_G159gat_2;
	wire [2:0] w_G165gat_0;
	wire [2:0] w_G165gat_1;
	wire [1:0] w_G165gat_2;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [1:0] w_G171gat_2;
	wire [2:0] w_G177gat_0;
	wire [2:0] w_G177gat_1;
	wire [1:0] w_G177gat_2;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G183gat_1;
	wire [1:0] w_G183gat_2;
	wire [2:0] w_G189gat_0;
	wire [2:0] w_G189gat_1;
	wire [1:0] w_G189gat_2;
	wire [2:0] w_G195gat_0;
	wire [2:0] w_G195gat_1;
	wire [1:0] w_G195gat_2;
	wire [2:0] w_G201gat_0;
	wire [2:0] w_G201gat_1;
	wire [2:0] w_G201gat_2;
	wire [2:0] w_G210gat_0;
	wire [2:0] w_G210gat_1;
	wire [2:0] w_G210gat_2;
	wire [1:0] w_G210gat_3;
	wire [2:0] w_G219gat_0;
	wire [2:0] w_G219gat_1;
	wire [2:0] w_G219gat_2;
	wire [1:0] w_G219gat_3;
	wire [2:0] w_G228gat_0;
	wire [2:0] w_G228gat_1;
	wire [2:0] w_G228gat_2;
	wire [1:0] w_G228gat_3;
	wire [2:0] w_G237gat_0;
	wire [2:0] w_G237gat_1;
	wire [2:0] w_G237gat_2;
	wire [1:0] w_G237gat_3;
	wire [2:0] w_G246gat_0;
	wire [2:0] w_G246gat_1;
	wire [2:0] w_G246gat_2;
	wire [1:0] w_G246gat_3;
	wire [2:0] w_G255gat_0;
	wire [2:0] w_G261gat_0;
	wire [1:0] w_G268gat_0;
	wire [1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire [2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire [1:0] w_n86_0;
	wire [1:0] w_n88_0;
	wire [2:0] w_n92_0;
	wire [1:0] w_n93_0;
	wire [1:0] w_n96_0;
	wire [1:0] w_n98_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n102_0;
	wire [1:0] w_n106_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n111_0;
	wire [2:0] w_n118_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n143_0;
	wire [1:0] w_n149_0;
	wire [2:0] w_n153_0;
	wire [2:0] w_n153_1;
	wire [2:0] w_n153_2;
	wire [1:0] w_n153_3;
	wire [1:0] w_n154_0;
	wire [1:0] w_n157_0;
	wire [2:0] w_n159_0;
	wire [1:0] w_n159_1;
	wire [1:0] w_n162_0;
	wire [1:0] w_n163_0;
	wire [2:0] w_n165_0;
	wire [2:0] w_n165_1;
	wire [2:0] w_n167_0;
	wire [1:0] w_n167_1;
	wire [2:0] w_n168_0;
	wire [2:0] w_n181_0;
	wire [2:0] w_n181_1;
	wire [2:0] w_n181_2;
	wire [1:0] w_n181_3;
	wire [2:0] w_n193_0;
	wire [1:0] w_n193_1;
	wire [2:0] w_n194_0;
	wire [1:0] w_n196_0;
	wire [1:0] w_n213_0;
	wire [2:0] w_n217_0;
	wire [1:0] w_n217_1;
	wire [1:0] w_n218_0;
	wire [2:0] w_n222_0;
	wire [1:0] w_n222_1;
	wire [1:0] w_n223_0;
	wire [1:0] w_n224_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n230_0;
	wire [1:0] w_n232_0;
	wire [2:0] w_n236_0;
	wire [1:0] w_n238_0;
	wire [2:0] w_n252_0;
	wire [1:0] w_n255_0;
	wire [2:0] w_n273_0;
	wire [2:0] w_n292_0;
	wire [1:0] w_n292_1;
	wire [2:0] w_n296_0;
	wire [1:0] w_n296_1;
	wire [2:0] w_n299_0;
	wire [1:0] w_n299_1;
	wire [1:0] w_n302_0;
	wire [1:0] w_n303_0;
	wire [2:0] w_n305_0;
	wire [1:0] w_n305_1;
	wire [2:0] w_n312_0;
	wire [1:0] w_n312_1;
	wire [1:0] w_n315_0;
	wire [2:0] w_n321_0;
	wire [1:0] w_n321_1;
	wire [1:0] w_n322_0;
	wire [2:0] w_n328_0;
	wire [1:0] w_n328_1;
	wire [2:0] w_n329_0;
	wire [2:0] w_n330_0;
	wire [1:0] w_n331_0;
	wire [2:0] w_n335_0;
	wire [2:0] w_n337_0;
	wire [1:0] w_n339_0;
	wire [1:0] w_n340_0;
	wire [2:0] w_n346_0;
	wire [1:0] w_n346_1;
	wire [2:0] w_n347_0;
	wire [2:0] w_n367_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n405_0;
	wire w_dff_B_BU45obMx4_2;
	wire w_dff_B_22qa2mCN4_1;
	wire w_dff_B_ZJ08p9kY6_1;
	wire w_dff_A_5uYtbCG08_1;
	wire w_dff_B_ceDN2Djk0_0;
	wire w_dff_B_HgsG02sy0_1;
	wire w_dff_B_JnfuJnBI7_1;
	wire w_dff_B_DkYoUwob4_0;
	wire w_dff_B_66ClkBp46_1;
	wire w_dff_B_d7QAY0mr7_0;
	wire w_dff_B_mlTGZ9UB3_0;
	wire w_dff_B_iUY5G3Q84_1;
	wire w_dff_B_d9aQ3Hsl2_0;
	wire w_dff_B_978t756o8_2;
	wire w_dff_B_eKCnf7nW4_0;
	wire w_dff_B_23MZzeTv0_0;
	wire w_dff_B_pPDGf0V36_0;
	wire w_dff_B_wuapAiYt0_0;
	wire w_dff_B_ylPBW2Nm7_0;
	wire w_dff_B_35T3dBtB9_0;
	wire w_dff_B_g769SKK74_0;
	wire w_dff_B_AVY1b9U14_0;
	wire w_dff_B_uM2M20Dq5_0;
	wire w_dff_B_5aExwmzQ1_0;
	wire w_dff_B_MnkDCOT22_0;
	wire w_dff_B_D401LXRg8_0;
	wire w_dff_B_df9p8KhU5_0;
	wire w_dff_A_wvNXrZLk3_1;
	wire w_dff_A_a7Hqmr399_1;
	wire w_dff_A_HA6vdDli5_1;
	wire w_dff_A_Eocuhlud6_1;
	wire w_dff_A_thWiTtzF7_1;
	wire w_dff_A_smmUMEVX2_1;
	wire w_dff_A_MD05oMil1_1;
	wire w_dff_A_AN8Xwk1H3_1;
	wire w_dff_B_A0jSQbd32_0;
	wire w_dff_B_ZelMu73y6_0;
	wire w_dff_B_khC0ug2t3_0;
	wire w_dff_B_DjfMI7uu4_0;
	wire w_dff_B_MFvsdWBy7_0;
	wire w_dff_B_5Bjpjaiq3_0;
	wire w_dff_B_VZlolp058_0;
	wire w_dff_B_zwv9qhOX5_0;
	wire w_dff_B_K5lGTDEM3_0;
	wire w_dff_B_53uxGn3G2_0;
	wire w_dff_B_YW3Yrrpb5_0;
	wire w_dff_B_gR5RYfHF0_0;
	wire w_dff_B_eBN9lLZU9_0;
	wire w_dff_B_8Q4QnE9a2_0;
	wire w_dff_B_yUhUZWtt3_0;
	wire w_dff_B_ydxMKmUe2_0;
	wire w_dff_B_EvIZxbTB2_0;
	wire w_dff_B_MxYrP5QC5_0;
	wire w_dff_A_dtsjmMvx8_0;
	wire w_dff_A_tlWR1w6w5_0;
	wire w_dff_A_53eI4pQg0_0;
	wire w_dff_A_EJDOXZUE8_0;
	wire w_dff_B_NAQTZAus9_1;
	wire w_dff_B_HmJUGg7H5_1;
	wire w_dff_B_vrgnYpuX7_1;
	wire w_dff_B_J7uiEXF66_1;
	wire w_dff_A_Mh1l4sjP7_1;
	wire w_dff_A_SkIorOFb3_1;
	wire w_dff_A_BGzuIdcz9_1;
	wire w_dff_A_mVPNFlTl0_1;
	wire w_dff_A_mqtz29nv3_0;
	wire w_dff_A_JVSnyORT2_0;
	wire w_dff_A_1JKA2zIv4_0;
	wire w_dff_A_oOzkPEPs5_0;
	wire w_dff_A_El0hZZmp6_0;
	wire w_dff_A_tiZ38Rkz4_0;
	wire w_dff_A_72Ud20aI9_0;
	wire w_dff_A_yvRtKMeT2_0;
	wire w_dff_B_ho6uvlZN0_0;
	wire w_dff_B_I6hY2S6W7_0;
	wire w_dff_B_tnQsj0tV8_0;
	wire w_dff_B_XHSx1ZBu3_0;
	wire w_dff_B_ZKSjb0ht7_0;
	wire w_dff_B_wfrQhoPj6_0;
	wire w_dff_B_nzPYfjuJ0_0;
	wire w_dff_B_IfB1r0h09_0;
	wire w_dff_B_hlTtz6bQ7_0;
	wire w_dff_B_Beu8LTgM6_0;
	wire w_dff_B_gKnj4rBG1_0;
	wire w_dff_B_Hk1vbXn17_0;
	wire w_dff_B_p4axHPQU7_0;
	wire w_dff_B_0JCT6MEU5_0;
	wire w_dff_B_BHnfWOY67_0;
	wire w_dff_B_r9j17qxj2_0;
	wire w_dff_B_iKCGrPsq2_0;
	wire w_dff_B_9PG3ojBh5_1;
	wire w_dff_B_Js87Eamr8_1;
	wire w_dff_B_QtNeyt9Z9_1;
	wire w_dff_B_C5AC7Cip1_1;
	wire w_dff_A_sTJD3KC79_1;
	wire w_dff_A_KIfhSZCt4_1;
	wire w_dff_A_Cp6SfsxI7_1;
	wire w_dff_A_IySSeJOx0_1;
	wire w_dff_B_Kcj0PMBs5_0;
	wire w_dff_B_RS7rAgY10_0;
	wire w_dff_B_KbnTInxV4_0;
	wire w_dff_B_3hReHb1S3_0;
	wire w_dff_B_7Ro2bqcZ9_0;
	wire w_dff_B_sDU7CWKL3_0;
	wire w_dff_B_MEe6xGvZ3_0;
	wire w_dff_B_39uTlUH40_0;
	wire w_dff_B_ccXQruad6_0;
	wire w_dff_B_4vc40hgv7_0;
	wire w_dff_B_L4UgJcEY6_0;
	wire w_dff_B_Rn4toji56_0;
	wire w_dff_B_JF5mahsl5_0;
	wire w_dff_B_01hQ1cwc4_0;
	wire w_dff_B_hIcihech9_0;
	wire w_dff_B_xsxlOgxW3_0;
	wire w_dff_B_eUvIE2o32_0;
	wire w_dff_A_T4dEj9Ob6_1;
	wire w_dff_A_DizNzasm0_1;
	wire w_dff_B_3YdSgdhR7_1;
	wire w_dff_B_LWTMNUNt7_1;
	wire w_dff_B_IIetBZfP8_1;
	wire w_dff_B_V9V0yxRE2_1;
	wire w_dff_B_AnPgj2KF8_1;
	wire w_dff_B_u8fZuA1f0_1;
	wire w_dff_B_83ceRUQp2_1;
	wire w_dff_B_tgHPkVDP5_1;
	wire w_dff_B_pzyD4PB77_1;
	wire w_dff_B_drA7A5wC2_1;
	wire w_dff_B_yykAJLWp3_1;
	wire w_dff_B_8izQVtUh2_1;
	wire w_dff_B_KDxHs3hd5_1;
	wire w_dff_B_DnY8NSN65_1;
	wire w_dff_B_NFWHi29h8_1;
	wire w_dff_B_dYeNWM4I5_1;
	wire w_dff_B_Dq2S9tTl5_1;
	wire w_dff_B_GFIofgPe5_1;
	wire w_dff_B_9x4JXOZc9_1;
	wire w_dff_A_1VeCIsG01_0;
	wire w_dff_A_6l3YBqOA0_0;
	wire w_dff_A_OUxX7aTZ4_0;
	wire w_dff_A_HMxZArqn0_0;
	wire w_dff_A_ueE7Fqvm8_0;
	wire w_dff_A_6NhCLcMG5_0;
	wire w_dff_A_T5wby41Q7_0;
	wire w_dff_B_NohDFIkr6_0;
	wire w_dff_B_g2q1NrVl8_0;
	wire w_dff_B_HupO2SMB8_0;
	wire w_dff_B_Awq6aRL81_0;
	wire w_dff_B_PS80H6pj5_0;
	wire w_dff_B_2jCX0utf5_0;
	wire w_dff_B_SHvCg2vu0_0;
	wire w_dff_B_ZvgTSLK49_0;
	wire w_dff_B_3cwJJFb74_0;
	wire w_dff_B_lE9VLwQq3_0;
	wire w_dff_B_dIKLuiks4_0;
	wire w_dff_B_PT4MfKwO1_0;
	wire w_dff_B_TuSVCqe91_0;
	wire w_dff_B_1iohtdfD7_0;
	wire w_dff_B_dEiiDR826_0;
	wire w_dff_B_eHewIdvm5_0;
	wire w_dff_B_dyuU603b1_0;
	wire w_dff_B_4S9IAbVG3_0;
	wire w_dff_B_58zR0n3s1_0;
	wire w_dff_A_iFem6Mhk9_1;
	wire w_dff_A_1u7JjUPF2_2;
	wire w_dff_A_iy772LK66_0;
	wire w_dff_A_RjFmsIgn2_0;
	wire w_dff_A_AHRPNo1Y6_0;
	wire w_dff_A_10DzDZaA4_0;
	wire w_dff_A_57hrO2Mz8_2;
	wire w_dff_A_qRXtUuAr5_2;
	wire w_dff_B_n7vBmzCc0_0;
	wire w_dff_B_W6AUlIsY8_0;
	wire w_dff_B_REeXiNpg3_0;
	wire w_dff_B_tdBjlrPr4_0;
	wire w_dff_B_MRBmsPZg6_0;
	wire w_dff_B_DduR3R5e2_0;
	wire w_dff_B_44poXEwj6_0;
	wire w_dff_A_023pSUSL8_1;
	wire w_dff_A_mQ522mJ64_1;
	wire w_dff_A_uWHcZJfe4_1;
	wire w_dff_A_wEDMyrs09_1;
	wire w_dff_A_mzoGyn4B0_1;
	wire w_dff_A_0u0C7DSN1_1;
	wire w_dff_A_382X31nZ2_1;
	wire w_dff_B_RbdGLSY84_0;
	wire w_dff_B_DCjs5pew3_0;
	wire w_dff_B_Qh2DSA8C9_0;
	wire w_dff_B_8MAWAhCN2_0;
	wire w_dff_B_3HOLFLU23_0;
	wire w_dff_B_UdIWA2le0_0;
	wire w_dff_B_K8L4snng6_0;
	wire w_dff_B_SV1T3fdX5_0;
	wire w_dff_B_6y7RmwYH6_0;
	wire w_dff_B_hfzIin7F9_0;
	wire w_dff_B_XsB5ta5w8_0;
	wire w_dff_B_HzuYTE3n4_0;
	wire w_dff_B_lGaIPzou0_0;
	wire w_dff_B_oxWpBES39_0;
	wire w_dff_B_O4iooApG8_0;
	wire w_dff_B_Ez5N4pDZ5_0;
	wire w_dff_B_BOETqyeV1_0;
	wire w_dff_B_CNQ7J28V6_0;
	wire w_dff_B_7kxTMH5k9_0;
	wire w_dff_B_Ypk3RyhC7_0;
	wire w_dff_B_Htl8yZ1Z7_0;
	wire w_dff_B_vlvA8ewb1_0;
	wire w_dff_B_PVg1L6ik6_0;
	wire w_dff_B_K9MJvytw5_0;
	wire w_dff_B_0vlXdP8K4_0;
	wire w_dff_B_jzB7yExU8_0;
	wire w_dff_B_iQYmiAqk8_0;
	wire w_dff_B_QxNk1A3N2_0;
	wire w_dff_B_UMThZjei6_0;
	wire w_dff_B_sABVbcuN3_0;
	wire w_dff_A_qMR68vi01_1;
	wire w_dff_A_moYjWur72_1;
	wire w_dff_A_zKQ21zr36_1;
	wire w_dff_A_sY73Bu0e0_1;
	wire w_dff_A_4bTtr4l67_1;
	wire w_dff_A_7YyEK7lJ1_1;
	wire w_dff_A_P6LhuJ0q7_1;
	wire w_dff_A_7lI4wPMX7_1;
	wire w_dff_A_kV4L7Rfy6_1;
	wire w_dff_B_CpyIbm2t2_1;
	wire w_dff_B_f4GQoigI6_1;
	wire w_dff_B_zCnyp4Y35_1;
	wire w_dff_A_nky78gyn8_1;
	wire w_dff_A_VyvMVabj5_1;
	wire w_dff_A_dZWcCDWf5_1;
	wire w_dff_A_oVl6N6Q58_1;
	wire w_dff_A_MLQumjyQ5_1;
	wire w_dff_A_TjKz3ELb1_1;
	wire w_dff_A_b8BjMrtc1_1;
	wire w_dff_A_4FtGxaiL4_2;
	wire w_dff_A_md4OBqlg8_2;
	wire w_dff_A_wHAWheAa9_2;
	wire w_dff_A_8yc16Ims3_2;
	wire w_dff_A_eulngWVQ4_2;
	wire w_dff_A_XILNzLwa2_2;
	wire w_dff_A_IeRBU1Vr6_2;
	wire w_dff_A_1K3pnApX4_2;
	wire w_dff_A_QYGY4fAK9_2;
	wire w_dff_A_JOkXOb1G4_2;
	wire w_dff_A_eE0L9O3I9_2;
	wire w_dff_B_E7Vdx2XL5_0;
	wire w_dff_B_qtI8Krpp6_0;
	wire w_dff_B_sn8D4Nq37_0;
	wire w_dff_B_qWOZGGdK5_0;
	wire w_dff_A_J7C3tMNX3_1;
	wire w_dff_A_HH4gkS7P9_1;
	wire w_dff_A_uUGfd9rD4_1;
	wire w_dff_A_bPtpMy9K0_1;
	wire w_dff_B_OzhusPhr2_1;
	wire w_dff_B_gVWJZjbU0_1;
	wire w_dff_B_53ySjMjh9_1;
	wire w_dff_B_FM5y4UtP8_0;
	wire w_dff_B_JILSaziY6_0;
	wire w_dff_B_JWZSHydl1_0;
	wire w_dff_B_mmHNanG33_0;
	wire w_dff_A_OH6QxyuU1_1;
	wire w_dff_A_q1zVOeYm6_1;
	wire w_dff_A_8PprXWsr3_1;
	wire w_dff_A_pWXqXzVN4_1;
	wire w_dff_B_KvBNEMRH7_1;
	wire w_dff_B_5Mqvhx6I2_1;
	wire w_dff_B_PRPPknrU4_1;
	wire w_dff_B_FSFvBsOb9_1;
	wire w_dff_B_Wrp2cw9V8_1;
	wire w_dff_B_lF2gqh2j1_1;
	wire w_dff_B_kHduTWwA0_1;
	wire w_dff_B_yl1X8NTG2_0;
	wire w_dff_B_3uw3lwSe7_0;
	wire w_dff_B_0xyM49Sd7_0;
	wire w_dff_B_zbB4NiyC9_0;
	wire w_dff_B_CPor4q7G2_0;
	wire w_dff_B_BY634uEU1_0;
	wire w_dff_B_yIo78zmx4_0;
	wire w_dff_B_9ET7sr8X5_0;
	wire w_dff_B_Cat0Iyhn9_0;
	wire w_dff_B_MStUdTdf6_0;
	wire w_dff_B_pMQMIh1e3_0;
	wire w_dff_B_WsR0QEeq2_0;
	wire w_dff_B_DVauISiy6_0;
	wire w_dff_B_jcMwPvpN9_0;
	wire w_dff_B_EEVJq2m21_0;
	wire w_dff_B_cWMBAM437_0;
	wire w_dff_A_huryzMfF8_1;
	wire w_dff_A_DgfzQoCX4_1;
	wire w_dff_A_4DlfPjRV8_1;
	wire w_dff_A_sdEtRUsN7_1;
	wire w_dff_A_bvAjlEZl6_1;
	wire w_dff_B_BW1dvTRe2_0;
	wire w_dff_B_xEHoGlVx5_0;
	wire w_dff_B_PKDxjfiw4_0;
	wire w_dff_B_HylNPQSS2_0;
	wire w_dff_B_3oznaR7T2_0;
	wire w_dff_B_ZZyaLcAX0_1;
	wire w_dff_B_EOmmUq8M2_1;
	wire w_dff_B_fc3ZsHN80_1;
	wire w_dff_B_xdlkKpp82_1;
	wire w_dff_B_ybFmn4pW7_1;
	wire w_dff_B_jupaB5j52_1;
	wire w_dff_B_j71rhLtx1_1;
	wire w_dff_B_HlHsTkUR3_1;
	wire w_dff_B_2sqQBAbT8_1;
	wire w_dff_B_pkhHLovh9_1;
	wire w_dff_B_2qkoVUpD3_1;
	wire w_dff_B_SMdlVIcZ8_1;
	wire w_dff_B_iKDwu7rb1_1;
	wire w_dff_B_ld0lXjEs6_1;
	wire w_dff_B_LMygMd880_1;
	wire w_dff_B_EIyeCtko2_0;
	wire w_dff_B_I3CFtX3L4_0;
	wire w_dff_B_UsUkjvnh0_0;
	wire w_dff_B_XZ6M5iqW0_0;
	wire w_dff_B_qVPQL56h8_0;
	wire w_dff_B_uubzqeWb6_0;
	wire w_dff_A_L2TC5P8y6_0;
	wire w_dff_A_TFkQEriz5_0;
	wire w_dff_A_rkDR5gqQ1_0;
	wire w_dff_A_UtsoPKga7_0;
	wire w_dff_A_Wx3p4QbY8_0;
	wire w_dff_A_qQw0GRV41_0;
	wire w_dff_A_DhhcOSpl4_2;
	wire w_dff_A_WpOXLQxj0_0;
	wire w_dff_A_InH4zSMu5_0;
	wire w_dff_A_KDppmavv5_0;
	wire w_dff_A_cjxMoRST6_0;
	wire w_dff_A_vKL0uEsy8_0;
	wire w_dff_A_pRnFC8hN5_0;
	wire w_dff_B_oNIztZJx2_1;
	wire w_dff_A_UiZv4fgH0_0;
	wire w_dff_A_EXWGyaFA6_0;
	wire w_dff_A_vrWLk6sg1_0;
	wire w_dff_A_aYU9cUQL8_0;
	wire w_dff_A_IqClEjgr2_0;
	wire w_dff_A_4EofUg327_0;
	wire w_dff_A_tZ4AwOED6_0;
	wire w_dff_A_pSwKBWbz1_1;
	wire w_dff_A_MW8qoubo6_1;
	wire w_dff_A_Xgz0D3YQ3_1;
	wire w_dff_A_SjYP66qU4_1;
	wire w_dff_A_thKKhcRZ4_1;
	wire w_dff_A_fh4unqz22_1;
	wire w_dff_A_f8xT1ohz1_1;
	wire w_dff_A_CIkqZ35X6_1;
	wire w_dff_A_sx4S7KWf4_1;
	wire w_dff_B_N8KTnB2I2_0;
	wire w_dff_B_uRv1tsp57_0;
	wire w_dff_B_vydm3phq2_0;
	wire w_dff_A_7U5ieRNk3_1;
	wire w_dff_A_uQWYk0R27_1;
	wire w_dff_A_T76Z3dAe3_1;
	wire w_dff_A_S6lMnYu62_1;
	wire w_dff_A_0YjlXqxJ8_1;
	wire w_dff_A_dEhNGnlV1_1;
	wire w_dff_A_aUqhprmc4_1;
	wire w_dff_A_KCQnRKxQ9_2;
	wire w_dff_A_q9IxyWtg4_2;
	wire w_dff_A_3SHusknK0_2;
	wire w_dff_A_q559sriz3_2;
	wire w_dff_A_OV83fcgm3_2;
	wire w_dff_A_2jpIlMhI6_2;
	wire w_dff_A_7TkqrJOl2_2;
	wire w_dff_A_0M2689PP2_2;
	wire w_dff_A_URQcZCMA3_2;
	wire w_dff_A_lkYp9Zpr5_2;
	wire w_dff_A_JxVtyyyi3_2;
	wire w_dff_B_yyFbo49d6_0;
	wire w_dff_B_TIXSsHnR0_0;
	wire w_dff_B_NXsse0kV1_0;
	wire w_dff_B_yWLP7EiH7_0;
	wire w_dff_B_4PMOP45N0_0;
	wire w_dff_B_e7gYZnl19_0;
	wire w_dff_B_BUdIGe8i6_0;
	wire w_dff_B_2UpF74z99_0;
	wire w_dff_B_oQziZTJD0_0;
	wire w_dff_B_WOXq1yvj3_0;
	wire w_dff_B_gSzxI1sk5_0;
	wire w_dff_B_Q750Mzc63_0;
	wire w_dff_B_gXQZt7qG0_0;
	wire w_dff_B_P88vgw3G7_0;
	wire w_dff_B_inUkwTzK7_0;
	wire w_dff_B_c16ODci74_0;
	wire w_dff_A_qUxQ9eR06_1;
	wire w_dff_A_p7GWrnAN8_1;
	wire w_dff_A_PS2cKhNH5_1;
	wire w_dff_A_pWyCPHBM6_1;
	wire w_dff_A_iJQF7wRB4_1;
	wire w_dff_B_ewaCWjXU5_1;
	wire w_dff_A_ziZeDzT31_0;
	wire w_dff_A_RaHkYuxw1_0;
	wire w_dff_B_ch065sgI9_0;
	wire w_dff_B_U00YQBUU1_0;
	wire w_dff_B_2VWT5c7e6_0;
	wire w_dff_B_8yeMtSAO4_0;
	wire w_dff_B_WmH6Gm1u3_0;
	wire w_dff_B_P18D2B739_3;
	wire w_dff_A_0DXRBDIX9_2;
	wire w_dff_B_Kz50rcue2_3;
	wire w_dff_B_LgDm6vuh4_3;
	wire w_dff_B_4HzdEsCK4_3;
	wire w_dff_B_4tMDYC4K9_3;
	wire w_dff_B_140s6vK56_3;
	wire w_dff_B_PH4bYPh99_3;
	wire w_dff_B_K03bJey14_3;
	wire w_dff_B_UjLH3mI44_3;
	wire w_dff_A_oQjb4of25_0;
	wire w_dff_A_KxGzhUvM7_0;
	wire w_dff_A_U5CWkvmu4_0;
	wire w_dff_A_dx2ZBOYL5_0;
	wire w_dff_A_7bI26hNa9_0;
	wire w_dff_A_pUS09l1f8_0;
	wire w_dff_A_TjJq9c1D9_0;
	wire w_dff_A_TFGMO4fp7_0;
	wire w_dff_A_KSFyXSy63_1;
	wire w_dff_A_m7XBoiE86_1;
	wire w_dff_B_qY9kZGth2_3;
	wire w_dff_B_OQbLd5zZ4_3;
	wire w_dff_B_G2UFY6Yt5_3;
	wire w_dff_B_SV42AhMi0_3;
	wire w_dff_B_qW1mf6b35_3;
	wire w_dff_B_YsUscIKX4_3;
	wire w_dff_B_Rxkon8iU2_3;
	wire w_dff_B_rYQCJwdT3_3;
	wire w_dff_B_nKAgiXkD0_3;
	wire w_dff_B_z2BH0hU70_3;
	wire w_dff_B_fJmceP214_1;
	wire w_dff_B_QmXyJxHM7_1;
	wire w_dff_B_eFDD5lIT6_1;
	wire w_dff_B_4EaAiSk57_1;
	wire w_dff_B_XcNkQ3955_1;
	wire w_dff_B_TVyze9Fy4_1;
	wire w_dff_B_ZF17TUEo5_1;
	wire w_dff_B_Ar3zaphe0_1;
	wire w_dff_B_zJD5ybiD5_1;
	wire w_dff_B_ZHTnix634_1;
	wire w_dff_B_4SqrJTfl3_1;
	wire w_dff_B_PFjDtg4p9_1;
	wire w_dff_B_umwW1L8p1_1;
	wire w_dff_B_aLqQkBwY6_1;
	wire w_dff_B_1NpAaQFN7_1;
	wire w_dff_B_iItLI2ul9_1;
	wire w_dff_B_2iVXjyDC6_1;
	wire w_dff_B_Ta0E71Dt8_0;
	wire w_dff_B_GiH63RCn7_0;
	wire w_dff_B_Oi1XeFGe5_0;
	wire w_dff_B_eZYDo9mQ2_0;
	wire w_dff_B_ysGrVblS0_0;
	wire w_dff_B_Mf2Gmwc63_0;
	wire w_dff_B_Zzqx5ko26_0;
	wire w_dff_A_kap8HMGd4_0;
	wire w_dff_A_uJK28g8t6_0;
	wire w_dff_A_hS4ktZtB8_0;
	wire w_dff_A_8i1GiwGN4_0;
	wire w_dff_A_Dq02Xrdc6_0;
	wire w_dff_A_gs9QbbYH8_0;
	wire w_dff_A_VNpFfYvM2_0;
	wire w_dff_A_R4JOrNwX5_0;
	wire w_dff_A_U6uXdiMU8_0;
	wire w_dff_A_RSAXALUE6_0;
	wire w_dff_A_o2mseczl8_0;
	wire w_dff_A_SEgK1xpa1_0;
	wire w_dff_A_s5KWcoQS1_0;
	wire w_dff_A_PTCrlAKa4_0;
	wire w_dff_B_8rJVeBf71_1;
	wire w_dff_B_j52NSK681_1;
	wire w_dff_B_i0BDKuiQ0_1;
	wire w_dff_B_4cjapgEs7_1;
	wire w_dff_B_TXmJT4UW2_1;
	wire w_dff_B_ZtESkSFn5_1;
	wire w_dff_B_PhMd6PAC4_1;
	wire w_dff_B_GqeoQfkK0_1;
	wire w_dff_B_VkeglazP1_1;
	wire w_dff_B_AGYNsHQ40_0;
	wire w_dff_A_QY1RKPjN8_0;
	wire w_dff_B_oKHxCJyl8_1;
	wire w_dff_A_gzShykAk1_0;
	wire w_dff_A_QMTfVDiR1_0;
	wire w_dff_A_9Lkwfsre6_0;
	wire w_dff_A_yEADm3ZI5_1;
	wire w_dff_A_s9XObmOD2_1;
	wire w_dff_A_UffxUXah3_1;
	wire w_dff_A_DJr3SYUW9_1;
	wire w_dff_A_Pu6abALy1_1;
	wire w_dff_A_ydeSI1L21_1;
	wire w_dff_A_ElakrV2A5_1;
	wire w_dff_A_2cjpNXO87_1;
	wire w_dff_A_mIwPmc5u6_2;
	wire w_dff_A_gOLB3rRu6_2;
	wire w_dff_A_sWud1j4Y0_2;
	wire w_dff_A_6QEMRrhw2_2;
	wire w_dff_A_yE7BqAgf8_2;
	wire w_dff_A_Aq3CPh3H7_2;
	wire w_dff_A_4GZ83DDk1_2;
	wire w_dff_A_Tk84Qdly2_2;
	wire w_dff_A_bUrEAGsK5_1;
	wire w_dff_A_ehd9gxtr1_1;
	wire w_dff_A_prgsGZBy1_1;
	wire w_dff_A_pEyQRMFm9_1;
	wire w_dff_A_uJTE1h3o9_1;
	wire w_dff_A_8ZlUDxPu3_1;
	wire w_dff_A_6o1fz2mx1_1;
	wire w_dff_A_5UNrjDdz5_1;
	wire w_dff_A_SyNsnOxU5_2;
	wire w_dff_A_V3fCSbYc7_2;
	wire w_dff_A_QwUCHtfL3_2;
	wire w_dff_A_eRq5pqKb6_2;
	wire w_dff_A_arRvqP0e4_2;
	wire w_dff_A_UuNH3cPQ9_2;
	wire w_dff_A_G37BWPzY1_2;
	wire w_dff_A_wLIgF7JD4_2;
	wire w_dff_B_NblQoCvy0_0;
	wire w_dff_A_P4A3xGbv7_0;
	wire w_dff_A_mARZLVck7_0;
	wire w_dff_A_xsDiUmav4_0;
	wire w_dff_B_Y91cRz3S3_1;
	wire w_dff_A_7v4YJTJZ3_0;
	wire w_dff_A_rD5nbX0R4_0;
	wire w_dff_A_leEiRrE34_0;
	wire w_dff_A_oB26pOZI7_0;
	wire w_dff_A_IsZfT29g9_0;
	wire w_dff_A_CRBlKU8z2_0;
	wire w_dff_A_6zm24qyD0_0;
	wire w_dff_A_Za1CKhsi4_0;
	wire w_dff_A_IjWelpfO1_0;
	wire w_dff_A_dJS1UTvR7_0;
	wire w_dff_A_Yz8mIEtH6_0;
	wire w_dff_A_FyBZqUeG8_0;
	wire w_dff_A_XMcUX3AP0_0;
	wire w_dff_A_dG0yYy4j0_2;
	wire w_dff_A_rQcTeXgG2_2;
	wire w_dff_A_4Kmdv6234_2;
	wire w_dff_A_8fG1lPkj0_2;
	wire w_dff_B_eenTpDDo4_1;
	wire w_dff_A_EcDp1A0e3_1;
	wire w_dff_A_BAnzpPqS4_1;
	wire w_dff_A_E7TWcOqN9_1;
	wire w_dff_A_ihDrd5km5_1;
	wire w_dff_A_s4lNmvvS8_1;
	wire w_dff_A_Utnvb7700_1;
	wire w_dff_B_T9mntcNv1_2;
	wire w_dff_B_wW0G0AWt7_2;
	wire w_dff_B_2S2tHoPe4_2;
	wire w_dff_B_RUCXEpUo8_2;
	wire w_dff_A_PBwWq9Ye3_0;
	wire w_dff_A_pHgR9PWW7_0;
	wire w_dff_A_tlyHrYGw4_0;
	wire w_dff_A_Tinws3kd7_0;
	wire w_dff_A_NmpuEUa86_0;
	wire w_dff_A_K3N3Zj0k7_0;
	wire w_dff_A_s1QoyaYE4_0;
	wire w_dff_A_F0P8hhOf4_0;
	wire w_dff_A_HuTQ1mql8_2;
	wire w_dff_A_jSXmu9qJ3_2;
	wire w_dff_A_ZEKpD2X67_2;
	wire w_dff_A_PhIG9if66_2;
	wire w_dff_B_rRFD66SL8_1;
	wire w_dff_B_23pPR6AI7_1;
	wire w_dff_B_FJZYVjBF8_1;
	wire w_dff_B_WdfitJyc1_1;
	wire w_dff_B_6xEaZtyY8_1;
	wire w_dff_B_yNef5tfK2_1;
	wire w_dff_B_heYskH6L4_1;
	wire w_dff_B_IJ6JFvqV3_1;
	wire w_dff_B_VhjGV70K6_1;
	wire w_dff_B_LtJRveWy4_1;
	wire w_dff_B_tp0AYuUa2_0;
	wire w_dff_B_GxaiRH1j7_0;
	wire w_dff_B_2LNkqAIQ2_1;
	wire w_dff_B_tDCpdrd55_1;
	wire w_dff_B_9Y1OM4CG8_1;
	wire w_dff_B_5ATfsu0t5_1;
	wire w_dff_B_yTizZ9lw6_1;
	wire w_dff_B_9Z2GTdBA3_1;
	wire w_dff_B_PIH3NLKl1_1;
	wire w_dff_B_QMDI3G081_1;
	wire w_dff_B_a3dEcDtW3_1;
	wire w_dff_B_FSuwRInr5_2;
	wire w_dff_B_rwbBHnH30_2;
	wire w_dff_B_uDz6Pol31_2;
	wire w_dff_B_bEuC7WNx2_2;
	wire w_dff_B_MzMoJbgy6_2;
	wire w_dff_B_TkhH7ngz6_2;
	wire w_dff_B_Ae9ugOcq8_2;
	wire w_dff_B_PUmuuksv1_2;
	wire w_dff_B_Ef3RQZoT8_2;
	wire w_dff_A_9oXkUTAz9_0;
	wire w_dff_A_wk1SUM0p8_0;
	wire w_dff_A_UEIPtOM79_0;
	wire w_dff_A_SVW2ApoK0_0;
	wire w_dff_A_hZAmTO0x5_0;
	wire w_dff_A_gfX8I5vR0_0;
	wire w_dff_A_qlmLcpAJ4_0;
	wire w_dff_A_b5D8cxwH4_0;
	wire w_dff_A_olrTfMMo1_0;
	wire w_dff_A_kPOlzqhg9_1;
	wire w_dff_A_CVsh6Tod2_1;
	wire w_dff_A_pHweGRNG9_1;
	wire w_dff_A_l3yf2L599_1;
	wire w_dff_A_GeyWpXcm2_1;
	wire w_dff_A_9032q7DC3_1;
	wire w_dff_A_Xu3zxC3c8_1;
	wire w_dff_A_yUHVYSVi6_1;
	wire w_dff_A_VDf97yrT4_1;
	wire w_dff_A_djOBsNTk8_0;
	wire w_dff_A_MeVNwU9y6_1;
	wire w_dff_A_W3FLjjEm2_0;
	wire w_dff_A_fUIRF1uh8_0;
	wire w_dff_A_jijkFqLL6_0;
	wire w_dff_A_SXSa9Abc2_0;
	wire w_dff_A_kj7LiY6u0_0;
	wire w_dff_A_Hjd5HB6V7_1;
	wire w_dff_A_1KrbjPmR9_1;
	wire w_dff_A_qM5UkkSD5_1;
	wire w_dff_A_QzOt0Dxq5_1;
	wire w_dff_A_9lvKOKTJ5_1;
	wire w_dff_A_nrpS9ytr7_1;
	wire w_dff_A_jUu6GTGU5_1;
	wire w_dff_A_zEIzOYzO8_1;
	wire w_dff_A_LWe7mISb3_2;
	wire w_dff_A_gI9avPq63_2;
	wire w_dff_A_anHXxQlP3_2;
	wire w_dff_A_L2PRPBEx7_2;
	wire w_dff_A_Jr0aNAZ54_2;
	wire w_dff_A_kgqIfa3Q5_2;
	wire w_dff_A_XzTdvpy37_2;
	wire w_dff_A_kSeB5CQy5_2;
	wire w_dff_A_jcTRIs114_2;
	wire w_dff_A_1GLIPFkh8_2;
	wire w_dff_A_DGiQDqBx1_2;
	wire w_dff_A_pdf0eo104_2;
	wire w_dff_A_mfbB0nMc5_1;
	wire w_dff_A_kbszwEzd6_1;
	wire w_dff_A_TOf5ODXz5_1;
	wire w_dff_A_YURtj78C0_1;
	wire w_dff_A_sZsdzTaB7_1;
	wire w_dff_A_0zPqIFrs3_1;
	wire w_dff_A_F9C2ZxEi1_1;
	wire w_dff_A_86cfAmWR2_1;
	wire w_dff_A_BCpoGdPS7_1;
	wire w_dff_B_rOE8WGvz2_1;
	wire w_dff_A_JZ7jqKdK4_1;
	wire w_dff_A_EjSzGy6S4_1;
	wire w_dff_A_7b2uoo306_1;
	wire w_dff_A_zjJiOsop4_1;
	wire w_dff_A_qrJOZv860_1;
	wire w_dff_A_oEzKJrnh1_1;
	wire w_dff_A_wJXMRtTS0_1;
	wire w_dff_A_VOkRqBMv5_2;
	wire w_dff_A_yK5wcWlf3_2;
	wire w_dff_A_N3VGMkfp7_1;
	wire w_dff_A_TypNUBOb1_1;
	wire w_dff_A_ND8Jvmt28_2;
	wire w_dff_A_OdzPs9rg2_2;
	wire w_dff_B_18olbLOP0_0;
	wire w_dff_A_KFfwWjQ50_0;
	wire w_dff_A_hIL54dP46_0;
	wire w_dff_A_P9EaKFnE3_0;
	wire w_dff_A_mLdU7aep6_1;
	wire w_dff_B_CFEopYXd6_2;
	wire w_dff_B_uU4fkVGW5_2;
	wire w_dff_B_8EmUAwgh0_2;
	wire w_dff_B_B0ihQo9d3_2;
	wire w_dff_A_QYu2gx179_0;
	wire w_dff_A_340dqXtv2_0;
	wire w_dff_A_D1NNrqd31_0;
	wire w_dff_A_FPNrMZMq6_0;
	wire w_dff_A_iXqca1Zk3_0;
	wire w_dff_A_aNX4dK6Y4_0;
	wire w_dff_A_JV25cchI2_0;
	wire w_dff_A_KKyrQJND4_0;
	wire w_dff_A_n8jyaAOY5_1;
	wire w_dff_A_pGiu4Gew8_1;
	wire w_dff_A_saBQNKzF6_1;
	wire w_dff_A_1QSSEYiG4_1;
	wire w_dff_A_RWnSet5j4_2;
	wire w_dff_A_LWWM06jf9_2;
	wire w_dff_A_dgh7e4WD9_2;
	wire w_dff_A_h6RLW3107_2;
	wire w_dff_A_6z70m9va4_2;
	wire w_dff_A_2Jj8F1tu7_2;
	wire w_dff_A_El1Nxp5O6_2;
	wire w_dff_A_Wr5l3qB80_2;
	wire w_dff_A_25Bq4v7R0_0;
	wire w_dff_A_MaDjIIkD6_0;
	wire w_dff_A_hsXq72MK2_0;
	wire w_dff_A_cOGD7dtu3_0;
	wire w_dff_A_dlplJRp08_0;
	wire w_dff_A_aCCnIhpQ0_0;
	wire w_dff_A_5anbM8rR4_0;
	wire w_dff_A_wYIkLhg66_0;
	wire w_dff_B_ij8LaE1r7_0;
	wire w_dff_B_byONNthQ6_0;
	wire w_dff_B_fkJQA9hn5_0;
	wire w_dff_A_vQFXgHor2_0;
	wire w_dff_A_xgh1ZQUf4_0;
	wire w_dff_A_pxaxEmwM6_0;
	wire w_dff_A_ehEewFN31_0;
	wire w_dff_A_CKg17ZEl4_2;
	wire w_dff_A_B3TbiyQQ6_2;
	wire w_dff_A_62hqqsVn3_2;
	wire w_dff_A_wlkSUAub8_2;
	wire w_dff_A_x5CwquCG5_2;
	wire w_dff_A_VquKTESQ3_0;
	wire w_dff_A_k9WQmgek1_0;
	wire w_dff_A_jssz4fDF0_0;
	wire w_dff_A_mV4frAKc3_0;
	wire w_dff_A_J5Vh6mSc0_0;
	wire w_dff_A_t1Rginlm8_1;
	wire w_dff_A_pWOIEiwN4_1;
	wire w_dff_A_edomZr5R7_1;
	wire w_dff_A_O5YKIHQ91_1;
	wire w_dff_A_XVL3MtqC0_1;
	wire w_dff_A_0A1pbHjQ5_1;
	wire w_dff_A_6sPlPBXq0_1;
	wire w_dff_A_F6E0aPbK6_2;
	wire w_dff_A_0SEFSqob5_2;
	wire w_dff_A_qCHLWT0n2_2;
	wire w_dff_A_DBtylpiE6_2;
	wire w_dff_A_0f6e43BR3_2;
	wire w_dff_A_L3hODdFd9_2;
	wire w_dff_A_VvwERKv35_2;
	wire w_dff_A_AgMBfGcu6_2;
	wire w_dff_A_98Ja3Kgg6_2;
	wire w_dff_A_3wT5SbGB2_2;
	wire w_dff_A_Hpxb2jRc1_2;
	wire w_dff_A_RUWEpb3u7_1;
	wire w_dff_A_NlhHi1S28_1;
	wire w_dff_A_J9JUekAm4_1;
	wire w_dff_A_SdNXbEZS2_1;
	wire w_dff_A_92ZoAiBn5_1;
	wire w_dff_A_L1hqvV9p8_1;
	wire w_dff_A_IfxB44gw2_1;
	wire w_dff_A_QL01JIBY2_1;
	wire w_dff_A_ndz4jTRC8_1;
	wire w_dff_B_AadmqBjn3_0;
	wire w_dff_B_8IsVf4RO3_0;
	wire w_dff_B_rzvQ8ikQ1_0;
	wire w_dff_B_jjjjMfHr1_0;
	wire w_dff_A_jI7X4yov3_0;
	wire w_dff_A_vCcubefC6_2;
	wire w_dff_A_bG7K8tIg9_2;
	wire w_dff_A_Om4YmTQj9_2;
	wire w_dff_A_meywaUyO7_0;
	wire w_dff_A_VxBXljXt1_2;
	wire w_dff_A_7gBdB4nI1_0;
	wire w_dff_A_g22o4OSZ5_0;
	wire w_dff_A_nCZDJcW77_0;
	wire w_dff_A_Xxz2xkIl5_1;
	wire w_dff_A_4JNFA8PX0_1;
	wire w_dff_B_ivJ2mVzD1_2;
	wire w_dff_B_Di0xFvKN4_2;
	wire w_dff_B_3xDweony9_2;
	wire w_dff_B_OZVGGOE57_2;
	wire w_dff_B_udpERRFX2_0;
	wire w_dff_A_Z8XJFfMx8_0;
	wire w_dff_A_tixy5xj33_0;
	wire w_dff_B_zETTW3TP2_0;
	wire w_dff_A_wQHYWXrg3_1;
	wire w_dff_A_mLhQAz6c5_1;
	wire w_dff_A_2nGZXnCE3_1;
	wire w_dff_A_DevPPZdC5_1;
	wire w_dff_A_YQB8dx4G5_1;
	wire w_dff_A_Mjm2LAJE6_1;
	wire w_dff_A_PGiJWcjm6_1;
	wire w_dff_A_w0p67XqF8_1;
	wire w_dff_A_dlIc9bHV9_1;
	wire w_dff_A_xkfjvA3f2_1;
	wire w_dff_A_HZUBRvl41_1;
	wire w_dff_A_Pa5fHq2F2_1;
	wire w_dff_A_YRAMphzX3_1;
	wire w_dff_A_36VyoqI13_1;
	wire w_dff_A_BZTn2BFP9_1;
	wire w_dff_A_MyGsg31O7_1;
	wire w_dff_A_8l8ryIwm9_1;
	wire w_dff_A_LYfBYSkL1_1;
	wire w_dff_A_x6DKqCwF4_1;
	wire w_dff_A_PSEKKTS35_1;
	wire w_dff_A_vxilYzBx3_2;
	wire w_dff_A_374xxYkZ3_2;
	wire w_dff_A_rGL5bg8K7_2;
	wire w_dff_A_mUtRlnah9_2;
	wire w_dff_A_LvBbnYVl7_2;
	wire w_dff_A_ksBnd4vT7_2;
	wire w_dff_A_GlMLFNvK1_2;
	wire w_dff_A_yKX2EfqP3_2;
	wire w_dff_A_6w2Q1Ity1_2;
	wire w_dff_A_ShPDGQPY9_2;
	wire w_dff_A_rs2z8Iys3_2;
	wire w_dff_A_Xntldy6t4_2;
	wire w_dff_A_KbI1O0Li6_0;
	wire w_dff_A_HwD9Gvsd8_0;
	wire w_dff_A_6RLNHJ3f8_0;
	wire w_dff_A_wzzlXE2A3_0;
	wire w_dff_A_OjMacc4E8_0;
	wire w_dff_A_iezIhc946_0;
	wire w_dff_A_fRI2OmYX3_0;
	wire w_dff_A_MbDeBTxb1_0;
	wire w_dff_A_dBKiL6a15_0;
	wire w_dff_A_L5orFgfL4_0;
	wire w_dff_A_joDeA7Tv2_0;
	wire w_dff_A_VPyLGf2T4_0;
	wire w_dff_A_dNkfhZNP1_0;
	wire w_dff_A_mwe0rlSt2_0;
	wire w_dff_A_kykKmry83_0;
	wire w_dff_A_fx5Guiuz6_0;
	wire w_dff_A_oDP3HgJm7_0;
	wire w_dff_A_MuDXKnsO6_0;
	wire w_dff_A_8q4hYZEa0_2;
	wire w_dff_A_xPTbtNGZ8_0;
	wire w_dff_A_wZm4wPkt0_0;
	wire w_dff_A_4UIBkS5G1_0;
	wire w_dff_A_l2vojIM87_0;
	wire w_dff_A_jV5KMfvS1_0;
	wire w_dff_A_T3vNj6o98_0;
	wire w_dff_A_OCkaEYu48_0;
	wire w_dff_A_zWRMz6nS0_0;
	wire w_dff_A_8zyTGUr33_0;
	wire w_dff_A_im91KOK28_0;
	wire w_dff_A_B2nULJo43_0;
	wire w_dff_A_BVUtzsI27_0;
	wire w_dff_A_RCIQiXpR9_0;
	wire w_dff_A_OfzcEk0X5_0;
	wire w_dff_A_ghzDh9FC4_0;
	wire w_dff_A_5evEE28F3_0;
	wire w_dff_A_IE8ejD1K8_0;
	wire w_dff_A_oq4UU4ah3_0;
	wire w_dff_A_LZkuzL3R5_2;
	wire w_dff_A_sTC6SooE5_0;
	wire w_dff_A_eo7wdQuK5_0;
	wire w_dff_A_pJscz6Kw9_0;
	wire w_dff_A_XrcXhGWw7_0;
	wire w_dff_A_JpPtK6Xf6_0;
	wire w_dff_A_bCngngao2_0;
	wire w_dff_A_z7vWbgRv5_0;
	wire w_dff_A_zwT3vDpk8_0;
	wire w_dff_A_RptEAGvp9_0;
	wire w_dff_A_Upvtfp5Y1_0;
	wire w_dff_A_ODUjvdJN6_0;
	wire w_dff_A_CoaYQUCE6_0;
	wire w_dff_A_sXex1YRa4_0;
	wire w_dff_A_JLiOVXCq5_0;
	wire w_dff_A_RJFpea0H9_0;
	wire w_dff_A_oXGKYB0N7_0;
	wire w_dff_A_izYa1v5x2_0;
	wire w_dff_A_AaRMdoEz8_0;
	wire w_dff_A_lNIUOv8Z3_2;
	wire w_dff_A_9QuSUTrw6_0;
	wire w_dff_A_s1sbIzuM7_0;
	wire w_dff_A_n8nz6vkt2_0;
	wire w_dff_A_JGm44D9l8_0;
	wire w_dff_A_QFMfETWL7_0;
	wire w_dff_A_9BQeGxpk9_0;
	wire w_dff_A_ZjoVzQfi6_0;
	wire w_dff_A_EfirJdH51_0;
	wire w_dff_A_GTAl8Tye4_0;
	wire w_dff_A_JFhCzmdc7_0;
	wire w_dff_A_q64hj3Sz5_0;
	wire w_dff_A_CuQ7muhK0_0;
	wire w_dff_A_PFSyVOOQ3_0;
	wire w_dff_A_FA5wy5YP7_0;
	wire w_dff_A_yd0fbcGO0_0;
	wire w_dff_A_jqhYfzFw6_0;
	wire w_dff_A_bCZxmP5L5_0;
	wire w_dff_A_7Ym21FOd6_0;
	wire w_dff_A_IyfHgiX69_0;
	wire w_dff_A_LcBxnPK44_2;
	wire w_dff_A_EVmSVshh4_0;
	wire w_dff_A_TAvlpuRY5_0;
	wire w_dff_A_Ng5jKy9L0_0;
	wire w_dff_A_oSDL6rJH2_0;
	wire w_dff_A_0CZpg5L10_0;
	wire w_dff_A_YTyortLz5_0;
	wire w_dff_A_eZia1YNg5_0;
	wire w_dff_A_jhD9kbtS6_0;
	wire w_dff_A_mgNjCEzV9_0;
	wire w_dff_A_4BTToW5j4_0;
	wire w_dff_A_UaT1PotL7_0;
	wire w_dff_A_6WAL0zSB2_0;
	wire w_dff_A_EXVPbxuf8_0;
	wire w_dff_A_65LjyrMF7_0;
	wire w_dff_A_vNuX6L9g4_0;
	wire w_dff_A_oblXIxF02_0;
	wire w_dff_A_FwO04bgL3_0;
	wire w_dff_A_JrWkhz5v5_0;
	wire w_dff_A_om5yfFJZ9_2;
	wire w_dff_A_wFkHDRkN0_0;
	wire w_dff_A_7DIPzXgA2_0;
	wire w_dff_A_kSQEXk5g5_0;
	wire w_dff_A_ca2QhFIc0_0;
	wire w_dff_A_6C7OKgw35_0;
	wire w_dff_A_Fp8rfe5R6_0;
	wire w_dff_A_8hsaQADq1_0;
	wire w_dff_A_zjvc2mYh4_0;
	wire w_dff_A_pgd1iREk3_0;
	wire w_dff_A_lbwzw8Zt0_0;
	wire w_dff_A_Mx92Rox19_0;
	wire w_dff_A_2jcBRt5V6_0;
	wire w_dff_A_u1Dr9DA03_0;
	wire w_dff_A_un9KlenZ7_0;
	wire w_dff_A_JZbjTR1k7_0;
	wire w_dff_A_fXPC6ktv8_0;
	wire w_dff_A_HeZ3jRFr2_2;
	wire w_dff_A_GWeUZ3Ph0_0;
	wire w_dff_A_BxQg5xdj5_0;
	wire w_dff_A_Lft3Zjlj3_0;
	wire w_dff_A_hRVzl9vg0_0;
	wire w_dff_A_vIGz3kAM3_0;
	wire w_dff_A_jKLSxyQb1_0;
	wire w_dff_A_eS3lpG7T6_0;
	wire w_dff_A_NA1xOXbL2_0;
	wire w_dff_A_9uZsmQkm2_0;
	wire w_dff_A_sb4fYoiv4_0;
	wire w_dff_A_fOJCMub76_0;
	wire w_dff_A_Y4gymV6T2_0;
	wire w_dff_A_IALfDD7n7_0;
	wire w_dff_A_VUkdmvpH5_0;
	wire w_dff_A_BN6dc5Vf5_0;
	wire w_dff_A_KC6954ZE3_0;
	wire w_dff_A_4BtlkvJK0_0;
	wire w_dff_A_fN7Sqhtz9_2;
	wire w_dff_A_X4vtqVKS5_0;
	wire w_dff_A_0V4AT2zD8_0;
	wire w_dff_A_AsYtUIVv9_0;
	wire w_dff_A_PtWdQm3q7_0;
	wire w_dff_A_2Ngi02M84_0;
	wire w_dff_A_mkmWWU8L8_0;
	wire w_dff_A_0GJzQxL10_0;
	wire w_dff_A_2xGe2Emd1_0;
	wire w_dff_A_EuNUbaaj2_0;
	wire w_dff_A_taDBZjTd4_0;
	wire w_dff_A_LFjYlNYn7_0;
	wire w_dff_A_R67gdMvw8_0;
	wire w_dff_A_m6nrYg2h5_0;
	wire w_dff_A_SaxFcQyt3_0;
	wire w_dff_A_9gk8OFil8_0;
	wire w_dff_A_tgQpqa4J2_0;
	wire w_dff_A_y9CJdFj68_0;
	wire w_dff_A_HLc1PW0D5_2;
	wire w_dff_A_xkvkgoy20_0;
	wire w_dff_A_NVy69MsY1_0;
	wire w_dff_A_BmKjPyn96_0;
	wire w_dff_A_CkY47CdA6_0;
	wire w_dff_A_eEf2ED1m7_0;
	wire w_dff_A_hmTwZ0ud4_0;
	wire w_dff_A_6e4D3hyf4_0;
	wire w_dff_A_ESJRskFL9_0;
	wire w_dff_A_tS4za1nY9_0;
	wire w_dff_A_1bBMaS7h7_0;
	wire w_dff_A_ywJAphae0_0;
	wire w_dff_A_ySyXdsmH1_0;
	wire w_dff_A_FNxxjxIv1_0;
	wire w_dff_A_IxHs60Sp0_0;
	wire w_dff_A_tcaDIE257_0;
	wire w_dff_A_ySiKg4xZ1_0;
	wire w_dff_A_ZpIgaS6M9_0;
	wire w_dff_A_iMewsF9N8_2;
	wire w_dff_A_vaSG4d708_0;
	wire w_dff_A_x4SuF3BL8_0;
	wire w_dff_A_szAv4nas4_0;
	wire w_dff_A_qtlPwTV65_0;
	wire w_dff_A_NiMiWQJ36_0;
	wire w_dff_A_sjNa6rfS2_0;
	wire w_dff_A_lmO4PdFJ0_0;
	wire w_dff_A_HaEKUkna8_0;
	wire w_dff_A_odmub6DX6_0;
	wire w_dff_A_jHBi5Bfo5_0;
	wire w_dff_A_toBZB2Nw6_0;
	wire w_dff_A_QIzUUu018_0;
	wire w_dff_A_H6to52x65_0;
	wire w_dff_A_SoN1Y4fW7_0;
	wire w_dff_A_GBXdkGzH7_0;
	wire w_dff_A_bNeRAaKI0_0;
	wire w_dff_A_YEhqLxN09_0;
	wire w_dff_A_SaCeGyxV2_0;
	wire w_dff_A_qRuj8HhM0_2;
	wire w_dff_A_71EuurKe6_0;
	wire w_dff_A_0RLeOXEr3_0;
	wire w_dff_A_JCDd51sk5_0;
	wire w_dff_A_cQ3UmHPN5_0;
	wire w_dff_A_3s5bnS9l2_0;
	wire w_dff_A_e48IVaOt7_0;
	wire w_dff_A_Pv9jvW6z7_0;
	wire w_dff_A_Cvz3BPRS8_0;
	wire w_dff_A_4NBxotBM5_0;
	wire w_dff_A_DA1vM29x0_0;
	wire w_dff_A_79i2WSZs8_0;
	wire w_dff_A_yTO5944o6_0;
	wire w_dff_A_L8zE4EKL6_0;
	wire w_dff_A_aeihurQx3_0;
	wire w_dff_A_rUFO2HwF2_0;
	wire w_dff_A_Te4VIOed3_0;
	wire w_dff_A_4xqBO2HF8_1;
	wire w_dff_A_somV81jX7_0;
	wire w_dff_A_eitVJNG94_0;
	wire w_dff_A_I2OjUYlH3_0;
	wire w_dff_A_oxdftX4d5_0;
	wire w_dff_A_bd3ws9tz4_0;
	wire w_dff_A_9Ojln7L75_0;
	wire w_dff_A_G878MytB8_0;
	wire w_dff_A_dScHZvv86_0;
	wire w_dff_A_MRbRN5f95_0;
	wire w_dff_A_B5ScHvZj1_0;
	wire w_dff_A_PAKlTkdn2_0;
	wire w_dff_A_Me6gvWQp7_0;
	wire w_dff_A_hS4DMq2w7_0;
	wire w_dff_A_1gFLst8r9_0;
	wire w_dff_A_a8ybMeff9_0;
	wire w_dff_A_yuPIEYgL9_0;
	wire w_dff_A_uee924xu4_0;
	wire w_dff_A_UKevBCaG4_0;
	wire w_dff_A_dO4Fam3e8_2;
	wire w_dff_A_uEPPxuz07_0;
	wire w_dff_A_rHzmUiJb4_0;
	wire w_dff_A_9R1MTHIf6_0;
	wire w_dff_A_dUecXQBk2_0;
	wire w_dff_A_05pOeuiE3_0;
	wire w_dff_A_5T3pQLEH4_0;
	wire w_dff_A_AD7lS7079_0;
	wire w_dff_A_zDJfbgFf2_0;
	wire w_dff_A_OD5qzNsb7_0;
	wire w_dff_A_P8ioZ82P7_0;
	wire w_dff_A_vGMP4ftZ9_0;
	wire w_dff_A_1BoVzjbG2_0;
	wire w_dff_A_i0PaspVa8_0;
	wire w_dff_A_KSkfFaDD8_0;
	wire w_dff_A_z1D2e0wE6_0;
	wire w_dff_A_AABn1yD90_0;
	wire w_dff_A_PWvanrdV6_0;
	wire w_dff_A_6MABsAz43_2;
	wire w_dff_A_oYESdbrw1_0;
	wire w_dff_A_JZxxlBLw0_0;
	wire w_dff_A_Ci9vNr2o4_0;
	wire w_dff_A_cqtx839A6_0;
	wire w_dff_A_QKyXmqNM5_0;
	wire w_dff_A_0SU8pNDo8_0;
	wire w_dff_A_meCZUS2W1_0;
	wire w_dff_A_xSsipH7N6_0;
	wire w_dff_A_1DriepDL8_0;
	wire w_dff_A_V19H7jzo8_0;
	wire w_dff_A_67hsqkPb6_0;
	wire w_dff_A_SNaqiekO6_0;
	wire w_dff_A_bZ2cGZRe5_0;
	wire w_dff_A_itEyNGxY3_0;
	wire w_dff_A_qg0kKzdK2_0;
	wire w_dff_A_bUch3oDI5_0;
	wire w_dff_A_CVZsVZfq1_0;
	wire w_dff_A_R1GJVanS7_2;
	wire w_dff_A_3v28Pjlo6_0;
	wire w_dff_A_b8K0qLE62_0;
	wire w_dff_A_BTi0qHKI5_0;
	wire w_dff_A_e3LTPdoj2_0;
	wire w_dff_A_2BCrTTh28_0;
	wire w_dff_A_uHLLDC1h5_0;
	wire w_dff_A_hHnDGNkM0_0;
	wire w_dff_A_atHNo8x77_0;
	wire w_dff_A_TjjxhGX70_0;
	wire w_dff_A_F7tNoc4t7_0;
	wire w_dff_A_02XtJSan5_0;
	wire w_dff_A_JRDzSJiE3_0;
	wire w_dff_A_RfVujGfb7_0;
	wire w_dff_A_PL7iiSe06_0;
	wire w_dff_A_NBRDja6d9_0;
	wire w_dff_A_9O6Idaah6_0;
	wire w_dff_A_H5TRvcPw8_0;
	wire w_dff_A_1mp9vioA7_0;
	wire w_dff_A_LvQP9xlj5_2;
	wire w_dff_A_tLfWjOPN7_0;
	wire w_dff_A_M8z8ftOG6_0;
	wire w_dff_A_lNhERKjM8_0;
	wire w_dff_A_tQKRItzr2_0;
	wire w_dff_A_RZKfr7rY2_0;
	wire w_dff_A_ssCfw2zJ8_0;
	wire w_dff_A_TvZkicBx4_0;
	wire w_dff_A_CSpgTGcP4_0;
	wire w_dff_A_b0r2iFMB7_0;
	wire w_dff_A_6dHyje1g9_0;
	wire w_dff_A_fepdQ3Ka4_0;
	wire w_dff_A_oe72zPQP5_0;
	wire w_dff_A_f40m703a5_0;
	wire w_dff_A_mZmqsYz20_0;
	wire w_dff_A_Pk8fqNE29_0;
	wire w_dff_A_hNmiyPSM6_0;
	wire w_dff_A_0r3C9dNv8_2;
	wire w_dff_A_Mc5hPslK9_0;
	wire w_dff_A_eH3k3LpP5_0;
	wire w_dff_A_ypaW0iCC9_0;
	wire w_dff_A_hkqX09064_0;
	wire w_dff_A_FDkR9MnI9_0;
	wire w_dff_A_TS5Kuw7M7_0;
	wire w_dff_A_pxVKceKG3_0;
	wire w_dff_A_8ofwVCIM1_0;
	wire w_dff_A_vOrzP7sF6_0;
	wire w_dff_A_ci6z7g5X6_0;
	wire w_dff_A_F19in5ad1_0;
	wire w_dff_A_LBMcHvg94_0;
	wire w_dff_A_QDsrD8c49_0;
	wire w_dff_A_VY2Sqll62_0;
	wire w_dff_A_TDRq9fEl1_0;
	wire w_dff_A_labbdHJQ5_0;
	wire w_dff_A_NdwaEkVp4_2;
	wire w_dff_A_iFhP6lex2_0;
	wire w_dff_A_wR1Kedpq4_0;
	wire w_dff_A_pB1RTRaH4_0;
	wire w_dff_A_qLrAg3sh5_0;
	wire w_dff_A_oZJQVz7Q7_0;
	wire w_dff_A_TyT9jA6O1_0;
	wire w_dff_A_9uLBxE1F1_0;
	wire w_dff_A_TtRDAdvq8_2;
	wire w_dff_A_Bj362FUu5_0;
	wire w_dff_A_DOjFwhZ78_0;
	wire w_dff_A_TBwLhrZr3_0;
	wire w_dff_A_rFZzsmmR5_2;
	wire w_dff_A_WqAF288w0_0;
	wire w_dff_A_s6veoO8B6_0;
	wire w_dff_A_Ea6N4bL97_0;
	wire w_dff_A_41kHcAp74_2;
	wire w_dff_A_BJkn4WKK8_0;
	wire w_dff_A_t3OCBdPy5_0;
	wire w_dff_A_bNeQcsHg1_0;
	wire w_dff_A_M5pyrNgW0_0;
	wire w_dff_A_HDpeWK6g8_0;
	wire w_dff_A_By0Ov4MX1_2;
	wire w_dff_A_Sp6MW25y5_0;
	wire w_dff_A_t7xpMCTX3_2;
	wire w_dff_A_Y6yi8leE7_0;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(w_dff_A_Xntldy6t4_2),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(w_dff_A_8q4hYZEa0_2),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(w_dff_A_lNIUOv8Z3_2),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_G17gat_2[2]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_n92_0[2]),.dout(w_dff_A_LcBxnPK44_2),.clk(gclk));
	jnot g009(.din(w_n93_0[0]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G1gat_1[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G26gat_0[1]),.dout(n97),.clk(gclk));
	jor g012(.dina(n97),.dinb(w_n96_0[1]),.dout(n98),.clk(gclk));
	jor g013(.dina(w_n98_0[1]),.dinb(n95),.dout(n99),.clk(gclk));
	jor g014(.dina(w_n99_0[1]),.dinb(w_G390gat_0[1]),.dout(w_dff_A_om5yfFJZ9_2),.clk(gclk));
	jnot g015(.din(w_G80gat_0[1]),.dout(n101),.clk(gclk));
	jand g016(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n102),.clk(gclk));
	jnot g017(.din(w_n102_0[1]),.dout(n103),.clk(gclk));
	jor g018(.dina(n103),.dinb(w_n101_0[1]),.dout(w_dff_A_HeZ3jRFr2_2),.clk(gclk));
	jnot g019(.din(w_G36gat_0[0]),.dout(n105),.clk(gclk));
	jnot g020(.din(w_G59gat_1[0]),.dout(n106),.clk(gclk));
	jor g021(.dina(w_n106_0[1]),.dinb(n105),.dout(n107),.clk(gclk));
	jor g022(.dina(w_n107_0[1]),.dinb(w_n101_0[0]),.dout(w_dff_A_fN7Sqhtz9_2),.clk(gclk));
	jnot g023(.din(w_G42gat_1[2]),.dout(n109),.clk(gclk));
	jor g024(.dina(w_n107_0[0]),.dinb(w_dff_B_22qa2mCN4_1),.dout(w_dff_A_HLc1PW0D5_2),.clk(gclk));
	jor g025(.dina(G88gat),.dinb(G87gat),.dout(n111),.clk(gclk));
	jand g026(.dina(w_n111_0[1]),.dinb(w_dff_B_ZJ08p9kY6_1),.dout(w_dff_A_iMewsF9N8_2),.clk(gclk));
	jnot g027(.din(w_G390gat_0[0]),.dout(n113),.clk(gclk));
	jor g028(.dina(w_n99_0[0]),.dinb(n113),.dout(w_dff_A_qRuj8HhM0_2),.clk(gclk));
	jand g029(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n115),.clk(gclk));
	jand g030(.dina(n115),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g031(.dina(w_G55gat_0[2]),.dinb(w_G13gat_0[0]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_n92_0[1]),.dout(n118),.clk(gclk));
	jand g033(.dina(w_G68gat_0[1]),.dinb(w_G29gat_0[0]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_dff_B_ceDN2Djk0_0),.dinb(w_n118_0[2]),.dout(w_dff_A_dO4Fam3e8_2),.clk(gclk));
	jand g035(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n121),.clk(gclk));
	jand g036(.dina(w_n121_0[1]),.dinb(w_dff_B_HgsG02sy0_1),.dout(n122),.clk(gclk));
	jand g037(.dina(n122),.dinb(w_n118_0[1]),.dout(w_dff_A_6MABsAz43_2),.clk(gclk));
	jand g038(.dina(w_n111_0[0]),.dinb(w_dff_B_JnfuJnBI7_1),.dout(w_dff_A_R1GJVanS7_2),.clk(gclk));
	jxor g039(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n125),.clk(gclk));
	jxor g040(.dina(n125),.dinb(w_G130gat_0[1]),.dout(n126),.clk(gclk));
	jxor g041(.dina(w_G126gat_0[1]),.dinb(w_G121gat_0[2]),.dout(n127),.clk(gclk));
	jxor g042(.dina(w_dff_B_d7QAY0mr7_0),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g043(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n129),.clk(gclk));
	jxor g044(.dina(n129),.dinb(w_dff_B_66ClkBp46_1),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(w_dff_B_DkYoUwob4_0),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n128),.dout(w_dff_A_LvQP9xlj5_2),.clk(gclk));
	jxor g048(.dina(w_G165gat_2[1]),.dinb(w_G159gat_2[1]),.dout(n134),.clk(gclk));
	jxor g049(.dina(n134),.dinb(w_G130gat_0[0]),.dout(n135),.clk(gclk));
	jxor g050(.dina(w_G201gat_2[2]),.dinb(w_G195gat_2[1]),.dout(n136),.clk(gclk));
	jxor g051(.dina(w_dff_B_d9aQ3Hsl2_0),.dinb(n135),.dout(n137),.clk(gclk));
	jxor g052(.dina(w_G189gat_2[1]),.dinb(w_G183gat_2[1]),.dout(n138),.clk(gclk));
	jxor g053(.dina(n138),.dinb(w_dff_B_iUY5G3Q84_1),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G177gat_2[1]),.dinb(w_G171gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(w_dff_B_mlTGZ9UB3_0),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n137),.dout(w_dff_A_0r3C9dNv8_2),.clk(gclk));
	jnot g057(.din(w_G261gat_0[2]),.dout(n143),.clk(gclk));
	jand g058(.dina(w_n102_0[0]),.dinb(w_G42gat_1[1]),.dout(n144),.clk(gclk));
	jnot g059(.din(n144),.dout(n145),.clk(gclk));
	jand g060(.dina(w_G51gat_1[0]),.dinb(w_G17gat_2[1]),.dout(n146),.clk(gclk));
	jand g061(.dina(n146),.dinb(w_n92_0[0]),.dout(n147),.clk(gclk));
	jand g062(.dina(w_dff_B_zETTW3TP2_0),.dinb(n145),.dout(n148),.clk(gclk));
	jand g063(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n149),.clk(gclk));
	jxor g064(.dina(w_G42gat_1[0]),.dinb(w_G17gat_2[0]),.dout(n150),.clk(gclk));
	jand g065(.dina(n150),.dinb(w_n149_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(n151),.dinb(w_G447gat_1),.dout(n152),.clk(gclk));
	jor g067(.dina(w_dff_B_udpERRFX2_0),.dinb(n148),.dout(n153),.clk(gclk));
	jand g068(.dina(w_n153_3[1]),.dinb(w_G126gat_0[0]),.dout(n154),.clk(gclk));
	jnot g069(.din(w_G156gat_0[0]),.dout(n155),.clk(gclk));
	jor g070(.dina(n155),.dinb(w_n106_0[0]),.dout(n156),.clk(gclk));
	jand g071(.dina(n156),.dinb(w_G447gat_0[2]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n157_0[1]),.dinb(w_G17gat_1[2]),.dout(n158),.clk(gclk));
	jor g073(.dina(n158),.dinb(w_n96_0[0]),.dout(n159),.clk(gclk));
	jand g074(.dina(w_n159_1[1]),.dinb(w_G153gat_0[2]),.dout(n160),.clk(gclk));
	jand g075(.dina(w_n86_0[0]),.dinb(w_G80gat_0[0]),.dout(n161),.clk(gclk));
	jand g076(.dina(n161),.dinb(w_G447gat_0[1]),.dout(n162),.clk(gclk));
	jnot g077(.din(w_G268gat_0[1]),.dout(n163),.clk(gclk));
	jand g078(.dina(w_n163_0[1]),.dinb(w_G55gat_0[1]),.dout(n164),.clk(gclk));
	jand g079(.dina(w_dff_B_18olbLOP0_0),.dinb(w_n162_0[1]),.dout(n165),.clk(gclk));
	jor g080(.dina(w_n165_1[2]),.dinb(n160),.dout(n166),.clk(gclk));
	jor g081(.dina(n166),.dinb(w_n154_0[1]),.dout(n167),.clk(gclk));
	jxor g082(.dina(w_n167_1[1]),.dinb(w_G201gat_2[1]),.dout(n168),.clk(gclk));
	jnot g083(.din(w_n168_0[2]),.dout(n169),.clk(gclk));
	jor g084(.dina(n169),.dinb(w_n143_0[1]),.dout(n170),.clk(gclk));
	jor g085(.dina(w_n168_0[1]),.dinb(w_G261gat_0[1]),.dout(n171),.clk(gclk));
	jand g086(.dina(n171),.dinb(w_G219gat_3[1]),.dout(n172),.clk(gclk));
	jand g087(.dina(n172),.dinb(n170),.dout(n173),.clk(gclk));
	jand g088(.dina(w_n168_0[0]),.dinb(w_G228gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_G237gat_3[1]),.dinb(w_G201gat_2[0]),.dout(n175),.clk(gclk));
	jor g090(.dina(n175),.dinb(w_G246gat_3[1]),.dout(n176),.clk(gclk));
	jand g091(.dina(w_dff_B_df9p8KhU5_0),.dinb(w_n167_1[0]),.dout(n177),.clk(gclk));
	jand g092(.dina(G72gat),.dinb(w_G42gat_0[2]),.dout(n178),.clk(gclk));
	jand g093(.dina(n178),.dinb(w_dff_B_ewaCWjXU5_1),.dout(n179),.clk(gclk));
	jand g094(.dina(n179),.dinb(w_n121_0[0]),.dout(n180),.clk(gclk));
	jand g095(.dina(n180),.dinb(w_n118_0[0]),.dout(n181),.clk(gclk));
	jand g096(.dina(w_n181_3[1]),.dinb(w_G201gat_1[2]),.dout(n182),.clk(gclk));
	jand g097(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n183),.clk(gclk));
	jand g098(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n184),.clk(gclk));
	jor g099(.dina(n184),.dinb(n183),.dout(n185),.clk(gclk));
	jor g100(.dina(w_dff_B_g769SKK74_0),.dinb(n182),.dout(n186),.clk(gclk));
	jor g101(.dina(w_dff_B_wuapAiYt0_0),.dinb(n177),.dout(n187),.clk(gclk));
	jor g102(.dina(n187),.dinb(n174),.dout(n188),.clk(gclk));
	jor g103(.dina(w_dff_B_eKCnf7nW4_0),.dinb(n173),.dout(w_dff_A_NdwaEkVp4_2),.clk(gclk));
	jand g104(.dina(w_n159_1[0]),.dinb(w_G143gat_0[1]),.dout(n190),.clk(gclk));
	jand g105(.dina(w_n153_3[0]),.dinb(w_G111gat_0[1]),.dout(n191),.clk(gclk));
	jor g106(.dina(n191),.dinb(w_n165_1[1]),.dout(n192),.clk(gclk));
	jor g107(.dina(n192),.dinb(w_dff_B_rOE8WGvz2_1),.dout(n193),.clk(gclk));
	jxor g108(.dina(w_n193_1[1]),.dinb(w_G183gat_2[0]),.dout(n194),.clk(gclk));
	jnot g109(.din(w_n194_0[2]),.dout(n195),.clk(gclk));
	jand g110(.dina(w_n167_0[2]),.dinb(w_G201gat_1[1]),.dout(n196),.clk(gclk));
	jnot g111(.din(w_n196_0[1]),.dout(n197),.clk(gclk));
	jnot g112(.din(w_G201gat_1[0]),.dout(n198),.clk(gclk));
	jnot g113(.din(w_n154_0[0]),.dout(n199),.clk(gclk));
	jnot g114(.din(w_G153gat_0[1]),.dout(n200),.clk(gclk));
	jnot g115(.din(w_G17gat_1[1]),.dout(n201),.clk(gclk));
	jnot g116(.din(w_G51gat_0[2]),.dout(n202),.clk(gclk));
	jor g117(.dina(w_n98_0[0]),.dinb(w_dff_B_a3dEcDtW3_1),.dout(n203),.clk(gclk));
	jor g118(.dina(w_n149_0[0]),.dinb(n203),.dout(n204),.clk(gclk));
	jor g119(.dina(n204),.dinb(w_dff_B_QMDI3G081_1),.dout(n205),.clk(gclk));
	jand g120(.dina(n205),.dinb(w_G1gat_0[1]),.dout(n206),.clk(gclk));
	jor g121(.dina(n206),.dinb(w_dff_B_yTizZ9lw6_1),.dout(n207),.clk(gclk));
	jnot g122(.din(w_n165_1[0]),.dout(n208),.clk(gclk));
	jand g123(.dina(w_dff_B_GxaiRH1j7_0),.dinb(n207),.dout(n209),.clk(gclk));
	jand g124(.dina(n209),.dinb(w_dff_B_LtJRveWy4_1),.dout(n210),.clk(gclk));
	jand g125(.dina(n210),.dinb(w_dff_B_VhjGV70K6_1),.dout(n211),.clk(gclk));
	jor g126(.dina(n211),.dinb(w_n143_0[0]),.dout(n212),.clk(gclk));
	jand g127(.dina(n212),.dinb(w_dff_B_rRFD66SL8_1),.dout(n213),.clk(gclk));
	jand g128(.dina(w_n159_0[2]),.dinb(w_G146gat_0[1]),.dout(n214),.clk(gclk));
	jand g129(.dina(w_n153_2[2]),.dinb(w_G116gat_0[1]),.dout(n215),.clk(gclk));
	jor g130(.dina(n215),.dinb(w_n165_0[2]),.dout(n216),.clk(gclk));
	jor g131(.dina(n216),.dinb(w_dff_B_eenTpDDo4_1),.dout(n217),.clk(gclk));
	jor g132(.dina(w_n217_1[1]),.dinb(w_G189gat_2[0]),.dout(n218),.clk(gclk));
	jand g133(.dina(w_n159_0[1]),.dinb(w_G149gat_0[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n153_2[1]),.dinb(w_G121gat_0[0]),.dout(n220),.clk(gclk));
	jor g135(.dina(n220),.dinb(w_n165_0[1]),.dout(n221),.clk(gclk));
	jor g136(.dina(n221),.dinb(w_dff_B_Y91cRz3S3_1),.dout(n222),.clk(gclk));
	jor g137(.dina(w_n222_1[1]),.dinb(w_G195gat_2[0]),.dout(n223),.clk(gclk));
	jand g138(.dina(w_n223_0[1]),.dinb(w_n218_0[1]),.dout(n224),.clk(gclk));
	jnot g139(.din(w_n224_0[1]),.dout(n225),.clk(gclk));
	jor g140(.dina(w_dff_B_NblQoCvy0_0),.dinb(w_n213_0[1]),.dout(n226),.clk(gclk));
	jand g141(.dina(w_n217_1[0]),.dinb(w_G189gat_1[2]),.dout(n227),.clk(gclk));
	jand g142(.dina(w_n222_1[0]),.dinb(w_G195gat_1[2]),.dout(n228),.clk(gclk));
	jand g143(.dina(w_n228_0[1]),.dinb(w_n218_0[0]),.dout(n229),.clk(gclk));
	jor g144(.dina(n229),.dinb(w_dff_B_oKHxCJyl8_1),.dout(n230),.clk(gclk));
	jnot g145(.din(w_n230_0[1]),.dout(n231),.clk(gclk));
	jand g146(.dina(w_dff_B_AGYNsHQ40_0),.dinb(n226),.dout(n232),.clk(gclk));
	jor g147(.dina(w_n232_0[1]),.dinb(w_dff_B_J7uiEXF66_1),.dout(n233),.clk(gclk));
	jor g148(.dina(w_n167_0[1]),.dinb(w_G201gat_0[2]),.dout(n234),.clk(gclk));
	jand g149(.dina(n234),.dinb(w_G261gat_0[0]),.dout(n235),.clk(gclk));
	jor g150(.dina(n235),.dinb(w_n196_0[0]),.dout(n236),.clk(gclk));
	jand g151(.dina(w_n224_0[0]),.dinb(w_n236_0[2]),.dout(n237),.clk(gclk));
	jor g152(.dina(w_n230_0[0]),.dinb(n237),.dout(n238),.clk(gclk));
	jor g153(.dina(w_n238_0[1]),.dinb(w_n194_0[1]),.dout(n239),.clk(gclk));
	jand g154(.dina(n239),.dinb(w_G219gat_3[0]),.dout(n240),.clk(gclk));
	jand g155(.dina(n240),.dinb(n233),.dout(n241),.clk(gclk));
	jand g156(.dina(w_n194_0[0]),.dinb(w_G228gat_3[0]),.dout(n242),.clk(gclk));
	jand g157(.dina(w_G237gat_3[0]),.dinb(w_G183gat_1[2]),.dout(n243),.clk(gclk));
	jor g158(.dina(n243),.dinb(w_G246gat_3[0]),.dout(n244),.clk(gclk));
	jand g159(.dina(w_dff_B_MxYrP5QC5_0),.dinb(w_n193_1[0]),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n181_3[0]),.dinb(w_G183gat_1[1]),.dout(n246),.clk(gclk));
	jand g161(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n247),.clk(gclk));
	jor g162(.dina(w_dff_B_gR5RYfHF0_0),.dinb(n246),.dout(n248),.clk(gclk));
	jor g163(.dina(w_dff_B_zwv9qhOX5_0),.dinb(n245),.dout(n249),.clk(gclk));
	jor g164(.dina(n249),.dinb(n242),.dout(n250),.clk(gclk));
	jor g165(.dina(w_dff_B_MFvsdWBy7_0),.dinb(n241),.dout(w_dff_A_TtRDAdvq8_2),.clk(gclk));
	jxor g166(.dina(w_n217_0[2]),.dinb(w_G189gat_1[1]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n252_0[2]),.dout(n253),.clk(gclk));
	jand g168(.dina(w_n223_0[0]),.dinb(w_n236_0[1]),.dout(n254),.clk(gclk));
	jor g169(.dina(n254),.dinb(w_n228_0[0]),.dout(n255),.clk(gclk));
	jnot g170(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jor g171(.dina(n256),.dinb(w_dff_B_C5AC7Cip1_1),.dout(n257),.clk(gclk));
	jor g172(.dina(w_n255_0[0]),.dinb(w_n252_0[1]),.dout(n258),.clk(gclk));
	jand g173(.dina(n258),.dinb(w_G219gat_2[2]),.dout(n259),.clk(gclk));
	jand g174(.dina(n259),.dinb(n257),.dout(n260),.clk(gclk));
	jand g175(.dina(w_n252_0[0]),.dinb(w_G228gat_2[2]),.dout(n261),.clk(gclk));
	jand g176(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n262),.clk(gclk));
	jor g177(.dina(n262),.dinb(w_G246gat_2[2]),.dout(n263),.clk(gclk));
	jand g178(.dina(w_dff_B_iKCGrPsq2_0),.dinb(w_n217_0[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(w_n181_2[2]),.dinb(w_G189gat_0[2]),.dout(n265),.clk(gclk));
	jand g180(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n266),.clk(gclk));
	jand g181(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n267),.clk(gclk));
	jor g182(.dina(n267),.dinb(n266),.dout(n268),.clk(gclk));
	jor g183(.dina(w_dff_B_gKnj4rBG1_0),.dinb(n265),.dout(n269),.clk(gclk));
	jor g184(.dina(w_dff_B_IfB1r0h09_0),.dinb(n264),.dout(n270),.clk(gclk));
	jor g185(.dina(n270),.dinb(n261),.dout(n271),.clk(gclk));
	jor g186(.dina(w_dff_B_ZKSjb0ht7_0),.dinb(n260),.dout(w_dff_A_rFZzsmmR5_2),.clk(gclk));
	jxor g187(.dina(w_n222_0[2]),.dinb(w_G195gat_1[1]),.dout(n273),.clk(gclk));
	jnot g188(.din(w_n273_0[2]),.dout(n274),.clk(gclk));
	jor g189(.dina(w_dff_B_eUvIE2o32_0),.dinb(w_n213_0[0]),.dout(n275),.clk(gclk));
	jor g190(.dina(w_n273_0[1]),.dinb(w_n236_0[0]),.dout(n276),.clk(gclk));
	jand g191(.dina(n276),.dinb(w_G219gat_2[1]),.dout(n277),.clk(gclk));
	jand g192(.dina(n277),.dinb(n275),.dout(n278),.clk(gclk));
	jand g193(.dina(w_n273_0[0]),.dinb(w_G228gat_2[1]),.dout(n279),.clk(gclk));
	jand g194(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n280),.clk(gclk));
	jor g195(.dina(n280),.dinb(w_G246gat_2[1]),.dout(n281),.clk(gclk));
	jand g196(.dina(w_dff_B_hIcihech9_0),.dinb(w_n222_0[1]),.dout(n282),.clk(gclk));
	jand g197(.dina(w_n181_2[1]),.dinb(w_G195gat_0[2]),.dout(n283),.clk(gclk));
	jand g198(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n284),.clk(gclk));
	jand g199(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n285),.clk(gclk));
	jor g200(.dina(n285),.dinb(n284),.dout(n286),.clk(gclk));
	jor g201(.dina(w_dff_B_ccXQruad6_0),.dinb(n283),.dout(n287),.clk(gclk));
	jor g202(.dina(w_dff_B_sDU7CWKL3_0),.dinb(n282),.dout(n288),.clk(gclk));
	jor g203(.dina(n288),.dinb(n279),.dout(n289),.clk(gclk));
	jor g204(.dina(w_dff_B_KbnTInxV4_0),.dinb(n278),.dout(w_dff_A_41kHcAp74_2),.clk(gclk));
	jand g205(.dina(w_n153_2[0]),.dinb(w_G91gat_0[1]),.dout(n291),.clk(gclk));
	jand g206(.dina(w_n157_0[0]),.dinb(w_G55gat_0[0]),.dout(n292),.clk(gclk));
	jand g207(.dina(w_n292_1[1]),.dinb(w_G143gat_0[0]),.dout(n293),.clk(gclk));
	jand g208(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n294),.clk(gclk));
	jand g209(.dina(w_n163_0[0]),.dinb(w_G17gat_1[0]),.dout(n295),.clk(gclk));
	jand g210(.dina(w_dff_B_jjjjMfHr1_0),.dinb(w_n162_0[0]),.dout(n296),.clk(gclk));
	jor g211(.dina(w_n296_1[1]),.dinb(w_dff_B_zCnyp4Y35_1),.dout(n297),.clk(gclk));
	jor g212(.dina(n297),.dinb(n293),.dout(n298),.clk(gclk));
	jor g213(.dina(n298),.dinb(n291),.dout(n299),.clk(gclk));
	jand g214(.dina(w_n299_1[1]),.dinb(w_G159gat_2[0]),.dout(n300),.clk(gclk));
	jor g215(.dina(w_n299_1[0]),.dinb(w_G159gat_1[2]),.dout(n301),.clk(gclk));
	jand g216(.dina(w_n193_0[2]),.dinb(w_G183gat_1[0]),.dout(n302),.clk(gclk));
	jor g217(.dina(w_n193_0[1]),.dinb(w_G183gat_0[2]),.dout(n303),.clk(gclk));
	jand g218(.dina(w_n238_0[0]),.dinb(w_n303_0[1]),.dout(n304),.clk(gclk));
	jor g219(.dina(n304),.dinb(w_n302_0[1]),.dout(n305),.clk(gclk));
	jnot g220(.din(w_G165gat_2[0]),.dout(n306),.clk(gclk));
	jand g221(.dina(w_n153_1[2]),.dinb(w_G96gat_0[1]),.dout(n307),.clk(gclk));
	jand g222(.dina(w_n292_1[0]),.dinb(w_G146gat_0[0]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n309),.clk(gclk));
	jor g224(.dina(w_dff_B_vydm3phq2_0),.dinb(w_n296_1[0]),.dout(n310),.clk(gclk));
	jor g225(.dina(n310),.dinb(n308),.dout(n311),.clk(gclk));
	jor g226(.dina(n311),.dinb(n307),.dout(n312),.clk(gclk));
	jnot g227(.din(w_n312_1[1]),.dout(n313),.clk(gclk));
	jand g228(.dina(n313),.dinb(w_dff_B_kHduTWwA0_1),.dout(n314),.clk(gclk));
	jnot g229(.din(n314),.dout(n315),.clk(gclk));
	jand g230(.dina(w_n153_1[1]),.dinb(w_G101gat_0[1]),.dout(n316),.clk(gclk));
	jand g231(.dina(w_n292_0[2]),.dinb(w_G149gat_0[0]),.dout(n317),.clk(gclk));
	jand g232(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n318),.clk(gclk));
	jor g233(.dina(w_dff_B_rzvQ8ikQ1_0),.dinb(w_n296_0[2]),.dout(n319),.clk(gclk));
	jor g234(.dina(n319),.dinb(n317),.dout(n320),.clk(gclk));
	jor g235(.dina(n320),.dinb(n316),.dout(n321),.clk(gclk));
	jor g236(.dina(w_n321_1[1]),.dinb(w_G171gat_2[0]),.dout(n322),.clk(gclk));
	jand g237(.dina(w_n153_1[0]),.dinb(w_G106gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_n292_0[1]),.dinb(w_G153gat_0[0]),.dout(n324),.clk(gclk));
	jand g239(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n325),.clk(gclk));
	jor g240(.dina(w_dff_B_fkJQA9hn5_0),.dinb(w_n296_0[1]),.dout(n326),.clk(gclk));
	jor g241(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jor g242(.dina(n327),.dinb(n323),.dout(n328),.clk(gclk));
	jor g243(.dina(w_n328_1[1]),.dinb(w_G177gat_2[0]),.dout(n329),.clk(gclk));
	jand g244(.dina(w_n329_0[2]),.dinb(w_n322_0[1]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n330_0[2]),.dinb(w_n315_0[1]),.dout(n331),.clk(gclk));
	jand g246(.dina(w_n331_0[1]),.dinb(w_n305_1[1]),.dout(n332),.clk(gclk));
	jand g247(.dina(w_n312_1[0]),.dinb(w_G165gat_1[2]),.dout(n333),.clk(gclk));
	jand g248(.dina(w_n321_1[0]),.dinb(w_G171gat_1[2]),.dout(n334),.clk(gclk));
	jand g249(.dina(w_n328_1[0]),.dinb(w_G177gat_1[2]),.dout(n335),.clk(gclk));
	jand g250(.dina(w_n335_0[2]),.dinb(w_n322_0[0]),.dout(n336),.clk(gclk));
	jor g251(.dina(n336),.dinb(w_dff_B_oNIztZJx2_1),.dout(n337),.clk(gclk));
	jand g252(.dina(w_n337_0[2]),.dinb(w_n315_0[0]),.dout(n338),.clk(gclk));
	jor g253(.dina(n338),.dinb(w_dff_B_53ySjMjh9_1),.dout(n339),.clk(gclk));
	jor g254(.dina(w_n339_0[1]),.dinb(n332),.dout(n340),.clk(gclk));
	jand g255(.dina(w_n340_0[1]),.dinb(w_dff_B_9x4JXOZc9_1),.dout(n341),.clk(gclk));
	jor g256(.dina(n341),.dinb(w_dff_B_drA7A5wC2_1),.dout(w_dff_A_By0Ov4MX1_2),.clk(gclk));
	jnot g257(.din(w_n302_0[0]),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n303_0[0]),.dout(n344),.clk(gclk));
	jor g259(.dina(w_n232_0[0]),.dinb(w_dff_B_VkeglazP1_1),.dout(n345),.clk(gclk));
	jand g260(.dina(n345),.dinb(w_dff_B_TXmJT4UW2_1),.dout(n346),.clk(gclk));
	jxor g261(.dina(w_n328_0[2]),.dinb(w_G177gat_1[1]),.dout(n347),.clk(gclk));
	jnot g262(.din(w_n347_0[2]),.dout(n348),.clk(gclk));
	jor g263(.dina(w_dff_B_44poXEwj6_0),.dinb(w_n346_1[1]),.dout(n349),.clk(gclk));
	jor g264(.dina(w_n347_0[1]),.dinb(w_n305_1[0]),.dout(n350),.clk(gclk));
	jand g265(.dina(n350),.dinb(w_G219gat_2[0]),.dout(n351),.clk(gclk));
	jand g266(.dina(n351),.dinb(n349),.dout(n352),.clk(gclk));
	jand g267(.dina(w_n347_0[0]),.dinb(w_G228gat_2[0]),.dout(n353),.clk(gclk));
	jand g268(.dina(w_G237gat_2[0]),.dinb(w_G177gat_1[0]),.dout(n354),.clk(gclk));
	jor g269(.dina(n354),.dinb(w_G246gat_2[0]),.dout(n355),.clk(gclk));
	jand g270(.dina(w_dff_B_58zR0n3s1_0),.dinb(w_n328_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n181_2[0]),.dinb(w_G177gat_0[2]),.dout(n357),.clk(gclk));
	jand g272(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n358),.clk(gclk));
	jor g273(.dina(w_dff_B_1iohtdfD7_0),.dinb(n357),.dout(n359),.clk(gclk));
	jor g274(.dina(w_dff_B_lE9VLwQq3_0),.dinb(n356),.dout(n360),.clk(gclk));
	jor g275(.dina(n360),.dinb(n353),.dout(n361),.clk(gclk));
	jor g276(.dina(w_dff_B_ZvgTSLK49_0),.dinb(n352),.dout(w_dff_A_t7xpMCTX3_2),.clk(gclk));
	jnot g277(.din(w_n331_0[0]),.dout(n363),.clk(gclk));
	jor g278(.dina(w_dff_B_mmHNanG33_0),.dinb(w_n346_1[0]),.dout(n364),.clk(gclk));
	jnot g279(.din(w_n339_0[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_dff_B_qWOZGGdK5_0),.dinb(n364),.dout(n366),.clk(gclk));
	jxor g281(.dina(w_n299_0[2]),.dinb(w_G159gat_1[1]),.dout(n367),.clk(gclk));
	jnot g282(.din(w_n367_0[2]),.dout(n368),.clk(gclk));
	jor g283(.dina(w_dff_B_sABVbcuN3_0),.dinb(n366),.dout(n369),.clk(gclk));
	jor g284(.dina(w_n367_0[1]),.dinb(w_n340_0[0]),.dout(n370),.clk(gclk));
	jand g285(.dina(n370),.dinb(w_G219gat_1[2]),.dout(n371),.clk(gclk));
	jand g286(.dina(n371),.dinb(n369),.dout(n372),.clk(gclk));
	jand g287(.dina(w_n367_0[0]),.dinb(w_G228gat_1[2]),.dout(n373),.clk(gclk));
	jand g288(.dina(w_G237gat_1[2]),.dinb(w_G159gat_1[0]),.dout(n374),.clk(gclk));
	jor g289(.dina(n374),.dinb(w_G246gat_1[2]),.dout(n375),.clk(gclk));
	jand g290(.dina(w_dff_B_Htl8yZ1Z7_0),.dinb(w_n299_0[1]),.dout(n376),.clk(gclk));
	jand g291(.dina(w_n181_1[2]),.dinb(w_G159gat_0[2]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n378),.clk(gclk));
	jor g293(.dina(w_dff_B_Ez5N4pDZ5_0),.dinb(n377),.dout(n379),.clk(gclk));
	jor g294(.dina(w_dff_B_HzuYTE3n4_0),.dinb(n376),.dout(n380),.clk(gclk));
	jor g295(.dina(n380),.dinb(n373),.dout(n381),.clk(gclk));
	jor g296(.dina(w_dff_B_hfzIin7F9_0),.dinb(n372),.dout(G878gat),.clk(gclk));
	jxor g297(.dina(w_n312_0[2]),.dinb(w_G165gat_1[1]),.dout(n383),.clk(gclk));
	jnot g298(.din(w_n383_0[2]),.dout(n384),.clk(gclk));
	jnot g299(.din(w_n337_0[1]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n330_0[1]),.dout(n386),.clk(gclk));
	jor g301(.dina(w_dff_B_uubzqeWb6_0),.dinb(w_n346_0[2]),.dout(n387),.clk(gclk));
	jand g302(.dina(n387),.dinb(w_dff_B_LMygMd880_1),.dout(n388),.clk(gclk));
	jor g303(.dina(n388),.dinb(w_dff_B_2sqQBAbT8_1),.dout(n389),.clk(gclk));
	jand g304(.dina(w_n330_0[0]),.dinb(w_n305_0[2]),.dout(n390),.clk(gclk));
	jor g305(.dina(n390),.dinb(w_n337_0[0]),.dout(n391),.clk(gclk));
	jor g306(.dina(n391),.dinb(w_n383_0[1]),.dout(n392),.clk(gclk));
	jand g307(.dina(n392),.dinb(w_G219gat_1[1]),.dout(n393),.clk(gclk));
	jand g308(.dina(n393),.dinb(n389),.dout(n394),.clk(gclk));
	jand g309(.dina(w_n383_0[0]),.dinb(w_G228gat_1[1]),.dout(n395),.clk(gclk));
	jand g310(.dina(w_G237gat_1[1]),.dinb(w_G165gat_1[0]),.dout(n396),.clk(gclk));
	jor g311(.dina(n396),.dinb(w_G246gat_1[1]),.dout(n397),.clk(gclk));
	jand g312(.dina(w_dff_B_3oznaR7T2_0),.dinb(w_n312_0[1]),.dout(n398),.clk(gclk));
	jand g313(.dina(w_n181_1[1]),.dinb(w_G165gat_0[2]),.dout(n399),.clk(gclk));
	jand g314(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n400),.clk(gclk));
	jor g315(.dina(w_dff_B_cWMBAM437_0),.dinb(n399),.dout(n401),.clk(gclk));
	jor g316(.dina(w_dff_B_WsR0QEeq2_0),.dinb(n398),.dout(n402),.clk(gclk));
	jor g317(.dina(n402),.dinb(n395),.dout(n403),.clk(gclk));
	jor g318(.dina(w_dff_B_MStUdTdf6_0),.dinb(n394),.dout(G879gat),.clk(gclk));
	jxor g319(.dina(w_n321_0[2]),.dinb(w_G171gat_1[1]),.dout(n405),.clk(gclk));
	jnot g320(.din(w_n405_0[2]),.dout(n406),.clk(gclk));
	jnot g321(.din(w_n335_0[1]),.dout(n407),.clk(gclk));
	jnot g322(.din(w_n329_0[1]),.dout(n408),.clk(gclk));
	jor g323(.dina(w_dff_B_Zzqx5ko26_0),.dinb(w_n346_0[1]),.dout(n409),.clk(gclk));
	jand g324(.dina(n409),.dinb(w_dff_B_2iVXjyDC6_1),.dout(n410),.clk(gclk));
	jor g325(.dina(n410),.dinb(w_dff_B_zJD5ybiD5_1),.dout(n411),.clk(gclk));
	jand g326(.dina(w_n329_0[0]),.dinb(w_n305_0[1]),.dout(n412),.clk(gclk));
	jor g327(.dina(n412),.dinb(w_n335_0[0]),.dout(n413),.clk(gclk));
	jor g328(.dina(n413),.dinb(w_n405_0[1]),.dout(n414),.clk(gclk));
	jand g329(.dina(n414),.dinb(w_G219gat_1[0]),.dout(n415),.clk(gclk));
	jand g330(.dina(n415),.dinb(n411),.dout(n416),.clk(gclk));
	jand g331(.dina(w_n405_0[0]),.dinb(w_G228gat_1[0]),.dout(n417),.clk(gclk));
	jand g332(.dina(w_G237gat_1[0]),.dinb(w_G171gat_1[0]),.dout(n418),.clk(gclk));
	jor g333(.dina(n418),.dinb(w_G246gat_1[0]),.dout(n419),.clk(gclk));
	jand g334(.dina(w_dff_B_WmH6Gm1u3_0),.dinb(w_n321_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n181_1[0]),.dinb(w_G171gat_0[2]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jor g337(.dina(w_dff_B_c16ODci74_0),.dinb(n421),.dout(n423),.clk(gclk));
	jor g338(.dina(w_dff_B_Q750Mzc63_0),.dinb(n420),.dout(n424),.clk(gclk));
	jor g339(.dina(n424),.dinb(n417),.dout(n425),.clk(gclk));
	jor g340(.dina(w_dff_B_WOXq1yvj3_0),.dinb(n416),.dout(G880gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_dff_A_Mjm2LAJE6_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_G13gat_0[1]),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_dff_A_jI7X4yov3_0),.doutb(w_G17gat_1[1]),.doutc(w_dff_A_Om4YmTQj9_2),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_G17gat_2[2]),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_G29gat_0[0]),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_dff_A_w0p67XqF8_1),.doutc(w_G42gat_0[2]),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_G42gat_1[0]),.doutb(w_dff_A_PGiJWcjm6_1),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_dff_A_wQHYWXrg3_1),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_dff_A_nCZDJcW77_0),.doutb(w_dff_A_Xxz2xkIl5_1),.doutc(w_G55gat_0[2]),.din(G55gat));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_G68gat_0[1]),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_dff_A_meywaUyO7_0),.doutb(w_G80gat_0[1]),.doutc(w_dff_A_VxBXljXt1_2),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_dff_A_bvAjlEZl6_1),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_dff_A_iJQF7wRB4_1),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_dff_A_YRAMphzX3_1),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_J5Vh6mSc0_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_dff_A_qrJOZv860_1),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_dff_A_s4lNmvvS8_1),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_dff_A_IsZfT29g9_0),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl jspl_w_G126gat_0(.douta(w_dff_A_kj7LiY6u0_0),.doutb(w_G126gat_0[1]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_G130gat_0[1]),.din(w_dff_B_978t756o8_2));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_dff_A_mLdU7aep6_1),.din(w_dff_B_B0ihQo9d3_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_dff_A_Utnvb7700_1),.din(w_dff_B_RUCXEpUo8_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_dff_A_4JNFA8PX0_1),.din(w_dff_B_OZVGGOE57_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_dff_A_ehEewFN31_0),.doutb(w_G153gat_0[1]),.doutc(w_dff_A_x5CwquCG5_2),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_G159gat_0[1]),.doutc(w_dff_A_eE0L9O3I9_2),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_G159gat_1[0]),.doutb(w_dff_A_b8BjMrtc1_1),.doutc(w_dff_A_IeRBU1Vr6_2),.din(w_G159gat_0[0]));
	jspl jspl_w_G159gat_2(.douta(w_dff_A_T5wby41Q7_0),.doutb(w_G159gat_2[1]),.din(w_G159gat_0[1]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_G165gat_0[1]),.doutc(w_dff_A_JxVtyyyi3_2),.din(G165gat));
	jspl3 jspl3_w_G165gat_1(.douta(w_G165gat_1[0]),.doutb(w_dff_A_aUqhprmc4_1),.doutc(w_dff_A_7TkqrJOl2_2),.din(w_G165gat_0[0]));
	jspl jspl_w_G165gat_2(.douta(w_G165gat_2[0]),.doutb(w_G165gat_2[1]),.din(w_G165gat_0[1]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_dff_A_rs2z8Iys3_2),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_dff_A_PSEKKTS35_1),.doutc(w_dff_A_GlMLFNvK1_2),.din(w_G171gat_0[0]));
	jspl jspl_w_G171gat_2(.douta(w_dff_A_tZ4AwOED6_0),.doutb(w_G171gat_2[1]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_G177gat_0[1]),.doutc(w_dff_A_Hpxb2jRc1_2),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_dff_A_6sPlPBXq0_1),.doutc(w_dff_A_VvwERKv35_2),.din(w_G177gat_0[0]));
	jspl jspl_w_G177gat_2(.douta(w_dff_A_PTCrlAKa4_0),.doutb(w_G177gat_2[1]),.din(w_G177gat_0[1]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_dff_A_Wr5l3qB80_2),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_dff_A_KKyrQJND4_0),.doutb(w_dff_A_1QSSEYiG4_1),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl jspl_w_G183gat_2(.douta(w_dff_A_yvRtKMeT2_0),.doutb(w_G183gat_2[1]),.din(w_G183gat_0[1]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_dff_A_PhIG9if66_2),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_dff_A_5UNrjDdz5_1),.doutc(w_dff_A_wLIgF7JD4_2),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_dff_A_F0P8hhOf4_0),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_dff_A_8fG1lPkj0_2),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_dff_A_2cjpNXO87_1),.doutc(w_dff_A_Tk84Qdly2_2),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_dff_A_XMcUX3AP0_0),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_G201gat_0[1]),.doutc(w_dff_A_pdf0eo104_2),.din(G201gat));
	jspl3 jspl3_w_G201gat_1(.douta(w_G201gat_1[0]),.doutb(w_dff_A_zEIzOYzO8_1),.doutc(w_dff_A_L2PRPBEx7_2),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G201gat_2(.douta(w_G201gat_2[0]),.doutb(w_dff_A_AN8Xwk1H3_1),.doutc(w_G201gat_2[2]),.din(w_G201gat_0[1]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_TFGMO4fp7_0),.doutb(w_dff_A_m7XBoiE86_1),.doutc(w_G219gat_0[2]),.din(w_dff_B_z2BH0hU70_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_G219gat_1[0]),.doutb(w_G219gat_1[1]),.doutc(w_G219gat_1[2]),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_10DzDZaA4_0),.doutb(w_G219gat_2[1]),.doutc(w_dff_A_qRXtUuAr5_2),.din(w_G219gat_0[1]));
	jspl jspl_w_G219gat_3(.douta(w_dff_A_EJDOXZUE8_0),.doutb(w_G219gat_3[1]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_G228gat_0[0]),.doutb(w_G228gat_0[1]),.doutc(w_dff_A_0DXRBDIX9_2),.din(w_dff_B_UjLH3mI44_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_G228gat_2[0]),.doutb(w_dff_A_iFem6Mhk9_1),.doutc(w_dff_A_1u7JjUPF2_2),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_G228gat_3[1]),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_G237gat_0[0]),.doutb(w_G237gat_0[1]),.doutc(w_G237gat_0[2]),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_G237gat_2[0]),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_G237gat_3[1]),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_G246gat_0[0]),.doutb(w_G246gat_0[1]),.doutc(w_G246gat_0[2]),.din(w_dff_B_P18D2B739_3));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_G246gat_2[0]),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_G246gat_3[1]),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_dff_A_olrTfMMo1_0),.doutb(w_dff_A_VDf97yrT4_1),.doutc(w_G261gat_0[2]),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_dff_A_5uYtbCG08_1),.doutc(w_dff_A_LZkuzL3R5_2),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_G447gat_0[2]),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(w_dff_A_4xqBO2HF8_1),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n96_0(.douta(w_dff_A_P9EaKFnE3_0),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(w_dff_B_BU45obMx4_2));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl jspl_w_n106_0(.douta(w_n106_0[0]),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n118_0(.douta(w_dff_A_RaHkYuxw1_0),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl jspl_w_n121_0(.douta(w_dff_A_ziZeDzT31_0),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(w_dff_B_Ef3RQZoT8_2));
	jspl jspl_w_n149_0(.douta(w_dff_A_tixy5xj33_0),.doutb(w_n149_0[1]),.din(n149));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.doutc(w_n153_1[2]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n153_2(.douta(w_n153_2[0]),.doutb(w_n153_2[1]),.doutc(w_n153_2[2]),.din(w_n153_0[1]));
	jspl jspl_w_n153_3(.douta(w_n153_3[0]),.doutb(w_n153_3[1]),.din(w_n153_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_dff_A_MeVNwU9y6_1),.din(n154));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_TypNUBOb1_1),.doutc(w_dff_A_OdzPs9rg2_2),.din(n165));
	jspl3 jspl3_w_n165_1(.douta(w_n165_1[0]),.doutb(w_dff_A_wJXMRtTS0_1),.doutc(w_dff_A_yK5wcWlf3_2),.din(w_n165_0[0]));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.doutc(w_n167_0[2]),.din(n167));
	jspl jspl_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n181_2(.douta(w_n181_2[0]),.doutb(w_n181_2[1]),.doutc(w_n181_2[2]),.din(w_n181_0[1]));
	jspl jspl_w_n181_3(.douta(w_n181_3[0]),.doutb(w_n181_3[1]),.din(w_n181_0[2]));
	jspl3 jspl3_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.doutc(w_n193_0[2]),.din(n193));
	jspl jspl_w_n193_1(.douta(w_n193_1[0]),.doutb(w_n193_1[1]),.din(w_n193_0[0]));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_dff_A_mVPNFlTl0_1),.doutc(w_n194_0[2]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_dff_A_djOBsNTk8_0),.doutb(w_n196_0[1]),.din(n196));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl jspl_w_n217_1(.douta(w_n217_1[0]),.doutb(w_n217_1[1]),.din(w_n217_0[0]));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.doutc(w_n222_0[2]),.din(n222));
	jspl jspl_w_n222_1(.douta(w_n222_1[0]),.doutb(w_n222_1[1]),.din(w_n222_0[0]));
	jspl jspl_w_n223_0(.douta(w_dff_A_xsDiUmav4_0),.doutb(w_n223_0[1]),.din(n223));
	jspl jspl_w_n224_0(.douta(w_dff_A_P4A3xGbv7_0),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n228_0(.douta(w_dff_A_9Lkwfsre6_0),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_dff_A_QY1RKPjN8_0),.doutb(w_n230_0[1]),.din(n230));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.doutc(w_n236_0[2]),.din(n236));
	jspl jspl_w_n238_0(.douta(w_n238_0[0]),.doutb(w_n238_0[1]),.din(n238));
	jspl3 jspl3_w_n252_0(.douta(w_n252_0[0]),.doutb(w_dff_A_IySSeJOx0_1),.doutc(w_n252_0[2]),.din(n252));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_dff_A_DizNzasm0_1),.doutc(w_n273_0[2]),.din(n273));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl jspl_w_n292_1(.douta(w_n292_1[0]),.doutb(w_n292_1[1]),.din(w_n292_0[0]));
	jspl3 jspl3_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.doutc(w_n296_0[2]),.din(n296));
	jspl jspl_w_n296_1(.douta(w_n296_1[0]),.doutb(w_n296_1[1]),.din(w_n296_0[0]));
	jspl3 jspl3_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.doutc(w_n299_0[2]),.din(n299));
	jspl jspl_w_n299_1(.douta(w_n299_1[0]),.doutb(w_n299_1[1]),.din(w_n299_0[0]));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_dff_A_BCpoGdPS7_1),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_YURtj78C0_1),.din(n303));
	jspl3 jspl3_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.doutc(w_n305_0[2]),.din(n305));
	jspl jspl_w_n305_1(.douta(w_n305_1[0]),.doutb(w_n305_1[1]),.din(w_n305_0[0]));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl3 jspl3_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.doutc(w_n321_0[2]),.din(n321));
	jspl jspl_w_n321_1(.douta(w_n321_1[0]),.doutb(w_n321_1[1]),.din(w_n321_0[0]));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n328_1(.douta(w_n328_1[0]),.doutb(w_n328_1[1]),.din(w_n328_0[0]));
	jspl3 jspl3_w_n329_0(.douta(w_dff_A_VNpFfYvM2_0),.doutb(w_n329_0[1]),.doutc(w_n329_0[2]),.din(n329));
	jspl3 jspl3_w_n330_0(.douta(w_dff_A_qQw0GRV41_0),.doutb(w_n330_0[1]),.doutc(w_dff_A_DhhcOSpl4_2),.din(n330));
	jspl jspl_w_n331_0(.douta(w_n331_0[0]),.doutb(w_dff_A_pWXqXzVN4_1),.din(n331));
	jspl3 jspl3_w_n335_0(.douta(w_dff_A_wYIkLhg66_0),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n337_0(.douta(w_dff_A_pRnFC8hN5_0),.doutb(w_n337_0[1]),.doutc(w_n337_0[2]),.din(n337));
	jspl jspl_w_n339_0(.douta(w_n339_0[0]),.doutb(w_dff_A_bPtpMy9K0_1),.din(n339));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n347_0(.douta(w_n347_0[0]),.doutb(w_dff_A_382X31nZ2_1),.doutc(w_n347_0[2]),.din(n347));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_dff_A_kV4L7Rfy6_1),.doutc(w_n367_0[2]),.din(n367));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_dff_A_sx4S7KWf4_1),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_dff_A_ndz4jTRC8_1),.doutc(w_n405_0[2]),.din(n405));
	jdff dff_B_BU45obMx4_2(.din(n101),.dout(w_dff_B_BU45obMx4_2),.clk(gclk));
	jdff dff_B_22qa2mCN4_1(.din(n109),.dout(w_dff_B_22qa2mCN4_1),.clk(gclk));
	jdff dff_B_ZJ08p9kY6_1(.din(G90gat),.dout(w_dff_B_ZJ08p9kY6_1),.clk(gclk));
	jdff dff_A_5uYtbCG08_1(.dout(w_G390gat_0[1]),.din(w_dff_A_5uYtbCG08_1),.clk(gclk));
	jdff dff_B_ceDN2Djk0_0(.din(n119),.dout(w_dff_B_ceDN2Djk0_0),.clk(gclk));
	jdff dff_B_HgsG02sy0_1(.din(G74gat),.dout(w_dff_B_HgsG02sy0_1),.clk(gclk));
	jdff dff_B_JnfuJnBI7_1(.din(G89gat),.dout(w_dff_B_JnfuJnBI7_1),.clk(gclk));
	jdff dff_B_DkYoUwob4_0(.din(n131),.dout(w_dff_B_DkYoUwob4_0),.clk(gclk));
	jdff dff_B_66ClkBp46_1(.din(G135gat),.dout(w_dff_B_66ClkBp46_1),.clk(gclk));
	jdff dff_B_d7QAY0mr7_0(.din(n127),.dout(w_dff_B_d7QAY0mr7_0),.clk(gclk));
	jdff dff_B_mlTGZ9UB3_0(.din(n140),.dout(w_dff_B_mlTGZ9UB3_0),.clk(gclk));
	jdff dff_B_iUY5G3Q84_1(.din(G207gat),.dout(w_dff_B_iUY5G3Q84_1),.clk(gclk));
	jdff dff_B_d9aQ3Hsl2_0(.din(n136),.dout(w_dff_B_d9aQ3Hsl2_0),.clk(gclk));
	jdff dff_B_978t756o8_2(.din(G130gat),.dout(w_dff_B_978t756o8_2),.clk(gclk));
	jdff dff_B_eKCnf7nW4_0(.din(n188),.dout(w_dff_B_eKCnf7nW4_0),.clk(gclk));
	jdff dff_B_23MZzeTv0_0(.din(n186),.dout(w_dff_B_23MZzeTv0_0),.clk(gclk));
	jdff dff_B_pPDGf0V36_0(.din(w_dff_B_23MZzeTv0_0),.dout(w_dff_B_pPDGf0V36_0),.clk(gclk));
	jdff dff_B_wuapAiYt0_0(.din(w_dff_B_pPDGf0V36_0),.dout(w_dff_B_wuapAiYt0_0),.clk(gclk));
	jdff dff_B_ylPBW2Nm7_0(.din(n185),.dout(w_dff_B_ylPBW2Nm7_0),.clk(gclk));
	jdff dff_B_35T3dBtB9_0(.din(w_dff_B_ylPBW2Nm7_0),.dout(w_dff_B_35T3dBtB9_0),.clk(gclk));
	jdff dff_B_g769SKK74_0(.din(w_dff_B_35T3dBtB9_0),.dout(w_dff_B_g769SKK74_0),.clk(gclk));
	jdff dff_B_AVY1b9U14_0(.din(n176),.dout(w_dff_B_AVY1b9U14_0),.clk(gclk));
	jdff dff_B_uM2M20Dq5_0(.din(w_dff_B_AVY1b9U14_0),.dout(w_dff_B_uM2M20Dq5_0),.clk(gclk));
	jdff dff_B_5aExwmzQ1_0(.din(w_dff_B_uM2M20Dq5_0),.dout(w_dff_B_5aExwmzQ1_0),.clk(gclk));
	jdff dff_B_MnkDCOT22_0(.din(w_dff_B_5aExwmzQ1_0),.dout(w_dff_B_MnkDCOT22_0),.clk(gclk));
	jdff dff_B_D401LXRg8_0(.din(w_dff_B_MnkDCOT22_0),.dout(w_dff_B_D401LXRg8_0),.clk(gclk));
	jdff dff_B_df9p8KhU5_0(.din(w_dff_B_D401LXRg8_0),.dout(w_dff_B_df9p8KhU5_0),.clk(gclk));
	jdff dff_A_wvNXrZLk3_1(.dout(w_G201gat_2[1]),.din(w_dff_A_wvNXrZLk3_1),.clk(gclk));
	jdff dff_A_a7Hqmr399_1(.dout(w_dff_A_wvNXrZLk3_1),.din(w_dff_A_a7Hqmr399_1),.clk(gclk));
	jdff dff_A_HA6vdDli5_1(.dout(w_dff_A_a7Hqmr399_1),.din(w_dff_A_HA6vdDli5_1),.clk(gclk));
	jdff dff_A_Eocuhlud6_1(.dout(w_dff_A_HA6vdDli5_1),.din(w_dff_A_Eocuhlud6_1),.clk(gclk));
	jdff dff_A_thWiTtzF7_1(.dout(w_dff_A_Eocuhlud6_1),.din(w_dff_A_thWiTtzF7_1),.clk(gclk));
	jdff dff_A_smmUMEVX2_1(.dout(w_dff_A_thWiTtzF7_1),.din(w_dff_A_smmUMEVX2_1),.clk(gclk));
	jdff dff_A_MD05oMil1_1(.dout(w_dff_A_smmUMEVX2_1),.din(w_dff_A_MD05oMil1_1),.clk(gclk));
	jdff dff_A_AN8Xwk1H3_1(.dout(w_dff_A_MD05oMil1_1),.din(w_dff_A_AN8Xwk1H3_1),.clk(gclk));
	jdff dff_B_A0jSQbd32_0(.din(n250),.dout(w_dff_B_A0jSQbd32_0),.clk(gclk));
	jdff dff_B_ZelMu73y6_0(.din(w_dff_B_A0jSQbd32_0),.dout(w_dff_B_ZelMu73y6_0),.clk(gclk));
	jdff dff_B_khC0ug2t3_0(.din(w_dff_B_ZelMu73y6_0),.dout(w_dff_B_khC0ug2t3_0),.clk(gclk));
	jdff dff_B_DjfMI7uu4_0(.din(w_dff_B_khC0ug2t3_0),.dout(w_dff_B_DjfMI7uu4_0),.clk(gclk));
	jdff dff_B_MFvsdWBy7_0(.din(w_dff_B_DjfMI7uu4_0),.dout(w_dff_B_MFvsdWBy7_0),.clk(gclk));
	jdff dff_B_5Bjpjaiq3_0(.din(n248),.dout(w_dff_B_5Bjpjaiq3_0),.clk(gclk));
	jdff dff_B_VZlolp058_0(.din(w_dff_B_5Bjpjaiq3_0),.dout(w_dff_B_VZlolp058_0),.clk(gclk));
	jdff dff_B_zwv9qhOX5_0(.din(w_dff_B_VZlolp058_0),.dout(w_dff_B_zwv9qhOX5_0),.clk(gclk));
	jdff dff_B_K5lGTDEM3_0(.din(n247),.dout(w_dff_B_K5lGTDEM3_0),.clk(gclk));
	jdff dff_B_53uxGn3G2_0(.din(w_dff_B_K5lGTDEM3_0),.dout(w_dff_B_53uxGn3G2_0),.clk(gclk));
	jdff dff_B_YW3Yrrpb5_0(.din(w_dff_B_53uxGn3G2_0),.dout(w_dff_B_YW3Yrrpb5_0),.clk(gclk));
	jdff dff_B_gR5RYfHF0_0(.din(w_dff_B_YW3Yrrpb5_0),.dout(w_dff_B_gR5RYfHF0_0),.clk(gclk));
	jdff dff_B_eBN9lLZU9_0(.din(n244),.dout(w_dff_B_eBN9lLZU9_0),.clk(gclk));
	jdff dff_B_8Q4QnE9a2_0(.din(w_dff_B_eBN9lLZU9_0),.dout(w_dff_B_8Q4QnE9a2_0),.clk(gclk));
	jdff dff_B_yUhUZWtt3_0(.din(w_dff_B_8Q4QnE9a2_0),.dout(w_dff_B_yUhUZWtt3_0),.clk(gclk));
	jdff dff_B_ydxMKmUe2_0(.din(w_dff_B_yUhUZWtt3_0),.dout(w_dff_B_ydxMKmUe2_0),.clk(gclk));
	jdff dff_B_EvIZxbTB2_0(.din(w_dff_B_ydxMKmUe2_0),.dout(w_dff_B_EvIZxbTB2_0),.clk(gclk));
	jdff dff_B_MxYrP5QC5_0(.din(w_dff_B_EvIZxbTB2_0),.dout(w_dff_B_MxYrP5QC5_0),.clk(gclk));
	jdff dff_A_dtsjmMvx8_0(.dout(w_G219gat_3[0]),.din(w_dff_A_dtsjmMvx8_0),.clk(gclk));
	jdff dff_A_tlWR1w6w5_0(.dout(w_dff_A_dtsjmMvx8_0),.din(w_dff_A_tlWR1w6w5_0),.clk(gclk));
	jdff dff_A_53eI4pQg0_0(.dout(w_dff_A_tlWR1w6w5_0),.din(w_dff_A_53eI4pQg0_0),.clk(gclk));
	jdff dff_A_EJDOXZUE8_0(.dout(w_dff_A_53eI4pQg0_0),.din(w_dff_A_EJDOXZUE8_0),.clk(gclk));
	jdff dff_B_NAQTZAus9_1(.din(n195),.dout(w_dff_B_NAQTZAus9_1),.clk(gclk));
	jdff dff_B_HmJUGg7H5_1(.din(w_dff_B_NAQTZAus9_1),.dout(w_dff_B_HmJUGg7H5_1),.clk(gclk));
	jdff dff_B_vrgnYpuX7_1(.din(w_dff_B_HmJUGg7H5_1),.dout(w_dff_B_vrgnYpuX7_1),.clk(gclk));
	jdff dff_B_J7uiEXF66_1(.din(w_dff_B_vrgnYpuX7_1),.dout(w_dff_B_J7uiEXF66_1),.clk(gclk));
	jdff dff_A_Mh1l4sjP7_1(.dout(w_n194_0[1]),.din(w_dff_A_Mh1l4sjP7_1),.clk(gclk));
	jdff dff_A_SkIorOFb3_1(.dout(w_dff_A_Mh1l4sjP7_1),.din(w_dff_A_SkIorOFb3_1),.clk(gclk));
	jdff dff_A_BGzuIdcz9_1(.dout(w_dff_A_SkIorOFb3_1),.din(w_dff_A_BGzuIdcz9_1),.clk(gclk));
	jdff dff_A_mVPNFlTl0_1(.dout(w_dff_A_BGzuIdcz9_1),.din(w_dff_A_mVPNFlTl0_1),.clk(gclk));
	jdff dff_A_mqtz29nv3_0(.dout(w_G183gat_2[0]),.din(w_dff_A_mqtz29nv3_0),.clk(gclk));
	jdff dff_A_JVSnyORT2_0(.dout(w_dff_A_mqtz29nv3_0),.din(w_dff_A_JVSnyORT2_0),.clk(gclk));
	jdff dff_A_1JKA2zIv4_0(.dout(w_dff_A_JVSnyORT2_0),.din(w_dff_A_1JKA2zIv4_0),.clk(gclk));
	jdff dff_A_oOzkPEPs5_0(.dout(w_dff_A_1JKA2zIv4_0),.din(w_dff_A_oOzkPEPs5_0),.clk(gclk));
	jdff dff_A_El0hZZmp6_0(.dout(w_dff_A_oOzkPEPs5_0),.din(w_dff_A_El0hZZmp6_0),.clk(gclk));
	jdff dff_A_tiZ38Rkz4_0(.dout(w_dff_A_El0hZZmp6_0),.din(w_dff_A_tiZ38Rkz4_0),.clk(gclk));
	jdff dff_A_72Ud20aI9_0(.dout(w_dff_A_tiZ38Rkz4_0),.din(w_dff_A_72Ud20aI9_0),.clk(gclk));
	jdff dff_A_yvRtKMeT2_0(.dout(w_dff_A_72Ud20aI9_0),.din(w_dff_A_yvRtKMeT2_0),.clk(gclk));
	jdff dff_B_ho6uvlZN0_0(.din(n271),.dout(w_dff_B_ho6uvlZN0_0),.clk(gclk));
	jdff dff_B_I6hY2S6W7_0(.din(w_dff_B_ho6uvlZN0_0),.dout(w_dff_B_I6hY2S6W7_0),.clk(gclk));
	jdff dff_B_tnQsj0tV8_0(.din(w_dff_B_I6hY2S6W7_0),.dout(w_dff_B_tnQsj0tV8_0),.clk(gclk));
	jdff dff_B_XHSx1ZBu3_0(.din(w_dff_B_tnQsj0tV8_0),.dout(w_dff_B_XHSx1ZBu3_0),.clk(gclk));
	jdff dff_B_ZKSjb0ht7_0(.din(w_dff_B_XHSx1ZBu3_0),.dout(w_dff_B_ZKSjb0ht7_0),.clk(gclk));
	jdff dff_B_wfrQhoPj6_0(.din(n269),.dout(w_dff_B_wfrQhoPj6_0),.clk(gclk));
	jdff dff_B_nzPYfjuJ0_0(.din(w_dff_B_wfrQhoPj6_0),.dout(w_dff_B_nzPYfjuJ0_0),.clk(gclk));
	jdff dff_B_IfB1r0h09_0(.din(w_dff_B_nzPYfjuJ0_0),.dout(w_dff_B_IfB1r0h09_0),.clk(gclk));
	jdff dff_B_hlTtz6bQ7_0(.din(n268),.dout(w_dff_B_hlTtz6bQ7_0),.clk(gclk));
	jdff dff_B_Beu8LTgM6_0(.din(w_dff_B_hlTtz6bQ7_0),.dout(w_dff_B_Beu8LTgM6_0),.clk(gclk));
	jdff dff_B_gKnj4rBG1_0(.din(w_dff_B_Beu8LTgM6_0),.dout(w_dff_B_gKnj4rBG1_0),.clk(gclk));
	jdff dff_B_Hk1vbXn17_0(.din(n263),.dout(w_dff_B_Hk1vbXn17_0),.clk(gclk));
	jdff dff_B_p4axHPQU7_0(.din(w_dff_B_Hk1vbXn17_0),.dout(w_dff_B_p4axHPQU7_0),.clk(gclk));
	jdff dff_B_0JCT6MEU5_0(.din(w_dff_B_p4axHPQU7_0),.dout(w_dff_B_0JCT6MEU5_0),.clk(gclk));
	jdff dff_B_BHnfWOY67_0(.din(w_dff_B_0JCT6MEU5_0),.dout(w_dff_B_BHnfWOY67_0),.clk(gclk));
	jdff dff_B_r9j17qxj2_0(.din(w_dff_B_BHnfWOY67_0),.dout(w_dff_B_r9j17qxj2_0),.clk(gclk));
	jdff dff_B_iKCGrPsq2_0(.din(w_dff_B_r9j17qxj2_0),.dout(w_dff_B_iKCGrPsq2_0),.clk(gclk));
	jdff dff_B_9PG3ojBh5_1(.din(n253),.dout(w_dff_B_9PG3ojBh5_1),.clk(gclk));
	jdff dff_B_Js87Eamr8_1(.din(w_dff_B_9PG3ojBh5_1),.dout(w_dff_B_Js87Eamr8_1),.clk(gclk));
	jdff dff_B_QtNeyt9Z9_1(.din(w_dff_B_Js87Eamr8_1),.dout(w_dff_B_QtNeyt9Z9_1),.clk(gclk));
	jdff dff_B_C5AC7Cip1_1(.din(w_dff_B_QtNeyt9Z9_1),.dout(w_dff_B_C5AC7Cip1_1),.clk(gclk));
	jdff dff_A_sTJD3KC79_1(.dout(w_n252_0[1]),.din(w_dff_A_sTJD3KC79_1),.clk(gclk));
	jdff dff_A_KIfhSZCt4_1(.dout(w_dff_A_sTJD3KC79_1),.din(w_dff_A_KIfhSZCt4_1),.clk(gclk));
	jdff dff_A_Cp6SfsxI7_1(.dout(w_dff_A_KIfhSZCt4_1),.din(w_dff_A_Cp6SfsxI7_1),.clk(gclk));
	jdff dff_A_IySSeJOx0_1(.dout(w_dff_A_Cp6SfsxI7_1),.din(w_dff_A_IySSeJOx0_1),.clk(gclk));
	jdff dff_B_Kcj0PMBs5_0(.din(n289),.dout(w_dff_B_Kcj0PMBs5_0),.clk(gclk));
	jdff dff_B_RS7rAgY10_0(.din(w_dff_B_Kcj0PMBs5_0),.dout(w_dff_B_RS7rAgY10_0),.clk(gclk));
	jdff dff_B_KbnTInxV4_0(.din(w_dff_B_RS7rAgY10_0),.dout(w_dff_B_KbnTInxV4_0),.clk(gclk));
	jdff dff_B_3hReHb1S3_0(.din(n287),.dout(w_dff_B_3hReHb1S3_0),.clk(gclk));
	jdff dff_B_7Ro2bqcZ9_0(.din(w_dff_B_3hReHb1S3_0),.dout(w_dff_B_7Ro2bqcZ9_0),.clk(gclk));
	jdff dff_B_sDU7CWKL3_0(.din(w_dff_B_7Ro2bqcZ9_0),.dout(w_dff_B_sDU7CWKL3_0),.clk(gclk));
	jdff dff_B_MEe6xGvZ3_0(.din(n286),.dout(w_dff_B_MEe6xGvZ3_0),.clk(gclk));
	jdff dff_B_39uTlUH40_0(.din(w_dff_B_MEe6xGvZ3_0),.dout(w_dff_B_39uTlUH40_0),.clk(gclk));
	jdff dff_B_ccXQruad6_0(.din(w_dff_B_39uTlUH40_0),.dout(w_dff_B_ccXQruad6_0),.clk(gclk));
	jdff dff_B_4vc40hgv7_0(.din(n281),.dout(w_dff_B_4vc40hgv7_0),.clk(gclk));
	jdff dff_B_L4UgJcEY6_0(.din(w_dff_B_4vc40hgv7_0),.dout(w_dff_B_L4UgJcEY6_0),.clk(gclk));
	jdff dff_B_Rn4toji56_0(.din(w_dff_B_L4UgJcEY6_0),.dout(w_dff_B_Rn4toji56_0),.clk(gclk));
	jdff dff_B_JF5mahsl5_0(.din(w_dff_B_Rn4toji56_0),.dout(w_dff_B_JF5mahsl5_0),.clk(gclk));
	jdff dff_B_01hQ1cwc4_0(.din(w_dff_B_JF5mahsl5_0),.dout(w_dff_B_01hQ1cwc4_0),.clk(gclk));
	jdff dff_B_hIcihech9_0(.din(w_dff_B_01hQ1cwc4_0),.dout(w_dff_B_hIcihech9_0),.clk(gclk));
	jdff dff_B_xsxlOgxW3_0(.din(n274),.dout(w_dff_B_xsxlOgxW3_0),.clk(gclk));
	jdff dff_B_eUvIE2o32_0(.din(w_dff_B_xsxlOgxW3_0),.dout(w_dff_B_eUvIE2o32_0),.clk(gclk));
	jdff dff_A_T4dEj9Ob6_1(.dout(w_n273_0[1]),.din(w_dff_A_T4dEj9Ob6_1),.clk(gclk));
	jdff dff_A_DizNzasm0_1(.dout(w_dff_A_T4dEj9Ob6_1),.din(w_dff_A_DizNzasm0_1),.clk(gclk));
	jdff dff_B_3YdSgdhR7_1(.din(n300),.dout(w_dff_B_3YdSgdhR7_1),.clk(gclk));
	jdff dff_B_LWTMNUNt7_1(.din(w_dff_B_3YdSgdhR7_1),.dout(w_dff_B_LWTMNUNt7_1),.clk(gclk));
	jdff dff_B_IIetBZfP8_1(.din(w_dff_B_LWTMNUNt7_1),.dout(w_dff_B_IIetBZfP8_1),.clk(gclk));
	jdff dff_B_V9V0yxRE2_1(.din(w_dff_B_IIetBZfP8_1),.dout(w_dff_B_V9V0yxRE2_1),.clk(gclk));
	jdff dff_B_AnPgj2KF8_1(.din(w_dff_B_V9V0yxRE2_1),.dout(w_dff_B_AnPgj2KF8_1),.clk(gclk));
	jdff dff_B_u8fZuA1f0_1(.din(w_dff_B_AnPgj2KF8_1),.dout(w_dff_B_u8fZuA1f0_1),.clk(gclk));
	jdff dff_B_83ceRUQp2_1(.din(w_dff_B_u8fZuA1f0_1),.dout(w_dff_B_83ceRUQp2_1),.clk(gclk));
	jdff dff_B_tgHPkVDP5_1(.din(w_dff_B_83ceRUQp2_1),.dout(w_dff_B_tgHPkVDP5_1),.clk(gclk));
	jdff dff_B_pzyD4PB77_1(.din(w_dff_B_tgHPkVDP5_1),.dout(w_dff_B_pzyD4PB77_1),.clk(gclk));
	jdff dff_B_drA7A5wC2_1(.din(w_dff_B_pzyD4PB77_1),.dout(w_dff_B_drA7A5wC2_1),.clk(gclk));
	jdff dff_B_yykAJLWp3_1(.din(n301),.dout(w_dff_B_yykAJLWp3_1),.clk(gclk));
	jdff dff_B_8izQVtUh2_1(.din(w_dff_B_yykAJLWp3_1),.dout(w_dff_B_8izQVtUh2_1),.clk(gclk));
	jdff dff_B_KDxHs3hd5_1(.din(w_dff_B_8izQVtUh2_1),.dout(w_dff_B_KDxHs3hd5_1),.clk(gclk));
	jdff dff_B_DnY8NSN65_1(.din(w_dff_B_KDxHs3hd5_1),.dout(w_dff_B_DnY8NSN65_1),.clk(gclk));
	jdff dff_B_NFWHi29h8_1(.din(w_dff_B_DnY8NSN65_1),.dout(w_dff_B_NFWHi29h8_1),.clk(gclk));
	jdff dff_B_dYeNWM4I5_1(.din(w_dff_B_NFWHi29h8_1),.dout(w_dff_B_dYeNWM4I5_1),.clk(gclk));
	jdff dff_B_Dq2S9tTl5_1(.din(w_dff_B_dYeNWM4I5_1),.dout(w_dff_B_Dq2S9tTl5_1),.clk(gclk));
	jdff dff_B_GFIofgPe5_1(.din(w_dff_B_Dq2S9tTl5_1),.dout(w_dff_B_GFIofgPe5_1),.clk(gclk));
	jdff dff_B_9x4JXOZc9_1(.din(w_dff_B_GFIofgPe5_1),.dout(w_dff_B_9x4JXOZc9_1),.clk(gclk));
	jdff dff_A_1VeCIsG01_0(.dout(w_G159gat_2[0]),.din(w_dff_A_1VeCIsG01_0),.clk(gclk));
	jdff dff_A_6l3YBqOA0_0(.dout(w_dff_A_1VeCIsG01_0),.din(w_dff_A_6l3YBqOA0_0),.clk(gclk));
	jdff dff_A_OUxX7aTZ4_0(.dout(w_dff_A_6l3YBqOA0_0),.din(w_dff_A_OUxX7aTZ4_0),.clk(gclk));
	jdff dff_A_HMxZArqn0_0(.dout(w_dff_A_OUxX7aTZ4_0),.din(w_dff_A_HMxZArqn0_0),.clk(gclk));
	jdff dff_A_ueE7Fqvm8_0(.dout(w_dff_A_HMxZArqn0_0),.din(w_dff_A_ueE7Fqvm8_0),.clk(gclk));
	jdff dff_A_6NhCLcMG5_0(.dout(w_dff_A_ueE7Fqvm8_0),.din(w_dff_A_6NhCLcMG5_0),.clk(gclk));
	jdff dff_A_T5wby41Q7_0(.dout(w_dff_A_6NhCLcMG5_0),.din(w_dff_A_T5wby41Q7_0),.clk(gclk));
	jdff dff_B_NohDFIkr6_0(.din(n361),.dout(w_dff_B_NohDFIkr6_0),.clk(gclk));
	jdff dff_B_g2q1NrVl8_0(.din(w_dff_B_NohDFIkr6_0),.dout(w_dff_B_g2q1NrVl8_0),.clk(gclk));
	jdff dff_B_HupO2SMB8_0(.din(w_dff_B_g2q1NrVl8_0),.dout(w_dff_B_HupO2SMB8_0),.clk(gclk));
	jdff dff_B_Awq6aRL81_0(.din(w_dff_B_HupO2SMB8_0),.dout(w_dff_B_Awq6aRL81_0),.clk(gclk));
	jdff dff_B_PS80H6pj5_0(.din(w_dff_B_Awq6aRL81_0),.dout(w_dff_B_PS80H6pj5_0),.clk(gclk));
	jdff dff_B_2jCX0utf5_0(.din(w_dff_B_PS80H6pj5_0),.dout(w_dff_B_2jCX0utf5_0),.clk(gclk));
	jdff dff_B_SHvCg2vu0_0(.din(w_dff_B_2jCX0utf5_0),.dout(w_dff_B_SHvCg2vu0_0),.clk(gclk));
	jdff dff_B_ZvgTSLK49_0(.din(w_dff_B_SHvCg2vu0_0),.dout(w_dff_B_ZvgTSLK49_0),.clk(gclk));
	jdff dff_B_3cwJJFb74_0(.din(n359),.dout(w_dff_B_3cwJJFb74_0),.clk(gclk));
	jdff dff_B_lE9VLwQq3_0(.din(w_dff_B_3cwJJFb74_0),.dout(w_dff_B_lE9VLwQq3_0),.clk(gclk));
	jdff dff_B_dIKLuiks4_0(.din(n358),.dout(w_dff_B_dIKLuiks4_0),.clk(gclk));
	jdff dff_B_PT4MfKwO1_0(.din(w_dff_B_dIKLuiks4_0),.dout(w_dff_B_PT4MfKwO1_0),.clk(gclk));
	jdff dff_B_TuSVCqe91_0(.din(w_dff_B_PT4MfKwO1_0),.dout(w_dff_B_TuSVCqe91_0),.clk(gclk));
	jdff dff_B_1iohtdfD7_0(.din(w_dff_B_TuSVCqe91_0),.dout(w_dff_B_1iohtdfD7_0),.clk(gclk));
	jdff dff_B_dEiiDR826_0(.din(n355),.dout(w_dff_B_dEiiDR826_0),.clk(gclk));
	jdff dff_B_eHewIdvm5_0(.din(w_dff_B_dEiiDR826_0),.dout(w_dff_B_eHewIdvm5_0),.clk(gclk));
	jdff dff_B_dyuU603b1_0(.din(w_dff_B_eHewIdvm5_0),.dout(w_dff_B_dyuU603b1_0),.clk(gclk));
	jdff dff_B_4S9IAbVG3_0(.din(w_dff_B_dyuU603b1_0),.dout(w_dff_B_4S9IAbVG3_0),.clk(gclk));
	jdff dff_B_58zR0n3s1_0(.din(w_dff_B_4S9IAbVG3_0),.dout(w_dff_B_58zR0n3s1_0),.clk(gclk));
	jdff dff_A_iFem6Mhk9_1(.dout(w_G228gat_2[1]),.din(w_dff_A_iFem6Mhk9_1),.clk(gclk));
	jdff dff_A_1u7JjUPF2_2(.dout(w_G228gat_2[2]),.din(w_dff_A_1u7JjUPF2_2),.clk(gclk));
	jdff dff_A_iy772LK66_0(.dout(w_G219gat_2[0]),.din(w_dff_A_iy772LK66_0),.clk(gclk));
	jdff dff_A_RjFmsIgn2_0(.dout(w_dff_A_iy772LK66_0),.din(w_dff_A_RjFmsIgn2_0),.clk(gclk));
	jdff dff_A_AHRPNo1Y6_0(.dout(w_dff_A_RjFmsIgn2_0),.din(w_dff_A_AHRPNo1Y6_0),.clk(gclk));
	jdff dff_A_10DzDZaA4_0(.dout(w_dff_A_AHRPNo1Y6_0),.din(w_dff_A_10DzDZaA4_0),.clk(gclk));
	jdff dff_A_57hrO2Mz8_2(.dout(w_G219gat_2[2]),.din(w_dff_A_57hrO2Mz8_2),.clk(gclk));
	jdff dff_A_qRXtUuAr5_2(.dout(w_dff_A_57hrO2Mz8_2),.din(w_dff_A_qRXtUuAr5_2),.clk(gclk));
	jdff dff_B_n7vBmzCc0_0(.din(n348),.dout(w_dff_B_n7vBmzCc0_0),.clk(gclk));
	jdff dff_B_W6AUlIsY8_0(.din(w_dff_B_n7vBmzCc0_0),.dout(w_dff_B_W6AUlIsY8_0),.clk(gclk));
	jdff dff_B_REeXiNpg3_0(.din(w_dff_B_W6AUlIsY8_0),.dout(w_dff_B_REeXiNpg3_0),.clk(gclk));
	jdff dff_B_tdBjlrPr4_0(.din(w_dff_B_REeXiNpg3_0),.dout(w_dff_B_tdBjlrPr4_0),.clk(gclk));
	jdff dff_B_MRBmsPZg6_0(.din(w_dff_B_tdBjlrPr4_0),.dout(w_dff_B_MRBmsPZg6_0),.clk(gclk));
	jdff dff_B_DduR3R5e2_0(.din(w_dff_B_MRBmsPZg6_0),.dout(w_dff_B_DduR3R5e2_0),.clk(gclk));
	jdff dff_B_44poXEwj6_0(.din(w_dff_B_DduR3R5e2_0),.dout(w_dff_B_44poXEwj6_0),.clk(gclk));
	jdff dff_A_023pSUSL8_1(.dout(w_n347_0[1]),.din(w_dff_A_023pSUSL8_1),.clk(gclk));
	jdff dff_A_mQ522mJ64_1(.dout(w_dff_A_023pSUSL8_1),.din(w_dff_A_mQ522mJ64_1),.clk(gclk));
	jdff dff_A_uWHcZJfe4_1(.dout(w_dff_A_mQ522mJ64_1),.din(w_dff_A_uWHcZJfe4_1),.clk(gclk));
	jdff dff_A_wEDMyrs09_1(.dout(w_dff_A_uWHcZJfe4_1),.din(w_dff_A_wEDMyrs09_1),.clk(gclk));
	jdff dff_A_mzoGyn4B0_1(.dout(w_dff_A_wEDMyrs09_1),.din(w_dff_A_mzoGyn4B0_1),.clk(gclk));
	jdff dff_A_0u0C7DSN1_1(.dout(w_dff_A_mzoGyn4B0_1),.din(w_dff_A_0u0C7DSN1_1),.clk(gclk));
	jdff dff_A_382X31nZ2_1(.dout(w_dff_A_0u0C7DSN1_1),.din(w_dff_A_382X31nZ2_1),.clk(gclk));
	jdff dff_B_RbdGLSY84_0(.din(n381),.dout(w_dff_B_RbdGLSY84_0),.clk(gclk));
	jdff dff_B_DCjs5pew3_0(.din(w_dff_B_RbdGLSY84_0),.dout(w_dff_B_DCjs5pew3_0),.clk(gclk));
	jdff dff_B_Qh2DSA8C9_0(.din(w_dff_B_DCjs5pew3_0),.dout(w_dff_B_Qh2DSA8C9_0),.clk(gclk));
	jdff dff_B_8MAWAhCN2_0(.din(w_dff_B_Qh2DSA8C9_0),.dout(w_dff_B_8MAWAhCN2_0),.clk(gclk));
	jdff dff_B_3HOLFLU23_0(.din(w_dff_B_8MAWAhCN2_0),.dout(w_dff_B_3HOLFLU23_0),.clk(gclk));
	jdff dff_B_UdIWA2le0_0(.din(w_dff_B_3HOLFLU23_0),.dout(w_dff_B_UdIWA2le0_0),.clk(gclk));
	jdff dff_B_K8L4snng6_0(.din(w_dff_B_UdIWA2le0_0),.dout(w_dff_B_K8L4snng6_0),.clk(gclk));
	jdff dff_B_SV1T3fdX5_0(.din(w_dff_B_K8L4snng6_0),.dout(w_dff_B_SV1T3fdX5_0),.clk(gclk));
	jdff dff_B_6y7RmwYH6_0(.din(w_dff_B_SV1T3fdX5_0),.dout(w_dff_B_6y7RmwYH6_0),.clk(gclk));
	jdff dff_B_hfzIin7F9_0(.din(w_dff_B_6y7RmwYH6_0),.dout(w_dff_B_hfzIin7F9_0),.clk(gclk));
	jdff dff_B_XsB5ta5w8_0(.din(n379),.dout(w_dff_B_XsB5ta5w8_0),.clk(gclk));
	jdff dff_B_HzuYTE3n4_0(.din(w_dff_B_XsB5ta5w8_0),.dout(w_dff_B_HzuYTE3n4_0),.clk(gclk));
	jdff dff_B_lGaIPzou0_0(.din(n378),.dout(w_dff_B_lGaIPzou0_0),.clk(gclk));
	jdff dff_B_oxWpBES39_0(.din(w_dff_B_lGaIPzou0_0),.dout(w_dff_B_oxWpBES39_0),.clk(gclk));
	jdff dff_B_O4iooApG8_0(.din(w_dff_B_oxWpBES39_0),.dout(w_dff_B_O4iooApG8_0),.clk(gclk));
	jdff dff_B_Ez5N4pDZ5_0(.din(w_dff_B_O4iooApG8_0),.dout(w_dff_B_Ez5N4pDZ5_0),.clk(gclk));
	jdff dff_B_BOETqyeV1_0(.din(n375),.dout(w_dff_B_BOETqyeV1_0),.clk(gclk));
	jdff dff_B_CNQ7J28V6_0(.din(w_dff_B_BOETqyeV1_0),.dout(w_dff_B_CNQ7J28V6_0),.clk(gclk));
	jdff dff_B_7kxTMH5k9_0(.din(w_dff_B_CNQ7J28V6_0),.dout(w_dff_B_7kxTMH5k9_0),.clk(gclk));
	jdff dff_B_Ypk3RyhC7_0(.din(w_dff_B_7kxTMH5k9_0),.dout(w_dff_B_Ypk3RyhC7_0),.clk(gclk));
	jdff dff_B_Htl8yZ1Z7_0(.din(w_dff_B_Ypk3RyhC7_0),.dout(w_dff_B_Htl8yZ1Z7_0),.clk(gclk));
	jdff dff_B_vlvA8ewb1_0(.din(n368),.dout(w_dff_B_vlvA8ewb1_0),.clk(gclk));
	jdff dff_B_PVg1L6ik6_0(.din(w_dff_B_vlvA8ewb1_0),.dout(w_dff_B_PVg1L6ik6_0),.clk(gclk));
	jdff dff_B_K9MJvytw5_0(.din(w_dff_B_PVg1L6ik6_0),.dout(w_dff_B_K9MJvytw5_0),.clk(gclk));
	jdff dff_B_0vlXdP8K4_0(.din(w_dff_B_K9MJvytw5_0),.dout(w_dff_B_0vlXdP8K4_0),.clk(gclk));
	jdff dff_B_jzB7yExU8_0(.din(w_dff_B_0vlXdP8K4_0),.dout(w_dff_B_jzB7yExU8_0),.clk(gclk));
	jdff dff_B_iQYmiAqk8_0(.din(w_dff_B_jzB7yExU8_0),.dout(w_dff_B_iQYmiAqk8_0),.clk(gclk));
	jdff dff_B_QxNk1A3N2_0(.din(w_dff_B_iQYmiAqk8_0),.dout(w_dff_B_QxNk1A3N2_0),.clk(gclk));
	jdff dff_B_UMThZjei6_0(.din(w_dff_B_QxNk1A3N2_0),.dout(w_dff_B_UMThZjei6_0),.clk(gclk));
	jdff dff_B_sABVbcuN3_0(.din(w_dff_B_UMThZjei6_0),.dout(w_dff_B_sABVbcuN3_0),.clk(gclk));
	jdff dff_A_qMR68vi01_1(.dout(w_n367_0[1]),.din(w_dff_A_qMR68vi01_1),.clk(gclk));
	jdff dff_A_moYjWur72_1(.dout(w_dff_A_qMR68vi01_1),.din(w_dff_A_moYjWur72_1),.clk(gclk));
	jdff dff_A_zKQ21zr36_1(.dout(w_dff_A_moYjWur72_1),.din(w_dff_A_zKQ21zr36_1),.clk(gclk));
	jdff dff_A_sY73Bu0e0_1(.dout(w_dff_A_zKQ21zr36_1),.din(w_dff_A_sY73Bu0e0_1),.clk(gclk));
	jdff dff_A_4bTtr4l67_1(.dout(w_dff_A_sY73Bu0e0_1),.din(w_dff_A_4bTtr4l67_1),.clk(gclk));
	jdff dff_A_7YyEK7lJ1_1(.dout(w_dff_A_4bTtr4l67_1),.din(w_dff_A_7YyEK7lJ1_1),.clk(gclk));
	jdff dff_A_P6LhuJ0q7_1(.dout(w_dff_A_7YyEK7lJ1_1),.din(w_dff_A_P6LhuJ0q7_1),.clk(gclk));
	jdff dff_A_7lI4wPMX7_1(.dout(w_dff_A_P6LhuJ0q7_1),.din(w_dff_A_7lI4wPMX7_1),.clk(gclk));
	jdff dff_A_kV4L7Rfy6_1(.dout(w_dff_A_7lI4wPMX7_1),.din(w_dff_A_kV4L7Rfy6_1),.clk(gclk));
	jdff dff_B_CpyIbm2t2_1(.din(n294),.dout(w_dff_B_CpyIbm2t2_1),.clk(gclk));
	jdff dff_B_f4GQoigI6_1(.din(w_dff_B_CpyIbm2t2_1),.dout(w_dff_B_f4GQoigI6_1),.clk(gclk));
	jdff dff_B_zCnyp4Y35_1(.din(w_dff_B_f4GQoigI6_1),.dout(w_dff_B_zCnyp4Y35_1),.clk(gclk));
	jdff dff_A_nky78gyn8_1(.dout(w_G159gat_1[1]),.din(w_dff_A_nky78gyn8_1),.clk(gclk));
	jdff dff_A_VyvMVabj5_1(.dout(w_dff_A_nky78gyn8_1),.din(w_dff_A_VyvMVabj5_1),.clk(gclk));
	jdff dff_A_dZWcCDWf5_1(.dout(w_dff_A_VyvMVabj5_1),.din(w_dff_A_dZWcCDWf5_1),.clk(gclk));
	jdff dff_A_oVl6N6Q58_1(.dout(w_dff_A_dZWcCDWf5_1),.din(w_dff_A_oVl6N6Q58_1),.clk(gclk));
	jdff dff_A_MLQumjyQ5_1(.dout(w_dff_A_oVl6N6Q58_1),.din(w_dff_A_MLQumjyQ5_1),.clk(gclk));
	jdff dff_A_TjKz3ELb1_1(.dout(w_dff_A_MLQumjyQ5_1),.din(w_dff_A_TjKz3ELb1_1),.clk(gclk));
	jdff dff_A_b8BjMrtc1_1(.dout(w_dff_A_TjKz3ELb1_1),.din(w_dff_A_b8BjMrtc1_1),.clk(gclk));
	jdff dff_A_4FtGxaiL4_2(.dout(w_G159gat_1[2]),.din(w_dff_A_4FtGxaiL4_2),.clk(gclk));
	jdff dff_A_md4OBqlg8_2(.dout(w_dff_A_4FtGxaiL4_2),.din(w_dff_A_md4OBqlg8_2),.clk(gclk));
	jdff dff_A_wHAWheAa9_2(.dout(w_dff_A_md4OBqlg8_2),.din(w_dff_A_wHAWheAa9_2),.clk(gclk));
	jdff dff_A_8yc16Ims3_2(.dout(w_dff_A_wHAWheAa9_2),.din(w_dff_A_8yc16Ims3_2),.clk(gclk));
	jdff dff_A_eulngWVQ4_2(.dout(w_dff_A_8yc16Ims3_2),.din(w_dff_A_eulngWVQ4_2),.clk(gclk));
	jdff dff_A_XILNzLwa2_2(.dout(w_dff_A_eulngWVQ4_2),.din(w_dff_A_XILNzLwa2_2),.clk(gclk));
	jdff dff_A_IeRBU1Vr6_2(.dout(w_dff_A_XILNzLwa2_2),.din(w_dff_A_IeRBU1Vr6_2),.clk(gclk));
	jdff dff_A_1K3pnApX4_2(.dout(w_G159gat_0[2]),.din(w_dff_A_1K3pnApX4_2),.clk(gclk));
	jdff dff_A_QYGY4fAK9_2(.dout(w_dff_A_1K3pnApX4_2),.din(w_dff_A_QYGY4fAK9_2),.clk(gclk));
	jdff dff_A_JOkXOb1G4_2(.dout(w_dff_A_QYGY4fAK9_2),.din(w_dff_A_JOkXOb1G4_2),.clk(gclk));
	jdff dff_A_eE0L9O3I9_2(.dout(w_dff_A_JOkXOb1G4_2),.din(w_dff_A_eE0L9O3I9_2),.clk(gclk));
	jdff dff_B_E7Vdx2XL5_0(.din(n365),.dout(w_dff_B_E7Vdx2XL5_0),.clk(gclk));
	jdff dff_B_qtI8Krpp6_0(.din(w_dff_B_E7Vdx2XL5_0),.dout(w_dff_B_qtI8Krpp6_0),.clk(gclk));
	jdff dff_B_sn8D4Nq37_0(.din(w_dff_B_qtI8Krpp6_0),.dout(w_dff_B_sn8D4Nq37_0),.clk(gclk));
	jdff dff_B_qWOZGGdK5_0(.din(w_dff_B_sn8D4Nq37_0),.dout(w_dff_B_qWOZGGdK5_0),.clk(gclk));
	jdff dff_A_J7C3tMNX3_1(.dout(w_n339_0[1]),.din(w_dff_A_J7C3tMNX3_1),.clk(gclk));
	jdff dff_A_HH4gkS7P9_1(.dout(w_dff_A_J7C3tMNX3_1),.din(w_dff_A_HH4gkS7P9_1),.clk(gclk));
	jdff dff_A_uUGfd9rD4_1(.dout(w_dff_A_HH4gkS7P9_1),.din(w_dff_A_uUGfd9rD4_1),.clk(gclk));
	jdff dff_A_bPtpMy9K0_1(.dout(w_dff_A_uUGfd9rD4_1),.din(w_dff_A_bPtpMy9K0_1),.clk(gclk));
	jdff dff_B_OzhusPhr2_1(.din(n333),.dout(w_dff_B_OzhusPhr2_1),.clk(gclk));
	jdff dff_B_gVWJZjbU0_1(.din(w_dff_B_OzhusPhr2_1),.dout(w_dff_B_gVWJZjbU0_1),.clk(gclk));
	jdff dff_B_53ySjMjh9_1(.din(w_dff_B_gVWJZjbU0_1),.dout(w_dff_B_53ySjMjh9_1),.clk(gclk));
	jdff dff_B_FM5y4UtP8_0(.din(n363),.dout(w_dff_B_FM5y4UtP8_0),.clk(gclk));
	jdff dff_B_JILSaziY6_0(.din(w_dff_B_FM5y4UtP8_0),.dout(w_dff_B_JILSaziY6_0),.clk(gclk));
	jdff dff_B_JWZSHydl1_0(.din(w_dff_B_JILSaziY6_0),.dout(w_dff_B_JWZSHydl1_0),.clk(gclk));
	jdff dff_B_mmHNanG33_0(.din(w_dff_B_JWZSHydl1_0),.dout(w_dff_B_mmHNanG33_0),.clk(gclk));
	jdff dff_A_OH6QxyuU1_1(.dout(w_n331_0[1]),.din(w_dff_A_OH6QxyuU1_1),.clk(gclk));
	jdff dff_A_q1zVOeYm6_1(.dout(w_dff_A_OH6QxyuU1_1),.din(w_dff_A_q1zVOeYm6_1),.clk(gclk));
	jdff dff_A_8PprXWsr3_1(.dout(w_dff_A_q1zVOeYm6_1),.din(w_dff_A_8PprXWsr3_1),.clk(gclk));
	jdff dff_A_pWXqXzVN4_1(.dout(w_dff_A_8PprXWsr3_1),.din(w_dff_A_pWXqXzVN4_1),.clk(gclk));
	jdff dff_B_KvBNEMRH7_1(.din(n306),.dout(w_dff_B_KvBNEMRH7_1),.clk(gclk));
	jdff dff_B_5Mqvhx6I2_1(.din(w_dff_B_KvBNEMRH7_1),.dout(w_dff_B_5Mqvhx6I2_1),.clk(gclk));
	jdff dff_B_PRPPknrU4_1(.din(w_dff_B_5Mqvhx6I2_1),.dout(w_dff_B_PRPPknrU4_1),.clk(gclk));
	jdff dff_B_FSFvBsOb9_1(.din(w_dff_B_PRPPknrU4_1),.dout(w_dff_B_FSFvBsOb9_1),.clk(gclk));
	jdff dff_B_Wrp2cw9V8_1(.din(w_dff_B_FSFvBsOb9_1),.dout(w_dff_B_Wrp2cw9V8_1),.clk(gclk));
	jdff dff_B_lF2gqh2j1_1(.din(w_dff_B_Wrp2cw9V8_1),.dout(w_dff_B_lF2gqh2j1_1),.clk(gclk));
	jdff dff_B_kHduTWwA0_1(.din(w_dff_B_lF2gqh2j1_1),.dout(w_dff_B_kHduTWwA0_1),.clk(gclk));
	jdff dff_B_yl1X8NTG2_0(.din(n403),.dout(w_dff_B_yl1X8NTG2_0),.clk(gclk));
	jdff dff_B_3uw3lwSe7_0(.din(w_dff_B_yl1X8NTG2_0),.dout(w_dff_B_3uw3lwSe7_0),.clk(gclk));
	jdff dff_B_0xyM49Sd7_0(.din(w_dff_B_3uw3lwSe7_0),.dout(w_dff_B_0xyM49Sd7_0),.clk(gclk));
	jdff dff_B_zbB4NiyC9_0(.din(w_dff_B_0xyM49Sd7_0),.dout(w_dff_B_zbB4NiyC9_0),.clk(gclk));
	jdff dff_B_CPor4q7G2_0(.din(w_dff_B_zbB4NiyC9_0),.dout(w_dff_B_CPor4q7G2_0),.clk(gclk));
	jdff dff_B_BY634uEU1_0(.din(w_dff_B_CPor4q7G2_0),.dout(w_dff_B_BY634uEU1_0),.clk(gclk));
	jdff dff_B_yIo78zmx4_0(.din(w_dff_B_BY634uEU1_0),.dout(w_dff_B_yIo78zmx4_0),.clk(gclk));
	jdff dff_B_9ET7sr8X5_0(.din(w_dff_B_yIo78zmx4_0),.dout(w_dff_B_9ET7sr8X5_0),.clk(gclk));
	jdff dff_B_Cat0Iyhn9_0(.din(w_dff_B_9ET7sr8X5_0),.dout(w_dff_B_Cat0Iyhn9_0),.clk(gclk));
	jdff dff_B_MStUdTdf6_0(.din(w_dff_B_Cat0Iyhn9_0),.dout(w_dff_B_MStUdTdf6_0),.clk(gclk));
	jdff dff_B_pMQMIh1e3_0(.din(n401),.dout(w_dff_B_pMQMIh1e3_0),.clk(gclk));
	jdff dff_B_WsR0QEeq2_0(.din(w_dff_B_pMQMIh1e3_0),.dout(w_dff_B_WsR0QEeq2_0),.clk(gclk));
	jdff dff_B_DVauISiy6_0(.din(n400),.dout(w_dff_B_DVauISiy6_0),.clk(gclk));
	jdff dff_B_jcMwPvpN9_0(.din(w_dff_B_DVauISiy6_0),.dout(w_dff_B_jcMwPvpN9_0),.clk(gclk));
	jdff dff_B_EEVJq2m21_0(.din(w_dff_B_jcMwPvpN9_0),.dout(w_dff_B_EEVJq2m21_0),.clk(gclk));
	jdff dff_B_cWMBAM437_0(.din(w_dff_B_EEVJq2m21_0),.dout(w_dff_B_cWMBAM437_0),.clk(gclk));
	jdff dff_A_huryzMfF8_1(.dout(w_G91gat_0[1]),.din(w_dff_A_huryzMfF8_1),.clk(gclk));
	jdff dff_A_DgfzQoCX4_1(.dout(w_dff_A_huryzMfF8_1),.din(w_dff_A_DgfzQoCX4_1),.clk(gclk));
	jdff dff_A_4DlfPjRV8_1(.dout(w_dff_A_DgfzQoCX4_1),.din(w_dff_A_4DlfPjRV8_1),.clk(gclk));
	jdff dff_A_sdEtRUsN7_1(.dout(w_dff_A_4DlfPjRV8_1),.din(w_dff_A_sdEtRUsN7_1),.clk(gclk));
	jdff dff_A_bvAjlEZl6_1(.dout(w_dff_A_sdEtRUsN7_1),.din(w_dff_A_bvAjlEZl6_1),.clk(gclk));
	jdff dff_B_BW1dvTRe2_0(.din(n397),.dout(w_dff_B_BW1dvTRe2_0),.clk(gclk));
	jdff dff_B_xEHoGlVx5_0(.din(w_dff_B_BW1dvTRe2_0),.dout(w_dff_B_xEHoGlVx5_0),.clk(gclk));
	jdff dff_B_PKDxjfiw4_0(.din(w_dff_B_xEHoGlVx5_0),.dout(w_dff_B_PKDxjfiw4_0),.clk(gclk));
	jdff dff_B_HylNPQSS2_0(.din(w_dff_B_PKDxjfiw4_0),.dout(w_dff_B_HylNPQSS2_0),.clk(gclk));
	jdff dff_B_3oznaR7T2_0(.din(w_dff_B_HylNPQSS2_0),.dout(w_dff_B_3oznaR7T2_0),.clk(gclk));
	jdff dff_B_ZZyaLcAX0_1(.din(n384),.dout(w_dff_B_ZZyaLcAX0_1),.clk(gclk));
	jdff dff_B_EOmmUq8M2_1(.din(w_dff_B_ZZyaLcAX0_1),.dout(w_dff_B_EOmmUq8M2_1),.clk(gclk));
	jdff dff_B_fc3ZsHN80_1(.din(w_dff_B_EOmmUq8M2_1),.dout(w_dff_B_fc3ZsHN80_1),.clk(gclk));
	jdff dff_B_xdlkKpp82_1(.din(w_dff_B_fc3ZsHN80_1),.dout(w_dff_B_xdlkKpp82_1),.clk(gclk));
	jdff dff_B_ybFmn4pW7_1(.din(w_dff_B_xdlkKpp82_1),.dout(w_dff_B_ybFmn4pW7_1),.clk(gclk));
	jdff dff_B_jupaB5j52_1(.din(w_dff_B_ybFmn4pW7_1),.dout(w_dff_B_jupaB5j52_1),.clk(gclk));
	jdff dff_B_j71rhLtx1_1(.din(w_dff_B_jupaB5j52_1),.dout(w_dff_B_j71rhLtx1_1),.clk(gclk));
	jdff dff_B_HlHsTkUR3_1(.din(w_dff_B_j71rhLtx1_1),.dout(w_dff_B_HlHsTkUR3_1),.clk(gclk));
	jdff dff_B_2sqQBAbT8_1(.din(w_dff_B_HlHsTkUR3_1),.dout(w_dff_B_2sqQBAbT8_1),.clk(gclk));
	jdff dff_B_pkhHLovh9_1(.din(n385),.dout(w_dff_B_pkhHLovh9_1),.clk(gclk));
	jdff dff_B_2qkoVUpD3_1(.din(w_dff_B_pkhHLovh9_1),.dout(w_dff_B_2qkoVUpD3_1),.clk(gclk));
	jdff dff_B_SMdlVIcZ8_1(.din(w_dff_B_2qkoVUpD3_1),.dout(w_dff_B_SMdlVIcZ8_1),.clk(gclk));
	jdff dff_B_iKDwu7rb1_1(.din(w_dff_B_SMdlVIcZ8_1),.dout(w_dff_B_iKDwu7rb1_1),.clk(gclk));
	jdff dff_B_ld0lXjEs6_1(.din(w_dff_B_iKDwu7rb1_1),.dout(w_dff_B_ld0lXjEs6_1),.clk(gclk));
	jdff dff_B_LMygMd880_1(.din(w_dff_B_ld0lXjEs6_1),.dout(w_dff_B_LMygMd880_1),.clk(gclk));
	jdff dff_B_EIyeCtko2_0(.din(n386),.dout(w_dff_B_EIyeCtko2_0),.clk(gclk));
	jdff dff_B_I3CFtX3L4_0(.din(w_dff_B_EIyeCtko2_0),.dout(w_dff_B_I3CFtX3L4_0),.clk(gclk));
	jdff dff_B_UsUkjvnh0_0(.din(w_dff_B_I3CFtX3L4_0),.dout(w_dff_B_UsUkjvnh0_0),.clk(gclk));
	jdff dff_B_XZ6M5iqW0_0(.din(w_dff_B_UsUkjvnh0_0),.dout(w_dff_B_XZ6M5iqW0_0),.clk(gclk));
	jdff dff_B_qVPQL56h8_0(.din(w_dff_B_XZ6M5iqW0_0),.dout(w_dff_B_qVPQL56h8_0),.clk(gclk));
	jdff dff_B_uubzqeWb6_0(.din(w_dff_B_qVPQL56h8_0),.dout(w_dff_B_uubzqeWb6_0),.clk(gclk));
	jdff dff_A_L2TC5P8y6_0(.dout(w_n330_0[0]),.din(w_dff_A_L2TC5P8y6_0),.clk(gclk));
	jdff dff_A_TFkQEriz5_0(.dout(w_dff_A_L2TC5P8y6_0),.din(w_dff_A_TFkQEriz5_0),.clk(gclk));
	jdff dff_A_rkDR5gqQ1_0(.dout(w_dff_A_TFkQEriz5_0),.din(w_dff_A_rkDR5gqQ1_0),.clk(gclk));
	jdff dff_A_UtsoPKga7_0(.dout(w_dff_A_rkDR5gqQ1_0),.din(w_dff_A_UtsoPKga7_0),.clk(gclk));
	jdff dff_A_Wx3p4QbY8_0(.dout(w_dff_A_UtsoPKga7_0),.din(w_dff_A_Wx3p4QbY8_0),.clk(gclk));
	jdff dff_A_qQw0GRV41_0(.dout(w_dff_A_Wx3p4QbY8_0),.din(w_dff_A_qQw0GRV41_0),.clk(gclk));
	jdff dff_A_DhhcOSpl4_2(.dout(w_n330_0[2]),.din(w_dff_A_DhhcOSpl4_2),.clk(gclk));
	jdff dff_A_WpOXLQxj0_0(.dout(w_n337_0[0]),.din(w_dff_A_WpOXLQxj0_0),.clk(gclk));
	jdff dff_A_InH4zSMu5_0(.dout(w_dff_A_WpOXLQxj0_0),.din(w_dff_A_InH4zSMu5_0),.clk(gclk));
	jdff dff_A_KDppmavv5_0(.dout(w_dff_A_InH4zSMu5_0),.din(w_dff_A_KDppmavv5_0),.clk(gclk));
	jdff dff_A_cjxMoRST6_0(.dout(w_dff_A_KDppmavv5_0),.din(w_dff_A_cjxMoRST6_0),.clk(gclk));
	jdff dff_A_vKL0uEsy8_0(.dout(w_dff_A_cjxMoRST6_0),.din(w_dff_A_vKL0uEsy8_0),.clk(gclk));
	jdff dff_A_pRnFC8hN5_0(.dout(w_dff_A_vKL0uEsy8_0),.din(w_dff_A_pRnFC8hN5_0),.clk(gclk));
	jdff dff_B_oNIztZJx2_1(.din(n334),.dout(w_dff_B_oNIztZJx2_1),.clk(gclk));
	jdff dff_A_UiZv4fgH0_0(.dout(w_G171gat_2[0]),.din(w_dff_A_UiZv4fgH0_0),.clk(gclk));
	jdff dff_A_EXWGyaFA6_0(.dout(w_dff_A_UiZv4fgH0_0),.din(w_dff_A_EXWGyaFA6_0),.clk(gclk));
	jdff dff_A_vrWLk6sg1_0(.dout(w_dff_A_EXWGyaFA6_0),.din(w_dff_A_vrWLk6sg1_0),.clk(gclk));
	jdff dff_A_aYU9cUQL8_0(.dout(w_dff_A_vrWLk6sg1_0),.din(w_dff_A_aYU9cUQL8_0),.clk(gclk));
	jdff dff_A_IqClEjgr2_0(.dout(w_dff_A_aYU9cUQL8_0),.din(w_dff_A_IqClEjgr2_0),.clk(gclk));
	jdff dff_A_4EofUg327_0(.dout(w_dff_A_IqClEjgr2_0),.din(w_dff_A_4EofUg327_0),.clk(gclk));
	jdff dff_A_tZ4AwOED6_0(.dout(w_dff_A_4EofUg327_0),.din(w_dff_A_tZ4AwOED6_0),.clk(gclk));
	jdff dff_A_pSwKBWbz1_1(.dout(w_n383_0[1]),.din(w_dff_A_pSwKBWbz1_1),.clk(gclk));
	jdff dff_A_MW8qoubo6_1(.dout(w_dff_A_pSwKBWbz1_1),.din(w_dff_A_MW8qoubo6_1),.clk(gclk));
	jdff dff_A_Xgz0D3YQ3_1(.dout(w_dff_A_MW8qoubo6_1),.din(w_dff_A_Xgz0D3YQ3_1),.clk(gclk));
	jdff dff_A_SjYP66qU4_1(.dout(w_dff_A_Xgz0D3YQ3_1),.din(w_dff_A_SjYP66qU4_1),.clk(gclk));
	jdff dff_A_thKKhcRZ4_1(.dout(w_dff_A_SjYP66qU4_1),.din(w_dff_A_thKKhcRZ4_1),.clk(gclk));
	jdff dff_A_fh4unqz22_1(.dout(w_dff_A_thKKhcRZ4_1),.din(w_dff_A_fh4unqz22_1),.clk(gclk));
	jdff dff_A_f8xT1ohz1_1(.dout(w_dff_A_fh4unqz22_1),.din(w_dff_A_f8xT1ohz1_1),.clk(gclk));
	jdff dff_A_CIkqZ35X6_1(.dout(w_dff_A_f8xT1ohz1_1),.din(w_dff_A_CIkqZ35X6_1),.clk(gclk));
	jdff dff_A_sx4S7KWf4_1(.dout(w_dff_A_CIkqZ35X6_1),.din(w_dff_A_sx4S7KWf4_1),.clk(gclk));
	jdff dff_B_N8KTnB2I2_0(.din(n309),.dout(w_dff_B_N8KTnB2I2_0),.clk(gclk));
	jdff dff_B_uRv1tsp57_0(.din(w_dff_B_N8KTnB2I2_0),.dout(w_dff_B_uRv1tsp57_0),.clk(gclk));
	jdff dff_B_vydm3phq2_0(.din(w_dff_B_uRv1tsp57_0),.dout(w_dff_B_vydm3phq2_0),.clk(gclk));
	jdff dff_A_7U5ieRNk3_1(.dout(w_G165gat_1[1]),.din(w_dff_A_7U5ieRNk3_1),.clk(gclk));
	jdff dff_A_uQWYk0R27_1(.dout(w_dff_A_7U5ieRNk3_1),.din(w_dff_A_uQWYk0R27_1),.clk(gclk));
	jdff dff_A_T76Z3dAe3_1(.dout(w_dff_A_uQWYk0R27_1),.din(w_dff_A_T76Z3dAe3_1),.clk(gclk));
	jdff dff_A_S6lMnYu62_1(.dout(w_dff_A_T76Z3dAe3_1),.din(w_dff_A_S6lMnYu62_1),.clk(gclk));
	jdff dff_A_0YjlXqxJ8_1(.dout(w_dff_A_S6lMnYu62_1),.din(w_dff_A_0YjlXqxJ8_1),.clk(gclk));
	jdff dff_A_dEhNGnlV1_1(.dout(w_dff_A_0YjlXqxJ8_1),.din(w_dff_A_dEhNGnlV1_1),.clk(gclk));
	jdff dff_A_aUqhprmc4_1(.dout(w_dff_A_dEhNGnlV1_1),.din(w_dff_A_aUqhprmc4_1),.clk(gclk));
	jdff dff_A_KCQnRKxQ9_2(.dout(w_G165gat_1[2]),.din(w_dff_A_KCQnRKxQ9_2),.clk(gclk));
	jdff dff_A_q9IxyWtg4_2(.dout(w_dff_A_KCQnRKxQ9_2),.din(w_dff_A_q9IxyWtg4_2),.clk(gclk));
	jdff dff_A_3SHusknK0_2(.dout(w_dff_A_q9IxyWtg4_2),.din(w_dff_A_3SHusknK0_2),.clk(gclk));
	jdff dff_A_q559sriz3_2(.dout(w_dff_A_3SHusknK0_2),.din(w_dff_A_q559sriz3_2),.clk(gclk));
	jdff dff_A_OV83fcgm3_2(.dout(w_dff_A_q559sriz3_2),.din(w_dff_A_OV83fcgm3_2),.clk(gclk));
	jdff dff_A_2jpIlMhI6_2(.dout(w_dff_A_OV83fcgm3_2),.din(w_dff_A_2jpIlMhI6_2),.clk(gclk));
	jdff dff_A_7TkqrJOl2_2(.dout(w_dff_A_2jpIlMhI6_2),.din(w_dff_A_7TkqrJOl2_2),.clk(gclk));
	jdff dff_A_0M2689PP2_2(.dout(w_G165gat_0[2]),.din(w_dff_A_0M2689PP2_2),.clk(gclk));
	jdff dff_A_URQcZCMA3_2(.dout(w_dff_A_0M2689PP2_2),.din(w_dff_A_URQcZCMA3_2),.clk(gclk));
	jdff dff_A_lkYp9Zpr5_2(.dout(w_dff_A_URQcZCMA3_2),.din(w_dff_A_lkYp9Zpr5_2),.clk(gclk));
	jdff dff_A_JxVtyyyi3_2(.dout(w_dff_A_lkYp9Zpr5_2),.din(w_dff_A_JxVtyyyi3_2),.clk(gclk));
	jdff dff_B_yyFbo49d6_0(.din(n425),.dout(w_dff_B_yyFbo49d6_0),.clk(gclk));
	jdff dff_B_TIXSsHnR0_0(.din(w_dff_B_yyFbo49d6_0),.dout(w_dff_B_TIXSsHnR0_0),.clk(gclk));
	jdff dff_B_NXsse0kV1_0(.din(w_dff_B_TIXSsHnR0_0),.dout(w_dff_B_NXsse0kV1_0),.clk(gclk));
	jdff dff_B_yWLP7EiH7_0(.din(w_dff_B_NXsse0kV1_0),.dout(w_dff_B_yWLP7EiH7_0),.clk(gclk));
	jdff dff_B_4PMOP45N0_0(.din(w_dff_B_yWLP7EiH7_0),.dout(w_dff_B_4PMOP45N0_0),.clk(gclk));
	jdff dff_B_e7gYZnl19_0(.din(w_dff_B_4PMOP45N0_0),.dout(w_dff_B_e7gYZnl19_0),.clk(gclk));
	jdff dff_B_BUdIGe8i6_0(.din(w_dff_B_e7gYZnl19_0),.dout(w_dff_B_BUdIGe8i6_0),.clk(gclk));
	jdff dff_B_2UpF74z99_0(.din(w_dff_B_BUdIGe8i6_0),.dout(w_dff_B_2UpF74z99_0),.clk(gclk));
	jdff dff_B_oQziZTJD0_0(.din(w_dff_B_2UpF74z99_0),.dout(w_dff_B_oQziZTJD0_0),.clk(gclk));
	jdff dff_B_WOXq1yvj3_0(.din(w_dff_B_oQziZTJD0_0),.dout(w_dff_B_WOXq1yvj3_0),.clk(gclk));
	jdff dff_B_gSzxI1sk5_0(.din(n423),.dout(w_dff_B_gSzxI1sk5_0),.clk(gclk));
	jdff dff_B_Q750Mzc63_0(.din(w_dff_B_gSzxI1sk5_0),.dout(w_dff_B_Q750Mzc63_0),.clk(gclk));
	jdff dff_B_gXQZt7qG0_0(.din(n422),.dout(w_dff_B_gXQZt7qG0_0),.clk(gclk));
	jdff dff_B_P88vgw3G7_0(.din(w_dff_B_gXQZt7qG0_0),.dout(w_dff_B_P88vgw3G7_0),.clk(gclk));
	jdff dff_B_inUkwTzK7_0(.din(w_dff_B_P88vgw3G7_0),.dout(w_dff_B_inUkwTzK7_0),.clk(gclk));
	jdff dff_B_c16ODci74_0(.din(w_dff_B_inUkwTzK7_0),.dout(w_dff_B_c16ODci74_0),.clk(gclk));
	jdff dff_A_qUxQ9eR06_1(.dout(w_G96gat_0[1]),.din(w_dff_A_qUxQ9eR06_1),.clk(gclk));
	jdff dff_A_p7GWrnAN8_1(.dout(w_dff_A_qUxQ9eR06_1),.din(w_dff_A_p7GWrnAN8_1),.clk(gclk));
	jdff dff_A_PS2cKhNH5_1(.dout(w_dff_A_p7GWrnAN8_1),.din(w_dff_A_PS2cKhNH5_1),.clk(gclk));
	jdff dff_A_pWyCPHBM6_1(.dout(w_dff_A_PS2cKhNH5_1),.din(w_dff_A_pWyCPHBM6_1),.clk(gclk));
	jdff dff_A_iJQF7wRB4_1(.dout(w_dff_A_pWyCPHBM6_1),.din(w_dff_A_iJQF7wRB4_1),.clk(gclk));
	jdff dff_B_ewaCWjXU5_1(.din(G73gat),.dout(w_dff_B_ewaCWjXU5_1),.clk(gclk));
	jdff dff_A_ziZeDzT31_0(.dout(w_n121_0[0]),.din(w_dff_A_ziZeDzT31_0),.clk(gclk));
	jdff dff_A_RaHkYuxw1_0(.dout(w_n118_0[0]),.din(w_dff_A_RaHkYuxw1_0),.clk(gclk));
	jdff dff_B_ch065sgI9_0(.din(n419),.dout(w_dff_B_ch065sgI9_0),.clk(gclk));
	jdff dff_B_U00YQBUU1_0(.din(w_dff_B_ch065sgI9_0),.dout(w_dff_B_U00YQBUU1_0),.clk(gclk));
	jdff dff_B_2VWT5c7e6_0(.din(w_dff_B_U00YQBUU1_0),.dout(w_dff_B_2VWT5c7e6_0),.clk(gclk));
	jdff dff_B_8yeMtSAO4_0(.din(w_dff_B_2VWT5c7e6_0),.dout(w_dff_B_8yeMtSAO4_0),.clk(gclk));
	jdff dff_B_WmH6Gm1u3_0(.din(w_dff_B_8yeMtSAO4_0),.dout(w_dff_B_WmH6Gm1u3_0),.clk(gclk));
	jdff dff_B_P18D2B739_3(.din(G246gat),.dout(w_dff_B_P18D2B739_3),.clk(gclk));
	jdff dff_A_0DXRBDIX9_2(.dout(w_G228gat_0[2]),.din(w_dff_A_0DXRBDIX9_2),.clk(gclk));
	jdff dff_B_Kz50rcue2_3(.din(G228gat),.dout(w_dff_B_Kz50rcue2_3),.clk(gclk));
	jdff dff_B_LgDm6vuh4_3(.din(w_dff_B_Kz50rcue2_3),.dout(w_dff_B_LgDm6vuh4_3),.clk(gclk));
	jdff dff_B_4HzdEsCK4_3(.din(w_dff_B_LgDm6vuh4_3),.dout(w_dff_B_4HzdEsCK4_3),.clk(gclk));
	jdff dff_B_4tMDYC4K9_3(.din(w_dff_B_4HzdEsCK4_3),.dout(w_dff_B_4tMDYC4K9_3),.clk(gclk));
	jdff dff_B_140s6vK56_3(.din(w_dff_B_4tMDYC4K9_3),.dout(w_dff_B_140s6vK56_3),.clk(gclk));
	jdff dff_B_PH4bYPh99_3(.din(w_dff_B_140s6vK56_3),.dout(w_dff_B_PH4bYPh99_3),.clk(gclk));
	jdff dff_B_K03bJey14_3(.din(w_dff_B_PH4bYPh99_3),.dout(w_dff_B_K03bJey14_3),.clk(gclk));
	jdff dff_B_UjLH3mI44_3(.din(w_dff_B_K03bJey14_3),.dout(w_dff_B_UjLH3mI44_3),.clk(gclk));
	jdff dff_A_oQjb4of25_0(.dout(w_G219gat_0[0]),.din(w_dff_A_oQjb4of25_0),.clk(gclk));
	jdff dff_A_KxGzhUvM7_0(.dout(w_dff_A_oQjb4of25_0),.din(w_dff_A_KxGzhUvM7_0),.clk(gclk));
	jdff dff_A_U5CWkvmu4_0(.dout(w_dff_A_KxGzhUvM7_0),.din(w_dff_A_U5CWkvmu4_0),.clk(gclk));
	jdff dff_A_dx2ZBOYL5_0(.dout(w_dff_A_U5CWkvmu4_0),.din(w_dff_A_dx2ZBOYL5_0),.clk(gclk));
	jdff dff_A_7bI26hNa9_0(.dout(w_dff_A_dx2ZBOYL5_0),.din(w_dff_A_7bI26hNa9_0),.clk(gclk));
	jdff dff_A_pUS09l1f8_0(.dout(w_dff_A_7bI26hNa9_0),.din(w_dff_A_pUS09l1f8_0),.clk(gclk));
	jdff dff_A_TjJq9c1D9_0(.dout(w_dff_A_pUS09l1f8_0),.din(w_dff_A_TjJq9c1D9_0),.clk(gclk));
	jdff dff_A_TFGMO4fp7_0(.dout(w_dff_A_TjJq9c1D9_0),.din(w_dff_A_TFGMO4fp7_0),.clk(gclk));
	jdff dff_A_KSFyXSy63_1(.dout(w_G219gat_0[1]),.din(w_dff_A_KSFyXSy63_1),.clk(gclk));
	jdff dff_A_m7XBoiE86_1(.dout(w_dff_A_KSFyXSy63_1),.din(w_dff_A_m7XBoiE86_1),.clk(gclk));
	jdff dff_B_qY9kZGth2_3(.din(G219gat),.dout(w_dff_B_qY9kZGth2_3),.clk(gclk));
	jdff dff_B_OQbLd5zZ4_3(.din(w_dff_B_qY9kZGth2_3),.dout(w_dff_B_OQbLd5zZ4_3),.clk(gclk));
	jdff dff_B_G2UFY6Yt5_3(.din(w_dff_B_OQbLd5zZ4_3),.dout(w_dff_B_G2UFY6Yt5_3),.clk(gclk));
	jdff dff_B_SV42AhMi0_3(.din(w_dff_B_G2UFY6Yt5_3),.dout(w_dff_B_SV42AhMi0_3),.clk(gclk));
	jdff dff_B_qW1mf6b35_3(.din(w_dff_B_SV42AhMi0_3),.dout(w_dff_B_qW1mf6b35_3),.clk(gclk));
	jdff dff_B_YsUscIKX4_3(.din(w_dff_B_qW1mf6b35_3),.dout(w_dff_B_YsUscIKX4_3),.clk(gclk));
	jdff dff_B_Rxkon8iU2_3(.din(w_dff_B_YsUscIKX4_3),.dout(w_dff_B_Rxkon8iU2_3),.clk(gclk));
	jdff dff_B_rYQCJwdT3_3(.din(w_dff_B_Rxkon8iU2_3),.dout(w_dff_B_rYQCJwdT3_3),.clk(gclk));
	jdff dff_B_nKAgiXkD0_3(.din(w_dff_B_rYQCJwdT3_3),.dout(w_dff_B_nKAgiXkD0_3),.clk(gclk));
	jdff dff_B_z2BH0hU70_3(.din(w_dff_B_nKAgiXkD0_3),.dout(w_dff_B_z2BH0hU70_3),.clk(gclk));
	jdff dff_B_fJmceP214_1(.din(n406),.dout(w_dff_B_fJmceP214_1),.clk(gclk));
	jdff dff_B_QmXyJxHM7_1(.din(w_dff_B_fJmceP214_1),.dout(w_dff_B_QmXyJxHM7_1),.clk(gclk));
	jdff dff_B_eFDD5lIT6_1(.din(w_dff_B_QmXyJxHM7_1),.dout(w_dff_B_eFDD5lIT6_1),.clk(gclk));
	jdff dff_B_4EaAiSk57_1(.din(w_dff_B_eFDD5lIT6_1),.dout(w_dff_B_4EaAiSk57_1),.clk(gclk));
	jdff dff_B_XcNkQ3955_1(.din(w_dff_B_4EaAiSk57_1),.dout(w_dff_B_XcNkQ3955_1),.clk(gclk));
	jdff dff_B_TVyze9Fy4_1(.din(w_dff_B_XcNkQ3955_1),.dout(w_dff_B_TVyze9Fy4_1),.clk(gclk));
	jdff dff_B_ZF17TUEo5_1(.din(w_dff_B_TVyze9Fy4_1),.dout(w_dff_B_ZF17TUEo5_1),.clk(gclk));
	jdff dff_B_Ar3zaphe0_1(.din(w_dff_B_ZF17TUEo5_1),.dout(w_dff_B_Ar3zaphe0_1),.clk(gclk));
	jdff dff_B_zJD5ybiD5_1(.din(w_dff_B_Ar3zaphe0_1),.dout(w_dff_B_zJD5ybiD5_1),.clk(gclk));
	jdff dff_B_ZHTnix634_1(.din(n407),.dout(w_dff_B_ZHTnix634_1),.clk(gclk));
	jdff dff_B_4SqrJTfl3_1(.din(w_dff_B_ZHTnix634_1),.dout(w_dff_B_4SqrJTfl3_1),.clk(gclk));
	jdff dff_B_PFjDtg4p9_1(.din(w_dff_B_4SqrJTfl3_1),.dout(w_dff_B_PFjDtg4p9_1),.clk(gclk));
	jdff dff_B_umwW1L8p1_1(.din(w_dff_B_PFjDtg4p9_1),.dout(w_dff_B_umwW1L8p1_1),.clk(gclk));
	jdff dff_B_aLqQkBwY6_1(.din(w_dff_B_umwW1L8p1_1),.dout(w_dff_B_aLqQkBwY6_1),.clk(gclk));
	jdff dff_B_1NpAaQFN7_1(.din(w_dff_B_aLqQkBwY6_1),.dout(w_dff_B_1NpAaQFN7_1),.clk(gclk));
	jdff dff_B_iItLI2ul9_1(.din(w_dff_B_1NpAaQFN7_1),.dout(w_dff_B_iItLI2ul9_1),.clk(gclk));
	jdff dff_B_2iVXjyDC6_1(.din(w_dff_B_iItLI2ul9_1),.dout(w_dff_B_2iVXjyDC6_1),.clk(gclk));
	jdff dff_B_Ta0E71Dt8_0(.din(n408),.dout(w_dff_B_Ta0E71Dt8_0),.clk(gclk));
	jdff dff_B_GiH63RCn7_0(.din(w_dff_B_Ta0E71Dt8_0),.dout(w_dff_B_GiH63RCn7_0),.clk(gclk));
	jdff dff_B_Oi1XeFGe5_0(.din(w_dff_B_GiH63RCn7_0),.dout(w_dff_B_Oi1XeFGe5_0),.clk(gclk));
	jdff dff_B_eZYDo9mQ2_0(.din(w_dff_B_Oi1XeFGe5_0),.dout(w_dff_B_eZYDo9mQ2_0),.clk(gclk));
	jdff dff_B_ysGrVblS0_0(.din(w_dff_B_eZYDo9mQ2_0),.dout(w_dff_B_ysGrVblS0_0),.clk(gclk));
	jdff dff_B_Mf2Gmwc63_0(.din(w_dff_B_ysGrVblS0_0),.dout(w_dff_B_Mf2Gmwc63_0),.clk(gclk));
	jdff dff_B_Zzqx5ko26_0(.din(w_dff_B_Mf2Gmwc63_0),.dout(w_dff_B_Zzqx5ko26_0),.clk(gclk));
	jdff dff_A_kap8HMGd4_0(.dout(w_n329_0[0]),.din(w_dff_A_kap8HMGd4_0),.clk(gclk));
	jdff dff_A_uJK28g8t6_0(.dout(w_dff_A_kap8HMGd4_0),.din(w_dff_A_uJK28g8t6_0),.clk(gclk));
	jdff dff_A_hS4ktZtB8_0(.dout(w_dff_A_uJK28g8t6_0),.din(w_dff_A_hS4ktZtB8_0),.clk(gclk));
	jdff dff_A_8i1GiwGN4_0(.dout(w_dff_A_hS4ktZtB8_0),.din(w_dff_A_8i1GiwGN4_0),.clk(gclk));
	jdff dff_A_Dq02Xrdc6_0(.dout(w_dff_A_8i1GiwGN4_0),.din(w_dff_A_Dq02Xrdc6_0),.clk(gclk));
	jdff dff_A_gs9QbbYH8_0(.dout(w_dff_A_Dq02Xrdc6_0),.din(w_dff_A_gs9QbbYH8_0),.clk(gclk));
	jdff dff_A_VNpFfYvM2_0(.dout(w_dff_A_gs9QbbYH8_0),.din(w_dff_A_VNpFfYvM2_0),.clk(gclk));
	jdff dff_A_R4JOrNwX5_0(.dout(w_G177gat_2[0]),.din(w_dff_A_R4JOrNwX5_0),.clk(gclk));
	jdff dff_A_U6uXdiMU8_0(.dout(w_dff_A_R4JOrNwX5_0),.din(w_dff_A_U6uXdiMU8_0),.clk(gclk));
	jdff dff_A_RSAXALUE6_0(.dout(w_dff_A_U6uXdiMU8_0),.din(w_dff_A_RSAXALUE6_0),.clk(gclk));
	jdff dff_A_o2mseczl8_0(.dout(w_dff_A_RSAXALUE6_0),.din(w_dff_A_o2mseczl8_0),.clk(gclk));
	jdff dff_A_SEgK1xpa1_0(.dout(w_dff_A_o2mseczl8_0),.din(w_dff_A_SEgK1xpa1_0),.clk(gclk));
	jdff dff_A_s5KWcoQS1_0(.dout(w_dff_A_SEgK1xpa1_0),.din(w_dff_A_s5KWcoQS1_0),.clk(gclk));
	jdff dff_A_PTCrlAKa4_0(.dout(w_dff_A_s5KWcoQS1_0),.din(w_dff_A_PTCrlAKa4_0),.clk(gclk));
	jdff dff_B_8rJVeBf71_1(.din(n343),.dout(w_dff_B_8rJVeBf71_1),.clk(gclk));
	jdff dff_B_j52NSK681_1(.din(w_dff_B_8rJVeBf71_1),.dout(w_dff_B_j52NSK681_1),.clk(gclk));
	jdff dff_B_i0BDKuiQ0_1(.din(w_dff_B_j52NSK681_1),.dout(w_dff_B_i0BDKuiQ0_1),.clk(gclk));
	jdff dff_B_4cjapgEs7_1(.din(w_dff_B_i0BDKuiQ0_1),.dout(w_dff_B_4cjapgEs7_1),.clk(gclk));
	jdff dff_B_TXmJT4UW2_1(.din(w_dff_B_4cjapgEs7_1),.dout(w_dff_B_TXmJT4UW2_1),.clk(gclk));
	jdff dff_B_ZtESkSFn5_1(.din(n344),.dout(w_dff_B_ZtESkSFn5_1),.clk(gclk));
	jdff dff_B_PhMd6PAC4_1(.din(w_dff_B_ZtESkSFn5_1),.dout(w_dff_B_PhMd6PAC4_1),.clk(gclk));
	jdff dff_B_GqeoQfkK0_1(.din(w_dff_B_PhMd6PAC4_1),.dout(w_dff_B_GqeoQfkK0_1),.clk(gclk));
	jdff dff_B_VkeglazP1_1(.din(w_dff_B_GqeoQfkK0_1),.dout(w_dff_B_VkeglazP1_1),.clk(gclk));
	jdff dff_B_AGYNsHQ40_0(.din(n231),.dout(w_dff_B_AGYNsHQ40_0),.clk(gclk));
	jdff dff_A_QY1RKPjN8_0(.dout(w_n230_0[0]),.din(w_dff_A_QY1RKPjN8_0),.clk(gclk));
	jdff dff_B_oKHxCJyl8_1(.din(n227),.dout(w_dff_B_oKHxCJyl8_1),.clk(gclk));
	jdff dff_A_gzShykAk1_0(.dout(w_n228_0[0]),.din(w_dff_A_gzShykAk1_0),.clk(gclk));
	jdff dff_A_QMTfVDiR1_0(.dout(w_dff_A_gzShykAk1_0),.din(w_dff_A_QMTfVDiR1_0),.clk(gclk));
	jdff dff_A_9Lkwfsre6_0(.dout(w_dff_A_QMTfVDiR1_0),.din(w_dff_A_9Lkwfsre6_0),.clk(gclk));
	jdff dff_A_yEADm3ZI5_1(.dout(w_G195gat_1[1]),.din(w_dff_A_yEADm3ZI5_1),.clk(gclk));
	jdff dff_A_s9XObmOD2_1(.dout(w_dff_A_yEADm3ZI5_1),.din(w_dff_A_s9XObmOD2_1),.clk(gclk));
	jdff dff_A_UffxUXah3_1(.dout(w_dff_A_s9XObmOD2_1),.din(w_dff_A_UffxUXah3_1),.clk(gclk));
	jdff dff_A_DJr3SYUW9_1(.dout(w_dff_A_UffxUXah3_1),.din(w_dff_A_DJr3SYUW9_1),.clk(gclk));
	jdff dff_A_Pu6abALy1_1(.dout(w_dff_A_DJr3SYUW9_1),.din(w_dff_A_Pu6abALy1_1),.clk(gclk));
	jdff dff_A_ydeSI1L21_1(.dout(w_dff_A_Pu6abALy1_1),.din(w_dff_A_ydeSI1L21_1),.clk(gclk));
	jdff dff_A_ElakrV2A5_1(.dout(w_dff_A_ydeSI1L21_1),.din(w_dff_A_ElakrV2A5_1),.clk(gclk));
	jdff dff_A_2cjpNXO87_1(.dout(w_dff_A_ElakrV2A5_1),.din(w_dff_A_2cjpNXO87_1),.clk(gclk));
	jdff dff_A_mIwPmc5u6_2(.dout(w_G195gat_1[2]),.din(w_dff_A_mIwPmc5u6_2),.clk(gclk));
	jdff dff_A_gOLB3rRu6_2(.dout(w_dff_A_mIwPmc5u6_2),.din(w_dff_A_gOLB3rRu6_2),.clk(gclk));
	jdff dff_A_sWud1j4Y0_2(.dout(w_dff_A_gOLB3rRu6_2),.din(w_dff_A_sWud1j4Y0_2),.clk(gclk));
	jdff dff_A_6QEMRrhw2_2(.dout(w_dff_A_sWud1j4Y0_2),.din(w_dff_A_6QEMRrhw2_2),.clk(gclk));
	jdff dff_A_yE7BqAgf8_2(.dout(w_dff_A_6QEMRrhw2_2),.din(w_dff_A_yE7BqAgf8_2),.clk(gclk));
	jdff dff_A_Aq3CPh3H7_2(.dout(w_dff_A_yE7BqAgf8_2),.din(w_dff_A_Aq3CPh3H7_2),.clk(gclk));
	jdff dff_A_4GZ83DDk1_2(.dout(w_dff_A_Aq3CPh3H7_2),.din(w_dff_A_4GZ83DDk1_2),.clk(gclk));
	jdff dff_A_Tk84Qdly2_2(.dout(w_dff_A_4GZ83DDk1_2),.din(w_dff_A_Tk84Qdly2_2),.clk(gclk));
	jdff dff_A_bUrEAGsK5_1(.dout(w_G189gat_1[1]),.din(w_dff_A_bUrEAGsK5_1),.clk(gclk));
	jdff dff_A_ehd9gxtr1_1(.dout(w_dff_A_bUrEAGsK5_1),.din(w_dff_A_ehd9gxtr1_1),.clk(gclk));
	jdff dff_A_prgsGZBy1_1(.dout(w_dff_A_ehd9gxtr1_1),.din(w_dff_A_prgsGZBy1_1),.clk(gclk));
	jdff dff_A_pEyQRMFm9_1(.dout(w_dff_A_prgsGZBy1_1),.din(w_dff_A_pEyQRMFm9_1),.clk(gclk));
	jdff dff_A_uJTE1h3o9_1(.dout(w_dff_A_pEyQRMFm9_1),.din(w_dff_A_uJTE1h3o9_1),.clk(gclk));
	jdff dff_A_8ZlUDxPu3_1(.dout(w_dff_A_uJTE1h3o9_1),.din(w_dff_A_8ZlUDxPu3_1),.clk(gclk));
	jdff dff_A_6o1fz2mx1_1(.dout(w_dff_A_8ZlUDxPu3_1),.din(w_dff_A_6o1fz2mx1_1),.clk(gclk));
	jdff dff_A_5UNrjDdz5_1(.dout(w_dff_A_6o1fz2mx1_1),.din(w_dff_A_5UNrjDdz5_1),.clk(gclk));
	jdff dff_A_SyNsnOxU5_2(.dout(w_G189gat_1[2]),.din(w_dff_A_SyNsnOxU5_2),.clk(gclk));
	jdff dff_A_V3fCSbYc7_2(.dout(w_dff_A_SyNsnOxU5_2),.din(w_dff_A_V3fCSbYc7_2),.clk(gclk));
	jdff dff_A_QwUCHtfL3_2(.dout(w_dff_A_V3fCSbYc7_2),.din(w_dff_A_QwUCHtfL3_2),.clk(gclk));
	jdff dff_A_eRq5pqKb6_2(.dout(w_dff_A_QwUCHtfL3_2),.din(w_dff_A_eRq5pqKb6_2),.clk(gclk));
	jdff dff_A_arRvqP0e4_2(.dout(w_dff_A_eRq5pqKb6_2),.din(w_dff_A_arRvqP0e4_2),.clk(gclk));
	jdff dff_A_UuNH3cPQ9_2(.dout(w_dff_A_arRvqP0e4_2),.din(w_dff_A_UuNH3cPQ9_2),.clk(gclk));
	jdff dff_A_G37BWPzY1_2(.dout(w_dff_A_UuNH3cPQ9_2),.din(w_dff_A_G37BWPzY1_2),.clk(gclk));
	jdff dff_A_wLIgF7JD4_2(.dout(w_dff_A_G37BWPzY1_2),.din(w_dff_A_wLIgF7JD4_2),.clk(gclk));
	jdff dff_B_NblQoCvy0_0(.din(n225),.dout(w_dff_B_NblQoCvy0_0),.clk(gclk));
	jdff dff_A_P4A3xGbv7_0(.dout(w_n224_0[0]),.din(w_dff_A_P4A3xGbv7_0),.clk(gclk));
	jdff dff_A_mARZLVck7_0(.dout(w_n223_0[0]),.din(w_dff_A_mARZLVck7_0),.clk(gclk));
	jdff dff_A_xsDiUmav4_0(.dout(w_dff_A_mARZLVck7_0),.din(w_dff_A_xsDiUmav4_0),.clk(gclk));
	jdff dff_B_Y91cRz3S3_1(.din(n219),.dout(w_dff_B_Y91cRz3S3_1),.clk(gclk));
	jdff dff_A_7v4YJTJZ3_0(.dout(w_G121gat_0[0]),.din(w_dff_A_7v4YJTJZ3_0),.clk(gclk));
	jdff dff_A_rD5nbX0R4_0(.dout(w_dff_A_7v4YJTJZ3_0),.din(w_dff_A_rD5nbX0R4_0),.clk(gclk));
	jdff dff_A_leEiRrE34_0(.dout(w_dff_A_rD5nbX0R4_0),.din(w_dff_A_leEiRrE34_0),.clk(gclk));
	jdff dff_A_oB26pOZI7_0(.dout(w_dff_A_leEiRrE34_0),.din(w_dff_A_oB26pOZI7_0),.clk(gclk));
	jdff dff_A_IsZfT29g9_0(.dout(w_dff_A_oB26pOZI7_0),.din(w_dff_A_IsZfT29g9_0),.clk(gclk));
	jdff dff_A_CRBlKU8z2_0(.dout(w_G195gat_2[0]),.din(w_dff_A_CRBlKU8z2_0),.clk(gclk));
	jdff dff_A_6zm24qyD0_0(.dout(w_dff_A_CRBlKU8z2_0),.din(w_dff_A_6zm24qyD0_0),.clk(gclk));
	jdff dff_A_Za1CKhsi4_0(.dout(w_dff_A_6zm24qyD0_0),.din(w_dff_A_Za1CKhsi4_0),.clk(gclk));
	jdff dff_A_IjWelpfO1_0(.dout(w_dff_A_Za1CKhsi4_0),.din(w_dff_A_IjWelpfO1_0),.clk(gclk));
	jdff dff_A_dJS1UTvR7_0(.dout(w_dff_A_IjWelpfO1_0),.din(w_dff_A_dJS1UTvR7_0),.clk(gclk));
	jdff dff_A_Yz8mIEtH6_0(.dout(w_dff_A_dJS1UTvR7_0),.din(w_dff_A_Yz8mIEtH6_0),.clk(gclk));
	jdff dff_A_FyBZqUeG8_0(.dout(w_dff_A_Yz8mIEtH6_0),.din(w_dff_A_FyBZqUeG8_0),.clk(gclk));
	jdff dff_A_XMcUX3AP0_0(.dout(w_dff_A_FyBZqUeG8_0),.din(w_dff_A_XMcUX3AP0_0),.clk(gclk));
	jdff dff_A_dG0yYy4j0_2(.dout(w_G195gat_0[2]),.din(w_dff_A_dG0yYy4j0_2),.clk(gclk));
	jdff dff_A_rQcTeXgG2_2(.dout(w_dff_A_dG0yYy4j0_2),.din(w_dff_A_rQcTeXgG2_2),.clk(gclk));
	jdff dff_A_4Kmdv6234_2(.dout(w_dff_A_rQcTeXgG2_2),.din(w_dff_A_4Kmdv6234_2),.clk(gclk));
	jdff dff_A_8fG1lPkj0_2(.dout(w_dff_A_4Kmdv6234_2),.din(w_dff_A_8fG1lPkj0_2),.clk(gclk));
	jdff dff_B_eenTpDDo4_1(.din(n214),.dout(w_dff_B_eenTpDDo4_1),.clk(gclk));
	jdff dff_A_EcDp1A0e3_1(.dout(w_G116gat_0[1]),.din(w_dff_A_EcDp1A0e3_1),.clk(gclk));
	jdff dff_A_BAnzpPqS4_1(.dout(w_dff_A_EcDp1A0e3_1),.din(w_dff_A_BAnzpPqS4_1),.clk(gclk));
	jdff dff_A_E7TWcOqN9_1(.dout(w_dff_A_BAnzpPqS4_1),.din(w_dff_A_E7TWcOqN9_1),.clk(gclk));
	jdff dff_A_ihDrd5km5_1(.dout(w_dff_A_E7TWcOqN9_1),.din(w_dff_A_ihDrd5km5_1),.clk(gclk));
	jdff dff_A_s4lNmvvS8_1(.dout(w_dff_A_ihDrd5km5_1),.din(w_dff_A_s4lNmvvS8_1),.clk(gclk));
	jdff dff_A_Utnvb7700_1(.dout(w_G146gat_0[1]),.din(w_dff_A_Utnvb7700_1),.clk(gclk));
	jdff dff_B_T9mntcNv1_2(.din(G146gat),.dout(w_dff_B_T9mntcNv1_2),.clk(gclk));
	jdff dff_B_wW0G0AWt7_2(.din(w_dff_B_T9mntcNv1_2),.dout(w_dff_B_wW0G0AWt7_2),.clk(gclk));
	jdff dff_B_2S2tHoPe4_2(.din(w_dff_B_wW0G0AWt7_2),.dout(w_dff_B_2S2tHoPe4_2),.clk(gclk));
	jdff dff_B_RUCXEpUo8_2(.din(w_dff_B_2S2tHoPe4_2),.dout(w_dff_B_RUCXEpUo8_2),.clk(gclk));
	jdff dff_A_PBwWq9Ye3_0(.dout(w_G189gat_2[0]),.din(w_dff_A_PBwWq9Ye3_0),.clk(gclk));
	jdff dff_A_pHgR9PWW7_0(.dout(w_dff_A_PBwWq9Ye3_0),.din(w_dff_A_pHgR9PWW7_0),.clk(gclk));
	jdff dff_A_tlyHrYGw4_0(.dout(w_dff_A_pHgR9PWW7_0),.din(w_dff_A_tlyHrYGw4_0),.clk(gclk));
	jdff dff_A_Tinws3kd7_0(.dout(w_dff_A_tlyHrYGw4_0),.din(w_dff_A_Tinws3kd7_0),.clk(gclk));
	jdff dff_A_NmpuEUa86_0(.dout(w_dff_A_Tinws3kd7_0),.din(w_dff_A_NmpuEUa86_0),.clk(gclk));
	jdff dff_A_K3N3Zj0k7_0(.dout(w_dff_A_NmpuEUa86_0),.din(w_dff_A_K3N3Zj0k7_0),.clk(gclk));
	jdff dff_A_s1QoyaYE4_0(.dout(w_dff_A_K3N3Zj0k7_0),.din(w_dff_A_s1QoyaYE4_0),.clk(gclk));
	jdff dff_A_F0P8hhOf4_0(.dout(w_dff_A_s1QoyaYE4_0),.din(w_dff_A_F0P8hhOf4_0),.clk(gclk));
	jdff dff_A_HuTQ1mql8_2(.dout(w_G189gat_0[2]),.din(w_dff_A_HuTQ1mql8_2),.clk(gclk));
	jdff dff_A_jSXmu9qJ3_2(.dout(w_dff_A_HuTQ1mql8_2),.din(w_dff_A_jSXmu9qJ3_2),.clk(gclk));
	jdff dff_A_ZEKpD2X67_2(.dout(w_dff_A_jSXmu9qJ3_2),.din(w_dff_A_ZEKpD2X67_2),.clk(gclk));
	jdff dff_A_PhIG9if66_2(.dout(w_dff_A_ZEKpD2X67_2),.din(w_dff_A_PhIG9if66_2),.clk(gclk));
	jdff dff_B_rRFD66SL8_1(.din(n197),.dout(w_dff_B_rRFD66SL8_1),.clk(gclk));
	jdff dff_B_23pPR6AI7_1(.din(n198),.dout(w_dff_B_23pPR6AI7_1),.clk(gclk));
	jdff dff_B_FJZYVjBF8_1(.din(w_dff_B_23pPR6AI7_1),.dout(w_dff_B_FJZYVjBF8_1),.clk(gclk));
	jdff dff_B_WdfitJyc1_1(.din(w_dff_B_FJZYVjBF8_1),.dout(w_dff_B_WdfitJyc1_1),.clk(gclk));
	jdff dff_B_6xEaZtyY8_1(.din(w_dff_B_WdfitJyc1_1),.dout(w_dff_B_6xEaZtyY8_1),.clk(gclk));
	jdff dff_B_yNef5tfK2_1(.din(w_dff_B_6xEaZtyY8_1),.dout(w_dff_B_yNef5tfK2_1),.clk(gclk));
	jdff dff_B_heYskH6L4_1(.din(w_dff_B_yNef5tfK2_1),.dout(w_dff_B_heYskH6L4_1),.clk(gclk));
	jdff dff_B_IJ6JFvqV3_1(.din(w_dff_B_heYskH6L4_1),.dout(w_dff_B_IJ6JFvqV3_1),.clk(gclk));
	jdff dff_B_VhjGV70K6_1(.din(w_dff_B_IJ6JFvqV3_1),.dout(w_dff_B_VhjGV70K6_1),.clk(gclk));
	jdff dff_B_LtJRveWy4_1(.din(n199),.dout(w_dff_B_LtJRveWy4_1),.clk(gclk));
	jdff dff_B_tp0AYuUa2_0(.din(n208),.dout(w_dff_B_tp0AYuUa2_0),.clk(gclk));
	jdff dff_B_GxaiRH1j7_0(.din(w_dff_B_tp0AYuUa2_0),.dout(w_dff_B_GxaiRH1j7_0),.clk(gclk));
	jdff dff_B_2LNkqAIQ2_1(.din(n200),.dout(w_dff_B_2LNkqAIQ2_1),.clk(gclk));
	jdff dff_B_tDCpdrd55_1(.din(w_dff_B_2LNkqAIQ2_1),.dout(w_dff_B_tDCpdrd55_1),.clk(gclk));
	jdff dff_B_9Y1OM4CG8_1(.din(w_dff_B_tDCpdrd55_1),.dout(w_dff_B_9Y1OM4CG8_1),.clk(gclk));
	jdff dff_B_5ATfsu0t5_1(.din(w_dff_B_9Y1OM4CG8_1),.dout(w_dff_B_5ATfsu0t5_1),.clk(gclk));
	jdff dff_B_yTizZ9lw6_1(.din(w_dff_B_5ATfsu0t5_1),.dout(w_dff_B_yTizZ9lw6_1),.clk(gclk));
	jdff dff_B_9Z2GTdBA3_1(.din(n201),.dout(w_dff_B_9Z2GTdBA3_1),.clk(gclk));
	jdff dff_B_PIH3NLKl1_1(.din(w_dff_B_9Z2GTdBA3_1),.dout(w_dff_B_PIH3NLKl1_1),.clk(gclk));
	jdff dff_B_QMDI3G081_1(.din(w_dff_B_PIH3NLKl1_1),.dout(w_dff_B_QMDI3G081_1),.clk(gclk));
	jdff dff_B_a3dEcDtW3_1(.din(n202),.dout(w_dff_B_a3dEcDtW3_1),.clk(gclk));
	jdff dff_B_FSuwRInr5_2(.din(n143),.dout(w_dff_B_FSuwRInr5_2),.clk(gclk));
	jdff dff_B_rwbBHnH30_2(.din(w_dff_B_FSuwRInr5_2),.dout(w_dff_B_rwbBHnH30_2),.clk(gclk));
	jdff dff_B_uDz6Pol31_2(.din(w_dff_B_rwbBHnH30_2),.dout(w_dff_B_uDz6Pol31_2),.clk(gclk));
	jdff dff_B_bEuC7WNx2_2(.din(w_dff_B_uDz6Pol31_2),.dout(w_dff_B_bEuC7WNx2_2),.clk(gclk));
	jdff dff_B_MzMoJbgy6_2(.din(w_dff_B_bEuC7WNx2_2),.dout(w_dff_B_MzMoJbgy6_2),.clk(gclk));
	jdff dff_B_TkhH7ngz6_2(.din(w_dff_B_MzMoJbgy6_2),.dout(w_dff_B_TkhH7ngz6_2),.clk(gclk));
	jdff dff_B_Ae9ugOcq8_2(.din(w_dff_B_TkhH7ngz6_2),.dout(w_dff_B_Ae9ugOcq8_2),.clk(gclk));
	jdff dff_B_PUmuuksv1_2(.din(w_dff_B_Ae9ugOcq8_2),.dout(w_dff_B_PUmuuksv1_2),.clk(gclk));
	jdff dff_B_Ef3RQZoT8_2(.din(w_dff_B_PUmuuksv1_2),.dout(w_dff_B_Ef3RQZoT8_2),.clk(gclk));
	jdff dff_A_9oXkUTAz9_0(.dout(w_G261gat_0[0]),.din(w_dff_A_9oXkUTAz9_0),.clk(gclk));
	jdff dff_A_wk1SUM0p8_0(.dout(w_dff_A_9oXkUTAz9_0),.din(w_dff_A_wk1SUM0p8_0),.clk(gclk));
	jdff dff_A_UEIPtOM79_0(.dout(w_dff_A_wk1SUM0p8_0),.din(w_dff_A_UEIPtOM79_0),.clk(gclk));
	jdff dff_A_SVW2ApoK0_0(.dout(w_dff_A_UEIPtOM79_0),.din(w_dff_A_SVW2ApoK0_0),.clk(gclk));
	jdff dff_A_hZAmTO0x5_0(.dout(w_dff_A_SVW2ApoK0_0),.din(w_dff_A_hZAmTO0x5_0),.clk(gclk));
	jdff dff_A_gfX8I5vR0_0(.dout(w_dff_A_hZAmTO0x5_0),.din(w_dff_A_gfX8I5vR0_0),.clk(gclk));
	jdff dff_A_qlmLcpAJ4_0(.dout(w_dff_A_gfX8I5vR0_0),.din(w_dff_A_qlmLcpAJ4_0),.clk(gclk));
	jdff dff_A_b5D8cxwH4_0(.dout(w_dff_A_qlmLcpAJ4_0),.din(w_dff_A_b5D8cxwH4_0),.clk(gclk));
	jdff dff_A_olrTfMMo1_0(.dout(w_dff_A_b5D8cxwH4_0),.din(w_dff_A_olrTfMMo1_0),.clk(gclk));
	jdff dff_A_kPOlzqhg9_1(.dout(w_G261gat_0[1]),.din(w_dff_A_kPOlzqhg9_1),.clk(gclk));
	jdff dff_A_CVsh6Tod2_1(.dout(w_dff_A_kPOlzqhg9_1),.din(w_dff_A_CVsh6Tod2_1),.clk(gclk));
	jdff dff_A_pHweGRNG9_1(.dout(w_dff_A_CVsh6Tod2_1),.din(w_dff_A_pHweGRNG9_1),.clk(gclk));
	jdff dff_A_l3yf2L599_1(.dout(w_dff_A_pHweGRNG9_1),.din(w_dff_A_l3yf2L599_1),.clk(gclk));
	jdff dff_A_GeyWpXcm2_1(.dout(w_dff_A_l3yf2L599_1),.din(w_dff_A_GeyWpXcm2_1),.clk(gclk));
	jdff dff_A_9032q7DC3_1(.dout(w_dff_A_GeyWpXcm2_1),.din(w_dff_A_9032q7DC3_1),.clk(gclk));
	jdff dff_A_Xu3zxC3c8_1(.dout(w_dff_A_9032q7DC3_1),.din(w_dff_A_Xu3zxC3c8_1),.clk(gclk));
	jdff dff_A_yUHVYSVi6_1(.dout(w_dff_A_Xu3zxC3c8_1),.din(w_dff_A_yUHVYSVi6_1),.clk(gclk));
	jdff dff_A_VDf97yrT4_1(.dout(w_dff_A_yUHVYSVi6_1),.din(w_dff_A_VDf97yrT4_1),.clk(gclk));
	jdff dff_A_djOBsNTk8_0(.dout(w_n196_0[0]),.din(w_dff_A_djOBsNTk8_0),.clk(gclk));
	jdff dff_A_MeVNwU9y6_1(.dout(w_n154_0[1]),.din(w_dff_A_MeVNwU9y6_1),.clk(gclk));
	jdff dff_A_W3FLjjEm2_0(.dout(w_G126gat_0[0]),.din(w_dff_A_W3FLjjEm2_0),.clk(gclk));
	jdff dff_A_fUIRF1uh8_0(.dout(w_dff_A_W3FLjjEm2_0),.din(w_dff_A_fUIRF1uh8_0),.clk(gclk));
	jdff dff_A_jijkFqLL6_0(.dout(w_dff_A_fUIRF1uh8_0),.din(w_dff_A_jijkFqLL6_0),.clk(gclk));
	jdff dff_A_SXSa9Abc2_0(.dout(w_dff_A_jijkFqLL6_0),.din(w_dff_A_SXSa9Abc2_0),.clk(gclk));
	jdff dff_A_kj7LiY6u0_0(.dout(w_dff_A_SXSa9Abc2_0),.din(w_dff_A_kj7LiY6u0_0),.clk(gclk));
	jdff dff_A_Hjd5HB6V7_1(.dout(w_G201gat_1[1]),.din(w_dff_A_Hjd5HB6V7_1),.clk(gclk));
	jdff dff_A_1KrbjPmR9_1(.dout(w_dff_A_Hjd5HB6V7_1),.din(w_dff_A_1KrbjPmR9_1),.clk(gclk));
	jdff dff_A_qM5UkkSD5_1(.dout(w_dff_A_1KrbjPmR9_1),.din(w_dff_A_qM5UkkSD5_1),.clk(gclk));
	jdff dff_A_QzOt0Dxq5_1(.dout(w_dff_A_qM5UkkSD5_1),.din(w_dff_A_QzOt0Dxq5_1),.clk(gclk));
	jdff dff_A_9lvKOKTJ5_1(.dout(w_dff_A_QzOt0Dxq5_1),.din(w_dff_A_9lvKOKTJ5_1),.clk(gclk));
	jdff dff_A_nrpS9ytr7_1(.dout(w_dff_A_9lvKOKTJ5_1),.din(w_dff_A_nrpS9ytr7_1),.clk(gclk));
	jdff dff_A_jUu6GTGU5_1(.dout(w_dff_A_nrpS9ytr7_1),.din(w_dff_A_jUu6GTGU5_1),.clk(gclk));
	jdff dff_A_zEIzOYzO8_1(.dout(w_dff_A_jUu6GTGU5_1),.din(w_dff_A_zEIzOYzO8_1),.clk(gclk));
	jdff dff_A_LWe7mISb3_2(.dout(w_G201gat_1[2]),.din(w_dff_A_LWe7mISb3_2),.clk(gclk));
	jdff dff_A_gI9avPq63_2(.dout(w_dff_A_LWe7mISb3_2),.din(w_dff_A_gI9avPq63_2),.clk(gclk));
	jdff dff_A_anHXxQlP3_2(.dout(w_dff_A_gI9avPq63_2),.din(w_dff_A_anHXxQlP3_2),.clk(gclk));
	jdff dff_A_L2PRPBEx7_2(.dout(w_dff_A_anHXxQlP3_2),.din(w_dff_A_L2PRPBEx7_2),.clk(gclk));
	jdff dff_A_Jr0aNAZ54_2(.dout(w_G201gat_0[2]),.din(w_dff_A_Jr0aNAZ54_2),.clk(gclk));
	jdff dff_A_kgqIfa3Q5_2(.dout(w_dff_A_Jr0aNAZ54_2),.din(w_dff_A_kgqIfa3Q5_2),.clk(gclk));
	jdff dff_A_XzTdvpy37_2(.dout(w_dff_A_kgqIfa3Q5_2),.din(w_dff_A_XzTdvpy37_2),.clk(gclk));
	jdff dff_A_kSeB5CQy5_2(.dout(w_dff_A_XzTdvpy37_2),.din(w_dff_A_kSeB5CQy5_2),.clk(gclk));
	jdff dff_A_jcTRIs114_2(.dout(w_dff_A_kSeB5CQy5_2),.din(w_dff_A_jcTRIs114_2),.clk(gclk));
	jdff dff_A_1GLIPFkh8_2(.dout(w_dff_A_jcTRIs114_2),.din(w_dff_A_1GLIPFkh8_2),.clk(gclk));
	jdff dff_A_DGiQDqBx1_2(.dout(w_dff_A_1GLIPFkh8_2),.din(w_dff_A_DGiQDqBx1_2),.clk(gclk));
	jdff dff_A_pdf0eo104_2(.dout(w_dff_A_DGiQDqBx1_2),.din(w_dff_A_pdf0eo104_2),.clk(gclk));
	jdff dff_A_mfbB0nMc5_1(.dout(w_n303_0[1]),.din(w_dff_A_mfbB0nMc5_1),.clk(gclk));
	jdff dff_A_kbszwEzd6_1(.dout(w_dff_A_mfbB0nMc5_1),.din(w_dff_A_kbszwEzd6_1),.clk(gclk));
	jdff dff_A_TOf5ODXz5_1(.dout(w_dff_A_kbszwEzd6_1),.din(w_dff_A_TOf5ODXz5_1),.clk(gclk));
	jdff dff_A_YURtj78C0_1(.dout(w_dff_A_TOf5ODXz5_1),.din(w_dff_A_YURtj78C0_1),.clk(gclk));
	jdff dff_A_sZsdzTaB7_1(.dout(w_n302_0[1]),.din(w_dff_A_sZsdzTaB7_1),.clk(gclk));
	jdff dff_A_0zPqIFrs3_1(.dout(w_dff_A_sZsdzTaB7_1),.din(w_dff_A_0zPqIFrs3_1),.clk(gclk));
	jdff dff_A_F9C2ZxEi1_1(.dout(w_dff_A_0zPqIFrs3_1),.din(w_dff_A_F9C2ZxEi1_1),.clk(gclk));
	jdff dff_A_86cfAmWR2_1(.dout(w_dff_A_F9C2ZxEi1_1),.din(w_dff_A_86cfAmWR2_1),.clk(gclk));
	jdff dff_A_BCpoGdPS7_1(.dout(w_dff_A_86cfAmWR2_1),.din(w_dff_A_BCpoGdPS7_1),.clk(gclk));
	jdff dff_B_rOE8WGvz2_1(.din(n190),.dout(w_dff_B_rOE8WGvz2_1),.clk(gclk));
	jdff dff_A_JZ7jqKdK4_1(.dout(w_G111gat_0[1]),.din(w_dff_A_JZ7jqKdK4_1),.clk(gclk));
	jdff dff_A_EjSzGy6S4_1(.dout(w_dff_A_JZ7jqKdK4_1),.din(w_dff_A_EjSzGy6S4_1),.clk(gclk));
	jdff dff_A_7b2uoo306_1(.dout(w_dff_A_EjSzGy6S4_1),.din(w_dff_A_7b2uoo306_1),.clk(gclk));
	jdff dff_A_zjJiOsop4_1(.dout(w_dff_A_7b2uoo306_1),.din(w_dff_A_zjJiOsop4_1),.clk(gclk));
	jdff dff_A_qrJOZv860_1(.dout(w_dff_A_zjJiOsop4_1),.din(w_dff_A_qrJOZv860_1),.clk(gclk));
	jdff dff_A_oEzKJrnh1_1(.dout(w_n165_1[1]),.din(w_dff_A_oEzKJrnh1_1),.clk(gclk));
	jdff dff_A_wJXMRtTS0_1(.dout(w_dff_A_oEzKJrnh1_1),.din(w_dff_A_wJXMRtTS0_1),.clk(gclk));
	jdff dff_A_VOkRqBMv5_2(.dout(w_n165_1[2]),.din(w_dff_A_VOkRqBMv5_2),.clk(gclk));
	jdff dff_A_yK5wcWlf3_2(.dout(w_dff_A_VOkRqBMv5_2),.din(w_dff_A_yK5wcWlf3_2),.clk(gclk));
	jdff dff_A_N3VGMkfp7_1(.dout(w_n165_0[1]),.din(w_dff_A_N3VGMkfp7_1),.clk(gclk));
	jdff dff_A_TypNUBOb1_1(.dout(w_dff_A_N3VGMkfp7_1),.din(w_dff_A_TypNUBOb1_1),.clk(gclk));
	jdff dff_A_ND8Jvmt28_2(.dout(w_n165_0[2]),.din(w_dff_A_ND8Jvmt28_2),.clk(gclk));
	jdff dff_A_OdzPs9rg2_2(.dout(w_dff_A_ND8Jvmt28_2),.din(w_dff_A_OdzPs9rg2_2),.clk(gclk));
	jdff dff_B_18olbLOP0_0(.din(n164),.dout(w_dff_B_18olbLOP0_0),.clk(gclk));
	jdff dff_A_KFfwWjQ50_0(.dout(w_n96_0[0]),.din(w_dff_A_KFfwWjQ50_0),.clk(gclk));
	jdff dff_A_hIL54dP46_0(.dout(w_dff_A_KFfwWjQ50_0),.din(w_dff_A_hIL54dP46_0),.clk(gclk));
	jdff dff_A_P9EaKFnE3_0(.dout(w_dff_A_hIL54dP46_0),.din(w_dff_A_P9EaKFnE3_0),.clk(gclk));
	jdff dff_A_mLdU7aep6_1(.dout(w_G143gat_0[1]),.din(w_dff_A_mLdU7aep6_1),.clk(gclk));
	jdff dff_B_CFEopYXd6_2(.din(G143gat),.dout(w_dff_B_CFEopYXd6_2),.clk(gclk));
	jdff dff_B_uU4fkVGW5_2(.din(w_dff_B_CFEopYXd6_2),.dout(w_dff_B_uU4fkVGW5_2),.clk(gclk));
	jdff dff_B_8EmUAwgh0_2(.din(w_dff_B_uU4fkVGW5_2),.dout(w_dff_B_8EmUAwgh0_2),.clk(gclk));
	jdff dff_B_B0ihQo9d3_2(.din(w_dff_B_8EmUAwgh0_2),.dout(w_dff_B_B0ihQo9d3_2),.clk(gclk));
	jdff dff_A_QYu2gx179_0(.dout(w_G183gat_1[0]),.din(w_dff_A_QYu2gx179_0),.clk(gclk));
	jdff dff_A_340dqXtv2_0(.dout(w_dff_A_QYu2gx179_0),.din(w_dff_A_340dqXtv2_0),.clk(gclk));
	jdff dff_A_D1NNrqd31_0(.dout(w_dff_A_340dqXtv2_0),.din(w_dff_A_D1NNrqd31_0),.clk(gclk));
	jdff dff_A_FPNrMZMq6_0(.dout(w_dff_A_D1NNrqd31_0),.din(w_dff_A_FPNrMZMq6_0),.clk(gclk));
	jdff dff_A_iXqca1Zk3_0(.dout(w_dff_A_FPNrMZMq6_0),.din(w_dff_A_iXqca1Zk3_0),.clk(gclk));
	jdff dff_A_aNX4dK6Y4_0(.dout(w_dff_A_iXqca1Zk3_0),.din(w_dff_A_aNX4dK6Y4_0),.clk(gclk));
	jdff dff_A_JV25cchI2_0(.dout(w_dff_A_aNX4dK6Y4_0),.din(w_dff_A_JV25cchI2_0),.clk(gclk));
	jdff dff_A_KKyrQJND4_0(.dout(w_dff_A_JV25cchI2_0),.din(w_dff_A_KKyrQJND4_0),.clk(gclk));
	jdff dff_A_n8jyaAOY5_1(.dout(w_G183gat_1[1]),.din(w_dff_A_n8jyaAOY5_1),.clk(gclk));
	jdff dff_A_pGiu4Gew8_1(.dout(w_dff_A_n8jyaAOY5_1),.din(w_dff_A_pGiu4Gew8_1),.clk(gclk));
	jdff dff_A_saBQNKzF6_1(.dout(w_dff_A_pGiu4Gew8_1),.din(w_dff_A_saBQNKzF6_1),.clk(gclk));
	jdff dff_A_1QSSEYiG4_1(.dout(w_dff_A_saBQNKzF6_1),.din(w_dff_A_1QSSEYiG4_1),.clk(gclk));
	jdff dff_A_RWnSet5j4_2(.dout(w_G183gat_0[2]),.din(w_dff_A_RWnSet5j4_2),.clk(gclk));
	jdff dff_A_LWWM06jf9_2(.dout(w_dff_A_RWnSet5j4_2),.din(w_dff_A_LWWM06jf9_2),.clk(gclk));
	jdff dff_A_dgh7e4WD9_2(.dout(w_dff_A_LWWM06jf9_2),.din(w_dff_A_dgh7e4WD9_2),.clk(gclk));
	jdff dff_A_h6RLW3107_2(.dout(w_dff_A_dgh7e4WD9_2),.din(w_dff_A_h6RLW3107_2),.clk(gclk));
	jdff dff_A_6z70m9va4_2(.dout(w_dff_A_h6RLW3107_2),.din(w_dff_A_6z70m9va4_2),.clk(gclk));
	jdff dff_A_2Jj8F1tu7_2(.dout(w_dff_A_6z70m9va4_2),.din(w_dff_A_2Jj8F1tu7_2),.clk(gclk));
	jdff dff_A_El1Nxp5O6_2(.dout(w_dff_A_2Jj8F1tu7_2),.din(w_dff_A_El1Nxp5O6_2),.clk(gclk));
	jdff dff_A_Wr5l3qB80_2(.dout(w_dff_A_El1Nxp5O6_2),.din(w_dff_A_Wr5l3qB80_2),.clk(gclk));
	jdff dff_A_25Bq4v7R0_0(.dout(w_n335_0[0]),.din(w_dff_A_25Bq4v7R0_0),.clk(gclk));
	jdff dff_A_MaDjIIkD6_0(.dout(w_dff_A_25Bq4v7R0_0),.din(w_dff_A_MaDjIIkD6_0),.clk(gclk));
	jdff dff_A_hsXq72MK2_0(.dout(w_dff_A_MaDjIIkD6_0),.din(w_dff_A_hsXq72MK2_0),.clk(gclk));
	jdff dff_A_cOGD7dtu3_0(.dout(w_dff_A_hsXq72MK2_0),.din(w_dff_A_cOGD7dtu3_0),.clk(gclk));
	jdff dff_A_dlplJRp08_0(.dout(w_dff_A_cOGD7dtu3_0),.din(w_dff_A_dlplJRp08_0),.clk(gclk));
	jdff dff_A_aCCnIhpQ0_0(.dout(w_dff_A_dlplJRp08_0),.din(w_dff_A_aCCnIhpQ0_0),.clk(gclk));
	jdff dff_A_5anbM8rR4_0(.dout(w_dff_A_aCCnIhpQ0_0),.din(w_dff_A_5anbM8rR4_0),.clk(gclk));
	jdff dff_A_wYIkLhg66_0(.dout(w_dff_A_5anbM8rR4_0),.din(w_dff_A_wYIkLhg66_0),.clk(gclk));
	jdff dff_B_ij8LaE1r7_0(.din(n325),.dout(w_dff_B_ij8LaE1r7_0),.clk(gclk));
	jdff dff_B_byONNthQ6_0(.din(w_dff_B_ij8LaE1r7_0),.dout(w_dff_B_byONNthQ6_0),.clk(gclk));
	jdff dff_B_fkJQA9hn5_0(.din(w_dff_B_byONNthQ6_0),.dout(w_dff_B_fkJQA9hn5_0),.clk(gclk));
	jdff dff_A_vQFXgHor2_0(.dout(w_G153gat_0[0]),.din(w_dff_A_vQFXgHor2_0),.clk(gclk));
	jdff dff_A_xgh1ZQUf4_0(.dout(w_dff_A_vQFXgHor2_0),.din(w_dff_A_xgh1ZQUf4_0),.clk(gclk));
	jdff dff_A_pxaxEmwM6_0(.dout(w_dff_A_xgh1ZQUf4_0),.din(w_dff_A_pxaxEmwM6_0),.clk(gclk));
	jdff dff_A_ehEewFN31_0(.dout(w_dff_A_pxaxEmwM6_0),.din(w_dff_A_ehEewFN31_0),.clk(gclk));
	jdff dff_A_CKg17ZEl4_2(.dout(w_G153gat_0[2]),.din(w_dff_A_CKg17ZEl4_2),.clk(gclk));
	jdff dff_A_B3TbiyQQ6_2(.dout(w_dff_A_CKg17ZEl4_2),.din(w_dff_A_B3TbiyQQ6_2),.clk(gclk));
	jdff dff_A_62hqqsVn3_2(.dout(w_dff_A_B3TbiyQQ6_2),.din(w_dff_A_62hqqsVn3_2),.clk(gclk));
	jdff dff_A_wlkSUAub8_2(.dout(w_dff_A_62hqqsVn3_2),.din(w_dff_A_wlkSUAub8_2),.clk(gclk));
	jdff dff_A_x5CwquCG5_2(.dout(w_dff_A_wlkSUAub8_2),.din(w_dff_A_x5CwquCG5_2),.clk(gclk));
	jdff dff_A_VquKTESQ3_0(.dout(w_G106gat_0[0]),.din(w_dff_A_VquKTESQ3_0),.clk(gclk));
	jdff dff_A_k9WQmgek1_0(.dout(w_dff_A_VquKTESQ3_0),.din(w_dff_A_k9WQmgek1_0),.clk(gclk));
	jdff dff_A_jssz4fDF0_0(.dout(w_dff_A_k9WQmgek1_0),.din(w_dff_A_jssz4fDF0_0),.clk(gclk));
	jdff dff_A_mV4frAKc3_0(.dout(w_dff_A_jssz4fDF0_0),.din(w_dff_A_mV4frAKc3_0),.clk(gclk));
	jdff dff_A_J5Vh6mSc0_0(.dout(w_dff_A_mV4frAKc3_0),.din(w_dff_A_J5Vh6mSc0_0),.clk(gclk));
	jdff dff_A_t1Rginlm8_1(.dout(w_G177gat_1[1]),.din(w_dff_A_t1Rginlm8_1),.clk(gclk));
	jdff dff_A_pWOIEiwN4_1(.dout(w_dff_A_t1Rginlm8_1),.din(w_dff_A_pWOIEiwN4_1),.clk(gclk));
	jdff dff_A_edomZr5R7_1(.dout(w_dff_A_pWOIEiwN4_1),.din(w_dff_A_edomZr5R7_1),.clk(gclk));
	jdff dff_A_O5YKIHQ91_1(.dout(w_dff_A_edomZr5R7_1),.din(w_dff_A_O5YKIHQ91_1),.clk(gclk));
	jdff dff_A_XVL3MtqC0_1(.dout(w_dff_A_O5YKIHQ91_1),.din(w_dff_A_XVL3MtqC0_1),.clk(gclk));
	jdff dff_A_0A1pbHjQ5_1(.dout(w_dff_A_XVL3MtqC0_1),.din(w_dff_A_0A1pbHjQ5_1),.clk(gclk));
	jdff dff_A_6sPlPBXq0_1(.dout(w_dff_A_0A1pbHjQ5_1),.din(w_dff_A_6sPlPBXq0_1),.clk(gclk));
	jdff dff_A_F6E0aPbK6_2(.dout(w_G177gat_1[2]),.din(w_dff_A_F6E0aPbK6_2),.clk(gclk));
	jdff dff_A_0SEFSqob5_2(.dout(w_dff_A_F6E0aPbK6_2),.din(w_dff_A_0SEFSqob5_2),.clk(gclk));
	jdff dff_A_qCHLWT0n2_2(.dout(w_dff_A_0SEFSqob5_2),.din(w_dff_A_qCHLWT0n2_2),.clk(gclk));
	jdff dff_A_DBtylpiE6_2(.dout(w_dff_A_qCHLWT0n2_2),.din(w_dff_A_DBtylpiE6_2),.clk(gclk));
	jdff dff_A_0f6e43BR3_2(.dout(w_dff_A_DBtylpiE6_2),.din(w_dff_A_0f6e43BR3_2),.clk(gclk));
	jdff dff_A_L3hODdFd9_2(.dout(w_dff_A_0f6e43BR3_2),.din(w_dff_A_L3hODdFd9_2),.clk(gclk));
	jdff dff_A_VvwERKv35_2(.dout(w_dff_A_L3hODdFd9_2),.din(w_dff_A_VvwERKv35_2),.clk(gclk));
	jdff dff_A_AgMBfGcu6_2(.dout(w_G177gat_0[2]),.din(w_dff_A_AgMBfGcu6_2),.clk(gclk));
	jdff dff_A_98Ja3Kgg6_2(.dout(w_dff_A_AgMBfGcu6_2),.din(w_dff_A_98Ja3Kgg6_2),.clk(gclk));
	jdff dff_A_3wT5SbGB2_2(.dout(w_dff_A_98Ja3Kgg6_2),.din(w_dff_A_3wT5SbGB2_2),.clk(gclk));
	jdff dff_A_Hpxb2jRc1_2(.dout(w_dff_A_3wT5SbGB2_2),.din(w_dff_A_Hpxb2jRc1_2),.clk(gclk));
	jdff dff_A_RUWEpb3u7_1(.dout(w_n405_0[1]),.din(w_dff_A_RUWEpb3u7_1),.clk(gclk));
	jdff dff_A_NlhHi1S28_1(.dout(w_dff_A_RUWEpb3u7_1),.din(w_dff_A_NlhHi1S28_1),.clk(gclk));
	jdff dff_A_J9JUekAm4_1(.dout(w_dff_A_NlhHi1S28_1),.din(w_dff_A_J9JUekAm4_1),.clk(gclk));
	jdff dff_A_SdNXbEZS2_1(.dout(w_dff_A_J9JUekAm4_1),.din(w_dff_A_SdNXbEZS2_1),.clk(gclk));
	jdff dff_A_92ZoAiBn5_1(.dout(w_dff_A_SdNXbEZS2_1),.din(w_dff_A_92ZoAiBn5_1),.clk(gclk));
	jdff dff_A_L1hqvV9p8_1(.dout(w_dff_A_92ZoAiBn5_1),.din(w_dff_A_L1hqvV9p8_1),.clk(gclk));
	jdff dff_A_IfxB44gw2_1(.dout(w_dff_A_L1hqvV9p8_1),.din(w_dff_A_IfxB44gw2_1),.clk(gclk));
	jdff dff_A_QL01JIBY2_1(.dout(w_dff_A_IfxB44gw2_1),.din(w_dff_A_QL01JIBY2_1),.clk(gclk));
	jdff dff_A_ndz4jTRC8_1(.dout(w_dff_A_QL01JIBY2_1),.din(w_dff_A_ndz4jTRC8_1),.clk(gclk));
	jdff dff_B_AadmqBjn3_0(.din(n318),.dout(w_dff_B_AadmqBjn3_0),.clk(gclk));
	jdff dff_B_8IsVf4RO3_0(.din(w_dff_B_AadmqBjn3_0),.dout(w_dff_B_8IsVf4RO3_0),.clk(gclk));
	jdff dff_B_rzvQ8ikQ1_0(.din(w_dff_B_8IsVf4RO3_0),.dout(w_dff_B_rzvQ8ikQ1_0),.clk(gclk));
	jdff dff_B_jjjjMfHr1_0(.din(n295),.dout(w_dff_B_jjjjMfHr1_0),.clk(gclk));
	jdff dff_A_jI7X4yov3_0(.dout(w_G17gat_1[0]),.din(w_dff_A_jI7X4yov3_0),.clk(gclk));
	jdff dff_A_vCcubefC6_2(.dout(w_G17gat_1[2]),.din(w_dff_A_vCcubefC6_2),.clk(gclk));
	jdff dff_A_bG7K8tIg9_2(.dout(w_dff_A_vCcubefC6_2),.din(w_dff_A_bG7K8tIg9_2),.clk(gclk));
	jdff dff_A_Om4YmTQj9_2(.dout(w_dff_A_bG7K8tIg9_2),.din(w_dff_A_Om4YmTQj9_2),.clk(gclk));
	jdff dff_A_meywaUyO7_0(.dout(w_G80gat_0[0]),.din(w_dff_A_meywaUyO7_0),.clk(gclk));
	jdff dff_A_VxBXljXt1_2(.dout(w_G80gat_0[2]),.din(w_dff_A_VxBXljXt1_2),.clk(gclk));
	jdff dff_A_7gBdB4nI1_0(.dout(w_G55gat_0[0]),.din(w_dff_A_7gBdB4nI1_0),.clk(gclk));
	jdff dff_A_g22o4OSZ5_0(.dout(w_dff_A_7gBdB4nI1_0),.din(w_dff_A_g22o4OSZ5_0),.clk(gclk));
	jdff dff_A_nCZDJcW77_0(.dout(w_dff_A_g22o4OSZ5_0),.din(w_dff_A_nCZDJcW77_0),.clk(gclk));
	jdff dff_A_Xxz2xkIl5_1(.dout(w_G55gat_0[1]),.din(w_dff_A_Xxz2xkIl5_1),.clk(gclk));
	jdff dff_A_4JNFA8PX0_1(.dout(w_G149gat_0[1]),.din(w_dff_A_4JNFA8PX0_1),.clk(gclk));
	jdff dff_B_ivJ2mVzD1_2(.din(G149gat),.dout(w_dff_B_ivJ2mVzD1_2),.clk(gclk));
	jdff dff_B_Di0xFvKN4_2(.din(w_dff_B_ivJ2mVzD1_2),.dout(w_dff_B_Di0xFvKN4_2),.clk(gclk));
	jdff dff_B_3xDweony9_2(.din(w_dff_B_Di0xFvKN4_2),.dout(w_dff_B_3xDweony9_2),.clk(gclk));
	jdff dff_B_OZVGGOE57_2(.din(w_dff_B_3xDweony9_2),.dout(w_dff_B_OZVGGOE57_2),.clk(gclk));
	jdff dff_B_udpERRFX2_0(.din(n152),.dout(w_dff_B_udpERRFX2_0),.clk(gclk));
	jdff dff_A_Z8XJFfMx8_0(.dout(w_n149_0[0]),.din(w_dff_A_Z8XJFfMx8_0),.clk(gclk));
	jdff dff_A_tixy5xj33_0(.dout(w_dff_A_Z8XJFfMx8_0),.din(w_dff_A_tixy5xj33_0),.clk(gclk));
	jdff dff_B_zETTW3TP2_0(.din(n147),.dout(w_dff_B_zETTW3TP2_0),.clk(gclk));
	jdff dff_A_wQHYWXrg3_1(.dout(w_G51gat_1[1]),.din(w_dff_A_wQHYWXrg3_1),.clk(gclk));
	jdff dff_A_mLhQAz6c5_1(.dout(w_G1gat_0[1]),.din(w_dff_A_mLhQAz6c5_1),.clk(gclk));
	jdff dff_A_2nGZXnCE3_1(.dout(w_dff_A_mLhQAz6c5_1),.din(w_dff_A_2nGZXnCE3_1),.clk(gclk));
	jdff dff_A_DevPPZdC5_1(.dout(w_dff_A_2nGZXnCE3_1),.din(w_dff_A_DevPPZdC5_1),.clk(gclk));
	jdff dff_A_YQB8dx4G5_1(.dout(w_dff_A_DevPPZdC5_1),.din(w_dff_A_YQB8dx4G5_1),.clk(gclk));
	jdff dff_A_Mjm2LAJE6_1(.dout(w_dff_A_YQB8dx4G5_1),.din(w_dff_A_Mjm2LAJE6_1),.clk(gclk));
	jdff dff_A_PGiJWcjm6_1(.dout(w_G42gat_1[1]),.din(w_dff_A_PGiJWcjm6_1),.clk(gclk));
	jdff dff_A_w0p67XqF8_1(.dout(w_G42gat_0[1]),.din(w_dff_A_w0p67XqF8_1),.clk(gclk));
	jdff dff_A_dlIc9bHV9_1(.dout(w_G101gat_0[1]),.din(w_dff_A_dlIc9bHV9_1),.clk(gclk));
	jdff dff_A_xkfjvA3f2_1(.dout(w_dff_A_dlIc9bHV9_1),.din(w_dff_A_xkfjvA3f2_1),.clk(gclk));
	jdff dff_A_HZUBRvl41_1(.dout(w_dff_A_xkfjvA3f2_1),.din(w_dff_A_HZUBRvl41_1),.clk(gclk));
	jdff dff_A_Pa5fHq2F2_1(.dout(w_dff_A_HZUBRvl41_1),.din(w_dff_A_Pa5fHq2F2_1),.clk(gclk));
	jdff dff_A_YRAMphzX3_1(.dout(w_dff_A_Pa5fHq2F2_1),.din(w_dff_A_YRAMphzX3_1),.clk(gclk));
	jdff dff_A_36VyoqI13_1(.dout(w_G171gat_1[1]),.din(w_dff_A_36VyoqI13_1),.clk(gclk));
	jdff dff_A_BZTn2BFP9_1(.dout(w_dff_A_36VyoqI13_1),.din(w_dff_A_BZTn2BFP9_1),.clk(gclk));
	jdff dff_A_MyGsg31O7_1(.dout(w_dff_A_BZTn2BFP9_1),.din(w_dff_A_MyGsg31O7_1),.clk(gclk));
	jdff dff_A_8l8ryIwm9_1(.dout(w_dff_A_MyGsg31O7_1),.din(w_dff_A_8l8ryIwm9_1),.clk(gclk));
	jdff dff_A_LYfBYSkL1_1(.dout(w_dff_A_8l8ryIwm9_1),.din(w_dff_A_LYfBYSkL1_1),.clk(gclk));
	jdff dff_A_x6DKqCwF4_1(.dout(w_dff_A_LYfBYSkL1_1),.din(w_dff_A_x6DKqCwF4_1),.clk(gclk));
	jdff dff_A_PSEKKTS35_1(.dout(w_dff_A_x6DKqCwF4_1),.din(w_dff_A_PSEKKTS35_1),.clk(gclk));
	jdff dff_A_vxilYzBx3_2(.dout(w_G171gat_1[2]),.din(w_dff_A_vxilYzBx3_2),.clk(gclk));
	jdff dff_A_374xxYkZ3_2(.dout(w_dff_A_vxilYzBx3_2),.din(w_dff_A_374xxYkZ3_2),.clk(gclk));
	jdff dff_A_rGL5bg8K7_2(.dout(w_dff_A_374xxYkZ3_2),.din(w_dff_A_rGL5bg8K7_2),.clk(gclk));
	jdff dff_A_mUtRlnah9_2(.dout(w_dff_A_rGL5bg8K7_2),.din(w_dff_A_mUtRlnah9_2),.clk(gclk));
	jdff dff_A_LvBbnYVl7_2(.dout(w_dff_A_mUtRlnah9_2),.din(w_dff_A_LvBbnYVl7_2),.clk(gclk));
	jdff dff_A_ksBnd4vT7_2(.dout(w_dff_A_LvBbnYVl7_2),.din(w_dff_A_ksBnd4vT7_2),.clk(gclk));
	jdff dff_A_GlMLFNvK1_2(.dout(w_dff_A_ksBnd4vT7_2),.din(w_dff_A_GlMLFNvK1_2),.clk(gclk));
	jdff dff_A_yKX2EfqP3_2(.dout(w_G171gat_0[2]),.din(w_dff_A_yKX2EfqP3_2),.clk(gclk));
	jdff dff_A_6w2Q1Ity1_2(.dout(w_dff_A_yKX2EfqP3_2),.din(w_dff_A_6w2Q1Ity1_2),.clk(gclk));
	jdff dff_A_ShPDGQPY9_2(.dout(w_dff_A_6w2Q1Ity1_2),.din(w_dff_A_ShPDGQPY9_2),.clk(gclk));
	jdff dff_A_rs2z8Iys3_2(.dout(w_dff_A_ShPDGQPY9_2),.din(w_dff_A_rs2z8Iys3_2),.clk(gclk));
	jdff dff_A_Xntldy6t4_2(.dout(w_dff_A_KbI1O0Li6_0),.din(w_dff_A_Xntldy6t4_2),.clk(gclk));
	jdff dff_A_KbI1O0Li6_0(.dout(w_dff_A_HwD9Gvsd8_0),.din(w_dff_A_KbI1O0Li6_0),.clk(gclk));
	jdff dff_A_HwD9Gvsd8_0(.dout(w_dff_A_6RLNHJ3f8_0),.din(w_dff_A_HwD9Gvsd8_0),.clk(gclk));
	jdff dff_A_6RLNHJ3f8_0(.dout(w_dff_A_wzzlXE2A3_0),.din(w_dff_A_6RLNHJ3f8_0),.clk(gclk));
	jdff dff_A_wzzlXE2A3_0(.dout(w_dff_A_OjMacc4E8_0),.din(w_dff_A_wzzlXE2A3_0),.clk(gclk));
	jdff dff_A_OjMacc4E8_0(.dout(w_dff_A_iezIhc946_0),.din(w_dff_A_OjMacc4E8_0),.clk(gclk));
	jdff dff_A_iezIhc946_0(.dout(w_dff_A_fRI2OmYX3_0),.din(w_dff_A_iezIhc946_0),.clk(gclk));
	jdff dff_A_fRI2OmYX3_0(.dout(w_dff_A_MbDeBTxb1_0),.din(w_dff_A_fRI2OmYX3_0),.clk(gclk));
	jdff dff_A_MbDeBTxb1_0(.dout(w_dff_A_dBKiL6a15_0),.din(w_dff_A_MbDeBTxb1_0),.clk(gclk));
	jdff dff_A_dBKiL6a15_0(.dout(w_dff_A_L5orFgfL4_0),.din(w_dff_A_dBKiL6a15_0),.clk(gclk));
	jdff dff_A_L5orFgfL4_0(.dout(w_dff_A_joDeA7Tv2_0),.din(w_dff_A_L5orFgfL4_0),.clk(gclk));
	jdff dff_A_joDeA7Tv2_0(.dout(w_dff_A_VPyLGf2T4_0),.din(w_dff_A_joDeA7Tv2_0),.clk(gclk));
	jdff dff_A_VPyLGf2T4_0(.dout(w_dff_A_dNkfhZNP1_0),.din(w_dff_A_VPyLGf2T4_0),.clk(gclk));
	jdff dff_A_dNkfhZNP1_0(.dout(w_dff_A_mwe0rlSt2_0),.din(w_dff_A_dNkfhZNP1_0),.clk(gclk));
	jdff dff_A_mwe0rlSt2_0(.dout(w_dff_A_kykKmry83_0),.din(w_dff_A_mwe0rlSt2_0),.clk(gclk));
	jdff dff_A_kykKmry83_0(.dout(w_dff_A_fx5Guiuz6_0),.din(w_dff_A_kykKmry83_0),.clk(gclk));
	jdff dff_A_fx5Guiuz6_0(.dout(w_dff_A_oDP3HgJm7_0),.din(w_dff_A_fx5Guiuz6_0),.clk(gclk));
	jdff dff_A_oDP3HgJm7_0(.dout(w_dff_A_MuDXKnsO6_0),.din(w_dff_A_oDP3HgJm7_0),.clk(gclk));
	jdff dff_A_MuDXKnsO6_0(.dout(G388gat),.din(w_dff_A_MuDXKnsO6_0),.clk(gclk));
	jdff dff_A_8q4hYZEa0_2(.dout(w_dff_A_xPTbtNGZ8_0),.din(w_dff_A_8q4hYZEa0_2),.clk(gclk));
	jdff dff_A_xPTbtNGZ8_0(.dout(w_dff_A_wZm4wPkt0_0),.din(w_dff_A_xPTbtNGZ8_0),.clk(gclk));
	jdff dff_A_wZm4wPkt0_0(.dout(w_dff_A_4UIBkS5G1_0),.din(w_dff_A_wZm4wPkt0_0),.clk(gclk));
	jdff dff_A_4UIBkS5G1_0(.dout(w_dff_A_l2vojIM87_0),.din(w_dff_A_4UIBkS5G1_0),.clk(gclk));
	jdff dff_A_l2vojIM87_0(.dout(w_dff_A_jV5KMfvS1_0),.din(w_dff_A_l2vojIM87_0),.clk(gclk));
	jdff dff_A_jV5KMfvS1_0(.dout(w_dff_A_T3vNj6o98_0),.din(w_dff_A_jV5KMfvS1_0),.clk(gclk));
	jdff dff_A_T3vNj6o98_0(.dout(w_dff_A_OCkaEYu48_0),.din(w_dff_A_T3vNj6o98_0),.clk(gclk));
	jdff dff_A_OCkaEYu48_0(.dout(w_dff_A_zWRMz6nS0_0),.din(w_dff_A_OCkaEYu48_0),.clk(gclk));
	jdff dff_A_zWRMz6nS0_0(.dout(w_dff_A_8zyTGUr33_0),.din(w_dff_A_zWRMz6nS0_0),.clk(gclk));
	jdff dff_A_8zyTGUr33_0(.dout(w_dff_A_im91KOK28_0),.din(w_dff_A_8zyTGUr33_0),.clk(gclk));
	jdff dff_A_im91KOK28_0(.dout(w_dff_A_B2nULJo43_0),.din(w_dff_A_im91KOK28_0),.clk(gclk));
	jdff dff_A_B2nULJo43_0(.dout(w_dff_A_BVUtzsI27_0),.din(w_dff_A_B2nULJo43_0),.clk(gclk));
	jdff dff_A_BVUtzsI27_0(.dout(w_dff_A_RCIQiXpR9_0),.din(w_dff_A_BVUtzsI27_0),.clk(gclk));
	jdff dff_A_RCIQiXpR9_0(.dout(w_dff_A_OfzcEk0X5_0),.din(w_dff_A_RCIQiXpR9_0),.clk(gclk));
	jdff dff_A_OfzcEk0X5_0(.dout(w_dff_A_ghzDh9FC4_0),.din(w_dff_A_OfzcEk0X5_0),.clk(gclk));
	jdff dff_A_ghzDh9FC4_0(.dout(w_dff_A_5evEE28F3_0),.din(w_dff_A_ghzDh9FC4_0),.clk(gclk));
	jdff dff_A_5evEE28F3_0(.dout(w_dff_A_IE8ejD1K8_0),.din(w_dff_A_5evEE28F3_0),.clk(gclk));
	jdff dff_A_IE8ejD1K8_0(.dout(w_dff_A_oq4UU4ah3_0),.din(w_dff_A_IE8ejD1K8_0),.clk(gclk));
	jdff dff_A_oq4UU4ah3_0(.dout(G389gat),.din(w_dff_A_oq4UU4ah3_0),.clk(gclk));
	jdff dff_A_LZkuzL3R5_2(.dout(w_dff_A_sTC6SooE5_0),.din(w_dff_A_LZkuzL3R5_2),.clk(gclk));
	jdff dff_A_sTC6SooE5_0(.dout(w_dff_A_eo7wdQuK5_0),.din(w_dff_A_sTC6SooE5_0),.clk(gclk));
	jdff dff_A_eo7wdQuK5_0(.dout(w_dff_A_pJscz6Kw9_0),.din(w_dff_A_eo7wdQuK5_0),.clk(gclk));
	jdff dff_A_pJscz6Kw9_0(.dout(w_dff_A_XrcXhGWw7_0),.din(w_dff_A_pJscz6Kw9_0),.clk(gclk));
	jdff dff_A_XrcXhGWw7_0(.dout(w_dff_A_JpPtK6Xf6_0),.din(w_dff_A_XrcXhGWw7_0),.clk(gclk));
	jdff dff_A_JpPtK6Xf6_0(.dout(w_dff_A_bCngngao2_0),.din(w_dff_A_JpPtK6Xf6_0),.clk(gclk));
	jdff dff_A_bCngngao2_0(.dout(w_dff_A_z7vWbgRv5_0),.din(w_dff_A_bCngngao2_0),.clk(gclk));
	jdff dff_A_z7vWbgRv5_0(.dout(w_dff_A_zwT3vDpk8_0),.din(w_dff_A_z7vWbgRv5_0),.clk(gclk));
	jdff dff_A_zwT3vDpk8_0(.dout(w_dff_A_RptEAGvp9_0),.din(w_dff_A_zwT3vDpk8_0),.clk(gclk));
	jdff dff_A_RptEAGvp9_0(.dout(w_dff_A_Upvtfp5Y1_0),.din(w_dff_A_RptEAGvp9_0),.clk(gclk));
	jdff dff_A_Upvtfp5Y1_0(.dout(w_dff_A_ODUjvdJN6_0),.din(w_dff_A_Upvtfp5Y1_0),.clk(gclk));
	jdff dff_A_ODUjvdJN6_0(.dout(w_dff_A_CoaYQUCE6_0),.din(w_dff_A_ODUjvdJN6_0),.clk(gclk));
	jdff dff_A_CoaYQUCE6_0(.dout(w_dff_A_sXex1YRa4_0),.din(w_dff_A_CoaYQUCE6_0),.clk(gclk));
	jdff dff_A_sXex1YRa4_0(.dout(w_dff_A_JLiOVXCq5_0),.din(w_dff_A_sXex1YRa4_0),.clk(gclk));
	jdff dff_A_JLiOVXCq5_0(.dout(w_dff_A_RJFpea0H9_0),.din(w_dff_A_JLiOVXCq5_0),.clk(gclk));
	jdff dff_A_RJFpea0H9_0(.dout(w_dff_A_oXGKYB0N7_0),.din(w_dff_A_RJFpea0H9_0),.clk(gclk));
	jdff dff_A_oXGKYB0N7_0(.dout(w_dff_A_izYa1v5x2_0),.din(w_dff_A_oXGKYB0N7_0),.clk(gclk));
	jdff dff_A_izYa1v5x2_0(.dout(w_dff_A_AaRMdoEz8_0),.din(w_dff_A_izYa1v5x2_0),.clk(gclk));
	jdff dff_A_AaRMdoEz8_0(.dout(G390gat),.din(w_dff_A_AaRMdoEz8_0),.clk(gclk));
	jdff dff_A_lNIUOv8Z3_2(.dout(w_dff_A_9QuSUTrw6_0),.din(w_dff_A_lNIUOv8Z3_2),.clk(gclk));
	jdff dff_A_9QuSUTrw6_0(.dout(w_dff_A_s1sbIzuM7_0),.din(w_dff_A_9QuSUTrw6_0),.clk(gclk));
	jdff dff_A_s1sbIzuM7_0(.dout(w_dff_A_n8nz6vkt2_0),.din(w_dff_A_s1sbIzuM7_0),.clk(gclk));
	jdff dff_A_n8nz6vkt2_0(.dout(w_dff_A_JGm44D9l8_0),.din(w_dff_A_n8nz6vkt2_0),.clk(gclk));
	jdff dff_A_JGm44D9l8_0(.dout(w_dff_A_QFMfETWL7_0),.din(w_dff_A_JGm44D9l8_0),.clk(gclk));
	jdff dff_A_QFMfETWL7_0(.dout(w_dff_A_9BQeGxpk9_0),.din(w_dff_A_QFMfETWL7_0),.clk(gclk));
	jdff dff_A_9BQeGxpk9_0(.dout(w_dff_A_ZjoVzQfi6_0),.din(w_dff_A_9BQeGxpk9_0),.clk(gclk));
	jdff dff_A_ZjoVzQfi6_0(.dout(w_dff_A_EfirJdH51_0),.din(w_dff_A_ZjoVzQfi6_0),.clk(gclk));
	jdff dff_A_EfirJdH51_0(.dout(w_dff_A_GTAl8Tye4_0),.din(w_dff_A_EfirJdH51_0),.clk(gclk));
	jdff dff_A_GTAl8Tye4_0(.dout(w_dff_A_JFhCzmdc7_0),.din(w_dff_A_GTAl8Tye4_0),.clk(gclk));
	jdff dff_A_JFhCzmdc7_0(.dout(w_dff_A_q64hj3Sz5_0),.din(w_dff_A_JFhCzmdc7_0),.clk(gclk));
	jdff dff_A_q64hj3Sz5_0(.dout(w_dff_A_CuQ7muhK0_0),.din(w_dff_A_q64hj3Sz5_0),.clk(gclk));
	jdff dff_A_CuQ7muhK0_0(.dout(w_dff_A_PFSyVOOQ3_0),.din(w_dff_A_CuQ7muhK0_0),.clk(gclk));
	jdff dff_A_PFSyVOOQ3_0(.dout(w_dff_A_FA5wy5YP7_0),.din(w_dff_A_PFSyVOOQ3_0),.clk(gclk));
	jdff dff_A_FA5wy5YP7_0(.dout(w_dff_A_yd0fbcGO0_0),.din(w_dff_A_FA5wy5YP7_0),.clk(gclk));
	jdff dff_A_yd0fbcGO0_0(.dout(w_dff_A_jqhYfzFw6_0),.din(w_dff_A_yd0fbcGO0_0),.clk(gclk));
	jdff dff_A_jqhYfzFw6_0(.dout(w_dff_A_bCZxmP5L5_0),.din(w_dff_A_jqhYfzFw6_0),.clk(gclk));
	jdff dff_A_bCZxmP5L5_0(.dout(w_dff_A_7Ym21FOd6_0),.din(w_dff_A_bCZxmP5L5_0),.clk(gclk));
	jdff dff_A_7Ym21FOd6_0(.dout(w_dff_A_IyfHgiX69_0),.din(w_dff_A_7Ym21FOd6_0),.clk(gclk));
	jdff dff_A_IyfHgiX69_0(.dout(G391gat),.din(w_dff_A_IyfHgiX69_0),.clk(gclk));
	jdff dff_A_LcBxnPK44_2(.dout(w_dff_A_EVmSVshh4_0),.din(w_dff_A_LcBxnPK44_2),.clk(gclk));
	jdff dff_A_EVmSVshh4_0(.dout(w_dff_A_TAvlpuRY5_0),.din(w_dff_A_EVmSVshh4_0),.clk(gclk));
	jdff dff_A_TAvlpuRY5_0(.dout(w_dff_A_Ng5jKy9L0_0),.din(w_dff_A_TAvlpuRY5_0),.clk(gclk));
	jdff dff_A_Ng5jKy9L0_0(.dout(w_dff_A_oSDL6rJH2_0),.din(w_dff_A_Ng5jKy9L0_0),.clk(gclk));
	jdff dff_A_oSDL6rJH2_0(.dout(w_dff_A_0CZpg5L10_0),.din(w_dff_A_oSDL6rJH2_0),.clk(gclk));
	jdff dff_A_0CZpg5L10_0(.dout(w_dff_A_YTyortLz5_0),.din(w_dff_A_0CZpg5L10_0),.clk(gclk));
	jdff dff_A_YTyortLz5_0(.dout(w_dff_A_eZia1YNg5_0),.din(w_dff_A_YTyortLz5_0),.clk(gclk));
	jdff dff_A_eZia1YNg5_0(.dout(w_dff_A_jhD9kbtS6_0),.din(w_dff_A_eZia1YNg5_0),.clk(gclk));
	jdff dff_A_jhD9kbtS6_0(.dout(w_dff_A_mgNjCEzV9_0),.din(w_dff_A_jhD9kbtS6_0),.clk(gclk));
	jdff dff_A_mgNjCEzV9_0(.dout(w_dff_A_4BTToW5j4_0),.din(w_dff_A_mgNjCEzV9_0),.clk(gclk));
	jdff dff_A_4BTToW5j4_0(.dout(w_dff_A_UaT1PotL7_0),.din(w_dff_A_4BTToW5j4_0),.clk(gclk));
	jdff dff_A_UaT1PotL7_0(.dout(w_dff_A_6WAL0zSB2_0),.din(w_dff_A_UaT1PotL7_0),.clk(gclk));
	jdff dff_A_6WAL0zSB2_0(.dout(w_dff_A_EXVPbxuf8_0),.din(w_dff_A_6WAL0zSB2_0),.clk(gclk));
	jdff dff_A_EXVPbxuf8_0(.dout(w_dff_A_65LjyrMF7_0),.din(w_dff_A_EXVPbxuf8_0),.clk(gclk));
	jdff dff_A_65LjyrMF7_0(.dout(w_dff_A_vNuX6L9g4_0),.din(w_dff_A_65LjyrMF7_0),.clk(gclk));
	jdff dff_A_vNuX6L9g4_0(.dout(w_dff_A_oblXIxF02_0),.din(w_dff_A_vNuX6L9g4_0),.clk(gclk));
	jdff dff_A_oblXIxF02_0(.dout(w_dff_A_FwO04bgL3_0),.din(w_dff_A_oblXIxF02_0),.clk(gclk));
	jdff dff_A_FwO04bgL3_0(.dout(w_dff_A_JrWkhz5v5_0),.din(w_dff_A_FwO04bgL3_0),.clk(gclk));
	jdff dff_A_JrWkhz5v5_0(.dout(G418gat),.din(w_dff_A_JrWkhz5v5_0),.clk(gclk));
	jdff dff_A_om5yfFJZ9_2(.dout(w_dff_A_wFkHDRkN0_0),.din(w_dff_A_om5yfFJZ9_2),.clk(gclk));
	jdff dff_A_wFkHDRkN0_0(.dout(w_dff_A_7DIPzXgA2_0),.din(w_dff_A_wFkHDRkN0_0),.clk(gclk));
	jdff dff_A_7DIPzXgA2_0(.dout(w_dff_A_kSQEXk5g5_0),.din(w_dff_A_7DIPzXgA2_0),.clk(gclk));
	jdff dff_A_kSQEXk5g5_0(.dout(w_dff_A_ca2QhFIc0_0),.din(w_dff_A_kSQEXk5g5_0),.clk(gclk));
	jdff dff_A_ca2QhFIc0_0(.dout(w_dff_A_6C7OKgw35_0),.din(w_dff_A_ca2QhFIc0_0),.clk(gclk));
	jdff dff_A_6C7OKgw35_0(.dout(w_dff_A_Fp8rfe5R6_0),.din(w_dff_A_6C7OKgw35_0),.clk(gclk));
	jdff dff_A_Fp8rfe5R6_0(.dout(w_dff_A_8hsaQADq1_0),.din(w_dff_A_Fp8rfe5R6_0),.clk(gclk));
	jdff dff_A_8hsaQADq1_0(.dout(w_dff_A_zjvc2mYh4_0),.din(w_dff_A_8hsaQADq1_0),.clk(gclk));
	jdff dff_A_zjvc2mYh4_0(.dout(w_dff_A_pgd1iREk3_0),.din(w_dff_A_zjvc2mYh4_0),.clk(gclk));
	jdff dff_A_pgd1iREk3_0(.dout(w_dff_A_lbwzw8Zt0_0),.din(w_dff_A_pgd1iREk3_0),.clk(gclk));
	jdff dff_A_lbwzw8Zt0_0(.dout(w_dff_A_Mx92Rox19_0),.din(w_dff_A_lbwzw8Zt0_0),.clk(gclk));
	jdff dff_A_Mx92Rox19_0(.dout(w_dff_A_2jcBRt5V6_0),.din(w_dff_A_Mx92Rox19_0),.clk(gclk));
	jdff dff_A_2jcBRt5V6_0(.dout(w_dff_A_u1Dr9DA03_0),.din(w_dff_A_2jcBRt5V6_0),.clk(gclk));
	jdff dff_A_u1Dr9DA03_0(.dout(w_dff_A_un9KlenZ7_0),.din(w_dff_A_u1Dr9DA03_0),.clk(gclk));
	jdff dff_A_un9KlenZ7_0(.dout(w_dff_A_JZbjTR1k7_0),.din(w_dff_A_un9KlenZ7_0),.clk(gclk));
	jdff dff_A_JZbjTR1k7_0(.dout(w_dff_A_fXPC6ktv8_0),.din(w_dff_A_JZbjTR1k7_0),.clk(gclk));
	jdff dff_A_fXPC6ktv8_0(.dout(G419gat),.din(w_dff_A_fXPC6ktv8_0),.clk(gclk));
	jdff dff_A_HeZ3jRFr2_2(.dout(w_dff_A_GWeUZ3Ph0_0),.din(w_dff_A_HeZ3jRFr2_2),.clk(gclk));
	jdff dff_A_GWeUZ3Ph0_0(.dout(w_dff_A_BxQg5xdj5_0),.din(w_dff_A_GWeUZ3Ph0_0),.clk(gclk));
	jdff dff_A_BxQg5xdj5_0(.dout(w_dff_A_Lft3Zjlj3_0),.din(w_dff_A_BxQg5xdj5_0),.clk(gclk));
	jdff dff_A_Lft3Zjlj3_0(.dout(w_dff_A_hRVzl9vg0_0),.din(w_dff_A_Lft3Zjlj3_0),.clk(gclk));
	jdff dff_A_hRVzl9vg0_0(.dout(w_dff_A_vIGz3kAM3_0),.din(w_dff_A_hRVzl9vg0_0),.clk(gclk));
	jdff dff_A_vIGz3kAM3_0(.dout(w_dff_A_jKLSxyQb1_0),.din(w_dff_A_vIGz3kAM3_0),.clk(gclk));
	jdff dff_A_jKLSxyQb1_0(.dout(w_dff_A_eS3lpG7T6_0),.din(w_dff_A_jKLSxyQb1_0),.clk(gclk));
	jdff dff_A_eS3lpG7T6_0(.dout(w_dff_A_NA1xOXbL2_0),.din(w_dff_A_eS3lpG7T6_0),.clk(gclk));
	jdff dff_A_NA1xOXbL2_0(.dout(w_dff_A_9uZsmQkm2_0),.din(w_dff_A_NA1xOXbL2_0),.clk(gclk));
	jdff dff_A_9uZsmQkm2_0(.dout(w_dff_A_sb4fYoiv4_0),.din(w_dff_A_9uZsmQkm2_0),.clk(gclk));
	jdff dff_A_sb4fYoiv4_0(.dout(w_dff_A_fOJCMub76_0),.din(w_dff_A_sb4fYoiv4_0),.clk(gclk));
	jdff dff_A_fOJCMub76_0(.dout(w_dff_A_Y4gymV6T2_0),.din(w_dff_A_fOJCMub76_0),.clk(gclk));
	jdff dff_A_Y4gymV6T2_0(.dout(w_dff_A_IALfDD7n7_0),.din(w_dff_A_Y4gymV6T2_0),.clk(gclk));
	jdff dff_A_IALfDD7n7_0(.dout(w_dff_A_VUkdmvpH5_0),.din(w_dff_A_IALfDD7n7_0),.clk(gclk));
	jdff dff_A_VUkdmvpH5_0(.dout(w_dff_A_BN6dc5Vf5_0),.din(w_dff_A_VUkdmvpH5_0),.clk(gclk));
	jdff dff_A_BN6dc5Vf5_0(.dout(w_dff_A_KC6954ZE3_0),.din(w_dff_A_BN6dc5Vf5_0),.clk(gclk));
	jdff dff_A_KC6954ZE3_0(.dout(w_dff_A_4BtlkvJK0_0),.din(w_dff_A_KC6954ZE3_0),.clk(gclk));
	jdff dff_A_4BtlkvJK0_0(.dout(G420gat),.din(w_dff_A_4BtlkvJK0_0),.clk(gclk));
	jdff dff_A_fN7Sqhtz9_2(.dout(w_dff_A_X4vtqVKS5_0),.din(w_dff_A_fN7Sqhtz9_2),.clk(gclk));
	jdff dff_A_X4vtqVKS5_0(.dout(w_dff_A_0V4AT2zD8_0),.din(w_dff_A_X4vtqVKS5_0),.clk(gclk));
	jdff dff_A_0V4AT2zD8_0(.dout(w_dff_A_AsYtUIVv9_0),.din(w_dff_A_0V4AT2zD8_0),.clk(gclk));
	jdff dff_A_AsYtUIVv9_0(.dout(w_dff_A_PtWdQm3q7_0),.din(w_dff_A_AsYtUIVv9_0),.clk(gclk));
	jdff dff_A_PtWdQm3q7_0(.dout(w_dff_A_2Ngi02M84_0),.din(w_dff_A_PtWdQm3q7_0),.clk(gclk));
	jdff dff_A_2Ngi02M84_0(.dout(w_dff_A_mkmWWU8L8_0),.din(w_dff_A_2Ngi02M84_0),.clk(gclk));
	jdff dff_A_mkmWWU8L8_0(.dout(w_dff_A_0GJzQxL10_0),.din(w_dff_A_mkmWWU8L8_0),.clk(gclk));
	jdff dff_A_0GJzQxL10_0(.dout(w_dff_A_2xGe2Emd1_0),.din(w_dff_A_0GJzQxL10_0),.clk(gclk));
	jdff dff_A_2xGe2Emd1_0(.dout(w_dff_A_EuNUbaaj2_0),.din(w_dff_A_2xGe2Emd1_0),.clk(gclk));
	jdff dff_A_EuNUbaaj2_0(.dout(w_dff_A_taDBZjTd4_0),.din(w_dff_A_EuNUbaaj2_0),.clk(gclk));
	jdff dff_A_taDBZjTd4_0(.dout(w_dff_A_LFjYlNYn7_0),.din(w_dff_A_taDBZjTd4_0),.clk(gclk));
	jdff dff_A_LFjYlNYn7_0(.dout(w_dff_A_R67gdMvw8_0),.din(w_dff_A_LFjYlNYn7_0),.clk(gclk));
	jdff dff_A_R67gdMvw8_0(.dout(w_dff_A_m6nrYg2h5_0),.din(w_dff_A_R67gdMvw8_0),.clk(gclk));
	jdff dff_A_m6nrYg2h5_0(.dout(w_dff_A_SaxFcQyt3_0),.din(w_dff_A_m6nrYg2h5_0),.clk(gclk));
	jdff dff_A_SaxFcQyt3_0(.dout(w_dff_A_9gk8OFil8_0),.din(w_dff_A_SaxFcQyt3_0),.clk(gclk));
	jdff dff_A_9gk8OFil8_0(.dout(w_dff_A_tgQpqa4J2_0),.din(w_dff_A_9gk8OFil8_0),.clk(gclk));
	jdff dff_A_tgQpqa4J2_0(.dout(w_dff_A_y9CJdFj68_0),.din(w_dff_A_tgQpqa4J2_0),.clk(gclk));
	jdff dff_A_y9CJdFj68_0(.dout(G421gat),.din(w_dff_A_y9CJdFj68_0),.clk(gclk));
	jdff dff_A_HLc1PW0D5_2(.dout(w_dff_A_xkvkgoy20_0),.din(w_dff_A_HLc1PW0D5_2),.clk(gclk));
	jdff dff_A_xkvkgoy20_0(.dout(w_dff_A_NVy69MsY1_0),.din(w_dff_A_xkvkgoy20_0),.clk(gclk));
	jdff dff_A_NVy69MsY1_0(.dout(w_dff_A_BmKjPyn96_0),.din(w_dff_A_NVy69MsY1_0),.clk(gclk));
	jdff dff_A_BmKjPyn96_0(.dout(w_dff_A_CkY47CdA6_0),.din(w_dff_A_BmKjPyn96_0),.clk(gclk));
	jdff dff_A_CkY47CdA6_0(.dout(w_dff_A_eEf2ED1m7_0),.din(w_dff_A_CkY47CdA6_0),.clk(gclk));
	jdff dff_A_eEf2ED1m7_0(.dout(w_dff_A_hmTwZ0ud4_0),.din(w_dff_A_eEf2ED1m7_0),.clk(gclk));
	jdff dff_A_hmTwZ0ud4_0(.dout(w_dff_A_6e4D3hyf4_0),.din(w_dff_A_hmTwZ0ud4_0),.clk(gclk));
	jdff dff_A_6e4D3hyf4_0(.dout(w_dff_A_ESJRskFL9_0),.din(w_dff_A_6e4D3hyf4_0),.clk(gclk));
	jdff dff_A_ESJRskFL9_0(.dout(w_dff_A_tS4za1nY9_0),.din(w_dff_A_ESJRskFL9_0),.clk(gclk));
	jdff dff_A_tS4za1nY9_0(.dout(w_dff_A_1bBMaS7h7_0),.din(w_dff_A_tS4za1nY9_0),.clk(gclk));
	jdff dff_A_1bBMaS7h7_0(.dout(w_dff_A_ywJAphae0_0),.din(w_dff_A_1bBMaS7h7_0),.clk(gclk));
	jdff dff_A_ywJAphae0_0(.dout(w_dff_A_ySyXdsmH1_0),.din(w_dff_A_ywJAphae0_0),.clk(gclk));
	jdff dff_A_ySyXdsmH1_0(.dout(w_dff_A_FNxxjxIv1_0),.din(w_dff_A_ySyXdsmH1_0),.clk(gclk));
	jdff dff_A_FNxxjxIv1_0(.dout(w_dff_A_IxHs60Sp0_0),.din(w_dff_A_FNxxjxIv1_0),.clk(gclk));
	jdff dff_A_IxHs60Sp0_0(.dout(w_dff_A_tcaDIE257_0),.din(w_dff_A_IxHs60Sp0_0),.clk(gclk));
	jdff dff_A_tcaDIE257_0(.dout(w_dff_A_ySiKg4xZ1_0),.din(w_dff_A_tcaDIE257_0),.clk(gclk));
	jdff dff_A_ySiKg4xZ1_0(.dout(w_dff_A_ZpIgaS6M9_0),.din(w_dff_A_ySiKg4xZ1_0),.clk(gclk));
	jdff dff_A_ZpIgaS6M9_0(.dout(G422gat),.din(w_dff_A_ZpIgaS6M9_0),.clk(gclk));
	jdff dff_A_iMewsF9N8_2(.dout(w_dff_A_vaSG4d708_0),.din(w_dff_A_iMewsF9N8_2),.clk(gclk));
	jdff dff_A_vaSG4d708_0(.dout(w_dff_A_x4SuF3BL8_0),.din(w_dff_A_vaSG4d708_0),.clk(gclk));
	jdff dff_A_x4SuF3BL8_0(.dout(w_dff_A_szAv4nas4_0),.din(w_dff_A_x4SuF3BL8_0),.clk(gclk));
	jdff dff_A_szAv4nas4_0(.dout(w_dff_A_qtlPwTV65_0),.din(w_dff_A_szAv4nas4_0),.clk(gclk));
	jdff dff_A_qtlPwTV65_0(.dout(w_dff_A_NiMiWQJ36_0),.din(w_dff_A_qtlPwTV65_0),.clk(gclk));
	jdff dff_A_NiMiWQJ36_0(.dout(w_dff_A_sjNa6rfS2_0),.din(w_dff_A_NiMiWQJ36_0),.clk(gclk));
	jdff dff_A_sjNa6rfS2_0(.dout(w_dff_A_lmO4PdFJ0_0),.din(w_dff_A_sjNa6rfS2_0),.clk(gclk));
	jdff dff_A_lmO4PdFJ0_0(.dout(w_dff_A_HaEKUkna8_0),.din(w_dff_A_lmO4PdFJ0_0),.clk(gclk));
	jdff dff_A_HaEKUkna8_0(.dout(w_dff_A_odmub6DX6_0),.din(w_dff_A_HaEKUkna8_0),.clk(gclk));
	jdff dff_A_odmub6DX6_0(.dout(w_dff_A_jHBi5Bfo5_0),.din(w_dff_A_odmub6DX6_0),.clk(gclk));
	jdff dff_A_jHBi5Bfo5_0(.dout(w_dff_A_toBZB2Nw6_0),.din(w_dff_A_jHBi5Bfo5_0),.clk(gclk));
	jdff dff_A_toBZB2Nw6_0(.dout(w_dff_A_QIzUUu018_0),.din(w_dff_A_toBZB2Nw6_0),.clk(gclk));
	jdff dff_A_QIzUUu018_0(.dout(w_dff_A_H6to52x65_0),.din(w_dff_A_QIzUUu018_0),.clk(gclk));
	jdff dff_A_H6to52x65_0(.dout(w_dff_A_SoN1Y4fW7_0),.din(w_dff_A_H6to52x65_0),.clk(gclk));
	jdff dff_A_SoN1Y4fW7_0(.dout(w_dff_A_GBXdkGzH7_0),.din(w_dff_A_SoN1Y4fW7_0),.clk(gclk));
	jdff dff_A_GBXdkGzH7_0(.dout(w_dff_A_bNeRAaKI0_0),.din(w_dff_A_GBXdkGzH7_0),.clk(gclk));
	jdff dff_A_bNeRAaKI0_0(.dout(w_dff_A_YEhqLxN09_0),.din(w_dff_A_bNeRAaKI0_0),.clk(gclk));
	jdff dff_A_YEhqLxN09_0(.dout(w_dff_A_SaCeGyxV2_0),.din(w_dff_A_YEhqLxN09_0),.clk(gclk));
	jdff dff_A_SaCeGyxV2_0(.dout(G423gat),.din(w_dff_A_SaCeGyxV2_0),.clk(gclk));
	jdff dff_A_qRuj8HhM0_2(.dout(w_dff_A_71EuurKe6_0),.din(w_dff_A_qRuj8HhM0_2),.clk(gclk));
	jdff dff_A_71EuurKe6_0(.dout(w_dff_A_0RLeOXEr3_0),.din(w_dff_A_71EuurKe6_0),.clk(gclk));
	jdff dff_A_0RLeOXEr3_0(.dout(w_dff_A_JCDd51sk5_0),.din(w_dff_A_0RLeOXEr3_0),.clk(gclk));
	jdff dff_A_JCDd51sk5_0(.dout(w_dff_A_cQ3UmHPN5_0),.din(w_dff_A_JCDd51sk5_0),.clk(gclk));
	jdff dff_A_cQ3UmHPN5_0(.dout(w_dff_A_3s5bnS9l2_0),.din(w_dff_A_cQ3UmHPN5_0),.clk(gclk));
	jdff dff_A_3s5bnS9l2_0(.dout(w_dff_A_e48IVaOt7_0),.din(w_dff_A_3s5bnS9l2_0),.clk(gclk));
	jdff dff_A_e48IVaOt7_0(.dout(w_dff_A_Pv9jvW6z7_0),.din(w_dff_A_e48IVaOt7_0),.clk(gclk));
	jdff dff_A_Pv9jvW6z7_0(.dout(w_dff_A_Cvz3BPRS8_0),.din(w_dff_A_Pv9jvW6z7_0),.clk(gclk));
	jdff dff_A_Cvz3BPRS8_0(.dout(w_dff_A_4NBxotBM5_0),.din(w_dff_A_Cvz3BPRS8_0),.clk(gclk));
	jdff dff_A_4NBxotBM5_0(.dout(w_dff_A_DA1vM29x0_0),.din(w_dff_A_4NBxotBM5_0),.clk(gclk));
	jdff dff_A_DA1vM29x0_0(.dout(w_dff_A_79i2WSZs8_0),.din(w_dff_A_DA1vM29x0_0),.clk(gclk));
	jdff dff_A_79i2WSZs8_0(.dout(w_dff_A_yTO5944o6_0),.din(w_dff_A_79i2WSZs8_0),.clk(gclk));
	jdff dff_A_yTO5944o6_0(.dout(w_dff_A_L8zE4EKL6_0),.din(w_dff_A_yTO5944o6_0),.clk(gclk));
	jdff dff_A_L8zE4EKL6_0(.dout(w_dff_A_aeihurQx3_0),.din(w_dff_A_L8zE4EKL6_0),.clk(gclk));
	jdff dff_A_aeihurQx3_0(.dout(w_dff_A_rUFO2HwF2_0),.din(w_dff_A_aeihurQx3_0),.clk(gclk));
	jdff dff_A_rUFO2HwF2_0(.dout(w_dff_A_Te4VIOed3_0),.din(w_dff_A_rUFO2HwF2_0),.clk(gclk));
	jdff dff_A_Te4VIOed3_0(.dout(G446gat),.din(w_dff_A_Te4VIOed3_0),.clk(gclk));
	jdff dff_A_4xqBO2HF8_1(.dout(w_dff_A_somV81jX7_0),.din(w_dff_A_4xqBO2HF8_1),.clk(gclk));
	jdff dff_A_somV81jX7_0(.dout(w_dff_A_eitVJNG94_0),.din(w_dff_A_somV81jX7_0),.clk(gclk));
	jdff dff_A_eitVJNG94_0(.dout(w_dff_A_I2OjUYlH3_0),.din(w_dff_A_eitVJNG94_0),.clk(gclk));
	jdff dff_A_I2OjUYlH3_0(.dout(w_dff_A_oxdftX4d5_0),.din(w_dff_A_I2OjUYlH3_0),.clk(gclk));
	jdff dff_A_oxdftX4d5_0(.dout(w_dff_A_bd3ws9tz4_0),.din(w_dff_A_oxdftX4d5_0),.clk(gclk));
	jdff dff_A_bd3ws9tz4_0(.dout(w_dff_A_9Ojln7L75_0),.din(w_dff_A_bd3ws9tz4_0),.clk(gclk));
	jdff dff_A_9Ojln7L75_0(.dout(w_dff_A_G878MytB8_0),.din(w_dff_A_9Ojln7L75_0),.clk(gclk));
	jdff dff_A_G878MytB8_0(.dout(w_dff_A_dScHZvv86_0),.din(w_dff_A_G878MytB8_0),.clk(gclk));
	jdff dff_A_dScHZvv86_0(.dout(w_dff_A_MRbRN5f95_0),.din(w_dff_A_dScHZvv86_0),.clk(gclk));
	jdff dff_A_MRbRN5f95_0(.dout(w_dff_A_B5ScHvZj1_0),.din(w_dff_A_MRbRN5f95_0),.clk(gclk));
	jdff dff_A_B5ScHvZj1_0(.dout(w_dff_A_PAKlTkdn2_0),.din(w_dff_A_B5ScHvZj1_0),.clk(gclk));
	jdff dff_A_PAKlTkdn2_0(.dout(w_dff_A_Me6gvWQp7_0),.din(w_dff_A_PAKlTkdn2_0),.clk(gclk));
	jdff dff_A_Me6gvWQp7_0(.dout(w_dff_A_hS4DMq2w7_0),.din(w_dff_A_Me6gvWQp7_0),.clk(gclk));
	jdff dff_A_hS4DMq2w7_0(.dout(w_dff_A_1gFLst8r9_0),.din(w_dff_A_hS4DMq2w7_0),.clk(gclk));
	jdff dff_A_1gFLst8r9_0(.dout(w_dff_A_a8ybMeff9_0),.din(w_dff_A_1gFLst8r9_0),.clk(gclk));
	jdff dff_A_a8ybMeff9_0(.dout(w_dff_A_yuPIEYgL9_0),.din(w_dff_A_a8ybMeff9_0),.clk(gclk));
	jdff dff_A_yuPIEYgL9_0(.dout(w_dff_A_uee924xu4_0),.din(w_dff_A_yuPIEYgL9_0),.clk(gclk));
	jdff dff_A_uee924xu4_0(.dout(w_dff_A_UKevBCaG4_0),.din(w_dff_A_uee924xu4_0),.clk(gclk));
	jdff dff_A_UKevBCaG4_0(.dout(G447gat),.din(w_dff_A_UKevBCaG4_0),.clk(gclk));
	jdff dff_A_dO4Fam3e8_2(.dout(w_dff_A_uEPPxuz07_0),.din(w_dff_A_dO4Fam3e8_2),.clk(gclk));
	jdff dff_A_uEPPxuz07_0(.dout(w_dff_A_rHzmUiJb4_0),.din(w_dff_A_uEPPxuz07_0),.clk(gclk));
	jdff dff_A_rHzmUiJb4_0(.dout(w_dff_A_9R1MTHIf6_0),.din(w_dff_A_rHzmUiJb4_0),.clk(gclk));
	jdff dff_A_9R1MTHIf6_0(.dout(w_dff_A_dUecXQBk2_0),.din(w_dff_A_9R1MTHIf6_0),.clk(gclk));
	jdff dff_A_dUecXQBk2_0(.dout(w_dff_A_05pOeuiE3_0),.din(w_dff_A_dUecXQBk2_0),.clk(gclk));
	jdff dff_A_05pOeuiE3_0(.dout(w_dff_A_5T3pQLEH4_0),.din(w_dff_A_05pOeuiE3_0),.clk(gclk));
	jdff dff_A_5T3pQLEH4_0(.dout(w_dff_A_AD7lS7079_0),.din(w_dff_A_5T3pQLEH4_0),.clk(gclk));
	jdff dff_A_AD7lS7079_0(.dout(w_dff_A_zDJfbgFf2_0),.din(w_dff_A_AD7lS7079_0),.clk(gclk));
	jdff dff_A_zDJfbgFf2_0(.dout(w_dff_A_OD5qzNsb7_0),.din(w_dff_A_zDJfbgFf2_0),.clk(gclk));
	jdff dff_A_OD5qzNsb7_0(.dout(w_dff_A_P8ioZ82P7_0),.din(w_dff_A_OD5qzNsb7_0),.clk(gclk));
	jdff dff_A_P8ioZ82P7_0(.dout(w_dff_A_vGMP4ftZ9_0),.din(w_dff_A_P8ioZ82P7_0),.clk(gclk));
	jdff dff_A_vGMP4ftZ9_0(.dout(w_dff_A_1BoVzjbG2_0),.din(w_dff_A_vGMP4ftZ9_0),.clk(gclk));
	jdff dff_A_1BoVzjbG2_0(.dout(w_dff_A_i0PaspVa8_0),.din(w_dff_A_1BoVzjbG2_0),.clk(gclk));
	jdff dff_A_i0PaspVa8_0(.dout(w_dff_A_KSkfFaDD8_0),.din(w_dff_A_i0PaspVa8_0),.clk(gclk));
	jdff dff_A_KSkfFaDD8_0(.dout(w_dff_A_z1D2e0wE6_0),.din(w_dff_A_KSkfFaDD8_0),.clk(gclk));
	jdff dff_A_z1D2e0wE6_0(.dout(w_dff_A_AABn1yD90_0),.din(w_dff_A_z1D2e0wE6_0),.clk(gclk));
	jdff dff_A_AABn1yD90_0(.dout(w_dff_A_PWvanrdV6_0),.din(w_dff_A_AABn1yD90_0),.clk(gclk));
	jdff dff_A_PWvanrdV6_0(.dout(G448gat),.din(w_dff_A_PWvanrdV6_0),.clk(gclk));
	jdff dff_A_6MABsAz43_2(.dout(w_dff_A_oYESdbrw1_0),.din(w_dff_A_6MABsAz43_2),.clk(gclk));
	jdff dff_A_oYESdbrw1_0(.dout(w_dff_A_JZxxlBLw0_0),.din(w_dff_A_oYESdbrw1_0),.clk(gclk));
	jdff dff_A_JZxxlBLw0_0(.dout(w_dff_A_Ci9vNr2o4_0),.din(w_dff_A_JZxxlBLw0_0),.clk(gclk));
	jdff dff_A_Ci9vNr2o4_0(.dout(w_dff_A_cqtx839A6_0),.din(w_dff_A_Ci9vNr2o4_0),.clk(gclk));
	jdff dff_A_cqtx839A6_0(.dout(w_dff_A_QKyXmqNM5_0),.din(w_dff_A_cqtx839A6_0),.clk(gclk));
	jdff dff_A_QKyXmqNM5_0(.dout(w_dff_A_0SU8pNDo8_0),.din(w_dff_A_QKyXmqNM5_0),.clk(gclk));
	jdff dff_A_0SU8pNDo8_0(.dout(w_dff_A_meCZUS2W1_0),.din(w_dff_A_0SU8pNDo8_0),.clk(gclk));
	jdff dff_A_meCZUS2W1_0(.dout(w_dff_A_xSsipH7N6_0),.din(w_dff_A_meCZUS2W1_0),.clk(gclk));
	jdff dff_A_xSsipH7N6_0(.dout(w_dff_A_1DriepDL8_0),.din(w_dff_A_xSsipH7N6_0),.clk(gclk));
	jdff dff_A_1DriepDL8_0(.dout(w_dff_A_V19H7jzo8_0),.din(w_dff_A_1DriepDL8_0),.clk(gclk));
	jdff dff_A_V19H7jzo8_0(.dout(w_dff_A_67hsqkPb6_0),.din(w_dff_A_V19H7jzo8_0),.clk(gclk));
	jdff dff_A_67hsqkPb6_0(.dout(w_dff_A_SNaqiekO6_0),.din(w_dff_A_67hsqkPb6_0),.clk(gclk));
	jdff dff_A_SNaqiekO6_0(.dout(w_dff_A_bZ2cGZRe5_0),.din(w_dff_A_SNaqiekO6_0),.clk(gclk));
	jdff dff_A_bZ2cGZRe5_0(.dout(w_dff_A_itEyNGxY3_0),.din(w_dff_A_bZ2cGZRe5_0),.clk(gclk));
	jdff dff_A_itEyNGxY3_0(.dout(w_dff_A_qg0kKzdK2_0),.din(w_dff_A_itEyNGxY3_0),.clk(gclk));
	jdff dff_A_qg0kKzdK2_0(.dout(w_dff_A_bUch3oDI5_0),.din(w_dff_A_qg0kKzdK2_0),.clk(gclk));
	jdff dff_A_bUch3oDI5_0(.dout(w_dff_A_CVZsVZfq1_0),.din(w_dff_A_bUch3oDI5_0),.clk(gclk));
	jdff dff_A_CVZsVZfq1_0(.dout(G449gat),.din(w_dff_A_CVZsVZfq1_0),.clk(gclk));
	jdff dff_A_R1GJVanS7_2(.dout(w_dff_A_3v28Pjlo6_0),.din(w_dff_A_R1GJVanS7_2),.clk(gclk));
	jdff dff_A_3v28Pjlo6_0(.dout(w_dff_A_b8K0qLE62_0),.din(w_dff_A_3v28Pjlo6_0),.clk(gclk));
	jdff dff_A_b8K0qLE62_0(.dout(w_dff_A_BTi0qHKI5_0),.din(w_dff_A_b8K0qLE62_0),.clk(gclk));
	jdff dff_A_BTi0qHKI5_0(.dout(w_dff_A_e3LTPdoj2_0),.din(w_dff_A_BTi0qHKI5_0),.clk(gclk));
	jdff dff_A_e3LTPdoj2_0(.dout(w_dff_A_2BCrTTh28_0),.din(w_dff_A_e3LTPdoj2_0),.clk(gclk));
	jdff dff_A_2BCrTTh28_0(.dout(w_dff_A_uHLLDC1h5_0),.din(w_dff_A_2BCrTTh28_0),.clk(gclk));
	jdff dff_A_uHLLDC1h5_0(.dout(w_dff_A_hHnDGNkM0_0),.din(w_dff_A_uHLLDC1h5_0),.clk(gclk));
	jdff dff_A_hHnDGNkM0_0(.dout(w_dff_A_atHNo8x77_0),.din(w_dff_A_hHnDGNkM0_0),.clk(gclk));
	jdff dff_A_atHNo8x77_0(.dout(w_dff_A_TjjxhGX70_0),.din(w_dff_A_atHNo8x77_0),.clk(gclk));
	jdff dff_A_TjjxhGX70_0(.dout(w_dff_A_F7tNoc4t7_0),.din(w_dff_A_TjjxhGX70_0),.clk(gclk));
	jdff dff_A_F7tNoc4t7_0(.dout(w_dff_A_02XtJSan5_0),.din(w_dff_A_F7tNoc4t7_0),.clk(gclk));
	jdff dff_A_02XtJSan5_0(.dout(w_dff_A_JRDzSJiE3_0),.din(w_dff_A_02XtJSan5_0),.clk(gclk));
	jdff dff_A_JRDzSJiE3_0(.dout(w_dff_A_RfVujGfb7_0),.din(w_dff_A_JRDzSJiE3_0),.clk(gclk));
	jdff dff_A_RfVujGfb7_0(.dout(w_dff_A_PL7iiSe06_0),.din(w_dff_A_RfVujGfb7_0),.clk(gclk));
	jdff dff_A_PL7iiSe06_0(.dout(w_dff_A_NBRDja6d9_0),.din(w_dff_A_PL7iiSe06_0),.clk(gclk));
	jdff dff_A_NBRDja6d9_0(.dout(w_dff_A_9O6Idaah6_0),.din(w_dff_A_NBRDja6d9_0),.clk(gclk));
	jdff dff_A_9O6Idaah6_0(.dout(w_dff_A_H5TRvcPw8_0),.din(w_dff_A_9O6Idaah6_0),.clk(gclk));
	jdff dff_A_H5TRvcPw8_0(.dout(w_dff_A_1mp9vioA7_0),.din(w_dff_A_H5TRvcPw8_0),.clk(gclk));
	jdff dff_A_1mp9vioA7_0(.dout(G450gat),.din(w_dff_A_1mp9vioA7_0),.clk(gclk));
	jdff dff_A_LvQP9xlj5_2(.dout(w_dff_A_tLfWjOPN7_0),.din(w_dff_A_LvQP9xlj5_2),.clk(gclk));
	jdff dff_A_tLfWjOPN7_0(.dout(w_dff_A_M8z8ftOG6_0),.din(w_dff_A_tLfWjOPN7_0),.clk(gclk));
	jdff dff_A_M8z8ftOG6_0(.dout(w_dff_A_lNhERKjM8_0),.din(w_dff_A_M8z8ftOG6_0),.clk(gclk));
	jdff dff_A_lNhERKjM8_0(.dout(w_dff_A_tQKRItzr2_0),.din(w_dff_A_lNhERKjM8_0),.clk(gclk));
	jdff dff_A_tQKRItzr2_0(.dout(w_dff_A_RZKfr7rY2_0),.din(w_dff_A_tQKRItzr2_0),.clk(gclk));
	jdff dff_A_RZKfr7rY2_0(.dout(w_dff_A_ssCfw2zJ8_0),.din(w_dff_A_RZKfr7rY2_0),.clk(gclk));
	jdff dff_A_ssCfw2zJ8_0(.dout(w_dff_A_TvZkicBx4_0),.din(w_dff_A_ssCfw2zJ8_0),.clk(gclk));
	jdff dff_A_TvZkicBx4_0(.dout(w_dff_A_CSpgTGcP4_0),.din(w_dff_A_TvZkicBx4_0),.clk(gclk));
	jdff dff_A_CSpgTGcP4_0(.dout(w_dff_A_b0r2iFMB7_0),.din(w_dff_A_CSpgTGcP4_0),.clk(gclk));
	jdff dff_A_b0r2iFMB7_0(.dout(w_dff_A_6dHyje1g9_0),.din(w_dff_A_b0r2iFMB7_0),.clk(gclk));
	jdff dff_A_6dHyje1g9_0(.dout(w_dff_A_fepdQ3Ka4_0),.din(w_dff_A_6dHyje1g9_0),.clk(gclk));
	jdff dff_A_fepdQ3Ka4_0(.dout(w_dff_A_oe72zPQP5_0),.din(w_dff_A_fepdQ3Ka4_0),.clk(gclk));
	jdff dff_A_oe72zPQP5_0(.dout(w_dff_A_f40m703a5_0),.din(w_dff_A_oe72zPQP5_0),.clk(gclk));
	jdff dff_A_f40m703a5_0(.dout(w_dff_A_mZmqsYz20_0),.din(w_dff_A_f40m703a5_0),.clk(gclk));
	jdff dff_A_mZmqsYz20_0(.dout(w_dff_A_Pk8fqNE29_0),.din(w_dff_A_mZmqsYz20_0),.clk(gclk));
	jdff dff_A_Pk8fqNE29_0(.dout(w_dff_A_hNmiyPSM6_0),.din(w_dff_A_Pk8fqNE29_0),.clk(gclk));
	jdff dff_A_hNmiyPSM6_0(.dout(G767gat),.din(w_dff_A_hNmiyPSM6_0),.clk(gclk));
	jdff dff_A_0r3C9dNv8_2(.dout(w_dff_A_Mc5hPslK9_0),.din(w_dff_A_0r3C9dNv8_2),.clk(gclk));
	jdff dff_A_Mc5hPslK9_0(.dout(w_dff_A_eH3k3LpP5_0),.din(w_dff_A_Mc5hPslK9_0),.clk(gclk));
	jdff dff_A_eH3k3LpP5_0(.dout(w_dff_A_ypaW0iCC9_0),.din(w_dff_A_eH3k3LpP5_0),.clk(gclk));
	jdff dff_A_ypaW0iCC9_0(.dout(w_dff_A_hkqX09064_0),.din(w_dff_A_ypaW0iCC9_0),.clk(gclk));
	jdff dff_A_hkqX09064_0(.dout(w_dff_A_FDkR9MnI9_0),.din(w_dff_A_hkqX09064_0),.clk(gclk));
	jdff dff_A_FDkR9MnI9_0(.dout(w_dff_A_TS5Kuw7M7_0),.din(w_dff_A_FDkR9MnI9_0),.clk(gclk));
	jdff dff_A_TS5Kuw7M7_0(.dout(w_dff_A_pxVKceKG3_0),.din(w_dff_A_TS5Kuw7M7_0),.clk(gclk));
	jdff dff_A_pxVKceKG3_0(.dout(w_dff_A_8ofwVCIM1_0),.din(w_dff_A_pxVKceKG3_0),.clk(gclk));
	jdff dff_A_8ofwVCIM1_0(.dout(w_dff_A_vOrzP7sF6_0),.din(w_dff_A_8ofwVCIM1_0),.clk(gclk));
	jdff dff_A_vOrzP7sF6_0(.dout(w_dff_A_ci6z7g5X6_0),.din(w_dff_A_vOrzP7sF6_0),.clk(gclk));
	jdff dff_A_ci6z7g5X6_0(.dout(w_dff_A_F19in5ad1_0),.din(w_dff_A_ci6z7g5X6_0),.clk(gclk));
	jdff dff_A_F19in5ad1_0(.dout(w_dff_A_LBMcHvg94_0),.din(w_dff_A_F19in5ad1_0),.clk(gclk));
	jdff dff_A_LBMcHvg94_0(.dout(w_dff_A_QDsrD8c49_0),.din(w_dff_A_LBMcHvg94_0),.clk(gclk));
	jdff dff_A_QDsrD8c49_0(.dout(w_dff_A_VY2Sqll62_0),.din(w_dff_A_QDsrD8c49_0),.clk(gclk));
	jdff dff_A_VY2Sqll62_0(.dout(w_dff_A_TDRq9fEl1_0),.din(w_dff_A_VY2Sqll62_0),.clk(gclk));
	jdff dff_A_TDRq9fEl1_0(.dout(w_dff_A_labbdHJQ5_0),.din(w_dff_A_TDRq9fEl1_0),.clk(gclk));
	jdff dff_A_labbdHJQ5_0(.dout(G768gat),.din(w_dff_A_labbdHJQ5_0),.clk(gclk));
	jdff dff_A_NdwaEkVp4_2(.dout(w_dff_A_iFhP6lex2_0),.din(w_dff_A_NdwaEkVp4_2),.clk(gclk));
	jdff dff_A_iFhP6lex2_0(.dout(w_dff_A_wR1Kedpq4_0),.din(w_dff_A_iFhP6lex2_0),.clk(gclk));
	jdff dff_A_wR1Kedpq4_0(.dout(w_dff_A_pB1RTRaH4_0),.din(w_dff_A_wR1Kedpq4_0),.clk(gclk));
	jdff dff_A_pB1RTRaH4_0(.dout(w_dff_A_qLrAg3sh5_0),.din(w_dff_A_pB1RTRaH4_0),.clk(gclk));
	jdff dff_A_qLrAg3sh5_0(.dout(w_dff_A_oZJQVz7Q7_0),.din(w_dff_A_qLrAg3sh5_0),.clk(gclk));
	jdff dff_A_oZJQVz7Q7_0(.dout(w_dff_A_TyT9jA6O1_0),.din(w_dff_A_oZJQVz7Q7_0),.clk(gclk));
	jdff dff_A_TyT9jA6O1_0(.dout(w_dff_A_9uLBxE1F1_0),.din(w_dff_A_TyT9jA6O1_0),.clk(gclk));
	jdff dff_A_9uLBxE1F1_0(.dout(G850gat),.din(w_dff_A_9uLBxE1F1_0),.clk(gclk));
	jdff dff_A_TtRDAdvq8_2(.dout(w_dff_A_Bj362FUu5_0),.din(w_dff_A_TtRDAdvq8_2),.clk(gclk));
	jdff dff_A_Bj362FUu5_0(.dout(w_dff_A_DOjFwhZ78_0),.din(w_dff_A_Bj362FUu5_0),.clk(gclk));
	jdff dff_A_DOjFwhZ78_0(.dout(w_dff_A_TBwLhrZr3_0),.din(w_dff_A_DOjFwhZ78_0),.clk(gclk));
	jdff dff_A_TBwLhrZr3_0(.dout(G863gat),.din(w_dff_A_TBwLhrZr3_0),.clk(gclk));
	jdff dff_A_rFZzsmmR5_2(.dout(w_dff_A_WqAF288w0_0),.din(w_dff_A_rFZzsmmR5_2),.clk(gclk));
	jdff dff_A_WqAF288w0_0(.dout(w_dff_A_s6veoO8B6_0),.din(w_dff_A_WqAF288w0_0),.clk(gclk));
	jdff dff_A_s6veoO8B6_0(.dout(w_dff_A_Ea6N4bL97_0),.din(w_dff_A_s6veoO8B6_0),.clk(gclk));
	jdff dff_A_Ea6N4bL97_0(.dout(G864gat),.din(w_dff_A_Ea6N4bL97_0),.clk(gclk));
	jdff dff_A_41kHcAp74_2(.dout(w_dff_A_BJkn4WKK8_0),.din(w_dff_A_41kHcAp74_2),.clk(gclk));
	jdff dff_A_BJkn4WKK8_0(.dout(w_dff_A_t3OCBdPy5_0),.din(w_dff_A_BJkn4WKK8_0),.clk(gclk));
	jdff dff_A_t3OCBdPy5_0(.dout(w_dff_A_bNeQcsHg1_0),.din(w_dff_A_t3OCBdPy5_0),.clk(gclk));
	jdff dff_A_bNeQcsHg1_0(.dout(w_dff_A_M5pyrNgW0_0),.din(w_dff_A_bNeQcsHg1_0),.clk(gclk));
	jdff dff_A_M5pyrNgW0_0(.dout(w_dff_A_HDpeWK6g8_0),.din(w_dff_A_M5pyrNgW0_0),.clk(gclk));
	jdff dff_A_HDpeWK6g8_0(.dout(G865gat),.din(w_dff_A_HDpeWK6g8_0),.clk(gclk));
	jdff dff_A_By0Ov4MX1_2(.dout(w_dff_A_Sp6MW25y5_0),.din(w_dff_A_By0Ov4MX1_2),.clk(gclk));
	jdff dff_A_Sp6MW25y5_0(.dout(G866gat),.din(w_dff_A_Sp6MW25y5_0),.clk(gclk));
	jdff dff_A_t7xpMCTX3_2(.dout(w_dff_A_Y6yi8leE7_0),.din(w_dff_A_t7xpMCTX3_2),.clk(gclk));
	jdff dff_A_Y6yi8leE7_0(.dout(G874gat),.din(w_dff_A_Y6yi8leE7_0),.clk(gclk));
endmodule

