/*

c880:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jdff: 1588
	jand: 151
	jor: 122

Summary:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jdff: 1588
	jand: 151
	jor: 122
*/

module c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n103;
	wire n104;
	wire n105;
	wire n107;
	wire n108;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n119;
	wire n120;
	wire n122;
	wire n123;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire [2:0] w_G1gat_0;
	wire [1:0] w_G1gat_1;
	wire [1:0] w_G8gat_0;
	wire [1:0] w_G13gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G17gat_1;
	wire [2:0] w_G17gat_2;
	wire [1:0] w_G26gat_0;
	wire [2:0] w_G29gat_0;
	wire [1:0] w_G36gat_0;
	wire [2:0] w_G42gat_0;
	wire [2:0] w_G42gat_1;
	wire [1:0] w_G42gat_2;
	wire [2:0] w_G51gat_0;
	wire [1:0] w_G51gat_1;
	wire [2:0] w_G55gat_0;
	wire [2:0] w_G59gat_0;
	wire [1:0] w_G59gat_1;
	wire [1:0] w_G68gat_0;
	wire [1:0] w_G75gat_0;
	wire [2:0] w_G80gat_0;
	wire [2:0] w_G91gat_0;
	wire [2:0] w_G96gat_0;
	wire [2:0] w_G101gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G111gat_0;
	wire [2:0] w_G116gat_0;
	wire [2:0] w_G121gat_0;
	wire [2:0] w_G126gat_0;
	wire [1:0] w_G130gat_0;
	wire [2:0] w_G138gat_0;
	wire [1:0] w_G138gat_1;
	wire [1:0] w_G143gat_0;
	wire [1:0] w_G146gat_0;
	wire [1:0] w_G149gat_0;
	wire [2:0] w_G153gat_0;
	wire [1:0] w_G156gat_0;
	wire [2:0] w_G159gat_0;
	wire [2:0] w_G159gat_1;
	wire [2:0] w_G165gat_0;
	wire [2:0] w_G165gat_1;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [2:0] w_G177gat_0;
	wire [2:0] w_G177gat_1;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G183gat_1;
	wire [2:0] w_G189gat_0;
	wire [2:0] w_G189gat_1;
	wire [1:0] w_G189gat_2;
	wire [2:0] w_G195gat_0;
	wire [2:0] w_G195gat_1;
	wire [1:0] w_G195gat_2;
	wire [2:0] w_G201gat_0;
	wire [1:0] w_G201gat_1;
	wire [2:0] w_G210gat_0;
	wire [2:0] w_G210gat_1;
	wire [2:0] w_G210gat_2;
	wire [1:0] w_G210gat_3;
	wire [2:0] w_G219gat_0;
	wire [2:0] w_G219gat_1;
	wire [2:0] w_G219gat_2;
	wire [2:0] w_G219gat_3;
	wire [2:0] w_G228gat_0;
	wire [2:0] w_G228gat_1;
	wire [2:0] w_G228gat_2;
	wire [1:0] w_G228gat_3;
	wire [2:0] w_G237gat_0;
	wire [2:0] w_G237gat_1;
	wire [2:0] w_G237gat_2;
	wire [1:0] w_G237gat_3;
	wire [2:0] w_G246gat_0;
	wire [2:0] w_G246gat_1;
	wire [2:0] w_G246gat_2;
	wire [1:0] w_G246gat_3;
	wire [2:0] w_G255gat_0;
	wire [2:0] w_G261gat_0;
	wire [1:0] w_G268gat_0;
	wire [1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire [2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire [1:0] w_n86_0;
	wire [1:0] w_n88_0;
	wire [1:0] w_n92_0;
	wire [1:0] w_n93_0;
	wire [2:0] w_n95_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n109_0;
	wire [1:0] w_n111_0;
	wire [1:0] w_n113_0;
	wire [2:0] w_n119_0;
	wire [1:0] w_n122_0;
	wire [1:0] w_n144_0;
	wire [1:0] w_n146_0;
	wire [2:0] w_n148_0;
	wire [2:0] w_n148_1;
	wire [1:0] w_n149_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n152_0;
	wire [1:0] w_n162_0;
	wire [2:0] w_n164_0;
	wire [2:0] w_n164_1;
	wire [2:0] w_n164_2;
	wire [1:0] w_n164_3;
	wire [1:0] w_n167_0;
	wire [1:0] w_n168_0;
	wire [2:0] w_n170_0;
	wire [1:0] w_n170_1;
	wire [1:0] w_n173_0;
	wire [2:0] w_n178_0;
	wire [2:0] w_n178_1;
	wire [2:0] w_n178_2;
	wire [1:0] w_n178_3;
	wire [2:0] w_n181_0;
	wire [1:0] w_n185_0;
	wire [2:0] w_n197_0;
	wire [2:0] w_n198_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n209_0;
	wire [2:0] w_n218_0;
	wire [1:0] w_n218_1;
	wire [2:0] w_n219_0;
	wire [2:0] w_n222_0;
	wire [2:0] w_n233_0;
	wire [1:0] w_n233_1;
	wire [1:0] w_n234_0;
	wire [1:0] w_n235_0;
	wire [2:0] w_n239_0;
	wire [1:0] w_n239_1;
	wire [1:0] w_n240_0;
	wire [1:0] w_n241_0;
	wire [1:0] w_n242_0;
	wire [1:0] w_n245_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n258_0;
	wire [1:0] w_n260_0;
	wire [1:0] w_n262_0;
	wire [2:0] w_n267_0;
	wire [2:0] w_n285_0;
	wire [2:0] w_n303_0;
	wire [1:0] w_n303_1;
	wire [2:0] w_n306_0;
	wire [1:0] w_n306_1;
	wire [2:0] w_n311_0;
	wire [2:0] w_n311_1;
	wire [2:0] w_n319_0;
	wire [2:0] w_n319_1;
	wire [1:0] w_n320_0;
	wire [1:0] w_n321_0;
	wire [2:0] w_n327_0;
	wire [2:0] w_n327_1;
	wire [1:0] w_n328_0;
	wire [1:0] w_n329_0;
	wire [2:0] w_n335_0;
	wire [1:0] w_n335_1;
	wire [2:0] w_n336_0;
	wire [1:0] w_n339_0;
	wire [1:0] w_n343_0;
	wire [1:0] w_n346_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n350_0;
	wire [1:0] w_n352_0;
	wire [1:0] w_n355_0;
	wire [1:0] w_n361_0;
	wire [2:0] w_n377_0;
	wire [1:0] w_n391_0;
	wire [1:0] w_n393_0;
	wire [2:0] w_n404_0;
	wire [2:0] w_n420_0;
	wire w_dff_B_xgt7oxkw4_2;
	wire w_dff_B_aBFOmxD08_1;
	wire w_dff_B_hW8Se1yu8_1;
	wire w_dff_B_owR0xsDs9_1;
	wire w_dff_A_oxB3695r7_1;
	wire w_dff_A_rew4hahm7_1;
	wire w_dff_B_Skdtk8Un0_1;
	wire w_dff_B_5UUizARO8_1;
	wire w_dff_B_aKz1ZNkd5_1;
	wire w_dff_B_JOj0NCKz0_1;
	wire w_dff_B_iA0hOQEb1_1;
	wire w_dff_B_EATIr7JD0_1;
	wire w_dff_B_znr3Y1ok4_1;
	wire w_dff_A_QyOVgLYl6_1;
	wire w_dff_B_R2xzlhF02_1;
	wire w_dff_B_JS1LUrZv1_1;
	wire w_dff_B_8VdP2dtW9_1;
	wire w_dff_B_CEQ0uHYm7_1;
	wire w_dff_B_xWZxn00B9_1;
	wire w_dff_B_B7wikmcL3_1;
	wire w_dff_B_KEyhOJQ37_0;
	wire w_dff_B_ZUokzprQ2_0;
	wire w_dff_B_ULczbqEV6_0;
	wire w_dff_B_Ac0ERhlf8_0;
	wire w_dff_B_6x74zz1B1_0;
	wire w_dff_B_x4rpQqzp7_0;
	wire w_dff_B_go5S0cmU4_0;
	wire w_dff_B_bZEgn9VB7_0;
	wire w_dff_B_8At1OGb22_0;
	wire w_dff_B_Ff6YlyyZ8_0;
	wire w_dff_B_hoMlVHfk7_0;
	wire w_dff_B_msmmgGy76_0;
	wire w_dff_B_93RQjyTa9_0;
	wire w_dff_B_rxaWXZwb5_0;
	wire w_dff_A_2qre1vtb0_0;
	wire w_dff_A_3sQMLgiR6_0;
	wire w_dff_A_S4nVfOFY5_0;
	wire w_dff_A_s18ggExM6_0;
	wire w_dff_B_adwAZrNl7_1;
	wire w_dff_B_9STfpRbb1_1;
	wire w_dff_B_XVpX5orf8_1;
	wire w_dff_B_Aj6bGocO9_1;
	wire w_dff_B_UuHxarYi1_1;
	wire w_dff_B_KIRMF6B32_1;
	wire w_dff_B_qxPgZkMo9_1;
	wire w_dff_B_D54inTRd9_1;
	wire w_dff_B_3r0BZzul0_1;
	wire w_dff_B_xOF3U8Xw3_1;
	wire w_dff_B_wQZuk2hL6_1;
	wire w_dff_B_XUaNJjtM9_1;
	wire w_dff_B_q38WAzoI3_1;
	wire w_dff_B_E03aGQNB0_1;
	wire w_dff_B_qB1Nkhzo7_1;
	wire w_dff_B_AOd4uBUG8_1;
	wire w_dff_B_GMQ21RxZ9_1;
	wire w_dff_B_MfxyW0mO9_1;
	wire w_dff_B_I2iIPerq3_1;
	wire w_dff_B_U9M9dbaP5_1;
	wire w_dff_B_fMTMlvDt8_1;
	wire w_dff_B_Rk0ofG141_0;
	wire w_dff_B_j7bbZSaO0_0;
	wire w_dff_B_HlYbTumq8_0;
	wire w_dff_B_9rO6rsWT1_0;
	wire w_dff_B_mlZQReuw7_0;
	wire w_dff_B_wrUscLWM9_0;
	wire w_dff_B_LdQumMHy9_0;
	wire w_dff_B_FfPcPOOZ2_0;
	wire w_dff_A_m9gDeRoh0_1;
	wire w_dff_A_4EqwaagK7_1;
	wire w_dff_A_jRK70mNr4_1;
	wire w_dff_A_f8WcpeTE4_1;
	wire w_dff_A_jrbqh4QO7_1;
	wire w_dff_A_643Jw5Qk2_1;
	wire w_dff_A_3G8nFk7W0_1;
	wire w_dff_A_YV6a4Gzn5_1;
	wire w_dff_A_WKAyP4vq4_1;
	wire w_dff_A_h6i5PYEH4_0;
	wire w_dff_A_7H5fcfOu9_0;
	wire w_dff_A_nFhN0sVP9_0;
	wire w_dff_A_5wvFnafV4_0;
	wire w_dff_A_LefcYNt21_1;
	wire w_dff_A_fbAfghFz1_1;
	wire w_dff_A_bdjxU63K5_1;
	wire w_dff_A_v4YiKeId8_1;
	wire w_dff_A_r9tAbfMX6_1;
	wire w_dff_A_ePi6SFEE7_1;
	wire w_dff_A_N7RiwQhL7_1;
	wire w_dff_A_Vael7ZcZ0_1;
	wire w_dff_A_Qw9v7Yie2_1;
	wire w_dff_B_sKPLjkxx7_1;
	wire w_dff_B_zvKx1LYf9_1;
	wire w_dff_B_QquYyicl0_1;
	wire w_dff_B_dDHrJEG72_1;
	wire w_dff_B_aisV8IiX3_1;
	wire w_dff_B_P64uaEJY4_1;
	wire w_dff_B_OdOP9BaB7_0;
	wire w_dff_B_o5XWamel1_0;
	wire w_dff_B_TKok4g8s0_0;
	wire w_dff_B_EckWqqYc5_0;
	wire w_dff_A_6ghpfoia9_0;
	wire w_dff_A_JzkKiM653_0;
	wire w_dff_A_ShCjBaep4_0;
	wire w_dff_A_hkrrthH71_1;
	wire w_dff_A_GPFa31IZ2_1;
	wire w_dff_A_DmJiZkl84_1;
	wire w_dff_A_ljdrSe2b7_1;
	wire w_dff_A_u2etzkMM4_1;
	wire w_dff_B_ip1O69zR9_1;
	wire w_dff_B_NF73eS3m0_0;
	wire w_dff_B_FgjDBKvU8_0;
	wire w_dff_B_pcuzcSUF9_0;
	wire w_dff_B_guoqX5rk6_0;
	wire w_dff_B_L9INqjsN8_1;
	wire w_dff_B_ZTZ7NpMe5_1;
	wire w_dff_B_oFAamp7l3_1;
	wire w_dff_B_6FXB3G1w8_1;
	wire w_dff_B_tbSerfKW1_1;
	wire w_dff_B_x36CsGqm2_1;
	wire w_dff_B_lBCbBLRQ2_1;
	wire w_dff_B_hb7M47we2_1;
	wire w_dff_B_xIvQHfp88_1;
	wire w_dff_B_BpUY3SjG5_1;
	wire w_dff_B_CcvYoYiK1_1;
	wire w_dff_B_doc87SNp3_1;
	wire w_dff_B_oHF4b3lP0_0;
	wire w_dff_B_8RYN9yIv4_0;
	wire w_dff_B_6cfMoPDX4_0;
	wire w_dff_B_fds7y00t6_0;
	wire w_dff_B_NDQPL4Cb3_0;
	wire w_dff_B_MwAU5TSD8_0;
	wire w_dff_A_G4FIs4pM6_1;
	wire w_dff_A_766102Ba8_1;
	wire w_dff_A_szlXohlj8_1;
	wire w_dff_A_em7gfIqr1_1;
	wire w_dff_A_oIwOpkCN4_1;
	wire w_dff_B_q38OqGB28_1;
	wire w_dff_B_dkizGsDs2_1;
	wire w_dff_B_sBXG36rQ5_1;
	wire w_dff_B_iNv189Yf9_1;
	wire w_dff_B_otlZuYIa1_0;
	wire w_dff_B_kH9ZOFXQ2_0;
	wire w_dff_B_ndu5LyJR1_1;
	wire w_dff_B_DTIFOlka2_0;
	wire w_dff_B_ezlAstUf3_0;
	wire w_dff_B_Zwr92fFJ9_0;
	wire w_dff_B_hXPlE1Gb5_0;
	wire w_dff_B_MCIkRQmJ4_0;
	wire w_dff_B_83HV8bV64_0;
	wire w_dff_B_i2P4lSKr4_0;
	wire w_dff_B_MyHsY2ym2_0;
	wire w_dff_B_0kDBjHJ52_1;
	wire w_dff_B_OUn71ubv4_1;
	wire w_dff_B_bYnvctjA7_1;
	wire w_dff_B_Cad6sX8N2_1;
	wire w_dff_B_G8BxU8L91_1;
	wire w_dff_B_HyOFN1pt4_1;
	wire w_dff_B_x0l3AsoL5_1;
	wire w_dff_B_vvj0HpDe2_1;
	wire w_dff_B_ckZOUTVT5_0;
	wire w_dff_B_VZfyjC3l4_0;
	wire w_dff_B_bHfCrVa15_0;
	wire w_dff_B_vTOh8UrP3_0;
	wire w_dff_B_BNahH4ob8_0;
	wire w_dff_B_FRm0f71R6_0;
	wire w_dff_A_z66bwLQm1_1;
	wire w_dff_A_FUPxMvZA0_1;
	wire w_dff_A_2sd0l6IR0_1;
	wire w_dff_B_GlXyYwwF9_1;
	wire w_dff_B_O50J3Kuq4_1;
	wire w_dff_B_xhdjv0j25_1;
	wire w_dff_B_T3bizIL53_1;
	wire w_dff_B_6o2QfV8Y8_1;
	wire w_dff_B_OnAOBO4L8_1;
	wire w_dff_B_WzVg6u1J8_1;
	wire w_dff_B_fQrFZnXJ4_1;
	wire w_dff_B_sijGcggi2_1;
	wire w_dff_B_So5b2yCD8_1;
	wire w_dff_B_UC0JnjnF7_1;
	wire w_dff_B_3I2iOSIa8_1;
	wire w_dff_B_uiLMbmCC7_1;
	wire w_dff_B_2qo0lXRl2_1;
	wire w_dff_B_YPDy7Iun2_1;
	wire w_dff_B_nSMC28Oa8_1;
	wire w_dff_B_xy6Fhd6t4_1;
	wire w_dff_B_EsqRNlVT9_1;
	wire w_dff_B_FI15eL6y1_1;
	wire w_dff_B_yfNz41jq9_1;
	wire w_dff_B_CDwawG0x0_1;
	wire w_dff_B_Kak8VqjB7_1;
	wire w_dff_B_jvMGe37M4_1;
	wire w_dff_B_QNnKLkjF5_1;
	wire w_dff_B_Jrd7GfwQ2_1;
	wire w_dff_B_NxdZk2vU0_1;
	wire w_dff_B_9ML7OhUv7_1;
	wire w_dff_B_Or1qyz1f0_1;
	wire w_dff_B_t1cU3XPa1_1;
	wire w_dff_A_xa2Lgavg6_0;
	wire w_dff_A_kGFG3yZG0_0;
	wire w_dff_A_PO5kjd967_0;
	wire w_dff_A_fLCaUrrJ5_0;
	wire w_dff_A_9ShXdnnB2_0;
	wire w_dff_A_IitPTuNO5_0;
	wire w_dff_A_n88HvGkE6_0;
	wire w_dff_A_J7UmDh821_0;
	wire w_dff_A_VPQapodH2_0;
	wire w_dff_A_FaO2ZNUX8_1;
	wire w_dff_A_atznSj4f2_1;
	wire w_dff_A_LveJbCk61_1;
	wire w_dff_A_10HSazra1_1;
	wire w_dff_A_FOzdQjo31_1;
	wire w_dff_A_XE1efOH42_1;
	wire w_dff_A_QMoXbwDy4_1;
	wire w_dff_A_YLv8NwLR8_1;
	wire w_dff_A_uXT30LP58_1;
	wire w_dff_B_DrWmOQ3G4_1;
	wire w_dff_B_SKllqSYH9_1;
	wire w_dff_B_m1586m9L8_0;
	wire w_dff_B_bLv1pV2j0_0;
	wire w_dff_B_93XyzLj32_0;
	wire w_dff_B_ctxjP86f9_0;
	wire w_dff_B_VpIXfvx32_0;
	wire w_dff_B_0GLwW4iA8_0;
	wire w_dff_B_Yk3VSakW1_0;
	wire w_dff_B_UDCLH5u87_0;
	wire w_dff_B_jrM5SpFM8_0;
	wire w_dff_B_T6ij8MWk3_0;
	wire w_dff_B_lq8hkTeu3_0;
	wire w_dff_B_orXl8P786_0;
	wire w_dff_B_wSRGaJsQ8_0;
	wire w_dff_B_kHaLqff29_1;
	wire w_dff_B_pRwP6pur1_1;
	wire w_dff_B_MjAmgKrD6_1;
	wire w_dff_B_q1deCKrm8_1;
	wire w_dff_A_2HqWG7O22_0;
	wire w_dff_A_kFtHrzAs3_0;
	wire w_dff_A_Gn4qwCi11_0;
	wire w_dff_A_yYwnJvjr0_0;
	wire w_dff_A_DZFSmrXP2_0;
	wire w_dff_A_bdFVGDSr6_0;
	wire w_dff_A_5hhDTQ4c6_0;
	wire w_dff_A_aSHbGEry9_0;
	wire w_dff_A_L8CM89wd5_0;
	wire w_dff_A_2mFXpMH17_0;
	wire w_dff_A_SL4FOWtT3_0;
	wire w_dff_A_ftrUmz822_0;
	wire w_dff_A_SFjHUcDx2_0;
	wire w_dff_A_nkTGWDF62_0;
	wire w_dff_A_b0gMc3W59_0;
	wire w_dff_A_eIovaeni1_0;
	wire w_dff_A_TfdjTBKt4_0;
	wire w_dff_A_NMD8Frsu5_0;
	wire w_dff_A_dfJLx5UD0_0;
	wire w_dff_A_dl7XLRC63_0;
	wire w_dff_A_OGL0MYyQ1_0;
	wire w_dff_A_5xc0eiyF9_0;
	wire w_dff_A_ZoeQule85_0;
	wire w_dff_A_ZNMvC3Ml1_0;
	wire w_dff_A_H1ADnFNM4_0;
	wire w_dff_A_RJJIUzRJ7_0;
	wire w_dff_A_qXgjvMms3_0;
	wire w_dff_A_cLdcIYs66_0;
	wire w_dff_B_Aq2UPSvS2_1;
	wire w_dff_B_YuDzUN6G6_1;
	wire w_dff_B_fBJRcelf6_1;
	wire w_dff_B_W4KZWh1j7_1;
	wire w_dff_B_shyw5PxS2_1;
	wire w_dff_B_euqnkUns6_1;
	wire w_dff_B_SLBiKYnm0_1;
	wire w_dff_B_6IKmdFBU2_1;
	wire w_dff_A_4bpxj24S7_0;
	wire w_dff_A_p5mQNXnX6_0;
	wire w_dff_A_rufeLn5R4_0;
	wire w_dff_A_Qtn3LZ9u7_0;
	wire w_dff_A_5bL57tID5_0;
	wire w_dff_A_cu6TzZTx5_1;
	wire w_dff_A_khgA3j7b9_1;
	wire w_dff_A_fcPCOdj53_1;
	wire w_dff_A_zr0Rae5B3_1;
	wire w_dff_A_wAl3WvJh8_1;
	wire w_dff_A_bEu2IV3Q4_0;
	wire w_dff_A_LtHueLH54_0;
	wire w_dff_A_uiMiqTwk7_0;
	wire w_dff_A_hxyWqPOB8_0;
	wire w_dff_A_7eLuDSf10_0;
	wire w_dff_A_Qb8ZzWj45_0;
	wire w_dff_A_92DFYHGG1_0;
	wire w_dff_A_50mAV60x7_0;
	wire w_dff_A_xHyMAU8u8_0;
	wire w_dff_A_FJFDQy9s7_0;
	wire w_dff_B_SXDplQRF6_1;
	wire w_dff_B_1eSM8wuX0_1;
	wire w_dff_B_ZKtxgBCx1_1;
	wire w_dff_B_ZPMoxhe70_1;
	wire w_dff_B_jASMbCkU1_1;
	wire w_dff_B_q4sDnhd28_1;
	wire w_dff_B_qnyZVeN43_1;
	wire w_dff_B_RhbtftjB8_1;
	wire w_dff_B_WJy5GkCG8_1;
	wire w_dff_B_jf9djXIB7_1;
	wire w_dff_B_5osexZ1Z7_1;
	wire w_dff_B_TMtZInnr4_1;
	wire w_dff_B_Eiyg7v3H6_1;
	wire w_dff_B_L92F2ZAH0_1;
	wire w_dff_B_jZOQOToS4_0;
	wire w_dff_B_1GT3auXp9_0;
	wire w_dff_B_AkeX8Jwn1_0;
	wire w_dff_B_6e3ZrFcL9_0;
	wire w_dff_B_GcvQsw8u4_0;
	wire w_dff_B_JC9M4Qdx4_0;
	wire w_dff_B_5Hfh4XDf6_0;
	wire w_dff_B_1mMqJSg65_0;
	wire w_dff_B_ufGA5QdL5_0;
	wire w_dff_B_9cY5hey30_0;
	wire w_dff_B_W8k17x5l3_0;
	wire w_dff_B_CvMGc4DV2_0;
	wire w_dff_B_zAgfXo5z3_0;
	wire w_dff_B_NYJdjsi79_1;
	wire w_dff_B_njk6QFK41_1;
	wire w_dff_B_rmPoUPLP4_1;
	wire w_dff_B_timix9rN1_1;
	wire w_dff_B_mrW6U2kI1_1;
	wire w_dff_B_YdvDzPAu6_1;
	wire w_dff_B_tvnE0rJr4_1;
	wire w_dff_B_tU4ZQYkN7_1;
	wire w_dff_B_nExStRYp5_1;
	wire w_dff_B_CpYOMRyJ5_1;
	wire w_dff_B_63BKISQi8_1;
	wire w_dff_B_a428seju5_1;
	wire w_dff_B_hMkxnIK09_1;
	wire w_dff_B_bCycd5jY6_1;
	wire w_dff_B_oAspcJrA0_1;
	wire w_dff_B_BPa9AnFI5_1;
	wire w_dff_B_G5PVtizS6_1;
	wire w_dff_B_AdIRQnOQ6_1;
	wire w_dff_B_3ao02iZo0_1;
	wire w_dff_B_vv7mdAgE4_1;
	wire w_dff_B_zEVtMg1H1_1;
	wire w_dff_B_dFp1mONK0_1;
	wire w_dff_B_Bo7oQoJK8_1;
	wire w_dff_A_Z22eqk216_1;
	wire w_dff_A_jiCiVtNY1_1;
	wire w_dff_A_NoLqKbR40_1;
	wire w_dff_A_j2w1C8PV1_1;
	wire w_dff_A_OEV2ulpJ1_1;
	wire w_dff_A_4lxNdACi7_1;
	wire w_dff_A_hPY5Y3Tl6_1;
	wire w_dff_A_XpHyiiBG8_1;
	wire w_dff_A_7qAWTxjC0_1;
	wire w_dff_A_lq6Ms2402_1;
	wire w_dff_A_c55AXmE41_1;
	wire w_dff_A_axQuh9PX7_1;
	wire w_dff_A_KbNxnfNW8_1;
	wire w_dff_A_Dbzozypn5_1;
	wire w_dff_A_EHVMy5Wb4_1;
	wire w_dff_A_BfUMS4cX4_1;
	wire w_dff_A_yVJlEyFT5_1;
	wire w_dff_A_Ej67evNU6_1;
	wire w_dff_A_Yzu5lBv14_1;
	wire w_dff_A_OdjLpzgq4_1;
	wire w_dff_A_WllzbeKy3_1;
	wire w_dff_A_VEBjHC828_1;
	wire w_dff_A_cKccF6vN3_1;
	wire w_dff_A_Dhk20cVU2_1;
	wire w_dff_A_40zSHeLb7_1;
	wire w_dff_A_JfZmhdgi8_0;
	wire w_dff_A_FnqWhfS72_0;
	wire w_dff_A_aYvGGn4P1_0;
	wire w_dff_A_N9KhBuqq0_0;
	wire w_dff_A_7umzxTUl5_0;
	wire w_dff_A_9ymrjDGK8_0;
	wire w_dff_A_NrX0Px4Y5_0;
	wire w_dff_A_aBmZ5SFr4_0;
	wire w_dff_A_8DVrXGV59_1;
	wire w_dff_A_3089IQFR8_1;
	wire w_dff_A_I3MyPCLg6_1;
	wire w_dff_A_1Maour7D0_1;
	wire w_dff_A_gutcIJ8Z5_1;
	wire w_dff_A_s4h5kpji8_1;
	wire w_dff_A_rxVNaLEr1_1;
	wire w_dff_A_20PT5cV23_1;
	wire w_dff_B_JdO4DSjG8_1;
	wire w_dff_B_JSqBN6F18_0;
	wire w_dff_B_vMeloIfP0_0;
	wire w_dff_B_u6fypIpY3_0;
	wire w_dff_B_RFArZE4m9_0;
	wire w_dff_B_aZLpfzCF1_0;
	wire w_dff_B_cePgMkB80_0;
	wire w_dff_B_jLU6SnWW2_0;
	wire w_dff_B_2DfuLQwR6_0;
	wire w_dff_B_mwbqMMFu7_0;
	wire w_dff_B_0NpV4Yn56_0;
	wire w_dff_B_jkVBsAco1_0;
	wire w_dff_B_lOKYu5SG3_0;
	wire w_dff_A_k0Uhqvpj9_1;
	wire w_dff_A_wv7Ex7Qj9_1;
	wire w_dff_A_k1HBqoWs4_1;
	wire w_dff_A_L5i2ieyX0_1;
	wire w_dff_A_gq88xnPb3_1;
	wire w_dff_A_8ni1nkcY5_1;
	wire w_dff_A_uoUUwTm15_1;
	wire w_dff_A_iwVYX3Zd3_1;
	wire w_dff_A_rODvyHfY2_1;
	wire w_dff_A_RNiQqSRT5_1;
	wire w_dff_A_e7zit8rx5_1;
	wire w_dff_A_SK0o8WK41_1;
	wire w_dff_A_beWY4Zs84_1;
	wire w_dff_A_kgIBAwiY8_1;
	wire w_dff_B_K8VI0lyJ8_1;
	wire w_dff_B_6jws5gbv6_0;
	wire w_dff_B_IK5EIIq12_0;
	wire w_dff_B_UDCo5pPR4_0;
	wire w_dff_B_Hjzc4SbF0_0;
	wire w_dff_B_hnrTEviD9_0;
	wire w_dff_B_dfoDyUwa0_0;
	wire w_dff_B_VTLnXASP2_1;
	wire w_dff_A_4Zj3AdZQ4_1;
	wire w_dff_A_tAxX9yhZ8_1;
	wire w_dff_A_vHOFF2l25_1;
	wire w_dff_A_TbPeTSzs7_1;
	wire w_dff_A_slZFUKBu2_1;
	wire w_dff_A_xEYgw5BB7_1;
	wire w_dff_A_uHBsdGeX2_1;
	wire w_dff_A_vnmmxkAC4_1;
	wire w_dff_A_Tf2lEuFd3_1;
	wire w_dff_A_kp3nSwIz2_2;
	wire w_dff_A_SeLWDs1C6_2;
	wire w_dff_A_OEU3F7TX7_2;
	wire w_dff_A_uo7l20Uw7_2;
	wire w_dff_A_8bO2taWJ8_2;
	wire w_dff_A_PHUy7fEB4_2;
	wire w_dff_A_ITrY2ZIz0_2;
	wire w_dff_A_omNB1vwN6_2;
	wire w_dff_A_uPQS5i6i4_2;
	wire w_dff_A_k1ee7xNV9_2;
	wire w_dff_A_R0RX7xce5_2;
	wire w_dff_B_eIirSXnc6_1;
	wire w_dff_B_Ky1FXVhY4_1;
	wire w_dff_B_eZTVX8EQ6_1;
	wire w_dff_B_XAbEllva5_1;
	wire w_dff_B_uJkrmF8P6_1;
	wire w_dff_B_roZd3Z9n4_1;
	wire w_dff_B_ycumxEgu4_1;
	wire w_dff_B_O4OyMdAz7_1;
	wire w_dff_B_qlpMLfen2_1;
	wire w_dff_B_X5uVtMo40_1;
	wire w_dff_B_qpsPCDeK3_1;
	wire w_dff_B_2eA68JVH7_1;
	wire w_dff_B_8KdJBbll1_0;
	wire w_dff_B_jxV3Q3h44_0;
	wire w_dff_B_msdHrvXn1_0;
	wire w_dff_B_pyf8G6p62_0;
	wire w_dff_B_qqWdOOx01_0;
	wire w_dff_B_WwYmBD714_0;
	wire w_dff_B_wQwNPLSZ5_0;
	wire w_dff_B_5oGhwwWM8_0;
	wire w_dff_B_eq2dpWGH8_0;
	wire w_dff_B_fOiOfrNH0_0;
	wire w_dff_B_hzZ3zAfb8_0;
	wire w_dff_B_1uRZtwzT1_1;
	wire w_dff_B_MglWwv2W7_1;
	wire w_dff_B_qEwBakl73_1;
	wire w_dff_B_DnLY0apf9_1;
	wire w_dff_B_vNEw1tAV8_1;
	wire w_dff_B_8x6CCG9t3_1;
	wire w_dff_B_19gMOpUe2_1;
	wire w_dff_B_uyb6QbQ87_1;
	wire w_dff_B_paBBHVNr4_1;
	wire w_dff_B_MLzv1ZkU1_1;
	wire w_dff_B_aEbuJ1zi8_1;
	wire w_dff_B_rcqBL7af9_1;
	wire w_dff_B_QQouUaOH4_1;
	wire w_dff_B_FNVWj71O0_1;
	wire w_dff_B_ZWPs6Pbv2_1;
	wire w_dff_B_TWjNr2ld3_1;
	wire w_dff_B_FZd1igRE1_1;
	wire w_dff_B_5ZNWOaTP6_1;
	wire w_dff_B_8w1OuQ7g3_1;
	wire w_dff_A_engRbXKT4_1;
	wire w_dff_A_3oFMPpWl3_1;
	wire w_dff_A_znlV3md30_1;
	wire w_dff_A_5XSnst9T3_1;
	wire w_dff_A_qASWQBJd9_1;
	wire w_dff_A_c4XqH9Jq6_1;
	wire w_dff_A_4p14Z57N8_1;
	wire w_dff_A_1LyHZ4gi4_1;
	wire w_dff_A_eXhgisLy9_1;
	wire w_dff_A_7tkxUkqg0_1;
	wire w_dff_A_wdomqhDh0_1;
	wire w_dff_A_J26MXrAT5_1;
	wire w_dff_A_dHegbbFb7_1;
	wire w_dff_A_v8NB6jfx4_1;
	wire w_dff_A_U98ulfnE3_1;
	wire w_dff_A_sOiJtSMu0_1;
	wire w_dff_A_my9Nsj4F8_1;
	wire w_dff_A_h68msO2v9_1;
	wire w_dff_A_wzvmsC068_1;
	wire w_dff_A_R1aCiAet8_1;
	wire w_dff_A_FTobAgMp7_1;
	wire w_dff_A_UU9iPBcA4_0;
	wire w_dff_A_9A9lp9Eb4_0;
	wire w_dff_A_INzUODqZ4_0;
	wire w_dff_A_xXRZk73L2_0;
	wire w_dff_A_KuLxciOz2_0;
	wire w_dff_A_ezwpn8W24_0;
	wire w_dff_A_cWtTiz9r3_0;
	wire w_dff_A_Q53lHbmZ0_0;
	wire w_dff_A_02D4fnOb6_0;
	wire w_dff_A_shllhsGN3_1;
	wire w_dff_A_InB01ckg0_1;
	wire w_dff_A_pKrmJp5H2_1;
	wire w_dff_A_9GVTtQD67_1;
	wire w_dff_A_EFqaIDSk5_1;
	wire w_dff_A_n6e7PoKP8_1;
	wire w_dff_A_pj5cndwv9_1;
	wire w_dff_A_UtSll5fY6_1;
	wire w_dff_A_g03eD6ey0_1;
	wire w_dff_B_dlwkneye3_1;
	wire w_dff_B_KIrQzHVz5_0;
	wire w_dff_B_uMvaqNZj5_0;
	wire w_dff_B_lpsEsrVg7_0;
	wire w_dff_B_agLkgqch1_0;
	wire w_dff_B_0ZiPLVHK9_0;
	wire w_dff_B_aBUg2K088_0;
	wire w_dff_B_9hUKfTx27_0;
	wire w_dff_B_AgCrDA4K5_0;
	wire w_dff_B_dUEFt5038_0;
	wire w_dff_B_HLQ7PiTf1_0;
	wire w_dff_B_6GizWAwk6_0;
	wire w_dff_B_L6Cx6YAe2_0;
	wire w_dff_A_bOHcy3SC2_1;
	wire w_dff_A_YvldfqGX2_1;
	wire w_dff_A_1tR2bwiQ8_1;
	wire w_dff_A_roJ5mBDn7_1;
	wire w_dff_A_WUrOF5Nu4_1;
	wire w_dff_A_oTpOBk6E7_1;
	wire w_dff_A_3vOBsTQw1_1;
	wire w_dff_A_AvNJqJvz7_1;
	wire w_dff_A_1tKKaC8p3_1;
	wire w_dff_A_F039WYSQ4_1;
	wire w_dff_A_Bc55XUFv9_1;
	wire w_dff_A_3Fd7i2wB9_1;
	wire w_dff_A_Sj0lpnoe4_1;
	wire w_dff_A_FoUjy6Ta5_1;
	wire w_dff_A_ooD3Ukf66_1;
	wire w_dff_A_gn18gln43_1;
	wire w_dff_A_otzWUpkS7_1;
	wire w_dff_A_Ye0keKFV5_1;
	wire w_dff_B_YIE4AI0Q3_0;
	wire w_dff_B_mLhkwnQJ8_0;
	wire w_dff_B_ehZpJYeN2_0;
	wire w_dff_B_FuEYpuSB1_0;
	wire w_dff_B_Lvdg5TNC7_0;
	wire w_dff_A_V5b14Wph3_0;
	wire w_dff_A_aZ5BSb7c0_0;
	wire w_dff_A_RSja8HpL9_1;
	wire w_dff_A_N6nQcjI13_1;
	wire w_dff_A_nP6MPk1y1_1;
	wire w_dff_A_LOCLfv7S9_1;
	wire w_dff_A_KwU262fS1_1;
	wire w_dff_A_9apxVu2V1_1;
	wire w_dff_A_iZ1Nq6986_1;
	wire w_dff_A_aaz0C0hF6_1;
	wire w_dff_A_In3Yvowm5_2;
	wire w_dff_A_1i6Plmm84_2;
	wire w_dff_A_x6FcYThh9_2;
	wire w_dff_A_ruisOMEA3_2;
	wire w_dff_A_8Yt1i2r50_2;
	wire w_dff_A_046Llune2_2;
	wire w_dff_A_Uv46jueQ6_2;
	wire w_dff_A_f8RbYu1F1_2;
	wire w_dff_A_UOV4zIC17_2;
	wire w_dff_A_47HpDG880_2;
	wire w_dff_B_zMkHJ0nj7_3;
	wire w_dff_B_vcx3oYgK1_1;
	wire w_dff_B_CnIApL732_1;
	wire w_dff_B_9yUJyxsw7_1;
	wire w_dff_B_92diCjO80_1;
	wire w_dff_B_zhrKKLg55_1;
	wire w_dff_B_rbfxAyFi3_1;
	wire w_dff_B_DdYGjlKf0_1;
	wire w_dff_B_eBRHz32i5_1;
	wire w_dff_B_TMxMNK401_1;
	wire w_dff_B_rAKNhPEe8_1;
	wire w_dff_B_QxlXhkmt8_1;
	wire w_dff_B_bhIKsTNy3_1;
	wire w_dff_B_3kgt0fwD0_1;
	wire w_dff_B_uIgVnf2l3_1;
	wire w_dff_B_a38qD3AE2_1;
	wire w_dff_B_LS8NEahk2_1;
	wire w_dff_B_RY4ui54r9_1;
	wire w_dff_B_xRzrSoIB5_1;
	wire w_dff_B_OlOPpOTr1_1;
	wire w_dff_B_7OCCR3vq1_1;
	wire w_dff_B_QKD3aOcz1_1;
	wire w_dff_B_QdPGDnfW5_0;
	wire w_dff_A_NcwZOuFP5_1;
	wire w_dff_A_dT4pKEOP1_1;
	wire w_dff_A_QW8NP6Ae8_2;
	wire w_dff_A_jFvzm0Ak7_2;
	wire w_dff_A_eNJeqv691_2;
	wire w_dff_A_Js3VHItE4_2;
	wire w_dff_A_GKozbHjS6_0;
	wire w_dff_A_q2edVvNo5_0;
	wire w_dff_A_dG4J56FL1_0;
	wire w_dff_A_JviPyOI71_0;
	wire w_dff_A_YVufY6Yn4_0;
	wire w_dff_A_MWxTom3X1_0;
	wire w_dff_A_9qNzPFPT4_0;
	wire w_dff_A_Ig8XvwYb0_0;
	wire w_dff_A_koVGwb1J7_0;
	wire w_dff_A_LIhv0HB99_1;
	wire w_dff_B_Jm7YAUIf8_3;
	wire w_dff_B_VTZ8uKpI5_3;
	wire w_dff_B_q9HzVpiH3_3;
	wire w_dff_B_KqeXf7Wc5_3;
	wire w_dff_B_HHSiVRuC2_3;
	wire w_dff_B_9mmNTlrJ0_3;
	wire w_dff_B_q0Ustjpx0_3;
	wire w_dff_B_oL5kaV4W9_3;
	wire w_dff_B_9W7BhV6T4_3;
	wire w_dff_B_gKD6Sfvu3_3;
	wire w_dff_B_DcB3BtP64_3;
	wire w_dff_B_m5Gj2lRU7_3;
	wire w_dff_B_1w4VTA2g9_0;
	wire w_dff_B_5fvz4Qhb5_0;
	wire w_dff_B_z9sdbC247_0;
	wire w_dff_B_CL48g2ma9_0;
	wire w_dff_B_dkBEa0IK9_0;
	wire w_dff_B_HDnOkxuC9_0;
	wire w_dff_B_DTepdAYK3_0;
	wire w_dff_B_T2h4Zyv13_0;
	wire w_dff_B_vuZe0bKa8_0;
	wire w_dff_B_qtxyYpw43_1;
	wire w_dff_B_EDaRfIjO0_1;
	wire w_dff_B_IuNQyzo01_1;
	wire w_dff_B_ThDmAcZc5_1;
	wire w_dff_B_RI333wRp4_1;
	wire w_dff_B_5O1U2irJ4_1;
	wire w_dff_B_dPoGyPpH7_1;
	wire w_dff_B_oP1zgrp35_1;
	wire w_dff_B_Msf3FSz51_1;
	wire w_dff_B_BCtGabV65_1;
	wire w_dff_B_D2FAKTIT6_1;
	wire w_dff_B_tGstGLdi9_1;
	wire w_dff_B_4NzgPSVU1_1;
	wire w_dff_B_aosymfRH9_1;
	wire w_dff_B_niR2iSyj5_1;
	wire w_dff_B_yqWbuv4n6_1;
	wire w_dff_B_12eFf1aX0_1;
	wire w_dff_B_2noeHm9M2_1;
	wire w_dff_B_EFKFLGYk2_1;
	wire w_dff_B_spIMZWyK8_1;
	wire w_dff_B_mCRnWzHO9_1;
	wire w_dff_B_cTamk3c79_1;
	wire w_dff_B_XDGuFuiR0_1;
	wire w_dff_B_19NGwPN46_1;
	wire w_dff_B_y38gfn5x8_1;
	wire w_dff_B_oKUvMmsd4_1;
	wire w_dff_B_xrz6Q3Nn9_1;
	wire w_dff_B_mOsoktAu8_1;
	wire w_dff_B_v3aEujkO0_1;
	wire w_dff_A_UVuRWb7K0_1;
	wire w_dff_B_CUGOx4Xa8_2;
	wire w_dff_B_u7wJvy8b2_2;
	wire w_dff_B_tNTHa7YL0_2;
	wire w_dff_B_MMHg49Z23_2;
	wire w_dff_B_xhveRNNy9_2;
	wire w_dff_B_VlAAHc3T9_2;
	wire w_dff_B_8LlkZY8y6_2;
	wire w_dff_B_dDtBeSFw6_2;
	wire w_dff_B_f1hnKObp1_2;
	wire w_dff_A_DqTnrhIl5_0;
	wire w_dff_A_nZeOoi1Q7_0;
	wire w_dff_A_0QlFjbiQ7_0;
	wire w_dff_A_1fi3r4ZL8_0;
	wire w_dff_A_S0v5LtTG4_0;
	wire w_dff_A_AH4XdhIQ4_0;
	wire w_dff_A_OZxINHqO5_0;
	wire w_dff_A_8H6jWBfK8_0;
	wire w_dff_A_o5Z5aBps6_0;
	wire w_dff_A_xvKkIVhB3_0;
	wire w_dff_A_XHiH6VLY5_2;
	wire w_dff_A_h3xHLoam6_2;
	wire w_dff_A_0ZzOJ9s41_2;
	wire w_dff_A_OkZcfFI15_2;
	wire w_dff_A_D94QmB3M0_2;
	wire w_dff_A_S3M3fRAn7_2;
	wire w_dff_A_P17HqdxI6_2;
	wire w_dff_A_qEG7kw0c2_2;
	wire w_dff_A_VYUcKGTx5_2;
	wire w_dff_A_tWLi3I009_2;
	wire w_dff_A_BR6IopgH9_0;
	wire w_dff_B_OPiSdhep1_1;
	wire w_dff_B_mA4MlP5C4_1;
	wire w_dff_B_x2lpgnGr9_1;
	wire w_dff_B_6nB9UQd83_1;
	wire w_dff_B_c070VwAL9_1;
	wire w_dff_B_GOhcr1J55_1;
	wire w_dff_B_Nj6Fttg42_1;
	wire w_dff_B_tDiisvgf9_1;
	wire w_dff_B_8loXTjO36_1;
	wire w_dff_B_o6S3j0gd1_1;
	wire w_dff_B_28qe7Luv9_1;
	wire w_dff_B_0l3hpL6U6_1;
	wire w_dff_A_2xfzd5o59_1;
	wire w_dff_A_pjMlJL7w5_1;
	wire w_dff_A_x2JRJvFm8_1;
	wire w_dff_A_0BM63biI3_1;
	wire w_dff_A_Kd4YlRlz3_1;
	wire w_dff_A_J9u0xkXT3_1;
	wire w_dff_B_zfKJ7N7m9_3;
	wire w_dff_B_SoYIK06C6_3;
	wire w_dff_B_wlzgIIT85_3;
	wire w_dff_B_A0QiUiGi9_3;
	wire w_dff_B_tAww97vC7_3;
	wire w_dff_B_AyP8ITd23_3;
	wire w_dff_B_u8o26h9M9_3;
	wire w_dff_B_04yVh3Ik9_3;
	wire w_dff_A_anwux2PY4_1;
	wire w_dff_A_QCsBnuU61_1;
	wire w_dff_A_BgmEGnbB8_1;
	wire w_dff_A_78llugOu7_1;
	wire w_dff_A_red26bU52_1;
	wire w_dff_A_YkBjhwvG7_1;
	wire w_dff_A_a1dYiDs89_1;
	wire w_dff_A_GmaYrDzu7_1;
	wire w_dff_A_ZBaVSZNC1_1;
	wire w_dff_A_nDGu6vTd3_1;
	wire w_dff_A_6uI5kzyr7_1;
	wire w_dff_A_quB8R3mO5_1;
	wire w_dff_A_W8te3zfr7_1;
	wire w_dff_A_UUMNC2K21_1;
	wire w_dff_A_1rbhOwR07_1;
	wire w_dff_A_8iTJRlCD9_1;
	wire w_dff_A_8IYVivLB2_1;
	wire w_dff_A_bIp7JPaB2_1;
	wire w_dff_A_TS8rg5tl1_1;
	wire w_dff_A_lU1z5EkX9_1;
	wire w_dff_A_M72P0FaF0_2;
	wire w_dff_A_An7VvAPD4_2;
	wire w_dff_A_2D24J6EF4_2;
	wire w_dff_A_uOUQTLOU8_2;
	wire w_dff_A_KkbhJVix4_2;
	wire w_dff_A_S69iXiTB7_2;
	wire w_dff_A_VeWXXP224_2;
	wire w_dff_A_C5Xdz3Bg2_2;
	wire w_dff_A_Qc9qz0su8_1;
	wire w_dff_A_mTCIWOxs1_1;
	wire w_dff_A_DybErGmq4_1;
	wire w_dff_A_9r8CxF4s7_1;
	wire w_dff_A_BTDMx0wS6_0;
	wire w_dff_A_1f5IhjJr9_0;
	wire w_dff_A_fEVCnXKE6_0;
	wire w_dff_A_zsvxAFX32_0;
	wire w_dff_A_4DZ0DHiw3_0;
	wire w_dff_A_FdI0WKCU2_0;
	wire w_dff_A_pn8SS0211_0;
	wire w_dff_A_cBbE321R9_0;
	wire w_dff_A_l7iNudkR1_0;
	wire w_dff_A_IFC4esab3_0;
	wire w_dff_A_Jl2E8xC86_0;
	wire w_dff_A_pHvtnFbZ5_0;
	wire w_dff_A_fSh8t9Nd7_0;
	wire w_dff_A_LuLFkDYT4_0;
	wire w_dff_A_e3J1pnr79_2;
	wire w_dff_A_T1EEyyyr8_2;
	wire w_dff_A_8WUbxf3m4_2;
	wire w_dff_A_kKqLSNdp8_2;
	wire w_dff_A_31DXj4Dq1_1;
	wire w_dff_A_b6EtOz573_1;
	wire w_dff_A_sq5ThnlK4_1;
	wire w_dff_A_P8WvbM3b1_1;
	wire w_dff_A_NQy8YkrC9_1;
	wire w_dff_A_v2Ylb1H41_1;
	wire w_dff_A_vz9pDDQx5_1;
	wire w_dff_A_seVjTeaD7_1;
	wire w_dff_A_ocRD18GY1_1;
	wire w_dff_A_H5c3FY6G9_1;
	wire w_dff_A_M5arLt3Z5_1;
	wire w_dff_A_o61HqWLd7_1;
	wire w_dff_A_gaObyY8W5_1;
	wire w_dff_A_ld2lwYjb7_2;
	wire w_dff_A_YYBLDlml1_2;
	wire w_dff_A_tYxlxKKx9_2;
	wire w_dff_A_396RtzK68_2;
	wire w_dff_A_zrFuKfsF3_2;
	wire w_dff_A_VNL9OsKT4_2;
	wire w_dff_A_whrbb0aH2_2;
	wire w_dff_A_WSQG2nQG3_2;
	wire w_dff_A_rLOKQHf29_1;
	wire w_dff_A_WGCtSMdN0_1;
	wire w_dff_A_Mv4oLQNj8_1;
	wire w_dff_A_Ha0CWY2D6_1;
	wire w_dff_A_mhs3MIuJ4_1;
	wire w_dff_A_iU1DSUeC9_1;
	wire w_dff_A_483dyFML3_1;
	wire w_dff_B_ezOcNm4t7_2;
	wire w_dff_B_CSmh3Je67_2;
	wire w_dff_B_bYRmQvUm5_2;
	wire w_dff_B_h0oRvhMQ9_2;
	wire w_dff_A_qHBl9uKS2_1;
	wire w_dff_A_6ZSykUXi2_1;
	wire w_dff_A_WhvCCJdA1_1;
	wire w_dff_A_Sy6TL7yt6_1;
	wire w_dff_A_dyRndxjG7_1;
	wire w_dff_A_a6m6ldqn7_1;
	wire w_dff_A_QQdI9oVS9_0;
	wire w_dff_A_oNEUMF918_0;
	wire w_dff_A_UzPspmBP3_0;
	wire w_dff_A_Aq8Fg3Xa2_0;
	wire w_dff_A_e9JCRNt20_0;
	wire w_dff_A_XUFsdvAL9_0;
	wire w_dff_A_fYzr3aT48_0;
	wire w_dff_A_14aERbys4_0;
	wire w_dff_A_oqx76kKr5_2;
	wire w_dff_A_DQ1Z1PfJ2_2;
	wire w_dff_A_eayyPNSI1_2;
	wire w_dff_A_MQ4ZGfIg5_2;
	wire w_dff_A_cYE7uU0K1_0;
	wire w_dff_A_99289PEm0_0;
	wire w_dff_A_ZKjimvXj0_0;
	wire w_dff_A_uynJ8NEj6_0;
	wire w_dff_A_w1PX75V02_0;
	wire w_dff_A_rxyxfakq4_0;
	wire w_dff_B_sSOx9gG42_1;
	wire w_dff_B_6AzZ1H1p5_1;
	wire w_dff_B_eXhev64l3_1;
	wire w_dff_B_3ls2tTbH4_1;
	wire w_dff_B_mWfgVQSe2_1;
	wire w_dff_B_mTKOuLs62_1;
	wire w_dff_B_8HHs6aWx1_1;
	wire w_dff_B_LDgTm4kC5_1;
	wire w_dff_A_IeXxQwRr4_1;
	wire w_dff_A_oDNK9dM52_1;
	wire w_dff_A_nsmsM7Vo0_1;
	wire w_dff_A_tA9KHJR77_1;
	wire w_dff_A_Cyhj0a630_1;
	wire w_dff_A_Z3H8oW8K2_1;
	wire w_dff_A_xNiTWMvz0_1;
	wire w_dff_A_4LfsyQc45_1;
	wire w_dff_A_hgne0GEA0_0;
	wire w_dff_A_5iBE1NWo9_0;
	wire w_dff_A_xEFdfxMG1_0;
	wire w_dff_A_wZPeJeD78_1;
	wire w_dff_B_H5rML4Bq6_2;
	wire w_dff_B_XUM3G9YB3_2;
	wire w_dff_B_GcG3CTAF9_2;
	wire w_dff_B_dot5MtOb6_2;
	wire w_dff_A_XteMjSZF9_2;
	wire w_dff_A_PlGa8xbR6_2;
	wire w_dff_A_8MOAOxRw6_1;
	wire w_dff_A_fN5ygeVL3_1;
	wire w_dff_A_JgVbIWJL5_1;
	wire w_dff_A_JglYVlhD9_1;
	wire w_dff_A_4mivqqko8_1;
	wire w_dff_A_8giyetID5_1;
	wire w_dff_A_VoTRGCWD8_2;
	wire w_dff_A_0P9PFKav6_2;
	wire w_dff_A_xjpJJIxn4_2;
	wire w_dff_A_Rg0lTCs67_2;
	wire w_dff_A_cZXvq4qV6_2;
	wire w_dff_A_UhbXes9l8_2;
	wire w_dff_A_IgmkuNQI7_2;
	wire w_dff_A_OWSYhHc90_2;
	wire w_dff_A_kNBxYv8t5_0;
	wire w_dff_A_7mb8LDXE0_0;
	wire w_dff_A_30AxGuti7_0;
	wire w_dff_A_U9PRKNo19_0;
	wire w_dff_A_Zn4YRXEX2_0;
	wire w_dff_A_a2PKnu931_0;
	wire w_dff_A_NxHilTNr9_0;
	wire w_dff_B_zKATrJC61_1;
	wire w_dff_B_tFzcNDQB6_1;
	wire w_dff_B_6w5U4doO2_1;
	wire w_dff_B_bR7s2PsI3_1;
	wire w_dff_B_qbjWD4IA1_1;
	wire w_dff_B_93zzVgNs4_1;
	wire w_dff_B_bGqRnnrb1_1;
	wire w_dff_B_glwFMbs99_1;
	wire w_dff_B_CsfeRIgW3_1;
	wire w_dff_A_jPfP6liW8_2;
	wire w_dff_A_ZqMaRV2H7_2;
	wire w_dff_A_bGJ9bNfQ5_2;
	wire w_dff_A_5dOh7JfE7_2;
	wire w_dff_A_4vBgFoIK6_2;
	wire w_dff_A_Nl4mGuNV9_2;
	wire w_dff_A_JOw5s2Eq2_2;
	wire w_dff_A_xK92jhr56_2;
	wire w_dff_A_ipW7HfAD2_2;
	wire w_dff_B_i9r3DG767_0;
	wire w_dff_B_ciqDUL263_0;
	wire w_dff_B_MvlAQtoZ1_0;
	wire w_dff_B_m3ntz6Ex2_0;
	wire w_dff_B_XIBcCA2F5_0;
	wire w_dff_A_y3mouBv03_0;
	wire w_dff_A_mRobThW06_0;
	wire w_dff_A_YFJmtlCU5_0;
	wire w_dff_A_kXQhz9PI4_0;
	wire w_dff_A_ax5WHUV90_2;
	wire w_dff_A_Ko2aLk6Z1_2;
	wire w_dff_A_8WT2TR5T9_2;
	wire w_dff_A_E94MrDL39_2;
	wire w_dff_A_26RT9joY1_2;
	wire w_dff_A_8UkbWSPV4_0;
	wire w_dff_A_jOc1Jrnr3_0;
	wire w_dff_A_McXe5nSs8_0;
	wire w_dff_A_fVWiohJz8_0;
	wire w_dff_A_glkzfi5T9_0;
	wire w_dff_A_B83qHL3A6_0;
	wire w_dff_A_334p8xQ43_1;
	wire w_dff_A_WAu5TI1a0_1;
	wire w_dff_A_maI4D0hJ8_1;
	wire w_dff_A_oJxUuxOI2_1;
	wire w_dff_A_KQyuikLw0_1;
	wire w_dff_A_Nba9897K8_1;
	wire w_dff_A_ajnsYlh83_1;
	wire w_dff_A_VKL9Ekpq5_1;
	wire w_dff_A_ZQhRPJSx0_1;
	wire w_dff_A_xm8pmE884_1;
	wire w_dff_A_i40jUrVr9_1;
	wire w_dff_A_PWeDNBPz6_1;
	wire w_dff_A_8z0yNlva8_1;
	wire w_dff_A_B3n3HVkC2_2;
	wire w_dff_A_mMsfJ8203_2;
	wire w_dff_A_MjWJOxc81_2;
	wire w_dff_A_8bcqVPPU3_2;
	wire w_dff_A_nWOC50gK2_2;
	wire w_dff_A_X3CsfTMx8_2;
	wire w_dff_A_4jtYmsgS6_2;
	wire w_dff_A_9dMYSdZK5_2;
	wire w_dff_A_fapqLrpq9_2;
	wire w_dff_B_yW24bOoj0_1;
	wire w_dff_B_PXIpsMDO0_0;
	wire w_dff_B_1lNdlfgg1_0;
	wire w_dff_A_J3TufkYU2_0;
	wire w_dff_A_0oS0ytmE4_0;
	wire w_dff_A_5EeMiH4l1_0;
	wire w_dff_A_nQrjMWle6_0;
	wire w_dff_A_8mjQFyAe5_0;
	wire w_dff_A_wpFHotuG2_0;
	wire w_dff_A_cYDbRQww9_0;
	wire w_dff_A_bJRktpWx4_0;
	wire w_dff_A_l59Oc1ZP9_2;
	wire w_dff_A_ZnS2gN058_2;
	wire w_dff_A_McmTfj3E8_2;
	wire w_dff_A_ENDYzWRt5_2;
	wire w_dff_A_MQjCafdt2_2;
	wire w_dff_A_INQieLpD8_2;
	wire w_dff_A_jUMdPeOn3_2;
	wire w_dff_B_FuEt0jiw2_3;
	wire w_dff_B_a8ZUsWrQ6_0;
	wire w_dff_B_7CxqC9hv5_0;
	wire w_dff_B_X2daWbQK3_0;
	wire w_dff_B_KR80YAfB2_0;
	wire w_dff_B_oFcLweFb0_0;
	wire w_dff_B_NmhCqco59_0;
	wire w_dff_B_DeNkSHNd1_0;
	wire w_dff_B_AWGhTw5V5_0;
	wire w_dff_B_HeOxiRsb9_0;
	wire w_dff_B_X1cVvvvP1_0;
	wire w_dff_A_l3dyGvki7_1;
	wire w_dff_A_5gSeBWFA1_1;
	wire w_dff_A_fuPD4Wj19_1;
	wire w_dff_A_GCysLHp14_1;
	wire w_dff_A_56i1vK9h4_1;
	wire w_dff_A_WHbkWSbK3_1;
	wire w_dff_A_mHazPNP62_0;
	wire w_dff_A_jRhd2ij34_0;
	wire w_dff_A_TWAme1XX3_0;
	wire w_dff_A_gw1ZNbC50_0;
	wire w_dff_A_uByAPhOX3_0;
	wire w_dff_A_9bIjw1zb2_0;
	wire w_dff_A_9snBwZOH6_0;
	wire w_dff_A_SpZ9MXzk7_0;
	wire w_dff_A_tt70Y21S8_0;
	wire w_dff_A_Jf5HE9pc1_0;
	wire w_dff_A_jpgYigNZ1_0;
	wire w_dff_B_jIOpMdkz7_3;
	wire w_dff_B_wEZAlOlh8_3;
	wire w_dff_B_0WCv3TLZ4_3;
	wire w_dff_B_cmbRQYD50_3;
	wire w_dff_B_eAxTthJk6_3;
	wire w_dff_B_KsX5GkW32_3;
	wire w_dff_B_UooiwDuE6_3;
	wire w_dff_B_XaUMzDJl3_3;
	wire w_dff_B_CFuqkUPg8_3;
	wire w_dff_B_WmpA10mb3_0;
	wire w_dff_B_9q0iVMlk8_0;
	wire w_dff_B_znw2Letk3_0;
	wire w_dff_B_2Xn32A0M5_0;
	wire w_dff_B_FNdWpG6L9_0;
	wire w_dff_A_DbDIXG4L9_1;
	wire w_dff_B_GMGR8vUN1_2;
	wire w_dff_B_4hxEKc4C6_2;
	wire w_dff_B_GKshyJAs5_2;
	wire w_dff_B_QQafkqky1_2;
	wire w_dff_A_o7YaiDDE6_0;
	wire w_dff_B_za8Oaqir8_1;
	wire w_dff_B_Bhc3yBAC4_1;
	wire w_dff_A_iD8pjJNg7_0;
	wire w_dff_A_7uVQtD3w3_0;
	wire w_dff_B_dvlmMZNO4_2;
	wire w_dff_A_cwhJZiCj7_0;
	wire w_dff_A_wiFWWXhH9_0;
	wire w_dff_A_xFSlZ5xQ9_1;
	wire w_dff_A_BQoxbgMb8_0;
	wire w_dff_A_QEZn7ZAO1_0;
	wire w_dff_A_rP2600wd7_0;
	wire w_dff_A_HbOCAKGA8_0;
	wire w_dff_A_LBtVcvM64_2;
	wire w_dff_A_B2NdSyJ34_2;
	wire w_dff_A_11kSvh163_2;
	wire w_dff_A_hUzUa7W96_2;
	wire w_dff_A_eHHhQ4o84_1;
	wire w_dff_A_01w6qS8Y7_1;
	wire w_dff_A_Dk4KRjiK0_1;
	wire w_dff_A_GXOmb7M46_1;
	wire w_dff_A_DGKLle9m8_1;
	wire w_dff_A_1ljbPany4_1;
	wire w_dff_A_vFeJ34va1_1;
	wire w_dff_A_PUuizGx86_1;
	wire w_dff_A_kvs579UK1_2;
	wire w_dff_A_MAiR4MzR9_2;
	wire w_dff_A_QWcMVJQJ4_2;
	wire w_dff_A_Gf9ahnaf0_1;
	wire w_dff_A_sZpEfjxm0_0;
	wire w_dff_A_jwJe59Ba3_0;
	wire w_dff_A_c5k75pdr7_2;
	wire w_dff_A_u03eq0JM0_0;
	wire w_dff_A_mQhW8Len8_0;
	wire w_dff_A_1QWScWbE0_0;
	wire w_dff_A_IB2i9IMQ5_0;
	wire w_dff_A_MKDZ5sdi8_0;
	wire w_dff_A_ksBqX5wI0_0;
	wire w_dff_A_K1eXx5hX9_0;
	wire w_dff_A_OEXtbVry9_0;
	wire w_dff_A_c58gNbtU5_0;
	wire w_dff_A_N2CFVJcF4_1;
	wire w_dff_A_MWMuOC8p1_1;
	wire w_dff_A_ILxZoKM10_1;
	wire w_dff_B_AN5zqfCe9_2;
	wire w_dff_B_YizhvhEt1_2;
	wire w_dff_B_11dJR2233_2;
	wire w_dff_B_P7cmgdDp0_2;
	wire w_dff_A_vzH8a5IH7_0;
	wire w_dff_A_2XlABTEg4_0;
	wire w_dff_A_dwxSv1RD3_0;
	wire w_dff_A_ia9jZOxB4_0;
	wire w_dff_A_BLBEEKtT3_0;
	wire w_dff_A_EWvd61zV2_0;
	wire w_dff_A_4VxHcluu1_0;
	wire w_dff_A_casShWez8_0;
	wire w_dff_A_pJ1fMVAp6_0;
	wire w_dff_A_zmkTIIpv0_2;
	wire w_dff_A_rfF6o2O05_2;
	wire w_dff_A_2c7NHnrQ1_2;
	wire w_dff_A_xQNw0OnY0_2;
	wire w_dff_A_gPeBrji92_2;
	wire w_dff_A_z8eXRr5A9_2;
	wire w_dff_A_2HEyaCAt9_2;
	wire w_dff_A_ZwDqmSz09_2;
	wire w_dff_A_8DAk1jc00_2;
	wire w_dff_A_u44msslo6_0;
	wire w_dff_A_AyCz4Zwr6_0;
	wire w_dff_A_IAfzXxZD6_0;
	wire w_dff_A_yoTihmYo6_0;
	wire w_dff_A_OX7Xvnjl4_0;
	wire w_dff_A_VzplXodn2_0;
	wire w_dff_B_fzp31Fxl5_0;
	wire w_dff_A_rMNiHgEZ7_1;
	wire w_dff_A_T8HV43pC6_1;
	wire w_dff_A_uDr2tGyW1_1;
	wire w_dff_A_KOJIDJab2_1;
	wire w_dff_A_OfANTNyH8_1;
	wire w_dff_A_NZCi6Slt0_1;
	wire w_dff_A_8SHFtRHc4_1;
	wire w_dff_A_LtKNNQCe6_1;
	wire w_dff_A_e94DEHcZ9_2;
	wire w_dff_A_BGG8C18W6_1;
	wire w_dff_A_2CGoF0uM9_1;
	wire w_dff_A_cgeT17iR4_1;
	wire w_dff_A_UMPOKdDL3_1;
	wire w_dff_A_0qB5OCiB0_1;
	wire w_dff_A_YZFSoUtL7_1;
	wire w_dff_A_o0FLiivG4_0;
	wire w_dff_A_ZQT4YDvQ5_1;
	wire w_dff_A_nKJDjkL34_1;
	wire w_dff_B_JujjifIW0_3;
	wire w_dff_B_xxKpXUDp7_3;
	wire w_dff_A_b32WYCJk1_1;
	wire w_dff_A_y9MYhpIM0_1;
	wire w_dff_A_cK461G5Q8_1;
	wire w_dff_A_YFSbislH0_1;
	wire w_dff_A_SXcLFPzC3_1;
	wire w_dff_A_2PfAN4md2_1;
	wire w_dff_A_Wf8QQ8nr5_1;
	wire w_dff_A_t5wWn38Z1_1;
	wire w_dff_A_cLI7CXP81_1;
	wire w_dff_A_abAoN42z4_2;
	wire w_dff_A_CxrZOvs51_2;
	wire w_dff_A_Sl3VTDFt4_2;
	wire w_dff_A_Ow6Vz5Bk2_2;
	wire w_dff_A_HnFtxZya6_2;
	wire w_dff_A_F5mEcLzK3_2;
	wire w_dff_A_6zpQ6MoK7_2;
	wire w_dff_A_BLh70akQ9_2;
	wire w_dff_A_GgjU2x5B7_2;
	wire w_dff_A_4Wk26QqG3_2;
	wire w_dff_A_SoV7oXqQ8_2;
	wire w_dff_A_GIQFJFMG3_2;
	wire w_dff_A_hNzUy3C26_0;
	wire w_dff_A_HYf2Kd3O9_0;
	wire w_dff_A_UdpQExC23_0;
	wire w_dff_A_9gIHhL6b2_0;
	wire w_dff_A_5xrj0h4v1_0;
	wire w_dff_A_ydi3PxeD3_0;
	wire w_dff_A_4YhMBPaD5_0;
	wire w_dff_A_CVIhwn9k7_0;
	wire w_dff_A_VtF0Vlih0_0;
	wire w_dff_A_COl9Ozh81_0;
	wire w_dff_A_yBQKFVk97_0;
	wire w_dff_A_jQWl3CYa9_0;
	wire w_dff_A_Bo2R4vhC6_0;
	wire w_dff_A_m23qoWUg7_0;
	wire w_dff_A_YHBTuddm7_0;
	wire w_dff_A_PWXCsM2V4_0;
	wire w_dff_A_Y795aTw98_0;
	wire w_dff_A_xtXY9Qgj6_0;
	wire w_dff_A_jyPsdBQa2_0;
	wire w_dff_A_IXkJs7qp0_0;
	wire w_dff_A_nAJ0ve2e5_0;
	wire w_dff_A_MWRKUUOo2_0;
	wire w_dff_A_PTVaSj3j8_0;
	wire w_dff_A_rryMQYmW9_0;
	wire w_dff_A_R3S5W4FU9_0;
	wire w_dff_A_fbbwZBC94_2;
	wire w_dff_A_jSaQN0AA1_0;
	wire w_dff_A_ve7dmZ7D2_0;
	wire w_dff_A_1hRV36Pn6_0;
	wire w_dff_A_PBm86oNA2_0;
	wire w_dff_A_2KRlKMh88_0;
	wire w_dff_A_uRl38xeF7_0;
	wire w_dff_A_6pObr9Ln7_0;
	wire w_dff_A_uMrqc91R6_0;
	wire w_dff_A_va78vqte5_0;
	wire w_dff_A_tPACDJAS1_0;
	wire w_dff_A_yoYm7YRD7_0;
	wire w_dff_A_IYLSHnMS1_0;
	wire w_dff_A_UdbzN5yS0_0;
	wire w_dff_A_F9RWbxcd9_0;
	wire w_dff_A_ZTbwGDAX5_0;
	wire w_dff_A_m8haK0v40_0;
	wire w_dff_A_zSKpGYeN9_0;
	wire w_dff_A_4eQtuMk60_0;
	wire w_dff_A_NIYwisdb9_0;
	wire w_dff_A_Ijs7conF8_0;
	wire w_dff_A_uwTdvjEV1_0;
	wire w_dff_A_x0aaxlvi6_0;
	wire w_dff_A_iuAo3Qz44_0;
	wire w_dff_A_XotlsMEW3_0;
	wire w_dff_A_QTpWsiND3_0;
	wire w_dff_A_B6Z4XMwz7_2;
	wire w_dff_A_wRmIRAMI0_0;
	wire w_dff_A_S3m42r8M6_0;
	wire w_dff_A_LZUfgs5F0_0;
	wire w_dff_A_yEjoW1Qk3_0;
	wire w_dff_A_OcKqlTmC9_0;
	wire w_dff_A_yW90sm0m6_0;
	wire w_dff_A_dP2rJuKa1_0;
	wire w_dff_A_sZzN5gI33_0;
	wire w_dff_A_Jo3KCtou0_0;
	wire w_dff_A_kgFX5hg30_0;
	wire w_dff_A_VUBk74w62_0;
	wire w_dff_A_eSqNkEQo7_0;
	wire w_dff_A_cYzay5hk4_0;
	wire w_dff_A_iO0Gkb0I3_0;
	wire w_dff_A_HuXGHdDg8_0;
	wire w_dff_A_NKwVIKgT5_0;
	wire w_dff_A_JDDW7R9A6_0;
	wire w_dff_A_ZANfmTyv5_0;
	wire w_dff_A_asSSJUnh0_0;
	wire w_dff_A_9Co9E0rq3_0;
	wire w_dff_A_4quQ58v91_0;
	wire w_dff_A_kJqkduKb7_0;
	wire w_dff_A_VpMAyCip6_0;
	wire w_dff_A_xi3aKtf99_0;
	wire w_dff_A_gSloLsBp0_0;
	wire w_dff_A_SfdgPlOZ3_2;
	wire w_dff_A_vBWDEs5c1_0;
	wire w_dff_A_KuiwLew39_0;
	wire w_dff_A_nyLFFR8d9_0;
	wire w_dff_A_k7ZNQdRN9_0;
	wire w_dff_A_hcdzESoJ0_0;
	wire w_dff_A_kggYYSB87_0;
	wire w_dff_A_HjgcAcXl8_0;
	wire w_dff_A_CUB2NcDZ0_0;
	wire w_dff_A_Ba809Wac7_0;
	wire w_dff_A_JxlBc8Sd7_0;
	wire w_dff_A_02TkcAql6_0;
	wire w_dff_A_7xwQTvFu0_0;
	wire w_dff_A_f3kPU7WM8_0;
	wire w_dff_A_NJtBqYph0_0;
	wire w_dff_A_KPZQvkGt3_0;
	wire w_dff_A_Qe8WeW3m9_0;
	wire w_dff_A_MeuYDjcY3_0;
	wire w_dff_A_6973Muxp3_0;
	wire w_dff_A_aVP18PBt1_0;
	wire w_dff_A_uBj7VEeD6_0;
	wire w_dff_A_A4ak95H22_0;
	wire w_dff_A_WGXjJkGa5_0;
	wire w_dff_A_HAdk9kq35_0;
	wire w_dff_A_lXsy4q6L0_0;
	wire w_dff_A_ymRDstN55_0;
	wire w_dff_A_XUrvf1oR3_0;
	wire w_dff_A_bkmCrY7r7_2;
	wire w_dff_A_hQPliWiR0_0;
	wire w_dff_A_WCCPC7mf8_0;
	wire w_dff_A_J46msa4H9_0;
	wire w_dff_A_JK3WZePZ1_0;
	wire w_dff_A_wVqMcpz18_0;
	wire w_dff_A_7dLJFCyl3_0;
	wire w_dff_A_Dj3KXIK08_0;
	wire w_dff_A_9IAYhGbG7_0;
	wire w_dff_A_ougHFFr31_0;
	wire w_dff_A_qTeYnMfb1_0;
	wire w_dff_A_aW7shEvn7_0;
	wire w_dff_A_VIQuqmzX1_0;
	wire w_dff_A_yvNuwgYP6_0;
	wire w_dff_A_bR1BvdoU1_0;
	wire w_dff_A_ZKtCFEUh6_0;
	wire w_dff_A_DBcX3uwA7_0;
	wire w_dff_A_tj90LY1N2_0;
	wire w_dff_A_HACOFh6N6_0;
	wire w_dff_A_Am9WZO1c8_0;
	wire w_dff_A_qKtCd8Ts5_0;
	wire w_dff_A_Y74HGvs07_0;
	wire w_dff_A_1RT2dsJt2_0;
	wire w_dff_A_hBxrswGj8_0;
	wire w_dff_A_9onCqjcb8_0;
	wire w_dff_A_1Qm6wZAT2_2;
	wire w_dff_A_fyU4uy8r8_0;
	wire w_dff_A_REviNEA89_0;
	wire w_dff_A_biMb3fA81_0;
	wire w_dff_A_e64spRBK1_0;
	wire w_dff_A_CuqN56HP9_0;
	wire w_dff_A_zUeRAHfu0_0;
	wire w_dff_A_QDRF8MyT5_0;
	wire w_dff_A_NwIKnT2t9_0;
	wire w_dff_A_OkbSKNTw9_0;
	wire w_dff_A_GIzN6gNR8_0;
	wire w_dff_A_iceEIwMC3_0;
	wire w_dff_A_JCj4zyd77_0;
	wire w_dff_A_TfrNrFBp0_0;
	wire w_dff_A_VjMYD0g27_0;
	wire w_dff_A_UXsqAlfR8_0;
	wire w_dff_A_Gig8wDLv7_0;
	wire w_dff_A_D8oX5u4W2_0;
	wire w_dff_A_1iPypINM9_0;
	wire w_dff_A_TGbE6zxt8_0;
	wire w_dff_A_9IgYhVHZ6_0;
	wire w_dff_A_4YkMIkOM9_0;
	wire w_dff_A_sEpUOhkm8_0;
	wire w_dff_A_9ZHzostQ4_2;
	wire w_dff_A_acBW3aA58_0;
	wire w_dff_A_wfNRpohp9_0;
	wire w_dff_A_KZUbdoto3_0;
	wire w_dff_A_wAsaG9s20_0;
	wire w_dff_A_beErWbUR7_0;
	wire w_dff_A_8ZaBReQ67_0;
	wire w_dff_A_0OxHTqHH2_0;
	wire w_dff_A_1Sm6ge9R7_0;
	wire w_dff_A_oFa3N5p55_0;
	wire w_dff_A_QphaYer82_0;
	wire w_dff_A_cGVdMqKs0_0;
	wire w_dff_A_2fAN20vg7_0;
	wire w_dff_A_7Up1IEB24_0;
	wire w_dff_A_Ga8YSLXj1_0;
	wire w_dff_A_2EC8B5CU6_0;
	wire w_dff_A_MviX3CIa3_0;
	wire w_dff_A_31fFjjjP5_0;
	wire w_dff_A_7JhZFazM7_0;
	wire w_dff_A_5ND675611_0;
	wire w_dff_A_VfkJ2ffF6_0;
	wire w_dff_A_7ZywvmuN4_0;
	wire w_dff_A_7ugerTbt5_0;
	wire w_dff_A_NbqsnwDp3_0;
	wire w_dff_A_zll0YeUD6_0;
	wire w_dff_A_SkEow26f5_2;
	wire w_dff_A_WTGvmPFJ6_0;
	wire w_dff_A_580p66MJ0_0;
	wire w_dff_A_HAe6mKe86_0;
	wire w_dff_A_8lztFpFF3_0;
	wire w_dff_A_whH2awry4_0;
	wire w_dff_A_pW0Tunmb3_0;
	wire w_dff_A_8FDJjDhL1_0;
	wire w_dff_A_1xpN1gvE0_0;
	wire w_dff_A_tjCnTYPO9_0;
	wire w_dff_A_q1RjnNjV2_0;
	wire w_dff_A_lGHzpP2K9_0;
	wire w_dff_A_8evsPL0x0_0;
	wire w_dff_A_mUrv24N39_0;
	wire w_dff_A_YUvPkBC11_0;
	wire w_dff_A_iy99ALRm4_0;
	wire w_dff_A_bquknk935_0;
	wire w_dff_A_ClWfCns00_0;
	wire w_dff_A_h6j1DMIR8_0;
	wire w_dff_A_Rd2m1PqP1_0;
	wire w_dff_A_W7Ta6o5n7_0;
	wire w_dff_A_QN1uYlrj0_0;
	wire w_dff_A_oK1GntID5_0;
	wire w_dff_A_2lJ3JvEA3_0;
	wire w_dff_A_4uussoog7_0;
	wire w_dff_A_I6hNTVIN6_2;
	wire w_dff_A_UWL0sjX75_0;
	wire w_dff_A_i3BAsUMv5_0;
	wire w_dff_A_IaZxsaC34_0;
	wire w_dff_A_LtjsvLjX6_0;
	wire w_dff_A_JP1jIevG1_0;
	wire w_dff_A_Nr1C3yTv3_0;
	wire w_dff_A_3f7IvP7f5_0;
	wire w_dff_A_U8xSx5Ew2_0;
	wire w_dff_A_FmgqqfDT6_0;
	wire w_dff_A_4T3mnRGm0_0;
	wire w_dff_A_rlDa8G7I0_0;
	wire w_dff_A_TrBUl0CH8_0;
	wire w_dff_A_cOteOzgK6_0;
	wire w_dff_A_agQG2JiC2_0;
	wire w_dff_A_Umkynk5O8_0;
	wire w_dff_A_gdtMSq9E0_0;
	wire w_dff_A_HEEfDagU7_0;
	wire w_dff_A_6iK7sCAt0_0;
	wire w_dff_A_0E8ukRdX8_0;
	wire w_dff_A_EEPdjaFa1_0;
	wire w_dff_A_3tBpD3Ub2_0;
	wire w_dff_A_HOKKmCWx5_0;
	wire w_dff_A_Wa24sCIH3_0;
	wire w_dff_A_F1ipmiP76_0;
	wire w_dff_A_T2sNp57Q1_2;
	wire w_dff_A_AViv2ydS4_0;
	wire w_dff_A_mOtVQSuK3_0;
	wire w_dff_A_QmUATijc3_0;
	wire w_dff_A_w06XInNC2_0;
	wire w_dff_A_kruvq9g07_0;
	wire w_dff_A_wXbxsZVw8_0;
	wire w_dff_A_lM2WTgx74_0;
	wire w_dff_A_lYK3QlDD8_0;
	wire w_dff_A_U8aXldGM7_0;
	wire w_dff_A_H09nZfvu1_0;
	wire w_dff_A_phD9twfj6_0;
	wire w_dff_A_yCaodL0W3_0;
	wire w_dff_A_B3C2OSum0_0;
	wire w_dff_A_eMjIMQTM2_0;
	wire w_dff_A_kQhVdl753_0;
	wire w_dff_A_XIIIajo33_0;
	wire w_dff_A_bfTbC6NH3_0;
	wire w_dff_A_Aj1U1yTI8_0;
	wire w_dff_A_ngAkVC322_0;
	wire w_dff_A_PBgaHB1v6_0;
	wire w_dff_A_rGjUSLxV1_0;
	wire w_dff_A_0bR3ugqN0_0;
	wire w_dff_A_em60hgpk7_0;
	wire w_dff_A_BLJyWh090_0;
	wire w_dff_A_Fusx2Vwr8_0;
	wire w_dff_A_kFfvaOFK5_2;
	wire w_dff_A_OzMqJS1k6_0;
	wire w_dff_A_RxOJXN9A2_0;
	wire w_dff_A_58wZptTP9_0;
	wire w_dff_A_7imoNw4O6_0;
	wire w_dff_A_NmI395vY1_0;
	wire w_dff_A_LaVAz5DS5_0;
	wire w_dff_A_wAGIcrs39_0;
	wire w_dff_A_Qtw4eZ4n9_0;
	wire w_dff_A_GUNwJM1d3_0;
	wire w_dff_A_tGLuDtpy5_0;
	wire w_dff_A_0O3iMY6p0_0;
	wire w_dff_A_AXd9OF3W7_0;
	wire w_dff_A_WYpEkHrg4_0;
	wire w_dff_A_rCjwCbZR5_0;
	wire w_dff_A_P2ceZMPk4_0;
	wire w_dff_A_Q4tJVLvs2_0;
	wire w_dff_A_gnCI5dYD0_0;
	wire w_dff_A_E1flEDp32_0;
	wire w_dff_A_4wahLqaV1_0;
	wire w_dff_A_uEZAeyGF3_0;
	wire w_dff_A_QtUIoXPa8_0;
	wire w_dff_A_gHXN3bwJ7_0;
	wire w_dff_A_lEJ8kvaV2_1;
	wire w_dff_A_QmD3fafN3_0;
	wire w_dff_A_FJLkcpR43_0;
	wire w_dff_A_PWAa442S8_0;
	wire w_dff_A_74lxLGlB1_0;
	wire w_dff_A_4Tzv2tcl6_0;
	wire w_dff_A_ayLFv6v43_0;
	wire w_dff_A_PS2K9Hhq2_0;
	wire w_dff_A_rZw7cAaJ6_0;
	wire w_dff_A_qXSm7VNz4_0;
	wire w_dff_A_btzlUGQO0_0;
	wire w_dff_A_2fwbiHCh5_0;
	wire w_dff_A_bpYxWGFP0_0;
	wire w_dff_A_wQLMnZ0d6_0;
	wire w_dff_A_J2d3jfCx5_0;
	wire w_dff_A_tgM0fDix1_0;
	wire w_dff_A_AKEwKhuf3_0;
	wire w_dff_A_vl5dJyz83_0;
	wire w_dff_A_ZOFqoI5P0_0;
	wire w_dff_A_iWxVOVxW1_0;
	wire w_dff_A_ZvXdbyex2_0;
	wire w_dff_A_ZUObxu8A1_0;
	wire w_dff_A_mt7vBhuX3_0;
	wire w_dff_A_GVyWvK378_0;
	wire w_dff_A_yDVVGrpt7_0;
	wire w_dff_A_mpN0foaq8_0;
	wire w_dff_A_oCZBiHiG0_2;
	wire w_dff_A_2JERXUrB0_0;
	wire w_dff_A_6NW6omcr6_0;
	wire w_dff_A_YHxMdtWv8_0;
	wire w_dff_A_ic6tqCU62_0;
	wire w_dff_A_kat0AlJe6_0;
	wire w_dff_A_wnUuWrXU7_0;
	wire w_dff_A_KaCbYYrN1_0;
	wire w_dff_A_YPj9QUrI7_0;
	wire w_dff_A_QaQMfFeL1_0;
	wire w_dff_A_zJRYce1J2_0;
	wire w_dff_A_dSx2ufSZ2_0;
	wire w_dff_A_CpT9y3rb1_0;
	wire w_dff_A_Hiz2JChW3_0;
	wire w_dff_A_VjdYfxEZ5_0;
	wire w_dff_A_1qbnn19P4_0;
	wire w_dff_A_oMvdRlKt5_0;
	wire w_dff_A_1wbfVwSH9_0;
	wire w_dff_A_nL2ZaUsE8_0;
	wire w_dff_A_bioNuumO7_0;
	wire w_dff_A_bJw0UQ8m2_0;
	wire w_dff_A_JFUxqJ0Y7_0;
	wire w_dff_A_pNAFHhct9_0;
	wire w_dff_A_WQugsFuT0_2;
	wire w_dff_A_XTcE3euz8_0;
	wire w_dff_A_waGQQAOv1_0;
	wire w_dff_A_rv02eS0u7_0;
	wire w_dff_A_F259Dxet0_0;
	wire w_dff_A_h86j0hNt3_0;
	wire w_dff_A_J9igMIAL8_0;
	wire w_dff_A_QIz5LeYD6_0;
	wire w_dff_A_u8g82CIV7_0;
	wire w_dff_A_dAaxuK4I1_0;
	wire w_dff_A_NijWWpc73_0;
	wire w_dff_A_xXt4BVmR5_0;
	wire w_dff_A_hTgsqFPi3_0;
	wire w_dff_A_rjO19pxN6_0;
	wire w_dff_A_Fuo5gRsU8_0;
	wire w_dff_A_NvxyFkI47_0;
	wire w_dff_A_D7AgZQwK1_0;
	wire w_dff_A_QmAyNK9p3_0;
	wire w_dff_A_eiV3VIfR3_0;
	wire w_dff_A_p4yhxYh72_0;
	wire w_dff_A_NiUnCLL54_0;
	wire w_dff_A_Is1bllA11_0;
	wire w_dff_A_OEwO9Xu70_0;
	wire w_dff_A_62IaO45P5_2;
	wire w_dff_A_ZxS6W6qB8_0;
	wire w_dff_A_ug4qJM6l3_0;
	wire w_dff_A_C7efjcvX5_0;
	wire w_dff_A_u88nR0RM1_0;
	wire w_dff_A_KCv2dHGN0_0;
	wire w_dff_A_UMGNC58v9_0;
	wire w_dff_A_72BmfYVd6_0;
	wire w_dff_A_BQWGDUTw9_0;
	wire w_dff_A_EIBhi0YZ6_0;
	wire w_dff_A_5fbcAUl66_0;
	wire w_dff_A_ddkWoOpC0_0;
	wire w_dff_A_vX8ioDB01_0;
	wire w_dff_A_ka0TKRWq7_0;
	wire w_dff_A_qOdIGPmS4_0;
	wire w_dff_A_Zt725Dud5_0;
	wire w_dff_A_ZAMa8JRO3_0;
	wire w_dff_A_7ZsLcK9Y2_0;
	wire w_dff_A_ICYRftez4_0;
	wire w_dff_A_ofPhop2v2_0;
	wire w_dff_A_95AUTe252_0;
	wire w_dff_A_tCMNmrpR3_0;
	wire w_dff_A_yk9RaUOh7_0;
	wire w_dff_A_0o7VBkEv9_0;
	wire w_dff_A_P26aDpeN7_0;
	wire w_dff_A_VOorZblU0_0;
	wire w_dff_A_OhvIt33J6_2;
	wire w_dff_A_AUMM5Vz60_0;
	wire w_dff_A_MuCpLdEp1_0;
	wire w_dff_A_aRuHzX8a2_0;
	wire w_dff_A_NbCZVsyv7_0;
	wire w_dff_A_XTyI7J1O0_0;
	wire w_dff_A_yVaoSb9n5_0;
	wire w_dff_A_1k7aEVIY2_0;
	wire w_dff_A_LC6fSsxW5_0;
	wire w_dff_A_OVKzfKEI9_0;
	wire w_dff_A_wFtQ1NoB3_0;
	wire w_dff_A_tUzFcp0y5_0;
	wire w_dff_A_8eD8pS870_0;
	wire w_dff_A_hIljqn2Y2_0;
	wire w_dff_A_BK98MWIm0_0;
	wire w_dff_A_0xWxjbdh4_0;
	wire w_dff_A_0Zl1UtQM3_0;
	wire w_dff_A_tvmBxap54_0;
	wire w_dff_A_S3mzQaB14_0;
	wire w_dff_A_g88LvIVh0_0;
	wire w_dff_A_tl4Y0fmj2_0;
	wire w_dff_A_mjJ7ijoY0_0;
	wire w_dff_A_hSRmfOOu2_0;
	wire w_dff_A_oSEqh7DY6_0;
	wire w_dff_A_ijyXFBE84_2;
	wire w_dff_A_KuZ0yOuE6_0;
	wire w_dff_A_aAAvfzJ80_0;
	wire w_dff_A_Pu6n5JId9_0;
	wire w_dff_A_AvgbYcVt5_0;
	wire w_dff_A_ZmfYtXFB7_0;
	wire w_dff_A_Pg91RuED2_0;
	wire w_dff_A_rMGvYZY82_0;
	wire w_dff_A_tmntGwPz8_0;
	wire w_dff_A_CsS5h76y1_0;
	wire w_dff_A_mma5k4kX1_0;
	wire w_dff_A_BnO6ZzXq4_0;
	wire w_dff_A_mgCwxtpr3_0;
	wire w_dff_A_rfpx7WkN7_0;
	wire w_dff_A_RW1mjh6D3_0;
	wire w_dff_A_qaVO5FQs0_0;
	wire w_dff_A_crGx4l1H3_0;
	wire w_dff_A_vUx8xaFD1_0;
	wire w_dff_A_gciaVF359_0;
	wire w_dff_A_HYVAJKsk6_0;
	wire w_dff_A_UJnDelxg1_0;
	wire w_dff_A_YKWzR1UF5_0;
	wire w_dff_A_FWpgesYV0_0;
	wire w_dff_A_LmQboStI7_0;
	wire w_dff_A_nh87JbUt4_2;
	wire w_dff_A_3HWwNyCh1_0;
	wire w_dff_A_8ewzlnrw4_0;
	wire w_dff_A_szbM88Hs5_0;
	wire w_dff_A_hh9atL544_0;
	wire w_dff_A_Iw8W4qYS5_0;
	wire w_dff_A_sk0xNoWH7_0;
	wire w_dff_A_0FE8NSYg9_0;
	wire w_dff_A_5KektUN41_0;
	wire w_dff_A_DiP8ilzB0_0;
	wire w_dff_A_EOaVoLqy9_0;
	wire w_dff_A_VM7UAmMV3_0;
	wire w_dff_A_77IM1GqG4_0;
	wire w_dff_A_83XL4cAE0_2;
	wire w_dff_A_bpe8gIj91_0;
	wire w_dff_A_We2goBjS7_0;
	wire w_dff_A_JsLojnvW6_0;
	wire w_dff_A_GFVDQyAf8_0;
	wire w_dff_A_SOw645RN6_0;
	wire w_dff_A_rjOJlnYr7_0;
	wire w_dff_A_SNdymnnu5_0;
	wire w_dff_A_QaPWEmmy9_2;
	wire w_dff_A_ValFc8q85_0;
	wire w_dff_A_kUTamCJQ5_0;
	wire w_dff_A_yxO3DTUZ5_0;
	wire w_dff_A_ZzVYyaWT0_0;
	wire w_dff_A_A8IE8g3U1_0;
	wire w_dff_A_bXBWkxwt4_0;
	wire w_dff_A_VXM6wOLH7_0;
	wire w_dff_A_cyP2e2Cq8_0;
	wire w_dff_A_3qCCnxzi9_0;
	wire w_dff_A_KtnSHZjt1_2;
	wire w_dff_A_eiJRXx2o6_0;
	wire w_dff_A_TmawjQ0z0_0;
	wire w_dff_A_wfClqdcP7_0;
	wire w_dff_A_bLZCEdsN7_0;
	wire w_dff_A_KUE60uwm4_0;
	wire w_dff_A_e5xMsPhh0_0;
	wire w_dff_A_ZksiIyXT7_0;
	wire w_dff_A_qif6j39L7_0;
	wire w_dff_A_470sFp8E4_0;
	wire w_dff_A_a42W2vVw9_0;
	wire w_dff_A_fbA61J2w0_0;
	wire w_dff_A_lxhkViEa1_2;
	wire w_dff_A_c67N0HXi9_0;
	wire w_dff_A_L5KrTId14_2;
	wire w_dff_A_x0qGp2kE0_0;
	wire w_dff_A_stx7Dq2G1_0;
	wire w_dff_A_EkudcTpl9_0;
	wire w_dff_A_1zwzZJkW2_0;
	wire w_dff_A_wWIeNAhW9_2;
	wire w_dff_A_rijtXIGe1_0;
	wire w_dff_A_vX37Lua63_2;
	wire w_dff_A_Txp4bkph8_0;
	wire w_dff_A_3hVaVjDW6_0;
	wire w_dff_A_vla4J1i82_0;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(w_dff_A_GIQFJFMG3_2),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(w_dff_A_fbbwZBC94_2),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(w_dff_A_SfdgPlOZ3_2),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_n92_0[1]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_G17gat_2[2]),.dout(w_dff_A_bkmCrY7r7_2),.clk(gclk));
	jnot g009(.din(w_G17gat_2[1]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G13gat_0[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G1gat_1[0]),.dout(n97),.clk(gclk));
	jnot g012(.din(w_G26gat_0[1]),.dout(n98),.clk(gclk));
	jor g013(.dina(n98),.dinb(w_n97_0[1]),.dout(n99),.clk(gclk));
	jor g014(.dina(w_n99_0[1]),.dinb(w_dff_B_owR0xsDs9_1),.dout(n100),.clk(gclk));
	jor g015(.dina(n100),.dinb(w_n95_0[2]),.dout(n101),.clk(gclk));
	jor g016(.dina(w_n101_0[1]),.dinb(w_G390gat_0[1]),.dout(w_dff_A_1Qm6wZAT2_2),.clk(gclk));
	jnot g017(.din(w_G80gat_0[1]),.dout(n103),.clk(gclk));
	jand g018(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n104),.clk(gclk));
	jnot g019(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jor g020(.dina(n105),.dinb(w_n103_0[1]),.dout(w_dff_A_9ZHzostQ4_2),.clk(gclk));
	jnot g021(.din(w_G36gat_0[0]),.dout(n107),.clk(gclk));
	jnot g022(.din(w_G59gat_1[0]),.dout(n108),.clk(gclk));
	jor g023(.dina(w_n108_0[1]),.dinb(n107),.dout(n109),.clk(gclk));
	jor g024(.dina(w_n109_0[1]),.dinb(w_n103_0[0]),.dout(w_dff_A_SkEow26f5_2),.clk(gclk));
	jnot g025(.din(w_G42gat_1[2]),.dout(n111),.clk(gclk));
	jor g026(.dina(w_n109_0[0]),.dinb(w_n111_0[1]),.dout(w_dff_A_I6hNTVIN6_2),.clk(gclk));
	jor g027(.dina(G88gat),.dinb(G87gat),.dout(n113),.clk(gclk));
	jand g028(.dina(w_n113_0[1]),.dinb(w_dff_B_aBFOmxD08_1),.dout(w_dff_A_T2sNp57Q1_2),.clk(gclk));
	jnot g029(.din(w_G390gat_0[0]),.dout(n115),.clk(gclk));
	jor g030(.dina(w_n101_0[0]),.dinb(w_dff_B_hW8Se1yu8_1),.dout(w_dff_A_kFfvaOFK5_2),.clk(gclk));
	jand g031(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g033(.dina(w_n93_0[0]),.dinb(w_G55gat_0[2]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_n119_0[2]),.dinb(w_G29gat_0[0]),.dout(n120),.clk(gclk));
	jand g035(.dina(n120),.dinb(w_G68gat_0[1]),.dout(w_dff_A_oCZBiHiG0_2),.clk(gclk));
	jand g036(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n122),.clk(gclk));
	jand g037(.dina(w_n119_0[1]),.dinb(w_dff_B_aKz1ZNkd5_1),.dout(n123),.clk(gclk));
	jand g038(.dina(n123),.dinb(w_n122_0[1]),.dout(w_dff_A_WQugsFuT0_2),.clk(gclk));
	jand g039(.dina(w_n113_0[0]),.dinb(w_dff_B_JOj0NCKz0_1),.dout(w_dff_A_62IaO45P5_2),.clk(gclk));
	jxor g040(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n126),.clk(gclk));
	jxor g041(.dina(n126),.dinb(w_dff_B_EATIr7JD0_1),.dout(n127),.clk(gclk));
	jxor g042(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n128),.clk(gclk));
	jxor g043(.dina(n128),.dinb(w_G130gat_0[1]),.dout(n129),.clk(gclk));
	jxor g044(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G126gat_0[2]),.dinb(w_G121gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(n131),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n129),.dout(n133),.clk(gclk));
	jxor g048(.dina(n133),.dinb(w_dff_B_iA0hOQEb1_1),.dout(w_dff_A_OhvIt33J6_2),.clk(gclk));
	jxor g049(.dina(w_G189gat_2[1]),.dinb(w_G183gat_1[2]),.dout(n135),.clk(gclk));
	jxor g050(.dina(n135),.dinb(w_dff_B_R2xzlhF02_1),.dout(n136),.clk(gclk));
	jxor g051(.dina(w_G159gat_1[2]),.dinb(w_G130gat_0[0]),.dout(n137),.clk(gclk));
	jxor g052(.dina(n137),.dinb(w_G165gat_1[2]),.dout(n138),.clk(gclk));
	jxor g053(.dina(w_G177gat_1[2]),.dinb(w_G171gat_1[2]),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G201gat_1[1]),.dinb(w_G195gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n138),.dout(n142),.clk(gclk));
	jxor g057(.dina(n142),.dinb(w_dff_B_znr3Y1ok4_1),.dout(w_dff_A_ijyXFBE84_2),.clk(gclk));
	jnot g058(.din(w_G268gat_0[1]),.dout(n144),.clk(gclk));
	jand g059(.dina(w_G447gat_1),.dinb(w_G80gat_0[0]),.dout(n145),.clk(gclk));
	jand g060(.dina(n145),.dinb(w_n86_0[0]),.dout(n146),.clk(gclk));
	jand g061(.dina(w_n146_0[1]),.dinb(w_G55gat_0[1]),.dout(n147),.clk(gclk));
	jand g062(.dina(n147),.dinb(w_n144_0[1]),.dout(n148),.clk(gclk));
	jand g063(.dina(w_n111_0[0]),.dinb(w_n95_0[1]),.dout(n149),.clk(gclk));
	jnot g064(.din(w_n149_0[1]),.dout(n150),.clk(gclk));
	jand g065(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(w_G42gat_1[1]),.dinb(w_G17gat_2[0]),.dout(n152),.clk(gclk));
	jnot g067(.din(w_n152_0[1]),.dout(n153),.clk(gclk));
	jand g068(.dina(n153),.dinb(w_n151_0[1]),.dout(n154),.clk(gclk));
	jand g069(.dina(n154),.dinb(w_G447gat_0[2]),.dout(n155),.clk(gclk));
	jand g070(.dina(n155),.dinb(w_dff_B_Bhc3yBAC4_1),.dout(n156),.clk(gclk));
	jnot g071(.din(w_n92_0[0]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n104_0[0]),.dinb(w_G42gat_1[0]),.dout(n158),.clk(gclk));
	jand g073(.dina(w_G51gat_1[0]),.dinb(w_G17gat_1[2]),.dout(n159),.clk(gclk));
	jnot g074(.din(n159),.dout(n160),.clk(gclk));
	jor g075(.dina(n160),.dinb(n158),.dout(n161),.clk(gclk));
	jor g076(.dina(n161),.dinb(w_dff_B_za8Oaqir8_1),.dout(n162),.clk(gclk));
	jnot g077(.din(w_n162_0[1]),.dout(n163),.clk(gclk));
	jor g078(.dina(n163),.dinb(n156),.dout(n164),.clk(gclk));
	jand g079(.dina(w_n164_3[1]),.dinb(w_G126gat_0[1]),.dout(n165),.clk(gclk));
	jnot g080(.din(w_G156gat_0[0]),.dout(n166),.clk(gclk));
	jor g081(.dina(n166),.dinb(w_n108_0[0]),.dout(n167),.clk(gclk));
	jand g082(.dina(w_n167_0[1]),.dinb(w_G447gat_0[1]),.dout(n168),.clk(gclk));
	jand g083(.dina(w_n168_0[1]),.dinb(w_G17gat_1[1]),.dout(n169),.clk(gclk));
	jor g084(.dina(n169),.dinb(w_n97_0[0]),.dout(n170),.clk(gclk));
	jand g085(.dina(w_n170_1[1]),.dinb(w_G153gat_0[2]),.dout(n171),.clk(gclk));
	jor g086(.dina(w_dff_B_QdPGDnfW5_0),.dinb(n165),.dout(n172),.clk(gclk));
	jor g087(.dina(n172),.dinb(w_n148_1[2]),.dout(n173),.clk(gclk));
	jand g088(.dina(w_n173_0[1]),.dinb(w_G246gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_n122_0[0]),.dinb(w_G42gat_0[2]),.dout(n175),.clk(gclk));
	jand g090(.dina(G73gat),.dinb(G72gat),.dout(n176),.clk(gclk));
	jand g091(.dina(w_dff_B_fzp31Fxl5_0),.dinb(n175),.dout(n177),.clk(gclk));
	jand g092(.dina(n177),.dinb(w_n119_0[0]),.dout(n178),.clk(gclk));
	jand g093(.dina(w_n178_3[1]),.dinb(w_G201gat_1[0]),.dout(n179),.clk(gclk));
	jor g094(.dina(w_dff_B_rxaWXZwb5_0),.dinb(n174),.dout(n180),.clk(gclk));
	jnot g095(.din(w_G201gat_0[2]),.dout(n181),.clk(gclk));
	jnot g096(.din(w_n148_1[1]),.dout(n182),.clk(gclk));
	jnot g097(.din(w_G126gat_0[0]),.dout(n183),.clk(gclk));
	jnot g098(.din(w_G51gat_0[2]),.dout(n184),.clk(gclk));
	jor g099(.dina(w_n99_0[0]),.dinb(w_dff_B_0l3hpL6U6_1),.dout(n185),.clk(gclk));
	jor g100(.dina(w_n152_0[0]),.dinb(w_n167_0[0]),.dout(n186),.clk(gclk));
	jor g101(.dina(n186),.dinb(w_n185_0[1]),.dout(n187),.clk(gclk));
	jor g102(.dina(n187),.dinb(w_n149_0[0]),.dout(n188),.clk(gclk));
	jand g103(.dina(w_n162_0[0]),.dinb(n188),.dout(n189),.clk(gclk));
	jor g104(.dina(n189),.dinb(w_dff_B_28qe7Luv9_1),.dout(n190),.clk(gclk));
	jnot g105(.din(w_G153gat_0[1]),.dout(n191),.clk(gclk));
	jor g106(.dina(w_n151_0[0]),.dinb(w_n185_0[0]),.dout(n192),.clk(gclk));
	jor g107(.dina(n192),.dinb(w_n95_0[0]),.dout(n193),.clk(gclk));
	jand g108(.dina(n193),.dinb(w_G1gat_0[1]),.dout(n194),.clk(gclk));
	jor g109(.dina(n194),.dinb(w_dff_B_GOhcr1J55_1),.dout(n195),.clk(gclk));
	jand g110(.dina(n195),.dinb(n190),.dout(n196),.clk(gclk));
	jand g111(.dina(n196),.dinb(w_dff_B_OPiSdhep1_1),.dout(n197),.clk(gclk));
	jxor g112(.dina(w_n197_0[2]),.dinb(w_n181_0[2]),.dout(n198),.clk(gclk));
	jand g113(.dina(w_n198_0[2]),.dinb(w_G228gat_3[1]),.dout(n199),.clk(gclk));
	jand g114(.dina(w_n173_0[0]),.dinb(w_G201gat_0[1]),.dout(n200),.clk(gclk));
	jand g115(.dina(w_n200_0[1]),.dinb(w_G237gat_3[1]),.dout(n201),.clk(gclk));
	jand g116(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n202),.clk(gclk));
	jand g117(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n203),.clk(gclk));
	jor g118(.dina(n203),.dinb(n202),.dout(n204),.clk(gclk));
	jor g119(.dina(w_dff_B_8At1OGb22_0),.dinb(n201),.dout(n205),.clk(gclk));
	jor g120(.dina(n205),.dinb(w_dff_B_B7wikmcL3_1),.dout(n206),.clk(gclk));
	jor g121(.dina(n206),.dinb(w_dff_B_xWZxn00B9_1),.dout(n207),.clk(gclk));
	jor g122(.dina(w_n198_0[1]),.dinb(w_G261gat_0[2]),.dout(n208),.clk(gclk));
	jnot g123(.din(w_G261gat_0[1]),.dout(n209),.clk(gclk));
	jnot g124(.din(w_n198_0[0]),.dout(n210),.clk(gclk));
	jor g125(.dina(n210),.dinb(w_n209_0[1]),.dout(n211),.clk(gclk));
	jand g126(.dina(n211),.dinb(w_G219gat_3[2]),.dout(n212),.clk(gclk));
	jand g127(.dina(n212),.dinb(w_dff_B_8VdP2dtW9_1),.dout(n213),.clk(gclk));
	jor g128(.dina(n213),.dinb(n207),.dout(w_dff_A_nh87JbUt4_2),.clk(gclk));
	jand g129(.dina(w_n164_3[0]),.dinb(w_G111gat_0[1]),.dout(n215),.clk(gclk));
	jand g130(.dina(w_n170_1[0]),.dinb(w_G143gat_0[1]),.dout(n216),.clk(gclk));
	jor g131(.dina(n216),.dinb(w_n148_1[0]),.dout(n217),.clk(gclk));
	jor g132(.dina(n217),.dinb(n215),.dout(n218),.clk(gclk));
	jxor g133(.dina(w_n218_1[1]),.dinb(w_G183gat_1[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n219_0[2]),.dinb(w_G228gat_3[0]),.dout(n220),.clk(gclk));
	jand g135(.dina(w_n178_3[0]),.dinb(w_G183gat_1[0]),.dout(n221),.clk(gclk));
	jand g136(.dina(w_n218_1[0]),.dinb(w_G183gat_0[2]),.dout(n222),.clk(gclk));
	jand g137(.dina(w_n222_0[2]),.dinb(w_G237gat_3[0]),.dout(n223),.clk(gclk));
	jand g138(.dina(w_n218_0[2]),.dinb(w_G246gat_3[0]),.dout(n224),.clk(gclk));
	jand g139(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n225),.clk(gclk));
	jor g140(.dina(w_dff_B_FfPcPOOZ2_0),.dinb(n224),.dout(n226),.clk(gclk));
	jor g141(.dina(n226),.dinb(n223),.dout(n227),.clk(gclk));
	jor g142(.dina(n227),.dinb(w_dff_B_fMTMlvDt8_1),.dout(n228),.clk(gclk));
	jor g143(.dina(n228),.dinb(w_dff_B_qB1Nkhzo7_1),.dout(n229),.clk(gclk));
	jand g144(.dina(w_n164_2[2]),.dinb(w_G116gat_0[1]),.dout(n230),.clk(gclk));
	jand g145(.dina(w_n170_0[2]),.dinb(w_G146gat_0[1]),.dout(n231),.clk(gclk));
	jor g146(.dina(n231),.dinb(w_n148_0[2]),.dout(n232),.clk(gclk));
	jor g147(.dina(n232),.dinb(n230),.dout(n233),.clk(gclk));
	jand g148(.dina(w_n233_1[1]),.dinb(w_G189gat_2[0]),.dout(n234),.clk(gclk));
	jor g149(.dina(w_n233_1[0]),.dinb(w_G189gat_1[2]),.dout(n235),.clk(gclk));
	jand g150(.dina(w_n164_2[1]),.dinb(w_G121gat_0[0]),.dout(n236),.clk(gclk));
	jand g151(.dina(w_n170_0[1]),.dinb(w_G149gat_0[1]),.dout(n237),.clk(gclk));
	jor g152(.dina(n237),.dinb(w_n148_0[1]),.dout(n238),.clk(gclk));
	jor g153(.dina(n238),.dinb(n236),.dout(n239),.clk(gclk));
	jand g154(.dina(w_n239_1[1]),.dinb(w_G195gat_2[0]),.dout(n240),.clk(gclk));
	jor g155(.dina(w_n239_1[0]),.dinb(w_G195gat_1[2]),.dout(n241),.clk(gclk));
	jand g156(.dina(w_n197_0[1]),.dinb(w_n181_0[1]),.dout(n242),.clk(gclk));
	jnot g157(.din(w_n242_0[1]),.dout(n243),.clk(gclk));
	jor g158(.dina(w_n200_0[0]),.dinb(w_G261gat_0[0]),.dout(n244),.clk(gclk));
	jand g159(.dina(n244),.dinb(n243),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n245_0[1]),.dinb(w_n241_0[1]),.dout(n246),.clk(gclk));
	jor g161(.dina(n246),.dinb(w_n240_0[1]),.dout(n247),.clk(gclk));
	jand g162(.dina(w_n247_0[1]),.dinb(w_n235_0[1]),.dout(n248),.clk(gclk));
	jor g163(.dina(n248),.dinb(w_n234_0[1]),.dout(n249),.clk(gclk));
	jor g164(.dina(w_n249_0[1]),.dinb(w_n219_0[1]),.dout(n250),.clk(gclk));
	jnot g165(.din(w_n219_0[0]),.dout(n251),.clk(gclk));
	jnot g166(.din(w_n234_0[0]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n235_0[0]),.dout(n253),.clk(gclk));
	jnot g168(.din(w_n240_0[0]),.dout(n254),.clk(gclk));
	jnot g169(.din(w_n241_0[0]),.dout(n255),.clk(gclk));
	jor g170(.dina(w_n197_0[0]),.dinb(w_n181_0[0]),.dout(n256),.clk(gclk));
	jand g171(.dina(n256),.dinb(w_n209_0[0]),.dout(n257),.clk(gclk));
	jor g172(.dina(n257),.dinb(w_n242_0[0]),.dout(n258),.clk(gclk));
	jor g173(.dina(w_n258_0[1]),.dinb(w_dff_B_v3aEujkO0_1),.dout(n259),.clk(gclk));
	jand g174(.dina(n259),.dinb(w_dff_B_xrz6Q3Nn9_1),.dout(n260),.clk(gclk));
	jor g175(.dina(w_n260_0[1]),.dinb(w_dff_B_19NGwPN46_1),.dout(n261),.clk(gclk));
	jand g176(.dina(n261),.dinb(w_dff_B_spIMZWyK8_1),.dout(n262),.clk(gclk));
	jor g177(.dina(w_n262_0[1]),.dinb(w_dff_B_q38WAzoI3_1),.dout(n263),.clk(gclk));
	jand g178(.dina(n263),.dinb(w_G219gat_3[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(n264),.dinb(w_dff_B_qxPgZkMo9_1),.dout(n265),.clk(gclk));
	jor g180(.dina(n265),.dinb(w_dff_B_KIRMF6B32_1),.dout(w_dff_A_83XL4cAE0_2),.clk(gclk));
	jxor g181(.dina(w_n233_0[2]),.dinb(w_G189gat_1[1]),.dout(n267),.clk(gclk));
	jand g182(.dina(w_n267_0[2]),.dinb(w_G228gat_2[2]),.dout(n268),.clk(gclk));
	jand g183(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n269),.clk(gclk));
	jand g184(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n270),.clk(gclk));
	jor g185(.dina(n270),.dinb(w_G246gat_2[2]),.dout(n271),.clk(gclk));
	jand g186(.dina(w_dff_B_MwAU5TSD8_0),.dinb(w_n233_0[1]),.dout(n272),.clk(gclk));
	jor g187(.dina(n272),.dinb(w_dff_B_doc87SNp3_1),.dout(n273),.clk(gclk));
	jand g188(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n274),.clk(gclk));
	jand g189(.dina(w_n178_2[2]),.dinb(w_G189gat_0[2]),.dout(n275),.clk(gclk));
	jor g190(.dina(n275),.dinb(w_dff_B_6FXB3G1w8_1),.dout(n276),.clk(gclk));
	jor g191(.dina(w_dff_B_guoqX5rk6_0),.dinb(n273),.dout(n277),.clk(gclk));
	jor g192(.dina(n277),.dinb(w_dff_B_ip1O69zR9_1),.dout(n278),.clk(gclk));
	jor g193(.dina(w_n267_0[1]),.dinb(w_n247_0[0]),.dout(n279),.clk(gclk));
	jnot g194(.din(w_n267_0[0]),.dout(n280),.clk(gclk));
	jor g195(.dina(w_dff_B_EckWqqYc5_0),.dinb(w_n260_0[0]),.dout(n281),.clk(gclk));
	jand g196(.dina(n281),.dinb(w_G219gat_3[0]),.dout(n282),.clk(gclk));
	jand g197(.dina(n282),.dinb(w_dff_B_P64uaEJY4_1),.dout(n283),.clk(gclk));
	jor g198(.dina(n283),.dinb(w_dff_B_aisV8IiX3_1),.dout(w_dff_A_QaPWEmmy9_2),.clk(gclk));
	jxor g199(.dina(w_n239_0[2]),.dinb(w_G195gat_1[1]),.dout(n285),.clk(gclk));
	jand g200(.dina(w_n285_0[2]),.dinb(w_G228gat_2[1]),.dout(n286),.clk(gclk));
	jand g201(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n287),.clk(gclk));
	jand g202(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n288),.clk(gclk));
	jor g203(.dina(n288),.dinb(w_G246gat_2[1]),.dout(n289),.clk(gclk));
	jand g204(.dina(w_dff_B_FRm0f71R6_0),.dinb(w_n239_0[1]),.dout(n290),.clk(gclk));
	jor g205(.dina(n290),.dinb(w_dff_B_vvj0HpDe2_1),.dout(n291),.clk(gclk));
	jand g206(.dina(w_n178_2[1]),.dinb(w_G195gat_0[2]),.dout(n292),.clk(gclk));
	jand g207(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n293),.clk(gclk));
	jor g208(.dina(w_dff_B_MyHsY2ym2_0),.dinb(n292),.dout(n294),.clk(gclk));
	jor g209(.dina(w_dff_B_hXPlE1Gb5_0),.dinb(n291),.dout(n295),.clk(gclk));
	jor g210(.dina(n295),.dinb(w_dff_B_ndu5LyJR1_1),.dout(n296),.clk(gclk));
	jor g211(.dina(w_n285_0[1]),.dinb(w_n245_0[0]),.dout(n297),.clk(gclk));
	jnot g212(.din(w_n285_0[0]),.dout(n298),.clk(gclk));
	jor g213(.dina(w_dff_B_kH9ZOFXQ2_0),.dinb(w_n258_0[0]),.dout(n299),.clk(gclk));
	jand g214(.dina(n299),.dinb(w_G219gat_2[2]),.dout(n300),.clk(gclk));
	jand g215(.dina(n300),.dinb(w_dff_B_iNv189Yf9_1),.dout(n301),.clk(gclk));
	jor g216(.dina(n301),.dinb(w_dff_B_sBXG36rQ5_1),.dout(w_dff_A_KtnSHZjt1_2),.clk(gclk));
	jand g217(.dina(w_n168_0[0]),.dinb(w_G55gat_0[0]),.dout(n303),.clk(gclk));
	jand g218(.dina(w_n303_1[1]),.dinb(w_G143gat_0[0]),.dout(n304),.clk(gclk));
	jand g219(.dina(w_n146_0[0]),.dinb(w_G17gat_1[0]),.dout(n305),.clk(gclk));
	jand g220(.dina(n305),.dinb(w_n144_0[0]),.dout(n306),.clk(gclk));
	jor g221(.dina(w_n306_1[1]),.dinb(w_dff_B_VTLnXASP2_1),.dout(n307),.clk(gclk));
	jand g222(.dina(w_n164_2[0]),.dinb(w_G91gat_0[1]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n309),.clk(gclk));
	jor g224(.dina(w_dff_B_dfoDyUwa0_0),.dinb(n308),.dout(n310),.clk(gclk));
	jor g225(.dina(n310),.dinb(w_dff_B_K8VI0lyJ8_1),.dout(n311),.clk(gclk));
	jand g226(.dina(w_n311_1[2]),.dinb(w_G159gat_1[1]),.dout(n312),.clk(gclk));
	jor g227(.dina(w_n311_1[1]),.dinb(w_G159gat_1[0]),.dout(n313),.clk(gclk));
	jand g228(.dina(w_n164_1[2]),.dinb(w_G96gat_0[1]),.dout(n314),.clk(gclk));
	jand g229(.dina(w_n303_1[0]),.dinb(w_G146gat_0[0]),.dout(n315),.clk(gclk));
	jand g230(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n316),.clk(gclk));
	jor g231(.dina(w_dff_B_Lvdg5TNC7_0),.dinb(n315),.dout(n317),.clk(gclk));
	jor g232(.dina(w_dff_B_YIE4AI0Q3_0),.dinb(n314),.dout(n318),.clk(gclk));
	jor g233(.dina(n318),.dinb(w_n306_1[0]),.dout(n319),.clk(gclk));
	jand g234(.dina(w_n319_1[2]),.dinb(w_G165gat_1[1]),.dout(n320),.clk(gclk));
	jor g235(.dina(w_n319_1[1]),.dinb(w_G165gat_1[0]),.dout(n321),.clk(gclk));
	jand g236(.dina(w_n164_1[1]),.dinb(w_G101gat_0[1]),.dout(n322),.clk(gclk));
	jand g237(.dina(w_n303_0[2]),.dinb(w_G149gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n324),.clk(gclk));
	jor g239(.dina(w_dff_B_FNdWpG6L9_0),.dinb(n323),.dout(n325),.clk(gclk));
	jor g240(.dina(w_dff_B_WmpA10mb3_0),.dinb(n322),.dout(n326),.clk(gclk));
	jor g241(.dina(n326),.dinb(w_n306_0[2]),.dout(n327),.clk(gclk));
	jand g242(.dina(w_n327_1[2]),.dinb(w_G171gat_1[1]),.dout(n328),.clk(gclk));
	jor g243(.dina(w_n327_1[1]),.dinb(w_G171gat_1[0]),.dout(n329),.clk(gclk));
	jand g244(.dina(w_n164_1[0]),.dinb(w_G106gat_0[0]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n303_0[1]),.dinb(w_G153gat_0[0]),.dout(n331),.clk(gclk));
	jand g246(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n332),.clk(gclk));
	jor g247(.dina(w_dff_B_XIBcCA2F5_0),.dinb(n331),.dout(n333),.clk(gclk));
	jor g248(.dina(w_dff_B_i9r3DG767_0),.dinb(n330),.dout(n334),.clk(gclk));
	jor g249(.dina(n334),.dinb(w_n306_0[1]),.dout(n335),.clk(gclk));
	jand g250(.dina(w_n335_1[1]),.dinb(w_G177gat_1[1]),.dout(n336),.clk(gclk));
	jnot g251(.din(w_G177gat_1[0]),.dout(n337),.clk(gclk));
	jnot g252(.din(w_n335_1[0]),.dout(n338),.clk(gclk));
	jand g253(.dina(n338),.dinb(w_dff_B_CsfeRIgW3_1),.dout(n339),.clk(gclk));
	jnot g254(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jnot g255(.din(w_G183gat_0[1]),.dout(n341),.clk(gclk));
	jnot g256(.din(w_n218_0[1]),.dout(n342),.clk(gclk));
	jand g257(.dina(n342),.dinb(w_dff_B_LDgTm4kC5_1),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n343_0[1]),.dout(n344),.clk(gclk));
	jand g259(.dina(w_n249_0[0]),.dinb(w_dff_B_QKD3aOcz1_1),.dout(n345),.clk(gclk));
	jor g260(.dina(n345),.dinb(w_n222_0[1]),.dout(n346),.clk(gclk));
	jand g261(.dina(w_n346_0[1]),.dinb(w_dff_B_LS8NEahk2_1),.dout(n347),.clk(gclk));
	jor g262(.dina(n347),.dinb(w_n336_0[2]),.dout(n348),.clk(gclk));
	jand g263(.dina(w_n348_0[1]),.dinb(w_n329_0[1]),.dout(n349),.clk(gclk));
	jor g264(.dina(n349),.dinb(w_n328_0[1]),.dout(n350),.clk(gclk));
	jand g265(.dina(w_n350_0[1]),.dinb(w_n321_0[1]),.dout(n351),.clk(gclk));
	jor g266(.dina(n351),.dinb(w_n320_0[1]),.dout(n352),.clk(gclk));
	jand g267(.dina(w_n352_0[1]),.dinb(w_dff_B_t1cU3XPa1_1),.dout(n353),.clk(gclk));
	jor g268(.dina(n353),.dinb(w_dff_B_YPDy7Iun2_1),.dout(w_dff_A_lxhkViEa1_2),.clk(gclk));
	jxor g269(.dina(w_n335_0[2]),.dinb(w_G177gat_0[2]),.dout(n355),.clk(gclk));
	jnot g270(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n346_0[0]),.dinb(w_G219gat_2[1]),.dout(n357),.clk(gclk));
	jand g272(.dina(n357),.dinb(w_dff_B_6IKmdFBU2_1),.dout(n358),.clk(gclk));
	jnot g273(.din(w_n222_0[0]),.dout(n359),.clk(gclk));
	jor g274(.dina(w_n262_0[0]),.dinb(w_n343_0[0]),.dout(n360),.clk(gclk));
	jand g275(.dina(n360),.dinb(w_dff_B_niR2iSyj5_1),.dout(n361),.clk(gclk));
	jand g276(.dina(w_n361_0[1]),.dinb(w_G219gat_2[0]),.dout(n362),.clk(gclk));
	jor g277(.dina(n362),.dinb(w_G228gat_2[0]),.dout(n363),.clk(gclk));
	jand g278(.dina(n363),.dinb(w_n355_0[0]),.dout(n364),.clk(gclk));
	jand g279(.dina(w_n336_0[1]),.dinb(w_G237gat_2[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_n335_0[1]),.dinb(w_G246gat_2[0]),.dout(n366),.clk(gclk));
	jand g281(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n367),.clk(gclk));
	jand g282(.dina(w_n178_2[0]),.dinb(w_G177gat_0[1]),.dout(n368),.clk(gclk));
	jor g283(.dina(n368),.dinb(w_dff_B_q1deCKrm8_1),.dout(n369),.clk(gclk));
	jor g284(.dina(w_dff_B_wSRGaJsQ8_0),.dinb(n366),.dout(n370),.clk(gclk));
	jor g285(.dina(n370),.dinb(n365),.dout(n371),.clk(gclk));
	jor g286(.dina(w_dff_B_jrM5SpFM8_0),.dinb(n364),.dout(n372),.clk(gclk));
	jor g287(.dina(n372),.dinb(w_dff_B_SKllqSYH9_1),.dout(w_dff_A_L5KrTId14_2),.clk(gclk));
	jand g288(.dina(w_n311_1[0]),.dinb(w_G237gat_1[2]),.dout(n374),.clk(gclk));
	jor g289(.dina(n374),.dinb(w_n178_1[2]),.dout(n375),.clk(gclk));
	jand g290(.dina(n375),.dinb(w_G159gat_0[2]),.dout(n376),.clk(gclk));
	jxor g291(.dina(w_n311_0[2]),.dinb(w_G159gat_0[1]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_n377_0[2]),.dinb(w_G228gat_1[2]),.dout(n378),.clk(gclk));
	jand g293(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n379),.clk(gclk));
	jor g294(.dina(w_dff_B_lOKYu5SG3_0),.dinb(n378),.dout(n380),.clk(gclk));
	jand g295(.dina(w_n311_0[1]),.dinb(w_G246gat_1[2]),.dout(n381),.clk(gclk));
	jor g296(.dina(w_dff_B_vMeloIfP0_0),.dinb(n380),.dout(n382),.clk(gclk));
	jor g297(.dina(n382),.dinb(w_dff_B_JdO4DSjG8_1),.dout(n383),.clk(gclk));
	jor g298(.dina(w_n377_0[1]),.dinb(w_n352_0[0]),.dout(n384),.clk(gclk));
	jnot g299(.din(w_n320_0[0]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n321_0[0]),.dout(n386),.clk(gclk));
	jnot g301(.din(w_n328_0[0]),.dout(n387),.clk(gclk));
	jnot g302(.din(w_n329_0[0]),.dout(n388),.clk(gclk));
	jnot g303(.din(w_n336_0[0]),.dout(n389),.clk(gclk));
	jor g304(.dina(w_n361_0[0]),.dinb(w_n339_0[0]),.dout(n390),.clk(gclk));
	jand g305(.dina(n390),.dinb(w_dff_B_oP1zgrp35_1),.dout(n391),.clk(gclk));
	jor g306(.dina(w_n391_0[1]),.dinb(w_dff_B_8w1OuQ7g3_1),.dout(n392),.clk(gclk));
	jand g307(.dina(n392),.dinb(w_dff_B_MLzv1ZkU1_1),.dout(n393),.clk(gclk));
	jor g308(.dina(w_n393_0[1]),.dinb(w_dff_B_Bo7oQoJK8_1),.dout(n394),.clk(gclk));
	jand g309(.dina(n394),.dinb(w_dff_B_a428seju5_1),.dout(n395),.clk(gclk));
	jnot g310(.din(w_n377_0[0]),.dout(n396),.clk(gclk));
	jor g311(.dina(w_dff_B_zAgfXo5z3_0),.dinb(n395),.dout(n397),.clk(gclk));
	jand g312(.dina(n397),.dinb(w_G219gat_1[2]),.dout(n398),.clk(gclk));
	jand g313(.dina(n398),.dinb(w_dff_B_L92F2ZAH0_1),.dout(n399),.clk(gclk));
	jor g314(.dina(n399),.dinb(w_dff_B_Eiyg7v3H6_1),.dout(G878gat),.clk(gclk));
	jand g315(.dina(w_n319_1[0]),.dinb(w_G237gat_1[1]),.dout(n401),.clk(gclk));
	jor g316(.dina(n401),.dinb(w_n178_1[1]),.dout(n402),.clk(gclk));
	jand g317(.dina(n402),.dinb(w_G165gat_0[2]),.dout(n403),.clk(gclk));
	jxor g318(.dina(w_n319_0[2]),.dinb(w_G165gat_0[1]),.dout(n404),.clk(gclk));
	jand g319(.dina(w_n404_0[2]),.dinb(w_G228gat_1[1]),.dout(n405),.clk(gclk));
	jand g320(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n406),.clk(gclk));
	jor g321(.dina(w_dff_B_L6Cx6YAe2_0),.dinb(n405),.dout(n407),.clk(gclk));
	jand g322(.dina(w_n319_0[1]),.dinb(w_G246gat_1[1]),.dout(n408),.clk(gclk));
	jor g323(.dina(w_dff_B_uMvaqNZj5_0),.dinb(n407),.dout(n409),.clk(gclk));
	jor g324(.dina(n409),.dinb(w_dff_B_dlwkneye3_1),.dout(n410),.clk(gclk));
	jor g325(.dina(w_n404_0[1]),.dinb(w_n350_0[0]),.dout(n411),.clk(gclk));
	jnot g326(.din(w_n404_0[0]),.dout(n412),.clk(gclk));
	jor g327(.dina(w_dff_B_hzZ3zAfb8_0),.dinb(w_n393_0[0]),.dout(n413),.clk(gclk));
	jand g328(.dina(n413),.dinb(w_G219gat_1[1]),.dout(n414),.clk(gclk));
	jand g329(.dina(n414),.dinb(w_dff_B_2eA68JVH7_1),.dout(n415),.clk(gclk));
	jor g330(.dina(n415),.dinb(w_dff_B_qpsPCDeK3_1),.dout(w_dff_A_wWIeNAhW9_2),.clk(gclk));
	jand g331(.dina(w_n327_1[0]),.dinb(w_G237gat_1[0]),.dout(n417),.clk(gclk));
	jor g332(.dina(n417),.dinb(w_n178_1[0]),.dout(n418),.clk(gclk));
	jand g333(.dina(n418),.dinb(w_G171gat_0[2]),.dout(n419),.clk(gclk));
	jxor g334(.dina(w_n327_0[2]),.dinb(w_G171gat_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n420_0[2]),.dinb(w_G228gat_1[0]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jor g337(.dina(w_dff_B_X1cVvvvP1_0),.dinb(n421),.dout(n423),.clk(gclk));
	jand g338(.dina(w_n327_0[1]),.dinb(w_G246gat_1[0]),.dout(n424),.clk(gclk));
	jor g339(.dina(w_dff_B_1lNdlfgg1_0),.dinb(n423),.dout(n425),.clk(gclk));
	jor g340(.dina(n425),.dinb(w_dff_B_yW24bOoj0_1),.dout(n426),.clk(gclk));
	jnot g341(.din(w_n420_0[1]),.dout(n427),.clk(gclk));
	jor g342(.dina(w_dff_B_vuZe0bKa8_0),.dinb(w_n391_0[0]),.dout(n428),.clk(gclk));
	jor g343(.dina(w_n420_0[0]),.dinb(w_n348_0[0]),.dout(n429),.clk(gclk));
	jand g344(.dina(n429),.dinb(w_G219gat_1[0]),.dout(n430),.clk(gclk));
	jand g345(.dina(n430),.dinb(w_dff_B_rAKNhPEe8_1),.dout(n431),.clk(gclk));
	jor g346(.dina(n431),.dinb(w_dff_B_TMxMNK401_1),.dout(w_dff_A_vX37Lua63_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_dff_A_0qB5OCiB0_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_dff_A_YZFSoUtL7_1),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_dff_A_c58gNbtU5_0),.doutb(w_dff_A_ILxZoKM10_1),.doutc(w_G17gat_1[2]),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_dff_A_hUzUa7W96_2),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_dff_A_MKDZ5sdi8_0),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_dff_A_LtKNNQCe6_1),.doutc(w_dff_A_e94DEHcZ9_2),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_dff_A_BQoxbgMb8_0),.doutb(w_G42gat_1[1]),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_dff_A_Gf9ahnaf0_1),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_dff_A_o0FLiivG4_0),.doutb(w_dff_A_nKJDjkL34_1),.doutc(w_G55gat_0[2]),.din(w_dff_B_xxKpXUDp7_3));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_dff_A_8SHFtRHc4_1),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_dff_A_jwJe59Ba3_0),.doutb(w_G80gat_0[1]),.doutc(w_dff_A_c5k75pdr7_2),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_dff_A_oTpOBk6E7_1),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_dff_A_WHbkWSbK3_1),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_dff_A_1ljbPany4_1),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_B83qHL3A6_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_dff_A_8giyetID5_1),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_dff_A_a6m6ldqn7_1),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_dff_A_FdI0WKCU2_0),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl3 jspl3_w_G126gat_0(.douta(w_G126gat_0[0]),.doutb(w_dff_A_J9u0xkXT3_1),.doutc(w_G126gat_0[2]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_dff_A_QyOVgLYl6_1),.din(G130gat));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_dff_A_wZPeJeD78_1),.din(w_dff_B_dot5MtOb6_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_dff_A_483dyFML3_1),.din(w_dff_B_h0oRvhMQ9_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_dff_A_DbDIXG4L9_1),.din(w_dff_B_QQafkqky1_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_dff_A_kXQhz9PI4_0),.doutb(w_G153gat_0[1]),.doutc(w_dff_A_26RT9joY1_2),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_dff_A_Tf2lEuFd3_1),.doutc(w_dff_A_R0RX7xce5_2),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_dff_A_VPQapodH2_0),.doutb(w_dff_A_uXT30LP58_1),.doutc(w_G159gat_1[2]),.din(w_G159gat_0[0]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_dff_A_aaz0C0hF6_1),.doutc(w_dff_A_47HpDG880_2),.din(w_dff_B_zMkHJ0nj7_3));
	jspl3 jspl3_w_G165gat_1(.douta(w_dff_A_aBmZ5SFr4_0),.doutb(w_dff_A_20PT5cV23_1),.doutc(w_G165gat_1[2]),.din(w_G165gat_0[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_dff_A_cLI7CXP81_1),.doutc(w_dff_A_SoV7oXqQ8_2),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_dff_A_02D4fnOb6_0),.doutb(w_dff_A_g03eD6ey0_1),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_dff_A_8z0yNlva8_1),.doutc(w_dff_A_fapqLrpq9_2),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_dff_A_ZQhRPJSx0_1),.doutc(w_G177gat_1[2]),.din(w_G177gat_0[0]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_dff_A_OWSYhHc90_2),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_dff_A_5wvFnafV4_0),.doutb(w_dff_A_Vael7ZcZ0_1),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_dff_A_MQ4ZGfIg5_2),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_dff_A_gaObyY8W5_1),.doutc(w_dff_A_WSQG2nQG3_2),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_dff_A_14aERbys4_0),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_dff_A_kKqLSNdp8_2),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_dff_A_lU1z5EkX9_1),.doutc(w_dff_A_C5Xdz3Bg2_2),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_dff_A_LuLFkDYT4_0),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_dff_A_ZBaVSZNC1_1),.doutc(w_G201gat_0[2]),.din(G201gat));
	jspl jspl_w_G201gat_1(.douta(w_dff_A_s18ggExM6_0),.doutb(w_G201gat_1[1]),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_koVGwb1J7_0),.doutb(w_dff_A_LIhv0HB99_1),.doutc(w_G219gat_0[2]),.din(w_dff_B_m5Gj2lRU7_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_G219gat_1[0]),.doutb(w_dff_A_dT4pKEOP1_1),.doutc(w_dff_A_Js3VHItE4_2),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_5bL57tID5_0),.doutb(w_dff_A_wAl3WvJh8_1),.doutc(w_G219gat_2[2]),.din(w_G219gat_0[1]));
	jspl3 jspl3_w_G219gat_3(.douta(w_dff_A_ShCjBaep4_0),.doutb(w_dff_A_u2etzkMM4_1),.doutc(w_G219gat_3[2]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_dff_A_jpgYigNZ1_0),.doutb(w_G228gat_0[1]),.doutc(w_G228gat_0[2]),.din(w_dff_B_CFuqkUPg8_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_dff_A_cLdcIYs66_0),.doutb(w_G228gat_2[1]),.doutc(w_G228gat_2[2]),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_dff_A_Qw9v7Yie2_1),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_dff_A_pJ1fMVAp6_0),.doutb(w_G237gat_0[1]),.doutc(w_dff_A_8DAk1jc00_2),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_dff_A_NMD8Frsu5_0),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_dff_A_4EqwaagK7_1),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_dff_A_bJRktpWx4_0),.doutb(w_G246gat_0[1]),.doutc(w_dff_A_jUMdPeOn3_2),.din(w_dff_B_FuEt0jiw2_3));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_dff_A_aSHbGEry9_0),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_dff_A_m9gDeRoh0_1),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_dff_A_xvKkIVhB3_0),.doutb(w_G261gat_0[1]),.doutc(w_dff_A_tWLi3I009_2),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_dff_A_rew4hahm7_1),.doutc(w_dff_A_B6Z4XMwz7_2),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_dff_A_QWcMVJQJ4_2),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(w_dff_A_lEJ8kvaV2_1),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_dff_A_mQhW8Len8_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n95_0(.douta(w_dff_A_HbOCAKGA8_0),.doutb(w_n95_0[1]),.doutc(w_dff_A_B2NdSyJ34_2),.din(n95));
	jspl jspl_w_n97_0(.douta(w_dff_A_xEFdfxMG1_0),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.din(w_dff_B_xgt7oxkw4_2));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_dff_A_xFSlZ5xQ9_1),.din(n111));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.din(n113));
	jspl3 jspl3_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.doutc(w_n119_0[2]),.din(n119));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_dff_A_uDr2tGyW1_1),.din(n122));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(w_dff_B_P7cmgdDp0_2));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_n148_1[0]),.doutb(w_n148_1[1]),.doutc(w_dff_A_PlGa8xbR6_2),.din(w_n148_0[0]));
	jspl jspl_w_n149_0(.douta(w_dff_A_wiFWWXhH9_0),.doutb(w_n149_0[1]),.din(n149));
	jspl jspl_w_n151_0(.douta(w_dff_A_7uVQtD3w3_0),.doutb(w_n151_0[1]),.din(w_dff_B_dvlmMZNO4_2));
	jspl jspl_w_n152_0(.douta(w_dff_A_iD8pjJNg7_0),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n162_0(.douta(w_dff_A_o7YaiDDE6_0),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_n164_0[2]),.din(n164));
	jspl3 jspl3_w_n164_1(.douta(w_n164_1[0]),.doutb(w_n164_1[1]),.doutc(w_n164_1[2]),.din(w_n164_0[0]));
	jspl3 jspl3_w_n164_2(.douta(w_n164_2[0]),.doutb(w_n164_2[1]),.doutc(w_n164_2[2]),.din(w_n164_0[1]));
	jspl jspl_w_n164_3(.douta(w_n164_3[0]),.doutb(w_n164_3[1]),.din(w_n164_0[2]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n170_1(.douta(w_n170_1[0]),.doutb(w_n170_1[1]),.din(w_n170_0[0]));
	jspl jspl_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.din(n173));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_VzplXodn2_0),.doutb(w_n178_0[1]),.doutc(w_n178_0[2]),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_n178_1[1]),.doutc(w_n178_1[2]),.din(w_n178_0[0]));
	jspl3 jspl3_w_n178_2(.douta(w_n178_2[0]),.doutb(w_n178_2[1]),.doutc(w_n178_2[2]),.din(w_n178_0[1]));
	jspl jspl_w_n178_3(.douta(w_n178_3[0]),.doutb(w_n178_3[1]),.din(w_n178_0[2]));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(w_dff_B_04yVh3Ik9_3));
	jspl jspl_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.din(n185));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_n198_0[2]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_dff_A_UVuRWb7K0_1),.din(w_dff_B_f1hnKObp1_2));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_n218_0[2]),.din(n218));
	jspl jspl_w_n218_1(.douta(w_n218_1[0]),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl3 jspl3_w_n219_0(.douta(w_n219_0[0]),.doutb(w_dff_A_WKAyP4vq4_1),.doutc(w_n219_0[2]),.din(n219));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_dff_A_4LfsyQc45_1),.doutc(w_n222_0[2]),.din(n222));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl jspl_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.din(w_n233_0[0]));
	jspl jspl_w_n234_0(.douta(w_n234_0[0]),.doutb(w_dff_A_iU1DSUeC9_1),.din(n234));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_dff_A_NQy8YkrC9_1),.din(n235));
	jspl3 jspl3_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.doutc(w_n239_0[2]),.din(n239));
	jspl jspl_w_n239_1(.douta(w_n239_1[0]),.doutb(w_n239_1[1]),.din(w_n239_0[0]));
	jspl jspl_w_n240_0(.douta(w_n240_0[0]),.doutb(w_dff_A_9r8CxF4s7_1),.din(n240));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_dff_A_quB8R3mO5_1),.din(n241));
	jspl jspl_w_n242_0(.douta(w_dff_A_BR6IopgH9_0),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.din(n258));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl jspl_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_dff_A_oIwOpkCN4_1),.doutc(w_n267_0[2]),.din(n267));
	jspl3 jspl3_w_n285_0(.douta(w_n285_0[0]),.doutb(w_dff_A_2sd0l6IR0_1),.doutc(w_n285_0[2]),.din(n285));
	jspl3 jspl3_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.doutc(w_n303_0[2]),.din(n303));
	jspl jspl_w_n303_1(.douta(w_n303_1[0]),.doutb(w_n303_1[1]),.din(w_n303_0[0]));
	jspl3 jspl3_w_n306_0(.douta(w_n306_0[0]),.doutb(w_dff_A_PUuizGx86_1),.doutc(w_dff_A_MAiR4MzR9_2),.din(n306));
	jspl jspl_w_n306_1(.douta(w_dff_A_aZ5BSb7c0_0),.doutb(w_n306_1[1]),.din(w_n306_0[0]));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.doutc(w_n311_0[2]),.din(n311));
	jspl3 jspl3_w_n311_1(.douta(w_n311_1[0]),.doutb(w_n311_1[1]),.doutc(w_n311_1[2]),.din(w_n311_0[0]));
	jspl3 jspl3_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.doutc(w_n319_0[2]),.din(n319));
	jspl3 jspl3_w_n319_1(.douta(w_n319_1[0]),.doutb(w_n319_1[1]),.doutc(w_n319_1[2]),.din(w_n319_0[0]));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_dff_A_40zSHeLb7_1),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_dff_A_axQuh9PX7_1),.din(n321));
	jspl3 jspl3_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.doutc(w_n327_0[2]),.din(n327));
	jspl3 jspl3_w_n327_1(.douta(w_n327_1[0]),.doutb(w_n327_1[1]),.doutc(w_n327_1[2]),.din(w_n327_0[0]));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_dff_A_FTobAgMp7_1),.din(n328));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_dff_A_7tkxUkqg0_1),.din(n329));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl jspl_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.din(w_n335_0[0]));
	jspl3 jspl3_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.doutc(w_dff_A_ipW7HfAD2_2),.din(n336));
	jspl jspl_w_n339_0(.douta(w_dff_A_NxHilTNr9_0),.doutb(w_n339_0[1]),.din(n339));
	jspl jspl_w_n343_0(.douta(w_dff_A_rxyxfakq4_0),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n352_0(.douta(w_n352_0[0]),.doutb(w_n352_0[1]),.din(n352));
	jspl jspl_w_n355_0(.douta(w_dff_A_FJFDQy9s7_0),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_dff_A_kgIBAwiY8_1),.doutc(w_n377_0[2]),.din(n377));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(n391));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_dff_A_Ye0keKFV5_1),.doutc(w_n404_0[2]),.din(n404));
	jspl3 jspl3_w_n420_0(.douta(w_dff_A_Jf5HE9pc1_0),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jdff dff_B_xgt7oxkw4_2(.din(n103),.dout(w_dff_B_xgt7oxkw4_2),.clk(gclk));
	jdff dff_B_aBFOmxD08_1(.din(G90gat),.dout(w_dff_B_aBFOmxD08_1),.clk(gclk));
	jdff dff_B_hW8Se1yu8_1(.din(n115),.dout(w_dff_B_hW8Se1yu8_1),.clk(gclk));
	jdff dff_B_owR0xsDs9_1(.din(n96),.dout(w_dff_B_owR0xsDs9_1),.clk(gclk));
	jdff dff_A_oxB3695r7_1(.dout(w_G390gat_0[1]),.din(w_dff_A_oxB3695r7_1),.clk(gclk));
	jdff dff_A_rew4hahm7_1(.dout(w_dff_A_oxB3695r7_1),.din(w_dff_A_rew4hahm7_1),.clk(gclk));
	jdff dff_B_Skdtk8Un0_1(.din(G74gat),.dout(w_dff_B_Skdtk8Un0_1),.clk(gclk));
	jdff dff_B_5UUizARO8_1(.din(w_dff_B_Skdtk8Un0_1),.dout(w_dff_B_5UUizARO8_1),.clk(gclk));
	jdff dff_B_aKz1ZNkd5_1(.din(w_dff_B_5UUizARO8_1),.dout(w_dff_B_aKz1ZNkd5_1),.clk(gclk));
	jdff dff_B_JOj0NCKz0_1(.din(G89gat),.dout(w_dff_B_JOj0NCKz0_1),.clk(gclk));
	jdff dff_B_iA0hOQEb1_1(.din(n127),.dout(w_dff_B_iA0hOQEb1_1),.clk(gclk));
	jdff dff_B_EATIr7JD0_1(.din(G135gat),.dout(w_dff_B_EATIr7JD0_1),.clk(gclk));
	jdff dff_B_znr3Y1ok4_1(.din(n136),.dout(w_dff_B_znr3Y1ok4_1),.clk(gclk));
	jdff dff_A_QyOVgLYl6_1(.dout(w_G130gat_0[1]),.din(w_dff_A_QyOVgLYl6_1),.clk(gclk));
	jdff dff_B_R2xzlhF02_1(.din(G207gat),.dout(w_dff_B_R2xzlhF02_1),.clk(gclk));
	jdff dff_B_JS1LUrZv1_1(.din(n208),.dout(w_dff_B_JS1LUrZv1_1),.clk(gclk));
	jdff dff_B_8VdP2dtW9_1(.din(w_dff_B_JS1LUrZv1_1),.dout(w_dff_B_8VdP2dtW9_1),.clk(gclk));
	jdff dff_B_CEQ0uHYm7_1(.din(n180),.dout(w_dff_B_CEQ0uHYm7_1),.clk(gclk));
	jdff dff_B_xWZxn00B9_1(.din(w_dff_B_CEQ0uHYm7_1),.dout(w_dff_B_xWZxn00B9_1),.clk(gclk));
	jdff dff_B_B7wikmcL3_1(.din(n199),.dout(w_dff_B_B7wikmcL3_1),.clk(gclk));
	jdff dff_B_KEyhOJQ37_0(.din(n204),.dout(w_dff_B_KEyhOJQ37_0),.clk(gclk));
	jdff dff_B_ZUokzprQ2_0(.din(w_dff_B_KEyhOJQ37_0),.dout(w_dff_B_ZUokzprQ2_0),.clk(gclk));
	jdff dff_B_ULczbqEV6_0(.din(w_dff_B_ZUokzprQ2_0),.dout(w_dff_B_ULczbqEV6_0),.clk(gclk));
	jdff dff_B_Ac0ERhlf8_0(.din(w_dff_B_ULczbqEV6_0),.dout(w_dff_B_Ac0ERhlf8_0),.clk(gclk));
	jdff dff_B_6x74zz1B1_0(.din(w_dff_B_Ac0ERhlf8_0),.dout(w_dff_B_6x74zz1B1_0),.clk(gclk));
	jdff dff_B_x4rpQqzp7_0(.din(w_dff_B_6x74zz1B1_0),.dout(w_dff_B_x4rpQqzp7_0),.clk(gclk));
	jdff dff_B_go5S0cmU4_0(.din(w_dff_B_x4rpQqzp7_0),.dout(w_dff_B_go5S0cmU4_0),.clk(gclk));
	jdff dff_B_bZEgn9VB7_0(.din(w_dff_B_go5S0cmU4_0),.dout(w_dff_B_bZEgn9VB7_0),.clk(gclk));
	jdff dff_B_8At1OGb22_0(.din(w_dff_B_bZEgn9VB7_0),.dout(w_dff_B_8At1OGb22_0),.clk(gclk));
	jdff dff_B_Ff6YlyyZ8_0(.din(n179),.dout(w_dff_B_Ff6YlyyZ8_0),.clk(gclk));
	jdff dff_B_hoMlVHfk7_0(.din(w_dff_B_Ff6YlyyZ8_0),.dout(w_dff_B_hoMlVHfk7_0),.clk(gclk));
	jdff dff_B_msmmgGy76_0(.din(w_dff_B_hoMlVHfk7_0),.dout(w_dff_B_msmmgGy76_0),.clk(gclk));
	jdff dff_B_93RQjyTa9_0(.din(w_dff_B_msmmgGy76_0),.dout(w_dff_B_93RQjyTa9_0),.clk(gclk));
	jdff dff_B_rxaWXZwb5_0(.din(w_dff_B_93RQjyTa9_0),.dout(w_dff_B_rxaWXZwb5_0),.clk(gclk));
	jdff dff_A_2qre1vtb0_0(.dout(w_G201gat_1[0]),.din(w_dff_A_2qre1vtb0_0),.clk(gclk));
	jdff dff_A_3sQMLgiR6_0(.dout(w_dff_A_2qre1vtb0_0),.din(w_dff_A_3sQMLgiR6_0),.clk(gclk));
	jdff dff_A_S4nVfOFY5_0(.dout(w_dff_A_3sQMLgiR6_0),.din(w_dff_A_S4nVfOFY5_0),.clk(gclk));
	jdff dff_A_s18ggExM6_0(.dout(w_dff_A_S4nVfOFY5_0),.din(w_dff_A_s18ggExM6_0),.clk(gclk));
	jdff dff_B_adwAZrNl7_1(.din(n229),.dout(w_dff_B_adwAZrNl7_1),.clk(gclk));
	jdff dff_B_9STfpRbb1_1(.din(w_dff_B_adwAZrNl7_1),.dout(w_dff_B_9STfpRbb1_1),.clk(gclk));
	jdff dff_B_XVpX5orf8_1(.din(w_dff_B_9STfpRbb1_1),.dout(w_dff_B_XVpX5orf8_1),.clk(gclk));
	jdff dff_B_Aj6bGocO9_1(.din(w_dff_B_XVpX5orf8_1),.dout(w_dff_B_Aj6bGocO9_1),.clk(gclk));
	jdff dff_B_UuHxarYi1_1(.din(w_dff_B_Aj6bGocO9_1),.dout(w_dff_B_UuHxarYi1_1),.clk(gclk));
	jdff dff_B_KIRMF6B32_1(.din(w_dff_B_UuHxarYi1_1),.dout(w_dff_B_KIRMF6B32_1),.clk(gclk));
	jdff dff_B_qxPgZkMo9_1(.din(n250),.dout(w_dff_B_qxPgZkMo9_1),.clk(gclk));
	jdff dff_B_D54inTRd9_1(.din(n251),.dout(w_dff_B_D54inTRd9_1),.clk(gclk));
	jdff dff_B_3r0BZzul0_1(.din(w_dff_B_D54inTRd9_1),.dout(w_dff_B_3r0BZzul0_1),.clk(gclk));
	jdff dff_B_xOF3U8Xw3_1(.din(w_dff_B_3r0BZzul0_1),.dout(w_dff_B_xOF3U8Xw3_1),.clk(gclk));
	jdff dff_B_wQZuk2hL6_1(.din(w_dff_B_xOF3U8Xw3_1),.dout(w_dff_B_wQZuk2hL6_1),.clk(gclk));
	jdff dff_B_XUaNJjtM9_1(.din(w_dff_B_wQZuk2hL6_1),.dout(w_dff_B_XUaNJjtM9_1),.clk(gclk));
	jdff dff_B_q38WAzoI3_1(.din(w_dff_B_XUaNJjtM9_1),.dout(w_dff_B_q38WAzoI3_1),.clk(gclk));
	jdff dff_B_E03aGQNB0_1(.din(n220),.dout(w_dff_B_E03aGQNB0_1),.clk(gclk));
	jdff dff_B_qB1Nkhzo7_1(.din(w_dff_B_E03aGQNB0_1),.dout(w_dff_B_qB1Nkhzo7_1),.clk(gclk));
	jdff dff_B_AOd4uBUG8_1(.din(n221),.dout(w_dff_B_AOd4uBUG8_1),.clk(gclk));
	jdff dff_B_GMQ21RxZ9_1(.din(w_dff_B_AOd4uBUG8_1),.dout(w_dff_B_GMQ21RxZ9_1),.clk(gclk));
	jdff dff_B_MfxyW0mO9_1(.din(w_dff_B_GMQ21RxZ9_1),.dout(w_dff_B_MfxyW0mO9_1),.clk(gclk));
	jdff dff_B_I2iIPerq3_1(.din(w_dff_B_MfxyW0mO9_1),.dout(w_dff_B_I2iIPerq3_1),.clk(gclk));
	jdff dff_B_U9M9dbaP5_1(.din(w_dff_B_I2iIPerq3_1),.dout(w_dff_B_U9M9dbaP5_1),.clk(gclk));
	jdff dff_B_fMTMlvDt8_1(.din(w_dff_B_U9M9dbaP5_1),.dout(w_dff_B_fMTMlvDt8_1),.clk(gclk));
	jdff dff_B_Rk0ofG141_0(.din(n225),.dout(w_dff_B_Rk0ofG141_0),.clk(gclk));
	jdff dff_B_j7bbZSaO0_0(.din(w_dff_B_Rk0ofG141_0),.dout(w_dff_B_j7bbZSaO0_0),.clk(gclk));
	jdff dff_B_HlYbTumq8_0(.din(w_dff_B_j7bbZSaO0_0),.dout(w_dff_B_HlYbTumq8_0),.clk(gclk));
	jdff dff_B_9rO6rsWT1_0(.din(w_dff_B_HlYbTumq8_0),.dout(w_dff_B_9rO6rsWT1_0),.clk(gclk));
	jdff dff_B_mlZQReuw7_0(.din(w_dff_B_9rO6rsWT1_0),.dout(w_dff_B_mlZQReuw7_0),.clk(gclk));
	jdff dff_B_wrUscLWM9_0(.din(w_dff_B_mlZQReuw7_0),.dout(w_dff_B_wrUscLWM9_0),.clk(gclk));
	jdff dff_B_LdQumMHy9_0(.din(w_dff_B_wrUscLWM9_0),.dout(w_dff_B_LdQumMHy9_0),.clk(gclk));
	jdff dff_B_FfPcPOOZ2_0(.din(w_dff_B_LdQumMHy9_0),.dout(w_dff_B_FfPcPOOZ2_0),.clk(gclk));
	jdff dff_A_m9gDeRoh0_1(.dout(w_G246gat_3[1]),.din(w_dff_A_m9gDeRoh0_1),.clk(gclk));
	jdff dff_A_4EqwaagK7_1(.dout(w_G237gat_3[1]),.din(w_dff_A_4EqwaagK7_1),.clk(gclk));
	jdff dff_A_jRK70mNr4_1(.dout(w_n219_0[1]),.din(w_dff_A_jRK70mNr4_1),.clk(gclk));
	jdff dff_A_f8WcpeTE4_1(.dout(w_dff_A_jRK70mNr4_1),.din(w_dff_A_f8WcpeTE4_1),.clk(gclk));
	jdff dff_A_jrbqh4QO7_1(.dout(w_dff_A_f8WcpeTE4_1),.din(w_dff_A_jrbqh4QO7_1),.clk(gclk));
	jdff dff_A_643Jw5Qk2_1(.dout(w_dff_A_jrbqh4QO7_1),.din(w_dff_A_643Jw5Qk2_1),.clk(gclk));
	jdff dff_A_3G8nFk7W0_1(.dout(w_dff_A_643Jw5Qk2_1),.din(w_dff_A_3G8nFk7W0_1),.clk(gclk));
	jdff dff_A_YV6a4Gzn5_1(.dout(w_dff_A_3G8nFk7W0_1),.din(w_dff_A_YV6a4Gzn5_1),.clk(gclk));
	jdff dff_A_WKAyP4vq4_1(.dout(w_dff_A_YV6a4Gzn5_1),.din(w_dff_A_WKAyP4vq4_1),.clk(gclk));
	jdff dff_A_h6i5PYEH4_0(.dout(w_G183gat_1[0]),.din(w_dff_A_h6i5PYEH4_0),.clk(gclk));
	jdff dff_A_7H5fcfOu9_0(.dout(w_dff_A_h6i5PYEH4_0),.din(w_dff_A_7H5fcfOu9_0),.clk(gclk));
	jdff dff_A_nFhN0sVP9_0(.dout(w_dff_A_7H5fcfOu9_0),.din(w_dff_A_nFhN0sVP9_0),.clk(gclk));
	jdff dff_A_5wvFnafV4_0(.dout(w_dff_A_nFhN0sVP9_0),.din(w_dff_A_5wvFnafV4_0),.clk(gclk));
	jdff dff_A_LefcYNt21_1(.dout(w_G183gat_1[1]),.din(w_dff_A_LefcYNt21_1),.clk(gclk));
	jdff dff_A_fbAfghFz1_1(.dout(w_dff_A_LefcYNt21_1),.din(w_dff_A_fbAfghFz1_1),.clk(gclk));
	jdff dff_A_bdjxU63K5_1(.dout(w_dff_A_fbAfghFz1_1),.din(w_dff_A_bdjxU63K5_1),.clk(gclk));
	jdff dff_A_v4YiKeId8_1(.dout(w_dff_A_bdjxU63K5_1),.din(w_dff_A_v4YiKeId8_1),.clk(gclk));
	jdff dff_A_r9tAbfMX6_1(.dout(w_dff_A_v4YiKeId8_1),.din(w_dff_A_r9tAbfMX6_1),.clk(gclk));
	jdff dff_A_ePi6SFEE7_1(.dout(w_dff_A_r9tAbfMX6_1),.din(w_dff_A_ePi6SFEE7_1),.clk(gclk));
	jdff dff_A_N7RiwQhL7_1(.dout(w_dff_A_ePi6SFEE7_1),.din(w_dff_A_N7RiwQhL7_1),.clk(gclk));
	jdff dff_A_Vael7ZcZ0_1(.dout(w_dff_A_N7RiwQhL7_1),.din(w_dff_A_Vael7ZcZ0_1),.clk(gclk));
	jdff dff_A_Qw9v7Yie2_1(.dout(w_G228gat_3[1]),.din(w_dff_A_Qw9v7Yie2_1),.clk(gclk));
	jdff dff_B_sKPLjkxx7_1(.din(n278),.dout(w_dff_B_sKPLjkxx7_1),.clk(gclk));
	jdff dff_B_zvKx1LYf9_1(.din(w_dff_B_sKPLjkxx7_1),.dout(w_dff_B_zvKx1LYf9_1),.clk(gclk));
	jdff dff_B_QquYyicl0_1(.din(w_dff_B_zvKx1LYf9_1),.dout(w_dff_B_QquYyicl0_1),.clk(gclk));
	jdff dff_B_dDHrJEG72_1(.din(w_dff_B_QquYyicl0_1),.dout(w_dff_B_dDHrJEG72_1),.clk(gclk));
	jdff dff_B_aisV8IiX3_1(.din(w_dff_B_dDHrJEG72_1),.dout(w_dff_B_aisV8IiX3_1),.clk(gclk));
	jdff dff_B_P64uaEJY4_1(.din(n279),.dout(w_dff_B_P64uaEJY4_1),.clk(gclk));
	jdff dff_B_OdOP9BaB7_0(.din(n280),.dout(w_dff_B_OdOP9BaB7_0),.clk(gclk));
	jdff dff_B_o5XWamel1_0(.din(w_dff_B_OdOP9BaB7_0),.dout(w_dff_B_o5XWamel1_0),.clk(gclk));
	jdff dff_B_TKok4g8s0_0(.din(w_dff_B_o5XWamel1_0),.dout(w_dff_B_TKok4g8s0_0),.clk(gclk));
	jdff dff_B_EckWqqYc5_0(.din(w_dff_B_TKok4g8s0_0),.dout(w_dff_B_EckWqqYc5_0),.clk(gclk));
	jdff dff_A_6ghpfoia9_0(.dout(w_G219gat_3[0]),.din(w_dff_A_6ghpfoia9_0),.clk(gclk));
	jdff dff_A_JzkKiM653_0(.dout(w_dff_A_6ghpfoia9_0),.din(w_dff_A_JzkKiM653_0),.clk(gclk));
	jdff dff_A_ShCjBaep4_0(.dout(w_dff_A_JzkKiM653_0),.din(w_dff_A_ShCjBaep4_0),.clk(gclk));
	jdff dff_A_hkrrthH71_1(.dout(w_G219gat_3[1]),.din(w_dff_A_hkrrthH71_1),.clk(gclk));
	jdff dff_A_GPFa31IZ2_1(.dout(w_dff_A_hkrrthH71_1),.din(w_dff_A_GPFa31IZ2_1),.clk(gclk));
	jdff dff_A_DmJiZkl84_1(.dout(w_dff_A_GPFa31IZ2_1),.din(w_dff_A_DmJiZkl84_1),.clk(gclk));
	jdff dff_A_ljdrSe2b7_1(.dout(w_dff_A_DmJiZkl84_1),.din(w_dff_A_ljdrSe2b7_1),.clk(gclk));
	jdff dff_A_u2etzkMM4_1(.dout(w_dff_A_ljdrSe2b7_1),.din(w_dff_A_u2etzkMM4_1),.clk(gclk));
	jdff dff_B_ip1O69zR9_1(.din(n268),.dout(w_dff_B_ip1O69zR9_1),.clk(gclk));
	jdff dff_B_NF73eS3m0_0(.din(n276),.dout(w_dff_B_NF73eS3m0_0),.clk(gclk));
	jdff dff_B_FgjDBKvU8_0(.din(w_dff_B_NF73eS3m0_0),.dout(w_dff_B_FgjDBKvU8_0),.clk(gclk));
	jdff dff_B_pcuzcSUF9_0(.din(w_dff_B_FgjDBKvU8_0),.dout(w_dff_B_pcuzcSUF9_0),.clk(gclk));
	jdff dff_B_guoqX5rk6_0(.din(w_dff_B_pcuzcSUF9_0),.dout(w_dff_B_guoqX5rk6_0),.clk(gclk));
	jdff dff_B_L9INqjsN8_1(.din(n274),.dout(w_dff_B_L9INqjsN8_1),.clk(gclk));
	jdff dff_B_ZTZ7NpMe5_1(.din(w_dff_B_L9INqjsN8_1),.dout(w_dff_B_ZTZ7NpMe5_1),.clk(gclk));
	jdff dff_B_oFAamp7l3_1(.din(w_dff_B_ZTZ7NpMe5_1),.dout(w_dff_B_oFAamp7l3_1),.clk(gclk));
	jdff dff_B_6FXB3G1w8_1(.din(w_dff_B_oFAamp7l3_1),.dout(w_dff_B_6FXB3G1w8_1),.clk(gclk));
	jdff dff_B_tbSerfKW1_1(.din(n269),.dout(w_dff_B_tbSerfKW1_1),.clk(gclk));
	jdff dff_B_x36CsGqm2_1(.din(w_dff_B_tbSerfKW1_1),.dout(w_dff_B_x36CsGqm2_1),.clk(gclk));
	jdff dff_B_lBCbBLRQ2_1(.din(w_dff_B_x36CsGqm2_1),.dout(w_dff_B_lBCbBLRQ2_1),.clk(gclk));
	jdff dff_B_hb7M47we2_1(.din(w_dff_B_lBCbBLRQ2_1),.dout(w_dff_B_hb7M47we2_1),.clk(gclk));
	jdff dff_B_xIvQHfp88_1(.din(w_dff_B_hb7M47we2_1),.dout(w_dff_B_xIvQHfp88_1),.clk(gclk));
	jdff dff_B_BpUY3SjG5_1(.din(w_dff_B_xIvQHfp88_1),.dout(w_dff_B_BpUY3SjG5_1),.clk(gclk));
	jdff dff_B_CcvYoYiK1_1(.din(w_dff_B_BpUY3SjG5_1),.dout(w_dff_B_CcvYoYiK1_1),.clk(gclk));
	jdff dff_B_doc87SNp3_1(.din(w_dff_B_CcvYoYiK1_1),.dout(w_dff_B_doc87SNp3_1),.clk(gclk));
	jdff dff_B_oHF4b3lP0_0(.din(n271),.dout(w_dff_B_oHF4b3lP0_0),.clk(gclk));
	jdff dff_B_8RYN9yIv4_0(.din(w_dff_B_oHF4b3lP0_0),.dout(w_dff_B_8RYN9yIv4_0),.clk(gclk));
	jdff dff_B_6cfMoPDX4_0(.din(w_dff_B_8RYN9yIv4_0),.dout(w_dff_B_6cfMoPDX4_0),.clk(gclk));
	jdff dff_B_fds7y00t6_0(.din(w_dff_B_6cfMoPDX4_0),.dout(w_dff_B_fds7y00t6_0),.clk(gclk));
	jdff dff_B_NDQPL4Cb3_0(.din(w_dff_B_fds7y00t6_0),.dout(w_dff_B_NDQPL4Cb3_0),.clk(gclk));
	jdff dff_B_MwAU5TSD8_0(.din(w_dff_B_NDQPL4Cb3_0),.dout(w_dff_B_MwAU5TSD8_0),.clk(gclk));
	jdff dff_A_G4FIs4pM6_1(.dout(w_n267_0[1]),.din(w_dff_A_G4FIs4pM6_1),.clk(gclk));
	jdff dff_A_766102Ba8_1(.dout(w_dff_A_G4FIs4pM6_1),.din(w_dff_A_766102Ba8_1),.clk(gclk));
	jdff dff_A_szlXohlj8_1(.dout(w_dff_A_766102Ba8_1),.din(w_dff_A_szlXohlj8_1),.clk(gclk));
	jdff dff_A_em7gfIqr1_1(.dout(w_dff_A_szlXohlj8_1),.din(w_dff_A_em7gfIqr1_1),.clk(gclk));
	jdff dff_A_oIwOpkCN4_1(.dout(w_dff_A_em7gfIqr1_1),.din(w_dff_A_oIwOpkCN4_1),.clk(gclk));
	jdff dff_B_q38OqGB28_1(.din(n296),.dout(w_dff_B_q38OqGB28_1),.clk(gclk));
	jdff dff_B_dkizGsDs2_1(.din(w_dff_B_q38OqGB28_1),.dout(w_dff_B_dkizGsDs2_1),.clk(gclk));
	jdff dff_B_sBXG36rQ5_1(.din(w_dff_B_dkizGsDs2_1),.dout(w_dff_B_sBXG36rQ5_1),.clk(gclk));
	jdff dff_B_iNv189Yf9_1(.din(n297),.dout(w_dff_B_iNv189Yf9_1),.clk(gclk));
	jdff dff_B_otlZuYIa1_0(.din(n298),.dout(w_dff_B_otlZuYIa1_0),.clk(gclk));
	jdff dff_B_kH9ZOFXQ2_0(.din(w_dff_B_otlZuYIa1_0),.dout(w_dff_B_kH9ZOFXQ2_0),.clk(gclk));
	jdff dff_B_ndu5LyJR1_1(.din(n286),.dout(w_dff_B_ndu5LyJR1_1),.clk(gclk));
	jdff dff_B_DTIFOlka2_0(.din(n294),.dout(w_dff_B_DTIFOlka2_0),.clk(gclk));
	jdff dff_B_ezlAstUf3_0(.din(w_dff_B_DTIFOlka2_0),.dout(w_dff_B_ezlAstUf3_0),.clk(gclk));
	jdff dff_B_Zwr92fFJ9_0(.din(w_dff_B_ezlAstUf3_0),.dout(w_dff_B_Zwr92fFJ9_0),.clk(gclk));
	jdff dff_B_hXPlE1Gb5_0(.din(w_dff_B_Zwr92fFJ9_0),.dout(w_dff_B_hXPlE1Gb5_0),.clk(gclk));
	jdff dff_B_MCIkRQmJ4_0(.din(n293),.dout(w_dff_B_MCIkRQmJ4_0),.clk(gclk));
	jdff dff_B_83HV8bV64_0(.din(w_dff_B_MCIkRQmJ4_0),.dout(w_dff_B_83HV8bV64_0),.clk(gclk));
	jdff dff_B_i2P4lSKr4_0(.din(w_dff_B_83HV8bV64_0),.dout(w_dff_B_i2P4lSKr4_0),.clk(gclk));
	jdff dff_B_MyHsY2ym2_0(.din(w_dff_B_i2P4lSKr4_0),.dout(w_dff_B_MyHsY2ym2_0),.clk(gclk));
	jdff dff_B_0kDBjHJ52_1(.din(n287),.dout(w_dff_B_0kDBjHJ52_1),.clk(gclk));
	jdff dff_B_OUn71ubv4_1(.din(w_dff_B_0kDBjHJ52_1),.dout(w_dff_B_OUn71ubv4_1),.clk(gclk));
	jdff dff_B_bYnvctjA7_1(.din(w_dff_B_OUn71ubv4_1),.dout(w_dff_B_bYnvctjA7_1),.clk(gclk));
	jdff dff_B_Cad6sX8N2_1(.din(w_dff_B_bYnvctjA7_1),.dout(w_dff_B_Cad6sX8N2_1),.clk(gclk));
	jdff dff_B_G8BxU8L91_1(.din(w_dff_B_Cad6sX8N2_1),.dout(w_dff_B_G8BxU8L91_1),.clk(gclk));
	jdff dff_B_HyOFN1pt4_1(.din(w_dff_B_G8BxU8L91_1),.dout(w_dff_B_HyOFN1pt4_1),.clk(gclk));
	jdff dff_B_x0l3AsoL5_1(.din(w_dff_B_HyOFN1pt4_1),.dout(w_dff_B_x0l3AsoL5_1),.clk(gclk));
	jdff dff_B_vvj0HpDe2_1(.din(w_dff_B_x0l3AsoL5_1),.dout(w_dff_B_vvj0HpDe2_1),.clk(gclk));
	jdff dff_B_ckZOUTVT5_0(.din(n289),.dout(w_dff_B_ckZOUTVT5_0),.clk(gclk));
	jdff dff_B_VZfyjC3l4_0(.din(w_dff_B_ckZOUTVT5_0),.dout(w_dff_B_VZfyjC3l4_0),.clk(gclk));
	jdff dff_B_bHfCrVa15_0(.din(w_dff_B_VZfyjC3l4_0),.dout(w_dff_B_bHfCrVa15_0),.clk(gclk));
	jdff dff_B_vTOh8UrP3_0(.din(w_dff_B_bHfCrVa15_0),.dout(w_dff_B_vTOh8UrP3_0),.clk(gclk));
	jdff dff_B_BNahH4ob8_0(.din(w_dff_B_vTOh8UrP3_0),.dout(w_dff_B_BNahH4ob8_0),.clk(gclk));
	jdff dff_B_FRm0f71R6_0(.din(w_dff_B_BNahH4ob8_0),.dout(w_dff_B_FRm0f71R6_0),.clk(gclk));
	jdff dff_A_z66bwLQm1_1(.dout(w_n285_0[1]),.din(w_dff_A_z66bwLQm1_1),.clk(gclk));
	jdff dff_A_FUPxMvZA0_1(.dout(w_dff_A_z66bwLQm1_1),.din(w_dff_A_FUPxMvZA0_1),.clk(gclk));
	jdff dff_A_2sd0l6IR0_1(.dout(w_dff_A_FUPxMvZA0_1),.din(w_dff_A_2sd0l6IR0_1),.clk(gclk));
	jdff dff_B_GlXyYwwF9_1(.din(n312),.dout(w_dff_B_GlXyYwwF9_1),.clk(gclk));
	jdff dff_B_O50J3Kuq4_1(.din(w_dff_B_GlXyYwwF9_1),.dout(w_dff_B_O50J3Kuq4_1),.clk(gclk));
	jdff dff_B_xhdjv0j25_1(.din(w_dff_B_O50J3Kuq4_1),.dout(w_dff_B_xhdjv0j25_1),.clk(gclk));
	jdff dff_B_T3bizIL53_1(.din(w_dff_B_xhdjv0j25_1),.dout(w_dff_B_T3bizIL53_1),.clk(gclk));
	jdff dff_B_6o2QfV8Y8_1(.din(w_dff_B_T3bizIL53_1),.dout(w_dff_B_6o2QfV8Y8_1),.clk(gclk));
	jdff dff_B_OnAOBO4L8_1(.din(w_dff_B_6o2QfV8Y8_1),.dout(w_dff_B_OnAOBO4L8_1),.clk(gclk));
	jdff dff_B_WzVg6u1J8_1(.din(w_dff_B_OnAOBO4L8_1),.dout(w_dff_B_WzVg6u1J8_1),.clk(gclk));
	jdff dff_B_fQrFZnXJ4_1(.din(w_dff_B_WzVg6u1J8_1),.dout(w_dff_B_fQrFZnXJ4_1),.clk(gclk));
	jdff dff_B_sijGcggi2_1(.din(w_dff_B_fQrFZnXJ4_1),.dout(w_dff_B_sijGcggi2_1),.clk(gclk));
	jdff dff_B_So5b2yCD8_1(.din(w_dff_B_sijGcggi2_1),.dout(w_dff_B_So5b2yCD8_1),.clk(gclk));
	jdff dff_B_UC0JnjnF7_1(.din(w_dff_B_So5b2yCD8_1),.dout(w_dff_B_UC0JnjnF7_1),.clk(gclk));
	jdff dff_B_3I2iOSIa8_1(.din(w_dff_B_UC0JnjnF7_1),.dout(w_dff_B_3I2iOSIa8_1),.clk(gclk));
	jdff dff_B_uiLMbmCC7_1(.din(w_dff_B_3I2iOSIa8_1),.dout(w_dff_B_uiLMbmCC7_1),.clk(gclk));
	jdff dff_B_2qo0lXRl2_1(.din(w_dff_B_uiLMbmCC7_1),.dout(w_dff_B_2qo0lXRl2_1),.clk(gclk));
	jdff dff_B_YPDy7Iun2_1(.din(w_dff_B_2qo0lXRl2_1),.dout(w_dff_B_YPDy7Iun2_1),.clk(gclk));
	jdff dff_B_nSMC28Oa8_1(.din(n313),.dout(w_dff_B_nSMC28Oa8_1),.clk(gclk));
	jdff dff_B_xy6Fhd6t4_1(.din(w_dff_B_nSMC28Oa8_1),.dout(w_dff_B_xy6Fhd6t4_1),.clk(gclk));
	jdff dff_B_EsqRNlVT9_1(.din(w_dff_B_xy6Fhd6t4_1),.dout(w_dff_B_EsqRNlVT9_1),.clk(gclk));
	jdff dff_B_FI15eL6y1_1(.din(w_dff_B_EsqRNlVT9_1),.dout(w_dff_B_FI15eL6y1_1),.clk(gclk));
	jdff dff_B_yfNz41jq9_1(.din(w_dff_B_FI15eL6y1_1),.dout(w_dff_B_yfNz41jq9_1),.clk(gclk));
	jdff dff_B_CDwawG0x0_1(.din(w_dff_B_yfNz41jq9_1),.dout(w_dff_B_CDwawG0x0_1),.clk(gclk));
	jdff dff_B_Kak8VqjB7_1(.din(w_dff_B_CDwawG0x0_1),.dout(w_dff_B_Kak8VqjB7_1),.clk(gclk));
	jdff dff_B_jvMGe37M4_1(.din(w_dff_B_Kak8VqjB7_1),.dout(w_dff_B_jvMGe37M4_1),.clk(gclk));
	jdff dff_B_QNnKLkjF5_1(.din(w_dff_B_jvMGe37M4_1),.dout(w_dff_B_QNnKLkjF5_1),.clk(gclk));
	jdff dff_B_Jrd7GfwQ2_1(.din(w_dff_B_QNnKLkjF5_1),.dout(w_dff_B_Jrd7GfwQ2_1),.clk(gclk));
	jdff dff_B_NxdZk2vU0_1(.din(w_dff_B_Jrd7GfwQ2_1),.dout(w_dff_B_NxdZk2vU0_1),.clk(gclk));
	jdff dff_B_9ML7OhUv7_1(.din(w_dff_B_NxdZk2vU0_1),.dout(w_dff_B_9ML7OhUv7_1),.clk(gclk));
	jdff dff_B_Or1qyz1f0_1(.din(w_dff_B_9ML7OhUv7_1),.dout(w_dff_B_Or1qyz1f0_1),.clk(gclk));
	jdff dff_B_t1cU3XPa1_1(.din(w_dff_B_Or1qyz1f0_1),.dout(w_dff_B_t1cU3XPa1_1),.clk(gclk));
	jdff dff_A_xa2Lgavg6_0(.dout(w_G159gat_1[0]),.din(w_dff_A_xa2Lgavg6_0),.clk(gclk));
	jdff dff_A_kGFG3yZG0_0(.dout(w_dff_A_xa2Lgavg6_0),.din(w_dff_A_kGFG3yZG0_0),.clk(gclk));
	jdff dff_A_PO5kjd967_0(.dout(w_dff_A_kGFG3yZG0_0),.din(w_dff_A_PO5kjd967_0),.clk(gclk));
	jdff dff_A_fLCaUrrJ5_0(.dout(w_dff_A_PO5kjd967_0),.din(w_dff_A_fLCaUrrJ5_0),.clk(gclk));
	jdff dff_A_9ShXdnnB2_0(.dout(w_dff_A_fLCaUrrJ5_0),.din(w_dff_A_9ShXdnnB2_0),.clk(gclk));
	jdff dff_A_IitPTuNO5_0(.dout(w_dff_A_9ShXdnnB2_0),.din(w_dff_A_IitPTuNO5_0),.clk(gclk));
	jdff dff_A_n88HvGkE6_0(.dout(w_dff_A_IitPTuNO5_0),.din(w_dff_A_n88HvGkE6_0),.clk(gclk));
	jdff dff_A_J7UmDh821_0(.dout(w_dff_A_n88HvGkE6_0),.din(w_dff_A_J7UmDh821_0),.clk(gclk));
	jdff dff_A_VPQapodH2_0(.dout(w_dff_A_J7UmDh821_0),.din(w_dff_A_VPQapodH2_0),.clk(gclk));
	jdff dff_A_FaO2ZNUX8_1(.dout(w_G159gat_1[1]),.din(w_dff_A_FaO2ZNUX8_1),.clk(gclk));
	jdff dff_A_atznSj4f2_1(.dout(w_dff_A_FaO2ZNUX8_1),.din(w_dff_A_atznSj4f2_1),.clk(gclk));
	jdff dff_A_LveJbCk61_1(.dout(w_dff_A_atznSj4f2_1),.din(w_dff_A_LveJbCk61_1),.clk(gclk));
	jdff dff_A_10HSazra1_1(.dout(w_dff_A_LveJbCk61_1),.din(w_dff_A_10HSazra1_1),.clk(gclk));
	jdff dff_A_FOzdQjo31_1(.dout(w_dff_A_10HSazra1_1),.din(w_dff_A_FOzdQjo31_1),.clk(gclk));
	jdff dff_A_XE1efOH42_1(.dout(w_dff_A_FOzdQjo31_1),.din(w_dff_A_XE1efOH42_1),.clk(gclk));
	jdff dff_A_QMoXbwDy4_1(.dout(w_dff_A_XE1efOH42_1),.din(w_dff_A_QMoXbwDy4_1),.clk(gclk));
	jdff dff_A_YLv8NwLR8_1(.dout(w_dff_A_QMoXbwDy4_1),.din(w_dff_A_YLv8NwLR8_1),.clk(gclk));
	jdff dff_A_uXT30LP58_1(.dout(w_dff_A_YLv8NwLR8_1),.din(w_dff_A_uXT30LP58_1),.clk(gclk));
	jdff dff_B_DrWmOQ3G4_1(.din(n358),.dout(w_dff_B_DrWmOQ3G4_1),.clk(gclk));
	jdff dff_B_SKllqSYH9_1(.din(w_dff_B_DrWmOQ3G4_1),.dout(w_dff_B_SKllqSYH9_1),.clk(gclk));
	jdff dff_B_m1586m9L8_0(.din(n371),.dout(w_dff_B_m1586m9L8_0),.clk(gclk));
	jdff dff_B_bLv1pV2j0_0(.din(w_dff_B_m1586m9L8_0),.dout(w_dff_B_bLv1pV2j0_0),.clk(gclk));
	jdff dff_B_93XyzLj32_0(.din(w_dff_B_bLv1pV2j0_0),.dout(w_dff_B_93XyzLj32_0),.clk(gclk));
	jdff dff_B_ctxjP86f9_0(.din(w_dff_B_93XyzLj32_0),.dout(w_dff_B_ctxjP86f9_0),.clk(gclk));
	jdff dff_B_VpIXfvx32_0(.din(w_dff_B_ctxjP86f9_0),.dout(w_dff_B_VpIXfvx32_0),.clk(gclk));
	jdff dff_B_0GLwW4iA8_0(.din(w_dff_B_VpIXfvx32_0),.dout(w_dff_B_0GLwW4iA8_0),.clk(gclk));
	jdff dff_B_Yk3VSakW1_0(.din(w_dff_B_0GLwW4iA8_0),.dout(w_dff_B_Yk3VSakW1_0),.clk(gclk));
	jdff dff_B_UDCLH5u87_0(.din(w_dff_B_Yk3VSakW1_0),.dout(w_dff_B_UDCLH5u87_0),.clk(gclk));
	jdff dff_B_jrM5SpFM8_0(.din(w_dff_B_UDCLH5u87_0),.dout(w_dff_B_jrM5SpFM8_0),.clk(gclk));
	jdff dff_B_T6ij8MWk3_0(.din(n369),.dout(w_dff_B_T6ij8MWk3_0),.clk(gclk));
	jdff dff_B_lq8hkTeu3_0(.din(w_dff_B_T6ij8MWk3_0),.dout(w_dff_B_lq8hkTeu3_0),.clk(gclk));
	jdff dff_B_orXl8P786_0(.din(w_dff_B_lq8hkTeu3_0),.dout(w_dff_B_orXl8P786_0),.clk(gclk));
	jdff dff_B_wSRGaJsQ8_0(.din(w_dff_B_orXl8P786_0),.dout(w_dff_B_wSRGaJsQ8_0),.clk(gclk));
	jdff dff_B_kHaLqff29_1(.din(n367),.dout(w_dff_B_kHaLqff29_1),.clk(gclk));
	jdff dff_B_pRwP6pur1_1(.din(w_dff_B_kHaLqff29_1),.dout(w_dff_B_pRwP6pur1_1),.clk(gclk));
	jdff dff_B_MjAmgKrD6_1(.din(w_dff_B_pRwP6pur1_1),.dout(w_dff_B_MjAmgKrD6_1),.clk(gclk));
	jdff dff_B_q1deCKrm8_1(.din(w_dff_B_MjAmgKrD6_1),.dout(w_dff_B_q1deCKrm8_1),.clk(gclk));
	jdff dff_A_2HqWG7O22_0(.dout(w_G246gat_2[0]),.din(w_dff_A_2HqWG7O22_0),.clk(gclk));
	jdff dff_A_kFtHrzAs3_0(.dout(w_dff_A_2HqWG7O22_0),.din(w_dff_A_kFtHrzAs3_0),.clk(gclk));
	jdff dff_A_Gn4qwCi11_0(.dout(w_dff_A_kFtHrzAs3_0),.din(w_dff_A_Gn4qwCi11_0),.clk(gclk));
	jdff dff_A_yYwnJvjr0_0(.dout(w_dff_A_Gn4qwCi11_0),.din(w_dff_A_yYwnJvjr0_0),.clk(gclk));
	jdff dff_A_DZFSmrXP2_0(.dout(w_dff_A_yYwnJvjr0_0),.din(w_dff_A_DZFSmrXP2_0),.clk(gclk));
	jdff dff_A_bdFVGDSr6_0(.dout(w_dff_A_DZFSmrXP2_0),.din(w_dff_A_bdFVGDSr6_0),.clk(gclk));
	jdff dff_A_5hhDTQ4c6_0(.dout(w_dff_A_bdFVGDSr6_0),.din(w_dff_A_5hhDTQ4c6_0),.clk(gclk));
	jdff dff_A_aSHbGEry9_0(.dout(w_dff_A_5hhDTQ4c6_0),.din(w_dff_A_aSHbGEry9_0),.clk(gclk));
	jdff dff_A_L8CM89wd5_0(.dout(w_G237gat_2[0]),.din(w_dff_A_L8CM89wd5_0),.clk(gclk));
	jdff dff_A_2mFXpMH17_0(.dout(w_dff_A_L8CM89wd5_0),.din(w_dff_A_2mFXpMH17_0),.clk(gclk));
	jdff dff_A_SL4FOWtT3_0(.dout(w_dff_A_2mFXpMH17_0),.din(w_dff_A_SL4FOWtT3_0),.clk(gclk));
	jdff dff_A_ftrUmz822_0(.dout(w_dff_A_SL4FOWtT3_0),.din(w_dff_A_ftrUmz822_0),.clk(gclk));
	jdff dff_A_SFjHUcDx2_0(.dout(w_dff_A_ftrUmz822_0),.din(w_dff_A_SFjHUcDx2_0),.clk(gclk));
	jdff dff_A_nkTGWDF62_0(.dout(w_dff_A_SFjHUcDx2_0),.din(w_dff_A_nkTGWDF62_0),.clk(gclk));
	jdff dff_A_b0gMc3W59_0(.dout(w_dff_A_nkTGWDF62_0),.din(w_dff_A_b0gMc3W59_0),.clk(gclk));
	jdff dff_A_eIovaeni1_0(.dout(w_dff_A_b0gMc3W59_0),.din(w_dff_A_eIovaeni1_0),.clk(gclk));
	jdff dff_A_TfdjTBKt4_0(.dout(w_dff_A_eIovaeni1_0),.din(w_dff_A_TfdjTBKt4_0),.clk(gclk));
	jdff dff_A_NMD8Frsu5_0(.dout(w_dff_A_TfdjTBKt4_0),.din(w_dff_A_NMD8Frsu5_0),.clk(gclk));
	jdff dff_A_dfJLx5UD0_0(.dout(w_G228gat_2[0]),.din(w_dff_A_dfJLx5UD0_0),.clk(gclk));
	jdff dff_A_dl7XLRC63_0(.dout(w_dff_A_dfJLx5UD0_0),.din(w_dff_A_dl7XLRC63_0),.clk(gclk));
	jdff dff_A_OGL0MYyQ1_0(.dout(w_dff_A_dl7XLRC63_0),.din(w_dff_A_OGL0MYyQ1_0),.clk(gclk));
	jdff dff_A_5xc0eiyF9_0(.dout(w_dff_A_OGL0MYyQ1_0),.din(w_dff_A_5xc0eiyF9_0),.clk(gclk));
	jdff dff_A_ZoeQule85_0(.dout(w_dff_A_5xc0eiyF9_0),.din(w_dff_A_ZoeQule85_0),.clk(gclk));
	jdff dff_A_ZNMvC3Ml1_0(.dout(w_dff_A_ZoeQule85_0),.din(w_dff_A_ZNMvC3Ml1_0),.clk(gclk));
	jdff dff_A_H1ADnFNM4_0(.dout(w_dff_A_ZNMvC3Ml1_0),.din(w_dff_A_H1ADnFNM4_0),.clk(gclk));
	jdff dff_A_RJJIUzRJ7_0(.dout(w_dff_A_H1ADnFNM4_0),.din(w_dff_A_RJJIUzRJ7_0),.clk(gclk));
	jdff dff_A_qXgjvMms3_0(.dout(w_dff_A_RJJIUzRJ7_0),.din(w_dff_A_qXgjvMms3_0),.clk(gclk));
	jdff dff_A_cLdcIYs66_0(.dout(w_dff_A_qXgjvMms3_0),.din(w_dff_A_cLdcIYs66_0),.clk(gclk));
	jdff dff_B_Aq2UPSvS2_1(.din(n356),.dout(w_dff_B_Aq2UPSvS2_1),.clk(gclk));
	jdff dff_B_YuDzUN6G6_1(.din(w_dff_B_Aq2UPSvS2_1),.dout(w_dff_B_YuDzUN6G6_1),.clk(gclk));
	jdff dff_B_fBJRcelf6_1(.din(w_dff_B_YuDzUN6G6_1),.dout(w_dff_B_fBJRcelf6_1),.clk(gclk));
	jdff dff_B_W4KZWh1j7_1(.din(w_dff_B_fBJRcelf6_1),.dout(w_dff_B_W4KZWh1j7_1),.clk(gclk));
	jdff dff_B_shyw5PxS2_1(.din(w_dff_B_W4KZWh1j7_1),.dout(w_dff_B_shyw5PxS2_1),.clk(gclk));
	jdff dff_B_euqnkUns6_1(.din(w_dff_B_shyw5PxS2_1),.dout(w_dff_B_euqnkUns6_1),.clk(gclk));
	jdff dff_B_SLBiKYnm0_1(.din(w_dff_B_euqnkUns6_1),.dout(w_dff_B_SLBiKYnm0_1),.clk(gclk));
	jdff dff_B_6IKmdFBU2_1(.din(w_dff_B_SLBiKYnm0_1),.dout(w_dff_B_6IKmdFBU2_1),.clk(gclk));
	jdff dff_A_4bpxj24S7_0(.dout(w_G219gat_2[0]),.din(w_dff_A_4bpxj24S7_0),.clk(gclk));
	jdff dff_A_p5mQNXnX6_0(.dout(w_dff_A_4bpxj24S7_0),.din(w_dff_A_p5mQNXnX6_0),.clk(gclk));
	jdff dff_A_rufeLn5R4_0(.dout(w_dff_A_p5mQNXnX6_0),.din(w_dff_A_rufeLn5R4_0),.clk(gclk));
	jdff dff_A_Qtn3LZ9u7_0(.dout(w_dff_A_rufeLn5R4_0),.din(w_dff_A_Qtn3LZ9u7_0),.clk(gclk));
	jdff dff_A_5bL57tID5_0(.dout(w_dff_A_Qtn3LZ9u7_0),.din(w_dff_A_5bL57tID5_0),.clk(gclk));
	jdff dff_A_cu6TzZTx5_1(.dout(w_G219gat_2[1]),.din(w_dff_A_cu6TzZTx5_1),.clk(gclk));
	jdff dff_A_khgA3j7b9_1(.dout(w_dff_A_cu6TzZTx5_1),.din(w_dff_A_khgA3j7b9_1),.clk(gclk));
	jdff dff_A_fcPCOdj53_1(.dout(w_dff_A_khgA3j7b9_1),.din(w_dff_A_fcPCOdj53_1),.clk(gclk));
	jdff dff_A_zr0Rae5B3_1(.dout(w_dff_A_fcPCOdj53_1),.din(w_dff_A_zr0Rae5B3_1),.clk(gclk));
	jdff dff_A_wAl3WvJh8_1(.dout(w_dff_A_zr0Rae5B3_1),.din(w_dff_A_wAl3WvJh8_1),.clk(gclk));
	jdff dff_A_bEu2IV3Q4_0(.dout(w_n355_0[0]),.din(w_dff_A_bEu2IV3Q4_0),.clk(gclk));
	jdff dff_A_LtHueLH54_0(.dout(w_dff_A_bEu2IV3Q4_0),.din(w_dff_A_LtHueLH54_0),.clk(gclk));
	jdff dff_A_uiMiqTwk7_0(.dout(w_dff_A_LtHueLH54_0),.din(w_dff_A_uiMiqTwk7_0),.clk(gclk));
	jdff dff_A_hxyWqPOB8_0(.dout(w_dff_A_uiMiqTwk7_0),.din(w_dff_A_hxyWqPOB8_0),.clk(gclk));
	jdff dff_A_7eLuDSf10_0(.dout(w_dff_A_hxyWqPOB8_0),.din(w_dff_A_7eLuDSf10_0),.clk(gclk));
	jdff dff_A_Qb8ZzWj45_0(.dout(w_dff_A_7eLuDSf10_0),.din(w_dff_A_Qb8ZzWj45_0),.clk(gclk));
	jdff dff_A_92DFYHGG1_0(.dout(w_dff_A_Qb8ZzWj45_0),.din(w_dff_A_92DFYHGG1_0),.clk(gclk));
	jdff dff_A_50mAV60x7_0(.dout(w_dff_A_92DFYHGG1_0),.din(w_dff_A_50mAV60x7_0),.clk(gclk));
	jdff dff_A_xHyMAU8u8_0(.dout(w_dff_A_50mAV60x7_0),.din(w_dff_A_xHyMAU8u8_0),.clk(gclk));
	jdff dff_A_FJFDQy9s7_0(.dout(w_dff_A_xHyMAU8u8_0),.din(w_dff_A_FJFDQy9s7_0),.clk(gclk));
	jdff dff_B_SXDplQRF6_1(.din(n383),.dout(w_dff_B_SXDplQRF6_1),.clk(gclk));
	jdff dff_B_1eSM8wuX0_1(.din(w_dff_B_SXDplQRF6_1),.dout(w_dff_B_1eSM8wuX0_1),.clk(gclk));
	jdff dff_B_ZKtxgBCx1_1(.din(w_dff_B_1eSM8wuX0_1),.dout(w_dff_B_ZKtxgBCx1_1),.clk(gclk));
	jdff dff_B_ZPMoxhe70_1(.din(w_dff_B_ZKtxgBCx1_1),.dout(w_dff_B_ZPMoxhe70_1),.clk(gclk));
	jdff dff_B_jASMbCkU1_1(.din(w_dff_B_ZPMoxhe70_1),.dout(w_dff_B_jASMbCkU1_1),.clk(gclk));
	jdff dff_B_q4sDnhd28_1(.din(w_dff_B_jASMbCkU1_1),.dout(w_dff_B_q4sDnhd28_1),.clk(gclk));
	jdff dff_B_qnyZVeN43_1(.din(w_dff_B_q4sDnhd28_1),.dout(w_dff_B_qnyZVeN43_1),.clk(gclk));
	jdff dff_B_RhbtftjB8_1(.din(w_dff_B_qnyZVeN43_1),.dout(w_dff_B_RhbtftjB8_1),.clk(gclk));
	jdff dff_B_WJy5GkCG8_1(.din(w_dff_B_RhbtftjB8_1),.dout(w_dff_B_WJy5GkCG8_1),.clk(gclk));
	jdff dff_B_jf9djXIB7_1(.din(w_dff_B_WJy5GkCG8_1),.dout(w_dff_B_jf9djXIB7_1),.clk(gclk));
	jdff dff_B_5osexZ1Z7_1(.din(w_dff_B_jf9djXIB7_1),.dout(w_dff_B_5osexZ1Z7_1),.clk(gclk));
	jdff dff_B_TMtZInnr4_1(.din(w_dff_B_5osexZ1Z7_1),.dout(w_dff_B_TMtZInnr4_1),.clk(gclk));
	jdff dff_B_Eiyg7v3H6_1(.din(w_dff_B_TMtZInnr4_1),.dout(w_dff_B_Eiyg7v3H6_1),.clk(gclk));
	jdff dff_B_L92F2ZAH0_1(.din(n384),.dout(w_dff_B_L92F2ZAH0_1),.clk(gclk));
	jdff dff_B_jZOQOToS4_0(.din(n396),.dout(w_dff_B_jZOQOToS4_0),.clk(gclk));
	jdff dff_B_1GT3auXp9_0(.din(w_dff_B_jZOQOToS4_0),.dout(w_dff_B_1GT3auXp9_0),.clk(gclk));
	jdff dff_B_AkeX8Jwn1_0(.din(w_dff_B_1GT3auXp9_0),.dout(w_dff_B_AkeX8Jwn1_0),.clk(gclk));
	jdff dff_B_6e3ZrFcL9_0(.din(w_dff_B_AkeX8Jwn1_0),.dout(w_dff_B_6e3ZrFcL9_0),.clk(gclk));
	jdff dff_B_GcvQsw8u4_0(.din(w_dff_B_6e3ZrFcL9_0),.dout(w_dff_B_GcvQsw8u4_0),.clk(gclk));
	jdff dff_B_JC9M4Qdx4_0(.din(w_dff_B_GcvQsw8u4_0),.dout(w_dff_B_JC9M4Qdx4_0),.clk(gclk));
	jdff dff_B_5Hfh4XDf6_0(.din(w_dff_B_JC9M4Qdx4_0),.dout(w_dff_B_5Hfh4XDf6_0),.clk(gclk));
	jdff dff_B_1mMqJSg65_0(.din(w_dff_B_5Hfh4XDf6_0),.dout(w_dff_B_1mMqJSg65_0),.clk(gclk));
	jdff dff_B_ufGA5QdL5_0(.din(w_dff_B_1mMqJSg65_0),.dout(w_dff_B_ufGA5QdL5_0),.clk(gclk));
	jdff dff_B_9cY5hey30_0(.din(w_dff_B_ufGA5QdL5_0),.dout(w_dff_B_9cY5hey30_0),.clk(gclk));
	jdff dff_B_W8k17x5l3_0(.din(w_dff_B_9cY5hey30_0),.dout(w_dff_B_W8k17x5l3_0),.clk(gclk));
	jdff dff_B_CvMGc4DV2_0(.din(w_dff_B_W8k17x5l3_0),.dout(w_dff_B_CvMGc4DV2_0),.clk(gclk));
	jdff dff_B_zAgfXo5z3_0(.din(w_dff_B_CvMGc4DV2_0),.dout(w_dff_B_zAgfXo5z3_0),.clk(gclk));
	jdff dff_B_NYJdjsi79_1(.din(n385),.dout(w_dff_B_NYJdjsi79_1),.clk(gclk));
	jdff dff_B_njk6QFK41_1(.din(w_dff_B_NYJdjsi79_1),.dout(w_dff_B_njk6QFK41_1),.clk(gclk));
	jdff dff_B_rmPoUPLP4_1(.din(w_dff_B_njk6QFK41_1),.dout(w_dff_B_rmPoUPLP4_1),.clk(gclk));
	jdff dff_B_timix9rN1_1(.din(w_dff_B_rmPoUPLP4_1),.dout(w_dff_B_timix9rN1_1),.clk(gclk));
	jdff dff_B_mrW6U2kI1_1(.din(w_dff_B_timix9rN1_1),.dout(w_dff_B_mrW6U2kI1_1),.clk(gclk));
	jdff dff_B_YdvDzPAu6_1(.din(w_dff_B_mrW6U2kI1_1),.dout(w_dff_B_YdvDzPAu6_1),.clk(gclk));
	jdff dff_B_tvnE0rJr4_1(.din(w_dff_B_YdvDzPAu6_1),.dout(w_dff_B_tvnE0rJr4_1),.clk(gclk));
	jdff dff_B_tU4ZQYkN7_1(.din(w_dff_B_tvnE0rJr4_1),.dout(w_dff_B_tU4ZQYkN7_1),.clk(gclk));
	jdff dff_B_nExStRYp5_1(.din(w_dff_B_tU4ZQYkN7_1),.dout(w_dff_B_nExStRYp5_1),.clk(gclk));
	jdff dff_B_CpYOMRyJ5_1(.din(w_dff_B_nExStRYp5_1),.dout(w_dff_B_CpYOMRyJ5_1),.clk(gclk));
	jdff dff_B_63BKISQi8_1(.din(w_dff_B_CpYOMRyJ5_1),.dout(w_dff_B_63BKISQi8_1),.clk(gclk));
	jdff dff_B_a428seju5_1(.din(w_dff_B_63BKISQi8_1),.dout(w_dff_B_a428seju5_1),.clk(gclk));
	jdff dff_B_hMkxnIK09_1(.din(n386),.dout(w_dff_B_hMkxnIK09_1),.clk(gclk));
	jdff dff_B_bCycd5jY6_1(.din(w_dff_B_hMkxnIK09_1),.dout(w_dff_B_bCycd5jY6_1),.clk(gclk));
	jdff dff_B_oAspcJrA0_1(.din(w_dff_B_bCycd5jY6_1),.dout(w_dff_B_oAspcJrA0_1),.clk(gclk));
	jdff dff_B_BPa9AnFI5_1(.din(w_dff_B_oAspcJrA0_1),.dout(w_dff_B_BPa9AnFI5_1),.clk(gclk));
	jdff dff_B_G5PVtizS6_1(.din(w_dff_B_BPa9AnFI5_1),.dout(w_dff_B_G5PVtizS6_1),.clk(gclk));
	jdff dff_B_AdIRQnOQ6_1(.din(w_dff_B_G5PVtizS6_1),.dout(w_dff_B_AdIRQnOQ6_1),.clk(gclk));
	jdff dff_B_3ao02iZo0_1(.din(w_dff_B_AdIRQnOQ6_1),.dout(w_dff_B_3ao02iZo0_1),.clk(gclk));
	jdff dff_B_vv7mdAgE4_1(.din(w_dff_B_3ao02iZo0_1),.dout(w_dff_B_vv7mdAgE4_1),.clk(gclk));
	jdff dff_B_zEVtMg1H1_1(.din(w_dff_B_vv7mdAgE4_1),.dout(w_dff_B_zEVtMg1H1_1),.clk(gclk));
	jdff dff_B_dFp1mONK0_1(.din(w_dff_B_zEVtMg1H1_1),.dout(w_dff_B_dFp1mONK0_1),.clk(gclk));
	jdff dff_B_Bo7oQoJK8_1(.din(w_dff_B_dFp1mONK0_1),.dout(w_dff_B_Bo7oQoJK8_1),.clk(gclk));
	jdff dff_A_Z22eqk216_1(.dout(w_n321_0[1]),.din(w_dff_A_Z22eqk216_1),.clk(gclk));
	jdff dff_A_jiCiVtNY1_1(.dout(w_dff_A_Z22eqk216_1),.din(w_dff_A_jiCiVtNY1_1),.clk(gclk));
	jdff dff_A_NoLqKbR40_1(.dout(w_dff_A_jiCiVtNY1_1),.din(w_dff_A_NoLqKbR40_1),.clk(gclk));
	jdff dff_A_j2w1C8PV1_1(.dout(w_dff_A_NoLqKbR40_1),.din(w_dff_A_j2w1C8PV1_1),.clk(gclk));
	jdff dff_A_OEV2ulpJ1_1(.dout(w_dff_A_j2w1C8PV1_1),.din(w_dff_A_OEV2ulpJ1_1),.clk(gclk));
	jdff dff_A_4lxNdACi7_1(.dout(w_dff_A_OEV2ulpJ1_1),.din(w_dff_A_4lxNdACi7_1),.clk(gclk));
	jdff dff_A_hPY5Y3Tl6_1(.dout(w_dff_A_4lxNdACi7_1),.din(w_dff_A_hPY5Y3Tl6_1),.clk(gclk));
	jdff dff_A_XpHyiiBG8_1(.dout(w_dff_A_hPY5Y3Tl6_1),.din(w_dff_A_XpHyiiBG8_1),.clk(gclk));
	jdff dff_A_7qAWTxjC0_1(.dout(w_dff_A_XpHyiiBG8_1),.din(w_dff_A_7qAWTxjC0_1),.clk(gclk));
	jdff dff_A_lq6Ms2402_1(.dout(w_dff_A_7qAWTxjC0_1),.din(w_dff_A_lq6Ms2402_1),.clk(gclk));
	jdff dff_A_c55AXmE41_1(.dout(w_dff_A_lq6Ms2402_1),.din(w_dff_A_c55AXmE41_1),.clk(gclk));
	jdff dff_A_axQuh9PX7_1(.dout(w_dff_A_c55AXmE41_1),.din(w_dff_A_axQuh9PX7_1),.clk(gclk));
	jdff dff_A_KbNxnfNW8_1(.dout(w_n320_0[1]),.din(w_dff_A_KbNxnfNW8_1),.clk(gclk));
	jdff dff_A_Dbzozypn5_1(.dout(w_dff_A_KbNxnfNW8_1),.din(w_dff_A_Dbzozypn5_1),.clk(gclk));
	jdff dff_A_EHVMy5Wb4_1(.dout(w_dff_A_Dbzozypn5_1),.din(w_dff_A_EHVMy5Wb4_1),.clk(gclk));
	jdff dff_A_BfUMS4cX4_1(.dout(w_dff_A_EHVMy5Wb4_1),.din(w_dff_A_BfUMS4cX4_1),.clk(gclk));
	jdff dff_A_yVJlEyFT5_1(.dout(w_dff_A_BfUMS4cX4_1),.din(w_dff_A_yVJlEyFT5_1),.clk(gclk));
	jdff dff_A_Ej67evNU6_1(.dout(w_dff_A_yVJlEyFT5_1),.din(w_dff_A_Ej67evNU6_1),.clk(gclk));
	jdff dff_A_Yzu5lBv14_1(.dout(w_dff_A_Ej67evNU6_1),.din(w_dff_A_Yzu5lBv14_1),.clk(gclk));
	jdff dff_A_OdjLpzgq4_1(.dout(w_dff_A_Yzu5lBv14_1),.din(w_dff_A_OdjLpzgq4_1),.clk(gclk));
	jdff dff_A_WllzbeKy3_1(.dout(w_dff_A_OdjLpzgq4_1),.din(w_dff_A_WllzbeKy3_1),.clk(gclk));
	jdff dff_A_VEBjHC828_1(.dout(w_dff_A_WllzbeKy3_1),.din(w_dff_A_VEBjHC828_1),.clk(gclk));
	jdff dff_A_cKccF6vN3_1(.dout(w_dff_A_VEBjHC828_1),.din(w_dff_A_cKccF6vN3_1),.clk(gclk));
	jdff dff_A_Dhk20cVU2_1(.dout(w_dff_A_cKccF6vN3_1),.din(w_dff_A_Dhk20cVU2_1),.clk(gclk));
	jdff dff_A_40zSHeLb7_1(.dout(w_dff_A_Dhk20cVU2_1),.din(w_dff_A_40zSHeLb7_1),.clk(gclk));
	jdff dff_A_JfZmhdgi8_0(.dout(w_G165gat_1[0]),.din(w_dff_A_JfZmhdgi8_0),.clk(gclk));
	jdff dff_A_FnqWhfS72_0(.dout(w_dff_A_JfZmhdgi8_0),.din(w_dff_A_FnqWhfS72_0),.clk(gclk));
	jdff dff_A_aYvGGn4P1_0(.dout(w_dff_A_FnqWhfS72_0),.din(w_dff_A_aYvGGn4P1_0),.clk(gclk));
	jdff dff_A_N9KhBuqq0_0(.dout(w_dff_A_aYvGGn4P1_0),.din(w_dff_A_N9KhBuqq0_0),.clk(gclk));
	jdff dff_A_7umzxTUl5_0(.dout(w_dff_A_N9KhBuqq0_0),.din(w_dff_A_7umzxTUl5_0),.clk(gclk));
	jdff dff_A_9ymrjDGK8_0(.dout(w_dff_A_7umzxTUl5_0),.din(w_dff_A_9ymrjDGK8_0),.clk(gclk));
	jdff dff_A_NrX0Px4Y5_0(.dout(w_dff_A_9ymrjDGK8_0),.din(w_dff_A_NrX0Px4Y5_0),.clk(gclk));
	jdff dff_A_aBmZ5SFr4_0(.dout(w_dff_A_NrX0Px4Y5_0),.din(w_dff_A_aBmZ5SFr4_0),.clk(gclk));
	jdff dff_A_8DVrXGV59_1(.dout(w_G165gat_1[1]),.din(w_dff_A_8DVrXGV59_1),.clk(gclk));
	jdff dff_A_3089IQFR8_1(.dout(w_dff_A_8DVrXGV59_1),.din(w_dff_A_3089IQFR8_1),.clk(gclk));
	jdff dff_A_I3MyPCLg6_1(.dout(w_dff_A_3089IQFR8_1),.din(w_dff_A_I3MyPCLg6_1),.clk(gclk));
	jdff dff_A_1Maour7D0_1(.dout(w_dff_A_I3MyPCLg6_1),.din(w_dff_A_1Maour7D0_1),.clk(gclk));
	jdff dff_A_gutcIJ8Z5_1(.dout(w_dff_A_1Maour7D0_1),.din(w_dff_A_gutcIJ8Z5_1),.clk(gclk));
	jdff dff_A_s4h5kpji8_1(.dout(w_dff_A_gutcIJ8Z5_1),.din(w_dff_A_s4h5kpji8_1),.clk(gclk));
	jdff dff_A_rxVNaLEr1_1(.dout(w_dff_A_s4h5kpji8_1),.din(w_dff_A_rxVNaLEr1_1),.clk(gclk));
	jdff dff_A_20PT5cV23_1(.dout(w_dff_A_rxVNaLEr1_1),.din(w_dff_A_20PT5cV23_1),.clk(gclk));
	jdff dff_B_JdO4DSjG8_1(.din(n376),.dout(w_dff_B_JdO4DSjG8_1),.clk(gclk));
	jdff dff_B_JSqBN6F18_0(.din(n381),.dout(w_dff_B_JSqBN6F18_0),.clk(gclk));
	jdff dff_B_vMeloIfP0_0(.din(w_dff_B_JSqBN6F18_0),.dout(w_dff_B_vMeloIfP0_0),.clk(gclk));
	jdff dff_B_u6fypIpY3_0(.din(n379),.dout(w_dff_B_u6fypIpY3_0),.clk(gclk));
	jdff dff_B_RFArZE4m9_0(.din(w_dff_B_u6fypIpY3_0),.dout(w_dff_B_RFArZE4m9_0),.clk(gclk));
	jdff dff_B_aZLpfzCF1_0(.din(w_dff_B_RFArZE4m9_0),.dout(w_dff_B_aZLpfzCF1_0),.clk(gclk));
	jdff dff_B_cePgMkB80_0(.din(w_dff_B_aZLpfzCF1_0),.dout(w_dff_B_cePgMkB80_0),.clk(gclk));
	jdff dff_B_jLU6SnWW2_0(.din(w_dff_B_cePgMkB80_0),.dout(w_dff_B_jLU6SnWW2_0),.clk(gclk));
	jdff dff_B_2DfuLQwR6_0(.din(w_dff_B_jLU6SnWW2_0),.dout(w_dff_B_2DfuLQwR6_0),.clk(gclk));
	jdff dff_B_mwbqMMFu7_0(.din(w_dff_B_2DfuLQwR6_0),.dout(w_dff_B_mwbqMMFu7_0),.clk(gclk));
	jdff dff_B_0NpV4Yn56_0(.din(w_dff_B_mwbqMMFu7_0),.dout(w_dff_B_0NpV4Yn56_0),.clk(gclk));
	jdff dff_B_jkVBsAco1_0(.din(w_dff_B_0NpV4Yn56_0),.dout(w_dff_B_jkVBsAco1_0),.clk(gclk));
	jdff dff_B_lOKYu5SG3_0(.din(w_dff_B_jkVBsAco1_0),.dout(w_dff_B_lOKYu5SG3_0),.clk(gclk));
	jdff dff_A_k0Uhqvpj9_1(.dout(w_n377_0[1]),.din(w_dff_A_k0Uhqvpj9_1),.clk(gclk));
	jdff dff_A_wv7Ex7Qj9_1(.dout(w_dff_A_k0Uhqvpj9_1),.din(w_dff_A_wv7Ex7Qj9_1),.clk(gclk));
	jdff dff_A_k1HBqoWs4_1(.dout(w_dff_A_wv7Ex7Qj9_1),.din(w_dff_A_k1HBqoWs4_1),.clk(gclk));
	jdff dff_A_L5i2ieyX0_1(.dout(w_dff_A_k1HBqoWs4_1),.din(w_dff_A_L5i2ieyX0_1),.clk(gclk));
	jdff dff_A_gq88xnPb3_1(.dout(w_dff_A_L5i2ieyX0_1),.din(w_dff_A_gq88xnPb3_1),.clk(gclk));
	jdff dff_A_8ni1nkcY5_1(.dout(w_dff_A_gq88xnPb3_1),.din(w_dff_A_8ni1nkcY5_1),.clk(gclk));
	jdff dff_A_uoUUwTm15_1(.dout(w_dff_A_8ni1nkcY5_1),.din(w_dff_A_uoUUwTm15_1),.clk(gclk));
	jdff dff_A_iwVYX3Zd3_1(.dout(w_dff_A_uoUUwTm15_1),.din(w_dff_A_iwVYX3Zd3_1),.clk(gclk));
	jdff dff_A_rODvyHfY2_1(.dout(w_dff_A_iwVYX3Zd3_1),.din(w_dff_A_rODvyHfY2_1),.clk(gclk));
	jdff dff_A_RNiQqSRT5_1(.dout(w_dff_A_rODvyHfY2_1),.din(w_dff_A_RNiQqSRT5_1),.clk(gclk));
	jdff dff_A_e7zit8rx5_1(.dout(w_dff_A_RNiQqSRT5_1),.din(w_dff_A_e7zit8rx5_1),.clk(gclk));
	jdff dff_A_SK0o8WK41_1(.dout(w_dff_A_e7zit8rx5_1),.din(w_dff_A_SK0o8WK41_1),.clk(gclk));
	jdff dff_A_beWY4Zs84_1(.dout(w_dff_A_SK0o8WK41_1),.din(w_dff_A_beWY4Zs84_1),.clk(gclk));
	jdff dff_A_kgIBAwiY8_1(.dout(w_dff_A_beWY4Zs84_1),.din(w_dff_A_kgIBAwiY8_1),.clk(gclk));
	jdff dff_B_K8VI0lyJ8_1(.din(n307),.dout(w_dff_B_K8VI0lyJ8_1),.clk(gclk));
	jdff dff_B_6jws5gbv6_0(.din(n309),.dout(w_dff_B_6jws5gbv6_0),.clk(gclk));
	jdff dff_B_IK5EIIq12_0(.din(w_dff_B_6jws5gbv6_0),.dout(w_dff_B_IK5EIIq12_0),.clk(gclk));
	jdff dff_B_UDCo5pPR4_0(.din(w_dff_B_IK5EIIq12_0),.dout(w_dff_B_UDCo5pPR4_0),.clk(gclk));
	jdff dff_B_Hjzc4SbF0_0(.din(w_dff_B_UDCo5pPR4_0),.dout(w_dff_B_Hjzc4SbF0_0),.clk(gclk));
	jdff dff_B_hnrTEviD9_0(.din(w_dff_B_Hjzc4SbF0_0),.dout(w_dff_B_hnrTEviD9_0),.clk(gclk));
	jdff dff_B_dfoDyUwa0_0(.din(w_dff_B_hnrTEviD9_0),.dout(w_dff_B_dfoDyUwa0_0),.clk(gclk));
	jdff dff_B_VTLnXASP2_1(.din(n304),.dout(w_dff_B_VTLnXASP2_1),.clk(gclk));
	jdff dff_A_4Zj3AdZQ4_1(.dout(w_G159gat_0[1]),.din(w_dff_A_4Zj3AdZQ4_1),.clk(gclk));
	jdff dff_A_tAxX9yhZ8_1(.dout(w_dff_A_4Zj3AdZQ4_1),.din(w_dff_A_tAxX9yhZ8_1),.clk(gclk));
	jdff dff_A_vHOFF2l25_1(.dout(w_dff_A_tAxX9yhZ8_1),.din(w_dff_A_vHOFF2l25_1),.clk(gclk));
	jdff dff_A_TbPeTSzs7_1(.dout(w_dff_A_vHOFF2l25_1),.din(w_dff_A_TbPeTSzs7_1),.clk(gclk));
	jdff dff_A_slZFUKBu2_1(.dout(w_dff_A_TbPeTSzs7_1),.din(w_dff_A_slZFUKBu2_1),.clk(gclk));
	jdff dff_A_xEYgw5BB7_1(.dout(w_dff_A_slZFUKBu2_1),.din(w_dff_A_xEYgw5BB7_1),.clk(gclk));
	jdff dff_A_uHBsdGeX2_1(.dout(w_dff_A_xEYgw5BB7_1),.din(w_dff_A_uHBsdGeX2_1),.clk(gclk));
	jdff dff_A_vnmmxkAC4_1(.dout(w_dff_A_uHBsdGeX2_1),.din(w_dff_A_vnmmxkAC4_1),.clk(gclk));
	jdff dff_A_Tf2lEuFd3_1(.dout(w_dff_A_vnmmxkAC4_1),.din(w_dff_A_Tf2lEuFd3_1),.clk(gclk));
	jdff dff_A_kp3nSwIz2_2(.dout(w_G159gat_0[2]),.din(w_dff_A_kp3nSwIz2_2),.clk(gclk));
	jdff dff_A_SeLWDs1C6_2(.dout(w_dff_A_kp3nSwIz2_2),.din(w_dff_A_SeLWDs1C6_2),.clk(gclk));
	jdff dff_A_OEU3F7TX7_2(.dout(w_dff_A_SeLWDs1C6_2),.din(w_dff_A_OEU3F7TX7_2),.clk(gclk));
	jdff dff_A_uo7l20Uw7_2(.dout(w_dff_A_OEU3F7TX7_2),.din(w_dff_A_uo7l20Uw7_2),.clk(gclk));
	jdff dff_A_8bO2taWJ8_2(.dout(w_dff_A_uo7l20Uw7_2),.din(w_dff_A_8bO2taWJ8_2),.clk(gclk));
	jdff dff_A_PHUy7fEB4_2(.dout(w_dff_A_8bO2taWJ8_2),.din(w_dff_A_PHUy7fEB4_2),.clk(gclk));
	jdff dff_A_ITrY2ZIz0_2(.dout(w_dff_A_PHUy7fEB4_2),.din(w_dff_A_ITrY2ZIz0_2),.clk(gclk));
	jdff dff_A_omNB1vwN6_2(.dout(w_dff_A_ITrY2ZIz0_2),.din(w_dff_A_omNB1vwN6_2),.clk(gclk));
	jdff dff_A_uPQS5i6i4_2(.dout(w_dff_A_omNB1vwN6_2),.din(w_dff_A_uPQS5i6i4_2),.clk(gclk));
	jdff dff_A_k1ee7xNV9_2(.dout(w_dff_A_uPQS5i6i4_2),.din(w_dff_A_k1ee7xNV9_2),.clk(gclk));
	jdff dff_A_R0RX7xce5_2(.dout(w_dff_A_k1ee7xNV9_2),.din(w_dff_A_R0RX7xce5_2),.clk(gclk));
	jdff dff_B_eIirSXnc6_1(.din(n410),.dout(w_dff_B_eIirSXnc6_1),.clk(gclk));
	jdff dff_B_Ky1FXVhY4_1(.din(w_dff_B_eIirSXnc6_1),.dout(w_dff_B_Ky1FXVhY4_1),.clk(gclk));
	jdff dff_B_eZTVX8EQ6_1(.din(w_dff_B_Ky1FXVhY4_1),.dout(w_dff_B_eZTVX8EQ6_1),.clk(gclk));
	jdff dff_B_XAbEllva5_1(.din(w_dff_B_eZTVX8EQ6_1),.dout(w_dff_B_XAbEllva5_1),.clk(gclk));
	jdff dff_B_uJkrmF8P6_1(.din(w_dff_B_XAbEllva5_1),.dout(w_dff_B_uJkrmF8P6_1),.clk(gclk));
	jdff dff_B_roZd3Z9n4_1(.din(w_dff_B_uJkrmF8P6_1),.dout(w_dff_B_roZd3Z9n4_1),.clk(gclk));
	jdff dff_B_ycumxEgu4_1(.din(w_dff_B_roZd3Z9n4_1),.dout(w_dff_B_ycumxEgu4_1),.clk(gclk));
	jdff dff_B_O4OyMdAz7_1(.din(w_dff_B_ycumxEgu4_1),.dout(w_dff_B_O4OyMdAz7_1),.clk(gclk));
	jdff dff_B_qlpMLfen2_1(.din(w_dff_B_O4OyMdAz7_1),.dout(w_dff_B_qlpMLfen2_1),.clk(gclk));
	jdff dff_B_X5uVtMo40_1(.din(w_dff_B_qlpMLfen2_1),.dout(w_dff_B_X5uVtMo40_1),.clk(gclk));
	jdff dff_B_qpsPCDeK3_1(.din(w_dff_B_X5uVtMo40_1),.dout(w_dff_B_qpsPCDeK3_1),.clk(gclk));
	jdff dff_B_2eA68JVH7_1(.din(n411),.dout(w_dff_B_2eA68JVH7_1),.clk(gclk));
	jdff dff_B_8KdJBbll1_0(.din(n412),.dout(w_dff_B_8KdJBbll1_0),.clk(gclk));
	jdff dff_B_jxV3Q3h44_0(.din(w_dff_B_8KdJBbll1_0),.dout(w_dff_B_jxV3Q3h44_0),.clk(gclk));
	jdff dff_B_msdHrvXn1_0(.din(w_dff_B_jxV3Q3h44_0),.dout(w_dff_B_msdHrvXn1_0),.clk(gclk));
	jdff dff_B_pyf8G6p62_0(.din(w_dff_B_msdHrvXn1_0),.dout(w_dff_B_pyf8G6p62_0),.clk(gclk));
	jdff dff_B_qqWdOOx01_0(.din(w_dff_B_pyf8G6p62_0),.dout(w_dff_B_qqWdOOx01_0),.clk(gclk));
	jdff dff_B_WwYmBD714_0(.din(w_dff_B_qqWdOOx01_0),.dout(w_dff_B_WwYmBD714_0),.clk(gclk));
	jdff dff_B_wQwNPLSZ5_0(.din(w_dff_B_WwYmBD714_0),.dout(w_dff_B_wQwNPLSZ5_0),.clk(gclk));
	jdff dff_B_5oGhwwWM8_0(.din(w_dff_B_wQwNPLSZ5_0),.dout(w_dff_B_5oGhwwWM8_0),.clk(gclk));
	jdff dff_B_eq2dpWGH8_0(.din(w_dff_B_5oGhwwWM8_0),.dout(w_dff_B_eq2dpWGH8_0),.clk(gclk));
	jdff dff_B_fOiOfrNH0_0(.din(w_dff_B_eq2dpWGH8_0),.dout(w_dff_B_fOiOfrNH0_0),.clk(gclk));
	jdff dff_B_hzZ3zAfb8_0(.din(w_dff_B_fOiOfrNH0_0),.dout(w_dff_B_hzZ3zAfb8_0),.clk(gclk));
	jdff dff_B_1uRZtwzT1_1(.din(n387),.dout(w_dff_B_1uRZtwzT1_1),.clk(gclk));
	jdff dff_B_MglWwv2W7_1(.din(w_dff_B_1uRZtwzT1_1),.dout(w_dff_B_MglWwv2W7_1),.clk(gclk));
	jdff dff_B_qEwBakl73_1(.din(w_dff_B_MglWwv2W7_1),.dout(w_dff_B_qEwBakl73_1),.clk(gclk));
	jdff dff_B_DnLY0apf9_1(.din(w_dff_B_qEwBakl73_1),.dout(w_dff_B_DnLY0apf9_1),.clk(gclk));
	jdff dff_B_vNEw1tAV8_1(.din(w_dff_B_DnLY0apf9_1),.dout(w_dff_B_vNEw1tAV8_1),.clk(gclk));
	jdff dff_B_8x6CCG9t3_1(.din(w_dff_B_vNEw1tAV8_1),.dout(w_dff_B_8x6CCG9t3_1),.clk(gclk));
	jdff dff_B_19gMOpUe2_1(.din(w_dff_B_8x6CCG9t3_1),.dout(w_dff_B_19gMOpUe2_1),.clk(gclk));
	jdff dff_B_uyb6QbQ87_1(.din(w_dff_B_19gMOpUe2_1),.dout(w_dff_B_uyb6QbQ87_1),.clk(gclk));
	jdff dff_B_paBBHVNr4_1(.din(w_dff_B_uyb6QbQ87_1),.dout(w_dff_B_paBBHVNr4_1),.clk(gclk));
	jdff dff_B_MLzv1ZkU1_1(.din(w_dff_B_paBBHVNr4_1),.dout(w_dff_B_MLzv1ZkU1_1),.clk(gclk));
	jdff dff_B_aEbuJ1zi8_1(.din(n388),.dout(w_dff_B_aEbuJ1zi8_1),.clk(gclk));
	jdff dff_B_rcqBL7af9_1(.din(w_dff_B_aEbuJ1zi8_1),.dout(w_dff_B_rcqBL7af9_1),.clk(gclk));
	jdff dff_B_QQouUaOH4_1(.din(w_dff_B_rcqBL7af9_1),.dout(w_dff_B_QQouUaOH4_1),.clk(gclk));
	jdff dff_B_FNVWj71O0_1(.din(w_dff_B_QQouUaOH4_1),.dout(w_dff_B_FNVWj71O0_1),.clk(gclk));
	jdff dff_B_ZWPs6Pbv2_1(.din(w_dff_B_FNVWj71O0_1),.dout(w_dff_B_ZWPs6Pbv2_1),.clk(gclk));
	jdff dff_B_TWjNr2ld3_1(.din(w_dff_B_ZWPs6Pbv2_1),.dout(w_dff_B_TWjNr2ld3_1),.clk(gclk));
	jdff dff_B_FZd1igRE1_1(.din(w_dff_B_TWjNr2ld3_1),.dout(w_dff_B_FZd1igRE1_1),.clk(gclk));
	jdff dff_B_5ZNWOaTP6_1(.din(w_dff_B_FZd1igRE1_1),.dout(w_dff_B_5ZNWOaTP6_1),.clk(gclk));
	jdff dff_B_8w1OuQ7g3_1(.din(w_dff_B_5ZNWOaTP6_1),.dout(w_dff_B_8w1OuQ7g3_1),.clk(gclk));
	jdff dff_A_engRbXKT4_1(.dout(w_n329_0[1]),.din(w_dff_A_engRbXKT4_1),.clk(gclk));
	jdff dff_A_3oFMPpWl3_1(.dout(w_dff_A_engRbXKT4_1),.din(w_dff_A_3oFMPpWl3_1),.clk(gclk));
	jdff dff_A_znlV3md30_1(.dout(w_dff_A_3oFMPpWl3_1),.din(w_dff_A_znlV3md30_1),.clk(gclk));
	jdff dff_A_5XSnst9T3_1(.dout(w_dff_A_znlV3md30_1),.din(w_dff_A_5XSnst9T3_1),.clk(gclk));
	jdff dff_A_qASWQBJd9_1(.dout(w_dff_A_5XSnst9T3_1),.din(w_dff_A_qASWQBJd9_1),.clk(gclk));
	jdff dff_A_c4XqH9Jq6_1(.dout(w_dff_A_qASWQBJd9_1),.din(w_dff_A_c4XqH9Jq6_1),.clk(gclk));
	jdff dff_A_4p14Z57N8_1(.dout(w_dff_A_c4XqH9Jq6_1),.din(w_dff_A_4p14Z57N8_1),.clk(gclk));
	jdff dff_A_1LyHZ4gi4_1(.dout(w_dff_A_4p14Z57N8_1),.din(w_dff_A_1LyHZ4gi4_1),.clk(gclk));
	jdff dff_A_eXhgisLy9_1(.dout(w_dff_A_1LyHZ4gi4_1),.din(w_dff_A_eXhgisLy9_1),.clk(gclk));
	jdff dff_A_7tkxUkqg0_1(.dout(w_dff_A_eXhgisLy9_1),.din(w_dff_A_7tkxUkqg0_1),.clk(gclk));
	jdff dff_A_wdomqhDh0_1(.dout(w_n328_0[1]),.din(w_dff_A_wdomqhDh0_1),.clk(gclk));
	jdff dff_A_J26MXrAT5_1(.dout(w_dff_A_wdomqhDh0_1),.din(w_dff_A_J26MXrAT5_1),.clk(gclk));
	jdff dff_A_dHegbbFb7_1(.dout(w_dff_A_J26MXrAT5_1),.din(w_dff_A_dHegbbFb7_1),.clk(gclk));
	jdff dff_A_v8NB6jfx4_1(.dout(w_dff_A_dHegbbFb7_1),.din(w_dff_A_v8NB6jfx4_1),.clk(gclk));
	jdff dff_A_U98ulfnE3_1(.dout(w_dff_A_v8NB6jfx4_1),.din(w_dff_A_U98ulfnE3_1),.clk(gclk));
	jdff dff_A_sOiJtSMu0_1(.dout(w_dff_A_U98ulfnE3_1),.din(w_dff_A_sOiJtSMu0_1),.clk(gclk));
	jdff dff_A_my9Nsj4F8_1(.dout(w_dff_A_sOiJtSMu0_1),.din(w_dff_A_my9Nsj4F8_1),.clk(gclk));
	jdff dff_A_h68msO2v9_1(.dout(w_dff_A_my9Nsj4F8_1),.din(w_dff_A_h68msO2v9_1),.clk(gclk));
	jdff dff_A_wzvmsC068_1(.dout(w_dff_A_h68msO2v9_1),.din(w_dff_A_wzvmsC068_1),.clk(gclk));
	jdff dff_A_R1aCiAet8_1(.dout(w_dff_A_wzvmsC068_1),.din(w_dff_A_R1aCiAet8_1),.clk(gclk));
	jdff dff_A_FTobAgMp7_1(.dout(w_dff_A_R1aCiAet8_1),.din(w_dff_A_FTobAgMp7_1),.clk(gclk));
	jdff dff_A_UU9iPBcA4_0(.dout(w_G171gat_1[0]),.din(w_dff_A_UU9iPBcA4_0),.clk(gclk));
	jdff dff_A_9A9lp9Eb4_0(.dout(w_dff_A_UU9iPBcA4_0),.din(w_dff_A_9A9lp9Eb4_0),.clk(gclk));
	jdff dff_A_INzUODqZ4_0(.dout(w_dff_A_9A9lp9Eb4_0),.din(w_dff_A_INzUODqZ4_0),.clk(gclk));
	jdff dff_A_xXRZk73L2_0(.dout(w_dff_A_INzUODqZ4_0),.din(w_dff_A_xXRZk73L2_0),.clk(gclk));
	jdff dff_A_KuLxciOz2_0(.dout(w_dff_A_xXRZk73L2_0),.din(w_dff_A_KuLxciOz2_0),.clk(gclk));
	jdff dff_A_ezwpn8W24_0(.dout(w_dff_A_KuLxciOz2_0),.din(w_dff_A_ezwpn8W24_0),.clk(gclk));
	jdff dff_A_cWtTiz9r3_0(.dout(w_dff_A_ezwpn8W24_0),.din(w_dff_A_cWtTiz9r3_0),.clk(gclk));
	jdff dff_A_Q53lHbmZ0_0(.dout(w_dff_A_cWtTiz9r3_0),.din(w_dff_A_Q53lHbmZ0_0),.clk(gclk));
	jdff dff_A_02D4fnOb6_0(.dout(w_dff_A_Q53lHbmZ0_0),.din(w_dff_A_02D4fnOb6_0),.clk(gclk));
	jdff dff_A_shllhsGN3_1(.dout(w_G171gat_1[1]),.din(w_dff_A_shllhsGN3_1),.clk(gclk));
	jdff dff_A_InB01ckg0_1(.dout(w_dff_A_shllhsGN3_1),.din(w_dff_A_InB01ckg0_1),.clk(gclk));
	jdff dff_A_pKrmJp5H2_1(.dout(w_dff_A_InB01ckg0_1),.din(w_dff_A_pKrmJp5H2_1),.clk(gclk));
	jdff dff_A_9GVTtQD67_1(.dout(w_dff_A_pKrmJp5H2_1),.din(w_dff_A_9GVTtQD67_1),.clk(gclk));
	jdff dff_A_EFqaIDSk5_1(.dout(w_dff_A_9GVTtQD67_1),.din(w_dff_A_EFqaIDSk5_1),.clk(gclk));
	jdff dff_A_n6e7PoKP8_1(.dout(w_dff_A_EFqaIDSk5_1),.din(w_dff_A_n6e7PoKP8_1),.clk(gclk));
	jdff dff_A_pj5cndwv9_1(.dout(w_dff_A_n6e7PoKP8_1),.din(w_dff_A_pj5cndwv9_1),.clk(gclk));
	jdff dff_A_UtSll5fY6_1(.dout(w_dff_A_pj5cndwv9_1),.din(w_dff_A_UtSll5fY6_1),.clk(gclk));
	jdff dff_A_g03eD6ey0_1(.dout(w_dff_A_UtSll5fY6_1),.din(w_dff_A_g03eD6ey0_1),.clk(gclk));
	jdff dff_B_dlwkneye3_1(.din(n403),.dout(w_dff_B_dlwkneye3_1),.clk(gclk));
	jdff dff_B_KIrQzHVz5_0(.din(n408),.dout(w_dff_B_KIrQzHVz5_0),.clk(gclk));
	jdff dff_B_uMvaqNZj5_0(.din(w_dff_B_KIrQzHVz5_0),.dout(w_dff_B_uMvaqNZj5_0),.clk(gclk));
	jdff dff_B_lpsEsrVg7_0(.din(n406),.dout(w_dff_B_lpsEsrVg7_0),.clk(gclk));
	jdff dff_B_agLkgqch1_0(.din(w_dff_B_lpsEsrVg7_0),.dout(w_dff_B_agLkgqch1_0),.clk(gclk));
	jdff dff_B_0ZiPLVHK9_0(.din(w_dff_B_agLkgqch1_0),.dout(w_dff_B_0ZiPLVHK9_0),.clk(gclk));
	jdff dff_B_aBUg2K088_0(.din(w_dff_B_0ZiPLVHK9_0),.dout(w_dff_B_aBUg2K088_0),.clk(gclk));
	jdff dff_B_9hUKfTx27_0(.din(w_dff_B_aBUg2K088_0),.dout(w_dff_B_9hUKfTx27_0),.clk(gclk));
	jdff dff_B_AgCrDA4K5_0(.din(w_dff_B_9hUKfTx27_0),.dout(w_dff_B_AgCrDA4K5_0),.clk(gclk));
	jdff dff_B_dUEFt5038_0(.din(w_dff_B_AgCrDA4K5_0),.dout(w_dff_B_dUEFt5038_0),.clk(gclk));
	jdff dff_B_HLQ7PiTf1_0(.din(w_dff_B_dUEFt5038_0),.dout(w_dff_B_HLQ7PiTf1_0),.clk(gclk));
	jdff dff_B_6GizWAwk6_0(.din(w_dff_B_HLQ7PiTf1_0),.dout(w_dff_B_6GizWAwk6_0),.clk(gclk));
	jdff dff_B_L6Cx6YAe2_0(.din(w_dff_B_6GizWAwk6_0),.dout(w_dff_B_L6Cx6YAe2_0),.clk(gclk));
	jdff dff_A_bOHcy3SC2_1(.dout(w_G91gat_0[1]),.din(w_dff_A_bOHcy3SC2_1),.clk(gclk));
	jdff dff_A_YvldfqGX2_1(.dout(w_dff_A_bOHcy3SC2_1),.din(w_dff_A_YvldfqGX2_1),.clk(gclk));
	jdff dff_A_1tR2bwiQ8_1(.dout(w_dff_A_YvldfqGX2_1),.din(w_dff_A_1tR2bwiQ8_1),.clk(gclk));
	jdff dff_A_roJ5mBDn7_1(.dout(w_dff_A_1tR2bwiQ8_1),.din(w_dff_A_roJ5mBDn7_1),.clk(gclk));
	jdff dff_A_WUrOF5Nu4_1(.dout(w_dff_A_roJ5mBDn7_1),.din(w_dff_A_WUrOF5Nu4_1),.clk(gclk));
	jdff dff_A_oTpOBk6E7_1(.dout(w_dff_A_WUrOF5Nu4_1),.din(w_dff_A_oTpOBk6E7_1),.clk(gclk));
	jdff dff_A_3vOBsTQw1_1(.dout(w_n404_0[1]),.din(w_dff_A_3vOBsTQw1_1),.clk(gclk));
	jdff dff_A_AvNJqJvz7_1(.dout(w_dff_A_3vOBsTQw1_1),.din(w_dff_A_AvNJqJvz7_1),.clk(gclk));
	jdff dff_A_1tKKaC8p3_1(.dout(w_dff_A_AvNJqJvz7_1),.din(w_dff_A_1tKKaC8p3_1),.clk(gclk));
	jdff dff_A_F039WYSQ4_1(.dout(w_dff_A_1tKKaC8p3_1),.din(w_dff_A_F039WYSQ4_1),.clk(gclk));
	jdff dff_A_Bc55XUFv9_1(.dout(w_dff_A_F039WYSQ4_1),.din(w_dff_A_Bc55XUFv9_1),.clk(gclk));
	jdff dff_A_3Fd7i2wB9_1(.dout(w_dff_A_Bc55XUFv9_1),.din(w_dff_A_3Fd7i2wB9_1),.clk(gclk));
	jdff dff_A_Sj0lpnoe4_1(.dout(w_dff_A_3Fd7i2wB9_1),.din(w_dff_A_Sj0lpnoe4_1),.clk(gclk));
	jdff dff_A_FoUjy6Ta5_1(.dout(w_dff_A_Sj0lpnoe4_1),.din(w_dff_A_FoUjy6Ta5_1),.clk(gclk));
	jdff dff_A_ooD3Ukf66_1(.dout(w_dff_A_FoUjy6Ta5_1),.din(w_dff_A_ooD3Ukf66_1),.clk(gclk));
	jdff dff_A_gn18gln43_1(.dout(w_dff_A_ooD3Ukf66_1),.din(w_dff_A_gn18gln43_1),.clk(gclk));
	jdff dff_A_otzWUpkS7_1(.dout(w_dff_A_gn18gln43_1),.din(w_dff_A_otzWUpkS7_1),.clk(gclk));
	jdff dff_A_Ye0keKFV5_1(.dout(w_dff_A_otzWUpkS7_1),.din(w_dff_A_Ye0keKFV5_1),.clk(gclk));
	jdff dff_B_YIE4AI0Q3_0(.din(n317),.dout(w_dff_B_YIE4AI0Q3_0),.clk(gclk));
	jdff dff_B_mLhkwnQJ8_0(.din(n316),.dout(w_dff_B_mLhkwnQJ8_0),.clk(gclk));
	jdff dff_B_ehZpJYeN2_0(.din(w_dff_B_mLhkwnQJ8_0),.dout(w_dff_B_ehZpJYeN2_0),.clk(gclk));
	jdff dff_B_FuEYpuSB1_0(.din(w_dff_B_ehZpJYeN2_0),.dout(w_dff_B_FuEYpuSB1_0),.clk(gclk));
	jdff dff_B_Lvdg5TNC7_0(.din(w_dff_B_FuEYpuSB1_0),.dout(w_dff_B_Lvdg5TNC7_0),.clk(gclk));
	jdff dff_A_V5b14Wph3_0(.dout(w_n306_1[0]),.din(w_dff_A_V5b14Wph3_0),.clk(gclk));
	jdff dff_A_aZ5BSb7c0_0(.dout(w_dff_A_V5b14Wph3_0),.din(w_dff_A_aZ5BSb7c0_0),.clk(gclk));
	jdff dff_A_RSja8HpL9_1(.dout(w_G165gat_0[1]),.din(w_dff_A_RSja8HpL9_1),.clk(gclk));
	jdff dff_A_N6nQcjI13_1(.dout(w_dff_A_RSja8HpL9_1),.din(w_dff_A_N6nQcjI13_1),.clk(gclk));
	jdff dff_A_nP6MPk1y1_1(.dout(w_dff_A_N6nQcjI13_1),.din(w_dff_A_nP6MPk1y1_1),.clk(gclk));
	jdff dff_A_LOCLfv7S9_1(.dout(w_dff_A_nP6MPk1y1_1),.din(w_dff_A_LOCLfv7S9_1),.clk(gclk));
	jdff dff_A_KwU262fS1_1(.dout(w_dff_A_LOCLfv7S9_1),.din(w_dff_A_KwU262fS1_1),.clk(gclk));
	jdff dff_A_9apxVu2V1_1(.dout(w_dff_A_KwU262fS1_1),.din(w_dff_A_9apxVu2V1_1),.clk(gclk));
	jdff dff_A_iZ1Nq6986_1(.dout(w_dff_A_9apxVu2V1_1),.din(w_dff_A_iZ1Nq6986_1),.clk(gclk));
	jdff dff_A_aaz0C0hF6_1(.dout(w_dff_A_iZ1Nq6986_1),.din(w_dff_A_aaz0C0hF6_1),.clk(gclk));
	jdff dff_A_In3Yvowm5_2(.dout(w_G165gat_0[2]),.din(w_dff_A_In3Yvowm5_2),.clk(gclk));
	jdff dff_A_1i6Plmm84_2(.dout(w_dff_A_In3Yvowm5_2),.din(w_dff_A_1i6Plmm84_2),.clk(gclk));
	jdff dff_A_x6FcYThh9_2(.dout(w_dff_A_1i6Plmm84_2),.din(w_dff_A_x6FcYThh9_2),.clk(gclk));
	jdff dff_A_ruisOMEA3_2(.dout(w_dff_A_x6FcYThh9_2),.din(w_dff_A_ruisOMEA3_2),.clk(gclk));
	jdff dff_A_8Yt1i2r50_2(.dout(w_dff_A_ruisOMEA3_2),.din(w_dff_A_8Yt1i2r50_2),.clk(gclk));
	jdff dff_A_046Llune2_2(.dout(w_dff_A_8Yt1i2r50_2),.din(w_dff_A_046Llune2_2),.clk(gclk));
	jdff dff_A_Uv46jueQ6_2(.dout(w_dff_A_046Llune2_2),.din(w_dff_A_Uv46jueQ6_2),.clk(gclk));
	jdff dff_A_f8RbYu1F1_2(.dout(w_dff_A_Uv46jueQ6_2),.din(w_dff_A_f8RbYu1F1_2),.clk(gclk));
	jdff dff_A_UOV4zIC17_2(.dout(w_dff_A_f8RbYu1F1_2),.din(w_dff_A_UOV4zIC17_2),.clk(gclk));
	jdff dff_A_47HpDG880_2(.dout(w_dff_A_UOV4zIC17_2),.din(w_dff_A_47HpDG880_2),.clk(gclk));
	jdff dff_B_zMkHJ0nj7_3(.din(G165gat),.dout(w_dff_B_zMkHJ0nj7_3),.clk(gclk));
	jdff dff_B_vcx3oYgK1_1(.din(n426),.dout(w_dff_B_vcx3oYgK1_1),.clk(gclk));
	jdff dff_B_CnIApL732_1(.din(w_dff_B_vcx3oYgK1_1),.dout(w_dff_B_CnIApL732_1),.clk(gclk));
	jdff dff_B_9yUJyxsw7_1(.din(w_dff_B_CnIApL732_1),.dout(w_dff_B_9yUJyxsw7_1),.clk(gclk));
	jdff dff_B_92diCjO80_1(.din(w_dff_B_9yUJyxsw7_1),.dout(w_dff_B_92diCjO80_1),.clk(gclk));
	jdff dff_B_zhrKKLg55_1(.din(w_dff_B_92diCjO80_1),.dout(w_dff_B_zhrKKLg55_1),.clk(gclk));
	jdff dff_B_rbfxAyFi3_1(.din(w_dff_B_zhrKKLg55_1),.dout(w_dff_B_rbfxAyFi3_1),.clk(gclk));
	jdff dff_B_DdYGjlKf0_1(.din(w_dff_B_rbfxAyFi3_1),.dout(w_dff_B_DdYGjlKf0_1),.clk(gclk));
	jdff dff_B_eBRHz32i5_1(.din(w_dff_B_DdYGjlKf0_1),.dout(w_dff_B_eBRHz32i5_1),.clk(gclk));
	jdff dff_B_TMxMNK401_1(.din(w_dff_B_eBRHz32i5_1),.dout(w_dff_B_TMxMNK401_1),.clk(gclk));
	jdff dff_B_rAKNhPEe8_1(.din(n428),.dout(w_dff_B_rAKNhPEe8_1),.clk(gclk));
	jdff dff_B_QxlXhkmt8_1(.din(n340),.dout(w_dff_B_QxlXhkmt8_1),.clk(gclk));
	jdff dff_B_bhIKsTNy3_1(.din(w_dff_B_QxlXhkmt8_1),.dout(w_dff_B_bhIKsTNy3_1),.clk(gclk));
	jdff dff_B_3kgt0fwD0_1(.din(w_dff_B_bhIKsTNy3_1),.dout(w_dff_B_3kgt0fwD0_1),.clk(gclk));
	jdff dff_B_uIgVnf2l3_1(.din(w_dff_B_3kgt0fwD0_1),.dout(w_dff_B_uIgVnf2l3_1),.clk(gclk));
	jdff dff_B_a38qD3AE2_1(.din(w_dff_B_uIgVnf2l3_1),.dout(w_dff_B_a38qD3AE2_1),.clk(gclk));
	jdff dff_B_LS8NEahk2_1(.din(w_dff_B_a38qD3AE2_1),.dout(w_dff_B_LS8NEahk2_1),.clk(gclk));
	jdff dff_B_RY4ui54r9_1(.din(n344),.dout(w_dff_B_RY4ui54r9_1),.clk(gclk));
	jdff dff_B_xRzrSoIB5_1(.din(w_dff_B_RY4ui54r9_1),.dout(w_dff_B_xRzrSoIB5_1),.clk(gclk));
	jdff dff_B_OlOPpOTr1_1(.din(w_dff_B_xRzrSoIB5_1),.dout(w_dff_B_OlOPpOTr1_1),.clk(gclk));
	jdff dff_B_7OCCR3vq1_1(.din(w_dff_B_OlOPpOTr1_1),.dout(w_dff_B_7OCCR3vq1_1),.clk(gclk));
	jdff dff_B_QKD3aOcz1_1(.din(w_dff_B_7OCCR3vq1_1),.dout(w_dff_B_QKD3aOcz1_1),.clk(gclk));
	jdff dff_B_QdPGDnfW5_0(.din(n171),.dout(w_dff_B_QdPGDnfW5_0),.clk(gclk));
	jdff dff_A_NcwZOuFP5_1(.dout(w_G219gat_1[1]),.din(w_dff_A_NcwZOuFP5_1),.clk(gclk));
	jdff dff_A_dT4pKEOP1_1(.dout(w_dff_A_NcwZOuFP5_1),.din(w_dff_A_dT4pKEOP1_1),.clk(gclk));
	jdff dff_A_QW8NP6Ae8_2(.dout(w_G219gat_1[2]),.din(w_dff_A_QW8NP6Ae8_2),.clk(gclk));
	jdff dff_A_jFvzm0Ak7_2(.dout(w_dff_A_QW8NP6Ae8_2),.din(w_dff_A_jFvzm0Ak7_2),.clk(gclk));
	jdff dff_A_eNJeqv691_2(.dout(w_dff_A_jFvzm0Ak7_2),.din(w_dff_A_eNJeqv691_2),.clk(gclk));
	jdff dff_A_Js3VHItE4_2(.dout(w_dff_A_eNJeqv691_2),.din(w_dff_A_Js3VHItE4_2),.clk(gclk));
	jdff dff_A_GKozbHjS6_0(.dout(w_G219gat_0[0]),.din(w_dff_A_GKozbHjS6_0),.clk(gclk));
	jdff dff_A_q2edVvNo5_0(.dout(w_dff_A_GKozbHjS6_0),.din(w_dff_A_q2edVvNo5_0),.clk(gclk));
	jdff dff_A_dG4J56FL1_0(.dout(w_dff_A_q2edVvNo5_0),.din(w_dff_A_dG4J56FL1_0),.clk(gclk));
	jdff dff_A_JviPyOI71_0(.dout(w_dff_A_dG4J56FL1_0),.din(w_dff_A_JviPyOI71_0),.clk(gclk));
	jdff dff_A_YVufY6Yn4_0(.dout(w_dff_A_JviPyOI71_0),.din(w_dff_A_YVufY6Yn4_0),.clk(gclk));
	jdff dff_A_MWxTom3X1_0(.dout(w_dff_A_YVufY6Yn4_0),.din(w_dff_A_MWxTom3X1_0),.clk(gclk));
	jdff dff_A_9qNzPFPT4_0(.dout(w_dff_A_MWxTom3X1_0),.din(w_dff_A_9qNzPFPT4_0),.clk(gclk));
	jdff dff_A_Ig8XvwYb0_0(.dout(w_dff_A_9qNzPFPT4_0),.din(w_dff_A_Ig8XvwYb0_0),.clk(gclk));
	jdff dff_A_koVGwb1J7_0(.dout(w_dff_A_Ig8XvwYb0_0),.din(w_dff_A_koVGwb1J7_0),.clk(gclk));
	jdff dff_A_LIhv0HB99_1(.dout(w_G219gat_0[1]),.din(w_dff_A_LIhv0HB99_1),.clk(gclk));
	jdff dff_B_Jm7YAUIf8_3(.din(G219gat),.dout(w_dff_B_Jm7YAUIf8_3),.clk(gclk));
	jdff dff_B_VTZ8uKpI5_3(.din(w_dff_B_Jm7YAUIf8_3),.dout(w_dff_B_VTZ8uKpI5_3),.clk(gclk));
	jdff dff_B_q9HzVpiH3_3(.din(w_dff_B_VTZ8uKpI5_3),.dout(w_dff_B_q9HzVpiH3_3),.clk(gclk));
	jdff dff_B_KqeXf7Wc5_3(.din(w_dff_B_q9HzVpiH3_3),.dout(w_dff_B_KqeXf7Wc5_3),.clk(gclk));
	jdff dff_B_HHSiVRuC2_3(.din(w_dff_B_KqeXf7Wc5_3),.dout(w_dff_B_HHSiVRuC2_3),.clk(gclk));
	jdff dff_B_9mmNTlrJ0_3(.din(w_dff_B_HHSiVRuC2_3),.dout(w_dff_B_9mmNTlrJ0_3),.clk(gclk));
	jdff dff_B_q0Ustjpx0_3(.din(w_dff_B_9mmNTlrJ0_3),.dout(w_dff_B_q0Ustjpx0_3),.clk(gclk));
	jdff dff_B_oL5kaV4W9_3(.din(w_dff_B_q0Ustjpx0_3),.dout(w_dff_B_oL5kaV4W9_3),.clk(gclk));
	jdff dff_B_9W7BhV6T4_3(.din(w_dff_B_oL5kaV4W9_3),.dout(w_dff_B_9W7BhV6T4_3),.clk(gclk));
	jdff dff_B_gKD6Sfvu3_3(.din(w_dff_B_9W7BhV6T4_3),.dout(w_dff_B_gKD6Sfvu3_3),.clk(gclk));
	jdff dff_B_DcB3BtP64_3(.din(w_dff_B_gKD6Sfvu3_3),.dout(w_dff_B_DcB3BtP64_3),.clk(gclk));
	jdff dff_B_m5Gj2lRU7_3(.din(w_dff_B_DcB3BtP64_3),.dout(w_dff_B_m5Gj2lRU7_3),.clk(gclk));
	jdff dff_B_1w4VTA2g9_0(.din(n427),.dout(w_dff_B_1w4VTA2g9_0),.clk(gclk));
	jdff dff_B_5fvz4Qhb5_0(.din(w_dff_B_1w4VTA2g9_0),.dout(w_dff_B_5fvz4Qhb5_0),.clk(gclk));
	jdff dff_B_z9sdbC247_0(.din(w_dff_B_5fvz4Qhb5_0),.dout(w_dff_B_z9sdbC247_0),.clk(gclk));
	jdff dff_B_CL48g2ma9_0(.din(w_dff_B_z9sdbC247_0),.dout(w_dff_B_CL48g2ma9_0),.clk(gclk));
	jdff dff_B_dkBEa0IK9_0(.din(w_dff_B_CL48g2ma9_0),.dout(w_dff_B_dkBEa0IK9_0),.clk(gclk));
	jdff dff_B_HDnOkxuC9_0(.din(w_dff_B_dkBEa0IK9_0),.dout(w_dff_B_HDnOkxuC9_0),.clk(gclk));
	jdff dff_B_DTepdAYK3_0(.din(w_dff_B_HDnOkxuC9_0),.dout(w_dff_B_DTepdAYK3_0),.clk(gclk));
	jdff dff_B_T2h4Zyv13_0(.din(w_dff_B_DTepdAYK3_0),.dout(w_dff_B_T2h4Zyv13_0),.clk(gclk));
	jdff dff_B_vuZe0bKa8_0(.din(w_dff_B_T2h4Zyv13_0),.dout(w_dff_B_vuZe0bKa8_0),.clk(gclk));
	jdff dff_B_qtxyYpw43_1(.din(n389),.dout(w_dff_B_qtxyYpw43_1),.clk(gclk));
	jdff dff_B_EDaRfIjO0_1(.din(w_dff_B_qtxyYpw43_1),.dout(w_dff_B_EDaRfIjO0_1),.clk(gclk));
	jdff dff_B_IuNQyzo01_1(.din(w_dff_B_EDaRfIjO0_1),.dout(w_dff_B_IuNQyzo01_1),.clk(gclk));
	jdff dff_B_ThDmAcZc5_1(.din(w_dff_B_IuNQyzo01_1),.dout(w_dff_B_ThDmAcZc5_1),.clk(gclk));
	jdff dff_B_RI333wRp4_1(.din(w_dff_B_ThDmAcZc5_1),.dout(w_dff_B_RI333wRp4_1),.clk(gclk));
	jdff dff_B_5O1U2irJ4_1(.din(w_dff_B_RI333wRp4_1),.dout(w_dff_B_5O1U2irJ4_1),.clk(gclk));
	jdff dff_B_dPoGyPpH7_1(.din(w_dff_B_5O1U2irJ4_1),.dout(w_dff_B_dPoGyPpH7_1),.clk(gclk));
	jdff dff_B_oP1zgrp35_1(.din(w_dff_B_dPoGyPpH7_1),.dout(w_dff_B_oP1zgrp35_1),.clk(gclk));
	jdff dff_B_Msf3FSz51_1(.din(n359),.dout(w_dff_B_Msf3FSz51_1),.clk(gclk));
	jdff dff_B_BCtGabV65_1(.din(w_dff_B_Msf3FSz51_1),.dout(w_dff_B_BCtGabV65_1),.clk(gclk));
	jdff dff_B_D2FAKTIT6_1(.din(w_dff_B_BCtGabV65_1),.dout(w_dff_B_D2FAKTIT6_1),.clk(gclk));
	jdff dff_B_tGstGLdi9_1(.din(w_dff_B_D2FAKTIT6_1),.dout(w_dff_B_tGstGLdi9_1),.clk(gclk));
	jdff dff_B_4NzgPSVU1_1(.din(w_dff_B_tGstGLdi9_1),.dout(w_dff_B_4NzgPSVU1_1),.clk(gclk));
	jdff dff_B_aosymfRH9_1(.din(w_dff_B_4NzgPSVU1_1),.dout(w_dff_B_aosymfRH9_1),.clk(gclk));
	jdff dff_B_niR2iSyj5_1(.din(w_dff_B_aosymfRH9_1),.dout(w_dff_B_niR2iSyj5_1),.clk(gclk));
	jdff dff_B_yqWbuv4n6_1(.din(n252),.dout(w_dff_B_yqWbuv4n6_1),.clk(gclk));
	jdff dff_B_12eFf1aX0_1(.din(w_dff_B_yqWbuv4n6_1),.dout(w_dff_B_12eFf1aX0_1),.clk(gclk));
	jdff dff_B_2noeHm9M2_1(.din(w_dff_B_12eFf1aX0_1),.dout(w_dff_B_2noeHm9M2_1),.clk(gclk));
	jdff dff_B_EFKFLGYk2_1(.din(w_dff_B_2noeHm9M2_1),.dout(w_dff_B_EFKFLGYk2_1),.clk(gclk));
	jdff dff_B_spIMZWyK8_1(.din(w_dff_B_EFKFLGYk2_1),.dout(w_dff_B_spIMZWyK8_1),.clk(gclk));
	jdff dff_B_mCRnWzHO9_1(.din(n253),.dout(w_dff_B_mCRnWzHO9_1),.clk(gclk));
	jdff dff_B_cTamk3c79_1(.din(w_dff_B_mCRnWzHO9_1),.dout(w_dff_B_cTamk3c79_1),.clk(gclk));
	jdff dff_B_XDGuFuiR0_1(.din(w_dff_B_cTamk3c79_1),.dout(w_dff_B_XDGuFuiR0_1),.clk(gclk));
	jdff dff_B_19NGwPN46_1(.din(w_dff_B_XDGuFuiR0_1),.dout(w_dff_B_19NGwPN46_1),.clk(gclk));
	jdff dff_B_y38gfn5x8_1(.din(n254),.dout(w_dff_B_y38gfn5x8_1),.clk(gclk));
	jdff dff_B_oKUvMmsd4_1(.din(w_dff_B_y38gfn5x8_1),.dout(w_dff_B_oKUvMmsd4_1),.clk(gclk));
	jdff dff_B_xrz6Q3Nn9_1(.din(w_dff_B_oKUvMmsd4_1),.dout(w_dff_B_xrz6Q3Nn9_1),.clk(gclk));
	jdff dff_B_mOsoktAu8_1(.din(n255),.dout(w_dff_B_mOsoktAu8_1),.clk(gclk));
	jdff dff_B_v3aEujkO0_1(.din(w_dff_B_mOsoktAu8_1),.dout(w_dff_B_v3aEujkO0_1),.clk(gclk));
	jdff dff_A_UVuRWb7K0_1(.dout(w_n209_0[1]),.din(w_dff_A_UVuRWb7K0_1),.clk(gclk));
	jdff dff_B_CUGOx4Xa8_2(.din(n209),.dout(w_dff_B_CUGOx4Xa8_2),.clk(gclk));
	jdff dff_B_u7wJvy8b2_2(.din(w_dff_B_CUGOx4Xa8_2),.dout(w_dff_B_u7wJvy8b2_2),.clk(gclk));
	jdff dff_B_tNTHa7YL0_2(.din(w_dff_B_u7wJvy8b2_2),.dout(w_dff_B_tNTHa7YL0_2),.clk(gclk));
	jdff dff_B_MMHg49Z23_2(.din(w_dff_B_tNTHa7YL0_2),.dout(w_dff_B_MMHg49Z23_2),.clk(gclk));
	jdff dff_B_xhveRNNy9_2(.din(w_dff_B_MMHg49Z23_2),.dout(w_dff_B_xhveRNNy9_2),.clk(gclk));
	jdff dff_B_VlAAHc3T9_2(.din(w_dff_B_xhveRNNy9_2),.dout(w_dff_B_VlAAHc3T9_2),.clk(gclk));
	jdff dff_B_8LlkZY8y6_2(.din(w_dff_B_VlAAHc3T9_2),.dout(w_dff_B_8LlkZY8y6_2),.clk(gclk));
	jdff dff_B_dDtBeSFw6_2(.din(w_dff_B_8LlkZY8y6_2),.dout(w_dff_B_dDtBeSFw6_2),.clk(gclk));
	jdff dff_B_f1hnKObp1_2(.din(w_dff_B_dDtBeSFw6_2),.dout(w_dff_B_f1hnKObp1_2),.clk(gclk));
	jdff dff_A_DqTnrhIl5_0(.dout(w_G261gat_0[0]),.din(w_dff_A_DqTnrhIl5_0),.clk(gclk));
	jdff dff_A_nZeOoi1Q7_0(.dout(w_dff_A_DqTnrhIl5_0),.din(w_dff_A_nZeOoi1Q7_0),.clk(gclk));
	jdff dff_A_0QlFjbiQ7_0(.dout(w_dff_A_nZeOoi1Q7_0),.din(w_dff_A_0QlFjbiQ7_0),.clk(gclk));
	jdff dff_A_1fi3r4ZL8_0(.dout(w_dff_A_0QlFjbiQ7_0),.din(w_dff_A_1fi3r4ZL8_0),.clk(gclk));
	jdff dff_A_S0v5LtTG4_0(.dout(w_dff_A_1fi3r4ZL8_0),.din(w_dff_A_S0v5LtTG4_0),.clk(gclk));
	jdff dff_A_AH4XdhIQ4_0(.dout(w_dff_A_S0v5LtTG4_0),.din(w_dff_A_AH4XdhIQ4_0),.clk(gclk));
	jdff dff_A_OZxINHqO5_0(.dout(w_dff_A_AH4XdhIQ4_0),.din(w_dff_A_OZxINHqO5_0),.clk(gclk));
	jdff dff_A_8H6jWBfK8_0(.dout(w_dff_A_OZxINHqO5_0),.din(w_dff_A_8H6jWBfK8_0),.clk(gclk));
	jdff dff_A_o5Z5aBps6_0(.dout(w_dff_A_8H6jWBfK8_0),.din(w_dff_A_o5Z5aBps6_0),.clk(gclk));
	jdff dff_A_xvKkIVhB3_0(.dout(w_dff_A_o5Z5aBps6_0),.din(w_dff_A_xvKkIVhB3_0),.clk(gclk));
	jdff dff_A_XHiH6VLY5_2(.dout(w_G261gat_0[2]),.din(w_dff_A_XHiH6VLY5_2),.clk(gclk));
	jdff dff_A_h3xHLoam6_2(.dout(w_dff_A_XHiH6VLY5_2),.din(w_dff_A_h3xHLoam6_2),.clk(gclk));
	jdff dff_A_0ZzOJ9s41_2(.dout(w_dff_A_h3xHLoam6_2),.din(w_dff_A_0ZzOJ9s41_2),.clk(gclk));
	jdff dff_A_OkZcfFI15_2(.dout(w_dff_A_0ZzOJ9s41_2),.din(w_dff_A_OkZcfFI15_2),.clk(gclk));
	jdff dff_A_D94QmB3M0_2(.dout(w_dff_A_OkZcfFI15_2),.din(w_dff_A_D94QmB3M0_2),.clk(gclk));
	jdff dff_A_S3M3fRAn7_2(.dout(w_dff_A_D94QmB3M0_2),.din(w_dff_A_S3M3fRAn7_2),.clk(gclk));
	jdff dff_A_P17HqdxI6_2(.dout(w_dff_A_S3M3fRAn7_2),.din(w_dff_A_P17HqdxI6_2),.clk(gclk));
	jdff dff_A_qEG7kw0c2_2(.dout(w_dff_A_P17HqdxI6_2),.din(w_dff_A_qEG7kw0c2_2),.clk(gclk));
	jdff dff_A_VYUcKGTx5_2(.dout(w_dff_A_qEG7kw0c2_2),.din(w_dff_A_VYUcKGTx5_2),.clk(gclk));
	jdff dff_A_tWLi3I009_2(.dout(w_dff_A_VYUcKGTx5_2),.din(w_dff_A_tWLi3I009_2),.clk(gclk));
	jdff dff_A_BR6IopgH9_0(.dout(w_n242_0[0]),.din(w_dff_A_BR6IopgH9_0),.clk(gclk));
	jdff dff_B_OPiSdhep1_1(.din(n182),.dout(w_dff_B_OPiSdhep1_1),.clk(gclk));
	jdff dff_B_mA4MlP5C4_1(.din(n191),.dout(w_dff_B_mA4MlP5C4_1),.clk(gclk));
	jdff dff_B_x2lpgnGr9_1(.din(w_dff_B_mA4MlP5C4_1),.dout(w_dff_B_x2lpgnGr9_1),.clk(gclk));
	jdff dff_B_6nB9UQd83_1(.din(w_dff_B_x2lpgnGr9_1),.dout(w_dff_B_6nB9UQd83_1),.clk(gclk));
	jdff dff_B_c070VwAL9_1(.din(w_dff_B_6nB9UQd83_1),.dout(w_dff_B_c070VwAL9_1),.clk(gclk));
	jdff dff_B_GOhcr1J55_1(.din(w_dff_B_c070VwAL9_1),.dout(w_dff_B_GOhcr1J55_1),.clk(gclk));
	jdff dff_B_Nj6Fttg42_1(.din(n183),.dout(w_dff_B_Nj6Fttg42_1),.clk(gclk));
	jdff dff_B_tDiisvgf9_1(.din(w_dff_B_Nj6Fttg42_1),.dout(w_dff_B_tDiisvgf9_1),.clk(gclk));
	jdff dff_B_8loXTjO36_1(.din(w_dff_B_tDiisvgf9_1),.dout(w_dff_B_8loXTjO36_1),.clk(gclk));
	jdff dff_B_o6S3j0gd1_1(.din(w_dff_B_8loXTjO36_1),.dout(w_dff_B_o6S3j0gd1_1),.clk(gclk));
	jdff dff_B_28qe7Luv9_1(.din(w_dff_B_o6S3j0gd1_1),.dout(w_dff_B_28qe7Luv9_1),.clk(gclk));
	jdff dff_B_0l3hpL6U6_1(.din(n184),.dout(w_dff_B_0l3hpL6U6_1),.clk(gclk));
	jdff dff_A_2xfzd5o59_1(.dout(w_G126gat_0[1]),.din(w_dff_A_2xfzd5o59_1),.clk(gclk));
	jdff dff_A_pjMlJL7w5_1(.dout(w_dff_A_2xfzd5o59_1),.din(w_dff_A_pjMlJL7w5_1),.clk(gclk));
	jdff dff_A_x2JRJvFm8_1(.dout(w_dff_A_pjMlJL7w5_1),.din(w_dff_A_x2JRJvFm8_1),.clk(gclk));
	jdff dff_A_0BM63biI3_1(.dout(w_dff_A_x2JRJvFm8_1),.din(w_dff_A_0BM63biI3_1),.clk(gclk));
	jdff dff_A_Kd4YlRlz3_1(.dout(w_dff_A_0BM63biI3_1),.din(w_dff_A_Kd4YlRlz3_1),.clk(gclk));
	jdff dff_A_J9u0xkXT3_1(.dout(w_dff_A_Kd4YlRlz3_1),.din(w_dff_A_J9u0xkXT3_1),.clk(gclk));
	jdff dff_B_zfKJ7N7m9_3(.din(n181),.dout(w_dff_B_zfKJ7N7m9_3),.clk(gclk));
	jdff dff_B_SoYIK06C6_3(.din(w_dff_B_zfKJ7N7m9_3),.dout(w_dff_B_SoYIK06C6_3),.clk(gclk));
	jdff dff_B_wlzgIIT85_3(.din(w_dff_B_SoYIK06C6_3),.dout(w_dff_B_wlzgIIT85_3),.clk(gclk));
	jdff dff_B_A0QiUiGi9_3(.din(w_dff_B_wlzgIIT85_3),.dout(w_dff_B_A0QiUiGi9_3),.clk(gclk));
	jdff dff_B_tAww97vC7_3(.din(w_dff_B_A0QiUiGi9_3),.dout(w_dff_B_tAww97vC7_3),.clk(gclk));
	jdff dff_B_AyP8ITd23_3(.din(w_dff_B_tAww97vC7_3),.dout(w_dff_B_AyP8ITd23_3),.clk(gclk));
	jdff dff_B_u8o26h9M9_3(.din(w_dff_B_AyP8ITd23_3),.dout(w_dff_B_u8o26h9M9_3),.clk(gclk));
	jdff dff_B_04yVh3Ik9_3(.din(w_dff_B_u8o26h9M9_3),.dout(w_dff_B_04yVh3Ik9_3),.clk(gclk));
	jdff dff_A_anwux2PY4_1(.dout(w_G201gat_0[1]),.din(w_dff_A_anwux2PY4_1),.clk(gclk));
	jdff dff_A_QCsBnuU61_1(.dout(w_dff_A_anwux2PY4_1),.din(w_dff_A_QCsBnuU61_1),.clk(gclk));
	jdff dff_A_BgmEGnbB8_1(.dout(w_dff_A_QCsBnuU61_1),.din(w_dff_A_BgmEGnbB8_1),.clk(gclk));
	jdff dff_A_78llugOu7_1(.dout(w_dff_A_BgmEGnbB8_1),.din(w_dff_A_78llugOu7_1),.clk(gclk));
	jdff dff_A_red26bU52_1(.dout(w_dff_A_78llugOu7_1),.din(w_dff_A_red26bU52_1),.clk(gclk));
	jdff dff_A_YkBjhwvG7_1(.dout(w_dff_A_red26bU52_1),.din(w_dff_A_YkBjhwvG7_1),.clk(gclk));
	jdff dff_A_a1dYiDs89_1(.dout(w_dff_A_YkBjhwvG7_1),.din(w_dff_A_a1dYiDs89_1),.clk(gclk));
	jdff dff_A_GmaYrDzu7_1(.dout(w_dff_A_a1dYiDs89_1),.din(w_dff_A_GmaYrDzu7_1),.clk(gclk));
	jdff dff_A_ZBaVSZNC1_1(.dout(w_dff_A_GmaYrDzu7_1),.din(w_dff_A_ZBaVSZNC1_1),.clk(gclk));
	jdff dff_A_nDGu6vTd3_1(.dout(w_n241_0[1]),.din(w_dff_A_nDGu6vTd3_1),.clk(gclk));
	jdff dff_A_6uI5kzyr7_1(.dout(w_dff_A_nDGu6vTd3_1),.din(w_dff_A_6uI5kzyr7_1),.clk(gclk));
	jdff dff_A_quB8R3mO5_1(.dout(w_dff_A_6uI5kzyr7_1),.din(w_dff_A_quB8R3mO5_1),.clk(gclk));
	jdff dff_A_W8te3zfr7_1(.dout(w_G195gat_1[1]),.din(w_dff_A_W8te3zfr7_1),.clk(gclk));
	jdff dff_A_UUMNC2K21_1(.dout(w_dff_A_W8te3zfr7_1),.din(w_dff_A_UUMNC2K21_1),.clk(gclk));
	jdff dff_A_1rbhOwR07_1(.dout(w_dff_A_UUMNC2K21_1),.din(w_dff_A_1rbhOwR07_1),.clk(gclk));
	jdff dff_A_8iTJRlCD9_1(.dout(w_dff_A_1rbhOwR07_1),.din(w_dff_A_8iTJRlCD9_1),.clk(gclk));
	jdff dff_A_8IYVivLB2_1(.dout(w_dff_A_8iTJRlCD9_1),.din(w_dff_A_8IYVivLB2_1),.clk(gclk));
	jdff dff_A_bIp7JPaB2_1(.dout(w_dff_A_8IYVivLB2_1),.din(w_dff_A_bIp7JPaB2_1),.clk(gclk));
	jdff dff_A_TS8rg5tl1_1(.dout(w_dff_A_bIp7JPaB2_1),.din(w_dff_A_TS8rg5tl1_1),.clk(gclk));
	jdff dff_A_lU1z5EkX9_1(.dout(w_dff_A_TS8rg5tl1_1),.din(w_dff_A_lU1z5EkX9_1),.clk(gclk));
	jdff dff_A_M72P0FaF0_2(.dout(w_G195gat_1[2]),.din(w_dff_A_M72P0FaF0_2),.clk(gclk));
	jdff dff_A_An7VvAPD4_2(.dout(w_dff_A_M72P0FaF0_2),.din(w_dff_A_An7VvAPD4_2),.clk(gclk));
	jdff dff_A_2D24J6EF4_2(.dout(w_dff_A_An7VvAPD4_2),.din(w_dff_A_2D24J6EF4_2),.clk(gclk));
	jdff dff_A_uOUQTLOU8_2(.dout(w_dff_A_2D24J6EF4_2),.din(w_dff_A_uOUQTLOU8_2),.clk(gclk));
	jdff dff_A_KkbhJVix4_2(.dout(w_dff_A_uOUQTLOU8_2),.din(w_dff_A_KkbhJVix4_2),.clk(gclk));
	jdff dff_A_S69iXiTB7_2(.dout(w_dff_A_KkbhJVix4_2),.din(w_dff_A_S69iXiTB7_2),.clk(gclk));
	jdff dff_A_VeWXXP224_2(.dout(w_dff_A_S69iXiTB7_2),.din(w_dff_A_VeWXXP224_2),.clk(gclk));
	jdff dff_A_C5Xdz3Bg2_2(.dout(w_dff_A_VeWXXP224_2),.din(w_dff_A_C5Xdz3Bg2_2),.clk(gclk));
	jdff dff_A_Qc9qz0su8_1(.dout(w_n240_0[1]),.din(w_dff_A_Qc9qz0su8_1),.clk(gclk));
	jdff dff_A_mTCIWOxs1_1(.dout(w_dff_A_Qc9qz0su8_1),.din(w_dff_A_mTCIWOxs1_1),.clk(gclk));
	jdff dff_A_DybErGmq4_1(.dout(w_dff_A_mTCIWOxs1_1),.din(w_dff_A_DybErGmq4_1),.clk(gclk));
	jdff dff_A_9r8CxF4s7_1(.dout(w_dff_A_DybErGmq4_1),.din(w_dff_A_9r8CxF4s7_1),.clk(gclk));
	jdff dff_A_BTDMx0wS6_0(.dout(w_G121gat_0[0]),.din(w_dff_A_BTDMx0wS6_0),.clk(gclk));
	jdff dff_A_1f5IhjJr9_0(.dout(w_dff_A_BTDMx0wS6_0),.din(w_dff_A_1f5IhjJr9_0),.clk(gclk));
	jdff dff_A_fEVCnXKE6_0(.dout(w_dff_A_1f5IhjJr9_0),.din(w_dff_A_fEVCnXKE6_0),.clk(gclk));
	jdff dff_A_zsvxAFX32_0(.dout(w_dff_A_fEVCnXKE6_0),.din(w_dff_A_zsvxAFX32_0),.clk(gclk));
	jdff dff_A_4DZ0DHiw3_0(.dout(w_dff_A_zsvxAFX32_0),.din(w_dff_A_4DZ0DHiw3_0),.clk(gclk));
	jdff dff_A_FdI0WKCU2_0(.dout(w_dff_A_4DZ0DHiw3_0),.din(w_dff_A_FdI0WKCU2_0),.clk(gclk));
	jdff dff_A_pn8SS0211_0(.dout(w_G195gat_2[0]),.din(w_dff_A_pn8SS0211_0),.clk(gclk));
	jdff dff_A_cBbE321R9_0(.dout(w_dff_A_pn8SS0211_0),.din(w_dff_A_cBbE321R9_0),.clk(gclk));
	jdff dff_A_l7iNudkR1_0(.dout(w_dff_A_cBbE321R9_0),.din(w_dff_A_l7iNudkR1_0),.clk(gclk));
	jdff dff_A_IFC4esab3_0(.dout(w_dff_A_l7iNudkR1_0),.din(w_dff_A_IFC4esab3_0),.clk(gclk));
	jdff dff_A_Jl2E8xC86_0(.dout(w_dff_A_IFC4esab3_0),.din(w_dff_A_Jl2E8xC86_0),.clk(gclk));
	jdff dff_A_pHvtnFbZ5_0(.dout(w_dff_A_Jl2E8xC86_0),.din(w_dff_A_pHvtnFbZ5_0),.clk(gclk));
	jdff dff_A_fSh8t9Nd7_0(.dout(w_dff_A_pHvtnFbZ5_0),.din(w_dff_A_fSh8t9Nd7_0),.clk(gclk));
	jdff dff_A_LuLFkDYT4_0(.dout(w_dff_A_fSh8t9Nd7_0),.din(w_dff_A_LuLFkDYT4_0),.clk(gclk));
	jdff dff_A_e3J1pnr79_2(.dout(w_G195gat_0[2]),.din(w_dff_A_e3J1pnr79_2),.clk(gclk));
	jdff dff_A_T1EEyyyr8_2(.dout(w_dff_A_e3J1pnr79_2),.din(w_dff_A_T1EEyyyr8_2),.clk(gclk));
	jdff dff_A_8WUbxf3m4_2(.dout(w_dff_A_T1EEyyyr8_2),.din(w_dff_A_8WUbxf3m4_2),.clk(gclk));
	jdff dff_A_kKqLSNdp8_2(.dout(w_dff_A_8WUbxf3m4_2),.din(w_dff_A_kKqLSNdp8_2),.clk(gclk));
	jdff dff_A_31DXj4Dq1_1(.dout(w_n235_0[1]),.din(w_dff_A_31DXj4Dq1_1),.clk(gclk));
	jdff dff_A_b6EtOz573_1(.dout(w_dff_A_31DXj4Dq1_1),.din(w_dff_A_b6EtOz573_1),.clk(gclk));
	jdff dff_A_sq5ThnlK4_1(.dout(w_dff_A_b6EtOz573_1),.din(w_dff_A_sq5ThnlK4_1),.clk(gclk));
	jdff dff_A_P8WvbM3b1_1(.dout(w_dff_A_sq5ThnlK4_1),.din(w_dff_A_P8WvbM3b1_1),.clk(gclk));
	jdff dff_A_NQy8YkrC9_1(.dout(w_dff_A_P8WvbM3b1_1),.din(w_dff_A_NQy8YkrC9_1),.clk(gclk));
	jdff dff_A_v2Ylb1H41_1(.dout(w_G189gat_1[1]),.din(w_dff_A_v2Ylb1H41_1),.clk(gclk));
	jdff dff_A_vz9pDDQx5_1(.dout(w_dff_A_v2Ylb1H41_1),.din(w_dff_A_vz9pDDQx5_1),.clk(gclk));
	jdff dff_A_seVjTeaD7_1(.dout(w_dff_A_vz9pDDQx5_1),.din(w_dff_A_seVjTeaD7_1),.clk(gclk));
	jdff dff_A_ocRD18GY1_1(.dout(w_dff_A_seVjTeaD7_1),.din(w_dff_A_ocRD18GY1_1),.clk(gclk));
	jdff dff_A_H5c3FY6G9_1(.dout(w_dff_A_ocRD18GY1_1),.din(w_dff_A_H5c3FY6G9_1),.clk(gclk));
	jdff dff_A_M5arLt3Z5_1(.dout(w_dff_A_H5c3FY6G9_1),.din(w_dff_A_M5arLt3Z5_1),.clk(gclk));
	jdff dff_A_o61HqWLd7_1(.dout(w_dff_A_M5arLt3Z5_1),.din(w_dff_A_o61HqWLd7_1),.clk(gclk));
	jdff dff_A_gaObyY8W5_1(.dout(w_dff_A_o61HqWLd7_1),.din(w_dff_A_gaObyY8W5_1),.clk(gclk));
	jdff dff_A_ld2lwYjb7_2(.dout(w_G189gat_1[2]),.din(w_dff_A_ld2lwYjb7_2),.clk(gclk));
	jdff dff_A_YYBLDlml1_2(.dout(w_dff_A_ld2lwYjb7_2),.din(w_dff_A_YYBLDlml1_2),.clk(gclk));
	jdff dff_A_tYxlxKKx9_2(.dout(w_dff_A_YYBLDlml1_2),.din(w_dff_A_tYxlxKKx9_2),.clk(gclk));
	jdff dff_A_396RtzK68_2(.dout(w_dff_A_tYxlxKKx9_2),.din(w_dff_A_396RtzK68_2),.clk(gclk));
	jdff dff_A_zrFuKfsF3_2(.dout(w_dff_A_396RtzK68_2),.din(w_dff_A_zrFuKfsF3_2),.clk(gclk));
	jdff dff_A_VNL9OsKT4_2(.dout(w_dff_A_zrFuKfsF3_2),.din(w_dff_A_VNL9OsKT4_2),.clk(gclk));
	jdff dff_A_whrbb0aH2_2(.dout(w_dff_A_VNL9OsKT4_2),.din(w_dff_A_whrbb0aH2_2),.clk(gclk));
	jdff dff_A_WSQG2nQG3_2(.dout(w_dff_A_whrbb0aH2_2),.din(w_dff_A_WSQG2nQG3_2),.clk(gclk));
	jdff dff_A_rLOKQHf29_1(.dout(w_n234_0[1]),.din(w_dff_A_rLOKQHf29_1),.clk(gclk));
	jdff dff_A_WGCtSMdN0_1(.dout(w_dff_A_rLOKQHf29_1),.din(w_dff_A_WGCtSMdN0_1),.clk(gclk));
	jdff dff_A_Mv4oLQNj8_1(.dout(w_dff_A_WGCtSMdN0_1),.din(w_dff_A_Mv4oLQNj8_1),.clk(gclk));
	jdff dff_A_Ha0CWY2D6_1(.dout(w_dff_A_Mv4oLQNj8_1),.din(w_dff_A_Ha0CWY2D6_1),.clk(gclk));
	jdff dff_A_mhs3MIuJ4_1(.dout(w_dff_A_Ha0CWY2D6_1),.din(w_dff_A_mhs3MIuJ4_1),.clk(gclk));
	jdff dff_A_iU1DSUeC9_1(.dout(w_dff_A_mhs3MIuJ4_1),.din(w_dff_A_iU1DSUeC9_1),.clk(gclk));
	jdff dff_A_483dyFML3_1(.dout(w_G146gat_0[1]),.din(w_dff_A_483dyFML3_1),.clk(gclk));
	jdff dff_B_ezOcNm4t7_2(.din(G146gat),.dout(w_dff_B_ezOcNm4t7_2),.clk(gclk));
	jdff dff_B_CSmh3Je67_2(.din(w_dff_B_ezOcNm4t7_2),.dout(w_dff_B_CSmh3Je67_2),.clk(gclk));
	jdff dff_B_bYRmQvUm5_2(.din(w_dff_B_CSmh3Je67_2),.dout(w_dff_B_bYRmQvUm5_2),.clk(gclk));
	jdff dff_B_h0oRvhMQ9_2(.din(w_dff_B_bYRmQvUm5_2),.dout(w_dff_B_h0oRvhMQ9_2),.clk(gclk));
	jdff dff_A_qHBl9uKS2_1(.dout(w_G116gat_0[1]),.din(w_dff_A_qHBl9uKS2_1),.clk(gclk));
	jdff dff_A_6ZSykUXi2_1(.dout(w_dff_A_qHBl9uKS2_1),.din(w_dff_A_6ZSykUXi2_1),.clk(gclk));
	jdff dff_A_WhvCCJdA1_1(.dout(w_dff_A_6ZSykUXi2_1),.din(w_dff_A_WhvCCJdA1_1),.clk(gclk));
	jdff dff_A_Sy6TL7yt6_1(.dout(w_dff_A_WhvCCJdA1_1),.din(w_dff_A_Sy6TL7yt6_1),.clk(gclk));
	jdff dff_A_dyRndxjG7_1(.dout(w_dff_A_Sy6TL7yt6_1),.din(w_dff_A_dyRndxjG7_1),.clk(gclk));
	jdff dff_A_a6m6ldqn7_1(.dout(w_dff_A_dyRndxjG7_1),.din(w_dff_A_a6m6ldqn7_1),.clk(gclk));
	jdff dff_A_QQdI9oVS9_0(.dout(w_G189gat_2[0]),.din(w_dff_A_QQdI9oVS9_0),.clk(gclk));
	jdff dff_A_oNEUMF918_0(.dout(w_dff_A_QQdI9oVS9_0),.din(w_dff_A_oNEUMF918_0),.clk(gclk));
	jdff dff_A_UzPspmBP3_0(.dout(w_dff_A_oNEUMF918_0),.din(w_dff_A_UzPspmBP3_0),.clk(gclk));
	jdff dff_A_Aq8Fg3Xa2_0(.dout(w_dff_A_UzPspmBP3_0),.din(w_dff_A_Aq8Fg3Xa2_0),.clk(gclk));
	jdff dff_A_e9JCRNt20_0(.dout(w_dff_A_Aq8Fg3Xa2_0),.din(w_dff_A_e9JCRNt20_0),.clk(gclk));
	jdff dff_A_XUFsdvAL9_0(.dout(w_dff_A_e9JCRNt20_0),.din(w_dff_A_XUFsdvAL9_0),.clk(gclk));
	jdff dff_A_fYzr3aT48_0(.dout(w_dff_A_XUFsdvAL9_0),.din(w_dff_A_fYzr3aT48_0),.clk(gclk));
	jdff dff_A_14aERbys4_0(.dout(w_dff_A_fYzr3aT48_0),.din(w_dff_A_14aERbys4_0),.clk(gclk));
	jdff dff_A_oqx76kKr5_2(.dout(w_G189gat_0[2]),.din(w_dff_A_oqx76kKr5_2),.clk(gclk));
	jdff dff_A_DQ1Z1PfJ2_2(.dout(w_dff_A_oqx76kKr5_2),.din(w_dff_A_DQ1Z1PfJ2_2),.clk(gclk));
	jdff dff_A_eayyPNSI1_2(.dout(w_dff_A_DQ1Z1PfJ2_2),.din(w_dff_A_eayyPNSI1_2),.clk(gclk));
	jdff dff_A_MQ4ZGfIg5_2(.dout(w_dff_A_eayyPNSI1_2),.din(w_dff_A_MQ4ZGfIg5_2),.clk(gclk));
	jdff dff_A_cYE7uU0K1_0(.dout(w_n343_0[0]),.din(w_dff_A_cYE7uU0K1_0),.clk(gclk));
	jdff dff_A_99289PEm0_0(.dout(w_dff_A_cYE7uU0K1_0),.din(w_dff_A_99289PEm0_0),.clk(gclk));
	jdff dff_A_ZKjimvXj0_0(.dout(w_dff_A_99289PEm0_0),.din(w_dff_A_ZKjimvXj0_0),.clk(gclk));
	jdff dff_A_uynJ8NEj6_0(.dout(w_dff_A_ZKjimvXj0_0),.din(w_dff_A_uynJ8NEj6_0),.clk(gclk));
	jdff dff_A_w1PX75V02_0(.dout(w_dff_A_uynJ8NEj6_0),.din(w_dff_A_w1PX75V02_0),.clk(gclk));
	jdff dff_A_rxyxfakq4_0(.dout(w_dff_A_w1PX75V02_0),.din(w_dff_A_rxyxfakq4_0),.clk(gclk));
	jdff dff_B_sSOx9gG42_1(.din(n341),.dout(w_dff_B_sSOx9gG42_1),.clk(gclk));
	jdff dff_B_6AzZ1H1p5_1(.din(w_dff_B_sSOx9gG42_1),.dout(w_dff_B_6AzZ1H1p5_1),.clk(gclk));
	jdff dff_B_eXhev64l3_1(.din(w_dff_B_6AzZ1H1p5_1),.dout(w_dff_B_eXhev64l3_1),.clk(gclk));
	jdff dff_B_3ls2tTbH4_1(.din(w_dff_B_eXhev64l3_1),.dout(w_dff_B_3ls2tTbH4_1),.clk(gclk));
	jdff dff_B_mWfgVQSe2_1(.din(w_dff_B_3ls2tTbH4_1),.dout(w_dff_B_mWfgVQSe2_1),.clk(gclk));
	jdff dff_B_mTKOuLs62_1(.din(w_dff_B_mWfgVQSe2_1),.dout(w_dff_B_mTKOuLs62_1),.clk(gclk));
	jdff dff_B_8HHs6aWx1_1(.din(w_dff_B_mTKOuLs62_1),.dout(w_dff_B_8HHs6aWx1_1),.clk(gclk));
	jdff dff_B_LDgTm4kC5_1(.din(w_dff_B_8HHs6aWx1_1),.dout(w_dff_B_LDgTm4kC5_1),.clk(gclk));
	jdff dff_A_IeXxQwRr4_1(.dout(w_n222_0[1]),.din(w_dff_A_IeXxQwRr4_1),.clk(gclk));
	jdff dff_A_oDNK9dM52_1(.dout(w_dff_A_IeXxQwRr4_1),.din(w_dff_A_oDNK9dM52_1),.clk(gclk));
	jdff dff_A_nsmsM7Vo0_1(.dout(w_dff_A_oDNK9dM52_1),.din(w_dff_A_nsmsM7Vo0_1),.clk(gclk));
	jdff dff_A_tA9KHJR77_1(.dout(w_dff_A_nsmsM7Vo0_1),.din(w_dff_A_tA9KHJR77_1),.clk(gclk));
	jdff dff_A_Cyhj0a630_1(.dout(w_dff_A_tA9KHJR77_1),.din(w_dff_A_Cyhj0a630_1),.clk(gclk));
	jdff dff_A_Z3H8oW8K2_1(.dout(w_dff_A_Cyhj0a630_1),.din(w_dff_A_Z3H8oW8K2_1),.clk(gclk));
	jdff dff_A_xNiTWMvz0_1(.dout(w_dff_A_Z3H8oW8K2_1),.din(w_dff_A_xNiTWMvz0_1),.clk(gclk));
	jdff dff_A_4LfsyQc45_1(.dout(w_dff_A_xNiTWMvz0_1),.din(w_dff_A_4LfsyQc45_1),.clk(gclk));
	jdff dff_A_hgne0GEA0_0(.dout(w_n97_0[0]),.din(w_dff_A_hgne0GEA0_0),.clk(gclk));
	jdff dff_A_5iBE1NWo9_0(.dout(w_dff_A_hgne0GEA0_0),.din(w_dff_A_5iBE1NWo9_0),.clk(gclk));
	jdff dff_A_xEFdfxMG1_0(.dout(w_dff_A_5iBE1NWo9_0),.din(w_dff_A_xEFdfxMG1_0),.clk(gclk));
	jdff dff_A_wZPeJeD78_1(.dout(w_G143gat_0[1]),.din(w_dff_A_wZPeJeD78_1),.clk(gclk));
	jdff dff_B_H5rML4Bq6_2(.din(G143gat),.dout(w_dff_B_H5rML4Bq6_2),.clk(gclk));
	jdff dff_B_XUM3G9YB3_2(.din(w_dff_B_H5rML4Bq6_2),.dout(w_dff_B_XUM3G9YB3_2),.clk(gclk));
	jdff dff_B_GcG3CTAF9_2(.din(w_dff_B_XUM3G9YB3_2),.dout(w_dff_B_GcG3CTAF9_2),.clk(gclk));
	jdff dff_B_dot5MtOb6_2(.din(w_dff_B_GcG3CTAF9_2),.dout(w_dff_B_dot5MtOb6_2),.clk(gclk));
	jdff dff_A_XteMjSZF9_2(.dout(w_n148_1[2]),.din(w_dff_A_XteMjSZF9_2),.clk(gclk));
	jdff dff_A_PlGa8xbR6_2(.dout(w_dff_A_XteMjSZF9_2),.din(w_dff_A_PlGa8xbR6_2),.clk(gclk));
	jdff dff_A_8MOAOxRw6_1(.dout(w_G111gat_0[1]),.din(w_dff_A_8MOAOxRw6_1),.clk(gclk));
	jdff dff_A_fN5ygeVL3_1(.dout(w_dff_A_8MOAOxRw6_1),.din(w_dff_A_fN5ygeVL3_1),.clk(gclk));
	jdff dff_A_JgVbIWJL5_1(.dout(w_dff_A_fN5ygeVL3_1),.din(w_dff_A_JgVbIWJL5_1),.clk(gclk));
	jdff dff_A_JglYVlhD9_1(.dout(w_dff_A_JgVbIWJL5_1),.din(w_dff_A_JglYVlhD9_1),.clk(gclk));
	jdff dff_A_4mivqqko8_1(.dout(w_dff_A_JglYVlhD9_1),.din(w_dff_A_4mivqqko8_1),.clk(gclk));
	jdff dff_A_8giyetID5_1(.dout(w_dff_A_4mivqqko8_1),.din(w_dff_A_8giyetID5_1),.clk(gclk));
	jdff dff_A_VoTRGCWD8_2(.dout(w_G183gat_0[2]),.din(w_dff_A_VoTRGCWD8_2),.clk(gclk));
	jdff dff_A_0P9PFKav6_2(.dout(w_dff_A_VoTRGCWD8_2),.din(w_dff_A_0P9PFKav6_2),.clk(gclk));
	jdff dff_A_xjpJJIxn4_2(.dout(w_dff_A_0P9PFKav6_2),.din(w_dff_A_xjpJJIxn4_2),.clk(gclk));
	jdff dff_A_Rg0lTCs67_2(.dout(w_dff_A_xjpJJIxn4_2),.din(w_dff_A_Rg0lTCs67_2),.clk(gclk));
	jdff dff_A_cZXvq4qV6_2(.dout(w_dff_A_Rg0lTCs67_2),.din(w_dff_A_cZXvq4qV6_2),.clk(gclk));
	jdff dff_A_UhbXes9l8_2(.dout(w_dff_A_cZXvq4qV6_2),.din(w_dff_A_UhbXes9l8_2),.clk(gclk));
	jdff dff_A_IgmkuNQI7_2(.dout(w_dff_A_UhbXes9l8_2),.din(w_dff_A_IgmkuNQI7_2),.clk(gclk));
	jdff dff_A_OWSYhHc90_2(.dout(w_dff_A_IgmkuNQI7_2),.din(w_dff_A_OWSYhHc90_2),.clk(gclk));
	jdff dff_A_kNBxYv8t5_0(.dout(w_n339_0[0]),.din(w_dff_A_kNBxYv8t5_0),.clk(gclk));
	jdff dff_A_7mb8LDXE0_0(.dout(w_dff_A_kNBxYv8t5_0),.din(w_dff_A_7mb8LDXE0_0),.clk(gclk));
	jdff dff_A_30AxGuti7_0(.dout(w_dff_A_7mb8LDXE0_0),.din(w_dff_A_30AxGuti7_0),.clk(gclk));
	jdff dff_A_U9PRKNo19_0(.dout(w_dff_A_30AxGuti7_0),.din(w_dff_A_U9PRKNo19_0),.clk(gclk));
	jdff dff_A_Zn4YRXEX2_0(.dout(w_dff_A_U9PRKNo19_0),.din(w_dff_A_Zn4YRXEX2_0),.clk(gclk));
	jdff dff_A_a2PKnu931_0(.dout(w_dff_A_Zn4YRXEX2_0),.din(w_dff_A_a2PKnu931_0),.clk(gclk));
	jdff dff_A_NxHilTNr9_0(.dout(w_dff_A_a2PKnu931_0),.din(w_dff_A_NxHilTNr9_0),.clk(gclk));
	jdff dff_B_zKATrJC61_1(.din(n337),.dout(w_dff_B_zKATrJC61_1),.clk(gclk));
	jdff dff_B_tFzcNDQB6_1(.din(w_dff_B_zKATrJC61_1),.dout(w_dff_B_tFzcNDQB6_1),.clk(gclk));
	jdff dff_B_6w5U4doO2_1(.din(w_dff_B_tFzcNDQB6_1),.dout(w_dff_B_6w5U4doO2_1),.clk(gclk));
	jdff dff_B_bR7s2PsI3_1(.din(w_dff_B_6w5U4doO2_1),.dout(w_dff_B_bR7s2PsI3_1),.clk(gclk));
	jdff dff_B_qbjWD4IA1_1(.din(w_dff_B_bR7s2PsI3_1),.dout(w_dff_B_qbjWD4IA1_1),.clk(gclk));
	jdff dff_B_93zzVgNs4_1(.din(w_dff_B_qbjWD4IA1_1),.dout(w_dff_B_93zzVgNs4_1),.clk(gclk));
	jdff dff_B_bGqRnnrb1_1(.din(w_dff_B_93zzVgNs4_1),.dout(w_dff_B_bGqRnnrb1_1),.clk(gclk));
	jdff dff_B_glwFMbs99_1(.din(w_dff_B_bGqRnnrb1_1),.dout(w_dff_B_glwFMbs99_1),.clk(gclk));
	jdff dff_B_CsfeRIgW3_1(.din(w_dff_B_glwFMbs99_1),.dout(w_dff_B_CsfeRIgW3_1),.clk(gclk));
	jdff dff_A_jPfP6liW8_2(.dout(w_n336_0[2]),.din(w_dff_A_jPfP6liW8_2),.clk(gclk));
	jdff dff_A_ZqMaRV2H7_2(.dout(w_dff_A_jPfP6liW8_2),.din(w_dff_A_ZqMaRV2H7_2),.clk(gclk));
	jdff dff_A_bGJ9bNfQ5_2(.dout(w_dff_A_ZqMaRV2H7_2),.din(w_dff_A_bGJ9bNfQ5_2),.clk(gclk));
	jdff dff_A_5dOh7JfE7_2(.dout(w_dff_A_bGJ9bNfQ5_2),.din(w_dff_A_5dOh7JfE7_2),.clk(gclk));
	jdff dff_A_4vBgFoIK6_2(.dout(w_dff_A_5dOh7JfE7_2),.din(w_dff_A_4vBgFoIK6_2),.clk(gclk));
	jdff dff_A_Nl4mGuNV9_2(.dout(w_dff_A_4vBgFoIK6_2),.din(w_dff_A_Nl4mGuNV9_2),.clk(gclk));
	jdff dff_A_JOw5s2Eq2_2(.dout(w_dff_A_Nl4mGuNV9_2),.din(w_dff_A_JOw5s2Eq2_2),.clk(gclk));
	jdff dff_A_xK92jhr56_2(.dout(w_dff_A_JOw5s2Eq2_2),.din(w_dff_A_xK92jhr56_2),.clk(gclk));
	jdff dff_A_ipW7HfAD2_2(.dout(w_dff_A_xK92jhr56_2),.din(w_dff_A_ipW7HfAD2_2),.clk(gclk));
	jdff dff_B_i9r3DG767_0(.din(n333),.dout(w_dff_B_i9r3DG767_0),.clk(gclk));
	jdff dff_B_ciqDUL263_0(.din(n332),.dout(w_dff_B_ciqDUL263_0),.clk(gclk));
	jdff dff_B_MvlAQtoZ1_0(.din(w_dff_B_ciqDUL263_0),.dout(w_dff_B_MvlAQtoZ1_0),.clk(gclk));
	jdff dff_B_m3ntz6Ex2_0(.din(w_dff_B_MvlAQtoZ1_0),.dout(w_dff_B_m3ntz6Ex2_0),.clk(gclk));
	jdff dff_B_XIBcCA2F5_0(.din(w_dff_B_m3ntz6Ex2_0),.dout(w_dff_B_XIBcCA2F5_0),.clk(gclk));
	jdff dff_A_y3mouBv03_0(.dout(w_G153gat_0[0]),.din(w_dff_A_y3mouBv03_0),.clk(gclk));
	jdff dff_A_mRobThW06_0(.dout(w_dff_A_y3mouBv03_0),.din(w_dff_A_mRobThW06_0),.clk(gclk));
	jdff dff_A_YFJmtlCU5_0(.dout(w_dff_A_mRobThW06_0),.din(w_dff_A_YFJmtlCU5_0),.clk(gclk));
	jdff dff_A_kXQhz9PI4_0(.dout(w_dff_A_YFJmtlCU5_0),.din(w_dff_A_kXQhz9PI4_0),.clk(gclk));
	jdff dff_A_ax5WHUV90_2(.dout(w_G153gat_0[2]),.din(w_dff_A_ax5WHUV90_2),.clk(gclk));
	jdff dff_A_Ko2aLk6Z1_2(.dout(w_dff_A_ax5WHUV90_2),.din(w_dff_A_Ko2aLk6Z1_2),.clk(gclk));
	jdff dff_A_8WT2TR5T9_2(.dout(w_dff_A_Ko2aLk6Z1_2),.din(w_dff_A_8WT2TR5T9_2),.clk(gclk));
	jdff dff_A_E94MrDL39_2(.dout(w_dff_A_8WT2TR5T9_2),.din(w_dff_A_E94MrDL39_2),.clk(gclk));
	jdff dff_A_26RT9joY1_2(.dout(w_dff_A_E94MrDL39_2),.din(w_dff_A_26RT9joY1_2),.clk(gclk));
	jdff dff_A_8UkbWSPV4_0(.dout(w_G106gat_0[0]),.din(w_dff_A_8UkbWSPV4_0),.clk(gclk));
	jdff dff_A_jOc1Jrnr3_0(.dout(w_dff_A_8UkbWSPV4_0),.din(w_dff_A_jOc1Jrnr3_0),.clk(gclk));
	jdff dff_A_McXe5nSs8_0(.dout(w_dff_A_jOc1Jrnr3_0),.din(w_dff_A_McXe5nSs8_0),.clk(gclk));
	jdff dff_A_fVWiohJz8_0(.dout(w_dff_A_McXe5nSs8_0),.din(w_dff_A_fVWiohJz8_0),.clk(gclk));
	jdff dff_A_glkzfi5T9_0(.dout(w_dff_A_fVWiohJz8_0),.din(w_dff_A_glkzfi5T9_0),.clk(gclk));
	jdff dff_A_B83qHL3A6_0(.dout(w_dff_A_glkzfi5T9_0),.din(w_dff_A_B83qHL3A6_0),.clk(gclk));
	jdff dff_A_334p8xQ43_1(.dout(w_G177gat_1[1]),.din(w_dff_A_334p8xQ43_1),.clk(gclk));
	jdff dff_A_WAu5TI1a0_1(.dout(w_dff_A_334p8xQ43_1),.din(w_dff_A_WAu5TI1a0_1),.clk(gclk));
	jdff dff_A_maI4D0hJ8_1(.dout(w_dff_A_WAu5TI1a0_1),.din(w_dff_A_maI4D0hJ8_1),.clk(gclk));
	jdff dff_A_oJxUuxOI2_1(.dout(w_dff_A_maI4D0hJ8_1),.din(w_dff_A_oJxUuxOI2_1),.clk(gclk));
	jdff dff_A_KQyuikLw0_1(.dout(w_dff_A_oJxUuxOI2_1),.din(w_dff_A_KQyuikLw0_1),.clk(gclk));
	jdff dff_A_Nba9897K8_1(.dout(w_dff_A_KQyuikLw0_1),.din(w_dff_A_Nba9897K8_1),.clk(gclk));
	jdff dff_A_ajnsYlh83_1(.dout(w_dff_A_Nba9897K8_1),.din(w_dff_A_ajnsYlh83_1),.clk(gclk));
	jdff dff_A_VKL9Ekpq5_1(.dout(w_dff_A_ajnsYlh83_1),.din(w_dff_A_VKL9Ekpq5_1),.clk(gclk));
	jdff dff_A_ZQhRPJSx0_1(.dout(w_dff_A_VKL9Ekpq5_1),.din(w_dff_A_ZQhRPJSx0_1),.clk(gclk));
	jdff dff_A_xm8pmE884_1(.dout(w_G177gat_0[1]),.din(w_dff_A_xm8pmE884_1),.clk(gclk));
	jdff dff_A_i40jUrVr9_1(.dout(w_dff_A_xm8pmE884_1),.din(w_dff_A_i40jUrVr9_1),.clk(gclk));
	jdff dff_A_PWeDNBPz6_1(.dout(w_dff_A_i40jUrVr9_1),.din(w_dff_A_PWeDNBPz6_1),.clk(gclk));
	jdff dff_A_8z0yNlva8_1(.dout(w_dff_A_PWeDNBPz6_1),.din(w_dff_A_8z0yNlva8_1),.clk(gclk));
	jdff dff_A_B3n3HVkC2_2(.dout(w_G177gat_0[2]),.din(w_dff_A_B3n3HVkC2_2),.clk(gclk));
	jdff dff_A_mMsfJ8203_2(.dout(w_dff_A_B3n3HVkC2_2),.din(w_dff_A_mMsfJ8203_2),.clk(gclk));
	jdff dff_A_MjWJOxc81_2(.dout(w_dff_A_mMsfJ8203_2),.din(w_dff_A_MjWJOxc81_2),.clk(gclk));
	jdff dff_A_8bcqVPPU3_2(.dout(w_dff_A_MjWJOxc81_2),.din(w_dff_A_8bcqVPPU3_2),.clk(gclk));
	jdff dff_A_nWOC50gK2_2(.dout(w_dff_A_8bcqVPPU3_2),.din(w_dff_A_nWOC50gK2_2),.clk(gclk));
	jdff dff_A_X3CsfTMx8_2(.dout(w_dff_A_nWOC50gK2_2),.din(w_dff_A_X3CsfTMx8_2),.clk(gclk));
	jdff dff_A_4jtYmsgS6_2(.dout(w_dff_A_X3CsfTMx8_2),.din(w_dff_A_4jtYmsgS6_2),.clk(gclk));
	jdff dff_A_9dMYSdZK5_2(.dout(w_dff_A_4jtYmsgS6_2),.din(w_dff_A_9dMYSdZK5_2),.clk(gclk));
	jdff dff_A_fapqLrpq9_2(.dout(w_dff_A_9dMYSdZK5_2),.din(w_dff_A_fapqLrpq9_2),.clk(gclk));
	jdff dff_B_yW24bOoj0_1(.din(n419),.dout(w_dff_B_yW24bOoj0_1),.clk(gclk));
	jdff dff_B_PXIpsMDO0_0(.din(n424),.dout(w_dff_B_PXIpsMDO0_0),.clk(gclk));
	jdff dff_B_1lNdlfgg1_0(.din(w_dff_B_PXIpsMDO0_0),.dout(w_dff_B_1lNdlfgg1_0),.clk(gclk));
	jdff dff_A_J3TufkYU2_0(.dout(w_G246gat_0[0]),.din(w_dff_A_J3TufkYU2_0),.clk(gclk));
	jdff dff_A_0oS0ytmE4_0(.dout(w_dff_A_J3TufkYU2_0),.din(w_dff_A_0oS0ytmE4_0),.clk(gclk));
	jdff dff_A_5EeMiH4l1_0(.dout(w_dff_A_0oS0ytmE4_0),.din(w_dff_A_5EeMiH4l1_0),.clk(gclk));
	jdff dff_A_nQrjMWle6_0(.dout(w_dff_A_5EeMiH4l1_0),.din(w_dff_A_nQrjMWle6_0),.clk(gclk));
	jdff dff_A_8mjQFyAe5_0(.dout(w_dff_A_nQrjMWle6_0),.din(w_dff_A_8mjQFyAe5_0),.clk(gclk));
	jdff dff_A_wpFHotuG2_0(.dout(w_dff_A_8mjQFyAe5_0),.din(w_dff_A_wpFHotuG2_0),.clk(gclk));
	jdff dff_A_cYDbRQww9_0(.dout(w_dff_A_wpFHotuG2_0),.din(w_dff_A_cYDbRQww9_0),.clk(gclk));
	jdff dff_A_bJRktpWx4_0(.dout(w_dff_A_cYDbRQww9_0),.din(w_dff_A_bJRktpWx4_0),.clk(gclk));
	jdff dff_A_l59Oc1ZP9_2(.dout(w_G246gat_0[2]),.din(w_dff_A_l59Oc1ZP9_2),.clk(gclk));
	jdff dff_A_ZnS2gN058_2(.dout(w_dff_A_l59Oc1ZP9_2),.din(w_dff_A_ZnS2gN058_2),.clk(gclk));
	jdff dff_A_McmTfj3E8_2(.dout(w_dff_A_ZnS2gN058_2),.din(w_dff_A_McmTfj3E8_2),.clk(gclk));
	jdff dff_A_ENDYzWRt5_2(.dout(w_dff_A_McmTfj3E8_2),.din(w_dff_A_ENDYzWRt5_2),.clk(gclk));
	jdff dff_A_MQjCafdt2_2(.dout(w_dff_A_ENDYzWRt5_2),.din(w_dff_A_MQjCafdt2_2),.clk(gclk));
	jdff dff_A_INQieLpD8_2(.dout(w_dff_A_MQjCafdt2_2),.din(w_dff_A_INQieLpD8_2),.clk(gclk));
	jdff dff_A_jUMdPeOn3_2(.dout(w_dff_A_INQieLpD8_2),.din(w_dff_A_jUMdPeOn3_2),.clk(gclk));
	jdff dff_B_FuEt0jiw2_3(.din(G246gat),.dout(w_dff_B_FuEt0jiw2_3),.clk(gclk));
	jdff dff_B_a8ZUsWrQ6_0(.din(n422),.dout(w_dff_B_a8ZUsWrQ6_0),.clk(gclk));
	jdff dff_B_7CxqC9hv5_0(.din(w_dff_B_a8ZUsWrQ6_0),.dout(w_dff_B_7CxqC9hv5_0),.clk(gclk));
	jdff dff_B_X2daWbQK3_0(.din(w_dff_B_7CxqC9hv5_0),.dout(w_dff_B_X2daWbQK3_0),.clk(gclk));
	jdff dff_B_KR80YAfB2_0(.din(w_dff_B_X2daWbQK3_0),.dout(w_dff_B_KR80YAfB2_0),.clk(gclk));
	jdff dff_B_oFcLweFb0_0(.din(w_dff_B_KR80YAfB2_0),.dout(w_dff_B_oFcLweFb0_0),.clk(gclk));
	jdff dff_B_NmhCqco59_0(.din(w_dff_B_oFcLweFb0_0),.dout(w_dff_B_NmhCqco59_0),.clk(gclk));
	jdff dff_B_DeNkSHNd1_0(.din(w_dff_B_NmhCqco59_0),.dout(w_dff_B_DeNkSHNd1_0),.clk(gclk));
	jdff dff_B_AWGhTw5V5_0(.din(w_dff_B_DeNkSHNd1_0),.dout(w_dff_B_AWGhTw5V5_0),.clk(gclk));
	jdff dff_B_HeOxiRsb9_0(.din(w_dff_B_AWGhTw5V5_0),.dout(w_dff_B_HeOxiRsb9_0),.clk(gclk));
	jdff dff_B_X1cVvvvP1_0(.din(w_dff_B_HeOxiRsb9_0),.dout(w_dff_B_X1cVvvvP1_0),.clk(gclk));
	jdff dff_A_l3dyGvki7_1(.dout(w_G96gat_0[1]),.din(w_dff_A_l3dyGvki7_1),.clk(gclk));
	jdff dff_A_5gSeBWFA1_1(.dout(w_dff_A_l3dyGvki7_1),.din(w_dff_A_5gSeBWFA1_1),.clk(gclk));
	jdff dff_A_fuPD4Wj19_1(.dout(w_dff_A_5gSeBWFA1_1),.din(w_dff_A_fuPD4Wj19_1),.clk(gclk));
	jdff dff_A_GCysLHp14_1(.dout(w_dff_A_fuPD4Wj19_1),.din(w_dff_A_GCysLHp14_1),.clk(gclk));
	jdff dff_A_56i1vK9h4_1(.dout(w_dff_A_GCysLHp14_1),.din(w_dff_A_56i1vK9h4_1),.clk(gclk));
	jdff dff_A_WHbkWSbK3_1(.dout(w_dff_A_56i1vK9h4_1),.din(w_dff_A_WHbkWSbK3_1),.clk(gclk));
	jdff dff_A_mHazPNP62_0(.dout(w_n420_0[0]),.din(w_dff_A_mHazPNP62_0),.clk(gclk));
	jdff dff_A_jRhd2ij34_0(.dout(w_dff_A_mHazPNP62_0),.din(w_dff_A_jRhd2ij34_0),.clk(gclk));
	jdff dff_A_TWAme1XX3_0(.dout(w_dff_A_jRhd2ij34_0),.din(w_dff_A_TWAme1XX3_0),.clk(gclk));
	jdff dff_A_gw1ZNbC50_0(.dout(w_dff_A_TWAme1XX3_0),.din(w_dff_A_gw1ZNbC50_0),.clk(gclk));
	jdff dff_A_uByAPhOX3_0(.dout(w_dff_A_gw1ZNbC50_0),.din(w_dff_A_uByAPhOX3_0),.clk(gclk));
	jdff dff_A_9bIjw1zb2_0(.dout(w_dff_A_uByAPhOX3_0),.din(w_dff_A_9bIjw1zb2_0),.clk(gclk));
	jdff dff_A_9snBwZOH6_0(.dout(w_dff_A_9bIjw1zb2_0),.din(w_dff_A_9snBwZOH6_0),.clk(gclk));
	jdff dff_A_SpZ9MXzk7_0(.dout(w_dff_A_9snBwZOH6_0),.din(w_dff_A_SpZ9MXzk7_0),.clk(gclk));
	jdff dff_A_tt70Y21S8_0(.dout(w_dff_A_SpZ9MXzk7_0),.din(w_dff_A_tt70Y21S8_0),.clk(gclk));
	jdff dff_A_Jf5HE9pc1_0(.dout(w_dff_A_tt70Y21S8_0),.din(w_dff_A_Jf5HE9pc1_0),.clk(gclk));
	jdff dff_A_jpgYigNZ1_0(.dout(w_G228gat_0[0]),.din(w_dff_A_jpgYigNZ1_0),.clk(gclk));
	jdff dff_B_jIOpMdkz7_3(.din(G228gat),.dout(w_dff_B_jIOpMdkz7_3),.clk(gclk));
	jdff dff_B_wEZAlOlh8_3(.din(w_dff_B_jIOpMdkz7_3),.dout(w_dff_B_wEZAlOlh8_3),.clk(gclk));
	jdff dff_B_0WCv3TLZ4_3(.din(w_dff_B_wEZAlOlh8_3),.dout(w_dff_B_0WCv3TLZ4_3),.clk(gclk));
	jdff dff_B_cmbRQYD50_3(.din(w_dff_B_0WCv3TLZ4_3),.dout(w_dff_B_cmbRQYD50_3),.clk(gclk));
	jdff dff_B_eAxTthJk6_3(.din(w_dff_B_cmbRQYD50_3),.dout(w_dff_B_eAxTthJk6_3),.clk(gclk));
	jdff dff_B_KsX5GkW32_3(.din(w_dff_B_eAxTthJk6_3),.dout(w_dff_B_KsX5GkW32_3),.clk(gclk));
	jdff dff_B_UooiwDuE6_3(.din(w_dff_B_KsX5GkW32_3),.dout(w_dff_B_UooiwDuE6_3),.clk(gclk));
	jdff dff_B_XaUMzDJl3_3(.din(w_dff_B_UooiwDuE6_3),.dout(w_dff_B_XaUMzDJl3_3),.clk(gclk));
	jdff dff_B_CFuqkUPg8_3(.din(w_dff_B_XaUMzDJl3_3),.dout(w_dff_B_CFuqkUPg8_3),.clk(gclk));
	jdff dff_B_WmpA10mb3_0(.din(n325),.dout(w_dff_B_WmpA10mb3_0),.clk(gclk));
	jdff dff_B_9q0iVMlk8_0(.din(n324),.dout(w_dff_B_9q0iVMlk8_0),.clk(gclk));
	jdff dff_B_znw2Letk3_0(.din(w_dff_B_9q0iVMlk8_0),.dout(w_dff_B_znw2Letk3_0),.clk(gclk));
	jdff dff_B_2Xn32A0M5_0(.din(w_dff_B_znw2Letk3_0),.dout(w_dff_B_2Xn32A0M5_0),.clk(gclk));
	jdff dff_B_FNdWpG6L9_0(.din(w_dff_B_2Xn32A0M5_0),.dout(w_dff_B_FNdWpG6L9_0),.clk(gclk));
	jdff dff_A_DbDIXG4L9_1(.dout(w_G149gat_0[1]),.din(w_dff_A_DbDIXG4L9_1),.clk(gclk));
	jdff dff_B_GMGR8vUN1_2(.din(G149gat),.dout(w_dff_B_GMGR8vUN1_2),.clk(gclk));
	jdff dff_B_4hxEKc4C6_2(.din(w_dff_B_GMGR8vUN1_2),.dout(w_dff_B_4hxEKc4C6_2),.clk(gclk));
	jdff dff_B_GKshyJAs5_2(.din(w_dff_B_4hxEKc4C6_2),.dout(w_dff_B_GKshyJAs5_2),.clk(gclk));
	jdff dff_B_QQafkqky1_2(.din(w_dff_B_GKshyJAs5_2),.dout(w_dff_B_QQafkqky1_2),.clk(gclk));
	jdff dff_A_o7YaiDDE6_0(.dout(w_n162_0[0]),.din(w_dff_A_o7YaiDDE6_0),.clk(gclk));
	jdff dff_B_za8Oaqir8_1(.din(n157),.dout(w_dff_B_za8Oaqir8_1),.clk(gclk));
	jdff dff_B_Bhc3yBAC4_1(.din(n150),.dout(w_dff_B_Bhc3yBAC4_1),.clk(gclk));
	jdff dff_A_iD8pjJNg7_0(.dout(w_n152_0[0]),.din(w_dff_A_iD8pjJNg7_0),.clk(gclk));
	jdff dff_A_7uVQtD3w3_0(.dout(w_n151_0[0]),.din(w_dff_A_7uVQtD3w3_0),.clk(gclk));
	jdff dff_B_dvlmMZNO4_2(.din(n151),.dout(w_dff_B_dvlmMZNO4_2),.clk(gclk));
	jdff dff_A_cwhJZiCj7_0(.dout(w_n149_0[0]),.din(w_dff_A_cwhJZiCj7_0),.clk(gclk));
	jdff dff_A_wiFWWXhH9_0(.dout(w_dff_A_cwhJZiCj7_0),.din(w_dff_A_wiFWWXhH9_0),.clk(gclk));
	jdff dff_A_xFSlZ5xQ9_1(.dout(w_n111_0[1]),.din(w_dff_A_xFSlZ5xQ9_1),.clk(gclk));
	jdff dff_A_BQoxbgMb8_0(.dout(w_G42gat_1[0]),.din(w_dff_A_BQoxbgMb8_0),.clk(gclk));
	jdff dff_A_QEZn7ZAO1_0(.dout(w_n95_0[0]),.din(w_dff_A_QEZn7ZAO1_0),.clk(gclk));
	jdff dff_A_rP2600wd7_0(.dout(w_dff_A_QEZn7ZAO1_0),.din(w_dff_A_rP2600wd7_0),.clk(gclk));
	jdff dff_A_HbOCAKGA8_0(.dout(w_dff_A_rP2600wd7_0),.din(w_dff_A_HbOCAKGA8_0),.clk(gclk));
	jdff dff_A_LBtVcvM64_2(.dout(w_n95_0[2]),.din(w_dff_A_LBtVcvM64_2),.clk(gclk));
	jdff dff_A_B2NdSyJ34_2(.dout(w_dff_A_LBtVcvM64_2),.din(w_dff_A_B2NdSyJ34_2),.clk(gclk));
	jdff dff_A_11kSvh163_2(.dout(w_G17gat_2[2]),.din(w_dff_A_11kSvh163_2),.clk(gclk));
	jdff dff_A_hUzUa7W96_2(.dout(w_dff_A_11kSvh163_2),.din(w_dff_A_hUzUa7W96_2),.clk(gclk));
	jdff dff_A_eHHhQ4o84_1(.dout(w_G101gat_0[1]),.din(w_dff_A_eHHhQ4o84_1),.clk(gclk));
	jdff dff_A_01w6qS8Y7_1(.dout(w_dff_A_eHHhQ4o84_1),.din(w_dff_A_01w6qS8Y7_1),.clk(gclk));
	jdff dff_A_Dk4KRjiK0_1(.dout(w_dff_A_01w6qS8Y7_1),.din(w_dff_A_Dk4KRjiK0_1),.clk(gclk));
	jdff dff_A_GXOmb7M46_1(.dout(w_dff_A_Dk4KRjiK0_1),.din(w_dff_A_GXOmb7M46_1),.clk(gclk));
	jdff dff_A_DGKLle9m8_1(.dout(w_dff_A_GXOmb7M46_1),.din(w_dff_A_DGKLle9m8_1),.clk(gclk));
	jdff dff_A_1ljbPany4_1(.dout(w_dff_A_DGKLle9m8_1),.din(w_dff_A_1ljbPany4_1),.clk(gclk));
	jdff dff_A_vFeJ34va1_1(.dout(w_n306_0[1]),.din(w_dff_A_vFeJ34va1_1),.clk(gclk));
	jdff dff_A_PUuizGx86_1(.dout(w_dff_A_vFeJ34va1_1),.din(w_dff_A_PUuizGx86_1),.clk(gclk));
	jdff dff_A_kvs579UK1_2(.dout(w_n306_0[2]),.din(w_dff_A_kvs579UK1_2),.clk(gclk));
	jdff dff_A_MAiR4MzR9_2(.dout(w_dff_A_kvs579UK1_2),.din(w_dff_A_MAiR4MzR9_2),.clk(gclk));
	jdff dff_A_QWcMVJQJ4_2(.dout(w_G447gat_0[2]),.din(w_dff_A_QWcMVJQJ4_2),.clk(gclk));
	jdff dff_A_Gf9ahnaf0_1(.dout(w_G51gat_1[1]),.din(w_dff_A_Gf9ahnaf0_1),.clk(gclk));
	jdff dff_A_sZpEfjxm0_0(.dout(w_G80gat_0[0]),.din(w_dff_A_sZpEfjxm0_0),.clk(gclk));
	jdff dff_A_jwJe59Ba3_0(.dout(w_dff_A_sZpEfjxm0_0),.din(w_dff_A_jwJe59Ba3_0),.clk(gclk));
	jdff dff_A_c5k75pdr7_2(.dout(w_G80gat_0[2]),.din(w_dff_A_c5k75pdr7_2),.clk(gclk));
	jdff dff_A_u03eq0JM0_0(.dout(w_n86_0[0]),.din(w_dff_A_u03eq0JM0_0),.clk(gclk));
	jdff dff_A_mQhW8Len8_0(.dout(w_dff_A_u03eq0JM0_0),.din(w_dff_A_mQhW8Len8_0),.clk(gclk));
	jdff dff_A_1QWScWbE0_0(.dout(w_G29gat_0[0]),.din(w_dff_A_1QWScWbE0_0),.clk(gclk));
	jdff dff_A_IB2i9IMQ5_0(.dout(w_dff_A_1QWScWbE0_0),.din(w_dff_A_IB2i9IMQ5_0),.clk(gclk));
	jdff dff_A_MKDZ5sdi8_0(.dout(w_dff_A_IB2i9IMQ5_0),.din(w_dff_A_MKDZ5sdi8_0),.clk(gclk));
	jdff dff_A_ksBqX5wI0_0(.dout(w_G17gat_1[0]),.din(w_dff_A_ksBqX5wI0_0),.clk(gclk));
	jdff dff_A_K1eXx5hX9_0(.dout(w_dff_A_ksBqX5wI0_0),.din(w_dff_A_K1eXx5hX9_0),.clk(gclk));
	jdff dff_A_OEXtbVry9_0(.dout(w_dff_A_K1eXx5hX9_0),.din(w_dff_A_OEXtbVry9_0),.clk(gclk));
	jdff dff_A_c58gNbtU5_0(.dout(w_dff_A_OEXtbVry9_0),.din(w_dff_A_c58gNbtU5_0),.clk(gclk));
	jdff dff_A_N2CFVJcF4_1(.dout(w_G17gat_1[1]),.din(w_dff_A_N2CFVJcF4_1),.clk(gclk));
	jdff dff_A_MWMuOC8p1_1(.dout(w_dff_A_N2CFVJcF4_1),.din(w_dff_A_MWMuOC8p1_1),.clk(gclk));
	jdff dff_A_ILxZoKM10_1(.dout(w_dff_A_MWMuOC8p1_1),.din(w_dff_A_ILxZoKM10_1),.clk(gclk));
	jdff dff_B_AN5zqfCe9_2(.din(n144),.dout(w_dff_B_AN5zqfCe9_2),.clk(gclk));
	jdff dff_B_YizhvhEt1_2(.din(w_dff_B_AN5zqfCe9_2),.dout(w_dff_B_YizhvhEt1_2),.clk(gclk));
	jdff dff_B_11dJR2233_2(.din(w_dff_B_YizhvhEt1_2),.dout(w_dff_B_11dJR2233_2),.clk(gclk));
	jdff dff_B_P7cmgdDp0_2(.din(w_dff_B_11dJR2233_2),.dout(w_dff_B_P7cmgdDp0_2),.clk(gclk));
	jdff dff_A_vzH8a5IH7_0(.dout(w_G237gat_0[0]),.din(w_dff_A_vzH8a5IH7_0),.clk(gclk));
	jdff dff_A_2XlABTEg4_0(.dout(w_dff_A_vzH8a5IH7_0),.din(w_dff_A_2XlABTEg4_0),.clk(gclk));
	jdff dff_A_dwxSv1RD3_0(.dout(w_dff_A_2XlABTEg4_0),.din(w_dff_A_dwxSv1RD3_0),.clk(gclk));
	jdff dff_A_ia9jZOxB4_0(.dout(w_dff_A_dwxSv1RD3_0),.din(w_dff_A_ia9jZOxB4_0),.clk(gclk));
	jdff dff_A_BLBEEKtT3_0(.dout(w_dff_A_ia9jZOxB4_0),.din(w_dff_A_BLBEEKtT3_0),.clk(gclk));
	jdff dff_A_EWvd61zV2_0(.dout(w_dff_A_BLBEEKtT3_0),.din(w_dff_A_EWvd61zV2_0),.clk(gclk));
	jdff dff_A_4VxHcluu1_0(.dout(w_dff_A_EWvd61zV2_0),.din(w_dff_A_4VxHcluu1_0),.clk(gclk));
	jdff dff_A_casShWez8_0(.dout(w_dff_A_4VxHcluu1_0),.din(w_dff_A_casShWez8_0),.clk(gclk));
	jdff dff_A_pJ1fMVAp6_0(.dout(w_dff_A_casShWez8_0),.din(w_dff_A_pJ1fMVAp6_0),.clk(gclk));
	jdff dff_A_zmkTIIpv0_2(.dout(w_G237gat_0[2]),.din(w_dff_A_zmkTIIpv0_2),.clk(gclk));
	jdff dff_A_rfF6o2O05_2(.dout(w_dff_A_zmkTIIpv0_2),.din(w_dff_A_rfF6o2O05_2),.clk(gclk));
	jdff dff_A_2c7NHnrQ1_2(.dout(w_dff_A_rfF6o2O05_2),.din(w_dff_A_2c7NHnrQ1_2),.clk(gclk));
	jdff dff_A_xQNw0OnY0_2(.dout(w_dff_A_2c7NHnrQ1_2),.din(w_dff_A_xQNw0OnY0_2),.clk(gclk));
	jdff dff_A_gPeBrji92_2(.dout(w_dff_A_xQNw0OnY0_2),.din(w_dff_A_gPeBrji92_2),.clk(gclk));
	jdff dff_A_z8eXRr5A9_2(.dout(w_dff_A_gPeBrji92_2),.din(w_dff_A_z8eXRr5A9_2),.clk(gclk));
	jdff dff_A_2HEyaCAt9_2(.dout(w_dff_A_z8eXRr5A9_2),.din(w_dff_A_2HEyaCAt9_2),.clk(gclk));
	jdff dff_A_ZwDqmSz09_2(.dout(w_dff_A_2HEyaCAt9_2),.din(w_dff_A_ZwDqmSz09_2),.clk(gclk));
	jdff dff_A_8DAk1jc00_2(.dout(w_dff_A_ZwDqmSz09_2),.din(w_dff_A_8DAk1jc00_2),.clk(gclk));
	jdff dff_A_u44msslo6_0(.dout(w_n178_0[0]),.din(w_dff_A_u44msslo6_0),.clk(gclk));
	jdff dff_A_AyCz4Zwr6_0(.dout(w_dff_A_u44msslo6_0),.din(w_dff_A_AyCz4Zwr6_0),.clk(gclk));
	jdff dff_A_IAfzXxZD6_0(.dout(w_dff_A_AyCz4Zwr6_0),.din(w_dff_A_IAfzXxZD6_0),.clk(gclk));
	jdff dff_A_yoTihmYo6_0(.dout(w_dff_A_IAfzXxZD6_0),.din(w_dff_A_yoTihmYo6_0),.clk(gclk));
	jdff dff_A_OX7Xvnjl4_0(.dout(w_dff_A_yoTihmYo6_0),.din(w_dff_A_OX7Xvnjl4_0),.clk(gclk));
	jdff dff_A_VzplXodn2_0(.dout(w_dff_A_OX7Xvnjl4_0),.din(w_dff_A_VzplXodn2_0),.clk(gclk));
	jdff dff_B_fzp31Fxl5_0(.din(n176),.dout(w_dff_B_fzp31Fxl5_0),.clk(gclk));
	jdff dff_A_rMNiHgEZ7_1(.dout(w_n122_0[1]),.din(w_dff_A_rMNiHgEZ7_1),.clk(gclk));
	jdff dff_A_T8HV43pC6_1(.dout(w_dff_A_rMNiHgEZ7_1),.din(w_dff_A_T8HV43pC6_1),.clk(gclk));
	jdff dff_A_uDr2tGyW1_1(.dout(w_dff_A_T8HV43pC6_1),.din(w_dff_A_uDr2tGyW1_1),.clk(gclk));
	jdff dff_A_KOJIDJab2_1(.dout(w_G68gat_0[1]),.din(w_dff_A_KOJIDJab2_1),.clk(gclk));
	jdff dff_A_OfANTNyH8_1(.dout(w_dff_A_KOJIDJab2_1),.din(w_dff_A_OfANTNyH8_1),.clk(gclk));
	jdff dff_A_NZCi6Slt0_1(.dout(w_dff_A_OfANTNyH8_1),.din(w_dff_A_NZCi6Slt0_1),.clk(gclk));
	jdff dff_A_8SHFtRHc4_1(.dout(w_dff_A_NZCi6Slt0_1),.din(w_dff_A_8SHFtRHc4_1),.clk(gclk));
	jdff dff_A_LtKNNQCe6_1(.dout(w_G42gat_0[1]),.din(w_dff_A_LtKNNQCe6_1),.clk(gclk));
	jdff dff_A_e94DEHcZ9_2(.dout(w_G42gat_0[2]),.din(w_dff_A_e94DEHcZ9_2),.clk(gclk));
	jdff dff_A_BGG8C18W6_1(.dout(w_G1gat_0[1]),.din(w_dff_A_BGG8C18W6_1),.clk(gclk));
	jdff dff_A_2CGoF0uM9_1(.dout(w_dff_A_BGG8C18W6_1),.din(w_dff_A_2CGoF0uM9_1),.clk(gclk));
	jdff dff_A_cgeT17iR4_1(.dout(w_dff_A_2CGoF0uM9_1),.din(w_dff_A_cgeT17iR4_1),.clk(gclk));
	jdff dff_A_UMPOKdDL3_1(.dout(w_dff_A_cgeT17iR4_1),.din(w_dff_A_UMPOKdDL3_1),.clk(gclk));
	jdff dff_A_0qB5OCiB0_1(.dout(w_dff_A_UMPOKdDL3_1),.din(w_dff_A_0qB5OCiB0_1),.clk(gclk));
	jdff dff_A_YZFSoUtL7_1(.dout(w_G13gat_0[1]),.din(w_dff_A_YZFSoUtL7_1),.clk(gclk));
	jdff dff_A_o0FLiivG4_0(.dout(w_G55gat_0[0]),.din(w_dff_A_o0FLiivG4_0),.clk(gclk));
	jdff dff_A_ZQT4YDvQ5_1(.dout(w_G55gat_0[1]),.din(w_dff_A_ZQT4YDvQ5_1),.clk(gclk));
	jdff dff_A_nKJDjkL34_1(.dout(w_dff_A_ZQT4YDvQ5_1),.din(w_dff_A_nKJDjkL34_1),.clk(gclk));
	jdff dff_B_JujjifIW0_3(.din(G55gat),.dout(w_dff_B_JujjifIW0_3),.clk(gclk));
	jdff dff_B_xxKpXUDp7_3(.din(w_dff_B_JujjifIW0_3),.dout(w_dff_B_xxKpXUDp7_3),.clk(gclk));
	jdff dff_A_b32WYCJk1_1(.dout(w_G171gat_0[1]),.din(w_dff_A_b32WYCJk1_1),.clk(gclk));
	jdff dff_A_y9MYhpIM0_1(.dout(w_dff_A_b32WYCJk1_1),.din(w_dff_A_y9MYhpIM0_1),.clk(gclk));
	jdff dff_A_cK461G5Q8_1(.dout(w_dff_A_y9MYhpIM0_1),.din(w_dff_A_cK461G5Q8_1),.clk(gclk));
	jdff dff_A_YFSbislH0_1(.dout(w_dff_A_cK461G5Q8_1),.din(w_dff_A_YFSbislH0_1),.clk(gclk));
	jdff dff_A_SXcLFPzC3_1(.dout(w_dff_A_YFSbislH0_1),.din(w_dff_A_SXcLFPzC3_1),.clk(gclk));
	jdff dff_A_2PfAN4md2_1(.dout(w_dff_A_SXcLFPzC3_1),.din(w_dff_A_2PfAN4md2_1),.clk(gclk));
	jdff dff_A_Wf8QQ8nr5_1(.dout(w_dff_A_2PfAN4md2_1),.din(w_dff_A_Wf8QQ8nr5_1),.clk(gclk));
	jdff dff_A_t5wWn38Z1_1(.dout(w_dff_A_Wf8QQ8nr5_1),.din(w_dff_A_t5wWn38Z1_1),.clk(gclk));
	jdff dff_A_cLI7CXP81_1(.dout(w_dff_A_t5wWn38Z1_1),.din(w_dff_A_cLI7CXP81_1),.clk(gclk));
	jdff dff_A_abAoN42z4_2(.dout(w_G171gat_0[2]),.din(w_dff_A_abAoN42z4_2),.clk(gclk));
	jdff dff_A_CxrZOvs51_2(.dout(w_dff_A_abAoN42z4_2),.din(w_dff_A_CxrZOvs51_2),.clk(gclk));
	jdff dff_A_Sl3VTDFt4_2(.dout(w_dff_A_CxrZOvs51_2),.din(w_dff_A_Sl3VTDFt4_2),.clk(gclk));
	jdff dff_A_Ow6Vz5Bk2_2(.dout(w_dff_A_Sl3VTDFt4_2),.din(w_dff_A_Ow6Vz5Bk2_2),.clk(gclk));
	jdff dff_A_HnFtxZya6_2(.dout(w_dff_A_Ow6Vz5Bk2_2),.din(w_dff_A_HnFtxZya6_2),.clk(gclk));
	jdff dff_A_F5mEcLzK3_2(.dout(w_dff_A_HnFtxZya6_2),.din(w_dff_A_F5mEcLzK3_2),.clk(gclk));
	jdff dff_A_6zpQ6MoK7_2(.dout(w_dff_A_F5mEcLzK3_2),.din(w_dff_A_6zpQ6MoK7_2),.clk(gclk));
	jdff dff_A_BLh70akQ9_2(.dout(w_dff_A_6zpQ6MoK7_2),.din(w_dff_A_BLh70akQ9_2),.clk(gclk));
	jdff dff_A_GgjU2x5B7_2(.dout(w_dff_A_BLh70akQ9_2),.din(w_dff_A_GgjU2x5B7_2),.clk(gclk));
	jdff dff_A_4Wk26QqG3_2(.dout(w_dff_A_GgjU2x5B7_2),.din(w_dff_A_4Wk26QqG3_2),.clk(gclk));
	jdff dff_A_SoV7oXqQ8_2(.dout(w_dff_A_4Wk26QqG3_2),.din(w_dff_A_SoV7oXqQ8_2),.clk(gclk));
	jdff dff_A_GIQFJFMG3_2(.dout(w_dff_A_hNzUy3C26_0),.din(w_dff_A_GIQFJFMG3_2),.clk(gclk));
	jdff dff_A_hNzUy3C26_0(.dout(w_dff_A_HYf2Kd3O9_0),.din(w_dff_A_hNzUy3C26_0),.clk(gclk));
	jdff dff_A_HYf2Kd3O9_0(.dout(w_dff_A_UdpQExC23_0),.din(w_dff_A_HYf2Kd3O9_0),.clk(gclk));
	jdff dff_A_UdpQExC23_0(.dout(w_dff_A_9gIHhL6b2_0),.din(w_dff_A_UdpQExC23_0),.clk(gclk));
	jdff dff_A_9gIHhL6b2_0(.dout(w_dff_A_5xrj0h4v1_0),.din(w_dff_A_9gIHhL6b2_0),.clk(gclk));
	jdff dff_A_5xrj0h4v1_0(.dout(w_dff_A_ydi3PxeD3_0),.din(w_dff_A_5xrj0h4v1_0),.clk(gclk));
	jdff dff_A_ydi3PxeD3_0(.dout(w_dff_A_4YhMBPaD5_0),.din(w_dff_A_ydi3PxeD3_0),.clk(gclk));
	jdff dff_A_4YhMBPaD5_0(.dout(w_dff_A_CVIhwn9k7_0),.din(w_dff_A_4YhMBPaD5_0),.clk(gclk));
	jdff dff_A_CVIhwn9k7_0(.dout(w_dff_A_VtF0Vlih0_0),.din(w_dff_A_CVIhwn9k7_0),.clk(gclk));
	jdff dff_A_VtF0Vlih0_0(.dout(w_dff_A_COl9Ozh81_0),.din(w_dff_A_VtF0Vlih0_0),.clk(gclk));
	jdff dff_A_COl9Ozh81_0(.dout(w_dff_A_yBQKFVk97_0),.din(w_dff_A_COl9Ozh81_0),.clk(gclk));
	jdff dff_A_yBQKFVk97_0(.dout(w_dff_A_jQWl3CYa9_0),.din(w_dff_A_yBQKFVk97_0),.clk(gclk));
	jdff dff_A_jQWl3CYa9_0(.dout(w_dff_A_Bo2R4vhC6_0),.din(w_dff_A_jQWl3CYa9_0),.clk(gclk));
	jdff dff_A_Bo2R4vhC6_0(.dout(w_dff_A_m23qoWUg7_0),.din(w_dff_A_Bo2R4vhC6_0),.clk(gclk));
	jdff dff_A_m23qoWUg7_0(.dout(w_dff_A_YHBTuddm7_0),.din(w_dff_A_m23qoWUg7_0),.clk(gclk));
	jdff dff_A_YHBTuddm7_0(.dout(w_dff_A_PWXCsM2V4_0),.din(w_dff_A_YHBTuddm7_0),.clk(gclk));
	jdff dff_A_PWXCsM2V4_0(.dout(w_dff_A_Y795aTw98_0),.din(w_dff_A_PWXCsM2V4_0),.clk(gclk));
	jdff dff_A_Y795aTw98_0(.dout(w_dff_A_xtXY9Qgj6_0),.din(w_dff_A_Y795aTw98_0),.clk(gclk));
	jdff dff_A_xtXY9Qgj6_0(.dout(w_dff_A_jyPsdBQa2_0),.din(w_dff_A_xtXY9Qgj6_0),.clk(gclk));
	jdff dff_A_jyPsdBQa2_0(.dout(w_dff_A_IXkJs7qp0_0),.din(w_dff_A_jyPsdBQa2_0),.clk(gclk));
	jdff dff_A_IXkJs7qp0_0(.dout(w_dff_A_nAJ0ve2e5_0),.din(w_dff_A_IXkJs7qp0_0),.clk(gclk));
	jdff dff_A_nAJ0ve2e5_0(.dout(w_dff_A_MWRKUUOo2_0),.din(w_dff_A_nAJ0ve2e5_0),.clk(gclk));
	jdff dff_A_MWRKUUOo2_0(.dout(w_dff_A_PTVaSj3j8_0),.din(w_dff_A_MWRKUUOo2_0),.clk(gclk));
	jdff dff_A_PTVaSj3j8_0(.dout(w_dff_A_rryMQYmW9_0),.din(w_dff_A_PTVaSj3j8_0),.clk(gclk));
	jdff dff_A_rryMQYmW9_0(.dout(w_dff_A_R3S5W4FU9_0),.din(w_dff_A_rryMQYmW9_0),.clk(gclk));
	jdff dff_A_R3S5W4FU9_0(.dout(G388gat),.din(w_dff_A_R3S5W4FU9_0),.clk(gclk));
	jdff dff_A_fbbwZBC94_2(.dout(w_dff_A_jSaQN0AA1_0),.din(w_dff_A_fbbwZBC94_2),.clk(gclk));
	jdff dff_A_jSaQN0AA1_0(.dout(w_dff_A_ve7dmZ7D2_0),.din(w_dff_A_jSaQN0AA1_0),.clk(gclk));
	jdff dff_A_ve7dmZ7D2_0(.dout(w_dff_A_1hRV36Pn6_0),.din(w_dff_A_ve7dmZ7D2_0),.clk(gclk));
	jdff dff_A_1hRV36Pn6_0(.dout(w_dff_A_PBm86oNA2_0),.din(w_dff_A_1hRV36Pn6_0),.clk(gclk));
	jdff dff_A_PBm86oNA2_0(.dout(w_dff_A_2KRlKMh88_0),.din(w_dff_A_PBm86oNA2_0),.clk(gclk));
	jdff dff_A_2KRlKMh88_0(.dout(w_dff_A_uRl38xeF7_0),.din(w_dff_A_2KRlKMh88_0),.clk(gclk));
	jdff dff_A_uRl38xeF7_0(.dout(w_dff_A_6pObr9Ln7_0),.din(w_dff_A_uRl38xeF7_0),.clk(gclk));
	jdff dff_A_6pObr9Ln7_0(.dout(w_dff_A_uMrqc91R6_0),.din(w_dff_A_6pObr9Ln7_0),.clk(gclk));
	jdff dff_A_uMrqc91R6_0(.dout(w_dff_A_va78vqte5_0),.din(w_dff_A_uMrqc91R6_0),.clk(gclk));
	jdff dff_A_va78vqte5_0(.dout(w_dff_A_tPACDJAS1_0),.din(w_dff_A_va78vqte5_0),.clk(gclk));
	jdff dff_A_tPACDJAS1_0(.dout(w_dff_A_yoYm7YRD7_0),.din(w_dff_A_tPACDJAS1_0),.clk(gclk));
	jdff dff_A_yoYm7YRD7_0(.dout(w_dff_A_IYLSHnMS1_0),.din(w_dff_A_yoYm7YRD7_0),.clk(gclk));
	jdff dff_A_IYLSHnMS1_0(.dout(w_dff_A_UdbzN5yS0_0),.din(w_dff_A_IYLSHnMS1_0),.clk(gclk));
	jdff dff_A_UdbzN5yS0_0(.dout(w_dff_A_F9RWbxcd9_0),.din(w_dff_A_UdbzN5yS0_0),.clk(gclk));
	jdff dff_A_F9RWbxcd9_0(.dout(w_dff_A_ZTbwGDAX5_0),.din(w_dff_A_F9RWbxcd9_0),.clk(gclk));
	jdff dff_A_ZTbwGDAX5_0(.dout(w_dff_A_m8haK0v40_0),.din(w_dff_A_ZTbwGDAX5_0),.clk(gclk));
	jdff dff_A_m8haK0v40_0(.dout(w_dff_A_zSKpGYeN9_0),.din(w_dff_A_m8haK0v40_0),.clk(gclk));
	jdff dff_A_zSKpGYeN9_0(.dout(w_dff_A_4eQtuMk60_0),.din(w_dff_A_zSKpGYeN9_0),.clk(gclk));
	jdff dff_A_4eQtuMk60_0(.dout(w_dff_A_NIYwisdb9_0),.din(w_dff_A_4eQtuMk60_0),.clk(gclk));
	jdff dff_A_NIYwisdb9_0(.dout(w_dff_A_Ijs7conF8_0),.din(w_dff_A_NIYwisdb9_0),.clk(gclk));
	jdff dff_A_Ijs7conF8_0(.dout(w_dff_A_uwTdvjEV1_0),.din(w_dff_A_Ijs7conF8_0),.clk(gclk));
	jdff dff_A_uwTdvjEV1_0(.dout(w_dff_A_x0aaxlvi6_0),.din(w_dff_A_uwTdvjEV1_0),.clk(gclk));
	jdff dff_A_x0aaxlvi6_0(.dout(w_dff_A_iuAo3Qz44_0),.din(w_dff_A_x0aaxlvi6_0),.clk(gclk));
	jdff dff_A_iuAo3Qz44_0(.dout(w_dff_A_XotlsMEW3_0),.din(w_dff_A_iuAo3Qz44_0),.clk(gclk));
	jdff dff_A_XotlsMEW3_0(.dout(w_dff_A_QTpWsiND3_0),.din(w_dff_A_XotlsMEW3_0),.clk(gclk));
	jdff dff_A_QTpWsiND3_0(.dout(G389gat),.din(w_dff_A_QTpWsiND3_0),.clk(gclk));
	jdff dff_A_B6Z4XMwz7_2(.dout(w_dff_A_wRmIRAMI0_0),.din(w_dff_A_B6Z4XMwz7_2),.clk(gclk));
	jdff dff_A_wRmIRAMI0_0(.dout(w_dff_A_S3m42r8M6_0),.din(w_dff_A_wRmIRAMI0_0),.clk(gclk));
	jdff dff_A_S3m42r8M6_0(.dout(w_dff_A_LZUfgs5F0_0),.din(w_dff_A_S3m42r8M6_0),.clk(gclk));
	jdff dff_A_LZUfgs5F0_0(.dout(w_dff_A_yEjoW1Qk3_0),.din(w_dff_A_LZUfgs5F0_0),.clk(gclk));
	jdff dff_A_yEjoW1Qk3_0(.dout(w_dff_A_OcKqlTmC9_0),.din(w_dff_A_yEjoW1Qk3_0),.clk(gclk));
	jdff dff_A_OcKqlTmC9_0(.dout(w_dff_A_yW90sm0m6_0),.din(w_dff_A_OcKqlTmC9_0),.clk(gclk));
	jdff dff_A_yW90sm0m6_0(.dout(w_dff_A_dP2rJuKa1_0),.din(w_dff_A_yW90sm0m6_0),.clk(gclk));
	jdff dff_A_dP2rJuKa1_0(.dout(w_dff_A_sZzN5gI33_0),.din(w_dff_A_dP2rJuKa1_0),.clk(gclk));
	jdff dff_A_sZzN5gI33_0(.dout(w_dff_A_Jo3KCtou0_0),.din(w_dff_A_sZzN5gI33_0),.clk(gclk));
	jdff dff_A_Jo3KCtou0_0(.dout(w_dff_A_kgFX5hg30_0),.din(w_dff_A_Jo3KCtou0_0),.clk(gclk));
	jdff dff_A_kgFX5hg30_0(.dout(w_dff_A_VUBk74w62_0),.din(w_dff_A_kgFX5hg30_0),.clk(gclk));
	jdff dff_A_VUBk74w62_0(.dout(w_dff_A_eSqNkEQo7_0),.din(w_dff_A_VUBk74w62_0),.clk(gclk));
	jdff dff_A_eSqNkEQo7_0(.dout(w_dff_A_cYzay5hk4_0),.din(w_dff_A_eSqNkEQo7_0),.clk(gclk));
	jdff dff_A_cYzay5hk4_0(.dout(w_dff_A_iO0Gkb0I3_0),.din(w_dff_A_cYzay5hk4_0),.clk(gclk));
	jdff dff_A_iO0Gkb0I3_0(.dout(w_dff_A_HuXGHdDg8_0),.din(w_dff_A_iO0Gkb0I3_0),.clk(gclk));
	jdff dff_A_HuXGHdDg8_0(.dout(w_dff_A_NKwVIKgT5_0),.din(w_dff_A_HuXGHdDg8_0),.clk(gclk));
	jdff dff_A_NKwVIKgT5_0(.dout(w_dff_A_JDDW7R9A6_0),.din(w_dff_A_NKwVIKgT5_0),.clk(gclk));
	jdff dff_A_JDDW7R9A6_0(.dout(w_dff_A_ZANfmTyv5_0),.din(w_dff_A_JDDW7R9A6_0),.clk(gclk));
	jdff dff_A_ZANfmTyv5_0(.dout(w_dff_A_asSSJUnh0_0),.din(w_dff_A_ZANfmTyv5_0),.clk(gclk));
	jdff dff_A_asSSJUnh0_0(.dout(w_dff_A_9Co9E0rq3_0),.din(w_dff_A_asSSJUnh0_0),.clk(gclk));
	jdff dff_A_9Co9E0rq3_0(.dout(w_dff_A_4quQ58v91_0),.din(w_dff_A_9Co9E0rq3_0),.clk(gclk));
	jdff dff_A_4quQ58v91_0(.dout(w_dff_A_kJqkduKb7_0),.din(w_dff_A_4quQ58v91_0),.clk(gclk));
	jdff dff_A_kJqkduKb7_0(.dout(w_dff_A_VpMAyCip6_0),.din(w_dff_A_kJqkduKb7_0),.clk(gclk));
	jdff dff_A_VpMAyCip6_0(.dout(w_dff_A_xi3aKtf99_0),.din(w_dff_A_VpMAyCip6_0),.clk(gclk));
	jdff dff_A_xi3aKtf99_0(.dout(w_dff_A_gSloLsBp0_0),.din(w_dff_A_xi3aKtf99_0),.clk(gclk));
	jdff dff_A_gSloLsBp0_0(.dout(G390gat),.din(w_dff_A_gSloLsBp0_0),.clk(gclk));
	jdff dff_A_SfdgPlOZ3_2(.dout(w_dff_A_vBWDEs5c1_0),.din(w_dff_A_SfdgPlOZ3_2),.clk(gclk));
	jdff dff_A_vBWDEs5c1_0(.dout(w_dff_A_KuiwLew39_0),.din(w_dff_A_vBWDEs5c1_0),.clk(gclk));
	jdff dff_A_KuiwLew39_0(.dout(w_dff_A_nyLFFR8d9_0),.din(w_dff_A_KuiwLew39_0),.clk(gclk));
	jdff dff_A_nyLFFR8d9_0(.dout(w_dff_A_k7ZNQdRN9_0),.din(w_dff_A_nyLFFR8d9_0),.clk(gclk));
	jdff dff_A_k7ZNQdRN9_0(.dout(w_dff_A_hcdzESoJ0_0),.din(w_dff_A_k7ZNQdRN9_0),.clk(gclk));
	jdff dff_A_hcdzESoJ0_0(.dout(w_dff_A_kggYYSB87_0),.din(w_dff_A_hcdzESoJ0_0),.clk(gclk));
	jdff dff_A_kggYYSB87_0(.dout(w_dff_A_HjgcAcXl8_0),.din(w_dff_A_kggYYSB87_0),.clk(gclk));
	jdff dff_A_HjgcAcXl8_0(.dout(w_dff_A_CUB2NcDZ0_0),.din(w_dff_A_HjgcAcXl8_0),.clk(gclk));
	jdff dff_A_CUB2NcDZ0_0(.dout(w_dff_A_Ba809Wac7_0),.din(w_dff_A_CUB2NcDZ0_0),.clk(gclk));
	jdff dff_A_Ba809Wac7_0(.dout(w_dff_A_JxlBc8Sd7_0),.din(w_dff_A_Ba809Wac7_0),.clk(gclk));
	jdff dff_A_JxlBc8Sd7_0(.dout(w_dff_A_02TkcAql6_0),.din(w_dff_A_JxlBc8Sd7_0),.clk(gclk));
	jdff dff_A_02TkcAql6_0(.dout(w_dff_A_7xwQTvFu0_0),.din(w_dff_A_02TkcAql6_0),.clk(gclk));
	jdff dff_A_7xwQTvFu0_0(.dout(w_dff_A_f3kPU7WM8_0),.din(w_dff_A_7xwQTvFu0_0),.clk(gclk));
	jdff dff_A_f3kPU7WM8_0(.dout(w_dff_A_NJtBqYph0_0),.din(w_dff_A_f3kPU7WM8_0),.clk(gclk));
	jdff dff_A_NJtBqYph0_0(.dout(w_dff_A_KPZQvkGt3_0),.din(w_dff_A_NJtBqYph0_0),.clk(gclk));
	jdff dff_A_KPZQvkGt3_0(.dout(w_dff_A_Qe8WeW3m9_0),.din(w_dff_A_KPZQvkGt3_0),.clk(gclk));
	jdff dff_A_Qe8WeW3m9_0(.dout(w_dff_A_MeuYDjcY3_0),.din(w_dff_A_Qe8WeW3m9_0),.clk(gclk));
	jdff dff_A_MeuYDjcY3_0(.dout(w_dff_A_6973Muxp3_0),.din(w_dff_A_MeuYDjcY3_0),.clk(gclk));
	jdff dff_A_6973Muxp3_0(.dout(w_dff_A_aVP18PBt1_0),.din(w_dff_A_6973Muxp3_0),.clk(gclk));
	jdff dff_A_aVP18PBt1_0(.dout(w_dff_A_uBj7VEeD6_0),.din(w_dff_A_aVP18PBt1_0),.clk(gclk));
	jdff dff_A_uBj7VEeD6_0(.dout(w_dff_A_A4ak95H22_0),.din(w_dff_A_uBj7VEeD6_0),.clk(gclk));
	jdff dff_A_A4ak95H22_0(.dout(w_dff_A_WGXjJkGa5_0),.din(w_dff_A_A4ak95H22_0),.clk(gclk));
	jdff dff_A_WGXjJkGa5_0(.dout(w_dff_A_HAdk9kq35_0),.din(w_dff_A_WGXjJkGa5_0),.clk(gclk));
	jdff dff_A_HAdk9kq35_0(.dout(w_dff_A_lXsy4q6L0_0),.din(w_dff_A_HAdk9kq35_0),.clk(gclk));
	jdff dff_A_lXsy4q6L0_0(.dout(w_dff_A_ymRDstN55_0),.din(w_dff_A_lXsy4q6L0_0),.clk(gclk));
	jdff dff_A_ymRDstN55_0(.dout(w_dff_A_XUrvf1oR3_0),.din(w_dff_A_ymRDstN55_0),.clk(gclk));
	jdff dff_A_XUrvf1oR3_0(.dout(G391gat),.din(w_dff_A_XUrvf1oR3_0),.clk(gclk));
	jdff dff_A_bkmCrY7r7_2(.dout(w_dff_A_hQPliWiR0_0),.din(w_dff_A_bkmCrY7r7_2),.clk(gclk));
	jdff dff_A_hQPliWiR0_0(.dout(w_dff_A_WCCPC7mf8_0),.din(w_dff_A_hQPliWiR0_0),.clk(gclk));
	jdff dff_A_WCCPC7mf8_0(.dout(w_dff_A_J46msa4H9_0),.din(w_dff_A_WCCPC7mf8_0),.clk(gclk));
	jdff dff_A_J46msa4H9_0(.dout(w_dff_A_JK3WZePZ1_0),.din(w_dff_A_J46msa4H9_0),.clk(gclk));
	jdff dff_A_JK3WZePZ1_0(.dout(w_dff_A_wVqMcpz18_0),.din(w_dff_A_JK3WZePZ1_0),.clk(gclk));
	jdff dff_A_wVqMcpz18_0(.dout(w_dff_A_7dLJFCyl3_0),.din(w_dff_A_wVqMcpz18_0),.clk(gclk));
	jdff dff_A_7dLJFCyl3_0(.dout(w_dff_A_Dj3KXIK08_0),.din(w_dff_A_7dLJFCyl3_0),.clk(gclk));
	jdff dff_A_Dj3KXIK08_0(.dout(w_dff_A_9IAYhGbG7_0),.din(w_dff_A_Dj3KXIK08_0),.clk(gclk));
	jdff dff_A_9IAYhGbG7_0(.dout(w_dff_A_ougHFFr31_0),.din(w_dff_A_9IAYhGbG7_0),.clk(gclk));
	jdff dff_A_ougHFFr31_0(.dout(w_dff_A_qTeYnMfb1_0),.din(w_dff_A_ougHFFr31_0),.clk(gclk));
	jdff dff_A_qTeYnMfb1_0(.dout(w_dff_A_aW7shEvn7_0),.din(w_dff_A_qTeYnMfb1_0),.clk(gclk));
	jdff dff_A_aW7shEvn7_0(.dout(w_dff_A_VIQuqmzX1_0),.din(w_dff_A_aW7shEvn7_0),.clk(gclk));
	jdff dff_A_VIQuqmzX1_0(.dout(w_dff_A_yvNuwgYP6_0),.din(w_dff_A_VIQuqmzX1_0),.clk(gclk));
	jdff dff_A_yvNuwgYP6_0(.dout(w_dff_A_bR1BvdoU1_0),.din(w_dff_A_yvNuwgYP6_0),.clk(gclk));
	jdff dff_A_bR1BvdoU1_0(.dout(w_dff_A_ZKtCFEUh6_0),.din(w_dff_A_bR1BvdoU1_0),.clk(gclk));
	jdff dff_A_ZKtCFEUh6_0(.dout(w_dff_A_DBcX3uwA7_0),.din(w_dff_A_ZKtCFEUh6_0),.clk(gclk));
	jdff dff_A_DBcX3uwA7_0(.dout(w_dff_A_tj90LY1N2_0),.din(w_dff_A_DBcX3uwA7_0),.clk(gclk));
	jdff dff_A_tj90LY1N2_0(.dout(w_dff_A_HACOFh6N6_0),.din(w_dff_A_tj90LY1N2_0),.clk(gclk));
	jdff dff_A_HACOFh6N6_0(.dout(w_dff_A_Am9WZO1c8_0),.din(w_dff_A_HACOFh6N6_0),.clk(gclk));
	jdff dff_A_Am9WZO1c8_0(.dout(w_dff_A_qKtCd8Ts5_0),.din(w_dff_A_Am9WZO1c8_0),.clk(gclk));
	jdff dff_A_qKtCd8Ts5_0(.dout(w_dff_A_Y74HGvs07_0),.din(w_dff_A_qKtCd8Ts5_0),.clk(gclk));
	jdff dff_A_Y74HGvs07_0(.dout(w_dff_A_1RT2dsJt2_0),.din(w_dff_A_Y74HGvs07_0),.clk(gclk));
	jdff dff_A_1RT2dsJt2_0(.dout(w_dff_A_hBxrswGj8_0),.din(w_dff_A_1RT2dsJt2_0),.clk(gclk));
	jdff dff_A_hBxrswGj8_0(.dout(w_dff_A_9onCqjcb8_0),.din(w_dff_A_hBxrswGj8_0),.clk(gclk));
	jdff dff_A_9onCqjcb8_0(.dout(G418gat),.din(w_dff_A_9onCqjcb8_0),.clk(gclk));
	jdff dff_A_1Qm6wZAT2_2(.dout(w_dff_A_fyU4uy8r8_0),.din(w_dff_A_1Qm6wZAT2_2),.clk(gclk));
	jdff dff_A_fyU4uy8r8_0(.dout(w_dff_A_REviNEA89_0),.din(w_dff_A_fyU4uy8r8_0),.clk(gclk));
	jdff dff_A_REviNEA89_0(.dout(w_dff_A_biMb3fA81_0),.din(w_dff_A_REviNEA89_0),.clk(gclk));
	jdff dff_A_biMb3fA81_0(.dout(w_dff_A_e64spRBK1_0),.din(w_dff_A_biMb3fA81_0),.clk(gclk));
	jdff dff_A_e64spRBK1_0(.dout(w_dff_A_CuqN56HP9_0),.din(w_dff_A_e64spRBK1_0),.clk(gclk));
	jdff dff_A_CuqN56HP9_0(.dout(w_dff_A_zUeRAHfu0_0),.din(w_dff_A_CuqN56HP9_0),.clk(gclk));
	jdff dff_A_zUeRAHfu0_0(.dout(w_dff_A_QDRF8MyT5_0),.din(w_dff_A_zUeRAHfu0_0),.clk(gclk));
	jdff dff_A_QDRF8MyT5_0(.dout(w_dff_A_NwIKnT2t9_0),.din(w_dff_A_QDRF8MyT5_0),.clk(gclk));
	jdff dff_A_NwIKnT2t9_0(.dout(w_dff_A_OkbSKNTw9_0),.din(w_dff_A_NwIKnT2t9_0),.clk(gclk));
	jdff dff_A_OkbSKNTw9_0(.dout(w_dff_A_GIzN6gNR8_0),.din(w_dff_A_OkbSKNTw9_0),.clk(gclk));
	jdff dff_A_GIzN6gNR8_0(.dout(w_dff_A_iceEIwMC3_0),.din(w_dff_A_GIzN6gNR8_0),.clk(gclk));
	jdff dff_A_iceEIwMC3_0(.dout(w_dff_A_JCj4zyd77_0),.din(w_dff_A_iceEIwMC3_0),.clk(gclk));
	jdff dff_A_JCj4zyd77_0(.dout(w_dff_A_TfrNrFBp0_0),.din(w_dff_A_JCj4zyd77_0),.clk(gclk));
	jdff dff_A_TfrNrFBp0_0(.dout(w_dff_A_VjMYD0g27_0),.din(w_dff_A_TfrNrFBp0_0),.clk(gclk));
	jdff dff_A_VjMYD0g27_0(.dout(w_dff_A_UXsqAlfR8_0),.din(w_dff_A_VjMYD0g27_0),.clk(gclk));
	jdff dff_A_UXsqAlfR8_0(.dout(w_dff_A_Gig8wDLv7_0),.din(w_dff_A_UXsqAlfR8_0),.clk(gclk));
	jdff dff_A_Gig8wDLv7_0(.dout(w_dff_A_D8oX5u4W2_0),.din(w_dff_A_Gig8wDLv7_0),.clk(gclk));
	jdff dff_A_D8oX5u4W2_0(.dout(w_dff_A_1iPypINM9_0),.din(w_dff_A_D8oX5u4W2_0),.clk(gclk));
	jdff dff_A_1iPypINM9_0(.dout(w_dff_A_TGbE6zxt8_0),.din(w_dff_A_1iPypINM9_0),.clk(gclk));
	jdff dff_A_TGbE6zxt8_0(.dout(w_dff_A_9IgYhVHZ6_0),.din(w_dff_A_TGbE6zxt8_0),.clk(gclk));
	jdff dff_A_9IgYhVHZ6_0(.dout(w_dff_A_4YkMIkOM9_0),.din(w_dff_A_9IgYhVHZ6_0),.clk(gclk));
	jdff dff_A_4YkMIkOM9_0(.dout(w_dff_A_sEpUOhkm8_0),.din(w_dff_A_4YkMIkOM9_0),.clk(gclk));
	jdff dff_A_sEpUOhkm8_0(.dout(G419gat),.din(w_dff_A_sEpUOhkm8_0),.clk(gclk));
	jdff dff_A_9ZHzostQ4_2(.dout(w_dff_A_acBW3aA58_0),.din(w_dff_A_9ZHzostQ4_2),.clk(gclk));
	jdff dff_A_acBW3aA58_0(.dout(w_dff_A_wfNRpohp9_0),.din(w_dff_A_acBW3aA58_0),.clk(gclk));
	jdff dff_A_wfNRpohp9_0(.dout(w_dff_A_KZUbdoto3_0),.din(w_dff_A_wfNRpohp9_0),.clk(gclk));
	jdff dff_A_KZUbdoto3_0(.dout(w_dff_A_wAsaG9s20_0),.din(w_dff_A_KZUbdoto3_0),.clk(gclk));
	jdff dff_A_wAsaG9s20_0(.dout(w_dff_A_beErWbUR7_0),.din(w_dff_A_wAsaG9s20_0),.clk(gclk));
	jdff dff_A_beErWbUR7_0(.dout(w_dff_A_8ZaBReQ67_0),.din(w_dff_A_beErWbUR7_0),.clk(gclk));
	jdff dff_A_8ZaBReQ67_0(.dout(w_dff_A_0OxHTqHH2_0),.din(w_dff_A_8ZaBReQ67_0),.clk(gclk));
	jdff dff_A_0OxHTqHH2_0(.dout(w_dff_A_1Sm6ge9R7_0),.din(w_dff_A_0OxHTqHH2_0),.clk(gclk));
	jdff dff_A_1Sm6ge9R7_0(.dout(w_dff_A_oFa3N5p55_0),.din(w_dff_A_1Sm6ge9R7_0),.clk(gclk));
	jdff dff_A_oFa3N5p55_0(.dout(w_dff_A_QphaYer82_0),.din(w_dff_A_oFa3N5p55_0),.clk(gclk));
	jdff dff_A_QphaYer82_0(.dout(w_dff_A_cGVdMqKs0_0),.din(w_dff_A_QphaYer82_0),.clk(gclk));
	jdff dff_A_cGVdMqKs0_0(.dout(w_dff_A_2fAN20vg7_0),.din(w_dff_A_cGVdMqKs0_0),.clk(gclk));
	jdff dff_A_2fAN20vg7_0(.dout(w_dff_A_7Up1IEB24_0),.din(w_dff_A_2fAN20vg7_0),.clk(gclk));
	jdff dff_A_7Up1IEB24_0(.dout(w_dff_A_Ga8YSLXj1_0),.din(w_dff_A_7Up1IEB24_0),.clk(gclk));
	jdff dff_A_Ga8YSLXj1_0(.dout(w_dff_A_2EC8B5CU6_0),.din(w_dff_A_Ga8YSLXj1_0),.clk(gclk));
	jdff dff_A_2EC8B5CU6_0(.dout(w_dff_A_MviX3CIa3_0),.din(w_dff_A_2EC8B5CU6_0),.clk(gclk));
	jdff dff_A_MviX3CIa3_0(.dout(w_dff_A_31fFjjjP5_0),.din(w_dff_A_MviX3CIa3_0),.clk(gclk));
	jdff dff_A_31fFjjjP5_0(.dout(w_dff_A_7JhZFazM7_0),.din(w_dff_A_31fFjjjP5_0),.clk(gclk));
	jdff dff_A_7JhZFazM7_0(.dout(w_dff_A_5ND675611_0),.din(w_dff_A_7JhZFazM7_0),.clk(gclk));
	jdff dff_A_5ND675611_0(.dout(w_dff_A_VfkJ2ffF6_0),.din(w_dff_A_5ND675611_0),.clk(gclk));
	jdff dff_A_VfkJ2ffF6_0(.dout(w_dff_A_7ZywvmuN4_0),.din(w_dff_A_VfkJ2ffF6_0),.clk(gclk));
	jdff dff_A_7ZywvmuN4_0(.dout(w_dff_A_7ugerTbt5_0),.din(w_dff_A_7ZywvmuN4_0),.clk(gclk));
	jdff dff_A_7ugerTbt5_0(.dout(w_dff_A_NbqsnwDp3_0),.din(w_dff_A_7ugerTbt5_0),.clk(gclk));
	jdff dff_A_NbqsnwDp3_0(.dout(w_dff_A_zll0YeUD6_0),.din(w_dff_A_NbqsnwDp3_0),.clk(gclk));
	jdff dff_A_zll0YeUD6_0(.dout(G420gat),.din(w_dff_A_zll0YeUD6_0),.clk(gclk));
	jdff dff_A_SkEow26f5_2(.dout(w_dff_A_WTGvmPFJ6_0),.din(w_dff_A_SkEow26f5_2),.clk(gclk));
	jdff dff_A_WTGvmPFJ6_0(.dout(w_dff_A_580p66MJ0_0),.din(w_dff_A_WTGvmPFJ6_0),.clk(gclk));
	jdff dff_A_580p66MJ0_0(.dout(w_dff_A_HAe6mKe86_0),.din(w_dff_A_580p66MJ0_0),.clk(gclk));
	jdff dff_A_HAe6mKe86_0(.dout(w_dff_A_8lztFpFF3_0),.din(w_dff_A_HAe6mKe86_0),.clk(gclk));
	jdff dff_A_8lztFpFF3_0(.dout(w_dff_A_whH2awry4_0),.din(w_dff_A_8lztFpFF3_0),.clk(gclk));
	jdff dff_A_whH2awry4_0(.dout(w_dff_A_pW0Tunmb3_0),.din(w_dff_A_whH2awry4_0),.clk(gclk));
	jdff dff_A_pW0Tunmb3_0(.dout(w_dff_A_8FDJjDhL1_0),.din(w_dff_A_pW0Tunmb3_0),.clk(gclk));
	jdff dff_A_8FDJjDhL1_0(.dout(w_dff_A_1xpN1gvE0_0),.din(w_dff_A_8FDJjDhL1_0),.clk(gclk));
	jdff dff_A_1xpN1gvE0_0(.dout(w_dff_A_tjCnTYPO9_0),.din(w_dff_A_1xpN1gvE0_0),.clk(gclk));
	jdff dff_A_tjCnTYPO9_0(.dout(w_dff_A_q1RjnNjV2_0),.din(w_dff_A_tjCnTYPO9_0),.clk(gclk));
	jdff dff_A_q1RjnNjV2_0(.dout(w_dff_A_lGHzpP2K9_0),.din(w_dff_A_q1RjnNjV2_0),.clk(gclk));
	jdff dff_A_lGHzpP2K9_0(.dout(w_dff_A_8evsPL0x0_0),.din(w_dff_A_lGHzpP2K9_0),.clk(gclk));
	jdff dff_A_8evsPL0x0_0(.dout(w_dff_A_mUrv24N39_0),.din(w_dff_A_8evsPL0x0_0),.clk(gclk));
	jdff dff_A_mUrv24N39_0(.dout(w_dff_A_YUvPkBC11_0),.din(w_dff_A_mUrv24N39_0),.clk(gclk));
	jdff dff_A_YUvPkBC11_0(.dout(w_dff_A_iy99ALRm4_0),.din(w_dff_A_YUvPkBC11_0),.clk(gclk));
	jdff dff_A_iy99ALRm4_0(.dout(w_dff_A_bquknk935_0),.din(w_dff_A_iy99ALRm4_0),.clk(gclk));
	jdff dff_A_bquknk935_0(.dout(w_dff_A_ClWfCns00_0),.din(w_dff_A_bquknk935_0),.clk(gclk));
	jdff dff_A_ClWfCns00_0(.dout(w_dff_A_h6j1DMIR8_0),.din(w_dff_A_ClWfCns00_0),.clk(gclk));
	jdff dff_A_h6j1DMIR8_0(.dout(w_dff_A_Rd2m1PqP1_0),.din(w_dff_A_h6j1DMIR8_0),.clk(gclk));
	jdff dff_A_Rd2m1PqP1_0(.dout(w_dff_A_W7Ta6o5n7_0),.din(w_dff_A_Rd2m1PqP1_0),.clk(gclk));
	jdff dff_A_W7Ta6o5n7_0(.dout(w_dff_A_QN1uYlrj0_0),.din(w_dff_A_W7Ta6o5n7_0),.clk(gclk));
	jdff dff_A_QN1uYlrj0_0(.dout(w_dff_A_oK1GntID5_0),.din(w_dff_A_QN1uYlrj0_0),.clk(gclk));
	jdff dff_A_oK1GntID5_0(.dout(w_dff_A_2lJ3JvEA3_0),.din(w_dff_A_oK1GntID5_0),.clk(gclk));
	jdff dff_A_2lJ3JvEA3_0(.dout(w_dff_A_4uussoog7_0),.din(w_dff_A_2lJ3JvEA3_0),.clk(gclk));
	jdff dff_A_4uussoog7_0(.dout(G421gat),.din(w_dff_A_4uussoog7_0),.clk(gclk));
	jdff dff_A_I6hNTVIN6_2(.dout(w_dff_A_UWL0sjX75_0),.din(w_dff_A_I6hNTVIN6_2),.clk(gclk));
	jdff dff_A_UWL0sjX75_0(.dout(w_dff_A_i3BAsUMv5_0),.din(w_dff_A_UWL0sjX75_0),.clk(gclk));
	jdff dff_A_i3BAsUMv5_0(.dout(w_dff_A_IaZxsaC34_0),.din(w_dff_A_i3BAsUMv5_0),.clk(gclk));
	jdff dff_A_IaZxsaC34_0(.dout(w_dff_A_LtjsvLjX6_0),.din(w_dff_A_IaZxsaC34_0),.clk(gclk));
	jdff dff_A_LtjsvLjX6_0(.dout(w_dff_A_JP1jIevG1_0),.din(w_dff_A_LtjsvLjX6_0),.clk(gclk));
	jdff dff_A_JP1jIevG1_0(.dout(w_dff_A_Nr1C3yTv3_0),.din(w_dff_A_JP1jIevG1_0),.clk(gclk));
	jdff dff_A_Nr1C3yTv3_0(.dout(w_dff_A_3f7IvP7f5_0),.din(w_dff_A_Nr1C3yTv3_0),.clk(gclk));
	jdff dff_A_3f7IvP7f5_0(.dout(w_dff_A_U8xSx5Ew2_0),.din(w_dff_A_3f7IvP7f5_0),.clk(gclk));
	jdff dff_A_U8xSx5Ew2_0(.dout(w_dff_A_FmgqqfDT6_0),.din(w_dff_A_U8xSx5Ew2_0),.clk(gclk));
	jdff dff_A_FmgqqfDT6_0(.dout(w_dff_A_4T3mnRGm0_0),.din(w_dff_A_FmgqqfDT6_0),.clk(gclk));
	jdff dff_A_4T3mnRGm0_0(.dout(w_dff_A_rlDa8G7I0_0),.din(w_dff_A_4T3mnRGm0_0),.clk(gclk));
	jdff dff_A_rlDa8G7I0_0(.dout(w_dff_A_TrBUl0CH8_0),.din(w_dff_A_rlDa8G7I0_0),.clk(gclk));
	jdff dff_A_TrBUl0CH8_0(.dout(w_dff_A_cOteOzgK6_0),.din(w_dff_A_TrBUl0CH8_0),.clk(gclk));
	jdff dff_A_cOteOzgK6_0(.dout(w_dff_A_agQG2JiC2_0),.din(w_dff_A_cOteOzgK6_0),.clk(gclk));
	jdff dff_A_agQG2JiC2_0(.dout(w_dff_A_Umkynk5O8_0),.din(w_dff_A_agQG2JiC2_0),.clk(gclk));
	jdff dff_A_Umkynk5O8_0(.dout(w_dff_A_gdtMSq9E0_0),.din(w_dff_A_Umkynk5O8_0),.clk(gclk));
	jdff dff_A_gdtMSq9E0_0(.dout(w_dff_A_HEEfDagU7_0),.din(w_dff_A_gdtMSq9E0_0),.clk(gclk));
	jdff dff_A_HEEfDagU7_0(.dout(w_dff_A_6iK7sCAt0_0),.din(w_dff_A_HEEfDagU7_0),.clk(gclk));
	jdff dff_A_6iK7sCAt0_0(.dout(w_dff_A_0E8ukRdX8_0),.din(w_dff_A_6iK7sCAt0_0),.clk(gclk));
	jdff dff_A_0E8ukRdX8_0(.dout(w_dff_A_EEPdjaFa1_0),.din(w_dff_A_0E8ukRdX8_0),.clk(gclk));
	jdff dff_A_EEPdjaFa1_0(.dout(w_dff_A_3tBpD3Ub2_0),.din(w_dff_A_EEPdjaFa1_0),.clk(gclk));
	jdff dff_A_3tBpD3Ub2_0(.dout(w_dff_A_HOKKmCWx5_0),.din(w_dff_A_3tBpD3Ub2_0),.clk(gclk));
	jdff dff_A_HOKKmCWx5_0(.dout(w_dff_A_Wa24sCIH3_0),.din(w_dff_A_HOKKmCWx5_0),.clk(gclk));
	jdff dff_A_Wa24sCIH3_0(.dout(w_dff_A_F1ipmiP76_0),.din(w_dff_A_Wa24sCIH3_0),.clk(gclk));
	jdff dff_A_F1ipmiP76_0(.dout(G422gat),.din(w_dff_A_F1ipmiP76_0),.clk(gclk));
	jdff dff_A_T2sNp57Q1_2(.dout(w_dff_A_AViv2ydS4_0),.din(w_dff_A_T2sNp57Q1_2),.clk(gclk));
	jdff dff_A_AViv2ydS4_0(.dout(w_dff_A_mOtVQSuK3_0),.din(w_dff_A_AViv2ydS4_0),.clk(gclk));
	jdff dff_A_mOtVQSuK3_0(.dout(w_dff_A_QmUATijc3_0),.din(w_dff_A_mOtVQSuK3_0),.clk(gclk));
	jdff dff_A_QmUATijc3_0(.dout(w_dff_A_w06XInNC2_0),.din(w_dff_A_QmUATijc3_0),.clk(gclk));
	jdff dff_A_w06XInNC2_0(.dout(w_dff_A_kruvq9g07_0),.din(w_dff_A_w06XInNC2_0),.clk(gclk));
	jdff dff_A_kruvq9g07_0(.dout(w_dff_A_wXbxsZVw8_0),.din(w_dff_A_kruvq9g07_0),.clk(gclk));
	jdff dff_A_wXbxsZVw8_0(.dout(w_dff_A_lM2WTgx74_0),.din(w_dff_A_wXbxsZVw8_0),.clk(gclk));
	jdff dff_A_lM2WTgx74_0(.dout(w_dff_A_lYK3QlDD8_0),.din(w_dff_A_lM2WTgx74_0),.clk(gclk));
	jdff dff_A_lYK3QlDD8_0(.dout(w_dff_A_U8aXldGM7_0),.din(w_dff_A_lYK3QlDD8_0),.clk(gclk));
	jdff dff_A_U8aXldGM7_0(.dout(w_dff_A_H09nZfvu1_0),.din(w_dff_A_U8aXldGM7_0),.clk(gclk));
	jdff dff_A_H09nZfvu1_0(.dout(w_dff_A_phD9twfj6_0),.din(w_dff_A_H09nZfvu1_0),.clk(gclk));
	jdff dff_A_phD9twfj6_0(.dout(w_dff_A_yCaodL0W3_0),.din(w_dff_A_phD9twfj6_0),.clk(gclk));
	jdff dff_A_yCaodL0W3_0(.dout(w_dff_A_B3C2OSum0_0),.din(w_dff_A_yCaodL0W3_0),.clk(gclk));
	jdff dff_A_B3C2OSum0_0(.dout(w_dff_A_eMjIMQTM2_0),.din(w_dff_A_B3C2OSum0_0),.clk(gclk));
	jdff dff_A_eMjIMQTM2_0(.dout(w_dff_A_kQhVdl753_0),.din(w_dff_A_eMjIMQTM2_0),.clk(gclk));
	jdff dff_A_kQhVdl753_0(.dout(w_dff_A_XIIIajo33_0),.din(w_dff_A_kQhVdl753_0),.clk(gclk));
	jdff dff_A_XIIIajo33_0(.dout(w_dff_A_bfTbC6NH3_0),.din(w_dff_A_XIIIajo33_0),.clk(gclk));
	jdff dff_A_bfTbC6NH3_0(.dout(w_dff_A_Aj1U1yTI8_0),.din(w_dff_A_bfTbC6NH3_0),.clk(gclk));
	jdff dff_A_Aj1U1yTI8_0(.dout(w_dff_A_ngAkVC322_0),.din(w_dff_A_Aj1U1yTI8_0),.clk(gclk));
	jdff dff_A_ngAkVC322_0(.dout(w_dff_A_PBgaHB1v6_0),.din(w_dff_A_ngAkVC322_0),.clk(gclk));
	jdff dff_A_PBgaHB1v6_0(.dout(w_dff_A_rGjUSLxV1_0),.din(w_dff_A_PBgaHB1v6_0),.clk(gclk));
	jdff dff_A_rGjUSLxV1_0(.dout(w_dff_A_0bR3ugqN0_0),.din(w_dff_A_rGjUSLxV1_0),.clk(gclk));
	jdff dff_A_0bR3ugqN0_0(.dout(w_dff_A_em60hgpk7_0),.din(w_dff_A_0bR3ugqN0_0),.clk(gclk));
	jdff dff_A_em60hgpk7_0(.dout(w_dff_A_BLJyWh090_0),.din(w_dff_A_em60hgpk7_0),.clk(gclk));
	jdff dff_A_BLJyWh090_0(.dout(w_dff_A_Fusx2Vwr8_0),.din(w_dff_A_BLJyWh090_0),.clk(gclk));
	jdff dff_A_Fusx2Vwr8_0(.dout(G423gat),.din(w_dff_A_Fusx2Vwr8_0),.clk(gclk));
	jdff dff_A_kFfvaOFK5_2(.dout(w_dff_A_OzMqJS1k6_0),.din(w_dff_A_kFfvaOFK5_2),.clk(gclk));
	jdff dff_A_OzMqJS1k6_0(.dout(w_dff_A_RxOJXN9A2_0),.din(w_dff_A_OzMqJS1k6_0),.clk(gclk));
	jdff dff_A_RxOJXN9A2_0(.dout(w_dff_A_58wZptTP9_0),.din(w_dff_A_RxOJXN9A2_0),.clk(gclk));
	jdff dff_A_58wZptTP9_0(.dout(w_dff_A_7imoNw4O6_0),.din(w_dff_A_58wZptTP9_0),.clk(gclk));
	jdff dff_A_7imoNw4O6_0(.dout(w_dff_A_NmI395vY1_0),.din(w_dff_A_7imoNw4O6_0),.clk(gclk));
	jdff dff_A_NmI395vY1_0(.dout(w_dff_A_LaVAz5DS5_0),.din(w_dff_A_NmI395vY1_0),.clk(gclk));
	jdff dff_A_LaVAz5DS5_0(.dout(w_dff_A_wAGIcrs39_0),.din(w_dff_A_LaVAz5DS5_0),.clk(gclk));
	jdff dff_A_wAGIcrs39_0(.dout(w_dff_A_Qtw4eZ4n9_0),.din(w_dff_A_wAGIcrs39_0),.clk(gclk));
	jdff dff_A_Qtw4eZ4n9_0(.dout(w_dff_A_GUNwJM1d3_0),.din(w_dff_A_Qtw4eZ4n9_0),.clk(gclk));
	jdff dff_A_GUNwJM1d3_0(.dout(w_dff_A_tGLuDtpy5_0),.din(w_dff_A_GUNwJM1d3_0),.clk(gclk));
	jdff dff_A_tGLuDtpy5_0(.dout(w_dff_A_0O3iMY6p0_0),.din(w_dff_A_tGLuDtpy5_0),.clk(gclk));
	jdff dff_A_0O3iMY6p0_0(.dout(w_dff_A_AXd9OF3W7_0),.din(w_dff_A_0O3iMY6p0_0),.clk(gclk));
	jdff dff_A_AXd9OF3W7_0(.dout(w_dff_A_WYpEkHrg4_0),.din(w_dff_A_AXd9OF3W7_0),.clk(gclk));
	jdff dff_A_WYpEkHrg4_0(.dout(w_dff_A_rCjwCbZR5_0),.din(w_dff_A_WYpEkHrg4_0),.clk(gclk));
	jdff dff_A_rCjwCbZR5_0(.dout(w_dff_A_P2ceZMPk4_0),.din(w_dff_A_rCjwCbZR5_0),.clk(gclk));
	jdff dff_A_P2ceZMPk4_0(.dout(w_dff_A_Q4tJVLvs2_0),.din(w_dff_A_P2ceZMPk4_0),.clk(gclk));
	jdff dff_A_Q4tJVLvs2_0(.dout(w_dff_A_gnCI5dYD0_0),.din(w_dff_A_Q4tJVLvs2_0),.clk(gclk));
	jdff dff_A_gnCI5dYD0_0(.dout(w_dff_A_E1flEDp32_0),.din(w_dff_A_gnCI5dYD0_0),.clk(gclk));
	jdff dff_A_E1flEDp32_0(.dout(w_dff_A_4wahLqaV1_0),.din(w_dff_A_E1flEDp32_0),.clk(gclk));
	jdff dff_A_4wahLqaV1_0(.dout(w_dff_A_uEZAeyGF3_0),.din(w_dff_A_4wahLqaV1_0),.clk(gclk));
	jdff dff_A_uEZAeyGF3_0(.dout(w_dff_A_QtUIoXPa8_0),.din(w_dff_A_uEZAeyGF3_0),.clk(gclk));
	jdff dff_A_QtUIoXPa8_0(.dout(w_dff_A_gHXN3bwJ7_0),.din(w_dff_A_QtUIoXPa8_0),.clk(gclk));
	jdff dff_A_gHXN3bwJ7_0(.dout(G446gat),.din(w_dff_A_gHXN3bwJ7_0),.clk(gclk));
	jdff dff_A_lEJ8kvaV2_1(.dout(w_dff_A_QmD3fafN3_0),.din(w_dff_A_lEJ8kvaV2_1),.clk(gclk));
	jdff dff_A_QmD3fafN3_0(.dout(w_dff_A_FJLkcpR43_0),.din(w_dff_A_QmD3fafN3_0),.clk(gclk));
	jdff dff_A_FJLkcpR43_0(.dout(w_dff_A_PWAa442S8_0),.din(w_dff_A_FJLkcpR43_0),.clk(gclk));
	jdff dff_A_PWAa442S8_0(.dout(w_dff_A_74lxLGlB1_0),.din(w_dff_A_PWAa442S8_0),.clk(gclk));
	jdff dff_A_74lxLGlB1_0(.dout(w_dff_A_4Tzv2tcl6_0),.din(w_dff_A_74lxLGlB1_0),.clk(gclk));
	jdff dff_A_4Tzv2tcl6_0(.dout(w_dff_A_ayLFv6v43_0),.din(w_dff_A_4Tzv2tcl6_0),.clk(gclk));
	jdff dff_A_ayLFv6v43_0(.dout(w_dff_A_PS2K9Hhq2_0),.din(w_dff_A_ayLFv6v43_0),.clk(gclk));
	jdff dff_A_PS2K9Hhq2_0(.dout(w_dff_A_rZw7cAaJ6_0),.din(w_dff_A_PS2K9Hhq2_0),.clk(gclk));
	jdff dff_A_rZw7cAaJ6_0(.dout(w_dff_A_qXSm7VNz4_0),.din(w_dff_A_rZw7cAaJ6_0),.clk(gclk));
	jdff dff_A_qXSm7VNz4_0(.dout(w_dff_A_btzlUGQO0_0),.din(w_dff_A_qXSm7VNz4_0),.clk(gclk));
	jdff dff_A_btzlUGQO0_0(.dout(w_dff_A_2fwbiHCh5_0),.din(w_dff_A_btzlUGQO0_0),.clk(gclk));
	jdff dff_A_2fwbiHCh5_0(.dout(w_dff_A_bpYxWGFP0_0),.din(w_dff_A_2fwbiHCh5_0),.clk(gclk));
	jdff dff_A_bpYxWGFP0_0(.dout(w_dff_A_wQLMnZ0d6_0),.din(w_dff_A_bpYxWGFP0_0),.clk(gclk));
	jdff dff_A_wQLMnZ0d6_0(.dout(w_dff_A_J2d3jfCx5_0),.din(w_dff_A_wQLMnZ0d6_0),.clk(gclk));
	jdff dff_A_J2d3jfCx5_0(.dout(w_dff_A_tgM0fDix1_0),.din(w_dff_A_J2d3jfCx5_0),.clk(gclk));
	jdff dff_A_tgM0fDix1_0(.dout(w_dff_A_AKEwKhuf3_0),.din(w_dff_A_tgM0fDix1_0),.clk(gclk));
	jdff dff_A_AKEwKhuf3_0(.dout(w_dff_A_vl5dJyz83_0),.din(w_dff_A_AKEwKhuf3_0),.clk(gclk));
	jdff dff_A_vl5dJyz83_0(.dout(w_dff_A_ZOFqoI5P0_0),.din(w_dff_A_vl5dJyz83_0),.clk(gclk));
	jdff dff_A_ZOFqoI5P0_0(.dout(w_dff_A_iWxVOVxW1_0),.din(w_dff_A_ZOFqoI5P0_0),.clk(gclk));
	jdff dff_A_iWxVOVxW1_0(.dout(w_dff_A_ZvXdbyex2_0),.din(w_dff_A_iWxVOVxW1_0),.clk(gclk));
	jdff dff_A_ZvXdbyex2_0(.dout(w_dff_A_ZUObxu8A1_0),.din(w_dff_A_ZvXdbyex2_0),.clk(gclk));
	jdff dff_A_ZUObxu8A1_0(.dout(w_dff_A_mt7vBhuX3_0),.din(w_dff_A_ZUObxu8A1_0),.clk(gclk));
	jdff dff_A_mt7vBhuX3_0(.dout(w_dff_A_GVyWvK378_0),.din(w_dff_A_mt7vBhuX3_0),.clk(gclk));
	jdff dff_A_GVyWvK378_0(.dout(w_dff_A_yDVVGrpt7_0),.din(w_dff_A_GVyWvK378_0),.clk(gclk));
	jdff dff_A_yDVVGrpt7_0(.dout(w_dff_A_mpN0foaq8_0),.din(w_dff_A_yDVVGrpt7_0),.clk(gclk));
	jdff dff_A_mpN0foaq8_0(.dout(G447gat),.din(w_dff_A_mpN0foaq8_0),.clk(gclk));
	jdff dff_A_oCZBiHiG0_2(.dout(w_dff_A_2JERXUrB0_0),.din(w_dff_A_oCZBiHiG0_2),.clk(gclk));
	jdff dff_A_2JERXUrB0_0(.dout(w_dff_A_6NW6omcr6_0),.din(w_dff_A_2JERXUrB0_0),.clk(gclk));
	jdff dff_A_6NW6omcr6_0(.dout(w_dff_A_YHxMdtWv8_0),.din(w_dff_A_6NW6omcr6_0),.clk(gclk));
	jdff dff_A_YHxMdtWv8_0(.dout(w_dff_A_ic6tqCU62_0),.din(w_dff_A_YHxMdtWv8_0),.clk(gclk));
	jdff dff_A_ic6tqCU62_0(.dout(w_dff_A_kat0AlJe6_0),.din(w_dff_A_ic6tqCU62_0),.clk(gclk));
	jdff dff_A_kat0AlJe6_0(.dout(w_dff_A_wnUuWrXU7_0),.din(w_dff_A_kat0AlJe6_0),.clk(gclk));
	jdff dff_A_wnUuWrXU7_0(.dout(w_dff_A_KaCbYYrN1_0),.din(w_dff_A_wnUuWrXU7_0),.clk(gclk));
	jdff dff_A_KaCbYYrN1_0(.dout(w_dff_A_YPj9QUrI7_0),.din(w_dff_A_KaCbYYrN1_0),.clk(gclk));
	jdff dff_A_YPj9QUrI7_0(.dout(w_dff_A_QaQMfFeL1_0),.din(w_dff_A_YPj9QUrI7_0),.clk(gclk));
	jdff dff_A_QaQMfFeL1_0(.dout(w_dff_A_zJRYce1J2_0),.din(w_dff_A_QaQMfFeL1_0),.clk(gclk));
	jdff dff_A_zJRYce1J2_0(.dout(w_dff_A_dSx2ufSZ2_0),.din(w_dff_A_zJRYce1J2_0),.clk(gclk));
	jdff dff_A_dSx2ufSZ2_0(.dout(w_dff_A_CpT9y3rb1_0),.din(w_dff_A_dSx2ufSZ2_0),.clk(gclk));
	jdff dff_A_CpT9y3rb1_0(.dout(w_dff_A_Hiz2JChW3_0),.din(w_dff_A_CpT9y3rb1_0),.clk(gclk));
	jdff dff_A_Hiz2JChW3_0(.dout(w_dff_A_VjdYfxEZ5_0),.din(w_dff_A_Hiz2JChW3_0),.clk(gclk));
	jdff dff_A_VjdYfxEZ5_0(.dout(w_dff_A_1qbnn19P4_0),.din(w_dff_A_VjdYfxEZ5_0),.clk(gclk));
	jdff dff_A_1qbnn19P4_0(.dout(w_dff_A_oMvdRlKt5_0),.din(w_dff_A_1qbnn19P4_0),.clk(gclk));
	jdff dff_A_oMvdRlKt5_0(.dout(w_dff_A_1wbfVwSH9_0),.din(w_dff_A_oMvdRlKt5_0),.clk(gclk));
	jdff dff_A_1wbfVwSH9_0(.dout(w_dff_A_nL2ZaUsE8_0),.din(w_dff_A_1wbfVwSH9_0),.clk(gclk));
	jdff dff_A_nL2ZaUsE8_0(.dout(w_dff_A_bioNuumO7_0),.din(w_dff_A_nL2ZaUsE8_0),.clk(gclk));
	jdff dff_A_bioNuumO7_0(.dout(w_dff_A_bJw0UQ8m2_0),.din(w_dff_A_bioNuumO7_0),.clk(gclk));
	jdff dff_A_bJw0UQ8m2_0(.dout(w_dff_A_JFUxqJ0Y7_0),.din(w_dff_A_bJw0UQ8m2_0),.clk(gclk));
	jdff dff_A_JFUxqJ0Y7_0(.dout(w_dff_A_pNAFHhct9_0),.din(w_dff_A_JFUxqJ0Y7_0),.clk(gclk));
	jdff dff_A_pNAFHhct9_0(.dout(G448gat),.din(w_dff_A_pNAFHhct9_0),.clk(gclk));
	jdff dff_A_WQugsFuT0_2(.dout(w_dff_A_XTcE3euz8_0),.din(w_dff_A_WQugsFuT0_2),.clk(gclk));
	jdff dff_A_XTcE3euz8_0(.dout(w_dff_A_waGQQAOv1_0),.din(w_dff_A_XTcE3euz8_0),.clk(gclk));
	jdff dff_A_waGQQAOv1_0(.dout(w_dff_A_rv02eS0u7_0),.din(w_dff_A_waGQQAOv1_0),.clk(gclk));
	jdff dff_A_rv02eS0u7_0(.dout(w_dff_A_F259Dxet0_0),.din(w_dff_A_rv02eS0u7_0),.clk(gclk));
	jdff dff_A_F259Dxet0_0(.dout(w_dff_A_h86j0hNt3_0),.din(w_dff_A_F259Dxet0_0),.clk(gclk));
	jdff dff_A_h86j0hNt3_0(.dout(w_dff_A_J9igMIAL8_0),.din(w_dff_A_h86j0hNt3_0),.clk(gclk));
	jdff dff_A_J9igMIAL8_0(.dout(w_dff_A_QIz5LeYD6_0),.din(w_dff_A_J9igMIAL8_0),.clk(gclk));
	jdff dff_A_QIz5LeYD6_0(.dout(w_dff_A_u8g82CIV7_0),.din(w_dff_A_QIz5LeYD6_0),.clk(gclk));
	jdff dff_A_u8g82CIV7_0(.dout(w_dff_A_dAaxuK4I1_0),.din(w_dff_A_u8g82CIV7_0),.clk(gclk));
	jdff dff_A_dAaxuK4I1_0(.dout(w_dff_A_NijWWpc73_0),.din(w_dff_A_dAaxuK4I1_0),.clk(gclk));
	jdff dff_A_NijWWpc73_0(.dout(w_dff_A_xXt4BVmR5_0),.din(w_dff_A_NijWWpc73_0),.clk(gclk));
	jdff dff_A_xXt4BVmR5_0(.dout(w_dff_A_hTgsqFPi3_0),.din(w_dff_A_xXt4BVmR5_0),.clk(gclk));
	jdff dff_A_hTgsqFPi3_0(.dout(w_dff_A_rjO19pxN6_0),.din(w_dff_A_hTgsqFPi3_0),.clk(gclk));
	jdff dff_A_rjO19pxN6_0(.dout(w_dff_A_Fuo5gRsU8_0),.din(w_dff_A_rjO19pxN6_0),.clk(gclk));
	jdff dff_A_Fuo5gRsU8_0(.dout(w_dff_A_NvxyFkI47_0),.din(w_dff_A_Fuo5gRsU8_0),.clk(gclk));
	jdff dff_A_NvxyFkI47_0(.dout(w_dff_A_D7AgZQwK1_0),.din(w_dff_A_NvxyFkI47_0),.clk(gclk));
	jdff dff_A_D7AgZQwK1_0(.dout(w_dff_A_QmAyNK9p3_0),.din(w_dff_A_D7AgZQwK1_0),.clk(gclk));
	jdff dff_A_QmAyNK9p3_0(.dout(w_dff_A_eiV3VIfR3_0),.din(w_dff_A_QmAyNK9p3_0),.clk(gclk));
	jdff dff_A_eiV3VIfR3_0(.dout(w_dff_A_p4yhxYh72_0),.din(w_dff_A_eiV3VIfR3_0),.clk(gclk));
	jdff dff_A_p4yhxYh72_0(.dout(w_dff_A_NiUnCLL54_0),.din(w_dff_A_p4yhxYh72_0),.clk(gclk));
	jdff dff_A_NiUnCLL54_0(.dout(w_dff_A_Is1bllA11_0),.din(w_dff_A_NiUnCLL54_0),.clk(gclk));
	jdff dff_A_Is1bllA11_0(.dout(w_dff_A_OEwO9Xu70_0),.din(w_dff_A_Is1bllA11_0),.clk(gclk));
	jdff dff_A_OEwO9Xu70_0(.dout(G449gat),.din(w_dff_A_OEwO9Xu70_0),.clk(gclk));
	jdff dff_A_62IaO45P5_2(.dout(w_dff_A_ZxS6W6qB8_0),.din(w_dff_A_62IaO45P5_2),.clk(gclk));
	jdff dff_A_ZxS6W6qB8_0(.dout(w_dff_A_ug4qJM6l3_0),.din(w_dff_A_ZxS6W6qB8_0),.clk(gclk));
	jdff dff_A_ug4qJM6l3_0(.dout(w_dff_A_C7efjcvX5_0),.din(w_dff_A_ug4qJM6l3_0),.clk(gclk));
	jdff dff_A_C7efjcvX5_0(.dout(w_dff_A_u88nR0RM1_0),.din(w_dff_A_C7efjcvX5_0),.clk(gclk));
	jdff dff_A_u88nR0RM1_0(.dout(w_dff_A_KCv2dHGN0_0),.din(w_dff_A_u88nR0RM1_0),.clk(gclk));
	jdff dff_A_KCv2dHGN0_0(.dout(w_dff_A_UMGNC58v9_0),.din(w_dff_A_KCv2dHGN0_0),.clk(gclk));
	jdff dff_A_UMGNC58v9_0(.dout(w_dff_A_72BmfYVd6_0),.din(w_dff_A_UMGNC58v9_0),.clk(gclk));
	jdff dff_A_72BmfYVd6_0(.dout(w_dff_A_BQWGDUTw9_0),.din(w_dff_A_72BmfYVd6_0),.clk(gclk));
	jdff dff_A_BQWGDUTw9_0(.dout(w_dff_A_EIBhi0YZ6_0),.din(w_dff_A_BQWGDUTw9_0),.clk(gclk));
	jdff dff_A_EIBhi0YZ6_0(.dout(w_dff_A_5fbcAUl66_0),.din(w_dff_A_EIBhi0YZ6_0),.clk(gclk));
	jdff dff_A_5fbcAUl66_0(.dout(w_dff_A_ddkWoOpC0_0),.din(w_dff_A_5fbcAUl66_0),.clk(gclk));
	jdff dff_A_ddkWoOpC0_0(.dout(w_dff_A_vX8ioDB01_0),.din(w_dff_A_ddkWoOpC0_0),.clk(gclk));
	jdff dff_A_vX8ioDB01_0(.dout(w_dff_A_ka0TKRWq7_0),.din(w_dff_A_vX8ioDB01_0),.clk(gclk));
	jdff dff_A_ka0TKRWq7_0(.dout(w_dff_A_qOdIGPmS4_0),.din(w_dff_A_ka0TKRWq7_0),.clk(gclk));
	jdff dff_A_qOdIGPmS4_0(.dout(w_dff_A_Zt725Dud5_0),.din(w_dff_A_qOdIGPmS4_0),.clk(gclk));
	jdff dff_A_Zt725Dud5_0(.dout(w_dff_A_ZAMa8JRO3_0),.din(w_dff_A_Zt725Dud5_0),.clk(gclk));
	jdff dff_A_ZAMa8JRO3_0(.dout(w_dff_A_7ZsLcK9Y2_0),.din(w_dff_A_ZAMa8JRO3_0),.clk(gclk));
	jdff dff_A_7ZsLcK9Y2_0(.dout(w_dff_A_ICYRftez4_0),.din(w_dff_A_7ZsLcK9Y2_0),.clk(gclk));
	jdff dff_A_ICYRftez4_0(.dout(w_dff_A_ofPhop2v2_0),.din(w_dff_A_ICYRftez4_0),.clk(gclk));
	jdff dff_A_ofPhop2v2_0(.dout(w_dff_A_95AUTe252_0),.din(w_dff_A_ofPhop2v2_0),.clk(gclk));
	jdff dff_A_95AUTe252_0(.dout(w_dff_A_tCMNmrpR3_0),.din(w_dff_A_95AUTe252_0),.clk(gclk));
	jdff dff_A_tCMNmrpR3_0(.dout(w_dff_A_yk9RaUOh7_0),.din(w_dff_A_tCMNmrpR3_0),.clk(gclk));
	jdff dff_A_yk9RaUOh7_0(.dout(w_dff_A_0o7VBkEv9_0),.din(w_dff_A_yk9RaUOh7_0),.clk(gclk));
	jdff dff_A_0o7VBkEv9_0(.dout(w_dff_A_P26aDpeN7_0),.din(w_dff_A_0o7VBkEv9_0),.clk(gclk));
	jdff dff_A_P26aDpeN7_0(.dout(w_dff_A_VOorZblU0_0),.din(w_dff_A_P26aDpeN7_0),.clk(gclk));
	jdff dff_A_VOorZblU0_0(.dout(G450gat),.din(w_dff_A_VOorZblU0_0),.clk(gclk));
	jdff dff_A_OhvIt33J6_2(.dout(w_dff_A_AUMM5Vz60_0),.din(w_dff_A_OhvIt33J6_2),.clk(gclk));
	jdff dff_A_AUMM5Vz60_0(.dout(w_dff_A_MuCpLdEp1_0),.din(w_dff_A_AUMM5Vz60_0),.clk(gclk));
	jdff dff_A_MuCpLdEp1_0(.dout(w_dff_A_aRuHzX8a2_0),.din(w_dff_A_MuCpLdEp1_0),.clk(gclk));
	jdff dff_A_aRuHzX8a2_0(.dout(w_dff_A_NbCZVsyv7_0),.din(w_dff_A_aRuHzX8a2_0),.clk(gclk));
	jdff dff_A_NbCZVsyv7_0(.dout(w_dff_A_XTyI7J1O0_0),.din(w_dff_A_NbCZVsyv7_0),.clk(gclk));
	jdff dff_A_XTyI7J1O0_0(.dout(w_dff_A_yVaoSb9n5_0),.din(w_dff_A_XTyI7J1O0_0),.clk(gclk));
	jdff dff_A_yVaoSb9n5_0(.dout(w_dff_A_1k7aEVIY2_0),.din(w_dff_A_yVaoSb9n5_0),.clk(gclk));
	jdff dff_A_1k7aEVIY2_0(.dout(w_dff_A_LC6fSsxW5_0),.din(w_dff_A_1k7aEVIY2_0),.clk(gclk));
	jdff dff_A_LC6fSsxW5_0(.dout(w_dff_A_OVKzfKEI9_0),.din(w_dff_A_LC6fSsxW5_0),.clk(gclk));
	jdff dff_A_OVKzfKEI9_0(.dout(w_dff_A_wFtQ1NoB3_0),.din(w_dff_A_OVKzfKEI9_0),.clk(gclk));
	jdff dff_A_wFtQ1NoB3_0(.dout(w_dff_A_tUzFcp0y5_0),.din(w_dff_A_wFtQ1NoB3_0),.clk(gclk));
	jdff dff_A_tUzFcp0y5_0(.dout(w_dff_A_8eD8pS870_0),.din(w_dff_A_tUzFcp0y5_0),.clk(gclk));
	jdff dff_A_8eD8pS870_0(.dout(w_dff_A_hIljqn2Y2_0),.din(w_dff_A_8eD8pS870_0),.clk(gclk));
	jdff dff_A_hIljqn2Y2_0(.dout(w_dff_A_BK98MWIm0_0),.din(w_dff_A_hIljqn2Y2_0),.clk(gclk));
	jdff dff_A_BK98MWIm0_0(.dout(w_dff_A_0xWxjbdh4_0),.din(w_dff_A_BK98MWIm0_0),.clk(gclk));
	jdff dff_A_0xWxjbdh4_0(.dout(w_dff_A_0Zl1UtQM3_0),.din(w_dff_A_0xWxjbdh4_0),.clk(gclk));
	jdff dff_A_0Zl1UtQM3_0(.dout(w_dff_A_tvmBxap54_0),.din(w_dff_A_0Zl1UtQM3_0),.clk(gclk));
	jdff dff_A_tvmBxap54_0(.dout(w_dff_A_S3mzQaB14_0),.din(w_dff_A_tvmBxap54_0),.clk(gclk));
	jdff dff_A_S3mzQaB14_0(.dout(w_dff_A_g88LvIVh0_0),.din(w_dff_A_S3mzQaB14_0),.clk(gclk));
	jdff dff_A_g88LvIVh0_0(.dout(w_dff_A_tl4Y0fmj2_0),.din(w_dff_A_g88LvIVh0_0),.clk(gclk));
	jdff dff_A_tl4Y0fmj2_0(.dout(w_dff_A_mjJ7ijoY0_0),.din(w_dff_A_tl4Y0fmj2_0),.clk(gclk));
	jdff dff_A_mjJ7ijoY0_0(.dout(w_dff_A_hSRmfOOu2_0),.din(w_dff_A_mjJ7ijoY0_0),.clk(gclk));
	jdff dff_A_hSRmfOOu2_0(.dout(w_dff_A_oSEqh7DY6_0),.din(w_dff_A_hSRmfOOu2_0),.clk(gclk));
	jdff dff_A_oSEqh7DY6_0(.dout(G767gat),.din(w_dff_A_oSEqh7DY6_0),.clk(gclk));
	jdff dff_A_ijyXFBE84_2(.dout(w_dff_A_KuZ0yOuE6_0),.din(w_dff_A_ijyXFBE84_2),.clk(gclk));
	jdff dff_A_KuZ0yOuE6_0(.dout(w_dff_A_aAAvfzJ80_0),.din(w_dff_A_KuZ0yOuE6_0),.clk(gclk));
	jdff dff_A_aAAvfzJ80_0(.dout(w_dff_A_Pu6n5JId9_0),.din(w_dff_A_aAAvfzJ80_0),.clk(gclk));
	jdff dff_A_Pu6n5JId9_0(.dout(w_dff_A_AvgbYcVt5_0),.din(w_dff_A_Pu6n5JId9_0),.clk(gclk));
	jdff dff_A_AvgbYcVt5_0(.dout(w_dff_A_ZmfYtXFB7_0),.din(w_dff_A_AvgbYcVt5_0),.clk(gclk));
	jdff dff_A_ZmfYtXFB7_0(.dout(w_dff_A_Pg91RuED2_0),.din(w_dff_A_ZmfYtXFB7_0),.clk(gclk));
	jdff dff_A_Pg91RuED2_0(.dout(w_dff_A_rMGvYZY82_0),.din(w_dff_A_Pg91RuED2_0),.clk(gclk));
	jdff dff_A_rMGvYZY82_0(.dout(w_dff_A_tmntGwPz8_0),.din(w_dff_A_rMGvYZY82_0),.clk(gclk));
	jdff dff_A_tmntGwPz8_0(.dout(w_dff_A_CsS5h76y1_0),.din(w_dff_A_tmntGwPz8_0),.clk(gclk));
	jdff dff_A_CsS5h76y1_0(.dout(w_dff_A_mma5k4kX1_0),.din(w_dff_A_CsS5h76y1_0),.clk(gclk));
	jdff dff_A_mma5k4kX1_0(.dout(w_dff_A_BnO6ZzXq4_0),.din(w_dff_A_mma5k4kX1_0),.clk(gclk));
	jdff dff_A_BnO6ZzXq4_0(.dout(w_dff_A_mgCwxtpr3_0),.din(w_dff_A_BnO6ZzXq4_0),.clk(gclk));
	jdff dff_A_mgCwxtpr3_0(.dout(w_dff_A_rfpx7WkN7_0),.din(w_dff_A_mgCwxtpr3_0),.clk(gclk));
	jdff dff_A_rfpx7WkN7_0(.dout(w_dff_A_RW1mjh6D3_0),.din(w_dff_A_rfpx7WkN7_0),.clk(gclk));
	jdff dff_A_RW1mjh6D3_0(.dout(w_dff_A_qaVO5FQs0_0),.din(w_dff_A_RW1mjh6D3_0),.clk(gclk));
	jdff dff_A_qaVO5FQs0_0(.dout(w_dff_A_crGx4l1H3_0),.din(w_dff_A_qaVO5FQs0_0),.clk(gclk));
	jdff dff_A_crGx4l1H3_0(.dout(w_dff_A_vUx8xaFD1_0),.din(w_dff_A_crGx4l1H3_0),.clk(gclk));
	jdff dff_A_vUx8xaFD1_0(.dout(w_dff_A_gciaVF359_0),.din(w_dff_A_vUx8xaFD1_0),.clk(gclk));
	jdff dff_A_gciaVF359_0(.dout(w_dff_A_HYVAJKsk6_0),.din(w_dff_A_gciaVF359_0),.clk(gclk));
	jdff dff_A_HYVAJKsk6_0(.dout(w_dff_A_UJnDelxg1_0),.din(w_dff_A_HYVAJKsk6_0),.clk(gclk));
	jdff dff_A_UJnDelxg1_0(.dout(w_dff_A_YKWzR1UF5_0),.din(w_dff_A_UJnDelxg1_0),.clk(gclk));
	jdff dff_A_YKWzR1UF5_0(.dout(w_dff_A_FWpgesYV0_0),.din(w_dff_A_YKWzR1UF5_0),.clk(gclk));
	jdff dff_A_FWpgesYV0_0(.dout(w_dff_A_LmQboStI7_0),.din(w_dff_A_FWpgesYV0_0),.clk(gclk));
	jdff dff_A_LmQboStI7_0(.dout(G768gat),.din(w_dff_A_LmQboStI7_0),.clk(gclk));
	jdff dff_A_nh87JbUt4_2(.dout(w_dff_A_3HWwNyCh1_0),.din(w_dff_A_nh87JbUt4_2),.clk(gclk));
	jdff dff_A_3HWwNyCh1_0(.dout(w_dff_A_8ewzlnrw4_0),.din(w_dff_A_3HWwNyCh1_0),.clk(gclk));
	jdff dff_A_8ewzlnrw4_0(.dout(w_dff_A_szbM88Hs5_0),.din(w_dff_A_8ewzlnrw4_0),.clk(gclk));
	jdff dff_A_szbM88Hs5_0(.dout(w_dff_A_hh9atL544_0),.din(w_dff_A_szbM88Hs5_0),.clk(gclk));
	jdff dff_A_hh9atL544_0(.dout(w_dff_A_Iw8W4qYS5_0),.din(w_dff_A_hh9atL544_0),.clk(gclk));
	jdff dff_A_Iw8W4qYS5_0(.dout(w_dff_A_sk0xNoWH7_0),.din(w_dff_A_Iw8W4qYS5_0),.clk(gclk));
	jdff dff_A_sk0xNoWH7_0(.dout(w_dff_A_0FE8NSYg9_0),.din(w_dff_A_sk0xNoWH7_0),.clk(gclk));
	jdff dff_A_0FE8NSYg9_0(.dout(w_dff_A_5KektUN41_0),.din(w_dff_A_0FE8NSYg9_0),.clk(gclk));
	jdff dff_A_5KektUN41_0(.dout(w_dff_A_DiP8ilzB0_0),.din(w_dff_A_5KektUN41_0),.clk(gclk));
	jdff dff_A_DiP8ilzB0_0(.dout(w_dff_A_EOaVoLqy9_0),.din(w_dff_A_DiP8ilzB0_0),.clk(gclk));
	jdff dff_A_EOaVoLqy9_0(.dout(w_dff_A_VM7UAmMV3_0),.din(w_dff_A_EOaVoLqy9_0),.clk(gclk));
	jdff dff_A_VM7UAmMV3_0(.dout(w_dff_A_77IM1GqG4_0),.din(w_dff_A_VM7UAmMV3_0),.clk(gclk));
	jdff dff_A_77IM1GqG4_0(.dout(G850gat),.din(w_dff_A_77IM1GqG4_0),.clk(gclk));
	jdff dff_A_83XL4cAE0_2(.dout(w_dff_A_bpe8gIj91_0),.din(w_dff_A_83XL4cAE0_2),.clk(gclk));
	jdff dff_A_bpe8gIj91_0(.dout(w_dff_A_We2goBjS7_0),.din(w_dff_A_bpe8gIj91_0),.clk(gclk));
	jdff dff_A_We2goBjS7_0(.dout(w_dff_A_JsLojnvW6_0),.din(w_dff_A_We2goBjS7_0),.clk(gclk));
	jdff dff_A_JsLojnvW6_0(.dout(w_dff_A_GFVDQyAf8_0),.din(w_dff_A_JsLojnvW6_0),.clk(gclk));
	jdff dff_A_GFVDQyAf8_0(.dout(w_dff_A_SOw645RN6_0),.din(w_dff_A_GFVDQyAf8_0),.clk(gclk));
	jdff dff_A_SOw645RN6_0(.dout(w_dff_A_rjOJlnYr7_0),.din(w_dff_A_SOw645RN6_0),.clk(gclk));
	jdff dff_A_rjOJlnYr7_0(.dout(w_dff_A_SNdymnnu5_0),.din(w_dff_A_rjOJlnYr7_0),.clk(gclk));
	jdff dff_A_SNdymnnu5_0(.dout(G863gat),.din(w_dff_A_SNdymnnu5_0),.clk(gclk));
	jdff dff_A_QaPWEmmy9_2(.dout(w_dff_A_ValFc8q85_0),.din(w_dff_A_QaPWEmmy9_2),.clk(gclk));
	jdff dff_A_ValFc8q85_0(.dout(w_dff_A_kUTamCJQ5_0),.din(w_dff_A_ValFc8q85_0),.clk(gclk));
	jdff dff_A_kUTamCJQ5_0(.dout(w_dff_A_yxO3DTUZ5_0),.din(w_dff_A_kUTamCJQ5_0),.clk(gclk));
	jdff dff_A_yxO3DTUZ5_0(.dout(w_dff_A_ZzVYyaWT0_0),.din(w_dff_A_yxO3DTUZ5_0),.clk(gclk));
	jdff dff_A_ZzVYyaWT0_0(.dout(w_dff_A_A8IE8g3U1_0),.din(w_dff_A_ZzVYyaWT0_0),.clk(gclk));
	jdff dff_A_A8IE8g3U1_0(.dout(w_dff_A_bXBWkxwt4_0),.din(w_dff_A_A8IE8g3U1_0),.clk(gclk));
	jdff dff_A_bXBWkxwt4_0(.dout(w_dff_A_VXM6wOLH7_0),.din(w_dff_A_bXBWkxwt4_0),.clk(gclk));
	jdff dff_A_VXM6wOLH7_0(.dout(w_dff_A_cyP2e2Cq8_0),.din(w_dff_A_VXM6wOLH7_0),.clk(gclk));
	jdff dff_A_cyP2e2Cq8_0(.dout(w_dff_A_3qCCnxzi9_0),.din(w_dff_A_cyP2e2Cq8_0),.clk(gclk));
	jdff dff_A_3qCCnxzi9_0(.dout(G864gat),.din(w_dff_A_3qCCnxzi9_0),.clk(gclk));
	jdff dff_A_KtnSHZjt1_2(.dout(w_dff_A_eiJRXx2o6_0),.din(w_dff_A_KtnSHZjt1_2),.clk(gclk));
	jdff dff_A_eiJRXx2o6_0(.dout(w_dff_A_TmawjQ0z0_0),.din(w_dff_A_eiJRXx2o6_0),.clk(gclk));
	jdff dff_A_TmawjQ0z0_0(.dout(w_dff_A_wfClqdcP7_0),.din(w_dff_A_TmawjQ0z0_0),.clk(gclk));
	jdff dff_A_wfClqdcP7_0(.dout(w_dff_A_bLZCEdsN7_0),.din(w_dff_A_wfClqdcP7_0),.clk(gclk));
	jdff dff_A_bLZCEdsN7_0(.dout(w_dff_A_KUE60uwm4_0),.din(w_dff_A_bLZCEdsN7_0),.clk(gclk));
	jdff dff_A_KUE60uwm4_0(.dout(w_dff_A_e5xMsPhh0_0),.din(w_dff_A_KUE60uwm4_0),.clk(gclk));
	jdff dff_A_e5xMsPhh0_0(.dout(w_dff_A_ZksiIyXT7_0),.din(w_dff_A_e5xMsPhh0_0),.clk(gclk));
	jdff dff_A_ZksiIyXT7_0(.dout(w_dff_A_qif6j39L7_0),.din(w_dff_A_ZksiIyXT7_0),.clk(gclk));
	jdff dff_A_qif6j39L7_0(.dout(w_dff_A_470sFp8E4_0),.din(w_dff_A_qif6j39L7_0),.clk(gclk));
	jdff dff_A_470sFp8E4_0(.dout(w_dff_A_a42W2vVw9_0),.din(w_dff_A_470sFp8E4_0),.clk(gclk));
	jdff dff_A_a42W2vVw9_0(.dout(w_dff_A_fbA61J2w0_0),.din(w_dff_A_a42W2vVw9_0),.clk(gclk));
	jdff dff_A_fbA61J2w0_0(.dout(G865gat),.din(w_dff_A_fbA61J2w0_0),.clk(gclk));
	jdff dff_A_lxhkViEa1_2(.dout(w_dff_A_c67N0HXi9_0),.din(w_dff_A_lxhkViEa1_2),.clk(gclk));
	jdff dff_A_c67N0HXi9_0(.dout(G866gat),.din(w_dff_A_c67N0HXi9_0),.clk(gclk));
	jdff dff_A_L5KrTId14_2(.dout(w_dff_A_x0qGp2kE0_0),.din(w_dff_A_L5KrTId14_2),.clk(gclk));
	jdff dff_A_x0qGp2kE0_0(.dout(w_dff_A_stx7Dq2G1_0),.din(w_dff_A_x0qGp2kE0_0),.clk(gclk));
	jdff dff_A_stx7Dq2G1_0(.dout(w_dff_A_EkudcTpl9_0),.din(w_dff_A_stx7Dq2G1_0),.clk(gclk));
	jdff dff_A_EkudcTpl9_0(.dout(w_dff_A_1zwzZJkW2_0),.din(w_dff_A_EkudcTpl9_0),.clk(gclk));
	jdff dff_A_1zwzZJkW2_0(.dout(G874gat),.din(w_dff_A_1zwzZJkW2_0),.clk(gclk));
	jdff dff_A_wWIeNAhW9_2(.dout(w_dff_A_rijtXIGe1_0),.din(w_dff_A_wWIeNAhW9_2),.clk(gclk));
	jdff dff_A_rijtXIGe1_0(.dout(G879gat),.din(w_dff_A_rijtXIGe1_0),.clk(gclk));
	jdff dff_A_vX37Lua63_2(.dout(w_dff_A_Txp4bkph8_0),.din(w_dff_A_vX37Lua63_2),.clk(gclk));
	jdff dff_A_Txp4bkph8_0(.dout(w_dff_A_3hVaVjDW6_0),.din(w_dff_A_Txp4bkph8_0),.clk(gclk));
	jdff dff_A_3hVaVjDW6_0(.dout(w_dff_A_vla4J1i82_0),.din(w_dff_A_3hVaVjDW6_0),.clk(gclk));
	jdff dff_A_vla4J1i82_0(.dout(G880gat),.din(w_dff_A_vla4J1i82_0),.clk(gclk));
endmodule

