/*

c6288:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jdff: 8046
	jand: 664
	jor: 312

Summary:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jdff: 8046
	jand: 664
	jor: 312
*/

module c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G1gat_1;
	wire[2:0] w_G1gat_2;
	wire[2:0] w_G1gat_3;
	wire[2:0] w_G1gat_4;
	wire[2:0] w_G1gat_5;
	wire[2:0] w_G1gat_6;
	wire[1:0] w_G1gat_7;
	wire[2:0] w_G18gat_0;
	wire[2:0] w_G18gat_1;
	wire[2:0] w_G18gat_2;
	wire[2:0] w_G18gat_3;
	wire[2:0] w_G18gat_4;
	wire[2:0] w_G18gat_5;
	wire[2:0] w_G18gat_6;
	wire[1:0] w_G18gat_7;
	wire[2:0] w_G35gat_0;
	wire[2:0] w_G35gat_1;
	wire[2:0] w_G35gat_2;
	wire[2:0] w_G35gat_3;
	wire[2:0] w_G35gat_4;
	wire[2:0] w_G35gat_5;
	wire[2:0] w_G35gat_6;
	wire[2:0] w_G35gat_7;
	wire[2:0] w_G52gat_0;
	wire[2:0] w_G52gat_1;
	wire[2:0] w_G52gat_2;
	wire[2:0] w_G52gat_3;
	wire[2:0] w_G52gat_4;
	wire[2:0] w_G52gat_5;
	wire[2:0] w_G52gat_6;
	wire[2:0] w_G52gat_7;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G69gat_1;
	wire[2:0] w_G69gat_2;
	wire[2:0] w_G69gat_3;
	wire[2:0] w_G69gat_4;
	wire[2:0] w_G69gat_5;
	wire[2:0] w_G69gat_6;
	wire[1:0] w_G69gat_7;
	wire[2:0] w_G86gat_0;
	wire[2:0] w_G86gat_1;
	wire[2:0] w_G86gat_2;
	wire[2:0] w_G86gat_3;
	wire[2:0] w_G86gat_4;
	wire[2:0] w_G86gat_5;
	wire[2:0] w_G86gat_6;
	wire[1:0] w_G86gat_7;
	wire[2:0] w_G103gat_0;
	wire[2:0] w_G103gat_1;
	wire[2:0] w_G103gat_2;
	wire[2:0] w_G103gat_3;
	wire[2:0] w_G103gat_4;
	wire[2:0] w_G103gat_5;
	wire[2:0] w_G103gat_6;
	wire[1:0] w_G103gat_7;
	wire[2:0] w_G120gat_0;
	wire[2:0] w_G120gat_1;
	wire[2:0] w_G120gat_2;
	wire[2:0] w_G120gat_3;
	wire[2:0] w_G120gat_4;
	wire[2:0] w_G120gat_5;
	wire[2:0] w_G120gat_6;
	wire[1:0] w_G120gat_7;
	wire[2:0] w_G137gat_0;
	wire[2:0] w_G137gat_1;
	wire[2:0] w_G137gat_2;
	wire[2:0] w_G137gat_3;
	wire[2:0] w_G137gat_4;
	wire[2:0] w_G137gat_5;
	wire[2:0] w_G137gat_6;
	wire[1:0] w_G137gat_7;
	wire[2:0] w_G154gat_0;
	wire[2:0] w_G154gat_1;
	wire[2:0] w_G154gat_2;
	wire[2:0] w_G154gat_3;
	wire[2:0] w_G154gat_4;
	wire[2:0] w_G154gat_5;
	wire[2:0] w_G154gat_6;
	wire[1:0] w_G154gat_7;
	wire[2:0] w_G171gat_0;
	wire[2:0] w_G171gat_1;
	wire[2:0] w_G171gat_2;
	wire[2:0] w_G171gat_3;
	wire[2:0] w_G171gat_4;
	wire[2:0] w_G171gat_5;
	wire[2:0] w_G171gat_6;
	wire[1:0] w_G171gat_7;
	wire[2:0] w_G188gat_0;
	wire[2:0] w_G188gat_1;
	wire[2:0] w_G188gat_2;
	wire[2:0] w_G188gat_3;
	wire[2:0] w_G188gat_4;
	wire[2:0] w_G188gat_5;
	wire[2:0] w_G188gat_6;
	wire[1:0] w_G188gat_7;
	wire[2:0] w_G205gat_0;
	wire[2:0] w_G205gat_1;
	wire[2:0] w_G205gat_2;
	wire[2:0] w_G205gat_3;
	wire[2:0] w_G205gat_4;
	wire[2:0] w_G205gat_5;
	wire[2:0] w_G205gat_6;
	wire[1:0] w_G205gat_7;
	wire[2:0] w_G222gat_0;
	wire[2:0] w_G222gat_1;
	wire[2:0] w_G222gat_2;
	wire[2:0] w_G222gat_3;
	wire[2:0] w_G222gat_4;
	wire[2:0] w_G222gat_5;
	wire[2:0] w_G222gat_6;
	wire[1:0] w_G222gat_7;
	wire[2:0] w_G239gat_0;
	wire[2:0] w_G239gat_1;
	wire[2:0] w_G239gat_2;
	wire[2:0] w_G239gat_3;
	wire[2:0] w_G239gat_4;
	wire[2:0] w_G239gat_5;
	wire[2:0] w_G239gat_6;
	wire[1:0] w_G239gat_7;
	wire[2:0] w_G256gat_0;
	wire[2:0] w_G256gat_1;
	wire[2:0] w_G256gat_2;
	wire[2:0] w_G256gat_3;
	wire[2:0] w_G256gat_4;
	wire[2:0] w_G256gat_5;
	wire[2:0] w_G256gat_6;
	wire[1:0] w_G256gat_7;
	wire[2:0] w_G273gat_0;
	wire[2:0] w_G273gat_1;
	wire[2:0] w_G273gat_2;
	wire[2:0] w_G273gat_3;
	wire[2:0] w_G273gat_4;
	wire[2:0] w_G273gat_5;
	wire[2:0] w_G273gat_6;
	wire[1:0] w_G273gat_7;
	wire[2:0] w_G290gat_0;
	wire[2:0] w_G290gat_1;
	wire[2:0] w_G290gat_2;
	wire[2:0] w_G290gat_3;
	wire[2:0] w_G290gat_4;
	wire[2:0] w_G290gat_5;
	wire[2:0] w_G290gat_6;
	wire[2:0] w_G290gat_7;
	wire[2:0] w_G307gat_0;
	wire[2:0] w_G307gat_1;
	wire[2:0] w_G307gat_2;
	wire[2:0] w_G307gat_3;
	wire[2:0] w_G307gat_4;
	wire[2:0] w_G307gat_5;
	wire[2:0] w_G307gat_6;
	wire[1:0] w_G307gat_7;
	wire[2:0] w_G324gat_0;
	wire[2:0] w_G324gat_1;
	wire[2:0] w_G324gat_2;
	wire[2:0] w_G324gat_3;
	wire[2:0] w_G324gat_4;
	wire[2:0] w_G324gat_5;
	wire[2:0] w_G324gat_6;
	wire[1:0] w_G324gat_7;
	wire[2:0] w_G341gat_0;
	wire[2:0] w_G341gat_1;
	wire[2:0] w_G341gat_2;
	wire[2:0] w_G341gat_3;
	wire[2:0] w_G341gat_4;
	wire[2:0] w_G341gat_5;
	wire[2:0] w_G341gat_6;
	wire[1:0] w_G341gat_7;
	wire[2:0] w_G358gat_0;
	wire[2:0] w_G358gat_1;
	wire[2:0] w_G358gat_2;
	wire[2:0] w_G358gat_3;
	wire[2:0] w_G358gat_4;
	wire[2:0] w_G358gat_5;
	wire[2:0] w_G358gat_6;
	wire[1:0] w_G358gat_7;
	wire[2:0] w_G375gat_0;
	wire[2:0] w_G375gat_1;
	wire[2:0] w_G375gat_2;
	wire[2:0] w_G375gat_3;
	wire[2:0] w_G375gat_4;
	wire[2:0] w_G375gat_5;
	wire[2:0] w_G375gat_6;
	wire[1:0] w_G375gat_7;
	wire[2:0] w_G392gat_0;
	wire[2:0] w_G392gat_1;
	wire[2:0] w_G392gat_2;
	wire[2:0] w_G392gat_3;
	wire[2:0] w_G392gat_4;
	wire[2:0] w_G392gat_5;
	wire[2:0] w_G392gat_6;
	wire[1:0] w_G392gat_7;
	wire[2:0] w_G409gat_0;
	wire[2:0] w_G409gat_1;
	wire[2:0] w_G409gat_2;
	wire[2:0] w_G409gat_3;
	wire[2:0] w_G409gat_4;
	wire[2:0] w_G409gat_5;
	wire[2:0] w_G409gat_6;
	wire[1:0] w_G409gat_7;
	wire[2:0] w_G426gat_0;
	wire[2:0] w_G426gat_1;
	wire[2:0] w_G426gat_2;
	wire[2:0] w_G426gat_3;
	wire[2:0] w_G426gat_4;
	wire[2:0] w_G426gat_5;
	wire[2:0] w_G426gat_6;
	wire[1:0] w_G426gat_7;
	wire[2:0] w_G443gat_0;
	wire[2:0] w_G443gat_1;
	wire[2:0] w_G443gat_2;
	wire[2:0] w_G443gat_3;
	wire[2:0] w_G443gat_4;
	wire[2:0] w_G443gat_5;
	wire[2:0] w_G443gat_6;
	wire[1:0] w_G443gat_7;
	wire[2:0] w_G460gat_0;
	wire[2:0] w_G460gat_1;
	wire[2:0] w_G460gat_2;
	wire[2:0] w_G460gat_3;
	wire[2:0] w_G460gat_4;
	wire[2:0] w_G460gat_5;
	wire[2:0] w_G460gat_6;
	wire[1:0] w_G460gat_7;
	wire[2:0] w_G477gat_0;
	wire[2:0] w_G477gat_1;
	wire[2:0] w_G477gat_2;
	wire[2:0] w_G477gat_3;
	wire[2:0] w_G477gat_4;
	wire[2:0] w_G477gat_5;
	wire[2:0] w_G477gat_6;
	wire[1:0] w_G477gat_7;
	wire[2:0] w_G494gat_0;
	wire[2:0] w_G494gat_1;
	wire[2:0] w_G494gat_2;
	wire[2:0] w_G494gat_3;
	wire[2:0] w_G494gat_4;
	wire[2:0] w_G494gat_5;
	wire[2:0] w_G494gat_6;
	wire[1:0] w_G494gat_7;
	wire[2:0] w_G511gat_0;
	wire[2:0] w_G511gat_1;
	wire[2:0] w_G511gat_2;
	wire[2:0] w_G511gat_3;
	wire[2:0] w_G511gat_4;
	wire[2:0] w_G511gat_5;
	wire[2:0] w_G511gat_6;
	wire[1:0] w_G511gat_7;
	wire[2:0] w_G528gat_0;
	wire[2:0] w_G528gat_1;
	wire[2:0] w_G528gat_2;
	wire[2:0] w_G528gat_3;
	wire[2:0] w_G528gat_4;
	wire[2:0] w_G528gat_5;
	wire[2:0] w_G528gat_6;
	wire[1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire[1:0] w_n65_0;
	wire[1:0] w_n66_0;
	wire[1:0] w_n67_0;
	wire[1:0] w_n69_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n75_0;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[2:0] w_n80_0;
	wire[1:0] w_n83_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[1:0] w_n90_0;
	wire[1:0] w_n91_0;
	wire[1:0] w_n93_0;
	wire[1:0] w_n97_0;
	wire[1:0] w_n99_0;
	wire[2:0] w_n101_0;
	wire[1:0] w_n103_0;
	wire[1:0] w_n104_0;
	wire[1:0] w_n106_0;
	wire[1:0] w_n111_0;
	wire[1:0] w_n112_0;
	wire[2:0] w_n117_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[1:0] w_n121_0;
	wire[1:0] w_n122_0;
	wire[1:0] w_n123_0;
	wire[1:0] w_n125_0;
	wire[1:0] w_n127_0;
	wire[1:0] w_n128_0;
	wire[1:0] w_n129_0;
	wire[1:0] w_n130_0;
	wire[1:0] w_n132_0;
	wire[1:0] w_n133_0;
	wire[1:0] w_n135_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n141_0;
	wire[2:0] w_n146_0;
	wire[1:0] w_n148_0;
	wire[1:0] w_n152_0;
	wire[1:0] w_n154_0;
	wire[1:0] w_n155_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n157_0;
	wire[1:0] w_n158_0;
	wire[1:0] w_n160_0;
	wire[1:0] w_n161_0;
	wire[1:0] w_n162_0;
	wire[1:0] w_n163_0;
	wire[1:0] w_n164_0;
	wire[1:0] w_n165_0;
	wire[1:0] w_n167_0;
	wire[1:0] w_n168_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n175_0;
	wire[1:0] w_n176_0;
	wire[2:0] w_n181_0;
	wire[1:0] w_n183_0;
	wire[1:0] w_n186_0;
	wire[1:0] w_n188_0;
	wire[1:0] w_n192_0;
	wire[1:0] w_n194_0;
	wire[1:0] w_n195_0;
	wire[2:0] w_n196_0;
	wire[1:0] w_n198_0;
	wire[1:0] w_n200_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n202_0;
	wire[1:0] w_n203_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n205_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n207_0;
	wire[1:0] w_n209_0;
	wire[1:0] w_n210_0;
	wire[1:0] w_n212_0;
	wire[1:0] w_n217_0;
	wire[1:0] w_n218_0;
	wire[2:0] w_n223_0;
	wire[1:0] w_n225_0;
	wire[1:0] w_n228_0;
	wire[1:0] w_n230_0;
	wire[1:0] w_n233_0;
	wire[1:0] w_n235_0;
	wire[1:0] w_n239_0;
	wire[1:0] w_n241_0;
	wire[1:0] w_n242_0;
	wire[2:0] w_n243_0;
	wire[1:0] w_n245_0;
	wire[1:0] w_n247_0;
	wire[1:0] w_n248_0;
	wire[1:0] w_n249_0;
	wire[1:0] w_n250_0;
	wire[1:0] w_n251_0;
	wire[1:0] w_n252_0;
	wire[1:0] w_n253_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n255_0;
	wire[1:0] w_n256_0;
	wire[1:0] w_n258_0;
	wire[1:0] w_n259_0;
	wire[1:0] w_n261_0;
	wire[1:0] w_n266_0;
	wire[1:0] w_n267_0;
	wire[2:0] w_n272_0;
	wire[1:0] w_n274_0;
	wire[1:0] w_n277_0;
	wire[1:0] w_n279_0;
	wire[1:0] w_n282_0;
	wire[1:0] w_n284_0;
	wire[1:0] w_n287_0;
	wire[1:0] w_n289_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n295_0;
	wire[1:0] w_n296_0;
	wire[2:0] w_n297_0;
	wire[1:0] w_n299_0;
	wire[1:0] w_n301_0;
	wire[1:0] w_n302_0;
	wire[1:0] w_n303_0;
	wire[1:0] w_n304_0;
	wire[1:0] w_n305_0;
	wire[1:0] w_n306_0;
	wire[1:0] w_n307_0;
	wire[1:0] w_n308_0;
	wire[1:0] w_n309_0;
	wire[1:0] w_n310_0;
	wire[1:0] w_n311_0;
	wire[1:0] w_n312_0;
	wire[1:0] w_n314_0;
	wire[1:0] w_n315_0;
	wire[1:0] w_n317_0;
	wire[1:0] w_n322_0;
	wire[1:0] w_n323_0;
	wire[2:0] w_n328_0;
	wire[1:0] w_n330_0;
	wire[1:0] w_n333_0;
	wire[1:0] w_n335_0;
	wire[1:0] w_n338_0;
	wire[1:0] w_n340_0;
	wire[1:0] w_n343_0;
	wire[1:0] w_n345_0;
	wire[1:0] w_n348_0;
	wire[1:0] w_n350_0;
	wire[1:0] w_n354_0;
	wire[1:0] w_n356_0;
	wire[1:0] w_n357_0;
	wire[2:0] w_n358_0;
	wire[1:0] w_n360_0;
	wire[1:0] w_n362_0;
	wire[1:0] w_n363_0;
	wire[1:0] w_n364_0;
	wire[1:0] w_n365_0;
	wire[1:0] w_n366_0;
	wire[1:0] w_n367_0;
	wire[1:0] w_n368_0;
	wire[1:0] w_n369_0;
	wire[1:0] w_n370_0;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n373_0;
	wire[1:0] w_n374_0;
	wire[1:0] w_n375_0;
	wire[1:0] w_n377_0;
	wire[1:0] w_n378_0;
	wire[1:0] w_n380_0;
	wire[1:0] w_n385_0;
	wire[1:0] w_n386_0;
	wire[2:0] w_n391_0;
	wire[1:0] w_n393_0;
	wire[1:0] w_n396_0;
	wire[1:0] w_n398_0;
	wire[1:0] w_n401_0;
	wire[1:0] w_n403_0;
	wire[1:0] w_n406_0;
	wire[1:0] w_n408_0;
	wire[1:0] w_n411_0;
	wire[1:0] w_n413_0;
	wire[1:0] w_n416_0;
	wire[1:0] w_n418_0;
	wire[1:0] w_n423_0;
	wire[1:0] w_n425_0;
	wire[1:0] w_n426_0;
	wire[2:0] w_n427_0;
	wire[1:0] w_n429_0;
	wire[1:0] w_n431_0;
	wire[1:0] w_n432_0;
	wire[1:0] w_n433_0;
	wire[1:0] w_n434_0;
	wire[1:0] w_n435_0;
	wire[1:0] w_n436_0;
	wire[1:0] w_n437_0;
	wire[1:0] w_n438_0;
	wire[1:0] w_n439_0;
	wire[1:0] w_n440_0;
	wire[1:0] w_n441_0;
	wire[1:0] w_n442_0;
	wire[1:0] w_n443_0;
	wire[1:0] w_n444_0;
	wire[1:0] w_n445_0;
	wire[1:0] w_n446_0;
	wire[1:0] w_n448_0;
	wire[1:0] w_n449_0;
	wire[1:0] w_n451_0;
	wire[1:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[2:0] w_n462_0;
	wire[1:0] w_n464_0;
	wire[1:0] w_n467_0;
	wire[1:0] w_n469_0;
	wire[1:0] w_n472_0;
	wire[1:0] w_n474_0;
	wire[1:0] w_n477_0;
	wire[1:0] w_n479_0;
	wire[1:0] w_n482_0;
	wire[1:0] w_n484_0;
	wire[1:0] w_n487_0;
	wire[1:0] w_n489_0;
	wire[1:0] w_n492_0;
	wire[1:0] w_n494_0;
	wire[1:0] w_n499_0;
	wire[1:0] w_n501_0;
	wire[1:0] w_n502_0;
	wire[2:0] w_n503_0;
	wire[1:0] w_n505_0;
	wire[1:0] w_n507_0;
	wire[1:0] w_n508_0;
	wire[1:0] w_n509_0;
	wire[1:0] w_n510_0;
	wire[1:0] w_n511_0;
	wire[1:0] w_n512_0;
	wire[1:0] w_n513_0;
	wire[1:0] w_n514_0;
	wire[1:0] w_n515_0;
	wire[1:0] w_n516_0;
	wire[1:0] w_n517_0;
	wire[1:0] w_n518_0;
	wire[1:0] w_n519_0;
	wire[1:0] w_n520_0;
	wire[1:0] w_n521_0;
	wire[1:0] w_n522_0;
	wire[1:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n526_0;
	wire[1:0] w_n527_0;
	wire[1:0] w_n529_0;
	wire[1:0] w_n534_0;
	wire[1:0] w_n535_0;
	wire[2:0] w_n540_0;
	wire[1:0] w_n542_0;
	wire[1:0] w_n545_0;
	wire[1:0] w_n547_0;
	wire[1:0] w_n550_0;
	wire[1:0] w_n552_0;
	wire[1:0] w_n555_0;
	wire[1:0] w_n557_0;
	wire[1:0] w_n560_0;
	wire[1:0] w_n562_0;
	wire[1:0] w_n565_0;
	wire[1:0] w_n567_0;
	wire[1:0] w_n570_0;
	wire[1:0] w_n572_0;
	wire[1:0] w_n575_0;
	wire[1:0] w_n577_0;
	wire[1:0] w_n582_0;
	wire[1:0] w_n584_0;
	wire[1:0] w_n585_0;
	wire[2:0] w_n586_0;
	wire[1:0] w_n588_0;
	wire[1:0] w_n590_0;
	wire[1:0] w_n591_0;
	wire[1:0] w_n592_0;
	wire[1:0] w_n593_0;
	wire[1:0] w_n594_0;
	wire[1:0] w_n595_0;
	wire[1:0] w_n596_0;
	wire[1:0] w_n597_0;
	wire[1:0] w_n598_0;
	wire[1:0] w_n599_0;
	wire[1:0] w_n600_0;
	wire[1:0] w_n601_0;
	wire[1:0] w_n602_0;
	wire[1:0] w_n603_0;
	wire[1:0] w_n604_0;
	wire[1:0] w_n605_0;
	wire[1:0] w_n606_0;
	wire[1:0] w_n607_0;
	wire[1:0] w_n608_0;
	wire[1:0] w_n609_0;
	wire[1:0] w_n611_0;
	wire[1:0] w_n612_0;
	wire[1:0] w_n614_0;
	wire[1:0] w_n619_0;
	wire[1:0] w_n620_0;
	wire[2:0] w_n625_0;
	wire[1:0] w_n627_0;
	wire[1:0] w_n630_0;
	wire[1:0] w_n632_0;
	wire[1:0] w_n635_0;
	wire[1:0] w_n637_0;
	wire[1:0] w_n640_0;
	wire[1:0] w_n642_0;
	wire[1:0] w_n645_0;
	wire[1:0] w_n647_0;
	wire[1:0] w_n650_0;
	wire[1:0] w_n652_0;
	wire[1:0] w_n655_0;
	wire[1:0] w_n657_0;
	wire[1:0] w_n660_0;
	wire[1:0] w_n662_0;
	wire[1:0] w_n665_0;
	wire[1:0] w_n667_0;
	wire[1:0] w_n672_0;
	wire[1:0] w_n674_0;
	wire[1:0] w_n675_0;
	wire[2:0] w_n676_0;
	wire[1:0] w_n678_0;
	wire[1:0] w_n680_0;
	wire[1:0] w_n681_0;
	wire[1:0] w_n682_0;
	wire[1:0] w_n683_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n685_0;
	wire[1:0] w_n686_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n688_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n691_0;
	wire[1:0] w_n692_0;
	wire[1:0] w_n693_0;
	wire[1:0] w_n694_0;
	wire[1:0] w_n695_0;
	wire[1:0] w_n696_0;
	wire[1:0] w_n697_0;
	wire[1:0] w_n698_0;
	wire[1:0] w_n699_0;
	wire[1:0] w_n700_0;
	wire[1:0] w_n701_0;
	wire[1:0] w_n703_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n706_0;
	wire[1:0] w_n711_0;
	wire[1:0] w_n712_0;
	wire[2:0] w_n717_0;
	wire[1:0] w_n719_0;
	wire[1:0] w_n722_0;
	wire[1:0] w_n724_0;
	wire[1:0] w_n727_0;
	wire[1:0] w_n729_0;
	wire[1:0] w_n732_0;
	wire[1:0] w_n734_0;
	wire[1:0] w_n737_0;
	wire[1:0] w_n739_0;
	wire[1:0] w_n742_0;
	wire[1:0] w_n744_0;
	wire[1:0] w_n747_0;
	wire[1:0] w_n749_0;
	wire[1:0] w_n752_0;
	wire[1:0] w_n754_0;
	wire[1:0] w_n757_0;
	wire[1:0] w_n759_0;
	wire[1:0] w_n762_0;
	wire[1:0] w_n764_0;
	wire[1:0] w_n769_0;
	wire[1:0] w_n771_0;
	wire[1:0] w_n772_0;
	wire[1:0] w_n773_0;
	wire[1:0] w_n774_0;
	wire[1:0] w_n775_0;
	wire[1:0] w_n777_0;
	wire[1:0] w_n778_0;
	wire[1:0] w_n779_0;
	wire[1:0] w_n780_0;
	wire[1:0] w_n781_0;
	wire[1:0] w_n782_0;
	wire[1:0] w_n783_0;
	wire[1:0] w_n784_0;
	wire[1:0] w_n785_0;
	wire[1:0] w_n786_0;
	wire[1:0] w_n787_0;
	wire[1:0] w_n788_0;
	wire[1:0] w_n789_0;
	wire[1:0] w_n790_0;
	wire[1:0] w_n791_0;
	wire[1:0] w_n792_0;
	wire[1:0] w_n793_0;
	wire[1:0] w_n794_0;
	wire[1:0] w_n795_0;
	wire[1:0] w_n796_0;
	wire[1:0] w_n797_0;
	wire[1:0] w_n798_0;
	wire[1:0] w_n799_0;
	wire[1:0] w_n800_0;
	wire[1:0] w_n802_0;
	wire[1:0] w_n803_0;
	wire[1:0] w_n805_0;
	wire[1:0] w_n810_0;
	wire[1:0] w_n811_0;
	wire[1:0] w_n815_0;
	wire[1:0] w_n816_0;
	wire[2:0] w_n820_0;
	wire[1:0] w_n822_0;
	wire[1:0] w_n825_0;
	wire[1:0] w_n827_0;
	wire[1:0] w_n830_0;
	wire[1:0] w_n832_0;
	wire[1:0] w_n835_0;
	wire[1:0] w_n837_0;
	wire[1:0] w_n840_0;
	wire[1:0] w_n842_0;
	wire[1:0] w_n845_0;
	wire[1:0] w_n847_0;
	wire[1:0] w_n850_0;
	wire[1:0] w_n852_0;
	wire[1:0] w_n855_0;
	wire[1:0] w_n857_0;
	wire[1:0] w_n860_0;
	wire[1:0] w_n862_0;
	wire[1:0] w_n865_0;
	wire[1:0] w_n867_0;
	wire[1:0] w_n872_0;
	wire[1:0] w_n874_0;
	wire[1:0] w_n875_0;
	wire[1:0] w_n877_0;
	wire[1:0] w_n879_0;
	wire[1:0] w_n880_0;
	wire[1:0] w_n881_0;
	wire[1:0] w_n882_0;
	wire[1:0] w_n883_0;
	wire[1:0] w_n884_0;
	wire[1:0] w_n885_0;
	wire[1:0] w_n886_0;
	wire[1:0] w_n887_0;
	wire[1:0] w_n888_0;
	wire[1:0] w_n889_0;
	wire[1:0] w_n890_0;
	wire[1:0] w_n891_0;
	wire[1:0] w_n892_0;
	wire[1:0] w_n893_0;
	wire[1:0] w_n894_0;
	wire[1:0] w_n895_0;
	wire[1:0] w_n896_0;
	wire[1:0] w_n897_0;
	wire[1:0] w_n898_0;
	wire[1:0] w_n899_0;
	wire[2:0] w_n900_0;
	wire[1:0] w_n902_0;
	wire[1:0] w_n903_0;
	wire[1:0] w_n904_0;
	wire[1:0] w_n905_0;
	wire[1:0] w_n910_0;
	wire[1:0] w_n911_0;
	wire[2:0] w_n915_0;
	wire[1:0] w_n916_0;
	wire[1:0] w_n922_0;
	wire[1:0] w_n924_0;
	wire[1:0] w_n927_0;
	wire[1:0] w_n929_0;
	wire[1:0] w_n932_0;
	wire[1:0] w_n934_0;
	wire[1:0] w_n937_0;
	wire[1:0] w_n939_0;
	wire[1:0] w_n942_0;
	wire[1:0] w_n944_0;
	wire[1:0] w_n947_0;
	wire[1:0] w_n949_0;
	wire[1:0] w_n952_0;
	wire[1:0] w_n954_0;
	wire[1:0] w_n957_0;
	wire[1:0] w_n959_0;
	wire[1:0] w_n962_0;
	wire[1:0] w_n964_0;
	wire[1:0] w_n967_0;
	wire[1:0] w_n969_0;
	wire[1:0] w_n972_0;
	wire[1:0] w_n974_0;
	wire[1:0] w_n978_0;
	wire[1:0] w_n980_0;
	wire[1:0] w_n982_0;
	wire[1:0] w_n983_0;
	wire[1:0] w_n984_0;
	wire[1:0] w_n985_0;
	wire[1:0] w_n986_0;
	wire[1:0] w_n987_0;
	wire[1:0] w_n988_0;
	wire[1:0] w_n989_0;
	wire[1:0] w_n990_0;
	wire[1:0] w_n991_0;
	wire[1:0] w_n992_0;
	wire[1:0] w_n993_0;
	wire[1:0] w_n994_0;
	wire[1:0] w_n995_0;
	wire[1:0] w_n996_0;
	wire[1:0] w_n997_0;
	wire[1:0] w_n998_0;
	wire[1:0] w_n999_0;
	wire[1:0] w_n1000_0;
	wire[1:0] w_n1001_0;
	wire[1:0] w_n1002_0;
	wire[1:0] w_n1003_0;
	wire[1:0] w_n1004_0;
	wire[1:0] w_n1005_0;
	wire[1:0] w_n1006_0;
	wire[1:0] w_n1007_0;
	wire[1:0] w_n1008_0;
	wire[1:0] w_n1009_0;
	wire[1:0] w_n1011_0;
	wire[1:0] w_n1013_0;
	wire[1:0] w_n1017_0;
	wire[1:0] w_n1018_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1023_0;
	wire[1:0] w_n1026_0;
	wire[1:0] w_n1028_0;
	wire[1:0] w_n1031_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1036_0;
	wire[1:0] w_n1038_0;
	wire[1:0] w_n1041_0;
	wire[1:0] w_n1043_0;
	wire[1:0] w_n1046_0;
	wire[1:0] w_n1048_0;
	wire[1:0] w_n1051_0;
	wire[1:0] w_n1053_0;
	wire[1:0] w_n1056_0;
	wire[1:0] w_n1058_0;
	wire[1:0] w_n1061_0;
	wire[1:0] w_n1063_0;
	wire[1:0] w_n1066_0;
	wire[1:0] w_n1068_0;
	wire[1:0] w_n1071_0;
	wire[1:0] w_n1073_0;
	wire[1:0] w_n1076_0;
	wire[1:0] w_n1077_0;
	wire[1:0] w_n1078_0;
	wire[1:0] w_n1080_0;
	wire[1:0] w_n1082_0;
	wire[1:0] w_n1083_0;
	wire[1:0] w_n1084_0;
	wire[1:0] w_n1085_0;
	wire[1:0] w_n1086_0;
	wire[1:0] w_n1087_0;
	wire[1:0] w_n1088_0;
	wire[1:0] w_n1089_0;
	wire[1:0] w_n1090_0;
	wire[1:0] w_n1091_0;
	wire[1:0] w_n1092_0;
	wire[1:0] w_n1093_0;
	wire[1:0] w_n1094_0;
	wire[1:0] w_n1095_0;
	wire[1:0] w_n1096_0;
	wire[1:0] w_n1097_0;
	wire[1:0] w_n1098_0;
	wire[1:0] w_n1099_0;
	wire[1:0] w_n1100_0;
	wire[1:0] w_n1101_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1103_0;
	wire[1:0] w_n1105_0;
	wire[1:0] w_n1106_0;
	wire[1:0] w_n1107_0;
	wire[1:0] w_n1108_0;
	wire[1:0] w_n1109_0;
	wire[1:0] w_n1115_0;
	wire[1:0] w_n1119_0;
	wire[1:0] w_n1120_0;
	wire[1:0] w_n1124_0;
	wire[1:0] w_n1126_0;
	wire[1:0] w_n1129_0;
	wire[1:0] w_n1131_0;
	wire[1:0] w_n1134_0;
	wire[1:0] w_n1136_0;
	wire[1:0] w_n1139_0;
	wire[1:0] w_n1141_0;
	wire[1:0] w_n1144_0;
	wire[1:0] w_n1146_0;
	wire[1:0] w_n1149_0;
	wire[1:0] w_n1151_0;
	wire[1:0] w_n1154_0;
	wire[1:0] w_n1156_0;
	wire[1:0] w_n1159_0;
	wire[1:0] w_n1161_0;
	wire[1:0] w_n1164_0;
	wire[1:0] w_n1166_0;
	wire[1:0] w_n1169_0;
	wire[1:0] w_n1171_0;
	wire[1:0] w_n1174_0;
	wire[1:0] w_n1175_0;
	wire[1:0] w_n1176_0;
	wire[1:0] w_n1179_0;
	wire[1:0] w_n1181_0;
	wire[1:0] w_n1182_0;
	wire[1:0] w_n1183_0;
	wire[1:0] w_n1184_0;
	wire[1:0] w_n1185_0;
	wire[1:0] w_n1186_0;
	wire[1:0] w_n1187_0;
	wire[1:0] w_n1188_0;
	wire[1:0] w_n1189_0;
	wire[1:0] w_n1190_0;
	wire[1:0] w_n1191_0;
	wire[1:0] w_n1192_0;
	wire[1:0] w_n1193_0;
	wire[1:0] w_n1194_0;
	wire[1:0] w_n1195_0;
	wire[1:0] w_n1196_0;
	wire[1:0] w_n1197_0;
	wire[1:0] w_n1198_0;
	wire[1:0] w_n1199_0;
	wire[1:0] w_n1200_0;
	wire[1:0] w_n1201_0;
	wire[1:0] w_n1203_0;
	wire[1:0] w_n1205_0;
	wire[1:0] w_n1206_0;
	wire[1:0] w_n1207_0;
	wire[1:0] w_n1213_0;
	wire[1:0] w_n1216_0;
	wire[1:0] w_n1217_0;
	wire[1:0] w_n1220_0;
	wire[1:0] w_n1222_0;
	wire[1:0] w_n1225_0;
	wire[1:0] w_n1227_0;
	wire[1:0] w_n1230_0;
	wire[1:0] w_n1232_0;
	wire[1:0] w_n1235_0;
	wire[1:0] w_n1237_0;
	wire[1:0] w_n1240_0;
	wire[1:0] w_n1242_0;
	wire[1:0] w_n1245_0;
	wire[1:0] w_n1247_0;
	wire[1:0] w_n1250_0;
	wire[1:0] w_n1252_0;
	wire[1:0] w_n1255_0;
	wire[1:0] w_n1257_0;
	wire[1:0] w_n1260_0;
	wire[1:0] w_n1262_0;
	wire[1:0] w_n1265_0;
	wire[1:0] w_n1266_0;
	wire[1:0] w_n1267_0;
	wire[1:0] w_n1270_0;
	wire[1:0] w_n1272_0;
	wire[1:0] w_n1273_0;
	wire[1:0] w_n1274_0;
	wire[1:0] w_n1275_0;
	wire[1:0] w_n1276_0;
	wire[1:0] w_n1277_0;
	wire[1:0] w_n1278_0;
	wire[1:0] w_n1279_0;
	wire[1:0] w_n1280_0;
	wire[1:0] w_n1281_0;
	wire[1:0] w_n1282_0;
	wire[1:0] w_n1283_0;
	wire[1:0] w_n1284_0;
	wire[1:0] w_n1285_0;
	wire[1:0] w_n1286_0;
	wire[1:0] w_n1287_0;
	wire[1:0] w_n1288_0;
	wire[1:0] w_n1289_0;
	wire[1:0] w_n1290_0;
	wire[1:0] w_n1291_0;
	wire[1:0] w_n1293_0;
	wire[1:0] w_n1294_0;
	wire[1:0] w_n1295_0;
	wire[1:0] w_n1301_0;
	wire[1:0] w_n1306_0;
	wire[1:0] w_n1307_0;
	wire[1:0] w_n1310_0;
	wire[1:0] w_n1312_0;
	wire[1:0] w_n1315_0;
	wire[1:0] w_n1317_0;
	wire[1:0] w_n1320_0;
	wire[1:0] w_n1322_0;
	wire[1:0] w_n1325_0;
	wire[1:0] w_n1327_0;
	wire[1:0] w_n1330_0;
	wire[1:0] w_n1332_0;
	wire[1:0] w_n1335_0;
	wire[1:0] w_n1337_0;
	wire[1:0] w_n1340_0;
	wire[1:0] w_n1342_0;
	wire[1:0] w_n1345_0;
	wire[1:0] w_n1347_0;
	wire[1:0] w_n1350_0;
	wire[1:0] w_n1351_0;
	wire[1:0] w_n1352_0;
	wire[1:0] w_n1355_0;
	wire[1:0] w_n1357_0;
	wire[1:0] w_n1358_0;
	wire[1:0] w_n1359_0;
	wire[1:0] w_n1360_0;
	wire[1:0] w_n1361_0;
	wire[1:0] w_n1362_0;
	wire[1:0] w_n1363_0;
	wire[1:0] w_n1364_0;
	wire[1:0] w_n1365_0;
	wire[1:0] w_n1366_0;
	wire[1:0] w_n1367_0;
	wire[1:0] w_n1368_0;
	wire[1:0] w_n1369_0;
	wire[1:0] w_n1370_0;
	wire[1:0] w_n1371_0;
	wire[1:0] w_n1372_0;
	wire[1:0] w_n1373_0;
	wire[1:0] w_n1374_0;
	wire[1:0] w_n1376_0;
	wire[1:0] w_n1378_0;
	wire[1:0] w_n1379_0;
	wire[1:0] w_n1384_0;
	wire[1:0] w_n1389_0;
	wire[1:0] w_n1390_0;
	wire[1:0] w_n1393_0;
	wire[1:0] w_n1395_0;
	wire[1:0] w_n1398_0;
	wire[1:0] w_n1400_0;
	wire[1:0] w_n1403_0;
	wire[1:0] w_n1405_0;
	wire[1:0] w_n1408_0;
	wire[1:0] w_n1410_0;
	wire[1:0] w_n1413_0;
	wire[1:0] w_n1415_0;
	wire[1:0] w_n1418_0;
	wire[1:0] w_n1420_0;
	wire[1:0] w_n1423_0;
	wire[1:0] w_n1425_0;
	wire[1:0] w_n1428_0;
	wire[1:0] w_n1429_0;
	wire[1:0] w_n1430_0;
	wire[1:0] w_n1433_0;
	wire[1:0] w_n1435_0;
	wire[1:0] w_n1436_0;
	wire[1:0] w_n1437_0;
	wire[1:0] w_n1438_0;
	wire[1:0] w_n1439_0;
	wire[1:0] w_n1440_0;
	wire[1:0] w_n1441_0;
	wire[1:0] w_n1442_0;
	wire[1:0] w_n1443_0;
	wire[1:0] w_n1444_0;
	wire[1:0] w_n1445_0;
	wire[1:0] w_n1446_0;
	wire[1:0] w_n1447_0;
	wire[1:0] w_n1448_0;
	wire[1:0] w_n1449_0;
	wire[1:0] w_n1450_0;
	wire[1:0] w_n1452_0;
	wire[1:0] w_n1454_0;
	wire[1:0] w_n1455_0;
	wire[1:0] w_n1460_0;
	wire[1:0] w_n1465_0;
	wire[1:0] w_n1466_0;
	wire[1:0] w_n1469_0;
	wire[1:0] w_n1471_0;
	wire[1:0] w_n1474_0;
	wire[1:0] w_n1476_0;
	wire[1:0] w_n1479_0;
	wire[1:0] w_n1481_0;
	wire[1:0] w_n1484_0;
	wire[1:0] w_n1486_0;
	wire[1:0] w_n1489_0;
	wire[1:0] w_n1491_0;
	wire[1:0] w_n1494_0;
	wire[1:0] w_n1496_0;
	wire[1:0] w_n1499_0;
	wire[1:0] w_n1500_0;
	wire[1:0] w_n1501_0;
	wire[1:0] w_n1504_0;
	wire[1:0] w_n1506_0;
	wire[1:0] w_n1507_0;
	wire[1:0] w_n1508_0;
	wire[1:0] w_n1509_0;
	wire[1:0] w_n1510_0;
	wire[1:0] w_n1511_0;
	wire[1:0] w_n1512_0;
	wire[1:0] w_n1513_0;
	wire[1:0] w_n1514_0;
	wire[1:0] w_n1515_0;
	wire[1:0] w_n1516_0;
	wire[1:0] w_n1517_0;
	wire[1:0] w_n1518_0;
	wire[1:0] w_n1519_0;
	wire[1:0] w_n1521_0;
	wire[1:0] w_n1523_0;
	wire[1:0] w_n1524_0;
	wire[1:0] w_n1529_0;
	wire[1:0] w_n1534_0;
	wire[1:0] w_n1535_0;
	wire[1:0] w_n1538_0;
	wire[1:0] w_n1540_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1545_0;
	wire[1:0] w_n1548_0;
	wire[1:0] w_n1550_0;
	wire[1:0] w_n1553_0;
	wire[1:0] w_n1555_0;
	wire[1:0] w_n1558_0;
	wire[1:0] w_n1560_0;
	wire[1:0] w_n1563_0;
	wire[1:0] w_n1564_0;
	wire[1:0] w_n1565_0;
	wire[1:0] w_n1568_0;
	wire[1:0] w_n1570_0;
	wire[1:0] w_n1571_0;
	wire[1:0] w_n1572_0;
	wire[1:0] w_n1573_0;
	wire[1:0] w_n1574_0;
	wire[1:0] w_n1575_0;
	wire[1:0] w_n1576_0;
	wire[1:0] w_n1577_0;
	wire[1:0] w_n1578_0;
	wire[1:0] w_n1579_0;
	wire[1:0] w_n1580_0;
	wire[1:0] w_n1581_0;
	wire[1:0] w_n1583_0;
	wire[1:0] w_n1585_0;
	wire[1:0] w_n1586_0;
	wire[1:0] w_n1591_0;
	wire[1:0] w_n1596_0;
	wire[1:0] w_n1597_0;
	wire[1:0] w_n1600_0;
	wire[1:0] w_n1602_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1607_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1612_0;
	wire[1:0] w_n1615_0;
	wire[1:0] w_n1617_0;
	wire[1:0] w_n1620_0;
	wire[1:0] w_n1621_0;
	wire[1:0] w_n1622_0;
	wire[1:0] w_n1625_0;
	wire[1:0] w_n1627_0;
	wire[1:0] w_n1628_0;
	wire[1:0] w_n1629_0;
	wire[1:0] w_n1630_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1632_0;
	wire[1:0] w_n1633_0;
	wire[1:0] w_n1634_0;
	wire[1:0] w_n1635_0;
	wire[1:0] w_n1636_0;
	wire[1:0] w_n1638_0;
	wire[1:0] w_n1640_0;
	wire[1:0] w_n1641_0;
	wire[1:0] w_n1646_0;
	wire[1:0] w_n1651_0;
	wire[1:0] w_n1653_0;
	wire[1:0] w_n1656_0;
	wire[1:0] w_n1658_0;
	wire[1:0] w_n1661_0;
	wire[1:0] w_n1663_0;
	wire[1:0] w_n1666_0;
	wire[1:0] w_n1668_0;
	wire[1:0] w_n1671_0;
	wire[1:0] w_n1672_0;
	wire[1:0] w_n1673_0;
	wire[1:0] w_n1676_0;
	wire[1:0] w_n1678_0;
	wire[1:0] w_n1679_0;
	wire[1:0] w_n1680_0;
	wire[1:0] w_n1681_0;
	wire[1:0] w_n1682_0;
	wire[1:0] w_n1683_0;
	wire[1:0] w_n1684_0;
	wire[1:0] w_n1685_0;
	wire[1:0] w_n1686_0;
	wire[1:0] w_n1688_0;
	wire[1:0] w_n1689_0;
	wire[1:0] w_n1694_0;
	wire[1:0] w_n1697_0;
	wire[1:0] w_n1699_0;
	wire[1:0] w_n1702_0;
	wire[1:0] w_n1704_0;
	wire[1:0] w_n1707_0;
	wire[1:0] w_n1709_0;
	wire[1:0] w_n1712_0;
	wire[1:0] w_n1713_0;
	wire[1:0] w_n1714_0;
	wire[1:0] w_n1717_0;
	wire[1:0] w_n1719_0;
	wire[1:0] w_n1720_0;
	wire[1:0] w_n1721_0;
	wire[1:0] w_n1722_0;
	wire[1:0] w_n1723_0;
	wire[1:0] w_n1724_0;
	wire[1:0] w_n1725_0;
	wire[1:0] w_n1726_0;
	wire[1:0] w_n1727_0;
	wire[1:0] w_n1734_0;
	wire[1:0] w_n1737_0;
	wire[1:0] w_n1739_0;
	wire[1:0] w_n1742_0;
	wire[1:0] w_n1744_0;
	wire[1:0] w_n1747_0;
	wire[1:0] w_n1748_0;
	wire[1:0] w_n1749_0;
	wire[1:0] w_n1752_0;
	wire[1:0] w_n1754_0;
	wire[1:0] w_n1755_0;
	wire[1:0] w_n1756_0;
	wire[1:0] w_n1757_0;
	wire[1:0] w_n1758_0;
	wire[1:0] w_n1759_0;
	wire[1:0] w_n1760_0;
	wire[1:0] w_n1767_0;
	wire[1:0] w_n1770_0;
	wire[1:0] w_n1772_0;
	wire[1:0] w_n1775_0;
	wire[1:0] w_n1776_0;
	wire[1:0] w_n1777_0;
	wire[1:0] w_n1780_0;
	wire[1:0] w_n1782_0;
	wire[1:0] w_n1783_0;
	wire[1:0] w_n1784_0;
	wire[1:0] w_n1785_0;
	wire[1:0] w_n1786_0;
	wire[1:0] w_n1793_0;
	wire[1:0] w_n1796_0;
	wire[1:0] w_n1797_0;
	wire[1:0] w_n1798_0;
	wire[1:0] w_n1801_0;
	wire[1:0] w_n1803_0;
	wire[1:0] w_n1804_0;
	wire[1:0] w_n1805_0;
	wire[1:0] w_n1807_0;
	wire[1:0] w_n1810_0;
	wire[1:0] w_n1817_0;
	wire[1:0] w_n1818_0;
	wire w_dff_B_vzvAZJxt5_0;
	wire w_dff_B_SUExNrn46_0;
	wire w_dff_B_QdpwnOgJ1_1;
	wire w_dff_B_gafEQwL95_1;
	wire w_dff_B_89v3w0f13_1;
	wire w_dff_B_InF7qtmv0_1;
	wire w_dff_B_1cqxJKRO6_1;
	wire w_dff_B_cP4vnAxd8_1;
	wire w_dff_B_Jcr8KLbV6_1;
	wire w_dff_B_6g4JKUI96_1;
	wire w_dff_B_yVHZgx371_1;
	wire w_dff_B_r6Cme3p80_1;
	wire w_dff_B_Ou6HbKVR3_1;
	wire w_dff_B_BqKy0Luv7_1;
	wire w_dff_B_mhYvGvOc6_1;
	wire w_dff_B_RZC5JMcr9_1;
	wire w_dff_B_bhnAR0OI2_1;
	wire w_dff_B_3prdParx6_1;
	wire w_dff_B_7lGMKzH84_1;
	wire w_dff_B_UWWTPYVO4_1;
	wire w_dff_B_Jj1iQ7xH1_1;
	wire w_dff_B_eEbaSphm0_1;
	wire w_dff_B_ClFCjDTN8_1;
	wire w_dff_B_7JIWZQuW2_1;
	wire w_dff_B_nT9vTHWR8_1;
	wire w_dff_B_4BbOqokv2_1;
	wire w_dff_B_Bpxv5lyf9_1;
	wire w_dff_B_8PSTu8Y33_1;
	wire w_dff_B_N4uXRTGa1_1;
	wire w_dff_B_fZ2jmcSn8_1;
	wire w_dff_B_yfPk977F3_1;
	wire w_dff_B_BnXbdPhm6_1;
	wire w_dff_B_V9VTPdn51_1;
	wire w_dff_B_X1hFynFU2_1;
	wire w_dff_B_teMGEn4P1_1;
	wire w_dff_B_jPKZdBkI7_1;
	wire w_dff_B_cmuusSQw1_1;
	wire w_dff_B_AoEMteKx4_1;
	wire w_dff_B_Ey3muK8q4_1;
	wire w_dff_B_yGHGyHBk9_1;
	wire w_dff_B_jKFyHFyH7_1;
	wire w_dff_B_IxjpZylU9_1;
	wire w_dff_B_cAlEFDav4_1;
	wire w_dff_B_awJm5IGm1_1;
	wire w_dff_B_ZpPlB2Wm0_1;
	wire w_dff_B_H6n3cIIX0_1;
	wire w_dff_B_DpFfkr0Y4_1;
	wire w_dff_B_m2ENnNou3_1;
	wire w_dff_B_6o123e5Y7_1;
	wire w_dff_B_VqpbOfil5_1;
	wire w_dff_B_7jW0raWj5_1;
	wire w_dff_B_tUSHvTyN0_1;
	wire w_dff_B_r7osvCbN1_1;
	wire w_dff_B_yrE90Xy56_1;
	wire w_dff_B_cIap07mj7_1;
	wire w_dff_B_3j8TDRSL8_1;
	wire w_dff_B_6s4IeKIh3_1;
	wire w_dff_B_hYLLQ15x6_1;
	wire w_dff_B_BAd2M8LT6_1;
	wire w_dff_B_DSoG4S084_1;
	wire w_dff_B_355LobdI0_1;
	wire w_dff_B_fukn4ltA0_1;
	wire w_dff_B_qgJReu1N7_1;
	wire w_dff_B_3N1B4Rtq0_1;
	wire w_dff_B_vJqVPxU03_1;
	wire w_dff_B_CwSRRwjN5_1;
	wire w_dff_B_GedtU0vi4_1;
	wire w_dff_B_oovehKht1_1;
	wire w_dff_B_iN5qnS8z5_1;
	wire w_dff_B_DL886yBF3_1;
	wire w_dff_B_SVAJzocY6_1;
	wire w_dff_B_urygT3bm1_1;
	wire w_dff_B_jORn2jGt1_1;
	wire w_dff_B_bZkIttkF1_1;
	wire w_dff_B_RfEAPgye7_1;
	wire w_dff_B_54bn7vVA8_1;
	wire w_dff_B_3v6pA5oI5_1;
	wire w_dff_B_v2VG6z1c8_1;
	wire w_dff_B_qxzwDn6E8_1;
	wire w_dff_B_XwVx16Ix4_1;
	wire w_dff_B_QyljmIj94_1;
	wire w_dff_B_1mmN5BzQ6_1;
	wire w_dff_B_3XoXNWDN7_1;
	wire w_dff_B_Q9fGXPqs0_1;
	wire w_dff_B_Wg3iCdZg8_1;
	wire w_dff_B_r3WimfWD0_1;
	wire w_dff_B_zFvfwIzp7_1;
	wire w_dff_B_qy1kQbUX1_1;
	wire w_dff_B_x69OOTQN3_1;
	wire w_dff_B_rCCDKrWU9_1;
	wire w_dff_B_Vxl0881H9_1;
	wire w_dff_B_3PWAp9Kk9_1;
	wire w_dff_B_7ClctyZ17_1;
	wire w_dff_B_tRLlBSwL4_1;
	wire w_dff_B_E8fVHq9U7_1;
	wire w_dff_B_rATvijCS6_1;
	wire w_dff_B_QHLHFRca2_1;
	wire w_dff_B_mSfyylXG9_1;
	wire w_dff_B_MBBrBup01_1;
	wire w_dff_B_B2o5QZKN3_1;
	wire w_dff_B_3411S7Qh3_1;
	wire w_dff_B_3D87MeEd7_1;
	wire w_dff_B_5BltfdqI3_1;
	wire w_dff_B_0rXH0pJp2_1;
	wire w_dff_B_GD49Hmfq1_1;
	wire w_dff_B_wSXpna8E5_1;
	wire w_dff_B_9xZoLqYk6_1;
	wire w_dff_B_NZoRyegg1_1;
	wire w_dff_B_c3me6WE41_1;
	wire w_dff_B_d7eeEngJ3_1;
	wire w_dff_B_kdsmAVtO7_1;
	wire w_dff_B_k1sgEzGa7_1;
	wire w_dff_B_j2EHEmno9_1;
	wire w_dff_B_bKpyVoNp3_1;
	wire w_dff_B_OecDV8788_1;
	wire w_dff_B_Y35OwnYU3_1;
	wire w_dff_B_JFNjBZFt9_1;
	wire w_dff_B_TL2bxGWf0_1;
	wire w_dff_B_axgoBAK62_1;
	wire w_dff_B_7FPtVNEg4_1;
	wire w_dff_B_ugwhrDwY8_1;
	wire w_dff_B_fLm8AuIN0_1;
	wire w_dff_B_GAM8RXKv7_1;
	wire w_dff_B_CUAIUGvI3_1;
	wire w_dff_B_hRB2htQv6_1;
	wire w_dff_B_om1Gq63v3_1;
	wire w_dff_B_cBM9Hzd33_1;
	wire w_dff_B_yPHyzvWq7_1;
	wire w_dff_B_1cTmXVId4_1;
	wire w_dff_B_6ID0EMhh4_1;
	wire w_dff_B_VSwwZBpj9_1;
	wire w_dff_B_UH1jfDFs6_1;
	wire w_dff_B_vAZaof7z0_1;
	wire w_dff_B_tRp9EaF18_1;
	wire w_dff_B_Ydftyv7r1_1;
	wire w_dff_B_nFLHIZA47_1;
	wire w_dff_B_ZlVotAqf9_1;
	wire w_dff_B_7lUb0BKv2_1;
	wire w_dff_B_QxQUFhzn0_1;
	wire w_dff_B_NJRF68sV5_1;
	wire w_dff_B_9SwlEMC75_1;
	wire w_dff_B_uaoz8z8P3_1;
	wire w_dff_B_fa9QVryM6_1;
	wire w_dff_B_YjoGX06V4_1;
	wire w_dff_B_spc827hJ4_1;
	wire w_dff_B_AfFkH6io8_1;
	wire w_dff_B_lROTlTqo4_1;
	wire w_dff_B_xu5w64Ol1_1;
	wire w_dff_B_e7S8QqC39_1;
	wire w_dff_B_UpOR4GE39_1;
	wire w_dff_B_5PwDEXba4_1;
	wire w_dff_B_0PhRkLP33_1;
	wire w_dff_B_l5aAVy7v5_1;
	wire w_dff_B_dpS8tZeW6_1;
	wire w_dff_B_aaOeSY6X0_1;
	wire w_dff_B_WL87fzhT6_1;
	wire w_dff_B_CDxtdfPQ8_1;
	wire w_dff_B_uJkSSJsU0_1;
	wire w_dff_B_K6dn33Fl4_1;
	wire w_dff_B_ZmREDV1C2_1;
	wire w_dff_B_wJpNu3ru1_1;
	wire w_dff_B_U6FlIi3u0_1;
	wire w_dff_B_OZaNzmmr6_1;
	wire w_dff_B_WvXoQYu74_1;
	wire w_dff_B_qsB6VOwN6_1;
	wire w_dff_B_yA7PwUM54_1;
	wire w_dff_B_YFRm4K5W1_1;
	wire w_dff_B_xBSuuJ7s4_1;
	wire w_dff_B_k5vWgTKx4_1;
	wire w_dff_B_y8g3ES8h6_1;
	wire w_dff_B_Tbgn4Dom7_1;
	wire w_dff_B_BHAnsAri8_1;
	wire w_dff_B_ldS3q1HM3_1;
	wire w_dff_B_we568uMK7_1;
	wire w_dff_B_5lwAKedS5_1;
	wire w_dff_B_10IAnLPV1_1;
	wire w_dff_B_QDjuZ69o9_1;
	wire w_dff_B_l3aIp33a0_1;
	wire w_dff_B_iNzi5dWU6_1;
	wire w_dff_B_E1qSF1qR7_1;
	wire w_dff_B_69kVTkT75_1;
	wire w_dff_B_aSayIanv6_1;
	wire w_dff_B_FyHTsubF8_1;
	wire w_dff_B_CLzBWEe19_1;
	wire w_dff_B_Ocbb6EEg2_1;
	wire w_dff_B_ryUpwBpC7_1;
	wire w_dff_B_9coZKIBA6_1;
	wire w_dff_B_ndGhYzjJ7_1;
	wire w_dff_B_sMzjXJOr7_1;
	wire w_dff_B_DGKZt9aO1_1;
	wire w_dff_B_bt0qO9ob1_1;
	wire w_dff_B_GvYmugE58_1;
	wire w_dff_B_Q3NRNJLN1_1;
	wire w_dff_B_DgvSxp4c5_1;
	wire w_dff_B_sX0C7uwN8_1;
	wire w_dff_B_KKdBTCpF4_1;
	wire w_dff_B_TZMF1tqX9_1;
	wire w_dff_B_J01r9X969_1;
	wire w_dff_B_B979yd3B0_1;
	wire w_dff_B_Hf4zsWZq2_1;
	wire w_dff_B_vqAjp3PQ7_1;
	wire w_dff_B_HRfTJ6D17_1;
	wire w_dff_B_0Xqp5hgY9_1;
	wire w_dff_B_kPTDKQsO5_1;
	wire w_dff_B_DQxuNFZS7_1;
	wire w_dff_B_Sg8ryoas8_1;
	wire w_dff_B_L378aHdO7_1;
	wire w_dff_B_6qm95FkR7_1;
	wire w_dff_B_m3tUgcO24_1;
	wire w_dff_B_ni4qlqbW4_1;
	wire w_dff_B_TWs3YKRW4_1;
	wire w_dff_B_QaDjQRqQ7_1;
	wire w_dff_B_tli5ftp98_1;
	wire w_dff_B_unw30J9S4_1;
	wire w_dff_B_m9JW1eFQ9_1;
	wire w_dff_B_rWDfYdle0_1;
	wire w_dff_B_wTGAELPA5_1;
	wire w_dff_B_4Qjncd7v3_1;
	wire w_dff_B_DLZ0O1FA3_1;
	wire w_dff_B_6wef0Zqj3_1;
	wire w_dff_B_ZwYgijw02_1;
	wire w_dff_B_yWI8v3Fj9_1;
	wire w_dff_B_XUlsDNFh9_1;
	wire w_dff_B_11YpHJLM3_1;
	wire w_dff_B_gJrbHuAA6_1;
	wire w_dff_B_1vaIfmbv3_1;
	wire w_dff_B_EccYk7iG1_1;
	wire w_dff_B_gVe4cBXl2_1;
	wire w_dff_B_4YUH2rzp4_1;
	wire w_dff_B_rjAx0b5z0_1;
	wire w_dff_B_j5znD4rJ2_1;
	wire w_dff_B_xbmNtxnL2_1;
	wire w_dff_B_gdt0f4fK9_1;
	wire w_dff_B_0EksrcoX7_1;
	wire w_dff_B_P8QCH00j3_1;
	wire w_dff_B_OLxsTluA8_1;
	wire w_dff_B_zPxi1Q6c6_1;
	wire w_dff_B_1R5NIVMX4_1;
	wire w_dff_B_CBGfoSOi5_1;
	wire w_dff_B_MSn1eXOV3_1;
	wire w_dff_B_w2aUY5463_1;
	wire w_dff_B_yKWRbLQF0_1;
	wire w_dff_B_lMS2eIjt1_1;
	wire w_dff_B_DywTu1qP2_1;
	wire w_dff_B_XXN3uC1g4_1;
	wire w_dff_B_TLdhMHVW7_1;
	wire w_dff_B_Rg8nneRf0_1;
	wire w_dff_B_nOjWZ9wV7_1;
	wire w_dff_B_dpM7eu7c6_1;
	wire w_dff_B_Rt0HQJTD1_1;
	wire w_dff_B_hBBOq6Yx8_1;
	wire w_dff_B_jtsEMNWB4_1;
	wire w_dff_B_HiLQJmiD4_1;
	wire w_dff_B_Z3o7y1ZP7_1;
	wire w_dff_B_awLXZavE6_1;
	wire w_dff_B_g7tV1r0n6_1;
	wire w_dff_B_78v9h3AL5_1;
	wire w_dff_B_cuAE0DiZ0_1;
	wire w_dff_B_VURBNHcq7_1;
	wire w_dff_B_Kbu1jCJ97_1;
	wire w_dff_B_VXsNt6IB4_1;
	wire w_dff_B_KmcaORtk9_1;
	wire w_dff_B_VoATBfvH2_1;
	wire w_dff_B_fc5rMa0k5_1;
	wire w_dff_B_ifhE0vC63_1;
	wire w_dff_B_H46xCC9P7_1;
	wire w_dff_B_07yO4O7s1_1;
	wire w_dff_B_Iplt7siZ5_1;
	wire w_dff_B_7XKU0PZ66_1;
	wire w_dff_B_50E9cy6U7_1;
	wire w_dff_B_oPcfGX5r3_1;
	wire w_dff_B_6Y6UIDei8_1;
	wire w_dff_B_fT11e3pk3_1;
	wire w_dff_B_7Isxlngi2_1;
	wire w_dff_B_aIJIHk8U5_1;
	wire w_dff_B_eUIL5prO2_1;
	wire w_dff_B_zsdwqWWC6_1;
	wire w_dff_B_AC70GyfJ3_1;
	wire w_dff_B_EQgIEvn86_1;
	wire w_dff_B_1pt4iQjB0_1;
	wire w_dff_B_5twYTAM69_1;
	wire w_dff_B_XvMQT9Em7_1;
	wire w_dff_B_oXsLUE7i9_1;
	wire w_dff_B_5Aqb1Bcf7_1;
	wire w_dff_B_3YEZUXHr3_1;
	wire w_dff_B_dN4Gl2Bi3_1;
	wire w_dff_B_v4on7eZH4_1;
	wire w_dff_B_lvLwZhrU5_1;
	wire w_dff_B_z2ltMgUF8_1;
	wire w_dff_B_eaYUr7tn3_1;
	wire w_dff_B_wjJ96IPJ7_1;
	wire w_dff_B_PHAmY9oJ3_1;
	wire w_dff_B_FFOYMaYX7_1;
	wire w_dff_B_OSzyPwEm5_1;
	wire w_dff_B_vLcq54tm9_1;
	wire w_dff_B_uNChc3vM8_1;
	wire w_dff_B_Yn94UJfX5_1;
	wire w_dff_B_GfkLe7Pa2_1;
	wire w_dff_B_q6t8fYaQ5_1;
	wire w_dff_B_DcliMkSo5_1;
	wire w_dff_B_Sz4aXa4Y8_1;
	wire w_dff_B_ygdhXT930_1;
	wire w_dff_B_FWnZsOR52_1;
	wire w_dff_B_lNEgrRaH7_1;
	wire w_dff_B_QbtBYitR4_1;
	wire w_dff_B_iwwBkjQF1_1;
	wire w_dff_B_VZFVd6Eo0_1;
	wire w_dff_B_A9yPP5Ju7_1;
	wire w_dff_B_4xBDN4SN7_1;
	wire w_dff_B_wGcbOP2r4_1;
	wire w_dff_B_UibN8WY33_1;
	wire w_dff_B_WhludnsO2_1;
	wire w_dff_B_kXwV66Zz5_1;
	wire w_dff_B_nWxQvpep3_1;
	wire w_dff_B_5xaIIYPo2_1;
	wire w_dff_B_HN3mt3dj6_1;
	wire w_dff_B_8uvPJXgT8_1;
	wire w_dff_B_4SLee9TS5_0;
	wire w_dff_B_fUcCcxHo9_1;
	wire w_dff_B_Bhe9K82J7_1;
	wire w_dff_B_dKSVDGQp3_1;
	wire w_dff_B_yANjRof44_1;
	wire w_dff_B_Q8RpNch32_1;
	wire w_dff_B_I7XTI24x6_1;
	wire w_dff_B_Q6uIvwn59_1;
	wire w_dff_B_LVUkFt7i7_1;
	wire w_dff_B_BS0EEH3O9_1;
	wire w_dff_B_YnSBBg2P9_1;
	wire w_dff_B_gUyNrNT92_1;
	wire w_dff_B_D2xwiLSQ8_1;
	wire w_dff_B_tpT1tXET2_1;
	wire w_dff_B_eSzynpin2_1;
	wire w_dff_B_DRCwA28l1_1;
	wire w_dff_B_mhfjPYd78_0;
	wire w_dff_B_EKGU0wum5_0;
	wire w_dff_B_HeNgJGVL0_0;
	wire w_dff_B_UfuBytbQ2_0;
	wire w_dff_B_KnsOjQ7V5_0;
	wire w_dff_B_niyCTkNf7_0;
	wire w_dff_B_2MIJS98l9_0;
	wire w_dff_B_odXVTPrx9_0;
	wire w_dff_B_SKacsID54_0;
	wire w_dff_B_2kJjINXo9_0;
	wire w_dff_B_2zAr0Qx19_0;
	wire w_dff_B_f7C5wsGT2_0;
	wire w_dff_B_JaAxITgE4_0;
	wire w_dff_A_rT3HLtX14_0;
	wire w_dff_A_47l8Pkz52_0;
	wire w_dff_A_V2w1ap1I2_0;
	wire w_dff_A_5Z5zWbGP6_0;
	wire w_dff_A_XSpZLn2a6_0;
	wire w_dff_A_VjqPeLEa6_0;
	wire w_dff_A_dzr5DIwN6_0;
	wire w_dff_A_WcFhi0pj7_0;
	wire w_dff_A_MC3QqYvh8_0;
	wire w_dff_A_ThkRr3Hp4_0;
	wire w_dff_A_r6U5jSWR8_0;
	wire w_dff_A_QHohHitX3_0;
	wire w_dff_A_eFMJw3St7_0;
	wire w_dff_A_MML1jZwp4_0;
	wire w_dff_B_6Ux8M5LD0_1;
	wire w_dff_B_iEasrwnB9_1;
	wire w_dff_B_uFHBApah4_2;
	wire w_dff_B_zCckU8lI1_2;
	wire w_dff_B_4z105Ir07_2;
	wire w_dff_B_Usdx7tpg4_2;
	wire w_dff_B_WGatuEiZ4_2;
	wire w_dff_B_BKypBA0d3_2;
	wire w_dff_B_BelfP1WG7_2;
	wire w_dff_B_AoPnHSzj8_2;
	wire w_dff_B_PzrcveSQ6_2;
	wire w_dff_B_zM4gup2S2_2;
	wire w_dff_B_HkVPkxYu2_2;
	wire w_dff_B_NrT46Yvb7_2;
	wire w_dff_B_wUhfrYwx9_2;
	wire w_dff_B_tR94esYr2_2;
	wire w_dff_B_2RxmWKIM2_2;
	wire w_dff_B_nlj7rfPb3_2;
	wire w_dff_B_9UJyqb441_2;
	wire w_dff_B_Olh2PG0B5_2;
	wire w_dff_B_D9t3yHs04_2;
	wire w_dff_B_o4tY4MSg9_2;
	wire w_dff_B_Q6QhPzwv5_2;
	wire w_dff_B_CWMSSikA9_2;
	wire w_dff_B_Rvw2hzp05_2;
	wire w_dff_B_xsjw2vsm1_2;
	wire w_dff_B_1ww1o8PK8_2;
	wire w_dff_B_FGEbX3AC1_2;
	wire w_dff_B_pycMZsDz7_2;
	wire w_dff_B_64JZRsGy3_2;
	wire w_dff_B_cwNudo3v4_2;
	wire w_dff_B_PH20KCtK0_2;
	wire w_dff_B_qOJ7SaTp7_2;
	wire w_dff_B_nl4spyBO7_2;
	wire w_dff_B_CZvtNbY69_2;
	wire w_dff_B_6mIumRbI5_2;
	wire w_dff_B_NogpHkaB5_2;
	wire w_dff_B_EFfczy0S8_2;
	wire w_dff_B_4WCADZEa8_2;
	wire w_dff_B_uNtaOoeT3_2;
	wire w_dff_B_OGu9jeuz7_2;
	wire w_dff_B_kM0ArLr20_2;
	wire w_dff_B_OtppCZaK9_2;
	wire w_dff_B_ruoBLLGk4_2;
	wire w_dff_B_Dhiqr7bm1_2;
	wire w_dff_B_5ZeXVluX2_2;
	wire w_dff_B_x0q1LzIb6_2;
	wire w_dff_B_qwAzB6TL7_2;
	wire w_dff_B_ZH0Ny7Zg1_2;
	wire w_dff_B_pH7VgZtv2_2;
	wire w_dff_B_r4thXlzw5_2;
	wire w_dff_B_urnONHy72_2;
	wire w_dff_B_nqeiPldB3_2;
	wire w_dff_B_wMGJ46wb7_2;
	wire w_dff_B_9ldd8rqJ0_2;
	wire w_dff_B_zTSUg7Xy3_2;
	wire w_dff_B_4885EH6h0_2;
	wire w_dff_B_6pA5vqom0_2;
	wire w_dff_B_lqpZejf25_2;
	wire w_dff_B_wlAl6BB07_1;
	wire w_dff_B_YOnoyAXq1_1;
	wire w_dff_B_MQVTQO0r6_1;
	wire w_dff_B_hMxpTDQX0_1;
	wire w_dff_B_oNFhpEqu3_1;
	wire w_dff_B_8BhzC5nv3_1;
	wire w_dff_B_D15VyJj03_1;
	wire w_dff_B_PQNzjg0H5_1;
	wire w_dff_B_oQ1WeUbe0_1;
	wire w_dff_B_hnCaVgjP7_1;
	wire w_dff_B_nK2CbcYs4_1;
	wire w_dff_B_vdbemxIZ8_1;
	wire w_dff_B_c6XrcEjR7_1;
	wire w_dff_B_GobpxdEP5_0;
	wire w_dff_B_xfahLXTG1_0;
	wire w_dff_B_mo2Mm79I4_0;
	wire w_dff_B_clHexbmH9_0;
	wire w_dff_B_7ChBB2AN8_0;
	wire w_dff_B_KABMMdis3_0;
	wire w_dff_B_04JWzxSZ9_0;
	wire w_dff_B_4wWzOLQK1_0;
	wire w_dff_B_BrDt18yw5_0;
	wire w_dff_B_4k14NuXX3_0;
	wire w_dff_B_MEBU3MHh5_0;
	wire w_dff_B_Zgspq9E55_0;
	wire w_dff_A_crPSyuO82_1;
	wire w_dff_A_WKuPtrmB4_1;
	wire w_dff_A_Zuk5bBdR2_1;
	wire w_dff_A_XmdMQl875_1;
	wire w_dff_A_fTGx2qLi0_1;
	wire w_dff_A_utYalneR2_1;
	wire w_dff_A_O3Ww4BRY8_1;
	wire w_dff_A_mKvn4gex2_1;
	wire w_dff_A_dLNERbTQ0_1;
	wire w_dff_A_f6YOuO1D5_1;
	wire w_dff_A_egaLtwEk4_1;
	wire w_dff_A_LUEqeTel1_1;
	wire w_dff_A_EijMotbY9_1;
	wire w_dff_B_JZFTKxDn2_1;
	wire w_dff_B_Q0BzWonC9_1;
	wire w_dff_B_pUELCfFY0_1;
	wire w_dff_B_qPzFQeqf9_1;
	wire w_dff_B_i7PfZVBg9_1;
	wire w_dff_B_OIjBg37i3_1;
	wire w_dff_B_qPt7sSKQ0_1;
	wire w_dff_B_7t4VlZ8f3_1;
	wire w_dff_B_5hOmHfHY5_1;
	wire w_dff_B_UzRMDacO5_1;
	wire w_dff_B_1h0hJmOv9_1;
	wire w_dff_B_40IKokeU0_1;
	wire w_dff_B_IpFzrpKs7_1;
	wire w_dff_B_IRhPFDK15_0;
	wire w_dff_B_DZZ7xxOB1_0;
	wire w_dff_B_Ms9m2RZg5_0;
	wire w_dff_B_Tf8hITD79_0;
	wire w_dff_B_VBqWJIOP3_0;
	wire w_dff_B_Q9Ep1u1e0_0;
	wire w_dff_B_RdanKSAU4_0;
	wire w_dff_B_zRxMcXDf4_0;
	wire w_dff_B_DZvr5bWe2_0;
	wire w_dff_B_8UlkmnOB0_0;
	wire w_dff_B_QyIv5YhC3_0;
	wire w_dff_B_Eax2j83u3_0;
	wire w_dff_A_T9KFEdex7_1;
	wire w_dff_A_thZzegve2_1;
	wire w_dff_A_NmoBlnr84_1;
	wire w_dff_A_YyDrITFP6_1;
	wire w_dff_A_u4u4lKZC1_1;
	wire w_dff_A_1khubOvS9_1;
	wire w_dff_A_cntyXHu83_1;
	wire w_dff_A_9fO0aOLe4_1;
	wire w_dff_A_00BVOmPM9_1;
	wire w_dff_A_PwVDHGN71_1;
	wire w_dff_A_Fge183R41_1;
	wire w_dff_A_KFt5GgIB4_1;
	wire w_dff_A_4KVlAlWx1_1;
	wire w_dff_B_7cx5V5OS2_1;
	wire w_dff_B_ReRrmSwX3_1;
	wire w_dff_B_NfX4C5BL4_1;
	wire w_dff_B_5r5z626r1_1;
	wire w_dff_B_COetow5J0_1;
	wire w_dff_B_pFK8Rx8K0_1;
	wire w_dff_B_8rAwLMxX9_1;
	wire w_dff_B_PrtGY1vA8_1;
	wire w_dff_B_l4sWRafE4_1;
	wire w_dff_B_W4LavJEj3_1;
	wire w_dff_B_nQ5eUGWD8_1;
	wire w_dff_B_Kp36zHGa5_1;
	wire w_dff_B_vZrwHUxD9_1;
	wire w_dff_B_jzMeZDf95_0;
	wire w_dff_B_5DhVa4wc8_0;
	wire w_dff_B_fVEdAqmM8_0;
	wire w_dff_B_5T5gmPkk3_0;
	wire w_dff_B_PZ3rIPaP9_0;
	wire w_dff_B_w6hWCenc1_0;
	wire w_dff_B_7Mf5edzX4_0;
	wire w_dff_B_RZvoK1t43_0;
	wire w_dff_B_b303HJ6h9_0;
	wire w_dff_B_G5rdZPoX8_0;
	wire w_dff_B_s6zas3fz4_0;
	wire w_dff_B_S9IxMMvX1_0;
	wire w_dff_A_Ug5KqzIZ5_1;
	wire w_dff_A_qO2T8b5F1_1;
	wire w_dff_A_TXgtV5ST9_1;
	wire w_dff_A_uKmyPLmp7_1;
	wire w_dff_A_KeylDWXq9_1;
	wire w_dff_A_KG7eG7Oz2_1;
	wire w_dff_A_U5LspV7W1_1;
	wire w_dff_A_kd3jYeLR4_1;
	wire w_dff_A_SwWRfXa71_1;
	wire w_dff_A_W4ClE6JB0_1;
	wire w_dff_A_qcyHLUih9_1;
	wire w_dff_A_W973r2Lm0_1;
	wire w_dff_A_2vTb8S2q8_1;
	wire w_dff_B_SLTue1W65_1;
	wire w_dff_B_wG7sHNVc7_1;
	wire w_dff_B_ba6ckuz21_1;
	wire w_dff_B_erD4iTHp1_1;
	wire w_dff_B_FvnSXbol5_1;
	wire w_dff_B_2IHLg49y6_1;
	wire w_dff_B_uyEcYBeg8_1;
	wire w_dff_B_rNQUTJS04_1;
	wire w_dff_B_1QXjkdFr7_1;
	wire w_dff_B_rQLgk7kU5_1;
	wire w_dff_B_PqH95pFh5_1;
	wire w_dff_B_QA0up3dU1_1;
	wire w_dff_B_GZ6FuMXH6_1;
	wire w_dff_B_Cb6IpgKB9_0;
	wire w_dff_B_ZdELOMLu5_0;
	wire w_dff_B_PF9u3AFH8_0;
	wire w_dff_B_S76kN2ap0_0;
	wire w_dff_B_ruAuqKJX9_0;
	wire w_dff_B_BLKp01f08_0;
	wire w_dff_B_PMavN43V1_0;
	wire w_dff_B_s64Hssp82_0;
	wire w_dff_B_pnyncAxt8_0;
	wire w_dff_B_zTtpbYN36_0;
	wire w_dff_B_XRCDyfgr8_0;
	wire w_dff_B_OqdGXR4B1_0;
	wire w_dff_A_JCm8jvZF4_1;
	wire w_dff_A_AhLKwjoj4_1;
	wire w_dff_A_lJae0g2f1_1;
	wire w_dff_A_vNbAUVf23_1;
	wire w_dff_A_yWsghXlF1_1;
	wire w_dff_A_hKMZwiL11_1;
	wire w_dff_A_DNxx7Crx3_1;
	wire w_dff_A_7lesqXUP2_1;
	wire w_dff_A_oWZPXYVD3_1;
	wire w_dff_A_pykIj7No3_1;
	wire w_dff_A_SeyeNzVn7_1;
	wire w_dff_A_xwhHnZWD3_1;
	wire w_dff_A_itjcwYbR2_1;
	wire w_dff_B_98i5q6i27_1;
	wire w_dff_B_Fh22ZAkX4_1;
	wire w_dff_B_FeHEPAxG1_1;
	wire w_dff_B_VdMhXcsq0_1;
	wire w_dff_B_O3wFpCtC9_1;
	wire w_dff_B_XAIlAHcE4_1;
	wire w_dff_B_Q9VHc7v35_1;
	wire w_dff_B_HXF8qjwB7_1;
	wire w_dff_B_Pqnhn7Bk7_1;
	wire w_dff_B_ITdeaySm6_1;
	wire w_dff_B_wSBEcLQg8_1;
	wire w_dff_B_KKewNWnA2_1;
	wire w_dff_B_uLOxlXOx2_1;
	wire w_dff_B_Wi4txK3w5_0;
	wire w_dff_B_CjUudyhj4_0;
	wire w_dff_B_GVUNx34g6_0;
	wire w_dff_B_Ld7x9OEn2_0;
	wire w_dff_B_qM2GOlFb8_0;
	wire w_dff_B_dVl6r7ub5_0;
	wire w_dff_B_WkKibG8O6_0;
	wire w_dff_B_LXJBMZb92_0;
	wire w_dff_B_b1Uc1eAx7_0;
	wire w_dff_B_9ji28POX1_0;
	wire w_dff_B_XuXI86Ur9_0;
	wire w_dff_A_gKVDurJ62_1;
	wire w_dff_A_1sc3yxxC3_1;
	wire w_dff_A_cu9ioHt23_1;
	wire w_dff_A_0mqTJW9U4_1;
	wire w_dff_A_EIqOoX1y5_1;
	wire w_dff_A_gRxDMbuh5_1;
	wire w_dff_A_dO0tdUbf9_1;
	wire w_dff_A_wO1vKqH19_1;
	wire w_dff_A_AlW3KyGb2_1;
	wire w_dff_A_cHmjjC4Q0_1;
	wire w_dff_A_ayZfOxte6_1;
	wire w_dff_A_hBr7Bvkn6_1;
	wire w_dff_B_xRqPyWT30_1;
	wire w_dff_B_7xCgBDri0_1;
	wire w_dff_B_3zrg0aoQ8_1;
	wire w_dff_B_R4DVJwf72_1;
	wire w_dff_B_WGzgPYBE1_1;
	wire w_dff_B_sf6Vy6wZ7_1;
	wire w_dff_B_mqIlxu2V0_1;
	wire w_dff_B_BeKu9XTA9_1;
	wire w_dff_B_J2xOxtYg1_1;
	wire w_dff_B_av4IUyOg2_1;
	wire w_dff_B_8W0lI1PT1_1;
	wire w_dff_B_UBMYoQfe2_1;
	wire w_dff_B_7QMxYCto9_0;
	wire w_dff_B_M5Yd0prC2_0;
	wire w_dff_B_Vx59Mf9W3_0;
	wire w_dff_B_iMYbj4g92_0;
	wire w_dff_B_DGejjhsJ7_0;
	wire w_dff_B_CxLbiHdJ0_0;
	wire w_dff_B_CoNQfLzc0_0;
	wire w_dff_B_5Qs5fN2D5_0;
	wire w_dff_B_lZtfl94T7_0;
	wire w_dff_B_AIWOmTrF2_0;
	wire w_dff_A_79xTRdAA4_1;
	wire w_dff_A_kH0vxITY7_1;
	wire w_dff_A_u570xPwX1_1;
	wire w_dff_A_dcjzw2mt2_1;
	wire w_dff_A_5uLvVhj20_1;
	wire w_dff_A_KvJKSr7d0_1;
	wire w_dff_A_sb1lZJCh5_1;
	wire w_dff_A_t3zvyWfM6_1;
	wire w_dff_A_vjISJLyS1_1;
	wire w_dff_A_rg0cV6kt8_1;
	wire w_dff_A_KvEs2OMJ1_1;
	wire w_dff_B_WWBzEK2t8_1;
	wire w_dff_B_jz9KcFHN7_1;
	wire w_dff_B_QwGmC3jj4_1;
	wire w_dff_B_DNqCeEMs2_1;
	wire w_dff_B_GIAzMXZK9_1;
	wire w_dff_B_sTdSgllS3_1;
	wire w_dff_B_bUz2w9d47_1;
	wire w_dff_B_g6IpYB3m0_1;
	wire w_dff_B_zsifSQsn5_1;
	wire w_dff_B_8ztmIV7a7_1;
	wire w_dff_B_cv02aKdX6_0;
	wire w_dff_B_Cl3RWvNn9_0;
	wire w_dff_B_QvEk66Jp5_0;
	wire w_dff_B_Dd3l0Fwh4_0;
	wire w_dff_B_HwVYhdoW9_0;
	wire w_dff_B_ywhYHoMz5_0;
	wire w_dff_B_3WLio9ZI0_0;
	wire w_dff_B_NWY9YSYe7_0;
	wire w_dff_A_Fk4Cu5155_1;
	wire w_dff_A_KZreOOdV9_1;
	wire w_dff_A_WGY0EMid1_1;
	wire w_dff_A_KFmSYE1H1_1;
	wire w_dff_A_uJ5HZv8s5_1;
	wire w_dff_A_1EExzx8z2_1;
	wire w_dff_A_do84FDrb8_1;
	wire w_dff_A_c7TN3Ezh7_1;
	wire w_dff_A_G80OTdUX1_1;
	wire w_dff_B_AA6gCB0m2_1;
	wire w_dff_B_UpwJJE7z9_1;
	wire w_dff_B_pUJ00lGB5_1;
	wire w_dff_B_rwfAv5aH8_1;
	wire w_dff_B_UuU8hRCC1_1;
	wire w_dff_B_HEkJ4m610_1;
	wire w_dff_B_pd6g6nrz3_1;
	wire w_dff_B_D3AzhsqY2_1;
	wire w_dff_B_611Z2rBw0_0;
	wire w_dff_B_F8XMhViI5_0;
	wire w_dff_B_mm7wYaZM8_0;
	wire w_dff_B_rNhRn8C72_0;
	wire w_dff_B_6qUBbKno5_0;
	wire w_dff_B_J0oQAQk06_0;
	wire w_dff_A_KrEMh2ET3_1;
	wire w_dff_A_qs22pyxv8_1;
	wire w_dff_A_yOIXtJdL9_1;
	wire w_dff_A_tRTdw8lN6_1;
	wire w_dff_A_pniuvVG98_1;
	wire w_dff_A_GVrYQgqz7_1;
	wire w_dff_A_FdAfEhwx6_1;
	wire w_dff_B_s5VMcwp71_1;
	wire w_dff_B_7181w4Jd4_1;
	wire w_dff_B_XLyrQERS0_1;
	wire w_dff_B_jQnhG3HK0_1;
	wire w_dff_B_q7HmttER1_1;
	wire w_dff_B_QfljtKyF7_1;
	wire w_dff_B_ubHAw9xw6_1;
	wire w_dff_B_A09hQSLQ0_0;
	wire w_dff_B_YJMp2cQO5_0;
	wire w_dff_B_D1ub6vNA8_0;
	wire w_dff_B_KZXJQL4Y4_0;
	wire w_dff_B_KxTD4Scz6_0;
	wire w_dff_A_cvJhLKV41_1;
	wire w_dff_A_9T6Ai5Ii2_1;
	wire w_dff_A_NmxiMzk67_1;
	wire w_dff_A_h258285L2_1;
	wire w_dff_A_peibwPQ52_1;
	wire w_dff_A_q7PYhXqR0_1;
	wire w_dff_B_SFLsw30A8_1;
	wire w_dff_B_CbvifFGY4_1;
	wire w_dff_B_HGeey1hP9_1;
	wire w_dff_B_mSLgcSV87_1;
	wire w_dff_B_NnlQCR6R8_1;
	wire w_dff_B_tmWz7Xxw0_1;
	wire w_dff_B_fKEZf45O2_0;
	wire w_dff_B_TW7vS4AY7_0;
	wire w_dff_B_oJtqagUn2_0;
	wire w_dff_B_cQ4vJJdm6_0;
	wire w_dff_A_xnWN3iB84_1;
	wire w_dff_A_pSshbNdD7_1;
	wire w_dff_A_xpEv0tNt5_1;
	wire w_dff_A_7FZ7qAsX5_1;
	wire w_dff_A_uVFeJtGu4_1;
	wire w_dff_B_3yIdB2n87_1;
	wire w_dff_B_ARe2uTSg8_1;
	wire w_dff_B_Koc5iBCH3_1;
	wire w_dff_A_hO5k5axH8_0;
	wire w_dff_A_J7L0F21u0_0;
	wire w_dff_B_ybojhGAX3_1;
	wire w_dff_A_kaFjA6Cr4_0;
	wire w_dff_B_fYgRh1hF7_1;
	wire w_dff_A_jiOGZly09_1;
	wire w_dff_B_CVkOlKTy6_2;
	wire w_dff_B_ZO5Jnt0Y5_1;
	wire w_dff_A_BHRY0G6L4_0;
	wire w_dff_A_wpcAzBN75_0;
	wire w_dff_A_P1kbRSS35_0;
	wire w_dff_A_RCxcO2ug9_0;
	wire w_dff_A_LRMM7CMf9_0;
	wire w_dff_A_GmkW7RrH2_0;
	wire w_dff_A_TrKXhuUI6_0;
	wire w_dff_A_0z2Gcrvs8_0;
	wire w_dff_A_Y6HhZCh19_0;
	wire w_dff_A_o3wO0o3u5_0;
	wire w_dff_A_LivJCd1u6_0;
	wire w_dff_A_Xe2cx39M6_0;
	wire w_dff_A_YIqSVSig2_0;
	wire w_dff_A_9wrzYiy57_0;
	wire w_dff_A_LFKxwgSu4_0;
	wire w_dff_A_g7wEpjmQ2_0;
	wire w_dff_A_IHC192zf5_0;
	wire w_dff_A_D7p12W4g6_0;
	wire w_dff_A_4FcbHW3v2_0;
	wire w_dff_A_0y68ajuR1_0;
	wire w_dff_A_6pzbKutD4_0;
	wire w_dff_A_EKGbOPrh9_0;
	wire w_dff_A_q1Gqd3m25_0;
	wire w_dff_A_8LyXd5j84_0;
	wire w_dff_A_3AOMD8TQ9_0;
	wire w_dff_A_vQbkMacA7_0;
	wire w_dff_A_hiFGNQmS1_0;
	wire w_dff_A_jCZtZdpQ0_0;
	wire w_dff_A_QE99YOKC2_0;
	wire w_dff_A_TSglZsyy4_0;
	wire w_dff_A_6f52oQ1b9_0;
	wire w_dff_A_JOYxbMpT4_0;
	wire w_dff_A_AhDiPKMt8_0;
	wire w_dff_A_kbLrsGem1_0;
	wire w_dff_A_0Hv1oFsx9_0;
	wire w_dff_A_RGXyUJYb4_0;
	wire w_dff_A_QIAOY69L9_0;
	wire w_dff_A_8MlR8qzX8_0;
	wire w_dff_A_suCZ3rK21_0;
	wire w_dff_A_gsJszbJZ1_0;
	wire w_dff_A_6fvcXd5l6_0;
	wire w_dff_A_gJAijCqu7_0;
	wire w_dff_A_QqOo8jfq1_0;
	wire w_dff_A_7cq0XO5c0_1;
	wire w_dff_B_2rNmKVuM2_1;
	wire w_dff_A_uoslVDBg8_0;
	wire w_dff_A_zWy9C9333_0;
	wire w_dff_A_lY29bOSw2_0;
	wire w_dff_A_gEdXHpU48_0;
	wire w_dff_A_0ky2T2yD0_0;
	wire w_dff_A_2UEEXuuF6_0;
	wire w_dff_A_nBI47ZtZ7_0;
	wire w_dff_A_5hDO9RcP7_0;
	wire w_dff_A_ho6tuuao7_0;
	wire w_dff_A_EfUSJx668_0;
	wire w_dff_A_LsyUGUE08_0;
	wire w_dff_A_jEAMMhjg7_0;
	wire w_dff_A_4QyU7vqQ7_0;
	wire w_dff_A_HfpsZWzC6_0;
	wire w_dff_A_xCvJr1wS9_0;
	wire w_dff_A_2AXeviiu6_0;
	wire w_dff_A_4OVFI3vb9_0;
	wire w_dff_A_fVwu7g6j9_0;
	wire w_dff_A_JnyOuQ9M1_0;
	wire w_dff_A_M4R8nM4p8_0;
	wire w_dff_A_Sr4zIyDc6_0;
	wire w_dff_A_rxkKefHw0_0;
	wire w_dff_A_OhoYsm5C6_0;
	wire w_dff_A_mEaqBEgc3_0;
	wire w_dff_A_Ojo1izpC9_0;
	wire w_dff_A_1WLY8Ti45_0;
	wire w_dff_A_IOv8kBW68_0;
	wire w_dff_A_5YeZap0Y0_0;
	wire w_dff_A_13EBlcFb1_0;
	wire w_dff_A_sotR9M5P8_0;
	wire w_dff_A_8Xlhih6v5_0;
	wire w_dff_A_0pmBw9Or1_0;
	wire w_dff_A_2YnWPVwZ1_0;
	wire w_dff_A_r9xvjQIv1_0;
	wire w_dff_A_DVBhDspW3_0;
	wire w_dff_A_bEXCFuCA2_0;
	wire w_dff_A_Dnaihokf7_0;
	wire w_dff_A_T6mgB7AE0_0;
	wire w_dff_A_Ob2Y3P6o2_0;
	wire w_dff_A_N18EMJBx6_0;
	wire w_dff_A_eo9lZxUw1_1;
	wire w_dff_B_KRtJVCPj7_1;
	wire w_dff_B_SkNhUAOP6_1;
	wire w_dff_B_Pt3fOwyy9_1;
	wire w_dff_B_5n8PwDHO6_1;
	wire w_dff_B_W9a4W4Wo1_1;
	wire w_dff_B_8OsFalwC3_1;
	wire w_dff_B_tzJsuKty0_1;
	wire w_dff_B_QlU18psY4_1;
	wire w_dff_B_cpNMblWV8_1;
	wire w_dff_B_mkqVkWJV9_1;
	wire w_dff_B_q58fuMNR0_1;
	wire w_dff_B_J0HIMT0P0_1;
	wire w_dff_B_zYfrQ9Hc6_1;
	wire w_dff_B_pdnRk0Ik7_1;
	wire w_dff_B_HhqsTWYQ0_1;
	wire w_dff_B_oFf4QXRh8_1;
	wire w_dff_B_PDqLJ4RM0_1;
	wire w_dff_B_jq8F6DXk1_1;
	wire w_dff_B_BvUPDUCv2_1;
	wire w_dff_B_MXakd8hJ1_1;
	wire w_dff_B_OTERYf4q8_1;
	wire w_dff_B_QehL6McB4_1;
	wire w_dff_B_tLCza84k3_1;
	wire w_dff_B_mXNHgVYp6_1;
	wire w_dff_B_9pNqoitb1_1;
	wire w_dff_B_hnLjxhIU1_1;
	wire w_dff_B_dQXMrhXN2_1;
	wire w_dff_B_1zxBwxWi4_1;
	wire w_dff_B_EH10RSXA9_1;
	wire w_dff_B_26zndpjw6_1;
	wire w_dff_B_ZA0QdNd89_1;
	wire w_dff_B_TMYzmnVo7_1;
	wire w_dff_B_FcazK6Hj8_1;
	wire w_dff_B_s9RCwLyC4_1;
	wire w_dff_B_O4Ixz7Ng6_1;
	wire w_dff_B_6wcSrPEr9_1;
	wire w_dff_B_Xym03pKl7_1;
	wire w_dff_A_FGwVRWCg9_0;
	wire w_dff_A_EJGcBJLE4_0;
	wire w_dff_A_RBoRpCHR1_0;
	wire w_dff_A_HHoIQMvM6_0;
	wire w_dff_A_r7T5RlNr6_0;
	wire w_dff_A_bmzqZhWS1_0;
	wire w_dff_A_JNPCvNGk0_0;
	wire w_dff_A_6kwrgV8p6_0;
	wire w_dff_A_IMdurQtH8_0;
	wire w_dff_A_CGN8djJ72_0;
	wire w_dff_A_ATty5JQI0_0;
	wire w_dff_A_PMALUlyS7_0;
	wire w_dff_A_8KLsGwWw6_0;
	wire w_dff_A_0YcmvCC04_0;
	wire w_dff_A_WgzJKzss6_0;
	wire w_dff_A_hSsYlydL9_0;
	wire w_dff_A_vIeHjNLH9_0;
	wire w_dff_A_SSQOAqDK9_0;
	wire w_dff_A_5rSlmiP55_0;
	wire w_dff_A_SLsPsEKY3_0;
	wire w_dff_A_RrwU77qV7_0;
	wire w_dff_A_ncFlE6jN3_0;
	wire w_dff_A_bHUUfagv2_0;
	wire w_dff_A_YsItLTIa6_0;
	wire w_dff_A_La0IhG493_0;
	wire w_dff_A_zyJjB6n00_0;
	wire w_dff_A_LTvM492u1_0;
	wire w_dff_A_lYeOZ6IH2_0;
	wire w_dff_A_WNnuKsmE2_0;
	wire w_dff_A_rNzVcCAP3_0;
	wire w_dff_A_vkFHbpTP2_0;
	wire w_dff_A_G6tQPmgk4_0;
	wire w_dff_A_TsaPcj4A5_0;
	wire w_dff_A_GbHM12Y08_0;
	wire w_dff_A_XqJgMGV55_0;
	wire w_dff_A_cPQU0PL80_0;
	wire w_dff_A_CEOAP1Il9_0;
	wire w_dff_A_WtcaqWte1_1;
	wire w_dff_B_6SyICT3r3_1;
	wire w_dff_B_zc7ZRKXU9_1;
	wire w_dff_B_0bzIwj9I4_1;
	wire w_dff_B_CpnOqE7C3_1;
	wire w_dff_B_pYBHqoFn1_1;
	wire w_dff_B_tAaFqgc84_1;
	wire w_dff_B_2xQqBtlx1_1;
	wire w_dff_B_uZet1faX3_1;
	wire w_dff_B_0SWNfy8y3_1;
	wire w_dff_B_CLQmzCwo2_1;
	wire w_dff_B_BPdERJ4A5_1;
	wire w_dff_B_Pa7lDxO18_1;
	wire w_dff_B_WssyBeGf5_1;
	wire w_dff_B_cTch3KW05_1;
	wire w_dff_B_J5E5CX8w7_1;
	wire w_dff_B_U47cGXxX3_1;
	wire w_dff_B_yy7jdFRp9_1;
	wire w_dff_B_2ZKnmGzf5_1;
	wire w_dff_B_2XQENLZS6_1;
	wire w_dff_B_7aU93EXp4_1;
	wire w_dff_B_VD49i5sc8_1;
	wire w_dff_B_xQ9J6wBl5_1;
	wire w_dff_B_WrYBGyXo8_1;
	wire w_dff_B_kGvVOY530_1;
	wire w_dff_B_p5LiN9Fo0_1;
	wire w_dff_B_XeT5F3Px7_1;
	wire w_dff_B_DOBIEwb76_1;
	wire w_dff_B_OTbd4oDl6_1;
	wire w_dff_B_I8bgpPvD4_1;
	wire w_dff_B_4AR1He6A7_1;
	wire w_dff_B_Uf638gyY1_1;
	wire w_dff_B_XRfW8VhR6_1;
	wire w_dff_B_GvGucZMJ3_1;
	wire w_dff_B_gDaYprKw4_1;
	wire w_dff_A_4JA57ErZ2_0;
	wire w_dff_A_4rijDBqq0_0;
	wire w_dff_A_xhNGnLFM1_0;
	wire w_dff_A_GZrW29ii7_0;
	wire w_dff_A_BAOEhlF92_0;
	wire w_dff_A_kRYDu1yu0_0;
	wire w_dff_A_Oi2TLuuA0_0;
	wire w_dff_A_fqhrYLO25_0;
	wire w_dff_A_w1NaCkg98_0;
	wire w_dff_A_jxxPaWK55_0;
	wire w_dff_A_0uN47Fnk6_0;
	wire w_dff_A_UXHYIZEl4_0;
	wire w_dff_A_w4iiWhvu1_0;
	wire w_dff_A_LpeGGcxZ3_0;
	wire w_dff_A_FWFJcQop7_0;
	wire w_dff_A_Ifu3STPv1_0;
	wire w_dff_A_4YkROka03_0;
	wire w_dff_A_iDS9mbmt7_0;
	wire w_dff_A_czW4u29l3_0;
	wire w_dff_A_l0799hok5_0;
	wire w_dff_A_iXQZhpRQ8_0;
	wire w_dff_A_DKSkIHZw6_0;
	wire w_dff_A_rUkZxJ0X8_0;
	wire w_dff_A_Ap06mBVh1_0;
	wire w_dff_A_66OlGLJO1_0;
	wire w_dff_A_z14vIt9g8_0;
	wire w_dff_A_RrB7piCl6_0;
	wire w_dff_A_D9IVdaYP7_0;
	wire w_dff_A_CfPw4iH52_0;
	wire w_dff_A_OWeJAIRQ9_0;
	wire w_dff_A_YAyVEApa5_0;
	wire w_dff_A_RSbttYl69_0;
	wire w_dff_A_MdNDT2Xl1_0;
	wire w_dff_A_mEqOSiLQ7_0;
	wire w_dff_A_ISeNVaNj6_1;
	wire w_dff_B_ne3tCZix4_1;
	wire w_dff_B_phupOrTO3_1;
	wire w_dff_B_7C3TQTWm9_1;
	wire w_dff_B_EtcckvmZ5_1;
	wire w_dff_B_G4U64aVO7_1;
	wire w_dff_B_sM15BQ009_1;
	wire w_dff_B_AzuYEjPK2_1;
	wire w_dff_B_JGkZPThU5_1;
	wire w_dff_B_23pPFu9Z4_1;
	wire w_dff_B_cQFhJUDS3_1;
	wire w_dff_B_p2mqKVMX0_1;
	wire w_dff_B_6tXR47171_1;
	wire w_dff_B_TUu0ZKo81_1;
	wire w_dff_B_kqQ9lN4g8_1;
	wire w_dff_B_d69QeIeX9_1;
	wire w_dff_B_NaqEPx3J0_1;
	wire w_dff_B_gp3UP3RY5_1;
	wire w_dff_B_ub8Uo2Id6_1;
	wire w_dff_B_PHXdFdkm2_1;
	wire w_dff_B_1OiyW2Kp0_1;
	wire w_dff_B_nW7ctQvP8_1;
	wire w_dff_B_A43KquRh1_1;
	wire w_dff_B_HbziTMfy1_1;
	wire w_dff_B_7O4IIOVB5_1;
	wire w_dff_B_f7HCLSeY0_1;
	wire w_dff_B_wjf1W34s0_1;
	wire w_dff_B_UOBfBc6k4_1;
	wire w_dff_B_QYZyfPO62_1;
	wire w_dff_B_Qw7lEFNL7_1;
	wire w_dff_B_NRDofYYa6_1;
	wire w_dff_B_7wRTG4kK2_1;
	wire w_dff_A_a8Fwb5RZ4_0;
	wire w_dff_A_TyAhhCyJ2_0;
	wire w_dff_A_wfj6IsTs4_0;
	wire w_dff_A_ITadPbkD3_0;
	wire w_dff_A_yPNTjDHC3_0;
	wire w_dff_A_PEkuYYf89_0;
	wire w_dff_A_z3YKOYsy5_0;
	wire w_dff_A_Nvfqj2z84_0;
	wire w_dff_A_l8qElnG82_0;
	wire w_dff_A_AfynoxTc3_0;
	wire w_dff_A_pTqbHSPV1_0;
	wire w_dff_A_VMEOnLgi9_0;
	wire w_dff_A_018a6RRB4_0;
	wire w_dff_A_nwjoImeu3_0;
	wire w_dff_A_qVk9fyOs2_0;
	wire w_dff_A_gK6cTBAU6_0;
	wire w_dff_A_fcRJirG81_0;
	wire w_dff_A_th70luBO7_0;
	wire w_dff_A_plS3fxfc6_0;
	wire w_dff_A_Oed7hk8V7_0;
	wire w_dff_A_zZPHYFOA2_0;
	wire w_dff_A_HEEn2e2t3_0;
	wire w_dff_A_8ajl39RZ5_0;
	wire w_dff_A_AZwe0iB83_0;
	wire w_dff_A_GgQ0PZpw2_0;
	wire w_dff_A_VbVH6lDI6_0;
	wire w_dff_A_un1r5UeO9_0;
	wire w_dff_A_L4UuEmJk4_0;
	wire w_dff_A_7j7km2QS2_0;
	wire w_dff_A_nYcqxPaO9_0;
	wire w_dff_A_YkPo2Xyi0_0;
	wire w_dff_A_SLB4Z28D3_1;
	wire w_dff_B_KVsXI5t10_1;
	wire w_dff_B_uhLZpc4R5_1;
	wire w_dff_B_TAReCawD2_1;
	wire w_dff_B_Hm4SJaXH4_1;
	wire w_dff_B_zJCXU40K9_1;
	wire w_dff_B_63lPQyr87_1;
	wire w_dff_B_VJHijFr08_1;
	wire w_dff_B_f2JXMnTy5_1;
	wire w_dff_B_zF69YUCj7_1;
	wire w_dff_B_oM0crne45_1;
	wire w_dff_B_HHSEyHm83_1;
	wire w_dff_B_2BYuB0uB1_1;
	wire w_dff_B_ZjYasMWt8_1;
	wire w_dff_B_B56FRRMA6_1;
	wire w_dff_B_KJAC98oo5_1;
	wire w_dff_B_DWT7UjjS2_1;
	wire w_dff_B_3k25Bayc1_1;
	wire w_dff_B_HaEkyVTz3_1;
	wire w_dff_B_lwac3JkV3_1;
	wire w_dff_B_WETmanAY0_1;
	wire w_dff_B_EjNMBUc71_1;
	wire w_dff_B_q9ZMHwLB5_1;
	wire w_dff_B_LGgs0VRt4_1;
	wire w_dff_B_mfJ2Qxfl4_1;
	wire w_dff_B_6E035ANg8_1;
	wire w_dff_B_bDqslVgs1_1;
	wire w_dff_B_KH04q8iw5_1;
	wire w_dff_B_yG4BhU3r1_1;
	wire w_dff_A_YmAFLElN3_0;
	wire w_dff_A_rCzgkMsT7_0;
	wire w_dff_A_MaXF1dXn4_0;
	wire w_dff_A_aKlxPGwU8_0;
	wire w_dff_A_GHNJICnn8_0;
	wire w_dff_A_fsfAiiJf9_0;
	wire w_dff_A_3OoPisMW8_0;
	wire w_dff_A_B69rtH2e2_0;
	wire w_dff_A_UyXZTCIt6_0;
	wire w_dff_A_jfWBjy941_0;
	wire w_dff_A_8MroAHsf3_0;
	wire w_dff_A_wpRmbtLm3_0;
	wire w_dff_A_mgEwifOG1_0;
	wire w_dff_A_dn9v5nAG5_0;
	wire w_dff_A_e3Fxy71B5_0;
	wire w_dff_A_WNTsDQSh0_0;
	wire w_dff_A_qBVO1gIB2_0;
	wire w_dff_A_9wPQLlci9_0;
	wire w_dff_A_TU7BpV7D4_0;
	wire w_dff_A_9c7n4xI33_0;
	wire w_dff_A_Ff3Shiyc3_0;
	wire w_dff_A_8qoe3A5D4_0;
	wire w_dff_A_aOXGokKK0_0;
	wire w_dff_A_5pXi0zUh1_0;
	wire w_dff_A_Ieuc4sDw6_0;
	wire w_dff_A_KJ01cv9u3_0;
	wire w_dff_A_L9gT24z83_0;
	wire w_dff_A_d3MCYPN24_0;
	wire w_dff_A_CXCuRGa09_1;
	wire w_dff_B_PtvS5JU96_1;
	wire w_dff_B_mbw1FOW70_1;
	wire w_dff_B_Nqg9vPeh8_1;
	wire w_dff_B_0MrTnKSn4_1;
	wire w_dff_B_ymdm0y3i6_1;
	wire w_dff_B_ynY3OOpW1_1;
	wire w_dff_B_YG9b6rev9_1;
	wire w_dff_B_vsmfJZEW6_1;
	wire w_dff_B_j9sUOswq7_1;
	wire w_dff_B_ACbfjm224_1;
	wire w_dff_B_Oju7GHiL1_1;
	wire w_dff_B_oOKxsGNp6_1;
	wire w_dff_B_McWBFlO55_1;
	wire w_dff_B_CkO3vphw4_1;
	wire w_dff_B_kvglClJI2_1;
	wire w_dff_B_xBQ5i8mo0_1;
	wire w_dff_B_90NTLAwQ7_1;
	wire w_dff_B_74P4vBwh1_1;
	wire w_dff_B_Pmorb9qW5_1;
	wire w_dff_B_cv4ZrcvC3_1;
	wire w_dff_B_PZphXTer8_1;
	wire w_dff_B_kZFmRd181_1;
	wire w_dff_B_YDqN3Te69_1;
	wire w_dff_B_qslerWkk7_1;
	wire w_dff_B_ZpA9JmNq8_1;
	wire w_dff_A_s5OHmhHg5_0;
	wire w_dff_A_SCFaBpoW3_0;
	wire w_dff_A_FghTPP2c3_0;
	wire w_dff_A_jbUXCWpC1_0;
	wire w_dff_A_WaOllnxS3_0;
	wire w_dff_A_NmYipz4U3_0;
	wire w_dff_A_1QXapqIj6_0;
	wire w_dff_A_SvPGsJvD4_0;
	wire w_dff_A_dqDgnsry8_0;
	wire w_dff_A_OOQilvVf2_0;
	wire w_dff_A_C59HJymX4_0;
	wire w_dff_A_WvzSRdQc3_0;
	wire w_dff_A_YVfE3w2d2_0;
	wire w_dff_A_RG13SCtY3_0;
	wire w_dff_A_M4fiS7nu5_0;
	wire w_dff_A_vGy1t0No1_0;
	wire w_dff_A_MSszrTlK3_0;
	wire w_dff_A_Xzih0xJN7_0;
	wire w_dff_A_pT8unBlS1_0;
	wire w_dff_A_4hT35RRM9_0;
	wire w_dff_A_X20zWPiF9_0;
	wire w_dff_A_iOu9PlQg8_0;
	wire w_dff_A_PdF60ZML1_0;
	wire w_dff_A_Hgv2ssJz7_0;
	wire w_dff_A_bZ4o1eNL3_0;
	wire w_dff_A_UNh2eDPN7_1;
	wire w_dff_B_446mc0tf3_1;
	wire w_dff_B_beI0umwh0_1;
	wire w_dff_B_diEnk7oY4_1;
	wire w_dff_B_6b2SGBvD7_1;
	wire w_dff_B_yMtqXUPN9_1;
	wire w_dff_B_MtD0yVFQ5_1;
	wire w_dff_B_DjsAcU4Y7_1;
	wire w_dff_B_GbhPqi6W5_1;
	wire w_dff_B_Eee7ff629_1;
	wire w_dff_B_mTMfebD38_1;
	wire w_dff_B_czrf5Jbs5_1;
	wire w_dff_B_6xEokzLD9_1;
	wire w_dff_B_cZZmQE5Q3_1;
	wire w_dff_B_HUTuF5Xa7_1;
	wire w_dff_B_WAakYAi93_1;
	wire w_dff_B_Snh2BeM71_1;
	wire w_dff_B_jQrVFQ9k5_1;
	wire w_dff_B_pjUBAyGf4_1;
	wire w_dff_B_QwwPHf2d4_1;
	wire w_dff_B_WkPDkMw68_1;
	wire w_dff_B_tbVrxYkZ0_1;
	wire w_dff_B_3wO4YlSX2_1;
	wire w_dff_A_4CNz0Ejq0_0;
	wire w_dff_A_obpJO30q9_0;
	wire w_dff_A_dZNstbAX2_0;
	wire w_dff_A_YkU4HKhe2_0;
	wire w_dff_A_ZOYfEGjf3_0;
	wire w_dff_A_j1eut0b90_0;
	wire w_dff_A_lHk6dL8F3_0;
	wire w_dff_A_Ad7PnX578_0;
	wire w_dff_A_bNdnQQHs9_0;
	wire w_dff_A_E7ZxRcSB1_0;
	wire w_dff_A_u10TAW412_0;
	wire w_dff_A_XCyAKAhL4_0;
	wire w_dff_A_ALQuVkGo2_0;
	wire w_dff_A_4CWDRDKO7_0;
	wire w_dff_A_XLKzj4l83_0;
	wire w_dff_A_bPCdQkeh4_0;
	wire w_dff_A_LsuONHZD2_0;
	wire w_dff_A_MN3hfL696_0;
	wire w_dff_A_vvbD3iRi9_0;
	wire w_dff_A_miFEZiZL9_0;
	wire w_dff_A_3vAgnj9q3_0;
	wire w_dff_A_xFr8Ne6S7_0;
	wire w_dff_A_iki1Wsv18_1;
	wire w_dff_B_oV4xYXZt9_1;
	wire w_dff_B_dvri7vgW5_1;
	wire w_dff_B_W5EZtmxx4_1;
	wire w_dff_B_CZsJfKZq6_1;
	wire w_dff_B_pnDOXqfT8_1;
	wire w_dff_B_aLpKKp8R1_1;
	wire w_dff_B_8RYHX3332_1;
	wire w_dff_B_p1Jo63Pu7_1;
	wire w_dff_B_6ykyMfno0_1;
	wire w_dff_B_Zl2tUOaP3_1;
	wire w_dff_B_GtgmVF3a7_1;
	wire w_dff_B_3mMvkFAu6_1;
	wire w_dff_B_QT86LUp77_1;
	wire w_dff_B_cnpNgyWw9_1;
	wire w_dff_B_2RZeftVy2_1;
	wire w_dff_B_IM95GAQg2_1;
	wire w_dff_B_r1CnYXuj2_1;
	wire w_dff_B_mPvqQbQg9_1;
	wire w_dff_B_cjBnXVB24_1;
	wire w_dff_A_96bRC0UK7_0;
	wire w_dff_A_kZEQKxM98_0;
	wire w_dff_A_sWdKdqXm3_0;
	wire w_dff_A_pCJ7f2W59_0;
	wire w_dff_A_PrBPUt7H2_0;
	wire w_dff_A_MGBfStTH7_0;
	wire w_dff_A_2n2Apw1D5_0;
	wire w_dff_A_8CJh9Ckb5_0;
	wire w_dff_A_RIAETzaY3_0;
	wire w_dff_A_543fqMmN2_0;
	wire w_dff_A_vK5bv9kC6_0;
	wire w_dff_A_CFUJTBnW1_0;
	wire w_dff_A_sErRkcCl4_0;
	wire w_dff_A_j6nAlm6e6_0;
	wire w_dff_A_57y9QFPw7_0;
	wire w_dff_A_3feiKSxl8_0;
	wire w_dff_A_w8zJmMbx2_0;
	wire w_dff_A_MbeXN5xh0_0;
	wire w_dff_A_hTpwivnN8_0;
	wire w_dff_A_T4cDbbGE9_1;
	wire w_dff_B_9KhjrN6S2_1;
	wire w_dff_B_QAm33Y5Q5_1;
	wire w_dff_B_r1jZANC11_1;
	wire w_dff_B_pCJkc8a62_1;
	wire w_dff_B_hLFgJVMM0_1;
	wire w_dff_B_KvRu4fax7_1;
	wire w_dff_B_RT4vUHdy6_1;
	wire w_dff_B_R2DSn46J8_1;
	wire w_dff_B_SL2Sb3oK8_1;
	wire w_dff_B_LbnUKm7O3_1;
	wire w_dff_B_ltJw6WsM4_1;
	wire w_dff_B_Nv1OoUv25_1;
	wire w_dff_B_cjOZ3a0d7_1;
	wire w_dff_B_2i1rmVbG7_1;
	wire w_dff_B_e1S54b0o3_1;
	wire w_dff_B_ARqMBHW71_1;
	wire w_dff_A_jN1yvcrQ3_0;
	wire w_dff_A_RaUhwoHn2_0;
	wire w_dff_A_HjnLsjbO2_0;
	wire w_dff_A_ToH3PObi3_0;
	wire w_dff_A_Oghdby3S3_0;
	wire w_dff_A_G8nSVk0x4_0;
	wire w_dff_A_YAxoQRoe4_0;
	wire w_dff_A_S6NMjrMg7_0;
	wire w_dff_A_WajgXwx04_0;
	wire w_dff_A_T6yBKPDw4_0;
	wire w_dff_A_kNDyUytj8_0;
	wire w_dff_A_LVPkdWoh0_0;
	wire w_dff_A_CICRyl5C9_0;
	wire w_dff_A_Hy7KfI5w8_0;
	wire w_dff_A_HRTrxZWu9_0;
	wire w_dff_A_qGBbdJg55_0;
	wire w_dff_A_uD5kYzFY7_1;
	wire w_dff_B_19xdoAS41_1;
	wire w_dff_B_0SFShaYm4_1;
	wire w_dff_B_cyx4Fo573_1;
	wire w_dff_B_Af8IFqgp2_1;
	wire w_dff_B_7rXxdFcr8_1;
	wire w_dff_B_flES295I5_1;
	wire w_dff_B_eMCIV4kl0_1;
	wire w_dff_B_HoYeT0Dg5_1;
	wire w_dff_B_E5Seo1lz6_1;
	wire w_dff_B_VevoZam20_1;
	wire w_dff_B_T019ONPG9_1;
	wire w_dff_B_OMTgwC4u0_1;
	wire w_dff_B_Sr0tDaY84_1;
	wire w_dff_A_Y8MDE0nn7_0;
	wire w_dff_A_y5Wih8TQ2_0;
	wire w_dff_A_R3EBK8zM4_0;
	wire w_dff_A_TKCT3uPW7_0;
	wire w_dff_A_AYHCPS5a0_0;
	wire w_dff_A_BW5oXrDJ0_0;
	wire w_dff_A_B2tNOhAu4_0;
	wire w_dff_A_GWCOKTZh8_0;
	wire w_dff_A_xYE3SDwP0_0;
	wire w_dff_A_7xIgJLIw6_0;
	wire w_dff_A_hzBWj4kg0_0;
	wire w_dff_A_2dQSuDDW1_0;
	wire w_dff_A_Kob3NXpf4_0;
	wire w_dff_A_MTOSucTE3_1;
	wire w_dff_B_TNm26uXl7_1;
	wire w_dff_B_vJUMpkoL3_1;
	wire w_dff_B_sZFoQiwo9_1;
	wire w_dff_B_hfrFw3Gl5_1;
	wire w_dff_B_FxCMNQb69_1;
	wire w_dff_B_moLoIsf50_1;
	wire w_dff_B_o2XwuzLU6_1;
	wire w_dff_B_8sbivfWl9_1;
	wire w_dff_B_UaMuF6AQ2_1;
	wire w_dff_B_UhHJoqrF3_1;
	wire w_dff_A_G8vsu7JU5_0;
	wire w_dff_A_UfYd6nfG4_0;
	wire w_dff_A_JLIULioC0_0;
	wire w_dff_A_95S42CIv1_0;
	wire w_dff_A_xJWFmSS82_0;
	wire w_dff_A_mI1FmnB74_0;
	wire w_dff_A_6yzDuOo62_0;
	wire w_dff_A_WeLQMx1r3_0;
	wire w_dff_A_V7osYO1T2_0;
	wire w_dff_A_qKRfbRCj6_0;
	wire w_dff_A_Hwo7FDkD5_1;
	wire w_dff_B_PjyqkwbN1_1;
	wire w_dff_B_lpuBoLUN7_1;
	wire w_dff_B_MFL0n9fK3_1;
	wire w_dff_B_gENoNltn3_1;
	wire w_dff_B_Z4EjBICu4_1;
	wire w_dff_B_VfglReMp4_1;
	wire w_dff_B_LscLupag7_1;
	wire w_dff_A_NR91Qro00_0;
	wire w_dff_A_tlL3Ex4Y2_0;
	wire w_dff_A_avBnkoxX8_0;
	wire w_dff_A_JVsq5GdX6_0;
	wire w_dff_A_hEoXENyr3_0;
	wire w_dff_A_6guS20r26_0;
	wire w_dff_A_zLcH8Jq08_0;
	wire w_dff_A_DRCi3GWz7_1;
	wire w_dff_B_XKBdWjFg5_1;
	wire w_dff_B_8WETelJ59_1;
	wire w_dff_B_x4Y6O9rC9_1;
	wire w_dff_B_QQCVQAKW5_1;
	wire w_dff_B_2dDyRXUu5_2;
	wire w_dff_A_KKIkw2iX1_0;
	wire w_dff_A_JvxhZenG3_0;
	wire w_dff_A_fDnV6WPg1_0;
	wire w_dff_A_fEHBPXtO2_0;
	wire w_dff_B_rhRcGDUD6_0;
	wire w_dff_A_TQJWSXqW0_0;
	wire w_dff_A_UFSzZaHP3_0;
	wire w_dff_A_yNR5ZAP00_1;
	wire w_dff_B_Hl1lC4wT5_1;
	wire w_dff_B_rZ8s8lDN4_2;
	wire w_dff_B_yp2wwtls7_2;
	wire w_dff_B_aM434uSq7_2;
	wire w_dff_B_ChjqsWof0_2;
	wire w_dff_B_bJtuTtBf9_2;
	wire w_dff_B_9iUe1dal3_2;
	wire w_dff_B_6Zp8lnp06_2;
	wire w_dff_B_CcrfbxCA1_2;
	wire w_dff_B_CSjfPYqI3_2;
	wire w_dff_B_vhrUB80L6_2;
	wire w_dff_B_7ZEVWyUE1_2;
	wire w_dff_B_iegYqkeL6_2;
	wire w_dff_B_jhQiMmtV6_2;
	wire w_dff_B_hs2IXzDu9_2;
	wire w_dff_B_h8C3J6dQ2_2;
	wire w_dff_B_Yj1TTTok5_2;
	wire w_dff_B_M4YbZoyE5_2;
	wire w_dff_B_9qkKWTqq3_2;
	wire w_dff_B_TUjygvcK5_2;
	wire w_dff_B_g6sxgFEa2_2;
	wire w_dff_B_5o3Niwzm4_2;
	wire w_dff_B_9ZriKGjR7_2;
	wire w_dff_B_ITnjLgFq3_2;
	wire w_dff_B_OTbk8dQe3_2;
	wire w_dff_B_vAy7nKbo6_2;
	wire w_dff_B_zko9G0EF9_2;
	wire w_dff_B_oewizM2L7_2;
	wire w_dff_B_18rLPyg92_2;
	wire w_dff_B_AznkhTSe5_2;
	wire w_dff_B_iRKK5uBZ5_2;
	wire w_dff_B_RDkpWgyC5_2;
	wire w_dff_B_IsAT5oNE5_2;
	wire w_dff_B_vD33Rv5p3_2;
	wire w_dff_B_rBUDOAro5_2;
	wire w_dff_B_xGeUXHEG8_2;
	wire w_dff_B_8YpdBS5l8_2;
	wire w_dff_B_GpO173Qt0_2;
	wire w_dff_B_jqf4z9hw4_2;
	wire w_dff_B_v8qrSDt55_2;
	wire w_dff_B_DqyOK3lR2_2;
	wire w_dff_B_dRj1MpAd3_2;
	wire w_dff_B_hwZ1OtS52_2;
	wire w_dff_B_uqtKeENz7_2;
	wire w_dff_A_SJbKKdsT3_0;
	wire w_dff_B_MBNG0AbL0_1;
	wire w_dff_B_3zDpu1uG9_2;
	wire w_dff_B_CHcGiAPZ2_2;
	wire w_dff_B_pJq9naAp7_2;
	wire w_dff_B_f3TDEalf0_2;
	wire w_dff_B_YHBt6OSN9_2;
	wire w_dff_B_okTx86I24_2;
	wire w_dff_B_eaiiPk1C6_2;
	wire w_dff_B_uWhg0wwL9_2;
	wire w_dff_B_p98dvSum8_2;
	wire w_dff_B_iF2JISr49_2;
	wire w_dff_B_ohKe0RqU3_2;
	wire w_dff_B_9l85lq9h1_2;
	wire w_dff_B_3lihAQWP4_2;
	wire w_dff_B_I9ogKqkI5_2;
	wire w_dff_B_okQiepVj7_2;
	wire w_dff_B_dwbuXAfJ5_2;
	wire w_dff_B_IX0RCoAP0_2;
	wire w_dff_B_3o8k60GS0_2;
	wire w_dff_B_3vCIXG629_2;
	wire w_dff_B_TrExfqNq4_2;
	wire w_dff_B_GRPf8g8Q0_2;
	wire w_dff_B_3dPtBbZp2_2;
	wire w_dff_B_Ye2pHaGy8_2;
	wire w_dff_B_Q0GEHBCq2_2;
	wire w_dff_B_9lFcFSz02_2;
	wire w_dff_B_IjHXEw4x1_2;
	wire w_dff_B_HGYISROJ9_2;
	wire w_dff_B_HJFbp7XU5_2;
	wire w_dff_B_oLNIsXrp1_2;
	wire w_dff_B_fJQXtMWB0_2;
	wire w_dff_B_fi0yePVZ9_2;
	wire w_dff_B_ZWF9xFTv5_2;
	wire w_dff_B_9mFRgacX9_2;
	wire w_dff_B_uhTGuTUp1_2;
	wire w_dff_B_yRDsDuK79_2;
	wire w_dff_B_KNAFYxlh8_2;
	wire w_dff_B_mnx6UzrJ5_2;
	wire w_dff_B_stdMvYqh0_2;
	wire w_dff_B_s9GJJHbZ7_2;
	wire w_dff_B_jdynKIxI1_2;
	wire w_dff_A_0J86BOMG3_1;
	wire w_dff_B_EdhNsq102_1;
	wire w_dff_B_IebQ4pk39_1;
	wire w_dff_B_NmxozeKk1_1;
	wire w_dff_B_K6QsIFnw8_1;
	wire w_dff_B_saJiN6wL6_1;
	wire w_dff_B_QGrHeXKe1_1;
	wire w_dff_B_7amMLWih9_1;
	wire w_dff_B_cX4LMgoZ7_1;
	wire w_dff_B_omE8ldRo9_1;
	wire w_dff_B_14GVMgo24_1;
	wire w_dff_B_CM2GwsrS9_1;
	wire w_dff_B_2OXlzZFR3_1;
	wire w_dff_B_vkoctqO24_1;
	wire w_dff_B_s0ZM7l6K6_1;
	wire w_dff_B_kAPEfvcS1_1;
	wire w_dff_B_4cMlSNKW0_1;
	wire w_dff_B_jCZPZeE45_1;
	wire w_dff_B_47NS7Vxr7_1;
	wire w_dff_B_z7yEQTDj7_1;
	wire w_dff_B_kZjTMcG31_1;
	wire w_dff_B_hX2jFXWD5_1;
	wire w_dff_B_z79omYr96_1;
	wire w_dff_B_P09nFvim3_1;
	wire w_dff_B_Q5WHh9rV8_1;
	wire w_dff_B_k9pIueEk0_1;
	wire w_dff_B_AFE9EtwD2_1;
	wire w_dff_B_m7e5fpkE5_1;
	wire w_dff_B_rBbUcQQm5_1;
	wire w_dff_B_5AqhTg7e1_1;
	wire w_dff_B_fjZHzyNI5_1;
	wire w_dff_B_fOafkO0e6_1;
	wire w_dff_B_RbOgAJPZ7_1;
	wire w_dff_B_EsJzeqQh8_1;
	wire w_dff_B_nTuVxjpI5_1;
	wire w_dff_B_WHfx4DNR3_1;
	wire w_dff_B_ANn0WTHP7_1;
	wire w_dff_B_XlmD80Zn1_1;
	wire w_dff_A_5YWEty9W9_0;
	wire w_dff_A_6XViArYY6_0;
	wire w_dff_A_D5A22Oee5_0;
	wire w_dff_A_Q2yIbwww6_0;
	wire w_dff_A_rRC4en4P9_0;
	wire w_dff_A_xj8eh06L0_0;
	wire w_dff_A_9UKn3HFl5_0;
	wire w_dff_A_o4Wctewa1_0;
	wire w_dff_A_DZnSOfM64_0;
	wire w_dff_A_wnia88V73_0;
	wire w_dff_A_W5URmVKc2_0;
	wire w_dff_A_aHOFvn8s4_0;
	wire w_dff_A_klRREsbW1_0;
	wire w_dff_A_o7ic6DTW2_0;
	wire w_dff_A_nvAytiyE1_0;
	wire w_dff_A_PHVMzs0Y3_0;
	wire w_dff_A_raQoTS7M3_0;
	wire w_dff_A_OGxE8JX77_0;
	wire w_dff_A_px31xyQS5_0;
	wire w_dff_A_YUgeAv468_0;
	wire w_dff_A_9QEbeaqf5_0;
	wire w_dff_A_zmXWwGoB8_0;
	wire w_dff_A_DJQN6eg72_0;
	wire w_dff_A_nbrH8tmC0_0;
	wire w_dff_A_ovVpdRfI5_0;
	wire w_dff_A_x2UNeOZM1_0;
	wire w_dff_A_lsJ0nEbo7_0;
	wire w_dff_A_pWtxQTJB2_0;
	wire w_dff_A_M473xJ4v7_0;
	wire w_dff_A_FZFd6F855_0;
	wire w_dff_A_udFgmkA59_0;
	wire w_dff_A_fWc4L2vd3_0;
	wire w_dff_A_jnF6Pakn5_0;
	wire w_dff_A_4FhdXpys8_0;
	wire w_dff_A_aX74ePjH3_0;
	wire w_dff_A_Zaf6Ilxr6_0;
	wire w_dff_A_4ptKqsnL1_0;
	wire w_dff_A_S6FwpfXP2_0;
	wire w_dff_B_pflvUWRu2_1;
	wire w_dff_A_BkMzg41H7_0;
	wire w_dff_A_874bzRIp1_0;
	wire w_dff_A_Pi9kDOzQ8_0;
	wire w_dff_A_FjrK4XQF9_0;
	wire w_dff_A_BD4R69X74_0;
	wire w_dff_A_5H5Mfybo4_0;
	wire w_dff_A_6Al7Lf9H1_0;
	wire w_dff_A_h45etCDT9_0;
	wire w_dff_A_yarTC1jo8_0;
	wire w_dff_A_pnXH4Ybz6_0;
	wire w_dff_A_xuWaMKId7_0;
	wire w_dff_A_TLnCxtf08_0;
	wire w_dff_A_hJupKqFd2_0;
	wire w_dff_A_wqnVDYpm4_0;
	wire w_dff_A_H6lXtifl8_0;
	wire w_dff_A_0o9ep4IJ2_0;
	wire w_dff_A_ngNl0rDB5_0;
	wire w_dff_A_MF5G3qvD7_0;
	wire w_dff_A_u91J4fVZ0_0;
	wire w_dff_A_SFzKZ4Af7_0;
	wire w_dff_A_omaWsmV62_0;
	wire w_dff_A_yzbQNLsX6_0;
	wire w_dff_A_dz7BvYCT4_0;
	wire w_dff_A_2RHVdoY11_0;
	wire w_dff_A_Gbvra4eQ6_0;
	wire w_dff_A_1ACIXW4Q5_0;
	wire w_dff_A_09Sa6nK39_0;
	wire w_dff_A_hUZRuwci2_0;
	wire w_dff_A_lzu8y0t96_0;
	wire w_dff_A_TZN8eWhu9_0;
	wire w_dff_A_RE0eJ62Y9_0;
	wire w_dff_A_zSfyDgec7_0;
	wire w_dff_A_ukLUEFGu4_0;
	wire w_dff_A_tq7qiosp1_0;
	wire w_dff_A_0YxJ5nxx6_0;
	wire w_dff_B_pjmkXbrx0_1;
	wire w_dff_A_hPP2WvLp3_0;
	wire w_dff_A_ZcpJgxuk2_0;
	wire w_dff_A_H7YS8Hq79_0;
	wire w_dff_A_RdgYIqt98_0;
	wire w_dff_A_UnLDxG4N4_0;
	wire w_dff_A_cwA9ZUkH5_0;
	wire w_dff_A_pVk3wPz71_0;
	wire w_dff_A_YgW0X4hY4_0;
	wire w_dff_A_uPymbpzY0_0;
	wire w_dff_A_nxYo3GfB3_0;
	wire w_dff_A_hys25FMj2_0;
	wire w_dff_A_xiTh05Q15_0;
	wire w_dff_A_5NdCmXGl7_0;
	wire w_dff_A_q5tHYBIt7_0;
	wire w_dff_A_I30KBgqn4_0;
	wire w_dff_A_eCCRbfEC2_0;
	wire w_dff_A_GzUIL9WD9_0;
	wire w_dff_A_Xhc8ANEq3_0;
	wire w_dff_A_aKybp6xT8_0;
	wire w_dff_A_amGNss0t3_0;
	wire w_dff_A_3NjSbybY7_0;
	wire w_dff_A_8mluqX3F5_0;
	wire w_dff_A_2JlJnlK45_0;
	wire w_dff_A_x2F3LTla3_0;
	wire w_dff_A_XxstEwhI9_0;
	wire w_dff_A_yMGypQkr1_0;
	wire w_dff_A_B9Q8kb3U8_0;
	wire w_dff_A_idSjjSXm6_0;
	wire w_dff_A_khsGPbNH3_0;
	wire w_dff_A_cZKhTl2L2_0;
	wire w_dff_A_fKn3qFcf1_0;
	wire w_dff_A_u6y9dCsG3_0;
	wire w_dff_B_NqzeNCcz1_1;
	wire w_dff_A_4xmEb0ep2_0;
	wire w_dff_A_IEYs6iOb1_0;
	wire w_dff_A_k9fkmrUQ1_0;
	wire w_dff_A_yYqPLQi00_0;
	wire w_dff_A_UTnePFQt5_0;
	wire w_dff_A_r34x6rcn3_0;
	wire w_dff_A_RhVxffoR6_0;
	wire w_dff_A_dUmpYrUh4_0;
	wire w_dff_A_psyDIvGL7_0;
	wire w_dff_A_lbgNL8dD1_0;
	wire w_dff_A_Bp7fFiIQ8_0;
	wire w_dff_A_PZTquga30_0;
	wire w_dff_A_kVWIOkab1_0;
	wire w_dff_A_fNLZtWMb5_0;
	wire w_dff_A_Q1hC4ogO9_0;
	wire w_dff_A_s0ukA6Jz5_0;
	wire w_dff_A_KuEc4sXA8_0;
	wire w_dff_A_qKHTRJsL6_0;
	wire w_dff_A_UuOZMD157_0;
	wire w_dff_A_crLqfn9P2_0;
	wire w_dff_A_nEeZKSXp7_0;
	wire w_dff_A_ehHhY8Ci6_0;
	wire w_dff_A_1HutRfl41_0;
	wire w_dff_A_t7R1ENKv3_0;
	wire w_dff_A_jPX4NgYz5_0;
	wire w_dff_A_PucVo6wk5_0;
	wire w_dff_A_lY6R6JyL6_0;
	wire w_dff_A_qmqeJ4rw5_0;
	wire w_dff_A_fQs3s16e9_0;
	wire w_dff_B_qGdEvmpm9_1;
	wire w_dff_A_vKobrcIW5_0;
	wire w_dff_A_vmQOtDJF2_0;
	wire w_dff_A_3gmszpDI1_0;
	wire w_dff_A_jt63r7Nx0_0;
	wire w_dff_A_RusFWgCS9_0;
	wire w_dff_A_ikiqNDu64_0;
	wire w_dff_A_hu30fkaM2_0;
	wire w_dff_A_CcKmnVpu3_0;
	wire w_dff_A_siJIrCQB3_0;
	wire w_dff_A_bnMv18Mk7_0;
	wire w_dff_A_anY4MMgQ7_0;
	wire w_dff_A_4wqqoZNz3_0;
	wire w_dff_A_y5FNnRqY6_0;
	wire w_dff_A_i3q8QPFv4_0;
	wire w_dff_A_yjZQIPzv6_0;
	wire w_dff_A_yp7xCUph3_0;
	wire w_dff_A_zAEsPfJ83_0;
	wire w_dff_A_0RY2ywOg5_0;
	wire w_dff_A_Nqp6xeQH0_0;
	wire w_dff_A_fGGLGsqf4_0;
	wire w_dff_A_nYBXpLvA8_0;
	wire w_dff_A_XW5iWM399_0;
	wire w_dff_A_ULGsBPMI9_0;
	wire w_dff_A_MUa2RZ6j8_0;
	wire w_dff_A_tCowXLRu0_0;
	wire w_dff_A_pU4uyEYh8_0;
	wire w_dff_B_jnPhVbWa4_1;
	wire w_dff_A_c9CUVApT3_0;
	wire w_dff_A_Wd4YsLYq3_0;
	wire w_dff_A_I1gyvQs00_0;
	wire w_dff_A_9YYawam92_0;
	wire w_dff_A_MK6i0Hfr3_0;
	wire w_dff_A_c5ArgNKk2_0;
	wire w_dff_A_YXKh3GUv6_0;
	wire w_dff_A_GG1B0wA87_0;
	wire w_dff_A_DdIj7Hqy1_0;
	wire w_dff_A_Pf1ejpuG9_0;
	wire w_dff_A_GibrthsK2_0;
	wire w_dff_A_47anQ0hc8_0;
	wire w_dff_A_x5WIydQU3_0;
	wire w_dff_A_VgvozxVI6_0;
	wire w_dff_A_qaKzyUob6_0;
	wire w_dff_A_ezOmsEHF8_0;
	wire w_dff_A_ZMOCpJGr0_0;
	wire w_dff_A_Ous7uqdB9_0;
	wire w_dff_A_yozDzvJL8_0;
	wire w_dff_A_vZC30y7j0_0;
	wire w_dff_A_QjGsalrL6_0;
	wire w_dff_A_RqtKQE7V3_0;
	wire w_dff_A_CDV3PFhs0_0;
	wire w_dff_B_s7OczH1C1_1;
	wire w_dff_A_EWcRos1r1_0;
	wire w_dff_A_Qppmjvlc5_0;
	wire w_dff_A_JTkS87u49_0;
	wire w_dff_A_EgBelY8x3_0;
	wire w_dff_A_ooDQBnt85_0;
	wire w_dff_A_OVkuv4Hf3_0;
	wire w_dff_A_WgdkfFkG3_0;
	wire w_dff_A_rYNFFamI9_0;
	wire w_dff_A_IhCktVbw2_0;
	wire w_dff_A_HTjec5nu6_0;
	wire w_dff_A_LCKHzrEY8_0;
	wire w_dff_A_gPa4Tju61_0;
	wire w_dff_A_DGqGTPOR1_0;
	wire w_dff_A_5V4KukZA8_0;
	wire w_dff_A_vlyGCtiS8_0;
	wire w_dff_A_x7l1k7f49_0;
	wire w_dff_A_3FW2y6830_0;
	wire w_dff_A_7bKFNt5E9_0;
	wire w_dff_A_Ob6ywave7_0;
	wire w_dff_A_WKLMPdYf9_0;
	wire w_dff_B_6xod8Z1X3_1;
	wire w_dff_A_gWXZKh5j0_0;
	wire w_dff_A_4ygwGMfm1_0;
	wire w_dff_A_jKOssVq52_0;
	wire w_dff_A_nXeguX2d5_0;
	wire w_dff_A_47b6gRoU0_0;
	wire w_dff_A_dlWJZGOb0_0;
	wire w_dff_A_Qp4jWFqG9_0;
	wire w_dff_A_34ICDyzh5_0;
	wire w_dff_A_VV5haM3s3_0;
	wire w_dff_A_Ab4P2APt8_0;
	wire w_dff_A_A7qlV5fJ8_0;
	wire w_dff_A_9NQH1Hck0_0;
	wire w_dff_A_Z3uEeiyT6_0;
	wire w_dff_A_mWdRIALO2_0;
	wire w_dff_A_r95HNJHx4_0;
	wire w_dff_A_f6h1wyU90_0;
	wire w_dff_A_Mw4tBpp83_0;
	wire w_dff_B_v4dJJxTg5_1;
	wire w_dff_A_v9ROwN3l1_0;
	wire w_dff_A_mlbnknNB5_0;
	wire w_dff_A_KHpYXwe94_0;
	wire w_dff_A_lc5GsPDE2_0;
	wire w_dff_A_Ax4HIcq91_0;
	wire w_dff_A_djrQjCzI8_0;
	wire w_dff_A_sJ0SeAbj8_0;
	wire w_dff_A_fQALokLp6_0;
	wire w_dff_A_FF16szPC6_0;
	wire w_dff_A_lbjjzWXB8_0;
	wire w_dff_A_otSeZaLP2_0;
	wire w_dff_A_M4KJUkD10_0;
	wire w_dff_A_NRNMucvL8_0;
	wire w_dff_A_w4z6xIvG0_0;
	wire w_dff_B_P5uHvnYR7_1;
	wire w_dff_A_9H74tyFG1_0;
	wire w_dff_A_vMII5KeB2_0;
	wire w_dff_A_JYeQomv10_0;
	wire w_dff_A_kDfU426D9_0;
	wire w_dff_A_onCYGSyy7_0;
	wire w_dff_A_Tr4czpk28_0;
	wire w_dff_A_HXgL8b5L6_0;
	wire w_dff_A_8u86IOad2_0;
	wire w_dff_A_Oi0d4Ul72_0;
	wire w_dff_A_cKR98tgH2_0;
	wire w_dff_A_kFA4SIdY6_0;
	wire w_dff_B_rLkhshyZ4_1;
	wire w_dff_A_w7t3SQ1H9_0;
	wire w_dff_A_j4jcI51m9_0;
	wire w_dff_A_ATAEXh6Y4_0;
	wire w_dff_A_iQIRmVPF3_0;
	wire w_dff_A_MDiL3YUI2_0;
	wire w_dff_A_xgwL2N8j9_0;
	wire w_dff_A_7Mzcdqd21_0;
	wire w_dff_A_HGFBKBQc8_0;
	wire w_dff_B_aDyFGiMl4_1;
	wire w_dff_A_XbFi8tcJ8_0;
	wire w_dff_A_KOTv3AcU0_0;
	wire w_dff_A_wwS2XDmP7_0;
	wire w_dff_A_LooSY29h1_0;
	wire w_dff_B_pauhNMKf4_0;
	wire w_dff_A_4Cr04xW87_0;
	wire w_dff_A_oD3ElxP60_0;
	wire w_dff_B_Bbcq3lRP1_2;
	wire w_dff_B_LgYTS43i4_2;
	wire w_dff_B_Oudw9POv2_2;
	wire w_dff_B_eJ0cDlGA4_2;
	wire w_dff_B_C2Pngclt1_2;
	wire w_dff_B_g2nK8mFz5_2;
	wire w_dff_B_xvgwsWYY3_2;
	wire w_dff_B_9BlIUzYT6_2;
	wire w_dff_B_UzWkzLDJ2_2;
	wire w_dff_B_Zden3azW1_2;
	wire w_dff_B_Xcp1Kz0p2_2;
	wire w_dff_B_ade9fVKS7_2;
	wire w_dff_B_BmnmFuhG8_2;
	wire w_dff_B_ngd7ZRpQ2_2;
	wire w_dff_B_ZmYg8W020_2;
	wire w_dff_B_BUex7L529_2;
	wire w_dff_B_JawP3uC30_2;
	wire w_dff_B_fH8IqvuM7_2;
	wire w_dff_B_WbbQwUMv3_2;
	wire w_dff_B_p5Bv42Nr6_2;
	wire w_dff_B_ycjaokEY0_2;
	wire w_dff_B_AOo7R1Bh7_2;
	wire w_dff_B_gQDPjm2r9_2;
	wire w_dff_B_HzEGZ5AM3_2;
	wire w_dff_B_YSkcUHKH6_2;
	wire w_dff_B_Z7Ma2Q4C4_2;
	wire w_dff_B_vKFnm0kb2_2;
	wire w_dff_B_jNXF6eTv5_2;
	wire w_dff_B_8ojo4nA36_2;
	wire w_dff_B_HbRJAvVw6_2;
	wire w_dff_B_mm3RPkfR6_2;
	wire w_dff_B_pEPvXgTw1_2;
	wire w_dff_B_gC6cCtvb2_2;
	wire w_dff_B_gEA4SDhR6_2;
	wire w_dff_B_iwPS3qqy2_2;
	wire w_dff_B_qPYFRTc24_2;
	wire w_dff_B_gPyMBkQI4_2;
	wire w_dff_B_c3u4iLAr3_2;
	wire w_dff_B_y6dDS9im9_2;
	wire w_dff_B_ZQB8hzz96_2;
	wire w_dff_B_IeLlsolF9_2;
	wire w_dff_B_qV3ZJGDP6_2;
	wire w_dff_B_wn7iVQvM7_2;
	wire w_dff_B_GkYwjBE79_2;
	wire w_dff_A_pgxmyIZO4_0;
	wire w_dff_B_AwXEy4nt7_1;
	wire w_dff_B_8BpXqk955_2;
	wire w_dff_B_5kaMtNpR5_2;
	wire w_dff_B_MsUm0t9m3_2;
	wire w_dff_B_30dGTRy01_2;
	wire w_dff_B_Gfa33qcr6_2;
	wire w_dff_B_7zo4x7nJ8_2;
	wire w_dff_B_QHDRsdIK2_2;
	wire w_dff_B_GV2dQea63_2;
	wire w_dff_B_zK2pMWOU6_2;
	wire w_dff_B_7jGyAMrY9_2;
	wire w_dff_B_0OKoFKiV5_2;
	wire w_dff_B_0B0WJbEs4_2;
	wire w_dff_B_x7uCCsQu0_2;
	wire w_dff_B_mGWQHK8e9_2;
	wire w_dff_B_CimIGaKH5_2;
	wire w_dff_B_bA1fIJzC5_2;
	wire w_dff_B_Kl2EFHPx5_2;
	wire w_dff_B_DPDyPAtr7_2;
	wire w_dff_B_V0FEB6WK2_2;
	wire w_dff_B_CntoOaCF0_2;
	wire w_dff_B_eB6f7E5r4_2;
	wire w_dff_B_LY4MKY2l8_2;
	wire w_dff_B_TVejp6KR9_2;
	wire w_dff_B_bE8Emp6j3_2;
	wire w_dff_B_KKlKOssP8_2;
	wire w_dff_B_b3jzkhOZ3_2;
	wire w_dff_B_nRt4USLP4_2;
	wire w_dff_B_Q7O5YwYF0_2;
	wire w_dff_B_ERabeJf06_2;
	wire w_dff_B_Gq7D5bBI7_2;
	wire w_dff_B_voqTkvNb5_2;
	wire w_dff_B_jRDmwexT9_2;
	wire w_dff_B_TeHlzT608_2;
	wire w_dff_B_tlyYCVOv9_2;
	wire w_dff_B_OofZ6gfh7_2;
	wire w_dff_B_B9TVCtWm2_2;
	wire w_dff_B_qTjXRTk78_2;
	wire w_dff_B_51vgnAj54_2;
	wire w_dff_B_RB89K6Gk5_2;
	wire w_dff_B_sNYQT0OB0_2;
	wire w_dff_A_Ig2IiMIV7_1;
	wire w_dff_A_S9PIOujp5_0;
	wire w_dff_A_xnh2ICtZ4_0;
	wire w_dff_A_O9TlwrpB7_0;
	wire w_dff_A_6awEeOUm7_0;
	wire w_dff_A_c7uzayFU0_0;
	wire w_dff_A_AcJlvA2K6_0;
	wire w_dff_A_tVpkZpNI1_0;
	wire w_dff_A_ltnxb5vx3_0;
	wire w_dff_A_2qeuCHrk9_0;
	wire w_dff_A_LxDgNnRa1_0;
	wire w_dff_A_HUxE6ItK3_0;
	wire w_dff_A_RUPJUt0V3_0;
	wire w_dff_A_XwqwnjGT3_0;
	wire w_dff_A_wyX1GCcq5_0;
	wire w_dff_A_mWlAdXdo8_0;
	wire w_dff_A_QWUW1Qou1_0;
	wire w_dff_A_IRijIAHQ0_0;
	wire w_dff_A_4acfb7WY5_0;
	wire w_dff_A_VjGgXz3y1_0;
	wire w_dff_A_5wSlEO0x5_0;
	wire w_dff_A_YloFWHmu7_0;
	wire w_dff_A_HgqSJjSE2_0;
	wire w_dff_A_M17ZIlp44_0;
	wire w_dff_A_wi1I0ai18_0;
	wire w_dff_A_qN1KMaIG3_0;
	wire w_dff_A_JKcFQTYX3_0;
	wire w_dff_A_7WdnC1v71_0;
	wire w_dff_A_IndqoNG13_0;
	wire w_dff_A_fC8iFi6T1_0;
	wire w_dff_A_WRQh3zLS5_0;
	wire w_dff_A_IsSXWxk38_0;
	wire w_dff_A_mWoYxURw9_0;
	wire w_dff_A_Muh60JkR9_0;
	wire w_dff_A_G9VXaPrw3_0;
	wire w_dff_A_xVDWveXm4_0;
	wire w_dff_A_CWzR1lEv6_0;
	wire w_dff_A_0TE8lFqx1_0;
	wire w_dff_A_l6lgNt926_1;
	wire w_dff_A_fTqCUQNZ9_2;
	wire w_dff_B_tjlHIzTL2_1;
	wire w_dff_B_hVtGoqtw7_2;
	wire w_dff_B_BGyenYGj6_2;
	wire w_dff_B_w4Lkn5jg6_2;
	wire w_dff_B_j9RLxeHL3_2;
	wire w_dff_B_HTSAbvKw5_2;
	wire w_dff_B_yFLPmvyQ9_2;
	wire w_dff_B_yuqETpIQ5_2;
	wire w_dff_B_C1xYgUPO6_2;
	wire w_dff_B_YnJXQg3j4_2;
	wire w_dff_B_VIqON7Z05_2;
	wire w_dff_B_72fmwJ2L9_2;
	wire w_dff_B_uNoHPmd20_2;
	wire w_dff_B_kZB5kuyT4_2;
	wire w_dff_B_uoAmyg234_2;
	wire w_dff_B_StdMDfwz9_2;
	wire w_dff_B_owRQFHUV4_2;
	wire w_dff_B_ubmCFz354_2;
	wire w_dff_B_ltVpqtfV1_2;
	wire w_dff_B_HojszjWL1_2;
	wire w_dff_B_VPB3AA0m8_2;
	wire w_dff_B_0AF2VxD82_2;
	wire w_dff_B_OI6G4csf5_2;
	wire w_dff_B_qP1jrZuS9_2;
	wire w_dff_B_jT2368OV1_2;
	wire w_dff_B_SvrTqzrS7_2;
	wire w_dff_B_uyGJBh3X2_2;
	wire w_dff_B_mtlYpPd84_2;
	wire w_dff_B_AY7Kt3ua7_2;
	wire w_dff_B_YGGkpzm89_2;
	wire w_dff_B_ZAwMDljP6_2;
	wire w_dff_B_IixtpD9V8_2;
	wire w_dff_B_ah4ViFEx7_2;
	wire w_dff_B_iI69Sy724_2;
	wire w_dff_B_jkAymBlt3_2;
	wire w_dff_B_qWDKSY1J5_1;
	wire w_dff_B_biP9Zti95_2;
	wire w_dff_B_8C4FMtFD3_2;
	wire w_dff_B_VYqPFXeF0_2;
	wire w_dff_B_4paEbKGf4_2;
	wire w_dff_B_nYpRnQdA2_2;
	wire w_dff_B_z9Of2kY57_2;
	wire w_dff_B_LdOO0mpp1_2;
	wire w_dff_B_GppeaWwv3_2;
	wire w_dff_B_3qosq3h65_2;
	wire w_dff_B_nGJuWHB58_2;
	wire w_dff_B_vcSlr4s27_2;
	wire w_dff_B_spNi7WVu3_2;
	wire w_dff_B_BvjI52qV9_2;
	wire w_dff_B_5gXu3jfi7_2;
	wire w_dff_B_MWhU6ZVS7_2;
	wire w_dff_B_YLTR9ZYY9_2;
	wire w_dff_B_GeVXzpm79_2;
	wire w_dff_B_fsAKEm1y8_2;
	wire w_dff_B_bHftqYYi0_2;
	wire w_dff_B_7vAgEoTV1_2;
	wire w_dff_B_ZWw8runF6_2;
	wire w_dff_B_Lmw2EkNw7_2;
	wire w_dff_B_lI7YnOhd9_2;
	wire w_dff_B_UzdgR5uo4_2;
	wire w_dff_B_7UhaOJkU0_2;
	wire w_dff_B_0WdFHa4f7_2;
	wire w_dff_B_ikGBUAgq8_2;
	wire w_dff_B_YA36SIE08_2;
	wire w_dff_B_k5xok1rj4_2;
	wire w_dff_B_l80K2F2M7_2;
	wire w_dff_B_mZTqKZKU0_2;
	wire w_dff_B_3fIFSjOP8_1;
	wire w_dff_B_69YsihiC8_2;
	wire w_dff_B_WkjculoG2_2;
	wire w_dff_B_9PjHFIgW2_2;
	wire w_dff_B_9QVii5Ix8_2;
	wire w_dff_B_2ZV56b0g1_2;
	wire w_dff_B_rMiGF1Qi9_2;
	wire w_dff_B_XfJFoGPi9_2;
	wire w_dff_B_cizMnaxg3_2;
	wire w_dff_B_BDw5m5AH8_2;
	wire w_dff_B_Y12UcpN05_2;
	wire w_dff_B_eaNrTYmG1_2;
	wire w_dff_B_x9n9wSfl5_2;
	wire w_dff_B_evK23eiy0_2;
	wire w_dff_B_jenYlyly2_2;
	wire w_dff_B_IbvcS0SH2_2;
	wire w_dff_B_9mRY4NJQ3_2;
	wire w_dff_B_cK2bwMb20_2;
	wire w_dff_B_ucru1cW17_2;
	wire w_dff_B_S687hQYd4_2;
	wire w_dff_B_09pPRDxc3_2;
	wire w_dff_B_Io5Mz4PT2_2;
	wire w_dff_B_rU7fOSqf7_2;
	wire w_dff_B_z4azcPV95_2;
	wire w_dff_B_RlRmQd2E9_2;
	wire w_dff_B_eALBBeqr7_2;
	wire w_dff_B_lscsfo6j1_2;
	wire w_dff_B_eR3Wb2sf5_2;
	wire w_dff_B_Q4Xb684L2_2;
	wire w_dff_B_KtEFl8uK2_1;
	wire w_dff_B_YOHpvLlj5_2;
	wire w_dff_B_c1sW522N2_2;
	wire w_dff_B_BXnsZxxL4_2;
	wire w_dff_B_HHnhWQfZ6_2;
	wire w_dff_B_ZvMJZtFk5_2;
	wire w_dff_B_NfSyGMGu5_2;
	wire w_dff_B_NvOE3LZD0_2;
	wire w_dff_B_vD9iUEHj6_2;
	wire w_dff_B_RRaTGuhc5_2;
	wire w_dff_B_VzDQvlwo3_2;
	wire w_dff_B_uquQkKXu1_2;
	wire w_dff_B_FXeKZdie9_2;
	wire w_dff_B_RB7PdyId3_2;
	wire w_dff_B_miIF4meo0_2;
	wire w_dff_B_DsbP680z0_2;
	wire w_dff_B_ZNhsVKBN3_2;
	wire w_dff_B_FMFjZmjJ5_2;
	wire w_dff_B_HkkgOSe64_2;
	wire w_dff_B_w6Ju8LO91_2;
	wire w_dff_B_RCpJbxQj1_2;
	wire w_dff_B_djHnKz494_2;
	wire w_dff_B_VrSQM04q7_2;
	wire w_dff_B_GT6xsgMZ8_2;
	wire w_dff_B_w7W1k9Hk6_2;
	wire w_dff_B_hZo4AJL16_2;
	wire w_dff_B_gOSBDxmP5_1;
	wire w_dff_B_MhdsDXXB8_2;
	wire w_dff_B_fwA2z8ik0_2;
	wire w_dff_B_IdyDmHs90_2;
	wire w_dff_B_H0cgRTLw6_2;
	wire w_dff_B_WxCVjQDi9_2;
	wire w_dff_B_MeEwdt0v6_2;
	wire w_dff_B_DZCKW1Al3_2;
	wire w_dff_B_MOxIcfym4_2;
	wire w_dff_B_ixAZpz546_2;
	wire w_dff_B_JJUzFS988_2;
	wire w_dff_B_ld838vVh5_2;
	wire w_dff_B_sxPuUwLJ7_2;
	wire w_dff_B_2YISQFJi4_2;
	wire w_dff_B_ELL9OwzR6_2;
	wire w_dff_B_0kEpU8ef5_2;
	wire w_dff_B_eQAYCGik0_2;
	wire w_dff_B_CopEqRwn1_2;
	wire w_dff_B_FVzKIRze0_2;
	wire w_dff_B_GlvoadhE4_2;
	wire w_dff_B_fyXt3Iiz2_2;
	wire w_dff_B_ZCDYx5Hp6_2;
	wire w_dff_B_VAUq4dSN9_2;
	wire w_dff_B_elABO3cg9_1;
	wire w_dff_B_hwLaWcnf6_2;
	wire w_dff_B_qEjWbzPN8_2;
	wire w_dff_B_2RNSW0dd4_2;
	wire w_dff_B_CFnm898Y0_2;
	wire w_dff_B_k77rVTrd2_2;
	wire w_dff_B_DA6fB0uE3_2;
	wire w_dff_B_4H64QbTv2_2;
	wire w_dff_B_5oAa4zcv6_2;
	wire w_dff_B_APU4c4Aq1_2;
	wire w_dff_B_3GT30ZCg7_2;
	wire w_dff_B_bELeBRCW3_2;
	wire w_dff_B_iE7qehjO7_2;
	wire w_dff_B_51i5gpmL9_2;
	wire w_dff_B_mF8Ej48u5_2;
	wire w_dff_B_HVnQXriL1_2;
	wire w_dff_B_28SrPSr41_2;
	wire w_dff_B_ioy2gMR02_2;
	wire w_dff_B_y67DCB5M1_2;
	wire w_dff_B_QEgq628n1_2;
	wire w_dff_B_01uMWL296_1;
	wire w_dff_B_a1T8jJQb3_2;
	wire w_dff_B_ZK8ndZg76_2;
	wire w_dff_B_kJ3DrL9d0_2;
	wire w_dff_B_rEJg5UC37_2;
	wire w_dff_B_AX0bdwf96_2;
	wire w_dff_B_garsuYDJ8_2;
	wire w_dff_B_7d4TyI5H9_2;
	wire w_dff_B_jYlutrkL3_2;
	wire w_dff_B_w3BqEHiK9_2;
	wire w_dff_B_21D6IUUz6_2;
	wire w_dff_B_SnbnlTq58_2;
	wire w_dff_B_dadRfedO6_2;
	wire w_dff_B_BI0V2RgV0_2;
	wire w_dff_B_fGx0M5r74_2;
	wire w_dff_B_4xzSKqT53_2;
	wire w_dff_B_O5DfBWIa0_2;
	wire w_dff_B_4NcILaiO4_1;
	wire w_dff_B_hWBQMU3w6_2;
	wire w_dff_B_I9RT2yjy3_2;
	wire w_dff_B_8mHZPK9a1_2;
	wire w_dff_B_DAN92S8r7_2;
	wire w_dff_B_V0YjDXYs4_2;
	wire w_dff_B_v98BEKwL6_2;
	wire w_dff_B_gYvV5HxF7_2;
	wire w_dff_B_6jVmbgM30_2;
	wire w_dff_B_5VJc7xDt7_2;
	wire w_dff_B_uzJH1FrF2_2;
	wire w_dff_B_cX0SYfVX4_2;
	wire w_dff_B_7od6T22O2_2;
	wire w_dff_B_gHhvR5im2_2;
	wire w_dff_B_awINEBjq5_1;
	wire w_dff_B_lJxH3CAW7_2;
	wire w_dff_B_R7uqlSYm0_2;
	wire w_dff_B_uC870PGZ9_2;
	wire w_dff_B_aoGuBHfk3_2;
	wire w_dff_B_hhSrjFqh1_2;
	wire w_dff_B_vZJGX8Ys3_2;
	wire w_dff_B_Qv5EgmYz6_2;
	wire w_dff_B_YsN32FRz8_2;
	wire w_dff_B_zjj0zFqA2_2;
	wire w_dff_B_OTekOYmC2_2;
	wire w_dff_B_Duh6237q9_1;
	wire w_dff_B_IfhUVmGC1_2;
	wire w_dff_B_LczE3Lmg0_2;
	wire w_dff_B_liEYByHO6_2;
	wire w_dff_B_QNxxOwXm4_2;
	wire w_dff_B_KefqDJAc4_2;
	wire w_dff_B_7T33LGME5_2;
	wire w_dff_B_My0VlJMI7_2;
	wire w_dff_B_TbGNR3Fo0_2;
	wire w_dff_B_YHLHf0045_2;
	wire w_dff_B_WUu4GHNc7_2;
	wire w_dff_B_ULWUSYyN0_0;
	wire w_dff_B_T7uFMeCt1_0;
	wire w_dff_A_0aHcLnK74_1;
	wire w_dff_A_vXmbbNVz1_1;
	wire w_dff_B_5cYZM5lH4_1;
	wire w_dff_B_dNEC8t638_1;
	wire w_dff_B_5FxeB74n6_2;
	wire w_dff_B_8eU6m3TK0_2;
	wire w_dff_B_aY7vb9RH3_2;
	wire w_dff_B_j3Y2cl8M0_2;
	wire w_dff_B_uQAWDbP54_2;
	wire w_dff_B_uLO0FDRf1_2;
	wire w_dff_B_nYY0mzsr5_2;
	wire w_dff_B_ojeGawvS1_2;
	wire w_dff_B_sDHPtxl30_2;
	wire w_dff_B_VcHc3vAx3_2;
	wire w_dff_B_zutsqV7m8_2;
	wire w_dff_B_wRJE5q9U3_2;
	wire w_dff_B_Oe9lUesJ4_2;
	wire w_dff_B_qkrpvotO8_2;
	wire w_dff_B_YM7dK0EM3_2;
	wire w_dff_B_X6WEpmbD5_2;
	wire w_dff_B_CQJ9m3qm2_2;
	wire w_dff_B_1PGOmBdS1_2;
	wire w_dff_B_HCSCg9zD9_2;
	wire w_dff_B_PqEYFeOp0_2;
	wire w_dff_B_DDibQBoL1_2;
	wire w_dff_B_2N9rZFQa5_2;
	wire w_dff_B_cZzXQ1nW6_2;
	wire w_dff_B_DrDDijPw6_2;
	wire w_dff_B_XVwnxa3E9_2;
	wire w_dff_B_ECwYTLId8_2;
	wire w_dff_B_NAQ7WFtU0_2;
	wire w_dff_B_kMFTsYbB8_2;
	wire w_dff_B_R1yWHHhj0_2;
	wire w_dff_B_aP5expyP3_2;
	wire w_dff_B_qWS2rGsJ2_2;
	wire w_dff_B_9dlO2y3O1_2;
	wire w_dff_B_lL2U8Set6_2;
	wire w_dff_B_RD5pl4S27_2;
	wire w_dff_B_vSTGKNJT7_2;
	wire w_dff_B_JHPmVqIP0_2;
	wire w_dff_B_D7ei4GmZ8_2;
	wire w_dff_B_gk4THjet9_2;
	wire w_dff_B_Aizn5nb75_2;
	wire w_dff_B_O4AsLtNS0_2;
	wire w_dff_B_7R6rw7q18_2;
	wire w_dff_B_lmnA66fG7_2;
	wire w_dff_B_IJ0Z0k6e4_2;
	wire w_dff_B_8V8XETCW6_2;
	wire w_dff_B_N6CcgjhU8_2;
	wire w_dff_B_g5qSM25j2_2;
	wire w_dff_B_dTWjquK89_1;
	wire w_dff_B_LaUlfFI53_2;
	wire w_dff_B_gMn8pWZ36_2;
	wire w_dff_B_xFQ39yQZ5_2;
	wire w_dff_B_uNDwr3PX4_2;
	wire w_dff_B_xpZFzXIR8_2;
	wire w_dff_B_C8qaNjaP0_2;
	wire w_dff_B_NLYtQFB73_2;
	wire w_dff_B_NE8sBkr32_2;
	wire w_dff_B_GclNvpcU8_2;
	wire w_dff_B_LRHHXjOn1_2;
	wire w_dff_B_rj4sTifu3_2;
	wire w_dff_B_qHMjqg013_2;
	wire w_dff_B_ghLWkcMT2_2;
	wire w_dff_B_KbVaCQiV0_2;
	wire w_dff_B_y5ZHfqiq0_2;
	wire w_dff_B_mXz8Kk2I4_2;
	wire w_dff_B_k5GTW3aM6_2;
	wire w_dff_B_R3VdjnQB9_2;
	wire w_dff_B_F5OGTpki4_2;
	wire w_dff_B_JjP8fJdZ6_2;
	wire w_dff_B_xH3nT4zI4_2;
	wire w_dff_B_I777N9s45_2;
	wire w_dff_B_OnC1kYJD0_2;
	wire w_dff_B_TQlTeIfE5_2;
	wire w_dff_B_IC9zf8wU6_2;
	wire w_dff_B_kotpLJaf9_2;
	wire w_dff_B_lC6K6ift0_2;
	wire w_dff_B_ZYwrdI9z7_2;
	wire w_dff_B_akkOtuSs1_2;
	wire w_dff_B_CJVmzvky6_2;
	wire w_dff_B_fvc3LnZ15_2;
	wire w_dff_B_GRWKdhPT1_2;
	wire w_dff_B_uiYizq8T8_2;
	wire w_dff_B_PxS9NFLH7_2;
	wire w_dff_B_jfCAjWSx2_2;
	wire w_dff_B_STRwvEif1_2;
	wire w_dff_B_6tlaWTFm4_2;
	wire w_dff_B_nB4hcta01_2;
	wire w_dff_B_Gd5v9ywR2_2;
	wire w_dff_B_gPTWyeiH9_2;
	wire w_dff_B_IcKyzXsc3_2;
	wire w_dff_B_LOO3qfnl6_2;
	wire w_dff_B_jSsFNk300_1;
	wire w_dff_B_0XkwwTlN3_2;
	wire w_dff_B_t0ZJEpMk9_2;
	wire w_dff_B_BaaxaJfV9_2;
	wire w_dff_B_1ZXBBSUE7_2;
	wire w_dff_B_DkTebevs3_2;
	wire w_dff_B_2snPNeIM4_2;
	wire w_dff_B_PQ6QK7BE4_2;
	wire w_dff_B_AaPCN2NS7_2;
	wire w_dff_B_ZpQbhU5f9_2;
	wire w_dff_B_XeU8s8Dm4_2;
	wire w_dff_B_NX8IPIdd2_2;
	wire w_dff_B_tkQr5MJK0_2;
	wire w_dff_B_50oh49lC2_2;
	wire w_dff_B_FTUJpMRK9_2;
	wire w_dff_B_GI3tVzFC1_2;
	wire w_dff_B_jigLqi2P8_2;
	wire w_dff_B_AjNQBBmb3_2;
	wire w_dff_B_2nesTlPu1_2;
	wire w_dff_B_zUy7i4RU1_2;
	wire w_dff_B_N0tbAMdL5_2;
	wire w_dff_B_8yFXKhmv1_2;
	wire w_dff_B_PwQOxcPN8_2;
	wire w_dff_B_1PR57Ky75_2;
	wire w_dff_B_DqTMZJTI9_2;
	wire w_dff_B_RwA7FrXB8_2;
	wire w_dff_B_ptrrO5bo4_2;
	wire w_dff_B_mAn2FqFP0_2;
	wire w_dff_B_uZhgiULn1_2;
	wire w_dff_B_bmx5x4EL3_2;
	wire w_dff_B_MxOZXmWe0_2;
	wire w_dff_B_tVDbwprB8_2;
	wire w_dff_B_zquJMwJE9_2;
	wire w_dff_B_6L2faNIN0_2;
	wire w_dff_B_nxNZdasy7_2;
	wire w_dff_B_iESR9fib1_2;
	wire w_dff_B_xChHUj2Q5_2;
	wire w_dff_B_ETjCxcFW4_2;
	wire w_dff_B_S5HypYcJ0_1;
	wire w_dff_B_BKIzaoqq7_2;
	wire w_dff_B_4efNMmNp7_2;
	wire w_dff_B_MQzKKLNi5_2;
	wire w_dff_B_kdiv25xZ1_2;
	wire w_dff_B_m3CTBBds8_2;
	wire w_dff_B_fwe6veCj2_2;
	wire w_dff_B_lzC79Yp17_2;
	wire w_dff_B_jmQrW7v43_2;
	wire w_dff_B_GStMJizB3_2;
	wire w_dff_B_jmCLi9nt9_2;
	wire w_dff_B_ZzAUrxgU7_2;
	wire w_dff_B_WWkUyhEj8_2;
	wire w_dff_B_a90X4dGt5_2;
	wire w_dff_B_BZAq3Vyx5_2;
	wire w_dff_B_WM7HKaPc4_2;
	wire w_dff_B_xvh14CFd3_2;
	wire w_dff_B_YODdw0mT7_2;
	wire w_dff_B_F9SR7Nmp0_2;
	wire w_dff_B_JcRg1OUE0_2;
	wire w_dff_B_FLaqh6SV7_2;
	wire w_dff_B_C9IZeMFD3_2;
	wire w_dff_B_WbwzmZ8a7_2;
	wire w_dff_B_B897gTyX3_2;
	wire w_dff_B_ZHXFM0Dt3_2;
	wire w_dff_B_cvNxBoHs4_2;
	wire w_dff_B_B7PPjqe50_2;
	wire w_dff_B_sSi7FJ9F2_2;
	wire w_dff_B_UHvERiTK3_2;
	wire w_dff_B_cC5oSMNd5_2;
	wire w_dff_B_KiCn9g8H1_2;
	wire w_dff_B_oPfQI8687_2;
	wire w_dff_B_Z7om9Y2Q4_2;
	wire w_dff_B_4qzbGwQl1_2;
	wire w_dff_B_UXHgDEAd7_2;
	wire w_dff_B_9fVbZpba6_1;
	wire w_dff_B_YEeYVfOJ1_2;
	wire w_dff_B_9njIobPw1_2;
	wire w_dff_B_4LVZACzC4_2;
	wire w_dff_B_5f5BNmE82_2;
	wire w_dff_B_sK8pOXa97_2;
	wire w_dff_B_ZiIp4TxA9_2;
	wire w_dff_B_6R4gMsf13_2;
	wire w_dff_B_a4fZc1ku5_2;
	wire w_dff_B_dUZ6XPSa6_2;
	wire w_dff_B_uCWOAT1R3_2;
	wire w_dff_B_69UFl0bE5_2;
	wire w_dff_B_Ojd71V7z6_2;
	wire w_dff_B_PJf9AxCq0_2;
	wire w_dff_B_QAdZL6ED1_2;
	wire w_dff_B_YI0NXY1Q5_2;
	wire w_dff_B_IehDabsF5_2;
	wire w_dff_B_lrvEgepr2_2;
	wire w_dff_B_lw8emsln6_2;
	wire w_dff_B_G7iQ1yfU2_2;
	wire w_dff_B_DUhNoIQU2_2;
	wire w_dff_B_G4K64gZg7_2;
	wire w_dff_B_PJs1L76p1_2;
	wire w_dff_B_ubGDez2D1_2;
	wire w_dff_B_hCeJSWaT6_2;
	wire w_dff_B_KUivg05M3_2;
	wire w_dff_B_g243iE7M3_2;
	wire w_dff_B_QJ2js2vY6_2;
	wire w_dff_B_ndrO8KCb4_2;
	wire w_dff_B_G9acgQ5R7_2;
	wire w_dff_B_slip2qC92_2;
	wire w_dff_B_AOXHx3Iw7_2;
	wire w_dff_B_K4OtTcjG8_1;
	wire w_dff_B_bTOkVMSv7_2;
	wire w_dff_B_wohXghU12_2;
	wire w_dff_B_JSNKy6jv4_2;
	wire w_dff_B_RTP7oSkr6_2;
	wire w_dff_B_Fvk8zEjL4_2;
	wire w_dff_B_lxmqH57C9_2;
	wire w_dff_B_RpME737s0_2;
	wire w_dff_B_L90nQbkT0_2;
	wire w_dff_B_hLXuRUF25_2;
	wire w_dff_B_NzuY3Hib3_2;
	wire w_dff_B_74JS0qwJ7_2;
	wire w_dff_B_s5zUVmvx7_2;
	wire w_dff_B_VXhF3oOD5_2;
	wire w_dff_B_MRDj5VZy9_2;
	wire w_dff_B_bUejtSQi4_2;
	wire w_dff_B_8KkOINzm9_2;
	wire w_dff_B_rxAcwCsf7_2;
	wire w_dff_B_Ow7OnWlN3_2;
	wire w_dff_B_A9AL2n199_2;
	wire w_dff_B_Zlob5Hhh8_2;
	wire w_dff_B_yHRWIc8f1_2;
	wire w_dff_B_hRDE12xl0_2;
	wire w_dff_B_e65a5p1x4_2;
	wire w_dff_B_Sm99qv2Q2_2;
	wire w_dff_B_qz9OmIKW8_2;
	wire w_dff_B_sVK3HWJo8_2;
	wire w_dff_B_XIPQYJju6_2;
	wire w_dff_B_9bFez3Sf8_2;
	wire w_dff_B_TNkzBPEQ1_1;
	wire w_dff_B_bBhkbszQ7_2;
	wire w_dff_B_f51oMVeo7_2;
	wire w_dff_B_UbNQtSth0_2;
	wire w_dff_B_FUkSvxAy3_2;
	wire w_dff_B_win2S9aE0_2;
	wire w_dff_B_UmyW3qT50_2;
	wire w_dff_B_yCmJTnyJ4_2;
	wire w_dff_B_Jt98ZZU86_2;
	wire w_dff_B_HvsZa83H6_2;
	wire w_dff_B_zTBHjKWh3_2;
	wire w_dff_B_t5yXvKYO9_2;
	wire w_dff_B_0HdcgnmU9_2;
	wire w_dff_B_sijVBhM94_2;
	wire w_dff_B_1PSw7WPZ5_2;
	wire w_dff_B_G2C2M3vD7_2;
	wire w_dff_B_u4S8Nntb1_2;
	wire w_dff_B_QKMMQkka4_2;
	wire w_dff_B_UQhP4lYA9_2;
	wire w_dff_B_XeM8pS0B5_2;
	wire w_dff_B_6ZeRMQGd4_2;
	wire w_dff_B_8kE73v0Q1_2;
	wire w_dff_B_M9GYRtXm4_2;
	wire w_dff_B_MR0lnAsI3_2;
	wire w_dff_B_jw7L1Y4g3_2;
	wire w_dff_B_fSPB99zU8_2;
	wire w_dff_B_uYM3roB00_1;
	wire w_dff_B_UeJKjEuo2_2;
	wire w_dff_B_M7SsA64h8_2;
	wire w_dff_B_Y3eAVrVf0_2;
	wire w_dff_B_oBiFGf9J4_2;
	wire w_dff_B_CPFMDieT8_2;
	wire w_dff_B_u7iQ1IHo5_2;
	wire w_dff_B_ndnpMWqP0_2;
	wire w_dff_B_vEgA1lS38_2;
	wire w_dff_B_bGn3YH7G4_2;
	wire w_dff_B_ysUq4Td77_2;
	wire w_dff_B_vE2VGbef5_2;
	wire w_dff_B_5Oiv5Ozn4_2;
	wire w_dff_B_mdVkEO9y0_2;
	wire w_dff_B_G6DwSyC76_2;
	wire w_dff_B_BACQ45Mw2_2;
	wire w_dff_B_WVecvOpA4_2;
	wire w_dff_B_qzelPbpo3_2;
	wire w_dff_B_y5X4O3hO9_2;
	wire w_dff_B_AuuQ60UU6_2;
	wire w_dff_B_zkTDCxtL2_2;
	wire w_dff_B_v1qq48ab4_2;
	wire w_dff_B_pYAEP80p8_2;
	wire w_dff_B_mVu63OJQ1_1;
	wire w_dff_B_WEWxMx065_2;
	wire w_dff_B_W1hpzVyU6_2;
	wire w_dff_B_8I3CbCaA9_2;
	wire w_dff_B_AWocKXOg8_2;
	wire w_dff_B_AIDr4X9M9_2;
	wire w_dff_B_NaQCEV502_2;
	wire w_dff_B_e08tTMd56_2;
	wire w_dff_B_1IUHKHOh2_2;
	wire w_dff_B_WTpAsNU15_2;
	wire w_dff_B_57uRIp4D6_2;
	wire w_dff_B_CCYEVUQR3_2;
	wire w_dff_B_fTfVusa95_2;
	wire w_dff_B_K6ainE281_2;
	wire w_dff_B_XaiHOww80_2;
	wire w_dff_B_jTyFb9U55_2;
	wire w_dff_B_2yqMtiOT6_2;
	wire w_dff_B_q5bQKJu14_2;
	wire w_dff_B_80hrZBpf0_2;
	wire w_dff_B_Dr1IrqGm8_2;
	wire w_dff_B_0rCHEG0m8_1;
	wire w_dff_B_Ys6VVuGu3_2;
	wire w_dff_B_0l6c51KU8_2;
	wire w_dff_B_Ty2zuga32_2;
	wire w_dff_B_uer5qByP8_2;
	wire w_dff_B_byXUke3X7_2;
	wire w_dff_B_4EfWPXMY9_2;
	wire w_dff_B_iYbmjNtZ7_2;
	wire w_dff_B_bvlS3ki57_2;
	wire w_dff_B_lezNhEqZ6_2;
	wire w_dff_B_aMd4yMz06_2;
	wire w_dff_B_7ixe8zJH6_2;
	wire w_dff_B_yeDuCsWG2_2;
	wire w_dff_B_QMujZxw62_2;
	wire w_dff_B_Ubl8n52K2_2;
	wire w_dff_B_Nzc0jN0X6_2;
	wire w_dff_B_ytpEQb7Q7_2;
	wire w_dff_B_1rtVAh7u6_1;
	wire w_dff_B_omdEaLWk4_2;
	wire w_dff_B_Fh3oMONb3_2;
	wire w_dff_B_JaeHTARs5_2;
	wire w_dff_B_arJq6s7v9_2;
	wire w_dff_B_RX7mPEjL1_2;
	wire w_dff_B_bZ6rfMWN6_2;
	wire w_dff_B_3wOjXPL01_2;
	wire w_dff_B_t9whI86T7_2;
	wire w_dff_B_Rf099flr7_2;
	wire w_dff_B_kjx61lNX5_2;
	wire w_dff_B_qlspWzHw1_2;
	wire w_dff_B_czwAcrTA5_2;
	wire w_dff_B_Xt3SxkYc6_2;
	wire w_dff_B_P2mKMjuP8_1;
	wire w_dff_B_5TdOO4dZ3_2;
	wire w_dff_B_3FucluDd3_2;
	wire w_dff_B_fgDT3QRk3_2;
	wire w_dff_B_UGXTrXMM9_2;
	wire w_dff_B_pj5D2l2T3_2;
	wire w_dff_B_cVccoivS0_2;
	wire w_dff_B_2evKtaZu4_2;
	wire w_dff_B_W6vCpGoW6_2;
	wire w_dff_B_dQEcMFM43_2;
	wire w_dff_B_VFWvjV9t5_2;
	wire w_dff_B_Zm1aESKy2_1;
	wire w_dff_B_nd94F0Wh0_2;
	wire w_dff_B_GfGcW0iz2_2;
	wire w_dff_B_8umv0ypU0_2;
	wire w_dff_B_NF4kGozM3_2;
	wire w_dff_B_a0SR0zze2_2;
	wire w_dff_B_kLH7gl653_2;
	wire w_dff_B_k8KuEIIu9_2;
	wire w_dff_B_SLOUeJJZ0_2;
	wire w_dff_B_UMrwSk2E5_2;
	wire w_dff_B_ICAcvj6l7_2;
	wire w_dff_B_fGZCObuk2_0;
	wire w_dff_A_CuJghATl4_0;
	wire w_dff_A_2DFVxxTq9_0;
	wire w_dff_A_FEWmkBeV4_0;
	wire w_dff_A_dYnoKGBq0_0;
	wire w_dff_B_SgiYHoB16_1;
	wire w_dff_B_PuYXf8Yd1_2;
	wire w_dff_B_mT5LsNOh5_2;
	wire w_dff_B_obQNMcPx1_2;
	wire w_dff_B_ZOnShia50_2;
	wire w_dff_B_y2vvH2jy3_2;
	wire w_dff_B_rwc7ZNq40_2;
	wire w_dff_B_1qeFN1HJ1_2;
	wire w_dff_B_R9MTpE0L0_2;
	wire w_dff_B_hh7WYfYd2_2;
	wire w_dff_B_scUmfuoJ4_2;
	wire w_dff_B_ebbtcAO11_2;
	wire w_dff_B_NbCVchy23_2;
	wire w_dff_B_56TI56UR8_2;
	wire w_dff_B_ffRliSXe4_2;
	wire w_dff_B_cFjqFrom6_2;
	wire w_dff_B_h3Z3iue59_2;
	wire w_dff_B_9Zyd006o1_2;
	wire w_dff_B_EQsHucWM1_2;
	wire w_dff_B_sWCLstXV1_2;
	wire w_dff_B_Gfgy7tTz8_2;
	wire w_dff_B_Twyo5fVA9_2;
	wire w_dff_B_gPVriFN42_2;
	wire w_dff_B_nmfKnA3F9_2;
	wire w_dff_B_K3HZopTd8_2;
	wire w_dff_B_Bya0IkSZ6_2;
	wire w_dff_B_WAHDLpkr5_2;
	wire w_dff_B_oJq5gcAZ4_2;
	wire w_dff_B_GdhzBQ3w5_2;
	wire w_dff_B_PvTZaMme2_2;
	wire w_dff_B_qkbJ1AV54_2;
	wire w_dff_B_3EWBsshh3_2;
	wire w_dff_B_mmDfA33w9_2;
	wire w_dff_B_EIMOwjdg0_2;
	wire w_dff_B_8Hfq9vft5_2;
	wire w_dff_B_zXPFMKne4_2;
	wire w_dff_B_4L7NdiLb8_2;
	wire w_dff_B_KeuXjNNN3_2;
	wire w_dff_B_85JFOAv87_2;
	wire w_dff_B_MMZQH4u04_2;
	wire w_dff_B_ohZ8VlNI6_2;
	wire w_dff_B_hcpIuflp3_2;
	wire w_dff_B_jLzE5Uwv9_2;
	wire w_dff_B_AN0KKKPE5_2;
	wire w_dff_B_plw1eKCA3_2;
	wire w_dff_B_WbgLpl9P7_0;
	wire w_dff_A_o830kju60_1;
	wire w_dff_B_I4hnYSxQ2_1;
	wire w_dff_B_jkJaKtAo0_2;
	wire w_dff_B_4ItMHm427_2;
	wire w_dff_B_nbYo9Rx48_2;
	wire w_dff_B_OwOa3Pot5_2;
	wire w_dff_B_f6MlyqXb1_2;
	wire w_dff_B_pzHWvknQ4_2;
	wire w_dff_B_AYkK0VcL3_2;
	wire w_dff_B_f7hrnO3D2_2;
	wire w_dff_B_4daHqpxM2_2;
	wire w_dff_B_ltOzQgEJ4_2;
	wire w_dff_B_vjG45HXm3_2;
	wire w_dff_B_m2FoSgTj2_2;
	wire w_dff_B_GEVloQc47_2;
	wire w_dff_B_B1ngRcMq1_2;
	wire w_dff_B_Zqxf87DJ3_2;
	wire w_dff_B_qey6le2O2_2;
	wire w_dff_B_8zS87Lyn8_2;
	wire w_dff_B_pbCY08Ci3_2;
	wire w_dff_B_vCleocnw7_2;
	wire w_dff_B_kgVGb8NU2_2;
	wire w_dff_B_Nh1Yluc92_2;
	wire w_dff_B_XidOhPvE0_2;
	wire w_dff_B_roFGmJYq1_2;
	wire w_dff_B_oR6ruBum6_2;
	wire w_dff_B_mnmNpu8t1_2;
	wire w_dff_B_OO6yCJeh7_2;
	wire w_dff_B_I1ZZlWbr4_2;
	wire w_dff_B_OOZZYZsv6_2;
	wire w_dff_B_JnnT4mFj7_2;
	wire w_dff_B_NjwGDvfe4_2;
	wire w_dff_B_IvMc5iTh9_2;
	wire w_dff_B_90Vlik5A7_2;
	wire w_dff_B_zj6kbofr7_2;
	wire w_dff_B_yPn4o7ol5_2;
	wire w_dff_B_Bk4DPF6d4_2;
	wire w_dff_B_QuiMGWJ42_2;
	wire w_dff_B_pqmtBimK2_2;
	wire w_dff_B_YHPlKlE47_2;
	wire w_dff_B_CofvUyBV3_2;
	wire w_dff_B_aV33VNxI7_2;
	wire w_dff_B_Y31JGknQ3_1;
	wire w_dff_B_acpUoPty5_2;
	wire w_dff_B_96J8h7BX2_2;
	wire w_dff_B_QTJ77WGC4_2;
	wire w_dff_B_ZnDgHNso0_2;
	wire w_dff_B_AqUB1R5v8_2;
	wire w_dff_B_wMyLZpig5_2;
	wire w_dff_B_TBntwDWV4_2;
	wire w_dff_B_1WpHUZwh8_2;
	wire w_dff_B_DpheNZBm7_2;
	wire w_dff_B_iIcWVjQf7_2;
	wire w_dff_B_uiRjDFcL5_2;
	wire w_dff_B_DL4b7u6b4_2;
	wire w_dff_B_AE5YTbSh3_2;
	wire w_dff_B_o0WHDeI58_2;
	wire w_dff_B_GTZxZd5X6_2;
	wire w_dff_B_NMJEzIe59_2;
	wire w_dff_B_1QPbR1Ov9_2;
	wire w_dff_B_ztOrIbZr8_2;
	wire w_dff_B_xrd6LqJy1_2;
	wire w_dff_B_dqkQ0NaF9_2;
	wire w_dff_B_w7AlJqd71_2;
	wire w_dff_B_dhmztLHM5_2;
	wire w_dff_B_itzEVHu35_2;
	wire w_dff_B_La0OAicv8_2;
	wire w_dff_B_VaBO4oAj2_2;
	wire w_dff_B_wYfqkKbE4_2;
	wire w_dff_B_6UegZdvZ1_2;
	wire w_dff_B_a1QEd8z56_2;
	wire w_dff_B_93QEYQGl0_2;
	wire w_dff_B_gbaybP8j8_2;
	wire w_dff_B_60rFZjMu3_2;
	wire w_dff_B_BtUXjWQK2_2;
	wire w_dff_B_hxDe64Qy8_2;
	wire w_dff_B_4nKzpZvV9_2;
	wire w_dff_B_oO3i39ic0_2;
	wire w_dff_B_yCfDalDw2_2;
	wire w_dff_B_bXXrmGpH8_2;
	wire w_dff_B_ldSAnnHy2_1;
	wire w_dff_B_EilGpvvI0_2;
	wire w_dff_B_1IqsQON04_2;
	wire w_dff_B_PiDytZrV8_2;
	wire w_dff_B_Vz7i4SA42_2;
	wire w_dff_B_bKIarbmF4_2;
	wire w_dff_B_6feI2gmN2_2;
	wire w_dff_B_K6i8BFwL1_2;
	wire w_dff_B_lIX68ivf3_2;
	wire w_dff_B_IN3iCCek4_2;
	wire w_dff_B_GEDQd7rQ3_2;
	wire w_dff_B_xiuvo8em2_2;
	wire w_dff_B_N615QvB30_2;
	wire w_dff_B_lLhgY6Ha1_2;
	wire w_dff_B_9lCWDov90_2;
	wire w_dff_B_lyH64LUT2_2;
	wire w_dff_B_Dos7dgYF2_2;
	wire w_dff_B_HMlrJCcl6_2;
	wire w_dff_B_3pc51oFf7_2;
	wire w_dff_B_HGvxUgeN8_2;
	wire w_dff_B_sLTAmdti4_2;
	wire w_dff_B_KNDHTW5v0_2;
	wire w_dff_B_SdOVWn6m8_2;
	wire w_dff_B_x18VzERf0_2;
	wire w_dff_B_Z8oWQsmm0_2;
	wire w_dff_B_YIvHtBNZ3_2;
	wire w_dff_B_CQnVwUjY2_2;
	wire w_dff_B_p0BB09JE1_2;
	wire w_dff_B_BU6hNa6v8_2;
	wire w_dff_B_JIHRhzCk2_2;
	wire w_dff_B_Gru3oGwW4_2;
	wire w_dff_B_Oe2IoQmu2_2;
	wire w_dff_B_QdykN0272_2;
	wire w_dff_B_XIQ0wdDi2_2;
	wire w_dff_B_hPP1DsNg0_2;
	wire w_dff_B_E7UF84ec7_1;
	wire w_dff_B_JJUTEcV79_2;
	wire w_dff_B_wb95uZfJ7_2;
	wire w_dff_B_LJKsoh0a8_2;
	wire w_dff_B_WQ639usY2_2;
	wire w_dff_B_khqkRhgq6_2;
	wire w_dff_B_N4a7jGat6_2;
	wire w_dff_B_9SDLVzEy2_2;
	wire w_dff_B_UlAGNrpR5_2;
	wire w_dff_B_m6luanHx8_2;
	wire w_dff_B_3KTBzRWX9_2;
	wire w_dff_B_00DuwbEL3_2;
	wire w_dff_B_oNuoyF3A7_2;
	wire w_dff_B_vPfTaCxx6_2;
	wire w_dff_B_eD3nbWwU9_2;
	wire w_dff_B_pBTxQ5713_2;
	wire w_dff_B_9ZZIiemO0_2;
	wire w_dff_B_9LB6HFc85_2;
	wire w_dff_B_7FaVvQxr1_2;
	wire w_dff_B_ycYhuZb70_2;
	wire w_dff_B_VqRdzQjE5_2;
	wire w_dff_B_hWqJidKw5_2;
	wire w_dff_B_iCB3jWab0_2;
	wire w_dff_B_m2v3M6pB1_2;
	wire w_dff_B_zD1LSr9q4_2;
	wire w_dff_B_LsO0OAbH8_2;
	wire w_dff_B_KUvefpuO2_2;
	wire w_dff_B_wQDQTwAC4_2;
	wire w_dff_B_RjcT4uXL9_2;
	wire w_dff_B_dhFdcFz57_2;
	wire w_dff_B_GT7w1IgP9_2;
	wire w_dff_B_3oDfo5a12_2;
	wire w_dff_B_xSfesVRc9_1;
	wire w_dff_B_ACgzCzzy6_2;
	wire w_dff_B_EpwGLWxt6_2;
	wire w_dff_B_0KCCAmmT6_2;
	wire w_dff_B_IaUUJVzR6_2;
	wire w_dff_B_p7n522pN3_2;
	wire w_dff_B_RemrzikY3_2;
	wire w_dff_B_noqfPgHG4_2;
	wire w_dff_B_ozmbDJWM2_2;
	wire w_dff_B_CxxdRRVv4_2;
	wire w_dff_B_wy24JjPb2_2;
	wire w_dff_B_3rOkTWP09_2;
	wire w_dff_B_brsTDgjn3_2;
	wire w_dff_B_JDBlXzAt8_2;
	wire w_dff_B_3QS68Yb67_2;
	wire w_dff_B_10428VuR9_2;
	wire w_dff_B_RUxOQRP63_2;
	wire w_dff_B_hhPxUJtY2_2;
	wire w_dff_B_9z4zqIHn4_2;
	wire w_dff_B_ZM71frwi0_2;
	wire w_dff_B_GANWOPY97_2;
	wire w_dff_B_EaXsR5ef7_2;
	wire w_dff_B_zBL5uHAf6_2;
	wire w_dff_B_lNTWVNJh3_2;
	wire w_dff_B_gvQiDGAg4_2;
	wire w_dff_B_jHwY5K0R5_2;
	wire w_dff_B_mXWLbgXM9_2;
	wire w_dff_B_FhOXP8Hs1_2;
	wire w_dff_B_hscgPvLM9_2;
	wire w_dff_B_mrmko7236_1;
	wire w_dff_B_ocB1jjbI3_2;
	wire w_dff_B_AUp4NN9Q9_2;
	wire w_dff_B_g3W2f0T00_2;
	wire w_dff_B_oFVbP1AG1_2;
	wire w_dff_B_XRTOGGnO0_2;
	wire w_dff_B_83PCAdnc1_2;
	wire w_dff_B_EAlun3y03_2;
	wire w_dff_B_C4Sp9jHK7_2;
	wire w_dff_B_wY7y3MAm8_2;
	wire w_dff_B_GNL0tK2o3_2;
	wire w_dff_B_BlglAkr03_2;
	wire w_dff_B_EN5gKSgN7_2;
	wire w_dff_B_JhTLyd5I4_2;
	wire w_dff_B_uqytermL2_2;
	wire w_dff_B_tm252inI4_2;
	wire w_dff_B_Z5Qox28V8_2;
	wire w_dff_B_wsCNFRPd8_2;
	wire w_dff_B_n0qtncWA4_2;
	wire w_dff_B_2LhLO1I82_2;
	wire w_dff_B_UJcDkIRb8_2;
	wire w_dff_B_HaJrmOX11_2;
	wire w_dff_B_fWLJ4b7X5_2;
	wire w_dff_B_w3HzIOnA0_2;
	wire w_dff_B_7cQ7JSZV7_2;
	wire w_dff_B_esxJIrZt0_2;
	wire w_dff_B_01Q6TyWu5_1;
	wire w_dff_B_Q0Vv8isl2_2;
	wire w_dff_B_qkTA4ZCi5_2;
	wire w_dff_B_YPgcGRzk3_2;
	wire w_dff_B_Fue7o7j42_2;
	wire w_dff_B_oMGLSwF08_2;
	wire w_dff_B_vw7MKNHx7_2;
	wire w_dff_B_OfZUjcP04_2;
	wire w_dff_B_QF3Mb0R18_2;
	wire w_dff_B_rRPojT5y0_2;
	wire w_dff_B_BqiFcAqp9_2;
	wire w_dff_B_262lAmYn2_2;
	wire w_dff_B_fj7uJlEA1_2;
	wire w_dff_B_vch0NsBX7_2;
	wire w_dff_B_Z1sKEGzN0_2;
	wire w_dff_B_2j8NJV3h3_2;
	wire w_dff_B_TjX9jPaj6_2;
	wire w_dff_B_X7LZ0EPa1_2;
	wire w_dff_B_rka0hyLL2_2;
	wire w_dff_B_1xmgAlz88_2;
	wire w_dff_B_26vWPJ9F8_2;
	wire w_dff_B_5X81MMu62_2;
	wire w_dff_B_BwJipq5t9_2;
	wire w_dff_B_bbmwRxcR6_1;
	wire w_dff_B_fq4m4c2V8_2;
	wire w_dff_B_ATKUlGrj4_2;
	wire w_dff_B_LuBiSRHd1_2;
	wire w_dff_B_jDPZHoBB1_2;
	wire w_dff_B_xiCAkGiy1_2;
	wire w_dff_B_01LedSxX2_2;
	wire w_dff_B_oBWK4tDx8_2;
	wire w_dff_B_1kqkdgZz1_2;
	wire w_dff_B_t5liWeGQ6_2;
	wire w_dff_B_93lIZMmJ3_2;
	wire w_dff_B_jeUgHtb47_2;
	wire w_dff_B_AgUTF43S0_2;
	wire w_dff_B_Hc59ebKa1_2;
	wire w_dff_B_tG8c4KYd0_2;
	wire w_dff_B_rIh6nSeB1_2;
	wire w_dff_B_yWq0szcb9_2;
	wire w_dff_B_qhsSym3h7_2;
	wire w_dff_B_mnwGxLnu0_2;
	wire w_dff_B_zuvg0Oqv6_2;
	wire w_dff_B_wgPc0zdc6_1;
	wire w_dff_B_VcL1Bh4P4_2;
	wire w_dff_B_ScNKj7PP7_2;
	wire w_dff_B_bROEBImR9_2;
	wire w_dff_B_SIamB0yQ1_2;
	wire w_dff_B_Xo46XUiJ2_2;
	wire w_dff_B_5YmWazk57_2;
	wire w_dff_B_NtzlXOCR4_2;
	wire w_dff_B_wuTxWuA16_2;
	wire w_dff_B_NQoEgRUb7_2;
	wire w_dff_B_UfutkyBZ8_2;
	wire w_dff_B_3DJ74Piq1_2;
	wire w_dff_B_9pP8DoTt6_2;
	wire w_dff_B_Zdifc1bG5_2;
	wire w_dff_B_Houm7mY63_2;
	wire w_dff_B_546d4bqi9_2;
	wire w_dff_B_1pHowUne4_2;
	wire w_dff_B_V1BaO2AM1_1;
	wire w_dff_B_6n5rAh3B4_2;
	wire w_dff_B_kmyotDWx4_2;
	wire w_dff_B_nNOGxE3k7_2;
	wire w_dff_B_ktjlnF2F2_2;
	wire w_dff_B_IojyvBFz0_2;
	wire w_dff_B_KcR8J3On6_2;
	wire w_dff_B_iZgEhadp4_2;
	wire w_dff_B_s7ibFKrE6_2;
	wire w_dff_B_l1Ufrj157_2;
	wire w_dff_B_4HYz8xk52_2;
	wire w_dff_B_MbPTzIlK1_2;
	wire w_dff_B_980k4pLA3_2;
	wire w_dff_B_AhFWDYpV0_2;
	wire w_dff_B_P4zG5qW56_1;
	wire w_dff_B_fEJ6gtzE9_2;
	wire w_dff_B_6uPCicR67_2;
	wire w_dff_B_Iu4Tv95D1_2;
	wire w_dff_B_wxtrgoak2_2;
	wire w_dff_B_ytWLxDEr9_2;
	wire w_dff_B_J9cF7xaz9_2;
	wire w_dff_B_EK5ZLz1L6_2;
	wire w_dff_B_ZY0becf17_2;
	wire w_dff_B_KI3bghAP8_2;
	wire w_dff_B_SUc5WIUE5_2;
	wire w_dff_B_9qhXiizZ6_1;
	wire w_dff_B_4R52ri585_2;
	wire w_dff_B_wwb2ZWi00_2;
	wire w_dff_B_qVa0tE9x1_2;
	wire w_dff_B_GlxKCXPs3_2;
	wire w_dff_B_iPgtyqG65_2;
	wire w_dff_B_r5l3dFb60_2;
	wire w_dff_B_F4vWvT7A0_2;
	wire w_dff_B_eTtxAsyR5_2;
	wire w_dff_B_qcV5ZJDx2_2;
	wire w_dff_B_HzLkcPRY1_2;
	wire w_dff_B_2jpNeUUR3_0;
	wire w_dff_A_71loFDDj1_0;
	wire w_dff_A_e5uR1iD21_0;
	wire w_dff_A_cW8jRnKE1_0;
	wire w_dff_A_DABRaDyw5_0;
	wire w_dff_B_63aFH6jf5_2;
	wire w_dff_B_NXjw3b0q3_1;
	wire w_dff_B_WvNCcHnA0_2;
	wire w_dff_B_f8kbonY97_2;
	wire w_dff_B_8NfIgwtA4_2;
	wire w_dff_B_2ZksKw4p4_2;
	wire w_dff_B_uJlInG0K5_2;
	wire w_dff_B_fBEpW50U9_2;
	wire w_dff_B_XYP0Xn6a7_2;
	wire w_dff_B_ZmOH45Qj1_2;
	wire w_dff_B_1xEWzVFg6_2;
	wire w_dff_B_IopllFTi0_2;
	wire w_dff_B_DNcvq4FG5_2;
	wire w_dff_B_vBptDxCp8_2;
	wire w_dff_B_JAgECIsB1_2;
	wire w_dff_B_iXRYG9OM9_2;
	wire w_dff_B_zigsYATG0_2;
	wire w_dff_B_BvKVLXxp5_2;
	wire w_dff_B_NlOVZJQk9_2;
	wire w_dff_B_jZSMzs900_2;
	wire w_dff_B_xae5irdm1_2;
	wire w_dff_B_pBanHuaK9_2;
	wire w_dff_B_tytTMAzz5_2;
	wire w_dff_B_2G6giiJ93_2;
	wire w_dff_B_pSwy0n4h3_2;
	wire w_dff_B_FQH5nr1b5_2;
	wire w_dff_B_AnmhUVRA9_2;
	wire w_dff_B_F2cpkg8H8_2;
	wire w_dff_B_pitjU4zR9_2;
	wire w_dff_B_uBkY3qeW1_2;
	wire w_dff_B_R2GrY3aD8_2;
	wire w_dff_B_Jl7i3bOb1_2;
	wire w_dff_B_zaYUQXuh4_2;
	wire w_dff_B_ubN5tJLJ2_2;
	wire w_dff_B_M092GrGo9_2;
	wire w_dff_B_WNO4BPVO5_2;
	wire w_dff_B_OmOUMwOM4_2;
	wire w_dff_B_kaNslhL44_2;
	wire w_dff_B_cqXn2RsE7_2;
	wire w_dff_B_1bs89Hry2_2;
	wire w_dff_B_kbo3ePki4_2;
	wire w_dff_B_g9IC65jP2_2;
	wire w_dff_B_vaMCqxmS3_2;
	wire w_dff_B_mYVREC2A6_2;
	wire w_dff_B_0x579tDP8_2;
	wire w_dff_B_bG0rai9o5_2;
	wire w_dff_B_IZi3Ndf67_1;
	wire w_dff_B_s0RBPDHg1_2;
	wire w_dff_B_HanLoImk7_2;
	wire w_dff_B_i0pgx0Z16_2;
	wire w_dff_B_iBy4ifVi2_2;
	wire w_dff_B_vvZ4gUhA0_2;
	wire w_dff_B_BJx4rVKg0_2;
	wire w_dff_B_qlJRZGE67_2;
	wire w_dff_B_G7W6kMJl5_2;
	wire w_dff_B_5MNwe50O3_2;
	wire w_dff_B_FTIZ3PTc0_2;
	wire w_dff_B_iJTd623c1_2;
	wire w_dff_B_wkqF6ASz4_2;
	wire w_dff_B_Lu7EvZan6_2;
	wire w_dff_B_mKMRxdbQ6_2;
	wire w_dff_B_d4f1OTzO1_2;
	wire w_dff_B_wkEdgNyA8_2;
	wire w_dff_B_qTliLYmf8_2;
	wire w_dff_B_bmAX0loh9_2;
	wire w_dff_B_I5evKUXl8_2;
	wire w_dff_B_cAl4t5yr7_2;
	wire w_dff_B_MAC51qts6_2;
	wire w_dff_B_L9WLI6E84_2;
	wire w_dff_B_e1YpAWm89_2;
	wire w_dff_B_fmkLYH6Y3_2;
	wire w_dff_B_f7nwM4HE0_2;
	wire w_dff_B_3DklKBKb4_2;
	wire w_dff_B_m7nhDawH8_2;
	wire w_dff_B_twoavS7N1_2;
	wire w_dff_B_1EZMyTPq3_2;
	wire w_dff_B_K3pDCnNB2_2;
	wire w_dff_B_YsxVunNc3_2;
	wire w_dff_B_TrjhvAcA3_2;
	wire w_dff_B_5o002yxn8_2;
	wire w_dff_B_0elspNfO9_2;
	wire w_dff_B_8DFGrMkU5_2;
	wire w_dff_B_rUGFPC6f3_2;
	wire w_dff_B_ex0Bfp8v6_2;
	wire w_dff_B_0Mw3Lr6J3_2;
	wire w_dff_B_xDLoDmzC7_2;
	wire w_dff_B_5a7iCyKw7_1;
	wire w_dff_B_xWuhoX1X7_2;
	wire w_dff_B_h95ajs822_2;
	wire w_dff_B_uMhWJFrQ3_2;
	wire w_dff_B_W4LQSCaJ2_2;
	wire w_dff_B_LM7e9pCe9_2;
	wire w_dff_B_pQb67gyp1_2;
	wire w_dff_B_nfUE4tXR6_2;
	wire w_dff_B_pUNhOJ6l1_2;
	wire w_dff_B_zbVRkb4F0_2;
	wire w_dff_B_olFUxNMp8_2;
	wire w_dff_B_BojOT41K0_2;
	wire w_dff_B_m0Q8sLYB5_2;
	wire w_dff_B_r7Mjqsdp4_2;
	wire w_dff_B_O6O25vXp3_2;
	wire w_dff_B_AoYe3P4t7_2;
	wire w_dff_B_EHDWu3SD6_2;
	wire w_dff_B_ZVfuvzi73_2;
	wire w_dff_B_9C29qdIr1_2;
	wire w_dff_B_X5MY2tUt9_2;
	wire w_dff_B_Ogz8plhk6_2;
	wire w_dff_B_UPlVshC21_2;
	wire w_dff_B_mvvDJxYs1_2;
	wire w_dff_B_oMYsIgpL8_2;
	wire w_dff_B_PreNpc8t8_2;
	wire w_dff_B_oG5d7WuC0_2;
	wire w_dff_B_vg6e87IX2_2;
	wire w_dff_B_RKLdNgBi0_2;
	wire w_dff_B_lofPN2A51_2;
	wire w_dff_B_iypVaiuf5_2;
	wire w_dff_B_sDLTB4A11_2;
	wire w_dff_B_OiK8AIAa3_2;
	wire w_dff_B_LzUwFY2H5_2;
	wire w_dff_B_k0tfvsBB0_2;
	wire w_dff_B_PzPgs8xv5_2;
	wire w_dff_B_NBnXsbqy3_2;
	wire w_dff_B_3asv6Oq43_2;
	wire w_dff_B_68zJrRQn6_1;
	wire w_dff_B_5OwEFkNk1_2;
	wire w_dff_B_6AfpDX0Q5_2;
	wire w_dff_B_26Pxisgh1_2;
	wire w_dff_B_JWMmyMSp1_2;
	wire w_dff_B_KLbaXe9X5_2;
	wire w_dff_B_zdqxO4HL0_2;
	wire w_dff_B_93Oe04y36_2;
	wire w_dff_B_jos6fRZi3_2;
	wire w_dff_B_6te7F88y9_2;
	wire w_dff_B_lsfY90UX1_2;
	wire w_dff_B_gLAVDZFi7_2;
	wire w_dff_B_h9r6XC8H2_2;
	wire w_dff_B_37yEnHBD8_2;
	wire w_dff_B_XQBSTqUz2_2;
	wire w_dff_B_xFo5YbXJ5_2;
	wire w_dff_B_eR3Rib7Z5_2;
	wire w_dff_B_VJN6Tcim2_2;
	wire w_dff_B_vJZdUpQX3_2;
	wire w_dff_B_V586TrTw1_2;
	wire w_dff_B_P5tkvkhM7_2;
	wire w_dff_B_BRKgUOf11_2;
	wire w_dff_B_yPMyfZje9_2;
	wire w_dff_B_ZIjmV4ZI3_2;
	wire w_dff_B_BoQb4wAr7_2;
	wire w_dff_B_j6wsByxZ4_2;
	wire w_dff_B_VjWvqrvv0_2;
	wire w_dff_B_GuVVIFjE3_2;
	wire w_dff_B_HFFPNWWF1_2;
	wire w_dff_B_N2o7P2Iu6_2;
	wire w_dff_B_JkOHAxqH1_2;
	wire w_dff_B_Vx0eqJSd2_2;
	wire w_dff_B_7SaKbanj4_2;
	wire w_dff_B_JxLDU3Sf6_2;
	wire w_dff_B_Nkz8yQSe9_1;
	wire w_dff_B_oPWwfmOW2_2;
	wire w_dff_B_PDRDQaFX9_2;
	wire w_dff_B_jHHJ8PDx1_2;
	wire w_dff_B_7Xo00ENa2_2;
	wire w_dff_B_i6tYNkW57_2;
	wire w_dff_B_4qVXhN027_2;
	wire w_dff_B_HLzOduDW4_2;
	wire w_dff_B_91Bkjm9r1_2;
	wire w_dff_B_pUeuR6Vw4_2;
	wire w_dff_B_44gx8QK28_2;
	wire w_dff_B_IBDQiS018_2;
	wire w_dff_B_ZBibaqdY2_2;
	wire w_dff_B_wSjEQpSB5_2;
	wire w_dff_B_Uzxdb5j56_2;
	wire w_dff_B_EIawDFfw6_2;
	wire w_dff_B_nrWNiFgD4_2;
	wire w_dff_B_Z87vWLnY3_2;
	wire w_dff_B_uUyHDpO56_2;
	wire w_dff_B_d5fzpVRe0_2;
	wire w_dff_B_rkYMmdb34_2;
	wire w_dff_B_Gnv8Uims4_2;
	wire w_dff_B_sds1cPBn4_2;
	wire w_dff_B_0CgY84cr6_2;
	wire w_dff_B_KFEh2fMa6_2;
	wire w_dff_B_KXruVjqQ3_2;
	wire w_dff_B_rXhW6QRZ7_2;
	wire w_dff_B_7d3MHg1i2_2;
	wire w_dff_B_5rJqiBB32_2;
	wire w_dff_B_mTaS2yNp5_2;
	wire w_dff_B_GETyUF4i3_2;
	wire w_dff_B_3xx9tJ5y5_1;
	wire w_dff_B_XQYEf3Bs7_2;
	wire w_dff_B_w2dm33815_2;
	wire w_dff_B_wnBR6JA50_2;
	wire w_dff_B_D8xKpJzf6_2;
	wire w_dff_B_XMZRe6bd6_2;
	wire w_dff_B_xMHIbwiF4_2;
	wire w_dff_B_x1pnD8RP4_2;
	wire w_dff_B_WQk8WZbI9_2;
	wire w_dff_B_9Z23VAxT0_2;
	wire w_dff_B_SDqwmYCU9_2;
	wire w_dff_B_pY0hJPWK9_2;
	wire w_dff_B_LTdyYCPM6_2;
	wire w_dff_B_HdBg7PPq7_2;
	wire w_dff_B_9byKDIrc7_2;
	wire w_dff_B_AHT48S058_2;
	wire w_dff_B_cB4Q6WJd3_2;
	wire w_dff_B_Z6V9HleY5_2;
	wire w_dff_B_xtNDmmBm2_2;
	wire w_dff_B_nrsyw6Nw7_2;
	wire w_dff_B_Frc572ea5_2;
	wire w_dff_B_1htllQC45_2;
	wire w_dff_B_XrFlQZ0f1_2;
	wire w_dff_B_CsaZPo1K9_2;
	wire w_dff_B_9mMRclRs6_2;
	wire w_dff_B_L1plQ7BJ1_2;
	wire w_dff_B_2ZzMFQ423_2;
	wire w_dff_B_1e5eJ58E4_2;
	wire w_dff_B_b0QFyRaJ4_1;
	wire w_dff_B_wH2FGRmR6_2;
	wire w_dff_B_7UsRrJa37_2;
	wire w_dff_B_qEwEU1VK5_2;
	wire w_dff_B_KrWbVi1o5_2;
	wire w_dff_B_OFj3II7e4_2;
	wire w_dff_B_wQuKQmho0_2;
	wire w_dff_B_rFM4KIgO3_2;
	wire w_dff_B_KwweXWJv6_2;
	wire w_dff_B_84x0jNk58_2;
	wire w_dff_B_wmXsjXrg8_2;
	wire w_dff_B_zpwBuqvP2_2;
	wire w_dff_B_sAQQOZ1Q3_2;
	wire w_dff_B_Dl3O1mtC9_2;
	wire w_dff_B_Yc9nggDa1_2;
	wire w_dff_B_4OP5NqJ49_2;
	wire w_dff_B_k4bqxa922_2;
	wire w_dff_B_daLnpbxA3_2;
	wire w_dff_B_S6m8QAh92_2;
	wire w_dff_B_MwqVd59X2_2;
	wire w_dff_B_2HiMGl5j1_2;
	wire w_dff_B_yemd9cAo9_2;
	wire w_dff_B_KrDsOy8L9_2;
	wire w_dff_B_6UDR1fBH9_2;
	wire w_dff_B_bTlMXmHN0_2;
	wire w_dff_B_a5hMvIXr4_1;
	wire w_dff_B_95TFH98x2_2;
	wire w_dff_B_FDB44I3s9_2;
	wire w_dff_B_ZRB8TWo86_2;
	wire w_dff_B_HuVF1xcf4_2;
	wire w_dff_B_5FPRP90C4_2;
	wire w_dff_B_qSveOskZ7_2;
	wire w_dff_B_IRLLnjOa4_2;
	wire w_dff_B_YxIoEKj84_2;
	wire w_dff_B_G6eUWOPl2_2;
	wire w_dff_B_RJY2uDu19_2;
	wire w_dff_B_mQhis6j15_2;
	wire w_dff_B_vk9FTMO82_2;
	wire w_dff_B_lLkldlYr8_2;
	wire w_dff_B_KmsgppnI8_2;
	wire w_dff_B_CVt3WYV58_2;
	wire w_dff_B_d5Ww78tP8_2;
	wire w_dff_B_51b1fma64_2;
	wire w_dff_B_m3qBvm096_2;
	wire w_dff_B_gWGqX1cA0_2;
	wire w_dff_B_9bJyjAPO7_2;
	wire w_dff_B_2KqAnSEU2_2;
	wire w_dff_B_SSFrj5Nk1_1;
	wire w_dff_B_qFoG6pek1_2;
	wire w_dff_B_BC4DsAIz2_2;
	wire w_dff_B_dyvud0fw6_2;
	wire w_dff_B_Z3gK0SMQ1_2;
	wire w_dff_B_8zz5iqBf0_2;
	wire w_dff_B_mCLqynJs3_2;
	wire w_dff_B_FBFMEVqD8_2;
	wire w_dff_B_SfHG0bQ89_2;
	wire w_dff_B_lzBz9qpK8_2;
	wire w_dff_B_zufUWRD91_2;
	wire w_dff_B_wLEgturd6_2;
	wire w_dff_B_orYTpMRz5_2;
	wire w_dff_B_n0Cmn7y92_2;
	wire w_dff_B_Y6FP9So05_2;
	wire w_dff_B_e38GIF168_2;
	wire w_dff_B_8W6mVw9a0_2;
	wire w_dff_B_lp1IivzI1_2;
	wire w_dff_B_PIUi5LCX0_2;
	wire w_dff_B_b6JibRo52_1;
	wire w_dff_B_uDq8J1XC0_2;
	wire w_dff_B_q9b7ZXoW7_2;
	wire w_dff_B_guXcKO6u4_2;
	wire w_dff_B_Jhv0cexv3_2;
	wire w_dff_B_SWTulCdI1_2;
	wire w_dff_B_V5JIIkF60_2;
	wire w_dff_B_P7aYFYCH8_2;
	wire w_dff_B_ETEoCqUj7_2;
	wire w_dff_B_9p4VykO81_2;
	wire w_dff_B_Nkvt1q1B3_2;
	wire w_dff_B_gVJ1WyDN5_2;
	wire w_dff_B_kNjXTNPM3_2;
	wire w_dff_B_17tYhwAN7_2;
	wire w_dff_B_sIc9ZKYP3_2;
	wire w_dff_B_74u6g0wf4_2;
	wire w_dff_B_HyF84s1z6_1;
	wire w_dff_B_QJgOlO5S3_2;
	wire w_dff_B_VC5AI2cE2_2;
	wire w_dff_B_6jvrfecC2_2;
	wire w_dff_B_LHqolNIR7_2;
	wire w_dff_B_Lc13rufq5_2;
	wire w_dff_B_0iV3cD4D1_2;
	wire w_dff_B_eslJJmNt6_2;
	wire w_dff_B_5Mytq3hu9_2;
	wire w_dff_B_15wlhsPs1_2;
	wire w_dff_B_ZadxiPV94_2;
	wire w_dff_B_kbKgaLLY7_2;
	wire w_dff_B_h9fjyNnY5_2;
	wire w_dff_B_MeQzjXfG9_1;
	wire w_dff_B_ZejeJu0H2_2;
	wire w_dff_B_9ommu0Cu8_2;
	wire w_dff_B_aXbMf3v88_2;
	wire w_dff_B_hRxqR5J26_2;
	wire w_dff_B_3wDR3Q5p8_2;
	wire w_dff_B_AhWySDnr8_2;
	wire w_dff_B_MHIfGEIW1_2;
	wire w_dff_B_TIHxiZXZ5_2;
	wire w_dff_B_UKDO5yzq0_2;
	wire w_dff_B_o71vjIz19_2;
	wire w_dff_B_d4C0Djht4_1;
	wire w_dff_B_QLmmHdBd3_2;
	wire w_dff_B_AD6FBGMr9_2;
	wire w_dff_B_yU97FjGZ8_2;
	wire w_dff_B_nQ8IACQD3_2;
	wire w_dff_B_aOg66IsC9_2;
	wire w_dff_B_nzEs7aAK5_2;
	wire w_dff_B_9ig1YyJM9_2;
	wire w_dff_B_PO4Y0hsc6_2;
	wire w_dff_B_PDaul29w4_2;
	wire w_dff_B_moe5ArhA2_2;
	wire w_dff_B_R06sGySs5_0;
	wire w_dff_A_avPaiqt82_0;
	wire w_dff_A_d0yTcVi09_0;
	wire w_dff_A_lmAUvAnN9_1;
	wire w_dff_A_Pm0Nd7zt9_1;
	wire w_dff_B_7IYrndFR5_2;
	wire w_dff_B_fcHIml3A7_1;
	wire w_dff_B_VByecPze9_2;
	wire w_dff_B_bnwwtrCn4_2;
	wire w_dff_B_qT3ZAFbp1_2;
	wire w_dff_B_uhMyfmmT5_2;
	wire w_dff_B_QEK7rfsY1_2;
	wire w_dff_B_9vpFs3On0_2;
	wire w_dff_B_YATb2Jj04_2;
	wire w_dff_B_EUSs6NCu4_2;
	wire w_dff_B_HoK8i75Z1_2;
	wire w_dff_B_QlNHCHsO0_2;
	wire w_dff_B_lzz0N8Uc5_2;
	wire w_dff_B_pPBQNrSV0_2;
	wire w_dff_B_Bs8SAgra7_2;
	wire w_dff_B_Q2eQFoDZ2_2;
	wire w_dff_B_4e4g0vIF9_2;
	wire w_dff_B_NIctntP14_2;
	wire w_dff_B_DPkKJCks4_2;
	wire w_dff_B_Sg6DnKlH5_2;
	wire w_dff_B_m6rfshPa9_2;
	wire w_dff_B_kv0gVde97_2;
	wire w_dff_B_LYAK9hG93_2;
	wire w_dff_B_3nU1rMaH3_2;
	wire w_dff_B_Yvk8M88Y8_2;
	wire w_dff_B_qow4P8zI1_2;
	wire w_dff_B_zy8II2T83_2;
	wire w_dff_B_hXMnjQfh8_2;
	wire w_dff_B_QkH2Hj617_2;
	wire w_dff_B_aBGDm4q65_2;
	wire w_dff_B_9YmMe76O7_2;
	wire w_dff_B_gtvk1xKi7_2;
	wire w_dff_B_SPqnErfz3_2;
	wire w_dff_B_iVZ44Ixp2_2;
	wire w_dff_B_a4Cj5tGN0_2;
	wire w_dff_B_gdkYer2Z1_2;
	wire w_dff_B_zJSwEd6f6_2;
	wire w_dff_B_OQ9pBsmO5_2;
	wire w_dff_B_vfvCQtii6_2;
	wire w_dff_B_N5nte4gK0_2;
	wire w_dff_B_vaU8AVxB7_2;
	wire w_dff_B_drAzDmhn5_2;
	wire w_dff_B_3tOTKcic8_2;
	wire w_dff_B_GSLVi2KG7_2;
	wire w_dff_B_0bc0jAd24_2;
	wire w_dff_B_fZkY1zIB6_2;
	wire w_dff_B_Pd21kpZx1_2;
	wire w_dff_B_xAz4mD5f3_1;
	wire w_dff_B_q6BFgqL85_2;
	wire w_dff_B_jigvGq0e2_2;
	wire w_dff_B_dVV9qFXZ5_2;
	wire w_dff_B_qssjqL4Q9_2;
	wire w_dff_B_sQ7DaFdy4_2;
	wire w_dff_B_6MDUZfcK1_2;
	wire w_dff_B_UruRfHuH3_2;
	wire w_dff_B_44iIadLG0_2;
	wire w_dff_B_pFGvHN1P6_2;
	wire w_dff_B_Jwm96ixk5_2;
	wire w_dff_B_MVuqNFAQ4_2;
	wire w_dff_B_LJ5MIyFT5_2;
	wire w_dff_B_olNavd7w7_2;
	wire w_dff_B_hnMyeiQQ8_2;
	wire w_dff_B_zB8CuPwy5_2;
	wire w_dff_B_DnGTPm9q1_2;
	wire w_dff_B_qWJRcS0Q2_2;
	wire w_dff_B_iqPujPyG7_2;
	wire w_dff_B_jAzmZZl82_2;
	wire w_dff_B_O6SonGJW2_2;
	wire w_dff_B_RPAuD1L04_2;
	wire w_dff_B_imRTaY8j3_2;
	wire w_dff_B_9Fyvj60o4_2;
	wire w_dff_B_aqEN59Os0_2;
	wire w_dff_B_2UUaVsUM1_2;
	wire w_dff_B_kfFmmocH7_2;
	wire w_dff_B_zFGf6PEK0_2;
	wire w_dff_B_YEw0aEIl7_2;
	wire w_dff_B_yIvWOSUj2_2;
	wire w_dff_B_Kplq0gJX7_2;
	wire w_dff_B_nkLYM3ov8_2;
	wire w_dff_B_Gwh5F2ak5_2;
	wire w_dff_B_mZJnrehT5_2;
	wire w_dff_B_WTzdh0vQ9_2;
	wire w_dff_B_oyip6Zpf3_2;
	wire w_dff_B_unzYtWQN5_2;
	wire w_dff_B_cvWtVvmy8_2;
	wire w_dff_B_RSoabqlo7_2;
	wire w_dff_B_SN2A4cA76_2;
	wire w_dff_B_tgvlIUag2_2;
	wire w_dff_B_p1ySQhIb4_1;
	wire w_dff_B_0jZhwfd52_2;
	wire w_dff_B_bwv6OI9X1_2;
	wire w_dff_B_w2r9OyeU9_2;
	wire w_dff_B_uJ3TkUiB6_2;
	wire w_dff_B_iQ6HjADO4_2;
	wire w_dff_B_oSJSHojw6_2;
	wire w_dff_B_8GMGOIep7_2;
	wire w_dff_B_WlWy4VaC6_2;
	wire w_dff_B_heGH44ag4_2;
	wire w_dff_B_4PqX7Zab3_2;
	wire w_dff_B_lpC4r68j0_2;
	wire w_dff_B_LXd1zZoD3_2;
	wire w_dff_B_BiXd18tC1_2;
	wire w_dff_B_CawyenJ93_2;
	wire w_dff_B_CFu21fDh7_2;
	wire w_dff_B_omETCELq1_2;
	wire w_dff_B_iUBFLVxG4_2;
	wire w_dff_B_IEFrqQnV0_2;
	wire w_dff_B_CdsExHPx0_2;
	wire w_dff_B_W8nbYeAN8_2;
	wire w_dff_B_Rwq1Dclc9_2;
	wire w_dff_B_Ja0QR4Ji5_2;
	wire w_dff_B_97D0QIxU7_2;
	wire w_dff_B_gqzqYgfg4_2;
	wire w_dff_B_Fx2RNUbk9_2;
	wire w_dff_B_XxquX4TF3_2;
	wire w_dff_B_DsH4y2Yt3_2;
	wire w_dff_B_UMuBHyn88_2;
	wire w_dff_B_erApfxOA6_2;
	wire w_dff_B_u2xWP5EJ2_2;
	wire w_dff_B_OvQo1C3o7_2;
	wire w_dff_B_Ogqofr107_2;
	wire w_dff_B_2nNPAo0D7_2;
	wire w_dff_B_Jd6l7w2P9_2;
	wire w_dff_B_qUd31gLq9_2;
	wire w_dff_B_gwwqRqOS0_2;
	wire w_dff_B_2TijpYi78_2;
	wire w_dff_B_Ncrix9Co4_1;
	wire w_dff_B_Y8wFsNR74_2;
	wire w_dff_B_Vg88ocSZ6_2;
	wire w_dff_B_zV0LuOs57_2;
	wire w_dff_B_hMxudX500_2;
	wire w_dff_B_s8ceWCYO4_2;
	wire w_dff_B_oyf71azQ6_2;
	wire w_dff_B_Hap07XHV0_2;
	wire w_dff_B_XAircJLx3_2;
	wire w_dff_B_2FoMNE2y9_2;
	wire w_dff_B_pY9HX9700_2;
	wire w_dff_B_7ZG8p6cb1_2;
	wire w_dff_B_txF6M97S4_2;
	wire w_dff_B_onCvetXI5_2;
	wire w_dff_B_DRd4W0KS2_2;
	wire w_dff_B_wHqNAGMY0_2;
	wire w_dff_B_opYE9eWC2_2;
	wire w_dff_B_sgkrrRGD7_2;
	wire w_dff_B_IVCPit3L1_2;
	wire w_dff_B_5KKygy3C9_2;
	wire w_dff_B_T2X5e5yQ8_2;
	wire w_dff_B_zKuZnUrH6_2;
	wire w_dff_B_Ef1DAYzs8_2;
	wire w_dff_B_Kpk2ZwEA6_2;
	wire w_dff_B_h7zqUyKf9_2;
	wire w_dff_B_FEBK82sH3_2;
	wire w_dff_B_K0zobonR7_2;
	wire w_dff_B_BEqFulR19_2;
	wire w_dff_B_C0fQjyRv5_2;
	wire w_dff_B_bVOlXeOK6_2;
	wire w_dff_B_2aCrStZ59_2;
	wire w_dff_B_VvNG1HuI7_2;
	wire w_dff_B_5EEBvNvP7_2;
	wire w_dff_B_lgYGEJcS8_2;
	wire w_dff_B_O7NpO5ou1_2;
	wire w_dff_B_mSgxvJiU9_1;
	wire w_dff_B_U1c0qcFe6_2;
	wire w_dff_B_dspjIlW31_2;
	wire w_dff_B_yqWxRizk1_2;
	wire w_dff_B_iAoyfUpp6_2;
	wire w_dff_B_71slUsZz2_2;
	wire w_dff_B_srbUcKaG7_2;
	wire w_dff_B_RBHC6Fcb4_2;
	wire w_dff_B_4J1vW2Yx1_2;
	wire w_dff_B_9kO19CQ53_2;
	wire w_dff_B_AdGsBN6o7_2;
	wire w_dff_B_A4wK2cUz5_2;
	wire w_dff_B_mY7vJ0G82_2;
	wire w_dff_B_WIL0UxPW3_2;
	wire w_dff_B_IV2gujoy4_2;
	wire w_dff_B_tMXdvZbI5_2;
	wire w_dff_B_nYp4JGmM8_2;
	wire w_dff_B_CHaodq9V6_2;
	wire w_dff_B_yJIvjSgk6_2;
	wire w_dff_B_6pcU0j1Q8_2;
	wire w_dff_B_sMRXcpsK7_2;
	wire w_dff_B_vtP9k1hW9_2;
	wire w_dff_B_cid6UOIn7_2;
	wire w_dff_B_UeWIvyM95_2;
	wire w_dff_B_Y5dPiKLC6_2;
	wire w_dff_B_Ue23enFQ0_2;
	wire w_dff_B_givJpf8v0_2;
	wire w_dff_B_hHa1j1AN3_2;
	wire w_dff_B_S5y9SNT34_2;
	wire w_dff_B_y6vpjOxy1_2;
	wire w_dff_B_xQciGphy7_2;
	wire w_dff_B_x2SPxzy90_2;
	wire w_dff_B_cqPJn0w51_1;
	wire w_dff_B_fq1BFHsr5_2;
	wire w_dff_B_cSzjWdue0_2;
	wire w_dff_B_JBEwOUys6_2;
	wire w_dff_B_mtfWq1CC7_2;
	wire w_dff_B_JQQkmHbq4_2;
	wire w_dff_B_4wTDaToZ7_2;
	wire w_dff_B_NmSPOJLx6_2;
	wire w_dff_B_eaefrATz8_2;
	wire w_dff_B_mtJULdaF2_2;
	wire w_dff_B_RiUjBtlv3_2;
	wire w_dff_B_CAOi4r8W1_2;
	wire w_dff_B_osF680Ms8_2;
	wire w_dff_B_uqs5i3tY6_2;
	wire w_dff_B_y8oaetqd4_2;
	wire w_dff_B_rQGcMrEs9_2;
	wire w_dff_B_BRNtNuXT4_2;
	wire w_dff_B_4Sx2gh6V7_2;
	wire w_dff_B_sBLIjZ9m4_2;
	wire w_dff_B_X4ong0Kj4_2;
	wire w_dff_B_rHnL7PN81_2;
	wire w_dff_B_uKCbPCPY7_2;
	wire w_dff_B_S02Bfd0r7_2;
	wire w_dff_B_nP7Fmwkm2_2;
	wire w_dff_B_dVGylOsn2_2;
	wire w_dff_B_hPuH5TjQ2_2;
	wire w_dff_B_5qNVlcW28_2;
	wire w_dff_B_1jpj3San1_2;
	wire w_dff_B_APlCJvM38_2;
	wire w_dff_B_oHrmig9b8_1;
	wire w_dff_B_rkfsy30s1_2;
	wire w_dff_B_Mxo3yYls4_2;
	wire w_dff_B_FqyUuTVD5_2;
	wire w_dff_B_SMxuUzVq0_2;
	wire w_dff_B_5dsBJsfb2_2;
	wire w_dff_B_Ty9VgCsB4_2;
	wire w_dff_B_F2dQohVp4_2;
	wire w_dff_B_DradSCFZ6_2;
	wire w_dff_B_jMoggx2e1_2;
	wire w_dff_B_BUhoAFux1_2;
	wire w_dff_B_m0OZvkKe2_2;
	wire w_dff_B_4t4LIWnU8_2;
	wire w_dff_B_48IWPnwM2_2;
	wire w_dff_B_LSjNWVPQ1_2;
	wire w_dff_B_fu1ZQUaY3_2;
	wire w_dff_B_yJfrJwUh2_2;
	wire w_dff_B_75uPTHOI5_2;
	wire w_dff_B_oZ2MO2l11_2;
	wire w_dff_B_hfvKoMDr7_2;
	wire w_dff_B_wyR6zR8Z8_2;
	wire w_dff_B_u2l2OQMG6_2;
	wire w_dff_B_BpOj8OnA6_2;
	wire w_dff_B_RaYknB3l7_2;
	wire w_dff_B_SunJ3O1y4_2;
	wire w_dff_B_UyzY5MlU4_2;
	wire w_dff_B_Ev4CQdpk0_1;
	wire w_dff_B_0pM1aYEb6_2;
	wire w_dff_B_3GWtVEYO3_2;
	wire w_dff_B_IX4X35ka6_2;
	wire w_dff_B_DVDEdXfi1_2;
	wire w_dff_B_kebgbYYS2_2;
	wire w_dff_B_s0jgHSUe3_2;
	wire w_dff_B_5M9CLjh65_2;
	wire w_dff_B_Uas4CeUS6_2;
	wire w_dff_B_Znvr1vFd2_2;
	wire w_dff_B_eKXQWiGV8_2;
	wire w_dff_B_NsFZQH9p6_2;
	wire w_dff_B_6E1N0qgj9_2;
	wire w_dff_B_ctiY2GBW2_2;
	wire w_dff_B_FSOn4wq39_2;
	wire w_dff_B_03w5wrtF0_2;
	wire w_dff_B_BXDoiOag6_2;
	wire w_dff_B_KujAZ5lW0_2;
	wire w_dff_B_SCiVOBJu5_2;
	wire w_dff_B_CjUmJcZb7_2;
	wire w_dff_B_dozsRspm0_2;
	wire w_dff_B_FD27LYtI0_2;
	wire w_dff_B_DgxOZg6R1_2;
	wire w_dff_B_uh9KG59w7_1;
	wire w_dff_B_khBAQAxY9_2;
	wire w_dff_B_1a3P04YC0_2;
	wire w_dff_B_1eVCw3IS4_2;
	wire w_dff_B_cXspYIdS7_2;
	wire w_dff_B_yOndADZW7_2;
	wire w_dff_B_aId95FVP0_2;
	wire w_dff_B_Zp74O74J9_2;
	wire w_dff_B_R2N939fv4_2;
	wire w_dff_B_m0DtOOQ88_2;
	wire w_dff_B_OKb7n73E7_2;
	wire w_dff_B_Knb5uX1Z5_2;
	wire w_dff_B_KGi53uo27_2;
	wire w_dff_B_hziZrZsd5_2;
	wire w_dff_B_bIXaZiWu4_2;
	wire w_dff_B_qscKhjSK6_2;
	wire w_dff_B_1grgBQC35_2;
	wire w_dff_B_mkGiDRUD8_2;
	wire w_dff_B_wVmiFhGN1_2;
	wire w_dff_B_cbKJmi6f7_2;
	wire w_dff_B_bPimEsZa9_1;
	wire w_dff_B_rWJETwad5_2;
	wire w_dff_B_RnOIm7mA1_2;
	wire w_dff_B_2XDlsdfZ8_2;
	wire w_dff_B_7hHJbMH16_2;
	wire w_dff_B_YL4rz5Oc4_2;
	wire w_dff_B_BBAL9Mm45_2;
	wire w_dff_B_4W6g83Ap5_2;
	wire w_dff_B_kbnzJNs73_2;
	wire w_dff_B_uiGck9g12_2;
	wire w_dff_B_w9vMPKL08_2;
	wire w_dff_B_NSeJwMri3_2;
	wire w_dff_B_TcPTESMx8_2;
	wire w_dff_B_T8WafdQk1_2;
	wire w_dff_B_8LVRvV5P4_2;
	wire w_dff_B_USbybAmP6_2;
	wire w_dff_B_NAIXv9WN7_2;
	wire w_dff_B_Op82aIIH5_1;
	wire w_dff_B_5fzhd01t4_2;
	wire w_dff_B_Q1EulNwY6_2;
	wire w_dff_B_AECID8ag8_2;
	wire w_dff_B_Chug2rJ45_2;
	wire w_dff_B_ZAKizlQK3_2;
	wire w_dff_B_K433J3Fj6_2;
	wire w_dff_B_iZsWPgul7_2;
	wire w_dff_B_fjdZW6g19_2;
	wire w_dff_B_enosXykL2_2;
	wire w_dff_B_sZrhq1Gf8_2;
	wire w_dff_B_z31PjNrX4_2;
	wire w_dff_B_ipLRqzef3_2;
	wire w_dff_B_hnVkheOv4_2;
	wire w_dff_B_vOu5VeOi2_1;
	wire w_dff_B_l59LYDJ84_2;
	wire w_dff_B_y8rb9ITS0_2;
	wire w_dff_B_SqeNrBCI9_2;
	wire w_dff_B_uOME5WZa9_2;
	wire w_dff_B_582O5wJe8_2;
	wire w_dff_B_9T145DRs4_2;
	wire w_dff_B_0O3cDWAy8_2;
	wire w_dff_B_m4MiRyCc2_2;
	wire w_dff_B_dH3500ym3_2;
	wire w_dff_B_jOYZKkVE5_2;
	wire w_dff_B_WbZgNx2W0_2;
	wire w_dff_B_HLZqCbhz3_1;
	wire w_dff_B_vdT1MCRY4_2;
	wire w_dff_B_n0IvnRvw2_2;
	wire w_dff_B_UhWQDQaU0_2;
	wire w_dff_B_cHuZeCJF9_2;
	wire w_dff_B_JiTexVVI6_2;
	wire w_dff_B_pKLuxngU2_2;
	wire w_dff_B_v1WaF1H94_2;
	wire w_dff_B_equHhrx92_2;
	wire w_dff_B_mP9gkpxo4_2;
	wire w_dff_B_xGVVmCvC2_2;
	wire w_dff_B_Nlus2vSY4_0;
	wire w_dff_A_UtJmcRHB7_0;
	wire w_dff_A_wPraWFFy9_0;
	wire w_dff_A_6eIcQALi3_1;
	wire w_dff_A_VyoFlOGM9_1;
	wire w_dff_B_Jk58wg5I9_1;
	wire w_dff_B_VswOaHDp8_2;
	wire w_dff_B_gyQuQIR00_2;
	wire w_dff_B_PWuIdnru6_2;
	wire w_dff_B_rrAS1YKE4_2;
	wire w_dff_B_jDGzIUPu7_2;
	wire w_dff_B_qAueXGVO4_2;
	wire w_dff_B_1wm2OyUI1_2;
	wire w_dff_B_otHU9EIX4_2;
	wire w_dff_B_i0R3tGtH7_2;
	wire w_dff_B_ysPxCx4m1_2;
	wire w_dff_B_JHLSWOjB5_2;
	wire w_dff_B_GHJNnxQR7_2;
	wire w_dff_B_Jb9rvoFV0_2;
	wire w_dff_B_wYKYUiNB6_2;
	wire w_dff_B_ijcB46EL8_2;
	wire w_dff_B_94t7fViY5_2;
	wire w_dff_B_jtTjHHDr1_2;
	wire w_dff_B_fjn5SRUZ0_2;
	wire w_dff_B_WSmMpNTo0_2;
	wire w_dff_B_9siyY3d93_2;
	wire w_dff_B_B2PypJQY7_2;
	wire w_dff_B_3CmrlFIu6_2;
	wire w_dff_B_fcglWAlY8_2;
	wire w_dff_B_aWnC45ll6_2;
	wire w_dff_B_KUFfFuAc8_2;
	wire w_dff_B_Mqyjql5n2_2;
	wire w_dff_B_MEQp75cg1_2;
	wire w_dff_B_5ligMp879_2;
	wire w_dff_B_mnZcbAnD2_2;
	wire w_dff_B_roI7RvcF0_2;
	wire w_dff_B_SFQP6Lyz8_2;
	wire w_dff_B_4Ba7yUbC7_2;
	wire w_dff_B_gdbDDKO17_2;
	wire w_dff_B_xDY6n8gT4_2;
	wire w_dff_B_kAAMWXrC9_2;
	wire w_dff_B_fe0Sx0cY3_2;
	wire w_dff_B_vVmjT4eL4_2;
	wire w_dff_B_UgcHleqv1_2;
	wire w_dff_B_4yxHmEsr7_2;
	wire w_dff_B_MO9xv4sd5_2;
	wire w_dff_B_FdfsJ2bu9_2;
	wire w_dff_B_KJgi9yBS9_2;
	wire w_dff_B_MmSVDjU50_2;
	wire w_dff_B_M7PjRRpN6_2;
	wire w_dff_B_2x6iD6hl6_2;
	wire w_dff_B_p3ZNSoEw1_2;
	wire w_dff_B_1ax3ECta3_0;
	wire w_dff_A_PxH1NRvU1_1;
	wire w_dff_B_1aMAG6Sh9_1;
	wire w_dff_B_inRuTdfA4_2;
	wire w_dff_B_AlyN7p6I0_2;
	wire w_dff_B_zAGxqyxT5_2;
	wire w_dff_B_wFlugMFi4_2;
	wire w_dff_B_TxlXRj5I9_2;
	wire w_dff_B_icdHhhTo6_2;
	wire w_dff_B_xi53Znlx0_2;
	wire w_dff_B_f7way87Z8_2;
	wire w_dff_B_WbFIrWsJ2_2;
	wire w_dff_B_A8ztJC4t9_2;
	wire w_dff_B_OyhKT9HT2_2;
	wire w_dff_B_MGtDrr1s5_2;
	wire w_dff_B_3YmYvg2T6_2;
	wire w_dff_B_fbiqLisC1_2;
	wire w_dff_B_6uFlHUwT1_2;
	wire w_dff_B_fwn4TuNY9_2;
	wire w_dff_B_d3Nai7tk8_2;
	wire w_dff_B_UJVtCxeN7_2;
	wire w_dff_B_FcJZjd6i2_2;
	wire w_dff_B_nMCAX8wY4_2;
	wire w_dff_B_tAKjTtwH1_2;
	wire w_dff_B_oAtIciFs5_2;
	wire w_dff_B_mmY24BI05_2;
	wire w_dff_B_GzKuMRKi2_2;
	wire w_dff_B_X82b9LiP9_2;
	wire w_dff_B_7bkMfmwt4_2;
	wire w_dff_B_qnyTeGld3_2;
	wire w_dff_B_qGC9KhU82_2;
	wire w_dff_B_ZvnobH0V6_2;
	wire w_dff_B_zZ9onDR59_2;
	wire w_dff_B_2Elc3VTP4_2;
	wire w_dff_B_xTZTmmn96_2;
	wire w_dff_B_v4KQNg9H3_2;
	wire w_dff_B_315ukMqs3_2;
	wire w_dff_B_I3NbLvJY0_2;
	wire w_dff_B_5QTuLfKd5_2;
	wire w_dff_B_r9hSc30U2_2;
	wire w_dff_B_y4IGddwb1_2;
	wire w_dff_B_ElXZYIa20_2;
	wire w_dff_B_M3LK1xzU2_2;
	wire w_dff_B_IbvucGwe3_2;
	wire w_dff_B_9qHtF55P1_2;
	wire w_dff_B_lZcZVzdw3_1;
	wire w_dff_B_XPhmulcQ5_2;
	wire w_dff_B_ODZG99Yp7_2;
	wire w_dff_B_bf3OVSsi8_2;
	wire w_dff_B_iqTgUew23_2;
	wire w_dff_B_m4v3d7Kv1_2;
	wire w_dff_B_neuP4lQ52_2;
	wire w_dff_B_TSUrgaKt8_2;
	wire w_dff_B_wD8Zr9vW6_2;
	wire w_dff_B_7Yfwf9aZ7_2;
	wire w_dff_B_RsgfZ2uu3_2;
	wire w_dff_B_K1KFsQ2u2_2;
	wire w_dff_B_i2KxM8Re5_2;
	wire w_dff_B_OlTIx4ce8_2;
	wire w_dff_B_mlj6Hy8p2_2;
	wire w_dff_B_OgCIYfPB8_2;
	wire w_dff_B_SnhMdyTp7_2;
	wire w_dff_B_cwGQd2xI4_2;
	wire w_dff_B_A9IIPvHv3_2;
	wire w_dff_B_4kjnqb1K6_2;
	wire w_dff_B_YZT9ddvX4_2;
	wire w_dff_B_JwZKP0fX2_2;
	wire w_dff_B_1CIVLKIj4_2;
	wire w_dff_B_Ld4rCjnd4_2;
	wire w_dff_B_kRSEWkmn0_2;
	wire w_dff_B_pepnupah9_2;
	wire w_dff_B_FOHMAXDs5_2;
	wire w_dff_B_Z74a6RK19_2;
	wire w_dff_B_J5YehL8a8_2;
	wire w_dff_B_yUuoIbTx8_2;
	wire w_dff_B_EvBpFlVv7_2;
	wire w_dff_B_JP0xAU0r3_2;
	wire w_dff_B_3FVv3jQY6_2;
	wire w_dff_B_pExHhlD19_2;
	wire w_dff_B_YVSvoF7J7_2;
	wire w_dff_B_WQ1WoQPh9_2;
	wire w_dff_B_0fI18B7O1_2;
	wire w_dff_B_GKDcWaz37_2;
	wire w_dff_B_Rp3ucYYc1_2;
	wire w_dff_B_MCd6ORrO0_2;
	wire w_dff_B_htxOHOD62_1;
	wire w_dff_B_1kv8LCsj3_2;
	wire w_dff_B_JcQK66OL1_2;
	wire w_dff_B_uaUhpf4s7_2;
	wire w_dff_B_G47l6X8V8_2;
	wire w_dff_B_Ro9KydpO7_2;
	wire w_dff_B_9SuPu77z6_2;
	wire w_dff_B_WrNEXcKN9_2;
	wire w_dff_B_43XMRe7j9_2;
	wire w_dff_B_s2cgr2AW3_2;
	wire w_dff_B_Ozkoba9W8_2;
	wire w_dff_B_yXxqEg2W1_2;
	wire w_dff_B_OAtSuQRO1_2;
	wire w_dff_B_mcp0dSs15_2;
	wire w_dff_B_6A6qlhvf4_2;
	wire w_dff_B_TnKfDes99_2;
	wire w_dff_B_cKDrpWUJ7_2;
	wire w_dff_B_vrDEH52I1_2;
	wire w_dff_B_0xICeWWk8_2;
	wire w_dff_B_2q53ClOO1_2;
	wire w_dff_B_Yk0RwQoZ2_2;
	wire w_dff_B_7HWmukWz4_2;
	wire w_dff_B_vskxeJnm5_2;
	wire w_dff_B_GliYpxA19_2;
	wire w_dff_B_ZcvSGS8T6_2;
	wire w_dff_B_mzHnQgh06_2;
	wire w_dff_B_iFYc1Zr22_2;
	wire w_dff_B_lFIs85bo3_2;
	wire w_dff_B_vRhkfnEJ5_2;
	wire w_dff_B_wle64HD04_2;
	wire w_dff_B_LybolC2y0_2;
	wire w_dff_B_Efvx2P9U3_2;
	wire w_dff_B_7J8XEpEw9_2;
	wire w_dff_B_cl5b4eIb2_2;
	wire w_dff_B_UnKdesTB9_2;
	wire w_dff_B_PCF5qNEU6_2;
	wire w_dff_B_JVkXs9h96_2;
	wire w_dff_B_rlehoPlh3_1;
	wire w_dff_B_qnRqOOAO4_2;
	wire w_dff_B_ZqoxD9Vg7_2;
	wire w_dff_B_xDle3Ej36_2;
	wire w_dff_B_AKAHyaMk5_2;
	wire w_dff_B_2mk9SXaj9_2;
	wire w_dff_B_Oa14ZuAL2_2;
	wire w_dff_B_r7CK5K8f0_2;
	wire w_dff_B_TP682LfF3_2;
	wire w_dff_B_t5S7MITs9_2;
	wire w_dff_B_8nU81K8n7_2;
	wire w_dff_B_T3GpPOQY2_2;
	wire w_dff_B_eF3Gpsp35_2;
	wire w_dff_B_ddrW5dNN3_2;
	wire w_dff_B_w4xr85qT5_2;
	wire w_dff_B_8pU5VBtd7_2;
	wire w_dff_B_GH8vwDxA0_2;
	wire w_dff_B_eKVAcyeV2_2;
	wire w_dff_B_mB3RxjI36_2;
	wire w_dff_B_CkRzwcqN2_2;
	wire w_dff_B_Pbp7yQOZ7_2;
	wire w_dff_B_NyT20UKI5_2;
	wire w_dff_B_3gwCqjJ39_2;
	wire w_dff_B_glm0SnPP8_2;
	wire w_dff_B_pti3UzU40_2;
	wire w_dff_B_FoFBl5Dz0_2;
	wire w_dff_B_yWvJUjzJ6_2;
	wire w_dff_B_SZlvdsNo7_2;
	wire w_dff_B_oDJxQXXZ3_2;
	wire w_dff_B_2lamB7ID9_2;
	wire w_dff_B_aggaVBfl3_2;
	wire w_dff_B_0vKqDatN5_2;
	wire w_dff_B_kuIpC0Vp4_2;
	wire w_dff_B_D3YZD5D76_2;
	wire w_dff_B_gg2FB3My6_1;
	wire w_dff_B_AnYtJzmb0_2;
	wire w_dff_B_CnCUs4fP3_2;
	wire w_dff_B_OE7PKV5v8_2;
	wire w_dff_B_boDm4h6Q6_2;
	wire w_dff_B_Cu9evJKv3_2;
	wire w_dff_B_KAXUlKk72_2;
	wire w_dff_B_SSStPbcG2_2;
	wire w_dff_B_H4pIjNWc0_2;
	wire w_dff_B_qtWiRgLX7_2;
	wire w_dff_B_tpxzfHba9_2;
	wire w_dff_B_LAEe8wqC0_2;
	wire w_dff_B_330shDWv3_2;
	wire w_dff_B_9DurIZci1_2;
	wire w_dff_B_BvuxMaUr8_2;
	wire w_dff_B_UrosZfpO2_2;
	wire w_dff_B_UKZvIUwg3_2;
	wire w_dff_B_wJxyiGT27_2;
	wire w_dff_B_5BjBczeA7_2;
	wire w_dff_B_5CNKYy1E9_2;
	wire w_dff_B_8b3QJ5jh9_2;
	wire w_dff_B_QckKYNf06_2;
	wire w_dff_B_cwz65iGh5_2;
	wire w_dff_B_wY0IsHG82_2;
	wire w_dff_B_klWKGcQv2_2;
	wire w_dff_B_3IaUNx172_2;
	wire w_dff_B_lEHS7Zak6_2;
	wire w_dff_B_K6D321cK1_2;
	wire w_dff_B_tYEhZjTJ3_2;
	wire w_dff_B_0et19v5d5_2;
	wire w_dff_B_SmpoGJ4N8_2;
	wire w_dff_B_7bnw41xC0_1;
	wire w_dff_B_p5YvcBGO7_2;
	wire w_dff_B_wSOusyKg6_2;
	wire w_dff_B_3vt0DaiS8_2;
	wire w_dff_B_wEcy0GZO6_2;
	wire w_dff_B_z4G4z7R83_2;
	wire w_dff_B_uUr8EfHm2_2;
	wire w_dff_B_TbXRX6eS1_2;
	wire w_dff_B_YmavrFzT1_2;
	wire w_dff_B_4bn01ozy2_2;
	wire w_dff_B_Ge5Cc4Kl6_2;
	wire w_dff_B_PimQafJy6_2;
	wire w_dff_B_ZEMII0Zt4_2;
	wire w_dff_B_DWDa9spu8_2;
	wire w_dff_B_voH1uFbB5_2;
	wire w_dff_B_d1tQvrDw6_2;
	wire w_dff_B_R0ygIqUD6_2;
	wire w_dff_B_U1dqrdTD5_2;
	wire w_dff_B_CKkttcAN6_2;
	wire w_dff_B_KGLorfy53_2;
	wire w_dff_B_RBtOME0j2_2;
	wire w_dff_B_TL7zEP7a7_2;
	wire w_dff_B_pzJHSiQL5_2;
	wire w_dff_B_gWArFEau1_2;
	wire w_dff_B_QtAs6B3W4_2;
	wire w_dff_B_PGbTllZq5_2;
	wire w_dff_B_ZaSiZtFw1_2;
	wire w_dff_B_hYJzon4O3_2;
	wire w_dff_B_OnoqUXsn8_1;
	wire w_dff_B_KefcasIe6_2;
	wire w_dff_B_HzG04r9G3_2;
	wire w_dff_B_fHjGnlhj5_2;
	wire w_dff_B_s6yqWXg95_2;
	wire w_dff_B_n1zXIAZP7_2;
	wire w_dff_B_yV6xjVtf5_2;
	wire w_dff_B_B7lOt4jv7_2;
	wire w_dff_B_htayxL4J3_2;
	wire w_dff_B_UpNnZp7M1_2;
	wire w_dff_B_hRxavixN3_2;
	wire w_dff_B_8VSF4nkX0_2;
	wire w_dff_B_Y3A3szwY8_2;
	wire w_dff_B_NRvHbfiu7_2;
	wire w_dff_B_Yp43ncj11_2;
	wire w_dff_B_mOXjGl9Q4_2;
	wire w_dff_B_Ik7mrRdj5_2;
	wire w_dff_B_yO9TkDke5_2;
	wire w_dff_B_MvEKXKAS1_2;
	wire w_dff_B_gYJCljrR4_2;
	wire w_dff_B_za8iUesw8_2;
	wire w_dff_B_u2NwlTMH0_2;
	wire w_dff_B_6Ah8I60j5_2;
	wire w_dff_B_cKWKrVXj8_2;
	wire w_dff_B_V85fjSlv9_2;
	wire w_dff_B_rB1nKRZA0_1;
	wire w_dff_B_B7KRyNZu6_2;
	wire w_dff_B_HMuKd9D11_2;
	wire w_dff_B_miT1FUoR1_2;
	wire w_dff_B_yMvNDoDM5_2;
	wire w_dff_B_sbJNVXe81_2;
	wire w_dff_B_eI9W4oGE3_2;
	wire w_dff_B_B8ee8iVP2_2;
	wire w_dff_B_PevLuJYF7_2;
	wire w_dff_B_5w3Av6GE3_2;
	wire w_dff_B_p0PG2wGQ8_2;
	wire w_dff_B_M8nokPFC0_2;
	wire w_dff_B_WZnKADMq0_2;
	wire w_dff_B_AZvMrFNO5_2;
	wire w_dff_B_xy8eEO6j9_2;
	wire w_dff_B_bMmjzMxZ7_2;
	wire w_dff_B_OerqAZ2r4_2;
	wire w_dff_B_jPKYSNFo1_2;
	wire w_dff_B_388w2Zga0_2;
	wire w_dff_B_kpIfSQFC1_2;
	wire w_dff_B_VA0c2Vd83_2;
	wire w_dff_B_iedO2Yhv8_2;
	wire w_dff_B_SLuxqxfn3_1;
	wire w_dff_B_3TAhVC4f7_2;
	wire w_dff_B_w3Yl70fm8_2;
	wire w_dff_B_L8n5hhGj3_2;
	wire w_dff_B_huCo1aGm2_2;
	wire w_dff_B_eoxFidYA3_2;
	wire w_dff_B_UZxZduZX0_2;
	wire w_dff_B_kOKqo6Ms2_2;
	wire w_dff_B_Rz7r1ZiV0_2;
	wire w_dff_B_xoXXaG8G1_2;
	wire w_dff_B_okcYbJYB4_2;
	wire w_dff_B_fsoFwImI9_2;
	wire w_dff_B_bYvR40qM9_2;
	wire w_dff_B_IjvRux7i0_2;
	wire w_dff_B_rBo1blwq5_2;
	wire w_dff_B_d9KG1JPN5_2;
	wire w_dff_B_lRAeVbAg5_2;
	wire w_dff_B_1d86I5RD5_2;
	wire w_dff_B_1w0Q7Pzv5_2;
	wire w_dff_B_9p2hFyFV9_1;
	wire w_dff_B_YSEJDdHr8_2;
	wire w_dff_B_7QtlJNFC1_2;
	wire w_dff_B_fecmAZju2_2;
	wire w_dff_B_T8h6c7c27_2;
	wire w_dff_B_o93ULIuq9_2;
	wire w_dff_B_ZTAuuj942_2;
	wire w_dff_B_ZR2rgU1e0_2;
	wire w_dff_B_wXvfAy4a7_2;
	wire w_dff_B_lkhQmSBd0_2;
	wire w_dff_B_E9KrE9Jw9_2;
	wire w_dff_B_T3444ETd4_2;
	wire w_dff_B_FMTujS1d9_2;
	wire w_dff_B_P8mzXKyo4_2;
	wire w_dff_B_yETXfUWg6_2;
	wire w_dff_B_Kuevk1gs9_2;
	wire w_dff_B_IdxXSTVP0_1;
	wire w_dff_B_Jdk1nkM12_2;
	wire w_dff_B_9bO056u13_2;
	wire w_dff_B_bmpZvaVQ5_2;
	wire w_dff_B_5yISK2Gy2_2;
	wire w_dff_B_REIWgtRT8_2;
	wire w_dff_B_NjLmuidY2_2;
	wire w_dff_B_IBGigjUL9_2;
	wire w_dff_B_2KEe7e9F6_2;
	wire w_dff_B_ELg0OH7J0_2;
	wire w_dff_B_qVefu5aa2_2;
	wire w_dff_B_dTMigAAZ6_2;
	wire w_dff_B_p2ZwLPy27_2;
	wire w_dff_B_4uHK7tHT0_1;
	wire w_dff_B_6jM7pCO53_2;
	wire w_dff_B_29AIBOeG6_2;
	wire w_dff_B_8jVsIgq90_2;
	wire w_dff_B_79Va2LeQ9_2;
	wire w_dff_B_4Jefg1ts2_2;
	wire w_dff_B_f97bKrLE2_2;
	wire w_dff_B_UNGCasGX6_2;
	wire w_dff_B_CuSaWmlk0_2;
	wire w_dff_B_KCgyCyz10_2;
	wire w_dff_B_4ORAqMPa0_2;
	wire w_dff_B_zrQ40S7o4_2;
	wire w_dff_B_XEg0eNsw0_1;
	wire w_dff_B_7jFsosD90_1;
	wire w_dff_B_APjeyntA5_2;
	wire w_dff_B_VzrCsoqi0_2;
	wire w_dff_B_a8u7jpK85_2;
	wire w_dff_B_PJsyqXJB2_0;
	wire w_dff_A_4mp05Umi5_0;
	wire w_dff_A_ErpNfXoR8_0;
	wire w_dff_A_4pv54OEY1_1;
	wire w_dff_A_dAKuKW9I4_1;
	wire w_dff_B_oYhPHKjl4_1;
	wire w_dff_B_2iX1qkJR9_2;
	wire w_dff_B_iPUBaDTI8_2;
	wire w_dff_B_kvLTVt0Z9_2;
	wire w_dff_B_4htIGfre7_2;
	wire w_dff_B_nd5vT7jX8_2;
	wire w_dff_B_rXjVEhCa5_2;
	wire w_dff_B_DkGFepT26_2;
	wire w_dff_B_BfvZLibs9_2;
	wire w_dff_B_zoPKMN4e8_2;
	wire w_dff_B_lJY29jr69_2;
	wire w_dff_B_ZYqT0wRN2_2;
	wire w_dff_B_n4tp6VBk4_2;
	wire w_dff_B_AAZ0HZk78_2;
	wire w_dff_B_jUZyEqdB8_2;
	wire w_dff_B_th0klIpv7_2;
	wire w_dff_B_76Gh53Sf5_2;
	wire w_dff_B_Z2dBzG2a3_2;
	wire w_dff_B_0qQCfqbM7_2;
	wire w_dff_B_3FCms8IU6_2;
	wire w_dff_B_ddgBhsn63_2;
	wire w_dff_B_Wn0haHJ42_2;
	wire w_dff_B_Qu2HyoT23_2;
	wire w_dff_B_kSgfh2fp8_2;
	wire w_dff_B_PSZTaUdt7_2;
	wire w_dff_B_nGPZtgZs5_2;
	wire w_dff_B_RZYqVgc03_2;
	wire w_dff_B_3MKWqkmm5_2;
	wire w_dff_B_Q3Z7tuAa4_2;
	wire w_dff_B_qRBu20oN3_2;
	wire w_dff_B_F6YZlYos5_2;
	wire w_dff_B_7MbxxquT9_2;
	wire w_dff_B_b2tvfak68_2;
	wire w_dff_B_2rWbq4s89_2;
	wire w_dff_B_aQIXke7N9_2;
	wire w_dff_B_isxosnJW5_2;
	wire w_dff_B_mnqzB8ou4_2;
	wire w_dff_B_aWtXyjR17_2;
	wire w_dff_B_2U4AEvCd8_2;
	wire w_dff_B_py8EmL695_2;
	wire w_dff_B_gHiaeyQm2_2;
	wire w_dff_B_r96ggMCF1_2;
	wire w_dff_B_bdbI5LpD7_2;
	wire w_dff_B_o10tMNDT3_2;
	wire w_dff_B_8FEdDFRe5_2;
	wire w_dff_B_XM4ocCmk3_2;
	wire w_dff_B_jZxX9Yif1_2;
	wire w_dff_B_BVI7x5lT3_0;
	wire w_dff_A_ZZHp1yH95_1;
	wire w_dff_B_zsNagZtx2_1;
	wire w_dff_B_KQN9dBK23_2;
	wire w_dff_B_eURYiopo0_2;
	wire w_dff_B_ccThDRwu2_2;
	wire w_dff_B_MA36lqUx7_2;
	wire w_dff_B_Oqy4fChH6_2;
	wire w_dff_B_ipOgdIF81_2;
	wire w_dff_B_HonmLwBS7_2;
	wire w_dff_B_KCJ4womP2_2;
	wire w_dff_B_tjDW81ES4_2;
	wire w_dff_B_7wyXYK1F8_2;
	wire w_dff_B_EMR9cLy91_2;
	wire w_dff_B_h9sf2DD17_2;
	wire w_dff_B_1QPeJpFK7_2;
	wire w_dff_B_HRpebVMQ4_2;
	wire w_dff_B_Vjz80nv38_2;
	wire w_dff_B_VwtcjlgE8_2;
	wire w_dff_B_8p9TZ9WH7_2;
	wire w_dff_B_GUQdrqMZ4_2;
	wire w_dff_B_dRuvbDyk6_2;
	wire w_dff_B_8izDSxvv1_2;
	wire w_dff_B_vW27K4gl9_2;
	wire w_dff_B_c8f8wfBy5_2;
	wire w_dff_B_akFMc7ZY1_2;
	wire w_dff_B_nVeiDsEe8_2;
	wire w_dff_B_SBu6N85x7_2;
	wire w_dff_B_BRxuSeMW6_2;
	wire w_dff_B_V2KEJ7W12_2;
	wire w_dff_B_7tv8BPpL8_2;
	wire w_dff_B_2WkUKoCC5_2;
	wire w_dff_B_kNuoio7N7_2;
	wire w_dff_B_PRzlvdY87_2;
	wire w_dff_B_SVSYuJBJ3_2;
	wire w_dff_B_jKfmhyGq3_2;
	wire w_dff_B_7itRnMKc8_2;
	wire w_dff_B_ZMHvjRCv7_2;
	wire w_dff_B_PcpCVi0w7_2;
	wire w_dff_B_XF04V13S3_2;
	wire w_dff_B_fQ5bDZ6e1_2;
	wire w_dff_B_MWkULhKK5_2;
	wire w_dff_B_yDVmqgXH7_2;
	wire w_dff_B_qRHni46W2_2;
	wire w_dff_B_FLkG0m4S9_2;
	wire w_dff_B_jJuYpWOA2_1;
	wire w_dff_B_5MebQy4y3_2;
	wire w_dff_B_tyil62C34_2;
	wire w_dff_B_wgyVInjP7_2;
	wire w_dff_B_EI2UErS63_2;
	wire w_dff_B_GaCBY2Zp1_2;
	wire w_dff_B_JShO2dtC3_2;
	wire w_dff_B_19s6xN4c4_2;
	wire w_dff_B_Tcm7HXuR9_2;
	wire w_dff_B_gfMISfdO3_2;
	wire w_dff_B_8DVVGD8C6_2;
	wire w_dff_B_Ff1yS4UM3_2;
	wire w_dff_B_wUmCV5oz1_2;
	wire w_dff_B_uLafZMRB4_2;
	wire w_dff_B_yo6FGxEx2_2;
	wire w_dff_B_utpluYEb2_2;
	wire w_dff_B_2qKwkANa9_2;
	wire w_dff_B_3YeARK4s5_2;
	wire w_dff_B_rxn99gtp8_2;
	wire w_dff_B_I15Z2ViY3_2;
	wire w_dff_B_yJylDi858_2;
	wire w_dff_B_3nJajgoy7_2;
	wire w_dff_B_bqEsBQLj2_2;
	wire w_dff_B_WdLbnMT72_2;
	wire w_dff_B_vPDYpPKz5_2;
	wire w_dff_B_R5vCPNJl1_2;
	wire w_dff_B_Mh8hxsIz2_2;
	wire w_dff_B_RhJvNJP53_2;
	wire w_dff_B_HDt627Dx1_2;
	wire w_dff_B_qHekgAvu2_2;
	wire w_dff_B_0CAk07Ti4_2;
	wire w_dff_B_t0QCoj4S8_2;
	wire w_dff_B_rdBYLdR77_2;
	wire w_dff_B_hASYa8Ly5_2;
	wire w_dff_B_fthatEhs0_2;
	wire w_dff_B_YcsuVGtl3_2;
	wire w_dff_B_c7dTpPDR9_2;
	wire w_dff_B_GZUGlUZm7_2;
	wire w_dff_B_o7k5VhFC6_2;
	wire w_dff_B_3LZA2KGF3_2;
	wire w_dff_B_mI1SzJPV7_1;
	wire w_dff_B_MS5RgPOK3_2;
	wire w_dff_B_qvjMcSCF3_2;
	wire w_dff_B_pAfmfhW22_2;
	wire w_dff_B_3ArIR8xx7_2;
	wire w_dff_B_4jukcp5a0_2;
	wire w_dff_B_xkjF5DsQ3_2;
	wire w_dff_B_nmFDYMGB6_2;
	wire w_dff_B_kdyF9wor8_2;
	wire w_dff_B_IjgkynGZ4_2;
	wire w_dff_B_ThGcIjRc9_2;
	wire w_dff_B_BjQXxbml7_2;
	wire w_dff_B_fN3cWTD72_2;
	wire w_dff_B_GlbVVF2m8_2;
	wire w_dff_B_KJzueAyN5_2;
	wire w_dff_B_UI78CJEv9_2;
	wire w_dff_B_XE56vBG73_2;
	wire w_dff_B_mDgqSqOO8_2;
	wire w_dff_B_bivT0ACb9_2;
	wire w_dff_B_ETGiKMWk9_2;
	wire w_dff_B_IgeJkEo30_2;
	wire w_dff_B_XEYGXgFd2_2;
	wire w_dff_B_0qo0iBGN2_2;
	wire w_dff_B_VbUsVrxV3_2;
	wire w_dff_B_00pExPWt1_2;
	wire w_dff_B_6cjjXCw71_2;
	wire w_dff_B_ZLEaQRx80_2;
	wire w_dff_B_VSx8nG8j7_2;
	wire w_dff_B_K4o352yn0_2;
	wire w_dff_B_4Bk24P1w5_2;
	wire w_dff_B_5awZzLdr3_2;
	wire w_dff_B_Bb8W7eVh7_2;
	wire w_dff_B_hDCKSB4k2_2;
	wire w_dff_B_GIw7g1rw3_2;
	wire w_dff_B_6q6Jk2e22_2;
	wire w_dff_B_l85Ij3Ye7_2;
	wire w_dff_B_Js1sOPgh7_2;
	wire w_dff_B_LbZi72ql7_1;
	wire w_dff_B_YD1atmkx4_2;
	wire w_dff_B_L9fRZkbE5_2;
	wire w_dff_B_IJfShoji8_2;
	wire w_dff_B_udOBCeIp6_2;
	wire w_dff_B_3A8ESZVg6_2;
	wire w_dff_B_fJ7DtA105_2;
	wire w_dff_B_5ZboEowH5_2;
	wire w_dff_B_zZyq1RD10_2;
	wire w_dff_B_QTtbc1qE5_2;
	wire w_dff_B_iBCncV6B3_2;
	wire w_dff_B_zYn8Ogo56_2;
	wire w_dff_B_wAP5mkC67_2;
	wire w_dff_B_4N4eDkzd6_2;
	wire w_dff_B_gy8SRj9I6_2;
	wire w_dff_B_hAVVkfDr8_2;
	wire w_dff_B_ZMha1dJU1_2;
	wire w_dff_B_n4xlXqnW0_2;
	wire w_dff_B_ozvO78aK6_2;
	wire w_dff_B_Z3pIL7yF1_2;
	wire w_dff_B_ncMAgAVV0_2;
	wire w_dff_B_GK5mYZBb3_2;
	wire w_dff_B_9L7cTObu3_2;
	wire w_dff_B_3ufLWbKX6_2;
	wire w_dff_B_uEG9OSjB3_2;
	wire w_dff_B_cRTjQz4a7_2;
	wire w_dff_B_SKMJ9imk3_2;
	wire w_dff_B_JJQPVFb56_2;
	wire w_dff_B_FGseNpCy1_2;
	wire w_dff_B_kVwVwxbL3_2;
	wire w_dff_B_I1W31Ccg7_2;
	wire w_dff_B_7q09bgBt4_2;
	wire w_dff_B_okKF1GY07_2;
	wire w_dff_B_6HhSHxWD4_2;
	wire w_dff_B_zIUS8s871_1;
	wire w_dff_B_NGDpqiWM6_2;
	wire w_dff_B_bJa4WDH61_2;
	wire w_dff_B_qaCn5nbH5_2;
	wire w_dff_B_HlsJiCPB2_2;
	wire w_dff_B_lY9gyQlw8_2;
	wire w_dff_B_8bHfZIRA7_2;
	wire w_dff_B_qanxPJZu4_2;
	wire w_dff_B_VG7ja1FN1_2;
	wire w_dff_B_krFEi6Am1_2;
	wire w_dff_B_yKbQhQDw4_2;
	wire w_dff_B_Hqvy0AWD3_2;
	wire w_dff_B_frCnMz7W3_2;
	wire w_dff_B_4iLs0C436_2;
	wire w_dff_B_CA29PapU9_2;
	wire w_dff_B_nNKIWlm17_2;
	wire w_dff_B_VkPwFpIc6_2;
	wire w_dff_B_ODiWUEgl9_2;
	wire w_dff_B_1ZayYYam8_2;
	wire w_dff_B_ftGECzqr9_2;
	wire w_dff_B_cuXEpZpm1_2;
	wire w_dff_B_XvSGN2c00_2;
	wire w_dff_B_jTdHultr4_2;
	wire w_dff_B_0ACKFj0z7_2;
	wire w_dff_B_hyn5HOFb7_2;
	wire w_dff_B_LIatZtMR5_2;
	wire w_dff_B_HSx2JnHT2_2;
	wire w_dff_B_6HZ8KgQp6_2;
	wire w_dff_B_DXGNdAQd6_2;
	wire w_dff_B_WHme5axn2_2;
	wire w_dff_B_8UoqdxrN9_2;
	wire w_dff_B_qGgjE1Rn5_1;
	wire w_dff_B_J6vRyHIx5_2;
	wire w_dff_B_LeAaHmsT5_2;
	wire w_dff_B_9ANxlNdu9_2;
	wire w_dff_B_OhayqCGm0_2;
	wire w_dff_B_WbQT8W073_2;
	wire w_dff_B_Kcb3axph0_2;
	wire w_dff_B_vEinAjQ44_2;
	wire w_dff_B_sNcA8fvc9_2;
	wire w_dff_B_G1W2vT0s2_2;
	wire w_dff_B_IYklaDxc3_2;
	wire w_dff_B_ySVQXHtq3_2;
	wire w_dff_B_edYN6leQ4_2;
	wire w_dff_B_zlpNHW0z1_2;
	wire w_dff_B_e1nUaIqS3_2;
	wire w_dff_B_cWzcx7Zj3_2;
	wire w_dff_B_o5Ssbzgm4_2;
	wire w_dff_B_ccHIVRvk7_2;
	wire w_dff_B_zsCqAjJ61_2;
	wire w_dff_B_1wUjJCab7_2;
	wire w_dff_B_ZoewvTH74_2;
	wire w_dff_B_6kQtoUCL0_2;
	wire w_dff_B_sswBTdAv5_2;
	wire w_dff_B_RijX5t8b1_2;
	wire w_dff_B_htjO9n1L6_2;
	wire w_dff_B_rPKIXgGq9_2;
	wire w_dff_B_CSNfWwZN2_2;
	wire w_dff_B_pravOeJa6_2;
	wire w_dff_B_NUJAPVTH1_1;
	wire w_dff_B_zRSG50vb3_2;
	wire w_dff_B_LdNbmbpL6_2;
	wire w_dff_B_eyJX0G1q9_2;
	wire w_dff_B_gSZYEKnZ8_2;
	wire w_dff_B_rtbX6WwV7_2;
	wire w_dff_B_G8fcrtJZ6_2;
	wire w_dff_B_kel6czC82_2;
	wire w_dff_B_wiPHTbKD7_2;
	wire w_dff_B_kWIfkf4A4_2;
	wire w_dff_B_QOdgpeCl9_2;
	wire w_dff_B_Z1pTSHl80_2;
	wire w_dff_B_M6u4jiNH0_2;
	wire w_dff_B_Uokl5F1z8_2;
	wire w_dff_B_DCjcOa3G1_2;
	wire w_dff_B_CmtaG9eP2_2;
	wire w_dff_B_R6a7cuxy8_2;
	wire w_dff_B_2dLhHX765_2;
	wire w_dff_B_M9dEtoLm5_2;
	wire w_dff_B_6vzcQcFf2_2;
	wire w_dff_B_nIqNbTDI6_2;
	wire w_dff_B_6gGDwck35_2;
	wire w_dff_B_iCMIOgkW8_2;
	wire w_dff_B_2WUixItf6_2;
	wire w_dff_B_EqvHgSLD6_2;
	wire w_dff_B_SY1dVtdg4_1;
	wire w_dff_B_fdLQXVQC8_2;
	wire w_dff_B_750sclDP4_2;
	wire w_dff_B_HYuka2wO9_2;
	wire w_dff_B_X6yIsHbD5_2;
	wire w_dff_B_19xtU5IV1_2;
	wire w_dff_B_KgMNJRlv7_2;
	wire w_dff_B_EXM3HdVp7_2;
	wire w_dff_B_QALLJNme5_2;
	wire w_dff_B_gNGT0SeE9_2;
	wire w_dff_B_lxa6Uaao8_2;
	wire w_dff_B_DoJYQiuo5_2;
	wire w_dff_B_4jkqOUvD3_2;
	wire w_dff_B_Y2u2Mk3D1_2;
	wire w_dff_B_xiZ4gCn92_2;
	wire w_dff_B_5q2KSaA64_2;
	wire w_dff_B_Uk2waCTi9_2;
	wire w_dff_B_YuRtDOMr4_2;
	wire w_dff_B_2FmEnAqX6_2;
	wire w_dff_B_qKnUK94u4_2;
	wire w_dff_B_xWjgITBo3_2;
	wire w_dff_B_YkoF4SCv4_2;
	wire w_dff_B_2GiWZanX5_1;
	wire w_dff_B_72qZHXs54_2;
	wire w_dff_B_aRivU5J29_2;
	wire w_dff_B_NfatX3m43_2;
	wire w_dff_B_aYOv1SLd6_2;
	wire w_dff_B_8aJc6ERt4_2;
	wire w_dff_B_7O0Zkyjx4_2;
	wire w_dff_B_Azy82fwj0_2;
	wire w_dff_B_gAWDaJPw5_2;
	wire w_dff_B_DXuin0ol9_2;
	wire w_dff_B_JZwvDQVf1_2;
	wire w_dff_B_TnlsbTit6_2;
	wire w_dff_B_57tzlzMX0_2;
	wire w_dff_B_Lvy2Z4Vx3_2;
	wire w_dff_B_LnA1wPUW8_2;
	wire w_dff_B_SbImryn38_2;
	wire w_dff_B_la7O5Nqs2_2;
	wire w_dff_B_28pqL9by1_2;
	wire w_dff_B_cF7Ixm6x1_2;
	wire w_dff_B_r9B0w8l35_1;
	wire w_dff_B_ZEwr4JXt5_2;
	wire w_dff_B_MesALP467_2;
	wire w_dff_B_UifpdZWV3_2;
	wire w_dff_B_M8txeVwG6_2;
	wire w_dff_B_oSMyBzXP0_2;
	wire w_dff_B_XBkNE5nj7_2;
	wire w_dff_B_mnpElBUh1_2;
	wire w_dff_B_7xLQkOa40_2;
	wire w_dff_B_fiMxtoMP6_2;
	wire w_dff_B_pCmurpbL1_2;
	wire w_dff_B_rYaauK352_2;
	wire w_dff_B_L9SLDhoh9_2;
	wire w_dff_B_u9nCgL5q5_2;
	wire w_dff_B_yuiA1Rrp4_2;
	wire w_dff_B_d8eQmLZH6_2;
	wire w_dff_B_m2Jk00NH5_1;
	wire w_dff_B_1epBzvRe8_2;
	wire w_dff_B_0rgXNger8_2;
	wire w_dff_B_sivrI2256_2;
	wire w_dff_B_hRnZjd0z4_2;
	wire w_dff_B_7J0qZQea2_2;
	wire w_dff_B_7CdF4jer7_2;
	wire w_dff_B_XObOW2hW1_2;
	wire w_dff_B_jBAZemRm5_2;
	wire w_dff_B_dINjm7Ft0_2;
	wire w_dff_B_JCuDsFxD7_2;
	wire w_dff_B_Bw3OsVie8_2;
	wire w_dff_B_iknV8gPt0_2;
	wire w_dff_B_akOY61NU1_1;
	wire w_dff_B_HtscdnlW7_2;
	wire w_dff_B_dVFGlK9i2_2;
	wire w_dff_B_a6qujakw4_2;
	wire w_dff_B_kb1pdHTW2_2;
	wire w_dff_B_5YBzyBpb5_2;
	wire w_dff_B_HonZBjHB0_2;
	wire w_dff_B_a37YOQbf1_2;
	wire w_dff_B_sW1vra5Q7_2;
	wire w_dff_B_ct0g8B0Q6_2;
	wire w_dff_B_7EClZ9OK6_2;
	wire w_dff_B_bSzKJyA47_2;
	wire w_dff_B_IxrNAbwX9_1;
	wire w_dff_B_9kJ7FV726_1;
	wire w_dff_B_MIJfWOow1_2;
	wire w_dff_B_UcTY9fRj4_2;
	wire w_dff_B_QGJTPq0i6_2;
	wire w_dff_B_CBpFB20e9_0;
	wire w_dff_A_CigddwwK4_0;
	wire w_dff_A_PN5thRrM1_0;
	wire w_dff_A_dB2hOinj9_1;
	wire w_dff_A_iBKlWHFh0_1;
	wire w_dff_B_PRuDwE9Y3_2;
	wire w_dff_B_fQdaedm32_1;
	wire w_dff_B_To1rGYVT8_2;
	wire w_dff_B_gOnr7dGR8_2;
	wire w_dff_B_rPV06Wdr9_2;
	wire w_dff_B_4yiI2Aek3_2;
	wire w_dff_B_gRBa6ZD10_2;
	wire w_dff_B_2FswoSkg0_2;
	wire w_dff_B_bBDIiziW4_2;
	wire w_dff_B_mb1cISqR2_2;
	wire w_dff_B_wJjhnMvt3_2;
	wire w_dff_B_93Fd7zLP2_2;
	wire w_dff_B_Wt3wfxyq9_2;
	wire w_dff_B_eG1fY8XZ7_2;
	wire w_dff_B_pMYxWNMv7_2;
	wire w_dff_B_aktjuSIn8_2;
	wire w_dff_B_0QUl3x8T0_2;
	wire w_dff_B_xN17xPVe2_2;
	wire w_dff_B_oI0bT2ii7_2;
	wire w_dff_B_3Jg0OAzJ5_2;
	wire w_dff_B_sVdn2fhy7_2;
	wire w_dff_B_fVGi4qnx7_2;
	wire w_dff_B_AMkpMV9r8_2;
	wire w_dff_B_K4u83C0p8_2;
	wire w_dff_B_ltjsJ0Mk8_2;
	wire w_dff_B_9sfKQkEq8_2;
	wire w_dff_B_8vH6OZhe0_2;
	wire w_dff_B_utd7gkqZ0_2;
	wire w_dff_B_wtuzRUED7_2;
	wire w_dff_B_2Seqvs3J0_2;
	wire w_dff_B_vFSIWNtd6_2;
	wire w_dff_B_qB5EOR3P9_2;
	wire w_dff_B_2C8aICjN2_2;
	wire w_dff_B_3JP1qNqk0_2;
	wire w_dff_B_9mcI6qZF7_2;
	wire w_dff_B_ikMCDLfs7_2;
	wire w_dff_B_vHHCFOAW5_2;
	wire w_dff_B_c2TpOike2_2;
	wire w_dff_B_IjOpXgSA9_2;
	wire w_dff_B_CsWSkPJk0_2;
	wire w_dff_B_bkPas9l87_2;
	wire w_dff_B_N84NUNze8_2;
	wire w_dff_B_5oPFgi4G2_2;
	wire w_dff_B_SbvijqDi9_2;
	wire w_dff_B_L5qjy5tn6_2;
	wire w_dff_B_6U8373391_2;
	wire w_dff_B_RZlwdoMm0_2;
	wire w_dff_B_vPvA7ghK4_2;
	wire w_dff_B_7wdXn7xq8_1;
	wire w_dff_B_MBaxzcXn6_2;
	wire w_dff_B_ffOzgL0A6_2;
	wire w_dff_B_DcaIJKdj8_2;
	wire w_dff_B_aKsbO9YB1_2;
	wire w_dff_B_vPkuSM7D9_2;
	wire w_dff_B_ri8K1K2j6_2;
	wire w_dff_B_NpVHOysA0_2;
	wire w_dff_B_rEtLTi0k3_2;
	wire w_dff_B_vZWYy1ZJ9_2;
	wire w_dff_B_TYm4E5dt4_2;
	wire w_dff_B_IITNda7D9_2;
	wire w_dff_B_aM3CxAwF5_2;
	wire w_dff_B_O6XAyyGO9_2;
	wire w_dff_B_yE6j8YpU0_2;
	wire w_dff_B_pmHyXNkc7_2;
	wire w_dff_B_jlVxlsF33_2;
	wire w_dff_B_Pd09L2yh1_2;
	wire w_dff_B_OPMTPTxp3_2;
	wire w_dff_B_IPZr3kO27_2;
	wire w_dff_B_Yf6Wlj752_2;
	wire w_dff_B_gdHjwZcI1_2;
	wire w_dff_B_2Vg8P0ca2_2;
	wire w_dff_B_cI4J6ngt3_2;
	wire w_dff_B_RNepMO3g6_2;
	wire w_dff_B_qnbjfDLL2_2;
	wire w_dff_B_vxXFrN1R4_2;
	wire w_dff_B_qGy1li6f4_2;
	wire w_dff_B_ZD39w16C8_2;
	wire w_dff_B_1dRbeTai0_2;
	wire w_dff_B_sS4TXpeF5_2;
	wire w_dff_B_w4QzL81w7_2;
	wire w_dff_B_8mFOqBu00_2;
	wire w_dff_B_PEGDJIF03_2;
	wire w_dff_B_hzKbM6lj2_2;
	wire w_dff_B_RKk958mT8_2;
	wire w_dff_B_cSgU2YQR8_2;
	wire w_dff_B_k67nTlFJ0_2;
	wire w_dff_B_j5ssqJ709_2;
	wire w_dff_B_KBP1Yr8X1_2;
	wire w_dff_B_10j4VEk86_2;
	wire w_dff_B_HCrwfOX29_2;
	wire w_dff_B_W50Qyrbw6_2;
	wire w_dff_B_rlviRy9l5_1;
	wire w_dff_B_tt85ceTp2_2;
	wire w_dff_B_YB6HQslk7_2;
	wire w_dff_B_UgTW4v2B1_2;
	wire w_dff_B_9UWUFGRU4_2;
	wire w_dff_B_SP0FId8K8_2;
	wire w_dff_B_ECITgqmX1_2;
	wire w_dff_B_pcVGBoLR6_2;
	wire w_dff_B_T3niKc1M2_2;
	wire w_dff_B_jX6oBj0i5_2;
	wire w_dff_B_MvHgLRx49_2;
	wire w_dff_B_VjrxxHLG7_2;
	wire w_dff_B_b6P5lV8Y8_2;
	wire w_dff_B_lo1Jo8NM4_2;
	wire w_dff_B_C7ztNqX31_2;
	wire w_dff_B_clW06KAT5_2;
	wire w_dff_B_NCBxeYwQ8_2;
	wire w_dff_B_PIUXLQ7r0_2;
	wire w_dff_B_c9Oqtcda7_2;
	wire w_dff_B_fOv2905U6_2;
	wire w_dff_B_BWvCBIQi6_2;
	wire w_dff_B_uhwLdBhe2_2;
	wire w_dff_B_eQQ9BNKv2_2;
	wire w_dff_B_HjkYvuQO4_2;
	wire w_dff_B_TMtBTEPy5_2;
	wire w_dff_B_jZRa4nPc3_2;
	wire w_dff_B_ASirHnKY8_2;
	wire w_dff_B_6SjSxr2G1_2;
	wire w_dff_B_COsSvsm94_2;
	wire w_dff_B_AJBXZuQz9_2;
	wire w_dff_B_qQGAcyMx7_2;
	wire w_dff_B_v2AbIQqE3_2;
	wire w_dff_B_Ldk91WU46_2;
	wire w_dff_B_A7d9UWtF9_2;
	wire w_dff_B_rzsEWZXU3_2;
	wire w_dff_B_M07pNaUx9_2;
	wire w_dff_B_nkLIFtgr7_2;
	wire w_dff_B_jAmeWmgd8_2;
	wire w_dff_B_SlMs5Ypt1_2;
	wire w_dff_B_EbZ9Y5HW1_2;
	wire w_dff_B_O45oxs1m1_1;
	wire w_dff_B_GIt6yQGw5_2;
	wire w_dff_B_uBdElKpA7_2;
	wire w_dff_B_jglgimgk5_2;
	wire w_dff_B_HNNBXJ0e3_2;
	wire w_dff_B_EUv7Pd5x5_2;
	wire w_dff_B_atYAZREb3_2;
	wire w_dff_B_OklQO3ti5_2;
	wire w_dff_B_51586D049_2;
	wire w_dff_B_RX6Unpp46_2;
	wire w_dff_B_L6jxg9U82_2;
	wire w_dff_B_ZqpAp6zJ1_2;
	wire w_dff_B_1YWDwpIV6_2;
	wire w_dff_B_zc2ww7O23_2;
	wire w_dff_B_sf3Z0jfs3_2;
	wire w_dff_B_og8ipIzG0_2;
	wire w_dff_B_pbacs4S92_2;
	wire w_dff_B_eQsyoHpB9_2;
	wire w_dff_B_copNBME19_2;
	wire w_dff_B_0U5qMBne2_2;
	wire w_dff_B_hhX7s2Gr4_2;
	wire w_dff_B_dlyx0Y127_2;
	wire w_dff_B_Wh8mMQl34_2;
	wire w_dff_B_pXcWmqzX7_2;
	wire w_dff_B_gj9jYQON2_2;
	wire w_dff_B_MdM0X7Ni8_2;
	wire w_dff_B_xD3kKjUQ0_2;
	wire w_dff_B_8bU7kZIR7_2;
	wire w_dff_B_B9dGR5wu0_2;
	wire w_dff_B_YVsFPeV26_2;
	wire w_dff_B_BrYF22Up2_2;
	wire w_dff_B_s7WC25b94_2;
	wire w_dff_B_1jKFPvBD8_2;
	wire w_dff_B_q5B90cfv0_2;
	wire w_dff_B_WhphCp273_2;
	wire w_dff_B_aWErp4ZT3_2;
	wire w_dff_B_T1ZHVrvU9_2;
	wire w_dff_B_Q0KMD2eo2_1;
	wire w_dff_B_3LotTdUk0_2;
	wire w_dff_B_9WChpInF5_2;
	wire w_dff_B_Av3Ax3GG9_2;
	wire w_dff_B_lAVYpExO7_2;
	wire w_dff_B_Skuahs6X6_2;
	wire w_dff_B_Kr0RdxBu4_2;
	wire w_dff_B_gRaHvrKl6_2;
	wire w_dff_B_w5jyNEoj4_2;
	wire w_dff_B_zbx9B9IZ0_2;
	wire w_dff_B_4iozQe248_2;
	wire w_dff_B_vAVO0Wtk5_2;
	wire w_dff_B_3VpJpqqL7_2;
	wire w_dff_B_pqCD6kKb8_2;
	wire w_dff_B_Ovd3VDzZ0_2;
	wire w_dff_B_R7Vb8WBB4_2;
	wire w_dff_B_Ui3t7buT2_2;
	wire w_dff_B_CEydjoAt0_2;
	wire w_dff_B_uAcEd9QB0_2;
	wire w_dff_B_3Q7Hm6xA9_2;
	wire w_dff_B_P0KwbxrD7_2;
	wire w_dff_B_3dwfZuv69_2;
	wire w_dff_B_KpchTjCI8_2;
	wire w_dff_B_zFYTX8CP8_2;
	wire w_dff_B_vXMzPBv28_2;
	wire w_dff_B_5DjJHNL86_2;
	wire w_dff_B_G2YbobsN1_2;
	wire w_dff_B_k7A2pZSS8_2;
	wire w_dff_B_h7gOn26C1_2;
	wire w_dff_B_5IOrGMpb5_2;
	wire w_dff_B_mJyNMxgk5_2;
	wire w_dff_B_9E7EO7PV7_2;
	wire w_dff_B_zoqa3g5I7_2;
	wire w_dff_B_LXPE0yOq1_2;
	wire w_dff_B_XsKObT771_1;
	wire w_dff_B_3FDkFYgy2_2;
	wire w_dff_B_DfyloW6U1_2;
	wire w_dff_B_WpmeYibs2_2;
	wire w_dff_B_ismQLkxc5_2;
	wire w_dff_B_f1dVwbxx3_2;
	wire w_dff_B_riePBStL7_2;
	wire w_dff_B_nOoUmHIE0_2;
	wire w_dff_B_VIEZRoua3_2;
	wire w_dff_B_A6ZGEqzY7_2;
	wire w_dff_B_lsQDhDfG6_2;
	wire w_dff_B_QPmYOZp32_2;
	wire w_dff_B_dfgWMsG67_2;
	wire w_dff_B_Oze0BHgY1_2;
	wire w_dff_B_sf5P6DNl2_2;
	wire w_dff_B_mjhS1ujV9_2;
	wire w_dff_B_Tz9mdE135_2;
	wire w_dff_B_qKmbLJQm9_2;
	wire w_dff_B_17SqajER6_2;
	wire w_dff_B_zTJ0d35B7_2;
	wire w_dff_B_tIJncfAq5_2;
	wire w_dff_B_9bg9qoa78_2;
	wire w_dff_B_qjZ2xRDk3_2;
	wire w_dff_B_T2f1wlHB5_2;
	wire w_dff_B_TQ6uh5ey7_2;
	wire w_dff_B_e7uPHoos3_2;
	wire w_dff_B_JB68xpvG4_2;
	wire w_dff_B_kH36B8Jr4_2;
	wire w_dff_B_cb5Lomwy8_2;
	wire w_dff_B_IVyUdDth9_2;
	wire w_dff_B_4unbKKyv2_2;
	wire w_dff_B_NTV0JpaY7_1;
	wire w_dff_B_M6MPbOP08_2;
	wire w_dff_B_HWIc7Vvh2_2;
	wire w_dff_B_X7ICUWdi5_2;
	wire w_dff_B_Us4ZMLs32_2;
	wire w_dff_B_EcnpEkef0_2;
	wire w_dff_B_usBG6r4L1_2;
	wire w_dff_B_qNQGmkJw9_2;
	wire w_dff_B_9E3q66NZ5_2;
	wire w_dff_B_wcSI2O9w3_2;
	wire w_dff_B_GBrbiIcZ4_2;
	wire w_dff_B_8UoTzZZQ5_2;
	wire w_dff_B_lng2jslR6_2;
	wire w_dff_B_ohyiPMzs1_2;
	wire w_dff_B_GcfzvsZZ4_2;
	wire w_dff_B_qyo95S2A8_2;
	wire w_dff_B_xWGnhoyp6_2;
	wire w_dff_B_xLVuIwOM2_2;
	wire w_dff_B_ABRvO3Gm6_2;
	wire w_dff_B_f2NoFdnG4_2;
	wire w_dff_B_F5XSCjvi4_2;
	wire w_dff_B_r5HJCcq01_2;
	wire w_dff_B_bR87hDVs3_2;
	wire w_dff_B_PdAB4Kf17_2;
	wire w_dff_B_5vVkkgl53_2;
	wire w_dff_B_PKyCj2292_2;
	wire w_dff_B_DANe89Pc6_2;
	wire w_dff_B_LVaaCOzx9_2;
	wire w_dff_B_6LIhDnGg7_1;
	wire w_dff_B_WoIHbr2B5_2;
	wire w_dff_B_AAN7k6AH0_2;
	wire w_dff_B_V6xVXnqP7_2;
	wire w_dff_B_IIkvho6D4_2;
	wire w_dff_B_Z9Z0fINg8_2;
	wire w_dff_B_1l5vlHV07_2;
	wire w_dff_B_4waNQHrE1_2;
	wire w_dff_B_xdniJO7t6_2;
	wire w_dff_B_N6wYs5GC1_2;
	wire w_dff_B_GStbbVmn4_2;
	wire w_dff_B_0nNUjlrC5_2;
	wire w_dff_B_uPr6GIUR6_2;
	wire w_dff_B_6q25G7C74_2;
	wire w_dff_B_ukJulgJa1_2;
	wire w_dff_B_yjmTH8IW6_2;
	wire w_dff_B_PQGRwwi04_2;
	wire w_dff_B_4rcKrpCa9_2;
	wire w_dff_B_GT3BDYVb2_2;
	wire w_dff_B_S6rGuAbY3_2;
	wire w_dff_B_GahVn0W57_2;
	wire w_dff_B_ln64X7KU1_2;
	wire w_dff_B_sMPMIBpe6_2;
	wire w_dff_B_M6F2BNcO5_2;
	wire w_dff_B_oht5QqZp1_2;
	wire w_dff_B_pX2KoYxw6_1;
	wire w_dff_B_0uFWQ1TT9_2;
	wire w_dff_B_jYMCYAoZ6_2;
	wire w_dff_B_lYYjqGL49_2;
	wire w_dff_B_Xoy6NoAW4_2;
	wire w_dff_B_IglZLohJ1_2;
	wire w_dff_B_6k9HpCEw6_2;
	wire w_dff_B_nw8Ev4eU7_2;
	wire w_dff_B_SlTpcpa97_2;
	wire w_dff_B_ZVNo4dll0_2;
	wire w_dff_B_K7ZoG8473_2;
	wire w_dff_B_bPzABTjK8_2;
	wire w_dff_B_ElpGkCPY9_2;
	wire w_dff_B_GK7pGRUK9_2;
	wire w_dff_B_LzD6n1ah9_2;
	wire w_dff_B_ue5rVFnc3_2;
	wire w_dff_B_D36rVPAI6_2;
	wire w_dff_B_b9G913cz9_2;
	wire w_dff_B_G7vm2dvU1_2;
	wire w_dff_B_Fl7mkeel8_2;
	wire w_dff_B_rYhzUowM4_2;
	wire w_dff_B_yMyjy5lP9_2;
	wire w_dff_B_TQIgVv3D2_1;
	wire w_dff_B_xKUoSrrP4_2;
	wire w_dff_B_nD9pGQkj7_2;
	wire w_dff_B_9DyghPPn3_2;
	wire w_dff_B_72R75wz33_2;
	wire w_dff_B_LQfYXBSY0_2;
	wire w_dff_B_LbFfgrF16_2;
	wire w_dff_B_rLCUsHLf5_2;
	wire w_dff_B_qyl61W6T4_2;
	wire w_dff_B_sFZEMTdJ3_2;
	wire w_dff_B_cZmosjrc7_2;
	wire w_dff_B_ROpFQ6wA0_2;
	wire w_dff_B_pF6zIYni9_2;
	wire w_dff_B_nnhxoa7W2_2;
	wire w_dff_B_AyeUgQ4M0_2;
	wire w_dff_B_SFfitdX00_2;
	wire w_dff_B_OOSPB0R73_2;
	wire w_dff_B_lOI0ErTq6_2;
	wire w_dff_B_e8521bL50_2;
	wire w_dff_B_CqXK098R2_1;
	wire w_dff_B_CPKbHixs6_2;
	wire w_dff_B_KODDDt5q0_2;
	wire w_dff_B_6PvG91yQ0_2;
	wire w_dff_B_woOb5ry74_2;
	wire w_dff_B_XY5MEbzx4_2;
	wire w_dff_B_2fCRdRov6_2;
	wire w_dff_B_Eg2j2r7n0_2;
	wire w_dff_B_J39YEIGX9_2;
	wire w_dff_B_AiEjmKEm2_2;
	wire w_dff_B_NGJH8CNT2_2;
	wire w_dff_B_aY6f32F14_2;
	wire w_dff_B_WTtcbrbp0_2;
	wire w_dff_B_Xto36zXd3_2;
	wire w_dff_B_6HXXvmvm1_2;
	wire w_dff_B_v1rhBZ8R9_2;
	wire w_dff_B_5jrER1x16_1;
	wire w_dff_B_2AYq0Bwy9_2;
	wire w_dff_B_H6BudrGj4_2;
	wire w_dff_B_3e6kCOJq3_2;
	wire w_dff_B_LUx15ufz7_2;
	wire w_dff_B_crrRVYAr6_2;
	wire w_dff_B_Y6t5K9Je2_2;
	wire w_dff_B_trGqSKB23_2;
	wire w_dff_B_9YpyBDd83_2;
	wire w_dff_B_uzlyiqiE0_2;
	wire w_dff_B_g63P4pV44_2;
	wire w_dff_B_yvjjMG5t8_2;
	wire w_dff_B_ntkPcTrO9_2;
	wire w_dff_B_TtpsuMRV5_1;
	wire w_dff_B_gRzaeMXP6_2;
	wire w_dff_B_Jytmd6hd1_2;
	wire w_dff_B_wgGQbVtJ3_2;
	wire w_dff_B_hwJsTtd18_2;
	wire w_dff_B_B9F1MYl50_2;
	wire w_dff_B_rdo5XgCz3_2;
	wire w_dff_B_IVmnjhSB0_2;
	wire w_dff_B_okQQNJjO8_2;
	wire w_dff_B_XyMDSPbS9_2;
	wire w_dff_B_Hm4uXY3R1_2;
	wire w_dff_B_rD2axpKL5_2;
	wire w_dff_B_xfeIIpLG8_1;
	wire w_dff_B_vue9wlNq3_1;
	wire w_dff_B_8Z4UK4ht2_2;
	wire w_dff_B_o3kYMXiw6_2;
	wire w_dff_B_a9yMZg6v9_2;
	wire w_dff_B_bGahM8op0_0;
	wire w_dff_A_dA4xiOw58_0;
	wire w_dff_A_pOvWQzFu1_0;
	wire w_dff_A_2yDzPjus9_1;
	wire w_dff_A_KrIQk1Yq0_1;
	wire w_dff_B_21KCN8U59_1;
	wire w_dff_A_FN7R7Wuv2_1;
	wire w_dff_B_l9V517vC0_1;
	wire w_dff_B_kDMst8ru0_2;
	wire w_dff_B_IswEgwWA0_2;
	wire w_dff_B_O5n8xANB5_2;
	wire w_dff_B_r5E6ob3k8_2;
	wire w_dff_B_Ra1N4xg39_2;
	wire w_dff_B_GVEJimHn8_2;
	wire w_dff_B_vIy9m4ZJ4_2;
	wire w_dff_B_bLhTxWf84_2;
	wire w_dff_B_TSGgaxC88_2;
	wire w_dff_B_O6AoPGDW7_2;
	wire w_dff_B_CyTUg9zY4_2;
	wire w_dff_B_R9hX5szf3_2;
	wire w_dff_B_4NvmlHSU1_2;
	wire w_dff_B_zLOVYjFV0_2;
	wire w_dff_B_Qw0EP8G27_2;
	wire w_dff_B_pG6bqBe88_2;
	wire w_dff_B_wHzXodWt3_2;
	wire w_dff_B_ZcHLUDGF3_2;
	wire w_dff_B_TPGh4hOh5_2;
	wire w_dff_B_2dfuuemb4_2;
	wire w_dff_B_srbJV4312_2;
	wire w_dff_B_v0HKAo3k6_2;
	wire w_dff_B_bWpJJRTS9_2;
	wire w_dff_B_1Z2HTE6W6_2;
	wire w_dff_B_MX2almsg4_2;
	wire w_dff_B_JtIv3EAd1_2;
	wire w_dff_B_XJXSJ4NN7_2;
	wire w_dff_B_obN1Fa2Y3_2;
	wire w_dff_B_zXAbX5OI6_2;
	wire w_dff_B_HWSRoIsS3_2;
	wire w_dff_B_U7LQDixK0_2;
	wire w_dff_B_U1gigY8K5_2;
	wire w_dff_B_Wk5qA5Vz4_2;
	wire w_dff_B_IjAhIE5b4_2;
	wire w_dff_B_uIwFxCoJ9_2;
	wire w_dff_B_vUmxW7Al8_2;
	wire w_dff_B_JF9L3uyX1_2;
	wire w_dff_B_9ma0up9x1_2;
	wire w_dff_B_oxLHPdvN3_2;
	wire w_dff_B_TdmzmMNp9_2;
	wire w_dff_B_P3OCRb2K7_2;
	wire w_dff_B_J1YjMSLR6_2;
	wire w_dff_B_FBIuk3mv6_2;
	wire w_dff_B_xfZV3ANG5_2;
	wire w_dff_B_tOaXRmgC1_2;
	wire w_dff_B_9eCQOicP7_2;
	wire w_dff_B_WrJ6V0nm5_2;
	wire w_dff_B_t9D5uTt80_1;
	wire w_dff_B_pNYOjhVC9_2;
	wire w_dff_B_5W9X6wvi3_2;
	wire w_dff_B_KHjqwb790_2;
	wire w_dff_B_dbEq4qeh2_2;
	wire w_dff_B_0hyjp00i9_2;
	wire w_dff_B_vZ2J4v7S5_2;
	wire w_dff_B_XUycLhxH7_2;
	wire w_dff_B_tCZoC5kF9_2;
	wire w_dff_B_wjaIMfrg1_2;
	wire w_dff_B_d6EuFWhm9_2;
	wire w_dff_B_SPKceGUe2_2;
	wire w_dff_B_YCDekAtL9_2;
	wire w_dff_B_JlT7ObC32_2;
	wire w_dff_B_S8NFVUaB2_2;
	wire w_dff_B_6X0kgRPa3_2;
	wire w_dff_B_mgBeuNHh3_2;
	wire w_dff_B_msd059e11_2;
	wire w_dff_B_HulELTYO0_2;
	wire w_dff_B_W0i79Icr6_2;
	wire w_dff_B_22ltXU1U5_2;
	wire w_dff_B_tY3PL4BS3_2;
	wire w_dff_B_glmeXJvf3_2;
	wire w_dff_B_BTCRbjOH4_2;
	wire w_dff_B_N1EjSTc73_2;
	wire w_dff_B_IGIG1Wu73_2;
	wire w_dff_B_874iPqy03_2;
	wire w_dff_B_DPySylyg0_2;
	wire w_dff_B_K6RHEaGa7_2;
	wire w_dff_B_IwEq0MXj4_2;
	wire w_dff_B_Ghr6fiuS3_2;
	wire w_dff_B_ybiFY6b38_2;
	wire w_dff_B_uZLDrLUz0_2;
	wire w_dff_B_ahSFkCHz7_2;
	wire w_dff_B_8QPG6n0H4_2;
	wire w_dff_B_sVk5CXUM7_2;
	wire w_dff_B_5L8wzYpj0_2;
	wire w_dff_B_5HqwWtqK8_2;
	wire w_dff_B_viTqWzlJ5_2;
	wire w_dff_B_5yoD2A4C2_2;
	wire w_dff_B_1xWcrS0v9_2;
	wire w_dff_B_2m7wddaq1_2;
	wire w_dff_B_o9zY27mx9_2;
	wire w_dff_B_0qTTQ4Ah9_2;
	wire w_dff_B_XFmAsQRz6_1;
	wire w_dff_B_fvwodyaw1_2;
	wire w_dff_B_gNgMs2UZ8_2;
	wire w_dff_B_syuvkTXI7_2;
	wire w_dff_B_A2vbns6u9_2;
	wire w_dff_B_WJ7efmps6_2;
	wire w_dff_B_C16YQgUm8_2;
	wire w_dff_B_t52tujzu6_2;
	wire w_dff_B_IkwsdRSm2_2;
	wire w_dff_B_JNrRfv6T2_2;
	wire w_dff_B_QzRvDUp34_2;
	wire w_dff_B_san3x6Xe1_2;
	wire w_dff_B_TiZUP3T61_2;
	wire w_dff_B_KYWjDAKY4_2;
	wire w_dff_B_hh3gpvA19_2;
	wire w_dff_B_EDB4rhT63_2;
	wire w_dff_B_ZdiTDCdE8_2;
	wire w_dff_B_6zdidnU93_2;
	wire w_dff_B_Pu5UpHsa0_2;
	wire w_dff_B_GTM5hGc03_2;
	wire w_dff_B_9jsokTcW3_2;
	wire w_dff_B_7cCbKGA89_2;
	wire w_dff_B_6XVx36N21_2;
	wire w_dff_B_0FfbOxez7_2;
	wire w_dff_B_4uYe4nTv3_2;
	wire w_dff_B_uhKaDYun1_2;
	wire w_dff_B_4kvG4O9I4_2;
	wire w_dff_B_zwY4jpUB0_2;
	wire w_dff_B_CRa0TBPZ1_2;
	wire w_dff_B_exNDzymW9_2;
	wire w_dff_B_lTc3NPak9_2;
	wire w_dff_B_c9qIiq8j2_2;
	wire w_dff_B_py3cDcPl0_2;
	wire w_dff_B_TcBjEos55_2;
	wire w_dff_B_FrGPuZe21_2;
	wire w_dff_B_6F0HSgVC7_2;
	wire w_dff_B_e4mtod7U1_2;
	wire w_dff_B_kAtuO9bV5_2;
	wire w_dff_B_PcSwCouR6_2;
	wire w_dff_B_16aT5zsN1_1;
	wire w_dff_B_3pLSN5CG3_2;
	wire w_dff_B_CazexgUy6_2;
	wire w_dff_B_8vyIbKAw5_2;
	wire w_dff_B_YnRnSAN96_2;
	wire w_dff_B_IveJ91e54_2;
	wire w_dff_B_OA9vheDX3_2;
	wire w_dff_B_w0gPgVsl0_2;
	wire w_dff_B_EnltlGRM5_2;
	wire w_dff_B_NtXKQfB58_2;
	wire w_dff_B_2E9D7a5M1_2;
	wire w_dff_B_uRJ3iyoj2_2;
	wire w_dff_B_ef8N4YWm2_2;
	wire w_dff_B_0dFP5lOF9_2;
	wire w_dff_B_6CkqVLE86_2;
	wire w_dff_B_jMVzD7GU2_2;
	wire w_dff_B_EzqaJBGg4_2;
	wire w_dff_B_HHpoGZCe5_2;
	wire w_dff_B_FyVQqYve0_2;
	wire w_dff_B_3MahnG3q5_2;
	wire w_dff_B_uGnD9CkP2_2;
	wire w_dff_B_AqOa60tT2_2;
	wire w_dff_B_SBy6zCVB8_2;
	wire w_dff_B_uhaj9Mai1_2;
	wire w_dff_B_uSF582VV1_2;
	wire w_dff_B_Z62PFuGl9_2;
	wire w_dff_B_Q8k6Skgy8_2;
	wire w_dff_B_7cNMhV7X9_2;
	wire w_dff_B_tHSvPa6A3_2;
	wire w_dff_B_V0Mg8WqM5_2;
	wire w_dff_B_gIZeW8nP4_2;
	wire w_dff_B_6bj8HGa52_2;
	wire w_dff_B_Qpys5LsV2_2;
	wire w_dff_B_Wd5rhdrX9_2;
	wire w_dff_B_3v7FLQP13_2;
	wire w_dff_B_5wq6JhJu8_2;
	wire w_dff_B_wnhFjLNo7_2;
	wire w_dff_B_1GGwFMXf4_1;
	wire w_dff_B_KVsQxj5R5_2;
	wire w_dff_B_avIcZMrb1_2;
	wire w_dff_B_iEXG9xPY9_2;
	wire w_dff_B_WkLhh7J52_2;
	wire w_dff_B_frBDfW6X0_2;
	wire w_dff_B_sLa1qN8a2_2;
	wire w_dff_B_pRjce0Ks8_2;
	wire w_dff_B_ytoBCoOm1_2;
	wire w_dff_B_sEyaELGB1_2;
	wire w_dff_B_i4n86loG1_2;
	wire w_dff_B_MH75h9N42_2;
	wire w_dff_B_ccx6fG382_2;
	wire w_dff_B_qErzRpsU7_2;
	wire w_dff_B_KnTHTJ6V6_2;
	wire w_dff_B_92WceIax7_2;
	wire w_dff_B_qgo46wpE7_2;
	wire w_dff_B_fXnTDbjO6_2;
	wire w_dff_B_eUYFIQY90_2;
	wire w_dff_B_NssLkWHN1_2;
	wire w_dff_B_zFHoNNH77_2;
	wire w_dff_B_V4VrACSw7_2;
	wire w_dff_B_GoZvDL4v5_2;
	wire w_dff_B_s9opWJOP0_2;
	wire w_dff_B_FW0RCixr1_2;
	wire w_dff_B_6uEMwGVI0_2;
	wire w_dff_B_7aWfhsmM8_2;
	wire w_dff_B_l7O45QNP2_2;
	wire w_dff_B_rswdLXD06_2;
	wire w_dff_B_R8TsZpYj4_2;
	wire w_dff_B_8gPLJpK13_2;
	wire w_dff_B_icy7nypp6_2;
	wire w_dff_B_kL36koVf8_2;
	wire w_dff_B_QSdI15m68_2;
	wire w_dff_B_03C4d0Nz5_1;
	wire w_dff_B_ZTRAGPzd5_2;
	wire w_dff_B_9mUIdDGm1_2;
	wire w_dff_B_sRiNvewp2_2;
	wire w_dff_B_SCk0ElQf8_2;
	wire w_dff_B_6Qw9lyRy7_2;
	wire w_dff_B_HcrkmSGr1_2;
	wire w_dff_B_PcIRYYr12_2;
	wire w_dff_B_IuBtgw9k2_2;
	wire w_dff_B_cCjUmUSv2_2;
	wire w_dff_B_mCgLaQyL4_2;
	wire w_dff_B_SvrCyC528_2;
	wire w_dff_B_LVEWAfhX3_2;
	wire w_dff_B_rfA7ybRF7_2;
	wire w_dff_B_6RdFhHoK9_2;
	wire w_dff_B_IMN8IZXh3_2;
	wire w_dff_B_i5BBpHps1_2;
	wire w_dff_B_EDWDpFGB3_2;
	wire w_dff_B_LG7Q3p3Z0_2;
	wire w_dff_B_ZIM0uiyb7_2;
	wire w_dff_B_NRyVUIUT4_2;
	wire w_dff_B_3bFWeXvq1_2;
	wire w_dff_B_fCgLx2Ab8_2;
	wire w_dff_B_Qy1bWVMt1_2;
	wire w_dff_B_TOdpPG1v6_2;
	wire w_dff_B_S0umS0Q60_2;
	wire w_dff_B_89mD8GuJ6_2;
	wire w_dff_B_vSKpSpCu6_2;
	wire w_dff_B_2AvGAdzv3_2;
	wire w_dff_B_B4idFpAm8_2;
	wire w_dff_B_FMdovfI97_2;
	wire w_dff_B_3YJs9FYL7_1;
	wire w_dff_B_O909kjOB6_2;
	wire w_dff_B_9cjHc9BA0_2;
	wire w_dff_B_MVX68V2I7_2;
	wire w_dff_B_JKNQFBoV8_2;
	wire w_dff_B_uKLSG0b28_2;
	wire w_dff_B_H9Dp2Wn96_2;
	wire w_dff_B_dFG8EpLY0_2;
	wire w_dff_B_kp039gr16_2;
	wire w_dff_B_3DKnH1Yz6_2;
	wire w_dff_B_YPKdWiKd3_2;
	wire w_dff_B_gwKTBcxk1_2;
	wire w_dff_B_VMQBcAm46_2;
	wire w_dff_B_hYocLxTP7_2;
	wire w_dff_B_dou3UOQX5_2;
	wire w_dff_B_OSju6Gw70_2;
	wire w_dff_B_PzPFNVaN8_2;
	wire w_dff_B_wdwGwaL93_2;
	wire w_dff_B_MeVbMxQn0_2;
	wire w_dff_B_XnuWoWXB9_2;
	wire w_dff_B_iLwZvHKa8_2;
	wire w_dff_B_R6KMT4Hv1_2;
	wire w_dff_B_wkF0Ap7w4_2;
	wire w_dff_B_VHx9nbKy2_2;
	wire w_dff_B_syeGgtK06_2;
	wire w_dff_B_8f5t40EH4_2;
	wire w_dff_B_vPZYQ9446_2;
	wire w_dff_B_Lm9mW8yr3_2;
	wire w_dff_B_r1b8WR3B7_1;
	wire w_dff_B_x3mFtPrJ8_2;
	wire w_dff_B_liXXXrSw7_2;
	wire w_dff_B_EUqn5DNy8_2;
	wire w_dff_B_L8DOvECq1_2;
	wire w_dff_B_GZwLpp811_2;
	wire w_dff_B_i7kLmSo80_2;
	wire w_dff_B_ziWRDt3A1_2;
	wire w_dff_B_zxyjUr9d6_2;
	wire w_dff_B_Iil3oNRz3_2;
	wire w_dff_B_9GIOokJC5_2;
	wire w_dff_B_SgO2pyAa9_2;
	wire w_dff_B_k6iOAHRL2_2;
	wire w_dff_B_qk8FC8x47_2;
	wire w_dff_B_wb14hT8h8_2;
	wire w_dff_B_PDZxi2Ag9_2;
	wire w_dff_B_IGOaujNL1_2;
	wire w_dff_B_91cugucc0_2;
	wire w_dff_B_PMNHLCSo4_2;
	wire w_dff_B_Nu2s07Qw3_2;
	wire w_dff_B_lIQmthI84_2;
	wire w_dff_B_osVDgbw17_2;
	wire w_dff_B_Z6oTmj7y9_2;
	wire w_dff_B_04xkvR896_2;
	wire w_dff_B_y33tYOu80_2;
	wire w_dff_B_dFvhUsMM4_1;
	wire w_dff_B_51y7hsma4_2;
	wire w_dff_B_f1KX6mMl1_2;
	wire w_dff_B_bIDddtaF4_2;
	wire w_dff_B_GwOFstOW2_2;
	wire w_dff_B_TmlORck29_2;
	wire w_dff_B_hbDt7uwv2_2;
	wire w_dff_B_fAU1TFqW5_2;
	wire w_dff_B_vnrKLf7b2_2;
	wire w_dff_B_pAnLs9fe8_2;
	wire w_dff_B_5eKEgA4p4_2;
	wire w_dff_B_Y3Aqfz2K4_2;
	wire w_dff_B_pcHUbSNj9_2;
	wire w_dff_B_Wf9ylcjt6_2;
	wire w_dff_B_KvGUxGQp0_2;
	wire w_dff_B_BeL5p8Pj2_2;
	wire w_dff_B_6Iu4fln07_2;
	wire w_dff_B_YvpQtGn88_2;
	wire w_dff_B_Qn9R1tgg8_2;
	wire w_dff_B_WTLmxP1M8_2;
	wire w_dff_B_7FGqqgOK4_2;
	wire w_dff_B_MV1nrUwB4_2;
	wire w_dff_B_cexRrHv16_1;
	wire w_dff_B_KWlvKiXB7_2;
	wire w_dff_B_oqHToH5b6_2;
	wire w_dff_B_sHph7eFO0_2;
	wire w_dff_B_tFYH2YVv9_2;
	wire w_dff_B_8WGE9fUd9_2;
	wire w_dff_B_iBJUXVJm7_2;
	wire w_dff_B_1e6Oejm25_2;
	wire w_dff_B_Tyy0JRCP1_2;
	wire w_dff_B_MD93t9ql0_2;
	wire w_dff_B_NYJavSmY3_2;
	wire w_dff_B_jQGM1Ts92_2;
	wire w_dff_B_hYmhH8Wz1_2;
	wire w_dff_B_0zZ2AAQo3_2;
	wire w_dff_B_Cxmen5VL8_2;
	wire w_dff_B_JzCAXZbT5_2;
	wire w_dff_B_z7HxxPCg7_2;
	wire w_dff_B_7uNOedha2_2;
	wire w_dff_B_UZquPyqL3_2;
	wire w_dff_B_RcaNpk1T7_1;
	wire w_dff_B_jyD9jlPS1_2;
	wire w_dff_B_M1MrszxR0_2;
	wire w_dff_B_be2rJyGh9_2;
	wire w_dff_B_l1sSRFEA6_2;
	wire w_dff_B_obOo6bfF4_2;
	wire w_dff_B_Auk0EMZ11_2;
	wire w_dff_B_pjGDfKvY6_2;
	wire w_dff_B_a3WcKyJ41_2;
	wire w_dff_B_6guXQXpl8_2;
	wire w_dff_B_iDqmTMMw8_2;
	wire w_dff_B_obKF3JNN7_2;
	wire w_dff_B_c7kGDYuK5_2;
	wire w_dff_B_2a9Kgfqe3_2;
	wire w_dff_B_6GItylHC3_2;
	wire w_dff_B_Wvs81bCN0_2;
	wire w_dff_B_3kdNpIDS2_1;
	wire w_dff_B_4UDEevnT5_2;
	wire w_dff_B_uz8Ib7D22_2;
	wire w_dff_B_qwaZHtGz0_2;
	wire w_dff_B_W3BAzdNv3_2;
	wire w_dff_B_ioPUdqXo0_2;
	wire w_dff_B_qJavXmVr2_2;
	wire w_dff_B_6MfAlA2I6_2;
	wire w_dff_B_pZG3zAAN2_2;
	wire w_dff_B_n3oivF5S0_2;
	wire w_dff_B_RjfTGN7b6_2;
	wire w_dff_B_XovSSTRy2_2;
	wire w_dff_B_1s3Leg2W0_2;
	wire w_dff_B_58V6RV5c9_1;
	wire w_dff_B_1DtK8UZq9_2;
	wire w_dff_B_hv0zbFXF1_2;
	wire w_dff_B_k0T8pjKR3_2;
	wire w_dff_B_JnbiRzxM6_2;
	wire w_dff_B_yve8NB3J4_2;
	wire w_dff_B_eJDvWjLt3_2;
	wire w_dff_B_aFnSAuSM5_2;
	wire w_dff_B_NcfWduB29_2;
	wire w_dff_B_uaazYh8H4_2;
	wire w_dff_B_FR9pN9Gn5_2;
	wire w_dff_B_NnRZQt6k9_2;
	wire w_dff_B_lctd7zUT2_1;
	wire w_dff_B_sNSkNFS63_1;
	wire w_dff_B_OxJMzRfB7_2;
	wire w_dff_B_Ms7VltmA1_2;
	wire w_dff_B_t8ZJcDmB0_2;
	wire w_dff_B_wGRbh8jc5_0;
	wire w_dff_A_io4gw1MZ2_0;
	wire w_dff_A_t6iX48tA8_0;
	wire w_dff_A_YF2EYJSt0_1;
	wire w_dff_A_qZksD9iJ4_1;
	wire w_dff_B_BKablcen2_1;
	wire w_dff_A_bsSlG3hO7_1;
	wire w_dff_B_FcTF5d0h3_1;
	wire w_dff_B_OUBhC1NO7_2;
	wire w_dff_B_fmJtwFIt2_2;
	wire w_dff_B_ItwRgNHp0_2;
	wire w_dff_B_Pw74HCmk5_2;
	wire w_dff_B_whysWFLh7_2;
	wire w_dff_B_vFHUHe1I6_2;
	wire w_dff_B_dNBzMi9l1_2;
	wire w_dff_B_t4aK7ddr9_2;
	wire w_dff_B_VRfdxMMV1_2;
	wire w_dff_B_PANLaeBs9_2;
	wire w_dff_B_lPWXXIzo8_2;
	wire w_dff_B_M36Y5qE90_2;
	wire w_dff_B_KfefUwkb1_2;
	wire w_dff_B_d71AzNVT2_2;
	wire w_dff_B_MMHvZwqM3_2;
	wire w_dff_B_0mPgEUwx9_2;
	wire w_dff_B_5VK78K6H1_2;
	wire w_dff_B_TP73D6c32_2;
	wire w_dff_B_lBaP8azp5_2;
	wire w_dff_B_Uvkgl5ZA7_2;
	wire w_dff_B_n4ysy3ao2_2;
	wire w_dff_B_g4XX9DeR3_2;
	wire w_dff_B_Ov3UanVv7_2;
	wire w_dff_B_FD0NL8Vi5_2;
	wire w_dff_B_VwtkVktY9_2;
	wire w_dff_B_ZRWJtusi2_2;
	wire w_dff_B_ipL11gTl0_2;
	wire w_dff_B_YJxHvJrQ8_2;
	wire w_dff_B_sFVwPFI35_2;
	wire w_dff_B_ZQKVMXdx0_2;
	wire w_dff_B_EAc4G7fo3_2;
	wire w_dff_B_QM6cG2iy0_2;
	wire w_dff_B_UkqzuT5k3_2;
	wire w_dff_B_J0lgCcYt9_2;
	wire w_dff_B_hQQo2If56_2;
	wire w_dff_B_2mlZENjF0_2;
	wire w_dff_B_khVW1U4E7_2;
	wire w_dff_B_26yFExap6_2;
	wire w_dff_B_gxIDlyg10_2;
	wire w_dff_B_HfKV2YGx6_2;
	wire w_dff_B_F85Oe1U58_2;
	wire w_dff_B_Dq8tn5gX4_2;
	wire w_dff_B_ude87cpT0_2;
	wire w_dff_B_T19x75My6_2;
	wire w_dff_B_QhLcJXdJ5_2;
	wire w_dff_B_VYjkvQDf1_2;
	wire w_dff_B_UTmKQY3Q3_2;
	wire w_dff_B_a2Kjpush8_2;
	wire w_dff_B_YwNIF9Vn6_2;
	wire w_dff_B_jjFo3b7d1_1;
	wire w_dff_B_eHB6nEBG0_2;
	wire w_dff_B_CHEiYN1l4_2;
	wire w_dff_B_72yhTXIg5_2;
	wire w_dff_B_4La54H0s1_2;
	wire w_dff_B_RtkH3Ulv6_2;
	wire w_dff_B_6Yrhcs9R7_2;
	wire w_dff_B_Sq5xUdzH9_2;
	wire w_dff_B_uMw4oF765_2;
	wire w_dff_B_kNMwuPsa4_2;
	wire w_dff_B_UHhjEkkI4_2;
	wire w_dff_B_9d4qtsyr5_2;
	wire w_dff_B_z06po0zU3_2;
	wire w_dff_B_VaWOY6TC8_2;
	wire w_dff_B_mwnjfS311_2;
	wire w_dff_B_ImxED3zz2_2;
	wire w_dff_B_UEAyJW5l1_2;
	wire w_dff_B_guwLKsvS8_2;
	wire w_dff_B_sHHvjsPS6_2;
	wire w_dff_B_qzHT2KNb3_2;
	wire w_dff_B_ocGRKwGS9_2;
	wire w_dff_B_rnd3yGtu5_2;
	wire w_dff_B_t7kK7vpJ3_2;
	wire w_dff_B_khTexeY66_2;
	wire w_dff_B_AP9FniQL4_2;
	wire w_dff_B_2CZ094Zn5_2;
	wire w_dff_B_g0ETjYvw9_2;
	wire w_dff_B_wGwYkgyp5_2;
	wire w_dff_B_TXFvDDTV0_2;
	wire w_dff_B_gnDsqmLA8_2;
	wire w_dff_B_lxBOVhXB5_2;
	wire w_dff_B_WrAUXnFC0_2;
	wire w_dff_B_E27KxMi70_2;
	wire w_dff_B_7zabKwqo9_2;
	wire w_dff_B_HeJAS2282_2;
	wire w_dff_B_7tKD9LPK4_2;
	wire w_dff_B_W9udXep88_2;
	wire w_dff_B_iMWVDoie5_2;
	wire w_dff_B_Gi4ooOp19_2;
	wire w_dff_B_UP7BAiTN3_2;
	wire w_dff_B_H4cSGW3E7_2;
	wire w_dff_B_46d62AYL0_2;
	wire w_dff_B_PL5uDZ9L5_2;
	wire w_dff_B_v7fAg0fD1_2;
	wire w_dff_B_9Pq9g6YL3_2;
	wire w_dff_B_mPJtTvrl4_2;
	wire w_dff_B_J1dXw1Si3_1;
	wire w_dff_B_DEXGpvSM7_2;
	wire w_dff_B_eFLJveyf3_2;
	wire w_dff_B_bOCPJfyW8_2;
	wire w_dff_B_36b6XdMD6_2;
	wire w_dff_B_pdwZLhvl3_2;
	wire w_dff_B_odG7Wl2P6_2;
	wire w_dff_B_2sxTNxK93_2;
	wire w_dff_B_5HARTNgB6_2;
	wire w_dff_B_YqYrLMvF8_2;
	wire w_dff_B_G9TyQWZW5_2;
	wire w_dff_B_JSaBwnQg6_2;
	wire w_dff_B_DbpJXVVX7_2;
	wire w_dff_B_fHojTLNq4_2;
	wire w_dff_B_5jDJJQiJ9_2;
	wire w_dff_B_N384otp13_2;
	wire w_dff_B_zWavUoES0_2;
	wire w_dff_B_eku0LzPZ7_2;
	wire w_dff_B_VFJ0Nj5D8_2;
	wire w_dff_B_lYXCGiOs8_2;
	wire w_dff_B_6ZsLZ4wK5_2;
	wire w_dff_B_LVfbHczP4_2;
	wire w_dff_B_0uX0iXsO9_2;
	wire w_dff_B_hNUFNmTL6_2;
	wire w_dff_B_nVotZP695_2;
	wire w_dff_B_p8pibRlP1_2;
	wire w_dff_B_5gPiEYGt8_2;
	wire w_dff_B_xHWM1olY6_2;
	wire w_dff_B_Si4HnNJr4_2;
	wire w_dff_B_vsiNTbZV0_2;
	wire w_dff_B_2mmrACs66_2;
	wire w_dff_B_Yd0GGByz4_2;
	wire w_dff_B_Lcm8LdNh2_2;
	wire w_dff_B_SAlxpB8D1_2;
	wire w_dff_B_x34HdRjl9_2;
	wire w_dff_B_XrvjAUW74_2;
	wire w_dff_B_fxaBQXP27_2;
	wire w_dff_B_MHLn6Nhr9_2;
	wire w_dff_B_pKNsPfbR9_2;
	wire w_dff_B_J5dSF4jh3_2;
	wire w_dff_B_NWclf5rq6_2;
	wire w_dff_B_s48Z0v4b3_2;
	wire w_dff_B_NToFGzAQ7_1;
	wire w_dff_B_vJXJgwPJ0_2;
	wire w_dff_B_CVcrzpfv7_2;
	wire w_dff_B_nQi6u14K6_2;
	wire w_dff_B_x120Z6yC1_2;
	wire w_dff_B_NM3kxtf45_2;
	wire w_dff_B_ATZybB8C1_2;
	wire w_dff_B_iIPdcsum9_2;
	wire w_dff_B_B2ObvuDJ1_2;
	wire w_dff_B_mB0evKK29_2;
	wire w_dff_B_z25aOPCP0_2;
	wire w_dff_B_mCc2ME7p8_2;
	wire w_dff_B_1UZJbKRA5_2;
	wire w_dff_B_4kijFdoW6_2;
	wire w_dff_B_l6Z6BXob2_2;
	wire w_dff_B_CZOEVuH90_2;
	wire w_dff_B_TY7LN03v8_2;
	wire w_dff_B_CYochupi6_2;
	wire w_dff_B_F2Boja8F4_2;
	wire w_dff_B_ssP6s4HK2_2;
	wire w_dff_B_t20TExDa2_2;
	wire w_dff_B_ClGlmacp8_2;
	wire w_dff_B_94sdIFXV0_2;
	wire w_dff_B_StdHmQqc6_2;
	wire w_dff_B_5yjgYhqu5_2;
	wire w_dff_B_fca5CBu10_2;
	wire w_dff_B_p3NBk60j6_2;
	wire w_dff_B_0ToTjtN56_2;
	wire w_dff_B_wn77oDMg1_2;
	wire w_dff_B_OwSITP280_2;
	wire w_dff_B_sjpAV16v1_2;
	wire w_dff_B_AfNT8kK71_2;
	wire w_dff_B_6h4ar9Ku6_2;
	wire w_dff_B_iJiDvakS7_2;
	wire w_dff_B_ZebamhUt0_2;
	wire w_dff_B_qgPNeUjA1_2;
	wire w_dff_B_7fjS4I5R0_2;
	wire w_dff_B_t8ZmUGWO1_2;
	wire w_dff_B_Q7YT2tXl2_1;
	wire w_dff_B_WYVJMJUn5_2;
	wire w_dff_B_ScVhj7am9_2;
	wire w_dff_B_ViNS0e246_2;
	wire w_dff_B_plE4owDJ0_2;
	wire w_dff_B_hfQVAflm3_2;
	wire w_dff_B_BhI42FS42_2;
	wire w_dff_B_npJAnwln5_2;
	wire w_dff_B_iRAuH4e56_2;
	wire w_dff_B_Y0uNT97w2_2;
	wire w_dff_B_c0z3FUhU2_2;
	wire w_dff_B_uNIK081t0_2;
	wire w_dff_B_6LMh9R2C2_2;
	wire w_dff_B_ZuJihfnl6_2;
	wire w_dff_B_yWFHp9fQ3_2;
	wire w_dff_B_vLvjLSms5_2;
	wire w_dff_B_iUJ8DrRb0_2;
	wire w_dff_B_cCIonvuG0_2;
	wire w_dff_B_EoGS1bbT2_2;
	wire w_dff_B_qRhLGgjD0_2;
	wire w_dff_B_BjXSP8lL4_2;
	wire w_dff_B_eA1aXsB79_2;
	wire w_dff_B_DnIDgaQK8_2;
	wire w_dff_B_2kSrcUO43_2;
	wire w_dff_B_E8yQ1OjJ7_2;
	wire w_dff_B_bSLruTOz6_2;
	wire w_dff_B_OJt0hsBe1_2;
	wire w_dff_B_eJJuzPRJ5_2;
	wire w_dff_B_CpjqXGqa7_2;
	wire w_dff_B_FhCzXo9Y4_2;
	wire w_dff_B_oCKEaP5c6_2;
	wire w_dff_B_FbhpoCpu2_2;
	wire w_dff_B_JzzDAZy18_2;
	wire w_dff_B_KqDwvtXB8_1;
	wire w_dff_B_4MW1dy5I3_2;
	wire w_dff_B_xBzRkKfh2_2;
	wire w_dff_B_tOcnGwwS4_2;
	wire w_dff_B_CuP3tzkD3_2;
	wire w_dff_B_ePe6b4s39_2;
	wire w_dff_B_KCEdPDOJ8_2;
	wire w_dff_B_kjyESEy86_2;
	wire w_dff_B_Cwx4TogP5_2;
	wire w_dff_B_XOyxlPop0_2;
	wire w_dff_B_SUnJpseU0_2;
	wire w_dff_B_Ad940SHD2_2;
	wire w_dff_B_sDMmGItq3_2;
	wire w_dff_B_xQwMSEmP7_2;
	wire w_dff_B_TZq1nyMg9_2;
	wire w_dff_B_GoF85LcZ0_2;
	wire w_dff_B_ArDhKMWe6_2;
	wire w_dff_B_FZWaVXJO4_2;
	wire w_dff_B_ldOADhiu5_2;
	wire w_dff_B_oaREJ4IR5_2;
	wire w_dff_B_8z27Dhzj8_2;
	wire w_dff_B_N2xtKETd9_2;
	wire w_dff_B_hbCXoDJi4_2;
	wire w_dff_B_tw11y9qt5_2;
	wire w_dff_B_F5wxppnt0_2;
	wire w_dff_B_m94nor1V1_2;
	wire w_dff_B_W4ymwp633_2;
	wire w_dff_B_axL7CF5E3_2;
	wire w_dff_B_ji4cfoxE8_2;
	wire w_dff_B_XU9zNzmb9_2;
	wire w_dff_B_7AmvrWmr2_2;
	wire w_dff_B_fhgkpsz11_1;
	wire w_dff_B_J0m5tXEJ0_2;
	wire w_dff_B_M7zkUsJD9_2;
	wire w_dff_B_0PW2za2H2_2;
	wire w_dff_B_sBefOyIN1_2;
	wire w_dff_B_WOqdT7zu6_2;
	wire w_dff_B_FYe3N1UV9_2;
	wire w_dff_B_u7h2gh5a1_2;
	wire w_dff_B_rL7bf5Xe0_2;
	wire w_dff_B_6e4h2Ofw5_2;
	wire w_dff_B_yyxgltEE0_2;
	wire w_dff_B_7iH8rB9v4_2;
	wire w_dff_B_KzE6huZh7_2;
	wire w_dff_B_mQY3A42h5_2;
	wire w_dff_B_kn0q0M0M4_2;
	wire w_dff_B_qzmXuNxB3_2;
	wire w_dff_B_LGULOmy35_2;
	wire w_dff_B_WYg5GW4C8_2;
	wire w_dff_B_9OEULCYx5_2;
	wire w_dff_B_qbHmGXhI1_2;
	wire w_dff_B_wOTDmG5X4_2;
	wire w_dff_B_IcJzz89m2_2;
	wire w_dff_B_9SsYb6J03_2;
	wire w_dff_B_VNRioU9r3_2;
	wire w_dff_B_ApGWT2H27_2;
	wire w_dff_B_PemKooQa6_2;
	wire w_dff_B_LDWxq2Tz1_2;
	wire w_dff_B_oXKCQvLj0_2;
	wire w_dff_B_RCvdprrW0_1;
	wire w_dff_B_K6oej78G5_2;
	wire w_dff_B_mbWKxVcy1_2;
	wire w_dff_B_UO3mjFJ69_2;
	wire w_dff_B_WtkGxZ4T0_2;
	wire w_dff_B_yQXfnlFn1_2;
	wire w_dff_B_AylUQdnU8_2;
	wire w_dff_B_RhSjcLl70_2;
	wire w_dff_B_UxqJJMzN7_2;
	wire w_dff_B_vwIjTXup1_2;
	wire w_dff_B_7Pjut8BE2_2;
	wire w_dff_B_0tfE0Zod5_2;
	wire w_dff_B_gzXi3Ktd1_2;
	wire w_dff_B_oVi7Px857_2;
	wire w_dff_B_IwYVabqU5_2;
	wire w_dff_B_t2pHHfU22_2;
	wire w_dff_B_AkPOQ7AW2_2;
	wire w_dff_B_ZTAd8W0A4_2;
	wire w_dff_B_JX6xhG9F6_2;
	wire w_dff_B_hhOQQPkJ8_2;
	wire w_dff_B_6uh1CL0c9_2;
	wire w_dff_B_07sf7OJa5_2;
	wire w_dff_B_Mg0dzEFw8_2;
	wire w_dff_B_rWoV4dyW9_2;
	wire w_dff_B_XFi4CKxd4_2;
	wire w_dff_B_XA6EwYAF0_1;
	wire w_dff_B_ZgFSeLE93_2;
	wire w_dff_B_4kXPqXZx7_2;
	wire w_dff_B_preJuuKJ6_2;
	wire w_dff_B_6JMv849W1_2;
	wire w_dff_B_nGeIk8gy3_2;
	wire w_dff_B_fsE8v4dZ8_2;
	wire w_dff_B_z9VJK7IZ7_2;
	wire w_dff_B_kQ3OXmrY2_2;
	wire w_dff_B_d14JP68W0_2;
	wire w_dff_B_sEJTVhfV8_2;
	wire w_dff_B_q7VaESVD2_2;
	wire w_dff_B_z3LdGgzA6_2;
	wire w_dff_B_s6Uw1iiy0_2;
	wire w_dff_B_AWaUS11O1_2;
	wire w_dff_B_UHC1K1kB7_2;
	wire w_dff_B_C3mduFv11_2;
	wire w_dff_B_NKA4irhU5_2;
	wire w_dff_B_aLmtdjwg7_2;
	wire w_dff_B_nV1wXi2P0_2;
	wire w_dff_B_2uCsVlcn6_2;
	wire w_dff_B_p4KQoNjV9_2;
	wire w_dff_B_Klmu89BJ8_1;
	wire w_dff_B_VhtQ0F8U1_2;
	wire w_dff_B_S41vNDXG9_2;
	wire w_dff_B_5FkHNdIs9_2;
	wire w_dff_B_DHaLOYlK7_2;
	wire w_dff_B_D0p5I5LU2_2;
	wire w_dff_B_s1sw8CgJ1_2;
	wire w_dff_B_Imy5NynV1_2;
	wire w_dff_B_nrLixpA81_2;
	wire w_dff_B_4yLsAD8X9_2;
	wire w_dff_B_ilrJxCb46_2;
	wire w_dff_B_ws29kss34_2;
	wire w_dff_B_3RbpLpql2_2;
	wire w_dff_B_bO280q4X1_2;
	wire w_dff_B_O3ciAwDl7_2;
	wire w_dff_B_XgTjRMOj1_2;
	wire w_dff_B_z8K4H9mD3_2;
	wire w_dff_B_UBQUdD8G3_2;
	wire w_dff_B_9dj6N0cZ0_2;
	wire w_dff_B_lElzpUqB8_1;
	wire w_dff_B_I99xRRJk7_2;
	wire w_dff_B_bRlAjyl20_2;
	wire w_dff_B_ihixATLA1_2;
	wire w_dff_B_hC0M6Dok5_2;
	wire w_dff_B_hq3ZFMDV9_2;
	wire w_dff_B_HD64EQci4_2;
	wire w_dff_B_xMu8lGfQ9_2;
	wire w_dff_B_aXNFyKXY9_2;
	wire w_dff_B_dXW1jjuC2_2;
	wire w_dff_B_9TMbwzxA3_2;
	wire w_dff_B_YY3jv06z6_2;
	wire w_dff_B_j0QtQlh04_2;
	wire w_dff_B_92GYoN5c6_2;
	wire w_dff_B_GpUGpCoU0_2;
	wire w_dff_B_FFyMfjKa9_2;
	wire w_dff_B_AEG78ezj7_1;
	wire w_dff_B_3pGNk0yz0_2;
	wire w_dff_B_FooUfOxn0_2;
	wire w_dff_B_pMR0IVFP0_2;
	wire w_dff_B_rRswQRFe0_2;
	wire w_dff_B_dzeX0QTt6_2;
	wire w_dff_B_YfGZtyco7_2;
	wire w_dff_B_yC0Dj2CN2_2;
	wire w_dff_B_YecMjM0H4_2;
	wire w_dff_B_SsgKgUyf4_2;
	wire w_dff_B_bIphNa268_2;
	wire w_dff_B_wSkPVZ5H8_2;
	wire w_dff_B_R921Ezfz5_2;
	wire w_dff_B_mHlV8etn5_1;
	wire w_dff_B_ybLsXfET3_2;
	wire w_dff_B_i7KImOju7_2;
	wire w_dff_B_P8FnVOW29_2;
	wire w_dff_B_cYHompDw4_2;
	wire w_dff_B_a0jShjwR1_2;
	wire w_dff_B_cSQmYooW7_2;
	wire w_dff_B_JQI5isGO9_2;
	wire w_dff_B_EXRxjeOL2_2;
	wire w_dff_B_pEsvVSsL5_2;
	wire w_dff_B_28L4XTPF9_2;
	wire w_dff_B_px5urLfF6_2;
	wire w_dff_B_ndMJxwyC9_1;
	wire w_dff_B_ny94K4xr4_1;
	wire w_dff_B_6OKlmBQJ6_2;
	wire w_dff_B_QDOksBRU7_2;
	wire w_dff_B_ymoeGeBM1_2;
	wire w_dff_B_2G8Dmrc76_0;
	wire w_dff_A_5u9AfVKa4_0;
	wire w_dff_A_lI9Tl6Ax2_0;
	wire w_dff_A_toJ3qaRi7_1;
	wire w_dff_A_SA268giF4_1;
	wire w_dff_B_gTft9evD3_1;
	wire w_dff_A_qYRAclYB1_1;
	wire w_dff_B_OVSklzkW6_1;
	wire w_dff_B_CBTpJeBU1_2;
	wire w_dff_B_cWF9zexF1_2;
	wire w_dff_B_LhDtNopF9_2;
	wire w_dff_B_e1VZUiPv8_2;
	wire w_dff_B_wE7C7L9t3_2;
	wire w_dff_B_CJ7gv1az3_2;
	wire w_dff_B_CybqY79d8_2;
	wire w_dff_B_NMnYLpWk7_2;
	wire w_dff_B_x8EaEdZO8_2;
	wire w_dff_B_VVrmtqHx5_2;
	wire w_dff_B_flKJsC0X0_2;
	wire w_dff_B_zJwt8dYs8_2;
	wire w_dff_B_czGG51lP5_2;
	wire w_dff_B_fT49r7xT1_2;
	wire w_dff_B_xxup8haT6_2;
	wire w_dff_B_ABDIfSrK3_2;
	wire w_dff_B_THITAzdv3_2;
	wire w_dff_B_6StuxNoU3_2;
	wire w_dff_B_hSJDsKhL3_2;
	wire w_dff_B_MqvlbyyA9_2;
	wire w_dff_B_5GRkqyut1_2;
	wire w_dff_B_z2AAoVie6_2;
	wire w_dff_B_xFmRr5hD8_2;
	wire w_dff_B_1EI6BfdN1_2;
	wire w_dff_B_rwsV5ITJ7_2;
	wire w_dff_B_i6TtNGgf4_2;
	wire w_dff_B_LVa7GPqN8_2;
	wire w_dff_B_S92yJVOM2_2;
	wire w_dff_B_BbrlAjXw0_2;
	wire w_dff_B_XmjbQ9ms5_2;
	wire w_dff_B_04cfFUiZ1_2;
	wire w_dff_B_dvjIDWEU1_2;
	wire w_dff_B_K3vfERUE5_2;
	wire w_dff_B_9P0P5iPE6_2;
	wire w_dff_B_g0v9ARu22_2;
	wire w_dff_B_79ohoplp4_2;
	wire w_dff_B_7kBKBRLV9_2;
	wire w_dff_B_3FU7fnm00_2;
	wire w_dff_B_JKUv5p9S3_2;
	wire w_dff_B_mNSbcnuv1_2;
	wire w_dff_B_PA4h3NaM5_2;
	wire w_dff_B_689Pt4u27_2;
	wire w_dff_B_aXoTpu649_2;
	wire w_dff_B_Pmw4J4Ih7_2;
	wire w_dff_B_krbNcL2i3_2;
	wire w_dff_B_8Dxmp4ON5_2;
	wire w_dff_B_B97tuTB35_2;
	wire w_dff_B_p5pi7sEK0_2;
	wire w_dff_B_7lIgAyzM7_2;
	wire w_dff_B_5eC0TGI62_2;
	wire w_dff_B_M75QlrxF7_2;
	wire w_dff_B_IJm0KGB21_1;
	wire w_dff_B_ewmSuU8E4_2;
	wire w_dff_B_se2OTqVx4_2;
	wire w_dff_B_xpCqhpgU5_2;
	wire w_dff_B_IOrp231l9_2;
	wire w_dff_B_z3XbKRlS4_2;
	wire w_dff_B_DfeeHPYi6_2;
	wire w_dff_B_tUQStImV2_2;
	wire w_dff_B_MuUMjhc89_2;
	wire w_dff_B_kFPuXkXY5_2;
	wire w_dff_B_KIpOZCrK4_2;
	wire w_dff_B_psENIpg98_2;
	wire w_dff_B_yzVsX0nW7_2;
	wire w_dff_B_Z50GMZMd8_2;
	wire w_dff_B_s2X1SFth1_2;
	wire w_dff_B_IPKxiNFC4_2;
	wire w_dff_B_pQXUsDfd1_2;
	wire w_dff_B_cukDzmpN0_2;
	wire w_dff_B_aX7gAgJ73_2;
	wire w_dff_B_iS20eu445_2;
	wire w_dff_B_4kMd7Gqp5_2;
	wire w_dff_B_V5lSAUpo3_2;
	wire w_dff_B_qIBPcK4C0_2;
	wire w_dff_B_BBE16eG26_2;
	wire w_dff_B_y9eYEcky2_2;
	wire w_dff_B_0roA5NhG1_2;
	wire w_dff_B_t4qJS2Tn9_2;
	wire w_dff_B_t34YdNge6_2;
	wire w_dff_B_XWIUAX9k0_2;
	wire w_dff_B_pKQkGmkS1_2;
	wire w_dff_B_I15EsNas6_2;
	wire w_dff_B_GenIUEX24_2;
	wire w_dff_B_rbVrT2E62_2;
	wire w_dff_B_KqmLfOlG6_2;
	wire w_dff_B_8aEYebXt9_2;
	wire w_dff_B_wc1wAwBc7_2;
	wire w_dff_B_lEmWHFXi5_2;
	wire w_dff_B_qCGAblvd4_2;
	wire w_dff_B_fmOeRQYn1_2;
	wire w_dff_B_m4o2AZ9N0_2;
	wire w_dff_B_fSG9SH0t3_2;
	wire w_dff_B_BZGSdULB3_2;
	wire w_dff_B_FSimbVGz8_2;
	wire w_dff_B_4TCVkJQQ4_2;
	wire w_dff_B_dywIAmWK6_2;
	wire w_dff_B_p4sLLeAm1_2;
	wire w_dff_B_oclFPpvi7_2;
	wire w_dff_B_RnJwT5Ck2_2;
	wire w_dff_B_xUhWQ7P78_1;
	wire w_dff_B_ZnUvd0pB6_2;
	wire w_dff_B_R1LkGii23_2;
	wire w_dff_B_ue6fJH8d2_2;
	wire w_dff_B_uaUI1tya2_2;
	wire w_dff_B_e0osTeAk0_2;
	wire w_dff_B_veltr0Mk4_2;
	wire w_dff_B_8I8ntM0i4_2;
	wire w_dff_B_H8gDoiJq2_2;
	wire w_dff_B_1ZXJWgzi7_2;
	wire w_dff_B_broJSCKl3_2;
	wire w_dff_B_AF3h5rwq0_2;
	wire w_dff_B_NnnaeN9S3_2;
	wire w_dff_B_jJnSiXcb6_2;
	wire w_dff_B_0a4Am7YK2_2;
	wire w_dff_B_8cipSeC47_2;
	wire w_dff_B_54lBBl5N7_2;
	wire w_dff_B_Ky4Z5DvP9_2;
	wire w_dff_B_2ATFLZSG5_2;
	wire w_dff_B_Ge13u8Ls4_2;
	wire w_dff_B_f1glNoIf6_2;
	wire w_dff_B_1NVNZibn5_2;
	wire w_dff_B_U5N9KqAq8_2;
	wire w_dff_B_0ukPKVr16_2;
	wire w_dff_B_Kk345oQU3_2;
	wire w_dff_B_6Y6NhmMw6_2;
	wire w_dff_B_wVowZGc66_2;
	wire w_dff_B_g9yUQ3sO8_2;
	wire w_dff_B_GZN7ssAe4_2;
	wire w_dff_B_GyvGxgWo0_2;
	wire w_dff_B_TO8no1gk0_2;
	wire w_dff_B_bzHPAJfm7_2;
	wire w_dff_B_kZDfj2IH8_2;
	wire w_dff_B_ZKZeaSGl1_2;
	wire w_dff_B_jWmgzRKY9_2;
	wire w_dff_B_9yQ7bBTg6_2;
	wire w_dff_B_0laUZmpq8_2;
	wire w_dff_B_VS1icB471_2;
	wire w_dff_B_7YdJci8z9_2;
	wire w_dff_B_VyMs4l4N2_2;
	wire w_dff_B_NJPxzKL28_2;
	wire w_dff_B_RVp14ZLk4_2;
	wire w_dff_B_LZLyJm3j4_2;
	wire w_dff_B_ja0mBXim9_2;
	wire w_dff_B_Z3kybcKC3_1;
	wire w_dff_B_OPVb36m03_2;
	wire w_dff_B_9kUpg01B3_2;
	wire w_dff_B_7YnxLA981_2;
	wire w_dff_B_32w9rWTP6_2;
	wire w_dff_B_MyQzIQD49_2;
	wire w_dff_B_3O83F5zh5_2;
	wire w_dff_B_086scwRj8_2;
	wire w_dff_B_zs3gKa1G6_2;
	wire w_dff_B_0Elg8Dxi0_2;
	wire w_dff_B_hBFSUMLP1_2;
	wire w_dff_B_qr1wgGro3_2;
	wire w_dff_B_R0e5yC4e2_2;
	wire w_dff_B_QIYXvTD87_2;
	wire w_dff_B_tjnddSiO0_2;
	wire w_dff_B_Cy7Xh06B4_2;
	wire w_dff_B_nEAQQnVQ1_2;
	wire w_dff_B_UwGJbpqU0_2;
	wire w_dff_B_KIZ64XxM0_2;
	wire w_dff_B_nAeiZhqK3_2;
	wire w_dff_B_5hnQ81NF1_2;
	wire w_dff_B_ddA0HavY3_2;
	wire w_dff_B_cChozTUg5_2;
	wire w_dff_B_nL861Zk87_2;
	wire w_dff_B_54Vr9SM96_2;
	wire w_dff_B_gKcCL3Xl1_2;
	wire w_dff_B_zIRcDqcF0_2;
	wire w_dff_B_ZWSCqcPd2_2;
	wire w_dff_B_ydOqIiGX8_2;
	wire w_dff_B_tqmGzePz4_2;
	wire w_dff_B_00CjC6pd0_2;
	wire w_dff_B_zNqGBlgz3_2;
	wire w_dff_B_mBDjjgkK8_2;
	wire w_dff_B_gLRzJdOx1_2;
	wire w_dff_B_5oC21Aiy7_2;
	wire w_dff_B_iGR8yivS8_2;
	wire w_dff_B_xOLGpIMd0_2;
	wire w_dff_B_JrgDec5g1_2;
	wire w_dff_B_xoIVA3GF0_2;
	wire w_dff_B_91rMqHuE3_2;
	wire w_dff_B_WCqwlkD57_1;
	wire w_dff_B_fPiuv2cm9_2;
	wire w_dff_B_RcopoAdc6_2;
	wire w_dff_B_AZlF2ya14_2;
	wire w_dff_B_fW15ihs65_2;
	wire w_dff_B_zn8AjPi58_2;
	wire w_dff_B_NRHqG14d8_2;
	wire w_dff_B_6WgsknMI6_2;
	wire w_dff_B_8sMMocFp3_2;
	wire w_dff_B_yktOetWv2_2;
	wire w_dff_B_bvoWQD3B5_2;
	wire w_dff_B_XFc5KKgL0_2;
	wire w_dff_B_rt4W2dJk9_2;
	wire w_dff_B_fY2z0SjK8_2;
	wire w_dff_B_P7Q2Tp9n5_2;
	wire w_dff_B_TdWZf15q6_2;
	wire w_dff_B_mpEPL3kk2_2;
	wire w_dff_B_4drblbfP0_2;
	wire w_dff_B_sIZefvHT4_2;
	wire w_dff_B_OsScXjat3_2;
	wire w_dff_B_gWnmwcgo4_2;
	wire w_dff_B_9TslwpQo4_2;
	wire w_dff_B_aOYXxL9T3_2;
	wire w_dff_B_aThpX9yG3_2;
	wire w_dff_B_2tr2JhNf2_2;
	wire w_dff_B_xdjcD8ek1_2;
	wire w_dff_B_ZUBg0cdR5_2;
	wire w_dff_B_enfe3FSn1_2;
	wire w_dff_B_lWoPGZ4f7_2;
	wire w_dff_B_yOe9LVJR5_2;
	wire w_dff_B_LIjf5T790_2;
	wire w_dff_B_lBz3PMqb0_2;
	wire w_dff_B_r7CUCfbe3_2;
	wire w_dff_B_TBk6PQ0Z0_2;
	wire w_dff_B_RkwElSTr3_2;
	wire w_dff_B_gP79HKPg5_2;
	wire w_dff_B_C2oGLTtB5_1;
	wire w_dff_B_av488jlZ9_2;
	wire w_dff_B_qXkxlrXA3_2;
	wire w_dff_B_zknPNhha5_2;
	wire w_dff_B_d1irbzPu0_2;
	wire w_dff_B_lRuSyQre1_2;
	wire w_dff_B_w5oOZ97R7_2;
	wire w_dff_B_Dgu7PPXC1_2;
	wire w_dff_B_uyoNLxOB3_2;
	wire w_dff_B_zzqO8dRf2_2;
	wire w_dff_B_R4IDc1Fl4_2;
	wire w_dff_B_9Q1NfQnx7_2;
	wire w_dff_B_XUEJ55j08_2;
	wire w_dff_B_IyDbQTbd1_2;
	wire w_dff_B_IhbNuhZ40_2;
	wire w_dff_B_LJ65Cxe72_2;
	wire w_dff_B_EsacYrXN3_2;
	wire w_dff_B_ScNGK3SD7_2;
	wire w_dff_B_lk13Ztqe3_2;
	wire w_dff_B_9GJa4h0v1_2;
	wire w_dff_B_VnAcH8bm7_2;
	wire w_dff_B_gxnA3I7a1_2;
	wire w_dff_B_jfJLPkd41_2;
	wire w_dff_B_FqDvi7Zh3_2;
	wire w_dff_B_AWigrkcm2_2;
	wire w_dff_B_49wzTS1w4_2;
	wire w_dff_B_3fSRVEIg5_2;
	wire w_dff_B_3WbzAvAo2_2;
	wire w_dff_B_ct5dX4hf7_2;
	wire w_dff_B_XnLifrND1_2;
	wire w_dff_B_88iN42Kq8_2;
	wire w_dff_B_cP8Rbmyk5_2;
	wire w_dff_B_I86KhtRw2_1;
	wire w_dff_B_ju7W2gGp6_2;
	wire w_dff_B_yIS7eXoJ0_2;
	wire w_dff_B_seK5TP5Z9_2;
	wire w_dff_B_GMiotzNZ0_2;
	wire w_dff_B_HxEAuNNN4_2;
	wire w_dff_B_D41Uv9zD2_2;
	wire w_dff_B_yO5d1ktJ2_2;
	wire w_dff_B_fGhgf1iw8_2;
	wire w_dff_B_8la4JtVp2_2;
	wire w_dff_B_jE1vvOdw8_2;
	wire w_dff_B_U47nJWp36_2;
	wire w_dff_B_pHgLMOTn8_2;
	wire w_dff_B_H8y7XJcP4_2;
	wire w_dff_B_yWJydMai0_2;
	wire w_dff_B_QtzlR6zi2_2;
	wire w_dff_B_OHufHraA4_2;
	wire w_dff_B_qfwGkaqB7_2;
	wire w_dff_B_noSn6UwS4_2;
	wire w_dff_B_8lQtiQRp3_2;
	wire w_dff_B_0wOwqwwg6_2;
	wire w_dff_B_ZsPoO47b0_2;
	wire w_dff_B_tlnucIfU0_2;
	wire w_dff_B_q8hU2th87_2;
	wire w_dff_B_lFseBrOB9_2;
	wire w_dff_B_UbOE9IND1_2;
	wire w_dff_B_3uQSKymP1_2;
	wire w_dff_B_LJDxjFoi4_1;
	wire w_dff_B_08VVXDkH0_2;
	wire w_dff_B_O4F29F054_2;
	wire w_dff_B_Dmc46R6q7_2;
	wire w_dff_B_S7GON89R7_2;
	wire w_dff_B_zSLUxsei5_2;
	wire w_dff_B_YDt6z6cg9_2;
	wire w_dff_B_M1yvTjJl5_2;
	wire w_dff_B_az8E3v9g6_2;
	wire w_dff_B_tAq2IbZl3_2;
	wire w_dff_B_J5e5KFVe2_2;
	wire w_dff_B_lTrmwefs6_2;
	wire w_dff_B_7AByAONw9_2;
	wire w_dff_B_ILkibUJj7_2;
	wire w_dff_B_WtOB8IT22_2;
	wire w_dff_B_ZzF7ou968_2;
	wire w_dff_B_V6qDCgDl4_2;
	wire w_dff_B_IoDUvnMM0_2;
	wire w_dff_B_CdBOnoWr5_2;
	wire w_dff_B_HA0nb6ci8_2;
	wire w_dff_B_rvlZNm1Z6_2;
	wire w_dff_B_K72b4cU16_2;
	wire w_dff_B_qNrSSy3u2_2;
	wire w_dff_B_QUpBqD0A6_2;
	wire w_dff_B_72tu2LAE3_2;
	wire w_dff_B_5mHjtuOZ5_1;
	wire w_dff_B_73sBYgZK7_2;
	wire w_dff_B_HXBvKebs7_2;
	wire w_dff_B_NmKTxOY83_2;
	wire w_dff_B_ZqNRnkbi7_2;
	wire w_dff_B_cBfevwWd8_2;
	wire w_dff_B_QR1ydtWC1_2;
	wire w_dff_B_eO9swGgq0_2;
	wire w_dff_B_2iXHiTP31_2;
	wire w_dff_B_VXM7YLfv8_2;
	wire w_dff_B_ythenOWD3_2;
	wire w_dff_B_Pdn9LChg6_2;
	wire w_dff_B_m4jRz59K9_2;
	wire w_dff_B_EAkevS0z0_2;
	wire w_dff_B_2kJUwQqd0_2;
	wire w_dff_B_NJbB9n1W7_2;
	wire w_dff_B_iSHyyvDm5_2;
	wire w_dff_B_8wbRfNYU4_2;
	wire w_dff_B_YVpeK3cy7_2;
	wire w_dff_B_h00hxkZJ6_2;
	wire w_dff_B_wQxdIANl7_2;
	wire w_dff_B_bXuZ2R9U2_2;
	wire w_dff_B_QNM7Qz8B1_1;
	wire w_dff_B_DxcT5UY99_2;
	wire w_dff_B_BTaoT8Xu8_2;
	wire w_dff_B_fGl5cl8s6_2;
	wire w_dff_B_7ppeqsrN5_2;
	wire w_dff_B_vj44D1I42_2;
	wire w_dff_B_0G1sA9Pt8_2;
	wire w_dff_B_DLbnZe7g7_2;
	wire w_dff_B_8VQDqMGD3_2;
	wire w_dff_B_tgA1Zv524_2;
	wire w_dff_B_bS3Fn67k7_2;
	wire w_dff_B_7gA6ZETQ1_2;
	wire w_dff_B_khCf8RYj8_2;
	wire w_dff_B_c0iKoziR7_2;
	wire w_dff_B_ZghivQ114_2;
	wire w_dff_B_5Z0tHiZu1_2;
	wire w_dff_B_iPUyH3sg7_2;
	wire w_dff_B_0fgYsl7M7_2;
	wire w_dff_B_FbDURwN55_2;
	wire w_dff_B_w6HJXtga9_1;
	wire w_dff_B_vtMewbRc0_2;
	wire w_dff_B_cX7EzFbw1_2;
	wire w_dff_B_oG3RKuPe3_2;
	wire w_dff_B_Uy5KFX1F9_2;
	wire w_dff_B_S6rwYapD8_2;
	wire w_dff_B_kzjhLKBF6_2;
	wire w_dff_B_92IMJ7ZM2_2;
	wire w_dff_B_iUbH7IrW8_2;
	wire w_dff_B_FvDLb4XM7_2;
	wire w_dff_B_qWN1ySMt7_2;
	wire w_dff_B_I145K9kq6_2;
	wire w_dff_B_2XSfBDqh9_2;
	wire w_dff_B_7BEK49uK1_2;
	wire w_dff_B_VfNDgjQa5_2;
	wire w_dff_B_bFThtfdB8_2;
	wire w_dff_B_zz5olJJm3_1;
	wire w_dff_B_mOWuvJG62_2;
	wire w_dff_B_WieyFUj92_2;
	wire w_dff_B_oJvtDd4k6_2;
	wire w_dff_B_VEVvxzre2_2;
	wire w_dff_B_IOgruZrP8_2;
	wire w_dff_B_cwBUrJLP2_2;
	wire w_dff_B_BERuTnDO0_2;
	wire w_dff_B_9RCoXGYh5_2;
	wire w_dff_B_cGp6XCah9_2;
	wire w_dff_B_dS5O7xwN9_2;
	wire w_dff_B_4ShqpVAq3_2;
	wire w_dff_B_5E2IGDSn9_2;
	wire w_dff_B_KaaAk79D5_1;
	wire w_dff_B_yF3ObJhE0_2;
	wire w_dff_B_BjUNqUy12_2;
	wire w_dff_B_NzqfFX740_2;
	wire w_dff_B_vte77m381_2;
	wire w_dff_B_HohZjWKK4_2;
	wire w_dff_B_7HnIj5zW7_2;
	wire w_dff_B_hQK9vWSi7_2;
	wire w_dff_B_AxdmzWHQ1_2;
	wire w_dff_B_iCsp48My5_2;
	wire w_dff_B_HA8qc1Lm5_2;
	wire w_dff_B_P00s8lh91_2;
	wire w_dff_B_dwgyX0h69_1;
	wire w_dff_B_B7jVbXwV8_1;
	wire w_dff_B_MJ3UurQN6_2;
	wire w_dff_B_OZfCZq0z4_2;
	wire w_dff_B_x2wZXyLI6_2;
	wire w_dff_B_CPt8EioO4_0;
	wire w_dff_A_WpIMPUUK4_0;
	wire w_dff_A_ddDRVV2g5_0;
	wire w_dff_A_Cvr6BZlL8_1;
	wire w_dff_A_u7HtRnIt1_1;
	wire w_dff_B_rnOokL9a0_1;
	wire w_dff_B_eemYFfZE1_1;
	wire w_dff_B_qoKI2Mw54_1;
	wire w_dff_B_fekuKRv69_2;
	wire w_dff_B_6o46UZoJ2_2;
	wire w_dff_B_ScWcUdbH1_2;
	wire w_dff_B_Fza23mTq3_2;
	wire w_dff_B_FKB9wtSE6_2;
	wire w_dff_B_pwQQ3Vxg0_2;
	wire w_dff_B_OSw2XQzE6_2;
	wire w_dff_B_8h2JOS4D1_2;
	wire w_dff_B_iSK38hw75_2;
	wire w_dff_B_SuNKY6o98_2;
	wire w_dff_B_WfFvJ3ds6_2;
	wire w_dff_B_YYfaUxtK7_2;
	wire w_dff_B_dYkhZAQ05_2;
	wire w_dff_B_UhWBAowR8_2;
	wire w_dff_B_3ogD9THR8_2;
	wire w_dff_B_1iM6xSUK3_2;
	wire w_dff_B_LbN90txj0_2;
	wire w_dff_B_HHx7ipqQ8_2;
	wire w_dff_B_V540786e0_2;
	wire w_dff_B_ylMcfni99_2;
	wire w_dff_B_cfL4g4H03_2;
	wire w_dff_B_waiXJdWJ2_2;
	wire w_dff_B_VjQ6fMhN5_2;
	wire w_dff_B_tpLpNfts2_2;
	wire w_dff_B_Et7EwVPd9_2;
	wire w_dff_B_UJCaMQ2l8_2;
	wire w_dff_B_54nb5RJS4_2;
	wire w_dff_B_ncsG6zO35_2;
	wire w_dff_B_AgJoGb7q0_2;
	wire w_dff_B_Dheq6hcl7_2;
	wire w_dff_B_EC1RA1He8_2;
	wire w_dff_B_i06ei0xs0_2;
	wire w_dff_B_32qNexT32_2;
	wire w_dff_B_A61xT71d8_2;
	wire w_dff_B_iepEY6QA4_2;
	wire w_dff_B_bfsOVy8W7_2;
	wire w_dff_B_F1O6xQX38_2;
	wire w_dff_B_XafBI5KU8_2;
	wire w_dff_B_V5ZrDsEz6_2;
	wire w_dff_B_fygMFRAS3_2;
	wire w_dff_B_BoMWUDut6_2;
	wire w_dff_B_VskeT8Gn3_2;
	wire w_dff_B_mfIE8pPi6_2;
	wire w_dff_B_oQAX6XgK2_2;
	wire w_dff_B_1tYcAu7d7_2;
	wire w_dff_B_iS8DQAJU4_2;
	wire w_dff_B_LD8x03BM6_2;
	wire w_dff_B_eiY4043F5_2;
	wire w_dff_B_yqGLUhTl0_2;
	wire w_dff_B_XsNfQcA90_2;
	wire w_dff_B_kHmAAaLS5_2;
	wire w_dff_B_GzkyVSpP2_2;
	wire w_dff_B_qbkifT6e7_2;
	wire w_dff_B_wHex4ErG5_2;
	wire w_dff_B_NRorvn3D1_2;
	wire w_dff_B_dnrhKfRz2_2;
	wire w_dff_B_iKSGlt2k2_2;
	wire w_dff_B_6KZtI9BN5_2;
	wire w_dff_B_BxohSfVY3_2;
	wire w_dff_B_hUDzoFWI9_2;
	wire w_dff_B_ISFZ6qAj6_2;
	wire w_dff_B_bZoKpMmg6_2;
	wire w_dff_B_ikxFmEcE1_2;
	wire w_dff_B_FcWayhaS9_2;
	wire w_dff_B_vQ8lOx3G1_2;
	wire w_dff_B_0dp8mov36_2;
	wire w_dff_B_sFdmXqkX9_2;
	wire w_dff_B_WF8y5fMJ1_2;
	wire w_dff_B_qq8b4wp45_2;
	wire w_dff_B_KQBaWEgq6_2;
	wire w_dff_B_euyVptgE5_2;
	wire w_dff_B_7pfLpn5v1_2;
	wire w_dff_B_fOGfCDcD5_2;
	wire w_dff_B_8hIqXpWi8_2;
	wire w_dff_B_9P8HEvje1_2;
	wire w_dff_B_HJ92Qrpr8_2;
	wire w_dff_B_e6rj65kD3_2;
	wire w_dff_B_4TqLvPoB2_2;
	wire w_dff_B_mXqIyH7B0_2;
	wire w_dff_B_rCTg4omV4_2;
	wire w_dff_B_6CKiChEE0_2;
	wire w_dff_B_J3iEX8oP7_2;
	wire w_dff_B_x11pYp299_2;
	wire w_dff_B_fqSX8xtR7_2;
	wire w_dff_B_aoLxrmVu7_2;
	wire w_dff_B_l2MwQBq36_2;
	wire w_dff_B_yWm41cbh2_2;
	wire w_dff_B_4ft1bbLm8_2;
	wire w_dff_B_SlnWQCht9_2;
	wire w_dff_B_aMCSR9bf3_2;
	wire w_dff_B_8GYIJnRQ1_2;
	wire w_dff_B_TJeub2rC8_2;
	wire w_dff_B_LlKDU5qL8_2;
	wire w_dff_B_3EcdPy3h2_2;
	wire w_dff_B_2MbxBxlc8_2;
	wire w_dff_B_47rlAOQB2_2;
	wire w_dff_B_oG65F0kM0_2;
	wire w_dff_B_PydkgQ309_2;
	wire w_dff_B_R0FdWsCi9_2;
	wire w_dff_B_PPUprleU2_2;
	wire w_dff_B_wCvOxZcE8_2;
	wire w_dff_B_qlLGs09n3_2;
	wire w_dff_B_J06WYYku7_2;
	wire w_dff_B_LYMiaIjV0_2;
	wire w_dff_B_3BcFTCck0_2;
	wire w_dff_B_24wYAHYp0_2;
	wire w_dff_B_w5zeJbcK1_2;
	wire w_dff_B_h5KCZ1I58_2;
	wire w_dff_A_AC3zetFj0_1;
	wire w_dff_B_85yW5gdO3_1;
	wire w_dff_B_8WF4KYqn5_2;
	wire w_dff_B_Jqn8uaQ92_2;
	wire w_dff_B_jy7C6HWf9_2;
	wire w_dff_B_Cy9GJQgW8_2;
	wire w_dff_B_CCiXw2dm0_2;
	wire w_dff_B_QMlT8fwp8_2;
	wire w_dff_B_UUOvCZ546_2;
	wire w_dff_B_uDvz2kqa7_2;
	wire w_dff_B_SsU40btC3_2;
	wire w_dff_B_a9aTANtB6_2;
	wire w_dff_B_vcyrLHtu7_2;
	wire w_dff_B_h5Efwqro5_2;
	wire w_dff_B_orAWzWoQ9_2;
	wire w_dff_B_CRQ6lrv31_2;
	wire w_dff_B_cDd7MEgJ8_2;
	wire w_dff_B_3HYPkTbX3_2;
	wire w_dff_B_BwZAt3Ko7_2;
	wire w_dff_B_ufmYqBUq7_2;
	wire w_dff_B_71L3SUDj8_2;
	wire w_dff_B_iAicqo8d6_2;
	wire w_dff_B_AM2GkTIl7_2;
	wire w_dff_B_zo6ENjUE4_2;
	wire w_dff_B_PD0ftZX28_2;
	wire w_dff_B_AUJz5OWt4_2;
	wire w_dff_B_VTBdWyW88_2;
	wire w_dff_B_nMBamYQy4_2;
	wire w_dff_B_9CqUlWIl8_2;
	wire w_dff_B_FM4MBQ361_2;
	wire w_dff_B_QoMGX0Ri1_2;
	wire w_dff_B_OJdxKCF99_2;
	wire w_dff_B_wS5SBU8a9_2;
	wire w_dff_B_Bs5Fozd86_2;
	wire w_dff_B_Gn2uyNUh3_2;
	wire w_dff_B_VQ9xYquK1_2;
	wire w_dff_B_lPksMeCS9_2;
	wire w_dff_B_MbFSliPR3_2;
	wire w_dff_B_yTXCb2XC6_2;
	wire w_dff_B_3ln4MD2j3_2;
	wire w_dff_B_57X8Wt5L5_2;
	wire w_dff_B_TBi551Nz5_2;
	wire w_dff_B_lHpg4irN2_2;
	wire w_dff_B_Eg0KSJP98_2;
	wire w_dff_B_2Jy3gg3s6_2;
	wire w_dff_B_o7E4ISy59_2;
	wire w_dff_B_ltad0Hjn0_2;
	wire w_dff_B_uJO1sXxd1_2;
	wire w_dff_B_T5uxMaiV8_2;
	wire w_dff_B_033E9Cvb2_2;
	wire w_dff_B_OHakaALJ9_2;
	wire w_dff_B_8vHTzRsX1_2;
	wire w_dff_B_gRltySca3_2;
	wire w_dff_B_2CXTIugB1_2;
	wire w_dff_B_HQF7bk0e2_1;
	wire w_dff_B_RPpjFPI81_1;
	wire w_dff_B_z32vzuen8_2;
	wire w_dff_B_2TxosvpK4_2;
	wire w_dff_B_2zP9rxji0_2;
	wire w_dff_B_tWO7PmSc9_2;
	wire w_dff_B_WlMbHSGw4_2;
	wire w_dff_B_FpxiYoBb8_2;
	wire w_dff_B_Dbvpant06_2;
	wire w_dff_B_0FjwZUAB1_2;
	wire w_dff_B_2ULonY1o0_2;
	wire w_dff_B_G8sLIlY88_2;
	wire w_dff_B_fcjllQOJ1_2;
	wire w_dff_B_yEW0P7HF4_2;
	wire w_dff_B_s8ylfpqX8_2;
	wire w_dff_B_MV29CfLk2_2;
	wire w_dff_B_DX3fr6qb6_2;
	wire w_dff_B_tlRlAHoH7_2;
	wire w_dff_B_9L95tK7M0_2;
	wire w_dff_B_QYeBX5YM1_2;
	wire w_dff_B_TCHWB0M38_2;
	wire w_dff_B_aVZyOHo32_2;
	wire w_dff_B_X8OHSapp3_2;
	wire w_dff_B_PYYePxEZ2_2;
	wire w_dff_B_0Zw2sFuo4_2;
	wire w_dff_B_hzZt9EVf5_2;
	wire w_dff_B_JvyXTsTy1_2;
	wire w_dff_B_5darSBRX8_2;
	wire w_dff_B_1GVf5QKc6_2;
	wire w_dff_B_5D241waB4_2;
	wire w_dff_B_cWtCDbYR5_2;
	wire w_dff_B_veMo1N1j1_2;
	wire w_dff_B_0iGAMoMH3_2;
	wire w_dff_B_OlQFWA1y7_2;
	wire w_dff_B_dkUO5tex3_2;
	wire w_dff_B_KHPZNq1z4_2;
	wire w_dff_B_uVHk9e7I4_2;
	wire w_dff_B_FFAQXH8y8_2;
	wire w_dff_B_HkgoVjKt2_2;
	wire w_dff_B_MS9o8qbU7_2;
	wire w_dff_B_rXqxLoeU5_2;
	wire w_dff_B_KHyzEeXE7_2;
	wire w_dff_B_k6RKacYf8_2;
	wire w_dff_B_kwa01AcH7_2;
	wire w_dff_B_iAwdxS9e9_2;
	wire w_dff_B_rWMhrAY43_2;
	wire w_dff_B_WDx2Oece0_2;
	wire w_dff_B_LHhYusnr3_2;
	wire w_dff_B_mG0hsKCn9_2;
	wire w_dff_B_1ULdHyqg5_2;
	wire w_dff_B_shCeCe4X9_2;
	wire w_dff_B_38XHFW1a0_2;
	wire w_dff_B_6l6LmxGh8_2;
	wire w_dff_B_pBxWMLd88_2;
	wire w_dff_B_VXmyVpwX6_2;
	wire w_dff_B_IdiO4bbN6_2;
	wire w_dff_B_NmtiALd18_2;
	wire w_dff_B_ao1mXhxw2_2;
	wire w_dff_B_ZbBMZt8j7_2;
	wire w_dff_B_kk0Uvfm58_2;
	wire w_dff_B_lZPcH5UB8_2;
	wire w_dff_B_ArcWtZyl0_2;
	wire w_dff_B_Ei18dZBy1_2;
	wire w_dff_B_mNppE8HK5_2;
	wire w_dff_B_1cqeLFF82_2;
	wire w_dff_B_gjrizHwI6_2;
	wire w_dff_B_Nr7qpHFG9_2;
	wire w_dff_B_Tp75y8Qm0_2;
	wire w_dff_B_uulUz8c12_2;
	wire w_dff_B_xBauWA2G6_2;
	wire w_dff_B_ueKq4WmA4_2;
	wire w_dff_B_nLC5pjLh4_2;
	wire w_dff_B_fNwM23435_2;
	wire w_dff_B_UoJcFxZb4_2;
	wire w_dff_B_hHUbooTL0_2;
	wire w_dff_B_t6v06zX06_2;
	wire w_dff_B_m4yMbSoz3_2;
	wire w_dff_B_p9bNeZhd7_2;
	wire w_dff_B_xDLC4G8i6_2;
	wire w_dff_B_Acwt59K28_2;
	wire w_dff_B_QQ75cPNx1_2;
	wire w_dff_B_BOTMtTsc3_2;
	wire w_dff_B_JwATBW8Q0_2;
	wire w_dff_B_l4CR5KVy8_2;
	wire w_dff_B_PVYLwQFE2_2;
	wire w_dff_B_1Epdjbom5_2;
	wire w_dff_B_L93FNHMi3_2;
	wire w_dff_B_EZ7VocIB0_2;
	wire w_dff_B_puR35NMM1_2;
	wire w_dff_B_5ePNdsAh0_2;
	wire w_dff_B_d7n0X0my4_2;
	wire w_dff_B_jWC2VfwL4_2;
	wire w_dff_B_HZj48SdY2_2;
	wire w_dff_B_49podTqW6_2;
	wire w_dff_B_XmgPat7m5_2;
	wire w_dff_B_uokwtuQD7_2;
	wire w_dff_B_OsJdbdGz5_2;
	wire w_dff_B_VPkaGOVS6_2;
	wire w_dff_B_deH8Th2h3_2;
	wire w_dff_B_UGOBmCau4_2;
	wire w_dff_B_7d4n6SbI0_2;
	wire w_dff_B_3OSCaDKz1_2;
	wire w_dff_B_8KA5KVCB4_2;
	wire w_dff_B_qWUxsDRZ7_1;
	wire w_dff_B_xD076iXe6_2;
	wire w_dff_B_kyesZ4rs8_2;
	wire w_dff_B_oik7KltN4_2;
	wire w_dff_B_e5tzgqE57_2;
	wire w_dff_B_oKcMerhe6_2;
	wire w_dff_B_Vryh36YB6_2;
	wire w_dff_B_6xBYqasI9_2;
	wire w_dff_B_19wc5L0r5_2;
	wire w_dff_B_aEX32HKi5_2;
	wire w_dff_B_sqvRMQzC6_2;
	wire w_dff_B_RSfjmcyd9_2;
	wire w_dff_B_gqbnx4fx0_2;
	wire w_dff_B_qJCpyv0l2_2;
	wire w_dff_B_M9aDvJwx7_2;
	wire w_dff_B_Y1ZmAn6a6_2;
	wire w_dff_B_9fo6GBzZ7_2;
	wire w_dff_B_82v8wYhk2_2;
	wire w_dff_B_um04Y1dA1_2;
	wire w_dff_B_fd7C7USc6_2;
	wire w_dff_B_G3UktORU8_2;
	wire w_dff_B_fH7pNbZu5_2;
	wire w_dff_B_WKNN1m8k1_2;
	wire w_dff_B_p3qWDmPL3_2;
	wire w_dff_B_lCPAivWe7_2;
	wire w_dff_B_DhRAhByB2_2;
	wire w_dff_B_VIdwCA4l9_2;
	wire w_dff_B_6MPY2VgM1_2;
	wire w_dff_B_zNWNzSBz5_2;
	wire w_dff_B_j9BTXpGQ8_2;
	wire w_dff_B_59sPQ6fC3_2;
	wire w_dff_B_GBHLQwtx8_2;
	wire w_dff_B_InKxkVFR3_2;
	wire w_dff_B_ow5G3P7x5_2;
	wire w_dff_B_XL2a7IEz7_2;
	wire w_dff_B_NGDDQFOp9_2;
	wire w_dff_B_sRVDEl1N3_2;
	wire w_dff_B_xrPVKBRL4_2;
	wire w_dff_B_qIUimjEC6_2;
	wire w_dff_B_LowstA8A8_2;
	wire w_dff_B_sC89UURm6_2;
	wire w_dff_B_yoHj2H7U8_2;
	wire w_dff_B_adlzWLRy3_2;
	wire w_dff_B_epf9saWp2_2;
	wire w_dff_B_Weh4jPJS0_2;
	wire w_dff_B_gRug1Bad9_2;
	wire w_dff_B_I6IYIYEb0_2;
	wire w_dff_B_DevLermn5_2;
	wire w_dff_B_12hr5EGl3_2;
	wire w_dff_B_CWGCbJ0w0_1;
	wire w_dff_B_d4ZAE1QM3_1;
	wire w_dff_B_faJ9xdeC4_2;
	wire w_dff_B_nF5ANBtQ5_2;
	wire w_dff_B_C0XUzrGO1_2;
	wire w_dff_B_yM3dHu371_2;
	wire w_dff_B_qsKw82EM9_2;
	wire w_dff_B_qY83BAly6_2;
	wire w_dff_B_Jwc7aw7h2_2;
	wire w_dff_B_8t6SukKM3_2;
	wire w_dff_B_lZXZY2CY6_2;
	wire w_dff_B_E6XZIp867_2;
	wire w_dff_B_ivekI5sQ4_2;
	wire w_dff_B_cqHO71de8_2;
	wire w_dff_B_QD0UR4Vz9_2;
	wire w_dff_B_RV1zZGpt4_2;
	wire w_dff_B_s7RlcEsX7_2;
	wire w_dff_B_J44t7Nwn4_2;
	wire w_dff_B_Y3jwTgdq1_2;
	wire w_dff_B_sbN9BVqF3_2;
	wire w_dff_B_hWWuQbSl0_2;
	wire w_dff_B_AphpyBUy8_2;
	wire w_dff_B_j50asqdf6_2;
	wire w_dff_B_HjQi7iLm1_2;
	wire w_dff_B_FGXlemH91_2;
	wire w_dff_B_Eb0oQOHA8_2;
	wire w_dff_B_abzWY0ir1_2;
	wire w_dff_B_hat5Xztu7_2;
	wire w_dff_B_NoUV1BRL3_2;
	wire w_dff_B_W50ncMDH3_2;
	wire w_dff_B_st73XXd01_2;
	wire w_dff_B_36MSZ6Yb8_2;
	wire w_dff_B_zVlBygQ15_2;
	wire w_dff_B_wFXBDUk77_2;
	wire w_dff_B_3R4mOfJH5_2;
	wire w_dff_B_wO8axMbp6_2;
	wire w_dff_B_MSlP7h3A3_2;
	wire w_dff_B_m21HxMrG0_2;
	wire w_dff_B_VhroFn5w0_2;
	wire w_dff_B_oBLqhJkX1_2;
	wire w_dff_B_HUoWclQQ1_2;
	wire w_dff_B_rrvRyZfs8_2;
	wire w_dff_B_cHFib2jT1_2;
	wire w_dff_B_C1kslyPO6_2;
	wire w_dff_B_mgDUfXp27_2;
	wire w_dff_B_fGsuuLXw7_2;
	wire w_dff_B_chfeBSJ11_2;
	wire w_dff_B_2EAVDkLl7_2;
	wire w_dff_B_ngLYd4XY5_2;
	wire w_dff_B_gzg6flQI8_2;
	wire w_dff_B_R4yFSMeE1_2;
	wire w_dff_B_YdBBbARr4_2;
	wire w_dff_B_avlYpuqv7_2;
	wire w_dff_B_bGdUGE8j5_2;
	wire w_dff_B_umVXL3Dw4_2;
	wire w_dff_B_jI5YRURc6_2;
	wire w_dff_B_7XKxpy8r3_2;
	wire w_dff_B_jKJ5sE8T3_2;
	wire w_dff_B_Hk7b3xWK1_2;
	wire w_dff_B_ew6PZ2WT2_2;
	wire w_dff_B_4eQudNhd7_2;
	wire w_dff_B_VrgPTmQO6_2;
	wire w_dff_B_GQEYkhqY1_2;
	wire w_dff_B_cVhU0I1q0_2;
	wire w_dff_B_ymzaI4fb8_2;
	wire w_dff_B_7iL8PC3L6_2;
	wire w_dff_B_OhBTwph58_2;
	wire w_dff_B_MIx31jh04_2;
	wire w_dff_B_9Qko8Pqy1_2;
	wire w_dff_B_IrmeGxQh5_2;
	wire w_dff_B_10HN8qt34_2;
	wire w_dff_B_FPoNjL1f0_2;
	wire w_dff_B_Ql9V8Nh02_2;
	wire w_dff_B_eZlUtsJ09_2;
	wire w_dff_B_GUQEn7xA6_2;
	wire w_dff_B_fWE6NGUT7_2;
	wire w_dff_B_7TruB4oG3_2;
	wire w_dff_B_0kioKlY41_2;
	wire w_dff_B_tJtqcomJ2_2;
	wire w_dff_B_0hdK8N0n6_2;
	wire w_dff_B_kuez1BPk2_2;
	wire w_dff_B_egoPkZ047_2;
	wire w_dff_B_e3ktsPK58_2;
	wire w_dff_B_yGNuGTbC4_2;
	wire w_dff_B_RO0r7OBj8_2;
	wire w_dff_B_1Z4GYRlm9_2;
	wire w_dff_B_apBpyLGa3_2;
	wire w_dff_B_1Kk16XHi5_2;
	wire w_dff_B_n1TXBwYX3_2;
	wire w_dff_B_LrNu2tmv7_2;
	wire w_dff_B_gvhiwkz56_2;
	wire w_dff_B_mJ3gr90N8_2;
	wire w_dff_B_srHe9ezn4_2;
	wire w_dff_B_t3UUnhQ63_2;
	wire w_dff_B_j4DIVSxT5_2;
	wire w_dff_B_1cUf0YGg3_1;
	wire w_dff_B_fYLZYovA4_2;
	wire w_dff_B_vSbmGcqz5_2;
	wire w_dff_B_jQbvSLKP1_2;
	wire w_dff_B_gszgBOQm4_2;
	wire w_dff_B_RuqD6PyM5_2;
	wire w_dff_B_52HjBxyi4_2;
	wire w_dff_B_NRd8nkEE1_2;
	wire w_dff_B_sN5CeOlZ1_2;
	wire w_dff_B_PIYKBRiq6_2;
	wire w_dff_B_VfWB5LxK4_2;
	wire w_dff_B_sKybOTp39_2;
	wire w_dff_B_ApqATlrs4_2;
	wire w_dff_B_mr0OaWUT2_2;
	wire w_dff_B_ARTueBT24_2;
	wire w_dff_B_6KuKY68J7_2;
	wire w_dff_B_hk87IMgY3_2;
	wire w_dff_B_887I8Jxa2_2;
	wire w_dff_B_yZjRqMe42_2;
	wire w_dff_B_NM0Y1hWn2_2;
	wire w_dff_B_CGQvG3yf8_2;
	wire w_dff_B_FBwPxAJx6_2;
	wire w_dff_B_Cd4ay4Wa8_2;
	wire w_dff_B_q8ta6jqp4_2;
	wire w_dff_B_iU8oq5SF4_2;
	wire w_dff_B_WcSJHpsH8_2;
	wire w_dff_B_sqHZn5su3_2;
	wire w_dff_B_6UbglX4O2_2;
	wire w_dff_B_UxQgDpqq2_2;
	wire w_dff_B_TYNlJLSn7_2;
	wire w_dff_B_HhpQE4kW9_2;
	wire w_dff_B_VVfQdY1B5_2;
	wire w_dff_B_Mf1IWDy81_2;
	wire w_dff_B_ZzQJFCZZ6_2;
	wire w_dff_B_UQ776D743_2;
	wire w_dff_B_VMc7Faea5_2;
	wire w_dff_B_xB2zWgPK7_2;
	wire w_dff_B_KjwqDgQE0_2;
	wire w_dff_B_UaOu27yt3_2;
	wire w_dff_B_E0t5ECdE0_2;
	wire w_dff_B_E1e5RC7n4_2;
	wire w_dff_B_B1p262JB2_2;
	wire w_dff_B_a4Ke2SEk4_2;
	wire w_dff_B_lRuyGLG24_2;
	wire w_dff_B_CBStuMlU2_2;
	wire w_dff_B_MOifhJCc8_1;
	wire w_dff_B_lVWo6LPI0_1;
	wire w_dff_B_W1fImlgg1_2;
	wire w_dff_B_gy0E2syy4_2;
	wire w_dff_B_8ILM1cof0_2;
	wire w_dff_B_XUi5sFrJ6_2;
	wire w_dff_B_kpE5Vyk67_2;
	wire w_dff_B_5qnMg1bU9_2;
	wire w_dff_B_ziY8UmGG3_2;
	wire w_dff_B_jXk44IW77_2;
	wire w_dff_B_xBNwlM3J6_2;
	wire w_dff_B_xhbjBwyY2_2;
	wire w_dff_B_QOnKBiC72_2;
	wire w_dff_B_GiLeXQaB9_2;
	wire w_dff_B_CbburaLq0_2;
	wire w_dff_B_7c29jQdE0_2;
	wire w_dff_B_KssGcenL7_2;
	wire w_dff_B_ujDKBUXA5_2;
	wire w_dff_B_Xq3z0dH93_2;
	wire w_dff_B_vWFAv8EE2_2;
	wire w_dff_B_D5Uwx2WR9_2;
	wire w_dff_B_7MqjbenK8_2;
	wire w_dff_B_cdfS37n29_2;
	wire w_dff_B_LH8nCjx98_2;
	wire w_dff_B_BA4Bn5JB6_2;
	wire w_dff_B_y1TIZDIi7_2;
	wire w_dff_B_hjIWMQYH1_2;
	wire w_dff_B_enC1StP34_2;
	wire w_dff_B_cVEEZnhd5_2;
	wire w_dff_B_6aTtpjm30_2;
	wire w_dff_B_59GPI1Sd1_2;
	wire w_dff_B_hhpnrpPS4_2;
	wire w_dff_B_HOyvwsa40_2;
	wire w_dff_B_9gvnNtA70_2;
	wire w_dff_B_2S7GHZ3H9_2;
	wire w_dff_B_owyP0Yx30_2;
	wire w_dff_B_tCP1VM0J5_2;
	wire w_dff_B_1gNVAssC9_2;
	wire w_dff_B_rZ9LUbfm1_2;
	wire w_dff_B_bELAnydM6_2;
	wire w_dff_B_kyT5jDZT2_2;
	wire w_dff_B_mWxr1naH6_2;
	wire w_dff_B_Cy9xGHOQ5_2;
	wire w_dff_B_NDQiaCOP5_2;
	wire w_dff_B_zte6Kcty8_2;
	wire w_dff_B_pLwJsyDp8_2;
	wire w_dff_B_n1SXt6eE9_2;
	wire w_dff_B_PYuac0zV5_2;
	wire w_dff_B_G83IlmWl6_2;
	wire w_dff_B_EHe0aV8Q0_2;
	wire w_dff_B_3IGIPZVt7_2;
	wire w_dff_B_jucUOgts6_2;
	wire w_dff_B_OxboZAsz4_2;
	wire w_dff_B_tUqE9xah2_2;
	wire w_dff_B_GyA2b7Tc5_2;
	wire w_dff_B_cogp0iZV3_2;
	wire w_dff_B_dfHMjl051_2;
	wire w_dff_B_N8NCNmHB5_2;
	wire w_dff_B_F6Vzk1BR9_2;
	wire w_dff_B_0aaFObD03_2;
	wire w_dff_B_ezSLIK7a4_2;
	wire w_dff_B_7MPW1RIy8_2;
	wire w_dff_B_k6dWuvBb1_2;
	wire w_dff_B_rI2td8W11_2;
	wire w_dff_B_NeLpJ9J22_2;
	wire w_dff_B_5i5q6OnL2_2;
	wire w_dff_B_Zc8aYGpA9_2;
	wire w_dff_B_lLdbZKoH9_2;
	wire w_dff_B_3eWry5JS6_2;
	wire w_dff_B_FLlRzHmu3_2;
	wire w_dff_B_EDf6ugCK0_2;
	wire w_dff_B_9wvPUEAv1_2;
	wire w_dff_B_yFTwmcv21_2;
	wire w_dff_B_anBSeP584_2;
	wire w_dff_B_PjVOV9nZ7_2;
	wire w_dff_B_6Ldbww9W2_2;
	wire w_dff_B_riiEll2j1_2;
	wire w_dff_B_mppRzF617_2;
	wire w_dff_B_Qseosek06_2;
	wire w_dff_B_J2fetmqx3_2;
	wire w_dff_B_S6MH5rPa7_2;
	wire w_dff_B_j7uGJMBe1_2;
	wire w_dff_B_MloNm4do6_2;
	wire w_dff_B_9KOoqiZj9_2;
	wire w_dff_B_rkl99rgz3_2;
	wire w_dff_B_hmcBy8Y75_2;
	wire w_dff_B_rttDH4w78_2;
	wire w_dff_B_SN63Z6ww0_1;
	wire w_dff_B_2w8MVoH53_2;
	wire w_dff_B_e46VTKop9_2;
	wire w_dff_B_LSisNa268_2;
	wire w_dff_B_oFCdudBJ2_2;
	wire w_dff_B_2DjnVYRp1_2;
	wire w_dff_B_ssWz4MEp5_2;
	wire w_dff_B_of32stQY3_2;
	wire w_dff_B_XHpujecB2_2;
	wire w_dff_B_zWPvtu2x9_2;
	wire w_dff_B_W2e9vhvR8_2;
	wire w_dff_B_8gKzIHv56_2;
	wire w_dff_B_ZFsO7iqZ2_2;
	wire w_dff_B_YON7aJgk8_2;
	wire w_dff_B_wC2KjiuU5_2;
	wire w_dff_B_b7JHQl2A4_2;
	wire w_dff_B_2kGRweaU6_2;
	wire w_dff_B_42bTzYJ90_2;
	wire w_dff_B_FxxJ7s439_2;
	wire w_dff_B_VGKt2nH15_2;
	wire w_dff_B_eWXal43W1_2;
	wire w_dff_B_czxxPufb9_2;
	wire w_dff_B_LQTbmUYy2_2;
	wire w_dff_B_nIXyuSJv5_2;
	wire w_dff_B_1Vojf63D9_2;
	wire w_dff_B_2z0zJWmN0_2;
	wire w_dff_B_1q4wkFhO8_2;
	wire w_dff_B_fm9r7YsV2_2;
	wire w_dff_B_BYvTr5Qp6_2;
	wire w_dff_B_WNFPVwXA5_2;
	wire w_dff_B_sUnW1Sx40_2;
	wire w_dff_B_kgzbo2OC7_2;
	wire w_dff_B_VZgp7J896_2;
	wire w_dff_B_cIbOwcwU2_2;
	wire w_dff_B_bKuJ5P6R3_2;
	wire w_dff_B_f1dZ6x8c1_2;
	wire w_dff_B_1DOe9Pgg1_2;
	wire w_dff_B_U28oDTfI7_2;
	wire w_dff_B_qBi4lIwq1_2;
	wire w_dff_B_ZjWGrG8E2_2;
	wire w_dff_B_hWflD2Rx4_2;
	wire w_dff_B_dQiY6pmy6_1;
	wire w_dff_B_O32QGbkt5_1;
	wire w_dff_B_RClOnliE9_2;
	wire w_dff_B_cz818Th53_2;
	wire w_dff_B_AgdktrfV4_2;
	wire w_dff_B_SyU2s1Sj8_2;
	wire w_dff_B_TmYQ4m1W4_2;
	wire w_dff_B_uVMWVjQb0_2;
	wire w_dff_B_uagxMc4J3_2;
	wire w_dff_B_nedMcWL41_2;
	wire w_dff_B_EJ602wVC7_2;
	wire w_dff_B_zNRMbOVC5_2;
	wire w_dff_B_O0XDEz0J2_2;
	wire w_dff_B_tMbhbP9K9_2;
	wire w_dff_B_GtMLA1TE7_2;
	wire w_dff_B_CfVVt80c6_2;
	wire w_dff_B_PNLk8pWd3_2;
	wire w_dff_B_amDPAmdF1_2;
	wire w_dff_B_zqrndod36_2;
	wire w_dff_B_fT7OgN7M8_2;
	wire w_dff_B_CG8ZfgVv1_2;
	wire w_dff_B_druNSZnM0_2;
	wire w_dff_B_wDy28X018_2;
	wire w_dff_B_VvoJFzTR3_2;
	wire w_dff_B_EB4uBugq0_2;
	wire w_dff_B_2T1XdtDl1_2;
	wire w_dff_B_BbgYCdJ65_2;
	wire w_dff_B_Kz6osrUH9_2;
	wire w_dff_B_J4nBOsCP7_2;
	wire w_dff_B_IQTdUg0M8_2;
	wire w_dff_B_vqVDl74n0_2;
	wire w_dff_B_s38a6tfY1_2;
	wire w_dff_B_HFPoG2LJ8_2;
	wire w_dff_B_nYTioUsq0_2;
	wire w_dff_B_gwJqSQnA4_2;
	wire w_dff_B_lBSLs1DI8_2;
	wire w_dff_B_NN8zJ1x25_2;
	wire w_dff_B_OZfqgxWB4_2;
	wire w_dff_B_6Y8cJT6S0_2;
	wire w_dff_B_gsjuqBPn0_2;
	wire w_dff_B_l7Sj046f1_2;
	wire w_dff_B_RZB5afjY7_2;
	wire w_dff_B_imRLAERZ0_2;
	wire w_dff_B_t5lxNJun8_2;
	wire w_dff_B_Z0BtaOVv9_2;
	wire w_dff_B_7ftk6shM5_2;
	wire w_dff_B_SJYor4cu9_2;
	wire w_dff_B_PYdspwWx5_2;
	wire w_dff_B_TdwCeMJV4_2;
	wire w_dff_B_r2JSgjXJ2_2;
	wire w_dff_B_vNvxmP1U6_2;
	wire w_dff_B_EJ1Pm7es9_2;
	wire w_dff_B_rQDUj1Vr9_2;
	wire w_dff_B_GNSPR3aJ4_2;
	wire w_dff_B_JI6uYzf38_2;
	wire w_dff_B_9C6Rr72o8_2;
	wire w_dff_B_aLlZACOc9_2;
	wire w_dff_B_RULpIXsq8_2;
	wire w_dff_B_Zsy0vRJv1_2;
	wire w_dff_B_IXMaCWHe2_2;
	wire w_dff_B_GA5bSx567_2;
	wire w_dff_B_8ZFvWMEG0_2;
	wire w_dff_B_2rgNDfTq6_2;
	wire w_dff_B_2Sgye0nx5_2;
	wire w_dff_B_CGz959fP4_2;
	wire w_dff_B_UMDIFo0e1_2;
	wire w_dff_B_YXTPGBjk7_2;
	wire w_dff_B_HdXbFFF26_2;
	wire w_dff_B_JAJzgZW73_2;
	wire w_dff_B_SlyuKEI28_2;
	wire w_dff_B_7gktJ1yw4_2;
	wire w_dff_B_Jns0gf7Z7_2;
	wire w_dff_B_Oky6VBgY6_2;
	wire w_dff_B_AZEJgdk93_2;
	wire w_dff_B_XYX6scPp4_2;
	wire w_dff_B_XK6G5zYL8_2;
	wire w_dff_B_cHEqulFX0_2;
	wire w_dff_B_kJbWkHSd9_2;
	wire w_dff_B_Gi5MsAd61_2;
	wire w_dff_B_df8nTyr38_1;
	wire w_dff_B_Kc3JxjFy3_2;
	wire w_dff_B_ab32jLiY5_2;
	wire w_dff_B_OdUybZNN6_2;
	wire w_dff_B_MahVShMK0_2;
	wire w_dff_B_WpV9de4t7_2;
	wire w_dff_B_neJ2wEdv6_2;
	wire w_dff_B_8bp1GZPb0_2;
	wire w_dff_B_bhOwstdk1_2;
	wire w_dff_B_HROPr6sp4_2;
	wire w_dff_B_udesApIZ9_2;
	wire w_dff_B_LDMCuwR39_2;
	wire w_dff_B_jFyLK0dc0_2;
	wire w_dff_B_uimemobK6_2;
	wire w_dff_B_vPCTWK6K1_2;
	wire w_dff_B_PGVuK9349_2;
	wire w_dff_B_9Ii5kWkm0_2;
	wire w_dff_B_3TsY9hxj0_2;
	wire w_dff_B_YSVlqAD68_2;
	wire w_dff_B_UI7fXv842_2;
	wire w_dff_B_ZvBh2sIL5_2;
	wire w_dff_B_dVzk8pWh9_2;
	wire w_dff_B_hgfIgNlB0_2;
	wire w_dff_B_GBdlN8tU1_2;
	wire w_dff_B_RryZuItE0_2;
	wire w_dff_B_yvTMCjiP7_2;
	wire w_dff_B_RkzM8Yi26_2;
	wire w_dff_B_NTPSMIke1_2;
	wire w_dff_B_eUYmdRU37_2;
	wire w_dff_B_MhSWmCHF2_2;
	wire w_dff_B_wqkcv9TC5_2;
	wire w_dff_B_doWquLHD6_2;
	wire w_dff_B_pA8vGTAg6_2;
	wire w_dff_B_0m6J8dqN9_2;
	wire w_dff_B_4MiELK345_2;
	wire w_dff_B_47ewNo307_2;
	wire w_dff_B_wjKxITkK3_2;
	wire w_dff_B_WJYGTsHj0_1;
	wire w_dff_B_Hip9cB0c0_1;
	wire w_dff_B_fqZYClF17_2;
	wire w_dff_B_XBTvMr9v1_2;
	wire w_dff_B_ghMS6MsN1_2;
	wire w_dff_B_59i6FpCy2_2;
	wire w_dff_B_moRsaybu7_2;
	wire w_dff_B_rcFslrCy7_2;
	wire w_dff_B_hSELKlPW8_2;
	wire w_dff_B_UG3916dJ5_2;
	wire w_dff_B_dZRTrxZB6_2;
	wire w_dff_B_b1N6H1r40_2;
	wire w_dff_B_5IbtYzTC1_2;
	wire w_dff_B_OCzzEgDC8_2;
	wire w_dff_B_ipgcKSCe3_2;
	wire w_dff_B_R4VJ3Sr68_2;
	wire w_dff_B_2wY2V7gg0_2;
	wire w_dff_B_1evDCg2j8_2;
	wire w_dff_B_t4L0GnZx2_2;
	wire w_dff_B_zFJza9Af3_2;
	wire w_dff_B_AZzzrBBw1_2;
	wire w_dff_B_VXIVymVf9_2;
	wire w_dff_B_uVoM8roE6_2;
	wire w_dff_B_ZhdP4AXv9_2;
	wire w_dff_B_3XsMJqFg2_2;
	wire w_dff_B_w0xk2gsv6_2;
	wire w_dff_B_93wGTiVo5_2;
	wire w_dff_B_V89d4gDM0_2;
	wire w_dff_B_ng2Se3Qv8_2;
	wire w_dff_B_7RSODiMM0_2;
	wire w_dff_B_xEekS89M6_2;
	wire w_dff_B_zJbCZklX8_2;
	wire w_dff_B_ipcv16086_2;
	wire w_dff_B_TTARY8Rj9_2;
	wire w_dff_B_a3zElpLN1_2;
	wire w_dff_B_KWKAVASx4_2;
	wire w_dff_B_P1kuuF9V8_2;
	wire w_dff_B_RGR5oJBC5_2;
	wire w_dff_B_Zd3O4XIk4_2;
	wire w_dff_B_xRXXHCDU5_2;
	wire w_dff_B_zNHXZvMf2_2;
	wire w_dff_B_BCyv68xR5_2;
	wire w_dff_B_znL5EFci3_2;
	wire w_dff_B_VZoOeUAS0_2;
	wire w_dff_B_su47rQAO5_2;
	wire w_dff_B_Vh8qAGoS0_2;
	wire w_dff_B_TDBdd1qY1_2;
	wire w_dff_B_3764zBtX5_2;
	wire w_dff_B_NnQj9aBl4_2;
	wire w_dff_B_nBeaxeVp2_2;
	wire w_dff_B_hWjvjyXJ5_2;
	wire w_dff_B_w6Yd3EN50_2;
	wire w_dff_B_uwE98vtO7_2;
	wire w_dff_B_dIrjrwRw6_2;
	wire w_dff_B_vlMeF1YR0_2;
	wire w_dff_B_GkYapuNh0_2;
	wire w_dff_B_Djwi7hZv2_2;
	wire w_dff_B_dlcXEriD3_2;
	wire w_dff_B_p1SbDHGp7_2;
	wire w_dff_B_YEAecKDB7_2;
	wire w_dff_B_agpdSzXV4_2;
	wire w_dff_B_7c1YjoS18_2;
	wire w_dff_B_Uyo0hUlD6_2;
	wire w_dff_B_lhHaqCbk2_2;
	wire w_dff_B_Jg0HP3nZ6_2;
	wire w_dff_B_r2J4KLyT0_2;
	wire w_dff_B_Q5bAYjee7_2;
	wire w_dff_B_APvONUqZ7_2;
	wire w_dff_B_5BiHwCAM0_2;
	wire w_dff_B_6V8zst9C7_2;
	wire w_dff_B_jQ8wPSVW4_2;
	wire w_dff_B_LwpMB43I2_1;
	wire w_dff_B_GugcLrnm6_2;
	wire w_dff_B_AbZlQYC56_2;
	wire w_dff_B_TZ8AIovi4_2;
	wire w_dff_B_RHITzt4v1_2;
	wire w_dff_B_NoDuwryF8_2;
	wire w_dff_B_wyoowKMJ2_2;
	wire w_dff_B_DjjCQl1h6_2;
	wire w_dff_B_OnTXUDJC7_2;
	wire w_dff_B_mWvhFxjm4_2;
	wire w_dff_B_j91NeEOV8_2;
	wire w_dff_B_ba1GqPRL1_2;
	wire w_dff_B_COn85NbT6_2;
	wire w_dff_B_F1bmglqz6_2;
	wire w_dff_B_rusZJjk15_2;
	wire w_dff_B_rjQ0MfK38_2;
	wire w_dff_B_uPzjkIAx0_2;
	wire w_dff_B_GVjPtiHJ5_2;
	wire w_dff_B_EWDpgouP8_2;
	wire w_dff_B_EYyV6B744_2;
	wire w_dff_B_SIrYyk2z7_2;
	wire w_dff_B_fXrWZS0D5_2;
	wire w_dff_B_SCO1RFWY4_2;
	wire w_dff_B_whHMKccd6_2;
	wire w_dff_B_qWG4D4Zx9_2;
	wire w_dff_B_uD3e3aUz3_2;
	wire w_dff_B_n9LNErZ02_2;
	wire w_dff_B_oQp4IJEg0_2;
	wire w_dff_B_2kZfCFYy1_2;
	wire w_dff_B_PUckGBek7_2;
	wire w_dff_B_63oH4BDt9_2;
	wire w_dff_B_7oxKpmbY9_2;
	wire w_dff_B_baoqdbM52_2;
	wire w_dff_B_c2yjbTwH0_1;
	wire w_dff_B_SlEBjpw15_1;
	wire w_dff_B_x7ZnNhe53_2;
	wire w_dff_B_8DnKZYTP2_2;
	wire w_dff_B_YkQjSEPa4_2;
	wire w_dff_B_SzWCiNbT8_2;
	wire w_dff_B_fN38XyAa7_2;
	wire w_dff_B_q4503rNP6_2;
	wire w_dff_B_gDkx0rSA9_2;
	wire w_dff_B_lsTORZFR4_2;
	wire w_dff_B_eMvivkk69_2;
	wire w_dff_B_2dOYPNCN6_2;
	wire w_dff_B_4lEFZheb6_2;
	wire w_dff_B_z5VFRaH92_2;
	wire w_dff_B_Bhhd5Y0G9_2;
	wire w_dff_B_pG3vB1Ii5_2;
	wire w_dff_B_FqJ8Xvwo0_2;
	wire w_dff_B_h1yJEpBM9_2;
	wire w_dff_B_A8eIH1ei6_2;
	wire w_dff_B_68fSbukW8_2;
	wire w_dff_B_gNwX56j45_2;
	wire w_dff_B_UNdv8N1s5_2;
	wire w_dff_B_ZI6kZ0CH1_2;
	wire w_dff_B_Xj80AD3f2_2;
	wire w_dff_B_ItotBtzo2_2;
	wire w_dff_B_zeBcSGFn5_2;
	wire w_dff_B_M96nUBHJ0_2;
	wire w_dff_B_aggZNkns5_2;
	wire w_dff_B_CwnYIZsQ2_2;
	wire w_dff_B_cKmGXSGE9_2;
	wire w_dff_B_BxO64W1V2_2;
	wire w_dff_B_vtUutOwt3_2;
	wire w_dff_B_7sTMXM465_2;
	wire w_dff_B_KKyuNzo66_2;
	wire w_dff_B_DDkdSG1i2_2;
	wire w_dff_B_mBhy0BFq7_2;
	wire w_dff_B_l7L0FhuG2_2;
	wire w_dff_B_u28Jy0qd1_2;
	wire w_dff_B_DRJyE8b40_2;
	wire w_dff_B_JiYLPRuo6_2;
	wire w_dff_B_5vuPtkq32_2;
	wire w_dff_B_UdjggULq0_2;
	wire w_dff_B_DNFsz12B0_2;
	wire w_dff_B_ny3lv2Jd9_2;
	wire w_dff_B_hhnvwzLR4_2;
	wire w_dff_B_gnsUch1D4_2;
	wire w_dff_B_0f9njkGx2_2;
	wire w_dff_B_fDmKdxwM5_2;
	wire w_dff_B_ELoFqzoL2_2;
	wire w_dff_B_hYN2DRpR5_2;
	wire w_dff_B_fEbKfBrj6_2;
	wire w_dff_B_98wTQw1G1_2;
	wire w_dff_B_GBiiiZej1_2;
	wire w_dff_B_lnUtt5NM5_2;
	wire w_dff_B_YNTsZpgP4_2;
	wire w_dff_B_UwOKQZCP9_2;
	wire w_dff_B_z27gR8kK1_2;
	wire w_dff_B_LMPaQdI47_2;
	wire w_dff_B_tXTTbGDF2_2;
	wire w_dff_B_YSqoSBQi6_2;
	wire w_dff_B_5TA3ku9h4_2;
	wire w_dff_B_oAJS2gxH9_2;
	wire w_dff_B_p4XeoJmg1_2;
	wire w_dff_B_eAljtyPM9_1;
	wire w_dff_B_dcRyaz0x3_2;
	wire w_dff_B_VfX6BxUF7_2;
	wire w_dff_B_innOVUcS8_2;
	wire w_dff_B_FaLf88IZ5_2;
	wire w_dff_B_edtbpbmp0_2;
	wire w_dff_B_H6OjrtMF1_2;
	wire w_dff_B_iTrgwVPV5_2;
	wire w_dff_B_S1rTYZ5R5_2;
	wire w_dff_B_GqmIozHi6_2;
	wire w_dff_B_PICjZBWz6_2;
	wire w_dff_B_FlKleEVC8_2;
	wire w_dff_B_hDozs50r1_2;
	wire w_dff_B_CNEgWOUT6_2;
	wire w_dff_B_Bn6sZ6mb0_2;
	wire w_dff_B_LYJCQMxE4_2;
	wire w_dff_B_wXJDgVuo0_2;
	wire w_dff_B_DZ0VPlyn8_2;
	wire w_dff_B_FegmY1Od9_2;
	wire w_dff_B_qTyaly0q4_2;
	wire w_dff_B_cQKEC7547_2;
	wire w_dff_B_uz5NnPzy5_2;
	wire w_dff_B_duFxJ8s00_2;
	wire w_dff_B_SC7R0snO2_2;
	wire w_dff_B_91KWYDUn6_2;
	wire w_dff_B_lCxN2mNQ5_2;
	wire w_dff_B_AuWPTUae7_2;
	wire w_dff_B_77y9GENH0_2;
	wire w_dff_B_3aHAWKT57_2;
	wire w_dff_B_c3bULSld1_1;
	wire w_dff_B_jkG7Gnh21_1;
	wire w_dff_B_3lm5RqDx4_2;
	wire w_dff_B_ZmTez0jb0_2;
	wire w_dff_B_QHzUqkc97_2;
	wire w_dff_B_6IBFZh2k8_2;
	wire w_dff_B_AuJfrlsY4_2;
	wire w_dff_B_8mW2OEhD4_2;
	wire w_dff_B_DfMVywnC4_2;
	wire w_dff_B_aOvUAm1s6_2;
	wire w_dff_B_ekBohHdc3_2;
	wire w_dff_B_M87LqWdH1_2;
	wire w_dff_B_JT8HwOxL6_2;
	wire w_dff_B_A3UkykDj6_2;
	wire w_dff_B_uNVEeAel7_2;
	wire w_dff_B_Phg1ej875_2;
	wire w_dff_B_bkF9Tx1m0_2;
	wire w_dff_B_FRuFpevk2_2;
	wire w_dff_B_9drKR0pB5_2;
	wire w_dff_B_OyvTpN4s8_2;
	wire w_dff_B_AycQ6MKX1_2;
	wire w_dff_B_cR2o2IGY3_2;
	wire w_dff_B_pfK1Zg7E2_2;
	wire w_dff_B_yFKj9PKM2_2;
	wire w_dff_B_SHUOJgeh1_2;
	wire w_dff_B_CC0YeSiT7_2;
	wire w_dff_B_0ytc6keY6_2;
	wire w_dff_B_kGcpJOVY7_2;
	wire w_dff_B_J4JWlldT8_2;
	wire w_dff_B_kObFjjDR0_2;
	wire w_dff_B_iED7qo193_2;
	wire w_dff_B_E8JasFAi5_2;
	wire w_dff_B_AvWwjkFq5_2;
	wire w_dff_B_M2709WEX8_2;
	wire w_dff_B_BgXFYNdH3_2;
	wire w_dff_B_Op3T7d9G6_2;
	wire w_dff_B_GGjH24kH3_2;
	wire w_dff_B_AJOeFvkt2_2;
	wire w_dff_B_JDPIXf858_2;
	wire w_dff_B_RcXo07651_2;
	wire w_dff_B_gasTXOml2_2;
	wire w_dff_B_FMzdovn09_2;
	wire w_dff_B_7kEQqkeJ4_2;
	wire w_dff_B_7Y8VCaGV4_2;
	wire w_dff_B_uZOvTSdZ3_2;
	wire w_dff_B_Q0GSHaYs1_2;
	wire w_dff_B_XAHFpnQC3_2;
	wire w_dff_B_ROfSh6Eo9_2;
	wire w_dff_B_HgsUEgEm5_2;
	wire w_dff_B_DQXPQeFA6_2;
	wire w_dff_B_GZgteWl33_2;
	wire w_dff_B_MkF20I2O9_2;
	wire w_dff_B_oDtEooSa4_2;
	wire w_dff_B_w3yWoLIG5_2;
	wire w_dff_B_1ZVbO9WY8_2;
	wire w_dff_B_Qgbz1cZp2_1;
	wire w_dff_B_piQY7FD69_2;
	wire w_dff_B_MjDz38Rb0_2;
	wire w_dff_B_NkNoymbq0_2;
	wire w_dff_B_kbq4Q1ix0_2;
	wire w_dff_B_GsCu1Mc82_2;
	wire w_dff_B_gsBRj3eu6_2;
	wire w_dff_B_GiL44ctW6_2;
	wire w_dff_B_t4jjJZ4n9_2;
	wire w_dff_B_8AMbdcLi9_2;
	wire w_dff_B_zuHQfkPo9_2;
	wire w_dff_B_2qWfIzGz7_2;
	wire w_dff_B_CdpdPQOS9_2;
	wire w_dff_B_2LbnHy5O1_2;
	wire w_dff_B_KejJAvHh6_2;
	wire w_dff_B_SV2YQmhc9_2;
	wire w_dff_B_N24Ub3J52_2;
	wire w_dff_B_zVqUjW0n6_2;
	wire w_dff_B_J71eQzl57_2;
	wire w_dff_B_HZDIJFTy6_2;
	wire w_dff_B_po3Xfo5O2_2;
	wire w_dff_B_um4wzFQ99_2;
	wire w_dff_B_CWHlLOav1_2;
	wire w_dff_B_95dXR3pb1_2;
	wire w_dff_B_EzliOta12_2;
	wire w_dff_B_OiPdZfzd9_1;
	wire w_dff_B_WWR6ioqC4_1;
	wire w_dff_B_doWhhhXj9_2;
	wire w_dff_B_NymjAeOs9_2;
	wire w_dff_B_lXDpwh3A1_2;
	wire w_dff_B_ER9wpk1s2_2;
	wire w_dff_B_580gmNBR1_2;
	wire w_dff_B_5XsftpV22_2;
	wire w_dff_B_DqEmxztK3_2;
	wire w_dff_B_fiR0a2pm3_2;
	wire w_dff_B_EGmb7ZUH8_2;
	wire w_dff_B_qKlxcxXJ3_2;
	wire w_dff_B_ArxJjXMQ5_2;
	wire w_dff_B_ZjEzips51_2;
	wire w_dff_B_pwy0Ktlq6_2;
	wire w_dff_B_gzqJSMd32_2;
	wire w_dff_B_gipH3PPL1_2;
	wire w_dff_B_hogzUncN2_2;
	wire w_dff_B_42pL21Zb0_2;
	wire w_dff_B_utlxdGBp8_2;
	wire w_dff_B_ONUyUNkJ2_2;
	wire w_dff_B_hE1OpSM45_2;
	wire w_dff_B_S3RGNprc3_2;
	wire w_dff_B_8v4kmHIr0_2;
	wire w_dff_B_oNAkpXc45_2;
	wire w_dff_B_J3Fv31er0_2;
	wire w_dff_B_sy6vPOu41_2;
	wire w_dff_B_pexyw1il9_2;
	wire w_dff_B_cQqQwQ7A9_2;
	wire w_dff_B_fKPmDFBN9_2;
	wire w_dff_B_UuNmlEi89_2;
	wire w_dff_B_GWOzs5ni6_2;
	wire w_dff_B_piPFD9aN1_2;
	wire w_dff_B_1Ph9KQoK7_2;
	wire w_dff_B_3nFcw1C58_2;
	wire w_dff_B_1t08g69X5_2;
	wire w_dff_B_ncdylhJS9_2;
	wire w_dff_B_VgY1Hdjs5_2;
	wire w_dff_B_rPA5s7yn8_2;
	wire w_dff_B_VjpRjuk45_2;
	wire w_dff_B_xasKGlYQ8_2;
	wire w_dff_B_felqBjNZ5_2;
	wire w_dff_B_ZPYw7DlJ2_2;
	wire w_dff_B_UV0Eixpq8_2;
	wire w_dff_B_HPnERQSg0_2;
	wire w_dff_B_P5aKcMzV6_2;
	wire w_dff_B_obud84Fq6_2;
	wire w_dff_B_xvrIb0mS9_1;
	wire w_dff_B_UZP12VuM1_2;
	wire w_dff_B_X46FJYec7_2;
	wire w_dff_B_hpqdlP1B8_2;
	wire w_dff_B_8oI7eOp77_2;
	wire w_dff_B_o6bquFzt8_2;
	wire w_dff_B_ckWZdXUX0_2;
	wire w_dff_B_5azc3tdZ1_2;
	wire w_dff_B_Dq587cjY0_2;
	wire w_dff_B_WYhCNK918_2;
	wire w_dff_B_OCoodkJc4_2;
	wire w_dff_B_UI7bWbGz9_2;
	wire w_dff_B_bGvhDLWC7_2;
	wire w_dff_B_RhCtjxKE0_2;
	wire w_dff_B_KvpPmaY98_2;
	wire w_dff_B_wof6xHnK4_2;
	wire w_dff_B_LKRcOnkX0_2;
	wire w_dff_B_op1iX8rY0_2;
	wire w_dff_B_OW6n44te8_2;
	wire w_dff_B_rpq5eHw38_2;
	wire w_dff_B_sIGu0EXt3_2;
	wire w_dff_B_Rauj33Hx7_1;
	wire w_dff_B_qLfpP2yC6_1;
	wire w_dff_B_ieZrxodV4_2;
	wire w_dff_B_h12KJgud2_2;
	wire w_dff_B_c8XFa7nk8_2;
	wire w_dff_B_DCEYz4Lr7_2;
	wire w_dff_B_BtuclDl46_2;
	wire w_dff_B_NOJpTwrO2_2;
	wire w_dff_B_Fe9Tkhlu7_2;
	wire w_dff_B_o8BBL3m74_2;
	wire w_dff_B_FFEWbkTz0_2;
	wire w_dff_B_FNwXay5i3_2;
	wire w_dff_B_Tt7NSMvs7_2;
	wire w_dff_B_snCwN42f3_2;
	wire w_dff_B_FZ8SdgGh0_2;
	wire w_dff_B_APAPQfSQ3_2;
	wire w_dff_B_3QZVNOAL8_2;
	wire w_dff_B_2JQWDic04_2;
	wire w_dff_B_FySL7aDB0_2;
	wire w_dff_B_Z8bmcoua3_2;
	wire w_dff_B_81FDSwIW1_2;
	wire w_dff_B_lWxB88oV9_2;
	wire w_dff_B_WGblt9En9_2;
	wire w_dff_B_xPNbKXED9_2;
	wire w_dff_B_lLgwbKra1_2;
	wire w_dff_B_CkXWAS8q2_2;
	wire w_dff_B_PywBbwpA8_2;
	wire w_dff_B_b4YVCQlx5_2;
	wire w_dff_B_QhXkmSDI0_2;
	wire w_dff_B_siap2Erl7_2;
	wire w_dff_B_ZDgohWOT2_2;
	wire w_dff_B_7DeUiXoB2_2;
	wire w_dff_B_kIZfLlmz3_2;
	wire w_dff_B_imIW2sWm4_2;
	wire w_dff_B_MFs6FmlM3_2;
	wire w_dff_B_X1CLj5ET8_2;
	wire w_dff_B_sOSGaqFI5_2;
	wire w_dff_B_4OFR99W31_2;
	wire w_dff_B_fF22xHZ72_1;
	wire w_dff_B_LpHrC3td5_2;
	wire w_dff_B_3bRU1I8S0_2;
	wire w_dff_B_mHldo0tM9_2;
	wire w_dff_B_OT2uoaZ40_2;
	wire w_dff_B_doxB9s1K8_2;
	wire w_dff_B_Oalguq2R5_2;
	wire w_dff_B_rsqeRcUk3_2;
	wire w_dff_B_WcySLL2d2_2;
	wire w_dff_B_rRChLAt44_2;
	wire w_dff_B_5oOxccy72_2;
	wire w_dff_B_A6Q4mzqB0_2;
	wire w_dff_B_qLh1rJOC9_2;
	wire w_dff_B_5TeLkKGR2_2;
	wire w_dff_B_EMvmhfn53_2;
	wire w_dff_B_h8AWiYyk6_2;
	wire w_dff_B_5D5Qzu784_2;
	wire w_dff_B_mp4WhI0R0_2;
	wire w_dff_B_4RzogzYx1_2;
	wire w_dff_B_YfxulAEM9_1;
	wire w_dff_B_DY66GdNE4_1;
	wire w_dff_B_6YIX5qiW0_2;
	wire w_dff_B_cFZ7vhnJ3_2;
	wire w_dff_B_LvMbsXMz4_2;
	wire w_dff_B_0afRMXRA5_2;
	wire w_dff_B_YbhA4pNj6_2;
	wire w_dff_B_PkWTiQfA4_2;
	wire w_dff_B_xOupLYoq8_2;
	wire w_dff_B_uKeiKftv8_2;
	wire w_dff_B_9vJRf5FY2_2;
	wire w_dff_B_HXqP3gBQ3_2;
	wire w_dff_B_EorAVzXZ9_2;
	wire w_dff_B_oivbJ5lx0_2;
	wire w_dff_B_1tzjXXiY8_2;
	wire w_dff_B_IIVSuTXM6_2;
	wire w_dff_B_qzKKlDqP2_2;
	wire w_dff_B_Qh1da2da3_2;
	wire w_dff_B_6e6bukUb7_2;
	wire w_dff_B_JzfdNGzG1_2;
	wire w_dff_B_XUaFS7bj0_2;
	wire w_dff_B_v4Nt48gh8_2;
	wire w_dff_B_jd1pvwFq1_2;
	wire w_dff_B_jHy9EOol7_2;
	wire w_dff_B_gH8pRmX97_2;
	wire w_dff_B_LfQ2JeJl7_2;
	wire w_dff_B_x8VQxSHb2_2;
	wire w_dff_B_8uHJxpYY7_2;
	wire w_dff_B_5YJDHX9f4_2;
	wire w_dff_B_wCNWPAxc6_2;
	wire w_dff_B_rMz0XjOQ0_1;
	wire w_dff_B_yh3oE8w74_2;
	wire w_dff_B_Kt4m0qyQ8_2;
	wire w_dff_B_0tysaLwm9_2;
	wire w_dff_B_soh2w2Vt2_2;
	wire w_dff_B_vHZeM2a86_2;
	wire w_dff_B_ZIxMueCJ2_2;
	wire w_dff_B_QHf1iKAe8_2;
	wire w_dff_B_L6B3r8fA2_2;
	wire w_dff_B_7UNYeD0A0_2;
	wire w_dff_B_JiOSGKO16_2;
	wire w_dff_B_n2uwMoUY0_2;
	wire w_dff_B_tlkm3Xnl4_2;
	wire w_dff_B_nXIyRATt2_2;
	wire w_dff_B_gsC6wqNH0_2;
	wire w_dff_B_LUhwgJYf1_2;
	wire w_dff_B_l1BIsj2K7_2;
	wire w_dff_B_FMMA80sR8_1;
	wire w_dff_B_T8VZlarh2_1;
	wire w_dff_B_sqZW4AaN1_2;
	wire w_dff_B_mB61WCyw8_2;
	wire w_dff_B_yG5hC4mr5_2;
	wire w_dff_B_rAP4h9PY5_2;
	wire w_dff_B_iYdgua2v5_2;
	wire w_dff_B_CHRacBht2_2;
	wire w_dff_B_tcyb7Ah26_2;
	wire w_dff_B_NqSMCDDU1_2;
	wire w_dff_B_bHlhii1X8_2;
	wire w_dff_B_tNYKdjia8_2;
	wire w_dff_B_lE9E1rrc1_2;
	wire w_dff_B_40Gezdqh1_2;
	wire w_dff_B_9Xzy9A743_2;
	wire w_dff_B_4Pdrrfuv6_2;
	wire w_dff_B_nKYygaBl3_2;
	wire w_dff_B_VgjF3Ddo0_2;
	wire w_dff_B_eNnSARLR1_2;
	wire w_dff_B_6JUHd4Uy0_2;
	wire w_dff_B_6EwDfvpH1_2;
	wire w_dff_B_3iHvH29H0_2;
	wire w_dff_B_EaFpkXqV1_1;
	wire w_dff_B_Y00VNV5P6_2;
	wire w_dff_B_tz2glaSP3_2;
	wire w_dff_B_OljZJaSS9_2;
	wire w_dff_B_IbXrYaYB1_2;
	wire w_dff_B_GWQHjMTX7_2;
	wire w_dff_B_hyat70PT0_2;
	wire w_dff_B_CSDHSm5r4_2;
	wire w_dff_B_ydb2yCIh5_2;
	wire w_dff_B_q3BEP2P83_2;
	wire w_dff_B_ScIGnvEV2_2;
	wire w_dff_B_vR19TmIW5_2;
	wire w_dff_B_iLqcGY7d8_2;
	wire w_dff_B_vTgByL8q6_2;
	wire w_dff_B_QBuWzmQu0_2;
	wire w_dff_B_NavRGwX05_2;
	wire w_dff_B_4rgkupxz3_2;
	wire w_dff_B_AgB7gdh96_2;
	wire w_dff_B_D0Rwz3jX7_2;
	wire w_dff_B_s8ukJ44q7_2;
	wire w_dff_B_t1JgZ43E2_2;
	wire w_dff_B_CGtPIEal5_2;
	wire w_dff_B_zMlyabps6_2;
	wire w_dff_B_YgOjHMXK5_2;
	wire w_dff_B_uAvbnW1L3_2;
	wire w_dff_B_9asOxlze8_2;
	wire w_dff_B_x50Fva0C5_2;
	wire w_dff_B_U2eEKYyt1_1;
	wire w_dff_B_B786o5QK3_2;
	wire w_dff_B_PnWj6IOu5_2;
	wire w_dff_B_y1XSpmK04_2;
	wire w_dff_B_enB6kYnQ0_2;
	wire w_dff_B_XIqwfjWb0_2;
	wire w_dff_B_RgoM6Jzc8_2;
	wire w_dff_B_6UsLvbar2_2;
	wire w_dff_B_c4z6oQvR5_2;
	wire w_dff_B_1XvQhRLC2_2;
	wire w_dff_B_HnC3DcPT0_2;
	wire w_dff_B_P6yanSA50_2;
	wire w_dff_B_1PruDQuf8_2;
	wire w_dff_B_lgtWnk074_2;
	wire w_dff_B_1aKC89GH2_2;
	wire w_dff_B_gu26uhNi2_2;
	wire w_dff_A_hWGiBTey5_0;
	wire w_dff_A_j2iJF3dD4_0;
	wire w_dff_A_cTYpb9Uc5_0;
	wire w_dff_B_0eI2STGI0_2;
	wire w_dff_A_Tj1mn60e8_0;
	wire w_dff_A_CHYnw0Mb4_0;
	wire w_dff_A_nVhSQM5i0_0;
	wire w_dff_B_91FhsFt05_2;
	wire w_dff_A_GSJ5BpHw4_0;
	wire w_dff_A_U3lV2lY70_0;
	wire w_dff_B_yVRLDYHI0_2;
	wire w_dff_B_wglqkA0O8_2;
	wire w_dff_B_sHzh34fk5_2;
	wire w_dff_A_Fe3KFXMD4_1;
	wire w_dff_A_spfPBIUn3_0;
	wire w_dff_A_95A7I1Kf9_0;
	wire w_dff_A_EqG0Wzs46_0;
	wire w_dff_A_uPVtwYRJ4_0;
	wire w_dff_A_C4CjRsh24_0;
	wire w_dff_A_V0en8nbW3_0;
	wire w_dff_A_ZjhSb9Oq4_0;
	wire w_dff_A_EvJcgQzi7_0;
	wire w_dff_A_6HaGyRM36_0;
	wire w_dff_A_gNoPZlNg0_0;
	wire w_dff_A_cfH63hYN2_0;
	wire w_dff_A_6D3v2Ycd2_0;
	wire w_dff_A_kgko3x4Q8_0;
	wire w_dff_A_jDHW5v3Q0_0;
	wire w_dff_A_L86RYP2Y6_0;
	wire w_dff_A_Bhzq0YMv5_0;
	wire w_dff_A_TbH3fasC7_0;
	wire w_dff_A_3gq02Vfb6_0;
	wire w_dff_A_hZKeKtNB7_0;
	wire w_dff_A_80GCqJf52_0;
	wire w_dff_A_AP83QNGI4_0;
	wire w_dff_A_46Jazfvb7_0;
	wire w_dff_A_8JMTCC4G7_0;
	wire w_dff_A_igBzCly85_0;
	wire w_dff_A_67uThCbv0_0;
	wire w_dff_A_BMfnBHBV9_0;
	wire w_dff_A_KH7iVs1y8_0;
	wire w_dff_A_5sBtDR4h7_0;
	wire w_dff_A_3TARjgSY8_0;
	wire w_dff_A_PXQYzuSd2_0;
	wire w_dff_A_A5UXe75s6_0;
	wire w_dff_A_VPlY73v35_0;
	wire w_dff_A_9wkwbeZy1_0;
	wire w_dff_A_4k9ggX7N0_0;
	wire w_dff_A_IJrmdSH98_0;
	wire w_dff_A_s9CQY1F47_0;
	wire w_dff_A_L4l8MKV24_0;
	wire w_dff_A_ep9F4Npv2_0;
	wire w_dff_A_s7o1HIsz7_0;
	wire w_dff_A_Ot1OUzNt5_0;
	wire w_dff_A_5OqTouOM2_0;
	wire w_dff_A_yjgt2cjq9_0;
	wire w_dff_A_FCyEI8Ij2_0;
	wire w_dff_A_XwTCm0QV6_0;
	wire w_dff_A_ib8Pv4T83_0;
	wire w_dff_A_IoObJSrG4_0;
	wire w_dff_A_i9lHLVO34_0;
	wire w_dff_A_8NAOYYnA8_0;
	wire w_dff_A_0yLf0eDj1_0;
	wire w_dff_A_eAGRm9zi7_0;
	wire w_dff_A_Yabd95VT8_0;
	wire w_dff_A_e21pVVJK5_0;
	wire w_dff_A_bCnAN8eK6_0;
	wire w_dff_A_jEjHb6RW0_0;
	wire w_dff_A_OTF0tl1Z2_0;
	wire w_dff_A_aA7Uiq1F0_0;
	wire w_dff_A_vqsK2C1f4_0;
	wire w_dff_A_14hF01UT8_0;
	wire w_dff_A_mFl9UivU7_0;
	wire w_dff_A_kOkCmNTa2_0;
	wire w_dff_A_BlFefluR4_0;
	wire w_dff_A_4TduGLqi5_0;
	wire w_dff_A_798Pic9G4_0;
	wire w_dff_A_90x6earD2_0;
	wire w_dff_A_EDcuu3vf3_0;
	wire w_dff_A_gTxKXYil8_0;
	wire w_dff_A_XQeKpwe45_0;
	wire w_dff_A_AlFKrb5A8_0;
	wire w_dff_A_l3ffOSui7_0;
	wire w_dff_A_K8tqUTVv5_0;
	wire w_dff_A_HNGQKIgh5_0;
	wire w_dff_A_sBFbWx9O6_0;
	wire w_dff_A_WB9YxVfw4_0;
	wire w_dff_A_NslXWg0x3_2;
	wire w_dff_A_I5WThFvY9_0;
	wire w_dff_A_5rbu215e2_0;
	wire w_dff_A_LPvp6EMm3_0;
	wire w_dff_A_pGhZ6fo68_0;
	wire w_dff_A_vFbWPHOG9_0;
	wire w_dff_A_Mr0aDnxi3_0;
	wire w_dff_A_jhmVoLMs2_0;
	wire w_dff_A_euC441m84_0;
	wire w_dff_A_F4hX5uHX8_0;
	wire w_dff_A_AI2F0nfn2_0;
	wire w_dff_A_f3mjBQUq4_0;
	wire w_dff_A_0WOiSrou4_0;
	wire w_dff_A_cYLQHQBX9_0;
	wire w_dff_A_eonTJ2wl7_0;
	wire w_dff_A_XeqP43tG6_0;
	wire w_dff_A_UOwWTtj39_0;
	wire w_dff_A_fIalWi3U6_0;
	wire w_dff_A_8wTPooyb8_0;
	wire w_dff_A_aZ5rjZAr3_0;
	wire w_dff_A_UPEs4K000_0;
	wire w_dff_A_axL163r37_0;
	wire w_dff_A_Jj1EUh8x7_0;
	wire w_dff_A_rh3nVGxM1_0;
	wire w_dff_A_eVuzDtIV0_0;
	wire w_dff_A_MzRNPNfU3_0;
	wire w_dff_A_YXKRck8f6_0;
	wire w_dff_A_88pVLx314_0;
	wire w_dff_A_3EdiyTJZ3_0;
	wire w_dff_A_qwSl4dj92_0;
	wire w_dff_A_lBMi7rQc6_0;
	wire w_dff_A_tPeRy6r72_0;
	wire w_dff_A_HR5LP9AX2_0;
	wire w_dff_A_7eglWOl51_0;
	wire w_dff_A_56AO8c590_0;
	wire w_dff_A_eVUbKRmL7_0;
	wire w_dff_A_QDLcDh6t8_0;
	wire w_dff_A_yPHr171L6_0;
	wire w_dff_A_ZZ4hvhWL9_0;
	wire w_dff_A_XvX4plDk1_0;
	wire w_dff_A_1a3VfOzx3_0;
	wire w_dff_A_75n9HyO70_0;
	wire w_dff_A_wQMs33ol9_0;
	wire w_dff_A_d51U9rm39_0;
	wire w_dff_A_xomWgcyQ5_0;
	wire w_dff_A_eutneaXU6_0;
	wire w_dff_A_9fKHYyrl0_0;
	wire w_dff_A_fyhr0Jde6_0;
	wire w_dff_A_tEs4guOG1_0;
	wire w_dff_A_dp3mvErr8_0;
	wire w_dff_A_wynkwt1E3_0;
	wire w_dff_A_y2v0RrB84_0;
	wire w_dff_A_eYPdsBSX3_0;
	wire w_dff_A_yV8RrRx57_0;
	wire w_dff_A_Q9puzdqY5_0;
	wire w_dff_A_05HWikCa1_0;
	wire w_dff_A_SuWjL1B27_0;
	wire w_dff_A_9KudURsQ1_0;
	wire w_dff_A_v5nks1rE4_0;
	wire w_dff_A_umQly1M49_0;
	wire w_dff_A_sk2oOwGJ4_0;
	wire w_dff_A_T6E2pNcF1_0;
	wire w_dff_A_uwSLX6KQ6_0;
	wire w_dff_A_6CYW7BgD0_0;
	wire w_dff_A_VrJxdA0N5_0;
	wire w_dff_A_mQuFLoBo3_0;
	wire w_dff_A_ypOMHuoY4_0;
	wire w_dff_A_ef3ofoF17_0;
	wire w_dff_A_CGlm3Azc7_0;
	wire w_dff_A_0EJiQWms3_0;
	wire w_dff_A_aqNNkNcQ8_2;
	wire w_dff_A_Bcadps6G9_0;
	wire w_dff_A_JngHxxGD0_0;
	wire w_dff_A_qnXymM9S5_0;
	wire w_dff_A_XFGSbv049_0;
	wire w_dff_A_iAPNqVDe6_0;
	wire w_dff_A_7JWiMhIr6_0;
	wire w_dff_A_DIApHEs70_0;
	wire w_dff_A_uqToj7HG0_0;
	wire w_dff_A_iRIcnbg91_0;
	wire w_dff_A_lXmb7PkR3_0;
	wire w_dff_A_ykG41ovV2_0;
	wire w_dff_A_0OoSYOW68_0;
	wire w_dff_A_p11g2EET9_0;
	wire w_dff_A_wR0RbipV7_0;
	wire w_dff_A_CuuGmkAA3_0;
	wire w_dff_A_x21qsiKw8_0;
	wire w_dff_A_U19Zw9DS5_0;
	wire w_dff_A_wTBy4Y314_0;
	wire w_dff_A_3ZPyqDpN0_0;
	wire w_dff_A_emNpalZw6_0;
	wire w_dff_A_JgSWAHOr3_0;
	wire w_dff_A_iENyi0Ou2_0;
	wire w_dff_A_l8YRJB5X1_0;
	wire w_dff_A_ngCzv0wq8_0;
	wire w_dff_A_7jrJ0Wn38_0;
	wire w_dff_A_vhVA9I2D5_0;
	wire w_dff_A_nGdAGcDr6_0;
	wire w_dff_A_MvXObyMj3_0;
	wire w_dff_A_Ge9b69P73_0;
	wire w_dff_A_ioWSYgyo1_0;
	wire w_dff_A_rDyev51K2_0;
	wire w_dff_A_KuPz8kQQ4_0;
	wire w_dff_A_086ab7BX0_0;
	wire w_dff_A_8d3JbXYl3_0;
	wire w_dff_A_XIdSLnhK1_0;
	wire w_dff_A_4C0Rxurq5_0;
	wire w_dff_A_YiMzQWIM0_0;
	wire w_dff_A_sBLe3Nxr3_0;
	wire w_dff_A_sK0OXaTN4_0;
	wire w_dff_A_kHePytj39_0;
	wire w_dff_A_XkN0OuQz6_0;
	wire w_dff_A_9CQ9uvkB1_0;
	wire w_dff_A_xFxhVMVn4_0;
	wire w_dff_A_p9jxaPIf0_0;
	wire w_dff_A_HMnq1jw19_0;
	wire w_dff_A_UdjTtzgm6_0;
	wire w_dff_A_mmcb6lT62_0;
	wire w_dff_A_sZBaC4AJ7_0;
	wire w_dff_A_6OPiAxXu3_0;
	wire w_dff_A_IgyQ1NGe8_0;
	wire w_dff_A_lHISZ7A64_0;
	wire w_dff_A_zV21c5Ja7_0;
	wire w_dff_A_QhYHca3w4_0;
	wire w_dff_A_dvsVWLrZ3_0;
	wire w_dff_A_MQ6t6Fq74_0;
	wire w_dff_A_rTDSSZh00_0;
	wire w_dff_A_ku56SRiv8_0;
	wire w_dff_A_Ui8RXGmf2_0;
	wire w_dff_A_jo8J4tIO0_0;
	wire w_dff_A_lhCUuOAq9_0;
	wire w_dff_A_9dS3Pf2z3_0;
	wire w_dff_A_D4LRZqVc4_0;
	wire w_dff_A_cG1P65du0_0;
	wire w_dff_A_jo7a9cxF6_0;
	wire w_dff_A_8AhaQ92M4_0;
	wire w_dff_A_2aFfJTxd9_0;
	wire w_dff_A_uyEcTvc40_0;
	wire w_dff_A_OdNAlUUY1_0;
	wire w_dff_A_ia5znL6j8_2;
	wire w_dff_A_Sil0NLgq3_0;
	wire w_dff_A_VT5zNKAv4_0;
	wire w_dff_A_ir5PzM1t9_0;
	wire w_dff_A_1WKU4g5p9_0;
	wire w_dff_A_1onpxYXY2_0;
	wire w_dff_A_1zanhRZy4_0;
	wire w_dff_A_3e91Gvn39_0;
	wire w_dff_A_006MIS991_0;
	wire w_dff_A_12b4hOkc4_0;
	wire w_dff_A_RaRIIDE68_0;
	wire w_dff_A_yaWVbUjb0_0;
	wire w_dff_A_kKb2a76c1_0;
	wire w_dff_A_a9hHyqNs9_0;
	wire w_dff_A_52yL5Oir8_0;
	wire w_dff_A_kMpLpclI6_0;
	wire w_dff_A_oucS8qp29_0;
	wire w_dff_A_ZYdeFAQq7_0;
	wire w_dff_A_sv5qDQit8_0;
	wire w_dff_A_cHT48gSs5_0;
	wire w_dff_A_Gzjyp4tK6_0;
	wire w_dff_A_8H9vCOIc4_0;
	wire w_dff_A_62FQUY7e9_0;
	wire w_dff_A_hrELfqsW8_0;
	wire w_dff_A_KDBF3E607_0;
	wire w_dff_A_ohHlkvwA4_0;
	wire w_dff_A_lVYVVi217_0;
	wire w_dff_A_ojj653AN2_0;
	wire w_dff_A_PzchLUhG1_0;
	wire w_dff_A_304jaEvm3_0;
	wire w_dff_A_8SnIt23R3_0;
	wire w_dff_A_2dkQMxX12_0;
	wire w_dff_A_sTkaVVIg9_0;
	wire w_dff_A_cQXSYRbY8_0;
	wire w_dff_A_zSo2aDVP3_0;
	wire w_dff_A_HPhFy2ab9_0;
	wire w_dff_A_3tdAzL8v3_0;
	wire w_dff_A_5FcrTReg5_0;
	wire w_dff_A_6eUgR59u9_0;
	wire w_dff_A_8CUDCYJB8_0;
	wire w_dff_A_nDsTolMs8_0;
	wire w_dff_A_R7vr0vRE3_0;
	wire w_dff_A_kgUuWbe53_0;
	wire w_dff_A_7NRKMlg45_0;
	wire w_dff_A_Y8H8L4Mh7_0;
	wire w_dff_A_9uTIdewM4_0;
	wire w_dff_A_5cH6oclo9_0;
	wire w_dff_A_VmwPEXiV7_0;
	wire w_dff_A_FmS0ciSa2_0;
	wire w_dff_A_RVgKvPYQ5_0;
	wire w_dff_A_1PDFdbZK4_0;
	wire w_dff_A_VMHJ3NcX1_0;
	wire w_dff_A_s5vgirpi1_0;
	wire w_dff_A_KozlldQB5_0;
	wire w_dff_A_fuQVxD3L5_0;
	wire w_dff_A_aO651zeA7_0;
	wire w_dff_A_mpVyZMfs2_0;
	wire w_dff_A_TjdUyd1m3_0;
	wire w_dff_A_hmaBXeqC7_0;
	wire w_dff_A_JhClA7XN6_0;
	wire w_dff_A_d1D5AJHx9_0;
	wire w_dff_A_R2OefjDr9_0;
	wire w_dff_A_2F0U9oUi3_0;
	wire w_dff_A_bCQyzGeO1_0;
	wire w_dff_A_EtvmkPLL6_0;
	wire w_dff_A_fnBrgqSm5_0;
	wire w_dff_A_aLbf6XPK1_2;
	wire w_dff_A_QaP3D5ZU3_0;
	wire w_dff_A_LjmKnrxD5_0;
	wire w_dff_A_ENeHB0fV4_0;
	wire w_dff_A_R54V7n3i8_0;
	wire w_dff_A_o52T4KMF8_0;
	wire w_dff_A_CvZlUgDk0_0;
	wire w_dff_A_GvQDGDh67_0;
	wire w_dff_A_bh2APSLp6_0;
	wire w_dff_A_DGYHpj5P7_0;
	wire w_dff_A_8TK6d1gG5_0;
	wire w_dff_A_sHry7NyT4_0;
	wire w_dff_A_IeOFZFFC1_0;
	wire w_dff_A_4eZgLYV21_0;
	wire w_dff_A_HXmEf8aN3_0;
	wire w_dff_A_KNF8iGyM1_0;
	wire w_dff_A_pPliMtAK0_0;
	wire w_dff_A_qSsHN3Ix4_0;
	wire w_dff_A_Ed2k6v438_0;
	wire w_dff_A_8rgolz4m2_0;
	wire w_dff_A_tLr9nbjR6_0;
	wire w_dff_A_x3AzODmj5_0;
	wire w_dff_A_QfUUn8bN6_0;
	wire w_dff_A_4HLVI9dQ5_0;
	wire w_dff_A_4s8PTElj1_0;
	wire w_dff_A_IAgpnSlD3_0;
	wire w_dff_A_yUAUJ1wR1_0;
	wire w_dff_A_xSNHOa6j7_0;
	wire w_dff_A_29fDN8L70_0;
	wire w_dff_A_tIPN73wT6_0;
	wire w_dff_A_Efcch7jW2_0;
	wire w_dff_A_xkCiVbQh7_0;
	wire w_dff_A_y6ohbpy86_0;
	wire w_dff_A_jQkCx8Dp7_0;
	wire w_dff_A_O4CF5uWf1_0;
	wire w_dff_A_yb2Ku54r4_0;
	wire w_dff_A_kEJvZqUP9_0;
	wire w_dff_A_YxJMjaIZ1_0;
	wire w_dff_A_JXwZ7n5C8_0;
	wire w_dff_A_GQ0A3ISV9_0;
	wire w_dff_A_PKYKLMPJ9_0;
	wire w_dff_A_w2qDXOxp3_0;
	wire w_dff_A_rhiqZhER5_0;
	wire w_dff_A_OaFrd7Qy4_0;
	wire w_dff_A_MB4GHscJ8_0;
	wire w_dff_A_RzZ07c8e1_0;
	wire w_dff_A_5Fx9KCuE9_0;
	wire w_dff_A_D37uXOCo7_0;
	wire w_dff_A_1nID5NdP6_0;
	wire w_dff_A_OoY8hnye1_0;
	wire w_dff_A_XUsa8Kup5_0;
	wire w_dff_A_DWsRDCbR6_0;
	wire w_dff_A_9gCRsJK16_0;
	wire w_dff_A_PzUR5csb4_0;
	wire w_dff_A_Qvmd2M0y3_0;
	wire w_dff_A_vBQUKRdX7_0;
	wire w_dff_A_cu0Bw0H98_0;
	wire w_dff_A_5IdgGGfG5_0;
	wire w_dff_A_8GlWDUqT0_0;
	wire w_dff_A_x1Lz4r392_0;
	wire w_dff_A_sjG6wrnR9_0;
	wire w_dff_A_K1mxTCAS4_0;
	wire w_dff_A_FNChFH696_0;
	wire w_dff_A_vopQHw7W8_2;
	wire w_dff_A_mFoBwehz9_0;
	wire w_dff_A_lpEAnQPX0_0;
	wire w_dff_A_k1XBAUvs0_0;
	wire w_dff_A_aDnyrkFj7_0;
	wire w_dff_A_8aONQoL34_0;
	wire w_dff_A_I6kKjmlw7_0;
	wire w_dff_A_9ddu3VGz6_0;
	wire w_dff_A_uFeY0ZwY9_0;
	wire w_dff_A_vrqJFr1D4_0;
	wire w_dff_A_mj9nnrBL8_0;
	wire w_dff_A_nAKHURSR4_0;
	wire w_dff_A_WAmUxhqR9_0;
	wire w_dff_A_iy2miqlv3_0;
	wire w_dff_A_31IDM0L67_0;
	wire w_dff_A_uUYaAqXH4_0;
	wire w_dff_A_yRdRrBuj7_0;
	wire w_dff_A_pWk8ihPO5_0;
	wire w_dff_A_SrPpZCxu8_0;
	wire w_dff_A_YxRUQL8A5_0;
	wire w_dff_A_xFDMzeuG3_0;
	wire w_dff_A_Wss4OJSK2_0;
	wire w_dff_A_tbOMpMK81_0;
	wire w_dff_A_dkf8Q8G94_0;
	wire w_dff_A_tKwFEqj33_0;
	wire w_dff_A_aDsSbgmo4_0;
	wire w_dff_A_EgsBPe6D2_0;
	wire w_dff_A_SZ00c0SZ2_0;
	wire w_dff_A_TwVRXF2y6_0;
	wire w_dff_A_jGUshw0S7_0;
	wire w_dff_A_BXzfYPKT0_0;
	wire w_dff_A_6M4fPLVj7_0;
	wire w_dff_A_DnJ8TZiW0_0;
	wire w_dff_A_iOdFmewz0_0;
	wire w_dff_A_OzQ2Ebdd0_0;
	wire w_dff_A_WOJr8laE8_0;
	wire w_dff_A_8AFyvlss7_0;
	wire w_dff_A_IpUk4VZL0_0;
	wire w_dff_A_z5vgm3J21_0;
	wire w_dff_A_jOe6T4Zy3_0;
	wire w_dff_A_uMbOQooM9_0;
	wire w_dff_A_6y1SwXfO1_0;
	wire w_dff_A_kI8w5MOE7_0;
	wire w_dff_A_b4Nm84XW8_0;
	wire w_dff_A_zRsSBkzh1_0;
	wire w_dff_A_Mg9D5fXL3_0;
	wire w_dff_A_kjm8Wqfw8_0;
	wire w_dff_A_b0En7ZcL2_0;
	wire w_dff_A_9vZ9g4sh5_0;
	wire w_dff_A_UFs2y91Z8_0;
	wire w_dff_A_4OtmtBbg9_0;
	wire w_dff_A_SGeC2zRk4_0;
	wire w_dff_A_Lo1pvlvF9_0;
	wire w_dff_A_jmE8YK7I1_0;
	wire w_dff_A_cPWEKegT1_0;
	wire w_dff_A_iWmkvgPp6_0;
	wire w_dff_A_0zhb5H5M3_0;
	wire w_dff_A_cfY3Mtns9_0;
	wire w_dff_A_9MDZ3hWf6_0;
	wire w_dff_A_6RkZudg36_0;
	wire w_dff_A_xPsKA8QQ4_2;
	wire w_dff_A_VtaktCyZ6_0;
	wire w_dff_A_TpZoPvat8_0;
	wire w_dff_A_tNbZIGhQ7_0;
	wire w_dff_A_HRd7yJal4_0;
	wire w_dff_A_zIfZ8yh84_0;
	wire w_dff_A_mHBE1IYC9_0;
	wire w_dff_A_IrB2qO3r4_0;
	wire w_dff_A_eJ66f0YT0_0;
	wire w_dff_A_nhzZEO2k6_0;
	wire w_dff_A_ddUKiAET7_0;
	wire w_dff_A_ZvWBmQti6_0;
	wire w_dff_A_0tMGJ2us5_0;
	wire w_dff_A_uuxNTB2n0_0;
	wire w_dff_A_dSX1gFKq9_0;
	wire w_dff_A_L4P54gpI0_0;
	wire w_dff_A_9uzdJkUP9_0;
	wire w_dff_A_yiuPU3LY2_0;
	wire w_dff_A_LQfmxIMN5_0;
	wire w_dff_A_1QeAzK8O0_0;
	wire w_dff_A_ZirUxbJy9_0;
	wire w_dff_A_a9z1lfKH1_0;
	wire w_dff_A_BCRZdo1t0_0;
	wire w_dff_A_y5odsYue8_0;
	wire w_dff_A_etjNtSsz3_0;
	wire w_dff_A_fsiO41dQ7_0;
	wire w_dff_A_SxwruHad3_0;
	wire w_dff_A_NLAVcwWt9_0;
	wire w_dff_A_21jvGW8Y0_0;
	wire w_dff_A_BjOUEZux0_0;
	wire w_dff_A_0euBjbWc6_0;
	wire w_dff_A_EKGJ3hDJ1_0;
	wire w_dff_A_WpFJcSxo9_0;
	wire w_dff_A_0DEEoLFt8_0;
	wire w_dff_A_3CxfT8b73_0;
	wire w_dff_A_fOrt9ejS3_0;
	wire w_dff_A_I3sMw07c3_0;
	wire w_dff_A_3yLcQN5i9_0;
	wire w_dff_A_goBP1uOm8_0;
	wire w_dff_A_9HQ5FCA44_0;
	wire w_dff_A_oqiLpstc0_0;
	wire w_dff_A_CxWcVPBl4_0;
	wire w_dff_A_SJkGpVdc0_0;
	wire w_dff_A_jmZeOd3P8_0;
	wire w_dff_A_PxTx5HK61_0;
	wire w_dff_A_aqfX5RqX1_0;
	wire w_dff_A_Ulav9pLt5_0;
	wire w_dff_A_UKs76Q702_0;
	wire w_dff_A_KQWdSDpY3_0;
	wire w_dff_A_RQzzZAYD7_0;
	wire w_dff_A_a41ksy7G6_0;
	wire w_dff_A_fn4jRplA1_0;
	wire w_dff_A_FChtwYNV6_0;
	wire w_dff_A_Km7j8Yhc0_0;
	wire w_dff_A_wF9lnkhh2_0;
	wire w_dff_A_hyne3PJx7_0;
	wire w_dff_A_r2P9juUz5_0;
	wire w_dff_A_ByNtDrk64_2;
	wire w_dff_A_MOy45Gta4_0;
	wire w_dff_A_5Tx3mpaO2_0;
	wire w_dff_A_8TC1SORo5_0;
	wire w_dff_A_onfZaWLE0_0;
	wire w_dff_A_aVugbHoH2_0;
	wire w_dff_A_ghdKFs9E3_0;
	wire w_dff_A_cOxkFxM15_0;
	wire w_dff_A_s1VdefxO8_0;
	wire w_dff_A_GqlkSCUu6_0;
	wire w_dff_A_y6rU666g2_0;
	wire w_dff_A_KqlqJ8e55_0;
	wire w_dff_A_BjBnoNwL7_0;
	wire w_dff_A_h9whmFh97_0;
	wire w_dff_A_pxFwMPUY1_0;
	wire w_dff_A_qeH9taZC0_0;
	wire w_dff_A_vmW6vxdh5_0;
	wire w_dff_A_Ayckzlpl6_0;
	wire w_dff_A_pIwsWaUa8_0;
	wire w_dff_A_O8hG4fWQ0_0;
	wire w_dff_A_Q5jClSu92_0;
	wire w_dff_A_Lns7Ijju7_0;
	wire w_dff_A_uWQ2yjvK6_0;
	wire w_dff_A_KMyGcg4b7_0;
	wire w_dff_A_G45DwoiU0_0;
	wire w_dff_A_9qtxAklF2_0;
	wire w_dff_A_qnEAhHQt3_0;
	wire w_dff_A_pIaS6yfF6_0;
	wire w_dff_A_y4X44ksk0_0;
	wire w_dff_A_RwLuFJSC5_0;
	wire w_dff_A_2PPGMt3j5_0;
	wire w_dff_A_FFA0ajUg8_0;
	wire w_dff_A_r9hNANWG7_0;
	wire w_dff_A_yB5jntl06_0;
	wire w_dff_A_vSW29hvO5_0;
	wire w_dff_A_ghCvYGAd8_0;
	wire w_dff_A_GbNOzueq6_0;
	wire w_dff_A_QJRJU3N02_0;
	wire w_dff_A_yXVuvWgT5_0;
	wire w_dff_A_9Qz7LQBP5_0;
	wire w_dff_A_TmM8lxpT3_0;
	wire w_dff_A_qLkWJwRB1_0;
	wire w_dff_A_krxee2Uc9_0;
	wire w_dff_A_UfKtTvOK1_0;
	wire w_dff_A_AWGoDzqR1_0;
	wire w_dff_A_vxcXAnTc6_0;
	wire w_dff_A_6902Kq5q3_0;
	wire w_dff_A_0zMcmGsi4_0;
	wire w_dff_A_mTmxVBjj2_0;
	wire w_dff_A_J4dk22Yl9_0;
	wire w_dff_A_4CdmSuGL9_0;
	wire w_dff_A_nHWK10bh2_0;
	wire w_dff_A_8VRwnKMI3_0;
	wire w_dff_A_MQl52QAR1_0;
	wire w_dff_A_nMXYqaCW1_2;
	wire w_dff_A_YYpgINDy3_0;
	wire w_dff_A_lwrrrB3p7_0;
	wire w_dff_A_B8fJ0ntx2_0;
	wire w_dff_A_YjvteGTd2_0;
	wire w_dff_A_yaTgu2VO1_0;
	wire w_dff_A_SEcWP5OR6_0;
	wire w_dff_A_D1OXEpw21_0;
	wire w_dff_A_v8GX5eHi7_0;
	wire w_dff_A_ZUHgF6Eb5_0;
	wire w_dff_A_u6QIqdzu5_0;
	wire w_dff_A_o5NFb3Ii8_0;
	wire w_dff_A_35zqimbM6_0;
	wire w_dff_A_kusZDYTx2_0;
	wire w_dff_A_cgnjCkye7_0;
	wire w_dff_A_Y0bRhwzn5_0;
	wire w_dff_A_JdIDhnLx5_0;
	wire w_dff_A_jsWGIM580_0;
	wire w_dff_A_Z9J2BnBh3_0;
	wire w_dff_A_izzOODcx7_0;
	wire w_dff_A_vyoYzxX94_0;
	wire w_dff_A_r4KHrzwQ1_0;
	wire w_dff_A_JrmBbtdJ8_0;
	wire w_dff_A_M6jBHEeD8_0;
	wire w_dff_A_y10g4YGS6_0;
	wire w_dff_A_nHcE0DUg9_0;
	wire w_dff_A_0BhYfPlQ7_0;
	wire w_dff_A_ywoydGKi4_0;
	wire w_dff_A_FeWTgB8k8_0;
	wire w_dff_A_yNnk6Uvw5_0;
	wire w_dff_A_9QLcHwXy2_0;
	wire w_dff_A_96No0DOe8_0;
	wire w_dff_A_TbQglCN53_0;
	wire w_dff_A_pI0ROOVO7_0;
	wire w_dff_A_19zbZyDP2_0;
	wire w_dff_A_wtQSMymi6_0;
	wire w_dff_A_pNM5oZap1_0;
	wire w_dff_A_OZvvVaKl1_0;
	wire w_dff_A_PzCWopPt7_0;
	wire w_dff_A_9S4vkzzc3_0;
	wire w_dff_A_Qi5Sacb09_0;
	wire w_dff_A_LLzdCRSK6_0;
	wire w_dff_A_8C7GdqWL1_0;
	wire w_dff_A_fcA96LoP8_0;
	wire w_dff_A_dTCWqSlQ2_0;
	wire w_dff_A_R0aARRQc7_0;
	wire w_dff_A_5Mm8Y8dt2_0;
	wire w_dff_A_Idj8UVp15_0;
	wire w_dff_A_Rdzpgkfa3_0;
	wire w_dff_A_ykGrHtUK1_0;
	wire w_dff_A_Er4tz4if6_0;
	wire w_dff_A_jS7LkhAz1_2;
	wire w_dff_A_rYdq5y3o6_0;
	wire w_dff_A_aNacdnhV0_0;
	wire w_dff_A_YpzLEucd6_0;
	wire w_dff_A_hGThfReO3_0;
	wire w_dff_A_qRNHv9At6_0;
	wire w_dff_A_11EZkWzy2_0;
	wire w_dff_A_95CyLDFD7_0;
	wire w_dff_A_L1mesjpJ0_0;
	wire w_dff_A_YbnuNaDi3_0;
	wire w_dff_A_D9Wqwrpl1_0;
	wire w_dff_A_Dmrc0wNa9_0;
	wire w_dff_A_9Vst5bMJ3_0;
	wire w_dff_A_btsBmhzI6_0;
	wire w_dff_A_P8hvuDZx6_0;
	wire w_dff_A_fpSGDsJV3_0;
	wire w_dff_A_JPcHcMZo9_0;
	wire w_dff_A_AHEyVeYx6_0;
	wire w_dff_A_CaUtmfT38_0;
	wire w_dff_A_OTz6aHL36_0;
	wire w_dff_A_7E1PTGuK9_0;
	wire w_dff_A_JxfX8zAx4_0;
	wire w_dff_A_4ogO21bK2_0;
	wire w_dff_A_mrEdarCm7_0;
	wire w_dff_A_e1XVe4sA1_0;
	wire w_dff_A_tH9kGI2s0_0;
	wire w_dff_A_L5zbAgZ49_0;
	wire w_dff_A_UbOOOFqZ1_0;
	wire w_dff_A_FKG7jUTr7_0;
	wire w_dff_A_fhSc2Xbt9_0;
	wire w_dff_A_bYyJYapF5_0;
	wire w_dff_A_bMoVnqGV3_0;
	wire w_dff_A_3fh4P4QS4_0;
	wire w_dff_A_aWvbuDCF3_0;
	wire w_dff_A_PFEd0Xos4_0;
	wire w_dff_A_e6iNcabG9_0;
	wire w_dff_A_eUgayTAz1_0;
	wire w_dff_A_FHm4QNY21_0;
	wire w_dff_A_0q13euX98_0;
	wire w_dff_A_IR2pIF1V0_0;
	wire w_dff_A_BPW7a3Os3_0;
	wire w_dff_A_dyBO7idN3_0;
	wire w_dff_A_fHtNZdYZ2_0;
	wire w_dff_A_x2JstJLm6_0;
	wire w_dff_A_KfmLhOCS4_0;
	wire w_dff_A_RqhStVCN8_0;
	wire w_dff_A_rfkhjkw56_0;
	wire w_dff_A_TsEFZypi0_0;
	wire w_dff_A_jXnwwKqc6_2;
	wire w_dff_A_EyhkW8kI9_0;
	wire w_dff_A_HHYTkiHh7_0;
	wire w_dff_A_pr4g7m6B6_0;
	wire w_dff_A_2sMFBNzG1_0;
	wire w_dff_A_YFyweRcv5_0;
	wire w_dff_A_3KCa8cg62_0;
	wire w_dff_A_dBclAjSs5_0;
	wire w_dff_A_OGYqzOkd6_0;
	wire w_dff_A_DlFXrXBO9_0;
	wire w_dff_A_lz2DAHkv1_0;
	wire w_dff_A_foRu15oU4_0;
	wire w_dff_A_N6AyBItT9_0;
	wire w_dff_A_jDlaZ5oN0_0;
	wire w_dff_A_4k5Arbv01_0;
	wire w_dff_A_wrJKIFmZ3_0;
	wire w_dff_A_eOHTfR564_0;
	wire w_dff_A_dpkBOj0d6_0;
	wire w_dff_A_zeFohYIq0_0;
	wire w_dff_A_m1RaIO4f8_0;
	wire w_dff_A_4sTr0x073_0;
	wire w_dff_A_lhDRANhY5_0;
	wire w_dff_A_U97lU8Df2_0;
	wire w_dff_A_cTpNyUj90_0;
	wire w_dff_A_85YsmSJS4_0;
	wire w_dff_A_Wi2L1H9b2_0;
	wire w_dff_A_32JurMhH5_0;
	wire w_dff_A_q6kNwUVp2_0;
	wire w_dff_A_VKwdWK2t8_0;
	wire w_dff_A_YCY0nPRx8_0;
	wire w_dff_A_DeD0Xxjt4_0;
	wire w_dff_A_aTOxYAW03_0;
	wire w_dff_A_5iGNlgD84_0;
	wire w_dff_A_LOCMHPqz1_0;
	wire w_dff_A_fuEUCixC4_0;
	wire w_dff_A_YcGhvpYK5_0;
	wire w_dff_A_Kq8QgNPy8_0;
	wire w_dff_A_IDge9Oud0_0;
	wire w_dff_A_NafXWdyD9_0;
	wire w_dff_A_moFZvKrK4_0;
	wire w_dff_A_jlJU8G6u5_0;
	wire w_dff_A_XEIVmxyX6_0;
	wire w_dff_A_J2NaBzCs1_0;
	wire w_dff_A_eYorYIE99_0;
	wire w_dff_A_0P7PXjZ73_0;
	wire w_dff_A_InJoAco86_2;
	wire w_dff_A_8tFjG5Nu4_0;
	wire w_dff_A_adZFhVWt3_0;
	wire w_dff_A_khQeFtbi2_0;
	wire w_dff_A_pawRfK1G2_0;
	wire w_dff_A_lHQnDnJv7_0;
	wire w_dff_A_kiy4hM7B1_0;
	wire w_dff_A_WZQwmKDJ9_0;
	wire w_dff_A_oeFFh1Qd8_0;
	wire w_dff_A_KNo4ep9N4_0;
	wire w_dff_A_LFG5QP5K3_0;
	wire w_dff_A_4wOkTt5C8_0;
	wire w_dff_A_7VtlChLr7_0;
	wire w_dff_A_VteV8FS84_0;
	wire w_dff_A_tlx0rhtQ9_0;
	wire w_dff_A_92ta0ssu8_0;
	wire w_dff_A_AEKKLIYV7_0;
	wire w_dff_A_0ixeKnDn9_0;
	wire w_dff_A_PqXnSlV98_0;
	wire w_dff_A_lgn9l7ch1_0;
	wire w_dff_A_KpNFLpMX4_0;
	wire w_dff_A_aWKhFH2m5_0;
	wire w_dff_A_VZdekvL53_0;
	wire w_dff_A_tAEldFgU2_0;
	wire w_dff_A_GUwmpE9s6_0;
	wire w_dff_A_AdUBg0mg6_0;
	wire w_dff_A_rP6G0iiV7_0;
	wire w_dff_A_kRm8IWAG9_0;
	wire w_dff_A_zknHFImh4_0;
	wire w_dff_A_bjuChTcd4_0;
	wire w_dff_A_Py5PRoml6_0;
	wire w_dff_A_XYMOkY597_0;
	wire w_dff_A_pgIJinxr2_0;
	wire w_dff_A_gR9x8sir8_0;
	wire w_dff_A_mTznjd3V1_0;
	wire w_dff_A_po6byZm51_0;
	wire w_dff_A_NkEXzxnV6_0;
	wire w_dff_A_bRrItFUZ7_0;
	wire w_dff_A_Z4r2umF19_0;
	wire w_dff_A_w9Y5PU9q1_0;
	wire w_dff_A_53xL7dgN4_0;
	wire w_dff_A_mocf161Y5_0;
	wire w_dff_A_XOoOUeVN7_2;
	wire w_dff_A_2XzYw5Sx7_0;
	wire w_dff_A_54or12fq0_0;
	wire w_dff_A_OWIeZrdq8_0;
	wire w_dff_A_3RK770oa1_0;
	wire w_dff_A_vMMXiNqg9_0;
	wire w_dff_A_ELqyL6p15_0;
	wire w_dff_A_ubsyBGdE0_0;
	wire w_dff_A_pHQzrwBN7_0;
	wire w_dff_A_X9yQ8z6n0_0;
	wire w_dff_A_xTgPQv3V5_0;
	wire w_dff_A_37HwXmjE4_0;
	wire w_dff_A_aNyO50tc7_0;
	wire w_dff_A_dRVfjY9J9_0;
	wire w_dff_A_OURD4cKj9_0;
	wire w_dff_A_tD30K2Zm8_0;
	wire w_dff_A_86Ws02WH4_0;
	wire w_dff_A_BWIjOuxE1_0;
	wire w_dff_A_GJAHJOxT4_0;
	wire w_dff_A_dyiAxvMi1_0;
	wire w_dff_A_cXVsAY8B3_0;
	wire w_dff_A_m1o9RK7j9_0;
	wire w_dff_A_G0pxffjw2_0;
	wire w_dff_A_vnjbYvWV6_0;
	wire w_dff_A_MSSxBnnR7_0;
	wire w_dff_A_u6Pp6xdQ7_0;
	wire w_dff_A_jFP94YyL3_0;
	wire w_dff_A_IrK5KcnO6_0;
	wire w_dff_A_0URgGxv48_0;
	wire w_dff_A_WCz3bCSs5_0;
	wire w_dff_A_Is2VsdUM2_0;
	wire w_dff_A_K1iWiehT4_0;
	wire w_dff_A_zA4Jzm3R2_0;
	wire w_dff_A_9AqNdbqI6_0;
	wire w_dff_A_ds57DFHj0_0;
	wire w_dff_A_AbnSA8Wv8_0;
	wire w_dff_A_fGrLnsBi1_0;
	wire w_dff_A_QCqrNgOf5_0;
	wire w_dff_A_DXzQ8kFL2_0;
	wire w_dff_A_2eploXL89_2;
	wire w_dff_A_UdC9gNAX3_0;
	wire w_dff_A_5FU17UXK0_0;
	wire w_dff_A_rXGbqFUD2_0;
	wire w_dff_A_JKUfwg6E9_0;
	wire w_dff_A_zJDzzZVk4_0;
	wire w_dff_A_raXzRdUI4_0;
	wire w_dff_A_P1LIRME81_0;
	wire w_dff_A_12yhYJn96_0;
	wire w_dff_A_R5faY6Ud2_0;
	wire w_dff_A_PzJMzCiL0_0;
	wire w_dff_A_8SeXCYUG5_0;
	wire w_dff_A_L3rDwbIB9_0;
	wire w_dff_A_VIsmJmRc0_0;
	wire w_dff_A_0qff5Z2H6_0;
	wire w_dff_A_mCB9qQjo0_0;
	wire w_dff_A_XSjJk7rX7_0;
	wire w_dff_A_1CRZe30o4_0;
	wire w_dff_A_QsA7PpOn5_0;
	wire w_dff_A_5UOx81rq2_0;
	wire w_dff_A_8Se1HEYT5_0;
	wire w_dff_A_BYiFPuHT0_0;
	wire w_dff_A_vEpqnFMt4_0;
	wire w_dff_A_vCxMsaqY4_0;
	wire w_dff_A_832snTKX6_0;
	wire w_dff_A_slnmOMLo7_0;
	wire w_dff_A_FxSLtNzd0_0;
	wire w_dff_A_y1ewrchc5_0;
	wire w_dff_A_wWB6wqIg1_0;
	wire w_dff_A_iTNRMvBc4_0;
	wire w_dff_A_U1rrjxAt8_0;
	wire w_dff_A_5AQSyvdS8_0;
	wire w_dff_A_wCpHk9zz9_0;
	wire w_dff_A_7g3GfLQ00_0;
	wire w_dff_A_LFKCZbbW1_0;
	wire w_dff_A_FbP4X9Z62_0;
	wire w_dff_A_Y7aiHoy19_2;
	wire w_dff_A_HJm9H9L25_0;
	wire w_dff_A_Xkr3vQ0J9_0;
	wire w_dff_A_L028gl8T8_0;
	wire w_dff_A_dfwW0gsq6_0;
	wire w_dff_A_Lv2BQzXU1_0;
	wire w_dff_A_6ZHXvjvc4_0;
	wire w_dff_A_auGLRn7K2_0;
	wire w_dff_A_R7GgadRq3_0;
	wire w_dff_A_9H7xgTXh8_0;
	wire w_dff_A_Z5YGKIa88_0;
	wire w_dff_A_7aUXMkwn7_0;
	wire w_dff_A_QGce68b84_0;
	wire w_dff_A_OVGBUYaL5_0;
	wire w_dff_A_9gXgKaXw0_0;
	wire w_dff_A_Ejheg2bu0_0;
	wire w_dff_A_NCiURC5E0_0;
	wire w_dff_A_BjBWmdEn8_0;
	wire w_dff_A_uPUZ9dsM6_0;
	wire w_dff_A_aYyvOcxe5_0;
	wire w_dff_A_Nct9yvsP4_0;
	wire w_dff_A_XGldcTk53_0;
	wire w_dff_A_jiqcNkw18_0;
	wire w_dff_A_VpvSj5dJ7_0;
	wire w_dff_A_ZtyUiTBv8_0;
	wire w_dff_A_cOrt3WrE8_0;
	wire w_dff_A_2ZSKEUyj8_0;
	wire w_dff_A_RqyyAWIx9_0;
	wire w_dff_A_wErVqJat2_0;
	wire w_dff_A_gPzvwB2F7_0;
	wire w_dff_A_zVweBWe90_0;
	wire w_dff_A_tqURTRsT5_0;
	wire w_dff_A_UyeQsIq00_0;
	wire w_dff_A_wIpjPOmp5_2;
	wire w_dff_A_AtNUbuPZ6_0;
	wire w_dff_A_BJinPbYE0_0;
	wire w_dff_A_m8BbU3kq9_0;
	wire w_dff_A_gYrjFtuP1_0;
	wire w_dff_A_qYnAGmuk8_0;
	wire w_dff_A_SjvbUbv44_0;
	wire w_dff_A_4HVpanFh3_0;
	wire w_dff_A_dOzpNVyM5_0;
	wire w_dff_A_oKk0otOe0_0;
	wire w_dff_A_z7oGsaG63_0;
	wire w_dff_A_S6k56uct6_0;
	wire w_dff_A_aazInrlM5_0;
	wire w_dff_A_GAW4iidl0_0;
	wire w_dff_A_dyvtR10S5_0;
	wire w_dff_A_S4sEj3uH1_0;
	wire w_dff_A_44n3h7Zq3_0;
	wire w_dff_A_i5zczjgk3_0;
	wire w_dff_A_YffjuMFx5_0;
	wire w_dff_A_LOi9yVsM4_0;
	wire w_dff_A_To8wRyRH4_0;
	wire w_dff_A_Raho7Dv51_0;
	wire w_dff_A_TgRyoHRk7_0;
	wire w_dff_A_xcMEHyMM7_0;
	wire w_dff_A_LR86UzAt5_0;
	wire w_dff_A_uLTMz8aG0_0;
	wire w_dff_A_9MW6V2Xb8_0;
	wire w_dff_A_DSmQh9sG8_0;
	wire w_dff_A_aRvqhXWD3_0;
	wire w_dff_A_ds6SS5sf0_0;
	wire w_dff_A_UloyOVAB2_2;
	wire w_dff_A_Ibwud07n3_0;
	wire w_dff_A_o2tDNQ8L1_0;
	wire w_dff_A_cYTGn0w85_0;
	wire w_dff_A_UFDwGYHv6_0;
	wire w_dff_A_hHgul19L0_0;
	wire w_dff_A_LxKvx0D30_0;
	wire w_dff_A_cVgx0giF9_0;
	wire w_dff_A_GJ77rgCE8_0;
	wire w_dff_A_qWSMzihb6_0;
	wire w_dff_A_gCAghKsR7_0;
	wire w_dff_A_fOl9z5zx4_0;
	wire w_dff_A_TsmY1Nzz1_0;
	wire w_dff_A_2FglyBmi3_0;
	wire w_dff_A_DREhNRDh2_0;
	wire w_dff_A_bE73Pfdf2_0;
	wire w_dff_A_jcKUJfu46_0;
	wire w_dff_A_GeOOR1Kw8_0;
	wire w_dff_A_lcIhxg9N3_0;
	wire w_dff_A_ElhITZKE8_0;
	wire w_dff_A_o2wrKTho2_0;
	wire w_dff_A_xOGH776w5_0;
	wire w_dff_A_9WEhy4VH4_0;
	wire w_dff_A_Ds88u79W7_0;
	wire w_dff_A_AJXQP84v1_0;
	wire w_dff_A_GTAKWQ9M5_0;
	wire w_dff_A_tWXmNiTj5_0;
	wire w_dff_A_NsXp71H74_0;
	wire w_dff_A_JVdXQdwf8_2;
	wire w_dff_A_1zH06zMy1_0;
	wire w_dff_A_x3873p1D6_0;
	wire w_dff_A_kmw9SK7V6_0;
	wire w_dff_A_PRf3HOJn2_0;
	wire w_dff_A_2KmzX7Ao7_0;
	wire w_dff_A_HmgcqW901_0;
	wire w_dff_A_gOZAnXRZ1_0;
	wire w_dff_A_wGEJkh7A6_0;
	wire w_dff_A_b388iv6w3_0;
	wire w_dff_A_GDfxKoOG2_0;
	wire w_dff_A_0yI39X0Y7_0;
	wire w_dff_A_T2NoHBtC4_0;
	wire w_dff_A_f2cnQIQF6_0;
	wire w_dff_A_NutVUu4T7_0;
	wire w_dff_A_1JVCAbvN6_0;
	wire w_dff_A_vlOyO0CB5_0;
	wire w_dff_A_UflzVYxz0_0;
	wire w_dff_A_H3lqwzVH4_0;
	wire w_dff_A_3NCNoKhF9_0;
	wire w_dff_A_kKO7wThK9_0;
	wire w_dff_A_7RolqyXH1_0;
	wire w_dff_A_2liRurwf0_0;
	wire w_dff_A_kvydyW6B5_0;
	wire w_dff_A_mEJGlNto5_0;
	wire w_dff_A_bu2MqwBY3_0;
	wire w_dff_A_CyfQuo9O5_2;
	wire w_dff_A_6QsmgJCT4_0;
	wire w_dff_A_QLgpwxGr1_0;
	wire w_dff_A_OhEcXmMH6_0;
	wire w_dff_A_f0sM1qhK3_0;
	wire w_dff_A_bKDVYeOx0_0;
	wire w_dff_A_7fgkbALf7_0;
	wire w_dff_A_TzUaa2e52_0;
	wire w_dff_A_pumQyfY82_0;
	wire w_dff_A_KTleP3A94_0;
	wire w_dff_A_67r9RmrV8_0;
	wire w_dff_A_LWKSoOGR7_0;
	wire w_dff_A_gzmOcQbw7_0;
	wire w_dff_A_o5JiHedi3_0;
	wire w_dff_A_F6Qgon7N7_0;
	wire w_dff_A_AKaExpA45_0;
	wire w_dff_A_rSedN8Au7_0;
	wire w_dff_A_c36Gp4Km5_0;
	wire w_dff_A_lSJDeB477_0;
	wire w_dff_A_Kahl07kv5_0;
	wire w_dff_A_w7zOwIuP6_0;
	wire w_dff_A_FM5DeNXp3_0;
	wire w_dff_A_2KiYTUpU1_0;
	wire w_dff_A_sD0cSjtY8_0;
	wire w_dff_A_PzmSJC3Q3_0;
	wire w_dff_A_MLPL8Tm53_2;
	wire w_dff_A_1cUE5gY61_0;
	wire w_dff_A_Nx2zFIdU0_0;
	wire w_dff_A_YbuSdF7k1_0;
	wire w_dff_A_PliTLY538_0;
	wire w_dff_A_IGbAi8d80_0;
	wire w_dff_A_g2HGkiKj8_0;
	wire w_dff_A_5tgjmMIm3_0;
	wire w_dff_A_SHFAsCLF7_0;
	wire w_dff_A_hGGFY9fF8_0;
	wire w_dff_A_R0UyvXsu2_0;
	wire w_dff_A_Dczdn4nl2_0;
	wire w_dff_A_QhXh7hU81_0;
	wire w_dff_A_Gv9ZysSp0_0;
	wire w_dff_A_gDevGOR13_0;
	wire w_dff_A_p0BmH3YN4_0;
	wire w_dff_A_VATKnVjT6_0;
	wire w_dff_A_h0gD6GjZ9_0;
	wire w_dff_A_vziCFJVO1_0;
	wire w_dff_A_Zy7WuMtb2_0;
	wire w_dff_A_aUNKkEc46_0;
	wire w_dff_A_PLHlw61x0_0;
	wire w_dff_A_OOLKuQoX2_0;
	wire w_dff_A_n713uqzH6_2;
	wire w_dff_A_1zyePD0k0_0;
	wire w_dff_A_8EkLrFWD9_0;
	wire w_dff_A_mkIIKsEY7_0;
	wire w_dff_A_VsZYpE2W6_0;
	wire w_dff_A_uG58UR1Y7_0;
	wire w_dff_A_37vdwpRh7_0;
	wire w_dff_A_2VlvsQ2N5_0;
	wire w_dff_A_G4rarnNb2_0;
	wire w_dff_A_bFGW1Aob9_0;
	wire w_dff_A_n1RWEHcT4_0;
	wire w_dff_A_Q1Hj46AI5_0;
	wire w_dff_A_2r7e5l4a2_0;
	wire w_dff_A_XKnSYu4M6_0;
	wire w_dff_A_K1QTPPHV9_0;
	wire w_dff_A_RRmvn2mA0_0;
	wire w_dff_A_Qp7kegdR0_0;
	wire w_dff_A_SxJHOqFh5_0;
	wire w_dff_A_7GqKYvYY1_0;
	wire w_dff_A_yCy4gWd84_0;
	wire w_dff_A_IR1hYRdO8_0;
	wire w_dff_A_uHImcr829_2;
	wire w_dff_A_PuntIyzd3_0;
	wire w_dff_A_9hC8YyDW0_0;
	wire w_dff_A_MAVKxQfy9_0;
	wire w_dff_A_OU1juCpu3_0;
	wire w_dff_A_vQsYsFQ84_0;
	wire w_dff_A_6JaZ3H5x0_0;
	wire w_dff_A_L0aAgzoy5_0;
	wire w_dff_A_YqFbGUtE6_0;
	wire w_dff_A_3chAuc6C7_0;
	wire w_dff_A_gJqYnwRf4_0;
	wire w_dff_A_HyR4pv8i8_0;
	wire w_dff_A_H31sQU3z4_0;
	wire w_dff_A_VXuuPWYE1_0;
	wire w_dff_A_cEQ7hE1d9_0;
	wire w_dff_A_fWBN7M7R5_0;
	wire w_dff_A_3IpZdmmt8_0;
	wire w_dff_A_fsnear8F0_0;
	wire w_dff_A_peG6gmsc2_0;
	wire w_dff_A_IVpIwNKv9_2;
	wire w_dff_A_6hil7dpQ8_0;
	wire w_dff_A_z9BO7XGP7_0;
	wire w_dff_A_iC1YrsCy7_0;
	wire w_dff_A_DvFndVcE9_0;
	wire w_dff_A_ODlpoHVs5_0;
	wire w_dff_A_XfuX7JNC6_0;
	wire w_dff_A_xbvxqzN21_0;
	wire w_dff_A_HqOzHMBf3_0;
	wire w_dff_A_qWw2ImB81_0;
	wire w_dff_A_MTKcdpiO3_0;
	wire w_dff_A_ybVgRRSY6_0;
	wire w_dff_A_iGfZIBto7_0;
	wire w_dff_A_EKf6nyf00_0;
	wire w_dff_A_3bgR5Esy3_0;
	wire w_dff_A_HgzcCpoD4_0;
	wire w_dff_A_qEnI3H503_0;
	wire w_dff_A_J9KkTH2x8_2;
	wire w_dff_A_3TFql5wV6_0;
	wire w_dff_A_Cg14zy3H6_0;
	wire w_dff_A_TKmPl4h12_0;
	wire w_dff_A_BMz3zrYF4_0;
	wire w_dff_A_xjsRzz3e0_0;
	wire w_dff_A_HPuBL4Zj8_0;
	wire w_dff_A_rAePVV5H4_0;
	wire w_dff_A_GC3C7Ipp8_0;
	wire w_dff_A_XICinNMW7_0;
	wire w_dff_A_jWnHqDMP3_0;
	wire w_dff_A_7YPS7KFr9_0;
	wire w_dff_A_vqTTAhJa6_0;
	wire w_dff_A_TI6FyUpQ0_0;
	wire w_dff_A_MzFxhQaF3_0;
	wire w_dff_A_SiAvJkIH2_2;
	wire w_dff_A_DMQvcXa57_0;
	wire w_dff_A_iaGQDlki6_0;
	wire w_dff_A_C5FUBbPf2_0;
	wire w_dff_A_Jirr21g67_0;
	wire w_dff_A_5cSz67HW5_0;
	wire w_dff_A_pVwqnoch6_0;
	wire w_dff_A_jPJSMjq68_0;
	wire w_dff_A_CzVrvDbH0_0;
	wire w_dff_A_sNlDG9Kl8_0;
	wire w_dff_A_CKVihfhb3_0;
	wire w_dff_A_OxoA2Dmw7_0;
	wire w_dff_A_MJmxjNUa6_0;
	wire w_dff_A_iPOTMMlN8_2;
	wire w_dff_A_Mcel7Ici0_0;
	wire w_dff_A_mLuGV0qZ8_0;
	wire w_dff_A_RTLILm7e3_0;
	wire w_dff_A_PguZKwg88_0;
	wire w_dff_A_NUqmzJqp4_0;
	wire w_dff_A_q8EXGjNW0_0;
	wire w_dff_A_z8DsJDDU7_0;
	wire w_dff_A_1SYlCHVO7_0;
	wire w_dff_A_KvCKM18V3_0;
	wire w_dff_A_HmcJ3q5s3_0;
	wire w_dff_A_ZynMqCJa0_2;
	wire w_dff_A_EfzsPbLb3_0;
	wire w_dff_A_lzkEW5DO4_0;
	wire w_dff_A_T3BcHT3C2_0;
	wire w_dff_A_hHw8iqDQ9_0;
	wire w_dff_A_LH6lzpir2_0;
	wire w_dff_A_Wl1wMhsX8_0;
	wire w_dff_A_O7PPRNrY9_0;
	wire w_dff_A_aqTIs5RT3_0;
	wire w_dff_A_DQBFPbwp8_2;
	wire w_dff_A_7Eum09t90_0;
	wire w_dff_A_1DK9Zo400_0;
	wire w_dff_A_u1PNOSYe3_0;
	wire w_dff_A_brfkCIms5_0;
	wire w_dff_A_GclQeXAU6_0;
	wire w_dff_A_Tyc7mDF21_0;
	wire w_dff_A_6HD4c7010_2;
	wire w_dff_A_H101jjJm2_0;
	wire w_dff_A_iCKC4Clq9_0;
	wire w_dff_A_NHm2bFxY2_0;
	wire w_dff_A_equOPP612_0;
	wire w_dff_A_onIovUsr0_2;
	wire w_dff_A_ghfVfWMO9_0;
	wire w_dff_A_SMJRn6R92_0;
	wire w_dff_A_mVaqxWQK4_2;
	jand g0000(.dina(w_G273gat_7[1]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G290gat_7[2]),.dinb(w_G18gat_7[1]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_n65_0[1]),.dinb(w_G545gat_0),.dout(n66),.clk(gclk));
	jnot g0003(.din(w_n66_0[1]),.dout(n67),.clk(gclk));
	jnot g0004(.din(w_G18gat_7[0]),.dout(n68),.clk(gclk));
	jnot g0005(.din(w_G273gat_7[0]),.dout(n69),.clk(gclk));
	jor g0006(.dina(w_n69_0[1]),.dinb(n68),.dout(n70),.clk(gclk));
	jnot g0007(.din(w_n70_0[1]),.dout(n71),.clk(gclk));
	jand g0008(.dina(w_G290gat_7[1]),.dinb(w_G1gat_7[0]),.dout(n72),.clk(gclk));
	jor g0009(.dina(w_dff_B_SUExNrn46_0),.dinb(n71),.dout(n73),.clk(gclk));
	jand g0010(.dina(n73),.dinb(w_n67_0[1]),.dout(w_dff_A_NslXWg0x3_2),.clk(gclk));
	jand g0011(.dina(w_G307gat_7[1]),.dinb(w_G1gat_6[2]),.dout(n75),.clk(gclk));
	jnot g0012(.din(w_n75_0[1]),.dout(n76),.clk(gclk));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G290gat_7[0]),.dout(n78),.clk(gclk));
	jor g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79),.clk(gclk));
	jor g0016(.dina(n79),.dinb(w_n70_0[0]),.dout(n80),.clk(gclk));
	jand g0017(.dina(w_G273gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jor g0018(.dina(n81),.dinb(w_n65_0[0]),.dout(n82),.clk(gclk));
	jand g0019(.dina(w_dff_B_rhRcGDUD6_0),.dinb(w_n80_0[2]),.dout(n83),.clk(gclk));
	jxor g0020(.dina(w_n83_0[1]),.dinb(w_n67_0[0]),.dout(n84),.clk(gclk));
	jxor g0021(.dina(w_n84_0[1]),.dinb(w_dff_B_89v3w0f13_1),.dout(w_dff_A_aqNNkNcQ8_2),.clk(gclk));
	jand g0022(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n86),.clk(gclk));
	jnot g0023(.din(w_n86_0[1]),.dout(n87),.clk(gclk));
	jor g0024(.dina(w_n83_0[0]),.dinb(w_n66_0[0]),.dout(n88),.clk(gclk));
	jor g0025(.dina(w_n84_0[0]),.dinb(w_n75_0[0]),.dout(n89),.clk(gclk));
	jand g0026(.dina(n89),.dinb(w_dff_B_QQCVQAKW5_1),.dout(n90),.clk(gclk));
	jand g0027(.dina(w_G307gat_7[0]),.dinb(w_G18gat_6[2]),.dout(n91),.clk(gclk));
	jnot g0028(.din(w_n91_0[1]),.dout(n92),.clk(gclk));
	jnot g0029(.din(w_n80_0[1]),.dout(n93),.clk(gclk));
	jor g0030(.dina(w_n69_0[0]),.dinb(w_n77_0[0]),.dout(n94),.clk(gclk));
	jnot g0031(.din(w_G52gat_7[2]),.dout(n95),.clk(gclk));
	jor g0032(.dina(w_n78_0[0]),.dinb(n95),.dout(n96),.clk(gclk));
	jor g0033(.dina(n96),.dinb(n94),.dout(n97),.clk(gclk));
	jand g0034(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G273gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jor g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100),.clk(gclk));
	jand g0037(.dina(w_dff_B_pauhNMKf4_0),.dinb(w_n97_0[1]),.dout(n101),.clk(gclk));
	jxor g0038(.dina(w_n101_0[2]),.dinb(w_n93_0[1]),.dout(n102),.clk(gclk));
	jxor g0039(.dina(n102),.dinb(w_dff_B_x4Y6O9rC9_1),.dout(n103),.clk(gclk));
	jxor g0040(.dina(w_n103_0[1]),.dinb(w_n90_0[1]),.dout(n104),.clk(gclk));
	jxor g0041(.dina(w_n104_0[1]),.dinb(w_dff_B_yVHZgx371_1),.dout(w_dff_A_ia5znL6j8_2),.clk(gclk));
	jand g0042(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n106),.clk(gclk));
	jnot g0043(.din(w_n106_0[1]),.dout(n107),.clk(gclk));
	jnot g0044(.din(w_n103_0[0]),.dout(n108),.clk(gclk));
	jor g0045(.dina(n108),.dinb(w_n90_0[0]),.dout(n109),.clk(gclk));
	jor g0046(.dina(w_n104_0[0]),.dinb(w_n86_0[0]),.dout(n110),.clk(gclk));
	jand g0047(.dina(n110),.dinb(w_dff_B_LscLupag7_1),.dout(n111),.clk(gclk));
	jand g0048(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n112),.clk(gclk));
	jnot g0049(.din(w_n112_0[1]),.dout(n113),.clk(gclk));
	jor g0050(.dina(w_n101_0[1]),.dinb(w_n93_0[0]),.dout(n114),.clk(gclk));
	jxor g0051(.dina(w_n101_0[0]),.dinb(w_n80_0[0]),.dout(n115),.clk(gclk));
	jor g0052(.dina(n115),.dinb(w_n91_0[0]),.dout(n116),.clk(gclk));
	jand g0053(.dina(n116),.dinb(w_dff_B_aDyFGiMl4_1),.dout(n117),.clk(gclk));
	jand g0054(.dina(w_G307gat_6[2]),.dinb(w_G35gat_6[2]),.dout(n118),.clk(gclk));
	jnot g0055(.din(n118),.dout(n119),.clk(gclk));
	jnot g0056(.din(w_n97_0[0]),.dout(n120),.clk(gclk));
	jand g0057(.dina(w_G290gat_6[1]),.dinb(w_G69gat_7[1]),.dout(n121),.clk(gclk));
	jand g0058(.dina(w_n121_0[1]),.dinb(w_n99_0[0]),.dout(n122),.clk(gclk));
	jnot g0059(.din(w_n122_0[1]),.dout(n123),.clk(gclk));
	jand g0060(.dina(w_G290gat_6[0]),.dinb(w_G52gat_7[0]),.dout(n124),.clk(gclk));
	jand g0061(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n125),.clk(gclk));
	jor g0062(.dina(w_n125_0[1]),.dinb(n124),.dout(n126),.clk(gclk));
	jand g0063(.dina(w_dff_B_ULWUSYyN0_0),.dinb(w_n123_0[1]),.dout(n127),.clk(gclk));
	jxor g0064(.dina(w_n127_0[1]),.dinb(w_n120_0[1]),.dout(n128),.clk(gclk));
	jxor g0065(.dina(w_n128_0[1]),.dinb(w_n119_0[1]),.dout(n129),.clk(gclk));
	jnot g0066(.din(w_n129_0[1]),.dout(n130),.clk(gclk));
	jxor g0067(.dina(w_n130_0[1]),.dinb(w_n117_0[2]),.dout(n131),.clk(gclk));
	jxor g0068(.dina(n131),.dinb(w_dff_B_VfglReMp4_1),.dout(n132),.clk(gclk));
	jxor g0069(.dina(w_n132_0[1]),.dinb(w_n111_0[1]),.dout(n133),.clk(gclk));
	jxor g0070(.dina(w_n133_0[1]),.dinb(w_dff_B_UWWTPYVO4_1),.dout(w_dff_A_aLbf6XPK1_2),.clk(gclk));
	jand g0071(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n135),.clk(gclk));
	jnot g0072(.din(w_n135_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(w_n132_0[0]),.dout(n137),.clk(gclk));
	jor g0074(.dina(n137),.dinb(w_n111_0[0]),.dout(n138),.clk(gclk));
	jor g0075(.dina(w_n133_0[0]),.dinb(w_n106_0[0]),.dout(n139),.clk(gclk));
	jand g0076(.dina(n139),.dinb(w_dff_B_UhHJoqrF3_1),.dout(n140),.clk(gclk));
	jand g0077(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n141),.clk(gclk));
	jnot g0078(.din(w_n141_0[1]),.dout(n142),.clk(gclk));
	jor g0079(.dina(w_n130_0[0]),.dinb(w_n117_0[1]),.dout(n143),.clk(gclk));
	jxor g0080(.dina(w_n129_0[0]),.dinb(w_n117_0[0]),.dout(n144),.clk(gclk));
	jor g0081(.dina(n144),.dinb(w_n112_0[0]),.dout(n145),.clk(gclk));
	jand g0082(.dina(n145),.dinb(w_dff_B_rLkhshyZ4_1),.dout(n146),.clk(gclk));
	jand g0083(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n147),.clk(gclk));
	jnot g0084(.din(n147),.dout(n148),.clk(gclk));
	jor g0085(.dina(w_n127_0[0]),.dinb(w_n120_0[0]),.dout(n149),.clk(gclk));
	jnot g0086(.din(n149),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_n128_0[0]),.dinb(w_n119_0[0]),.dout(n151),.clk(gclk));
	jor g0088(.dina(n151),.dinb(n150),.dout(n152),.clk(gclk));
	jand g0089(.dina(w_G307gat_6[1]),.dinb(w_G52gat_6[2]),.dout(n153),.clk(gclk));
	jnot g0090(.din(n153),.dout(n154),.clk(gclk));
	jand g0091(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n155),.clk(gclk));
	jand g0092(.dina(w_n155_0[1]),.dinb(w_n125_0[0]),.dout(n156),.clk(gclk));
	jnot g0093(.din(w_n156_0[1]),.dout(n157),.clk(gclk));
	jand g0094(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n158),.clk(gclk));
	jor g0095(.dina(w_n158_0[1]),.dinb(w_n121_0[0]),.dout(n159),.clk(gclk));
	jand g0096(.dina(w_dff_B_fGZCObuk2_0),.dinb(w_n157_0[1]),.dout(n160),.clk(gclk));
	jxor g0097(.dina(w_n160_0[1]),.dinb(w_n122_0[0]),.dout(n161),.clk(gclk));
	jxor g0098(.dina(w_n161_0[1]),.dinb(w_n154_0[1]),.dout(n162),.clk(gclk));
	jxor g0099(.dina(w_n162_0[1]),.dinb(w_n152_0[1]),.dout(n163),.clk(gclk));
	jxor g0100(.dina(w_n163_0[1]),.dinb(w_n148_0[1]),.dout(n164),.clk(gclk));
	jnot g0101(.din(w_n164_0[1]),.dout(n165),.clk(gclk));
	jxor g0102(.dina(w_n165_0[1]),.dinb(w_n146_0[2]),.dout(n166),.clk(gclk));
	jxor g0103(.dina(n166),.dinb(w_dff_B_UaMuF6AQ2_1),.dout(n167),.clk(gclk));
	jxor g0104(.dina(w_n167_0[1]),.dinb(w_n140_0[1]),.dout(n168),.clk(gclk));
	jxor g0105(.dina(w_n168_0[1]),.dinb(w_dff_B_BnXbdPhm6_1),.dout(w_dff_A_vopQHw7W8_2),.clk(gclk));
	jand g0106(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n170),.clk(gclk));
	jnot g0107(.din(w_n170_0[1]),.dout(n171),.clk(gclk));
	jnot g0108(.din(w_n167_0[0]),.dout(n172),.clk(gclk));
	jor g0109(.dina(n172),.dinb(w_n140_0[0]),.dout(n173),.clk(gclk));
	jor g0110(.dina(w_n168_0[0]),.dinb(w_n135_0[0]),.dout(n174),.clk(gclk));
	jand g0111(.dina(n174),.dinb(w_dff_B_Sr0tDaY84_1),.dout(n175),.clk(gclk));
	jand g0112(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n176),.clk(gclk));
	jnot g0113(.din(w_n176_0[1]),.dout(n177),.clk(gclk));
	jor g0114(.dina(w_n165_0[0]),.dinb(w_n146_0[1]),.dout(n178),.clk(gclk));
	jxor g0115(.dina(w_n164_0[0]),.dinb(w_n146_0[0]),.dout(n179),.clk(gclk));
	jor g0116(.dina(n179),.dinb(w_n141_0[0]),.dout(n180),.clk(gclk));
	jand g0117(.dina(n180),.dinb(w_dff_B_P5uHvnYR7_1),.dout(n181),.clk(gclk));
	jand g0118(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n182),.clk(gclk));
	jnot g0119(.din(n182),.dout(n183),.clk(gclk));
	jand g0120(.dina(w_n162_0[0]),.dinb(w_n152_0[0]),.dout(n184),.clk(gclk));
	jand g0121(.dina(w_n163_0[0]),.dinb(w_n148_0[0]),.dout(n185),.clk(gclk));
	jor g0122(.dina(n185),.dinb(w_dff_B_Duh6237q9_1),.dout(n186),.clk(gclk));
	jand g0123(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n187),.clk(gclk));
	jnot g0124(.din(n187),.dout(n188),.clk(gclk));
	jnot g0125(.din(w_n160_0[0]),.dout(n189),.clk(gclk));
	jand g0126(.dina(n189),.dinb(w_n123_0[0]),.dout(n190),.clk(gclk));
	jand g0127(.dina(w_n161_0[0]),.dinb(w_n154_0[0]),.dout(n191),.clk(gclk));
	jor g0128(.dina(n191),.dinb(n190),.dout(n192),.clk(gclk));
	jand g0129(.dina(w_G307gat_6[0]),.dinb(w_G69gat_6[2]),.dout(n193),.clk(gclk));
	jnot g0130(.din(n193),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n195),.clk(gclk));
	jand g0132(.dina(w_n195_0[1]),.dinb(w_n158_0[0]),.dout(n196),.clk(gclk));
	jnot g0133(.din(w_n196_0[2]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n198),.clk(gclk));
	jor g0135(.dina(w_n198_0[1]),.dinb(w_n155_0[0]),.dout(n199),.clk(gclk));
	jand g0136(.dina(w_dff_B_2jpNeUUR3_0),.dinb(n197),.dout(n200),.clk(gclk));
	jxor g0137(.dina(w_n200_0[1]),.dinb(w_n156_0[0]),.dout(n201),.clk(gclk));
	jxor g0138(.dina(w_n201_0[1]),.dinb(w_n194_0[1]),.dout(n202),.clk(gclk));
	jxor g0139(.dina(w_n202_0[1]),.dinb(w_n192_0[1]),.dout(n203),.clk(gclk));
	jxor g0140(.dina(w_n203_0[1]),.dinb(w_n188_0[1]),.dout(n204),.clk(gclk));
	jxor g0141(.dina(w_n204_0[1]),.dinb(w_n186_0[1]),.dout(n205),.clk(gclk));
	jxor g0142(.dina(w_n205_0[1]),.dinb(w_n183_0[1]),.dout(n206),.clk(gclk));
	jnot g0143(.din(w_n206_0[1]),.dout(n207),.clk(gclk));
	jxor g0144(.dina(w_n207_0[1]),.dinb(w_n181_0[2]),.dout(n208),.clk(gclk));
	jxor g0145(.dina(n208),.dinb(w_dff_B_OMTgwC4u0_1),.dout(n209),.clk(gclk));
	jxor g0146(.dina(w_n209_0[1]),.dinb(w_n175_0[1]),.dout(n210),.clk(gclk));
	jxor g0147(.dina(w_n210_0[1]),.dinb(w_dff_B_DpFfkr0Y4_1),.dout(w_dff_A_xPsKA8QQ4_2),.clk(gclk));
	jand g0148(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n212),.clk(gclk));
	jnot g0149(.din(w_n212_0[1]),.dout(n213),.clk(gclk));
	jnot g0150(.din(w_n209_0[0]),.dout(n214),.clk(gclk));
	jor g0151(.dina(n214),.dinb(w_n175_0[0]),.dout(n215),.clk(gclk));
	jor g0152(.dina(w_n210_0[0]),.dinb(w_n170_0[0]),.dout(n216),.clk(gclk));
	jand g0153(.dina(n216),.dinb(w_dff_B_ARqMBHW71_1),.dout(n217),.clk(gclk));
	jand g0154(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n218),.clk(gclk));
	jnot g0155(.din(w_n218_0[1]),.dout(n219),.clk(gclk));
	jor g0156(.dina(w_n207_0[0]),.dinb(w_n181_0[1]),.dout(n220),.clk(gclk));
	jxor g0157(.dina(w_n206_0[0]),.dinb(w_n181_0[0]),.dout(n221),.clk(gclk));
	jor g0158(.dina(n221),.dinb(w_n176_0[0]),.dout(n222),.clk(gclk));
	jand g0159(.dina(n222),.dinb(w_dff_B_v4dJJxTg5_1),.dout(n223),.clk(gclk));
	jand g0160(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n224),.clk(gclk));
	jnot g0161(.din(n224),.dout(n225),.clk(gclk));
	jand g0162(.dina(w_n204_0[0]),.dinb(w_n186_0[0]),.dout(n226),.clk(gclk));
	jand g0163(.dina(w_n205_0[0]),.dinb(w_n183_0[0]),.dout(n227),.clk(gclk));
	jor g0164(.dina(n227),.dinb(w_dff_B_awINEBjq5_1),.dout(n228),.clk(gclk));
	jand g0165(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n229),.clk(gclk));
	jnot g0166(.din(n229),.dout(n230),.clk(gclk));
	jand g0167(.dina(w_n202_0[0]),.dinb(w_n192_0[0]),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_n203_0[0]),.dinb(w_n188_0[0]),.dout(n232),.clk(gclk));
	jor g0169(.dina(n232),.dinb(w_dff_B_Zm1aESKy2_1),.dout(n233),.clk(gclk));
	jand g0170(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n234),.clk(gclk));
	jnot g0171(.din(n234),.dout(n235),.clk(gclk));
	jnot g0172(.din(w_n200_0[0]),.dout(n236),.clk(gclk));
	jand g0173(.dina(n236),.dinb(w_n157_0[0]),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_n201_0[0]),.dinb(w_n194_0[0]),.dout(n238),.clk(gclk));
	jor g0175(.dina(n238),.dinb(n237),.dout(n239),.clk(gclk));
	jand g0176(.dina(w_G307gat_5[2]),.dinb(w_G86gat_6[2]),.dout(n240),.clk(gclk));
	jnot g0177(.din(n240),.dout(n241),.clk(gclk));
	jand g0178(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n242),.clk(gclk));
	jand g0179(.dina(w_n242_0[1]),.dinb(w_n198_0[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(w_n243_0[2]),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n245),.clk(gclk));
	jor g0182(.dina(w_n245_0[1]),.dinb(w_n195_0[0]),.dout(n246),.clk(gclk));
	jand g0183(.dina(w_dff_B_R06sGySs5_0),.dinb(n244),.dout(n247),.clk(gclk));
	jxor g0184(.dina(w_n247_0[1]),.dinb(w_n196_0[1]),.dout(n248),.clk(gclk));
	jxor g0185(.dina(w_n248_0[1]),.dinb(w_n241_0[1]),.dout(n249),.clk(gclk));
	jxor g0186(.dina(w_n249_0[1]),.dinb(w_n239_0[1]),.dout(n250),.clk(gclk));
	jxor g0187(.dina(w_n250_0[1]),.dinb(w_n235_0[1]),.dout(n251),.clk(gclk));
	jxor g0188(.dina(w_n251_0[1]),.dinb(w_n233_0[1]),.dout(n252),.clk(gclk));
	jxor g0189(.dina(w_n252_0[1]),.dinb(w_n230_0[1]),.dout(n253),.clk(gclk));
	jxor g0190(.dina(w_n253_0[1]),.dinb(w_n228_0[1]),.dout(n254),.clk(gclk));
	jxor g0191(.dina(w_n254_0[1]),.dinb(w_n225_0[1]),.dout(n255),.clk(gclk));
	jnot g0192(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jxor g0193(.dina(w_n256_0[1]),.dinb(w_n223_0[2]),.dout(n257),.clk(gclk));
	jxor g0194(.dina(n257),.dinb(w_dff_B_e1S54b0o3_1),.dout(n258),.clk(gclk));
	jxor g0195(.dina(w_n258_0[1]),.dinb(w_n217_0[1]),.dout(n259),.clk(gclk));
	jxor g0196(.dina(w_n259_0[1]),.dinb(w_dff_B_vJqVPxU03_1),.dout(w_dff_A_ByNtDrk64_2),.clk(gclk));
	jand g0197(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n261),.clk(gclk));
	jnot g0198(.din(w_n261_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(w_n258_0[0]),.dout(n263),.clk(gclk));
	jor g0200(.dina(n263),.dinb(w_n217_0[0]),.dout(n264),.clk(gclk));
	jor g0201(.dina(w_n259_0[0]),.dinb(w_n212_0[0]),.dout(n265),.clk(gclk));
	jand g0202(.dina(n265),.dinb(w_dff_B_cjBnXVB24_1),.dout(n266),.clk(gclk));
	jand g0203(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n267),.clk(gclk));
	jnot g0204(.din(w_n267_0[1]),.dout(n268),.clk(gclk));
	jor g0205(.dina(w_n256_0[0]),.dinb(w_n223_0[1]),.dout(n269),.clk(gclk));
	jxor g0206(.dina(w_n255_0[0]),.dinb(w_n223_0[0]),.dout(n270),.clk(gclk));
	jor g0207(.dina(n270),.dinb(w_n218_0[0]),.dout(n271),.clk(gclk));
	jand g0208(.dina(n271),.dinb(w_dff_B_6xod8Z1X3_1),.dout(n272),.clk(gclk));
	jand g0209(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n273),.clk(gclk));
	jnot g0210(.din(n273),.dout(n274),.clk(gclk));
	jand g0211(.dina(w_n253_0[0]),.dinb(w_n228_0[0]),.dout(n275),.clk(gclk));
	jand g0212(.dina(w_n254_0[0]),.dinb(w_n225_0[0]),.dout(n276),.clk(gclk));
	jor g0213(.dina(n276),.dinb(w_dff_B_4NcILaiO4_1),.dout(n277),.clk(gclk));
	jand g0214(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n278),.clk(gclk));
	jnot g0215(.din(n278),.dout(n279),.clk(gclk));
	jand g0216(.dina(w_n251_0[0]),.dinb(w_n233_0[0]),.dout(n280),.clk(gclk));
	jand g0217(.dina(w_n252_0[0]),.dinb(w_n230_0[0]),.dout(n281),.clk(gclk));
	jor g0218(.dina(n281),.dinb(w_dff_B_P2mKMjuP8_1),.dout(n282),.clk(gclk));
	jand g0219(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(n283),.dout(n284),.clk(gclk));
	jand g0221(.dina(w_n249_0[0]),.dinb(w_n239_0[0]),.dout(n285),.clk(gclk));
	jand g0222(.dina(w_n250_0[0]),.dinb(w_n235_0[0]),.dout(n286),.clk(gclk));
	jor g0223(.dina(n286),.dinb(w_dff_B_9qhXiizZ6_1),.dout(n287),.clk(gclk));
	jand g0224(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n288),.clk(gclk));
	jnot g0225(.din(n288),.dout(n289),.clk(gclk));
	jor g0226(.dina(w_n247_0[0]),.dinb(w_n196_0[0]),.dout(n290),.clk(gclk));
	jnot g0227(.din(n290),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n248_0[0]),.dinb(w_n241_0[0]),.dout(n292),.clk(gclk));
	jor g0229(.dina(n292),.dinb(n291),.dout(n293),.clk(gclk));
	jand g0230(.dina(w_G307gat_5[1]),.dinb(w_G103gat_6[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n296_0[1]),.dinb(w_n245_0[0]),.dout(n297),.clk(gclk));
	jnot g0234(.din(w_n297_0[2]),.dout(n298),.clk(gclk));
	jand g0235(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n299),.clk(gclk));
	jor g0236(.dina(w_n299_0[1]),.dinb(w_n242_0[0]),.dout(n300),.clk(gclk));
	jand g0237(.dina(w_dff_B_Nlus2vSY4_0),.dinb(n298),.dout(n301),.clk(gclk));
	jxor g0238(.dina(w_n301_0[1]),.dinb(w_n243_0[1]),.dout(n302),.clk(gclk));
	jxor g0239(.dina(w_n302_0[1]),.dinb(w_n295_0[1]),.dout(n303),.clk(gclk));
	jxor g0240(.dina(w_n303_0[1]),.dinb(w_n293_0[1]),.dout(n304),.clk(gclk));
	jxor g0241(.dina(w_n304_0[1]),.dinb(w_n289_0[1]),.dout(n305),.clk(gclk));
	jxor g0242(.dina(w_n305_0[1]),.dinb(w_n287_0[1]),.dout(n306),.clk(gclk));
	jxor g0243(.dina(w_n306_0[1]),.dinb(w_n284_0[1]),.dout(n307),.clk(gclk));
	jxor g0244(.dina(w_n307_0[1]),.dinb(w_n282_0[1]),.dout(n308),.clk(gclk));
	jxor g0245(.dina(w_n308_0[1]),.dinb(w_n279_0[1]),.dout(n309),.clk(gclk));
	jxor g0246(.dina(w_n309_0[1]),.dinb(w_n277_0[1]),.dout(n310),.clk(gclk));
	jxor g0247(.dina(w_n310_0[1]),.dinb(w_n274_0[1]),.dout(n311),.clk(gclk));
	jnot g0248(.din(w_n311_0[1]),.dout(n312),.clk(gclk));
	jxor g0249(.dina(w_n312_0[1]),.dinb(w_n272_0[2]),.dout(n313),.clk(gclk));
	jxor g0250(.dina(n313),.dinb(w_dff_B_mPvqQbQg9_1),.dout(n314),.clk(gclk));
	jxor g0251(.dina(w_n314_0[1]),.dinb(w_n266_0[1]),.dout(n315),.clk(gclk));
	jxor g0252(.dina(w_n315_0[1]),.dinb(w_dff_B_r3WimfWD0_1),.dout(w_dff_A_nMXYqaCW1_2),.clk(gclk));
	jand g0253(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n317),.clk(gclk));
	jnot g0254(.din(w_n317_0[1]),.dout(n318),.clk(gclk));
	jnot g0255(.din(w_n314_0[0]),.dout(n319),.clk(gclk));
	jor g0256(.dina(n319),.dinb(w_n266_0[0]),.dout(n320),.clk(gclk));
	jor g0257(.dina(w_n315_0[0]),.dinb(w_n261_0[0]),.dout(n321),.clk(gclk));
	jand g0258(.dina(n321),.dinb(w_dff_B_3wO4YlSX2_1),.dout(n322),.clk(gclk));
	jand g0259(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n323),.clk(gclk));
	jnot g0260(.din(w_n323_0[1]),.dout(n324),.clk(gclk));
	jor g0261(.dina(w_n312_0[0]),.dinb(w_n272_0[1]),.dout(n325),.clk(gclk));
	jxor g0262(.dina(w_n311_0[0]),.dinb(w_n272_0[0]),.dout(n326),.clk(gclk));
	jor g0263(.dina(n326),.dinb(w_n267_0[0]),.dout(n327),.clk(gclk));
	jand g0264(.dina(n327),.dinb(w_dff_B_s7OczH1C1_1),.dout(n328),.clk(gclk));
	jand g0265(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n329),.clk(gclk));
	jnot g0266(.din(n329),.dout(n330),.clk(gclk));
	jand g0267(.dina(w_n309_0[0]),.dinb(w_n277_0[0]),.dout(n331),.clk(gclk));
	jand g0268(.dina(w_n310_0[0]),.dinb(w_n274_0[0]),.dout(n332),.clk(gclk));
	jor g0269(.dina(n332),.dinb(w_dff_B_01uMWL296_1),.dout(n333),.clk(gclk));
	jand g0270(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n334),.clk(gclk));
	jnot g0271(.din(n334),.dout(n335),.clk(gclk));
	jand g0272(.dina(w_n307_0[0]),.dinb(w_n282_0[0]),.dout(n336),.clk(gclk));
	jand g0273(.dina(w_n308_0[0]),.dinb(w_n279_0[0]),.dout(n337),.clk(gclk));
	jor g0274(.dina(n337),.dinb(w_dff_B_1rtVAh7u6_1),.dout(n338),.clk(gclk));
	jand g0275(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n339),.clk(gclk));
	jnot g0276(.din(n339),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_n305_0[0]),.dinb(w_n287_0[0]),.dout(n341),.clk(gclk));
	jand g0278(.dina(w_n306_0[0]),.dinb(w_n284_0[0]),.dout(n342),.clk(gclk));
	jor g0279(.dina(n342),.dinb(w_dff_B_P4zG5qW56_1),.dout(n343),.clk(gclk));
	jand g0280(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n344),.clk(gclk));
	jnot g0281(.din(n344),.dout(n345),.clk(gclk));
	jand g0282(.dina(w_n303_0[0]),.dinb(w_n293_0[0]),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_n304_0[0]),.dinb(w_n289_0[0]),.dout(n347),.clk(gclk));
	jor g0284(.dina(n347),.dinb(w_dff_B_d4C0Djht4_1),.dout(n348),.clk(gclk));
	jand g0285(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n349),.clk(gclk));
	jnot g0286(.din(n349),.dout(n350),.clk(gclk));
	jor g0287(.dina(w_n301_0[0]),.dinb(w_n243_0[0]),.dout(n351),.clk(gclk));
	jnot g0288(.din(n351),.dout(n352),.clk(gclk));
	jand g0289(.dina(w_n302_0[0]),.dinb(w_n295_0[0]),.dout(n353),.clk(gclk));
	jor g0290(.dina(n353),.dinb(n352),.dout(n354),.clk(gclk));
	jand g0291(.dina(w_G307gat_5[0]),.dinb(w_G120gat_6[2]),.dout(n355),.clk(gclk));
	jnot g0292(.din(n355),.dout(n356),.clk(gclk));
	jand g0293(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n357),.clk(gclk));
	jand g0294(.dina(w_n357_0[1]),.dinb(w_n299_0[0]),.dout(n358),.clk(gclk));
	jnot g0295(.din(w_n358_0[2]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n360),.clk(gclk));
	jor g0297(.dina(w_n360_0[1]),.dinb(w_n296_0[0]),.dout(n361),.clk(gclk));
	jand g0298(.dina(w_dff_B_PJsyqXJB2_0),.dinb(n359),.dout(n362),.clk(gclk));
	jxor g0299(.dina(w_n362_0[1]),.dinb(w_n297_0[1]),.dout(n363),.clk(gclk));
	jxor g0300(.dina(w_n363_0[1]),.dinb(w_n356_0[1]),.dout(n364),.clk(gclk));
	jxor g0301(.dina(w_n364_0[1]),.dinb(w_n354_0[1]),.dout(n365),.clk(gclk));
	jxor g0302(.dina(w_n365_0[1]),.dinb(w_n350_0[1]),.dout(n366),.clk(gclk));
	jxor g0303(.dina(w_n366_0[1]),.dinb(w_n348_0[1]),.dout(n367),.clk(gclk));
	jxor g0304(.dina(w_n367_0[1]),.dinb(w_n345_0[1]),.dout(n368),.clk(gclk));
	jxor g0305(.dina(w_n368_0[1]),.dinb(w_n343_0[1]),.dout(n369),.clk(gclk));
	jxor g0306(.dina(w_n369_0[1]),.dinb(w_n340_0[1]),.dout(n370),.clk(gclk));
	jxor g0307(.dina(w_n370_0[1]),.dinb(w_n338_0[1]),.dout(n371),.clk(gclk));
	jxor g0308(.dina(w_n371_0[1]),.dinb(w_n335_0[1]),.dout(n372),.clk(gclk));
	jxor g0309(.dina(w_n372_0[1]),.dinb(w_n333_0[1]),.dout(n373),.clk(gclk));
	jxor g0310(.dina(w_n373_0[1]),.dinb(w_n330_0[1]),.dout(n374),.clk(gclk));
	jnot g0311(.din(w_n374_0[1]),.dout(n375),.clk(gclk));
	jxor g0312(.dina(w_n375_0[1]),.dinb(w_n328_0[2]),.dout(n376),.clk(gclk));
	jxor g0313(.dina(n376),.dinb(w_dff_B_tbVrxYkZ0_1),.dout(n377),.clk(gclk));
	jxor g0314(.dina(w_n377_0[1]),.dinb(w_n322_0[1]),.dout(n378),.clk(gclk));
	jxor g0315(.dina(w_n378_0[1]),.dinb(w_dff_B_d7eeEngJ3_1),.dout(w_dff_A_jS7LkhAz1_2),.clk(gclk));
	jand g0316(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n380),.clk(gclk));
	jnot g0317(.din(w_n380_0[1]),.dout(n381),.clk(gclk));
	jnot g0318(.din(w_n377_0[0]),.dout(n382),.clk(gclk));
	jor g0319(.dina(n382),.dinb(w_n322_0[0]),.dout(n383),.clk(gclk));
	jor g0320(.dina(w_n378_0[0]),.dinb(w_n317_0[0]),.dout(n384),.clk(gclk));
	jand g0321(.dina(n384),.dinb(w_dff_B_ZpA9JmNq8_1),.dout(n385),.clk(gclk));
	jand g0322(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n386),.clk(gclk));
	jnot g0323(.din(w_n386_0[1]),.dout(n387),.clk(gclk));
	jor g0324(.dina(w_n375_0[0]),.dinb(w_n328_0[1]),.dout(n388),.clk(gclk));
	jxor g0325(.dina(w_n374_0[0]),.dinb(w_n328_0[0]),.dout(n389),.clk(gclk));
	jor g0326(.dina(n389),.dinb(w_n323_0[0]),.dout(n390),.clk(gclk));
	jand g0327(.dina(n390),.dinb(w_dff_B_jnPhVbWa4_1),.dout(n391),.clk(gclk));
	jand g0328(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n392),.clk(gclk));
	jnot g0329(.din(n392),.dout(n393),.clk(gclk));
	jand g0330(.dina(w_n372_0[0]),.dinb(w_n333_0[0]),.dout(n394),.clk(gclk));
	jand g0331(.dina(w_n373_0[0]),.dinb(w_n330_0[0]),.dout(n395),.clk(gclk));
	jor g0332(.dina(n395),.dinb(w_dff_B_elABO3cg9_1),.dout(n396),.clk(gclk));
	jand g0333(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n397),.clk(gclk));
	jnot g0334(.din(n397),.dout(n398),.clk(gclk));
	jand g0335(.dina(w_n370_0[0]),.dinb(w_n338_0[0]),.dout(n399),.clk(gclk));
	jand g0336(.dina(w_n371_0[0]),.dinb(w_n335_0[0]),.dout(n400),.clk(gclk));
	jor g0337(.dina(n400),.dinb(w_dff_B_0rCHEG0m8_1),.dout(n401),.clk(gclk));
	jand g0338(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n402),.clk(gclk));
	jnot g0339(.din(n402),.dout(n403),.clk(gclk));
	jand g0340(.dina(w_n368_0[0]),.dinb(w_n343_0[0]),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_n369_0[0]),.dinb(w_n340_0[0]),.dout(n405),.clk(gclk));
	jor g0342(.dina(n405),.dinb(w_dff_B_V1BaO2AM1_1),.dout(n406),.clk(gclk));
	jand g0343(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n407),.clk(gclk));
	jnot g0344(.din(n407),.dout(n408),.clk(gclk));
	jand g0345(.dina(w_n366_0[0]),.dinb(w_n348_0[0]),.dout(n409),.clk(gclk));
	jand g0346(.dina(w_n367_0[0]),.dinb(w_n345_0[0]),.dout(n410),.clk(gclk));
	jor g0347(.dina(n410),.dinb(w_dff_B_MeQzjXfG9_1),.dout(n411),.clk(gclk));
	jand g0348(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n412),.clk(gclk));
	jnot g0349(.din(n412),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n364_0[0]),.dinb(w_n354_0[0]),.dout(n414),.clk(gclk));
	jand g0351(.dina(w_n365_0[0]),.dinb(w_n350_0[0]),.dout(n415),.clk(gclk));
	jor g0352(.dina(n415),.dinb(w_dff_B_HLZqCbhz3_1),.dout(n416),.clk(gclk));
	jand g0353(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n417),.clk(gclk));
	jnot g0354(.din(n417),.dout(n418),.clk(gclk));
	jor g0355(.dina(w_n362_0[0]),.dinb(w_n297_0[0]),.dout(n419),.clk(gclk));
	jand g0356(.dina(w_n363_0[0]),.dinb(w_n356_0[0]),.dout(n420),.clk(gclk));
	jnot g0357(.din(n420),.dout(n421),.clk(gclk));
	jand g0358(.dina(n421),.dinb(w_dff_B_7jFsosD90_1),.dout(n422),.clk(gclk));
	jnot g0359(.din(n422),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_G307gat_4[2]),.dinb(w_G137gat_6[2]),.dout(n424),.clk(gclk));
	jnot g0361(.din(n424),.dout(n425),.clk(gclk));
	jand g0362(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n426),.clk(gclk));
	jand g0363(.dina(w_n426_0[1]),.dinb(w_n360_0[0]),.dout(n427),.clk(gclk));
	jnot g0364(.din(w_n427_0[2]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n429),.clk(gclk));
	jor g0366(.dina(w_n429_0[1]),.dinb(w_n357_0[0]),.dout(n430),.clk(gclk));
	jand g0367(.dina(w_dff_B_CBpFB20e9_0),.dinb(n428),.dout(n431),.clk(gclk));
	jxor g0368(.dina(w_n431_0[1]),.dinb(w_n358_0[1]),.dout(n432),.clk(gclk));
	jxor g0369(.dina(w_n432_0[1]),.dinb(w_n425_0[1]),.dout(n433),.clk(gclk));
	jxor g0370(.dina(w_n433_0[1]),.dinb(w_n423_0[1]),.dout(n434),.clk(gclk));
	jxor g0371(.dina(w_n434_0[1]),.dinb(w_n418_0[1]),.dout(n435),.clk(gclk));
	jxor g0372(.dina(w_n435_0[1]),.dinb(w_n416_0[1]),.dout(n436),.clk(gclk));
	jxor g0373(.dina(w_n436_0[1]),.dinb(w_n413_0[1]),.dout(n437),.clk(gclk));
	jxor g0374(.dina(w_n437_0[1]),.dinb(w_n411_0[1]),.dout(n438),.clk(gclk));
	jxor g0375(.dina(w_n438_0[1]),.dinb(w_n408_0[1]),.dout(n439),.clk(gclk));
	jxor g0376(.dina(w_n439_0[1]),.dinb(w_n406_0[1]),.dout(n440),.clk(gclk));
	jxor g0377(.dina(w_n440_0[1]),.dinb(w_n403_0[1]),.dout(n441),.clk(gclk));
	jxor g0378(.dina(w_n441_0[1]),.dinb(w_n401_0[1]),.dout(n442),.clk(gclk));
	jxor g0379(.dina(w_n442_0[1]),.dinb(w_n398_0[1]),.dout(n443),.clk(gclk));
	jxor g0380(.dina(w_n443_0[1]),.dinb(w_n396_0[1]),.dout(n444),.clk(gclk));
	jxor g0381(.dina(w_n444_0[1]),.dinb(w_n393_0[1]),.dout(n445),.clk(gclk));
	jnot g0382(.din(w_n445_0[1]),.dout(n446),.clk(gclk));
	jxor g0383(.dina(w_n446_0[1]),.dinb(w_n391_0[2]),.dout(n447),.clk(gclk));
	jxor g0384(.dina(n447),.dinb(w_dff_B_qslerWkk7_1),.dout(n448),.clk(gclk));
	jxor g0385(.dina(w_n448_0[1]),.dinb(w_n385_0[1]),.dout(n449),.clk(gclk));
	jxor g0386(.dina(w_n449_0[1]),.dinb(w_dff_B_ZlVotAqf9_1),.dout(w_dff_A_jXnwwKqc6_2),.clk(gclk));
	jand g0387(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n451),.clk(gclk));
	jnot g0388(.din(w_n451_0[1]),.dout(n452),.clk(gclk));
	jnot g0389(.din(w_n448_0[0]),.dout(n453),.clk(gclk));
	jor g0390(.dina(n453),.dinb(w_n385_0[0]),.dout(n454),.clk(gclk));
	jor g0391(.dina(w_n449_0[0]),.dinb(w_n380_0[0]),.dout(n455),.clk(gclk));
	jand g0392(.dina(n455),.dinb(w_dff_B_yG4BhU3r1_1),.dout(n456),.clk(gclk));
	jand g0393(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n457),.clk(gclk));
	jnot g0394(.din(w_n457_0[1]),.dout(n458),.clk(gclk));
	jor g0395(.dina(w_n446_0[0]),.dinb(w_n391_0[1]),.dout(n459),.clk(gclk));
	jxor g0396(.dina(w_n445_0[0]),.dinb(w_n391_0[0]),.dout(n460),.clk(gclk));
	jor g0397(.dina(n460),.dinb(w_n386_0[0]),.dout(n461),.clk(gclk));
	jand g0398(.dina(n461),.dinb(w_dff_B_qGdEvmpm9_1),.dout(n462),.clk(gclk));
	jand g0399(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n463),.clk(gclk));
	jnot g0400(.din(n463),.dout(n464),.clk(gclk));
	jand g0401(.dina(w_n443_0[0]),.dinb(w_n396_0[0]),.dout(n465),.clk(gclk));
	jand g0402(.dina(w_n444_0[0]),.dinb(w_n393_0[0]),.dout(n466),.clk(gclk));
	jor g0403(.dina(n466),.dinb(w_dff_B_gOSBDxmP5_1),.dout(n467),.clk(gclk));
	jand g0404(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n468),.clk(gclk));
	jnot g0405(.din(n468),.dout(n469),.clk(gclk));
	jand g0406(.dina(w_n441_0[0]),.dinb(w_n401_0[0]),.dout(n470),.clk(gclk));
	jand g0407(.dina(w_n442_0[0]),.dinb(w_n398_0[0]),.dout(n471),.clk(gclk));
	jor g0408(.dina(n471),.dinb(w_dff_B_mVu63OJQ1_1),.dout(n472),.clk(gclk));
	jand g0409(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n473),.clk(gclk));
	jnot g0410(.din(n473),.dout(n474),.clk(gclk));
	jand g0411(.dina(w_n439_0[0]),.dinb(w_n406_0[0]),.dout(n475),.clk(gclk));
	jand g0412(.dina(w_n440_0[0]),.dinb(w_n403_0[0]),.dout(n476),.clk(gclk));
	jor g0413(.dina(n476),.dinb(w_dff_B_wgPc0zdc6_1),.dout(n477),.clk(gclk));
	jand g0414(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n478),.clk(gclk));
	jnot g0415(.din(n478),.dout(n479),.clk(gclk));
	jand g0416(.dina(w_n437_0[0]),.dinb(w_n411_0[0]),.dout(n480),.clk(gclk));
	jand g0417(.dina(w_n438_0[0]),.dinb(w_n408_0[0]),.dout(n481),.clk(gclk));
	jor g0418(.dina(n481),.dinb(w_dff_B_HyF84s1z6_1),.dout(n482),.clk(gclk));
	jand g0419(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n435_0[0]),.dinb(w_n416_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n436_0[0]),.dinb(w_n413_0[0]),.dout(n486),.clk(gclk));
	jor g0423(.dina(n486),.dinb(w_dff_B_vOu5VeOi2_1),.dout(n487),.clk(gclk));
	jand g0424(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n433_0[0]),.dinb(w_n423_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n434_0[0]),.dinb(w_n418_0[0]),.dout(n491),.clk(gclk));
	jor g0428(.dina(n491),.dinb(w_dff_B_4uHK7tHT0_1),.dout(n492),.clk(gclk));
	jand g0429(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jor g0431(.dina(w_n431_0[0]),.dinb(w_n358_0[0]),.dout(n495),.clk(gclk));
	jand g0432(.dina(w_n432_0[0]),.dinb(w_n425_0[0]),.dout(n496),.clk(gclk));
	jnot g0433(.din(n496),.dout(n497),.clk(gclk));
	jand g0434(.dina(n497),.dinb(w_dff_B_9kJ7FV726_1),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_G307gat_4[1]),.dinb(w_G154gat_6[2]),.dout(n500),.clk(gclk));
	jnot g0437(.din(n500),.dout(n501),.clk(gclk));
	jand g0438(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n502),.clk(gclk));
	jand g0439(.dina(w_n502_0[1]),.dinb(w_n429_0[0]),.dout(n503),.clk(gclk));
	jnot g0440(.din(w_n503_0[2]),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n505),.clk(gclk));
	jor g0442(.dina(w_n505_0[1]),.dinb(w_n426_0[0]),.dout(n506),.clk(gclk));
	jand g0443(.dina(w_dff_B_bGahM8op0_0),.dinb(n504),.dout(n507),.clk(gclk));
	jxor g0444(.dina(w_n507_0[1]),.dinb(w_n427_0[1]),.dout(n508),.clk(gclk));
	jxor g0445(.dina(w_n508_0[1]),.dinb(w_n501_0[1]),.dout(n509),.clk(gclk));
	jxor g0446(.dina(w_n509_0[1]),.dinb(w_n499_0[1]),.dout(n510),.clk(gclk));
	jxor g0447(.dina(w_n510_0[1]),.dinb(w_n494_0[1]),.dout(n511),.clk(gclk));
	jxor g0448(.dina(w_n511_0[1]),.dinb(w_n492_0[1]),.dout(n512),.clk(gclk));
	jxor g0449(.dina(w_n512_0[1]),.dinb(w_n489_0[1]),.dout(n513),.clk(gclk));
	jxor g0450(.dina(w_n513_0[1]),.dinb(w_n487_0[1]),.dout(n514),.clk(gclk));
	jxor g0451(.dina(w_n514_0[1]),.dinb(w_n484_0[1]),.dout(n515),.clk(gclk));
	jxor g0452(.dina(w_n515_0[1]),.dinb(w_n482_0[1]),.dout(n516),.clk(gclk));
	jxor g0453(.dina(w_n516_0[1]),.dinb(w_n479_0[1]),.dout(n517),.clk(gclk));
	jxor g0454(.dina(w_n517_0[1]),.dinb(w_n477_0[1]),.dout(n518),.clk(gclk));
	jxor g0455(.dina(w_n518_0[1]),.dinb(w_n474_0[1]),.dout(n519),.clk(gclk));
	jxor g0456(.dina(w_n519_0[1]),.dinb(w_n472_0[1]),.dout(n520),.clk(gclk));
	jxor g0457(.dina(w_n520_0[1]),.dinb(w_n469_0[1]),.dout(n521),.clk(gclk));
	jxor g0458(.dina(w_n521_0[1]),.dinb(w_n467_0[1]),.dout(n522),.clk(gclk));
	jxor g0459(.dina(w_n522_0[1]),.dinb(w_n464_0[1]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[1]),.dout(n524),.clk(gclk));
	jxor g0461(.dina(w_n524_0[1]),.dinb(w_n462_0[2]),.dout(n525),.clk(gclk));
	jxor g0462(.dina(n525),.dinb(w_dff_B_KH04q8iw5_1),.dout(n526),.clk(gclk));
	jxor g0463(.dina(w_n526_0[1]),.dinb(w_n456_0[1]),.dout(n527),.clk(gclk));
	jxor g0464(.dina(w_n527_0[1]),.dinb(w_dff_B_YFRm4K5W1_1),.dout(w_dff_A_InJoAco86_2),.clk(gclk));
	jand g0465(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n529),.clk(gclk));
	jnot g0466(.din(w_n529_0[1]),.dout(n530),.clk(gclk));
	jnot g0467(.din(w_n526_0[0]),.dout(n531),.clk(gclk));
	jor g0468(.dina(n531),.dinb(w_n456_0[0]),.dout(n532),.clk(gclk));
	jor g0469(.dina(w_n527_0[0]),.dinb(w_n451_0[0]),.dout(n533),.clk(gclk));
	jand g0470(.dina(n533),.dinb(w_dff_B_7wRTG4kK2_1),.dout(n534),.clk(gclk));
	jand g0471(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n535),.clk(gclk));
	jnot g0472(.din(w_n535_0[1]),.dout(n536),.clk(gclk));
	jor g0473(.dina(w_n524_0[0]),.dinb(w_n462_0[1]),.dout(n537),.clk(gclk));
	jxor g0474(.dina(w_n523_0[0]),.dinb(w_n462_0[0]),.dout(n538),.clk(gclk));
	jor g0475(.dina(n538),.dinb(w_n457_0[0]),.dout(n539),.clk(gclk));
	jand g0476(.dina(n539),.dinb(w_dff_B_NqzeNCcz1_1),.dout(n540),.clk(gclk));
	jand g0477(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n541),.clk(gclk));
	jnot g0478(.din(n541),.dout(n542),.clk(gclk));
	jand g0479(.dina(w_n521_0[0]),.dinb(w_n467_0[0]),.dout(n543),.clk(gclk));
	jand g0480(.dina(w_n522_0[0]),.dinb(w_n464_0[0]),.dout(n544),.clk(gclk));
	jor g0481(.dina(n544),.dinb(w_dff_B_KtEFl8uK2_1),.dout(n545),.clk(gclk));
	jand g0482(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n546),.clk(gclk));
	jnot g0483(.din(n546),.dout(n547),.clk(gclk));
	jand g0484(.dina(w_n519_0[0]),.dinb(w_n472_0[0]),.dout(n548),.clk(gclk));
	jand g0485(.dina(w_n520_0[0]),.dinb(w_n469_0[0]),.dout(n549),.clk(gclk));
	jor g0486(.dina(n549),.dinb(w_dff_B_uYM3roB00_1),.dout(n550),.clk(gclk));
	jand g0487(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n551),.clk(gclk));
	jnot g0488(.din(n551),.dout(n552),.clk(gclk));
	jand g0489(.dina(w_n517_0[0]),.dinb(w_n477_0[0]),.dout(n553),.clk(gclk));
	jand g0490(.dina(w_n518_0[0]),.dinb(w_n474_0[0]),.dout(n554),.clk(gclk));
	jor g0491(.dina(n554),.dinb(w_dff_B_bbmwRxcR6_1),.dout(n555),.clk(gclk));
	jand g0492(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n556),.clk(gclk));
	jnot g0493(.din(n556),.dout(n557),.clk(gclk));
	jand g0494(.dina(w_n515_0[0]),.dinb(w_n482_0[0]),.dout(n558),.clk(gclk));
	jand g0495(.dina(w_n516_0[0]),.dinb(w_n479_0[0]),.dout(n559),.clk(gclk));
	jor g0496(.dina(n559),.dinb(w_dff_B_b6JibRo52_1),.dout(n560),.clk(gclk));
	jand g0497(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n561),.clk(gclk));
	jnot g0498(.din(n561),.dout(n562),.clk(gclk));
	jand g0499(.dina(w_n513_0[0]),.dinb(w_n487_0[0]),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n514_0[0]),.dinb(w_n484_0[0]),.dout(n564),.clk(gclk));
	jor g0501(.dina(n564),.dinb(w_dff_B_Op82aIIH5_1),.dout(n565),.clk(gclk));
	jand g0502(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n566),.clk(gclk));
	jnot g0503(.din(n566),.dout(n567),.clk(gclk));
	jand g0504(.dina(w_n511_0[0]),.dinb(w_n492_0[0]),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n512_0[0]),.dinb(w_n489_0[0]),.dout(n569),.clk(gclk));
	jor g0506(.dina(n569),.dinb(w_dff_B_IdxXSTVP0_1),.dout(n570),.clk(gclk));
	jand g0507(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n571),.clk(gclk));
	jnot g0508(.din(n571),.dout(n572),.clk(gclk));
	jand g0509(.dina(w_n509_0[0]),.dinb(w_n499_0[0]),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n510_0[0]),.dinb(w_n494_0[0]),.dout(n574),.clk(gclk));
	jor g0511(.dina(n574),.dinb(w_dff_B_akOY61NU1_1),.dout(n575),.clk(gclk));
	jand g0512(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n576),.clk(gclk));
	jnot g0513(.din(n576),.dout(n577),.clk(gclk));
	jor g0514(.dina(w_n507_0[0]),.dinb(w_n427_0[0]),.dout(n578),.clk(gclk));
	jand g0515(.dina(w_n508_0[0]),.dinb(w_n501_0[0]),.dout(n579),.clk(gclk));
	jnot g0516(.din(n579),.dout(n580),.clk(gclk));
	jand g0517(.dina(n580),.dinb(w_dff_B_vue9wlNq3_1),.dout(n581),.clk(gclk));
	jnot g0518(.din(n581),.dout(n582),.clk(gclk));
	jand g0519(.dina(w_G307gat_4[0]),.dinb(w_G171gat_6[2]),.dout(n583),.clk(gclk));
	jnot g0520(.din(n583),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n585),.clk(gclk));
	jand g0522(.dina(w_n585_0[1]),.dinb(w_n505_0[0]),.dout(n586),.clk(gclk));
	jnot g0523(.din(w_n586_0[2]),.dout(n587),.clk(gclk));
	jand g0524(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n588),.clk(gclk));
	jor g0525(.dina(w_n588_0[1]),.dinb(w_n502_0[0]),.dout(n589),.clk(gclk));
	jand g0526(.dina(w_dff_B_wGRbh8jc5_0),.dinb(n587),.dout(n590),.clk(gclk));
	jxor g0527(.dina(w_n590_0[1]),.dinb(w_n503_0[1]),.dout(n591),.clk(gclk));
	jxor g0528(.dina(w_n591_0[1]),.dinb(w_n584_0[1]),.dout(n592),.clk(gclk));
	jxor g0529(.dina(w_n592_0[1]),.dinb(w_n582_0[1]),.dout(n593),.clk(gclk));
	jxor g0530(.dina(w_n593_0[1]),.dinb(w_n577_0[1]),.dout(n594),.clk(gclk));
	jxor g0531(.dina(w_n594_0[1]),.dinb(w_n575_0[1]),.dout(n595),.clk(gclk));
	jxor g0532(.dina(w_n595_0[1]),.dinb(w_n572_0[1]),.dout(n596),.clk(gclk));
	jxor g0533(.dina(w_n596_0[1]),.dinb(w_n570_0[1]),.dout(n597),.clk(gclk));
	jxor g0534(.dina(w_n597_0[1]),.dinb(w_n567_0[1]),.dout(n598),.clk(gclk));
	jxor g0535(.dina(w_n598_0[1]),.dinb(w_n565_0[1]),.dout(n599),.clk(gclk));
	jxor g0536(.dina(w_n599_0[1]),.dinb(w_n562_0[1]),.dout(n600),.clk(gclk));
	jxor g0537(.dina(w_n600_0[1]),.dinb(w_n560_0[1]),.dout(n601),.clk(gclk));
	jxor g0538(.dina(w_n601_0[1]),.dinb(w_n557_0[1]),.dout(n602),.clk(gclk));
	jxor g0539(.dina(w_n602_0[1]),.dinb(w_n555_0[1]),.dout(n603),.clk(gclk));
	jxor g0540(.dina(w_n603_0[1]),.dinb(w_n552_0[1]),.dout(n604),.clk(gclk));
	jxor g0541(.dina(w_n604_0[1]),.dinb(w_n550_0[1]),.dout(n605),.clk(gclk));
	jxor g0542(.dina(w_n605_0[1]),.dinb(w_n547_0[1]),.dout(n606),.clk(gclk));
	jxor g0543(.dina(w_n606_0[1]),.dinb(w_n545_0[1]),.dout(n607),.clk(gclk));
	jxor g0544(.dina(w_n607_0[1]),.dinb(w_n542_0[1]),.dout(n608),.clk(gclk));
	jnot g0545(.din(w_n608_0[1]),.dout(n609),.clk(gclk));
	jxor g0546(.dina(w_n609_0[1]),.dinb(w_n540_0[2]),.dout(n610),.clk(gclk));
	jxor g0547(.dina(n610),.dinb(w_dff_B_NRDofYYa6_1),.dout(n611),.clk(gclk));
	jxor g0548(.dina(w_n611_0[1]),.dinb(w_n534_0[1]),.dout(n612),.clk(gclk));
	jxor g0549(.dina(w_n612_0[1]),.dinb(w_dff_B_Hf4zsWZq2_1),.dout(w_dff_A_XOoOUeVN7_2),.clk(gclk));
	jand g0550(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n614),.clk(gclk));
	jnot g0551(.din(w_n614_0[1]),.dout(n615),.clk(gclk));
	jnot g0552(.din(w_n611_0[0]),.dout(n616),.clk(gclk));
	jor g0553(.dina(n616),.dinb(w_n534_0[0]),.dout(n617),.clk(gclk));
	jor g0554(.dina(w_n612_0[0]),.dinb(w_n529_0[0]),.dout(n618),.clk(gclk));
	jand g0555(.dina(n618),.dinb(w_dff_B_gDaYprKw4_1),.dout(n619),.clk(gclk));
	jand g0556(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n620),.clk(gclk));
	jnot g0557(.din(w_n620_0[1]),.dout(n621),.clk(gclk));
	jor g0558(.dina(w_n609_0[0]),.dinb(w_n540_0[1]),.dout(n622),.clk(gclk));
	jxor g0559(.dina(w_n608_0[0]),.dinb(w_n540_0[0]),.dout(n623),.clk(gclk));
	jor g0560(.dina(n623),.dinb(w_n535_0[0]),.dout(n624),.clk(gclk));
	jand g0561(.dina(n624),.dinb(w_dff_B_pjmkXbrx0_1),.dout(n625),.clk(gclk));
	jand g0562(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n626),.clk(gclk));
	jnot g0563(.din(n626),.dout(n627),.clk(gclk));
	jand g0564(.dina(w_n606_0[0]),.dinb(w_n545_0[0]),.dout(n628),.clk(gclk));
	jand g0565(.dina(w_n607_0[0]),.dinb(w_n542_0[0]),.dout(n629),.clk(gclk));
	jor g0566(.dina(n629),.dinb(w_dff_B_3fIFSjOP8_1),.dout(n630),.clk(gclk));
	jand g0567(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n631),.clk(gclk));
	jnot g0568(.din(n631),.dout(n632),.clk(gclk));
	jand g0569(.dina(w_n604_0[0]),.dinb(w_n550_0[0]),.dout(n633),.clk(gclk));
	jand g0570(.dina(w_n605_0[0]),.dinb(w_n547_0[0]),.dout(n634),.clk(gclk));
	jor g0571(.dina(n634),.dinb(w_dff_B_TNkzBPEQ1_1),.dout(n635),.clk(gclk));
	jand g0572(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n636),.clk(gclk));
	jnot g0573(.din(n636),.dout(n637),.clk(gclk));
	jand g0574(.dina(w_n602_0[0]),.dinb(w_n555_0[0]),.dout(n638),.clk(gclk));
	jand g0575(.dina(w_n603_0[0]),.dinb(w_n552_0[0]),.dout(n639),.clk(gclk));
	jor g0576(.dina(n639),.dinb(w_dff_B_01Q6TyWu5_1),.dout(n640),.clk(gclk));
	jand g0577(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n641),.clk(gclk));
	jnot g0578(.din(n641),.dout(n642),.clk(gclk));
	jand g0579(.dina(w_n600_0[0]),.dinb(w_n560_0[0]),.dout(n643),.clk(gclk));
	jand g0580(.dina(w_n601_0[0]),.dinb(w_n557_0[0]),.dout(n644),.clk(gclk));
	jor g0581(.dina(n644),.dinb(w_dff_B_SSFrj5Nk1_1),.dout(n645),.clk(gclk));
	jand g0582(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n646),.clk(gclk));
	jnot g0583(.din(n646),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_n598_0[0]),.dinb(w_n565_0[0]),.dout(n648),.clk(gclk));
	jand g0585(.dina(w_n599_0[0]),.dinb(w_n562_0[0]),.dout(n649),.clk(gclk));
	jor g0586(.dina(n649),.dinb(w_dff_B_bPimEsZa9_1),.dout(n650),.clk(gclk));
	jand g0587(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n651),.clk(gclk));
	jnot g0588(.din(n651),.dout(n652),.clk(gclk));
	jand g0589(.dina(w_n596_0[0]),.dinb(w_n570_0[0]),.dout(n653),.clk(gclk));
	jand g0590(.dina(w_n597_0[0]),.dinb(w_n567_0[0]),.dout(n654),.clk(gclk));
	jor g0591(.dina(n654),.dinb(w_dff_B_9p2hFyFV9_1),.dout(n655),.clk(gclk));
	jand g0592(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n656),.clk(gclk));
	jnot g0593(.din(n656),.dout(n657),.clk(gclk));
	jand g0594(.dina(w_n594_0[0]),.dinb(w_n575_0[0]),.dout(n658),.clk(gclk));
	jand g0595(.dina(w_n595_0[0]),.dinb(w_n572_0[0]),.dout(n659),.clk(gclk));
	jor g0596(.dina(n659),.dinb(w_dff_B_m2Jk00NH5_1),.dout(n660),.clk(gclk));
	jand g0597(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n661),.clk(gclk));
	jnot g0598(.din(n661),.dout(n662),.clk(gclk));
	jand g0599(.dina(w_n592_0[0]),.dinb(w_n582_0[0]),.dout(n663),.clk(gclk));
	jand g0600(.dina(w_n593_0[0]),.dinb(w_n577_0[0]),.dout(n664),.clk(gclk));
	jor g0601(.dina(n664),.dinb(w_dff_B_TtpsuMRV5_1),.dout(n665),.clk(gclk));
	jand g0602(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n666),.clk(gclk));
	jnot g0603(.din(n666),.dout(n667),.clk(gclk));
	jor g0604(.dina(w_n590_0[0]),.dinb(w_n503_0[0]),.dout(n668),.clk(gclk));
	jand g0605(.dina(w_n591_0[0]),.dinb(w_n584_0[0]),.dout(n669),.clk(gclk));
	jnot g0606(.din(n669),.dout(n670),.clk(gclk));
	jand g0607(.dina(n670),.dinb(w_dff_B_sNSkNFS63_1),.dout(n671),.clk(gclk));
	jnot g0608(.din(n671),.dout(n672),.clk(gclk));
	jand g0609(.dina(w_G307gat_3[2]),.dinb(w_G188gat_6[2]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n675_0[1]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jnot g0613(.din(w_n676_0[2]),.dout(n677),.clk(gclk));
	jand g0614(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n678),.clk(gclk));
	jor g0615(.dina(w_n678_0[1]),.dinb(w_n585_0[0]),.dout(n679),.clk(gclk));
	jand g0616(.dina(w_dff_B_2G8Dmrc76_0),.dinb(n677),.dout(n680),.clk(gclk));
	jxor g0617(.dina(w_n680_0[1]),.dinb(w_n586_0[1]),.dout(n681),.clk(gclk));
	jxor g0618(.dina(w_n681_0[1]),.dinb(w_n674_0[1]),.dout(n682),.clk(gclk));
	jxor g0619(.dina(w_n682_0[1]),.dinb(w_n672_0[1]),.dout(n683),.clk(gclk));
	jxor g0620(.dina(w_n683_0[1]),.dinb(w_n667_0[1]),.dout(n684),.clk(gclk));
	jxor g0621(.dina(w_n684_0[1]),.dinb(w_n665_0[1]),.dout(n685),.clk(gclk));
	jxor g0622(.dina(w_n685_0[1]),.dinb(w_n662_0[1]),.dout(n686),.clk(gclk));
	jxor g0623(.dina(w_n686_0[1]),.dinb(w_n660_0[1]),.dout(n687),.clk(gclk));
	jxor g0624(.dina(w_n687_0[1]),.dinb(w_n657_0[1]),.dout(n688),.clk(gclk));
	jxor g0625(.dina(w_n688_0[1]),.dinb(w_n655_0[1]),.dout(n689),.clk(gclk));
	jxor g0626(.dina(w_n689_0[1]),.dinb(w_n652_0[1]),.dout(n690),.clk(gclk));
	jxor g0627(.dina(w_n690_0[1]),.dinb(w_n650_0[1]),.dout(n691),.clk(gclk));
	jxor g0628(.dina(w_n691_0[1]),.dinb(w_n647_0[1]),.dout(n692),.clk(gclk));
	jxor g0629(.dina(w_n692_0[1]),.dinb(w_n645_0[1]),.dout(n693),.clk(gclk));
	jxor g0630(.dina(w_n693_0[1]),.dinb(w_n642_0[1]),.dout(n694),.clk(gclk));
	jxor g0631(.dina(w_n694_0[1]),.dinb(w_n640_0[1]),.dout(n695),.clk(gclk));
	jxor g0632(.dina(w_n695_0[1]),.dinb(w_n637_0[1]),.dout(n696),.clk(gclk));
	jxor g0633(.dina(w_n696_0[1]),.dinb(w_n635_0[1]),.dout(n697),.clk(gclk));
	jxor g0634(.dina(w_n697_0[1]),.dinb(w_n632_0[1]),.dout(n698),.clk(gclk));
	jxor g0635(.dina(w_n698_0[1]),.dinb(w_n630_0[1]),.dout(n699),.clk(gclk));
	jxor g0636(.dina(w_n699_0[1]),.dinb(w_n627_0[1]),.dout(n700),.clk(gclk));
	jnot g0637(.din(w_n700_0[1]),.dout(n701),.clk(gclk));
	jxor g0638(.dina(w_n701_0[1]),.dinb(w_n625_0[2]),.dout(n702),.clk(gclk));
	jxor g0639(.dina(n702),.dinb(w_dff_B_GvGucZMJ3_1),.dout(n703),.clk(gclk));
	jxor g0640(.dina(w_n703_0[1]),.dinb(w_n619_0[1]),.dout(n704),.clk(gclk));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_dff_B_OLxsTluA8_1),.dout(w_dff_A_2eploXL89_2),.clk(gclk));
	jand g0642(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n706),.clk(gclk));
	jnot g0643(.din(w_n706_0[1]),.dout(n707),.clk(gclk));
	jnot g0644(.din(w_n703_0[0]),.dout(n708),.clk(gclk));
	jor g0645(.dina(n708),.dinb(w_n619_0[0]),.dout(n709),.clk(gclk));
	jor g0646(.dina(w_n704_0[0]),.dinb(w_n614_0[0]),.dout(n710),.clk(gclk));
	jand g0647(.dina(n710),.dinb(w_dff_B_Xym03pKl7_1),.dout(n711),.clk(gclk));
	jand g0648(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n712),.clk(gclk));
	jnot g0649(.din(w_n712_0[1]),.dout(n713),.clk(gclk));
	jor g0650(.dina(w_n701_0[0]),.dinb(w_n625_0[1]),.dout(n714),.clk(gclk));
	jxor g0651(.dina(w_n700_0[0]),.dinb(w_n625_0[0]),.dout(n715),.clk(gclk));
	jor g0652(.dina(n715),.dinb(w_n620_0[0]),.dout(n716),.clk(gclk));
	jand g0653(.dina(n716),.dinb(w_dff_B_pflvUWRu2_1),.dout(n717),.clk(gclk));
	jand g0654(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n718),.clk(gclk));
	jnot g0655(.din(n718),.dout(n719),.clk(gclk));
	jand g0656(.dina(w_n698_0[0]),.dinb(w_n630_0[0]),.dout(n720),.clk(gclk));
	jand g0657(.dina(w_n699_0[0]),.dinb(w_n627_0[0]),.dout(n721),.clk(gclk));
	jor g0658(.dina(n721),.dinb(w_dff_B_qWDKSY1J5_1),.dout(n722),.clk(gclk));
	jand g0659(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n723),.clk(gclk));
	jnot g0660(.din(n723),.dout(n724),.clk(gclk));
	jand g0661(.dina(w_n696_0[0]),.dinb(w_n635_0[0]),.dout(n725),.clk(gclk));
	jand g0662(.dina(w_n697_0[0]),.dinb(w_n632_0[0]),.dout(n726),.clk(gclk));
	jor g0663(.dina(n726),.dinb(w_dff_B_K4OtTcjG8_1),.dout(n727),.clk(gclk));
	jand g0664(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n728),.clk(gclk));
	jnot g0665(.din(n728),.dout(n729),.clk(gclk));
	jand g0666(.dina(w_n694_0[0]),.dinb(w_n640_0[0]),.dout(n730),.clk(gclk));
	jand g0667(.dina(w_n695_0[0]),.dinb(w_n637_0[0]),.dout(n731),.clk(gclk));
	jor g0668(.dina(n731),.dinb(w_dff_B_mrmko7236_1),.dout(n732),.clk(gclk));
	jand g0669(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n733),.clk(gclk));
	jnot g0670(.din(n733),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_n692_0[0]),.dinb(w_n645_0[0]),.dout(n735),.clk(gclk));
	jand g0672(.dina(w_n693_0[0]),.dinb(w_n642_0[0]),.dout(n736),.clk(gclk));
	jor g0673(.dina(n736),.dinb(w_dff_B_a5hMvIXr4_1),.dout(n737),.clk(gclk));
	jand g0674(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n738),.clk(gclk));
	jnot g0675(.din(n738),.dout(n739),.clk(gclk));
	jand g0676(.dina(w_n690_0[0]),.dinb(w_n650_0[0]),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_n691_0[0]),.dinb(w_n647_0[0]),.dout(n741),.clk(gclk));
	jor g0678(.dina(n741),.dinb(w_dff_B_uh9KG59w7_1),.dout(n742),.clk(gclk));
	jand g0679(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n743),.clk(gclk));
	jnot g0680(.din(n743),.dout(n744),.clk(gclk));
	jand g0681(.dina(w_n688_0[0]),.dinb(w_n655_0[0]),.dout(n745),.clk(gclk));
	jand g0682(.dina(w_n689_0[0]),.dinb(w_n652_0[0]),.dout(n746),.clk(gclk));
	jor g0683(.dina(n746),.dinb(w_dff_B_SLuxqxfn3_1),.dout(n747),.clk(gclk));
	jand g0684(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n748),.clk(gclk));
	jnot g0685(.din(n748),.dout(n749),.clk(gclk));
	jand g0686(.dina(w_n686_0[0]),.dinb(w_n660_0[0]),.dout(n750),.clk(gclk));
	jand g0687(.dina(w_n687_0[0]),.dinb(w_n657_0[0]),.dout(n751),.clk(gclk));
	jor g0688(.dina(n751),.dinb(w_dff_B_r9B0w8l35_1),.dout(n752),.clk(gclk));
	jand g0689(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n753),.clk(gclk));
	jnot g0690(.din(n753),.dout(n754),.clk(gclk));
	jand g0691(.dina(w_n684_0[0]),.dinb(w_n665_0[0]),.dout(n755),.clk(gclk));
	jand g0692(.dina(w_n685_0[0]),.dinb(w_n662_0[0]),.dout(n756),.clk(gclk));
	jor g0693(.dina(n756),.dinb(w_dff_B_5jrER1x16_1),.dout(n757),.clk(gclk));
	jand g0694(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n758),.clk(gclk));
	jnot g0695(.din(n758),.dout(n759),.clk(gclk));
	jand g0696(.dina(w_n682_0[0]),.dinb(w_n672_0[0]),.dout(n760),.clk(gclk));
	jand g0697(.dina(w_n683_0[0]),.dinb(w_n667_0[0]),.dout(n761),.clk(gclk));
	jor g0698(.dina(n761),.dinb(w_dff_B_58V6RV5c9_1),.dout(n762),.clk(gclk));
	jand g0699(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n763),.clk(gclk));
	jnot g0700(.din(n763),.dout(n764),.clk(gclk));
	jor g0701(.dina(w_n680_0[0]),.dinb(w_n586_0[0]),.dout(n765),.clk(gclk));
	jand g0702(.dina(w_n681_0[0]),.dinb(w_n674_0[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(n767),.dinb(w_dff_B_ny94K4xr4_1),.dout(n768),.clk(gclk));
	jnot g0705(.din(n768),.dout(n769),.clk(gclk));
	jand g0706(.dina(w_G307gat_3[1]),.dinb(w_G205gat_6[2]),.dout(n770),.clk(gclk));
	jnot g0707(.din(n770),.dout(n771),.clk(gclk));
	jand g0708(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n772_0[1]),.dinb(w_n678_0[0]),.dout(n773),.clk(gclk));
	jnot g0710(.din(w_n773_0[1]),.dout(n774),.clk(gclk));
	jand g0711(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n775),.clk(gclk));
	jor g0712(.dina(w_n775_0[1]),.dinb(w_n675_0[0]),.dout(n776),.clk(gclk));
	jand g0713(.dina(w_dff_B_CPt8EioO4_0),.dinb(w_n774_0[1]),.dout(n777),.clk(gclk));
	jxor g0714(.dina(w_n777_0[1]),.dinb(w_n676_0[1]),.dout(n778),.clk(gclk));
	jxor g0715(.dina(w_n778_0[1]),.dinb(w_n771_0[1]),.dout(n779),.clk(gclk));
	jxor g0716(.dina(w_n779_0[1]),.dinb(w_n769_0[1]),.dout(n780),.clk(gclk));
	jxor g0717(.dina(w_n780_0[1]),.dinb(w_n764_0[1]),.dout(n781),.clk(gclk));
	jxor g0718(.dina(w_n781_0[1]),.dinb(w_n762_0[1]),.dout(n782),.clk(gclk));
	jxor g0719(.dina(w_n782_0[1]),.dinb(w_n759_0[1]),.dout(n783),.clk(gclk));
	jxor g0720(.dina(w_n783_0[1]),.dinb(w_n757_0[1]),.dout(n784),.clk(gclk));
	jxor g0721(.dina(w_n784_0[1]),.dinb(w_n754_0[1]),.dout(n785),.clk(gclk));
	jxor g0722(.dina(w_n785_0[1]),.dinb(w_n752_0[1]),.dout(n786),.clk(gclk));
	jxor g0723(.dina(w_n786_0[1]),.dinb(w_n749_0[1]),.dout(n787),.clk(gclk));
	jxor g0724(.dina(w_n787_0[1]),.dinb(w_n747_0[1]),.dout(n788),.clk(gclk));
	jxor g0725(.dina(w_n788_0[1]),.dinb(w_n744_0[1]),.dout(n789),.clk(gclk));
	jxor g0726(.dina(w_n789_0[1]),.dinb(w_n742_0[1]),.dout(n790),.clk(gclk));
	jxor g0727(.dina(w_n790_0[1]),.dinb(w_n739_0[1]),.dout(n791),.clk(gclk));
	jxor g0728(.dina(w_n791_0[1]),.dinb(w_n737_0[1]),.dout(n792),.clk(gclk));
	jxor g0729(.dina(w_n792_0[1]),.dinb(w_n734_0[1]),.dout(n793),.clk(gclk));
	jxor g0730(.dina(w_n793_0[1]),.dinb(w_n732_0[1]),.dout(n794),.clk(gclk));
	jxor g0731(.dina(w_n794_0[1]),.dinb(w_n729_0[1]),.dout(n795),.clk(gclk));
	jxor g0732(.dina(w_n795_0[1]),.dinb(w_n727_0[1]),.dout(n796),.clk(gclk));
	jxor g0733(.dina(w_n796_0[1]),.dinb(w_n724_0[1]),.dout(n797),.clk(gclk));
	jxor g0734(.dina(w_n797_0[1]),.dinb(w_n722_0[1]),.dout(n798),.clk(gclk));
	jxor g0735(.dina(w_n798_0[1]),.dinb(w_n719_0[1]),.dout(n799),.clk(gclk));
	jnot g0736(.din(w_n799_0[1]),.dout(n800),.clk(gclk));
	jxor g0737(.dina(w_n800_0[1]),.dinb(w_n717_0[2]),.dout(n801),.clk(gclk));
	jxor g0738(.dina(n801),.dinb(w_dff_B_6wcSrPEr9_1),.dout(n802),.clk(gclk));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n711_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_dff_B_aIJIHk8U5_1),.dout(w_dff_A_Y7aiHoy19_2),.clk(gclk));
	jand g0741(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n805),.clk(gclk));
	jnot g0742(.din(w_n805_0[1]),.dout(n806),.clk(gclk));
	jnot g0743(.din(w_n802_0[0]),.dout(n807),.clk(gclk));
	jor g0744(.dina(n807),.dinb(w_n711_0[0]),.dout(n808),.clk(gclk));
	jor g0745(.dina(w_n803_0[0]),.dinb(w_n706_0[0]),.dout(n809),.clk(gclk));
	jand g0746(.dina(n809),.dinb(w_dff_B_2rNmKVuM2_1),.dout(n810),.clk(gclk));
	jand g0747(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n811),.clk(gclk));
	jor g0748(.dina(w_n800_0[0]),.dinb(w_n717_0[1]),.dout(n812),.clk(gclk));
	jxor g0749(.dina(w_n799_0[0]),.dinb(w_n717_0[0]),.dout(n813),.clk(gclk));
	jor g0750(.dina(n813),.dinb(w_n712_0[0]),.dout(n814),.clk(gclk));
	jand g0751(.dina(n814),.dinb(w_dff_B_XlmD80Zn1_1),.dout(n815),.clk(gclk));
	jand g0752(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n816),.clk(gclk));
	jnot g0753(.din(w_n816_0[1]),.dout(n817),.clk(gclk));
	jand g0754(.dina(w_n797_0[0]),.dinb(w_n722_0[0]),.dout(n818),.clk(gclk));
	jand g0755(.dina(w_n798_0[0]),.dinb(w_n719_0[0]),.dout(n819),.clk(gclk));
	jor g0756(.dina(n819),.dinb(w_dff_B_tjlHIzTL2_1),.dout(n820),.clk(gclk));
	jand g0757(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n821),.clk(gclk));
	jnot g0758(.din(n821),.dout(n822),.clk(gclk));
	jand g0759(.dina(w_n795_0[0]),.dinb(w_n727_0[0]),.dout(n823),.clk(gclk));
	jand g0760(.dina(w_n796_0[0]),.dinb(w_n724_0[0]),.dout(n824),.clk(gclk));
	jor g0761(.dina(n824),.dinb(w_dff_B_9fVbZpba6_1),.dout(n825),.clk(gclk));
	jand g0762(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n826),.clk(gclk));
	jnot g0763(.din(n826),.dout(n827),.clk(gclk));
	jand g0764(.dina(w_n793_0[0]),.dinb(w_n732_0[0]),.dout(n828),.clk(gclk));
	jand g0765(.dina(w_n794_0[0]),.dinb(w_n729_0[0]),.dout(n829),.clk(gclk));
	jor g0766(.dina(n829),.dinb(w_dff_B_xSfesVRc9_1),.dout(n830),.clk(gclk));
	jand g0767(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n831),.clk(gclk));
	jnot g0768(.din(n831),.dout(n832),.clk(gclk));
	jand g0769(.dina(w_n791_0[0]),.dinb(w_n737_0[0]),.dout(n833),.clk(gclk));
	jand g0770(.dina(w_n792_0[0]),.dinb(w_n734_0[0]),.dout(n834),.clk(gclk));
	jor g0771(.dina(n834),.dinb(w_dff_B_b0QFyRaJ4_1),.dout(n835),.clk(gclk));
	jand g0772(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n836),.clk(gclk));
	jnot g0773(.din(n836),.dout(n837),.clk(gclk));
	jand g0774(.dina(w_n789_0[0]),.dinb(w_n742_0[0]),.dout(n838),.clk(gclk));
	jand g0775(.dina(w_n790_0[0]),.dinb(w_n739_0[0]),.dout(n839),.clk(gclk));
	jor g0776(.dina(n839),.dinb(w_dff_B_Ev4CQdpk0_1),.dout(n840),.clk(gclk));
	jand g0777(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n841),.clk(gclk));
	jnot g0778(.din(n841),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n787_0[0]),.dinb(w_n747_0[0]),.dout(n843),.clk(gclk));
	jand g0780(.dina(w_n788_0[0]),.dinb(w_n744_0[0]),.dout(n844),.clk(gclk));
	jor g0781(.dina(n844),.dinb(w_dff_B_rB1nKRZA0_1),.dout(n845),.clk(gclk));
	jand g0782(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n846),.clk(gclk));
	jnot g0783(.din(n846),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n785_0[0]),.dinb(w_n752_0[0]),.dout(n848),.clk(gclk));
	jand g0785(.dina(w_n786_0[0]),.dinb(w_n749_0[0]),.dout(n849),.clk(gclk));
	jor g0786(.dina(n849),.dinb(w_dff_B_2GiWZanX5_1),.dout(n850),.clk(gclk));
	jand g0787(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n851),.clk(gclk));
	jnot g0788(.din(n851),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n783_0[0]),.dinb(w_n757_0[0]),.dout(n853),.clk(gclk));
	jand g0790(.dina(w_n784_0[0]),.dinb(w_n754_0[0]),.dout(n854),.clk(gclk));
	jor g0791(.dina(n854),.dinb(w_dff_B_CqXK098R2_1),.dout(n855),.clk(gclk));
	jand g0792(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n856),.clk(gclk));
	jnot g0793(.din(n856),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n781_0[0]),.dinb(w_n762_0[0]),.dout(n858),.clk(gclk));
	jand g0795(.dina(w_n782_0[0]),.dinb(w_n759_0[0]),.dout(n859),.clk(gclk));
	jor g0796(.dina(n859),.dinb(w_dff_B_3kdNpIDS2_1),.dout(n860),.clk(gclk));
	jand g0797(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n861),.clk(gclk));
	jnot g0798(.din(n861),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n779_0[0]),.dinb(w_n769_0[0]),.dout(n863),.clk(gclk));
	jand g0800(.dina(w_n780_0[0]),.dinb(w_n764_0[0]),.dout(n864),.clk(gclk));
	jor g0801(.dina(n864),.dinb(w_dff_B_mHlV8etn5_1),.dout(n865),.clk(gclk));
	jand g0802(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n866),.clk(gclk));
	jnot g0803(.din(n866),.dout(n867),.clk(gclk));
	jor g0804(.dina(w_n777_0[0]),.dinb(w_n676_0[0]),.dout(n868),.clk(gclk));
	jand g0805(.dina(w_n778_0[0]),.dinb(w_n771_0[0]),.dout(n869),.clk(gclk));
	jnot g0806(.din(n869),.dout(n870),.clk(gclk));
	jand g0807(.dina(n870),.dinb(w_dff_B_B7jVbXwV8_1),.dout(n871),.clk(gclk));
	jnot g0808(.din(n871),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_G307gat_3[0]),.dinb(w_G222gat_6[2]),.dout(n873),.clk(gclk));
	jnot g0810(.din(n873),.dout(n874),.clk(gclk));
	jand g0811(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n875),.clk(gclk));
	jxor g0812(.dina(w_n875_0[1]),.dinb(w_n772_0[0]),.dout(n876),.clk(gclk));
	jor g0813(.dina(n876),.dinb(w_n773_0[0]),.dout(n877),.clk(gclk));
	jor g0814(.dina(w_n875_0[0]),.dinb(w_n774_0[0]),.dout(n878),.clk(gclk));
	jand g0815(.dina(n878),.dinb(w_n877_0[1]),.dout(n879),.clk(gclk));
	jxor g0816(.dina(w_n879_0[1]),.dinb(w_n874_0[1]),.dout(n880),.clk(gclk));
	jxor g0817(.dina(w_n880_0[1]),.dinb(w_n872_0[1]),.dout(n881),.clk(gclk));
	jxor g0818(.dina(w_n881_0[1]),.dinb(w_n867_0[1]),.dout(n882),.clk(gclk));
	jxor g0819(.dina(w_n882_0[1]),.dinb(w_n865_0[1]),.dout(n883),.clk(gclk));
	jxor g0820(.dina(w_n883_0[1]),.dinb(w_n862_0[1]),.dout(n884),.clk(gclk));
	jxor g0821(.dina(w_n884_0[1]),.dinb(w_n860_0[1]),.dout(n885),.clk(gclk));
	jxor g0822(.dina(w_n885_0[1]),.dinb(w_n857_0[1]),.dout(n886),.clk(gclk));
	jxor g0823(.dina(w_n886_0[1]),.dinb(w_n855_0[1]),.dout(n887),.clk(gclk));
	jxor g0824(.dina(w_n887_0[1]),.dinb(w_n852_0[1]),.dout(n888),.clk(gclk));
	jxor g0825(.dina(w_n888_0[1]),.dinb(w_n850_0[1]),.dout(n889),.clk(gclk));
	jxor g0826(.dina(w_n889_0[1]),.dinb(w_n847_0[1]),.dout(n890),.clk(gclk));
	jxor g0827(.dina(w_n890_0[1]),.dinb(w_n845_0[1]),.dout(n891),.clk(gclk));
	jxor g0828(.dina(w_n891_0[1]),.dinb(w_n842_0[1]),.dout(n892),.clk(gclk));
	jxor g0829(.dina(w_n892_0[1]),.dinb(w_n840_0[1]),.dout(n893),.clk(gclk));
	jxor g0830(.dina(w_n893_0[1]),.dinb(w_n837_0[1]),.dout(n894),.clk(gclk));
	jxor g0831(.dina(w_n894_0[1]),.dinb(w_n835_0[1]),.dout(n895),.clk(gclk));
	jxor g0832(.dina(w_n895_0[1]),.dinb(w_n832_0[1]),.dout(n896),.clk(gclk));
	jxor g0833(.dina(w_n896_0[1]),.dinb(w_n830_0[1]),.dout(n897),.clk(gclk));
	jxor g0834(.dina(w_n897_0[1]),.dinb(w_n827_0[1]),.dout(n898),.clk(gclk));
	jxor g0835(.dina(w_n898_0[1]),.dinb(w_n825_0[1]),.dout(n899),.clk(gclk));
	jxor g0836(.dina(w_n899_0[1]),.dinb(w_n822_0[1]),.dout(n900),.clk(gclk));
	jxor g0837(.dina(w_n900_0[2]),.dinb(w_n820_0[2]),.dout(n901),.clk(gclk));
	jxor g0838(.dina(n901),.dinb(w_dff_B_ANn0WTHP7_1),.dout(n902),.clk(gclk));
	jxor g0839(.dina(w_n902_0[1]),.dinb(w_n815_0[1]),.dout(n903),.clk(gclk));
	jxor g0840(.dina(w_n903_0[1]),.dinb(w_n811_0[1]),.dout(n904),.clk(gclk));
	jxor g0841(.dina(w_n904_0[1]),.dinb(w_n810_0[1]),.dout(n905),.clk(gclk));
	jxor g0842(.dina(w_n905_0[1]),.dinb(w_dff_B_8uvPJXgT8_1),.dout(w_dff_A_wIpjPOmp5_2),.clk(gclk));
	jnot g0843(.din(w_n904_0[0]),.dout(n907),.clk(gclk));
	jor g0844(.dina(n907),.dinb(w_n810_0[0]),.dout(n908),.clk(gclk));
	jor g0845(.dina(w_n905_0[0]),.dinb(w_n805_0[0]),.dout(n909),.clk(gclk));
	jand g0846(.dina(n909),.dinb(w_dff_B_ZO5Jnt0Y5_1),.dout(n910),.clk(gclk));
	jand g0847(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n911),.clk(gclk));
	jnot g0848(.din(w_n902_0[0]),.dout(n912),.clk(gclk));
	jor g0849(.dina(n912),.dinb(w_n815_0[0]),.dout(n913),.clk(gclk));
	jor g0850(.dina(w_n903_0[0]),.dinb(w_n811_0[0]),.dout(n914),.clk(gclk));
	jand g0851(.dina(n914),.dinb(w_dff_B_MBNG0AbL0_1),.dout(n915),.clk(gclk));
	jand g0852(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n916),.clk(gclk));
	jand g0853(.dina(w_n900_0[1]),.dinb(w_n820_0[1]),.dout(n917),.clk(gclk));
	jnot g0854(.din(n917),.dout(n918),.clk(gclk));
	jnot g0855(.din(w_n900_0[0]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(n919),.dinb(w_n820_0[0]),.dout(n920),.clk(gclk));
	jor g0857(.dina(n920),.dinb(w_n816_0[0]),.dout(n921),.clk(gclk));
	jand g0858(.dina(n921),.dinb(n918),.dout(n922),.clk(gclk));
	jand g0859(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n923),.clk(gclk));
	jnot g0860(.din(n923),.dout(n924),.clk(gclk));
	jand g0861(.dina(w_n898_0[0]),.dinb(w_n825_0[0]),.dout(n925),.clk(gclk));
	jand g0862(.dina(w_n899_0[0]),.dinb(w_n822_0[0]),.dout(n926),.clk(gclk));
	jor g0863(.dina(n926),.dinb(w_dff_B_S5HypYcJ0_1),.dout(n927),.clk(gclk));
	jand g0864(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n928),.clk(gclk));
	jnot g0865(.din(n928),.dout(n929),.clk(gclk));
	jand g0866(.dina(w_n896_0[0]),.dinb(w_n830_0[0]),.dout(n930),.clk(gclk));
	jand g0867(.dina(w_n897_0[0]),.dinb(w_n827_0[0]),.dout(n931),.clk(gclk));
	jor g0868(.dina(n931),.dinb(w_dff_B_E7UF84ec7_1),.dout(n932),.clk(gclk));
	jand g0869(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n933),.clk(gclk));
	jnot g0870(.din(n933),.dout(n934),.clk(gclk));
	jand g0871(.dina(w_n894_0[0]),.dinb(w_n835_0[0]),.dout(n935),.clk(gclk));
	jand g0872(.dina(w_n895_0[0]),.dinb(w_n832_0[0]),.dout(n936),.clk(gclk));
	jor g0873(.dina(n936),.dinb(w_dff_B_3xx9tJ5y5_1),.dout(n937),.clk(gclk));
	jand g0874(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n938),.clk(gclk));
	jnot g0875(.din(n938),.dout(n939),.clk(gclk));
	jand g0876(.dina(w_n892_0[0]),.dinb(w_n840_0[0]),.dout(n940),.clk(gclk));
	jand g0877(.dina(w_n893_0[0]),.dinb(w_n837_0[0]),.dout(n941),.clk(gclk));
	jor g0878(.dina(n941),.dinb(w_dff_B_oHrmig9b8_1),.dout(n942),.clk(gclk));
	jand g0879(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n943),.clk(gclk));
	jnot g0880(.din(n943),.dout(n944),.clk(gclk));
	jand g0881(.dina(w_n890_0[0]),.dinb(w_n845_0[0]),.dout(n945),.clk(gclk));
	jand g0882(.dina(w_n891_0[0]),.dinb(w_n842_0[0]),.dout(n946),.clk(gclk));
	jor g0883(.dina(n946),.dinb(w_dff_B_OnoqUXsn8_1),.dout(n947),.clk(gclk));
	jand g0884(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n948),.clk(gclk));
	jnot g0885(.din(n948),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_n888_0[0]),.dinb(w_n850_0[0]),.dout(n950),.clk(gclk));
	jand g0887(.dina(w_n889_0[0]),.dinb(w_n847_0[0]),.dout(n951),.clk(gclk));
	jor g0888(.dina(n951),.dinb(w_dff_B_SY1dVtdg4_1),.dout(n952),.clk(gclk));
	jand g0889(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n953),.clk(gclk));
	jnot g0890(.din(n953),.dout(n954),.clk(gclk));
	jand g0891(.dina(w_n886_0[0]),.dinb(w_n855_0[0]),.dout(n955),.clk(gclk));
	jand g0892(.dina(w_n887_0[0]),.dinb(w_n852_0[0]),.dout(n956),.clk(gclk));
	jor g0893(.dina(n956),.dinb(w_dff_B_TQIgVv3D2_1),.dout(n957),.clk(gclk));
	jand g0894(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n958),.clk(gclk));
	jnot g0895(.din(n958),.dout(n959),.clk(gclk));
	jand g0896(.dina(w_n884_0[0]),.dinb(w_n860_0[0]),.dout(n960),.clk(gclk));
	jand g0897(.dina(w_n885_0[0]),.dinb(w_n857_0[0]),.dout(n961),.clk(gclk));
	jor g0898(.dina(n961),.dinb(w_dff_B_RcaNpk1T7_1),.dout(n962),.clk(gclk));
	jand g0899(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n963),.clk(gclk));
	jnot g0900(.din(n963),.dout(n964),.clk(gclk));
	jand g0901(.dina(w_n882_0[0]),.dinb(w_n865_0[0]),.dout(n965),.clk(gclk));
	jand g0902(.dina(w_n883_0[0]),.dinb(w_n862_0[0]),.dout(n966),.clk(gclk));
	jor g0903(.dina(n966),.dinb(w_dff_B_AEG78ezj7_1),.dout(n967),.clk(gclk));
	jand g0904(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n968),.clk(gclk));
	jnot g0905(.din(n968),.dout(n969),.clk(gclk));
	jand g0906(.dina(w_n880_0[0]),.dinb(w_n872_0[0]),.dout(n970),.clk(gclk));
	jand g0907(.dina(w_n881_0[0]),.dinb(w_n867_0[0]),.dout(n971),.clk(gclk));
	jor g0908(.dina(n971),.dinb(w_dff_B_KaaAk79D5_1),.dout(n972),.clk(gclk));
	jand g0909(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n973),.clk(gclk));
	jnot g0910(.din(n973),.dout(n974),.clk(gclk));
	jand g0911(.dina(w_n879_0[0]),.dinb(w_n874_0[0]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(n976),.dinb(w_n877_0[0]),.dout(n977),.clk(gclk));
	jnot g0914(.din(n977),.dout(n978),.clk(gclk));
	jnot g0915(.din(w_n775_0[0]),.dout(n979),.clk(gclk));
	jand g0916(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n980),.clk(gclk));
	jand g0917(.dina(w_n980_0[1]),.dinb(n979),.dout(n981),.clk(gclk));
	jnot g0918(.din(n981),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_G307gat_2[2]),.dinb(w_G239gat_6[2]),.dout(n983),.clk(gclk));
	jxor g0920(.dina(w_n983_0[1]),.dinb(w_n982_0[1]),.dout(n984),.clk(gclk));
	jxor g0921(.dina(w_n984_0[1]),.dinb(w_n978_0[1]),.dout(n985),.clk(gclk));
	jxor g0922(.dina(w_n985_0[1]),.dinb(w_n974_0[1]),.dout(n986),.clk(gclk));
	jxor g0923(.dina(w_n986_0[1]),.dinb(w_n972_0[1]),.dout(n987),.clk(gclk));
	jxor g0924(.dina(w_n987_0[1]),.dinb(w_n969_0[1]),.dout(n988),.clk(gclk));
	jxor g0925(.dina(w_n988_0[1]),.dinb(w_n967_0[1]),.dout(n989),.clk(gclk));
	jxor g0926(.dina(w_n989_0[1]),.dinb(w_n964_0[1]),.dout(n990),.clk(gclk));
	jxor g0927(.dina(w_n990_0[1]),.dinb(w_n962_0[1]),.dout(n991),.clk(gclk));
	jxor g0928(.dina(w_n991_0[1]),.dinb(w_n959_0[1]),.dout(n992),.clk(gclk));
	jxor g0929(.dina(w_n992_0[1]),.dinb(w_n957_0[1]),.dout(n993),.clk(gclk));
	jxor g0930(.dina(w_n993_0[1]),.dinb(w_n954_0[1]),.dout(n994),.clk(gclk));
	jxor g0931(.dina(w_n994_0[1]),.dinb(w_n952_0[1]),.dout(n995),.clk(gclk));
	jxor g0932(.dina(w_n995_0[1]),.dinb(w_n949_0[1]),.dout(n996),.clk(gclk));
	jxor g0933(.dina(w_n996_0[1]),.dinb(w_n947_0[1]),.dout(n997),.clk(gclk));
	jxor g0934(.dina(w_n997_0[1]),.dinb(w_n944_0[1]),.dout(n998),.clk(gclk));
	jxor g0935(.dina(w_n998_0[1]),.dinb(w_n942_0[1]),.dout(n999),.clk(gclk));
	jxor g0936(.dina(w_n999_0[1]),.dinb(w_n939_0[1]),.dout(n1000),.clk(gclk));
	jxor g0937(.dina(w_n1000_0[1]),.dinb(w_n937_0[1]),.dout(n1001),.clk(gclk));
	jxor g0938(.dina(w_n1001_0[1]),.dinb(w_n934_0[1]),.dout(n1002),.clk(gclk));
	jxor g0939(.dina(w_n1002_0[1]),.dinb(w_n932_0[1]),.dout(n1003),.clk(gclk));
	jxor g0940(.dina(w_n1003_0[1]),.dinb(w_n929_0[1]),.dout(n1004),.clk(gclk));
	jxor g0941(.dina(w_n1004_0[1]),.dinb(w_n927_0[1]),.dout(n1005),.clk(gclk));
	jxor g0942(.dina(w_n1005_0[1]),.dinb(w_n924_0[1]),.dout(n1006),.clk(gclk));
	jxor g0943(.dina(w_n1006_0[1]),.dinb(w_n922_0[1]),.dout(n1007),.clk(gclk));
	jxor g0944(.dina(w_n1007_0[1]),.dinb(w_n916_0[1]),.dout(n1008),.clk(gclk));
	jnot g0945(.din(w_n1008_0[1]),.dout(n1009),.clk(gclk));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n915_0[2]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(n1010),.dinb(w_n911_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n910_0[1]),.dout(w_dff_A_UloyOVAB2_2),.clk(gclk));
	jand g0949(.dina(w_n1011_0[0]),.dinb(w_n910_0[0]),.dout(n1013),.clk(gclk));
	jor g0950(.dina(w_n1009_0[0]),.dinb(w_n915_0[1]),.dout(n1014),.clk(gclk));
	jxor g0951(.dina(w_n1008_0[0]),.dinb(w_n915_0[0]),.dout(n1015),.clk(gclk));
	jor g0952(.dina(n1015),.dinb(w_n911_0[0]),.dout(n1016),.clk(gclk));
	jand g0953(.dina(n1016),.dinb(w_dff_B_Hl1lC4wT5_1),.dout(n1017),.clk(gclk));
	jand g0954(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1018),.clk(gclk));
	jnot g0955(.din(w_n1006_0[0]),.dout(n1019),.clk(gclk));
	jor g0956(.dina(n1019),.dinb(w_n922_0[0]),.dout(n1020),.clk(gclk));
	jor g0957(.dina(w_n1007_0[0]),.dinb(w_n916_0[0]),.dout(n1021),.clk(gclk));
	jand g0958(.dina(n1021),.dinb(w_dff_B_AwXEy4nt7_1),.dout(n1022),.clk(gclk));
	jand g0959(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1023),.clk(gclk));
	jand g0960(.dina(w_n1004_0[0]),.dinb(w_n927_0[0]),.dout(n1024),.clk(gclk));
	jand g0961(.dina(w_n1005_0[0]),.dinb(w_n924_0[0]),.dout(n1025),.clk(gclk));
	jor g0962(.dina(n1025),.dinb(w_dff_B_jSsFNk300_1),.dout(n1026),.clk(gclk));
	jand g0963(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1027),.clk(gclk));
	jnot g0964(.din(n1027),.dout(n1028),.clk(gclk));
	jand g0965(.dina(w_n1002_0[0]),.dinb(w_n932_0[0]),.dout(n1029),.clk(gclk));
	jand g0966(.dina(w_n1003_0[0]),.dinb(w_n929_0[0]),.dout(n1030),.clk(gclk));
	jor g0967(.dina(n1030),.dinb(w_dff_B_ldSAnnHy2_1),.dout(n1031),.clk(gclk));
	jand g0968(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1032),.clk(gclk));
	jnot g0969(.din(n1032),.dout(n1033),.clk(gclk));
	jand g0970(.dina(w_n1000_0[0]),.dinb(w_n937_0[0]),.dout(n1034),.clk(gclk));
	jand g0971(.dina(w_n1001_0[0]),.dinb(w_n934_0[0]),.dout(n1035),.clk(gclk));
	jor g0972(.dina(n1035),.dinb(w_dff_B_Nkz8yQSe9_1),.dout(n1036),.clk(gclk));
	jand g0973(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1037),.clk(gclk));
	jnot g0974(.din(n1037),.dout(n1038),.clk(gclk));
	jand g0975(.dina(w_n998_0[0]),.dinb(w_n942_0[0]),.dout(n1039),.clk(gclk));
	jand g0976(.dina(w_n999_0[0]),.dinb(w_n939_0[0]),.dout(n1040),.clk(gclk));
	jor g0977(.dina(n1040),.dinb(w_dff_B_cqPJn0w51_1),.dout(n1041),.clk(gclk));
	jand g0978(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1042),.clk(gclk));
	jnot g0979(.din(n1042),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_n996_0[0]),.dinb(w_n947_0[0]),.dout(n1044),.clk(gclk));
	jand g0981(.dina(w_n997_0[0]),.dinb(w_n944_0[0]),.dout(n1045),.clk(gclk));
	jor g0982(.dina(n1045),.dinb(w_dff_B_7bnw41xC0_1),.dout(n1046),.clk(gclk));
	jand g0983(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1047),.clk(gclk));
	jnot g0984(.din(n1047),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_n994_0[0]),.dinb(w_n952_0[0]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n995_0[0]),.dinb(w_n949_0[0]),.dout(n1050),.clk(gclk));
	jor g0987(.dina(n1050),.dinb(w_dff_B_NUJAPVTH1_1),.dout(n1051),.clk(gclk));
	jand g0988(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1052),.clk(gclk));
	jnot g0989(.din(n1052),.dout(n1053),.clk(gclk));
	jand g0990(.dina(w_n992_0[0]),.dinb(w_n957_0[0]),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n993_0[0]),.dinb(w_n954_0[0]),.dout(n1055),.clk(gclk));
	jor g0992(.dina(n1055),.dinb(w_dff_B_pX2KoYxw6_1),.dout(n1056),.clk(gclk));
	jand g0993(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1057),.clk(gclk));
	jnot g0994(.din(n1057),.dout(n1058),.clk(gclk));
	jand g0995(.dina(w_n990_0[0]),.dinb(w_n962_0[0]),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n991_0[0]),.dinb(w_n959_0[0]),.dout(n1060),.clk(gclk));
	jor g0997(.dina(n1060),.dinb(w_dff_B_cexRrHv16_1),.dout(n1061),.clk(gclk));
	jand g0998(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1062),.clk(gclk));
	jnot g0999(.din(n1062),.dout(n1063),.clk(gclk));
	jand g1000(.dina(w_n988_0[0]),.dinb(w_n967_0[0]),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n989_0[0]),.dinb(w_n964_0[0]),.dout(n1065),.clk(gclk));
	jor g1002(.dina(n1065),.dinb(w_dff_B_lElzpUqB8_1),.dout(n1066),.clk(gclk));
	jand g1003(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1067),.clk(gclk));
	jnot g1004(.din(n1067),.dout(n1068),.clk(gclk));
	jand g1005(.dina(w_n986_0[0]),.dinb(w_n972_0[0]),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n987_0[0]),.dinb(w_n969_0[0]),.dout(n1070),.clk(gclk));
	jor g1007(.dina(n1070),.dinb(w_dff_B_zz5olJJm3_1),.dout(n1071),.clk(gclk));
	jand g1008(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1072),.clk(gclk));
	jnot g1009(.din(n1072),.dout(n1073),.clk(gclk));
	jand g1010(.dina(w_n984_0[0]),.dinb(w_n978_0[0]),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n985_0[0]),.dinb(w_n974_0[0]),.dout(n1075),.clk(gclk));
	jor g1012(.dina(n1075),.dinb(w_dff_B_U2eEKYyt1_1),.dout(n1076),.clk(gclk));
	jand g1013(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1077),.clk(gclk));
	jand g1014(.dina(w_G307gat_2[1]),.dinb(w_G256gat_6[2]),.dout(n1078),.clk(gclk));
	jor g1015(.dina(w_n983_0[0]),.dinb(w_n982_0[0]),.dout(n1079),.clk(gclk));
	jand g1016(.dina(n1079),.dinb(w_n980_0[0]),.dout(n1080),.clk(gclk));
	jxor g1017(.dina(w_n1080_0[1]),.dinb(w_n1078_0[1]),.dout(n1081),.clk(gclk));
	jnot g1018(.din(n1081),.dout(n1082),.clk(gclk));
	jxor g1019(.dina(w_n1082_0[1]),.dinb(w_n1077_0[1]),.dout(n1083),.clk(gclk));
	jxor g1020(.dina(w_n1083_0[1]),.dinb(w_n1076_0[1]),.dout(n1084),.clk(gclk));
	jxor g1021(.dina(w_n1084_0[1]),.dinb(w_n1073_0[1]),.dout(n1085),.clk(gclk));
	jxor g1022(.dina(w_n1085_0[1]),.dinb(w_n1071_0[1]),.dout(n1086),.clk(gclk));
	jxor g1023(.dina(w_n1086_0[1]),.dinb(w_n1068_0[1]),.dout(n1087),.clk(gclk));
	jxor g1024(.dina(w_n1087_0[1]),.dinb(w_n1066_0[1]),.dout(n1088),.clk(gclk));
	jxor g1025(.dina(w_n1088_0[1]),.dinb(w_n1063_0[1]),.dout(n1089),.clk(gclk));
	jxor g1026(.dina(w_n1089_0[1]),.dinb(w_n1061_0[1]),.dout(n1090),.clk(gclk));
	jxor g1027(.dina(w_n1090_0[1]),.dinb(w_n1058_0[1]),.dout(n1091),.clk(gclk));
	jxor g1028(.dina(w_n1091_0[1]),.dinb(w_n1056_0[1]),.dout(n1092),.clk(gclk));
	jxor g1029(.dina(w_n1092_0[1]),.dinb(w_n1053_0[1]),.dout(n1093),.clk(gclk));
	jxor g1030(.dina(w_n1093_0[1]),.dinb(w_n1051_0[1]),.dout(n1094),.clk(gclk));
	jxor g1031(.dina(w_n1094_0[1]),.dinb(w_n1048_0[1]),.dout(n1095),.clk(gclk));
	jxor g1032(.dina(w_n1095_0[1]),.dinb(w_n1046_0[1]),.dout(n1096),.clk(gclk));
	jxor g1033(.dina(w_n1096_0[1]),.dinb(w_n1043_0[1]),.dout(n1097),.clk(gclk));
	jxor g1034(.dina(w_n1097_0[1]),.dinb(w_n1041_0[1]),.dout(n1098),.clk(gclk));
	jxor g1035(.dina(w_n1098_0[1]),.dinb(w_n1038_0[1]),.dout(n1099),.clk(gclk));
	jxor g1036(.dina(w_n1099_0[1]),.dinb(w_n1036_0[1]),.dout(n1100),.clk(gclk));
	jxor g1037(.dina(w_n1100_0[1]),.dinb(w_n1033_0[1]),.dout(n1101),.clk(gclk));
	jxor g1038(.dina(w_n1101_0[1]),.dinb(w_n1031_0[1]),.dout(n1102),.clk(gclk));
	jxor g1039(.dina(w_n1102_0[1]),.dinb(w_n1028_0[1]),.dout(n1103),.clk(gclk));
	jxor g1040(.dina(w_n1103_0[1]),.dinb(w_n1026_0[1]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(n1104),.dout(n1105),.clk(gclk));
	jxor g1042(.dina(w_n1105_0[1]),.dinb(w_n1023_0[1]),.dout(n1106),.clk(gclk));
	jxor g1043(.dina(w_n1106_0[1]),.dinb(w_n1022_0[1]),.dout(n1107),.clk(gclk));
	jxor g1044(.dina(w_n1107_0[1]),.dinb(w_n1018_0[1]),.dout(n1108),.clk(gclk));
	jxor g1045(.dina(w_n1108_0[1]),.dinb(w_n1017_0[1]),.dout(n1109),.clk(gclk));
	jnot g1046(.din(w_n1109_0[1]),.dout(n1110),.clk(gclk));
	jxor g1047(.dina(n1110),.dinb(w_n1013_0[1]),.dout(w_dff_A_JVdXQdwf8_2),.clk(gclk));
	jnot g1048(.din(w_n1108_0[0]),.dout(n1112),.clk(gclk));
	jor g1049(.dina(n1112),.dinb(w_n1017_0[0]),.dout(n1113),.clk(gclk));
	jor g1050(.dina(w_n1109_0[0]),.dinb(w_n1013_0[0]),.dout(n1114),.clk(gclk));
	jand g1051(.dina(n1114),.dinb(w_dff_B_fYgRh1hF7_1),.dout(n1115),.clk(gclk));
	jnot g1052(.din(w_n1106_0[0]),.dout(n1116),.clk(gclk));
	jor g1053(.dina(n1116),.dinb(w_n1022_0[0]),.dout(n1117),.clk(gclk));
	jor g1054(.dina(w_n1107_0[0]),.dinb(w_n1018_0[0]),.dout(n1118),.clk(gclk));
	jand g1055(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jand g1056(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1120),.clk(gclk));
	jand g1057(.dina(w_n1103_0[0]),.dinb(w_n1026_0[0]),.dout(n1121),.clk(gclk));
	jnot g1058(.din(n1121),.dout(n1122),.clk(gclk));
	jor g1059(.dina(w_n1105_0[0]),.dinb(w_n1023_0[0]),.dout(n1123),.clk(gclk));
	jand g1060(.dina(n1123),.dinb(w_dff_B_dTWjquK89_1),.dout(n1124),.clk(gclk));
	jand g1061(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1125),.clk(gclk));
	jnot g1062(.din(n1125),.dout(n1126),.clk(gclk));
	jand g1063(.dina(w_n1101_0[0]),.dinb(w_n1031_0[0]),.dout(n1127),.clk(gclk));
	jand g1064(.dina(w_n1102_0[0]),.dinb(w_n1028_0[0]),.dout(n1128),.clk(gclk));
	jor g1065(.dina(n1128),.dinb(w_dff_B_Y31JGknQ3_1),.dout(n1129),.clk(gclk));
	jand g1066(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1130),.clk(gclk));
	jnot g1067(.din(n1130),.dout(n1131),.clk(gclk));
	jand g1068(.dina(w_n1099_0[0]),.dinb(w_n1036_0[0]),.dout(n1132),.clk(gclk));
	jand g1069(.dina(w_n1100_0[0]),.dinb(w_n1033_0[0]),.dout(n1133),.clk(gclk));
	jor g1070(.dina(n1133),.dinb(w_dff_B_68zJrRQn6_1),.dout(n1134),.clk(gclk));
	jand g1071(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1135),.clk(gclk));
	jnot g1072(.din(n1135),.dout(n1136),.clk(gclk));
	jand g1073(.dina(w_n1097_0[0]),.dinb(w_n1041_0[0]),.dout(n1137),.clk(gclk));
	jand g1074(.dina(w_n1098_0[0]),.dinb(w_n1038_0[0]),.dout(n1138),.clk(gclk));
	jor g1075(.dina(n1138),.dinb(w_dff_B_mSgxvJiU9_1),.dout(n1139),.clk(gclk));
	jand g1076(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1140),.clk(gclk));
	jnot g1077(.din(n1140),.dout(n1141),.clk(gclk));
	jand g1078(.dina(w_n1095_0[0]),.dinb(w_n1046_0[0]),.dout(n1142),.clk(gclk));
	jand g1079(.dina(w_n1096_0[0]),.dinb(w_n1043_0[0]),.dout(n1143),.clk(gclk));
	jor g1080(.dina(n1143),.dinb(w_dff_B_gg2FB3My6_1),.dout(n1144),.clk(gclk));
	jand g1081(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1145),.clk(gclk));
	jnot g1082(.din(n1145),.dout(n1146),.clk(gclk));
	jand g1083(.dina(w_n1093_0[0]),.dinb(w_n1051_0[0]),.dout(n1147),.clk(gclk));
	jand g1084(.dina(w_n1094_0[0]),.dinb(w_n1048_0[0]),.dout(n1148),.clk(gclk));
	jor g1085(.dina(n1148),.dinb(w_dff_B_qGgjE1Rn5_1),.dout(n1149),.clk(gclk));
	jand g1086(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1150),.clk(gclk));
	jnot g1087(.din(n1150),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_n1091_0[0]),.dinb(w_n1056_0[0]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1092_0[0]),.dinb(w_n1053_0[0]),.dout(n1153),.clk(gclk));
	jor g1090(.dina(n1153),.dinb(w_dff_B_6LIhDnGg7_1),.dout(n1154),.clk(gclk));
	jand g1091(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1155),.clk(gclk));
	jnot g1092(.din(n1155),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_n1089_0[0]),.dinb(w_n1061_0[0]),.dout(n1157),.clk(gclk));
	jand g1094(.dina(w_n1090_0[0]),.dinb(w_n1058_0[0]),.dout(n1158),.clk(gclk));
	jor g1095(.dina(n1158),.dinb(w_dff_B_dFvhUsMM4_1),.dout(n1159),.clk(gclk));
	jand g1096(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1160),.clk(gclk));
	jnot g1097(.din(n1160),.dout(n1161),.clk(gclk));
	jand g1098(.dina(w_n1087_0[0]),.dinb(w_n1066_0[0]),.dout(n1162),.clk(gclk));
	jand g1099(.dina(w_n1088_0[0]),.dinb(w_n1063_0[0]),.dout(n1163),.clk(gclk));
	jor g1100(.dina(n1163),.dinb(w_dff_B_Klmu89BJ8_1),.dout(n1164),.clk(gclk));
	jand g1101(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1165),.clk(gclk));
	jnot g1102(.din(n1165),.dout(n1166),.clk(gclk));
	jand g1103(.dina(w_n1085_0[0]),.dinb(w_n1071_0[0]),.dout(n1167),.clk(gclk));
	jand g1104(.dina(w_n1086_0[0]),.dinb(w_n1068_0[0]),.dout(n1168),.clk(gclk));
	jor g1105(.dina(n1168),.dinb(w_dff_B_w6HJXtga9_1),.dout(n1169),.clk(gclk));
	jand g1106(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1170),.clk(gclk));
	jnot g1107(.din(n1170),.dout(n1171),.clk(gclk));
	jand g1108(.dina(w_n1083_0[0]),.dinb(w_n1076_0[0]),.dout(n1172),.clk(gclk));
	jand g1109(.dina(w_n1084_0[0]),.dinb(w_n1073_0[0]),.dout(n1173),.clk(gclk));
	jor g1110(.dina(n1173),.dinb(w_dff_B_EaFpkXqV1_1),.dout(n1174),.clk(gclk));
	jand g1111(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1175),.clk(gclk));
	jand g1112(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1176),.clk(gclk));
	jor g1113(.dina(w_n1080_0[0]),.dinb(w_n1078_0[0]),.dout(n1177),.clk(gclk));
	jor g1114(.dina(w_n1082_0[0]),.dinb(w_n1077_0[0]),.dout(n1178),.clk(gclk));
	jand g1115(.dina(n1178),.dinb(w_dff_B_T8VZlarh2_1),.dout(n1179),.clk(gclk));
	jxor g1116(.dina(w_n1179_0[1]),.dinb(w_n1176_0[1]),.dout(n1180),.clk(gclk));
	jnot g1117(.din(n1180),.dout(n1181),.clk(gclk));
	jxor g1118(.dina(w_n1181_0[1]),.dinb(w_n1175_0[1]),.dout(n1182),.clk(gclk));
	jxor g1119(.dina(w_n1182_0[1]),.dinb(w_n1174_0[1]),.dout(n1183),.clk(gclk));
	jxor g1120(.dina(w_n1183_0[1]),.dinb(w_n1171_0[1]),.dout(n1184),.clk(gclk));
	jxor g1121(.dina(w_n1184_0[1]),.dinb(w_n1169_0[1]),.dout(n1185),.clk(gclk));
	jxor g1122(.dina(w_n1185_0[1]),.dinb(w_n1166_0[1]),.dout(n1186),.clk(gclk));
	jxor g1123(.dina(w_n1186_0[1]),.dinb(w_n1164_0[1]),.dout(n1187),.clk(gclk));
	jxor g1124(.dina(w_n1187_0[1]),.dinb(w_n1161_0[1]),.dout(n1188),.clk(gclk));
	jxor g1125(.dina(w_n1188_0[1]),.dinb(w_n1159_0[1]),.dout(n1189),.clk(gclk));
	jxor g1126(.dina(w_n1189_0[1]),.dinb(w_n1156_0[1]),.dout(n1190),.clk(gclk));
	jxor g1127(.dina(w_n1190_0[1]),.dinb(w_n1154_0[1]),.dout(n1191),.clk(gclk));
	jxor g1128(.dina(w_n1191_0[1]),.dinb(w_n1151_0[1]),.dout(n1192),.clk(gclk));
	jxor g1129(.dina(w_n1192_0[1]),.dinb(w_n1149_0[1]),.dout(n1193),.clk(gclk));
	jxor g1130(.dina(w_n1193_0[1]),.dinb(w_n1146_0[1]),.dout(n1194),.clk(gclk));
	jxor g1131(.dina(w_n1194_0[1]),.dinb(w_n1144_0[1]),.dout(n1195),.clk(gclk));
	jxor g1132(.dina(w_n1195_0[1]),.dinb(w_n1141_0[1]),.dout(n1196),.clk(gclk));
	jxor g1133(.dina(w_n1196_0[1]),.dinb(w_n1139_0[1]),.dout(n1197),.clk(gclk));
	jxor g1134(.dina(w_n1197_0[1]),.dinb(w_n1136_0[1]),.dout(n1198),.clk(gclk));
	jxor g1135(.dina(w_n1198_0[1]),.dinb(w_n1134_0[1]),.dout(n1199),.clk(gclk));
	jxor g1136(.dina(w_n1199_0[1]),.dinb(w_n1131_0[1]),.dout(n1200),.clk(gclk));
	jxor g1137(.dina(w_n1200_0[1]),.dinb(w_n1129_0[1]),.dout(n1201),.clk(gclk));
	jxor g1138(.dina(w_n1201_0[1]),.dinb(w_n1126_0[1]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jxor g1140(.dina(w_n1203_0[1]),.dinb(w_n1124_0[1]),.dout(n1204),.clk(gclk));
	jnot g1141(.din(n1204),.dout(n1205),.clk(gclk));
	jxor g1142(.dina(w_n1205_0[1]),.dinb(w_n1120_0[1]),.dout(n1206),.clk(gclk));
	jxor g1143(.dina(w_n1206_0[1]),.dinb(w_n1119_0[1]),.dout(n1207),.clk(gclk));
	jnot g1144(.din(w_n1207_0[1]),.dout(n1208),.clk(gclk));
	jxor g1145(.dina(n1208),.dinb(w_n1115_0[1]),.dout(w_dff_A_CyfQuo9O5_2),.clk(gclk));
	jnot g1146(.din(w_n1206_0[0]),.dout(n1210),.clk(gclk));
	jor g1147(.dina(n1210),.dinb(w_n1119_0[0]),.dout(n1211),.clk(gclk));
	jor g1148(.dina(w_n1207_0[0]),.dinb(w_n1115_0[0]),.dout(n1212),.clk(gclk));
	jand g1149(.dina(n1212),.dinb(w_dff_B_ybojhGAX3_1),.dout(n1213),.clk(gclk));
	jor g1150(.dina(w_n1203_0[0]),.dinb(w_n1124_0[0]),.dout(n1214),.clk(gclk));
	jor g1151(.dina(w_n1205_0[0]),.dinb(w_n1120_0[0]),.dout(n1215),.clk(gclk));
	jand g1152(.dina(n1215),.dinb(w_dff_B_dNEC8t638_1),.dout(n1216),.clk(gclk));
	jand g1153(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1217),.clk(gclk));
	jand g1154(.dina(w_n1200_0[0]),.dinb(w_n1129_0[0]),.dout(n1218),.clk(gclk));
	jand g1155(.dina(w_n1201_0[0]),.dinb(w_n1126_0[0]),.dout(n1219),.clk(gclk));
	jor g1156(.dina(n1219),.dinb(w_dff_B_I4hnYSxQ2_1),.dout(n1220),.clk(gclk));
	jand g1157(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1221),.clk(gclk));
	jnot g1158(.din(n1221),.dout(n1222),.clk(gclk));
	jand g1159(.dina(w_n1198_0[0]),.dinb(w_n1134_0[0]),.dout(n1223),.clk(gclk));
	jand g1160(.dina(w_n1199_0[0]),.dinb(w_n1131_0[0]),.dout(n1224),.clk(gclk));
	jor g1161(.dina(n1224),.dinb(w_dff_B_5a7iCyKw7_1),.dout(n1225),.clk(gclk));
	jand g1162(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1226),.clk(gclk));
	jnot g1163(.din(n1226),.dout(n1227),.clk(gclk));
	jand g1164(.dina(w_n1196_0[0]),.dinb(w_n1139_0[0]),.dout(n1228),.clk(gclk));
	jand g1165(.dina(w_n1197_0[0]),.dinb(w_n1136_0[0]),.dout(n1229),.clk(gclk));
	jor g1166(.dina(n1229),.dinb(w_dff_B_Ncrix9Co4_1),.dout(n1230),.clk(gclk));
	jand g1167(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1231),.clk(gclk));
	jnot g1168(.din(n1231),.dout(n1232),.clk(gclk));
	jand g1169(.dina(w_n1194_0[0]),.dinb(w_n1144_0[0]),.dout(n1233),.clk(gclk));
	jand g1170(.dina(w_n1195_0[0]),.dinb(w_n1141_0[0]),.dout(n1234),.clk(gclk));
	jor g1171(.dina(n1234),.dinb(w_dff_B_rlehoPlh3_1),.dout(n1235),.clk(gclk));
	jand g1172(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1236),.clk(gclk));
	jnot g1173(.din(n1236),.dout(n1237),.clk(gclk));
	jand g1174(.dina(w_n1192_0[0]),.dinb(w_n1149_0[0]),.dout(n1238),.clk(gclk));
	jand g1175(.dina(w_n1193_0[0]),.dinb(w_n1146_0[0]),.dout(n1239),.clk(gclk));
	jor g1176(.dina(n1239),.dinb(w_dff_B_zIUS8s871_1),.dout(n1240),.clk(gclk));
	jand g1177(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1241),.clk(gclk));
	jnot g1178(.din(n1241),.dout(n1242),.clk(gclk));
	jand g1179(.dina(w_n1190_0[0]),.dinb(w_n1154_0[0]),.dout(n1243),.clk(gclk));
	jand g1180(.dina(w_n1191_0[0]),.dinb(w_n1151_0[0]),.dout(n1244),.clk(gclk));
	jor g1181(.dina(n1244),.dinb(w_dff_B_NTV0JpaY7_1),.dout(n1245),.clk(gclk));
	jand g1182(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1246),.clk(gclk));
	jnot g1183(.din(n1246),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_n1188_0[0]),.dinb(w_n1159_0[0]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1189_0[0]),.dinb(w_n1156_0[0]),.dout(n1249),.clk(gclk));
	jor g1186(.dina(n1249),.dinb(w_dff_B_r1b8WR3B7_1),.dout(n1250),.clk(gclk));
	jand g1187(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1251),.clk(gclk));
	jnot g1188(.din(n1251),.dout(n1252),.clk(gclk));
	jand g1189(.dina(w_n1186_0[0]),.dinb(w_n1164_0[0]),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1187_0[0]),.dinb(w_n1161_0[0]),.dout(n1254),.clk(gclk));
	jor g1191(.dina(n1254),.dinb(w_dff_B_XA6EwYAF0_1),.dout(n1255),.clk(gclk));
	jand g1192(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1256),.clk(gclk));
	jnot g1193(.din(n1256),.dout(n1257),.clk(gclk));
	jand g1194(.dina(w_n1184_0[0]),.dinb(w_n1169_0[0]),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1185_0[0]),.dinb(w_n1166_0[0]),.dout(n1259),.clk(gclk));
	jor g1196(.dina(n1259),.dinb(w_dff_B_QNM7Qz8B1_1),.dout(n1260),.clk(gclk));
	jand g1197(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1261),.clk(gclk));
	jnot g1198(.din(n1261),.dout(n1262),.clk(gclk));
	jand g1199(.dina(w_n1182_0[0]),.dinb(w_n1174_0[0]),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1183_0[0]),.dinb(w_n1171_0[0]),.dout(n1264),.clk(gclk));
	jor g1201(.dina(n1264),.dinb(w_dff_B_rMz0XjOQ0_1),.dout(n1265),.clk(gclk));
	jand g1202(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1266),.clk(gclk));
	jand g1203(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1267),.clk(gclk));
	jor g1204(.dina(w_n1179_0[0]),.dinb(w_n1176_0[0]),.dout(n1268),.clk(gclk));
	jor g1205(.dina(w_n1181_0[0]),.dinb(w_n1175_0[0]),.dout(n1269),.clk(gclk));
	jand g1206(.dina(n1269),.dinb(w_dff_B_DY66GdNE4_1),.dout(n1270),.clk(gclk));
	jxor g1207(.dina(w_n1270_0[1]),.dinb(w_n1267_0[1]),.dout(n1271),.clk(gclk));
	jnot g1208(.din(n1271),.dout(n1272),.clk(gclk));
	jxor g1209(.dina(w_n1272_0[1]),.dinb(w_n1266_0[1]),.dout(n1273),.clk(gclk));
	jxor g1210(.dina(w_n1273_0[1]),.dinb(w_n1265_0[1]),.dout(n1274),.clk(gclk));
	jxor g1211(.dina(w_n1274_0[1]),.dinb(w_n1262_0[1]),.dout(n1275),.clk(gclk));
	jxor g1212(.dina(w_n1275_0[1]),.dinb(w_n1260_0[1]),.dout(n1276),.clk(gclk));
	jxor g1213(.dina(w_n1276_0[1]),.dinb(w_n1257_0[1]),.dout(n1277),.clk(gclk));
	jxor g1214(.dina(w_n1277_0[1]),.dinb(w_n1255_0[1]),.dout(n1278),.clk(gclk));
	jxor g1215(.dina(w_n1278_0[1]),.dinb(w_n1252_0[1]),.dout(n1279),.clk(gclk));
	jxor g1216(.dina(w_n1279_0[1]),.dinb(w_n1250_0[1]),.dout(n1280),.clk(gclk));
	jxor g1217(.dina(w_n1280_0[1]),.dinb(w_n1247_0[1]),.dout(n1281),.clk(gclk));
	jxor g1218(.dina(w_n1281_0[1]),.dinb(w_n1245_0[1]),.dout(n1282),.clk(gclk));
	jxor g1219(.dina(w_n1282_0[1]),.dinb(w_n1242_0[1]),.dout(n1283),.clk(gclk));
	jxor g1220(.dina(w_n1283_0[1]),.dinb(w_n1240_0[1]),.dout(n1284),.clk(gclk));
	jxor g1221(.dina(w_n1284_0[1]),.dinb(w_n1237_0[1]),.dout(n1285),.clk(gclk));
	jxor g1222(.dina(w_n1285_0[1]),.dinb(w_n1235_0[1]),.dout(n1286),.clk(gclk));
	jxor g1223(.dina(w_n1286_0[1]),.dinb(w_n1232_0[1]),.dout(n1287),.clk(gclk));
	jxor g1224(.dina(w_n1287_0[1]),.dinb(w_n1230_0[1]),.dout(n1288),.clk(gclk));
	jxor g1225(.dina(w_n1288_0[1]),.dinb(w_n1227_0[1]),.dout(n1289),.clk(gclk));
	jxor g1226(.dina(w_n1289_0[1]),.dinb(w_n1225_0[1]),.dout(n1290),.clk(gclk));
	jxor g1227(.dina(w_n1290_0[1]),.dinb(w_n1222_0[1]),.dout(n1291),.clk(gclk));
	jxor g1228(.dina(w_n1291_0[1]),.dinb(w_n1220_0[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jxor g1230(.dina(w_n1293_0[1]),.dinb(w_n1217_0[1]),.dout(n1294),.clk(gclk));
	jxor g1231(.dina(w_n1294_0[1]),.dinb(w_n1216_0[1]),.dout(n1295),.clk(gclk));
	jnot g1232(.din(w_n1295_0[1]),.dout(n1296),.clk(gclk));
	jxor g1233(.dina(w_dff_B_4SLee9TS5_0),.dinb(w_n1213_0[1]),.dout(w_dff_A_MLPL8Tm53_2),.clk(gclk));
	jnot g1234(.din(w_n1294_0[0]),.dout(n1298),.clk(gclk));
	jor g1235(.dina(w_dff_B_T7uFMeCt1_0),.dinb(w_n1216_0[0]),.dout(n1299),.clk(gclk));
	jor g1236(.dina(w_n1295_0[0]),.dinb(w_n1213_0[0]),.dout(n1300),.clk(gclk));
	jand g1237(.dina(n1300),.dinb(w_dff_B_Koc5iBCH3_1),.dout(n1301),.clk(gclk));
	jnot g1238(.din(w_n1220_0[0]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(w_n1291_0[0]),.dout(n1303),.clk(gclk));
	jor g1240(.dina(w_dff_B_WbgLpl9P7_0),.dinb(n1302),.dout(n1304),.clk(gclk));
	jor g1241(.dina(w_n1293_0[0]),.dinb(w_n1217_0[0]),.dout(n1305),.clk(gclk));
	jand g1242(.dina(n1305),.dinb(w_dff_B_SgiYHoB16_1),.dout(n1306),.clk(gclk));
	jand g1243(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1307),.clk(gclk));
	jand g1244(.dina(w_n1289_0[0]),.dinb(w_n1225_0[0]),.dout(n1308),.clk(gclk));
	jand g1245(.dina(w_n1290_0[0]),.dinb(w_n1222_0[0]),.dout(n1309),.clk(gclk));
	jor g1246(.dina(n1309),.dinb(w_dff_B_IZi3Ndf67_1),.dout(n1310),.clk(gclk));
	jand g1247(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1311),.clk(gclk));
	jnot g1248(.din(n1311),.dout(n1312),.clk(gclk));
	jand g1249(.dina(w_n1287_0[0]),.dinb(w_n1230_0[0]),.dout(n1313),.clk(gclk));
	jand g1250(.dina(w_n1288_0[0]),.dinb(w_n1227_0[0]),.dout(n1314),.clk(gclk));
	jor g1251(.dina(n1314),.dinb(w_dff_B_p1ySQhIb4_1),.dout(n1315),.clk(gclk));
	jand g1252(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1316),.clk(gclk));
	jnot g1253(.din(n1316),.dout(n1317),.clk(gclk));
	jand g1254(.dina(w_n1285_0[0]),.dinb(w_n1235_0[0]),.dout(n1318),.clk(gclk));
	jand g1255(.dina(w_n1286_0[0]),.dinb(w_n1232_0[0]),.dout(n1319),.clk(gclk));
	jor g1256(.dina(n1319),.dinb(w_dff_B_htxOHOD62_1),.dout(n1320),.clk(gclk));
	jand g1257(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1321),.clk(gclk));
	jnot g1258(.din(n1321),.dout(n1322),.clk(gclk));
	jand g1259(.dina(w_n1283_0[0]),.dinb(w_n1240_0[0]),.dout(n1323),.clk(gclk));
	jand g1260(.dina(w_n1284_0[0]),.dinb(w_n1237_0[0]),.dout(n1324),.clk(gclk));
	jor g1261(.dina(n1324),.dinb(w_dff_B_LbZi72ql7_1),.dout(n1325),.clk(gclk));
	jand g1262(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(n1326),.dout(n1327),.clk(gclk));
	jand g1264(.dina(w_n1281_0[0]),.dinb(w_n1245_0[0]),.dout(n1328),.clk(gclk));
	jand g1265(.dina(w_n1282_0[0]),.dinb(w_n1242_0[0]),.dout(n1329),.clk(gclk));
	jor g1266(.dina(n1329),.dinb(w_dff_B_XsKObT771_1),.dout(n1330),.clk(gclk));
	jand g1267(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1331),.clk(gclk));
	jnot g1268(.din(n1331),.dout(n1332),.clk(gclk));
	jand g1269(.dina(w_n1279_0[0]),.dinb(w_n1250_0[0]),.dout(n1333),.clk(gclk));
	jand g1270(.dina(w_n1280_0[0]),.dinb(w_n1247_0[0]),.dout(n1334),.clk(gclk));
	jor g1271(.dina(n1334),.dinb(w_dff_B_3YJs9FYL7_1),.dout(n1335),.clk(gclk));
	jand g1272(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1336),.clk(gclk));
	jnot g1273(.din(n1336),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_n1277_0[0]),.dinb(w_n1255_0[0]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1278_0[0]),.dinb(w_n1252_0[0]),.dout(n1339),.clk(gclk));
	jor g1276(.dina(n1339),.dinb(w_dff_B_RCvdprrW0_1),.dout(n1340),.clk(gclk));
	jand g1277(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1341),.clk(gclk));
	jnot g1278(.din(n1341),.dout(n1342),.clk(gclk));
	jand g1279(.dina(w_n1275_0[0]),.dinb(w_n1260_0[0]),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1276_0[0]),.dinb(w_n1257_0[0]),.dout(n1344),.clk(gclk));
	jor g1281(.dina(n1344),.dinb(w_dff_B_5mHjtuOZ5_1),.dout(n1345),.clk(gclk));
	jand g1282(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1346),.clk(gclk));
	jnot g1283(.din(n1346),.dout(n1347),.clk(gclk));
	jand g1284(.dina(w_n1273_0[0]),.dinb(w_n1265_0[0]),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1274_0[0]),.dinb(w_n1262_0[0]),.dout(n1349),.clk(gclk));
	jor g1286(.dina(n1349),.dinb(w_dff_B_fF22xHZ72_1),.dout(n1350),.clk(gclk));
	jand g1287(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1351),.clk(gclk));
	jand g1288(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1352),.clk(gclk));
	jor g1289(.dina(w_n1270_0[0]),.dinb(w_n1267_0[0]),.dout(n1353),.clk(gclk));
	jor g1290(.dina(w_n1272_0[0]),.dinb(w_n1266_0[0]),.dout(n1354),.clk(gclk));
	jand g1291(.dina(n1354),.dinb(w_dff_B_qLfpP2yC6_1),.dout(n1355),.clk(gclk));
	jxor g1292(.dina(w_n1355_0[1]),.dinb(w_n1352_0[1]),.dout(n1356),.clk(gclk));
	jnot g1293(.din(n1356),.dout(n1357),.clk(gclk));
	jxor g1294(.dina(w_n1357_0[1]),.dinb(w_n1351_0[1]),.dout(n1358),.clk(gclk));
	jxor g1295(.dina(w_n1358_0[1]),.dinb(w_n1350_0[1]),.dout(n1359),.clk(gclk));
	jxor g1296(.dina(w_n1359_0[1]),.dinb(w_n1347_0[1]),.dout(n1360),.clk(gclk));
	jxor g1297(.dina(w_n1360_0[1]),.dinb(w_n1345_0[1]),.dout(n1361),.clk(gclk));
	jxor g1298(.dina(w_n1361_0[1]),.dinb(w_n1342_0[1]),.dout(n1362),.clk(gclk));
	jxor g1299(.dina(w_n1362_0[1]),.dinb(w_n1340_0[1]),.dout(n1363),.clk(gclk));
	jxor g1300(.dina(w_n1363_0[1]),.dinb(w_n1337_0[1]),.dout(n1364),.clk(gclk));
	jxor g1301(.dina(w_n1364_0[1]),.dinb(w_n1335_0[1]),.dout(n1365),.clk(gclk));
	jxor g1302(.dina(w_n1365_0[1]),.dinb(w_n1332_0[1]),.dout(n1366),.clk(gclk));
	jxor g1303(.dina(w_n1366_0[1]),.dinb(w_n1330_0[1]),.dout(n1367),.clk(gclk));
	jxor g1304(.dina(w_n1367_0[1]),.dinb(w_n1327_0[1]),.dout(n1368),.clk(gclk));
	jxor g1305(.dina(w_n1368_0[1]),.dinb(w_n1325_0[1]),.dout(n1369),.clk(gclk));
	jxor g1306(.dina(w_n1369_0[1]),.dinb(w_n1322_0[1]),.dout(n1370),.clk(gclk));
	jxor g1307(.dina(w_n1370_0[1]),.dinb(w_n1320_0[1]),.dout(n1371),.clk(gclk));
	jxor g1308(.dina(w_n1371_0[1]),.dinb(w_n1317_0[1]),.dout(n1372),.clk(gclk));
	jxor g1309(.dina(w_n1372_0[1]),.dinb(w_n1315_0[1]),.dout(n1373),.clk(gclk));
	jxor g1310(.dina(w_n1373_0[1]),.dinb(w_n1312_0[1]),.dout(n1374),.clk(gclk));
	jxor g1311(.dina(w_n1374_0[1]),.dinb(w_n1310_0[1]),.dout(n1375),.clk(gclk));
	jnot g1312(.din(n1375),.dout(n1376),.clk(gclk));
	jxor g1313(.dina(w_n1376_0[1]),.dinb(w_n1307_0[1]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jxor g1315(.dina(w_n1378_0[1]),.dinb(w_n1306_0[1]),.dout(n1379),.clk(gclk));
	jxor g1316(.dina(w_n1379_0[1]),.dinb(w_n1301_0[1]),.dout(w_dff_A_n713uqzH6_2),.clk(gclk));
	jor g1317(.dina(w_n1378_0[0]),.dinb(w_n1306_0[0]),.dout(n1381),.clk(gclk));
	jnot g1318(.din(w_n1379_0[0]),.dout(n1382),.clk(gclk));
	jor g1319(.dina(w_dff_B_cQ4vJJdm6_0),.dinb(w_n1301_0[0]),.dout(n1383),.clk(gclk));
	jand g1320(.dina(n1383),.dinb(w_dff_B_tmWz7Xxw0_1),.dout(n1384),.clk(gclk));
	jnot g1321(.din(w_n1310_0[0]),.dout(n1385),.clk(gclk));
	jnot g1322(.din(w_n1374_0[0]),.dout(n1386),.clk(gclk));
	jor g1323(.dina(n1386),.dinb(n1385),.dout(n1387),.clk(gclk));
	jor g1324(.dina(w_n1376_0[0]),.dinb(w_n1307_0[0]),.dout(n1388),.clk(gclk));
	jand g1325(.dina(n1388),.dinb(w_dff_B_NXjw3b0q3_1),.dout(n1389),.clk(gclk));
	jand g1326(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1390),.clk(gclk));
	jand g1327(.dina(w_n1372_0[0]),.dinb(w_n1315_0[0]),.dout(n1391),.clk(gclk));
	jand g1328(.dina(w_n1373_0[0]),.dinb(w_n1312_0[0]),.dout(n1392),.clk(gclk));
	jor g1329(.dina(n1392),.dinb(w_dff_B_xAz4mD5f3_1),.dout(n1393),.clk(gclk));
	jand g1330(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1394),.clk(gclk));
	jnot g1331(.din(n1394),.dout(n1395),.clk(gclk));
	jand g1332(.dina(w_n1370_0[0]),.dinb(w_n1320_0[0]),.dout(n1396),.clk(gclk));
	jand g1333(.dina(w_n1371_0[0]),.dinb(w_n1317_0[0]),.dout(n1397),.clk(gclk));
	jor g1334(.dina(n1397),.dinb(w_dff_B_lZcZVzdw3_1),.dout(n1398),.clk(gclk));
	jand g1335(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1399),.clk(gclk));
	jnot g1336(.din(n1399),.dout(n1400),.clk(gclk));
	jand g1337(.dina(w_n1368_0[0]),.dinb(w_n1325_0[0]),.dout(n1401),.clk(gclk));
	jand g1338(.dina(w_n1369_0[0]),.dinb(w_n1322_0[0]),.dout(n1402),.clk(gclk));
	jor g1339(.dina(n1402),.dinb(w_dff_B_mI1SzJPV7_1),.dout(n1403),.clk(gclk));
	jand g1340(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1404),.clk(gclk));
	jnot g1341(.din(n1404),.dout(n1405),.clk(gclk));
	jand g1342(.dina(w_n1366_0[0]),.dinb(w_n1330_0[0]),.dout(n1406),.clk(gclk));
	jand g1343(.dina(w_n1367_0[0]),.dinb(w_n1327_0[0]),.dout(n1407),.clk(gclk));
	jor g1344(.dina(n1407),.dinb(w_dff_B_Q0KMD2eo2_1),.dout(n1408),.clk(gclk));
	jand g1345(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1409),.clk(gclk));
	jnot g1346(.din(n1409),.dout(n1410),.clk(gclk));
	jand g1347(.dina(w_n1364_0[0]),.dinb(w_n1335_0[0]),.dout(n1411),.clk(gclk));
	jand g1348(.dina(w_n1365_0[0]),.dinb(w_n1332_0[0]),.dout(n1412),.clk(gclk));
	jor g1349(.dina(n1412),.dinb(w_dff_B_03C4d0Nz5_1),.dout(n1413),.clk(gclk));
	jand g1350(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1414),.clk(gclk));
	jnot g1351(.din(n1414),.dout(n1415),.clk(gclk));
	jand g1352(.dina(w_n1362_0[0]),.dinb(w_n1340_0[0]),.dout(n1416),.clk(gclk));
	jand g1353(.dina(w_n1363_0[0]),.dinb(w_n1337_0[0]),.dout(n1417),.clk(gclk));
	jor g1354(.dina(n1417),.dinb(w_dff_B_fhgkpsz11_1),.dout(n1418),.clk(gclk));
	jand g1355(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1419),.clk(gclk));
	jnot g1356(.din(n1419),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_n1360_0[0]),.dinb(w_n1345_0[0]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1361_0[0]),.dinb(w_n1342_0[0]),.dout(n1422),.clk(gclk));
	jor g1359(.dina(n1422),.dinb(w_dff_B_LJDxjFoi4_1),.dout(n1423),.clk(gclk));
	jand g1360(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1424),.clk(gclk));
	jnot g1361(.din(n1424),.dout(n1425),.clk(gclk));
	jand g1362(.dina(w_n1358_0[0]),.dinb(w_n1350_0[0]),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1359_0[0]),.dinb(w_n1347_0[0]),.dout(n1427),.clk(gclk));
	jor g1364(.dina(n1427),.dinb(w_dff_B_xvrIb0mS9_1),.dout(n1428),.clk(gclk));
	jand g1365(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1429),.clk(gclk));
	jand g1366(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1430),.clk(gclk));
	jor g1367(.dina(w_n1355_0[0]),.dinb(w_n1352_0[0]),.dout(n1431),.clk(gclk));
	jor g1368(.dina(w_n1357_0[0]),.dinb(w_n1351_0[0]),.dout(n1432),.clk(gclk));
	jand g1369(.dina(n1432),.dinb(w_dff_B_WWR6ioqC4_1),.dout(n1433),.clk(gclk));
	jxor g1370(.dina(w_n1433_0[1]),.dinb(w_n1430_0[1]),.dout(n1434),.clk(gclk));
	jnot g1371(.din(n1434),.dout(n1435),.clk(gclk));
	jxor g1372(.dina(w_n1435_0[1]),.dinb(w_n1429_0[1]),.dout(n1436),.clk(gclk));
	jxor g1373(.dina(w_n1436_0[1]),.dinb(w_n1428_0[1]),.dout(n1437),.clk(gclk));
	jxor g1374(.dina(w_n1437_0[1]),.dinb(w_n1425_0[1]),.dout(n1438),.clk(gclk));
	jxor g1375(.dina(w_n1438_0[1]),.dinb(w_n1423_0[1]),.dout(n1439),.clk(gclk));
	jxor g1376(.dina(w_n1439_0[1]),.dinb(w_n1420_0[1]),.dout(n1440),.clk(gclk));
	jxor g1377(.dina(w_n1440_0[1]),.dinb(w_n1418_0[1]),.dout(n1441),.clk(gclk));
	jxor g1378(.dina(w_n1441_0[1]),.dinb(w_n1415_0[1]),.dout(n1442),.clk(gclk));
	jxor g1379(.dina(w_n1442_0[1]),.dinb(w_n1413_0[1]),.dout(n1443),.clk(gclk));
	jxor g1380(.dina(w_n1443_0[1]),.dinb(w_n1410_0[1]),.dout(n1444),.clk(gclk));
	jxor g1381(.dina(w_n1444_0[1]),.dinb(w_n1408_0[1]),.dout(n1445),.clk(gclk));
	jxor g1382(.dina(w_n1445_0[1]),.dinb(w_n1405_0[1]),.dout(n1446),.clk(gclk));
	jxor g1383(.dina(w_n1446_0[1]),.dinb(w_n1403_0[1]),.dout(n1447),.clk(gclk));
	jxor g1384(.dina(w_n1447_0[1]),.dinb(w_n1400_0[1]),.dout(n1448),.clk(gclk));
	jxor g1385(.dina(w_n1448_0[1]),.dinb(w_n1398_0[1]),.dout(n1449),.clk(gclk));
	jxor g1386(.dina(w_n1449_0[1]),.dinb(w_n1395_0[1]),.dout(n1450),.clk(gclk));
	jxor g1387(.dina(w_n1450_0[1]),.dinb(w_n1393_0[1]),.dout(n1451),.clk(gclk));
	jnot g1388(.din(n1451),.dout(n1452),.clk(gclk));
	jxor g1389(.dina(w_n1452_0[1]),.dinb(w_n1390_0[1]),.dout(n1453),.clk(gclk));
	jnot g1390(.din(n1453),.dout(n1454),.clk(gclk));
	jxor g1391(.dina(w_n1454_0[1]),.dinb(w_n1389_0[1]),.dout(n1455),.clk(gclk));
	jxor g1392(.dina(w_n1455_0[1]),.dinb(w_n1384_0[1]),.dout(w_dff_A_uHImcr829_2),.clk(gclk));
	jor g1393(.dina(w_n1454_0[0]),.dinb(w_n1389_0[0]),.dout(n1457),.clk(gclk));
	jnot g1394(.din(w_n1455_0[0]),.dout(n1458),.clk(gclk));
	jor g1395(.dina(w_dff_B_KxTD4Scz6_0),.dinb(w_n1384_0[0]),.dout(n1459),.clk(gclk));
	jand g1396(.dina(n1459),.dinb(w_dff_B_ubHAw9xw6_1),.dout(n1460),.clk(gclk));
	jnot g1397(.din(w_n1393_0[0]),.dout(n1461),.clk(gclk));
	jnot g1398(.din(w_n1450_0[0]),.dout(n1462),.clk(gclk));
	jor g1399(.dina(n1462),.dinb(n1461),.dout(n1463),.clk(gclk));
	jor g1400(.dina(w_n1452_0[0]),.dinb(w_n1390_0[0]),.dout(n1464),.clk(gclk));
	jand g1401(.dina(n1464),.dinb(w_dff_B_fcHIml3A7_1),.dout(n1465),.clk(gclk));
	jand g1402(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1466),.clk(gclk));
	jand g1403(.dina(w_n1448_0[0]),.dinb(w_n1398_0[0]),.dout(n1467),.clk(gclk));
	jand g1404(.dina(w_n1449_0[0]),.dinb(w_n1395_0[0]),.dout(n1468),.clk(gclk));
	jor g1405(.dina(n1468),.dinb(w_dff_B_1aMAG6Sh9_1),.dout(n1469),.clk(gclk));
	jand g1406(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1470),.clk(gclk));
	jnot g1407(.din(n1470),.dout(n1471),.clk(gclk));
	jand g1408(.dina(w_n1446_0[0]),.dinb(w_n1403_0[0]),.dout(n1472),.clk(gclk));
	jand g1409(.dina(w_n1447_0[0]),.dinb(w_n1400_0[0]),.dout(n1473),.clk(gclk));
	jor g1410(.dina(n1473),.dinb(w_dff_B_jJuYpWOA2_1),.dout(n1474),.clk(gclk));
	jand g1411(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1475),.clk(gclk));
	jnot g1412(.din(n1475),.dout(n1476),.clk(gclk));
	jand g1413(.dina(w_n1444_0[0]),.dinb(w_n1408_0[0]),.dout(n1477),.clk(gclk));
	jand g1414(.dina(w_n1445_0[0]),.dinb(w_n1405_0[0]),.dout(n1478),.clk(gclk));
	jor g1415(.dina(n1478),.dinb(w_dff_B_O45oxs1m1_1),.dout(n1479),.clk(gclk));
	jand g1416(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1480),.clk(gclk));
	jnot g1417(.din(n1480),.dout(n1481),.clk(gclk));
	jand g1418(.dina(w_n1442_0[0]),.dinb(w_n1413_0[0]),.dout(n1482),.clk(gclk));
	jand g1419(.dina(w_n1443_0[0]),.dinb(w_n1410_0[0]),.dout(n1483),.clk(gclk));
	jor g1420(.dina(n1483),.dinb(w_dff_B_1GGwFMXf4_1),.dout(n1484),.clk(gclk));
	jand g1421(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1485),.clk(gclk));
	jnot g1422(.din(n1485),.dout(n1486),.clk(gclk));
	jand g1423(.dina(w_n1440_0[0]),.dinb(w_n1418_0[0]),.dout(n1487),.clk(gclk));
	jand g1424(.dina(w_n1441_0[0]),.dinb(w_n1415_0[0]),.dout(n1488),.clk(gclk));
	jor g1425(.dina(n1488),.dinb(w_dff_B_KqDwvtXB8_1),.dout(n1489),.clk(gclk));
	jand g1426(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1490),.clk(gclk));
	jnot g1427(.din(n1490),.dout(n1491),.clk(gclk));
	jand g1428(.dina(w_n1438_0[0]),.dinb(w_n1423_0[0]),.dout(n1492),.clk(gclk));
	jand g1429(.dina(w_n1439_0[0]),.dinb(w_n1420_0[0]),.dout(n1493),.clk(gclk));
	jor g1430(.dina(n1493),.dinb(w_dff_B_I86KhtRw2_1),.dout(n1494),.clk(gclk));
	jand g1431(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1495),.clk(gclk));
	jnot g1432(.din(n1495),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_n1436_0[0]),.dinb(w_n1428_0[0]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1437_0[0]),.dinb(w_n1425_0[0]),.dout(n1498),.clk(gclk));
	jor g1435(.dina(n1498),.dinb(w_dff_B_Qgbz1cZp2_1),.dout(n1499),.clk(gclk));
	jand g1436(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1500),.clk(gclk));
	jand g1437(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1501),.clk(gclk));
	jor g1438(.dina(w_n1433_0[0]),.dinb(w_n1430_0[0]),.dout(n1502),.clk(gclk));
	jor g1439(.dina(w_n1435_0[0]),.dinb(w_n1429_0[0]),.dout(n1503),.clk(gclk));
	jand g1440(.dina(n1503),.dinb(w_dff_B_jkG7Gnh21_1),.dout(n1504),.clk(gclk));
	jxor g1441(.dina(w_n1504_0[1]),.dinb(w_n1501_0[1]),.dout(n1505),.clk(gclk));
	jnot g1442(.din(n1505),.dout(n1506),.clk(gclk));
	jxor g1443(.dina(w_n1506_0[1]),.dinb(w_n1500_0[1]),.dout(n1507),.clk(gclk));
	jxor g1444(.dina(w_n1507_0[1]),.dinb(w_n1499_0[1]),.dout(n1508),.clk(gclk));
	jxor g1445(.dina(w_n1508_0[1]),.dinb(w_n1496_0[1]),.dout(n1509),.clk(gclk));
	jxor g1446(.dina(w_n1509_0[1]),.dinb(w_n1494_0[1]),.dout(n1510),.clk(gclk));
	jxor g1447(.dina(w_n1510_0[1]),.dinb(w_n1491_0[1]),.dout(n1511),.clk(gclk));
	jxor g1448(.dina(w_n1511_0[1]),.dinb(w_n1489_0[1]),.dout(n1512),.clk(gclk));
	jxor g1449(.dina(w_n1512_0[1]),.dinb(w_n1486_0[1]),.dout(n1513),.clk(gclk));
	jxor g1450(.dina(w_n1513_0[1]),.dinb(w_n1484_0[1]),.dout(n1514),.clk(gclk));
	jxor g1451(.dina(w_n1514_0[1]),.dinb(w_n1481_0[1]),.dout(n1515),.clk(gclk));
	jxor g1452(.dina(w_n1515_0[1]),.dinb(w_n1479_0[1]),.dout(n1516),.clk(gclk));
	jxor g1453(.dina(w_n1516_0[1]),.dinb(w_n1476_0[1]),.dout(n1517),.clk(gclk));
	jxor g1454(.dina(w_n1517_0[1]),.dinb(w_n1474_0[1]),.dout(n1518),.clk(gclk));
	jxor g1455(.dina(w_n1518_0[1]),.dinb(w_n1471_0[1]),.dout(n1519),.clk(gclk));
	jxor g1456(.dina(w_n1519_0[1]),.dinb(w_n1469_0[1]),.dout(n1520),.clk(gclk));
	jnot g1457(.din(n1520),.dout(n1521),.clk(gclk));
	jxor g1458(.dina(w_n1521_0[1]),.dinb(w_n1466_0[1]),.dout(n1522),.clk(gclk));
	jnot g1459(.din(n1522),.dout(n1523),.clk(gclk));
	jxor g1460(.dina(w_n1523_0[1]),.dinb(w_n1465_0[1]),.dout(n1524),.clk(gclk));
	jxor g1461(.dina(w_n1524_0[1]),.dinb(w_n1460_0[1]),.dout(w_dff_A_IVpIwNKv9_2),.clk(gclk));
	jor g1462(.dina(w_n1523_0[0]),.dinb(w_n1465_0[0]),.dout(n1526),.clk(gclk));
	jnot g1463(.din(w_n1524_0[0]),.dout(n1527),.clk(gclk));
	jor g1464(.dina(w_dff_B_J0oQAQk06_0),.dinb(w_n1460_0[0]),.dout(n1528),.clk(gclk));
	jand g1465(.dina(n1528),.dinb(w_dff_B_D3AzhsqY2_1),.dout(n1529),.clk(gclk));
	jnot g1466(.din(w_n1469_0[0]),.dout(n1530),.clk(gclk));
	jnot g1467(.din(w_n1519_0[0]),.dout(n1531),.clk(gclk));
	jor g1468(.dina(w_dff_B_1ax3ECta3_0),.dinb(n1530),.dout(n1532),.clk(gclk));
	jor g1469(.dina(w_n1521_0[0]),.dinb(w_n1466_0[0]),.dout(n1533),.clk(gclk));
	jand g1470(.dina(n1533),.dinb(w_dff_B_Jk58wg5I9_1),.dout(n1534),.clk(gclk));
	jand g1471(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1535),.clk(gclk));
	jand g1472(.dina(w_n1517_0[0]),.dinb(w_n1474_0[0]),.dout(n1536),.clk(gclk));
	jand g1473(.dina(w_n1518_0[0]),.dinb(w_n1471_0[0]),.dout(n1537),.clk(gclk));
	jor g1474(.dina(n1537),.dinb(w_dff_B_zsNagZtx2_1),.dout(n1538),.clk(gclk));
	jand g1475(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1539),.clk(gclk));
	jnot g1476(.din(n1539),.dout(n1540),.clk(gclk));
	jand g1477(.dina(w_n1515_0[0]),.dinb(w_n1479_0[0]),.dout(n1541),.clk(gclk));
	jand g1478(.dina(w_n1516_0[0]),.dinb(w_n1476_0[0]),.dout(n1542),.clk(gclk));
	jor g1479(.dina(n1542),.dinb(w_dff_B_rlviRy9l5_1),.dout(n1543),.clk(gclk));
	jand g1480(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1544),.clk(gclk));
	jnot g1481(.din(n1544),.dout(n1545),.clk(gclk));
	jand g1482(.dina(w_n1513_0[0]),.dinb(w_n1484_0[0]),.dout(n1546),.clk(gclk));
	jand g1483(.dina(w_n1514_0[0]),.dinb(w_n1481_0[0]),.dout(n1547),.clk(gclk));
	jor g1484(.dina(n1547),.dinb(w_dff_B_16aT5zsN1_1),.dout(n1548),.clk(gclk));
	jand g1485(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1549),.clk(gclk));
	jnot g1486(.din(n1549),.dout(n1550),.clk(gclk));
	jand g1487(.dina(w_n1511_0[0]),.dinb(w_n1489_0[0]),.dout(n1551),.clk(gclk));
	jand g1488(.dina(w_n1512_0[0]),.dinb(w_n1486_0[0]),.dout(n1552),.clk(gclk));
	jor g1489(.dina(n1552),.dinb(w_dff_B_Q7YT2tXl2_1),.dout(n1553),.clk(gclk));
	jand g1490(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1554),.clk(gclk));
	jnot g1491(.din(n1554),.dout(n1555),.clk(gclk));
	jand g1492(.dina(w_n1509_0[0]),.dinb(w_n1494_0[0]),.dout(n1556),.clk(gclk));
	jand g1493(.dina(w_n1510_0[0]),.dinb(w_n1491_0[0]),.dout(n1557),.clk(gclk));
	jor g1494(.dina(n1557),.dinb(w_dff_B_C2oGLTtB5_1),.dout(n1558),.clk(gclk));
	jand g1495(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1559),.clk(gclk));
	jnot g1496(.din(n1559),.dout(n1560),.clk(gclk));
	jand g1497(.dina(w_n1507_0[0]),.dinb(w_n1499_0[0]),.dout(n1561),.clk(gclk));
	jand g1498(.dina(w_n1508_0[0]),.dinb(w_n1496_0[0]),.dout(n1562),.clk(gclk));
	jor g1499(.dina(n1562),.dinb(w_dff_B_eAljtyPM9_1),.dout(n1563),.clk(gclk));
	jand g1500(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1564),.clk(gclk));
	jand g1501(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1565),.clk(gclk));
	jor g1502(.dina(w_n1504_0[0]),.dinb(w_n1501_0[0]),.dout(n1566),.clk(gclk));
	jor g1503(.dina(w_n1506_0[0]),.dinb(w_n1500_0[0]),.dout(n1567),.clk(gclk));
	jand g1504(.dina(n1567),.dinb(w_dff_B_SlEBjpw15_1),.dout(n1568),.clk(gclk));
	jxor g1505(.dina(w_n1568_0[1]),.dinb(w_n1565_0[1]),.dout(n1569),.clk(gclk));
	jnot g1506(.din(n1569),.dout(n1570),.clk(gclk));
	jxor g1507(.dina(w_n1570_0[1]),.dinb(w_n1564_0[1]),.dout(n1571),.clk(gclk));
	jxor g1508(.dina(w_n1571_0[1]),.dinb(w_n1563_0[1]),.dout(n1572),.clk(gclk));
	jxor g1509(.dina(w_n1572_0[1]),.dinb(w_n1560_0[1]),.dout(n1573),.clk(gclk));
	jxor g1510(.dina(w_n1573_0[1]),.dinb(w_n1558_0[1]),.dout(n1574),.clk(gclk));
	jxor g1511(.dina(w_n1574_0[1]),.dinb(w_n1555_0[1]),.dout(n1575),.clk(gclk));
	jxor g1512(.dina(w_n1575_0[1]),.dinb(w_n1553_0[1]),.dout(n1576),.clk(gclk));
	jxor g1513(.dina(w_n1576_0[1]),.dinb(w_n1550_0[1]),.dout(n1577),.clk(gclk));
	jxor g1514(.dina(w_n1577_0[1]),.dinb(w_n1548_0[1]),.dout(n1578),.clk(gclk));
	jxor g1515(.dina(w_n1578_0[1]),.dinb(w_n1545_0[1]),.dout(n1579),.clk(gclk));
	jxor g1516(.dina(w_n1579_0[1]),.dinb(w_n1543_0[1]),.dout(n1580),.clk(gclk));
	jxor g1517(.dina(w_n1580_0[1]),.dinb(w_n1540_0[1]),.dout(n1581),.clk(gclk));
	jxor g1518(.dina(w_n1581_0[1]),.dinb(w_n1538_0[1]),.dout(n1582),.clk(gclk));
	jnot g1519(.din(n1582),.dout(n1583),.clk(gclk));
	jxor g1520(.dina(w_n1583_0[1]),.dinb(w_n1535_0[1]),.dout(n1584),.clk(gclk));
	jnot g1521(.din(n1584),.dout(n1585),.clk(gclk));
	jxor g1522(.dina(w_n1585_0[1]),.dinb(w_n1534_0[1]),.dout(n1586),.clk(gclk));
	jxor g1523(.dina(w_n1586_0[1]),.dinb(w_n1529_0[1]),.dout(w_dff_A_J9KkTH2x8_2),.clk(gclk));
	jor g1524(.dina(w_n1585_0[0]),.dinb(w_n1534_0[0]),.dout(n1588),.clk(gclk));
	jnot g1525(.din(w_n1586_0[0]),.dout(n1589),.clk(gclk));
	jor g1526(.dina(w_dff_B_NWY9YSYe7_0),.dinb(w_n1529_0[0]),.dout(n1590),.clk(gclk));
	jand g1527(.dina(n1590),.dinb(w_dff_B_8ztmIV7a7_1),.dout(n1591),.clk(gclk));
	jnot g1528(.din(w_n1538_0[0]),.dout(n1592),.clk(gclk));
	jnot g1529(.din(w_n1581_0[0]),.dout(n1593),.clk(gclk));
	jor g1530(.dina(w_dff_B_BVI7x5lT3_0),.dinb(n1592),.dout(n1594),.clk(gclk));
	jor g1531(.dina(w_n1583_0[0]),.dinb(w_n1535_0[0]),.dout(n1595),.clk(gclk));
	jand g1532(.dina(n1595),.dinb(w_dff_B_oYhPHKjl4_1),.dout(n1596),.clk(gclk));
	jand g1533(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1597),.clk(gclk));
	jand g1534(.dina(w_n1579_0[0]),.dinb(w_n1543_0[0]),.dout(n1598),.clk(gclk));
	jand g1535(.dina(w_n1580_0[0]),.dinb(w_n1540_0[0]),.dout(n1599),.clk(gclk));
	jor g1536(.dina(n1599),.dinb(w_dff_B_7wdXn7xq8_1),.dout(n1600),.clk(gclk));
	jand g1537(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1601),.clk(gclk));
	jnot g1538(.din(n1601),.dout(n1602),.clk(gclk));
	jand g1539(.dina(w_n1577_0[0]),.dinb(w_n1548_0[0]),.dout(n1603),.clk(gclk));
	jand g1540(.dina(w_n1578_0[0]),.dinb(w_n1545_0[0]),.dout(n1604),.clk(gclk));
	jor g1541(.dina(n1604),.dinb(w_dff_B_XFmAsQRz6_1),.dout(n1605),.clk(gclk));
	jand g1542(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1606),.clk(gclk));
	jnot g1543(.din(n1606),.dout(n1607),.clk(gclk));
	jand g1544(.dina(w_n1575_0[0]),.dinb(w_n1553_0[0]),.dout(n1608),.clk(gclk));
	jand g1545(.dina(w_n1576_0[0]),.dinb(w_n1550_0[0]),.dout(n1609),.clk(gclk));
	jor g1546(.dina(n1609),.dinb(w_dff_B_NToFGzAQ7_1),.dout(n1610),.clk(gclk));
	jand g1547(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1611),.clk(gclk));
	jnot g1548(.din(n1611),.dout(n1612),.clk(gclk));
	jand g1549(.dina(w_n1573_0[0]),.dinb(w_n1558_0[0]),.dout(n1613),.clk(gclk));
	jand g1550(.dina(w_n1574_0[0]),.dinb(w_n1555_0[0]),.dout(n1614),.clk(gclk));
	jor g1551(.dina(n1614),.dinb(w_dff_B_WCqwlkD57_1),.dout(n1615),.clk(gclk));
	jand g1552(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1616),.clk(gclk));
	jnot g1553(.din(n1616),.dout(n1617),.clk(gclk));
	jand g1554(.dina(w_n1571_0[0]),.dinb(w_n1563_0[0]),.dout(n1618),.clk(gclk));
	jand g1555(.dina(w_n1572_0[0]),.dinb(w_n1560_0[0]),.dout(n1619),.clk(gclk));
	jor g1556(.dina(n1619),.dinb(w_dff_B_LwpMB43I2_1),.dout(n1620),.clk(gclk));
	jand g1557(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1621),.clk(gclk));
	jand g1558(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1622),.clk(gclk));
	jor g1559(.dina(w_n1568_0[0]),.dinb(w_n1565_0[0]),.dout(n1623),.clk(gclk));
	jor g1560(.dina(w_n1570_0[0]),.dinb(w_n1564_0[0]),.dout(n1624),.clk(gclk));
	jand g1561(.dina(n1624),.dinb(w_dff_B_Hip9cB0c0_1),.dout(n1625),.clk(gclk));
	jxor g1562(.dina(w_n1625_0[1]),.dinb(w_n1622_0[1]),.dout(n1626),.clk(gclk));
	jnot g1563(.din(n1626),.dout(n1627),.clk(gclk));
	jxor g1564(.dina(w_n1627_0[1]),.dinb(w_n1621_0[1]),.dout(n1628),.clk(gclk));
	jxor g1565(.dina(w_n1628_0[1]),.dinb(w_n1620_0[1]),.dout(n1629),.clk(gclk));
	jxor g1566(.dina(w_n1629_0[1]),.dinb(w_n1617_0[1]),.dout(n1630),.clk(gclk));
	jxor g1567(.dina(w_n1630_0[1]),.dinb(w_n1615_0[1]),.dout(n1631),.clk(gclk));
	jxor g1568(.dina(w_n1631_0[1]),.dinb(w_n1612_0[1]),.dout(n1632),.clk(gclk));
	jxor g1569(.dina(w_n1632_0[1]),.dinb(w_n1610_0[1]),.dout(n1633),.clk(gclk));
	jxor g1570(.dina(w_n1633_0[1]),.dinb(w_n1607_0[1]),.dout(n1634),.clk(gclk));
	jxor g1571(.dina(w_n1634_0[1]),.dinb(w_n1605_0[1]),.dout(n1635),.clk(gclk));
	jxor g1572(.dina(w_n1635_0[1]),.dinb(w_n1602_0[1]),.dout(n1636),.clk(gclk));
	jxor g1573(.dina(w_n1636_0[1]),.dinb(w_n1600_0[1]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jxor g1575(.dina(w_n1638_0[1]),.dinb(w_n1597_0[1]),.dout(n1639),.clk(gclk));
	jnot g1576(.din(n1639),.dout(n1640),.clk(gclk));
	jxor g1577(.dina(w_n1640_0[1]),.dinb(w_n1596_0[1]),.dout(n1641),.clk(gclk));
	jxor g1578(.dina(w_n1641_0[1]),.dinb(w_n1591_0[1]),.dout(w_dff_A_SiAvJkIH2_2),.clk(gclk));
	jor g1579(.dina(w_n1640_0[0]),.dinb(w_n1596_0[0]),.dout(n1643),.clk(gclk));
	jnot g1580(.din(w_n1641_0[0]),.dout(n1644),.clk(gclk));
	jor g1581(.dina(w_dff_B_AIWOmTrF2_0),.dinb(w_n1591_0[0]),.dout(n1645),.clk(gclk));
	jand g1582(.dina(n1645),.dinb(w_dff_B_UBMYoQfe2_1),.dout(n1646),.clk(gclk));
	jnot g1583(.din(w_n1600_0[0]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(w_n1636_0[0]),.dout(n1648),.clk(gclk));
	jor g1585(.dina(n1648),.dinb(n1647),.dout(n1649),.clk(gclk));
	jor g1586(.dina(w_n1638_0[0]),.dinb(w_n1597_0[0]),.dout(n1650),.clk(gclk));
	jand g1587(.dina(n1650),.dinb(w_dff_B_fQdaedm32_1),.dout(n1651),.clk(gclk));
	jand g1588(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1652),.clk(gclk));
	jnot g1589(.din(n1652),.dout(n1653),.clk(gclk));
	jand g1590(.dina(w_n1634_0[0]),.dinb(w_n1605_0[0]),.dout(n1654),.clk(gclk));
	jand g1591(.dina(w_n1635_0[0]),.dinb(w_n1602_0[0]),.dout(n1655),.clk(gclk));
	jor g1592(.dina(n1655),.dinb(w_dff_B_t9D5uTt80_1),.dout(n1656),.clk(gclk));
	jand g1593(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jand g1595(.dina(w_n1632_0[0]),.dinb(w_n1610_0[0]),.dout(n1659),.clk(gclk));
	jand g1596(.dina(w_n1633_0[0]),.dinb(w_n1607_0[0]),.dout(n1660),.clk(gclk));
	jor g1597(.dina(n1660),.dinb(w_dff_B_J1dXw1Si3_1),.dout(n1661),.clk(gclk));
	jand g1598(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1662),.clk(gclk));
	jnot g1599(.din(n1662),.dout(n1663),.clk(gclk));
	jand g1600(.dina(w_n1630_0[0]),.dinb(w_n1615_0[0]),.dout(n1664),.clk(gclk));
	jand g1601(.dina(w_n1631_0[0]),.dinb(w_n1612_0[0]),.dout(n1665),.clk(gclk));
	jor g1602(.dina(n1665),.dinb(w_dff_B_Z3kybcKC3_1),.dout(n1666),.clk(gclk));
	jand g1603(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1667),.clk(gclk));
	jnot g1604(.din(n1667),.dout(n1668),.clk(gclk));
	jand g1605(.dina(w_n1628_0[0]),.dinb(w_n1620_0[0]),.dout(n1669),.clk(gclk));
	jand g1606(.dina(w_n1629_0[0]),.dinb(w_n1617_0[0]),.dout(n1670),.clk(gclk));
	jor g1607(.dina(n1670),.dinb(w_dff_B_df8nTyr38_1),.dout(n1671),.clk(gclk));
	jand g1608(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1672),.clk(gclk));
	jand g1609(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1673),.clk(gclk));
	jor g1610(.dina(w_n1625_0[0]),.dinb(w_n1622_0[0]),.dout(n1674),.clk(gclk));
	jor g1611(.dina(w_n1627_0[0]),.dinb(w_n1621_0[0]),.dout(n1675),.clk(gclk));
	jand g1612(.dina(n1675),.dinb(w_dff_B_O32QGbkt5_1),.dout(n1676),.clk(gclk));
	jxor g1613(.dina(w_n1676_0[1]),.dinb(w_n1673_0[1]),.dout(n1677),.clk(gclk));
	jnot g1614(.din(n1677),.dout(n1678),.clk(gclk));
	jxor g1615(.dina(w_n1678_0[1]),.dinb(w_n1672_0[1]),.dout(n1679),.clk(gclk));
	jxor g1616(.dina(w_n1679_0[1]),.dinb(w_n1671_0[1]),.dout(n1680),.clk(gclk));
	jxor g1617(.dina(w_n1680_0[1]),.dinb(w_n1668_0[1]),.dout(n1681),.clk(gclk));
	jxor g1618(.dina(w_n1681_0[1]),.dinb(w_n1666_0[1]),.dout(n1682),.clk(gclk));
	jxor g1619(.dina(w_n1682_0[1]),.dinb(w_n1663_0[1]),.dout(n1683),.clk(gclk));
	jxor g1620(.dina(w_n1683_0[1]),.dinb(w_n1661_0[1]),.dout(n1684),.clk(gclk));
	jxor g1621(.dina(w_n1684_0[1]),.dinb(w_n1658_0[1]),.dout(n1685),.clk(gclk));
	jxor g1622(.dina(w_n1685_0[1]),.dinb(w_n1656_0[1]),.dout(n1686),.clk(gclk));
	jxor g1623(.dina(w_n1686_0[1]),.dinb(w_n1653_0[1]),.dout(n1687),.clk(gclk));
	jnot g1624(.din(n1687),.dout(n1688),.clk(gclk));
	jxor g1625(.dina(w_n1688_0[1]),.dinb(w_n1651_0[1]),.dout(n1689),.clk(gclk));
	jxor g1626(.dina(w_n1689_0[1]),.dinb(w_n1646_0[1]),.dout(w_dff_A_iPOTMMlN8_2),.clk(gclk));
	jor g1627(.dina(w_n1688_0[0]),.dinb(w_n1651_0[0]),.dout(n1691),.clk(gclk));
	jnot g1628(.din(w_n1689_0[0]),.dout(n1692),.clk(gclk));
	jor g1629(.dina(w_dff_B_XuXI86Ur9_0),.dinb(w_n1646_0[0]),.dout(n1693),.clk(gclk));
	jand g1630(.dina(n1693),.dinb(w_dff_B_uLOxlXOx2_1),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1685_0[0]),.dinb(w_n1656_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1686_0[0]),.dinb(w_n1653_0[0]),.dout(n1696),.clk(gclk));
	jor g1633(.dina(n1696),.dinb(w_dff_B_l9V517vC0_1),.dout(n1697),.clk(gclk));
	jand g1634(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1683_0[0]),.dinb(w_n1661_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1684_0[0]),.dinb(w_n1658_0[0]),.dout(n1701),.clk(gclk));
	jor g1638(.dina(n1701),.dinb(w_dff_B_jjFo3b7d1_1),.dout(n1702),.clk(gclk));
	jand g1639(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1703),.clk(gclk));
	jnot g1640(.din(n1703),.dout(n1704),.clk(gclk));
	jand g1641(.dina(w_n1681_0[0]),.dinb(w_n1666_0[0]),.dout(n1705),.clk(gclk));
	jand g1642(.dina(w_n1682_0[0]),.dinb(w_n1663_0[0]),.dout(n1706),.clk(gclk));
	jor g1643(.dina(n1706),.dinb(w_dff_B_xUhWQ7P78_1),.dout(n1707),.clk(gclk));
	jand g1644(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jand g1646(.dina(w_n1679_0[0]),.dinb(w_n1671_0[0]),.dout(n1710),.clk(gclk));
	jand g1647(.dina(w_n1680_0[0]),.dinb(w_n1668_0[0]),.dout(n1711),.clk(gclk));
	jor g1648(.dina(n1711),.dinb(w_dff_B_SN63Z6ww0_1),.dout(n1712),.clk(gclk));
	jand g1649(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1713),.clk(gclk));
	jand g1650(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1714),.clk(gclk));
	jor g1651(.dina(w_n1676_0[0]),.dinb(w_n1673_0[0]),.dout(n1715),.clk(gclk));
	jor g1652(.dina(w_n1678_0[0]),.dinb(w_n1672_0[0]),.dout(n1716),.clk(gclk));
	jand g1653(.dina(n1716),.dinb(w_dff_B_lVWo6LPI0_1),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1714_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1713_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1712_0[1]),.dout(n1721),.clk(gclk));
	jxor g1658(.dina(w_n1721_0[1]),.dinb(w_n1709_0[1]),.dout(n1722),.clk(gclk));
	jxor g1659(.dina(w_n1722_0[1]),.dinb(w_n1707_0[1]),.dout(n1723),.clk(gclk));
	jxor g1660(.dina(w_n1723_0[1]),.dinb(w_n1704_0[1]),.dout(n1724),.clk(gclk));
	jxor g1661(.dina(w_n1724_0[1]),.dinb(w_n1702_0[1]),.dout(n1725),.clk(gclk));
	jxor g1662(.dina(w_n1725_0[1]),.dinb(w_n1699_0[1]),.dout(n1726),.clk(gclk));
	jxor g1663(.dina(w_n1726_0[1]),.dinb(w_n1697_0[1]),.dout(n1727),.clk(gclk));
	jxor g1664(.dina(w_n1727_0[1]),.dinb(w_n1694_0[1]),.dout(w_dff_A_ZynMqCJa0_2),.clk(gclk));
	jnot g1665(.din(w_n1697_0[0]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(w_n1726_0[0]),.dout(n1730),.clk(gclk));
	jor g1667(.dina(n1730),.dinb(w_dff_B_21KCN8U59_1),.dout(n1731),.clk(gclk));
	jnot g1668(.din(w_n1727_0[0]),.dout(n1732),.clk(gclk));
	jor g1669(.dina(w_dff_B_OqdGXR4B1_0),.dinb(w_n1694_0[0]),.dout(n1733),.clk(gclk));
	jand g1670(.dina(n1733),.dinb(w_dff_B_GZ6FuMXH6_1),.dout(n1734),.clk(gclk));
	jand g1671(.dina(w_n1724_0[0]),.dinb(w_n1702_0[0]),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1725_0[0]),.dinb(w_n1699_0[0]),.dout(n1736),.clk(gclk));
	jor g1673(.dina(n1736),.dinb(w_dff_B_FcTF5d0h3_1),.dout(n1737),.clk(gclk));
	jand g1674(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1738),.clk(gclk));
	jnot g1675(.din(n1738),.dout(n1739),.clk(gclk));
	jand g1676(.dina(w_n1722_0[0]),.dinb(w_n1707_0[0]),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1723_0[0]),.dinb(w_n1704_0[0]),.dout(n1741),.clk(gclk));
	jor g1678(.dina(n1741),.dinb(w_dff_B_IJm0KGB21_1),.dout(n1742),.clk(gclk));
	jand g1679(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1743),.clk(gclk));
	jnot g1680(.din(n1743),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_n1720_0[0]),.dinb(w_n1712_0[0]),.dout(n1745),.clk(gclk));
	jand g1682(.dina(w_n1721_0[0]),.dinb(w_n1709_0[0]),.dout(n1746),.clk(gclk));
	jor g1683(.dina(n1746),.dinb(w_dff_B_1cUf0YGg3_1),.dout(n1747),.clk(gclk));
	jand g1684(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1748),.clk(gclk));
	jand g1685(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1749),.clk(gclk));
	jor g1686(.dina(w_n1717_0[0]),.dinb(w_n1714_0[0]),.dout(n1750),.clk(gclk));
	jor g1687(.dina(w_n1719_0[0]),.dinb(w_n1713_0[0]),.dout(n1751),.clk(gclk));
	jand g1688(.dina(n1751),.dinb(w_dff_B_d4ZAE1QM3_1),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1749_0[1]),.dout(n1753),.clk(gclk));
	jnot g1690(.din(n1753),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1748_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1747_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1744_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1742_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1739_0[1]),.dout(n1759),.clk(gclk));
	jxor g1696(.dina(w_n1759_0[1]),.dinb(w_n1737_0[1]),.dout(n1760),.clk(gclk));
	jxor g1697(.dina(w_n1760_0[1]),.dinb(w_n1734_0[1]),.dout(w_dff_A_DQBFPbwp8_2),.clk(gclk));
	jnot g1698(.din(w_n1737_0[0]),.dout(n1762),.clk(gclk));
	jnot g1699(.din(w_n1759_0[0]),.dout(n1763),.clk(gclk));
	jor g1700(.dina(n1763),.dinb(w_dff_B_BKablcen2_1),.dout(n1764),.clk(gclk));
	jnot g1701(.din(w_n1760_0[0]),.dout(n1765),.clk(gclk));
	jor g1702(.dina(w_dff_B_S9IxMMvX1_0),.dinb(w_n1734_0[0]),.dout(n1766),.clk(gclk));
	jand g1703(.dina(n1766),.dinb(w_dff_B_vZrwHUxD9_1),.dout(n1767),.clk(gclk));
	jand g1704(.dina(w_n1757_0[0]),.dinb(w_n1742_0[0]),.dout(n1768),.clk(gclk));
	jand g1705(.dina(w_n1758_0[0]),.dinb(w_n1739_0[0]),.dout(n1769),.clk(gclk));
	jor g1706(.dina(n1769),.dinb(w_dff_B_OVSklzkW6_1),.dout(n1770),.clk(gclk));
	jand g1707(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1771),.clk(gclk));
	jnot g1708(.din(n1771),.dout(n1772),.clk(gclk));
	jand g1709(.dina(w_n1755_0[0]),.dinb(w_n1747_0[0]),.dout(n1773),.clk(gclk));
	jand g1710(.dina(w_n1756_0[0]),.dinb(w_n1744_0[0]),.dout(n1774),.clk(gclk));
	jor g1711(.dina(n1774),.dinb(w_dff_B_qWUxsDRZ7_1),.dout(n1775),.clk(gclk));
	jand g1712(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1777),.clk(gclk));
	jor g1714(.dina(w_n1752_0[0]),.dinb(w_n1749_0[0]),.dout(n1778),.clk(gclk));
	jor g1715(.dina(w_n1754_0[0]),.dinb(w_n1748_0[0]),.dout(n1779),.clk(gclk));
	jand g1716(.dina(n1779),.dinb(w_dff_B_RPpjFPI81_1),.dout(n1780),.clk(gclk));
	jxor g1717(.dina(w_n1780_0[1]),.dinb(w_n1777_0[1]),.dout(n1781),.clk(gclk));
	jnot g1718(.din(n1781),.dout(n1782),.clk(gclk));
	jxor g1719(.dina(w_n1782_0[1]),.dinb(w_n1776_0[1]),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1775_0[1]),.dout(n1784),.clk(gclk));
	jxor g1721(.dina(w_n1784_0[1]),.dinb(w_n1772_0[1]),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1770_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1767_0[1]),.dout(w_dff_A_6HD4c7010_2),.clk(gclk));
	jnot g1724(.din(w_n1770_0[0]),.dout(n1788),.clk(gclk));
	jnot g1725(.din(w_n1785_0[0]),.dout(n1789),.clk(gclk));
	jor g1726(.dina(n1789),.dinb(w_dff_B_gTft9evD3_1),.dout(n1790),.clk(gclk));
	jnot g1727(.din(w_n1786_0[0]),.dout(n1791),.clk(gclk));
	jor g1728(.dina(w_dff_B_Eax2j83u3_0),.dinb(w_n1767_0[0]),.dout(n1792),.clk(gclk));
	jand g1729(.dina(n1792),.dinb(w_dff_B_IpFzrpKs7_1),.dout(n1793),.clk(gclk));
	jand g1730(.dina(w_n1783_0[0]),.dinb(w_n1775_0[0]),.dout(n1794),.clk(gclk));
	jand g1731(.dina(w_n1784_0[0]),.dinb(w_n1772_0[0]),.dout(n1795),.clk(gclk));
	jor g1732(.dina(n1795),.dinb(w_dff_B_85yW5gdO3_1),.dout(n1796),.clk(gclk));
	jand g1733(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1797),.clk(gclk));
	jand g1734(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1798),.clk(gclk));
	jor g1735(.dina(w_n1780_0[0]),.dinb(w_n1777_0[0]),.dout(n1799),.clk(gclk));
	jor g1736(.dina(w_n1782_0[0]),.dinb(w_n1776_0[0]),.dout(n1800),.clk(gclk));
	jand g1737(.dina(n1800),.dinb(w_dff_B_qoKI2Mw54_1),.dout(n1801),.clk(gclk));
	jxor g1738(.dina(w_n1801_0[1]),.dinb(w_n1798_0[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jxor g1740(.dina(w_n1803_0[1]),.dinb(w_n1797_0[1]),.dout(n1804),.clk(gclk));
	jxor g1741(.dina(w_n1804_0[1]),.dinb(w_n1796_0[1]),.dout(n1805),.clk(gclk));
	jxor g1742(.dina(w_n1805_0[1]),.dinb(w_n1793_0[1]),.dout(w_dff_A_onIovUsr0_2),.clk(gclk));
	jand g1743(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1807),.clk(gclk));
	jor g1744(.dina(w_n1801_0[0]),.dinb(w_n1798_0[0]),.dout(n1808),.clk(gclk));
	jor g1745(.dina(w_n1803_0[0]),.dinb(w_n1797_0[0]),.dout(n1809),.clk(gclk));
	jand g1746(.dina(n1809),.dinb(w_dff_B_iEasrwnB9_1),.dout(n1810),.clk(gclk));
	jor g1747(.dina(w_n1810_0[1]),.dinb(w_n1807_0[1]),.dout(n1811),.clk(gclk));
	jnot g1748(.din(w_n1796_0[0]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(w_n1804_0[0]),.dout(n1813),.clk(gclk));
	jor g1750(.dina(n1813),.dinb(w_dff_B_rnOokL9a0_1),.dout(n1814),.clk(gclk));
	jnot g1751(.din(w_n1805_0[0]),.dout(n1815),.clk(gclk));
	jor g1752(.dina(w_dff_B_Zgspq9E55_0),.dinb(w_n1793_0[0]),.dout(n1816),.clk(gclk));
	jand g1753(.dina(n1816),.dinb(w_dff_B_c6XrcEjR7_1),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1810_0[0]),.dinb(w_n1807_0[0]),.dout(n1818),.clk(gclk));
	jnot g1755(.din(w_n1818_0[1]),.dout(n1819),.clk(gclk));
	jor g1756(.dina(w_dff_B_JaAxITgE4_0),.dinb(w_n1817_0[1]),.dout(n1820),.clk(gclk));
	jand g1757(.dina(n1820),.dinb(w_dff_B_DRCwA28l1_1),.dout(G6287gat),.clk(gclk));
	jxor g1758(.dina(w_n1818_0[0]),.dinb(w_n1817_0[0]),.dout(w_dff_A_mVaqxWQK4_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl jspl_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl jspl_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_G307gat_2[1]),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl jspl_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(w_dff_A_Fe3KFXMD4_1),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n66_0(.douta(w_dff_A_UFSzZaHP3_0),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(w_dff_B_2dDyRXUu5_2));
	jspl jspl_w_n69_0(.douta(w_n69_0[0]),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n75_0(.douta(w_dff_A_fEHBPXtO2_0),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl3 jspl3_w_n80_0(.douta(w_dff_A_4Cr04xW87_0),.doutb(w_n80_0[1]),.doutc(w_n80_0[2]),.din(n80));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_dff_A_zLcH8Jq08_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_dff_A_LooSY29h1_0),.doutb(w_n91_0[1]),.din(n91));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_DRCi3GWz7_1),.din(n103));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n106_0(.douta(w_dff_A_qKRfbRCj6_0),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl jspl_w_n112_0(.douta(w_dff_A_7Mzcdqd21_0),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(w_dff_B_WUu4GHNc7_2));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n122_0(.douta(w_dff_A_dYnoKGBq0_0),.doutb(w_n122_0[1]),.din(n122));
	jspl jspl_w_n123_0(.douta(w_dff_A_2DFVxxTq9_0),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n129_0(.douta(w_dff_A_HGFBKBQc8_0),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.din(n130));
	jspl jspl_w_n132_0(.douta(w_n132_0[0]),.doutb(w_dff_A_Hwo7FDkD5_1),.din(n132));
	jspl jspl_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.din(n133));
	jspl jspl_w_n135_0(.douta(w_dff_A_Kob3NXpf4_0),.doutb(w_n135_0[1]),.din(n135));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n141_0(.douta(w_dff_A_cKR98tgH2_0),.doutb(w_n141_0[1]),.din(n141));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.doutc(w_n146_0[2]),.din(n146));
	jspl jspl_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.din(w_dff_B_7T33LGME5_2));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(w_dff_B_ICAcvj6l7_2));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_dff_A_DABRaDyw5_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n157_0(.douta(w_dff_A_e5uR1iD21_0),.doutb(w_n157_0[1]),.din(n157));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(n158));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl jspl_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(w_dff_B_My0VlJMI7_2));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n164_0(.douta(w_dff_A_kFA4SIdY6_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(n165));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_dff_A_MTOSucTE3_1),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl jspl_w_n170_0(.douta(w_dff_A_qGBbdJg55_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n176_0(.douta(w_dff_A_NRNMucvL8_0),.doutb(w_n176_0[1]),.din(n176));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl jspl_w_n183_0(.douta(w_n183_0[0]),.doutb(w_n183_0[1]),.din(w_dff_B_zjj0zFqA2_2));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(w_dff_B_kLH7gl653_2));
	jspl jspl_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.din(n192));
	jspl jspl_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.din(w_dff_B_HzLkcPRY1_2));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_dff_A_d0yTcVi09_0),.doutb(w_dff_A_Pm0Nd7zt9_1),.doutc(w_n196_0[2]),.din(n196));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(w_dff_B_k8KuEIIu9_2));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(n203));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(w_dff_B_OTekOYmC2_2));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n206_0(.douta(w_dff_A_w4z6xIvG0_0),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_dff_A_uD5kYzFY7_1),.din(n209));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_dff_A_hTpwivnN8_0),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_dff_A_f6h1wyU90_0),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.doutc(w_n223_0[2]),.din(n223));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(w_dff_B_7od6T22O2_2));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.din(w_dff_B_dQEcMFM43_2));
	jspl jspl_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.din(n233));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_n235_0[1]),.din(w_dff_B_r5l3dFb60_2));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(n239));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(w_dff_B_moe5ArhA2_2));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_dff_A_wPraWFFy9_0),.doutb(w_dff_A_VyoFlOGM9_1),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n248_0(.douta(w_n248_0[0]),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_F4vWvT7A0_2));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.din(w_dff_B_VFWvjV9t5_2));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.din(w_dff_B_gHhvR5im2_2));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n255_0(.douta(w_dff_A_Mw4tBpp83_0),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n256_0(.douta(w_n256_0[0]),.doutb(w_n256_0[1]),.din(n256));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_dff_A_T4cDbbGE9_1),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_dff_A_xFr8Ne6S7_0),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_dff_A_Ob6ywave7_0),.doutb(w_n267_0[1]),.din(n267));
	jspl3 jspl3_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.doutc(w_n272_0[2]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(w_dff_B_4xzSKqT53_2));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(w_dff_B_czwAcrTA5_2));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n284_0(.douta(w_n284_0[0]),.doutb(w_n284_0[1]),.din(w_dff_B_KI3bghAP8_2));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl jspl_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.din(w_dff_B_nzEs7aAK5_2));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(w_dff_B_xGVVmCvC2_2));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl3 jspl3_w_n297_0(.douta(w_dff_A_ErpNfXoR8_0),.doutb(w_dff_A_dAKuKW9I4_1),.doutc(w_n297_0[2]),.din(n297));
	jspl jspl_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.din(n299));
	jspl jspl_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.din(n301));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_n302_0[1]),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(w_dff_B_9ig1YyJM9_2));
	jspl jspl_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.din(n304));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(w_dff_B_SUc5WIUE5_2));
	jspl jspl_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.din(n306));
	jspl jspl_w_n307_0(.douta(w_n307_0[0]),.doutb(w_n307_0[1]),.din(w_dff_B_Xt3SxkYc6_2));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(w_dff_B_O5DfBWIa0_2));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(n310));
	jspl jspl_w_n311_0(.douta(w_dff_A_WKLMPdYf9_0),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.din(n312));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_dff_A_iki1Wsv18_1),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_dff_A_bZ4o1eNL3_0),.doutb(w_n317_0[1]),.din(n317));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_dff_A_RqtKQE7V3_0),.doutb(w_n323_0[1]),.din(n323));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(w_dff_B_y67DCB5M1_2));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.din(w_dff_B_Nzc0jN0X6_2));
	jspl jspl_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.din(n338));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(w_dff_B_980k4pLA3_2));
	jspl jspl_w_n343_0(.douta(w_n343_0[0]),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(w_dff_B_UKDO5yzq0_2));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(w_dff_B_pKLuxngU2_2));
	jspl jspl_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.din(n354));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(w_dff_B_a8u7jpK85_2));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl3 jspl3_w_n358_0(.douta(w_dff_A_PN5thRrM1_0),.doutb(w_dff_A_iBKlWHFh0_1),.doutc(w_n358_0[2]),.din(n358));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(n363));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(w_dff_B_v1WaF1H94_2));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(w_dff_B_o71vjIz19_2));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(w_dff_B_AhFWDYpV0_2));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(w_dff_B_ytpEQb7Q7_2));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(w_dff_B_QEgq628n1_2));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n374_0(.douta(w_dff_A_CDV3PFhs0_0),.doutb(w_n374_0[1]),.din(n374));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_dff_A_UNh2eDPN7_1),.din(n377));
	jspl jspl_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.din(n378));
	jspl jspl_w_n380_0(.douta(w_dff_A_d3MCYPN24_0),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl jspl_w_n386_0(.douta(w_dff_A_tCowXLRu0_0),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.doutc(w_n391_0[2]),.din(n391));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(w_dff_B_ZCDYx5Hp6_2));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.din(n396));
	jspl jspl_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.din(w_dff_B_80hrZBpf0_2));
	jspl jspl_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.din(n401));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(w_dff_B_546d4bqi9_2));
	jspl jspl_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.din(n406));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(w_dff_B_h9fjyNnY5_2));
	jspl jspl_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.din(n411));
	jspl jspl_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.din(w_dff_B_jOYZKkVE5_2));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(w_dff_B_WbZgNx2W0_2));
	jspl jspl_w_n418_0(.douta(w_n418_0[0]),.doutb(w_n418_0[1]),.din(w_dff_B_CuSaWmlk0_2));
	jspl jspl_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.din(n423));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(w_dff_B_QGJTPq0i6_2));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl3 jspl3_w_n427_0(.douta(w_dff_A_pOvWQzFu1_0),.doutb(w_dff_A_KrIQk1Yq0_1),.doutc(w_n427_0[2]),.din(n427));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl jspl_w_n431_0(.douta(w_n431_0[0]),.doutb(w_n431_0[1]),.din(n431));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(n432));
	jspl jspl_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.din(w_dff_B_zrQ40S7o4_2));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl jspl_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.din(n436));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl jspl_w_n438_0(.douta(w_n438_0[0]),.doutb(w_n438_0[1]),.din(n438));
	jspl jspl_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.din(w_dff_B_1pHowUne4_2));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(w_dff_B_Dr1IrqGm8_2));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_n442_0[1]),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(w_dff_B_VAUq4dSN9_2));
	jspl jspl_w_n444_0(.douta(w_n444_0[0]),.doutb(w_n444_0[1]),.din(n444));
	jspl jspl_w_n445_0(.douta(w_dff_A_pU4uyEYh8_0),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_dff_A_CXCuRGa09_1),.din(n448));
	jspl jspl_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.din(n449));
	jspl jspl_w_n451_0(.douta(w_dff_A_YkPo2Xyi0_0),.doutb(w_n451_0[1]),.din(n451));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_dff_A_qmqeJ4rw5_0),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(w_dff_B_w7W1k9Hk6_2));
	jspl jspl_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.din(n467));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(w_dff_B_v1qq48ab4_2));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(w_dff_B_mnwGxLnu0_2));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(w_dff_B_74u6g0wf4_2));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(w_dff_B_hnVkheOv4_2));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(w_dff_B_dTMigAAZ6_2));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(w_dff_B_sW1vra5Q7_2));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(n499));
	jspl jspl_w_n501_0(.douta(w_n501_0[0]),.doutb(w_n501_0[1]),.din(w_dff_B_a9yMZg6v9_2));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl3 jspl3_w_n503_0(.douta(w_dff_A_t6iX48tA8_0),.doutb(w_dff_A_qZksD9iJ4_1),.doutc(w_n503_0[2]),.din(n503));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_bSzKJyA47_2));
	jspl jspl_w_n510_0(.douta(w_n510_0[0]),.doutb(w_n510_0[1]),.din(n510));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(w_dff_B_p2ZwLPy27_2));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.din(n513));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n515_0(.douta(w_n515_0[0]),.doutb(w_n515_0[1]),.din(n515));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(w_dff_B_zuvg0Oqv6_2));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(w_dff_B_pYAEP80p8_2));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n521_0(.douta(w_n521_0[0]),.doutb(w_n521_0[1]),.din(w_dff_B_hZo4AJL16_2));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl jspl_w_n523_0(.douta(w_dff_A_fQs3s16e9_0),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n526_0(.douta(w_n526_0[0]),.doutb(w_dff_A_SLB4Z28D3_1),.din(n526));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_dff_A_mEqOSiLQ7_0),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_dff_A_fKn3qFcf1_0),.doutb(w_n535_0[1]),.din(n535));
	jspl3 jspl3_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.doutc(w_n540_0[2]),.din(n540));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(w_dff_B_eR3Wb2sf5_2));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(w_dff_B_jw7L1Y4g3_2));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(w_dff_B_5X81MMu62_2));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(w_dff_B_PIUi5LCX0_2));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(w_dff_B_NAIXv9WN7_2));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(w_dff_B_yETXfUWg6_2));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl jspl_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.din(w_dff_B_Bw3OsVie8_2));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(w_dff_B_okQQNJjO8_2));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(w_dff_B_t8ZJcDmB0_2));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n586_0(.douta(w_dff_A_lI9Tl6Ax2_0),.doutb(w_dff_A_SA268giF4_1),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(n588));
	jspl jspl_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.din(n590));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(w_dff_B_rD2axpKL5_2));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl jspl_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.din(w_dff_B_iknV8gPt0_2));
	jspl jspl_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.din(n595));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(w_dff_B_Kuevk1gs9_2));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl jspl_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.din(n599));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(n600));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(w_dff_B_BwJipq5t9_2));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(w_dff_B_fSPB99zU8_2));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(w_dff_B_Q4Xb684L2_2));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_dff_A_u6y9dCsG3_0),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.din(n609));
	jspl jspl_w_n611_0(.douta(w_n611_0[0]),.doutb(w_dff_A_ISeNVaNj6_1),.din(n611));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl jspl_w_n614_0(.douta(w_dff_A_CEOAP1Il9_0),.doutb(w_n614_0[1]),.din(n614));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_dff_A_tq7qiosp1_0),.doutb(w_n620_0[1]),.din(n620));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(w_dff_B_l80K2F2M7_2));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(w_dff_B_XIPQYJju6_2));
	jspl jspl_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.din(n635));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(w_dff_B_7cQ7JSZV7_2));
	jspl jspl_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.din(n640));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(w_dff_B_2KqAnSEU2_2));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(w_dff_B_cbKJmi6f7_2));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(w_dff_B_1d86I5RD5_2));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(w_dff_B_yuiA1Rrp4_2));
	jspl jspl_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.din(n660));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(w_dff_B_yvjjMG5t8_2));
	jspl jspl_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.din(n665));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(w_dff_B_NcfWduB29_2));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(w_dff_B_ymoeGeBM1_2));
	jspl jspl_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.din(n675));
	jspl3 jspl3_w_n676_0(.douta(w_dff_A_ddDRVV2g5_0),.doutb(w_dff_A_u7HtRnIt1_1),.doutc(w_n676_0[2]),.din(n676));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl jspl_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.din(n681));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(w_dff_B_NnRZQt6k9_2));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(w_dff_B_ntkPcTrO9_2));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(w_dff_B_d8eQmLZH6_2));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n688_0(.douta(w_n688_0[0]),.doutb(w_n688_0[1]),.din(w_dff_B_1w0Q7Pzv5_2));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.din(n691));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.din(n692));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.din(w_dff_B_esxJIrZt0_2));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.din(w_dff_B_9bFez3Sf8_2));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(w_dff_B_mZTqKZKU0_2));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n700_0(.douta(w_dff_A_0YxJ5nxx6_0),.doutb(w_n700_0[1]),.din(n700));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_dff_A_WtcaqWte1_1),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n706_0(.douta(w_dff_A_N18EMJBx6_0),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_dff_A_4ptKqsnL1_0),.doutb(w_n712_0[1]),.din(n712));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.doutc(w_n717_0[2]),.din(n717));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(w_dff_B_iI69Sy724_2));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(w_dff_B_slip2qC92_2));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.din(w_dff_B_FhOXP8Hs1_2));
	jspl jspl_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.din(n732));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(w_dff_B_bTlMXmHN0_2));
	jspl jspl_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.din(n737));
	jspl jspl_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.din(w_dff_B_DgxOZg6R1_2));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl jspl_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.din(w_dff_B_VA0c2Vd83_2));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(n747));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(w_dff_B_28pqL9by1_2));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(w_dff_B_6HXXvmvm1_2));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(w_dff_B_XovSSTRy2_2));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(n762));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(w_dff_B_EXRxjeOL2_2));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(w_dff_B_x2wZXyLI6_2));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.din(n774));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.din(w_dff_B_px5urLfF6_2));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.din(w_dff_B_1s3Leg2W0_2));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.din(w_dff_B_v1rhBZ8R9_2));
	jspl jspl_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.din(n784));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(w_dff_B_cF7Ixm6x1_2));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_iedO2Yhv8_2));
	jspl jspl_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.din(n788));
	jspl jspl_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.din(n789));
	jspl jspl_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.din(n790));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl jspl_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.din(w_dff_B_hscgPvLM9_2));
	jspl jspl_w_n794_0(.douta(w_n794_0[0]),.doutb(w_n794_0[1]),.din(n794));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(w_dff_B_AOXHx3Iw7_2));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl jspl_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.din(w_dff_B_jkAymBlt3_2));
	jspl jspl_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.din(n798));
	jspl jspl_w_n799_0(.douta(w_dff_A_S6FwpfXP2_0),.doutb(w_n799_0[1]),.din(n799));
	jspl jspl_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_dff_A_eo9lZxUw1_1),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(n803));
	jspl jspl_w_n805_0(.douta(w_dff_A_QqOo8jfq1_0),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(w_dff_B_jdynKIxI1_2));
	jspl jspl_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_dff_A_0TE8lFqx1_0),.doutb(w_n816_0[1]),.din(n816));
	jspl3 jspl3_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.doutc(w_n820_0[2]),.din(n820));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(w_dff_B_4qzbGwQl1_2));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(w_dff_B_GT7w1IgP9_2));
	jspl jspl_w_n830_0(.douta(w_n830_0[0]),.doutb(w_n830_0[1]),.din(n830));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(w_dff_B_1e5eJ58E4_2));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl jspl_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.din(w_dff_B_UyzY5MlU4_2));
	jspl jspl_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.din(n840));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(w_dff_B_cKWKrVXj8_2));
	jspl jspl_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.din(n845));
	jspl jspl_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.din(w_dff_B_xWjgITBo3_2));
	jspl jspl_w_n850_0(.douta(w_n850_0[0]),.doutb(w_n850_0[1]),.din(n850));
	jspl jspl_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.din(w_dff_B_lOI0ErTq6_2));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(w_dff_B_6GItylHC3_2));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(w_dff_B_wSkPVZ5H8_2));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(w_dff_B_AxdmzWHQ1_2));
	jspl jspl_w_n872_0(.douta(w_n872_0[0]),.doutb(w_n872_0[1]),.din(n872));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(w_dff_B_sHzh34fk5_2));
	jspl jspl_w_n875_0(.douta(w_dff_A_U3lV2lY70_0),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n877_0(.douta(w_dff_A_nVhSQM5i0_0),.doutb(w_n877_0[1]),.din(w_dff_B_91FhsFt05_2));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.din(w_dff_B_P00s8lh91_2));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n882_0(.douta(w_n882_0[0]),.doutb(w_n882_0[1]),.din(w_dff_B_R921Ezfz5_2));
	jspl jspl_w_n883_0(.douta(w_n883_0[0]),.doutb(w_n883_0[1]),.din(n883));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(w_dff_B_Wvs81bCN0_2));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(w_dff_B_e8521bL50_2));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.din(n887));
	jspl jspl_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.din(w_dff_B_YkoF4SCv4_2));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(w_dff_B_V85fjSlv9_2));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(n891));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n893_0(.douta(w_n893_0[0]),.doutb(w_n893_0[1]),.din(n893));
	jspl jspl_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(w_dff_B_3oDfo5a12_2));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(w_dff_B_UXHgDEAd7_2));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.din(n899));
	jspl3 jspl3_w_n900_0(.douta(w_n900_0[0]),.doutb(w_dff_A_l6lgNt926_1),.doutc(w_dff_A_fTqCUQNZ9_2),.din(n900));
	jspl jspl_w_n902_0(.douta(w_n902_0[0]),.doutb(w_dff_A_0J86BOMG3_1),.din(n902));
	jspl jspl_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n904_0(.douta(w_n904_0[0]),.doutb(w_dff_A_7cq0XO5c0_1),.din(n904));
	jspl jspl_w_n905_0(.douta(w_n905_0[0]),.doutb(w_n905_0[1]),.din(n905));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(n910));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(w_dff_B_uqtKeENz7_2));
	jspl3 jspl3_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.doutc(w_n915_0[2]),.din(n915));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(w_dff_B_sNYQT0OB0_2));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(w_dff_B_xChHUj2Q5_2));
	jspl jspl_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(w_dff_B_XIQ0wdDi2_2));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n934_0(.douta(w_n934_0[0]),.doutb(w_n934_0[1]),.din(w_dff_B_GETyUF4i3_2));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n939_0(.douta(w_n939_0[0]),.doutb(w_n939_0[1]),.din(w_dff_B_APlCJvM38_2));
	jspl jspl_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.din(n942));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(w_dff_B_ZaSiZtFw1_2));
	jspl jspl_w_n947_0(.douta(w_n947_0[0]),.doutb(w_n947_0[1]),.din(n947));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(w_dff_B_2WUixItf6_2));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(w_dff_B_rYhzUowM4_2));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(w_dff_B_7uNOedha2_2));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(w_dff_B_GpUGpCoU0_2));
	jspl jspl_w_n967_0(.douta(w_n967_0[0]),.doutb(w_n967_0[1]),.din(n967));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(w_dff_B_4ShqpVAq3_2));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(w_dff_B_c4z6oQvR5_2));
	jspl jspl_w_n978_0(.douta(w_n978_0[0]),.doutb(w_n978_0[1]),.din(n978));
	jspl jspl_w_n980_0(.douta(w_dff_A_cTYpb9Uc5_0),.doutb(w_n980_0[1]),.din(w_dff_B_0eI2STGI0_2));
	jspl jspl_w_n982_0(.douta(w_n982_0[0]),.doutb(w_n982_0[1]),.din(n982));
	jspl jspl_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.din(w_dff_B_gu26uhNi2_2));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(w_dff_B_1PruDQuf8_2));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(w_dff_B_5E2IGDSn9_2));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl jspl_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.din(w_dff_B_FFyMfjKa9_2));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.din(w_dff_B_UZquPyqL3_2));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(w_dff_B_yMyjy5lP9_2));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(w_dff_B_EqvHgSLD6_2));
	jspl jspl_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.din(n995));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(w_dff_B_hYJzon4O3_2));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl jspl_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.din(w_dff_B_hPP1DsNg0_2));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.din(w_dff_B_ETjCxcFW4_2));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_dff_A_Ig2IiMIV7_1),.din(n1006));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_dff_A_SJbKKdsT3_0),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(w_dff_B_CVkOlKTy6_2));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_dff_A_jiOGZly09_1),.din(n1013));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(w_dff_B_GkYwjBE79_2));
	jspl jspl_w_n1022_0(.douta(w_dff_A_pgxmyIZO4_0),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(w_dff_B_IcKyzXsc3_2));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(w_dff_B_yCfDalDw2_2));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(w_dff_B_JxLDU3Sf6_2));
	jspl jspl_w_n1036_0(.douta(w_n1036_0[0]),.doutb(w_n1036_0[1]),.din(n1036));
	jspl jspl_w_n1038_0(.douta(w_n1038_0[0]),.doutb(w_n1038_0[1]),.din(w_dff_B_x2SPxzy90_2));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(w_dff_B_0et19v5d5_2));
	jspl jspl_w_n1046_0(.douta(w_n1046_0[0]),.doutb(w_n1046_0[1]),.din(n1046));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(w_dff_B_CSNfWwZN2_2));
	jspl jspl_w_n1051_0(.douta(w_n1051_0[0]),.doutb(w_n1051_0[1]),.din(n1051));
	jspl jspl_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.din(w_dff_B_M6F2BNcO5_2));
	jspl jspl_w_n1056_0(.douta(w_n1056_0[0]),.doutb(w_n1056_0[1]),.din(n1056));
	jspl jspl_w_n1058_0(.douta(w_n1058_0[0]),.doutb(w_n1058_0[1]),.din(w_dff_B_7FGqqgOK4_2));
	jspl jspl_w_n1061_0(.douta(w_n1061_0[0]),.doutb(w_n1061_0[1]),.din(n1061));
	jspl jspl_w_n1063_0(.douta(w_n1063_0[0]),.doutb(w_n1063_0[1]),.din(w_dff_B_UBQUdD8G3_2));
	jspl jspl_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.din(n1066));
	jspl jspl_w_n1068_0(.douta(w_n1068_0[0]),.doutb(w_n1068_0[1]),.din(w_dff_B_VfNDgjQa5_2));
	jspl jspl_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.din(n1071));
	jspl jspl_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.din(w_dff_B_vR19TmIW5_2));
	jspl jspl_w_n1076_0(.douta(w_n1076_0[0]),.doutb(w_n1076_0[1]),.din(n1076));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(w_dff_B_x50Fva0C5_2));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(w_dff_B_s8ukJ44q7_2));
	jspl jspl_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.din(n1080));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl jspl_w_n1083_0(.douta(w_n1083_0[0]),.doutb(w_n1083_0[1]),.din(w_dff_B_QBuWzmQu0_2));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(n1084));
	jspl jspl_w_n1085_0(.douta(w_n1085_0[0]),.doutb(w_n1085_0[1]),.din(w_dff_B_bFThtfdB8_2));
	jspl jspl_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.din(n1086));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(w_dff_B_9dj6N0cZ0_2));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(w_dff_B_MV1nrUwB4_2));
	jspl jspl_w_n1090_0(.douta(w_n1090_0[0]),.doutb(w_n1090_0[1]),.din(n1090));
	jspl jspl_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.din(w_dff_B_oht5QqZp1_2));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1093_0(.douta(w_n1093_0[0]),.doutb(w_n1093_0[1]),.din(w_dff_B_pravOeJa6_2));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(n1094));
	jspl jspl_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.din(w_dff_B_SmpoGJ4N8_2));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1098_0(.douta(w_n1098_0[0]),.doutb(w_n1098_0[1]),.din(n1098));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1100_0(.douta(w_n1100_0[0]),.doutb(w_n1100_0[1]),.din(n1100));
	jspl jspl_w_n1101_0(.douta(w_n1101_0[0]),.doutb(w_n1101_0[1]),.din(w_dff_B_bXXrmGpH8_2));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(w_dff_B_LOO3qfnl6_2));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.din(n1105));
	jspl jspl_w_n1106_0(.douta(w_n1106_0[0]),.doutb(w_n1106_0[1]),.din(n1106));
	jspl jspl_w_n1107_0(.douta(w_n1107_0[0]),.doutb(w_n1107_0[1]),.din(n1107));
	jspl jspl_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_dff_A_yNR5ZAP00_1),.din(n1108));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1119_0(.douta(w_dff_A_oD3ElxP60_0),.doutb(w_n1119_0[1]),.din(w_dff_B_Bbcq3lRP1_2));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(w_dff_B_N6CcgjhU8_2));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(w_dff_B_CofvUyBV3_2));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(w_dff_B_3asv6Oq43_2));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1136_0(.douta(w_n1136_0[0]),.doutb(w_n1136_0[1]),.din(w_dff_B_O7NpO5ou1_2));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(w_dff_B_kuIpC0Vp4_2));
	jspl jspl_w_n1144_0(.douta(w_n1144_0[0]),.doutb(w_n1144_0[1]),.din(n1144));
	jspl jspl_w_n1146_0(.douta(w_n1146_0[0]),.doutb(w_n1146_0[1]),.din(w_dff_B_WHme5axn2_2));
	jspl jspl_w_n1149_0(.douta(w_n1149_0[0]),.doutb(w_n1149_0[1]),.din(n1149));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(w_dff_B_DANe89Pc6_2));
	jspl jspl_w_n1154_0(.douta(w_n1154_0[0]),.doutb(w_n1154_0[1]),.din(n1154));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(w_dff_B_04xkvR896_2));
	jspl jspl_w_n1159_0(.douta(w_n1159_0[0]),.doutb(w_n1159_0[1]),.din(n1159));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(w_dff_B_2uCsVlcn6_2));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(n1164));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(w_dff_B_0fgYsl7M7_2));
	jspl jspl_w_n1169_0(.douta(w_n1169_0[0]),.doutb(w_n1169_0[1]),.din(n1169));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(w_dff_B_gsC6wqNH0_2));
	jspl jspl_w_n1174_0(.douta(w_n1174_0[0]),.doutb(w_n1174_0[1]),.din(n1174));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_n1175_0[1]),.din(w_dff_B_3iHvH29H0_2));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(w_dff_B_bHlhii1X8_2));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1182_0(.douta(w_n1182_0[0]),.doutb(w_n1182_0[1]),.din(w_dff_B_l1BIsj2K7_2));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.din(w_dff_B_FbDURwN55_2));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(w_dff_B_p4KQoNjV9_2));
	jspl jspl_w_n1187_0(.douta(w_n1187_0[0]),.doutb(w_n1187_0[1]),.din(n1187));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(w_dff_B_y33tYOu80_2));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1190_0(.douta(w_n1190_0[0]),.doutb(w_n1190_0[1]),.din(w_dff_B_LVaaCOzx9_2));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(n1191));
	jspl jspl_w_n1192_0(.douta(w_n1192_0[0]),.doutb(w_n1192_0[1]),.din(w_dff_B_8UoqdxrN9_2));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(n1193));
	jspl jspl_w_n1194_0(.douta(w_n1194_0[0]),.doutb(w_n1194_0[1]),.din(w_dff_B_D3YZD5D76_2));
	jspl jspl_w_n1195_0(.douta(w_n1195_0[0]),.doutb(w_n1195_0[1]),.din(n1195));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.din(n1197));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(n1198));
	jspl jspl_w_n1199_0(.douta(w_n1199_0[0]),.doutb(w_n1199_0[1]),.din(n1199));
	jspl jspl_w_n1200_0(.douta(w_n1200_0[0]),.doutb(w_n1200_0[1]),.din(w_dff_B_aV33VNxI7_2));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(w_dff_B_g5qSM25j2_2));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(n1206));
	jspl jspl_w_n1207_0(.douta(w_dff_A_kaFjA6Cr4_0),.doutb(w_n1207_0[1]),.din(n1207));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(w_dff_B_plw1eKCA3_2));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(w_dff_B_xDLoDmzC7_2));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(n1225));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(w_dff_B_2TijpYi78_2));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(w_dff_B_PCF5qNEU6_2));
	jspl jspl_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.din(n1235));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(w_dff_B_okKF1GY07_2));
	jspl jspl_w_n1240_0(.douta(w_n1240_0[0]),.doutb(w_n1240_0[1]),.din(n1240));
	jspl jspl_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.din(w_dff_B_IVyUdDth9_2));
	jspl jspl_w_n1245_0(.douta(w_n1245_0[0]),.doutb(w_n1245_0[1]),.din(n1245));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(w_dff_B_vPZYQ9446_2));
	jspl jspl_w_n1250_0(.douta(w_n1250_0[0]),.doutb(w_n1250_0[1]),.din(n1250));
	jspl jspl_w_n1252_0(.douta(w_n1252_0[0]),.doutb(w_n1252_0[1]),.din(w_dff_B_rWoV4dyW9_2));
	jspl jspl_w_n1255_0(.douta(w_n1255_0[0]),.doutb(w_n1255_0[1]),.din(n1255));
	jspl jspl_w_n1257_0(.douta(w_n1257_0[0]),.doutb(w_n1257_0[1]),.din(w_dff_B_wQxdIANl7_2));
	jspl jspl_w_n1260_0(.douta(w_n1260_0[0]),.doutb(w_n1260_0[1]),.din(n1260));
	jspl jspl_w_n1262_0(.douta(w_n1262_0[0]),.doutb(w_n1262_0[1]),.din(w_dff_B_mp4WhI0R0_2));
	jspl jspl_w_n1265_0(.douta(w_n1265_0[0]),.doutb(w_n1265_0[1]),.din(n1265));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(w_dff_B_wCNWPAxc6_2));
	jspl jspl_w_n1267_0(.douta(w_n1267_0[0]),.doutb(w_n1267_0[1]),.din(w_dff_B_1tzjXXiY8_2));
	jspl jspl_w_n1270_0(.douta(w_n1270_0[0]),.doutb(w_n1270_0[1]),.din(n1270));
	jspl jspl_w_n1272_0(.douta(w_n1272_0[0]),.doutb(w_n1272_0[1]),.din(n1272));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(w_dff_B_4RzogzYx1_2));
	jspl jspl_w_n1274_0(.douta(w_n1274_0[0]),.doutb(w_n1274_0[1]),.din(n1274));
	jspl jspl_w_n1275_0(.douta(w_n1275_0[0]),.doutb(w_n1275_0[1]),.din(w_dff_B_bXuZ2R9U2_2));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(n1276));
	jspl jspl_w_n1277_0(.douta(w_n1277_0[0]),.doutb(w_n1277_0[1]),.din(w_dff_B_XFi4CKxd4_2));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(n1278));
	jspl jspl_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.din(w_dff_B_Lm9mW8yr3_2));
	jspl jspl_w_n1280_0(.douta(w_n1280_0[0]),.doutb(w_n1280_0[1]),.din(n1280));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(w_dff_B_4unbKKyv2_2));
	jspl jspl_w_n1282_0(.douta(w_n1282_0[0]),.doutb(w_n1282_0[1]),.din(n1282));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(w_dff_B_6HhSHxWD4_2));
	jspl jspl_w_n1284_0(.douta(w_n1284_0[0]),.doutb(w_n1284_0[1]),.din(n1284));
	jspl jspl_w_n1285_0(.douta(w_n1285_0[0]),.doutb(w_n1285_0[1]),.din(w_dff_B_JVkXs9h96_2));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(n1286));
	jspl jspl_w_n1287_0(.douta(w_n1287_0[0]),.doutb(w_n1287_0[1]),.din(n1287));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(n1288));
	jspl jspl_w_n1289_0(.douta(w_n1289_0[0]),.doutb(w_n1289_0[1]),.din(n1289));
	jspl jspl_w_n1290_0(.douta(w_n1290_0[0]),.doutb(w_n1290_0[1]),.din(n1290));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_dff_A_o830kju60_1),.din(n1291));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(n1293));
	jspl jspl_w_n1294_0(.douta(w_n1294_0[0]),.doutb(w_dff_A_vXmbbNVz1_1),.din(n1294));
	jspl jspl_w_n1295_0(.douta(w_dff_A_J7L0F21u0_0),.doutb(w_n1295_0[1]),.din(n1295));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(w_dff_B_bG0rai9o5_2));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(w_dff_B_tgvlIUag2_2));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(w_dff_B_Rp3ucYYc1_2));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.din(w_dff_B_l85Ij3Ye7_2));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl jspl_w_n1327_0(.douta(w_n1327_0[0]),.doutb(w_n1327_0[1]),.din(w_dff_B_zoqa3g5I7_2));
	jspl jspl_w_n1330_0(.douta(w_n1330_0[0]),.doutb(w_n1330_0[1]),.din(n1330));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(w_dff_B_B4idFpAm8_2));
	jspl jspl_w_n1335_0(.douta(w_n1335_0[0]),.doutb(w_n1335_0[1]),.din(n1335));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(w_dff_B_LDWxq2Tz1_2));
	jspl jspl_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_n1340_0[1]),.din(n1340));
	jspl jspl_w_n1342_0(.douta(w_n1342_0[0]),.doutb(w_n1342_0[1]),.din(w_dff_B_QUpBqD0A6_2));
	jspl jspl_w_n1345_0(.douta(w_n1345_0[0]),.doutb(w_n1345_0[1]),.din(n1345));
	jspl jspl_w_n1347_0(.douta(w_n1347_0[0]),.doutb(w_n1347_0[1]),.din(w_dff_B_sIGu0EXt3_2));
	jspl jspl_w_n1350_0(.douta(w_n1350_0[0]),.doutb(w_n1350_0[1]),.din(n1350));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(w_dff_B_4OFR99W31_2));
	jspl jspl_w_n1352_0(.douta(w_n1352_0[0]),.doutb(w_n1352_0[1]),.din(w_dff_B_FySL7aDB0_2));
	jspl jspl_w_n1355_0(.douta(w_n1355_0[0]),.doutb(w_n1355_0[1]),.din(n1355));
	jspl jspl_w_n1357_0(.douta(w_n1357_0[0]),.doutb(w_n1357_0[1]),.din(n1357));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.din(n1359));
	jspl jspl_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.din(w_dff_B_72tu2LAE3_2));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1362_0(.douta(w_n1362_0[0]),.doutb(w_n1362_0[1]),.din(w_dff_B_oXKCQvLj0_2));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(n1363));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_n1364_0[1]),.din(w_dff_B_FMdovfI97_2));
	jspl jspl_w_n1365_0(.douta(w_n1365_0[0]),.doutb(w_n1365_0[1]),.din(n1365));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(w_dff_B_LXPE0yOq1_2));
	jspl jspl_w_n1367_0(.douta(w_n1367_0[0]),.doutb(w_n1367_0[1]),.din(n1367));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(w_dff_B_Js1sOPgh7_2));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(n1369));
	jspl jspl_w_n1370_0(.douta(w_n1370_0[0]),.doutb(w_n1370_0[1]),.din(w_dff_B_MCd6ORrO0_2));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(n1373));
	jspl jspl_w_n1374_0(.douta(w_n1374_0[0]),.doutb(w_n1374_0[1]),.din(n1374));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(n1376));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(n1378));
	jspl jspl_w_n1379_0(.douta(w_n1379_0[0]),.doutb(w_dff_A_uVFeJtGu4_1),.din(n1379));
	jspl jspl_w_n1384_0(.douta(w_n1384_0[0]),.doutb(w_n1384_0[1]),.din(n1384));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(w_dff_B_63aFH6jf5_2));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(w_dff_B_Pd21kpZx1_2));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(w_dff_B_IbvucGwe3_2));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(w_dff_B_o7k5VhFC6_2));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(w_dff_B_aWErp4ZT3_2));
	jspl jspl_w_n1408_0(.douta(w_n1408_0[0]),.doutb(w_n1408_0[1]),.din(n1408));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(w_dff_B_kL36koVf8_2));
	jspl jspl_w_n1413_0(.douta(w_n1413_0[0]),.doutb(w_n1413_0[1]),.din(n1413));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(w_dff_B_XU9zNzmb9_2));
	jspl jspl_w_n1418_0(.douta(w_n1418_0[0]),.doutb(w_n1418_0[1]),.din(n1418));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(w_dff_B_3uQSKymP1_2));
	jspl jspl_w_n1423_0(.douta(w_n1423_0[0]),.doutb(w_n1423_0[1]),.din(n1423));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(w_dff_B_EzliOta12_2));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(w_dff_B_obud84Fq6_2));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(w_dff_B_P5aKcMzV6_2));
	jspl jspl_w_n1430_0(.douta(w_n1430_0[0]),.doutb(w_n1430_0[1]),.din(w_dff_B_S3RGNprc3_2));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1435_0(.douta(w_n1435_0[0]),.doutb(w_n1435_0[1]),.din(n1435));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(n1436));
	jspl jspl_w_n1437_0(.douta(w_n1437_0[0]),.doutb(w_n1437_0[1]),.din(n1437));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_n1438_0[1]),.din(n1438));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.din(w_dff_B_7AmvrWmr2_2));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl jspl_w_n1442_0(.douta(w_n1442_0[0]),.doutb(w_n1442_0[1]),.din(w_dff_B_QSdI15m68_2));
	jspl jspl_w_n1443_0(.douta(w_n1443_0[0]),.doutb(w_n1443_0[1]),.din(n1443));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(w_dff_B_T1ZHVrvU9_2));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(w_dff_B_3LZA2KGF3_2));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1448_0(.douta(w_n1448_0[0]),.doutb(w_n1448_0[1]),.din(w_dff_B_9qHtF55P1_2));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(n1449));
	jspl jspl_w_n1450_0(.douta(w_n1450_0[0]),.doutb(w_n1450_0[1]),.din(n1450));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(n1454));
	jspl jspl_w_n1455_0(.douta(w_n1455_0[0]),.doutb(w_dff_A_q7PYhXqR0_1),.din(n1455));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(n1460));
	jspl jspl_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.din(w_dff_B_7IYrndFR5_2));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(w_dff_B_p3ZNSoEw1_2));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(w_dff_B_qRHni46W2_2));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(n1474));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(w_dff_B_SlMs5Ypt1_2));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(n1479));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(w_dff_B_5wq6JhJu8_2));
	jspl jspl_w_n1484_0(.douta(w_n1484_0[0]),.doutb(w_n1484_0[1]),.din(n1484));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(w_dff_B_JzzDAZy18_2));
	jspl jspl_w_n1489_0(.douta(w_n1489_0[0]),.doutb(w_n1489_0[1]),.din(n1489));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(w_dff_B_88iN42Kq8_2));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(w_dff_B_cP8Rbmyk5_2));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(w_dff_B_3aHAWKT57_2));
	jspl jspl_w_n1499_0(.douta(w_n1499_0[0]),.doutb(w_n1499_0[1]),.din(w_dff_B_1ZVbO9WY8_2));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(w_dff_B_w3yWoLIG5_2));
	jspl jspl_w_n1501_0(.douta(w_n1501_0[0]),.doutb(w_n1501_0[1]),.din(w_dff_B_0ytc6keY6_2));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.din(n1506));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(n1507));
	jspl jspl_w_n1508_0(.douta(w_n1508_0[0]),.doutb(w_n1508_0[1]),.din(n1508));
	jspl jspl_w_n1509_0(.douta(w_n1509_0[0]),.doutb(w_n1509_0[1]),.din(n1509));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1511_0(.douta(w_n1511_0[0]),.doutb(w_n1511_0[1]),.din(n1511));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(n1512));
	jspl jspl_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.din(w_dff_B_wnhFjLNo7_2));
	jspl jspl_w_n1514_0(.douta(w_n1514_0[0]),.doutb(w_n1514_0[1]),.din(n1514));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(w_dff_B_EbZ9Y5HW1_2));
	jspl jspl_w_n1516_0(.douta(w_n1516_0[0]),.doutb(w_n1516_0[1]),.din(n1516));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(w_dff_B_FLkG0m4S9_2));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1519_0(.douta(w_n1519_0[0]),.doutb(w_dff_A_PxH1NRvU1_1),.din(n1519));
	jspl jspl_w_n1521_0(.douta(w_n1521_0[0]),.doutb(w_n1521_0[1]),.din(n1521));
	jspl jspl_w_n1523_0(.douta(w_n1523_0[0]),.doutb(w_n1523_0[1]),.din(n1523));
	jspl jspl_w_n1524_0(.douta(w_n1524_0[0]),.doutb(w_dff_A_FdAfEhwx6_1),.din(n1524));
	jspl jspl_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.din(n1529));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(n1534));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(w_dff_B_jZxX9Yif1_2));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(w_dff_B_HCrwfOX29_2));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(w_dff_B_PcSwCouR6_2));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(n1548));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_n1550_0[1]),.din(w_dff_B_7fjS4I5R0_2));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(w_dff_B_t8ZmUGWO1_2));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(w_dff_B_RkwElSTr3_2));
	jspl jspl_w_n1558_0(.douta(w_n1558_0[0]),.doutb(w_n1558_0[1]),.din(w_dff_B_gP79HKPg5_2));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(w_dff_B_baoqdbM52_2));
	jspl jspl_w_n1563_0(.douta(w_n1563_0[0]),.doutb(w_n1563_0[1]),.din(w_dff_B_p4XeoJmg1_2));
	jspl jspl_w_n1564_0(.douta(w_n1564_0[0]),.doutb(w_n1564_0[1]),.din(w_dff_B_oAJS2gxH9_2));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(w_dff_B_BxO64W1V2_2));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_n1568_0[1]),.din(n1568));
	jspl jspl_w_n1570_0(.douta(w_n1570_0[0]),.doutb(w_n1570_0[1]),.din(n1570));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(n1571));
	jspl jspl_w_n1572_0(.douta(w_n1572_0[0]),.doutb(w_n1572_0[1]),.din(n1572));
	jspl jspl_w_n1573_0(.douta(w_n1573_0[0]),.doutb(w_n1573_0[1]),.din(n1573));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(n1574));
	jspl jspl_w_n1575_0(.douta(w_n1575_0[0]),.doutb(w_n1575_0[1]),.din(n1575));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(n1576));
	jspl jspl_w_n1577_0(.douta(w_n1577_0[0]),.doutb(w_n1577_0[1]),.din(n1577));
	jspl jspl_w_n1578_0(.douta(w_n1578_0[0]),.doutb(w_n1578_0[1]),.din(n1578));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(w_dff_B_W50Qyrbw6_2));
	jspl jspl_w_n1580_0(.douta(w_n1580_0[0]),.doutb(w_n1580_0[1]),.din(n1580));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_dff_A_ZZHp1yH95_1),.din(n1581));
	jspl jspl_w_n1583_0(.douta(w_n1583_0[0]),.doutb(w_n1583_0[1]),.din(n1583));
	jspl jspl_w_n1585_0(.douta(w_n1585_0[0]),.doutb(w_n1585_0[1]),.din(n1585));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_dff_A_G80OTdUX1_1),.din(n1586));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(w_dff_B_vPvA7ghK4_2));
	jspl jspl_w_n1600_0(.douta(w_n1600_0[0]),.doutb(w_n1600_0[1]),.din(n1600));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(w_dff_B_o9zY27mx9_2));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(w_dff_B_0qTTQ4Ah9_2));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(w_dff_B_NWclf5rq6_2));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(w_dff_B_s48Z0v4b3_2));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(w_dff_B_xoIVA3GF0_2));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(w_dff_B_91rMqHuE3_2));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_n1617_0[1]),.din(w_dff_B_wjKxITkK3_2));
	jspl jspl_w_n1620_0(.douta(w_n1620_0[0]),.doutb(w_n1620_0[1]),.din(w_dff_B_jQ8wPSVW4_2));
	jspl jspl_w_n1621_0(.douta(w_n1621_0[0]),.doutb(w_n1621_0[1]),.din(w_dff_B_6V8zst9C7_2));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(w_dff_B_a3zElpLN1_2));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(n1628));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1630_0(.douta(w_n1630_0[0]),.doutb(w_n1630_0[1]),.din(n1630));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(n1631));
	jspl jspl_w_n1632_0(.douta(w_n1632_0[0]),.doutb(w_n1632_0[1]),.din(n1632));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(n1633));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(n1634));
	jspl jspl_w_n1635_0(.douta(w_n1635_0[0]),.doutb(w_n1635_0[1]),.din(n1635));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(n1636));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(n1638));
	jspl jspl_w_n1640_0(.douta(w_n1640_0[0]),.doutb(w_n1640_0[1]),.din(n1640));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_dff_A_KvEs2OMJ1_1),.din(n1641));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(n1646));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(w_dff_B_PRuDwE9Y3_2));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(w_dff_B_9eCQOicP7_2));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(w_dff_B_WrJ6V0nm5_2));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(w_dff_B_9Pq9g6YL3_2));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(w_dff_B_mPJtTvrl4_2));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(w_dff_B_LZLyJm3j4_2));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(w_dff_B_ja0mBXim9_2));
	jspl jspl_w_n1668_0(.douta(w_n1668_0[0]),.doutb(w_n1668_0[1]),.din(w_dff_B_hWflD2Rx4_2));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(w_dff_B_Gi5MsAd61_2));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(w_dff_B_kJbWkHSd9_2));
	jspl jspl_w_n1673_0(.douta(w_n1673_0[0]),.doutb(w_n1673_0[1]),.din(w_dff_B_6Y8cJT6S0_2));
	jspl jspl_w_n1676_0(.douta(w_n1676_0[0]),.doutb(w_n1676_0[1]),.din(n1676));
	jspl jspl_w_n1678_0(.douta(w_n1678_0[0]),.doutb(w_n1678_0[1]),.din(n1678));
	jspl jspl_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1681_0(.douta(w_n1681_0[0]),.doutb(w_n1681_0[1]),.din(n1681));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(n1682));
	jspl jspl_w_n1683_0(.douta(w_n1683_0[0]),.doutb(w_n1683_0[1]),.din(n1683));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(n1684));
	jspl jspl_w_n1685_0(.douta(w_n1685_0[0]),.doutb(w_n1685_0[1]),.din(n1685));
	jspl jspl_w_n1686_0(.douta(w_n1686_0[0]),.doutb(w_n1686_0[1]),.din(n1686));
	jspl jspl_w_n1688_0(.douta(w_n1688_0[0]),.doutb(w_n1688_0[1]),.din(n1688));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_dff_A_hBr7Bvkn6_1),.din(n1689));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(n1694));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_dff_A_FN7R7Wuv2_1),.din(n1697));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(w_dff_B_a2Kjpush8_2));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(w_dff_B_YwNIF9Vn6_2));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(w_dff_B_oclFPpvi7_2));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(w_dff_B_RnJwT5Ck2_2));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(w_dff_B_CBStuMlU2_2));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(w_dff_B_rttDH4w78_2));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(w_dff_B_hmcBy8Y75_2));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(w_dff_B_Cy9xGHOQ5_2));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_n1720_0[1]),.din(n1720));
	jspl jspl_w_n1721_0(.douta(w_n1721_0[0]),.doutb(w_n1721_0[1]),.din(n1721));
	jspl jspl_w_n1722_0(.douta(w_n1722_0[0]),.doutb(w_n1722_0[1]),.din(n1722));
	jspl jspl_w_n1723_0(.douta(w_n1723_0[0]),.doutb(w_n1723_0[1]),.din(n1723));
	jspl jspl_w_n1724_0(.douta(w_n1724_0[0]),.doutb(w_n1724_0[1]),.din(n1724));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1726_0(.douta(w_n1726_0[0]),.doutb(w_n1726_0[1]),.din(n1726));
	jspl jspl_w_n1727_0(.douta(w_n1727_0[0]),.doutb(w_dff_A_itjcwYbR2_1),.din(n1727));
	jspl jspl_w_n1734_0(.douta(w_n1734_0[0]),.doutb(w_n1734_0[1]),.din(n1734));
	jspl jspl_w_n1737_0(.douta(w_n1737_0[0]),.doutb(w_dff_A_bsSlG3hO7_1),.din(n1737));
	jspl jspl_w_n1739_0(.douta(w_n1739_0[0]),.doutb(w_n1739_0[1]),.din(w_dff_B_5eC0TGI62_2));
	jspl jspl_w_n1742_0(.douta(w_n1742_0[0]),.doutb(w_n1742_0[1]),.din(w_dff_B_M75QlrxF7_2));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(w_dff_B_12hr5EGl3_2));
	jspl jspl_w_n1747_0(.douta(w_n1747_0[0]),.doutb(w_n1747_0[1]),.din(w_dff_B_j4DIVSxT5_2));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(w_dff_B_t3UUnhQ63_2));
	jspl jspl_w_n1749_0(.douta(w_n1749_0[0]),.doutb(w_n1749_0[1]),.din(w_dff_B_chfeBSJ11_2));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_n1758_0[1]),.din(n1758));
	jspl jspl_w_n1759_0(.douta(w_n1759_0[0]),.doutb(w_n1759_0[1]),.din(n1759));
	jspl jspl_w_n1760_0(.douta(w_n1760_0[0]),.doutb(w_dff_A_2vTb8S2q8_1),.din(n1760));
	jspl jspl_w_n1767_0(.douta(w_n1767_0[0]),.doutb(w_n1767_0[1]),.din(n1767));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_dff_A_qYRAclYB1_1),.din(n1770));
	jspl jspl_w_n1772_0(.douta(w_n1772_0[0]),.doutb(w_n1772_0[1]),.din(w_dff_B_2CXTIugB1_2));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(w_dff_B_8KA5KVCB4_2));
	jspl jspl_w_n1776_0(.douta(w_n1776_0[0]),.doutb(w_n1776_0[1]),.din(w_dff_B_3OSCaDKz1_2));
	jspl jspl_w_n1777_0(.douta(w_n1777_0[0]),.doutb(w_n1777_0[1]),.din(w_dff_B_shCeCe4X9_2));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(n1780));
	jspl jspl_w_n1782_0(.douta(w_n1782_0[0]),.doutb(w_n1782_0[1]),.din(n1782));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1784_0(.douta(w_n1784_0[0]),.doutb(w_n1784_0[1]),.din(n1784));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_dff_A_4KVlAlWx1_1),.din(n1786));
	jspl jspl_w_n1793_0(.douta(w_n1793_0[0]),.doutb(w_n1793_0[1]),.din(n1793));
	jspl jspl_w_n1796_0(.douta(w_n1796_0[0]),.doutb(w_dff_A_AC3zetFj0_1),.din(n1796));
	jspl jspl_w_n1797_0(.douta(w_n1797_0[0]),.doutb(w_n1797_0[1]),.din(w_dff_B_h5KCZ1I58_2));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(w_dff_B_qbkifT6e7_2));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_n1801_0[1]),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(n1803));
	jspl jspl_w_n1804_0(.douta(w_n1804_0[0]),.doutb(w_n1804_0[1]),.din(n1804));
	jspl jspl_w_n1805_0(.douta(w_n1805_0[0]),.doutb(w_dff_A_EijMotbY9_1),.din(n1805));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(w_dff_B_lqpZejf25_2));
	jspl jspl_w_n1810_0(.douta(w_n1810_0[0]),.doutb(w_n1810_0[1]),.din(n1810));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_n1817_0[1]),.din(n1817));
	jspl jspl_w_n1818_0(.douta(w_dff_A_MML1jZwp4_0),.doutb(w_n1818_0[1]),.din(n1818));
	jdff dff_B_vzvAZJxt5_0(.din(n72),.dout(w_dff_B_vzvAZJxt5_0),.clk(gclk));
	jdff dff_B_SUExNrn46_0(.din(w_dff_B_vzvAZJxt5_0),.dout(w_dff_B_SUExNrn46_0),.clk(gclk));
	jdff dff_B_QdpwnOgJ1_1(.din(n76),.dout(w_dff_B_QdpwnOgJ1_1),.clk(gclk));
	jdff dff_B_gafEQwL95_1(.din(w_dff_B_QdpwnOgJ1_1),.dout(w_dff_B_gafEQwL95_1),.clk(gclk));
	jdff dff_B_89v3w0f13_1(.din(w_dff_B_gafEQwL95_1),.dout(w_dff_B_89v3w0f13_1),.clk(gclk));
	jdff dff_B_InF7qtmv0_1(.din(n87),.dout(w_dff_B_InF7qtmv0_1),.clk(gclk));
	jdff dff_B_1cqxJKRO6_1(.din(w_dff_B_InF7qtmv0_1),.dout(w_dff_B_1cqxJKRO6_1),.clk(gclk));
	jdff dff_B_cP4vnAxd8_1(.din(w_dff_B_1cqxJKRO6_1),.dout(w_dff_B_cP4vnAxd8_1),.clk(gclk));
	jdff dff_B_Jcr8KLbV6_1(.din(w_dff_B_cP4vnAxd8_1),.dout(w_dff_B_Jcr8KLbV6_1),.clk(gclk));
	jdff dff_B_6g4JKUI96_1(.din(w_dff_B_Jcr8KLbV6_1),.dout(w_dff_B_6g4JKUI96_1),.clk(gclk));
	jdff dff_B_yVHZgx371_1(.din(w_dff_B_6g4JKUI96_1),.dout(w_dff_B_yVHZgx371_1),.clk(gclk));
	jdff dff_B_r6Cme3p80_1(.din(n107),.dout(w_dff_B_r6Cme3p80_1),.clk(gclk));
	jdff dff_B_Ou6HbKVR3_1(.din(w_dff_B_r6Cme3p80_1),.dout(w_dff_B_Ou6HbKVR3_1),.clk(gclk));
	jdff dff_B_BqKy0Luv7_1(.din(w_dff_B_Ou6HbKVR3_1),.dout(w_dff_B_BqKy0Luv7_1),.clk(gclk));
	jdff dff_B_mhYvGvOc6_1(.din(w_dff_B_BqKy0Luv7_1),.dout(w_dff_B_mhYvGvOc6_1),.clk(gclk));
	jdff dff_B_RZC5JMcr9_1(.din(w_dff_B_mhYvGvOc6_1),.dout(w_dff_B_RZC5JMcr9_1),.clk(gclk));
	jdff dff_B_bhnAR0OI2_1(.din(w_dff_B_RZC5JMcr9_1),.dout(w_dff_B_bhnAR0OI2_1),.clk(gclk));
	jdff dff_B_3prdParx6_1(.din(w_dff_B_bhnAR0OI2_1),.dout(w_dff_B_3prdParx6_1),.clk(gclk));
	jdff dff_B_7lGMKzH84_1(.din(w_dff_B_3prdParx6_1),.dout(w_dff_B_7lGMKzH84_1),.clk(gclk));
	jdff dff_B_UWWTPYVO4_1(.din(w_dff_B_7lGMKzH84_1),.dout(w_dff_B_UWWTPYVO4_1),.clk(gclk));
	jdff dff_B_Jj1iQ7xH1_1(.din(n136),.dout(w_dff_B_Jj1iQ7xH1_1),.clk(gclk));
	jdff dff_B_eEbaSphm0_1(.din(w_dff_B_Jj1iQ7xH1_1),.dout(w_dff_B_eEbaSphm0_1),.clk(gclk));
	jdff dff_B_ClFCjDTN8_1(.din(w_dff_B_eEbaSphm0_1),.dout(w_dff_B_ClFCjDTN8_1),.clk(gclk));
	jdff dff_B_7JIWZQuW2_1(.din(w_dff_B_ClFCjDTN8_1),.dout(w_dff_B_7JIWZQuW2_1),.clk(gclk));
	jdff dff_B_nT9vTHWR8_1(.din(w_dff_B_7JIWZQuW2_1),.dout(w_dff_B_nT9vTHWR8_1),.clk(gclk));
	jdff dff_B_4BbOqokv2_1(.din(w_dff_B_nT9vTHWR8_1),.dout(w_dff_B_4BbOqokv2_1),.clk(gclk));
	jdff dff_B_Bpxv5lyf9_1(.din(w_dff_B_4BbOqokv2_1),.dout(w_dff_B_Bpxv5lyf9_1),.clk(gclk));
	jdff dff_B_8PSTu8Y33_1(.din(w_dff_B_Bpxv5lyf9_1),.dout(w_dff_B_8PSTu8Y33_1),.clk(gclk));
	jdff dff_B_N4uXRTGa1_1(.din(w_dff_B_8PSTu8Y33_1),.dout(w_dff_B_N4uXRTGa1_1),.clk(gclk));
	jdff dff_B_fZ2jmcSn8_1(.din(w_dff_B_N4uXRTGa1_1),.dout(w_dff_B_fZ2jmcSn8_1),.clk(gclk));
	jdff dff_B_yfPk977F3_1(.din(w_dff_B_fZ2jmcSn8_1),.dout(w_dff_B_yfPk977F3_1),.clk(gclk));
	jdff dff_B_BnXbdPhm6_1(.din(w_dff_B_yfPk977F3_1),.dout(w_dff_B_BnXbdPhm6_1),.clk(gclk));
	jdff dff_B_V9VTPdn51_1(.din(n171),.dout(w_dff_B_V9VTPdn51_1),.clk(gclk));
	jdff dff_B_X1hFynFU2_1(.din(w_dff_B_V9VTPdn51_1),.dout(w_dff_B_X1hFynFU2_1),.clk(gclk));
	jdff dff_B_teMGEn4P1_1(.din(w_dff_B_X1hFynFU2_1),.dout(w_dff_B_teMGEn4P1_1),.clk(gclk));
	jdff dff_B_jPKZdBkI7_1(.din(w_dff_B_teMGEn4P1_1),.dout(w_dff_B_jPKZdBkI7_1),.clk(gclk));
	jdff dff_B_cmuusSQw1_1(.din(w_dff_B_jPKZdBkI7_1),.dout(w_dff_B_cmuusSQw1_1),.clk(gclk));
	jdff dff_B_AoEMteKx4_1(.din(w_dff_B_cmuusSQw1_1),.dout(w_dff_B_AoEMteKx4_1),.clk(gclk));
	jdff dff_B_Ey3muK8q4_1(.din(w_dff_B_AoEMteKx4_1),.dout(w_dff_B_Ey3muK8q4_1),.clk(gclk));
	jdff dff_B_yGHGyHBk9_1(.din(w_dff_B_Ey3muK8q4_1),.dout(w_dff_B_yGHGyHBk9_1),.clk(gclk));
	jdff dff_B_jKFyHFyH7_1(.din(w_dff_B_yGHGyHBk9_1),.dout(w_dff_B_jKFyHFyH7_1),.clk(gclk));
	jdff dff_B_IxjpZylU9_1(.din(w_dff_B_jKFyHFyH7_1),.dout(w_dff_B_IxjpZylU9_1),.clk(gclk));
	jdff dff_B_cAlEFDav4_1(.din(w_dff_B_IxjpZylU9_1),.dout(w_dff_B_cAlEFDav4_1),.clk(gclk));
	jdff dff_B_awJm5IGm1_1(.din(w_dff_B_cAlEFDav4_1),.dout(w_dff_B_awJm5IGm1_1),.clk(gclk));
	jdff dff_B_ZpPlB2Wm0_1(.din(w_dff_B_awJm5IGm1_1),.dout(w_dff_B_ZpPlB2Wm0_1),.clk(gclk));
	jdff dff_B_H6n3cIIX0_1(.din(w_dff_B_ZpPlB2Wm0_1),.dout(w_dff_B_H6n3cIIX0_1),.clk(gclk));
	jdff dff_B_DpFfkr0Y4_1(.din(w_dff_B_H6n3cIIX0_1),.dout(w_dff_B_DpFfkr0Y4_1),.clk(gclk));
	jdff dff_B_m2ENnNou3_1(.din(n213),.dout(w_dff_B_m2ENnNou3_1),.clk(gclk));
	jdff dff_B_6o123e5Y7_1(.din(w_dff_B_m2ENnNou3_1),.dout(w_dff_B_6o123e5Y7_1),.clk(gclk));
	jdff dff_B_VqpbOfil5_1(.din(w_dff_B_6o123e5Y7_1),.dout(w_dff_B_VqpbOfil5_1),.clk(gclk));
	jdff dff_B_7jW0raWj5_1(.din(w_dff_B_VqpbOfil5_1),.dout(w_dff_B_7jW0raWj5_1),.clk(gclk));
	jdff dff_B_tUSHvTyN0_1(.din(w_dff_B_7jW0raWj5_1),.dout(w_dff_B_tUSHvTyN0_1),.clk(gclk));
	jdff dff_B_r7osvCbN1_1(.din(w_dff_B_tUSHvTyN0_1),.dout(w_dff_B_r7osvCbN1_1),.clk(gclk));
	jdff dff_B_yrE90Xy56_1(.din(w_dff_B_r7osvCbN1_1),.dout(w_dff_B_yrE90Xy56_1),.clk(gclk));
	jdff dff_B_cIap07mj7_1(.din(w_dff_B_yrE90Xy56_1),.dout(w_dff_B_cIap07mj7_1),.clk(gclk));
	jdff dff_B_3j8TDRSL8_1(.din(w_dff_B_cIap07mj7_1),.dout(w_dff_B_3j8TDRSL8_1),.clk(gclk));
	jdff dff_B_6s4IeKIh3_1(.din(w_dff_B_3j8TDRSL8_1),.dout(w_dff_B_6s4IeKIh3_1),.clk(gclk));
	jdff dff_B_hYLLQ15x6_1(.din(w_dff_B_6s4IeKIh3_1),.dout(w_dff_B_hYLLQ15x6_1),.clk(gclk));
	jdff dff_B_BAd2M8LT6_1(.din(w_dff_B_hYLLQ15x6_1),.dout(w_dff_B_BAd2M8LT6_1),.clk(gclk));
	jdff dff_B_DSoG4S084_1(.din(w_dff_B_BAd2M8LT6_1),.dout(w_dff_B_DSoG4S084_1),.clk(gclk));
	jdff dff_B_355LobdI0_1(.din(w_dff_B_DSoG4S084_1),.dout(w_dff_B_355LobdI0_1),.clk(gclk));
	jdff dff_B_fukn4ltA0_1(.din(w_dff_B_355LobdI0_1),.dout(w_dff_B_fukn4ltA0_1),.clk(gclk));
	jdff dff_B_qgJReu1N7_1(.din(w_dff_B_fukn4ltA0_1),.dout(w_dff_B_qgJReu1N7_1),.clk(gclk));
	jdff dff_B_3N1B4Rtq0_1(.din(w_dff_B_qgJReu1N7_1),.dout(w_dff_B_3N1B4Rtq0_1),.clk(gclk));
	jdff dff_B_vJqVPxU03_1(.din(w_dff_B_3N1B4Rtq0_1),.dout(w_dff_B_vJqVPxU03_1),.clk(gclk));
	jdff dff_B_CwSRRwjN5_1(.din(n262),.dout(w_dff_B_CwSRRwjN5_1),.clk(gclk));
	jdff dff_B_GedtU0vi4_1(.din(w_dff_B_CwSRRwjN5_1),.dout(w_dff_B_GedtU0vi4_1),.clk(gclk));
	jdff dff_B_oovehKht1_1(.din(w_dff_B_GedtU0vi4_1),.dout(w_dff_B_oovehKht1_1),.clk(gclk));
	jdff dff_B_iN5qnS8z5_1(.din(w_dff_B_oovehKht1_1),.dout(w_dff_B_iN5qnS8z5_1),.clk(gclk));
	jdff dff_B_DL886yBF3_1(.din(w_dff_B_iN5qnS8z5_1),.dout(w_dff_B_DL886yBF3_1),.clk(gclk));
	jdff dff_B_SVAJzocY6_1(.din(w_dff_B_DL886yBF3_1),.dout(w_dff_B_SVAJzocY6_1),.clk(gclk));
	jdff dff_B_urygT3bm1_1(.din(w_dff_B_SVAJzocY6_1),.dout(w_dff_B_urygT3bm1_1),.clk(gclk));
	jdff dff_B_jORn2jGt1_1(.din(w_dff_B_urygT3bm1_1),.dout(w_dff_B_jORn2jGt1_1),.clk(gclk));
	jdff dff_B_bZkIttkF1_1(.din(w_dff_B_jORn2jGt1_1),.dout(w_dff_B_bZkIttkF1_1),.clk(gclk));
	jdff dff_B_RfEAPgye7_1(.din(w_dff_B_bZkIttkF1_1),.dout(w_dff_B_RfEAPgye7_1),.clk(gclk));
	jdff dff_B_54bn7vVA8_1(.din(w_dff_B_RfEAPgye7_1),.dout(w_dff_B_54bn7vVA8_1),.clk(gclk));
	jdff dff_B_3v6pA5oI5_1(.din(w_dff_B_54bn7vVA8_1),.dout(w_dff_B_3v6pA5oI5_1),.clk(gclk));
	jdff dff_B_v2VG6z1c8_1(.din(w_dff_B_3v6pA5oI5_1),.dout(w_dff_B_v2VG6z1c8_1),.clk(gclk));
	jdff dff_B_qxzwDn6E8_1(.din(w_dff_B_v2VG6z1c8_1),.dout(w_dff_B_qxzwDn6E8_1),.clk(gclk));
	jdff dff_B_XwVx16Ix4_1(.din(w_dff_B_qxzwDn6E8_1),.dout(w_dff_B_XwVx16Ix4_1),.clk(gclk));
	jdff dff_B_QyljmIj94_1(.din(w_dff_B_XwVx16Ix4_1),.dout(w_dff_B_QyljmIj94_1),.clk(gclk));
	jdff dff_B_1mmN5BzQ6_1(.din(w_dff_B_QyljmIj94_1),.dout(w_dff_B_1mmN5BzQ6_1),.clk(gclk));
	jdff dff_B_3XoXNWDN7_1(.din(w_dff_B_1mmN5BzQ6_1),.dout(w_dff_B_3XoXNWDN7_1),.clk(gclk));
	jdff dff_B_Q9fGXPqs0_1(.din(w_dff_B_3XoXNWDN7_1),.dout(w_dff_B_Q9fGXPqs0_1),.clk(gclk));
	jdff dff_B_Wg3iCdZg8_1(.din(w_dff_B_Q9fGXPqs0_1),.dout(w_dff_B_Wg3iCdZg8_1),.clk(gclk));
	jdff dff_B_r3WimfWD0_1(.din(w_dff_B_Wg3iCdZg8_1),.dout(w_dff_B_r3WimfWD0_1),.clk(gclk));
	jdff dff_B_zFvfwIzp7_1(.din(n318),.dout(w_dff_B_zFvfwIzp7_1),.clk(gclk));
	jdff dff_B_qy1kQbUX1_1(.din(w_dff_B_zFvfwIzp7_1),.dout(w_dff_B_qy1kQbUX1_1),.clk(gclk));
	jdff dff_B_x69OOTQN3_1(.din(w_dff_B_qy1kQbUX1_1),.dout(w_dff_B_x69OOTQN3_1),.clk(gclk));
	jdff dff_B_rCCDKrWU9_1(.din(w_dff_B_x69OOTQN3_1),.dout(w_dff_B_rCCDKrWU9_1),.clk(gclk));
	jdff dff_B_Vxl0881H9_1(.din(w_dff_B_rCCDKrWU9_1),.dout(w_dff_B_Vxl0881H9_1),.clk(gclk));
	jdff dff_B_3PWAp9Kk9_1(.din(w_dff_B_Vxl0881H9_1),.dout(w_dff_B_3PWAp9Kk9_1),.clk(gclk));
	jdff dff_B_7ClctyZ17_1(.din(w_dff_B_3PWAp9Kk9_1),.dout(w_dff_B_7ClctyZ17_1),.clk(gclk));
	jdff dff_B_tRLlBSwL4_1(.din(w_dff_B_7ClctyZ17_1),.dout(w_dff_B_tRLlBSwL4_1),.clk(gclk));
	jdff dff_B_E8fVHq9U7_1(.din(w_dff_B_tRLlBSwL4_1),.dout(w_dff_B_E8fVHq9U7_1),.clk(gclk));
	jdff dff_B_rATvijCS6_1(.din(w_dff_B_E8fVHq9U7_1),.dout(w_dff_B_rATvijCS6_1),.clk(gclk));
	jdff dff_B_QHLHFRca2_1(.din(w_dff_B_rATvijCS6_1),.dout(w_dff_B_QHLHFRca2_1),.clk(gclk));
	jdff dff_B_mSfyylXG9_1(.din(w_dff_B_QHLHFRca2_1),.dout(w_dff_B_mSfyylXG9_1),.clk(gclk));
	jdff dff_B_MBBrBup01_1(.din(w_dff_B_mSfyylXG9_1),.dout(w_dff_B_MBBrBup01_1),.clk(gclk));
	jdff dff_B_B2o5QZKN3_1(.din(w_dff_B_MBBrBup01_1),.dout(w_dff_B_B2o5QZKN3_1),.clk(gclk));
	jdff dff_B_3411S7Qh3_1(.din(w_dff_B_B2o5QZKN3_1),.dout(w_dff_B_3411S7Qh3_1),.clk(gclk));
	jdff dff_B_3D87MeEd7_1(.din(w_dff_B_3411S7Qh3_1),.dout(w_dff_B_3D87MeEd7_1),.clk(gclk));
	jdff dff_B_5BltfdqI3_1(.din(w_dff_B_3D87MeEd7_1),.dout(w_dff_B_5BltfdqI3_1),.clk(gclk));
	jdff dff_B_0rXH0pJp2_1(.din(w_dff_B_5BltfdqI3_1),.dout(w_dff_B_0rXH0pJp2_1),.clk(gclk));
	jdff dff_B_GD49Hmfq1_1(.din(w_dff_B_0rXH0pJp2_1),.dout(w_dff_B_GD49Hmfq1_1),.clk(gclk));
	jdff dff_B_wSXpna8E5_1(.din(w_dff_B_GD49Hmfq1_1),.dout(w_dff_B_wSXpna8E5_1),.clk(gclk));
	jdff dff_B_9xZoLqYk6_1(.din(w_dff_B_wSXpna8E5_1),.dout(w_dff_B_9xZoLqYk6_1),.clk(gclk));
	jdff dff_B_NZoRyegg1_1(.din(w_dff_B_9xZoLqYk6_1),.dout(w_dff_B_NZoRyegg1_1),.clk(gclk));
	jdff dff_B_c3me6WE41_1(.din(w_dff_B_NZoRyegg1_1),.dout(w_dff_B_c3me6WE41_1),.clk(gclk));
	jdff dff_B_d7eeEngJ3_1(.din(w_dff_B_c3me6WE41_1),.dout(w_dff_B_d7eeEngJ3_1),.clk(gclk));
	jdff dff_B_kdsmAVtO7_1(.din(n381),.dout(w_dff_B_kdsmAVtO7_1),.clk(gclk));
	jdff dff_B_k1sgEzGa7_1(.din(w_dff_B_kdsmAVtO7_1),.dout(w_dff_B_k1sgEzGa7_1),.clk(gclk));
	jdff dff_B_j2EHEmno9_1(.din(w_dff_B_k1sgEzGa7_1),.dout(w_dff_B_j2EHEmno9_1),.clk(gclk));
	jdff dff_B_bKpyVoNp3_1(.din(w_dff_B_j2EHEmno9_1),.dout(w_dff_B_bKpyVoNp3_1),.clk(gclk));
	jdff dff_B_OecDV8788_1(.din(w_dff_B_bKpyVoNp3_1),.dout(w_dff_B_OecDV8788_1),.clk(gclk));
	jdff dff_B_Y35OwnYU3_1(.din(w_dff_B_OecDV8788_1),.dout(w_dff_B_Y35OwnYU3_1),.clk(gclk));
	jdff dff_B_JFNjBZFt9_1(.din(w_dff_B_Y35OwnYU3_1),.dout(w_dff_B_JFNjBZFt9_1),.clk(gclk));
	jdff dff_B_TL2bxGWf0_1(.din(w_dff_B_JFNjBZFt9_1),.dout(w_dff_B_TL2bxGWf0_1),.clk(gclk));
	jdff dff_B_axgoBAK62_1(.din(w_dff_B_TL2bxGWf0_1),.dout(w_dff_B_axgoBAK62_1),.clk(gclk));
	jdff dff_B_7FPtVNEg4_1(.din(w_dff_B_axgoBAK62_1),.dout(w_dff_B_7FPtVNEg4_1),.clk(gclk));
	jdff dff_B_ugwhrDwY8_1(.din(w_dff_B_7FPtVNEg4_1),.dout(w_dff_B_ugwhrDwY8_1),.clk(gclk));
	jdff dff_B_fLm8AuIN0_1(.din(w_dff_B_ugwhrDwY8_1),.dout(w_dff_B_fLm8AuIN0_1),.clk(gclk));
	jdff dff_B_GAM8RXKv7_1(.din(w_dff_B_fLm8AuIN0_1),.dout(w_dff_B_GAM8RXKv7_1),.clk(gclk));
	jdff dff_B_CUAIUGvI3_1(.din(w_dff_B_GAM8RXKv7_1),.dout(w_dff_B_CUAIUGvI3_1),.clk(gclk));
	jdff dff_B_hRB2htQv6_1(.din(w_dff_B_CUAIUGvI3_1),.dout(w_dff_B_hRB2htQv6_1),.clk(gclk));
	jdff dff_B_om1Gq63v3_1(.din(w_dff_B_hRB2htQv6_1),.dout(w_dff_B_om1Gq63v3_1),.clk(gclk));
	jdff dff_B_cBM9Hzd33_1(.din(w_dff_B_om1Gq63v3_1),.dout(w_dff_B_cBM9Hzd33_1),.clk(gclk));
	jdff dff_B_yPHyzvWq7_1(.din(w_dff_B_cBM9Hzd33_1),.dout(w_dff_B_yPHyzvWq7_1),.clk(gclk));
	jdff dff_B_1cTmXVId4_1(.din(w_dff_B_yPHyzvWq7_1),.dout(w_dff_B_1cTmXVId4_1),.clk(gclk));
	jdff dff_B_6ID0EMhh4_1(.din(w_dff_B_1cTmXVId4_1),.dout(w_dff_B_6ID0EMhh4_1),.clk(gclk));
	jdff dff_B_VSwwZBpj9_1(.din(w_dff_B_6ID0EMhh4_1),.dout(w_dff_B_VSwwZBpj9_1),.clk(gclk));
	jdff dff_B_UH1jfDFs6_1(.din(w_dff_B_VSwwZBpj9_1),.dout(w_dff_B_UH1jfDFs6_1),.clk(gclk));
	jdff dff_B_vAZaof7z0_1(.din(w_dff_B_UH1jfDFs6_1),.dout(w_dff_B_vAZaof7z0_1),.clk(gclk));
	jdff dff_B_tRp9EaF18_1(.din(w_dff_B_vAZaof7z0_1),.dout(w_dff_B_tRp9EaF18_1),.clk(gclk));
	jdff dff_B_Ydftyv7r1_1(.din(w_dff_B_tRp9EaF18_1),.dout(w_dff_B_Ydftyv7r1_1),.clk(gclk));
	jdff dff_B_nFLHIZA47_1(.din(w_dff_B_Ydftyv7r1_1),.dout(w_dff_B_nFLHIZA47_1),.clk(gclk));
	jdff dff_B_ZlVotAqf9_1(.din(w_dff_B_nFLHIZA47_1),.dout(w_dff_B_ZlVotAqf9_1),.clk(gclk));
	jdff dff_B_7lUb0BKv2_1(.din(n452),.dout(w_dff_B_7lUb0BKv2_1),.clk(gclk));
	jdff dff_B_QxQUFhzn0_1(.din(w_dff_B_7lUb0BKv2_1),.dout(w_dff_B_QxQUFhzn0_1),.clk(gclk));
	jdff dff_B_NJRF68sV5_1(.din(w_dff_B_QxQUFhzn0_1),.dout(w_dff_B_NJRF68sV5_1),.clk(gclk));
	jdff dff_B_9SwlEMC75_1(.din(w_dff_B_NJRF68sV5_1),.dout(w_dff_B_9SwlEMC75_1),.clk(gclk));
	jdff dff_B_uaoz8z8P3_1(.din(w_dff_B_9SwlEMC75_1),.dout(w_dff_B_uaoz8z8P3_1),.clk(gclk));
	jdff dff_B_fa9QVryM6_1(.din(w_dff_B_uaoz8z8P3_1),.dout(w_dff_B_fa9QVryM6_1),.clk(gclk));
	jdff dff_B_YjoGX06V4_1(.din(w_dff_B_fa9QVryM6_1),.dout(w_dff_B_YjoGX06V4_1),.clk(gclk));
	jdff dff_B_spc827hJ4_1(.din(w_dff_B_YjoGX06V4_1),.dout(w_dff_B_spc827hJ4_1),.clk(gclk));
	jdff dff_B_AfFkH6io8_1(.din(w_dff_B_spc827hJ4_1),.dout(w_dff_B_AfFkH6io8_1),.clk(gclk));
	jdff dff_B_lROTlTqo4_1(.din(w_dff_B_AfFkH6io8_1),.dout(w_dff_B_lROTlTqo4_1),.clk(gclk));
	jdff dff_B_xu5w64Ol1_1(.din(w_dff_B_lROTlTqo4_1),.dout(w_dff_B_xu5w64Ol1_1),.clk(gclk));
	jdff dff_B_e7S8QqC39_1(.din(w_dff_B_xu5w64Ol1_1),.dout(w_dff_B_e7S8QqC39_1),.clk(gclk));
	jdff dff_B_UpOR4GE39_1(.din(w_dff_B_e7S8QqC39_1),.dout(w_dff_B_UpOR4GE39_1),.clk(gclk));
	jdff dff_B_5PwDEXba4_1(.din(w_dff_B_UpOR4GE39_1),.dout(w_dff_B_5PwDEXba4_1),.clk(gclk));
	jdff dff_B_0PhRkLP33_1(.din(w_dff_B_5PwDEXba4_1),.dout(w_dff_B_0PhRkLP33_1),.clk(gclk));
	jdff dff_B_l5aAVy7v5_1(.din(w_dff_B_0PhRkLP33_1),.dout(w_dff_B_l5aAVy7v5_1),.clk(gclk));
	jdff dff_B_dpS8tZeW6_1(.din(w_dff_B_l5aAVy7v5_1),.dout(w_dff_B_dpS8tZeW6_1),.clk(gclk));
	jdff dff_B_aaOeSY6X0_1(.din(w_dff_B_dpS8tZeW6_1),.dout(w_dff_B_aaOeSY6X0_1),.clk(gclk));
	jdff dff_B_WL87fzhT6_1(.din(w_dff_B_aaOeSY6X0_1),.dout(w_dff_B_WL87fzhT6_1),.clk(gclk));
	jdff dff_B_CDxtdfPQ8_1(.din(w_dff_B_WL87fzhT6_1),.dout(w_dff_B_CDxtdfPQ8_1),.clk(gclk));
	jdff dff_B_uJkSSJsU0_1(.din(w_dff_B_CDxtdfPQ8_1),.dout(w_dff_B_uJkSSJsU0_1),.clk(gclk));
	jdff dff_B_K6dn33Fl4_1(.din(w_dff_B_uJkSSJsU0_1),.dout(w_dff_B_K6dn33Fl4_1),.clk(gclk));
	jdff dff_B_ZmREDV1C2_1(.din(w_dff_B_K6dn33Fl4_1),.dout(w_dff_B_ZmREDV1C2_1),.clk(gclk));
	jdff dff_B_wJpNu3ru1_1(.din(w_dff_B_ZmREDV1C2_1),.dout(w_dff_B_wJpNu3ru1_1),.clk(gclk));
	jdff dff_B_U6FlIi3u0_1(.din(w_dff_B_wJpNu3ru1_1),.dout(w_dff_B_U6FlIi3u0_1),.clk(gclk));
	jdff dff_B_OZaNzmmr6_1(.din(w_dff_B_U6FlIi3u0_1),.dout(w_dff_B_OZaNzmmr6_1),.clk(gclk));
	jdff dff_B_WvXoQYu74_1(.din(w_dff_B_OZaNzmmr6_1),.dout(w_dff_B_WvXoQYu74_1),.clk(gclk));
	jdff dff_B_qsB6VOwN6_1(.din(w_dff_B_WvXoQYu74_1),.dout(w_dff_B_qsB6VOwN6_1),.clk(gclk));
	jdff dff_B_yA7PwUM54_1(.din(w_dff_B_qsB6VOwN6_1),.dout(w_dff_B_yA7PwUM54_1),.clk(gclk));
	jdff dff_B_YFRm4K5W1_1(.din(w_dff_B_yA7PwUM54_1),.dout(w_dff_B_YFRm4K5W1_1),.clk(gclk));
	jdff dff_B_xBSuuJ7s4_1(.din(n530),.dout(w_dff_B_xBSuuJ7s4_1),.clk(gclk));
	jdff dff_B_k5vWgTKx4_1(.din(w_dff_B_xBSuuJ7s4_1),.dout(w_dff_B_k5vWgTKx4_1),.clk(gclk));
	jdff dff_B_y8g3ES8h6_1(.din(w_dff_B_k5vWgTKx4_1),.dout(w_dff_B_y8g3ES8h6_1),.clk(gclk));
	jdff dff_B_Tbgn4Dom7_1(.din(w_dff_B_y8g3ES8h6_1),.dout(w_dff_B_Tbgn4Dom7_1),.clk(gclk));
	jdff dff_B_BHAnsAri8_1(.din(w_dff_B_Tbgn4Dom7_1),.dout(w_dff_B_BHAnsAri8_1),.clk(gclk));
	jdff dff_B_ldS3q1HM3_1(.din(w_dff_B_BHAnsAri8_1),.dout(w_dff_B_ldS3q1HM3_1),.clk(gclk));
	jdff dff_B_we568uMK7_1(.din(w_dff_B_ldS3q1HM3_1),.dout(w_dff_B_we568uMK7_1),.clk(gclk));
	jdff dff_B_5lwAKedS5_1(.din(w_dff_B_we568uMK7_1),.dout(w_dff_B_5lwAKedS5_1),.clk(gclk));
	jdff dff_B_10IAnLPV1_1(.din(w_dff_B_5lwAKedS5_1),.dout(w_dff_B_10IAnLPV1_1),.clk(gclk));
	jdff dff_B_QDjuZ69o9_1(.din(w_dff_B_10IAnLPV1_1),.dout(w_dff_B_QDjuZ69o9_1),.clk(gclk));
	jdff dff_B_l3aIp33a0_1(.din(w_dff_B_QDjuZ69o9_1),.dout(w_dff_B_l3aIp33a0_1),.clk(gclk));
	jdff dff_B_iNzi5dWU6_1(.din(w_dff_B_l3aIp33a0_1),.dout(w_dff_B_iNzi5dWU6_1),.clk(gclk));
	jdff dff_B_E1qSF1qR7_1(.din(w_dff_B_iNzi5dWU6_1),.dout(w_dff_B_E1qSF1qR7_1),.clk(gclk));
	jdff dff_B_69kVTkT75_1(.din(w_dff_B_E1qSF1qR7_1),.dout(w_dff_B_69kVTkT75_1),.clk(gclk));
	jdff dff_B_aSayIanv6_1(.din(w_dff_B_69kVTkT75_1),.dout(w_dff_B_aSayIanv6_1),.clk(gclk));
	jdff dff_B_FyHTsubF8_1(.din(w_dff_B_aSayIanv6_1),.dout(w_dff_B_FyHTsubF8_1),.clk(gclk));
	jdff dff_B_CLzBWEe19_1(.din(w_dff_B_FyHTsubF8_1),.dout(w_dff_B_CLzBWEe19_1),.clk(gclk));
	jdff dff_B_Ocbb6EEg2_1(.din(w_dff_B_CLzBWEe19_1),.dout(w_dff_B_Ocbb6EEg2_1),.clk(gclk));
	jdff dff_B_ryUpwBpC7_1(.din(w_dff_B_Ocbb6EEg2_1),.dout(w_dff_B_ryUpwBpC7_1),.clk(gclk));
	jdff dff_B_9coZKIBA6_1(.din(w_dff_B_ryUpwBpC7_1),.dout(w_dff_B_9coZKIBA6_1),.clk(gclk));
	jdff dff_B_ndGhYzjJ7_1(.din(w_dff_B_9coZKIBA6_1),.dout(w_dff_B_ndGhYzjJ7_1),.clk(gclk));
	jdff dff_B_sMzjXJOr7_1(.din(w_dff_B_ndGhYzjJ7_1),.dout(w_dff_B_sMzjXJOr7_1),.clk(gclk));
	jdff dff_B_DGKZt9aO1_1(.din(w_dff_B_sMzjXJOr7_1),.dout(w_dff_B_DGKZt9aO1_1),.clk(gclk));
	jdff dff_B_bt0qO9ob1_1(.din(w_dff_B_DGKZt9aO1_1),.dout(w_dff_B_bt0qO9ob1_1),.clk(gclk));
	jdff dff_B_GvYmugE58_1(.din(w_dff_B_bt0qO9ob1_1),.dout(w_dff_B_GvYmugE58_1),.clk(gclk));
	jdff dff_B_Q3NRNJLN1_1(.din(w_dff_B_GvYmugE58_1),.dout(w_dff_B_Q3NRNJLN1_1),.clk(gclk));
	jdff dff_B_DgvSxp4c5_1(.din(w_dff_B_Q3NRNJLN1_1),.dout(w_dff_B_DgvSxp4c5_1),.clk(gclk));
	jdff dff_B_sX0C7uwN8_1(.din(w_dff_B_DgvSxp4c5_1),.dout(w_dff_B_sX0C7uwN8_1),.clk(gclk));
	jdff dff_B_KKdBTCpF4_1(.din(w_dff_B_sX0C7uwN8_1),.dout(w_dff_B_KKdBTCpF4_1),.clk(gclk));
	jdff dff_B_TZMF1tqX9_1(.din(w_dff_B_KKdBTCpF4_1),.dout(w_dff_B_TZMF1tqX9_1),.clk(gclk));
	jdff dff_B_J01r9X969_1(.din(w_dff_B_TZMF1tqX9_1),.dout(w_dff_B_J01r9X969_1),.clk(gclk));
	jdff dff_B_B979yd3B0_1(.din(w_dff_B_J01r9X969_1),.dout(w_dff_B_B979yd3B0_1),.clk(gclk));
	jdff dff_B_Hf4zsWZq2_1(.din(w_dff_B_B979yd3B0_1),.dout(w_dff_B_Hf4zsWZq2_1),.clk(gclk));
	jdff dff_B_vqAjp3PQ7_1(.din(n615),.dout(w_dff_B_vqAjp3PQ7_1),.clk(gclk));
	jdff dff_B_HRfTJ6D17_1(.din(w_dff_B_vqAjp3PQ7_1),.dout(w_dff_B_HRfTJ6D17_1),.clk(gclk));
	jdff dff_B_0Xqp5hgY9_1(.din(w_dff_B_HRfTJ6D17_1),.dout(w_dff_B_0Xqp5hgY9_1),.clk(gclk));
	jdff dff_B_kPTDKQsO5_1(.din(w_dff_B_0Xqp5hgY9_1),.dout(w_dff_B_kPTDKQsO5_1),.clk(gclk));
	jdff dff_B_DQxuNFZS7_1(.din(w_dff_B_kPTDKQsO5_1),.dout(w_dff_B_DQxuNFZS7_1),.clk(gclk));
	jdff dff_B_Sg8ryoas8_1(.din(w_dff_B_DQxuNFZS7_1),.dout(w_dff_B_Sg8ryoas8_1),.clk(gclk));
	jdff dff_B_L378aHdO7_1(.din(w_dff_B_Sg8ryoas8_1),.dout(w_dff_B_L378aHdO7_1),.clk(gclk));
	jdff dff_B_6qm95FkR7_1(.din(w_dff_B_L378aHdO7_1),.dout(w_dff_B_6qm95FkR7_1),.clk(gclk));
	jdff dff_B_m3tUgcO24_1(.din(w_dff_B_6qm95FkR7_1),.dout(w_dff_B_m3tUgcO24_1),.clk(gclk));
	jdff dff_B_ni4qlqbW4_1(.din(w_dff_B_m3tUgcO24_1),.dout(w_dff_B_ni4qlqbW4_1),.clk(gclk));
	jdff dff_B_TWs3YKRW4_1(.din(w_dff_B_ni4qlqbW4_1),.dout(w_dff_B_TWs3YKRW4_1),.clk(gclk));
	jdff dff_B_QaDjQRqQ7_1(.din(w_dff_B_TWs3YKRW4_1),.dout(w_dff_B_QaDjQRqQ7_1),.clk(gclk));
	jdff dff_B_tli5ftp98_1(.din(w_dff_B_QaDjQRqQ7_1),.dout(w_dff_B_tli5ftp98_1),.clk(gclk));
	jdff dff_B_unw30J9S4_1(.din(w_dff_B_tli5ftp98_1),.dout(w_dff_B_unw30J9S4_1),.clk(gclk));
	jdff dff_B_m9JW1eFQ9_1(.din(w_dff_B_unw30J9S4_1),.dout(w_dff_B_m9JW1eFQ9_1),.clk(gclk));
	jdff dff_B_rWDfYdle0_1(.din(w_dff_B_m9JW1eFQ9_1),.dout(w_dff_B_rWDfYdle0_1),.clk(gclk));
	jdff dff_B_wTGAELPA5_1(.din(w_dff_B_rWDfYdle0_1),.dout(w_dff_B_wTGAELPA5_1),.clk(gclk));
	jdff dff_B_4Qjncd7v3_1(.din(w_dff_B_wTGAELPA5_1),.dout(w_dff_B_4Qjncd7v3_1),.clk(gclk));
	jdff dff_B_DLZ0O1FA3_1(.din(w_dff_B_4Qjncd7v3_1),.dout(w_dff_B_DLZ0O1FA3_1),.clk(gclk));
	jdff dff_B_6wef0Zqj3_1(.din(w_dff_B_DLZ0O1FA3_1),.dout(w_dff_B_6wef0Zqj3_1),.clk(gclk));
	jdff dff_B_ZwYgijw02_1(.din(w_dff_B_6wef0Zqj3_1),.dout(w_dff_B_ZwYgijw02_1),.clk(gclk));
	jdff dff_B_yWI8v3Fj9_1(.din(w_dff_B_ZwYgijw02_1),.dout(w_dff_B_yWI8v3Fj9_1),.clk(gclk));
	jdff dff_B_XUlsDNFh9_1(.din(w_dff_B_yWI8v3Fj9_1),.dout(w_dff_B_XUlsDNFh9_1),.clk(gclk));
	jdff dff_B_11YpHJLM3_1(.din(w_dff_B_XUlsDNFh9_1),.dout(w_dff_B_11YpHJLM3_1),.clk(gclk));
	jdff dff_B_gJrbHuAA6_1(.din(w_dff_B_11YpHJLM3_1),.dout(w_dff_B_gJrbHuAA6_1),.clk(gclk));
	jdff dff_B_1vaIfmbv3_1(.din(w_dff_B_gJrbHuAA6_1),.dout(w_dff_B_1vaIfmbv3_1),.clk(gclk));
	jdff dff_B_EccYk7iG1_1(.din(w_dff_B_1vaIfmbv3_1),.dout(w_dff_B_EccYk7iG1_1),.clk(gclk));
	jdff dff_B_gVe4cBXl2_1(.din(w_dff_B_EccYk7iG1_1),.dout(w_dff_B_gVe4cBXl2_1),.clk(gclk));
	jdff dff_B_4YUH2rzp4_1(.din(w_dff_B_gVe4cBXl2_1),.dout(w_dff_B_4YUH2rzp4_1),.clk(gclk));
	jdff dff_B_rjAx0b5z0_1(.din(w_dff_B_4YUH2rzp4_1),.dout(w_dff_B_rjAx0b5z0_1),.clk(gclk));
	jdff dff_B_j5znD4rJ2_1(.din(w_dff_B_rjAx0b5z0_1),.dout(w_dff_B_j5znD4rJ2_1),.clk(gclk));
	jdff dff_B_xbmNtxnL2_1(.din(w_dff_B_j5znD4rJ2_1),.dout(w_dff_B_xbmNtxnL2_1),.clk(gclk));
	jdff dff_B_gdt0f4fK9_1(.din(w_dff_B_xbmNtxnL2_1),.dout(w_dff_B_gdt0f4fK9_1),.clk(gclk));
	jdff dff_B_0EksrcoX7_1(.din(w_dff_B_gdt0f4fK9_1),.dout(w_dff_B_0EksrcoX7_1),.clk(gclk));
	jdff dff_B_P8QCH00j3_1(.din(w_dff_B_0EksrcoX7_1),.dout(w_dff_B_P8QCH00j3_1),.clk(gclk));
	jdff dff_B_OLxsTluA8_1(.din(w_dff_B_P8QCH00j3_1),.dout(w_dff_B_OLxsTluA8_1),.clk(gclk));
	jdff dff_B_zPxi1Q6c6_1(.din(n707),.dout(w_dff_B_zPxi1Q6c6_1),.clk(gclk));
	jdff dff_B_1R5NIVMX4_1(.din(w_dff_B_zPxi1Q6c6_1),.dout(w_dff_B_1R5NIVMX4_1),.clk(gclk));
	jdff dff_B_CBGfoSOi5_1(.din(w_dff_B_1R5NIVMX4_1),.dout(w_dff_B_CBGfoSOi5_1),.clk(gclk));
	jdff dff_B_MSn1eXOV3_1(.din(w_dff_B_CBGfoSOi5_1),.dout(w_dff_B_MSn1eXOV3_1),.clk(gclk));
	jdff dff_B_w2aUY5463_1(.din(w_dff_B_MSn1eXOV3_1),.dout(w_dff_B_w2aUY5463_1),.clk(gclk));
	jdff dff_B_yKWRbLQF0_1(.din(w_dff_B_w2aUY5463_1),.dout(w_dff_B_yKWRbLQF0_1),.clk(gclk));
	jdff dff_B_lMS2eIjt1_1(.din(w_dff_B_yKWRbLQF0_1),.dout(w_dff_B_lMS2eIjt1_1),.clk(gclk));
	jdff dff_B_DywTu1qP2_1(.din(w_dff_B_lMS2eIjt1_1),.dout(w_dff_B_DywTu1qP2_1),.clk(gclk));
	jdff dff_B_XXN3uC1g4_1(.din(w_dff_B_DywTu1qP2_1),.dout(w_dff_B_XXN3uC1g4_1),.clk(gclk));
	jdff dff_B_TLdhMHVW7_1(.din(w_dff_B_XXN3uC1g4_1),.dout(w_dff_B_TLdhMHVW7_1),.clk(gclk));
	jdff dff_B_Rg8nneRf0_1(.din(w_dff_B_TLdhMHVW7_1),.dout(w_dff_B_Rg8nneRf0_1),.clk(gclk));
	jdff dff_B_nOjWZ9wV7_1(.din(w_dff_B_Rg8nneRf0_1),.dout(w_dff_B_nOjWZ9wV7_1),.clk(gclk));
	jdff dff_B_dpM7eu7c6_1(.din(w_dff_B_nOjWZ9wV7_1),.dout(w_dff_B_dpM7eu7c6_1),.clk(gclk));
	jdff dff_B_Rt0HQJTD1_1(.din(w_dff_B_dpM7eu7c6_1),.dout(w_dff_B_Rt0HQJTD1_1),.clk(gclk));
	jdff dff_B_hBBOq6Yx8_1(.din(w_dff_B_Rt0HQJTD1_1),.dout(w_dff_B_hBBOq6Yx8_1),.clk(gclk));
	jdff dff_B_jtsEMNWB4_1(.din(w_dff_B_hBBOq6Yx8_1),.dout(w_dff_B_jtsEMNWB4_1),.clk(gclk));
	jdff dff_B_HiLQJmiD4_1(.din(w_dff_B_jtsEMNWB4_1),.dout(w_dff_B_HiLQJmiD4_1),.clk(gclk));
	jdff dff_B_Z3o7y1ZP7_1(.din(w_dff_B_HiLQJmiD4_1),.dout(w_dff_B_Z3o7y1ZP7_1),.clk(gclk));
	jdff dff_B_awLXZavE6_1(.din(w_dff_B_Z3o7y1ZP7_1),.dout(w_dff_B_awLXZavE6_1),.clk(gclk));
	jdff dff_B_g7tV1r0n6_1(.din(w_dff_B_awLXZavE6_1),.dout(w_dff_B_g7tV1r0n6_1),.clk(gclk));
	jdff dff_B_78v9h3AL5_1(.din(w_dff_B_g7tV1r0n6_1),.dout(w_dff_B_78v9h3AL5_1),.clk(gclk));
	jdff dff_B_cuAE0DiZ0_1(.din(w_dff_B_78v9h3AL5_1),.dout(w_dff_B_cuAE0DiZ0_1),.clk(gclk));
	jdff dff_B_VURBNHcq7_1(.din(w_dff_B_cuAE0DiZ0_1),.dout(w_dff_B_VURBNHcq7_1),.clk(gclk));
	jdff dff_B_Kbu1jCJ97_1(.din(w_dff_B_VURBNHcq7_1),.dout(w_dff_B_Kbu1jCJ97_1),.clk(gclk));
	jdff dff_B_VXsNt6IB4_1(.din(w_dff_B_Kbu1jCJ97_1),.dout(w_dff_B_VXsNt6IB4_1),.clk(gclk));
	jdff dff_B_KmcaORtk9_1(.din(w_dff_B_VXsNt6IB4_1),.dout(w_dff_B_KmcaORtk9_1),.clk(gclk));
	jdff dff_B_VoATBfvH2_1(.din(w_dff_B_KmcaORtk9_1),.dout(w_dff_B_VoATBfvH2_1),.clk(gclk));
	jdff dff_B_fc5rMa0k5_1(.din(w_dff_B_VoATBfvH2_1),.dout(w_dff_B_fc5rMa0k5_1),.clk(gclk));
	jdff dff_B_ifhE0vC63_1(.din(w_dff_B_fc5rMa0k5_1),.dout(w_dff_B_ifhE0vC63_1),.clk(gclk));
	jdff dff_B_H46xCC9P7_1(.din(w_dff_B_ifhE0vC63_1),.dout(w_dff_B_H46xCC9P7_1),.clk(gclk));
	jdff dff_B_07yO4O7s1_1(.din(w_dff_B_H46xCC9P7_1),.dout(w_dff_B_07yO4O7s1_1),.clk(gclk));
	jdff dff_B_Iplt7siZ5_1(.din(w_dff_B_07yO4O7s1_1),.dout(w_dff_B_Iplt7siZ5_1),.clk(gclk));
	jdff dff_B_7XKU0PZ66_1(.din(w_dff_B_Iplt7siZ5_1),.dout(w_dff_B_7XKU0PZ66_1),.clk(gclk));
	jdff dff_B_50E9cy6U7_1(.din(w_dff_B_7XKU0PZ66_1),.dout(w_dff_B_50E9cy6U7_1),.clk(gclk));
	jdff dff_B_oPcfGX5r3_1(.din(w_dff_B_50E9cy6U7_1),.dout(w_dff_B_oPcfGX5r3_1),.clk(gclk));
	jdff dff_B_6Y6UIDei8_1(.din(w_dff_B_oPcfGX5r3_1),.dout(w_dff_B_6Y6UIDei8_1),.clk(gclk));
	jdff dff_B_fT11e3pk3_1(.din(w_dff_B_6Y6UIDei8_1),.dout(w_dff_B_fT11e3pk3_1),.clk(gclk));
	jdff dff_B_7Isxlngi2_1(.din(w_dff_B_fT11e3pk3_1),.dout(w_dff_B_7Isxlngi2_1),.clk(gclk));
	jdff dff_B_aIJIHk8U5_1(.din(w_dff_B_7Isxlngi2_1),.dout(w_dff_B_aIJIHk8U5_1),.clk(gclk));
	jdff dff_B_eUIL5prO2_1(.din(n806),.dout(w_dff_B_eUIL5prO2_1),.clk(gclk));
	jdff dff_B_zsdwqWWC6_1(.din(w_dff_B_eUIL5prO2_1),.dout(w_dff_B_zsdwqWWC6_1),.clk(gclk));
	jdff dff_B_AC70GyfJ3_1(.din(w_dff_B_zsdwqWWC6_1),.dout(w_dff_B_AC70GyfJ3_1),.clk(gclk));
	jdff dff_B_EQgIEvn86_1(.din(w_dff_B_AC70GyfJ3_1),.dout(w_dff_B_EQgIEvn86_1),.clk(gclk));
	jdff dff_B_1pt4iQjB0_1(.din(w_dff_B_EQgIEvn86_1),.dout(w_dff_B_1pt4iQjB0_1),.clk(gclk));
	jdff dff_B_5twYTAM69_1(.din(w_dff_B_1pt4iQjB0_1),.dout(w_dff_B_5twYTAM69_1),.clk(gclk));
	jdff dff_B_XvMQT9Em7_1(.din(w_dff_B_5twYTAM69_1),.dout(w_dff_B_XvMQT9Em7_1),.clk(gclk));
	jdff dff_B_oXsLUE7i9_1(.din(w_dff_B_XvMQT9Em7_1),.dout(w_dff_B_oXsLUE7i9_1),.clk(gclk));
	jdff dff_B_5Aqb1Bcf7_1(.din(w_dff_B_oXsLUE7i9_1),.dout(w_dff_B_5Aqb1Bcf7_1),.clk(gclk));
	jdff dff_B_3YEZUXHr3_1(.din(w_dff_B_5Aqb1Bcf7_1),.dout(w_dff_B_3YEZUXHr3_1),.clk(gclk));
	jdff dff_B_dN4Gl2Bi3_1(.din(w_dff_B_3YEZUXHr3_1),.dout(w_dff_B_dN4Gl2Bi3_1),.clk(gclk));
	jdff dff_B_v4on7eZH4_1(.din(w_dff_B_dN4Gl2Bi3_1),.dout(w_dff_B_v4on7eZH4_1),.clk(gclk));
	jdff dff_B_lvLwZhrU5_1(.din(w_dff_B_v4on7eZH4_1),.dout(w_dff_B_lvLwZhrU5_1),.clk(gclk));
	jdff dff_B_z2ltMgUF8_1(.din(w_dff_B_lvLwZhrU5_1),.dout(w_dff_B_z2ltMgUF8_1),.clk(gclk));
	jdff dff_B_eaYUr7tn3_1(.din(w_dff_B_z2ltMgUF8_1),.dout(w_dff_B_eaYUr7tn3_1),.clk(gclk));
	jdff dff_B_wjJ96IPJ7_1(.din(w_dff_B_eaYUr7tn3_1),.dout(w_dff_B_wjJ96IPJ7_1),.clk(gclk));
	jdff dff_B_PHAmY9oJ3_1(.din(w_dff_B_wjJ96IPJ7_1),.dout(w_dff_B_PHAmY9oJ3_1),.clk(gclk));
	jdff dff_B_FFOYMaYX7_1(.din(w_dff_B_PHAmY9oJ3_1),.dout(w_dff_B_FFOYMaYX7_1),.clk(gclk));
	jdff dff_B_OSzyPwEm5_1(.din(w_dff_B_FFOYMaYX7_1),.dout(w_dff_B_OSzyPwEm5_1),.clk(gclk));
	jdff dff_B_vLcq54tm9_1(.din(w_dff_B_OSzyPwEm5_1),.dout(w_dff_B_vLcq54tm9_1),.clk(gclk));
	jdff dff_B_uNChc3vM8_1(.din(w_dff_B_vLcq54tm9_1),.dout(w_dff_B_uNChc3vM8_1),.clk(gclk));
	jdff dff_B_Yn94UJfX5_1(.din(w_dff_B_uNChc3vM8_1),.dout(w_dff_B_Yn94UJfX5_1),.clk(gclk));
	jdff dff_B_GfkLe7Pa2_1(.din(w_dff_B_Yn94UJfX5_1),.dout(w_dff_B_GfkLe7Pa2_1),.clk(gclk));
	jdff dff_B_q6t8fYaQ5_1(.din(w_dff_B_GfkLe7Pa2_1),.dout(w_dff_B_q6t8fYaQ5_1),.clk(gclk));
	jdff dff_B_DcliMkSo5_1(.din(w_dff_B_q6t8fYaQ5_1),.dout(w_dff_B_DcliMkSo5_1),.clk(gclk));
	jdff dff_B_Sz4aXa4Y8_1(.din(w_dff_B_DcliMkSo5_1),.dout(w_dff_B_Sz4aXa4Y8_1),.clk(gclk));
	jdff dff_B_ygdhXT930_1(.din(w_dff_B_Sz4aXa4Y8_1),.dout(w_dff_B_ygdhXT930_1),.clk(gclk));
	jdff dff_B_FWnZsOR52_1(.din(w_dff_B_ygdhXT930_1),.dout(w_dff_B_FWnZsOR52_1),.clk(gclk));
	jdff dff_B_lNEgrRaH7_1(.din(w_dff_B_FWnZsOR52_1),.dout(w_dff_B_lNEgrRaH7_1),.clk(gclk));
	jdff dff_B_QbtBYitR4_1(.din(w_dff_B_lNEgrRaH7_1),.dout(w_dff_B_QbtBYitR4_1),.clk(gclk));
	jdff dff_B_iwwBkjQF1_1(.din(w_dff_B_QbtBYitR4_1),.dout(w_dff_B_iwwBkjQF1_1),.clk(gclk));
	jdff dff_B_VZFVd6Eo0_1(.din(w_dff_B_iwwBkjQF1_1),.dout(w_dff_B_VZFVd6Eo0_1),.clk(gclk));
	jdff dff_B_A9yPP5Ju7_1(.din(w_dff_B_VZFVd6Eo0_1),.dout(w_dff_B_A9yPP5Ju7_1),.clk(gclk));
	jdff dff_B_4xBDN4SN7_1(.din(w_dff_B_A9yPP5Ju7_1),.dout(w_dff_B_4xBDN4SN7_1),.clk(gclk));
	jdff dff_B_wGcbOP2r4_1(.din(w_dff_B_4xBDN4SN7_1),.dout(w_dff_B_wGcbOP2r4_1),.clk(gclk));
	jdff dff_B_UibN8WY33_1(.din(w_dff_B_wGcbOP2r4_1),.dout(w_dff_B_UibN8WY33_1),.clk(gclk));
	jdff dff_B_WhludnsO2_1(.din(w_dff_B_UibN8WY33_1),.dout(w_dff_B_WhludnsO2_1),.clk(gclk));
	jdff dff_B_kXwV66Zz5_1(.din(w_dff_B_WhludnsO2_1),.dout(w_dff_B_kXwV66Zz5_1),.clk(gclk));
	jdff dff_B_nWxQvpep3_1(.din(w_dff_B_kXwV66Zz5_1),.dout(w_dff_B_nWxQvpep3_1),.clk(gclk));
	jdff dff_B_5xaIIYPo2_1(.din(w_dff_B_nWxQvpep3_1),.dout(w_dff_B_5xaIIYPo2_1),.clk(gclk));
	jdff dff_B_HN3mt3dj6_1(.din(w_dff_B_5xaIIYPo2_1),.dout(w_dff_B_HN3mt3dj6_1),.clk(gclk));
	jdff dff_B_8uvPJXgT8_1(.din(w_dff_B_HN3mt3dj6_1),.dout(w_dff_B_8uvPJXgT8_1),.clk(gclk));
	jdff dff_B_4SLee9TS5_0(.din(n1296),.dout(w_dff_B_4SLee9TS5_0),.clk(gclk));
	jdff dff_B_fUcCcxHo9_1(.din(n1811),.dout(w_dff_B_fUcCcxHo9_1),.clk(gclk));
	jdff dff_B_Bhe9K82J7_1(.din(w_dff_B_fUcCcxHo9_1),.dout(w_dff_B_Bhe9K82J7_1),.clk(gclk));
	jdff dff_B_dKSVDGQp3_1(.din(w_dff_B_Bhe9K82J7_1),.dout(w_dff_B_dKSVDGQp3_1),.clk(gclk));
	jdff dff_B_yANjRof44_1(.din(w_dff_B_dKSVDGQp3_1),.dout(w_dff_B_yANjRof44_1),.clk(gclk));
	jdff dff_B_Q8RpNch32_1(.din(w_dff_B_yANjRof44_1),.dout(w_dff_B_Q8RpNch32_1),.clk(gclk));
	jdff dff_B_I7XTI24x6_1(.din(w_dff_B_Q8RpNch32_1),.dout(w_dff_B_I7XTI24x6_1),.clk(gclk));
	jdff dff_B_Q6uIvwn59_1(.din(w_dff_B_I7XTI24x6_1),.dout(w_dff_B_Q6uIvwn59_1),.clk(gclk));
	jdff dff_B_LVUkFt7i7_1(.din(w_dff_B_Q6uIvwn59_1),.dout(w_dff_B_LVUkFt7i7_1),.clk(gclk));
	jdff dff_B_BS0EEH3O9_1(.din(w_dff_B_LVUkFt7i7_1),.dout(w_dff_B_BS0EEH3O9_1),.clk(gclk));
	jdff dff_B_YnSBBg2P9_1(.din(w_dff_B_BS0EEH3O9_1),.dout(w_dff_B_YnSBBg2P9_1),.clk(gclk));
	jdff dff_B_gUyNrNT92_1(.din(w_dff_B_YnSBBg2P9_1),.dout(w_dff_B_gUyNrNT92_1),.clk(gclk));
	jdff dff_B_D2xwiLSQ8_1(.din(w_dff_B_gUyNrNT92_1),.dout(w_dff_B_D2xwiLSQ8_1),.clk(gclk));
	jdff dff_B_tpT1tXET2_1(.din(w_dff_B_D2xwiLSQ8_1),.dout(w_dff_B_tpT1tXET2_1),.clk(gclk));
	jdff dff_B_eSzynpin2_1(.din(w_dff_B_tpT1tXET2_1),.dout(w_dff_B_eSzynpin2_1),.clk(gclk));
	jdff dff_B_DRCwA28l1_1(.din(w_dff_B_eSzynpin2_1),.dout(w_dff_B_DRCwA28l1_1),.clk(gclk));
	jdff dff_B_mhfjPYd78_0(.din(n1819),.dout(w_dff_B_mhfjPYd78_0),.clk(gclk));
	jdff dff_B_EKGU0wum5_0(.din(w_dff_B_mhfjPYd78_0),.dout(w_dff_B_EKGU0wum5_0),.clk(gclk));
	jdff dff_B_HeNgJGVL0_0(.din(w_dff_B_EKGU0wum5_0),.dout(w_dff_B_HeNgJGVL0_0),.clk(gclk));
	jdff dff_B_UfuBytbQ2_0(.din(w_dff_B_HeNgJGVL0_0),.dout(w_dff_B_UfuBytbQ2_0),.clk(gclk));
	jdff dff_B_KnsOjQ7V5_0(.din(w_dff_B_UfuBytbQ2_0),.dout(w_dff_B_KnsOjQ7V5_0),.clk(gclk));
	jdff dff_B_niyCTkNf7_0(.din(w_dff_B_KnsOjQ7V5_0),.dout(w_dff_B_niyCTkNf7_0),.clk(gclk));
	jdff dff_B_2MIJS98l9_0(.din(w_dff_B_niyCTkNf7_0),.dout(w_dff_B_2MIJS98l9_0),.clk(gclk));
	jdff dff_B_odXVTPrx9_0(.din(w_dff_B_2MIJS98l9_0),.dout(w_dff_B_odXVTPrx9_0),.clk(gclk));
	jdff dff_B_SKacsID54_0(.din(w_dff_B_odXVTPrx9_0),.dout(w_dff_B_SKacsID54_0),.clk(gclk));
	jdff dff_B_2kJjINXo9_0(.din(w_dff_B_SKacsID54_0),.dout(w_dff_B_2kJjINXo9_0),.clk(gclk));
	jdff dff_B_2zAr0Qx19_0(.din(w_dff_B_2kJjINXo9_0),.dout(w_dff_B_2zAr0Qx19_0),.clk(gclk));
	jdff dff_B_f7C5wsGT2_0(.din(w_dff_B_2zAr0Qx19_0),.dout(w_dff_B_f7C5wsGT2_0),.clk(gclk));
	jdff dff_B_JaAxITgE4_0(.din(w_dff_B_f7C5wsGT2_0),.dout(w_dff_B_JaAxITgE4_0),.clk(gclk));
	jdff dff_A_rT3HLtX14_0(.dout(w_n1818_0[0]),.din(w_dff_A_rT3HLtX14_0),.clk(gclk));
	jdff dff_A_47l8Pkz52_0(.dout(w_dff_A_rT3HLtX14_0),.din(w_dff_A_47l8Pkz52_0),.clk(gclk));
	jdff dff_A_V2w1ap1I2_0(.dout(w_dff_A_47l8Pkz52_0),.din(w_dff_A_V2w1ap1I2_0),.clk(gclk));
	jdff dff_A_5Z5zWbGP6_0(.dout(w_dff_A_V2w1ap1I2_0),.din(w_dff_A_5Z5zWbGP6_0),.clk(gclk));
	jdff dff_A_XSpZLn2a6_0(.dout(w_dff_A_5Z5zWbGP6_0),.din(w_dff_A_XSpZLn2a6_0),.clk(gclk));
	jdff dff_A_VjqPeLEa6_0(.dout(w_dff_A_XSpZLn2a6_0),.din(w_dff_A_VjqPeLEa6_0),.clk(gclk));
	jdff dff_A_dzr5DIwN6_0(.dout(w_dff_A_VjqPeLEa6_0),.din(w_dff_A_dzr5DIwN6_0),.clk(gclk));
	jdff dff_A_WcFhi0pj7_0(.dout(w_dff_A_dzr5DIwN6_0),.din(w_dff_A_WcFhi0pj7_0),.clk(gclk));
	jdff dff_A_MC3QqYvh8_0(.dout(w_dff_A_WcFhi0pj7_0),.din(w_dff_A_MC3QqYvh8_0),.clk(gclk));
	jdff dff_A_ThkRr3Hp4_0(.dout(w_dff_A_MC3QqYvh8_0),.din(w_dff_A_ThkRr3Hp4_0),.clk(gclk));
	jdff dff_A_r6U5jSWR8_0(.dout(w_dff_A_ThkRr3Hp4_0),.din(w_dff_A_r6U5jSWR8_0),.clk(gclk));
	jdff dff_A_QHohHitX3_0(.dout(w_dff_A_r6U5jSWR8_0),.din(w_dff_A_QHohHitX3_0),.clk(gclk));
	jdff dff_A_eFMJw3St7_0(.dout(w_dff_A_QHohHitX3_0),.din(w_dff_A_eFMJw3St7_0),.clk(gclk));
	jdff dff_A_MML1jZwp4_0(.dout(w_dff_A_eFMJw3St7_0),.din(w_dff_A_MML1jZwp4_0),.clk(gclk));
	jdff dff_B_6Ux8M5LD0_1(.din(n1808),.dout(w_dff_B_6Ux8M5LD0_1),.clk(gclk));
	jdff dff_B_iEasrwnB9_1(.din(w_dff_B_6Ux8M5LD0_1),.dout(w_dff_B_iEasrwnB9_1),.clk(gclk));
	jdff dff_B_uFHBApah4_2(.din(n1807),.dout(w_dff_B_uFHBApah4_2),.clk(gclk));
	jdff dff_B_zCckU8lI1_2(.din(w_dff_B_uFHBApah4_2),.dout(w_dff_B_zCckU8lI1_2),.clk(gclk));
	jdff dff_B_4z105Ir07_2(.din(w_dff_B_zCckU8lI1_2),.dout(w_dff_B_4z105Ir07_2),.clk(gclk));
	jdff dff_B_Usdx7tpg4_2(.din(w_dff_B_4z105Ir07_2),.dout(w_dff_B_Usdx7tpg4_2),.clk(gclk));
	jdff dff_B_WGatuEiZ4_2(.din(w_dff_B_Usdx7tpg4_2),.dout(w_dff_B_WGatuEiZ4_2),.clk(gclk));
	jdff dff_B_BKypBA0d3_2(.din(w_dff_B_WGatuEiZ4_2),.dout(w_dff_B_BKypBA0d3_2),.clk(gclk));
	jdff dff_B_BelfP1WG7_2(.din(w_dff_B_BKypBA0d3_2),.dout(w_dff_B_BelfP1WG7_2),.clk(gclk));
	jdff dff_B_AoPnHSzj8_2(.din(w_dff_B_BelfP1WG7_2),.dout(w_dff_B_AoPnHSzj8_2),.clk(gclk));
	jdff dff_B_PzrcveSQ6_2(.din(w_dff_B_AoPnHSzj8_2),.dout(w_dff_B_PzrcveSQ6_2),.clk(gclk));
	jdff dff_B_zM4gup2S2_2(.din(w_dff_B_PzrcveSQ6_2),.dout(w_dff_B_zM4gup2S2_2),.clk(gclk));
	jdff dff_B_HkVPkxYu2_2(.din(w_dff_B_zM4gup2S2_2),.dout(w_dff_B_HkVPkxYu2_2),.clk(gclk));
	jdff dff_B_NrT46Yvb7_2(.din(w_dff_B_HkVPkxYu2_2),.dout(w_dff_B_NrT46Yvb7_2),.clk(gclk));
	jdff dff_B_wUhfrYwx9_2(.din(w_dff_B_NrT46Yvb7_2),.dout(w_dff_B_wUhfrYwx9_2),.clk(gclk));
	jdff dff_B_tR94esYr2_2(.din(w_dff_B_wUhfrYwx9_2),.dout(w_dff_B_tR94esYr2_2),.clk(gclk));
	jdff dff_B_2RxmWKIM2_2(.din(w_dff_B_tR94esYr2_2),.dout(w_dff_B_2RxmWKIM2_2),.clk(gclk));
	jdff dff_B_nlj7rfPb3_2(.din(w_dff_B_2RxmWKIM2_2),.dout(w_dff_B_nlj7rfPb3_2),.clk(gclk));
	jdff dff_B_9UJyqb441_2(.din(w_dff_B_nlj7rfPb3_2),.dout(w_dff_B_9UJyqb441_2),.clk(gclk));
	jdff dff_B_Olh2PG0B5_2(.din(w_dff_B_9UJyqb441_2),.dout(w_dff_B_Olh2PG0B5_2),.clk(gclk));
	jdff dff_B_D9t3yHs04_2(.din(w_dff_B_Olh2PG0B5_2),.dout(w_dff_B_D9t3yHs04_2),.clk(gclk));
	jdff dff_B_o4tY4MSg9_2(.din(w_dff_B_D9t3yHs04_2),.dout(w_dff_B_o4tY4MSg9_2),.clk(gclk));
	jdff dff_B_Q6QhPzwv5_2(.din(w_dff_B_o4tY4MSg9_2),.dout(w_dff_B_Q6QhPzwv5_2),.clk(gclk));
	jdff dff_B_CWMSSikA9_2(.din(w_dff_B_Q6QhPzwv5_2),.dout(w_dff_B_CWMSSikA9_2),.clk(gclk));
	jdff dff_B_Rvw2hzp05_2(.din(w_dff_B_CWMSSikA9_2),.dout(w_dff_B_Rvw2hzp05_2),.clk(gclk));
	jdff dff_B_xsjw2vsm1_2(.din(w_dff_B_Rvw2hzp05_2),.dout(w_dff_B_xsjw2vsm1_2),.clk(gclk));
	jdff dff_B_1ww1o8PK8_2(.din(w_dff_B_xsjw2vsm1_2),.dout(w_dff_B_1ww1o8PK8_2),.clk(gclk));
	jdff dff_B_FGEbX3AC1_2(.din(w_dff_B_1ww1o8PK8_2),.dout(w_dff_B_FGEbX3AC1_2),.clk(gclk));
	jdff dff_B_pycMZsDz7_2(.din(w_dff_B_FGEbX3AC1_2),.dout(w_dff_B_pycMZsDz7_2),.clk(gclk));
	jdff dff_B_64JZRsGy3_2(.din(w_dff_B_pycMZsDz7_2),.dout(w_dff_B_64JZRsGy3_2),.clk(gclk));
	jdff dff_B_cwNudo3v4_2(.din(w_dff_B_64JZRsGy3_2),.dout(w_dff_B_cwNudo3v4_2),.clk(gclk));
	jdff dff_B_PH20KCtK0_2(.din(w_dff_B_cwNudo3v4_2),.dout(w_dff_B_PH20KCtK0_2),.clk(gclk));
	jdff dff_B_qOJ7SaTp7_2(.din(w_dff_B_PH20KCtK0_2),.dout(w_dff_B_qOJ7SaTp7_2),.clk(gclk));
	jdff dff_B_nl4spyBO7_2(.din(w_dff_B_qOJ7SaTp7_2),.dout(w_dff_B_nl4spyBO7_2),.clk(gclk));
	jdff dff_B_CZvtNbY69_2(.din(w_dff_B_nl4spyBO7_2),.dout(w_dff_B_CZvtNbY69_2),.clk(gclk));
	jdff dff_B_6mIumRbI5_2(.din(w_dff_B_CZvtNbY69_2),.dout(w_dff_B_6mIumRbI5_2),.clk(gclk));
	jdff dff_B_NogpHkaB5_2(.din(w_dff_B_6mIumRbI5_2),.dout(w_dff_B_NogpHkaB5_2),.clk(gclk));
	jdff dff_B_EFfczy0S8_2(.din(w_dff_B_NogpHkaB5_2),.dout(w_dff_B_EFfczy0S8_2),.clk(gclk));
	jdff dff_B_4WCADZEa8_2(.din(w_dff_B_EFfczy0S8_2),.dout(w_dff_B_4WCADZEa8_2),.clk(gclk));
	jdff dff_B_uNtaOoeT3_2(.din(w_dff_B_4WCADZEa8_2),.dout(w_dff_B_uNtaOoeT3_2),.clk(gclk));
	jdff dff_B_OGu9jeuz7_2(.din(w_dff_B_uNtaOoeT3_2),.dout(w_dff_B_OGu9jeuz7_2),.clk(gclk));
	jdff dff_B_kM0ArLr20_2(.din(w_dff_B_OGu9jeuz7_2),.dout(w_dff_B_kM0ArLr20_2),.clk(gclk));
	jdff dff_B_OtppCZaK9_2(.din(w_dff_B_kM0ArLr20_2),.dout(w_dff_B_OtppCZaK9_2),.clk(gclk));
	jdff dff_B_ruoBLLGk4_2(.din(w_dff_B_OtppCZaK9_2),.dout(w_dff_B_ruoBLLGk4_2),.clk(gclk));
	jdff dff_B_Dhiqr7bm1_2(.din(w_dff_B_ruoBLLGk4_2),.dout(w_dff_B_Dhiqr7bm1_2),.clk(gclk));
	jdff dff_B_5ZeXVluX2_2(.din(w_dff_B_Dhiqr7bm1_2),.dout(w_dff_B_5ZeXVluX2_2),.clk(gclk));
	jdff dff_B_x0q1LzIb6_2(.din(w_dff_B_5ZeXVluX2_2),.dout(w_dff_B_x0q1LzIb6_2),.clk(gclk));
	jdff dff_B_qwAzB6TL7_2(.din(w_dff_B_x0q1LzIb6_2),.dout(w_dff_B_qwAzB6TL7_2),.clk(gclk));
	jdff dff_B_ZH0Ny7Zg1_2(.din(w_dff_B_qwAzB6TL7_2),.dout(w_dff_B_ZH0Ny7Zg1_2),.clk(gclk));
	jdff dff_B_pH7VgZtv2_2(.din(w_dff_B_ZH0Ny7Zg1_2),.dout(w_dff_B_pH7VgZtv2_2),.clk(gclk));
	jdff dff_B_r4thXlzw5_2(.din(w_dff_B_pH7VgZtv2_2),.dout(w_dff_B_r4thXlzw5_2),.clk(gclk));
	jdff dff_B_urnONHy72_2(.din(w_dff_B_r4thXlzw5_2),.dout(w_dff_B_urnONHy72_2),.clk(gclk));
	jdff dff_B_nqeiPldB3_2(.din(w_dff_B_urnONHy72_2),.dout(w_dff_B_nqeiPldB3_2),.clk(gclk));
	jdff dff_B_wMGJ46wb7_2(.din(w_dff_B_nqeiPldB3_2),.dout(w_dff_B_wMGJ46wb7_2),.clk(gclk));
	jdff dff_B_9ldd8rqJ0_2(.din(w_dff_B_wMGJ46wb7_2),.dout(w_dff_B_9ldd8rqJ0_2),.clk(gclk));
	jdff dff_B_zTSUg7Xy3_2(.din(w_dff_B_9ldd8rqJ0_2),.dout(w_dff_B_zTSUg7Xy3_2),.clk(gclk));
	jdff dff_B_4885EH6h0_2(.din(w_dff_B_zTSUg7Xy3_2),.dout(w_dff_B_4885EH6h0_2),.clk(gclk));
	jdff dff_B_6pA5vqom0_2(.din(w_dff_B_4885EH6h0_2),.dout(w_dff_B_6pA5vqom0_2),.clk(gclk));
	jdff dff_B_lqpZejf25_2(.din(w_dff_B_6pA5vqom0_2),.dout(w_dff_B_lqpZejf25_2),.clk(gclk));
	jdff dff_B_wlAl6BB07_1(.din(n1814),.dout(w_dff_B_wlAl6BB07_1),.clk(gclk));
	jdff dff_B_YOnoyAXq1_1(.din(w_dff_B_wlAl6BB07_1),.dout(w_dff_B_YOnoyAXq1_1),.clk(gclk));
	jdff dff_B_MQVTQO0r6_1(.din(w_dff_B_YOnoyAXq1_1),.dout(w_dff_B_MQVTQO0r6_1),.clk(gclk));
	jdff dff_B_hMxpTDQX0_1(.din(w_dff_B_MQVTQO0r6_1),.dout(w_dff_B_hMxpTDQX0_1),.clk(gclk));
	jdff dff_B_oNFhpEqu3_1(.din(w_dff_B_hMxpTDQX0_1),.dout(w_dff_B_oNFhpEqu3_1),.clk(gclk));
	jdff dff_B_8BhzC5nv3_1(.din(w_dff_B_oNFhpEqu3_1),.dout(w_dff_B_8BhzC5nv3_1),.clk(gclk));
	jdff dff_B_D15VyJj03_1(.din(w_dff_B_8BhzC5nv3_1),.dout(w_dff_B_D15VyJj03_1),.clk(gclk));
	jdff dff_B_PQNzjg0H5_1(.din(w_dff_B_D15VyJj03_1),.dout(w_dff_B_PQNzjg0H5_1),.clk(gclk));
	jdff dff_B_oQ1WeUbe0_1(.din(w_dff_B_PQNzjg0H5_1),.dout(w_dff_B_oQ1WeUbe0_1),.clk(gclk));
	jdff dff_B_hnCaVgjP7_1(.din(w_dff_B_oQ1WeUbe0_1),.dout(w_dff_B_hnCaVgjP7_1),.clk(gclk));
	jdff dff_B_nK2CbcYs4_1(.din(w_dff_B_hnCaVgjP7_1),.dout(w_dff_B_nK2CbcYs4_1),.clk(gclk));
	jdff dff_B_vdbemxIZ8_1(.din(w_dff_B_nK2CbcYs4_1),.dout(w_dff_B_vdbemxIZ8_1),.clk(gclk));
	jdff dff_B_c6XrcEjR7_1(.din(w_dff_B_vdbemxIZ8_1),.dout(w_dff_B_c6XrcEjR7_1),.clk(gclk));
	jdff dff_B_GobpxdEP5_0(.din(n1815),.dout(w_dff_B_GobpxdEP5_0),.clk(gclk));
	jdff dff_B_xfahLXTG1_0(.din(w_dff_B_GobpxdEP5_0),.dout(w_dff_B_xfahLXTG1_0),.clk(gclk));
	jdff dff_B_mo2Mm79I4_0(.din(w_dff_B_xfahLXTG1_0),.dout(w_dff_B_mo2Mm79I4_0),.clk(gclk));
	jdff dff_B_clHexbmH9_0(.din(w_dff_B_mo2Mm79I4_0),.dout(w_dff_B_clHexbmH9_0),.clk(gclk));
	jdff dff_B_7ChBB2AN8_0(.din(w_dff_B_clHexbmH9_0),.dout(w_dff_B_7ChBB2AN8_0),.clk(gclk));
	jdff dff_B_KABMMdis3_0(.din(w_dff_B_7ChBB2AN8_0),.dout(w_dff_B_KABMMdis3_0),.clk(gclk));
	jdff dff_B_04JWzxSZ9_0(.din(w_dff_B_KABMMdis3_0),.dout(w_dff_B_04JWzxSZ9_0),.clk(gclk));
	jdff dff_B_4wWzOLQK1_0(.din(w_dff_B_04JWzxSZ9_0),.dout(w_dff_B_4wWzOLQK1_0),.clk(gclk));
	jdff dff_B_BrDt18yw5_0(.din(w_dff_B_4wWzOLQK1_0),.dout(w_dff_B_BrDt18yw5_0),.clk(gclk));
	jdff dff_B_4k14NuXX3_0(.din(w_dff_B_BrDt18yw5_0),.dout(w_dff_B_4k14NuXX3_0),.clk(gclk));
	jdff dff_B_MEBU3MHh5_0(.din(w_dff_B_4k14NuXX3_0),.dout(w_dff_B_MEBU3MHh5_0),.clk(gclk));
	jdff dff_B_Zgspq9E55_0(.din(w_dff_B_MEBU3MHh5_0),.dout(w_dff_B_Zgspq9E55_0),.clk(gclk));
	jdff dff_A_crPSyuO82_1(.dout(w_n1805_0[1]),.din(w_dff_A_crPSyuO82_1),.clk(gclk));
	jdff dff_A_WKuPtrmB4_1(.dout(w_dff_A_crPSyuO82_1),.din(w_dff_A_WKuPtrmB4_1),.clk(gclk));
	jdff dff_A_Zuk5bBdR2_1(.dout(w_dff_A_WKuPtrmB4_1),.din(w_dff_A_Zuk5bBdR2_1),.clk(gclk));
	jdff dff_A_XmdMQl875_1(.dout(w_dff_A_Zuk5bBdR2_1),.din(w_dff_A_XmdMQl875_1),.clk(gclk));
	jdff dff_A_fTGx2qLi0_1(.dout(w_dff_A_XmdMQl875_1),.din(w_dff_A_fTGx2qLi0_1),.clk(gclk));
	jdff dff_A_utYalneR2_1(.dout(w_dff_A_fTGx2qLi0_1),.din(w_dff_A_utYalneR2_1),.clk(gclk));
	jdff dff_A_O3Ww4BRY8_1(.dout(w_dff_A_utYalneR2_1),.din(w_dff_A_O3Ww4BRY8_1),.clk(gclk));
	jdff dff_A_mKvn4gex2_1(.dout(w_dff_A_O3Ww4BRY8_1),.din(w_dff_A_mKvn4gex2_1),.clk(gclk));
	jdff dff_A_dLNERbTQ0_1(.dout(w_dff_A_mKvn4gex2_1),.din(w_dff_A_dLNERbTQ0_1),.clk(gclk));
	jdff dff_A_f6YOuO1D5_1(.dout(w_dff_A_dLNERbTQ0_1),.din(w_dff_A_f6YOuO1D5_1),.clk(gclk));
	jdff dff_A_egaLtwEk4_1(.dout(w_dff_A_f6YOuO1D5_1),.din(w_dff_A_egaLtwEk4_1),.clk(gclk));
	jdff dff_A_LUEqeTel1_1(.dout(w_dff_A_egaLtwEk4_1),.din(w_dff_A_LUEqeTel1_1),.clk(gclk));
	jdff dff_A_EijMotbY9_1(.dout(w_dff_A_LUEqeTel1_1),.din(w_dff_A_EijMotbY9_1),.clk(gclk));
	jdff dff_B_JZFTKxDn2_1(.din(n1790),.dout(w_dff_B_JZFTKxDn2_1),.clk(gclk));
	jdff dff_B_Q0BzWonC9_1(.din(w_dff_B_JZFTKxDn2_1),.dout(w_dff_B_Q0BzWonC9_1),.clk(gclk));
	jdff dff_B_pUELCfFY0_1(.din(w_dff_B_Q0BzWonC9_1),.dout(w_dff_B_pUELCfFY0_1),.clk(gclk));
	jdff dff_B_qPzFQeqf9_1(.din(w_dff_B_pUELCfFY0_1),.dout(w_dff_B_qPzFQeqf9_1),.clk(gclk));
	jdff dff_B_i7PfZVBg9_1(.din(w_dff_B_qPzFQeqf9_1),.dout(w_dff_B_i7PfZVBg9_1),.clk(gclk));
	jdff dff_B_OIjBg37i3_1(.din(w_dff_B_i7PfZVBg9_1),.dout(w_dff_B_OIjBg37i3_1),.clk(gclk));
	jdff dff_B_qPt7sSKQ0_1(.din(w_dff_B_OIjBg37i3_1),.dout(w_dff_B_qPt7sSKQ0_1),.clk(gclk));
	jdff dff_B_7t4VlZ8f3_1(.din(w_dff_B_qPt7sSKQ0_1),.dout(w_dff_B_7t4VlZ8f3_1),.clk(gclk));
	jdff dff_B_5hOmHfHY5_1(.din(w_dff_B_7t4VlZ8f3_1),.dout(w_dff_B_5hOmHfHY5_1),.clk(gclk));
	jdff dff_B_UzRMDacO5_1(.din(w_dff_B_5hOmHfHY5_1),.dout(w_dff_B_UzRMDacO5_1),.clk(gclk));
	jdff dff_B_1h0hJmOv9_1(.din(w_dff_B_UzRMDacO5_1),.dout(w_dff_B_1h0hJmOv9_1),.clk(gclk));
	jdff dff_B_40IKokeU0_1(.din(w_dff_B_1h0hJmOv9_1),.dout(w_dff_B_40IKokeU0_1),.clk(gclk));
	jdff dff_B_IpFzrpKs7_1(.din(w_dff_B_40IKokeU0_1),.dout(w_dff_B_IpFzrpKs7_1),.clk(gclk));
	jdff dff_B_IRhPFDK15_0(.din(n1791),.dout(w_dff_B_IRhPFDK15_0),.clk(gclk));
	jdff dff_B_DZZ7xxOB1_0(.din(w_dff_B_IRhPFDK15_0),.dout(w_dff_B_DZZ7xxOB1_0),.clk(gclk));
	jdff dff_B_Ms9m2RZg5_0(.din(w_dff_B_DZZ7xxOB1_0),.dout(w_dff_B_Ms9m2RZg5_0),.clk(gclk));
	jdff dff_B_Tf8hITD79_0(.din(w_dff_B_Ms9m2RZg5_0),.dout(w_dff_B_Tf8hITD79_0),.clk(gclk));
	jdff dff_B_VBqWJIOP3_0(.din(w_dff_B_Tf8hITD79_0),.dout(w_dff_B_VBqWJIOP3_0),.clk(gclk));
	jdff dff_B_Q9Ep1u1e0_0(.din(w_dff_B_VBqWJIOP3_0),.dout(w_dff_B_Q9Ep1u1e0_0),.clk(gclk));
	jdff dff_B_RdanKSAU4_0(.din(w_dff_B_Q9Ep1u1e0_0),.dout(w_dff_B_RdanKSAU4_0),.clk(gclk));
	jdff dff_B_zRxMcXDf4_0(.din(w_dff_B_RdanKSAU4_0),.dout(w_dff_B_zRxMcXDf4_0),.clk(gclk));
	jdff dff_B_DZvr5bWe2_0(.din(w_dff_B_zRxMcXDf4_0),.dout(w_dff_B_DZvr5bWe2_0),.clk(gclk));
	jdff dff_B_8UlkmnOB0_0(.din(w_dff_B_DZvr5bWe2_0),.dout(w_dff_B_8UlkmnOB0_0),.clk(gclk));
	jdff dff_B_QyIv5YhC3_0(.din(w_dff_B_8UlkmnOB0_0),.dout(w_dff_B_QyIv5YhC3_0),.clk(gclk));
	jdff dff_B_Eax2j83u3_0(.din(w_dff_B_QyIv5YhC3_0),.dout(w_dff_B_Eax2j83u3_0),.clk(gclk));
	jdff dff_A_T9KFEdex7_1(.dout(w_n1786_0[1]),.din(w_dff_A_T9KFEdex7_1),.clk(gclk));
	jdff dff_A_thZzegve2_1(.dout(w_dff_A_T9KFEdex7_1),.din(w_dff_A_thZzegve2_1),.clk(gclk));
	jdff dff_A_NmoBlnr84_1(.dout(w_dff_A_thZzegve2_1),.din(w_dff_A_NmoBlnr84_1),.clk(gclk));
	jdff dff_A_YyDrITFP6_1(.dout(w_dff_A_NmoBlnr84_1),.din(w_dff_A_YyDrITFP6_1),.clk(gclk));
	jdff dff_A_u4u4lKZC1_1(.dout(w_dff_A_YyDrITFP6_1),.din(w_dff_A_u4u4lKZC1_1),.clk(gclk));
	jdff dff_A_1khubOvS9_1(.dout(w_dff_A_u4u4lKZC1_1),.din(w_dff_A_1khubOvS9_1),.clk(gclk));
	jdff dff_A_cntyXHu83_1(.dout(w_dff_A_1khubOvS9_1),.din(w_dff_A_cntyXHu83_1),.clk(gclk));
	jdff dff_A_9fO0aOLe4_1(.dout(w_dff_A_cntyXHu83_1),.din(w_dff_A_9fO0aOLe4_1),.clk(gclk));
	jdff dff_A_00BVOmPM9_1(.dout(w_dff_A_9fO0aOLe4_1),.din(w_dff_A_00BVOmPM9_1),.clk(gclk));
	jdff dff_A_PwVDHGN71_1(.dout(w_dff_A_00BVOmPM9_1),.din(w_dff_A_PwVDHGN71_1),.clk(gclk));
	jdff dff_A_Fge183R41_1(.dout(w_dff_A_PwVDHGN71_1),.din(w_dff_A_Fge183R41_1),.clk(gclk));
	jdff dff_A_KFt5GgIB4_1(.dout(w_dff_A_Fge183R41_1),.din(w_dff_A_KFt5GgIB4_1),.clk(gclk));
	jdff dff_A_4KVlAlWx1_1(.dout(w_dff_A_KFt5GgIB4_1),.din(w_dff_A_4KVlAlWx1_1),.clk(gclk));
	jdff dff_B_7cx5V5OS2_1(.din(n1764),.dout(w_dff_B_7cx5V5OS2_1),.clk(gclk));
	jdff dff_B_ReRrmSwX3_1(.din(w_dff_B_7cx5V5OS2_1),.dout(w_dff_B_ReRrmSwX3_1),.clk(gclk));
	jdff dff_B_NfX4C5BL4_1(.din(w_dff_B_ReRrmSwX3_1),.dout(w_dff_B_NfX4C5BL4_1),.clk(gclk));
	jdff dff_B_5r5z626r1_1(.din(w_dff_B_NfX4C5BL4_1),.dout(w_dff_B_5r5z626r1_1),.clk(gclk));
	jdff dff_B_COetow5J0_1(.din(w_dff_B_5r5z626r1_1),.dout(w_dff_B_COetow5J0_1),.clk(gclk));
	jdff dff_B_pFK8Rx8K0_1(.din(w_dff_B_COetow5J0_1),.dout(w_dff_B_pFK8Rx8K0_1),.clk(gclk));
	jdff dff_B_8rAwLMxX9_1(.din(w_dff_B_pFK8Rx8K0_1),.dout(w_dff_B_8rAwLMxX9_1),.clk(gclk));
	jdff dff_B_PrtGY1vA8_1(.din(w_dff_B_8rAwLMxX9_1),.dout(w_dff_B_PrtGY1vA8_1),.clk(gclk));
	jdff dff_B_l4sWRafE4_1(.din(w_dff_B_PrtGY1vA8_1),.dout(w_dff_B_l4sWRafE4_1),.clk(gclk));
	jdff dff_B_W4LavJEj3_1(.din(w_dff_B_l4sWRafE4_1),.dout(w_dff_B_W4LavJEj3_1),.clk(gclk));
	jdff dff_B_nQ5eUGWD8_1(.din(w_dff_B_W4LavJEj3_1),.dout(w_dff_B_nQ5eUGWD8_1),.clk(gclk));
	jdff dff_B_Kp36zHGa5_1(.din(w_dff_B_nQ5eUGWD8_1),.dout(w_dff_B_Kp36zHGa5_1),.clk(gclk));
	jdff dff_B_vZrwHUxD9_1(.din(w_dff_B_Kp36zHGa5_1),.dout(w_dff_B_vZrwHUxD9_1),.clk(gclk));
	jdff dff_B_jzMeZDf95_0(.din(n1765),.dout(w_dff_B_jzMeZDf95_0),.clk(gclk));
	jdff dff_B_5DhVa4wc8_0(.din(w_dff_B_jzMeZDf95_0),.dout(w_dff_B_5DhVa4wc8_0),.clk(gclk));
	jdff dff_B_fVEdAqmM8_0(.din(w_dff_B_5DhVa4wc8_0),.dout(w_dff_B_fVEdAqmM8_0),.clk(gclk));
	jdff dff_B_5T5gmPkk3_0(.din(w_dff_B_fVEdAqmM8_0),.dout(w_dff_B_5T5gmPkk3_0),.clk(gclk));
	jdff dff_B_PZ3rIPaP9_0(.din(w_dff_B_5T5gmPkk3_0),.dout(w_dff_B_PZ3rIPaP9_0),.clk(gclk));
	jdff dff_B_w6hWCenc1_0(.din(w_dff_B_PZ3rIPaP9_0),.dout(w_dff_B_w6hWCenc1_0),.clk(gclk));
	jdff dff_B_7Mf5edzX4_0(.din(w_dff_B_w6hWCenc1_0),.dout(w_dff_B_7Mf5edzX4_0),.clk(gclk));
	jdff dff_B_RZvoK1t43_0(.din(w_dff_B_7Mf5edzX4_0),.dout(w_dff_B_RZvoK1t43_0),.clk(gclk));
	jdff dff_B_b303HJ6h9_0(.din(w_dff_B_RZvoK1t43_0),.dout(w_dff_B_b303HJ6h9_0),.clk(gclk));
	jdff dff_B_G5rdZPoX8_0(.din(w_dff_B_b303HJ6h9_0),.dout(w_dff_B_G5rdZPoX8_0),.clk(gclk));
	jdff dff_B_s6zas3fz4_0(.din(w_dff_B_G5rdZPoX8_0),.dout(w_dff_B_s6zas3fz4_0),.clk(gclk));
	jdff dff_B_S9IxMMvX1_0(.din(w_dff_B_s6zas3fz4_0),.dout(w_dff_B_S9IxMMvX1_0),.clk(gclk));
	jdff dff_A_Ug5KqzIZ5_1(.dout(w_n1760_0[1]),.din(w_dff_A_Ug5KqzIZ5_1),.clk(gclk));
	jdff dff_A_qO2T8b5F1_1(.dout(w_dff_A_Ug5KqzIZ5_1),.din(w_dff_A_qO2T8b5F1_1),.clk(gclk));
	jdff dff_A_TXgtV5ST9_1(.dout(w_dff_A_qO2T8b5F1_1),.din(w_dff_A_TXgtV5ST9_1),.clk(gclk));
	jdff dff_A_uKmyPLmp7_1(.dout(w_dff_A_TXgtV5ST9_1),.din(w_dff_A_uKmyPLmp7_1),.clk(gclk));
	jdff dff_A_KeylDWXq9_1(.dout(w_dff_A_uKmyPLmp7_1),.din(w_dff_A_KeylDWXq9_1),.clk(gclk));
	jdff dff_A_KG7eG7Oz2_1(.dout(w_dff_A_KeylDWXq9_1),.din(w_dff_A_KG7eG7Oz2_1),.clk(gclk));
	jdff dff_A_U5LspV7W1_1(.dout(w_dff_A_KG7eG7Oz2_1),.din(w_dff_A_U5LspV7W1_1),.clk(gclk));
	jdff dff_A_kd3jYeLR4_1(.dout(w_dff_A_U5LspV7W1_1),.din(w_dff_A_kd3jYeLR4_1),.clk(gclk));
	jdff dff_A_SwWRfXa71_1(.dout(w_dff_A_kd3jYeLR4_1),.din(w_dff_A_SwWRfXa71_1),.clk(gclk));
	jdff dff_A_W4ClE6JB0_1(.dout(w_dff_A_SwWRfXa71_1),.din(w_dff_A_W4ClE6JB0_1),.clk(gclk));
	jdff dff_A_qcyHLUih9_1(.dout(w_dff_A_W4ClE6JB0_1),.din(w_dff_A_qcyHLUih9_1),.clk(gclk));
	jdff dff_A_W973r2Lm0_1(.dout(w_dff_A_qcyHLUih9_1),.din(w_dff_A_W973r2Lm0_1),.clk(gclk));
	jdff dff_A_2vTb8S2q8_1(.dout(w_dff_A_W973r2Lm0_1),.din(w_dff_A_2vTb8S2q8_1),.clk(gclk));
	jdff dff_B_SLTue1W65_1(.din(n1731),.dout(w_dff_B_SLTue1W65_1),.clk(gclk));
	jdff dff_B_wG7sHNVc7_1(.din(w_dff_B_SLTue1W65_1),.dout(w_dff_B_wG7sHNVc7_1),.clk(gclk));
	jdff dff_B_ba6ckuz21_1(.din(w_dff_B_wG7sHNVc7_1),.dout(w_dff_B_ba6ckuz21_1),.clk(gclk));
	jdff dff_B_erD4iTHp1_1(.din(w_dff_B_ba6ckuz21_1),.dout(w_dff_B_erD4iTHp1_1),.clk(gclk));
	jdff dff_B_FvnSXbol5_1(.din(w_dff_B_erD4iTHp1_1),.dout(w_dff_B_FvnSXbol5_1),.clk(gclk));
	jdff dff_B_2IHLg49y6_1(.din(w_dff_B_FvnSXbol5_1),.dout(w_dff_B_2IHLg49y6_1),.clk(gclk));
	jdff dff_B_uyEcYBeg8_1(.din(w_dff_B_2IHLg49y6_1),.dout(w_dff_B_uyEcYBeg8_1),.clk(gclk));
	jdff dff_B_rNQUTJS04_1(.din(w_dff_B_uyEcYBeg8_1),.dout(w_dff_B_rNQUTJS04_1),.clk(gclk));
	jdff dff_B_1QXjkdFr7_1(.din(w_dff_B_rNQUTJS04_1),.dout(w_dff_B_1QXjkdFr7_1),.clk(gclk));
	jdff dff_B_rQLgk7kU5_1(.din(w_dff_B_1QXjkdFr7_1),.dout(w_dff_B_rQLgk7kU5_1),.clk(gclk));
	jdff dff_B_PqH95pFh5_1(.din(w_dff_B_rQLgk7kU5_1),.dout(w_dff_B_PqH95pFh5_1),.clk(gclk));
	jdff dff_B_QA0up3dU1_1(.din(w_dff_B_PqH95pFh5_1),.dout(w_dff_B_QA0up3dU1_1),.clk(gclk));
	jdff dff_B_GZ6FuMXH6_1(.din(w_dff_B_QA0up3dU1_1),.dout(w_dff_B_GZ6FuMXH6_1),.clk(gclk));
	jdff dff_B_Cb6IpgKB9_0(.din(n1732),.dout(w_dff_B_Cb6IpgKB9_0),.clk(gclk));
	jdff dff_B_ZdELOMLu5_0(.din(w_dff_B_Cb6IpgKB9_0),.dout(w_dff_B_ZdELOMLu5_0),.clk(gclk));
	jdff dff_B_PF9u3AFH8_0(.din(w_dff_B_ZdELOMLu5_0),.dout(w_dff_B_PF9u3AFH8_0),.clk(gclk));
	jdff dff_B_S76kN2ap0_0(.din(w_dff_B_PF9u3AFH8_0),.dout(w_dff_B_S76kN2ap0_0),.clk(gclk));
	jdff dff_B_ruAuqKJX9_0(.din(w_dff_B_S76kN2ap0_0),.dout(w_dff_B_ruAuqKJX9_0),.clk(gclk));
	jdff dff_B_BLKp01f08_0(.din(w_dff_B_ruAuqKJX9_0),.dout(w_dff_B_BLKp01f08_0),.clk(gclk));
	jdff dff_B_PMavN43V1_0(.din(w_dff_B_BLKp01f08_0),.dout(w_dff_B_PMavN43V1_0),.clk(gclk));
	jdff dff_B_s64Hssp82_0(.din(w_dff_B_PMavN43V1_0),.dout(w_dff_B_s64Hssp82_0),.clk(gclk));
	jdff dff_B_pnyncAxt8_0(.din(w_dff_B_s64Hssp82_0),.dout(w_dff_B_pnyncAxt8_0),.clk(gclk));
	jdff dff_B_zTtpbYN36_0(.din(w_dff_B_pnyncAxt8_0),.dout(w_dff_B_zTtpbYN36_0),.clk(gclk));
	jdff dff_B_XRCDyfgr8_0(.din(w_dff_B_zTtpbYN36_0),.dout(w_dff_B_XRCDyfgr8_0),.clk(gclk));
	jdff dff_B_OqdGXR4B1_0(.din(w_dff_B_XRCDyfgr8_0),.dout(w_dff_B_OqdGXR4B1_0),.clk(gclk));
	jdff dff_A_JCm8jvZF4_1(.dout(w_n1727_0[1]),.din(w_dff_A_JCm8jvZF4_1),.clk(gclk));
	jdff dff_A_AhLKwjoj4_1(.dout(w_dff_A_JCm8jvZF4_1),.din(w_dff_A_AhLKwjoj4_1),.clk(gclk));
	jdff dff_A_lJae0g2f1_1(.dout(w_dff_A_AhLKwjoj4_1),.din(w_dff_A_lJae0g2f1_1),.clk(gclk));
	jdff dff_A_vNbAUVf23_1(.dout(w_dff_A_lJae0g2f1_1),.din(w_dff_A_vNbAUVf23_1),.clk(gclk));
	jdff dff_A_yWsghXlF1_1(.dout(w_dff_A_vNbAUVf23_1),.din(w_dff_A_yWsghXlF1_1),.clk(gclk));
	jdff dff_A_hKMZwiL11_1(.dout(w_dff_A_yWsghXlF1_1),.din(w_dff_A_hKMZwiL11_1),.clk(gclk));
	jdff dff_A_DNxx7Crx3_1(.dout(w_dff_A_hKMZwiL11_1),.din(w_dff_A_DNxx7Crx3_1),.clk(gclk));
	jdff dff_A_7lesqXUP2_1(.dout(w_dff_A_DNxx7Crx3_1),.din(w_dff_A_7lesqXUP2_1),.clk(gclk));
	jdff dff_A_oWZPXYVD3_1(.dout(w_dff_A_7lesqXUP2_1),.din(w_dff_A_oWZPXYVD3_1),.clk(gclk));
	jdff dff_A_pykIj7No3_1(.dout(w_dff_A_oWZPXYVD3_1),.din(w_dff_A_pykIj7No3_1),.clk(gclk));
	jdff dff_A_SeyeNzVn7_1(.dout(w_dff_A_pykIj7No3_1),.din(w_dff_A_SeyeNzVn7_1),.clk(gclk));
	jdff dff_A_xwhHnZWD3_1(.dout(w_dff_A_SeyeNzVn7_1),.din(w_dff_A_xwhHnZWD3_1),.clk(gclk));
	jdff dff_A_itjcwYbR2_1(.dout(w_dff_A_xwhHnZWD3_1),.din(w_dff_A_itjcwYbR2_1),.clk(gclk));
	jdff dff_B_98i5q6i27_1(.din(n1691),.dout(w_dff_B_98i5q6i27_1),.clk(gclk));
	jdff dff_B_Fh22ZAkX4_1(.din(w_dff_B_98i5q6i27_1),.dout(w_dff_B_Fh22ZAkX4_1),.clk(gclk));
	jdff dff_B_FeHEPAxG1_1(.din(w_dff_B_Fh22ZAkX4_1),.dout(w_dff_B_FeHEPAxG1_1),.clk(gclk));
	jdff dff_B_VdMhXcsq0_1(.din(w_dff_B_FeHEPAxG1_1),.dout(w_dff_B_VdMhXcsq0_1),.clk(gclk));
	jdff dff_B_O3wFpCtC9_1(.din(w_dff_B_VdMhXcsq0_1),.dout(w_dff_B_O3wFpCtC9_1),.clk(gclk));
	jdff dff_B_XAIlAHcE4_1(.din(w_dff_B_O3wFpCtC9_1),.dout(w_dff_B_XAIlAHcE4_1),.clk(gclk));
	jdff dff_B_Q9VHc7v35_1(.din(w_dff_B_XAIlAHcE4_1),.dout(w_dff_B_Q9VHc7v35_1),.clk(gclk));
	jdff dff_B_HXF8qjwB7_1(.din(w_dff_B_Q9VHc7v35_1),.dout(w_dff_B_HXF8qjwB7_1),.clk(gclk));
	jdff dff_B_Pqnhn7Bk7_1(.din(w_dff_B_HXF8qjwB7_1),.dout(w_dff_B_Pqnhn7Bk7_1),.clk(gclk));
	jdff dff_B_ITdeaySm6_1(.din(w_dff_B_Pqnhn7Bk7_1),.dout(w_dff_B_ITdeaySm6_1),.clk(gclk));
	jdff dff_B_wSBEcLQg8_1(.din(w_dff_B_ITdeaySm6_1),.dout(w_dff_B_wSBEcLQg8_1),.clk(gclk));
	jdff dff_B_KKewNWnA2_1(.din(w_dff_B_wSBEcLQg8_1),.dout(w_dff_B_KKewNWnA2_1),.clk(gclk));
	jdff dff_B_uLOxlXOx2_1(.din(w_dff_B_KKewNWnA2_1),.dout(w_dff_B_uLOxlXOx2_1),.clk(gclk));
	jdff dff_B_Wi4txK3w5_0(.din(n1692),.dout(w_dff_B_Wi4txK3w5_0),.clk(gclk));
	jdff dff_B_CjUudyhj4_0(.din(w_dff_B_Wi4txK3w5_0),.dout(w_dff_B_CjUudyhj4_0),.clk(gclk));
	jdff dff_B_GVUNx34g6_0(.din(w_dff_B_CjUudyhj4_0),.dout(w_dff_B_GVUNx34g6_0),.clk(gclk));
	jdff dff_B_Ld7x9OEn2_0(.din(w_dff_B_GVUNx34g6_0),.dout(w_dff_B_Ld7x9OEn2_0),.clk(gclk));
	jdff dff_B_qM2GOlFb8_0(.din(w_dff_B_Ld7x9OEn2_0),.dout(w_dff_B_qM2GOlFb8_0),.clk(gclk));
	jdff dff_B_dVl6r7ub5_0(.din(w_dff_B_qM2GOlFb8_0),.dout(w_dff_B_dVl6r7ub5_0),.clk(gclk));
	jdff dff_B_WkKibG8O6_0(.din(w_dff_B_dVl6r7ub5_0),.dout(w_dff_B_WkKibG8O6_0),.clk(gclk));
	jdff dff_B_LXJBMZb92_0(.din(w_dff_B_WkKibG8O6_0),.dout(w_dff_B_LXJBMZb92_0),.clk(gclk));
	jdff dff_B_b1Uc1eAx7_0(.din(w_dff_B_LXJBMZb92_0),.dout(w_dff_B_b1Uc1eAx7_0),.clk(gclk));
	jdff dff_B_9ji28POX1_0(.din(w_dff_B_b1Uc1eAx7_0),.dout(w_dff_B_9ji28POX1_0),.clk(gclk));
	jdff dff_B_XuXI86Ur9_0(.din(w_dff_B_9ji28POX1_0),.dout(w_dff_B_XuXI86Ur9_0),.clk(gclk));
	jdff dff_A_gKVDurJ62_1(.dout(w_n1689_0[1]),.din(w_dff_A_gKVDurJ62_1),.clk(gclk));
	jdff dff_A_1sc3yxxC3_1(.dout(w_dff_A_gKVDurJ62_1),.din(w_dff_A_1sc3yxxC3_1),.clk(gclk));
	jdff dff_A_cu9ioHt23_1(.dout(w_dff_A_1sc3yxxC3_1),.din(w_dff_A_cu9ioHt23_1),.clk(gclk));
	jdff dff_A_0mqTJW9U4_1(.dout(w_dff_A_cu9ioHt23_1),.din(w_dff_A_0mqTJW9U4_1),.clk(gclk));
	jdff dff_A_EIqOoX1y5_1(.dout(w_dff_A_0mqTJW9U4_1),.din(w_dff_A_EIqOoX1y5_1),.clk(gclk));
	jdff dff_A_gRxDMbuh5_1(.dout(w_dff_A_EIqOoX1y5_1),.din(w_dff_A_gRxDMbuh5_1),.clk(gclk));
	jdff dff_A_dO0tdUbf9_1(.dout(w_dff_A_gRxDMbuh5_1),.din(w_dff_A_dO0tdUbf9_1),.clk(gclk));
	jdff dff_A_wO1vKqH19_1(.dout(w_dff_A_dO0tdUbf9_1),.din(w_dff_A_wO1vKqH19_1),.clk(gclk));
	jdff dff_A_AlW3KyGb2_1(.dout(w_dff_A_wO1vKqH19_1),.din(w_dff_A_AlW3KyGb2_1),.clk(gclk));
	jdff dff_A_cHmjjC4Q0_1(.dout(w_dff_A_AlW3KyGb2_1),.din(w_dff_A_cHmjjC4Q0_1),.clk(gclk));
	jdff dff_A_ayZfOxte6_1(.dout(w_dff_A_cHmjjC4Q0_1),.din(w_dff_A_ayZfOxte6_1),.clk(gclk));
	jdff dff_A_hBr7Bvkn6_1(.dout(w_dff_A_ayZfOxte6_1),.din(w_dff_A_hBr7Bvkn6_1),.clk(gclk));
	jdff dff_B_xRqPyWT30_1(.din(n1643),.dout(w_dff_B_xRqPyWT30_1),.clk(gclk));
	jdff dff_B_7xCgBDri0_1(.din(w_dff_B_xRqPyWT30_1),.dout(w_dff_B_7xCgBDri0_1),.clk(gclk));
	jdff dff_B_3zrg0aoQ8_1(.din(w_dff_B_7xCgBDri0_1),.dout(w_dff_B_3zrg0aoQ8_1),.clk(gclk));
	jdff dff_B_R4DVJwf72_1(.din(w_dff_B_3zrg0aoQ8_1),.dout(w_dff_B_R4DVJwf72_1),.clk(gclk));
	jdff dff_B_WGzgPYBE1_1(.din(w_dff_B_R4DVJwf72_1),.dout(w_dff_B_WGzgPYBE1_1),.clk(gclk));
	jdff dff_B_sf6Vy6wZ7_1(.din(w_dff_B_WGzgPYBE1_1),.dout(w_dff_B_sf6Vy6wZ7_1),.clk(gclk));
	jdff dff_B_mqIlxu2V0_1(.din(w_dff_B_sf6Vy6wZ7_1),.dout(w_dff_B_mqIlxu2V0_1),.clk(gclk));
	jdff dff_B_BeKu9XTA9_1(.din(w_dff_B_mqIlxu2V0_1),.dout(w_dff_B_BeKu9XTA9_1),.clk(gclk));
	jdff dff_B_J2xOxtYg1_1(.din(w_dff_B_BeKu9XTA9_1),.dout(w_dff_B_J2xOxtYg1_1),.clk(gclk));
	jdff dff_B_av4IUyOg2_1(.din(w_dff_B_J2xOxtYg1_1),.dout(w_dff_B_av4IUyOg2_1),.clk(gclk));
	jdff dff_B_8W0lI1PT1_1(.din(w_dff_B_av4IUyOg2_1),.dout(w_dff_B_8W0lI1PT1_1),.clk(gclk));
	jdff dff_B_UBMYoQfe2_1(.din(w_dff_B_8W0lI1PT1_1),.dout(w_dff_B_UBMYoQfe2_1),.clk(gclk));
	jdff dff_B_7QMxYCto9_0(.din(n1644),.dout(w_dff_B_7QMxYCto9_0),.clk(gclk));
	jdff dff_B_M5Yd0prC2_0(.din(w_dff_B_7QMxYCto9_0),.dout(w_dff_B_M5Yd0prC2_0),.clk(gclk));
	jdff dff_B_Vx59Mf9W3_0(.din(w_dff_B_M5Yd0prC2_0),.dout(w_dff_B_Vx59Mf9W3_0),.clk(gclk));
	jdff dff_B_iMYbj4g92_0(.din(w_dff_B_Vx59Mf9W3_0),.dout(w_dff_B_iMYbj4g92_0),.clk(gclk));
	jdff dff_B_DGejjhsJ7_0(.din(w_dff_B_iMYbj4g92_0),.dout(w_dff_B_DGejjhsJ7_0),.clk(gclk));
	jdff dff_B_CxLbiHdJ0_0(.din(w_dff_B_DGejjhsJ7_0),.dout(w_dff_B_CxLbiHdJ0_0),.clk(gclk));
	jdff dff_B_CoNQfLzc0_0(.din(w_dff_B_CxLbiHdJ0_0),.dout(w_dff_B_CoNQfLzc0_0),.clk(gclk));
	jdff dff_B_5Qs5fN2D5_0(.din(w_dff_B_CoNQfLzc0_0),.dout(w_dff_B_5Qs5fN2D5_0),.clk(gclk));
	jdff dff_B_lZtfl94T7_0(.din(w_dff_B_5Qs5fN2D5_0),.dout(w_dff_B_lZtfl94T7_0),.clk(gclk));
	jdff dff_B_AIWOmTrF2_0(.din(w_dff_B_lZtfl94T7_0),.dout(w_dff_B_AIWOmTrF2_0),.clk(gclk));
	jdff dff_A_79xTRdAA4_1(.dout(w_n1641_0[1]),.din(w_dff_A_79xTRdAA4_1),.clk(gclk));
	jdff dff_A_kH0vxITY7_1(.dout(w_dff_A_79xTRdAA4_1),.din(w_dff_A_kH0vxITY7_1),.clk(gclk));
	jdff dff_A_u570xPwX1_1(.dout(w_dff_A_kH0vxITY7_1),.din(w_dff_A_u570xPwX1_1),.clk(gclk));
	jdff dff_A_dcjzw2mt2_1(.dout(w_dff_A_u570xPwX1_1),.din(w_dff_A_dcjzw2mt2_1),.clk(gclk));
	jdff dff_A_5uLvVhj20_1(.dout(w_dff_A_dcjzw2mt2_1),.din(w_dff_A_5uLvVhj20_1),.clk(gclk));
	jdff dff_A_KvJKSr7d0_1(.dout(w_dff_A_5uLvVhj20_1),.din(w_dff_A_KvJKSr7d0_1),.clk(gclk));
	jdff dff_A_sb1lZJCh5_1(.dout(w_dff_A_KvJKSr7d0_1),.din(w_dff_A_sb1lZJCh5_1),.clk(gclk));
	jdff dff_A_t3zvyWfM6_1(.dout(w_dff_A_sb1lZJCh5_1),.din(w_dff_A_t3zvyWfM6_1),.clk(gclk));
	jdff dff_A_vjISJLyS1_1(.dout(w_dff_A_t3zvyWfM6_1),.din(w_dff_A_vjISJLyS1_1),.clk(gclk));
	jdff dff_A_rg0cV6kt8_1(.dout(w_dff_A_vjISJLyS1_1),.din(w_dff_A_rg0cV6kt8_1),.clk(gclk));
	jdff dff_A_KvEs2OMJ1_1(.dout(w_dff_A_rg0cV6kt8_1),.din(w_dff_A_KvEs2OMJ1_1),.clk(gclk));
	jdff dff_B_WWBzEK2t8_1(.din(n1588),.dout(w_dff_B_WWBzEK2t8_1),.clk(gclk));
	jdff dff_B_jz9KcFHN7_1(.din(w_dff_B_WWBzEK2t8_1),.dout(w_dff_B_jz9KcFHN7_1),.clk(gclk));
	jdff dff_B_QwGmC3jj4_1(.din(w_dff_B_jz9KcFHN7_1),.dout(w_dff_B_QwGmC3jj4_1),.clk(gclk));
	jdff dff_B_DNqCeEMs2_1(.din(w_dff_B_QwGmC3jj4_1),.dout(w_dff_B_DNqCeEMs2_1),.clk(gclk));
	jdff dff_B_GIAzMXZK9_1(.din(w_dff_B_DNqCeEMs2_1),.dout(w_dff_B_GIAzMXZK9_1),.clk(gclk));
	jdff dff_B_sTdSgllS3_1(.din(w_dff_B_GIAzMXZK9_1),.dout(w_dff_B_sTdSgllS3_1),.clk(gclk));
	jdff dff_B_bUz2w9d47_1(.din(w_dff_B_sTdSgllS3_1),.dout(w_dff_B_bUz2w9d47_1),.clk(gclk));
	jdff dff_B_g6IpYB3m0_1(.din(w_dff_B_bUz2w9d47_1),.dout(w_dff_B_g6IpYB3m0_1),.clk(gclk));
	jdff dff_B_zsifSQsn5_1(.din(w_dff_B_g6IpYB3m0_1),.dout(w_dff_B_zsifSQsn5_1),.clk(gclk));
	jdff dff_B_8ztmIV7a7_1(.din(w_dff_B_zsifSQsn5_1),.dout(w_dff_B_8ztmIV7a7_1),.clk(gclk));
	jdff dff_B_cv02aKdX6_0(.din(n1589),.dout(w_dff_B_cv02aKdX6_0),.clk(gclk));
	jdff dff_B_Cl3RWvNn9_0(.din(w_dff_B_cv02aKdX6_0),.dout(w_dff_B_Cl3RWvNn9_0),.clk(gclk));
	jdff dff_B_QvEk66Jp5_0(.din(w_dff_B_Cl3RWvNn9_0),.dout(w_dff_B_QvEk66Jp5_0),.clk(gclk));
	jdff dff_B_Dd3l0Fwh4_0(.din(w_dff_B_QvEk66Jp5_0),.dout(w_dff_B_Dd3l0Fwh4_0),.clk(gclk));
	jdff dff_B_HwVYhdoW9_0(.din(w_dff_B_Dd3l0Fwh4_0),.dout(w_dff_B_HwVYhdoW9_0),.clk(gclk));
	jdff dff_B_ywhYHoMz5_0(.din(w_dff_B_HwVYhdoW9_0),.dout(w_dff_B_ywhYHoMz5_0),.clk(gclk));
	jdff dff_B_3WLio9ZI0_0(.din(w_dff_B_ywhYHoMz5_0),.dout(w_dff_B_3WLio9ZI0_0),.clk(gclk));
	jdff dff_B_NWY9YSYe7_0(.din(w_dff_B_3WLio9ZI0_0),.dout(w_dff_B_NWY9YSYe7_0),.clk(gclk));
	jdff dff_A_Fk4Cu5155_1(.dout(w_n1586_0[1]),.din(w_dff_A_Fk4Cu5155_1),.clk(gclk));
	jdff dff_A_KZreOOdV9_1(.dout(w_dff_A_Fk4Cu5155_1),.din(w_dff_A_KZreOOdV9_1),.clk(gclk));
	jdff dff_A_WGY0EMid1_1(.dout(w_dff_A_KZreOOdV9_1),.din(w_dff_A_WGY0EMid1_1),.clk(gclk));
	jdff dff_A_KFmSYE1H1_1(.dout(w_dff_A_WGY0EMid1_1),.din(w_dff_A_KFmSYE1H1_1),.clk(gclk));
	jdff dff_A_uJ5HZv8s5_1(.dout(w_dff_A_KFmSYE1H1_1),.din(w_dff_A_uJ5HZv8s5_1),.clk(gclk));
	jdff dff_A_1EExzx8z2_1(.dout(w_dff_A_uJ5HZv8s5_1),.din(w_dff_A_1EExzx8z2_1),.clk(gclk));
	jdff dff_A_do84FDrb8_1(.dout(w_dff_A_1EExzx8z2_1),.din(w_dff_A_do84FDrb8_1),.clk(gclk));
	jdff dff_A_c7TN3Ezh7_1(.dout(w_dff_A_do84FDrb8_1),.din(w_dff_A_c7TN3Ezh7_1),.clk(gclk));
	jdff dff_A_G80OTdUX1_1(.dout(w_dff_A_c7TN3Ezh7_1),.din(w_dff_A_G80OTdUX1_1),.clk(gclk));
	jdff dff_B_AA6gCB0m2_1(.din(n1526),.dout(w_dff_B_AA6gCB0m2_1),.clk(gclk));
	jdff dff_B_UpwJJE7z9_1(.din(w_dff_B_AA6gCB0m2_1),.dout(w_dff_B_UpwJJE7z9_1),.clk(gclk));
	jdff dff_B_pUJ00lGB5_1(.din(w_dff_B_UpwJJE7z9_1),.dout(w_dff_B_pUJ00lGB5_1),.clk(gclk));
	jdff dff_B_rwfAv5aH8_1(.din(w_dff_B_pUJ00lGB5_1),.dout(w_dff_B_rwfAv5aH8_1),.clk(gclk));
	jdff dff_B_UuU8hRCC1_1(.din(w_dff_B_rwfAv5aH8_1),.dout(w_dff_B_UuU8hRCC1_1),.clk(gclk));
	jdff dff_B_HEkJ4m610_1(.din(w_dff_B_UuU8hRCC1_1),.dout(w_dff_B_HEkJ4m610_1),.clk(gclk));
	jdff dff_B_pd6g6nrz3_1(.din(w_dff_B_HEkJ4m610_1),.dout(w_dff_B_pd6g6nrz3_1),.clk(gclk));
	jdff dff_B_D3AzhsqY2_1(.din(w_dff_B_pd6g6nrz3_1),.dout(w_dff_B_D3AzhsqY2_1),.clk(gclk));
	jdff dff_B_611Z2rBw0_0(.din(n1527),.dout(w_dff_B_611Z2rBw0_0),.clk(gclk));
	jdff dff_B_F8XMhViI5_0(.din(w_dff_B_611Z2rBw0_0),.dout(w_dff_B_F8XMhViI5_0),.clk(gclk));
	jdff dff_B_mm7wYaZM8_0(.din(w_dff_B_F8XMhViI5_0),.dout(w_dff_B_mm7wYaZM8_0),.clk(gclk));
	jdff dff_B_rNhRn8C72_0(.din(w_dff_B_mm7wYaZM8_0),.dout(w_dff_B_rNhRn8C72_0),.clk(gclk));
	jdff dff_B_6qUBbKno5_0(.din(w_dff_B_rNhRn8C72_0),.dout(w_dff_B_6qUBbKno5_0),.clk(gclk));
	jdff dff_B_J0oQAQk06_0(.din(w_dff_B_6qUBbKno5_0),.dout(w_dff_B_J0oQAQk06_0),.clk(gclk));
	jdff dff_A_KrEMh2ET3_1(.dout(w_n1524_0[1]),.din(w_dff_A_KrEMh2ET3_1),.clk(gclk));
	jdff dff_A_qs22pyxv8_1(.dout(w_dff_A_KrEMh2ET3_1),.din(w_dff_A_qs22pyxv8_1),.clk(gclk));
	jdff dff_A_yOIXtJdL9_1(.dout(w_dff_A_qs22pyxv8_1),.din(w_dff_A_yOIXtJdL9_1),.clk(gclk));
	jdff dff_A_tRTdw8lN6_1(.dout(w_dff_A_yOIXtJdL9_1),.din(w_dff_A_tRTdw8lN6_1),.clk(gclk));
	jdff dff_A_pniuvVG98_1(.dout(w_dff_A_tRTdw8lN6_1),.din(w_dff_A_pniuvVG98_1),.clk(gclk));
	jdff dff_A_GVrYQgqz7_1(.dout(w_dff_A_pniuvVG98_1),.din(w_dff_A_GVrYQgqz7_1),.clk(gclk));
	jdff dff_A_FdAfEhwx6_1(.dout(w_dff_A_GVrYQgqz7_1),.din(w_dff_A_FdAfEhwx6_1),.clk(gclk));
	jdff dff_B_s5VMcwp71_1(.din(n1457),.dout(w_dff_B_s5VMcwp71_1),.clk(gclk));
	jdff dff_B_7181w4Jd4_1(.din(w_dff_B_s5VMcwp71_1),.dout(w_dff_B_7181w4Jd4_1),.clk(gclk));
	jdff dff_B_XLyrQERS0_1(.din(w_dff_B_7181w4Jd4_1),.dout(w_dff_B_XLyrQERS0_1),.clk(gclk));
	jdff dff_B_jQnhG3HK0_1(.din(w_dff_B_XLyrQERS0_1),.dout(w_dff_B_jQnhG3HK0_1),.clk(gclk));
	jdff dff_B_q7HmttER1_1(.din(w_dff_B_jQnhG3HK0_1),.dout(w_dff_B_q7HmttER1_1),.clk(gclk));
	jdff dff_B_QfljtKyF7_1(.din(w_dff_B_q7HmttER1_1),.dout(w_dff_B_QfljtKyF7_1),.clk(gclk));
	jdff dff_B_ubHAw9xw6_1(.din(w_dff_B_QfljtKyF7_1),.dout(w_dff_B_ubHAw9xw6_1),.clk(gclk));
	jdff dff_B_A09hQSLQ0_0(.din(n1458),.dout(w_dff_B_A09hQSLQ0_0),.clk(gclk));
	jdff dff_B_YJMp2cQO5_0(.din(w_dff_B_A09hQSLQ0_0),.dout(w_dff_B_YJMp2cQO5_0),.clk(gclk));
	jdff dff_B_D1ub6vNA8_0(.din(w_dff_B_YJMp2cQO5_0),.dout(w_dff_B_D1ub6vNA8_0),.clk(gclk));
	jdff dff_B_KZXJQL4Y4_0(.din(w_dff_B_D1ub6vNA8_0),.dout(w_dff_B_KZXJQL4Y4_0),.clk(gclk));
	jdff dff_B_KxTD4Scz6_0(.din(w_dff_B_KZXJQL4Y4_0),.dout(w_dff_B_KxTD4Scz6_0),.clk(gclk));
	jdff dff_A_cvJhLKV41_1(.dout(w_n1455_0[1]),.din(w_dff_A_cvJhLKV41_1),.clk(gclk));
	jdff dff_A_9T6Ai5Ii2_1(.dout(w_dff_A_cvJhLKV41_1),.din(w_dff_A_9T6Ai5Ii2_1),.clk(gclk));
	jdff dff_A_NmxiMzk67_1(.dout(w_dff_A_9T6Ai5Ii2_1),.din(w_dff_A_NmxiMzk67_1),.clk(gclk));
	jdff dff_A_h258285L2_1(.dout(w_dff_A_NmxiMzk67_1),.din(w_dff_A_h258285L2_1),.clk(gclk));
	jdff dff_A_peibwPQ52_1(.dout(w_dff_A_h258285L2_1),.din(w_dff_A_peibwPQ52_1),.clk(gclk));
	jdff dff_A_q7PYhXqR0_1(.dout(w_dff_A_peibwPQ52_1),.din(w_dff_A_q7PYhXqR0_1),.clk(gclk));
	jdff dff_B_SFLsw30A8_1(.din(n1381),.dout(w_dff_B_SFLsw30A8_1),.clk(gclk));
	jdff dff_B_CbvifFGY4_1(.din(w_dff_B_SFLsw30A8_1),.dout(w_dff_B_CbvifFGY4_1),.clk(gclk));
	jdff dff_B_HGeey1hP9_1(.din(w_dff_B_CbvifFGY4_1),.dout(w_dff_B_HGeey1hP9_1),.clk(gclk));
	jdff dff_B_mSLgcSV87_1(.din(w_dff_B_HGeey1hP9_1),.dout(w_dff_B_mSLgcSV87_1),.clk(gclk));
	jdff dff_B_NnlQCR6R8_1(.din(w_dff_B_mSLgcSV87_1),.dout(w_dff_B_NnlQCR6R8_1),.clk(gclk));
	jdff dff_B_tmWz7Xxw0_1(.din(w_dff_B_NnlQCR6R8_1),.dout(w_dff_B_tmWz7Xxw0_1),.clk(gclk));
	jdff dff_B_fKEZf45O2_0(.din(n1382),.dout(w_dff_B_fKEZf45O2_0),.clk(gclk));
	jdff dff_B_TW7vS4AY7_0(.din(w_dff_B_fKEZf45O2_0),.dout(w_dff_B_TW7vS4AY7_0),.clk(gclk));
	jdff dff_B_oJtqagUn2_0(.din(w_dff_B_TW7vS4AY7_0),.dout(w_dff_B_oJtqagUn2_0),.clk(gclk));
	jdff dff_B_cQ4vJJdm6_0(.din(w_dff_B_oJtqagUn2_0),.dout(w_dff_B_cQ4vJJdm6_0),.clk(gclk));
	jdff dff_A_xnWN3iB84_1(.dout(w_n1379_0[1]),.din(w_dff_A_xnWN3iB84_1),.clk(gclk));
	jdff dff_A_pSshbNdD7_1(.dout(w_dff_A_xnWN3iB84_1),.din(w_dff_A_pSshbNdD7_1),.clk(gclk));
	jdff dff_A_xpEv0tNt5_1(.dout(w_dff_A_pSshbNdD7_1),.din(w_dff_A_xpEv0tNt5_1),.clk(gclk));
	jdff dff_A_7FZ7qAsX5_1(.dout(w_dff_A_xpEv0tNt5_1),.din(w_dff_A_7FZ7qAsX5_1),.clk(gclk));
	jdff dff_A_uVFeJtGu4_1(.dout(w_dff_A_7FZ7qAsX5_1),.din(w_dff_A_uVFeJtGu4_1),.clk(gclk));
	jdff dff_B_3yIdB2n87_1(.din(n1299),.dout(w_dff_B_3yIdB2n87_1),.clk(gclk));
	jdff dff_B_ARe2uTSg8_1(.din(w_dff_B_3yIdB2n87_1),.dout(w_dff_B_ARe2uTSg8_1),.clk(gclk));
	jdff dff_B_Koc5iBCH3_1(.din(w_dff_B_ARe2uTSg8_1),.dout(w_dff_B_Koc5iBCH3_1),.clk(gclk));
	jdff dff_A_hO5k5axH8_0(.dout(w_n1295_0[0]),.din(w_dff_A_hO5k5axH8_0),.clk(gclk));
	jdff dff_A_J7L0F21u0_0(.dout(w_dff_A_hO5k5axH8_0),.din(w_dff_A_J7L0F21u0_0),.clk(gclk));
	jdff dff_B_ybojhGAX3_1(.din(n1211),.dout(w_dff_B_ybojhGAX3_1),.clk(gclk));
	jdff dff_A_kaFjA6Cr4_0(.dout(w_n1207_0[0]),.din(w_dff_A_kaFjA6Cr4_0),.clk(gclk));
	jdff dff_B_fYgRh1hF7_1(.din(n1113),.dout(w_dff_B_fYgRh1hF7_1),.clk(gclk));
	jdff dff_A_jiOGZly09_1(.dout(w_n1013_0[1]),.din(w_dff_A_jiOGZly09_1),.clk(gclk));
	jdff dff_B_CVkOlKTy6_2(.din(n1011),.dout(w_dff_B_CVkOlKTy6_2),.clk(gclk));
	jdff dff_B_ZO5Jnt0Y5_1(.din(n908),.dout(w_dff_B_ZO5Jnt0Y5_1),.clk(gclk));
	jdff dff_A_BHRY0G6L4_0(.dout(w_n805_0[0]),.din(w_dff_A_BHRY0G6L4_0),.clk(gclk));
	jdff dff_A_wpcAzBN75_0(.dout(w_dff_A_BHRY0G6L4_0),.din(w_dff_A_wpcAzBN75_0),.clk(gclk));
	jdff dff_A_P1kbRSS35_0(.dout(w_dff_A_wpcAzBN75_0),.din(w_dff_A_P1kbRSS35_0),.clk(gclk));
	jdff dff_A_RCxcO2ug9_0(.dout(w_dff_A_P1kbRSS35_0),.din(w_dff_A_RCxcO2ug9_0),.clk(gclk));
	jdff dff_A_LRMM7CMf9_0(.dout(w_dff_A_RCxcO2ug9_0),.din(w_dff_A_LRMM7CMf9_0),.clk(gclk));
	jdff dff_A_GmkW7RrH2_0(.dout(w_dff_A_LRMM7CMf9_0),.din(w_dff_A_GmkW7RrH2_0),.clk(gclk));
	jdff dff_A_TrKXhuUI6_0(.dout(w_dff_A_GmkW7RrH2_0),.din(w_dff_A_TrKXhuUI6_0),.clk(gclk));
	jdff dff_A_0z2Gcrvs8_0(.dout(w_dff_A_TrKXhuUI6_0),.din(w_dff_A_0z2Gcrvs8_0),.clk(gclk));
	jdff dff_A_Y6HhZCh19_0(.dout(w_dff_A_0z2Gcrvs8_0),.din(w_dff_A_Y6HhZCh19_0),.clk(gclk));
	jdff dff_A_o3wO0o3u5_0(.dout(w_dff_A_Y6HhZCh19_0),.din(w_dff_A_o3wO0o3u5_0),.clk(gclk));
	jdff dff_A_LivJCd1u6_0(.dout(w_dff_A_o3wO0o3u5_0),.din(w_dff_A_LivJCd1u6_0),.clk(gclk));
	jdff dff_A_Xe2cx39M6_0(.dout(w_dff_A_LivJCd1u6_0),.din(w_dff_A_Xe2cx39M6_0),.clk(gclk));
	jdff dff_A_YIqSVSig2_0(.dout(w_dff_A_Xe2cx39M6_0),.din(w_dff_A_YIqSVSig2_0),.clk(gclk));
	jdff dff_A_9wrzYiy57_0(.dout(w_dff_A_YIqSVSig2_0),.din(w_dff_A_9wrzYiy57_0),.clk(gclk));
	jdff dff_A_LFKxwgSu4_0(.dout(w_dff_A_9wrzYiy57_0),.din(w_dff_A_LFKxwgSu4_0),.clk(gclk));
	jdff dff_A_g7wEpjmQ2_0(.dout(w_dff_A_LFKxwgSu4_0),.din(w_dff_A_g7wEpjmQ2_0),.clk(gclk));
	jdff dff_A_IHC192zf5_0(.dout(w_dff_A_g7wEpjmQ2_0),.din(w_dff_A_IHC192zf5_0),.clk(gclk));
	jdff dff_A_D7p12W4g6_0(.dout(w_dff_A_IHC192zf5_0),.din(w_dff_A_D7p12W4g6_0),.clk(gclk));
	jdff dff_A_4FcbHW3v2_0(.dout(w_dff_A_D7p12W4g6_0),.din(w_dff_A_4FcbHW3v2_0),.clk(gclk));
	jdff dff_A_0y68ajuR1_0(.dout(w_dff_A_4FcbHW3v2_0),.din(w_dff_A_0y68ajuR1_0),.clk(gclk));
	jdff dff_A_6pzbKutD4_0(.dout(w_dff_A_0y68ajuR1_0),.din(w_dff_A_6pzbKutD4_0),.clk(gclk));
	jdff dff_A_EKGbOPrh9_0(.dout(w_dff_A_6pzbKutD4_0),.din(w_dff_A_EKGbOPrh9_0),.clk(gclk));
	jdff dff_A_q1Gqd3m25_0(.dout(w_dff_A_EKGbOPrh9_0),.din(w_dff_A_q1Gqd3m25_0),.clk(gclk));
	jdff dff_A_8LyXd5j84_0(.dout(w_dff_A_q1Gqd3m25_0),.din(w_dff_A_8LyXd5j84_0),.clk(gclk));
	jdff dff_A_3AOMD8TQ9_0(.dout(w_dff_A_8LyXd5j84_0),.din(w_dff_A_3AOMD8TQ9_0),.clk(gclk));
	jdff dff_A_vQbkMacA7_0(.dout(w_dff_A_3AOMD8TQ9_0),.din(w_dff_A_vQbkMacA7_0),.clk(gclk));
	jdff dff_A_hiFGNQmS1_0(.dout(w_dff_A_vQbkMacA7_0),.din(w_dff_A_hiFGNQmS1_0),.clk(gclk));
	jdff dff_A_jCZtZdpQ0_0(.dout(w_dff_A_hiFGNQmS1_0),.din(w_dff_A_jCZtZdpQ0_0),.clk(gclk));
	jdff dff_A_QE99YOKC2_0(.dout(w_dff_A_jCZtZdpQ0_0),.din(w_dff_A_QE99YOKC2_0),.clk(gclk));
	jdff dff_A_TSglZsyy4_0(.dout(w_dff_A_QE99YOKC2_0),.din(w_dff_A_TSglZsyy4_0),.clk(gclk));
	jdff dff_A_6f52oQ1b9_0(.dout(w_dff_A_TSglZsyy4_0),.din(w_dff_A_6f52oQ1b9_0),.clk(gclk));
	jdff dff_A_JOYxbMpT4_0(.dout(w_dff_A_6f52oQ1b9_0),.din(w_dff_A_JOYxbMpT4_0),.clk(gclk));
	jdff dff_A_AhDiPKMt8_0(.dout(w_dff_A_JOYxbMpT4_0),.din(w_dff_A_AhDiPKMt8_0),.clk(gclk));
	jdff dff_A_kbLrsGem1_0(.dout(w_dff_A_AhDiPKMt8_0),.din(w_dff_A_kbLrsGem1_0),.clk(gclk));
	jdff dff_A_0Hv1oFsx9_0(.dout(w_dff_A_kbLrsGem1_0),.din(w_dff_A_0Hv1oFsx9_0),.clk(gclk));
	jdff dff_A_RGXyUJYb4_0(.dout(w_dff_A_0Hv1oFsx9_0),.din(w_dff_A_RGXyUJYb4_0),.clk(gclk));
	jdff dff_A_QIAOY69L9_0(.dout(w_dff_A_RGXyUJYb4_0),.din(w_dff_A_QIAOY69L9_0),.clk(gclk));
	jdff dff_A_8MlR8qzX8_0(.dout(w_dff_A_QIAOY69L9_0),.din(w_dff_A_8MlR8qzX8_0),.clk(gclk));
	jdff dff_A_suCZ3rK21_0(.dout(w_dff_A_8MlR8qzX8_0),.din(w_dff_A_suCZ3rK21_0),.clk(gclk));
	jdff dff_A_gsJszbJZ1_0(.dout(w_dff_A_suCZ3rK21_0),.din(w_dff_A_gsJszbJZ1_0),.clk(gclk));
	jdff dff_A_6fvcXd5l6_0(.dout(w_dff_A_gsJszbJZ1_0),.din(w_dff_A_6fvcXd5l6_0),.clk(gclk));
	jdff dff_A_gJAijCqu7_0(.dout(w_dff_A_6fvcXd5l6_0),.din(w_dff_A_gJAijCqu7_0),.clk(gclk));
	jdff dff_A_QqOo8jfq1_0(.dout(w_dff_A_gJAijCqu7_0),.din(w_dff_A_QqOo8jfq1_0),.clk(gclk));
	jdff dff_A_7cq0XO5c0_1(.dout(w_n904_0[1]),.din(w_dff_A_7cq0XO5c0_1),.clk(gclk));
	jdff dff_B_2rNmKVuM2_1(.din(n808),.dout(w_dff_B_2rNmKVuM2_1),.clk(gclk));
	jdff dff_A_uoslVDBg8_0(.dout(w_n706_0[0]),.din(w_dff_A_uoslVDBg8_0),.clk(gclk));
	jdff dff_A_zWy9C9333_0(.dout(w_dff_A_uoslVDBg8_0),.din(w_dff_A_zWy9C9333_0),.clk(gclk));
	jdff dff_A_lY29bOSw2_0(.dout(w_dff_A_zWy9C9333_0),.din(w_dff_A_lY29bOSw2_0),.clk(gclk));
	jdff dff_A_gEdXHpU48_0(.dout(w_dff_A_lY29bOSw2_0),.din(w_dff_A_gEdXHpU48_0),.clk(gclk));
	jdff dff_A_0ky2T2yD0_0(.dout(w_dff_A_gEdXHpU48_0),.din(w_dff_A_0ky2T2yD0_0),.clk(gclk));
	jdff dff_A_2UEEXuuF6_0(.dout(w_dff_A_0ky2T2yD0_0),.din(w_dff_A_2UEEXuuF6_0),.clk(gclk));
	jdff dff_A_nBI47ZtZ7_0(.dout(w_dff_A_2UEEXuuF6_0),.din(w_dff_A_nBI47ZtZ7_0),.clk(gclk));
	jdff dff_A_5hDO9RcP7_0(.dout(w_dff_A_nBI47ZtZ7_0),.din(w_dff_A_5hDO9RcP7_0),.clk(gclk));
	jdff dff_A_ho6tuuao7_0(.dout(w_dff_A_5hDO9RcP7_0),.din(w_dff_A_ho6tuuao7_0),.clk(gclk));
	jdff dff_A_EfUSJx668_0(.dout(w_dff_A_ho6tuuao7_0),.din(w_dff_A_EfUSJx668_0),.clk(gclk));
	jdff dff_A_LsyUGUE08_0(.dout(w_dff_A_EfUSJx668_0),.din(w_dff_A_LsyUGUE08_0),.clk(gclk));
	jdff dff_A_jEAMMhjg7_0(.dout(w_dff_A_LsyUGUE08_0),.din(w_dff_A_jEAMMhjg7_0),.clk(gclk));
	jdff dff_A_4QyU7vqQ7_0(.dout(w_dff_A_jEAMMhjg7_0),.din(w_dff_A_4QyU7vqQ7_0),.clk(gclk));
	jdff dff_A_HfpsZWzC6_0(.dout(w_dff_A_4QyU7vqQ7_0),.din(w_dff_A_HfpsZWzC6_0),.clk(gclk));
	jdff dff_A_xCvJr1wS9_0(.dout(w_dff_A_HfpsZWzC6_0),.din(w_dff_A_xCvJr1wS9_0),.clk(gclk));
	jdff dff_A_2AXeviiu6_0(.dout(w_dff_A_xCvJr1wS9_0),.din(w_dff_A_2AXeviiu6_0),.clk(gclk));
	jdff dff_A_4OVFI3vb9_0(.dout(w_dff_A_2AXeviiu6_0),.din(w_dff_A_4OVFI3vb9_0),.clk(gclk));
	jdff dff_A_fVwu7g6j9_0(.dout(w_dff_A_4OVFI3vb9_0),.din(w_dff_A_fVwu7g6j9_0),.clk(gclk));
	jdff dff_A_JnyOuQ9M1_0(.dout(w_dff_A_fVwu7g6j9_0),.din(w_dff_A_JnyOuQ9M1_0),.clk(gclk));
	jdff dff_A_M4R8nM4p8_0(.dout(w_dff_A_JnyOuQ9M1_0),.din(w_dff_A_M4R8nM4p8_0),.clk(gclk));
	jdff dff_A_Sr4zIyDc6_0(.dout(w_dff_A_M4R8nM4p8_0),.din(w_dff_A_Sr4zIyDc6_0),.clk(gclk));
	jdff dff_A_rxkKefHw0_0(.dout(w_dff_A_Sr4zIyDc6_0),.din(w_dff_A_rxkKefHw0_0),.clk(gclk));
	jdff dff_A_OhoYsm5C6_0(.dout(w_dff_A_rxkKefHw0_0),.din(w_dff_A_OhoYsm5C6_0),.clk(gclk));
	jdff dff_A_mEaqBEgc3_0(.dout(w_dff_A_OhoYsm5C6_0),.din(w_dff_A_mEaqBEgc3_0),.clk(gclk));
	jdff dff_A_Ojo1izpC9_0(.dout(w_dff_A_mEaqBEgc3_0),.din(w_dff_A_Ojo1izpC9_0),.clk(gclk));
	jdff dff_A_1WLY8Ti45_0(.dout(w_dff_A_Ojo1izpC9_0),.din(w_dff_A_1WLY8Ti45_0),.clk(gclk));
	jdff dff_A_IOv8kBW68_0(.dout(w_dff_A_1WLY8Ti45_0),.din(w_dff_A_IOv8kBW68_0),.clk(gclk));
	jdff dff_A_5YeZap0Y0_0(.dout(w_dff_A_IOv8kBW68_0),.din(w_dff_A_5YeZap0Y0_0),.clk(gclk));
	jdff dff_A_13EBlcFb1_0(.dout(w_dff_A_5YeZap0Y0_0),.din(w_dff_A_13EBlcFb1_0),.clk(gclk));
	jdff dff_A_sotR9M5P8_0(.dout(w_dff_A_13EBlcFb1_0),.din(w_dff_A_sotR9M5P8_0),.clk(gclk));
	jdff dff_A_8Xlhih6v5_0(.dout(w_dff_A_sotR9M5P8_0),.din(w_dff_A_8Xlhih6v5_0),.clk(gclk));
	jdff dff_A_0pmBw9Or1_0(.dout(w_dff_A_8Xlhih6v5_0),.din(w_dff_A_0pmBw9Or1_0),.clk(gclk));
	jdff dff_A_2YnWPVwZ1_0(.dout(w_dff_A_0pmBw9Or1_0),.din(w_dff_A_2YnWPVwZ1_0),.clk(gclk));
	jdff dff_A_r9xvjQIv1_0(.dout(w_dff_A_2YnWPVwZ1_0),.din(w_dff_A_r9xvjQIv1_0),.clk(gclk));
	jdff dff_A_DVBhDspW3_0(.dout(w_dff_A_r9xvjQIv1_0),.din(w_dff_A_DVBhDspW3_0),.clk(gclk));
	jdff dff_A_bEXCFuCA2_0(.dout(w_dff_A_DVBhDspW3_0),.din(w_dff_A_bEXCFuCA2_0),.clk(gclk));
	jdff dff_A_Dnaihokf7_0(.dout(w_dff_A_bEXCFuCA2_0),.din(w_dff_A_Dnaihokf7_0),.clk(gclk));
	jdff dff_A_T6mgB7AE0_0(.dout(w_dff_A_Dnaihokf7_0),.din(w_dff_A_T6mgB7AE0_0),.clk(gclk));
	jdff dff_A_Ob2Y3P6o2_0(.dout(w_dff_A_T6mgB7AE0_0),.din(w_dff_A_Ob2Y3P6o2_0),.clk(gclk));
	jdff dff_A_N18EMJBx6_0(.dout(w_dff_A_Ob2Y3P6o2_0),.din(w_dff_A_N18EMJBx6_0),.clk(gclk));
	jdff dff_A_eo9lZxUw1_1(.dout(w_n802_0[1]),.din(w_dff_A_eo9lZxUw1_1),.clk(gclk));
	jdff dff_B_KRtJVCPj7_1(.din(n713),.dout(w_dff_B_KRtJVCPj7_1),.clk(gclk));
	jdff dff_B_SkNhUAOP6_1(.din(w_dff_B_KRtJVCPj7_1),.dout(w_dff_B_SkNhUAOP6_1),.clk(gclk));
	jdff dff_B_Pt3fOwyy9_1(.din(w_dff_B_SkNhUAOP6_1),.dout(w_dff_B_Pt3fOwyy9_1),.clk(gclk));
	jdff dff_B_5n8PwDHO6_1(.din(w_dff_B_Pt3fOwyy9_1),.dout(w_dff_B_5n8PwDHO6_1),.clk(gclk));
	jdff dff_B_W9a4W4Wo1_1(.din(w_dff_B_5n8PwDHO6_1),.dout(w_dff_B_W9a4W4Wo1_1),.clk(gclk));
	jdff dff_B_8OsFalwC3_1(.din(w_dff_B_W9a4W4Wo1_1),.dout(w_dff_B_8OsFalwC3_1),.clk(gclk));
	jdff dff_B_tzJsuKty0_1(.din(w_dff_B_8OsFalwC3_1),.dout(w_dff_B_tzJsuKty0_1),.clk(gclk));
	jdff dff_B_QlU18psY4_1(.din(w_dff_B_tzJsuKty0_1),.dout(w_dff_B_QlU18psY4_1),.clk(gclk));
	jdff dff_B_cpNMblWV8_1(.din(w_dff_B_QlU18psY4_1),.dout(w_dff_B_cpNMblWV8_1),.clk(gclk));
	jdff dff_B_mkqVkWJV9_1(.din(w_dff_B_cpNMblWV8_1),.dout(w_dff_B_mkqVkWJV9_1),.clk(gclk));
	jdff dff_B_q58fuMNR0_1(.din(w_dff_B_mkqVkWJV9_1),.dout(w_dff_B_q58fuMNR0_1),.clk(gclk));
	jdff dff_B_J0HIMT0P0_1(.din(w_dff_B_q58fuMNR0_1),.dout(w_dff_B_J0HIMT0P0_1),.clk(gclk));
	jdff dff_B_zYfrQ9Hc6_1(.din(w_dff_B_J0HIMT0P0_1),.dout(w_dff_B_zYfrQ9Hc6_1),.clk(gclk));
	jdff dff_B_pdnRk0Ik7_1(.din(w_dff_B_zYfrQ9Hc6_1),.dout(w_dff_B_pdnRk0Ik7_1),.clk(gclk));
	jdff dff_B_HhqsTWYQ0_1(.din(w_dff_B_pdnRk0Ik7_1),.dout(w_dff_B_HhqsTWYQ0_1),.clk(gclk));
	jdff dff_B_oFf4QXRh8_1(.din(w_dff_B_HhqsTWYQ0_1),.dout(w_dff_B_oFf4QXRh8_1),.clk(gclk));
	jdff dff_B_PDqLJ4RM0_1(.din(w_dff_B_oFf4QXRh8_1),.dout(w_dff_B_PDqLJ4RM0_1),.clk(gclk));
	jdff dff_B_jq8F6DXk1_1(.din(w_dff_B_PDqLJ4RM0_1),.dout(w_dff_B_jq8F6DXk1_1),.clk(gclk));
	jdff dff_B_BvUPDUCv2_1(.din(w_dff_B_jq8F6DXk1_1),.dout(w_dff_B_BvUPDUCv2_1),.clk(gclk));
	jdff dff_B_MXakd8hJ1_1(.din(w_dff_B_BvUPDUCv2_1),.dout(w_dff_B_MXakd8hJ1_1),.clk(gclk));
	jdff dff_B_OTERYf4q8_1(.din(w_dff_B_MXakd8hJ1_1),.dout(w_dff_B_OTERYf4q8_1),.clk(gclk));
	jdff dff_B_QehL6McB4_1(.din(w_dff_B_OTERYf4q8_1),.dout(w_dff_B_QehL6McB4_1),.clk(gclk));
	jdff dff_B_tLCza84k3_1(.din(w_dff_B_QehL6McB4_1),.dout(w_dff_B_tLCza84k3_1),.clk(gclk));
	jdff dff_B_mXNHgVYp6_1(.din(w_dff_B_tLCza84k3_1),.dout(w_dff_B_mXNHgVYp6_1),.clk(gclk));
	jdff dff_B_9pNqoitb1_1(.din(w_dff_B_mXNHgVYp6_1),.dout(w_dff_B_9pNqoitb1_1),.clk(gclk));
	jdff dff_B_hnLjxhIU1_1(.din(w_dff_B_9pNqoitb1_1),.dout(w_dff_B_hnLjxhIU1_1),.clk(gclk));
	jdff dff_B_dQXMrhXN2_1(.din(w_dff_B_hnLjxhIU1_1),.dout(w_dff_B_dQXMrhXN2_1),.clk(gclk));
	jdff dff_B_1zxBwxWi4_1(.din(w_dff_B_dQXMrhXN2_1),.dout(w_dff_B_1zxBwxWi4_1),.clk(gclk));
	jdff dff_B_EH10RSXA9_1(.din(w_dff_B_1zxBwxWi4_1),.dout(w_dff_B_EH10RSXA9_1),.clk(gclk));
	jdff dff_B_26zndpjw6_1(.din(w_dff_B_EH10RSXA9_1),.dout(w_dff_B_26zndpjw6_1),.clk(gclk));
	jdff dff_B_ZA0QdNd89_1(.din(w_dff_B_26zndpjw6_1),.dout(w_dff_B_ZA0QdNd89_1),.clk(gclk));
	jdff dff_B_TMYzmnVo7_1(.din(w_dff_B_ZA0QdNd89_1),.dout(w_dff_B_TMYzmnVo7_1),.clk(gclk));
	jdff dff_B_FcazK6Hj8_1(.din(w_dff_B_TMYzmnVo7_1),.dout(w_dff_B_FcazK6Hj8_1),.clk(gclk));
	jdff dff_B_s9RCwLyC4_1(.din(w_dff_B_FcazK6Hj8_1),.dout(w_dff_B_s9RCwLyC4_1),.clk(gclk));
	jdff dff_B_O4Ixz7Ng6_1(.din(w_dff_B_s9RCwLyC4_1),.dout(w_dff_B_O4Ixz7Ng6_1),.clk(gclk));
	jdff dff_B_6wcSrPEr9_1(.din(w_dff_B_O4Ixz7Ng6_1),.dout(w_dff_B_6wcSrPEr9_1),.clk(gclk));
	jdff dff_B_Xym03pKl7_1(.din(n709),.dout(w_dff_B_Xym03pKl7_1),.clk(gclk));
	jdff dff_A_FGwVRWCg9_0(.dout(w_n614_0[0]),.din(w_dff_A_FGwVRWCg9_0),.clk(gclk));
	jdff dff_A_EJGcBJLE4_0(.dout(w_dff_A_FGwVRWCg9_0),.din(w_dff_A_EJGcBJLE4_0),.clk(gclk));
	jdff dff_A_RBoRpCHR1_0(.dout(w_dff_A_EJGcBJLE4_0),.din(w_dff_A_RBoRpCHR1_0),.clk(gclk));
	jdff dff_A_HHoIQMvM6_0(.dout(w_dff_A_RBoRpCHR1_0),.din(w_dff_A_HHoIQMvM6_0),.clk(gclk));
	jdff dff_A_r7T5RlNr6_0(.dout(w_dff_A_HHoIQMvM6_0),.din(w_dff_A_r7T5RlNr6_0),.clk(gclk));
	jdff dff_A_bmzqZhWS1_0(.dout(w_dff_A_r7T5RlNr6_0),.din(w_dff_A_bmzqZhWS1_0),.clk(gclk));
	jdff dff_A_JNPCvNGk0_0(.dout(w_dff_A_bmzqZhWS1_0),.din(w_dff_A_JNPCvNGk0_0),.clk(gclk));
	jdff dff_A_6kwrgV8p6_0(.dout(w_dff_A_JNPCvNGk0_0),.din(w_dff_A_6kwrgV8p6_0),.clk(gclk));
	jdff dff_A_IMdurQtH8_0(.dout(w_dff_A_6kwrgV8p6_0),.din(w_dff_A_IMdurQtH8_0),.clk(gclk));
	jdff dff_A_CGN8djJ72_0(.dout(w_dff_A_IMdurQtH8_0),.din(w_dff_A_CGN8djJ72_0),.clk(gclk));
	jdff dff_A_ATty5JQI0_0(.dout(w_dff_A_CGN8djJ72_0),.din(w_dff_A_ATty5JQI0_0),.clk(gclk));
	jdff dff_A_PMALUlyS7_0(.dout(w_dff_A_ATty5JQI0_0),.din(w_dff_A_PMALUlyS7_0),.clk(gclk));
	jdff dff_A_8KLsGwWw6_0(.dout(w_dff_A_PMALUlyS7_0),.din(w_dff_A_8KLsGwWw6_0),.clk(gclk));
	jdff dff_A_0YcmvCC04_0(.dout(w_dff_A_8KLsGwWw6_0),.din(w_dff_A_0YcmvCC04_0),.clk(gclk));
	jdff dff_A_WgzJKzss6_0(.dout(w_dff_A_0YcmvCC04_0),.din(w_dff_A_WgzJKzss6_0),.clk(gclk));
	jdff dff_A_hSsYlydL9_0(.dout(w_dff_A_WgzJKzss6_0),.din(w_dff_A_hSsYlydL9_0),.clk(gclk));
	jdff dff_A_vIeHjNLH9_0(.dout(w_dff_A_hSsYlydL9_0),.din(w_dff_A_vIeHjNLH9_0),.clk(gclk));
	jdff dff_A_SSQOAqDK9_0(.dout(w_dff_A_vIeHjNLH9_0),.din(w_dff_A_SSQOAqDK9_0),.clk(gclk));
	jdff dff_A_5rSlmiP55_0(.dout(w_dff_A_SSQOAqDK9_0),.din(w_dff_A_5rSlmiP55_0),.clk(gclk));
	jdff dff_A_SLsPsEKY3_0(.dout(w_dff_A_5rSlmiP55_0),.din(w_dff_A_SLsPsEKY3_0),.clk(gclk));
	jdff dff_A_RrwU77qV7_0(.dout(w_dff_A_SLsPsEKY3_0),.din(w_dff_A_RrwU77qV7_0),.clk(gclk));
	jdff dff_A_ncFlE6jN3_0(.dout(w_dff_A_RrwU77qV7_0),.din(w_dff_A_ncFlE6jN3_0),.clk(gclk));
	jdff dff_A_bHUUfagv2_0(.dout(w_dff_A_ncFlE6jN3_0),.din(w_dff_A_bHUUfagv2_0),.clk(gclk));
	jdff dff_A_YsItLTIa6_0(.dout(w_dff_A_bHUUfagv2_0),.din(w_dff_A_YsItLTIa6_0),.clk(gclk));
	jdff dff_A_La0IhG493_0(.dout(w_dff_A_YsItLTIa6_0),.din(w_dff_A_La0IhG493_0),.clk(gclk));
	jdff dff_A_zyJjB6n00_0(.dout(w_dff_A_La0IhG493_0),.din(w_dff_A_zyJjB6n00_0),.clk(gclk));
	jdff dff_A_LTvM492u1_0(.dout(w_dff_A_zyJjB6n00_0),.din(w_dff_A_LTvM492u1_0),.clk(gclk));
	jdff dff_A_lYeOZ6IH2_0(.dout(w_dff_A_LTvM492u1_0),.din(w_dff_A_lYeOZ6IH2_0),.clk(gclk));
	jdff dff_A_WNnuKsmE2_0(.dout(w_dff_A_lYeOZ6IH2_0),.din(w_dff_A_WNnuKsmE2_0),.clk(gclk));
	jdff dff_A_rNzVcCAP3_0(.dout(w_dff_A_WNnuKsmE2_0),.din(w_dff_A_rNzVcCAP3_0),.clk(gclk));
	jdff dff_A_vkFHbpTP2_0(.dout(w_dff_A_rNzVcCAP3_0),.din(w_dff_A_vkFHbpTP2_0),.clk(gclk));
	jdff dff_A_G6tQPmgk4_0(.dout(w_dff_A_vkFHbpTP2_0),.din(w_dff_A_G6tQPmgk4_0),.clk(gclk));
	jdff dff_A_TsaPcj4A5_0(.dout(w_dff_A_G6tQPmgk4_0),.din(w_dff_A_TsaPcj4A5_0),.clk(gclk));
	jdff dff_A_GbHM12Y08_0(.dout(w_dff_A_TsaPcj4A5_0),.din(w_dff_A_GbHM12Y08_0),.clk(gclk));
	jdff dff_A_XqJgMGV55_0(.dout(w_dff_A_GbHM12Y08_0),.din(w_dff_A_XqJgMGV55_0),.clk(gclk));
	jdff dff_A_cPQU0PL80_0(.dout(w_dff_A_XqJgMGV55_0),.din(w_dff_A_cPQU0PL80_0),.clk(gclk));
	jdff dff_A_CEOAP1Il9_0(.dout(w_dff_A_cPQU0PL80_0),.din(w_dff_A_CEOAP1Il9_0),.clk(gclk));
	jdff dff_A_WtcaqWte1_1(.dout(w_n703_0[1]),.din(w_dff_A_WtcaqWte1_1),.clk(gclk));
	jdff dff_B_6SyICT3r3_1(.din(n621),.dout(w_dff_B_6SyICT3r3_1),.clk(gclk));
	jdff dff_B_zc7ZRKXU9_1(.din(w_dff_B_6SyICT3r3_1),.dout(w_dff_B_zc7ZRKXU9_1),.clk(gclk));
	jdff dff_B_0bzIwj9I4_1(.din(w_dff_B_zc7ZRKXU9_1),.dout(w_dff_B_0bzIwj9I4_1),.clk(gclk));
	jdff dff_B_CpnOqE7C3_1(.din(w_dff_B_0bzIwj9I4_1),.dout(w_dff_B_CpnOqE7C3_1),.clk(gclk));
	jdff dff_B_pYBHqoFn1_1(.din(w_dff_B_CpnOqE7C3_1),.dout(w_dff_B_pYBHqoFn1_1),.clk(gclk));
	jdff dff_B_tAaFqgc84_1(.din(w_dff_B_pYBHqoFn1_1),.dout(w_dff_B_tAaFqgc84_1),.clk(gclk));
	jdff dff_B_2xQqBtlx1_1(.din(w_dff_B_tAaFqgc84_1),.dout(w_dff_B_2xQqBtlx1_1),.clk(gclk));
	jdff dff_B_uZet1faX3_1(.din(w_dff_B_2xQqBtlx1_1),.dout(w_dff_B_uZet1faX3_1),.clk(gclk));
	jdff dff_B_0SWNfy8y3_1(.din(w_dff_B_uZet1faX3_1),.dout(w_dff_B_0SWNfy8y3_1),.clk(gclk));
	jdff dff_B_CLQmzCwo2_1(.din(w_dff_B_0SWNfy8y3_1),.dout(w_dff_B_CLQmzCwo2_1),.clk(gclk));
	jdff dff_B_BPdERJ4A5_1(.din(w_dff_B_CLQmzCwo2_1),.dout(w_dff_B_BPdERJ4A5_1),.clk(gclk));
	jdff dff_B_Pa7lDxO18_1(.din(w_dff_B_BPdERJ4A5_1),.dout(w_dff_B_Pa7lDxO18_1),.clk(gclk));
	jdff dff_B_WssyBeGf5_1(.din(w_dff_B_Pa7lDxO18_1),.dout(w_dff_B_WssyBeGf5_1),.clk(gclk));
	jdff dff_B_cTch3KW05_1(.din(w_dff_B_WssyBeGf5_1),.dout(w_dff_B_cTch3KW05_1),.clk(gclk));
	jdff dff_B_J5E5CX8w7_1(.din(w_dff_B_cTch3KW05_1),.dout(w_dff_B_J5E5CX8w7_1),.clk(gclk));
	jdff dff_B_U47cGXxX3_1(.din(w_dff_B_J5E5CX8w7_1),.dout(w_dff_B_U47cGXxX3_1),.clk(gclk));
	jdff dff_B_yy7jdFRp9_1(.din(w_dff_B_U47cGXxX3_1),.dout(w_dff_B_yy7jdFRp9_1),.clk(gclk));
	jdff dff_B_2ZKnmGzf5_1(.din(w_dff_B_yy7jdFRp9_1),.dout(w_dff_B_2ZKnmGzf5_1),.clk(gclk));
	jdff dff_B_2XQENLZS6_1(.din(w_dff_B_2ZKnmGzf5_1),.dout(w_dff_B_2XQENLZS6_1),.clk(gclk));
	jdff dff_B_7aU93EXp4_1(.din(w_dff_B_2XQENLZS6_1),.dout(w_dff_B_7aU93EXp4_1),.clk(gclk));
	jdff dff_B_VD49i5sc8_1(.din(w_dff_B_7aU93EXp4_1),.dout(w_dff_B_VD49i5sc8_1),.clk(gclk));
	jdff dff_B_xQ9J6wBl5_1(.din(w_dff_B_VD49i5sc8_1),.dout(w_dff_B_xQ9J6wBl5_1),.clk(gclk));
	jdff dff_B_WrYBGyXo8_1(.din(w_dff_B_xQ9J6wBl5_1),.dout(w_dff_B_WrYBGyXo8_1),.clk(gclk));
	jdff dff_B_kGvVOY530_1(.din(w_dff_B_WrYBGyXo8_1),.dout(w_dff_B_kGvVOY530_1),.clk(gclk));
	jdff dff_B_p5LiN9Fo0_1(.din(w_dff_B_kGvVOY530_1),.dout(w_dff_B_p5LiN9Fo0_1),.clk(gclk));
	jdff dff_B_XeT5F3Px7_1(.din(w_dff_B_p5LiN9Fo0_1),.dout(w_dff_B_XeT5F3Px7_1),.clk(gclk));
	jdff dff_B_DOBIEwb76_1(.din(w_dff_B_XeT5F3Px7_1),.dout(w_dff_B_DOBIEwb76_1),.clk(gclk));
	jdff dff_B_OTbd4oDl6_1(.din(w_dff_B_DOBIEwb76_1),.dout(w_dff_B_OTbd4oDl6_1),.clk(gclk));
	jdff dff_B_I8bgpPvD4_1(.din(w_dff_B_OTbd4oDl6_1),.dout(w_dff_B_I8bgpPvD4_1),.clk(gclk));
	jdff dff_B_4AR1He6A7_1(.din(w_dff_B_I8bgpPvD4_1),.dout(w_dff_B_4AR1He6A7_1),.clk(gclk));
	jdff dff_B_Uf638gyY1_1(.din(w_dff_B_4AR1He6A7_1),.dout(w_dff_B_Uf638gyY1_1),.clk(gclk));
	jdff dff_B_XRfW8VhR6_1(.din(w_dff_B_Uf638gyY1_1),.dout(w_dff_B_XRfW8VhR6_1),.clk(gclk));
	jdff dff_B_GvGucZMJ3_1(.din(w_dff_B_XRfW8VhR6_1),.dout(w_dff_B_GvGucZMJ3_1),.clk(gclk));
	jdff dff_B_gDaYprKw4_1(.din(n617),.dout(w_dff_B_gDaYprKw4_1),.clk(gclk));
	jdff dff_A_4JA57ErZ2_0(.dout(w_n529_0[0]),.din(w_dff_A_4JA57ErZ2_0),.clk(gclk));
	jdff dff_A_4rijDBqq0_0(.dout(w_dff_A_4JA57ErZ2_0),.din(w_dff_A_4rijDBqq0_0),.clk(gclk));
	jdff dff_A_xhNGnLFM1_0(.dout(w_dff_A_4rijDBqq0_0),.din(w_dff_A_xhNGnLFM1_0),.clk(gclk));
	jdff dff_A_GZrW29ii7_0(.dout(w_dff_A_xhNGnLFM1_0),.din(w_dff_A_GZrW29ii7_0),.clk(gclk));
	jdff dff_A_BAOEhlF92_0(.dout(w_dff_A_GZrW29ii7_0),.din(w_dff_A_BAOEhlF92_0),.clk(gclk));
	jdff dff_A_kRYDu1yu0_0(.dout(w_dff_A_BAOEhlF92_0),.din(w_dff_A_kRYDu1yu0_0),.clk(gclk));
	jdff dff_A_Oi2TLuuA0_0(.dout(w_dff_A_kRYDu1yu0_0),.din(w_dff_A_Oi2TLuuA0_0),.clk(gclk));
	jdff dff_A_fqhrYLO25_0(.dout(w_dff_A_Oi2TLuuA0_0),.din(w_dff_A_fqhrYLO25_0),.clk(gclk));
	jdff dff_A_w1NaCkg98_0(.dout(w_dff_A_fqhrYLO25_0),.din(w_dff_A_w1NaCkg98_0),.clk(gclk));
	jdff dff_A_jxxPaWK55_0(.dout(w_dff_A_w1NaCkg98_0),.din(w_dff_A_jxxPaWK55_0),.clk(gclk));
	jdff dff_A_0uN47Fnk6_0(.dout(w_dff_A_jxxPaWK55_0),.din(w_dff_A_0uN47Fnk6_0),.clk(gclk));
	jdff dff_A_UXHYIZEl4_0(.dout(w_dff_A_0uN47Fnk6_0),.din(w_dff_A_UXHYIZEl4_0),.clk(gclk));
	jdff dff_A_w4iiWhvu1_0(.dout(w_dff_A_UXHYIZEl4_0),.din(w_dff_A_w4iiWhvu1_0),.clk(gclk));
	jdff dff_A_LpeGGcxZ3_0(.dout(w_dff_A_w4iiWhvu1_0),.din(w_dff_A_LpeGGcxZ3_0),.clk(gclk));
	jdff dff_A_FWFJcQop7_0(.dout(w_dff_A_LpeGGcxZ3_0),.din(w_dff_A_FWFJcQop7_0),.clk(gclk));
	jdff dff_A_Ifu3STPv1_0(.dout(w_dff_A_FWFJcQop7_0),.din(w_dff_A_Ifu3STPv1_0),.clk(gclk));
	jdff dff_A_4YkROka03_0(.dout(w_dff_A_Ifu3STPv1_0),.din(w_dff_A_4YkROka03_0),.clk(gclk));
	jdff dff_A_iDS9mbmt7_0(.dout(w_dff_A_4YkROka03_0),.din(w_dff_A_iDS9mbmt7_0),.clk(gclk));
	jdff dff_A_czW4u29l3_0(.dout(w_dff_A_iDS9mbmt7_0),.din(w_dff_A_czW4u29l3_0),.clk(gclk));
	jdff dff_A_l0799hok5_0(.dout(w_dff_A_czW4u29l3_0),.din(w_dff_A_l0799hok5_0),.clk(gclk));
	jdff dff_A_iXQZhpRQ8_0(.dout(w_dff_A_l0799hok5_0),.din(w_dff_A_iXQZhpRQ8_0),.clk(gclk));
	jdff dff_A_DKSkIHZw6_0(.dout(w_dff_A_iXQZhpRQ8_0),.din(w_dff_A_DKSkIHZw6_0),.clk(gclk));
	jdff dff_A_rUkZxJ0X8_0(.dout(w_dff_A_DKSkIHZw6_0),.din(w_dff_A_rUkZxJ0X8_0),.clk(gclk));
	jdff dff_A_Ap06mBVh1_0(.dout(w_dff_A_rUkZxJ0X8_0),.din(w_dff_A_Ap06mBVh1_0),.clk(gclk));
	jdff dff_A_66OlGLJO1_0(.dout(w_dff_A_Ap06mBVh1_0),.din(w_dff_A_66OlGLJO1_0),.clk(gclk));
	jdff dff_A_z14vIt9g8_0(.dout(w_dff_A_66OlGLJO1_0),.din(w_dff_A_z14vIt9g8_0),.clk(gclk));
	jdff dff_A_RrB7piCl6_0(.dout(w_dff_A_z14vIt9g8_0),.din(w_dff_A_RrB7piCl6_0),.clk(gclk));
	jdff dff_A_D9IVdaYP7_0(.dout(w_dff_A_RrB7piCl6_0),.din(w_dff_A_D9IVdaYP7_0),.clk(gclk));
	jdff dff_A_CfPw4iH52_0(.dout(w_dff_A_D9IVdaYP7_0),.din(w_dff_A_CfPw4iH52_0),.clk(gclk));
	jdff dff_A_OWeJAIRQ9_0(.dout(w_dff_A_CfPw4iH52_0),.din(w_dff_A_OWeJAIRQ9_0),.clk(gclk));
	jdff dff_A_YAyVEApa5_0(.dout(w_dff_A_OWeJAIRQ9_0),.din(w_dff_A_YAyVEApa5_0),.clk(gclk));
	jdff dff_A_RSbttYl69_0(.dout(w_dff_A_YAyVEApa5_0),.din(w_dff_A_RSbttYl69_0),.clk(gclk));
	jdff dff_A_MdNDT2Xl1_0(.dout(w_dff_A_RSbttYl69_0),.din(w_dff_A_MdNDT2Xl1_0),.clk(gclk));
	jdff dff_A_mEqOSiLQ7_0(.dout(w_dff_A_MdNDT2Xl1_0),.din(w_dff_A_mEqOSiLQ7_0),.clk(gclk));
	jdff dff_A_ISeNVaNj6_1(.dout(w_n611_0[1]),.din(w_dff_A_ISeNVaNj6_1),.clk(gclk));
	jdff dff_B_ne3tCZix4_1(.din(n536),.dout(w_dff_B_ne3tCZix4_1),.clk(gclk));
	jdff dff_B_phupOrTO3_1(.din(w_dff_B_ne3tCZix4_1),.dout(w_dff_B_phupOrTO3_1),.clk(gclk));
	jdff dff_B_7C3TQTWm9_1(.din(w_dff_B_phupOrTO3_1),.dout(w_dff_B_7C3TQTWm9_1),.clk(gclk));
	jdff dff_B_EtcckvmZ5_1(.din(w_dff_B_7C3TQTWm9_1),.dout(w_dff_B_EtcckvmZ5_1),.clk(gclk));
	jdff dff_B_G4U64aVO7_1(.din(w_dff_B_EtcckvmZ5_1),.dout(w_dff_B_G4U64aVO7_1),.clk(gclk));
	jdff dff_B_sM15BQ009_1(.din(w_dff_B_G4U64aVO7_1),.dout(w_dff_B_sM15BQ009_1),.clk(gclk));
	jdff dff_B_AzuYEjPK2_1(.din(w_dff_B_sM15BQ009_1),.dout(w_dff_B_AzuYEjPK2_1),.clk(gclk));
	jdff dff_B_JGkZPThU5_1(.din(w_dff_B_AzuYEjPK2_1),.dout(w_dff_B_JGkZPThU5_1),.clk(gclk));
	jdff dff_B_23pPFu9Z4_1(.din(w_dff_B_JGkZPThU5_1),.dout(w_dff_B_23pPFu9Z4_1),.clk(gclk));
	jdff dff_B_cQFhJUDS3_1(.din(w_dff_B_23pPFu9Z4_1),.dout(w_dff_B_cQFhJUDS3_1),.clk(gclk));
	jdff dff_B_p2mqKVMX0_1(.din(w_dff_B_cQFhJUDS3_1),.dout(w_dff_B_p2mqKVMX0_1),.clk(gclk));
	jdff dff_B_6tXR47171_1(.din(w_dff_B_p2mqKVMX0_1),.dout(w_dff_B_6tXR47171_1),.clk(gclk));
	jdff dff_B_TUu0ZKo81_1(.din(w_dff_B_6tXR47171_1),.dout(w_dff_B_TUu0ZKo81_1),.clk(gclk));
	jdff dff_B_kqQ9lN4g8_1(.din(w_dff_B_TUu0ZKo81_1),.dout(w_dff_B_kqQ9lN4g8_1),.clk(gclk));
	jdff dff_B_d69QeIeX9_1(.din(w_dff_B_kqQ9lN4g8_1),.dout(w_dff_B_d69QeIeX9_1),.clk(gclk));
	jdff dff_B_NaqEPx3J0_1(.din(w_dff_B_d69QeIeX9_1),.dout(w_dff_B_NaqEPx3J0_1),.clk(gclk));
	jdff dff_B_gp3UP3RY5_1(.din(w_dff_B_NaqEPx3J0_1),.dout(w_dff_B_gp3UP3RY5_1),.clk(gclk));
	jdff dff_B_ub8Uo2Id6_1(.din(w_dff_B_gp3UP3RY5_1),.dout(w_dff_B_ub8Uo2Id6_1),.clk(gclk));
	jdff dff_B_PHXdFdkm2_1(.din(w_dff_B_ub8Uo2Id6_1),.dout(w_dff_B_PHXdFdkm2_1),.clk(gclk));
	jdff dff_B_1OiyW2Kp0_1(.din(w_dff_B_PHXdFdkm2_1),.dout(w_dff_B_1OiyW2Kp0_1),.clk(gclk));
	jdff dff_B_nW7ctQvP8_1(.din(w_dff_B_1OiyW2Kp0_1),.dout(w_dff_B_nW7ctQvP8_1),.clk(gclk));
	jdff dff_B_A43KquRh1_1(.din(w_dff_B_nW7ctQvP8_1),.dout(w_dff_B_A43KquRh1_1),.clk(gclk));
	jdff dff_B_HbziTMfy1_1(.din(w_dff_B_A43KquRh1_1),.dout(w_dff_B_HbziTMfy1_1),.clk(gclk));
	jdff dff_B_7O4IIOVB5_1(.din(w_dff_B_HbziTMfy1_1),.dout(w_dff_B_7O4IIOVB5_1),.clk(gclk));
	jdff dff_B_f7HCLSeY0_1(.din(w_dff_B_7O4IIOVB5_1),.dout(w_dff_B_f7HCLSeY0_1),.clk(gclk));
	jdff dff_B_wjf1W34s0_1(.din(w_dff_B_f7HCLSeY0_1),.dout(w_dff_B_wjf1W34s0_1),.clk(gclk));
	jdff dff_B_UOBfBc6k4_1(.din(w_dff_B_wjf1W34s0_1),.dout(w_dff_B_UOBfBc6k4_1),.clk(gclk));
	jdff dff_B_QYZyfPO62_1(.din(w_dff_B_UOBfBc6k4_1),.dout(w_dff_B_QYZyfPO62_1),.clk(gclk));
	jdff dff_B_Qw7lEFNL7_1(.din(w_dff_B_QYZyfPO62_1),.dout(w_dff_B_Qw7lEFNL7_1),.clk(gclk));
	jdff dff_B_NRDofYYa6_1(.din(w_dff_B_Qw7lEFNL7_1),.dout(w_dff_B_NRDofYYa6_1),.clk(gclk));
	jdff dff_B_7wRTG4kK2_1(.din(n532),.dout(w_dff_B_7wRTG4kK2_1),.clk(gclk));
	jdff dff_A_a8Fwb5RZ4_0(.dout(w_n451_0[0]),.din(w_dff_A_a8Fwb5RZ4_0),.clk(gclk));
	jdff dff_A_TyAhhCyJ2_0(.dout(w_dff_A_a8Fwb5RZ4_0),.din(w_dff_A_TyAhhCyJ2_0),.clk(gclk));
	jdff dff_A_wfj6IsTs4_0(.dout(w_dff_A_TyAhhCyJ2_0),.din(w_dff_A_wfj6IsTs4_0),.clk(gclk));
	jdff dff_A_ITadPbkD3_0(.dout(w_dff_A_wfj6IsTs4_0),.din(w_dff_A_ITadPbkD3_0),.clk(gclk));
	jdff dff_A_yPNTjDHC3_0(.dout(w_dff_A_ITadPbkD3_0),.din(w_dff_A_yPNTjDHC3_0),.clk(gclk));
	jdff dff_A_PEkuYYf89_0(.dout(w_dff_A_yPNTjDHC3_0),.din(w_dff_A_PEkuYYf89_0),.clk(gclk));
	jdff dff_A_z3YKOYsy5_0(.dout(w_dff_A_PEkuYYf89_0),.din(w_dff_A_z3YKOYsy5_0),.clk(gclk));
	jdff dff_A_Nvfqj2z84_0(.dout(w_dff_A_z3YKOYsy5_0),.din(w_dff_A_Nvfqj2z84_0),.clk(gclk));
	jdff dff_A_l8qElnG82_0(.dout(w_dff_A_Nvfqj2z84_0),.din(w_dff_A_l8qElnG82_0),.clk(gclk));
	jdff dff_A_AfynoxTc3_0(.dout(w_dff_A_l8qElnG82_0),.din(w_dff_A_AfynoxTc3_0),.clk(gclk));
	jdff dff_A_pTqbHSPV1_0(.dout(w_dff_A_AfynoxTc3_0),.din(w_dff_A_pTqbHSPV1_0),.clk(gclk));
	jdff dff_A_VMEOnLgi9_0(.dout(w_dff_A_pTqbHSPV1_0),.din(w_dff_A_VMEOnLgi9_0),.clk(gclk));
	jdff dff_A_018a6RRB4_0(.dout(w_dff_A_VMEOnLgi9_0),.din(w_dff_A_018a6RRB4_0),.clk(gclk));
	jdff dff_A_nwjoImeu3_0(.dout(w_dff_A_018a6RRB4_0),.din(w_dff_A_nwjoImeu3_0),.clk(gclk));
	jdff dff_A_qVk9fyOs2_0(.dout(w_dff_A_nwjoImeu3_0),.din(w_dff_A_qVk9fyOs2_0),.clk(gclk));
	jdff dff_A_gK6cTBAU6_0(.dout(w_dff_A_qVk9fyOs2_0),.din(w_dff_A_gK6cTBAU6_0),.clk(gclk));
	jdff dff_A_fcRJirG81_0(.dout(w_dff_A_gK6cTBAU6_0),.din(w_dff_A_fcRJirG81_0),.clk(gclk));
	jdff dff_A_th70luBO7_0(.dout(w_dff_A_fcRJirG81_0),.din(w_dff_A_th70luBO7_0),.clk(gclk));
	jdff dff_A_plS3fxfc6_0(.dout(w_dff_A_th70luBO7_0),.din(w_dff_A_plS3fxfc6_0),.clk(gclk));
	jdff dff_A_Oed7hk8V7_0(.dout(w_dff_A_plS3fxfc6_0),.din(w_dff_A_Oed7hk8V7_0),.clk(gclk));
	jdff dff_A_zZPHYFOA2_0(.dout(w_dff_A_Oed7hk8V7_0),.din(w_dff_A_zZPHYFOA2_0),.clk(gclk));
	jdff dff_A_HEEn2e2t3_0(.dout(w_dff_A_zZPHYFOA2_0),.din(w_dff_A_HEEn2e2t3_0),.clk(gclk));
	jdff dff_A_8ajl39RZ5_0(.dout(w_dff_A_HEEn2e2t3_0),.din(w_dff_A_8ajl39RZ5_0),.clk(gclk));
	jdff dff_A_AZwe0iB83_0(.dout(w_dff_A_8ajl39RZ5_0),.din(w_dff_A_AZwe0iB83_0),.clk(gclk));
	jdff dff_A_GgQ0PZpw2_0(.dout(w_dff_A_AZwe0iB83_0),.din(w_dff_A_GgQ0PZpw2_0),.clk(gclk));
	jdff dff_A_VbVH6lDI6_0(.dout(w_dff_A_GgQ0PZpw2_0),.din(w_dff_A_VbVH6lDI6_0),.clk(gclk));
	jdff dff_A_un1r5UeO9_0(.dout(w_dff_A_VbVH6lDI6_0),.din(w_dff_A_un1r5UeO9_0),.clk(gclk));
	jdff dff_A_L4UuEmJk4_0(.dout(w_dff_A_un1r5UeO9_0),.din(w_dff_A_L4UuEmJk4_0),.clk(gclk));
	jdff dff_A_7j7km2QS2_0(.dout(w_dff_A_L4UuEmJk4_0),.din(w_dff_A_7j7km2QS2_0),.clk(gclk));
	jdff dff_A_nYcqxPaO9_0(.dout(w_dff_A_7j7km2QS2_0),.din(w_dff_A_nYcqxPaO9_0),.clk(gclk));
	jdff dff_A_YkPo2Xyi0_0(.dout(w_dff_A_nYcqxPaO9_0),.din(w_dff_A_YkPo2Xyi0_0),.clk(gclk));
	jdff dff_A_SLB4Z28D3_1(.dout(w_n526_0[1]),.din(w_dff_A_SLB4Z28D3_1),.clk(gclk));
	jdff dff_B_KVsXI5t10_1(.din(n458),.dout(w_dff_B_KVsXI5t10_1),.clk(gclk));
	jdff dff_B_uhLZpc4R5_1(.din(w_dff_B_KVsXI5t10_1),.dout(w_dff_B_uhLZpc4R5_1),.clk(gclk));
	jdff dff_B_TAReCawD2_1(.din(w_dff_B_uhLZpc4R5_1),.dout(w_dff_B_TAReCawD2_1),.clk(gclk));
	jdff dff_B_Hm4SJaXH4_1(.din(w_dff_B_TAReCawD2_1),.dout(w_dff_B_Hm4SJaXH4_1),.clk(gclk));
	jdff dff_B_zJCXU40K9_1(.din(w_dff_B_Hm4SJaXH4_1),.dout(w_dff_B_zJCXU40K9_1),.clk(gclk));
	jdff dff_B_63lPQyr87_1(.din(w_dff_B_zJCXU40K9_1),.dout(w_dff_B_63lPQyr87_1),.clk(gclk));
	jdff dff_B_VJHijFr08_1(.din(w_dff_B_63lPQyr87_1),.dout(w_dff_B_VJHijFr08_1),.clk(gclk));
	jdff dff_B_f2JXMnTy5_1(.din(w_dff_B_VJHijFr08_1),.dout(w_dff_B_f2JXMnTy5_1),.clk(gclk));
	jdff dff_B_zF69YUCj7_1(.din(w_dff_B_f2JXMnTy5_1),.dout(w_dff_B_zF69YUCj7_1),.clk(gclk));
	jdff dff_B_oM0crne45_1(.din(w_dff_B_zF69YUCj7_1),.dout(w_dff_B_oM0crne45_1),.clk(gclk));
	jdff dff_B_HHSEyHm83_1(.din(w_dff_B_oM0crne45_1),.dout(w_dff_B_HHSEyHm83_1),.clk(gclk));
	jdff dff_B_2BYuB0uB1_1(.din(w_dff_B_HHSEyHm83_1),.dout(w_dff_B_2BYuB0uB1_1),.clk(gclk));
	jdff dff_B_ZjYasMWt8_1(.din(w_dff_B_2BYuB0uB1_1),.dout(w_dff_B_ZjYasMWt8_1),.clk(gclk));
	jdff dff_B_B56FRRMA6_1(.din(w_dff_B_ZjYasMWt8_1),.dout(w_dff_B_B56FRRMA6_1),.clk(gclk));
	jdff dff_B_KJAC98oo5_1(.din(w_dff_B_B56FRRMA6_1),.dout(w_dff_B_KJAC98oo5_1),.clk(gclk));
	jdff dff_B_DWT7UjjS2_1(.din(w_dff_B_KJAC98oo5_1),.dout(w_dff_B_DWT7UjjS2_1),.clk(gclk));
	jdff dff_B_3k25Bayc1_1(.din(w_dff_B_DWT7UjjS2_1),.dout(w_dff_B_3k25Bayc1_1),.clk(gclk));
	jdff dff_B_HaEkyVTz3_1(.din(w_dff_B_3k25Bayc1_1),.dout(w_dff_B_HaEkyVTz3_1),.clk(gclk));
	jdff dff_B_lwac3JkV3_1(.din(w_dff_B_HaEkyVTz3_1),.dout(w_dff_B_lwac3JkV3_1),.clk(gclk));
	jdff dff_B_WETmanAY0_1(.din(w_dff_B_lwac3JkV3_1),.dout(w_dff_B_WETmanAY0_1),.clk(gclk));
	jdff dff_B_EjNMBUc71_1(.din(w_dff_B_WETmanAY0_1),.dout(w_dff_B_EjNMBUc71_1),.clk(gclk));
	jdff dff_B_q9ZMHwLB5_1(.din(w_dff_B_EjNMBUc71_1),.dout(w_dff_B_q9ZMHwLB5_1),.clk(gclk));
	jdff dff_B_LGgs0VRt4_1(.din(w_dff_B_q9ZMHwLB5_1),.dout(w_dff_B_LGgs0VRt4_1),.clk(gclk));
	jdff dff_B_mfJ2Qxfl4_1(.din(w_dff_B_LGgs0VRt4_1),.dout(w_dff_B_mfJ2Qxfl4_1),.clk(gclk));
	jdff dff_B_6E035ANg8_1(.din(w_dff_B_mfJ2Qxfl4_1),.dout(w_dff_B_6E035ANg8_1),.clk(gclk));
	jdff dff_B_bDqslVgs1_1(.din(w_dff_B_6E035ANg8_1),.dout(w_dff_B_bDqslVgs1_1),.clk(gclk));
	jdff dff_B_KH04q8iw5_1(.din(w_dff_B_bDqslVgs1_1),.dout(w_dff_B_KH04q8iw5_1),.clk(gclk));
	jdff dff_B_yG4BhU3r1_1(.din(n454),.dout(w_dff_B_yG4BhU3r1_1),.clk(gclk));
	jdff dff_A_YmAFLElN3_0(.dout(w_n380_0[0]),.din(w_dff_A_YmAFLElN3_0),.clk(gclk));
	jdff dff_A_rCzgkMsT7_0(.dout(w_dff_A_YmAFLElN3_0),.din(w_dff_A_rCzgkMsT7_0),.clk(gclk));
	jdff dff_A_MaXF1dXn4_0(.dout(w_dff_A_rCzgkMsT7_0),.din(w_dff_A_MaXF1dXn4_0),.clk(gclk));
	jdff dff_A_aKlxPGwU8_0(.dout(w_dff_A_MaXF1dXn4_0),.din(w_dff_A_aKlxPGwU8_0),.clk(gclk));
	jdff dff_A_GHNJICnn8_0(.dout(w_dff_A_aKlxPGwU8_0),.din(w_dff_A_GHNJICnn8_0),.clk(gclk));
	jdff dff_A_fsfAiiJf9_0(.dout(w_dff_A_GHNJICnn8_0),.din(w_dff_A_fsfAiiJf9_0),.clk(gclk));
	jdff dff_A_3OoPisMW8_0(.dout(w_dff_A_fsfAiiJf9_0),.din(w_dff_A_3OoPisMW8_0),.clk(gclk));
	jdff dff_A_B69rtH2e2_0(.dout(w_dff_A_3OoPisMW8_0),.din(w_dff_A_B69rtH2e2_0),.clk(gclk));
	jdff dff_A_UyXZTCIt6_0(.dout(w_dff_A_B69rtH2e2_0),.din(w_dff_A_UyXZTCIt6_0),.clk(gclk));
	jdff dff_A_jfWBjy941_0(.dout(w_dff_A_UyXZTCIt6_0),.din(w_dff_A_jfWBjy941_0),.clk(gclk));
	jdff dff_A_8MroAHsf3_0(.dout(w_dff_A_jfWBjy941_0),.din(w_dff_A_8MroAHsf3_0),.clk(gclk));
	jdff dff_A_wpRmbtLm3_0(.dout(w_dff_A_8MroAHsf3_0),.din(w_dff_A_wpRmbtLm3_0),.clk(gclk));
	jdff dff_A_mgEwifOG1_0(.dout(w_dff_A_wpRmbtLm3_0),.din(w_dff_A_mgEwifOG1_0),.clk(gclk));
	jdff dff_A_dn9v5nAG5_0(.dout(w_dff_A_mgEwifOG1_0),.din(w_dff_A_dn9v5nAG5_0),.clk(gclk));
	jdff dff_A_e3Fxy71B5_0(.dout(w_dff_A_dn9v5nAG5_0),.din(w_dff_A_e3Fxy71B5_0),.clk(gclk));
	jdff dff_A_WNTsDQSh0_0(.dout(w_dff_A_e3Fxy71B5_0),.din(w_dff_A_WNTsDQSh0_0),.clk(gclk));
	jdff dff_A_qBVO1gIB2_0(.dout(w_dff_A_WNTsDQSh0_0),.din(w_dff_A_qBVO1gIB2_0),.clk(gclk));
	jdff dff_A_9wPQLlci9_0(.dout(w_dff_A_qBVO1gIB2_0),.din(w_dff_A_9wPQLlci9_0),.clk(gclk));
	jdff dff_A_TU7BpV7D4_0(.dout(w_dff_A_9wPQLlci9_0),.din(w_dff_A_TU7BpV7D4_0),.clk(gclk));
	jdff dff_A_9c7n4xI33_0(.dout(w_dff_A_TU7BpV7D4_0),.din(w_dff_A_9c7n4xI33_0),.clk(gclk));
	jdff dff_A_Ff3Shiyc3_0(.dout(w_dff_A_9c7n4xI33_0),.din(w_dff_A_Ff3Shiyc3_0),.clk(gclk));
	jdff dff_A_8qoe3A5D4_0(.dout(w_dff_A_Ff3Shiyc3_0),.din(w_dff_A_8qoe3A5D4_0),.clk(gclk));
	jdff dff_A_aOXGokKK0_0(.dout(w_dff_A_8qoe3A5D4_0),.din(w_dff_A_aOXGokKK0_0),.clk(gclk));
	jdff dff_A_5pXi0zUh1_0(.dout(w_dff_A_aOXGokKK0_0),.din(w_dff_A_5pXi0zUh1_0),.clk(gclk));
	jdff dff_A_Ieuc4sDw6_0(.dout(w_dff_A_5pXi0zUh1_0),.din(w_dff_A_Ieuc4sDw6_0),.clk(gclk));
	jdff dff_A_KJ01cv9u3_0(.dout(w_dff_A_Ieuc4sDw6_0),.din(w_dff_A_KJ01cv9u3_0),.clk(gclk));
	jdff dff_A_L9gT24z83_0(.dout(w_dff_A_KJ01cv9u3_0),.din(w_dff_A_L9gT24z83_0),.clk(gclk));
	jdff dff_A_d3MCYPN24_0(.dout(w_dff_A_L9gT24z83_0),.din(w_dff_A_d3MCYPN24_0),.clk(gclk));
	jdff dff_A_CXCuRGa09_1(.dout(w_n448_0[1]),.din(w_dff_A_CXCuRGa09_1),.clk(gclk));
	jdff dff_B_PtvS5JU96_1(.din(n387),.dout(w_dff_B_PtvS5JU96_1),.clk(gclk));
	jdff dff_B_mbw1FOW70_1(.din(w_dff_B_PtvS5JU96_1),.dout(w_dff_B_mbw1FOW70_1),.clk(gclk));
	jdff dff_B_Nqg9vPeh8_1(.din(w_dff_B_mbw1FOW70_1),.dout(w_dff_B_Nqg9vPeh8_1),.clk(gclk));
	jdff dff_B_0MrTnKSn4_1(.din(w_dff_B_Nqg9vPeh8_1),.dout(w_dff_B_0MrTnKSn4_1),.clk(gclk));
	jdff dff_B_ymdm0y3i6_1(.din(w_dff_B_0MrTnKSn4_1),.dout(w_dff_B_ymdm0y3i6_1),.clk(gclk));
	jdff dff_B_ynY3OOpW1_1(.din(w_dff_B_ymdm0y3i6_1),.dout(w_dff_B_ynY3OOpW1_1),.clk(gclk));
	jdff dff_B_YG9b6rev9_1(.din(w_dff_B_ynY3OOpW1_1),.dout(w_dff_B_YG9b6rev9_1),.clk(gclk));
	jdff dff_B_vsmfJZEW6_1(.din(w_dff_B_YG9b6rev9_1),.dout(w_dff_B_vsmfJZEW6_1),.clk(gclk));
	jdff dff_B_j9sUOswq7_1(.din(w_dff_B_vsmfJZEW6_1),.dout(w_dff_B_j9sUOswq7_1),.clk(gclk));
	jdff dff_B_ACbfjm224_1(.din(w_dff_B_j9sUOswq7_1),.dout(w_dff_B_ACbfjm224_1),.clk(gclk));
	jdff dff_B_Oju7GHiL1_1(.din(w_dff_B_ACbfjm224_1),.dout(w_dff_B_Oju7GHiL1_1),.clk(gclk));
	jdff dff_B_oOKxsGNp6_1(.din(w_dff_B_Oju7GHiL1_1),.dout(w_dff_B_oOKxsGNp6_1),.clk(gclk));
	jdff dff_B_McWBFlO55_1(.din(w_dff_B_oOKxsGNp6_1),.dout(w_dff_B_McWBFlO55_1),.clk(gclk));
	jdff dff_B_CkO3vphw4_1(.din(w_dff_B_McWBFlO55_1),.dout(w_dff_B_CkO3vphw4_1),.clk(gclk));
	jdff dff_B_kvglClJI2_1(.din(w_dff_B_CkO3vphw4_1),.dout(w_dff_B_kvglClJI2_1),.clk(gclk));
	jdff dff_B_xBQ5i8mo0_1(.din(w_dff_B_kvglClJI2_1),.dout(w_dff_B_xBQ5i8mo0_1),.clk(gclk));
	jdff dff_B_90NTLAwQ7_1(.din(w_dff_B_xBQ5i8mo0_1),.dout(w_dff_B_90NTLAwQ7_1),.clk(gclk));
	jdff dff_B_74P4vBwh1_1(.din(w_dff_B_90NTLAwQ7_1),.dout(w_dff_B_74P4vBwh1_1),.clk(gclk));
	jdff dff_B_Pmorb9qW5_1(.din(w_dff_B_74P4vBwh1_1),.dout(w_dff_B_Pmorb9qW5_1),.clk(gclk));
	jdff dff_B_cv4ZrcvC3_1(.din(w_dff_B_Pmorb9qW5_1),.dout(w_dff_B_cv4ZrcvC3_1),.clk(gclk));
	jdff dff_B_PZphXTer8_1(.din(w_dff_B_cv4ZrcvC3_1),.dout(w_dff_B_PZphXTer8_1),.clk(gclk));
	jdff dff_B_kZFmRd181_1(.din(w_dff_B_PZphXTer8_1),.dout(w_dff_B_kZFmRd181_1),.clk(gclk));
	jdff dff_B_YDqN3Te69_1(.din(w_dff_B_kZFmRd181_1),.dout(w_dff_B_YDqN3Te69_1),.clk(gclk));
	jdff dff_B_qslerWkk7_1(.din(w_dff_B_YDqN3Te69_1),.dout(w_dff_B_qslerWkk7_1),.clk(gclk));
	jdff dff_B_ZpA9JmNq8_1(.din(n383),.dout(w_dff_B_ZpA9JmNq8_1),.clk(gclk));
	jdff dff_A_s5OHmhHg5_0(.dout(w_n317_0[0]),.din(w_dff_A_s5OHmhHg5_0),.clk(gclk));
	jdff dff_A_SCFaBpoW3_0(.dout(w_dff_A_s5OHmhHg5_0),.din(w_dff_A_SCFaBpoW3_0),.clk(gclk));
	jdff dff_A_FghTPP2c3_0(.dout(w_dff_A_SCFaBpoW3_0),.din(w_dff_A_FghTPP2c3_0),.clk(gclk));
	jdff dff_A_jbUXCWpC1_0(.dout(w_dff_A_FghTPP2c3_0),.din(w_dff_A_jbUXCWpC1_0),.clk(gclk));
	jdff dff_A_WaOllnxS3_0(.dout(w_dff_A_jbUXCWpC1_0),.din(w_dff_A_WaOllnxS3_0),.clk(gclk));
	jdff dff_A_NmYipz4U3_0(.dout(w_dff_A_WaOllnxS3_0),.din(w_dff_A_NmYipz4U3_0),.clk(gclk));
	jdff dff_A_1QXapqIj6_0(.dout(w_dff_A_NmYipz4U3_0),.din(w_dff_A_1QXapqIj6_0),.clk(gclk));
	jdff dff_A_SvPGsJvD4_0(.dout(w_dff_A_1QXapqIj6_0),.din(w_dff_A_SvPGsJvD4_0),.clk(gclk));
	jdff dff_A_dqDgnsry8_0(.dout(w_dff_A_SvPGsJvD4_0),.din(w_dff_A_dqDgnsry8_0),.clk(gclk));
	jdff dff_A_OOQilvVf2_0(.dout(w_dff_A_dqDgnsry8_0),.din(w_dff_A_OOQilvVf2_0),.clk(gclk));
	jdff dff_A_C59HJymX4_0(.dout(w_dff_A_OOQilvVf2_0),.din(w_dff_A_C59HJymX4_0),.clk(gclk));
	jdff dff_A_WvzSRdQc3_0(.dout(w_dff_A_C59HJymX4_0),.din(w_dff_A_WvzSRdQc3_0),.clk(gclk));
	jdff dff_A_YVfE3w2d2_0(.dout(w_dff_A_WvzSRdQc3_0),.din(w_dff_A_YVfE3w2d2_0),.clk(gclk));
	jdff dff_A_RG13SCtY3_0(.dout(w_dff_A_YVfE3w2d2_0),.din(w_dff_A_RG13SCtY3_0),.clk(gclk));
	jdff dff_A_M4fiS7nu5_0(.dout(w_dff_A_RG13SCtY3_0),.din(w_dff_A_M4fiS7nu5_0),.clk(gclk));
	jdff dff_A_vGy1t0No1_0(.dout(w_dff_A_M4fiS7nu5_0),.din(w_dff_A_vGy1t0No1_0),.clk(gclk));
	jdff dff_A_MSszrTlK3_0(.dout(w_dff_A_vGy1t0No1_0),.din(w_dff_A_MSszrTlK3_0),.clk(gclk));
	jdff dff_A_Xzih0xJN7_0(.dout(w_dff_A_MSszrTlK3_0),.din(w_dff_A_Xzih0xJN7_0),.clk(gclk));
	jdff dff_A_pT8unBlS1_0(.dout(w_dff_A_Xzih0xJN7_0),.din(w_dff_A_pT8unBlS1_0),.clk(gclk));
	jdff dff_A_4hT35RRM9_0(.dout(w_dff_A_pT8unBlS1_0),.din(w_dff_A_4hT35RRM9_0),.clk(gclk));
	jdff dff_A_X20zWPiF9_0(.dout(w_dff_A_4hT35RRM9_0),.din(w_dff_A_X20zWPiF9_0),.clk(gclk));
	jdff dff_A_iOu9PlQg8_0(.dout(w_dff_A_X20zWPiF9_0),.din(w_dff_A_iOu9PlQg8_0),.clk(gclk));
	jdff dff_A_PdF60ZML1_0(.dout(w_dff_A_iOu9PlQg8_0),.din(w_dff_A_PdF60ZML1_0),.clk(gclk));
	jdff dff_A_Hgv2ssJz7_0(.dout(w_dff_A_PdF60ZML1_0),.din(w_dff_A_Hgv2ssJz7_0),.clk(gclk));
	jdff dff_A_bZ4o1eNL3_0(.dout(w_dff_A_Hgv2ssJz7_0),.din(w_dff_A_bZ4o1eNL3_0),.clk(gclk));
	jdff dff_A_UNh2eDPN7_1(.dout(w_n377_0[1]),.din(w_dff_A_UNh2eDPN7_1),.clk(gclk));
	jdff dff_B_446mc0tf3_1(.din(n324),.dout(w_dff_B_446mc0tf3_1),.clk(gclk));
	jdff dff_B_beI0umwh0_1(.din(w_dff_B_446mc0tf3_1),.dout(w_dff_B_beI0umwh0_1),.clk(gclk));
	jdff dff_B_diEnk7oY4_1(.din(w_dff_B_beI0umwh0_1),.dout(w_dff_B_diEnk7oY4_1),.clk(gclk));
	jdff dff_B_6b2SGBvD7_1(.din(w_dff_B_diEnk7oY4_1),.dout(w_dff_B_6b2SGBvD7_1),.clk(gclk));
	jdff dff_B_yMtqXUPN9_1(.din(w_dff_B_6b2SGBvD7_1),.dout(w_dff_B_yMtqXUPN9_1),.clk(gclk));
	jdff dff_B_MtD0yVFQ5_1(.din(w_dff_B_yMtqXUPN9_1),.dout(w_dff_B_MtD0yVFQ5_1),.clk(gclk));
	jdff dff_B_DjsAcU4Y7_1(.din(w_dff_B_MtD0yVFQ5_1),.dout(w_dff_B_DjsAcU4Y7_1),.clk(gclk));
	jdff dff_B_GbhPqi6W5_1(.din(w_dff_B_DjsAcU4Y7_1),.dout(w_dff_B_GbhPqi6W5_1),.clk(gclk));
	jdff dff_B_Eee7ff629_1(.din(w_dff_B_GbhPqi6W5_1),.dout(w_dff_B_Eee7ff629_1),.clk(gclk));
	jdff dff_B_mTMfebD38_1(.din(w_dff_B_Eee7ff629_1),.dout(w_dff_B_mTMfebD38_1),.clk(gclk));
	jdff dff_B_czrf5Jbs5_1(.din(w_dff_B_mTMfebD38_1),.dout(w_dff_B_czrf5Jbs5_1),.clk(gclk));
	jdff dff_B_6xEokzLD9_1(.din(w_dff_B_czrf5Jbs5_1),.dout(w_dff_B_6xEokzLD9_1),.clk(gclk));
	jdff dff_B_cZZmQE5Q3_1(.din(w_dff_B_6xEokzLD9_1),.dout(w_dff_B_cZZmQE5Q3_1),.clk(gclk));
	jdff dff_B_HUTuF5Xa7_1(.din(w_dff_B_cZZmQE5Q3_1),.dout(w_dff_B_HUTuF5Xa7_1),.clk(gclk));
	jdff dff_B_WAakYAi93_1(.din(w_dff_B_HUTuF5Xa7_1),.dout(w_dff_B_WAakYAi93_1),.clk(gclk));
	jdff dff_B_Snh2BeM71_1(.din(w_dff_B_WAakYAi93_1),.dout(w_dff_B_Snh2BeM71_1),.clk(gclk));
	jdff dff_B_jQrVFQ9k5_1(.din(w_dff_B_Snh2BeM71_1),.dout(w_dff_B_jQrVFQ9k5_1),.clk(gclk));
	jdff dff_B_pjUBAyGf4_1(.din(w_dff_B_jQrVFQ9k5_1),.dout(w_dff_B_pjUBAyGf4_1),.clk(gclk));
	jdff dff_B_QwwPHf2d4_1(.din(w_dff_B_pjUBAyGf4_1),.dout(w_dff_B_QwwPHf2d4_1),.clk(gclk));
	jdff dff_B_WkPDkMw68_1(.din(w_dff_B_QwwPHf2d4_1),.dout(w_dff_B_WkPDkMw68_1),.clk(gclk));
	jdff dff_B_tbVrxYkZ0_1(.din(w_dff_B_WkPDkMw68_1),.dout(w_dff_B_tbVrxYkZ0_1),.clk(gclk));
	jdff dff_B_3wO4YlSX2_1(.din(n320),.dout(w_dff_B_3wO4YlSX2_1),.clk(gclk));
	jdff dff_A_4CNz0Ejq0_0(.dout(w_n261_0[0]),.din(w_dff_A_4CNz0Ejq0_0),.clk(gclk));
	jdff dff_A_obpJO30q9_0(.dout(w_dff_A_4CNz0Ejq0_0),.din(w_dff_A_obpJO30q9_0),.clk(gclk));
	jdff dff_A_dZNstbAX2_0(.dout(w_dff_A_obpJO30q9_0),.din(w_dff_A_dZNstbAX2_0),.clk(gclk));
	jdff dff_A_YkU4HKhe2_0(.dout(w_dff_A_dZNstbAX2_0),.din(w_dff_A_YkU4HKhe2_0),.clk(gclk));
	jdff dff_A_ZOYfEGjf3_0(.dout(w_dff_A_YkU4HKhe2_0),.din(w_dff_A_ZOYfEGjf3_0),.clk(gclk));
	jdff dff_A_j1eut0b90_0(.dout(w_dff_A_ZOYfEGjf3_0),.din(w_dff_A_j1eut0b90_0),.clk(gclk));
	jdff dff_A_lHk6dL8F3_0(.dout(w_dff_A_j1eut0b90_0),.din(w_dff_A_lHk6dL8F3_0),.clk(gclk));
	jdff dff_A_Ad7PnX578_0(.dout(w_dff_A_lHk6dL8F3_0),.din(w_dff_A_Ad7PnX578_0),.clk(gclk));
	jdff dff_A_bNdnQQHs9_0(.dout(w_dff_A_Ad7PnX578_0),.din(w_dff_A_bNdnQQHs9_0),.clk(gclk));
	jdff dff_A_E7ZxRcSB1_0(.dout(w_dff_A_bNdnQQHs9_0),.din(w_dff_A_E7ZxRcSB1_0),.clk(gclk));
	jdff dff_A_u10TAW412_0(.dout(w_dff_A_E7ZxRcSB1_0),.din(w_dff_A_u10TAW412_0),.clk(gclk));
	jdff dff_A_XCyAKAhL4_0(.dout(w_dff_A_u10TAW412_0),.din(w_dff_A_XCyAKAhL4_0),.clk(gclk));
	jdff dff_A_ALQuVkGo2_0(.dout(w_dff_A_XCyAKAhL4_0),.din(w_dff_A_ALQuVkGo2_0),.clk(gclk));
	jdff dff_A_4CWDRDKO7_0(.dout(w_dff_A_ALQuVkGo2_0),.din(w_dff_A_4CWDRDKO7_0),.clk(gclk));
	jdff dff_A_XLKzj4l83_0(.dout(w_dff_A_4CWDRDKO7_0),.din(w_dff_A_XLKzj4l83_0),.clk(gclk));
	jdff dff_A_bPCdQkeh4_0(.dout(w_dff_A_XLKzj4l83_0),.din(w_dff_A_bPCdQkeh4_0),.clk(gclk));
	jdff dff_A_LsuONHZD2_0(.dout(w_dff_A_bPCdQkeh4_0),.din(w_dff_A_LsuONHZD2_0),.clk(gclk));
	jdff dff_A_MN3hfL696_0(.dout(w_dff_A_LsuONHZD2_0),.din(w_dff_A_MN3hfL696_0),.clk(gclk));
	jdff dff_A_vvbD3iRi9_0(.dout(w_dff_A_MN3hfL696_0),.din(w_dff_A_vvbD3iRi9_0),.clk(gclk));
	jdff dff_A_miFEZiZL9_0(.dout(w_dff_A_vvbD3iRi9_0),.din(w_dff_A_miFEZiZL9_0),.clk(gclk));
	jdff dff_A_3vAgnj9q3_0(.dout(w_dff_A_miFEZiZL9_0),.din(w_dff_A_3vAgnj9q3_0),.clk(gclk));
	jdff dff_A_xFr8Ne6S7_0(.dout(w_dff_A_3vAgnj9q3_0),.din(w_dff_A_xFr8Ne6S7_0),.clk(gclk));
	jdff dff_A_iki1Wsv18_1(.dout(w_n314_0[1]),.din(w_dff_A_iki1Wsv18_1),.clk(gclk));
	jdff dff_B_oV4xYXZt9_1(.din(n268),.dout(w_dff_B_oV4xYXZt9_1),.clk(gclk));
	jdff dff_B_dvri7vgW5_1(.din(w_dff_B_oV4xYXZt9_1),.dout(w_dff_B_dvri7vgW5_1),.clk(gclk));
	jdff dff_B_W5EZtmxx4_1(.din(w_dff_B_dvri7vgW5_1),.dout(w_dff_B_W5EZtmxx4_1),.clk(gclk));
	jdff dff_B_CZsJfKZq6_1(.din(w_dff_B_W5EZtmxx4_1),.dout(w_dff_B_CZsJfKZq6_1),.clk(gclk));
	jdff dff_B_pnDOXqfT8_1(.din(w_dff_B_CZsJfKZq6_1),.dout(w_dff_B_pnDOXqfT8_1),.clk(gclk));
	jdff dff_B_aLpKKp8R1_1(.din(w_dff_B_pnDOXqfT8_1),.dout(w_dff_B_aLpKKp8R1_1),.clk(gclk));
	jdff dff_B_8RYHX3332_1(.din(w_dff_B_aLpKKp8R1_1),.dout(w_dff_B_8RYHX3332_1),.clk(gclk));
	jdff dff_B_p1Jo63Pu7_1(.din(w_dff_B_8RYHX3332_1),.dout(w_dff_B_p1Jo63Pu7_1),.clk(gclk));
	jdff dff_B_6ykyMfno0_1(.din(w_dff_B_p1Jo63Pu7_1),.dout(w_dff_B_6ykyMfno0_1),.clk(gclk));
	jdff dff_B_Zl2tUOaP3_1(.din(w_dff_B_6ykyMfno0_1),.dout(w_dff_B_Zl2tUOaP3_1),.clk(gclk));
	jdff dff_B_GtgmVF3a7_1(.din(w_dff_B_Zl2tUOaP3_1),.dout(w_dff_B_GtgmVF3a7_1),.clk(gclk));
	jdff dff_B_3mMvkFAu6_1(.din(w_dff_B_GtgmVF3a7_1),.dout(w_dff_B_3mMvkFAu6_1),.clk(gclk));
	jdff dff_B_QT86LUp77_1(.din(w_dff_B_3mMvkFAu6_1),.dout(w_dff_B_QT86LUp77_1),.clk(gclk));
	jdff dff_B_cnpNgyWw9_1(.din(w_dff_B_QT86LUp77_1),.dout(w_dff_B_cnpNgyWw9_1),.clk(gclk));
	jdff dff_B_2RZeftVy2_1(.din(w_dff_B_cnpNgyWw9_1),.dout(w_dff_B_2RZeftVy2_1),.clk(gclk));
	jdff dff_B_IM95GAQg2_1(.din(w_dff_B_2RZeftVy2_1),.dout(w_dff_B_IM95GAQg2_1),.clk(gclk));
	jdff dff_B_r1CnYXuj2_1(.din(w_dff_B_IM95GAQg2_1),.dout(w_dff_B_r1CnYXuj2_1),.clk(gclk));
	jdff dff_B_mPvqQbQg9_1(.din(w_dff_B_r1CnYXuj2_1),.dout(w_dff_B_mPvqQbQg9_1),.clk(gclk));
	jdff dff_B_cjBnXVB24_1(.din(n264),.dout(w_dff_B_cjBnXVB24_1),.clk(gclk));
	jdff dff_A_96bRC0UK7_0(.dout(w_n212_0[0]),.din(w_dff_A_96bRC0UK7_0),.clk(gclk));
	jdff dff_A_kZEQKxM98_0(.dout(w_dff_A_96bRC0UK7_0),.din(w_dff_A_kZEQKxM98_0),.clk(gclk));
	jdff dff_A_sWdKdqXm3_0(.dout(w_dff_A_kZEQKxM98_0),.din(w_dff_A_sWdKdqXm3_0),.clk(gclk));
	jdff dff_A_pCJ7f2W59_0(.dout(w_dff_A_sWdKdqXm3_0),.din(w_dff_A_pCJ7f2W59_0),.clk(gclk));
	jdff dff_A_PrBPUt7H2_0(.dout(w_dff_A_pCJ7f2W59_0),.din(w_dff_A_PrBPUt7H2_0),.clk(gclk));
	jdff dff_A_MGBfStTH7_0(.dout(w_dff_A_PrBPUt7H2_0),.din(w_dff_A_MGBfStTH7_0),.clk(gclk));
	jdff dff_A_2n2Apw1D5_0(.dout(w_dff_A_MGBfStTH7_0),.din(w_dff_A_2n2Apw1D5_0),.clk(gclk));
	jdff dff_A_8CJh9Ckb5_0(.dout(w_dff_A_2n2Apw1D5_0),.din(w_dff_A_8CJh9Ckb5_0),.clk(gclk));
	jdff dff_A_RIAETzaY3_0(.dout(w_dff_A_8CJh9Ckb5_0),.din(w_dff_A_RIAETzaY3_0),.clk(gclk));
	jdff dff_A_543fqMmN2_0(.dout(w_dff_A_RIAETzaY3_0),.din(w_dff_A_543fqMmN2_0),.clk(gclk));
	jdff dff_A_vK5bv9kC6_0(.dout(w_dff_A_543fqMmN2_0),.din(w_dff_A_vK5bv9kC6_0),.clk(gclk));
	jdff dff_A_CFUJTBnW1_0(.dout(w_dff_A_vK5bv9kC6_0),.din(w_dff_A_CFUJTBnW1_0),.clk(gclk));
	jdff dff_A_sErRkcCl4_0(.dout(w_dff_A_CFUJTBnW1_0),.din(w_dff_A_sErRkcCl4_0),.clk(gclk));
	jdff dff_A_j6nAlm6e6_0(.dout(w_dff_A_sErRkcCl4_0),.din(w_dff_A_j6nAlm6e6_0),.clk(gclk));
	jdff dff_A_57y9QFPw7_0(.dout(w_dff_A_j6nAlm6e6_0),.din(w_dff_A_57y9QFPw7_0),.clk(gclk));
	jdff dff_A_3feiKSxl8_0(.dout(w_dff_A_57y9QFPw7_0),.din(w_dff_A_3feiKSxl8_0),.clk(gclk));
	jdff dff_A_w8zJmMbx2_0(.dout(w_dff_A_3feiKSxl8_0),.din(w_dff_A_w8zJmMbx2_0),.clk(gclk));
	jdff dff_A_MbeXN5xh0_0(.dout(w_dff_A_w8zJmMbx2_0),.din(w_dff_A_MbeXN5xh0_0),.clk(gclk));
	jdff dff_A_hTpwivnN8_0(.dout(w_dff_A_MbeXN5xh0_0),.din(w_dff_A_hTpwivnN8_0),.clk(gclk));
	jdff dff_A_T4cDbbGE9_1(.dout(w_n258_0[1]),.din(w_dff_A_T4cDbbGE9_1),.clk(gclk));
	jdff dff_B_9KhjrN6S2_1(.din(n219),.dout(w_dff_B_9KhjrN6S2_1),.clk(gclk));
	jdff dff_B_QAm33Y5Q5_1(.din(w_dff_B_9KhjrN6S2_1),.dout(w_dff_B_QAm33Y5Q5_1),.clk(gclk));
	jdff dff_B_r1jZANC11_1(.din(w_dff_B_QAm33Y5Q5_1),.dout(w_dff_B_r1jZANC11_1),.clk(gclk));
	jdff dff_B_pCJkc8a62_1(.din(w_dff_B_r1jZANC11_1),.dout(w_dff_B_pCJkc8a62_1),.clk(gclk));
	jdff dff_B_hLFgJVMM0_1(.din(w_dff_B_pCJkc8a62_1),.dout(w_dff_B_hLFgJVMM0_1),.clk(gclk));
	jdff dff_B_KvRu4fax7_1(.din(w_dff_B_hLFgJVMM0_1),.dout(w_dff_B_KvRu4fax7_1),.clk(gclk));
	jdff dff_B_RT4vUHdy6_1(.din(w_dff_B_KvRu4fax7_1),.dout(w_dff_B_RT4vUHdy6_1),.clk(gclk));
	jdff dff_B_R2DSn46J8_1(.din(w_dff_B_RT4vUHdy6_1),.dout(w_dff_B_R2DSn46J8_1),.clk(gclk));
	jdff dff_B_SL2Sb3oK8_1(.din(w_dff_B_R2DSn46J8_1),.dout(w_dff_B_SL2Sb3oK8_1),.clk(gclk));
	jdff dff_B_LbnUKm7O3_1(.din(w_dff_B_SL2Sb3oK8_1),.dout(w_dff_B_LbnUKm7O3_1),.clk(gclk));
	jdff dff_B_ltJw6WsM4_1(.din(w_dff_B_LbnUKm7O3_1),.dout(w_dff_B_ltJw6WsM4_1),.clk(gclk));
	jdff dff_B_Nv1OoUv25_1(.din(w_dff_B_ltJw6WsM4_1),.dout(w_dff_B_Nv1OoUv25_1),.clk(gclk));
	jdff dff_B_cjOZ3a0d7_1(.din(w_dff_B_Nv1OoUv25_1),.dout(w_dff_B_cjOZ3a0d7_1),.clk(gclk));
	jdff dff_B_2i1rmVbG7_1(.din(w_dff_B_cjOZ3a0d7_1),.dout(w_dff_B_2i1rmVbG7_1),.clk(gclk));
	jdff dff_B_e1S54b0o3_1(.din(w_dff_B_2i1rmVbG7_1),.dout(w_dff_B_e1S54b0o3_1),.clk(gclk));
	jdff dff_B_ARqMBHW71_1(.din(n215),.dout(w_dff_B_ARqMBHW71_1),.clk(gclk));
	jdff dff_A_jN1yvcrQ3_0(.dout(w_n170_0[0]),.din(w_dff_A_jN1yvcrQ3_0),.clk(gclk));
	jdff dff_A_RaUhwoHn2_0(.dout(w_dff_A_jN1yvcrQ3_0),.din(w_dff_A_RaUhwoHn2_0),.clk(gclk));
	jdff dff_A_HjnLsjbO2_0(.dout(w_dff_A_RaUhwoHn2_0),.din(w_dff_A_HjnLsjbO2_0),.clk(gclk));
	jdff dff_A_ToH3PObi3_0(.dout(w_dff_A_HjnLsjbO2_0),.din(w_dff_A_ToH3PObi3_0),.clk(gclk));
	jdff dff_A_Oghdby3S3_0(.dout(w_dff_A_ToH3PObi3_0),.din(w_dff_A_Oghdby3S3_0),.clk(gclk));
	jdff dff_A_G8nSVk0x4_0(.dout(w_dff_A_Oghdby3S3_0),.din(w_dff_A_G8nSVk0x4_0),.clk(gclk));
	jdff dff_A_YAxoQRoe4_0(.dout(w_dff_A_G8nSVk0x4_0),.din(w_dff_A_YAxoQRoe4_0),.clk(gclk));
	jdff dff_A_S6NMjrMg7_0(.dout(w_dff_A_YAxoQRoe4_0),.din(w_dff_A_S6NMjrMg7_0),.clk(gclk));
	jdff dff_A_WajgXwx04_0(.dout(w_dff_A_S6NMjrMg7_0),.din(w_dff_A_WajgXwx04_0),.clk(gclk));
	jdff dff_A_T6yBKPDw4_0(.dout(w_dff_A_WajgXwx04_0),.din(w_dff_A_T6yBKPDw4_0),.clk(gclk));
	jdff dff_A_kNDyUytj8_0(.dout(w_dff_A_T6yBKPDw4_0),.din(w_dff_A_kNDyUytj8_0),.clk(gclk));
	jdff dff_A_LVPkdWoh0_0(.dout(w_dff_A_kNDyUytj8_0),.din(w_dff_A_LVPkdWoh0_0),.clk(gclk));
	jdff dff_A_CICRyl5C9_0(.dout(w_dff_A_LVPkdWoh0_0),.din(w_dff_A_CICRyl5C9_0),.clk(gclk));
	jdff dff_A_Hy7KfI5w8_0(.dout(w_dff_A_CICRyl5C9_0),.din(w_dff_A_Hy7KfI5w8_0),.clk(gclk));
	jdff dff_A_HRTrxZWu9_0(.dout(w_dff_A_Hy7KfI5w8_0),.din(w_dff_A_HRTrxZWu9_0),.clk(gclk));
	jdff dff_A_qGBbdJg55_0(.dout(w_dff_A_HRTrxZWu9_0),.din(w_dff_A_qGBbdJg55_0),.clk(gclk));
	jdff dff_A_uD5kYzFY7_1(.dout(w_n209_0[1]),.din(w_dff_A_uD5kYzFY7_1),.clk(gclk));
	jdff dff_B_19xdoAS41_1(.din(n177),.dout(w_dff_B_19xdoAS41_1),.clk(gclk));
	jdff dff_B_0SFShaYm4_1(.din(w_dff_B_19xdoAS41_1),.dout(w_dff_B_0SFShaYm4_1),.clk(gclk));
	jdff dff_B_cyx4Fo573_1(.din(w_dff_B_0SFShaYm4_1),.dout(w_dff_B_cyx4Fo573_1),.clk(gclk));
	jdff dff_B_Af8IFqgp2_1(.din(w_dff_B_cyx4Fo573_1),.dout(w_dff_B_Af8IFqgp2_1),.clk(gclk));
	jdff dff_B_7rXxdFcr8_1(.din(w_dff_B_Af8IFqgp2_1),.dout(w_dff_B_7rXxdFcr8_1),.clk(gclk));
	jdff dff_B_flES295I5_1(.din(w_dff_B_7rXxdFcr8_1),.dout(w_dff_B_flES295I5_1),.clk(gclk));
	jdff dff_B_eMCIV4kl0_1(.din(w_dff_B_flES295I5_1),.dout(w_dff_B_eMCIV4kl0_1),.clk(gclk));
	jdff dff_B_HoYeT0Dg5_1(.din(w_dff_B_eMCIV4kl0_1),.dout(w_dff_B_HoYeT0Dg5_1),.clk(gclk));
	jdff dff_B_E5Seo1lz6_1(.din(w_dff_B_HoYeT0Dg5_1),.dout(w_dff_B_E5Seo1lz6_1),.clk(gclk));
	jdff dff_B_VevoZam20_1(.din(w_dff_B_E5Seo1lz6_1),.dout(w_dff_B_VevoZam20_1),.clk(gclk));
	jdff dff_B_T019ONPG9_1(.din(w_dff_B_VevoZam20_1),.dout(w_dff_B_T019ONPG9_1),.clk(gclk));
	jdff dff_B_OMTgwC4u0_1(.din(w_dff_B_T019ONPG9_1),.dout(w_dff_B_OMTgwC4u0_1),.clk(gclk));
	jdff dff_B_Sr0tDaY84_1(.din(n173),.dout(w_dff_B_Sr0tDaY84_1),.clk(gclk));
	jdff dff_A_Y8MDE0nn7_0(.dout(w_n135_0[0]),.din(w_dff_A_Y8MDE0nn7_0),.clk(gclk));
	jdff dff_A_y5Wih8TQ2_0(.dout(w_dff_A_Y8MDE0nn7_0),.din(w_dff_A_y5Wih8TQ2_0),.clk(gclk));
	jdff dff_A_R3EBK8zM4_0(.dout(w_dff_A_y5Wih8TQ2_0),.din(w_dff_A_R3EBK8zM4_0),.clk(gclk));
	jdff dff_A_TKCT3uPW7_0(.dout(w_dff_A_R3EBK8zM4_0),.din(w_dff_A_TKCT3uPW7_0),.clk(gclk));
	jdff dff_A_AYHCPS5a0_0(.dout(w_dff_A_TKCT3uPW7_0),.din(w_dff_A_AYHCPS5a0_0),.clk(gclk));
	jdff dff_A_BW5oXrDJ0_0(.dout(w_dff_A_AYHCPS5a0_0),.din(w_dff_A_BW5oXrDJ0_0),.clk(gclk));
	jdff dff_A_B2tNOhAu4_0(.dout(w_dff_A_BW5oXrDJ0_0),.din(w_dff_A_B2tNOhAu4_0),.clk(gclk));
	jdff dff_A_GWCOKTZh8_0(.dout(w_dff_A_B2tNOhAu4_0),.din(w_dff_A_GWCOKTZh8_0),.clk(gclk));
	jdff dff_A_xYE3SDwP0_0(.dout(w_dff_A_GWCOKTZh8_0),.din(w_dff_A_xYE3SDwP0_0),.clk(gclk));
	jdff dff_A_7xIgJLIw6_0(.dout(w_dff_A_xYE3SDwP0_0),.din(w_dff_A_7xIgJLIw6_0),.clk(gclk));
	jdff dff_A_hzBWj4kg0_0(.dout(w_dff_A_7xIgJLIw6_0),.din(w_dff_A_hzBWj4kg0_0),.clk(gclk));
	jdff dff_A_2dQSuDDW1_0(.dout(w_dff_A_hzBWj4kg0_0),.din(w_dff_A_2dQSuDDW1_0),.clk(gclk));
	jdff dff_A_Kob3NXpf4_0(.dout(w_dff_A_2dQSuDDW1_0),.din(w_dff_A_Kob3NXpf4_0),.clk(gclk));
	jdff dff_A_MTOSucTE3_1(.dout(w_n167_0[1]),.din(w_dff_A_MTOSucTE3_1),.clk(gclk));
	jdff dff_B_TNm26uXl7_1(.din(n142),.dout(w_dff_B_TNm26uXl7_1),.clk(gclk));
	jdff dff_B_vJUMpkoL3_1(.din(w_dff_B_TNm26uXl7_1),.dout(w_dff_B_vJUMpkoL3_1),.clk(gclk));
	jdff dff_B_sZFoQiwo9_1(.din(w_dff_B_vJUMpkoL3_1),.dout(w_dff_B_sZFoQiwo9_1),.clk(gclk));
	jdff dff_B_hfrFw3Gl5_1(.din(w_dff_B_sZFoQiwo9_1),.dout(w_dff_B_hfrFw3Gl5_1),.clk(gclk));
	jdff dff_B_FxCMNQb69_1(.din(w_dff_B_hfrFw3Gl5_1),.dout(w_dff_B_FxCMNQb69_1),.clk(gclk));
	jdff dff_B_moLoIsf50_1(.din(w_dff_B_FxCMNQb69_1),.dout(w_dff_B_moLoIsf50_1),.clk(gclk));
	jdff dff_B_o2XwuzLU6_1(.din(w_dff_B_moLoIsf50_1),.dout(w_dff_B_o2XwuzLU6_1),.clk(gclk));
	jdff dff_B_8sbivfWl9_1(.din(w_dff_B_o2XwuzLU6_1),.dout(w_dff_B_8sbivfWl9_1),.clk(gclk));
	jdff dff_B_UaMuF6AQ2_1(.din(w_dff_B_8sbivfWl9_1),.dout(w_dff_B_UaMuF6AQ2_1),.clk(gclk));
	jdff dff_B_UhHJoqrF3_1(.din(n138),.dout(w_dff_B_UhHJoqrF3_1),.clk(gclk));
	jdff dff_A_G8vsu7JU5_0(.dout(w_n106_0[0]),.din(w_dff_A_G8vsu7JU5_0),.clk(gclk));
	jdff dff_A_UfYd6nfG4_0(.dout(w_dff_A_G8vsu7JU5_0),.din(w_dff_A_UfYd6nfG4_0),.clk(gclk));
	jdff dff_A_JLIULioC0_0(.dout(w_dff_A_UfYd6nfG4_0),.din(w_dff_A_JLIULioC0_0),.clk(gclk));
	jdff dff_A_95S42CIv1_0(.dout(w_dff_A_JLIULioC0_0),.din(w_dff_A_95S42CIv1_0),.clk(gclk));
	jdff dff_A_xJWFmSS82_0(.dout(w_dff_A_95S42CIv1_0),.din(w_dff_A_xJWFmSS82_0),.clk(gclk));
	jdff dff_A_mI1FmnB74_0(.dout(w_dff_A_xJWFmSS82_0),.din(w_dff_A_mI1FmnB74_0),.clk(gclk));
	jdff dff_A_6yzDuOo62_0(.dout(w_dff_A_mI1FmnB74_0),.din(w_dff_A_6yzDuOo62_0),.clk(gclk));
	jdff dff_A_WeLQMx1r3_0(.dout(w_dff_A_6yzDuOo62_0),.din(w_dff_A_WeLQMx1r3_0),.clk(gclk));
	jdff dff_A_V7osYO1T2_0(.dout(w_dff_A_WeLQMx1r3_0),.din(w_dff_A_V7osYO1T2_0),.clk(gclk));
	jdff dff_A_qKRfbRCj6_0(.dout(w_dff_A_V7osYO1T2_0),.din(w_dff_A_qKRfbRCj6_0),.clk(gclk));
	jdff dff_A_Hwo7FDkD5_1(.dout(w_n132_0[1]),.din(w_dff_A_Hwo7FDkD5_1),.clk(gclk));
	jdff dff_B_PjyqkwbN1_1(.din(n113),.dout(w_dff_B_PjyqkwbN1_1),.clk(gclk));
	jdff dff_B_lpuBoLUN7_1(.din(w_dff_B_PjyqkwbN1_1),.dout(w_dff_B_lpuBoLUN7_1),.clk(gclk));
	jdff dff_B_MFL0n9fK3_1(.din(w_dff_B_lpuBoLUN7_1),.dout(w_dff_B_MFL0n9fK3_1),.clk(gclk));
	jdff dff_B_gENoNltn3_1(.din(w_dff_B_MFL0n9fK3_1),.dout(w_dff_B_gENoNltn3_1),.clk(gclk));
	jdff dff_B_Z4EjBICu4_1(.din(w_dff_B_gENoNltn3_1),.dout(w_dff_B_Z4EjBICu4_1),.clk(gclk));
	jdff dff_B_VfglReMp4_1(.din(w_dff_B_Z4EjBICu4_1),.dout(w_dff_B_VfglReMp4_1),.clk(gclk));
	jdff dff_B_LscLupag7_1(.din(n109),.dout(w_dff_B_LscLupag7_1),.clk(gclk));
	jdff dff_A_NR91Qro00_0(.dout(w_n86_0[0]),.din(w_dff_A_NR91Qro00_0),.clk(gclk));
	jdff dff_A_tlL3Ex4Y2_0(.dout(w_dff_A_NR91Qro00_0),.din(w_dff_A_tlL3Ex4Y2_0),.clk(gclk));
	jdff dff_A_avBnkoxX8_0(.dout(w_dff_A_tlL3Ex4Y2_0),.din(w_dff_A_avBnkoxX8_0),.clk(gclk));
	jdff dff_A_JVsq5GdX6_0(.dout(w_dff_A_avBnkoxX8_0),.din(w_dff_A_JVsq5GdX6_0),.clk(gclk));
	jdff dff_A_hEoXENyr3_0(.dout(w_dff_A_JVsq5GdX6_0),.din(w_dff_A_hEoXENyr3_0),.clk(gclk));
	jdff dff_A_6guS20r26_0(.dout(w_dff_A_hEoXENyr3_0),.din(w_dff_A_6guS20r26_0),.clk(gclk));
	jdff dff_A_zLcH8Jq08_0(.dout(w_dff_A_6guS20r26_0),.din(w_dff_A_zLcH8Jq08_0),.clk(gclk));
	jdff dff_A_DRCi3GWz7_1(.dout(w_n103_0[1]),.din(w_dff_A_DRCi3GWz7_1),.clk(gclk));
	jdff dff_B_XKBdWjFg5_1(.din(n92),.dout(w_dff_B_XKBdWjFg5_1),.clk(gclk));
	jdff dff_B_8WETelJ59_1(.din(w_dff_B_XKBdWjFg5_1),.dout(w_dff_B_8WETelJ59_1),.clk(gclk));
	jdff dff_B_x4Y6O9rC9_1(.din(w_dff_B_8WETelJ59_1),.dout(w_dff_B_x4Y6O9rC9_1),.clk(gclk));
	jdff dff_B_QQCVQAKW5_1(.din(n88),.dout(w_dff_B_QQCVQAKW5_1),.clk(gclk));
	jdff dff_B_2dDyRXUu5_2(.din(n67),.dout(w_dff_B_2dDyRXUu5_2),.clk(gclk));
	jdff dff_A_KKIkw2iX1_0(.dout(w_n75_0[0]),.din(w_dff_A_KKIkw2iX1_0),.clk(gclk));
	jdff dff_A_JvxhZenG3_0(.dout(w_dff_A_KKIkw2iX1_0),.din(w_dff_A_JvxhZenG3_0),.clk(gclk));
	jdff dff_A_fDnV6WPg1_0(.dout(w_dff_A_JvxhZenG3_0),.din(w_dff_A_fDnV6WPg1_0),.clk(gclk));
	jdff dff_A_fEHBPXtO2_0(.dout(w_dff_A_fDnV6WPg1_0),.din(w_dff_A_fEHBPXtO2_0),.clk(gclk));
	jdff dff_B_rhRcGDUD6_0(.din(n82),.dout(w_dff_B_rhRcGDUD6_0),.clk(gclk));
	jdff dff_A_TQJWSXqW0_0(.dout(w_n66_0[0]),.din(w_dff_A_TQJWSXqW0_0),.clk(gclk));
	jdff dff_A_UFSzZaHP3_0(.dout(w_dff_A_TQJWSXqW0_0),.din(w_dff_A_UFSzZaHP3_0),.clk(gclk));
	jdff dff_A_yNR5ZAP00_1(.dout(w_n1108_0[1]),.din(w_dff_A_yNR5ZAP00_1),.clk(gclk));
	jdff dff_B_Hl1lC4wT5_1(.din(n1014),.dout(w_dff_B_Hl1lC4wT5_1),.clk(gclk));
	jdff dff_B_rZ8s8lDN4_2(.din(n911),.dout(w_dff_B_rZ8s8lDN4_2),.clk(gclk));
	jdff dff_B_yp2wwtls7_2(.din(w_dff_B_rZ8s8lDN4_2),.dout(w_dff_B_yp2wwtls7_2),.clk(gclk));
	jdff dff_B_aM434uSq7_2(.din(w_dff_B_yp2wwtls7_2),.dout(w_dff_B_aM434uSq7_2),.clk(gclk));
	jdff dff_B_ChjqsWof0_2(.din(w_dff_B_aM434uSq7_2),.dout(w_dff_B_ChjqsWof0_2),.clk(gclk));
	jdff dff_B_bJtuTtBf9_2(.din(w_dff_B_ChjqsWof0_2),.dout(w_dff_B_bJtuTtBf9_2),.clk(gclk));
	jdff dff_B_9iUe1dal3_2(.din(w_dff_B_bJtuTtBf9_2),.dout(w_dff_B_9iUe1dal3_2),.clk(gclk));
	jdff dff_B_6Zp8lnp06_2(.din(w_dff_B_9iUe1dal3_2),.dout(w_dff_B_6Zp8lnp06_2),.clk(gclk));
	jdff dff_B_CcrfbxCA1_2(.din(w_dff_B_6Zp8lnp06_2),.dout(w_dff_B_CcrfbxCA1_2),.clk(gclk));
	jdff dff_B_CSjfPYqI3_2(.din(w_dff_B_CcrfbxCA1_2),.dout(w_dff_B_CSjfPYqI3_2),.clk(gclk));
	jdff dff_B_vhrUB80L6_2(.din(w_dff_B_CSjfPYqI3_2),.dout(w_dff_B_vhrUB80L6_2),.clk(gclk));
	jdff dff_B_7ZEVWyUE1_2(.din(w_dff_B_vhrUB80L6_2),.dout(w_dff_B_7ZEVWyUE1_2),.clk(gclk));
	jdff dff_B_iegYqkeL6_2(.din(w_dff_B_7ZEVWyUE1_2),.dout(w_dff_B_iegYqkeL6_2),.clk(gclk));
	jdff dff_B_jhQiMmtV6_2(.din(w_dff_B_iegYqkeL6_2),.dout(w_dff_B_jhQiMmtV6_2),.clk(gclk));
	jdff dff_B_hs2IXzDu9_2(.din(w_dff_B_jhQiMmtV6_2),.dout(w_dff_B_hs2IXzDu9_2),.clk(gclk));
	jdff dff_B_h8C3J6dQ2_2(.din(w_dff_B_hs2IXzDu9_2),.dout(w_dff_B_h8C3J6dQ2_2),.clk(gclk));
	jdff dff_B_Yj1TTTok5_2(.din(w_dff_B_h8C3J6dQ2_2),.dout(w_dff_B_Yj1TTTok5_2),.clk(gclk));
	jdff dff_B_M4YbZoyE5_2(.din(w_dff_B_Yj1TTTok5_2),.dout(w_dff_B_M4YbZoyE5_2),.clk(gclk));
	jdff dff_B_9qkKWTqq3_2(.din(w_dff_B_M4YbZoyE5_2),.dout(w_dff_B_9qkKWTqq3_2),.clk(gclk));
	jdff dff_B_TUjygvcK5_2(.din(w_dff_B_9qkKWTqq3_2),.dout(w_dff_B_TUjygvcK5_2),.clk(gclk));
	jdff dff_B_g6sxgFEa2_2(.din(w_dff_B_TUjygvcK5_2),.dout(w_dff_B_g6sxgFEa2_2),.clk(gclk));
	jdff dff_B_5o3Niwzm4_2(.din(w_dff_B_g6sxgFEa2_2),.dout(w_dff_B_5o3Niwzm4_2),.clk(gclk));
	jdff dff_B_9ZriKGjR7_2(.din(w_dff_B_5o3Niwzm4_2),.dout(w_dff_B_9ZriKGjR7_2),.clk(gclk));
	jdff dff_B_ITnjLgFq3_2(.din(w_dff_B_9ZriKGjR7_2),.dout(w_dff_B_ITnjLgFq3_2),.clk(gclk));
	jdff dff_B_OTbk8dQe3_2(.din(w_dff_B_ITnjLgFq3_2),.dout(w_dff_B_OTbk8dQe3_2),.clk(gclk));
	jdff dff_B_vAy7nKbo6_2(.din(w_dff_B_OTbk8dQe3_2),.dout(w_dff_B_vAy7nKbo6_2),.clk(gclk));
	jdff dff_B_zko9G0EF9_2(.din(w_dff_B_vAy7nKbo6_2),.dout(w_dff_B_zko9G0EF9_2),.clk(gclk));
	jdff dff_B_oewizM2L7_2(.din(w_dff_B_zko9G0EF9_2),.dout(w_dff_B_oewizM2L7_2),.clk(gclk));
	jdff dff_B_18rLPyg92_2(.din(w_dff_B_oewizM2L7_2),.dout(w_dff_B_18rLPyg92_2),.clk(gclk));
	jdff dff_B_AznkhTSe5_2(.din(w_dff_B_18rLPyg92_2),.dout(w_dff_B_AznkhTSe5_2),.clk(gclk));
	jdff dff_B_iRKK5uBZ5_2(.din(w_dff_B_AznkhTSe5_2),.dout(w_dff_B_iRKK5uBZ5_2),.clk(gclk));
	jdff dff_B_RDkpWgyC5_2(.din(w_dff_B_iRKK5uBZ5_2),.dout(w_dff_B_RDkpWgyC5_2),.clk(gclk));
	jdff dff_B_IsAT5oNE5_2(.din(w_dff_B_RDkpWgyC5_2),.dout(w_dff_B_IsAT5oNE5_2),.clk(gclk));
	jdff dff_B_vD33Rv5p3_2(.din(w_dff_B_IsAT5oNE5_2),.dout(w_dff_B_vD33Rv5p3_2),.clk(gclk));
	jdff dff_B_rBUDOAro5_2(.din(w_dff_B_vD33Rv5p3_2),.dout(w_dff_B_rBUDOAro5_2),.clk(gclk));
	jdff dff_B_xGeUXHEG8_2(.din(w_dff_B_rBUDOAro5_2),.dout(w_dff_B_xGeUXHEG8_2),.clk(gclk));
	jdff dff_B_8YpdBS5l8_2(.din(w_dff_B_xGeUXHEG8_2),.dout(w_dff_B_8YpdBS5l8_2),.clk(gclk));
	jdff dff_B_GpO173Qt0_2(.din(w_dff_B_8YpdBS5l8_2),.dout(w_dff_B_GpO173Qt0_2),.clk(gclk));
	jdff dff_B_jqf4z9hw4_2(.din(w_dff_B_GpO173Qt0_2),.dout(w_dff_B_jqf4z9hw4_2),.clk(gclk));
	jdff dff_B_v8qrSDt55_2(.din(w_dff_B_jqf4z9hw4_2),.dout(w_dff_B_v8qrSDt55_2),.clk(gclk));
	jdff dff_B_DqyOK3lR2_2(.din(w_dff_B_v8qrSDt55_2),.dout(w_dff_B_DqyOK3lR2_2),.clk(gclk));
	jdff dff_B_dRj1MpAd3_2(.din(w_dff_B_DqyOK3lR2_2),.dout(w_dff_B_dRj1MpAd3_2),.clk(gclk));
	jdff dff_B_hwZ1OtS52_2(.din(w_dff_B_dRj1MpAd3_2),.dout(w_dff_B_hwZ1OtS52_2),.clk(gclk));
	jdff dff_B_uqtKeENz7_2(.din(w_dff_B_hwZ1OtS52_2),.dout(w_dff_B_uqtKeENz7_2),.clk(gclk));
	jdff dff_A_SJbKKdsT3_0(.dout(w_n1008_0[0]),.din(w_dff_A_SJbKKdsT3_0),.clk(gclk));
	jdff dff_B_MBNG0AbL0_1(.din(n913),.dout(w_dff_B_MBNG0AbL0_1),.clk(gclk));
	jdff dff_B_3zDpu1uG9_2(.din(n811),.dout(w_dff_B_3zDpu1uG9_2),.clk(gclk));
	jdff dff_B_CHcGiAPZ2_2(.din(w_dff_B_3zDpu1uG9_2),.dout(w_dff_B_CHcGiAPZ2_2),.clk(gclk));
	jdff dff_B_pJq9naAp7_2(.din(w_dff_B_CHcGiAPZ2_2),.dout(w_dff_B_pJq9naAp7_2),.clk(gclk));
	jdff dff_B_f3TDEalf0_2(.din(w_dff_B_pJq9naAp7_2),.dout(w_dff_B_f3TDEalf0_2),.clk(gclk));
	jdff dff_B_YHBt6OSN9_2(.din(w_dff_B_f3TDEalf0_2),.dout(w_dff_B_YHBt6OSN9_2),.clk(gclk));
	jdff dff_B_okTx86I24_2(.din(w_dff_B_YHBt6OSN9_2),.dout(w_dff_B_okTx86I24_2),.clk(gclk));
	jdff dff_B_eaiiPk1C6_2(.din(w_dff_B_okTx86I24_2),.dout(w_dff_B_eaiiPk1C6_2),.clk(gclk));
	jdff dff_B_uWhg0wwL9_2(.din(w_dff_B_eaiiPk1C6_2),.dout(w_dff_B_uWhg0wwL9_2),.clk(gclk));
	jdff dff_B_p98dvSum8_2(.din(w_dff_B_uWhg0wwL9_2),.dout(w_dff_B_p98dvSum8_2),.clk(gclk));
	jdff dff_B_iF2JISr49_2(.din(w_dff_B_p98dvSum8_2),.dout(w_dff_B_iF2JISr49_2),.clk(gclk));
	jdff dff_B_ohKe0RqU3_2(.din(w_dff_B_iF2JISr49_2),.dout(w_dff_B_ohKe0RqU3_2),.clk(gclk));
	jdff dff_B_9l85lq9h1_2(.din(w_dff_B_ohKe0RqU3_2),.dout(w_dff_B_9l85lq9h1_2),.clk(gclk));
	jdff dff_B_3lihAQWP4_2(.din(w_dff_B_9l85lq9h1_2),.dout(w_dff_B_3lihAQWP4_2),.clk(gclk));
	jdff dff_B_I9ogKqkI5_2(.din(w_dff_B_3lihAQWP4_2),.dout(w_dff_B_I9ogKqkI5_2),.clk(gclk));
	jdff dff_B_okQiepVj7_2(.din(w_dff_B_I9ogKqkI5_2),.dout(w_dff_B_okQiepVj7_2),.clk(gclk));
	jdff dff_B_dwbuXAfJ5_2(.din(w_dff_B_okQiepVj7_2),.dout(w_dff_B_dwbuXAfJ5_2),.clk(gclk));
	jdff dff_B_IX0RCoAP0_2(.din(w_dff_B_dwbuXAfJ5_2),.dout(w_dff_B_IX0RCoAP0_2),.clk(gclk));
	jdff dff_B_3o8k60GS0_2(.din(w_dff_B_IX0RCoAP0_2),.dout(w_dff_B_3o8k60GS0_2),.clk(gclk));
	jdff dff_B_3vCIXG629_2(.din(w_dff_B_3o8k60GS0_2),.dout(w_dff_B_3vCIXG629_2),.clk(gclk));
	jdff dff_B_TrExfqNq4_2(.din(w_dff_B_3vCIXG629_2),.dout(w_dff_B_TrExfqNq4_2),.clk(gclk));
	jdff dff_B_GRPf8g8Q0_2(.din(w_dff_B_TrExfqNq4_2),.dout(w_dff_B_GRPf8g8Q0_2),.clk(gclk));
	jdff dff_B_3dPtBbZp2_2(.din(w_dff_B_GRPf8g8Q0_2),.dout(w_dff_B_3dPtBbZp2_2),.clk(gclk));
	jdff dff_B_Ye2pHaGy8_2(.din(w_dff_B_3dPtBbZp2_2),.dout(w_dff_B_Ye2pHaGy8_2),.clk(gclk));
	jdff dff_B_Q0GEHBCq2_2(.din(w_dff_B_Ye2pHaGy8_2),.dout(w_dff_B_Q0GEHBCq2_2),.clk(gclk));
	jdff dff_B_9lFcFSz02_2(.din(w_dff_B_Q0GEHBCq2_2),.dout(w_dff_B_9lFcFSz02_2),.clk(gclk));
	jdff dff_B_IjHXEw4x1_2(.din(w_dff_B_9lFcFSz02_2),.dout(w_dff_B_IjHXEw4x1_2),.clk(gclk));
	jdff dff_B_HGYISROJ9_2(.din(w_dff_B_IjHXEw4x1_2),.dout(w_dff_B_HGYISROJ9_2),.clk(gclk));
	jdff dff_B_HJFbp7XU5_2(.din(w_dff_B_HGYISROJ9_2),.dout(w_dff_B_HJFbp7XU5_2),.clk(gclk));
	jdff dff_B_oLNIsXrp1_2(.din(w_dff_B_HJFbp7XU5_2),.dout(w_dff_B_oLNIsXrp1_2),.clk(gclk));
	jdff dff_B_fJQXtMWB0_2(.din(w_dff_B_oLNIsXrp1_2),.dout(w_dff_B_fJQXtMWB0_2),.clk(gclk));
	jdff dff_B_fi0yePVZ9_2(.din(w_dff_B_fJQXtMWB0_2),.dout(w_dff_B_fi0yePVZ9_2),.clk(gclk));
	jdff dff_B_ZWF9xFTv5_2(.din(w_dff_B_fi0yePVZ9_2),.dout(w_dff_B_ZWF9xFTv5_2),.clk(gclk));
	jdff dff_B_9mFRgacX9_2(.din(w_dff_B_ZWF9xFTv5_2),.dout(w_dff_B_9mFRgacX9_2),.clk(gclk));
	jdff dff_B_uhTGuTUp1_2(.din(w_dff_B_9mFRgacX9_2),.dout(w_dff_B_uhTGuTUp1_2),.clk(gclk));
	jdff dff_B_yRDsDuK79_2(.din(w_dff_B_uhTGuTUp1_2),.dout(w_dff_B_yRDsDuK79_2),.clk(gclk));
	jdff dff_B_KNAFYxlh8_2(.din(w_dff_B_yRDsDuK79_2),.dout(w_dff_B_KNAFYxlh8_2),.clk(gclk));
	jdff dff_B_mnx6UzrJ5_2(.din(w_dff_B_KNAFYxlh8_2),.dout(w_dff_B_mnx6UzrJ5_2),.clk(gclk));
	jdff dff_B_stdMvYqh0_2(.din(w_dff_B_mnx6UzrJ5_2),.dout(w_dff_B_stdMvYqh0_2),.clk(gclk));
	jdff dff_B_s9GJJHbZ7_2(.din(w_dff_B_stdMvYqh0_2),.dout(w_dff_B_s9GJJHbZ7_2),.clk(gclk));
	jdff dff_B_jdynKIxI1_2(.din(w_dff_B_s9GJJHbZ7_2),.dout(w_dff_B_jdynKIxI1_2),.clk(gclk));
	jdff dff_A_0J86BOMG3_1(.dout(w_n902_0[1]),.din(w_dff_A_0J86BOMG3_1),.clk(gclk));
	jdff dff_B_EdhNsq102_1(.din(n817),.dout(w_dff_B_EdhNsq102_1),.clk(gclk));
	jdff dff_B_IebQ4pk39_1(.din(w_dff_B_EdhNsq102_1),.dout(w_dff_B_IebQ4pk39_1),.clk(gclk));
	jdff dff_B_NmxozeKk1_1(.din(w_dff_B_IebQ4pk39_1),.dout(w_dff_B_NmxozeKk1_1),.clk(gclk));
	jdff dff_B_K6QsIFnw8_1(.din(w_dff_B_NmxozeKk1_1),.dout(w_dff_B_K6QsIFnw8_1),.clk(gclk));
	jdff dff_B_saJiN6wL6_1(.din(w_dff_B_K6QsIFnw8_1),.dout(w_dff_B_saJiN6wL6_1),.clk(gclk));
	jdff dff_B_QGrHeXKe1_1(.din(w_dff_B_saJiN6wL6_1),.dout(w_dff_B_QGrHeXKe1_1),.clk(gclk));
	jdff dff_B_7amMLWih9_1(.din(w_dff_B_QGrHeXKe1_1),.dout(w_dff_B_7amMLWih9_1),.clk(gclk));
	jdff dff_B_cX4LMgoZ7_1(.din(w_dff_B_7amMLWih9_1),.dout(w_dff_B_cX4LMgoZ7_1),.clk(gclk));
	jdff dff_B_omE8ldRo9_1(.din(w_dff_B_cX4LMgoZ7_1),.dout(w_dff_B_omE8ldRo9_1),.clk(gclk));
	jdff dff_B_14GVMgo24_1(.din(w_dff_B_omE8ldRo9_1),.dout(w_dff_B_14GVMgo24_1),.clk(gclk));
	jdff dff_B_CM2GwsrS9_1(.din(w_dff_B_14GVMgo24_1),.dout(w_dff_B_CM2GwsrS9_1),.clk(gclk));
	jdff dff_B_2OXlzZFR3_1(.din(w_dff_B_CM2GwsrS9_1),.dout(w_dff_B_2OXlzZFR3_1),.clk(gclk));
	jdff dff_B_vkoctqO24_1(.din(w_dff_B_2OXlzZFR3_1),.dout(w_dff_B_vkoctqO24_1),.clk(gclk));
	jdff dff_B_s0ZM7l6K6_1(.din(w_dff_B_vkoctqO24_1),.dout(w_dff_B_s0ZM7l6K6_1),.clk(gclk));
	jdff dff_B_kAPEfvcS1_1(.din(w_dff_B_s0ZM7l6K6_1),.dout(w_dff_B_kAPEfvcS1_1),.clk(gclk));
	jdff dff_B_4cMlSNKW0_1(.din(w_dff_B_kAPEfvcS1_1),.dout(w_dff_B_4cMlSNKW0_1),.clk(gclk));
	jdff dff_B_jCZPZeE45_1(.din(w_dff_B_4cMlSNKW0_1),.dout(w_dff_B_jCZPZeE45_1),.clk(gclk));
	jdff dff_B_47NS7Vxr7_1(.din(w_dff_B_jCZPZeE45_1),.dout(w_dff_B_47NS7Vxr7_1),.clk(gclk));
	jdff dff_B_z7yEQTDj7_1(.din(w_dff_B_47NS7Vxr7_1),.dout(w_dff_B_z7yEQTDj7_1),.clk(gclk));
	jdff dff_B_kZjTMcG31_1(.din(w_dff_B_z7yEQTDj7_1),.dout(w_dff_B_kZjTMcG31_1),.clk(gclk));
	jdff dff_B_hX2jFXWD5_1(.din(w_dff_B_kZjTMcG31_1),.dout(w_dff_B_hX2jFXWD5_1),.clk(gclk));
	jdff dff_B_z79omYr96_1(.din(w_dff_B_hX2jFXWD5_1),.dout(w_dff_B_z79omYr96_1),.clk(gclk));
	jdff dff_B_P09nFvim3_1(.din(w_dff_B_z79omYr96_1),.dout(w_dff_B_P09nFvim3_1),.clk(gclk));
	jdff dff_B_Q5WHh9rV8_1(.din(w_dff_B_P09nFvim3_1),.dout(w_dff_B_Q5WHh9rV8_1),.clk(gclk));
	jdff dff_B_k9pIueEk0_1(.din(w_dff_B_Q5WHh9rV8_1),.dout(w_dff_B_k9pIueEk0_1),.clk(gclk));
	jdff dff_B_AFE9EtwD2_1(.din(w_dff_B_k9pIueEk0_1),.dout(w_dff_B_AFE9EtwD2_1),.clk(gclk));
	jdff dff_B_m7e5fpkE5_1(.din(w_dff_B_AFE9EtwD2_1),.dout(w_dff_B_m7e5fpkE5_1),.clk(gclk));
	jdff dff_B_rBbUcQQm5_1(.din(w_dff_B_m7e5fpkE5_1),.dout(w_dff_B_rBbUcQQm5_1),.clk(gclk));
	jdff dff_B_5AqhTg7e1_1(.din(w_dff_B_rBbUcQQm5_1),.dout(w_dff_B_5AqhTg7e1_1),.clk(gclk));
	jdff dff_B_fjZHzyNI5_1(.din(w_dff_B_5AqhTg7e1_1),.dout(w_dff_B_fjZHzyNI5_1),.clk(gclk));
	jdff dff_B_fOafkO0e6_1(.din(w_dff_B_fjZHzyNI5_1),.dout(w_dff_B_fOafkO0e6_1),.clk(gclk));
	jdff dff_B_RbOgAJPZ7_1(.din(w_dff_B_fOafkO0e6_1),.dout(w_dff_B_RbOgAJPZ7_1),.clk(gclk));
	jdff dff_B_EsJzeqQh8_1(.din(w_dff_B_RbOgAJPZ7_1),.dout(w_dff_B_EsJzeqQh8_1),.clk(gclk));
	jdff dff_B_nTuVxjpI5_1(.din(w_dff_B_EsJzeqQh8_1),.dout(w_dff_B_nTuVxjpI5_1),.clk(gclk));
	jdff dff_B_WHfx4DNR3_1(.din(w_dff_B_nTuVxjpI5_1),.dout(w_dff_B_WHfx4DNR3_1),.clk(gclk));
	jdff dff_B_ANn0WTHP7_1(.din(w_dff_B_WHfx4DNR3_1),.dout(w_dff_B_ANn0WTHP7_1),.clk(gclk));
	jdff dff_B_XlmD80Zn1_1(.din(n812),.dout(w_dff_B_XlmD80Zn1_1),.clk(gclk));
	jdff dff_A_5YWEty9W9_0(.dout(w_n712_0[0]),.din(w_dff_A_5YWEty9W9_0),.clk(gclk));
	jdff dff_A_6XViArYY6_0(.dout(w_dff_A_5YWEty9W9_0),.din(w_dff_A_6XViArYY6_0),.clk(gclk));
	jdff dff_A_D5A22Oee5_0(.dout(w_dff_A_6XViArYY6_0),.din(w_dff_A_D5A22Oee5_0),.clk(gclk));
	jdff dff_A_Q2yIbwww6_0(.dout(w_dff_A_D5A22Oee5_0),.din(w_dff_A_Q2yIbwww6_0),.clk(gclk));
	jdff dff_A_rRC4en4P9_0(.dout(w_dff_A_Q2yIbwww6_0),.din(w_dff_A_rRC4en4P9_0),.clk(gclk));
	jdff dff_A_xj8eh06L0_0(.dout(w_dff_A_rRC4en4P9_0),.din(w_dff_A_xj8eh06L0_0),.clk(gclk));
	jdff dff_A_9UKn3HFl5_0(.dout(w_dff_A_xj8eh06L0_0),.din(w_dff_A_9UKn3HFl5_0),.clk(gclk));
	jdff dff_A_o4Wctewa1_0(.dout(w_dff_A_9UKn3HFl5_0),.din(w_dff_A_o4Wctewa1_0),.clk(gclk));
	jdff dff_A_DZnSOfM64_0(.dout(w_dff_A_o4Wctewa1_0),.din(w_dff_A_DZnSOfM64_0),.clk(gclk));
	jdff dff_A_wnia88V73_0(.dout(w_dff_A_DZnSOfM64_0),.din(w_dff_A_wnia88V73_0),.clk(gclk));
	jdff dff_A_W5URmVKc2_0(.dout(w_dff_A_wnia88V73_0),.din(w_dff_A_W5URmVKc2_0),.clk(gclk));
	jdff dff_A_aHOFvn8s4_0(.dout(w_dff_A_W5URmVKc2_0),.din(w_dff_A_aHOFvn8s4_0),.clk(gclk));
	jdff dff_A_klRREsbW1_0(.dout(w_dff_A_aHOFvn8s4_0),.din(w_dff_A_klRREsbW1_0),.clk(gclk));
	jdff dff_A_o7ic6DTW2_0(.dout(w_dff_A_klRREsbW1_0),.din(w_dff_A_o7ic6DTW2_0),.clk(gclk));
	jdff dff_A_nvAytiyE1_0(.dout(w_dff_A_o7ic6DTW2_0),.din(w_dff_A_nvAytiyE1_0),.clk(gclk));
	jdff dff_A_PHVMzs0Y3_0(.dout(w_dff_A_nvAytiyE1_0),.din(w_dff_A_PHVMzs0Y3_0),.clk(gclk));
	jdff dff_A_raQoTS7M3_0(.dout(w_dff_A_PHVMzs0Y3_0),.din(w_dff_A_raQoTS7M3_0),.clk(gclk));
	jdff dff_A_OGxE8JX77_0(.dout(w_dff_A_raQoTS7M3_0),.din(w_dff_A_OGxE8JX77_0),.clk(gclk));
	jdff dff_A_px31xyQS5_0(.dout(w_dff_A_OGxE8JX77_0),.din(w_dff_A_px31xyQS5_0),.clk(gclk));
	jdff dff_A_YUgeAv468_0(.dout(w_dff_A_px31xyQS5_0),.din(w_dff_A_YUgeAv468_0),.clk(gclk));
	jdff dff_A_9QEbeaqf5_0(.dout(w_dff_A_YUgeAv468_0),.din(w_dff_A_9QEbeaqf5_0),.clk(gclk));
	jdff dff_A_zmXWwGoB8_0(.dout(w_dff_A_9QEbeaqf5_0),.din(w_dff_A_zmXWwGoB8_0),.clk(gclk));
	jdff dff_A_DJQN6eg72_0(.dout(w_dff_A_zmXWwGoB8_0),.din(w_dff_A_DJQN6eg72_0),.clk(gclk));
	jdff dff_A_nbrH8tmC0_0(.dout(w_dff_A_DJQN6eg72_0),.din(w_dff_A_nbrH8tmC0_0),.clk(gclk));
	jdff dff_A_ovVpdRfI5_0(.dout(w_dff_A_nbrH8tmC0_0),.din(w_dff_A_ovVpdRfI5_0),.clk(gclk));
	jdff dff_A_x2UNeOZM1_0(.dout(w_dff_A_ovVpdRfI5_0),.din(w_dff_A_x2UNeOZM1_0),.clk(gclk));
	jdff dff_A_lsJ0nEbo7_0(.dout(w_dff_A_x2UNeOZM1_0),.din(w_dff_A_lsJ0nEbo7_0),.clk(gclk));
	jdff dff_A_pWtxQTJB2_0(.dout(w_dff_A_lsJ0nEbo7_0),.din(w_dff_A_pWtxQTJB2_0),.clk(gclk));
	jdff dff_A_M473xJ4v7_0(.dout(w_dff_A_pWtxQTJB2_0),.din(w_dff_A_M473xJ4v7_0),.clk(gclk));
	jdff dff_A_FZFd6F855_0(.dout(w_dff_A_M473xJ4v7_0),.din(w_dff_A_FZFd6F855_0),.clk(gclk));
	jdff dff_A_udFgmkA59_0(.dout(w_dff_A_FZFd6F855_0),.din(w_dff_A_udFgmkA59_0),.clk(gclk));
	jdff dff_A_fWc4L2vd3_0(.dout(w_dff_A_udFgmkA59_0),.din(w_dff_A_fWc4L2vd3_0),.clk(gclk));
	jdff dff_A_jnF6Pakn5_0(.dout(w_dff_A_fWc4L2vd3_0),.din(w_dff_A_jnF6Pakn5_0),.clk(gclk));
	jdff dff_A_4FhdXpys8_0(.dout(w_dff_A_jnF6Pakn5_0),.din(w_dff_A_4FhdXpys8_0),.clk(gclk));
	jdff dff_A_aX74ePjH3_0(.dout(w_dff_A_4FhdXpys8_0),.din(w_dff_A_aX74ePjH3_0),.clk(gclk));
	jdff dff_A_Zaf6Ilxr6_0(.dout(w_dff_A_aX74ePjH3_0),.din(w_dff_A_Zaf6Ilxr6_0),.clk(gclk));
	jdff dff_A_4ptKqsnL1_0(.dout(w_dff_A_Zaf6Ilxr6_0),.din(w_dff_A_4ptKqsnL1_0),.clk(gclk));
	jdff dff_A_S6FwpfXP2_0(.dout(w_n799_0[0]),.din(w_dff_A_S6FwpfXP2_0),.clk(gclk));
	jdff dff_B_pflvUWRu2_1(.din(n714),.dout(w_dff_B_pflvUWRu2_1),.clk(gclk));
	jdff dff_A_BkMzg41H7_0(.dout(w_n620_0[0]),.din(w_dff_A_BkMzg41H7_0),.clk(gclk));
	jdff dff_A_874bzRIp1_0(.dout(w_dff_A_BkMzg41H7_0),.din(w_dff_A_874bzRIp1_0),.clk(gclk));
	jdff dff_A_Pi9kDOzQ8_0(.dout(w_dff_A_874bzRIp1_0),.din(w_dff_A_Pi9kDOzQ8_0),.clk(gclk));
	jdff dff_A_FjrK4XQF9_0(.dout(w_dff_A_Pi9kDOzQ8_0),.din(w_dff_A_FjrK4XQF9_0),.clk(gclk));
	jdff dff_A_BD4R69X74_0(.dout(w_dff_A_FjrK4XQF9_0),.din(w_dff_A_BD4R69X74_0),.clk(gclk));
	jdff dff_A_5H5Mfybo4_0(.dout(w_dff_A_BD4R69X74_0),.din(w_dff_A_5H5Mfybo4_0),.clk(gclk));
	jdff dff_A_6Al7Lf9H1_0(.dout(w_dff_A_5H5Mfybo4_0),.din(w_dff_A_6Al7Lf9H1_0),.clk(gclk));
	jdff dff_A_h45etCDT9_0(.dout(w_dff_A_6Al7Lf9H1_0),.din(w_dff_A_h45etCDT9_0),.clk(gclk));
	jdff dff_A_yarTC1jo8_0(.dout(w_dff_A_h45etCDT9_0),.din(w_dff_A_yarTC1jo8_0),.clk(gclk));
	jdff dff_A_pnXH4Ybz6_0(.dout(w_dff_A_yarTC1jo8_0),.din(w_dff_A_pnXH4Ybz6_0),.clk(gclk));
	jdff dff_A_xuWaMKId7_0(.dout(w_dff_A_pnXH4Ybz6_0),.din(w_dff_A_xuWaMKId7_0),.clk(gclk));
	jdff dff_A_TLnCxtf08_0(.dout(w_dff_A_xuWaMKId7_0),.din(w_dff_A_TLnCxtf08_0),.clk(gclk));
	jdff dff_A_hJupKqFd2_0(.dout(w_dff_A_TLnCxtf08_0),.din(w_dff_A_hJupKqFd2_0),.clk(gclk));
	jdff dff_A_wqnVDYpm4_0(.dout(w_dff_A_hJupKqFd2_0),.din(w_dff_A_wqnVDYpm4_0),.clk(gclk));
	jdff dff_A_H6lXtifl8_0(.dout(w_dff_A_wqnVDYpm4_0),.din(w_dff_A_H6lXtifl8_0),.clk(gclk));
	jdff dff_A_0o9ep4IJ2_0(.dout(w_dff_A_H6lXtifl8_0),.din(w_dff_A_0o9ep4IJ2_0),.clk(gclk));
	jdff dff_A_ngNl0rDB5_0(.dout(w_dff_A_0o9ep4IJ2_0),.din(w_dff_A_ngNl0rDB5_0),.clk(gclk));
	jdff dff_A_MF5G3qvD7_0(.dout(w_dff_A_ngNl0rDB5_0),.din(w_dff_A_MF5G3qvD7_0),.clk(gclk));
	jdff dff_A_u91J4fVZ0_0(.dout(w_dff_A_MF5G3qvD7_0),.din(w_dff_A_u91J4fVZ0_0),.clk(gclk));
	jdff dff_A_SFzKZ4Af7_0(.dout(w_dff_A_u91J4fVZ0_0),.din(w_dff_A_SFzKZ4Af7_0),.clk(gclk));
	jdff dff_A_omaWsmV62_0(.dout(w_dff_A_SFzKZ4Af7_0),.din(w_dff_A_omaWsmV62_0),.clk(gclk));
	jdff dff_A_yzbQNLsX6_0(.dout(w_dff_A_omaWsmV62_0),.din(w_dff_A_yzbQNLsX6_0),.clk(gclk));
	jdff dff_A_dz7BvYCT4_0(.dout(w_dff_A_yzbQNLsX6_0),.din(w_dff_A_dz7BvYCT4_0),.clk(gclk));
	jdff dff_A_2RHVdoY11_0(.dout(w_dff_A_dz7BvYCT4_0),.din(w_dff_A_2RHVdoY11_0),.clk(gclk));
	jdff dff_A_Gbvra4eQ6_0(.dout(w_dff_A_2RHVdoY11_0),.din(w_dff_A_Gbvra4eQ6_0),.clk(gclk));
	jdff dff_A_1ACIXW4Q5_0(.dout(w_dff_A_Gbvra4eQ6_0),.din(w_dff_A_1ACIXW4Q5_0),.clk(gclk));
	jdff dff_A_09Sa6nK39_0(.dout(w_dff_A_1ACIXW4Q5_0),.din(w_dff_A_09Sa6nK39_0),.clk(gclk));
	jdff dff_A_hUZRuwci2_0(.dout(w_dff_A_09Sa6nK39_0),.din(w_dff_A_hUZRuwci2_0),.clk(gclk));
	jdff dff_A_lzu8y0t96_0(.dout(w_dff_A_hUZRuwci2_0),.din(w_dff_A_lzu8y0t96_0),.clk(gclk));
	jdff dff_A_TZN8eWhu9_0(.dout(w_dff_A_lzu8y0t96_0),.din(w_dff_A_TZN8eWhu9_0),.clk(gclk));
	jdff dff_A_RE0eJ62Y9_0(.dout(w_dff_A_TZN8eWhu9_0),.din(w_dff_A_RE0eJ62Y9_0),.clk(gclk));
	jdff dff_A_zSfyDgec7_0(.dout(w_dff_A_RE0eJ62Y9_0),.din(w_dff_A_zSfyDgec7_0),.clk(gclk));
	jdff dff_A_ukLUEFGu4_0(.dout(w_dff_A_zSfyDgec7_0),.din(w_dff_A_ukLUEFGu4_0),.clk(gclk));
	jdff dff_A_tq7qiosp1_0(.dout(w_dff_A_ukLUEFGu4_0),.din(w_dff_A_tq7qiosp1_0),.clk(gclk));
	jdff dff_A_0YxJ5nxx6_0(.dout(w_n700_0[0]),.din(w_dff_A_0YxJ5nxx6_0),.clk(gclk));
	jdff dff_B_pjmkXbrx0_1(.din(n622),.dout(w_dff_B_pjmkXbrx0_1),.clk(gclk));
	jdff dff_A_hPP2WvLp3_0(.dout(w_n535_0[0]),.din(w_dff_A_hPP2WvLp3_0),.clk(gclk));
	jdff dff_A_ZcpJgxuk2_0(.dout(w_dff_A_hPP2WvLp3_0),.din(w_dff_A_ZcpJgxuk2_0),.clk(gclk));
	jdff dff_A_H7YS8Hq79_0(.dout(w_dff_A_ZcpJgxuk2_0),.din(w_dff_A_H7YS8Hq79_0),.clk(gclk));
	jdff dff_A_RdgYIqt98_0(.dout(w_dff_A_H7YS8Hq79_0),.din(w_dff_A_RdgYIqt98_0),.clk(gclk));
	jdff dff_A_UnLDxG4N4_0(.dout(w_dff_A_RdgYIqt98_0),.din(w_dff_A_UnLDxG4N4_0),.clk(gclk));
	jdff dff_A_cwA9ZUkH5_0(.dout(w_dff_A_UnLDxG4N4_0),.din(w_dff_A_cwA9ZUkH5_0),.clk(gclk));
	jdff dff_A_pVk3wPz71_0(.dout(w_dff_A_cwA9ZUkH5_0),.din(w_dff_A_pVk3wPz71_0),.clk(gclk));
	jdff dff_A_YgW0X4hY4_0(.dout(w_dff_A_pVk3wPz71_0),.din(w_dff_A_YgW0X4hY4_0),.clk(gclk));
	jdff dff_A_uPymbpzY0_0(.dout(w_dff_A_YgW0X4hY4_0),.din(w_dff_A_uPymbpzY0_0),.clk(gclk));
	jdff dff_A_nxYo3GfB3_0(.dout(w_dff_A_uPymbpzY0_0),.din(w_dff_A_nxYo3GfB3_0),.clk(gclk));
	jdff dff_A_hys25FMj2_0(.dout(w_dff_A_nxYo3GfB3_0),.din(w_dff_A_hys25FMj2_0),.clk(gclk));
	jdff dff_A_xiTh05Q15_0(.dout(w_dff_A_hys25FMj2_0),.din(w_dff_A_xiTh05Q15_0),.clk(gclk));
	jdff dff_A_5NdCmXGl7_0(.dout(w_dff_A_xiTh05Q15_0),.din(w_dff_A_5NdCmXGl7_0),.clk(gclk));
	jdff dff_A_q5tHYBIt7_0(.dout(w_dff_A_5NdCmXGl7_0),.din(w_dff_A_q5tHYBIt7_0),.clk(gclk));
	jdff dff_A_I30KBgqn4_0(.dout(w_dff_A_q5tHYBIt7_0),.din(w_dff_A_I30KBgqn4_0),.clk(gclk));
	jdff dff_A_eCCRbfEC2_0(.dout(w_dff_A_I30KBgqn4_0),.din(w_dff_A_eCCRbfEC2_0),.clk(gclk));
	jdff dff_A_GzUIL9WD9_0(.dout(w_dff_A_eCCRbfEC2_0),.din(w_dff_A_GzUIL9WD9_0),.clk(gclk));
	jdff dff_A_Xhc8ANEq3_0(.dout(w_dff_A_GzUIL9WD9_0),.din(w_dff_A_Xhc8ANEq3_0),.clk(gclk));
	jdff dff_A_aKybp6xT8_0(.dout(w_dff_A_Xhc8ANEq3_0),.din(w_dff_A_aKybp6xT8_0),.clk(gclk));
	jdff dff_A_amGNss0t3_0(.dout(w_dff_A_aKybp6xT8_0),.din(w_dff_A_amGNss0t3_0),.clk(gclk));
	jdff dff_A_3NjSbybY7_0(.dout(w_dff_A_amGNss0t3_0),.din(w_dff_A_3NjSbybY7_0),.clk(gclk));
	jdff dff_A_8mluqX3F5_0(.dout(w_dff_A_3NjSbybY7_0),.din(w_dff_A_8mluqX3F5_0),.clk(gclk));
	jdff dff_A_2JlJnlK45_0(.dout(w_dff_A_8mluqX3F5_0),.din(w_dff_A_2JlJnlK45_0),.clk(gclk));
	jdff dff_A_x2F3LTla3_0(.dout(w_dff_A_2JlJnlK45_0),.din(w_dff_A_x2F3LTla3_0),.clk(gclk));
	jdff dff_A_XxstEwhI9_0(.dout(w_dff_A_x2F3LTla3_0),.din(w_dff_A_XxstEwhI9_0),.clk(gclk));
	jdff dff_A_yMGypQkr1_0(.dout(w_dff_A_XxstEwhI9_0),.din(w_dff_A_yMGypQkr1_0),.clk(gclk));
	jdff dff_A_B9Q8kb3U8_0(.dout(w_dff_A_yMGypQkr1_0),.din(w_dff_A_B9Q8kb3U8_0),.clk(gclk));
	jdff dff_A_idSjjSXm6_0(.dout(w_dff_A_B9Q8kb3U8_0),.din(w_dff_A_idSjjSXm6_0),.clk(gclk));
	jdff dff_A_khsGPbNH3_0(.dout(w_dff_A_idSjjSXm6_0),.din(w_dff_A_khsGPbNH3_0),.clk(gclk));
	jdff dff_A_cZKhTl2L2_0(.dout(w_dff_A_khsGPbNH3_0),.din(w_dff_A_cZKhTl2L2_0),.clk(gclk));
	jdff dff_A_fKn3qFcf1_0(.dout(w_dff_A_cZKhTl2L2_0),.din(w_dff_A_fKn3qFcf1_0),.clk(gclk));
	jdff dff_A_u6y9dCsG3_0(.dout(w_n608_0[0]),.din(w_dff_A_u6y9dCsG3_0),.clk(gclk));
	jdff dff_B_NqzeNCcz1_1(.din(n537),.dout(w_dff_B_NqzeNCcz1_1),.clk(gclk));
	jdff dff_A_4xmEb0ep2_0(.dout(w_n457_0[0]),.din(w_dff_A_4xmEb0ep2_0),.clk(gclk));
	jdff dff_A_IEYs6iOb1_0(.dout(w_dff_A_4xmEb0ep2_0),.din(w_dff_A_IEYs6iOb1_0),.clk(gclk));
	jdff dff_A_k9fkmrUQ1_0(.dout(w_dff_A_IEYs6iOb1_0),.din(w_dff_A_k9fkmrUQ1_0),.clk(gclk));
	jdff dff_A_yYqPLQi00_0(.dout(w_dff_A_k9fkmrUQ1_0),.din(w_dff_A_yYqPLQi00_0),.clk(gclk));
	jdff dff_A_UTnePFQt5_0(.dout(w_dff_A_yYqPLQi00_0),.din(w_dff_A_UTnePFQt5_0),.clk(gclk));
	jdff dff_A_r34x6rcn3_0(.dout(w_dff_A_UTnePFQt5_0),.din(w_dff_A_r34x6rcn3_0),.clk(gclk));
	jdff dff_A_RhVxffoR6_0(.dout(w_dff_A_r34x6rcn3_0),.din(w_dff_A_RhVxffoR6_0),.clk(gclk));
	jdff dff_A_dUmpYrUh4_0(.dout(w_dff_A_RhVxffoR6_0),.din(w_dff_A_dUmpYrUh4_0),.clk(gclk));
	jdff dff_A_psyDIvGL7_0(.dout(w_dff_A_dUmpYrUh4_0),.din(w_dff_A_psyDIvGL7_0),.clk(gclk));
	jdff dff_A_lbgNL8dD1_0(.dout(w_dff_A_psyDIvGL7_0),.din(w_dff_A_lbgNL8dD1_0),.clk(gclk));
	jdff dff_A_Bp7fFiIQ8_0(.dout(w_dff_A_lbgNL8dD1_0),.din(w_dff_A_Bp7fFiIQ8_0),.clk(gclk));
	jdff dff_A_PZTquga30_0(.dout(w_dff_A_Bp7fFiIQ8_0),.din(w_dff_A_PZTquga30_0),.clk(gclk));
	jdff dff_A_kVWIOkab1_0(.dout(w_dff_A_PZTquga30_0),.din(w_dff_A_kVWIOkab1_0),.clk(gclk));
	jdff dff_A_fNLZtWMb5_0(.dout(w_dff_A_kVWIOkab1_0),.din(w_dff_A_fNLZtWMb5_0),.clk(gclk));
	jdff dff_A_Q1hC4ogO9_0(.dout(w_dff_A_fNLZtWMb5_0),.din(w_dff_A_Q1hC4ogO9_0),.clk(gclk));
	jdff dff_A_s0ukA6Jz5_0(.dout(w_dff_A_Q1hC4ogO9_0),.din(w_dff_A_s0ukA6Jz5_0),.clk(gclk));
	jdff dff_A_KuEc4sXA8_0(.dout(w_dff_A_s0ukA6Jz5_0),.din(w_dff_A_KuEc4sXA8_0),.clk(gclk));
	jdff dff_A_qKHTRJsL6_0(.dout(w_dff_A_KuEc4sXA8_0),.din(w_dff_A_qKHTRJsL6_0),.clk(gclk));
	jdff dff_A_UuOZMD157_0(.dout(w_dff_A_qKHTRJsL6_0),.din(w_dff_A_UuOZMD157_0),.clk(gclk));
	jdff dff_A_crLqfn9P2_0(.dout(w_dff_A_UuOZMD157_0),.din(w_dff_A_crLqfn9P2_0),.clk(gclk));
	jdff dff_A_nEeZKSXp7_0(.dout(w_dff_A_crLqfn9P2_0),.din(w_dff_A_nEeZKSXp7_0),.clk(gclk));
	jdff dff_A_ehHhY8Ci6_0(.dout(w_dff_A_nEeZKSXp7_0),.din(w_dff_A_ehHhY8Ci6_0),.clk(gclk));
	jdff dff_A_1HutRfl41_0(.dout(w_dff_A_ehHhY8Ci6_0),.din(w_dff_A_1HutRfl41_0),.clk(gclk));
	jdff dff_A_t7R1ENKv3_0(.dout(w_dff_A_1HutRfl41_0),.din(w_dff_A_t7R1ENKv3_0),.clk(gclk));
	jdff dff_A_jPX4NgYz5_0(.dout(w_dff_A_t7R1ENKv3_0),.din(w_dff_A_jPX4NgYz5_0),.clk(gclk));
	jdff dff_A_PucVo6wk5_0(.dout(w_dff_A_jPX4NgYz5_0),.din(w_dff_A_PucVo6wk5_0),.clk(gclk));
	jdff dff_A_lY6R6JyL6_0(.dout(w_dff_A_PucVo6wk5_0),.din(w_dff_A_lY6R6JyL6_0),.clk(gclk));
	jdff dff_A_qmqeJ4rw5_0(.dout(w_dff_A_lY6R6JyL6_0),.din(w_dff_A_qmqeJ4rw5_0),.clk(gclk));
	jdff dff_A_fQs3s16e9_0(.dout(w_n523_0[0]),.din(w_dff_A_fQs3s16e9_0),.clk(gclk));
	jdff dff_B_qGdEvmpm9_1(.din(n459),.dout(w_dff_B_qGdEvmpm9_1),.clk(gclk));
	jdff dff_A_vKobrcIW5_0(.dout(w_n386_0[0]),.din(w_dff_A_vKobrcIW5_0),.clk(gclk));
	jdff dff_A_vmQOtDJF2_0(.dout(w_dff_A_vKobrcIW5_0),.din(w_dff_A_vmQOtDJF2_0),.clk(gclk));
	jdff dff_A_3gmszpDI1_0(.dout(w_dff_A_vmQOtDJF2_0),.din(w_dff_A_3gmszpDI1_0),.clk(gclk));
	jdff dff_A_jt63r7Nx0_0(.dout(w_dff_A_3gmszpDI1_0),.din(w_dff_A_jt63r7Nx0_0),.clk(gclk));
	jdff dff_A_RusFWgCS9_0(.dout(w_dff_A_jt63r7Nx0_0),.din(w_dff_A_RusFWgCS9_0),.clk(gclk));
	jdff dff_A_ikiqNDu64_0(.dout(w_dff_A_RusFWgCS9_0),.din(w_dff_A_ikiqNDu64_0),.clk(gclk));
	jdff dff_A_hu30fkaM2_0(.dout(w_dff_A_ikiqNDu64_0),.din(w_dff_A_hu30fkaM2_0),.clk(gclk));
	jdff dff_A_CcKmnVpu3_0(.dout(w_dff_A_hu30fkaM2_0),.din(w_dff_A_CcKmnVpu3_0),.clk(gclk));
	jdff dff_A_siJIrCQB3_0(.dout(w_dff_A_CcKmnVpu3_0),.din(w_dff_A_siJIrCQB3_0),.clk(gclk));
	jdff dff_A_bnMv18Mk7_0(.dout(w_dff_A_siJIrCQB3_0),.din(w_dff_A_bnMv18Mk7_0),.clk(gclk));
	jdff dff_A_anY4MMgQ7_0(.dout(w_dff_A_bnMv18Mk7_0),.din(w_dff_A_anY4MMgQ7_0),.clk(gclk));
	jdff dff_A_4wqqoZNz3_0(.dout(w_dff_A_anY4MMgQ7_0),.din(w_dff_A_4wqqoZNz3_0),.clk(gclk));
	jdff dff_A_y5FNnRqY6_0(.dout(w_dff_A_4wqqoZNz3_0),.din(w_dff_A_y5FNnRqY6_0),.clk(gclk));
	jdff dff_A_i3q8QPFv4_0(.dout(w_dff_A_y5FNnRqY6_0),.din(w_dff_A_i3q8QPFv4_0),.clk(gclk));
	jdff dff_A_yjZQIPzv6_0(.dout(w_dff_A_i3q8QPFv4_0),.din(w_dff_A_yjZQIPzv6_0),.clk(gclk));
	jdff dff_A_yp7xCUph3_0(.dout(w_dff_A_yjZQIPzv6_0),.din(w_dff_A_yp7xCUph3_0),.clk(gclk));
	jdff dff_A_zAEsPfJ83_0(.dout(w_dff_A_yp7xCUph3_0),.din(w_dff_A_zAEsPfJ83_0),.clk(gclk));
	jdff dff_A_0RY2ywOg5_0(.dout(w_dff_A_zAEsPfJ83_0),.din(w_dff_A_0RY2ywOg5_0),.clk(gclk));
	jdff dff_A_Nqp6xeQH0_0(.dout(w_dff_A_0RY2ywOg5_0),.din(w_dff_A_Nqp6xeQH0_0),.clk(gclk));
	jdff dff_A_fGGLGsqf4_0(.dout(w_dff_A_Nqp6xeQH0_0),.din(w_dff_A_fGGLGsqf4_0),.clk(gclk));
	jdff dff_A_nYBXpLvA8_0(.dout(w_dff_A_fGGLGsqf4_0),.din(w_dff_A_nYBXpLvA8_0),.clk(gclk));
	jdff dff_A_XW5iWM399_0(.dout(w_dff_A_nYBXpLvA8_0),.din(w_dff_A_XW5iWM399_0),.clk(gclk));
	jdff dff_A_ULGsBPMI9_0(.dout(w_dff_A_XW5iWM399_0),.din(w_dff_A_ULGsBPMI9_0),.clk(gclk));
	jdff dff_A_MUa2RZ6j8_0(.dout(w_dff_A_ULGsBPMI9_0),.din(w_dff_A_MUa2RZ6j8_0),.clk(gclk));
	jdff dff_A_tCowXLRu0_0(.dout(w_dff_A_MUa2RZ6j8_0),.din(w_dff_A_tCowXLRu0_0),.clk(gclk));
	jdff dff_A_pU4uyEYh8_0(.dout(w_n445_0[0]),.din(w_dff_A_pU4uyEYh8_0),.clk(gclk));
	jdff dff_B_jnPhVbWa4_1(.din(n388),.dout(w_dff_B_jnPhVbWa4_1),.clk(gclk));
	jdff dff_A_c9CUVApT3_0(.dout(w_n323_0[0]),.din(w_dff_A_c9CUVApT3_0),.clk(gclk));
	jdff dff_A_Wd4YsLYq3_0(.dout(w_dff_A_c9CUVApT3_0),.din(w_dff_A_Wd4YsLYq3_0),.clk(gclk));
	jdff dff_A_I1gyvQs00_0(.dout(w_dff_A_Wd4YsLYq3_0),.din(w_dff_A_I1gyvQs00_0),.clk(gclk));
	jdff dff_A_9YYawam92_0(.dout(w_dff_A_I1gyvQs00_0),.din(w_dff_A_9YYawam92_0),.clk(gclk));
	jdff dff_A_MK6i0Hfr3_0(.dout(w_dff_A_9YYawam92_0),.din(w_dff_A_MK6i0Hfr3_0),.clk(gclk));
	jdff dff_A_c5ArgNKk2_0(.dout(w_dff_A_MK6i0Hfr3_0),.din(w_dff_A_c5ArgNKk2_0),.clk(gclk));
	jdff dff_A_YXKh3GUv6_0(.dout(w_dff_A_c5ArgNKk2_0),.din(w_dff_A_YXKh3GUv6_0),.clk(gclk));
	jdff dff_A_GG1B0wA87_0(.dout(w_dff_A_YXKh3GUv6_0),.din(w_dff_A_GG1B0wA87_0),.clk(gclk));
	jdff dff_A_DdIj7Hqy1_0(.dout(w_dff_A_GG1B0wA87_0),.din(w_dff_A_DdIj7Hqy1_0),.clk(gclk));
	jdff dff_A_Pf1ejpuG9_0(.dout(w_dff_A_DdIj7Hqy1_0),.din(w_dff_A_Pf1ejpuG9_0),.clk(gclk));
	jdff dff_A_GibrthsK2_0(.dout(w_dff_A_Pf1ejpuG9_0),.din(w_dff_A_GibrthsK2_0),.clk(gclk));
	jdff dff_A_47anQ0hc8_0(.dout(w_dff_A_GibrthsK2_0),.din(w_dff_A_47anQ0hc8_0),.clk(gclk));
	jdff dff_A_x5WIydQU3_0(.dout(w_dff_A_47anQ0hc8_0),.din(w_dff_A_x5WIydQU3_0),.clk(gclk));
	jdff dff_A_VgvozxVI6_0(.dout(w_dff_A_x5WIydQU3_0),.din(w_dff_A_VgvozxVI6_0),.clk(gclk));
	jdff dff_A_qaKzyUob6_0(.dout(w_dff_A_VgvozxVI6_0),.din(w_dff_A_qaKzyUob6_0),.clk(gclk));
	jdff dff_A_ezOmsEHF8_0(.dout(w_dff_A_qaKzyUob6_0),.din(w_dff_A_ezOmsEHF8_0),.clk(gclk));
	jdff dff_A_ZMOCpJGr0_0(.dout(w_dff_A_ezOmsEHF8_0),.din(w_dff_A_ZMOCpJGr0_0),.clk(gclk));
	jdff dff_A_Ous7uqdB9_0(.dout(w_dff_A_ZMOCpJGr0_0),.din(w_dff_A_Ous7uqdB9_0),.clk(gclk));
	jdff dff_A_yozDzvJL8_0(.dout(w_dff_A_Ous7uqdB9_0),.din(w_dff_A_yozDzvJL8_0),.clk(gclk));
	jdff dff_A_vZC30y7j0_0(.dout(w_dff_A_yozDzvJL8_0),.din(w_dff_A_vZC30y7j0_0),.clk(gclk));
	jdff dff_A_QjGsalrL6_0(.dout(w_dff_A_vZC30y7j0_0),.din(w_dff_A_QjGsalrL6_0),.clk(gclk));
	jdff dff_A_RqtKQE7V3_0(.dout(w_dff_A_QjGsalrL6_0),.din(w_dff_A_RqtKQE7V3_0),.clk(gclk));
	jdff dff_A_CDV3PFhs0_0(.dout(w_n374_0[0]),.din(w_dff_A_CDV3PFhs0_0),.clk(gclk));
	jdff dff_B_s7OczH1C1_1(.din(n325),.dout(w_dff_B_s7OczH1C1_1),.clk(gclk));
	jdff dff_A_EWcRos1r1_0(.dout(w_n267_0[0]),.din(w_dff_A_EWcRos1r1_0),.clk(gclk));
	jdff dff_A_Qppmjvlc5_0(.dout(w_dff_A_EWcRos1r1_0),.din(w_dff_A_Qppmjvlc5_0),.clk(gclk));
	jdff dff_A_JTkS87u49_0(.dout(w_dff_A_Qppmjvlc5_0),.din(w_dff_A_JTkS87u49_0),.clk(gclk));
	jdff dff_A_EgBelY8x3_0(.dout(w_dff_A_JTkS87u49_0),.din(w_dff_A_EgBelY8x3_0),.clk(gclk));
	jdff dff_A_ooDQBnt85_0(.dout(w_dff_A_EgBelY8x3_0),.din(w_dff_A_ooDQBnt85_0),.clk(gclk));
	jdff dff_A_OVkuv4Hf3_0(.dout(w_dff_A_ooDQBnt85_0),.din(w_dff_A_OVkuv4Hf3_0),.clk(gclk));
	jdff dff_A_WgdkfFkG3_0(.dout(w_dff_A_OVkuv4Hf3_0),.din(w_dff_A_WgdkfFkG3_0),.clk(gclk));
	jdff dff_A_rYNFFamI9_0(.dout(w_dff_A_WgdkfFkG3_0),.din(w_dff_A_rYNFFamI9_0),.clk(gclk));
	jdff dff_A_IhCktVbw2_0(.dout(w_dff_A_rYNFFamI9_0),.din(w_dff_A_IhCktVbw2_0),.clk(gclk));
	jdff dff_A_HTjec5nu6_0(.dout(w_dff_A_IhCktVbw2_0),.din(w_dff_A_HTjec5nu6_0),.clk(gclk));
	jdff dff_A_LCKHzrEY8_0(.dout(w_dff_A_HTjec5nu6_0),.din(w_dff_A_LCKHzrEY8_0),.clk(gclk));
	jdff dff_A_gPa4Tju61_0(.dout(w_dff_A_LCKHzrEY8_0),.din(w_dff_A_gPa4Tju61_0),.clk(gclk));
	jdff dff_A_DGqGTPOR1_0(.dout(w_dff_A_gPa4Tju61_0),.din(w_dff_A_DGqGTPOR1_0),.clk(gclk));
	jdff dff_A_5V4KukZA8_0(.dout(w_dff_A_DGqGTPOR1_0),.din(w_dff_A_5V4KukZA8_0),.clk(gclk));
	jdff dff_A_vlyGCtiS8_0(.dout(w_dff_A_5V4KukZA8_0),.din(w_dff_A_vlyGCtiS8_0),.clk(gclk));
	jdff dff_A_x7l1k7f49_0(.dout(w_dff_A_vlyGCtiS8_0),.din(w_dff_A_x7l1k7f49_0),.clk(gclk));
	jdff dff_A_3FW2y6830_0(.dout(w_dff_A_x7l1k7f49_0),.din(w_dff_A_3FW2y6830_0),.clk(gclk));
	jdff dff_A_7bKFNt5E9_0(.dout(w_dff_A_3FW2y6830_0),.din(w_dff_A_7bKFNt5E9_0),.clk(gclk));
	jdff dff_A_Ob6ywave7_0(.dout(w_dff_A_7bKFNt5E9_0),.din(w_dff_A_Ob6ywave7_0),.clk(gclk));
	jdff dff_A_WKLMPdYf9_0(.dout(w_n311_0[0]),.din(w_dff_A_WKLMPdYf9_0),.clk(gclk));
	jdff dff_B_6xod8Z1X3_1(.din(n269),.dout(w_dff_B_6xod8Z1X3_1),.clk(gclk));
	jdff dff_A_gWXZKh5j0_0(.dout(w_n218_0[0]),.din(w_dff_A_gWXZKh5j0_0),.clk(gclk));
	jdff dff_A_4ygwGMfm1_0(.dout(w_dff_A_gWXZKh5j0_0),.din(w_dff_A_4ygwGMfm1_0),.clk(gclk));
	jdff dff_A_jKOssVq52_0(.dout(w_dff_A_4ygwGMfm1_0),.din(w_dff_A_jKOssVq52_0),.clk(gclk));
	jdff dff_A_nXeguX2d5_0(.dout(w_dff_A_jKOssVq52_0),.din(w_dff_A_nXeguX2d5_0),.clk(gclk));
	jdff dff_A_47b6gRoU0_0(.dout(w_dff_A_nXeguX2d5_0),.din(w_dff_A_47b6gRoU0_0),.clk(gclk));
	jdff dff_A_dlWJZGOb0_0(.dout(w_dff_A_47b6gRoU0_0),.din(w_dff_A_dlWJZGOb0_0),.clk(gclk));
	jdff dff_A_Qp4jWFqG9_0(.dout(w_dff_A_dlWJZGOb0_0),.din(w_dff_A_Qp4jWFqG9_0),.clk(gclk));
	jdff dff_A_34ICDyzh5_0(.dout(w_dff_A_Qp4jWFqG9_0),.din(w_dff_A_34ICDyzh5_0),.clk(gclk));
	jdff dff_A_VV5haM3s3_0(.dout(w_dff_A_34ICDyzh5_0),.din(w_dff_A_VV5haM3s3_0),.clk(gclk));
	jdff dff_A_Ab4P2APt8_0(.dout(w_dff_A_VV5haM3s3_0),.din(w_dff_A_Ab4P2APt8_0),.clk(gclk));
	jdff dff_A_A7qlV5fJ8_0(.dout(w_dff_A_Ab4P2APt8_0),.din(w_dff_A_A7qlV5fJ8_0),.clk(gclk));
	jdff dff_A_9NQH1Hck0_0(.dout(w_dff_A_A7qlV5fJ8_0),.din(w_dff_A_9NQH1Hck0_0),.clk(gclk));
	jdff dff_A_Z3uEeiyT6_0(.dout(w_dff_A_9NQH1Hck0_0),.din(w_dff_A_Z3uEeiyT6_0),.clk(gclk));
	jdff dff_A_mWdRIALO2_0(.dout(w_dff_A_Z3uEeiyT6_0),.din(w_dff_A_mWdRIALO2_0),.clk(gclk));
	jdff dff_A_r95HNJHx4_0(.dout(w_dff_A_mWdRIALO2_0),.din(w_dff_A_r95HNJHx4_0),.clk(gclk));
	jdff dff_A_f6h1wyU90_0(.dout(w_dff_A_r95HNJHx4_0),.din(w_dff_A_f6h1wyU90_0),.clk(gclk));
	jdff dff_A_Mw4tBpp83_0(.dout(w_n255_0[0]),.din(w_dff_A_Mw4tBpp83_0),.clk(gclk));
	jdff dff_B_v4dJJxTg5_1(.din(n220),.dout(w_dff_B_v4dJJxTg5_1),.clk(gclk));
	jdff dff_A_v9ROwN3l1_0(.dout(w_n176_0[0]),.din(w_dff_A_v9ROwN3l1_0),.clk(gclk));
	jdff dff_A_mlbnknNB5_0(.dout(w_dff_A_v9ROwN3l1_0),.din(w_dff_A_mlbnknNB5_0),.clk(gclk));
	jdff dff_A_KHpYXwe94_0(.dout(w_dff_A_mlbnknNB5_0),.din(w_dff_A_KHpYXwe94_0),.clk(gclk));
	jdff dff_A_lc5GsPDE2_0(.dout(w_dff_A_KHpYXwe94_0),.din(w_dff_A_lc5GsPDE2_0),.clk(gclk));
	jdff dff_A_Ax4HIcq91_0(.dout(w_dff_A_lc5GsPDE2_0),.din(w_dff_A_Ax4HIcq91_0),.clk(gclk));
	jdff dff_A_djrQjCzI8_0(.dout(w_dff_A_Ax4HIcq91_0),.din(w_dff_A_djrQjCzI8_0),.clk(gclk));
	jdff dff_A_sJ0SeAbj8_0(.dout(w_dff_A_djrQjCzI8_0),.din(w_dff_A_sJ0SeAbj8_0),.clk(gclk));
	jdff dff_A_fQALokLp6_0(.dout(w_dff_A_sJ0SeAbj8_0),.din(w_dff_A_fQALokLp6_0),.clk(gclk));
	jdff dff_A_FF16szPC6_0(.dout(w_dff_A_fQALokLp6_0),.din(w_dff_A_FF16szPC6_0),.clk(gclk));
	jdff dff_A_lbjjzWXB8_0(.dout(w_dff_A_FF16szPC6_0),.din(w_dff_A_lbjjzWXB8_0),.clk(gclk));
	jdff dff_A_otSeZaLP2_0(.dout(w_dff_A_lbjjzWXB8_0),.din(w_dff_A_otSeZaLP2_0),.clk(gclk));
	jdff dff_A_M4KJUkD10_0(.dout(w_dff_A_otSeZaLP2_0),.din(w_dff_A_M4KJUkD10_0),.clk(gclk));
	jdff dff_A_NRNMucvL8_0(.dout(w_dff_A_M4KJUkD10_0),.din(w_dff_A_NRNMucvL8_0),.clk(gclk));
	jdff dff_A_w4z6xIvG0_0(.dout(w_n206_0[0]),.din(w_dff_A_w4z6xIvG0_0),.clk(gclk));
	jdff dff_B_P5uHvnYR7_1(.din(n178),.dout(w_dff_B_P5uHvnYR7_1),.clk(gclk));
	jdff dff_A_9H74tyFG1_0(.dout(w_n141_0[0]),.din(w_dff_A_9H74tyFG1_0),.clk(gclk));
	jdff dff_A_vMII5KeB2_0(.dout(w_dff_A_9H74tyFG1_0),.din(w_dff_A_vMII5KeB2_0),.clk(gclk));
	jdff dff_A_JYeQomv10_0(.dout(w_dff_A_vMII5KeB2_0),.din(w_dff_A_JYeQomv10_0),.clk(gclk));
	jdff dff_A_kDfU426D9_0(.dout(w_dff_A_JYeQomv10_0),.din(w_dff_A_kDfU426D9_0),.clk(gclk));
	jdff dff_A_onCYGSyy7_0(.dout(w_dff_A_kDfU426D9_0),.din(w_dff_A_onCYGSyy7_0),.clk(gclk));
	jdff dff_A_Tr4czpk28_0(.dout(w_dff_A_onCYGSyy7_0),.din(w_dff_A_Tr4czpk28_0),.clk(gclk));
	jdff dff_A_HXgL8b5L6_0(.dout(w_dff_A_Tr4czpk28_0),.din(w_dff_A_HXgL8b5L6_0),.clk(gclk));
	jdff dff_A_8u86IOad2_0(.dout(w_dff_A_HXgL8b5L6_0),.din(w_dff_A_8u86IOad2_0),.clk(gclk));
	jdff dff_A_Oi0d4Ul72_0(.dout(w_dff_A_8u86IOad2_0),.din(w_dff_A_Oi0d4Ul72_0),.clk(gclk));
	jdff dff_A_cKR98tgH2_0(.dout(w_dff_A_Oi0d4Ul72_0),.din(w_dff_A_cKR98tgH2_0),.clk(gclk));
	jdff dff_A_kFA4SIdY6_0(.dout(w_n164_0[0]),.din(w_dff_A_kFA4SIdY6_0),.clk(gclk));
	jdff dff_B_rLkhshyZ4_1(.din(n143),.dout(w_dff_B_rLkhshyZ4_1),.clk(gclk));
	jdff dff_A_w7t3SQ1H9_0(.dout(w_n112_0[0]),.din(w_dff_A_w7t3SQ1H9_0),.clk(gclk));
	jdff dff_A_j4jcI51m9_0(.dout(w_dff_A_w7t3SQ1H9_0),.din(w_dff_A_j4jcI51m9_0),.clk(gclk));
	jdff dff_A_ATAEXh6Y4_0(.dout(w_dff_A_j4jcI51m9_0),.din(w_dff_A_ATAEXh6Y4_0),.clk(gclk));
	jdff dff_A_iQIRmVPF3_0(.dout(w_dff_A_ATAEXh6Y4_0),.din(w_dff_A_iQIRmVPF3_0),.clk(gclk));
	jdff dff_A_MDiL3YUI2_0(.dout(w_dff_A_iQIRmVPF3_0),.din(w_dff_A_MDiL3YUI2_0),.clk(gclk));
	jdff dff_A_xgwL2N8j9_0(.dout(w_dff_A_MDiL3YUI2_0),.din(w_dff_A_xgwL2N8j9_0),.clk(gclk));
	jdff dff_A_7Mzcdqd21_0(.dout(w_dff_A_xgwL2N8j9_0),.din(w_dff_A_7Mzcdqd21_0),.clk(gclk));
	jdff dff_A_HGFBKBQc8_0(.dout(w_n129_0[0]),.din(w_dff_A_HGFBKBQc8_0),.clk(gclk));
	jdff dff_B_aDyFGiMl4_1(.din(n114),.dout(w_dff_B_aDyFGiMl4_1),.clk(gclk));
	jdff dff_A_XbFi8tcJ8_0(.dout(w_n91_0[0]),.din(w_dff_A_XbFi8tcJ8_0),.clk(gclk));
	jdff dff_A_KOTv3AcU0_0(.dout(w_dff_A_XbFi8tcJ8_0),.din(w_dff_A_KOTv3AcU0_0),.clk(gclk));
	jdff dff_A_wwS2XDmP7_0(.dout(w_dff_A_KOTv3AcU0_0),.din(w_dff_A_wwS2XDmP7_0),.clk(gclk));
	jdff dff_A_LooSY29h1_0(.dout(w_dff_A_wwS2XDmP7_0),.din(w_dff_A_LooSY29h1_0),.clk(gclk));
	jdff dff_B_pauhNMKf4_0(.din(n100),.dout(w_dff_B_pauhNMKf4_0),.clk(gclk));
	jdff dff_A_4Cr04xW87_0(.dout(w_n80_0[0]),.din(w_dff_A_4Cr04xW87_0),.clk(gclk));
	jdff dff_A_oD3ElxP60_0(.dout(w_n1119_0[0]),.din(w_dff_A_oD3ElxP60_0),.clk(gclk));
	jdff dff_B_Bbcq3lRP1_2(.din(n1119),.dout(w_dff_B_Bbcq3lRP1_2),.clk(gclk));
	jdff dff_B_LgYTS43i4_2(.din(n1018),.dout(w_dff_B_LgYTS43i4_2),.clk(gclk));
	jdff dff_B_Oudw9POv2_2(.din(w_dff_B_LgYTS43i4_2),.dout(w_dff_B_Oudw9POv2_2),.clk(gclk));
	jdff dff_B_eJ0cDlGA4_2(.din(w_dff_B_Oudw9POv2_2),.dout(w_dff_B_eJ0cDlGA4_2),.clk(gclk));
	jdff dff_B_C2Pngclt1_2(.din(w_dff_B_eJ0cDlGA4_2),.dout(w_dff_B_C2Pngclt1_2),.clk(gclk));
	jdff dff_B_g2nK8mFz5_2(.din(w_dff_B_C2Pngclt1_2),.dout(w_dff_B_g2nK8mFz5_2),.clk(gclk));
	jdff dff_B_xvgwsWYY3_2(.din(w_dff_B_g2nK8mFz5_2),.dout(w_dff_B_xvgwsWYY3_2),.clk(gclk));
	jdff dff_B_9BlIUzYT6_2(.din(w_dff_B_xvgwsWYY3_2),.dout(w_dff_B_9BlIUzYT6_2),.clk(gclk));
	jdff dff_B_UzWkzLDJ2_2(.din(w_dff_B_9BlIUzYT6_2),.dout(w_dff_B_UzWkzLDJ2_2),.clk(gclk));
	jdff dff_B_Zden3azW1_2(.din(w_dff_B_UzWkzLDJ2_2),.dout(w_dff_B_Zden3azW1_2),.clk(gclk));
	jdff dff_B_Xcp1Kz0p2_2(.din(w_dff_B_Zden3azW1_2),.dout(w_dff_B_Xcp1Kz0p2_2),.clk(gclk));
	jdff dff_B_ade9fVKS7_2(.din(w_dff_B_Xcp1Kz0p2_2),.dout(w_dff_B_ade9fVKS7_2),.clk(gclk));
	jdff dff_B_BmnmFuhG8_2(.din(w_dff_B_ade9fVKS7_2),.dout(w_dff_B_BmnmFuhG8_2),.clk(gclk));
	jdff dff_B_ngd7ZRpQ2_2(.din(w_dff_B_BmnmFuhG8_2),.dout(w_dff_B_ngd7ZRpQ2_2),.clk(gclk));
	jdff dff_B_ZmYg8W020_2(.din(w_dff_B_ngd7ZRpQ2_2),.dout(w_dff_B_ZmYg8W020_2),.clk(gclk));
	jdff dff_B_BUex7L529_2(.din(w_dff_B_ZmYg8W020_2),.dout(w_dff_B_BUex7L529_2),.clk(gclk));
	jdff dff_B_JawP3uC30_2(.din(w_dff_B_BUex7L529_2),.dout(w_dff_B_JawP3uC30_2),.clk(gclk));
	jdff dff_B_fH8IqvuM7_2(.din(w_dff_B_JawP3uC30_2),.dout(w_dff_B_fH8IqvuM7_2),.clk(gclk));
	jdff dff_B_WbbQwUMv3_2(.din(w_dff_B_fH8IqvuM7_2),.dout(w_dff_B_WbbQwUMv3_2),.clk(gclk));
	jdff dff_B_p5Bv42Nr6_2(.din(w_dff_B_WbbQwUMv3_2),.dout(w_dff_B_p5Bv42Nr6_2),.clk(gclk));
	jdff dff_B_ycjaokEY0_2(.din(w_dff_B_p5Bv42Nr6_2),.dout(w_dff_B_ycjaokEY0_2),.clk(gclk));
	jdff dff_B_AOo7R1Bh7_2(.din(w_dff_B_ycjaokEY0_2),.dout(w_dff_B_AOo7R1Bh7_2),.clk(gclk));
	jdff dff_B_gQDPjm2r9_2(.din(w_dff_B_AOo7R1Bh7_2),.dout(w_dff_B_gQDPjm2r9_2),.clk(gclk));
	jdff dff_B_HzEGZ5AM3_2(.din(w_dff_B_gQDPjm2r9_2),.dout(w_dff_B_HzEGZ5AM3_2),.clk(gclk));
	jdff dff_B_YSkcUHKH6_2(.din(w_dff_B_HzEGZ5AM3_2),.dout(w_dff_B_YSkcUHKH6_2),.clk(gclk));
	jdff dff_B_Z7Ma2Q4C4_2(.din(w_dff_B_YSkcUHKH6_2),.dout(w_dff_B_Z7Ma2Q4C4_2),.clk(gclk));
	jdff dff_B_vKFnm0kb2_2(.din(w_dff_B_Z7Ma2Q4C4_2),.dout(w_dff_B_vKFnm0kb2_2),.clk(gclk));
	jdff dff_B_jNXF6eTv5_2(.din(w_dff_B_vKFnm0kb2_2),.dout(w_dff_B_jNXF6eTv5_2),.clk(gclk));
	jdff dff_B_8ojo4nA36_2(.din(w_dff_B_jNXF6eTv5_2),.dout(w_dff_B_8ojo4nA36_2),.clk(gclk));
	jdff dff_B_HbRJAvVw6_2(.din(w_dff_B_8ojo4nA36_2),.dout(w_dff_B_HbRJAvVw6_2),.clk(gclk));
	jdff dff_B_mm3RPkfR6_2(.din(w_dff_B_HbRJAvVw6_2),.dout(w_dff_B_mm3RPkfR6_2),.clk(gclk));
	jdff dff_B_pEPvXgTw1_2(.din(w_dff_B_mm3RPkfR6_2),.dout(w_dff_B_pEPvXgTw1_2),.clk(gclk));
	jdff dff_B_gC6cCtvb2_2(.din(w_dff_B_pEPvXgTw1_2),.dout(w_dff_B_gC6cCtvb2_2),.clk(gclk));
	jdff dff_B_gEA4SDhR6_2(.din(w_dff_B_gC6cCtvb2_2),.dout(w_dff_B_gEA4SDhR6_2),.clk(gclk));
	jdff dff_B_iwPS3qqy2_2(.din(w_dff_B_gEA4SDhR6_2),.dout(w_dff_B_iwPS3qqy2_2),.clk(gclk));
	jdff dff_B_qPYFRTc24_2(.din(w_dff_B_iwPS3qqy2_2),.dout(w_dff_B_qPYFRTc24_2),.clk(gclk));
	jdff dff_B_gPyMBkQI4_2(.din(w_dff_B_qPYFRTc24_2),.dout(w_dff_B_gPyMBkQI4_2),.clk(gclk));
	jdff dff_B_c3u4iLAr3_2(.din(w_dff_B_gPyMBkQI4_2),.dout(w_dff_B_c3u4iLAr3_2),.clk(gclk));
	jdff dff_B_y6dDS9im9_2(.din(w_dff_B_c3u4iLAr3_2),.dout(w_dff_B_y6dDS9im9_2),.clk(gclk));
	jdff dff_B_ZQB8hzz96_2(.din(w_dff_B_y6dDS9im9_2),.dout(w_dff_B_ZQB8hzz96_2),.clk(gclk));
	jdff dff_B_IeLlsolF9_2(.din(w_dff_B_ZQB8hzz96_2),.dout(w_dff_B_IeLlsolF9_2),.clk(gclk));
	jdff dff_B_qV3ZJGDP6_2(.din(w_dff_B_IeLlsolF9_2),.dout(w_dff_B_qV3ZJGDP6_2),.clk(gclk));
	jdff dff_B_wn7iVQvM7_2(.din(w_dff_B_qV3ZJGDP6_2),.dout(w_dff_B_wn7iVQvM7_2),.clk(gclk));
	jdff dff_B_GkYwjBE79_2(.din(w_dff_B_wn7iVQvM7_2),.dout(w_dff_B_GkYwjBE79_2),.clk(gclk));
	jdff dff_A_pgxmyIZO4_0(.dout(w_n1022_0[0]),.din(w_dff_A_pgxmyIZO4_0),.clk(gclk));
	jdff dff_B_AwXEy4nt7_1(.din(n1020),.dout(w_dff_B_AwXEy4nt7_1),.clk(gclk));
	jdff dff_B_8BpXqk955_2(.din(n916),.dout(w_dff_B_8BpXqk955_2),.clk(gclk));
	jdff dff_B_5kaMtNpR5_2(.din(w_dff_B_8BpXqk955_2),.dout(w_dff_B_5kaMtNpR5_2),.clk(gclk));
	jdff dff_B_MsUm0t9m3_2(.din(w_dff_B_5kaMtNpR5_2),.dout(w_dff_B_MsUm0t9m3_2),.clk(gclk));
	jdff dff_B_30dGTRy01_2(.din(w_dff_B_MsUm0t9m3_2),.dout(w_dff_B_30dGTRy01_2),.clk(gclk));
	jdff dff_B_Gfa33qcr6_2(.din(w_dff_B_30dGTRy01_2),.dout(w_dff_B_Gfa33qcr6_2),.clk(gclk));
	jdff dff_B_7zo4x7nJ8_2(.din(w_dff_B_Gfa33qcr6_2),.dout(w_dff_B_7zo4x7nJ8_2),.clk(gclk));
	jdff dff_B_QHDRsdIK2_2(.din(w_dff_B_7zo4x7nJ8_2),.dout(w_dff_B_QHDRsdIK2_2),.clk(gclk));
	jdff dff_B_GV2dQea63_2(.din(w_dff_B_QHDRsdIK2_2),.dout(w_dff_B_GV2dQea63_2),.clk(gclk));
	jdff dff_B_zK2pMWOU6_2(.din(w_dff_B_GV2dQea63_2),.dout(w_dff_B_zK2pMWOU6_2),.clk(gclk));
	jdff dff_B_7jGyAMrY9_2(.din(w_dff_B_zK2pMWOU6_2),.dout(w_dff_B_7jGyAMrY9_2),.clk(gclk));
	jdff dff_B_0OKoFKiV5_2(.din(w_dff_B_7jGyAMrY9_2),.dout(w_dff_B_0OKoFKiV5_2),.clk(gclk));
	jdff dff_B_0B0WJbEs4_2(.din(w_dff_B_0OKoFKiV5_2),.dout(w_dff_B_0B0WJbEs4_2),.clk(gclk));
	jdff dff_B_x7uCCsQu0_2(.din(w_dff_B_0B0WJbEs4_2),.dout(w_dff_B_x7uCCsQu0_2),.clk(gclk));
	jdff dff_B_mGWQHK8e9_2(.din(w_dff_B_x7uCCsQu0_2),.dout(w_dff_B_mGWQHK8e9_2),.clk(gclk));
	jdff dff_B_CimIGaKH5_2(.din(w_dff_B_mGWQHK8e9_2),.dout(w_dff_B_CimIGaKH5_2),.clk(gclk));
	jdff dff_B_bA1fIJzC5_2(.din(w_dff_B_CimIGaKH5_2),.dout(w_dff_B_bA1fIJzC5_2),.clk(gclk));
	jdff dff_B_Kl2EFHPx5_2(.din(w_dff_B_bA1fIJzC5_2),.dout(w_dff_B_Kl2EFHPx5_2),.clk(gclk));
	jdff dff_B_DPDyPAtr7_2(.din(w_dff_B_Kl2EFHPx5_2),.dout(w_dff_B_DPDyPAtr7_2),.clk(gclk));
	jdff dff_B_V0FEB6WK2_2(.din(w_dff_B_DPDyPAtr7_2),.dout(w_dff_B_V0FEB6WK2_2),.clk(gclk));
	jdff dff_B_CntoOaCF0_2(.din(w_dff_B_V0FEB6WK2_2),.dout(w_dff_B_CntoOaCF0_2),.clk(gclk));
	jdff dff_B_eB6f7E5r4_2(.din(w_dff_B_CntoOaCF0_2),.dout(w_dff_B_eB6f7E5r4_2),.clk(gclk));
	jdff dff_B_LY4MKY2l8_2(.din(w_dff_B_eB6f7E5r4_2),.dout(w_dff_B_LY4MKY2l8_2),.clk(gclk));
	jdff dff_B_TVejp6KR9_2(.din(w_dff_B_LY4MKY2l8_2),.dout(w_dff_B_TVejp6KR9_2),.clk(gclk));
	jdff dff_B_bE8Emp6j3_2(.din(w_dff_B_TVejp6KR9_2),.dout(w_dff_B_bE8Emp6j3_2),.clk(gclk));
	jdff dff_B_KKlKOssP8_2(.din(w_dff_B_bE8Emp6j3_2),.dout(w_dff_B_KKlKOssP8_2),.clk(gclk));
	jdff dff_B_b3jzkhOZ3_2(.din(w_dff_B_KKlKOssP8_2),.dout(w_dff_B_b3jzkhOZ3_2),.clk(gclk));
	jdff dff_B_nRt4USLP4_2(.din(w_dff_B_b3jzkhOZ3_2),.dout(w_dff_B_nRt4USLP4_2),.clk(gclk));
	jdff dff_B_Q7O5YwYF0_2(.din(w_dff_B_nRt4USLP4_2),.dout(w_dff_B_Q7O5YwYF0_2),.clk(gclk));
	jdff dff_B_ERabeJf06_2(.din(w_dff_B_Q7O5YwYF0_2),.dout(w_dff_B_ERabeJf06_2),.clk(gclk));
	jdff dff_B_Gq7D5bBI7_2(.din(w_dff_B_ERabeJf06_2),.dout(w_dff_B_Gq7D5bBI7_2),.clk(gclk));
	jdff dff_B_voqTkvNb5_2(.din(w_dff_B_Gq7D5bBI7_2),.dout(w_dff_B_voqTkvNb5_2),.clk(gclk));
	jdff dff_B_jRDmwexT9_2(.din(w_dff_B_voqTkvNb5_2),.dout(w_dff_B_jRDmwexT9_2),.clk(gclk));
	jdff dff_B_TeHlzT608_2(.din(w_dff_B_jRDmwexT9_2),.dout(w_dff_B_TeHlzT608_2),.clk(gclk));
	jdff dff_B_tlyYCVOv9_2(.din(w_dff_B_TeHlzT608_2),.dout(w_dff_B_tlyYCVOv9_2),.clk(gclk));
	jdff dff_B_OofZ6gfh7_2(.din(w_dff_B_tlyYCVOv9_2),.dout(w_dff_B_OofZ6gfh7_2),.clk(gclk));
	jdff dff_B_B9TVCtWm2_2(.din(w_dff_B_OofZ6gfh7_2),.dout(w_dff_B_B9TVCtWm2_2),.clk(gclk));
	jdff dff_B_qTjXRTk78_2(.din(w_dff_B_B9TVCtWm2_2),.dout(w_dff_B_qTjXRTk78_2),.clk(gclk));
	jdff dff_B_51vgnAj54_2(.din(w_dff_B_qTjXRTk78_2),.dout(w_dff_B_51vgnAj54_2),.clk(gclk));
	jdff dff_B_RB89K6Gk5_2(.din(w_dff_B_51vgnAj54_2),.dout(w_dff_B_RB89K6Gk5_2),.clk(gclk));
	jdff dff_B_sNYQT0OB0_2(.din(w_dff_B_RB89K6Gk5_2),.dout(w_dff_B_sNYQT0OB0_2),.clk(gclk));
	jdff dff_A_Ig2IiMIV7_1(.dout(w_n1006_0[1]),.din(w_dff_A_Ig2IiMIV7_1),.clk(gclk));
	jdff dff_A_S9PIOujp5_0(.dout(w_n816_0[0]),.din(w_dff_A_S9PIOujp5_0),.clk(gclk));
	jdff dff_A_xnh2ICtZ4_0(.dout(w_dff_A_S9PIOujp5_0),.din(w_dff_A_xnh2ICtZ4_0),.clk(gclk));
	jdff dff_A_O9TlwrpB7_0(.dout(w_dff_A_xnh2ICtZ4_0),.din(w_dff_A_O9TlwrpB7_0),.clk(gclk));
	jdff dff_A_6awEeOUm7_0(.dout(w_dff_A_O9TlwrpB7_0),.din(w_dff_A_6awEeOUm7_0),.clk(gclk));
	jdff dff_A_c7uzayFU0_0(.dout(w_dff_A_6awEeOUm7_0),.din(w_dff_A_c7uzayFU0_0),.clk(gclk));
	jdff dff_A_AcJlvA2K6_0(.dout(w_dff_A_c7uzayFU0_0),.din(w_dff_A_AcJlvA2K6_0),.clk(gclk));
	jdff dff_A_tVpkZpNI1_0(.dout(w_dff_A_AcJlvA2K6_0),.din(w_dff_A_tVpkZpNI1_0),.clk(gclk));
	jdff dff_A_ltnxb5vx3_0(.dout(w_dff_A_tVpkZpNI1_0),.din(w_dff_A_ltnxb5vx3_0),.clk(gclk));
	jdff dff_A_2qeuCHrk9_0(.dout(w_dff_A_ltnxb5vx3_0),.din(w_dff_A_2qeuCHrk9_0),.clk(gclk));
	jdff dff_A_LxDgNnRa1_0(.dout(w_dff_A_2qeuCHrk9_0),.din(w_dff_A_LxDgNnRa1_0),.clk(gclk));
	jdff dff_A_HUxE6ItK3_0(.dout(w_dff_A_LxDgNnRa1_0),.din(w_dff_A_HUxE6ItK3_0),.clk(gclk));
	jdff dff_A_RUPJUt0V3_0(.dout(w_dff_A_HUxE6ItK3_0),.din(w_dff_A_RUPJUt0V3_0),.clk(gclk));
	jdff dff_A_XwqwnjGT3_0(.dout(w_dff_A_RUPJUt0V3_0),.din(w_dff_A_XwqwnjGT3_0),.clk(gclk));
	jdff dff_A_wyX1GCcq5_0(.dout(w_dff_A_XwqwnjGT3_0),.din(w_dff_A_wyX1GCcq5_0),.clk(gclk));
	jdff dff_A_mWlAdXdo8_0(.dout(w_dff_A_wyX1GCcq5_0),.din(w_dff_A_mWlAdXdo8_0),.clk(gclk));
	jdff dff_A_QWUW1Qou1_0(.dout(w_dff_A_mWlAdXdo8_0),.din(w_dff_A_QWUW1Qou1_0),.clk(gclk));
	jdff dff_A_IRijIAHQ0_0(.dout(w_dff_A_QWUW1Qou1_0),.din(w_dff_A_IRijIAHQ0_0),.clk(gclk));
	jdff dff_A_4acfb7WY5_0(.dout(w_dff_A_IRijIAHQ0_0),.din(w_dff_A_4acfb7WY5_0),.clk(gclk));
	jdff dff_A_VjGgXz3y1_0(.dout(w_dff_A_4acfb7WY5_0),.din(w_dff_A_VjGgXz3y1_0),.clk(gclk));
	jdff dff_A_5wSlEO0x5_0(.dout(w_dff_A_VjGgXz3y1_0),.din(w_dff_A_5wSlEO0x5_0),.clk(gclk));
	jdff dff_A_YloFWHmu7_0(.dout(w_dff_A_5wSlEO0x5_0),.din(w_dff_A_YloFWHmu7_0),.clk(gclk));
	jdff dff_A_HgqSJjSE2_0(.dout(w_dff_A_YloFWHmu7_0),.din(w_dff_A_HgqSJjSE2_0),.clk(gclk));
	jdff dff_A_M17ZIlp44_0(.dout(w_dff_A_HgqSJjSE2_0),.din(w_dff_A_M17ZIlp44_0),.clk(gclk));
	jdff dff_A_wi1I0ai18_0(.dout(w_dff_A_M17ZIlp44_0),.din(w_dff_A_wi1I0ai18_0),.clk(gclk));
	jdff dff_A_qN1KMaIG3_0(.dout(w_dff_A_wi1I0ai18_0),.din(w_dff_A_qN1KMaIG3_0),.clk(gclk));
	jdff dff_A_JKcFQTYX3_0(.dout(w_dff_A_qN1KMaIG3_0),.din(w_dff_A_JKcFQTYX3_0),.clk(gclk));
	jdff dff_A_7WdnC1v71_0(.dout(w_dff_A_JKcFQTYX3_0),.din(w_dff_A_7WdnC1v71_0),.clk(gclk));
	jdff dff_A_IndqoNG13_0(.dout(w_dff_A_7WdnC1v71_0),.din(w_dff_A_IndqoNG13_0),.clk(gclk));
	jdff dff_A_fC8iFi6T1_0(.dout(w_dff_A_IndqoNG13_0),.din(w_dff_A_fC8iFi6T1_0),.clk(gclk));
	jdff dff_A_WRQh3zLS5_0(.dout(w_dff_A_fC8iFi6T1_0),.din(w_dff_A_WRQh3zLS5_0),.clk(gclk));
	jdff dff_A_IsSXWxk38_0(.dout(w_dff_A_WRQh3zLS5_0),.din(w_dff_A_IsSXWxk38_0),.clk(gclk));
	jdff dff_A_mWoYxURw9_0(.dout(w_dff_A_IsSXWxk38_0),.din(w_dff_A_mWoYxURw9_0),.clk(gclk));
	jdff dff_A_Muh60JkR9_0(.dout(w_dff_A_mWoYxURw9_0),.din(w_dff_A_Muh60JkR9_0),.clk(gclk));
	jdff dff_A_G9VXaPrw3_0(.dout(w_dff_A_Muh60JkR9_0),.din(w_dff_A_G9VXaPrw3_0),.clk(gclk));
	jdff dff_A_xVDWveXm4_0(.dout(w_dff_A_G9VXaPrw3_0),.din(w_dff_A_xVDWveXm4_0),.clk(gclk));
	jdff dff_A_CWzR1lEv6_0(.dout(w_dff_A_xVDWveXm4_0),.din(w_dff_A_CWzR1lEv6_0),.clk(gclk));
	jdff dff_A_0TE8lFqx1_0(.dout(w_dff_A_CWzR1lEv6_0),.din(w_dff_A_0TE8lFqx1_0),.clk(gclk));
	jdff dff_A_l6lgNt926_1(.dout(w_n900_0[1]),.din(w_dff_A_l6lgNt926_1),.clk(gclk));
	jdff dff_A_fTqCUQNZ9_2(.dout(w_n900_0[2]),.din(w_dff_A_fTqCUQNZ9_2),.clk(gclk));
	jdff dff_B_tjlHIzTL2_1(.din(n818),.dout(w_dff_B_tjlHIzTL2_1),.clk(gclk));
	jdff dff_B_hVtGoqtw7_2(.din(n719),.dout(w_dff_B_hVtGoqtw7_2),.clk(gclk));
	jdff dff_B_BGyenYGj6_2(.din(w_dff_B_hVtGoqtw7_2),.dout(w_dff_B_BGyenYGj6_2),.clk(gclk));
	jdff dff_B_w4Lkn5jg6_2(.din(w_dff_B_BGyenYGj6_2),.dout(w_dff_B_w4Lkn5jg6_2),.clk(gclk));
	jdff dff_B_j9RLxeHL3_2(.din(w_dff_B_w4Lkn5jg6_2),.dout(w_dff_B_j9RLxeHL3_2),.clk(gclk));
	jdff dff_B_HTSAbvKw5_2(.din(w_dff_B_j9RLxeHL3_2),.dout(w_dff_B_HTSAbvKw5_2),.clk(gclk));
	jdff dff_B_yFLPmvyQ9_2(.din(w_dff_B_HTSAbvKw5_2),.dout(w_dff_B_yFLPmvyQ9_2),.clk(gclk));
	jdff dff_B_yuqETpIQ5_2(.din(w_dff_B_yFLPmvyQ9_2),.dout(w_dff_B_yuqETpIQ5_2),.clk(gclk));
	jdff dff_B_C1xYgUPO6_2(.din(w_dff_B_yuqETpIQ5_2),.dout(w_dff_B_C1xYgUPO6_2),.clk(gclk));
	jdff dff_B_YnJXQg3j4_2(.din(w_dff_B_C1xYgUPO6_2),.dout(w_dff_B_YnJXQg3j4_2),.clk(gclk));
	jdff dff_B_VIqON7Z05_2(.din(w_dff_B_YnJXQg3j4_2),.dout(w_dff_B_VIqON7Z05_2),.clk(gclk));
	jdff dff_B_72fmwJ2L9_2(.din(w_dff_B_VIqON7Z05_2),.dout(w_dff_B_72fmwJ2L9_2),.clk(gclk));
	jdff dff_B_uNoHPmd20_2(.din(w_dff_B_72fmwJ2L9_2),.dout(w_dff_B_uNoHPmd20_2),.clk(gclk));
	jdff dff_B_kZB5kuyT4_2(.din(w_dff_B_uNoHPmd20_2),.dout(w_dff_B_kZB5kuyT4_2),.clk(gclk));
	jdff dff_B_uoAmyg234_2(.din(w_dff_B_kZB5kuyT4_2),.dout(w_dff_B_uoAmyg234_2),.clk(gclk));
	jdff dff_B_StdMDfwz9_2(.din(w_dff_B_uoAmyg234_2),.dout(w_dff_B_StdMDfwz9_2),.clk(gclk));
	jdff dff_B_owRQFHUV4_2(.din(w_dff_B_StdMDfwz9_2),.dout(w_dff_B_owRQFHUV4_2),.clk(gclk));
	jdff dff_B_ubmCFz354_2(.din(w_dff_B_owRQFHUV4_2),.dout(w_dff_B_ubmCFz354_2),.clk(gclk));
	jdff dff_B_ltVpqtfV1_2(.din(w_dff_B_ubmCFz354_2),.dout(w_dff_B_ltVpqtfV1_2),.clk(gclk));
	jdff dff_B_HojszjWL1_2(.din(w_dff_B_ltVpqtfV1_2),.dout(w_dff_B_HojszjWL1_2),.clk(gclk));
	jdff dff_B_VPB3AA0m8_2(.din(w_dff_B_HojszjWL1_2),.dout(w_dff_B_VPB3AA0m8_2),.clk(gclk));
	jdff dff_B_0AF2VxD82_2(.din(w_dff_B_VPB3AA0m8_2),.dout(w_dff_B_0AF2VxD82_2),.clk(gclk));
	jdff dff_B_OI6G4csf5_2(.din(w_dff_B_0AF2VxD82_2),.dout(w_dff_B_OI6G4csf5_2),.clk(gclk));
	jdff dff_B_qP1jrZuS9_2(.din(w_dff_B_OI6G4csf5_2),.dout(w_dff_B_qP1jrZuS9_2),.clk(gclk));
	jdff dff_B_jT2368OV1_2(.din(w_dff_B_qP1jrZuS9_2),.dout(w_dff_B_jT2368OV1_2),.clk(gclk));
	jdff dff_B_SvrTqzrS7_2(.din(w_dff_B_jT2368OV1_2),.dout(w_dff_B_SvrTqzrS7_2),.clk(gclk));
	jdff dff_B_uyGJBh3X2_2(.din(w_dff_B_SvrTqzrS7_2),.dout(w_dff_B_uyGJBh3X2_2),.clk(gclk));
	jdff dff_B_mtlYpPd84_2(.din(w_dff_B_uyGJBh3X2_2),.dout(w_dff_B_mtlYpPd84_2),.clk(gclk));
	jdff dff_B_AY7Kt3ua7_2(.din(w_dff_B_mtlYpPd84_2),.dout(w_dff_B_AY7Kt3ua7_2),.clk(gclk));
	jdff dff_B_YGGkpzm89_2(.din(w_dff_B_AY7Kt3ua7_2),.dout(w_dff_B_YGGkpzm89_2),.clk(gclk));
	jdff dff_B_ZAwMDljP6_2(.din(w_dff_B_YGGkpzm89_2),.dout(w_dff_B_ZAwMDljP6_2),.clk(gclk));
	jdff dff_B_IixtpD9V8_2(.din(w_dff_B_ZAwMDljP6_2),.dout(w_dff_B_IixtpD9V8_2),.clk(gclk));
	jdff dff_B_ah4ViFEx7_2(.din(w_dff_B_IixtpD9V8_2),.dout(w_dff_B_ah4ViFEx7_2),.clk(gclk));
	jdff dff_B_iI69Sy724_2(.din(w_dff_B_ah4ViFEx7_2),.dout(w_dff_B_iI69Sy724_2),.clk(gclk));
	jdff dff_B_jkAymBlt3_2(.din(n797),.dout(w_dff_B_jkAymBlt3_2),.clk(gclk));
	jdff dff_B_qWDKSY1J5_1(.din(n720),.dout(w_dff_B_qWDKSY1J5_1),.clk(gclk));
	jdff dff_B_biP9Zti95_2(.din(n627),.dout(w_dff_B_biP9Zti95_2),.clk(gclk));
	jdff dff_B_8C4FMtFD3_2(.din(w_dff_B_biP9Zti95_2),.dout(w_dff_B_8C4FMtFD3_2),.clk(gclk));
	jdff dff_B_VYqPFXeF0_2(.din(w_dff_B_8C4FMtFD3_2),.dout(w_dff_B_VYqPFXeF0_2),.clk(gclk));
	jdff dff_B_4paEbKGf4_2(.din(w_dff_B_VYqPFXeF0_2),.dout(w_dff_B_4paEbKGf4_2),.clk(gclk));
	jdff dff_B_nYpRnQdA2_2(.din(w_dff_B_4paEbKGf4_2),.dout(w_dff_B_nYpRnQdA2_2),.clk(gclk));
	jdff dff_B_z9Of2kY57_2(.din(w_dff_B_nYpRnQdA2_2),.dout(w_dff_B_z9Of2kY57_2),.clk(gclk));
	jdff dff_B_LdOO0mpp1_2(.din(w_dff_B_z9Of2kY57_2),.dout(w_dff_B_LdOO0mpp1_2),.clk(gclk));
	jdff dff_B_GppeaWwv3_2(.din(w_dff_B_LdOO0mpp1_2),.dout(w_dff_B_GppeaWwv3_2),.clk(gclk));
	jdff dff_B_3qosq3h65_2(.din(w_dff_B_GppeaWwv3_2),.dout(w_dff_B_3qosq3h65_2),.clk(gclk));
	jdff dff_B_nGJuWHB58_2(.din(w_dff_B_3qosq3h65_2),.dout(w_dff_B_nGJuWHB58_2),.clk(gclk));
	jdff dff_B_vcSlr4s27_2(.din(w_dff_B_nGJuWHB58_2),.dout(w_dff_B_vcSlr4s27_2),.clk(gclk));
	jdff dff_B_spNi7WVu3_2(.din(w_dff_B_vcSlr4s27_2),.dout(w_dff_B_spNi7WVu3_2),.clk(gclk));
	jdff dff_B_BvjI52qV9_2(.din(w_dff_B_spNi7WVu3_2),.dout(w_dff_B_BvjI52qV9_2),.clk(gclk));
	jdff dff_B_5gXu3jfi7_2(.din(w_dff_B_BvjI52qV9_2),.dout(w_dff_B_5gXu3jfi7_2),.clk(gclk));
	jdff dff_B_MWhU6ZVS7_2(.din(w_dff_B_5gXu3jfi7_2),.dout(w_dff_B_MWhU6ZVS7_2),.clk(gclk));
	jdff dff_B_YLTR9ZYY9_2(.din(w_dff_B_MWhU6ZVS7_2),.dout(w_dff_B_YLTR9ZYY9_2),.clk(gclk));
	jdff dff_B_GeVXzpm79_2(.din(w_dff_B_YLTR9ZYY9_2),.dout(w_dff_B_GeVXzpm79_2),.clk(gclk));
	jdff dff_B_fsAKEm1y8_2(.din(w_dff_B_GeVXzpm79_2),.dout(w_dff_B_fsAKEm1y8_2),.clk(gclk));
	jdff dff_B_bHftqYYi0_2(.din(w_dff_B_fsAKEm1y8_2),.dout(w_dff_B_bHftqYYi0_2),.clk(gclk));
	jdff dff_B_7vAgEoTV1_2(.din(w_dff_B_bHftqYYi0_2),.dout(w_dff_B_7vAgEoTV1_2),.clk(gclk));
	jdff dff_B_ZWw8runF6_2(.din(w_dff_B_7vAgEoTV1_2),.dout(w_dff_B_ZWw8runF6_2),.clk(gclk));
	jdff dff_B_Lmw2EkNw7_2(.din(w_dff_B_ZWw8runF6_2),.dout(w_dff_B_Lmw2EkNw7_2),.clk(gclk));
	jdff dff_B_lI7YnOhd9_2(.din(w_dff_B_Lmw2EkNw7_2),.dout(w_dff_B_lI7YnOhd9_2),.clk(gclk));
	jdff dff_B_UzdgR5uo4_2(.din(w_dff_B_lI7YnOhd9_2),.dout(w_dff_B_UzdgR5uo4_2),.clk(gclk));
	jdff dff_B_7UhaOJkU0_2(.din(w_dff_B_UzdgR5uo4_2),.dout(w_dff_B_7UhaOJkU0_2),.clk(gclk));
	jdff dff_B_0WdFHa4f7_2(.din(w_dff_B_7UhaOJkU0_2),.dout(w_dff_B_0WdFHa4f7_2),.clk(gclk));
	jdff dff_B_ikGBUAgq8_2(.din(w_dff_B_0WdFHa4f7_2),.dout(w_dff_B_ikGBUAgq8_2),.clk(gclk));
	jdff dff_B_YA36SIE08_2(.din(w_dff_B_ikGBUAgq8_2),.dout(w_dff_B_YA36SIE08_2),.clk(gclk));
	jdff dff_B_k5xok1rj4_2(.din(w_dff_B_YA36SIE08_2),.dout(w_dff_B_k5xok1rj4_2),.clk(gclk));
	jdff dff_B_l80K2F2M7_2(.din(w_dff_B_k5xok1rj4_2),.dout(w_dff_B_l80K2F2M7_2),.clk(gclk));
	jdff dff_B_mZTqKZKU0_2(.din(n698),.dout(w_dff_B_mZTqKZKU0_2),.clk(gclk));
	jdff dff_B_3fIFSjOP8_1(.din(n628),.dout(w_dff_B_3fIFSjOP8_1),.clk(gclk));
	jdff dff_B_69YsihiC8_2(.din(n542),.dout(w_dff_B_69YsihiC8_2),.clk(gclk));
	jdff dff_B_WkjculoG2_2(.din(w_dff_B_69YsihiC8_2),.dout(w_dff_B_WkjculoG2_2),.clk(gclk));
	jdff dff_B_9PjHFIgW2_2(.din(w_dff_B_WkjculoG2_2),.dout(w_dff_B_9PjHFIgW2_2),.clk(gclk));
	jdff dff_B_9QVii5Ix8_2(.din(w_dff_B_9PjHFIgW2_2),.dout(w_dff_B_9QVii5Ix8_2),.clk(gclk));
	jdff dff_B_2ZV56b0g1_2(.din(w_dff_B_9QVii5Ix8_2),.dout(w_dff_B_2ZV56b0g1_2),.clk(gclk));
	jdff dff_B_rMiGF1Qi9_2(.din(w_dff_B_2ZV56b0g1_2),.dout(w_dff_B_rMiGF1Qi9_2),.clk(gclk));
	jdff dff_B_XfJFoGPi9_2(.din(w_dff_B_rMiGF1Qi9_2),.dout(w_dff_B_XfJFoGPi9_2),.clk(gclk));
	jdff dff_B_cizMnaxg3_2(.din(w_dff_B_XfJFoGPi9_2),.dout(w_dff_B_cizMnaxg3_2),.clk(gclk));
	jdff dff_B_BDw5m5AH8_2(.din(w_dff_B_cizMnaxg3_2),.dout(w_dff_B_BDw5m5AH8_2),.clk(gclk));
	jdff dff_B_Y12UcpN05_2(.din(w_dff_B_BDw5m5AH8_2),.dout(w_dff_B_Y12UcpN05_2),.clk(gclk));
	jdff dff_B_eaNrTYmG1_2(.din(w_dff_B_Y12UcpN05_2),.dout(w_dff_B_eaNrTYmG1_2),.clk(gclk));
	jdff dff_B_x9n9wSfl5_2(.din(w_dff_B_eaNrTYmG1_2),.dout(w_dff_B_x9n9wSfl5_2),.clk(gclk));
	jdff dff_B_evK23eiy0_2(.din(w_dff_B_x9n9wSfl5_2),.dout(w_dff_B_evK23eiy0_2),.clk(gclk));
	jdff dff_B_jenYlyly2_2(.din(w_dff_B_evK23eiy0_2),.dout(w_dff_B_jenYlyly2_2),.clk(gclk));
	jdff dff_B_IbvcS0SH2_2(.din(w_dff_B_jenYlyly2_2),.dout(w_dff_B_IbvcS0SH2_2),.clk(gclk));
	jdff dff_B_9mRY4NJQ3_2(.din(w_dff_B_IbvcS0SH2_2),.dout(w_dff_B_9mRY4NJQ3_2),.clk(gclk));
	jdff dff_B_cK2bwMb20_2(.din(w_dff_B_9mRY4NJQ3_2),.dout(w_dff_B_cK2bwMb20_2),.clk(gclk));
	jdff dff_B_ucru1cW17_2(.din(w_dff_B_cK2bwMb20_2),.dout(w_dff_B_ucru1cW17_2),.clk(gclk));
	jdff dff_B_S687hQYd4_2(.din(w_dff_B_ucru1cW17_2),.dout(w_dff_B_S687hQYd4_2),.clk(gclk));
	jdff dff_B_09pPRDxc3_2(.din(w_dff_B_S687hQYd4_2),.dout(w_dff_B_09pPRDxc3_2),.clk(gclk));
	jdff dff_B_Io5Mz4PT2_2(.din(w_dff_B_09pPRDxc3_2),.dout(w_dff_B_Io5Mz4PT2_2),.clk(gclk));
	jdff dff_B_rU7fOSqf7_2(.din(w_dff_B_Io5Mz4PT2_2),.dout(w_dff_B_rU7fOSqf7_2),.clk(gclk));
	jdff dff_B_z4azcPV95_2(.din(w_dff_B_rU7fOSqf7_2),.dout(w_dff_B_z4azcPV95_2),.clk(gclk));
	jdff dff_B_RlRmQd2E9_2(.din(w_dff_B_z4azcPV95_2),.dout(w_dff_B_RlRmQd2E9_2),.clk(gclk));
	jdff dff_B_eALBBeqr7_2(.din(w_dff_B_RlRmQd2E9_2),.dout(w_dff_B_eALBBeqr7_2),.clk(gclk));
	jdff dff_B_lscsfo6j1_2(.din(w_dff_B_eALBBeqr7_2),.dout(w_dff_B_lscsfo6j1_2),.clk(gclk));
	jdff dff_B_eR3Wb2sf5_2(.din(w_dff_B_lscsfo6j1_2),.dout(w_dff_B_eR3Wb2sf5_2),.clk(gclk));
	jdff dff_B_Q4Xb684L2_2(.din(n606),.dout(w_dff_B_Q4Xb684L2_2),.clk(gclk));
	jdff dff_B_KtEFl8uK2_1(.din(n543),.dout(w_dff_B_KtEFl8uK2_1),.clk(gclk));
	jdff dff_B_YOHpvLlj5_2(.din(n464),.dout(w_dff_B_YOHpvLlj5_2),.clk(gclk));
	jdff dff_B_c1sW522N2_2(.din(w_dff_B_YOHpvLlj5_2),.dout(w_dff_B_c1sW522N2_2),.clk(gclk));
	jdff dff_B_BXnsZxxL4_2(.din(w_dff_B_c1sW522N2_2),.dout(w_dff_B_BXnsZxxL4_2),.clk(gclk));
	jdff dff_B_HHnhWQfZ6_2(.din(w_dff_B_BXnsZxxL4_2),.dout(w_dff_B_HHnhWQfZ6_2),.clk(gclk));
	jdff dff_B_ZvMJZtFk5_2(.din(w_dff_B_HHnhWQfZ6_2),.dout(w_dff_B_ZvMJZtFk5_2),.clk(gclk));
	jdff dff_B_NfSyGMGu5_2(.din(w_dff_B_ZvMJZtFk5_2),.dout(w_dff_B_NfSyGMGu5_2),.clk(gclk));
	jdff dff_B_NvOE3LZD0_2(.din(w_dff_B_NfSyGMGu5_2),.dout(w_dff_B_NvOE3LZD0_2),.clk(gclk));
	jdff dff_B_vD9iUEHj6_2(.din(w_dff_B_NvOE3LZD0_2),.dout(w_dff_B_vD9iUEHj6_2),.clk(gclk));
	jdff dff_B_RRaTGuhc5_2(.din(w_dff_B_vD9iUEHj6_2),.dout(w_dff_B_RRaTGuhc5_2),.clk(gclk));
	jdff dff_B_VzDQvlwo3_2(.din(w_dff_B_RRaTGuhc5_2),.dout(w_dff_B_VzDQvlwo3_2),.clk(gclk));
	jdff dff_B_uquQkKXu1_2(.din(w_dff_B_VzDQvlwo3_2),.dout(w_dff_B_uquQkKXu1_2),.clk(gclk));
	jdff dff_B_FXeKZdie9_2(.din(w_dff_B_uquQkKXu1_2),.dout(w_dff_B_FXeKZdie9_2),.clk(gclk));
	jdff dff_B_RB7PdyId3_2(.din(w_dff_B_FXeKZdie9_2),.dout(w_dff_B_RB7PdyId3_2),.clk(gclk));
	jdff dff_B_miIF4meo0_2(.din(w_dff_B_RB7PdyId3_2),.dout(w_dff_B_miIF4meo0_2),.clk(gclk));
	jdff dff_B_DsbP680z0_2(.din(w_dff_B_miIF4meo0_2),.dout(w_dff_B_DsbP680z0_2),.clk(gclk));
	jdff dff_B_ZNhsVKBN3_2(.din(w_dff_B_DsbP680z0_2),.dout(w_dff_B_ZNhsVKBN3_2),.clk(gclk));
	jdff dff_B_FMFjZmjJ5_2(.din(w_dff_B_ZNhsVKBN3_2),.dout(w_dff_B_FMFjZmjJ5_2),.clk(gclk));
	jdff dff_B_HkkgOSe64_2(.din(w_dff_B_FMFjZmjJ5_2),.dout(w_dff_B_HkkgOSe64_2),.clk(gclk));
	jdff dff_B_w6Ju8LO91_2(.din(w_dff_B_HkkgOSe64_2),.dout(w_dff_B_w6Ju8LO91_2),.clk(gclk));
	jdff dff_B_RCpJbxQj1_2(.din(w_dff_B_w6Ju8LO91_2),.dout(w_dff_B_RCpJbxQj1_2),.clk(gclk));
	jdff dff_B_djHnKz494_2(.din(w_dff_B_RCpJbxQj1_2),.dout(w_dff_B_djHnKz494_2),.clk(gclk));
	jdff dff_B_VrSQM04q7_2(.din(w_dff_B_djHnKz494_2),.dout(w_dff_B_VrSQM04q7_2),.clk(gclk));
	jdff dff_B_GT6xsgMZ8_2(.din(w_dff_B_VrSQM04q7_2),.dout(w_dff_B_GT6xsgMZ8_2),.clk(gclk));
	jdff dff_B_w7W1k9Hk6_2(.din(w_dff_B_GT6xsgMZ8_2),.dout(w_dff_B_w7W1k9Hk6_2),.clk(gclk));
	jdff dff_B_hZo4AJL16_2(.din(n521),.dout(w_dff_B_hZo4AJL16_2),.clk(gclk));
	jdff dff_B_gOSBDxmP5_1(.din(n465),.dout(w_dff_B_gOSBDxmP5_1),.clk(gclk));
	jdff dff_B_MhdsDXXB8_2(.din(n393),.dout(w_dff_B_MhdsDXXB8_2),.clk(gclk));
	jdff dff_B_fwA2z8ik0_2(.din(w_dff_B_MhdsDXXB8_2),.dout(w_dff_B_fwA2z8ik0_2),.clk(gclk));
	jdff dff_B_IdyDmHs90_2(.din(w_dff_B_fwA2z8ik0_2),.dout(w_dff_B_IdyDmHs90_2),.clk(gclk));
	jdff dff_B_H0cgRTLw6_2(.din(w_dff_B_IdyDmHs90_2),.dout(w_dff_B_H0cgRTLw6_2),.clk(gclk));
	jdff dff_B_WxCVjQDi9_2(.din(w_dff_B_H0cgRTLw6_2),.dout(w_dff_B_WxCVjQDi9_2),.clk(gclk));
	jdff dff_B_MeEwdt0v6_2(.din(w_dff_B_WxCVjQDi9_2),.dout(w_dff_B_MeEwdt0v6_2),.clk(gclk));
	jdff dff_B_DZCKW1Al3_2(.din(w_dff_B_MeEwdt0v6_2),.dout(w_dff_B_DZCKW1Al3_2),.clk(gclk));
	jdff dff_B_MOxIcfym4_2(.din(w_dff_B_DZCKW1Al3_2),.dout(w_dff_B_MOxIcfym4_2),.clk(gclk));
	jdff dff_B_ixAZpz546_2(.din(w_dff_B_MOxIcfym4_2),.dout(w_dff_B_ixAZpz546_2),.clk(gclk));
	jdff dff_B_JJUzFS988_2(.din(w_dff_B_ixAZpz546_2),.dout(w_dff_B_JJUzFS988_2),.clk(gclk));
	jdff dff_B_ld838vVh5_2(.din(w_dff_B_JJUzFS988_2),.dout(w_dff_B_ld838vVh5_2),.clk(gclk));
	jdff dff_B_sxPuUwLJ7_2(.din(w_dff_B_ld838vVh5_2),.dout(w_dff_B_sxPuUwLJ7_2),.clk(gclk));
	jdff dff_B_2YISQFJi4_2(.din(w_dff_B_sxPuUwLJ7_2),.dout(w_dff_B_2YISQFJi4_2),.clk(gclk));
	jdff dff_B_ELL9OwzR6_2(.din(w_dff_B_2YISQFJi4_2),.dout(w_dff_B_ELL9OwzR6_2),.clk(gclk));
	jdff dff_B_0kEpU8ef5_2(.din(w_dff_B_ELL9OwzR6_2),.dout(w_dff_B_0kEpU8ef5_2),.clk(gclk));
	jdff dff_B_eQAYCGik0_2(.din(w_dff_B_0kEpU8ef5_2),.dout(w_dff_B_eQAYCGik0_2),.clk(gclk));
	jdff dff_B_CopEqRwn1_2(.din(w_dff_B_eQAYCGik0_2),.dout(w_dff_B_CopEqRwn1_2),.clk(gclk));
	jdff dff_B_FVzKIRze0_2(.din(w_dff_B_CopEqRwn1_2),.dout(w_dff_B_FVzKIRze0_2),.clk(gclk));
	jdff dff_B_GlvoadhE4_2(.din(w_dff_B_FVzKIRze0_2),.dout(w_dff_B_GlvoadhE4_2),.clk(gclk));
	jdff dff_B_fyXt3Iiz2_2(.din(w_dff_B_GlvoadhE4_2),.dout(w_dff_B_fyXt3Iiz2_2),.clk(gclk));
	jdff dff_B_ZCDYx5Hp6_2(.din(w_dff_B_fyXt3Iiz2_2),.dout(w_dff_B_ZCDYx5Hp6_2),.clk(gclk));
	jdff dff_B_VAUq4dSN9_2(.din(n443),.dout(w_dff_B_VAUq4dSN9_2),.clk(gclk));
	jdff dff_B_elABO3cg9_1(.din(n394),.dout(w_dff_B_elABO3cg9_1),.clk(gclk));
	jdff dff_B_hwLaWcnf6_2(.din(n330),.dout(w_dff_B_hwLaWcnf6_2),.clk(gclk));
	jdff dff_B_qEjWbzPN8_2(.din(w_dff_B_hwLaWcnf6_2),.dout(w_dff_B_qEjWbzPN8_2),.clk(gclk));
	jdff dff_B_2RNSW0dd4_2(.din(w_dff_B_qEjWbzPN8_2),.dout(w_dff_B_2RNSW0dd4_2),.clk(gclk));
	jdff dff_B_CFnm898Y0_2(.din(w_dff_B_2RNSW0dd4_2),.dout(w_dff_B_CFnm898Y0_2),.clk(gclk));
	jdff dff_B_k77rVTrd2_2(.din(w_dff_B_CFnm898Y0_2),.dout(w_dff_B_k77rVTrd2_2),.clk(gclk));
	jdff dff_B_DA6fB0uE3_2(.din(w_dff_B_k77rVTrd2_2),.dout(w_dff_B_DA6fB0uE3_2),.clk(gclk));
	jdff dff_B_4H64QbTv2_2(.din(w_dff_B_DA6fB0uE3_2),.dout(w_dff_B_4H64QbTv2_2),.clk(gclk));
	jdff dff_B_5oAa4zcv6_2(.din(w_dff_B_4H64QbTv2_2),.dout(w_dff_B_5oAa4zcv6_2),.clk(gclk));
	jdff dff_B_APU4c4Aq1_2(.din(w_dff_B_5oAa4zcv6_2),.dout(w_dff_B_APU4c4Aq1_2),.clk(gclk));
	jdff dff_B_3GT30ZCg7_2(.din(w_dff_B_APU4c4Aq1_2),.dout(w_dff_B_3GT30ZCg7_2),.clk(gclk));
	jdff dff_B_bELeBRCW3_2(.din(w_dff_B_3GT30ZCg7_2),.dout(w_dff_B_bELeBRCW3_2),.clk(gclk));
	jdff dff_B_iE7qehjO7_2(.din(w_dff_B_bELeBRCW3_2),.dout(w_dff_B_iE7qehjO7_2),.clk(gclk));
	jdff dff_B_51i5gpmL9_2(.din(w_dff_B_iE7qehjO7_2),.dout(w_dff_B_51i5gpmL9_2),.clk(gclk));
	jdff dff_B_mF8Ej48u5_2(.din(w_dff_B_51i5gpmL9_2),.dout(w_dff_B_mF8Ej48u5_2),.clk(gclk));
	jdff dff_B_HVnQXriL1_2(.din(w_dff_B_mF8Ej48u5_2),.dout(w_dff_B_HVnQXriL1_2),.clk(gclk));
	jdff dff_B_28SrPSr41_2(.din(w_dff_B_HVnQXriL1_2),.dout(w_dff_B_28SrPSr41_2),.clk(gclk));
	jdff dff_B_ioy2gMR02_2(.din(w_dff_B_28SrPSr41_2),.dout(w_dff_B_ioy2gMR02_2),.clk(gclk));
	jdff dff_B_y67DCB5M1_2(.din(w_dff_B_ioy2gMR02_2),.dout(w_dff_B_y67DCB5M1_2),.clk(gclk));
	jdff dff_B_QEgq628n1_2(.din(n372),.dout(w_dff_B_QEgq628n1_2),.clk(gclk));
	jdff dff_B_01uMWL296_1(.din(n331),.dout(w_dff_B_01uMWL296_1),.clk(gclk));
	jdff dff_B_a1T8jJQb3_2(.din(n274),.dout(w_dff_B_a1T8jJQb3_2),.clk(gclk));
	jdff dff_B_ZK8ndZg76_2(.din(w_dff_B_a1T8jJQb3_2),.dout(w_dff_B_ZK8ndZg76_2),.clk(gclk));
	jdff dff_B_kJ3DrL9d0_2(.din(w_dff_B_ZK8ndZg76_2),.dout(w_dff_B_kJ3DrL9d0_2),.clk(gclk));
	jdff dff_B_rEJg5UC37_2(.din(w_dff_B_kJ3DrL9d0_2),.dout(w_dff_B_rEJg5UC37_2),.clk(gclk));
	jdff dff_B_AX0bdwf96_2(.din(w_dff_B_rEJg5UC37_2),.dout(w_dff_B_AX0bdwf96_2),.clk(gclk));
	jdff dff_B_garsuYDJ8_2(.din(w_dff_B_AX0bdwf96_2),.dout(w_dff_B_garsuYDJ8_2),.clk(gclk));
	jdff dff_B_7d4TyI5H9_2(.din(w_dff_B_garsuYDJ8_2),.dout(w_dff_B_7d4TyI5H9_2),.clk(gclk));
	jdff dff_B_jYlutrkL3_2(.din(w_dff_B_7d4TyI5H9_2),.dout(w_dff_B_jYlutrkL3_2),.clk(gclk));
	jdff dff_B_w3BqEHiK9_2(.din(w_dff_B_jYlutrkL3_2),.dout(w_dff_B_w3BqEHiK9_2),.clk(gclk));
	jdff dff_B_21D6IUUz6_2(.din(w_dff_B_w3BqEHiK9_2),.dout(w_dff_B_21D6IUUz6_2),.clk(gclk));
	jdff dff_B_SnbnlTq58_2(.din(w_dff_B_21D6IUUz6_2),.dout(w_dff_B_SnbnlTq58_2),.clk(gclk));
	jdff dff_B_dadRfedO6_2(.din(w_dff_B_SnbnlTq58_2),.dout(w_dff_B_dadRfedO6_2),.clk(gclk));
	jdff dff_B_BI0V2RgV0_2(.din(w_dff_B_dadRfedO6_2),.dout(w_dff_B_BI0V2RgV0_2),.clk(gclk));
	jdff dff_B_fGx0M5r74_2(.din(w_dff_B_BI0V2RgV0_2),.dout(w_dff_B_fGx0M5r74_2),.clk(gclk));
	jdff dff_B_4xzSKqT53_2(.din(w_dff_B_fGx0M5r74_2),.dout(w_dff_B_4xzSKqT53_2),.clk(gclk));
	jdff dff_B_O5DfBWIa0_2(.din(n309),.dout(w_dff_B_O5DfBWIa0_2),.clk(gclk));
	jdff dff_B_4NcILaiO4_1(.din(n275),.dout(w_dff_B_4NcILaiO4_1),.clk(gclk));
	jdff dff_B_hWBQMU3w6_2(.din(n225),.dout(w_dff_B_hWBQMU3w6_2),.clk(gclk));
	jdff dff_B_I9RT2yjy3_2(.din(w_dff_B_hWBQMU3w6_2),.dout(w_dff_B_I9RT2yjy3_2),.clk(gclk));
	jdff dff_B_8mHZPK9a1_2(.din(w_dff_B_I9RT2yjy3_2),.dout(w_dff_B_8mHZPK9a1_2),.clk(gclk));
	jdff dff_B_DAN92S8r7_2(.din(w_dff_B_8mHZPK9a1_2),.dout(w_dff_B_DAN92S8r7_2),.clk(gclk));
	jdff dff_B_V0YjDXYs4_2(.din(w_dff_B_DAN92S8r7_2),.dout(w_dff_B_V0YjDXYs4_2),.clk(gclk));
	jdff dff_B_v98BEKwL6_2(.din(w_dff_B_V0YjDXYs4_2),.dout(w_dff_B_v98BEKwL6_2),.clk(gclk));
	jdff dff_B_gYvV5HxF7_2(.din(w_dff_B_v98BEKwL6_2),.dout(w_dff_B_gYvV5HxF7_2),.clk(gclk));
	jdff dff_B_6jVmbgM30_2(.din(w_dff_B_gYvV5HxF7_2),.dout(w_dff_B_6jVmbgM30_2),.clk(gclk));
	jdff dff_B_5VJc7xDt7_2(.din(w_dff_B_6jVmbgM30_2),.dout(w_dff_B_5VJc7xDt7_2),.clk(gclk));
	jdff dff_B_uzJH1FrF2_2(.din(w_dff_B_5VJc7xDt7_2),.dout(w_dff_B_uzJH1FrF2_2),.clk(gclk));
	jdff dff_B_cX0SYfVX4_2(.din(w_dff_B_uzJH1FrF2_2),.dout(w_dff_B_cX0SYfVX4_2),.clk(gclk));
	jdff dff_B_7od6T22O2_2(.din(w_dff_B_cX0SYfVX4_2),.dout(w_dff_B_7od6T22O2_2),.clk(gclk));
	jdff dff_B_gHhvR5im2_2(.din(n253),.dout(w_dff_B_gHhvR5im2_2),.clk(gclk));
	jdff dff_B_awINEBjq5_1(.din(n226),.dout(w_dff_B_awINEBjq5_1),.clk(gclk));
	jdff dff_B_lJxH3CAW7_2(.din(n183),.dout(w_dff_B_lJxH3CAW7_2),.clk(gclk));
	jdff dff_B_R7uqlSYm0_2(.din(w_dff_B_lJxH3CAW7_2),.dout(w_dff_B_R7uqlSYm0_2),.clk(gclk));
	jdff dff_B_uC870PGZ9_2(.din(w_dff_B_R7uqlSYm0_2),.dout(w_dff_B_uC870PGZ9_2),.clk(gclk));
	jdff dff_B_aoGuBHfk3_2(.din(w_dff_B_uC870PGZ9_2),.dout(w_dff_B_aoGuBHfk3_2),.clk(gclk));
	jdff dff_B_hhSrjFqh1_2(.din(w_dff_B_aoGuBHfk3_2),.dout(w_dff_B_hhSrjFqh1_2),.clk(gclk));
	jdff dff_B_vZJGX8Ys3_2(.din(w_dff_B_hhSrjFqh1_2),.dout(w_dff_B_vZJGX8Ys3_2),.clk(gclk));
	jdff dff_B_Qv5EgmYz6_2(.din(w_dff_B_vZJGX8Ys3_2),.dout(w_dff_B_Qv5EgmYz6_2),.clk(gclk));
	jdff dff_B_YsN32FRz8_2(.din(w_dff_B_Qv5EgmYz6_2),.dout(w_dff_B_YsN32FRz8_2),.clk(gclk));
	jdff dff_B_zjj0zFqA2_2(.din(w_dff_B_YsN32FRz8_2),.dout(w_dff_B_zjj0zFqA2_2),.clk(gclk));
	jdff dff_B_OTekOYmC2_2(.din(n204),.dout(w_dff_B_OTekOYmC2_2),.clk(gclk));
	jdff dff_B_Duh6237q9_1(.din(n184),.dout(w_dff_B_Duh6237q9_1),.clk(gclk));
	jdff dff_B_IfhUVmGC1_2(.din(n148),.dout(w_dff_B_IfhUVmGC1_2),.clk(gclk));
	jdff dff_B_LczE3Lmg0_2(.din(w_dff_B_IfhUVmGC1_2),.dout(w_dff_B_LczE3Lmg0_2),.clk(gclk));
	jdff dff_B_liEYByHO6_2(.din(w_dff_B_LczE3Lmg0_2),.dout(w_dff_B_liEYByHO6_2),.clk(gclk));
	jdff dff_B_QNxxOwXm4_2(.din(w_dff_B_liEYByHO6_2),.dout(w_dff_B_QNxxOwXm4_2),.clk(gclk));
	jdff dff_B_KefqDJAc4_2(.din(w_dff_B_QNxxOwXm4_2),.dout(w_dff_B_KefqDJAc4_2),.clk(gclk));
	jdff dff_B_7T33LGME5_2(.din(w_dff_B_KefqDJAc4_2),.dout(w_dff_B_7T33LGME5_2),.clk(gclk));
	jdff dff_B_My0VlJMI7_2(.din(n162),.dout(w_dff_B_My0VlJMI7_2),.clk(gclk));
	jdff dff_B_TbGNR3Fo0_2(.din(n119),.dout(w_dff_B_TbGNR3Fo0_2),.clk(gclk));
	jdff dff_B_YHLHf0045_2(.din(w_dff_B_TbGNR3Fo0_2),.dout(w_dff_B_YHLHf0045_2),.clk(gclk));
	jdff dff_B_WUu4GHNc7_2(.din(w_dff_B_YHLHf0045_2),.dout(w_dff_B_WUu4GHNc7_2),.clk(gclk));
	jdff dff_B_ULWUSYyN0_0(.din(n126),.dout(w_dff_B_ULWUSYyN0_0),.clk(gclk));
	jdff dff_B_T7uFMeCt1_0(.din(n1298),.dout(w_dff_B_T7uFMeCt1_0),.clk(gclk));
	jdff dff_A_0aHcLnK74_1(.dout(w_n1294_0[1]),.din(w_dff_A_0aHcLnK74_1),.clk(gclk));
	jdff dff_A_vXmbbNVz1_1(.dout(w_dff_A_0aHcLnK74_1),.din(w_dff_A_vXmbbNVz1_1),.clk(gclk));
	jdff dff_B_5cYZM5lH4_1(.din(n1214),.dout(w_dff_B_5cYZM5lH4_1),.clk(gclk));
	jdff dff_B_dNEC8t638_1(.din(w_dff_B_5cYZM5lH4_1),.dout(w_dff_B_dNEC8t638_1),.clk(gclk));
	jdff dff_B_5FxeB74n6_2(.din(n1120),.dout(w_dff_B_5FxeB74n6_2),.clk(gclk));
	jdff dff_B_8eU6m3TK0_2(.din(w_dff_B_5FxeB74n6_2),.dout(w_dff_B_8eU6m3TK0_2),.clk(gclk));
	jdff dff_B_aY7vb9RH3_2(.din(w_dff_B_8eU6m3TK0_2),.dout(w_dff_B_aY7vb9RH3_2),.clk(gclk));
	jdff dff_B_j3Y2cl8M0_2(.din(w_dff_B_aY7vb9RH3_2),.dout(w_dff_B_j3Y2cl8M0_2),.clk(gclk));
	jdff dff_B_uQAWDbP54_2(.din(w_dff_B_j3Y2cl8M0_2),.dout(w_dff_B_uQAWDbP54_2),.clk(gclk));
	jdff dff_B_uLO0FDRf1_2(.din(w_dff_B_uQAWDbP54_2),.dout(w_dff_B_uLO0FDRf1_2),.clk(gclk));
	jdff dff_B_nYY0mzsr5_2(.din(w_dff_B_uLO0FDRf1_2),.dout(w_dff_B_nYY0mzsr5_2),.clk(gclk));
	jdff dff_B_ojeGawvS1_2(.din(w_dff_B_nYY0mzsr5_2),.dout(w_dff_B_ojeGawvS1_2),.clk(gclk));
	jdff dff_B_sDHPtxl30_2(.din(w_dff_B_ojeGawvS1_2),.dout(w_dff_B_sDHPtxl30_2),.clk(gclk));
	jdff dff_B_VcHc3vAx3_2(.din(w_dff_B_sDHPtxl30_2),.dout(w_dff_B_VcHc3vAx3_2),.clk(gclk));
	jdff dff_B_zutsqV7m8_2(.din(w_dff_B_VcHc3vAx3_2),.dout(w_dff_B_zutsqV7m8_2),.clk(gclk));
	jdff dff_B_wRJE5q9U3_2(.din(w_dff_B_zutsqV7m8_2),.dout(w_dff_B_wRJE5q9U3_2),.clk(gclk));
	jdff dff_B_Oe9lUesJ4_2(.din(w_dff_B_wRJE5q9U3_2),.dout(w_dff_B_Oe9lUesJ4_2),.clk(gclk));
	jdff dff_B_qkrpvotO8_2(.din(w_dff_B_Oe9lUesJ4_2),.dout(w_dff_B_qkrpvotO8_2),.clk(gclk));
	jdff dff_B_YM7dK0EM3_2(.din(w_dff_B_qkrpvotO8_2),.dout(w_dff_B_YM7dK0EM3_2),.clk(gclk));
	jdff dff_B_X6WEpmbD5_2(.din(w_dff_B_YM7dK0EM3_2),.dout(w_dff_B_X6WEpmbD5_2),.clk(gclk));
	jdff dff_B_CQJ9m3qm2_2(.din(w_dff_B_X6WEpmbD5_2),.dout(w_dff_B_CQJ9m3qm2_2),.clk(gclk));
	jdff dff_B_1PGOmBdS1_2(.din(w_dff_B_CQJ9m3qm2_2),.dout(w_dff_B_1PGOmBdS1_2),.clk(gclk));
	jdff dff_B_HCSCg9zD9_2(.din(w_dff_B_1PGOmBdS1_2),.dout(w_dff_B_HCSCg9zD9_2),.clk(gclk));
	jdff dff_B_PqEYFeOp0_2(.din(w_dff_B_HCSCg9zD9_2),.dout(w_dff_B_PqEYFeOp0_2),.clk(gclk));
	jdff dff_B_DDibQBoL1_2(.din(w_dff_B_PqEYFeOp0_2),.dout(w_dff_B_DDibQBoL1_2),.clk(gclk));
	jdff dff_B_2N9rZFQa5_2(.din(w_dff_B_DDibQBoL1_2),.dout(w_dff_B_2N9rZFQa5_2),.clk(gclk));
	jdff dff_B_cZzXQ1nW6_2(.din(w_dff_B_2N9rZFQa5_2),.dout(w_dff_B_cZzXQ1nW6_2),.clk(gclk));
	jdff dff_B_DrDDijPw6_2(.din(w_dff_B_cZzXQ1nW6_2),.dout(w_dff_B_DrDDijPw6_2),.clk(gclk));
	jdff dff_B_XVwnxa3E9_2(.din(w_dff_B_DrDDijPw6_2),.dout(w_dff_B_XVwnxa3E9_2),.clk(gclk));
	jdff dff_B_ECwYTLId8_2(.din(w_dff_B_XVwnxa3E9_2),.dout(w_dff_B_ECwYTLId8_2),.clk(gclk));
	jdff dff_B_NAQ7WFtU0_2(.din(w_dff_B_ECwYTLId8_2),.dout(w_dff_B_NAQ7WFtU0_2),.clk(gclk));
	jdff dff_B_kMFTsYbB8_2(.din(w_dff_B_NAQ7WFtU0_2),.dout(w_dff_B_kMFTsYbB8_2),.clk(gclk));
	jdff dff_B_R1yWHHhj0_2(.din(w_dff_B_kMFTsYbB8_2),.dout(w_dff_B_R1yWHHhj0_2),.clk(gclk));
	jdff dff_B_aP5expyP3_2(.din(w_dff_B_R1yWHHhj0_2),.dout(w_dff_B_aP5expyP3_2),.clk(gclk));
	jdff dff_B_qWS2rGsJ2_2(.din(w_dff_B_aP5expyP3_2),.dout(w_dff_B_qWS2rGsJ2_2),.clk(gclk));
	jdff dff_B_9dlO2y3O1_2(.din(w_dff_B_qWS2rGsJ2_2),.dout(w_dff_B_9dlO2y3O1_2),.clk(gclk));
	jdff dff_B_lL2U8Set6_2(.din(w_dff_B_9dlO2y3O1_2),.dout(w_dff_B_lL2U8Set6_2),.clk(gclk));
	jdff dff_B_RD5pl4S27_2(.din(w_dff_B_lL2U8Set6_2),.dout(w_dff_B_RD5pl4S27_2),.clk(gclk));
	jdff dff_B_vSTGKNJT7_2(.din(w_dff_B_RD5pl4S27_2),.dout(w_dff_B_vSTGKNJT7_2),.clk(gclk));
	jdff dff_B_JHPmVqIP0_2(.din(w_dff_B_vSTGKNJT7_2),.dout(w_dff_B_JHPmVqIP0_2),.clk(gclk));
	jdff dff_B_D7ei4GmZ8_2(.din(w_dff_B_JHPmVqIP0_2),.dout(w_dff_B_D7ei4GmZ8_2),.clk(gclk));
	jdff dff_B_gk4THjet9_2(.din(w_dff_B_D7ei4GmZ8_2),.dout(w_dff_B_gk4THjet9_2),.clk(gclk));
	jdff dff_B_Aizn5nb75_2(.din(w_dff_B_gk4THjet9_2),.dout(w_dff_B_Aizn5nb75_2),.clk(gclk));
	jdff dff_B_O4AsLtNS0_2(.din(w_dff_B_Aizn5nb75_2),.dout(w_dff_B_O4AsLtNS0_2),.clk(gclk));
	jdff dff_B_7R6rw7q18_2(.din(w_dff_B_O4AsLtNS0_2),.dout(w_dff_B_7R6rw7q18_2),.clk(gclk));
	jdff dff_B_lmnA66fG7_2(.din(w_dff_B_7R6rw7q18_2),.dout(w_dff_B_lmnA66fG7_2),.clk(gclk));
	jdff dff_B_IJ0Z0k6e4_2(.din(w_dff_B_lmnA66fG7_2),.dout(w_dff_B_IJ0Z0k6e4_2),.clk(gclk));
	jdff dff_B_8V8XETCW6_2(.din(w_dff_B_IJ0Z0k6e4_2),.dout(w_dff_B_8V8XETCW6_2),.clk(gclk));
	jdff dff_B_N6CcgjhU8_2(.din(w_dff_B_8V8XETCW6_2),.dout(w_dff_B_N6CcgjhU8_2),.clk(gclk));
	jdff dff_B_g5qSM25j2_2(.din(n1203),.dout(w_dff_B_g5qSM25j2_2),.clk(gclk));
	jdff dff_B_dTWjquK89_1(.din(n1122),.dout(w_dff_B_dTWjquK89_1),.clk(gclk));
	jdff dff_B_LaUlfFI53_2(.din(n1023),.dout(w_dff_B_LaUlfFI53_2),.clk(gclk));
	jdff dff_B_gMn8pWZ36_2(.din(w_dff_B_LaUlfFI53_2),.dout(w_dff_B_gMn8pWZ36_2),.clk(gclk));
	jdff dff_B_xFQ39yQZ5_2(.din(w_dff_B_gMn8pWZ36_2),.dout(w_dff_B_xFQ39yQZ5_2),.clk(gclk));
	jdff dff_B_uNDwr3PX4_2(.din(w_dff_B_xFQ39yQZ5_2),.dout(w_dff_B_uNDwr3PX4_2),.clk(gclk));
	jdff dff_B_xpZFzXIR8_2(.din(w_dff_B_uNDwr3PX4_2),.dout(w_dff_B_xpZFzXIR8_2),.clk(gclk));
	jdff dff_B_C8qaNjaP0_2(.din(w_dff_B_xpZFzXIR8_2),.dout(w_dff_B_C8qaNjaP0_2),.clk(gclk));
	jdff dff_B_NLYtQFB73_2(.din(w_dff_B_C8qaNjaP0_2),.dout(w_dff_B_NLYtQFB73_2),.clk(gclk));
	jdff dff_B_NE8sBkr32_2(.din(w_dff_B_NLYtQFB73_2),.dout(w_dff_B_NE8sBkr32_2),.clk(gclk));
	jdff dff_B_GclNvpcU8_2(.din(w_dff_B_NE8sBkr32_2),.dout(w_dff_B_GclNvpcU8_2),.clk(gclk));
	jdff dff_B_LRHHXjOn1_2(.din(w_dff_B_GclNvpcU8_2),.dout(w_dff_B_LRHHXjOn1_2),.clk(gclk));
	jdff dff_B_rj4sTifu3_2(.din(w_dff_B_LRHHXjOn1_2),.dout(w_dff_B_rj4sTifu3_2),.clk(gclk));
	jdff dff_B_qHMjqg013_2(.din(w_dff_B_rj4sTifu3_2),.dout(w_dff_B_qHMjqg013_2),.clk(gclk));
	jdff dff_B_ghLWkcMT2_2(.din(w_dff_B_qHMjqg013_2),.dout(w_dff_B_ghLWkcMT2_2),.clk(gclk));
	jdff dff_B_KbVaCQiV0_2(.din(w_dff_B_ghLWkcMT2_2),.dout(w_dff_B_KbVaCQiV0_2),.clk(gclk));
	jdff dff_B_y5ZHfqiq0_2(.din(w_dff_B_KbVaCQiV0_2),.dout(w_dff_B_y5ZHfqiq0_2),.clk(gclk));
	jdff dff_B_mXz8Kk2I4_2(.din(w_dff_B_y5ZHfqiq0_2),.dout(w_dff_B_mXz8Kk2I4_2),.clk(gclk));
	jdff dff_B_k5GTW3aM6_2(.din(w_dff_B_mXz8Kk2I4_2),.dout(w_dff_B_k5GTW3aM6_2),.clk(gclk));
	jdff dff_B_R3VdjnQB9_2(.din(w_dff_B_k5GTW3aM6_2),.dout(w_dff_B_R3VdjnQB9_2),.clk(gclk));
	jdff dff_B_F5OGTpki4_2(.din(w_dff_B_R3VdjnQB9_2),.dout(w_dff_B_F5OGTpki4_2),.clk(gclk));
	jdff dff_B_JjP8fJdZ6_2(.din(w_dff_B_F5OGTpki4_2),.dout(w_dff_B_JjP8fJdZ6_2),.clk(gclk));
	jdff dff_B_xH3nT4zI4_2(.din(w_dff_B_JjP8fJdZ6_2),.dout(w_dff_B_xH3nT4zI4_2),.clk(gclk));
	jdff dff_B_I777N9s45_2(.din(w_dff_B_xH3nT4zI4_2),.dout(w_dff_B_I777N9s45_2),.clk(gclk));
	jdff dff_B_OnC1kYJD0_2(.din(w_dff_B_I777N9s45_2),.dout(w_dff_B_OnC1kYJD0_2),.clk(gclk));
	jdff dff_B_TQlTeIfE5_2(.din(w_dff_B_OnC1kYJD0_2),.dout(w_dff_B_TQlTeIfE5_2),.clk(gclk));
	jdff dff_B_IC9zf8wU6_2(.din(w_dff_B_TQlTeIfE5_2),.dout(w_dff_B_IC9zf8wU6_2),.clk(gclk));
	jdff dff_B_kotpLJaf9_2(.din(w_dff_B_IC9zf8wU6_2),.dout(w_dff_B_kotpLJaf9_2),.clk(gclk));
	jdff dff_B_lC6K6ift0_2(.din(w_dff_B_kotpLJaf9_2),.dout(w_dff_B_lC6K6ift0_2),.clk(gclk));
	jdff dff_B_ZYwrdI9z7_2(.din(w_dff_B_lC6K6ift0_2),.dout(w_dff_B_ZYwrdI9z7_2),.clk(gclk));
	jdff dff_B_akkOtuSs1_2(.din(w_dff_B_ZYwrdI9z7_2),.dout(w_dff_B_akkOtuSs1_2),.clk(gclk));
	jdff dff_B_CJVmzvky6_2(.din(w_dff_B_akkOtuSs1_2),.dout(w_dff_B_CJVmzvky6_2),.clk(gclk));
	jdff dff_B_fvc3LnZ15_2(.din(w_dff_B_CJVmzvky6_2),.dout(w_dff_B_fvc3LnZ15_2),.clk(gclk));
	jdff dff_B_GRWKdhPT1_2(.din(w_dff_B_fvc3LnZ15_2),.dout(w_dff_B_GRWKdhPT1_2),.clk(gclk));
	jdff dff_B_uiYizq8T8_2(.din(w_dff_B_GRWKdhPT1_2),.dout(w_dff_B_uiYizq8T8_2),.clk(gclk));
	jdff dff_B_PxS9NFLH7_2(.din(w_dff_B_uiYizq8T8_2),.dout(w_dff_B_PxS9NFLH7_2),.clk(gclk));
	jdff dff_B_jfCAjWSx2_2(.din(w_dff_B_PxS9NFLH7_2),.dout(w_dff_B_jfCAjWSx2_2),.clk(gclk));
	jdff dff_B_STRwvEif1_2(.din(w_dff_B_jfCAjWSx2_2),.dout(w_dff_B_STRwvEif1_2),.clk(gclk));
	jdff dff_B_6tlaWTFm4_2(.din(w_dff_B_STRwvEif1_2),.dout(w_dff_B_6tlaWTFm4_2),.clk(gclk));
	jdff dff_B_nB4hcta01_2(.din(w_dff_B_6tlaWTFm4_2),.dout(w_dff_B_nB4hcta01_2),.clk(gclk));
	jdff dff_B_Gd5v9ywR2_2(.din(w_dff_B_nB4hcta01_2),.dout(w_dff_B_Gd5v9ywR2_2),.clk(gclk));
	jdff dff_B_gPTWyeiH9_2(.din(w_dff_B_Gd5v9ywR2_2),.dout(w_dff_B_gPTWyeiH9_2),.clk(gclk));
	jdff dff_B_IcKyzXsc3_2(.din(w_dff_B_gPTWyeiH9_2),.dout(w_dff_B_IcKyzXsc3_2),.clk(gclk));
	jdff dff_B_LOO3qfnl6_2(.din(n1103),.dout(w_dff_B_LOO3qfnl6_2),.clk(gclk));
	jdff dff_B_jSsFNk300_1(.din(n1024),.dout(w_dff_B_jSsFNk300_1),.clk(gclk));
	jdff dff_B_0XkwwTlN3_2(.din(n924),.dout(w_dff_B_0XkwwTlN3_2),.clk(gclk));
	jdff dff_B_t0ZJEpMk9_2(.din(w_dff_B_0XkwwTlN3_2),.dout(w_dff_B_t0ZJEpMk9_2),.clk(gclk));
	jdff dff_B_BaaxaJfV9_2(.din(w_dff_B_t0ZJEpMk9_2),.dout(w_dff_B_BaaxaJfV9_2),.clk(gclk));
	jdff dff_B_1ZXBBSUE7_2(.din(w_dff_B_BaaxaJfV9_2),.dout(w_dff_B_1ZXBBSUE7_2),.clk(gclk));
	jdff dff_B_DkTebevs3_2(.din(w_dff_B_1ZXBBSUE7_2),.dout(w_dff_B_DkTebevs3_2),.clk(gclk));
	jdff dff_B_2snPNeIM4_2(.din(w_dff_B_DkTebevs3_2),.dout(w_dff_B_2snPNeIM4_2),.clk(gclk));
	jdff dff_B_PQ6QK7BE4_2(.din(w_dff_B_2snPNeIM4_2),.dout(w_dff_B_PQ6QK7BE4_2),.clk(gclk));
	jdff dff_B_AaPCN2NS7_2(.din(w_dff_B_PQ6QK7BE4_2),.dout(w_dff_B_AaPCN2NS7_2),.clk(gclk));
	jdff dff_B_ZpQbhU5f9_2(.din(w_dff_B_AaPCN2NS7_2),.dout(w_dff_B_ZpQbhU5f9_2),.clk(gclk));
	jdff dff_B_XeU8s8Dm4_2(.din(w_dff_B_ZpQbhU5f9_2),.dout(w_dff_B_XeU8s8Dm4_2),.clk(gclk));
	jdff dff_B_NX8IPIdd2_2(.din(w_dff_B_XeU8s8Dm4_2),.dout(w_dff_B_NX8IPIdd2_2),.clk(gclk));
	jdff dff_B_tkQr5MJK0_2(.din(w_dff_B_NX8IPIdd2_2),.dout(w_dff_B_tkQr5MJK0_2),.clk(gclk));
	jdff dff_B_50oh49lC2_2(.din(w_dff_B_tkQr5MJK0_2),.dout(w_dff_B_50oh49lC2_2),.clk(gclk));
	jdff dff_B_FTUJpMRK9_2(.din(w_dff_B_50oh49lC2_2),.dout(w_dff_B_FTUJpMRK9_2),.clk(gclk));
	jdff dff_B_GI3tVzFC1_2(.din(w_dff_B_FTUJpMRK9_2),.dout(w_dff_B_GI3tVzFC1_2),.clk(gclk));
	jdff dff_B_jigLqi2P8_2(.din(w_dff_B_GI3tVzFC1_2),.dout(w_dff_B_jigLqi2P8_2),.clk(gclk));
	jdff dff_B_AjNQBBmb3_2(.din(w_dff_B_jigLqi2P8_2),.dout(w_dff_B_AjNQBBmb3_2),.clk(gclk));
	jdff dff_B_2nesTlPu1_2(.din(w_dff_B_AjNQBBmb3_2),.dout(w_dff_B_2nesTlPu1_2),.clk(gclk));
	jdff dff_B_zUy7i4RU1_2(.din(w_dff_B_2nesTlPu1_2),.dout(w_dff_B_zUy7i4RU1_2),.clk(gclk));
	jdff dff_B_N0tbAMdL5_2(.din(w_dff_B_zUy7i4RU1_2),.dout(w_dff_B_N0tbAMdL5_2),.clk(gclk));
	jdff dff_B_8yFXKhmv1_2(.din(w_dff_B_N0tbAMdL5_2),.dout(w_dff_B_8yFXKhmv1_2),.clk(gclk));
	jdff dff_B_PwQOxcPN8_2(.din(w_dff_B_8yFXKhmv1_2),.dout(w_dff_B_PwQOxcPN8_2),.clk(gclk));
	jdff dff_B_1PR57Ky75_2(.din(w_dff_B_PwQOxcPN8_2),.dout(w_dff_B_1PR57Ky75_2),.clk(gclk));
	jdff dff_B_DqTMZJTI9_2(.din(w_dff_B_1PR57Ky75_2),.dout(w_dff_B_DqTMZJTI9_2),.clk(gclk));
	jdff dff_B_RwA7FrXB8_2(.din(w_dff_B_DqTMZJTI9_2),.dout(w_dff_B_RwA7FrXB8_2),.clk(gclk));
	jdff dff_B_ptrrO5bo4_2(.din(w_dff_B_RwA7FrXB8_2),.dout(w_dff_B_ptrrO5bo4_2),.clk(gclk));
	jdff dff_B_mAn2FqFP0_2(.din(w_dff_B_ptrrO5bo4_2),.dout(w_dff_B_mAn2FqFP0_2),.clk(gclk));
	jdff dff_B_uZhgiULn1_2(.din(w_dff_B_mAn2FqFP0_2),.dout(w_dff_B_uZhgiULn1_2),.clk(gclk));
	jdff dff_B_bmx5x4EL3_2(.din(w_dff_B_uZhgiULn1_2),.dout(w_dff_B_bmx5x4EL3_2),.clk(gclk));
	jdff dff_B_MxOZXmWe0_2(.din(w_dff_B_bmx5x4EL3_2),.dout(w_dff_B_MxOZXmWe0_2),.clk(gclk));
	jdff dff_B_tVDbwprB8_2(.din(w_dff_B_MxOZXmWe0_2),.dout(w_dff_B_tVDbwprB8_2),.clk(gclk));
	jdff dff_B_zquJMwJE9_2(.din(w_dff_B_tVDbwprB8_2),.dout(w_dff_B_zquJMwJE9_2),.clk(gclk));
	jdff dff_B_6L2faNIN0_2(.din(w_dff_B_zquJMwJE9_2),.dout(w_dff_B_6L2faNIN0_2),.clk(gclk));
	jdff dff_B_nxNZdasy7_2(.din(w_dff_B_6L2faNIN0_2),.dout(w_dff_B_nxNZdasy7_2),.clk(gclk));
	jdff dff_B_iESR9fib1_2(.din(w_dff_B_nxNZdasy7_2),.dout(w_dff_B_iESR9fib1_2),.clk(gclk));
	jdff dff_B_xChHUj2Q5_2(.din(w_dff_B_iESR9fib1_2),.dout(w_dff_B_xChHUj2Q5_2),.clk(gclk));
	jdff dff_B_ETjCxcFW4_2(.din(n1004),.dout(w_dff_B_ETjCxcFW4_2),.clk(gclk));
	jdff dff_B_S5HypYcJ0_1(.din(n925),.dout(w_dff_B_S5HypYcJ0_1),.clk(gclk));
	jdff dff_B_BKIzaoqq7_2(.din(n822),.dout(w_dff_B_BKIzaoqq7_2),.clk(gclk));
	jdff dff_B_4efNMmNp7_2(.din(w_dff_B_BKIzaoqq7_2),.dout(w_dff_B_4efNMmNp7_2),.clk(gclk));
	jdff dff_B_MQzKKLNi5_2(.din(w_dff_B_4efNMmNp7_2),.dout(w_dff_B_MQzKKLNi5_2),.clk(gclk));
	jdff dff_B_kdiv25xZ1_2(.din(w_dff_B_MQzKKLNi5_2),.dout(w_dff_B_kdiv25xZ1_2),.clk(gclk));
	jdff dff_B_m3CTBBds8_2(.din(w_dff_B_kdiv25xZ1_2),.dout(w_dff_B_m3CTBBds8_2),.clk(gclk));
	jdff dff_B_fwe6veCj2_2(.din(w_dff_B_m3CTBBds8_2),.dout(w_dff_B_fwe6veCj2_2),.clk(gclk));
	jdff dff_B_lzC79Yp17_2(.din(w_dff_B_fwe6veCj2_2),.dout(w_dff_B_lzC79Yp17_2),.clk(gclk));
	jdff dff_B_jmQrW7v43_2(.din(w_dff_B_lzC79Yp17_2),.dout(w_dff_B_jmQrW7v43_2),.clk(gclk));
	jdff dff_B_GStMJizB3_2(.din(w_dff_B_jmQrW7v43_2),.dout(w_dff_B_GStMJizB3_2),.clk(gclk));
	jdff dff_B_jmCLi9nt9_2(.din(w_dff_B_GStMJizB3_2),.dout(w_dff_B_jmCLi9nt9_2),.clk(gclk));
	jdff dff_B_ZzAUrxgU7_2(.din(w_dff_B_jmCLi9nt9_2),.dout(w_dff_B_ZzAUrxgU7_2),.clk(gclk));
	jdff dff_B_WWkUyhEj8_2(.din(w_dff_B_ZzAUrxgU7_2),.dout(w_dff_B_WWkUyhEj8_2),.clk(gclk));
	jdff dff_B_a90X4dGt5_2(.din(w_dff_B_WWkUyhEj8_2),.dout(w_dff_B_a90X4dGt5_2),.clk(gclk));
	jdff dff_B_BZAq3Vyx5_2(.din(w_dff_B_a90X4dGt5_2),.dout(w_dff_B_BZAq3Vyx5_2),.clk(gclk));
	jdff dff_B_WM7HKaPc4_2(.din(w_dff_B_BZAq3Vyx5_2),.dout(w_dff_B_WM7HKaPc4_2),.clk(gclk));
	jdff dff_B_xvh14CFd3_2(.din(w_dff_B_WM7HKaPc4_2),.dout(w_dff_B_xvh14CFd3_2),.clk(gclk));
	jdff dff_B_YODdw0mT7_2(.din(w_dff_B_xvh14CFd3_2),.dout(w_dff_B_YODdw0mT7_2),.clk(gclk));
	jdff dff_B_F9SR7Nmp0_2(.din(w_dff_B_YODdw0mT7_2),.dout(w_dff_B_F9SR7Nmp0_2),.clk(gclk));
	jdff dff_B_JcRg1OUE0_2(.din(w_dff_B_F9SR7Nmp0_2),.dout(w_dff_B_JcRg1OUE0_2),.clk(gclk));
	jdff dff_B_FLaqh6SV7_2(.din(w_dff_B_JcRg1OUE0_2),.dout(w_dff_B_FLaqh6SV7_2),.clk(gclk));
	jdff dff_B_C9IZeMFD3_2(.din(w_dff_B_FLaqh6SV7_2),.dout(w_dff_B_C9IZeMFD3_2),.clk(gclk));
	jdff dff_B_WbwzmZ8a7_2(.din(w_dff_B_C9IZeMFD3_2),.dout(w_dff_B_WbwzmZ8a7_2),.clk(gclk));
	jdff dff_B_B897gTyX3_2(.din(w_dff_B_WbwzmZ8a7_2),.dout(w_dff_B_B897gTyX3_2),.clk(gclk));
	jdff dff_B_ZHXFM0Dt3_2(.din(w_dff_B_B897gTyX3_2),.dout(w_dff_B_ZHXFM0Dt3_2),.clk(gclk));
	jdff dff_B_cvNxBoHs4_2(.din(w_dff_B_ZHXFM0Dt3_2),.dout(w_dff_B_cvNxBoHs4_2),.clk(gclk));
	jdff dff_B_B7PPjqe50_2(.din(w_dff_B_cvNxBoHs4_2),.dout(w_dff_B_B7PPjqe50_2),.clk(gclk));
	jdff dff_B_sSi7FJ9F2_2(.din(w_dff_B_B7PPjqe50_2),.dout(w_dff_B_sSi7FJ9F2_2),.clk(gclk));
	jdff dff_B_UHvERiTK3_2(.din(w_dff_B_sSi7FJ9F2_2),.dout(w_dff_B_UHvERiTK3_2),.clk(gclk));
	jdff dff_B_cC5oSMNd5_2(.din(w_dff_B_UHvERiTK3_2),.dout(w_dff_B_cC5oSMNd5_2),.clk(gclk));
	jdff dff_B_KiCn9g8H1_2(.din(w_dff_B_cC5oSMNd5_2),.dout(w_dff_B_KiCn9g8H1_2),.clk(gclk));
	jdff dff_B_oPfQI8687_2(.din(w_dff_B_KiCn9g8H1_2),.dout(w_dff_B_oPfQI8687_2),.clk(gclk));
	jdff dff_B_Z7om9Y2Q4_2(.din(w_dff_B_oPfQI8687_2),.dout(w_dff_B_Z7om9Y2Q4_2),.clk(gclk));
	jdff dff_B_4qzbGwQl1_2(.din(w_dff_B_Z7om9Y2Q4_2),.dout(w_dff_B_4qzbGwQl1_2),.clk(gclk));
	jdff dff_B_UXHgDEAd7_2(.din(n898),.dout(w_dff_B_UXHgDEAd7_2),.clk(gclk));
	jdff dff_B_9fVbZpba6_1(.din(n823),.dout(w_dff_B_9fVbZpba6_1),.clk(gclk));
	jdff dff_B_YEeYVfOJ1_2(.din(n724),.dout(w_dff_B_YEeYVfOJ1_2),.clk(gclk));
	jdff dff_B_9njIobPw1_2(.din(w_dff_B_YEeYVfOJ1_2),.dout(w_dff_B_9njIobPw1_2),.clk(gclk));
	jdff dff_B_4LVZACzC4_2(.din(w_dff_B_9njIobPw1_2),.dout(w_dff_B_4LVZACzC4_2),.clk(gclk));
	jdff dff_B_5f5BNmE82_2(.din(w_dff_B_4LVZACzC4_2),.dout(w_dff_B_5f5BNmE82_2),.clk(gclk));
	jdff dff_B_sK8pOXa97_2(.din(w_dff_B_5f5BNmE82_2),.dout(w_dff_B_sK8pOXa97_2),.clk(gclk));
	jdff dff_B_ZiIp4TxA9_2(.din(w_dff_B_sK8pOXa97_2),.dout(w_dff_B_ZiIp4TxA9_2),.clk(gclk));
	jdff dff_B_6R4gMsf13_2(.din(w_dff_B_ZiIp4TxA9_2),.dout(w_dff_B_6R4gMsf13_2),.clk(gclk));
	jdff dff_B_a4fZc1ku5_2(.din(w_dff_B_6R4gMsf13_2),.dout(w_dff_B_a4fZc1ku5_2),.clk(gclk));
	jdff dff_B_dUZ6XPSa6_2(.din(w_dff_B_a4fZc1ku5_2),.dout(w_dff_B_dUZ6XPSa6_2),.clk(gclk));
	jdff dff_B_uCWOAT1R3_2(.din(w_dff_B_dUZ6XPSa6_2),.dout(w_dff_B_uCWOAT1R3_2),.clk(gclk));
	jdff dff_B_69UFl0bE5_2(.din(w_dff_B_uCWOAT1R3_2),.dout(w_dff_B_69UFl0bE5_2),.clk(gclk));
	jdff dff_B_Ojd71V7z6_2(.din(w_dff_B_69UFl0bE5_2),.dout(w_dff_B_Ojd71V7z6_2),.clk(gclk));
	jdff dff_B_PJf9AxCq0_2(.din(w_dff_B_Ojd71V7z6_2),.dout(w_dff_B_PJf9AxCq0_2),.clk(gclk));
	jdff dff_B_QAdZL6ED1_2(.din(w_dff_B_PJf9AxCq0_2),.dout(w_dff_B_QAdZL6ED1_2),.clk(gclk));
	jdff dff_B_YI0NXY1Q5_2(.din(w_dff_B_QAdZL6ED1_2),.dout(w_dff_B_YI0NXY1Q5_2),.clk(gclk));
	jdff dff_B_IehDabsF5_2(.din(w_dff_B_YI0NXY1Q5_2),.dout(w_dff_B_IehDabsF5_2),.clk(gclk));
	jdff dff_B_lrvEgepr2_2(.din(w_dff_B_IehDabsF5_2),.dout(w_dff_B_lrvEgepr2_2),.clk(gclk));
	jdff dff_B_lw8emsln6_2(.din(w_dff_B_lrvEgepr2_2),.dout(w_dff_B_lw8emsln6_2),.clk(gclk));
	jdff dff_B_G7iQ1yfU2_2(.din(w_dff_B_lw8emsln6_2),.dout(w_dff_B_G7iQ1yfU2_2),.clk(gclk));
	jdff dff_B_DUhNoIQU2_2(.din(w_dff_B_G7iQ1yfU2_2),.dout(w_dff_B_DUhNoIQU2_2),.clk(gclk));
	jdff dff_B_G4K64gZg7_2(.din(w_dff_B_DUhNoIQU2_2),.dout(w_dff_B_G4K64gZg7_2),.clk(gclk));
	jdff dff_B_PJs1L76p1_2(.din(w_dff_B_G4K64gZg7_2),.dout(w_dff_B_PJs1L76p1_2),.clk(gclk));
	jdff dff_B_ubGDez2D1_2(.din(w_dff_B_PJs1L76p1_2),.dout(w_dff_B_ubGDez2D1_2),.clk(gclk));
	jdff dff_B_hCeJSWaT6_2(.din(w_dff_B_ubGDez2D1_2),.dout(w_dff_B_hCeJSWaT6_2),.clk(gclk));
	jdff dff_B_KUivg05M3_2(.din(w_dff_B_hCeJSWaT6_2),.dout(w_dff_B_KUivg05M3_2),.clk(gclk));
	jdff dff_B_g243iE7M3_2(.din(w_dff_B_KUivg05M3_2),.dout(w_dff_B_g243iE7M3_2),.clk(gclk));
	jdff dff_B_QJ2js2vY6_2(.din(w_dff_B_g243iE7M3_2),.dout(w_dff_B_QJ2js2vY6_2),.clk(gclk));
	jdff dff_B_ndrO8KCb4_2(.din(w_dff_B_QJ2js2vY6_2),.dout(w_dff_B_ndrO8KCb4_2),.clk(gclk));
	jdff dff_B_G9acgQ5R7_2(.din(w_dff_B_ndrO8KCb4_2),.dout(w_dff_B_G9acgQ5R7_2),.clk(gclk));
	jdff dff_B_slip2qC92_2(.din(w_dff_B_G9acgQ5R7_2),.dout(w_dff_B_slip2qC92_2),.clk(gclk));
	jdff dff_B_AOXHx3Iw7_2(.din(n795),.dout(w_dff_B_AOXHx3Iw7_2),.clk(gclk));
	jdff dff_B_K4OtTcjG8_1(.din(n725),.dout(w_dff_B_K4OtTcjG8_1),.clk(gclk));
	jdff dff_B_bTOkVMSv7_2(.din(n632),.dout(w_dff_B_bTOkVMSv7_2),.clk(gclk));
	jdff dff_B_wohXghU12_2(.din(w_dff_B_bTOkVMSv7_2),.dout(w_dff_B_wohXghU12_2),.clk(gclk));
	jdff dff_B_JSNKy6jv4_2(.din(w_dff_B_wohXghU12_2),.dout(w_dff_B_JSNKy6jv4_2),.clk(gclk));
	jdff dff_B_RTP7oSkr6_2(.din(w_dff_B_JSNKy6jv4_2),.dout(w_dff_B_RTP7oSkr6_2),.clk(gclk));
	jdff dff_B_Fvk8zEjL4_2(.din(w_dff_B_RTP7oSkr6_2),.dout(w_dff_B_Fvk8zEjL4_2),.clk(gclk));
	jdff dff_B_lxmqH57C9_2(.din(w_dff_B_Fvk8zEjL4_2),.dout(w_dff_B_lxmqH57C9_2),.clk(gclk));
	jdff dff_B_RpME737s0_2(.din(w_dff_B_lxmqH57C9_2),.dout(w_dff_B_RpME737s0_2),.clk(gclk));
	jdff dff_B_L90nQbkT0_2(.din(w_dff_B_RpME737s0_2),.dout(w_dff_B_L90nQbkT0_2),.clk(gclk));
	jdff dff_B_hLXuRUF25_2(.din(w_dff_B_L90nQbkT0_2),.dout(w_dff_B_hLXuRUF25_2),.clk(gclk));
	jdff dff_B_NzuY3Hib3_2(.din(w_dff_B_hLXuRUF25_2),.dout(w_dff_B_NzuY3Hib3_2),.clk(gclk));
	jdff dff_B_74JS0qwJ7_2(.din(w_dff_B_NzuY3Hib3_2),.dout(w_dff_B_74JS0qwJ7_2),.clk(gclk));
	jdff dff_B_s5zUVmvx7_2(.din(w_dff_B_74JS0qwJ7_2),.dout(w_dff_B_s5zUVmvx7_2),.clk(gclk));
	jdff dff_B_VXhF3oOD5_2(.din(w_dff_B_s5zUVmvx7_2),.dout(w_dff_B_VXhF3oOD5_2),.clk(gclk));
	jdff dff_B_MRDj5VZy9_2(.din(w_dff_B_VXhF3oOD5_2),.dout(w_dff_B_MRDj5VZy9_2),.clk(gclk));
	jdff dff_B_bUejtSQi4_2(.din(w_dff_B_MRDj5VZy9_2),.dout(w_dff_B_bUejtSQi4_2),.clk(gclk));
	jdff dff_B_8KkOINzm9_2(.din(w_dff_B_bUejtSQi4_2),.dout(w_dff_B_8KkOINzm9_2),.clk(gclk));
	jdff dff_B_rxAcwCsf7_2(.din(w_dff_B_8KkOINzm9_2),.dout(w_dff_B_rxAcwCsf7_2),.clk(gclk));
	jdff dff_B_Ow7OnWlN3_2(.din(w_dff_B_rxAcwCsf7_2),.dout(w_dff_B_Ow7OnWlN3_2),.clk(gclk));
	jdff dff_B_A9AL2n199_2(.din(w_dff_B_Ow7OnWlN3_2),.dout(w_dff_B_A9AL2n199_2),.clk(gclk));
	jdff dff_B_Zlob5Hhh8_2(.din(w_dff_B_A9AL2n199_2),.dout(w_dff_B_Zlob5Hhh8_2),.clk(gclk));
	jdff dff_B_yHRWIc8f1_2(.din(w_dff_B_Zlob5Hhh8_2),.dout(w_dff_B_yHRWIc8f1_2),.clk(gclk));
	jdff dff_B_hRDE12xl0_2(.din(w_dff_B_yHRWIc8f1_2),.dout(w_dff_B_hRDE12xl0_2),.clk(gclk));
	jdff dff_B_e65a5p1x4_2(.din(w_dff_B_hRDE12xl0_2),.dout(w_dff_B_e65a5p1x4_2),.clk(gclk));
	jdff dff_B_Sm99qv2Q2_2(.din(w_dff_B_e65a5p1x4_2),.dout(w_dff_B_Sm99qv2Q2_2),.clk(gclk));
	jdff dff_B_qz9OmIKW8_2(.din(w_dff_B_Sm99qv2Q2_2),.dout(w_dff_B_qz9OmIKW8_2),.clk(gclk));
	jdff dff_B_sVK3HWJo8_2(.din(w_dff_B_qz9OmIKW8_2),.dout(w_dff_B_sVK3HWJo8_2),.clk(gclk));
	jdff dff_B_XIPQYJju6_2(.din(w_dff_B_sVK3HWJo8_2),.dout(w_dff_B_XIPQYJju6_2),.clk(gclk));
	jdff dff_B_9bFez3Sf8_2(.din(n696),.dout(w_dff_B_9bFez3Sf8_2),.clk(gclk));
	jdff dff_B_TNkzBPEQ1_1(.din(n633),.dout(w_dff_B_TNkzBPEQ1_1),.clk(gclk));
	jdff dff_B_bBhkbszQ7_2(.din(n547),.dout(w_dff_B_bBhkbszQ7_2),.clk(gclk));
	jdff dff_B_f51oMVeo7_2(.din(w_dff_B_bBhkbszQ7_2),.dout(w_dff_B_f51oMVeo7_2),.clk(gclk));
	jdff dff_B_UbNQtSth0_2(.din(w_dff_B_f51oMVeo7_2),.dout(w_dff_B_UbNQtSth0_2),.clk(gclk));
	jdff dff_B_FUkSvxAy3_2(.din(w_dff_B_UbNQtSth0_2),.dout(w_dff_B_FUkSvxAy3_2),.clk(gclk));
	jdff dff_B_win2S9aE0_2(.din(w_dff_B_FUkSvxAy3_2),.dout(w_dff_B_win2S9aE0_2),.clk(gclk));
	jdff dff_B_UmyW3qT50_2(.din(w_dff_B_win2S9aE0_2),.dout(w_dff_B_UmyW3qT50_2),.clk(gclk));
	jdff dff_B_yCmJTnyJ4_2(.din(w_dff_B_UmyW3qT50_2),.dout(w_dff_B_yCmJTnyJ4_2),.clk(gclk));
	jdff dff_B_Jt98ZZU86_2(.din(w_dff_B_yCmJTnyJ4_2),.dout(w_dff_B_Jt98ZZU86_2),.clk(gclk));
	jdff dff_B_HvsZa83H6_2(.din(w_dff_B_Jt98ZZU86_2),.dout(w_dff_B_HvsZa83H6_2),.clk(gclk));
	jdff dff_B_zTBHjKWh3_2(.din(w_dff_B_HvsZa83H6_2),.dout(w_dff_B_zTBHjKWh3_2),.clk(gclk));
	jdff dff_B_t5yXvKYO9_2(.din(w_dff_B_zTBHjKWh3_2),.dout(w_dff_B_t5yXvKYO9_2),.clk(gclk));
	jdff dff_B_0HdcgnmU9_2(.din(w_dff_B_t5yXvKYO9_2),.dout(w_dff_B_0HdcgnmU9_2),.clk(gclk));
	jdff dff_B_sijVBhM94_2(.din(w_dff_B_0HdcgnmU9_2),.dout(w_dff_B_sijVBhM94_2),.clk(gclk));
	jdff dff_B_1PSw7WPZ5_2(.din(w_dff_B_sijVBhM94_2),.dout(w_dff_B_1PSw7WPZ5_2),.clk(gclk));
	jdff dff_B_G2C2M3vD7_2(.din(w_dff_B_1PSw7WPZ5_2),.dout(w_dff_B_G2C2M3vD7_2),.clk(gclk));
	jdff dff_B_u4S8Nntb1_2(.din(w_dff_B_G2C2M3vD7_2),.dout(w_dff_B_u4S8Nntb1_2),.clk(gclk));
	jdff dff_B_QKMMQkka4_2(.din(w_dff_B_u4S8Nntb1_2),.dout(w_dff_B_QKMMQkka4_2),.clk(gclk));
	jdff dff_B_UQhP4lYA9_2(.din(w_dff_B_QKMMQkka4_2),.dout(w_dff_B_UQhP4lYA9_2),.clk(gclk));
	jdff dff_B_XeM8pS0B5_2(.din(w_dff_B_UQhP4lYA9_2),.dout(w_dff_B_XeM8pS0B5_2),.clk(gclk));
	jdff dff_B_6ZeRMQGd4_2(.din(w_dff_B_XeM8pS0B5_2),.dout(w_dff_B_6ZeRMQGd4_2),.clk(gclk));
	jdff dff_B_8kE73v0Q1_2(.din(w_dff_B_6ZeRMQGd4_2),.dout(w_dff_B_8kE73v0Q1_2),.clk(gclk));
	jdff dff_B_M9GYRtXm4_2(.din(w_dff_B_8kE73v0Q1_2),.dout(w_dff_B_M9GYRtXm4_2),.clk(gclk));
	jdff dff_B_MR0lnAsI3_2(.din(w_dff_B_M9GYRtXm4_2),.dout(w_dff_B_MR0lnAsI3_2),.clk(gclk));
	jdff dff_B_jw7L1Y4g3_2(.din(w_dff_B_MR0lnAsI3_2),.dout(w_dff_B_jw7L1Y4g3_2),.clk(gclk));
	jdff dff_B_fSPB99zU8_2(.din(n604),.dout(w_dff_B_fSPB99zU8_2),.clk(gclk));
	jdff dff_B_uYM3roB00_1(.din(n548),.dout(w_dff_B_uYM3roB00_1),.clk(gclk));
	jdff dff_B_UeJKjEuo2_2(.din(n469),.dout(w_dff_B_UeJKjEuo2_2),.clk(gclk));
	jdff dff_B_M7SsA64h8_2(.din(w_dff_B_UeJKjEuo2_2),.dout(w_dff_B_M7SsA64h8_2),.clk(gclk));
	jdff dff_B_Y3eAVrVf0_2(.din(w_dff_B_M7SsA64h8_2),.dout(w_dff_B_Y3eAVrVf0_2),.clk(gclk));
	jdff dff_B_oBiFGf9J4_2(.din(w_dff_B_Y3eAVrVf0_2),.dout(w_dff_B_oBiFGf9J4_2),.clk(gclk));
	jdff dff_B_CPFMDieT8_2(.din(w_dff_B_oBiFGf9J4_2),.dout(w_dff_B_CPFMDieT8_2),.clk(gclk));
	jdff dff_B_u7iQ1IHo5_2(.din(w_dff_B_CPFMDieT8_2),.dout(w_dff_B_u7iQ1IHo5_2),.clk(gclk));
	jdff dff_B_ndnpMWqP0_2(.din(w_dff_B_u7iQ1IHo5_2),.dout(w_dff_B_ndnpMWqP0_2),.clk(gclk));
	jdff dff_B_vEgA1lS38_2(.din(w_dff_B_ndnpMWqP0_2),.dout(w_dff_B_vEgA1lS38_2),.clk(gclk));
	jdff dff_B_bGn3YH7G4_2(.din(w_dff_B_vEgA1lS38_2),.dout(w_dff_B_bGn3YH7G4_2),.clk(gclk));
	jdff dff_B_ysUq4Td77_2(.din(w_dff_B_bGn3YH7G4_2),.dout(w_dff_B_ysUq4Td77_2),.clk(gclk));
	jdff dff_B_vE2VGbef5_2(.din(w_dff_B_ysUq4Td77_2),.dout(w_dff_B_vE2VGbef5_2),.clk(gclk));
	jdff dff_B_5Oiv5Ozn4_2(.din(w_dff_B_vE2VGbef5_2),.dout(w_dff_B_5Oiv5Ozn4_2),.clk(gclk));
	jdff dff_B_mdVkEO9y0_2(.din(w_dff_B_5Oiv5Ozn4_2),.dout(w_dff_B_mdVkEO9y0_2),.clk(gclk));
	jdff dff_B_G6DwSyC76_2(.din(w_dff_B_mdVkEO9y0_2),.dout(w_dff_B_G6DwSyC76_2),.clk(gclk));
	jdff dff_B_BACQ45Mw2_2(.din(w_dff_B_G6DwSyC76_2),.dout(w_dff_B_BACQ45Mw2_2),.clk(gclk));
	jdff dff_B_WVecvOpA4_2(.din(w_dff_B_BACQ45Mw2_2),.dout(w_dff_B_WVecvOpA4_2),.clk(gclk));
	jdff dff_B_qzelPbpo3_2(.din(w_dff_B_WVecvOpA4_2),.dout(w_dff_B_qzelPbpo3_2),.clk(gclk));
	jdff dff_B_y5X4O3hO9_2(.din(w_dff_B_qzelPbpo3_2),.dout(w_dff_B_y5X4O3hO9_2),.clk(gclk));
	jdff dff_B_AuuQ60UU6_2(.din(w_dff_B_y5X4O3hO9_2),.dout(w_dff_B_AuuQ60UU6_2),.clk(gclk));
	jdff dff_B_zkTDCxtL2_2(.din(w_dff_B_AuuQ60UU6_2),.dout(w_dff_B_zkTDCxtL2_2),.clk(gclk));
	jdff dff_B_v1qq48ab4_2(.din(w_dff_B_zkTDCxtL2_2),.dout(w_dff_B_v1qq48ab4_2),.clk(gclk));
	jdff dff_B_pYAEP80p8_2(.din(n519),.dout(w_dff_B_pYAEP80p8_2),.clk(gclk));
	jdff dff_B_mVu63OJQ1_1(.din(n470),.dout(w_dff_B_mVu63OJQ1_1),.clk(gclk));
	jdff dff_B_WEWxMx065_2(.din(n398),.dout(w_dff_B_WEWxMx065_2),.clk(gclk));
	jdff dff_B_W1hpzVyU6_2(.din(w_dff_B_WEWxMx065_2),.dout(w_dff_B_W1hpzVyU6_2),.clk(gclk));
	jdff dff_B_8I3CbCaA9_2(.din(w_dff_B_W1hpzVyU6_2),.dout(w_dff_B_8I3CbCaA9_2),.clk(gclk));
	jdff dff_B_AWocKXOg8_2(.din(w_dff_B_8I3CbCaA9_2),.dout(w_dff_B_AWocKXOg8_2),.clk(gclk));
	jdff dff_B_AIDr4X9M9_2(.din(w_dff_B_AWocKXOg8_2),.dout(w_dff_B_AIDr4X9M9_2),.clk(gclk));
	jdff dff_B_NaQCEV502_2(.din(w_dff_B_AIDr4X9M9_2),.dout(w_dff_B_NaQCEV502_2),.clk(gclk));
	jdff dff_B_e08tTMd56_2(.din(w_dff_B_NaQCEV502_2),.dout(w_dff_B_e08tTMd56_2),.clk(gclk));
	jdff dff_B_1IUHKHOh2_2(.din(w_dff_B_e08tTMd56_2),.dout(w_dff_B_1IUHKHOh2_2),.clk(gclk));
	jdff dff_B_WTpAsNU15_2(.din(w_dff_B_1IUHKHOh2_2),.dout(w_dff_B_WTpAsNU15_2),.clk(gclk));
	jdff dff_B_57uRIp4D6_2(.din(w_dff_B_WTpAsNU15_2),.dout(w_dff_B_57uRIp4D6_2),.clk(gclk));
	jdff dff_B_CCYEVUQR3_2(.din(w_dff_B_57uRIp4D6_2),.dout(w_dff_B_CCYEVUQR3_2),.clk(gclk));
	jdff dff_B_fTfVusa95_2(.din(w_dff_B_CCYEVUQR3_2),.dout(w_dff_B_fTfVusa95_2),.clk(gclk));
	jdff dff_B_K6ainE281_2(.din(w_dff_B_fTfVusa95_2),.dout(w_dff_B_K6ainE281_2),.clk(gclk));
	jdff dff_B_XaiHOww80_2(.din(w_dff_B_K6ainE281_2),.dout(w_dff_B_XaiHOww80_2),.clk(gclk));
	jdff dff_B_jTyFb9U55_2(.din(w_dff_B_XaiHOww80_2),.dout(w_dff_B_jTyFb9U55_2),.clk(gclk));
	jdff dff_B_2yqMtiOT6_2(.din(w_dff_B_jTyFb9U55_2),.dout(w_dff_B_2yqMtiOT6_2),.clk(gclk));
	jdff dff_B_q5bQKJu14_2(.din(w_dff_B_2yqMtiOT6_2),.dout(w_dff_B_q5bQKJu14_2),.clk(gclk));
	jdff dff_B_80hrZBpf0_2(.din(w_dff_B_q5bQKJu14_2),.dout(w_dff_B_80hrZBpf0_2),.clk(gclk));
	jdff dff_B_Dr1IrqGm8_2(.din(n441),.dout(w_dff_B_Dr1IrqGm8_2),.clk(gclk));
	jdff dff_B_0rCHEG0m8_1(.din(n399),.dout(w_dff_B_0rCHEG0m8_1),.clk(gclk));
	jdff dff_B_Ys6VVuGu3_2(.din(n335),.dout(w_dff_B_Ys6VVuGu3_2),.clk(gclk));
	jdff dff_B_0l6c51KU8_2(.din(w_dff_B_Ys6VVuGu3_2),.dout(w_dff_B_0l6c51KU8_2),.clk(gclk));
	jdff dff_B_Ty2zuga32_2(.din(w_dff_B_0l6c51KU8_2),.dout(w_dff_B_Ty2zuga32_2),.clk(gclk));
	jdff dff_B_uer5qByP8_2(.din(w_dff_B_Ty2zuga32_2),.dout(w_dff_B_uer5qByP8_2),.clk(gclk));
	jdff dff_B_byXUke3X7_2(.din(w_dff_B_uer5qByP8_2),.dout(w_dff_B_byXUke3X7_2),.clk(gclk));
	jdff dff_B_4EfWPXMY9_2(.din(w_dff_B_byXUke3X7_2),.dout(w_dff_B_4EfWPXMY9_2),.clk(gclk));
	jdff dff_B_iYbmjNtZ7_2(.din(w_dff_B_4EfWPXMY9_2),.dout(w_dff_B_iYbmjNtZ7_2),.clk(gclk));
	jdff dff_B_bvlS3ki57_2(.din(w_dff_B_iYbmjNtZ7_2),.dout(w_dff_B_bvlS3ki57_2),.clk(gclk));
	jdff dff_B_lezNhEqZ6_2(.din(w_dff_B_bvlS3ki57_2),.dout(w_dff_B_lezNhEqZ6_2),.clk(gclk));
	jdff dff_B_aMd4yMz06_2(.din(w_dff_B_lezNhEqZ6_2),.dout(w_dff_B_aMd4yMz06_2),.clk(gclk));
	jdff dff_B_7ixe8zJH6_2(.din(w_dff_B_aMd4yMz06_2),.dout(w_dff_B_7ixe8zJH6_2),.clk(gclk));
	jdff dff_B_yeDuCsWG2_2(.din(w_dff_B_7ixe8zJH6_2),.dout(w_dff_B_yeDuCsWG2_2),.clk(gclk));
	jdff dff_B_QMujZxw62_2(.din(w_dff_B_yeDuCsWG2_2),.dout(w_dff_B_QMujZxw62_2),.clk(gclk));
	jdff dff_B_Ubl8n52K2_2(.din(w_dff_B_QMujZxw62_2),.dout(w_dff_B_Ubl8n52K2_2),.clk(gclk));
	jdff dff_B_Nzc0jN0X6_2(.din(w_dff_B_Ubl8n52K2_2),.dout(w_dff_B_Nzc0jN0X6_2),.clk(gclk));
	jdff dff_B_ytpEQb7Q7_2(.din(n370),.dout(w_dff_B_ytpEQb7Q7_2),.clk(gclk));
	jdff dff_B_1rtVAh7u6_1(.din(n336),.dout(w_dff_B_1rtVAh7u6_1),.clk(gclk));
	jdff dff_B_omdEaLWk4_2(.din(n279),.dout(w_dff_B_omdEaLWk4_2),.clk(gclk));
	jdff dff_B_Fh3oMONb3_2(.din(w_dff_B_omdEaLWk4_2),.dout(w_dff_B_Fh3oMONb3_2),.clk(gclk));
	jdff dff_B_JaeHTARs5_2(.din(w_dff_B_Fh3oMONb3_2),.dout(w_dff_B_JaeHTARs5_2),.clk(gclk));
	jdff dff_B_arJq6s7v9_2(.din(w_dff_B_JaeHTARs5_2),.dout(w_dff_B_arJq6s7v9_2),.clk(gclk));
	jdff dff_B_RX7mPEjL1_2(.din(w_dff_B_arJq6s7v9_2),.dout(w_dff_B_RX7mPEjL1_2),.clk(gclk));
	jdff dff_B_bZ6rfMWN6_2(.din(w_dff_B_RX7mPEjL1_2),.dout(w_dff_B_bZ6rfMWN6_2),.clk(gclk));
	jdff dff_B_3wOjXPL01_2(.din(w_dff_B_bZ6rfMWN6_2),.dout(w_dff_B_3wOjXPL01_2),.clk(gclk));
	jdff dff_B_t9whI86T7_2(.din(w_dff_B_3wOjXPL01_2),.dout(w_dff_B_t9whI86T7_2),.clk(gclk));
	jdff dff_B_Rf099flr7_2(.din(w_dff_B_t9whI86T7_2),.dout(w_dff_B_Rf099flr7_2),.clk(gclk));
	jdff dff_B_kjx61lNX5_2(.din(w_dff_B_Rf099flr7_2),.dout(w_dff_B_kjx61lNX5_2),.clk(gclk));
	jdff dff_B_qlspWzHw1_2(.din(w_dff_B_kjx61lNX5_2),.dout(w_dff_B_qlspWzHw1_2),.clk(gclk));
	jdff dff_B_czwAcrTA5_2(.din(w_dff_B_qlspWzHw1_2),.dout(w_dff_B_czwAcrTA5_2),.clk(gclk));
	jdff dff_B_Xt3SxkYc6_2(.din(n307),.dout(w_dff_B_Xt3SxkYc6_2),.clk(gclk));
	jdff dff_B_P2mKMjuP8_1(.din(n280),.dout(w_dff_B_P2mKMjuP8_1),.clk(gclk));
	jdff dff_B_5TdOO4dZ3_2(.din(n230),.dout(w_dff_B_5TdOO4dZ3_2),.clk(gclk));
	jdff dff_B_3FucluDd3_2(.din(w_dff_B_5TdOO4dZ3_2),.dout(w_dff_B_3FucluDd3_2),.clk(gclk));
	jdff dff_B_fgDT3QRk3_2(.din(w_dff_B_3FucluDd3_2),.dout(w_dff_B_fgDT3QRk3_2),.clk(gclk));
	jdff dff_B_UGXTrXMM9_2(.din(w_dff_B_fgDT3QRk3_2),.dout(w_dff_B_UGXTrXMM9_2),.clk(gclk));
	jdff dff_B_pj5D2l2T3_2(.din(w_dff_B_UGXTrXMM9_2),.dout(w_dff_B_pj5D2l2T3_2),.clk(gclk));
	jdff dff_B_cVccoivS0_2(.din(w_dff_B_pj5D2l2T3_2),.dout(w_dff_B_cVccoivS0_2),.clk(gclk));
	jdff dff_B_2evKtaZu4_2(.din(w_dff_B_cVccoivS0_2),.dout(w_dff_B_2evKtaZu4_2),.clk(gclk));
	jdff dff_B_W6vCpGoW6_2(.din(w_dff_B_2evKtaZu4_2),.dout(w_dff_B_W6vCpGoW6_2),.clk(gclk));
	jdff dff_B_dQEcMFM43_2(.din(w_dff_B_W6vCpGoW6_2),.dout(w_dff_B_dQEcMFM43_2),.clk(gclk));
	jdff dff_B_VFWvjV9t5_2(.din(n251),.dout(w_dff_B_VFWvjV9t5_2),.clk(gclk));
	jdff dff_B_Zm1aESKy2_1(.din(n231),.dout(w_dff_B_Zm1aESKy2_1),.clk(gclk));
	jdff dff_B_nd94F0Wh0_2(.din(n188),.dout(w_dff_B_nd94F0Wh0_2),.clk(gclk));
	jdff dff_B_GfGcW0iz2_2(.din(w_dff_B_nd94F0Wh0_2),.dout(w_dff_B_GfGcW0iz2_2),.clk(gclk));
	jdff dff_B_8umv0ypU0_2(.din(w_dff_B_GfGcW0iz2_2),.dout(w_dff_B_8umv0ypU0_2),.clk(gclk));
	jdff dff_B_NF4kGozM3_2(.din(w_dff_B_8umv0ypU0_2),.dout(w_dff_B_NF4kGozM3_2),.clk(gclk));
	jdff dff_B_a0SR0zze2_2(.din(w_dff_B_NF4kGozM3_2),.dout(w_dff_B_a0SR0zze2_2),.clk(gclk));
	jdff dff_B_kLH7gl653_2(.din(w_dff_B_a0SR0zze2_2),.dout(w_dff_B_kLH7gl653_2),.clk(gclk));
	jdff dff_B_k8KuEIIu9_2(.din(n202),.dout(w_dff_B_k8KuEIIu9_2),.clk(gclk));
	jdff dff_B_SLOUeJJZ0_2(.din(n154),.dout(w_dff_B_SLOUeJJZ0_2),.clk(gclk));
	jdff dff_B_UMrwSk2E5_2(.din(w_dff_B_SLOUeJJZ0_2),.dout(w_dff_B_UMrwSk2E5_2),.clk(gclk));
	jdff dff_B_ICAcvj6l7_2(.din(w_dff_B_UMrwSk2E5_2),.dout(w_dff_B_ICAcvj6l7_2),.clk(gclk));
	jdff dff_B_fGZCObuk2_0(.din(n159),.dout(w_dff_B_fGZCObuk2_0),.clk(gclk));
	jdff dff_A_CuJghATl4_0(.dout(w_n123_0[0]),.din(w_dff_A_CuJghATl4_0),.clk(gclk));
	jdff dff_A_2DFVxxTq9_0(.dout(w_dff_A_CuJghATl4_0),.din(w_dff_A_2DFVxxTq9_0),.clk(gclk));
	jdff dff_A_FEWmkBeV4_0(.dout(w_n122_0[0]),.din(w_dff_A_FEWmkBeV4_0),.clk(gclk));
	jdff dff_A_dYnoKGBq0_0(.dout(w_dff_A_FEWmkBeV4_0),.din(w_dff_A_dYnoKGBq0_0),.clk(gclk));
	jdff dff_B_SgiYHoB16_1(.din(n1304),.dout(w_dff_B_SgiYHoB16_1),.clk(gclk));
	jdff dff_B_PuYXf8Yd1_2(.din(n1217),.dout(w_dff_B_PuYXf8Yd1_2),.clk(gclk));
	jdff dff_B_mT5LsNOh5_2(.din(w_dff_B_PuYXf8Yd1_2),.dout(w_dff_B_mT5LsNOh5_2),.clk(gclk));
	jdff dff_B_obQNMcPx1_2(.din(w_dff_B_mT5LsNOh5_2),.dout(w_dff_B_obQNMcPx1_2),.clk(gclk));
	jdff dff_B_ZOnShia50_2(.din(w_dff_B_obQNMcPx1_2),.dout(w_dff_B_ZOnShia50_2),.clk(gclk));
	jdff dff_B_y2vvH2jy3_2(.din(w_dff_B_ZOnShia50_2),.dout(w_dff_B_y2vvH2jy3_2),.clk(gclk));
	jdff dff_B_rwc7ZNq40_2(.din(w_dff_B_y2vvH2jy3_2),.dout(w_dff_B_rwc7ZNq40_2),.clk(gclk));
	jdff dff_B_1qeFN1HJ1_2(.din(w_dff_B_rwc7ZNq40_2),.dout(w_dff_B_1qeFN1HJ1_2),.clk(gclk));
	jdff dff_B_R9MTpE0L0_2(.din(w_dff_B_1qeFN1HJ1_2),.dout(w_dff_B_R9MTpE0L0_2),.clk(gclk));
	jdff dff_B_hh7WYfYd2_2(.din(w_dff_B_R9MTpE0L0_2),.dout(w_dff_B_hh7WYfYd2_2),.clk(gclk));
	jdff dff_B_scUmfuoJ4_2(.din(w_dff_B_hh7WYfYd2_2),.dout(w_dff_B_scUmfuoJ4_2),.clk(gclk));
	jdff dff_B_ebbtcAO11_2(.din(w_dff_B_scUmfuoJ4_2),.dout(w_dff_B_ebbtcAO11_2),.clk(gclk));
	jdff dff_B_NbCVchy23_2(.din(w_dff_B_ebbtcAO11_2),.dout(w_dff_B_NbCVchy23_2),.clk(gclk));
	jdff dff_B_56TI56UR8_2(.din(w_dff_B_NbCVchy23_2),.dout(w_dff_B_56TI56UR8_2),.clk(gclk));
	jdff dff_B_ffRliSXe4_2(.din(w_dff_B_56TI56UR8_2),.dout(w_dff_B_ffRliSXe4_2),.clk(gclk));
	jdff dff_B_cFjqFrom6_2(.din(w_dff_B_ffRliSXe4_2),.dout(w_dff_B_cFjqFrom6_2),.clk(gclk));
	jdff dff_B_h3Z3iue59_2(.din(w_dff_B_cFjqFrom6_2),.dout(w_dff_B_h3Z3iue59_2),.clk(gclk));
	jdff dff_B_9Zyd006o1_2(.din(w_dff_B_h3Z3iue59_2),.dout(w_dff_B_9Zyd006o1_2),.clk(gclk));
	jdff dff_B_EQsHucWM1_2(.din(w_dff_B_9Zyd006o1_2),.dout(w_dff_B_EQsHucWM1_2),.clk(gclk));
	jdff dff_B_sWCLstXV1_2(.din(w_dff_B_EQsHucWM1_2),.dout(w_dff_B_sWCLstXV1_2),.clk(gclk));
	jdff dff_B_Gfgy7tTz8_2(.din(w_dff_B_sWCLstXV1_2),.dout(w_dff_B_Gfgy7tTz8_2),.clk(gclk));
	jdff dff_B_Twyo5fVA9_2(.din(w_dff_B_Gfgy7tTz8_2),.dout(w_dff_B_Twyo5fVA9_2),.clk(gclk));
	jdff dff_B_gPVriFN42_2(.din(w_dff_B_Twyo5fVA9_2),.dout(w_dff_B_gPVriFN42_2),.clk(gclk));
	jdff dff_B_nmfKnA3F9_2(.din(w_dff_B_gPVriFN42_2),.dout(w_dff_B_nmfKnA3F9_2),.clk(gclk));
	jdff dff_B_K3HZopTd8_2(.din(w_dff_B_nmfKnA3F9_2),.dout(w_dff_B_K3HZopTd8_2),.clk(gclk));
	jdff dff_B_Bya0IkSZ6_2(.din(w_dff_B_K3HZopTd8_2),.dout(w_dff_B_Bya0IkSZ6_2),.clk(gclk));
	jdff dff_B_WAHDLpkr5_2(.din(w_dff_B_Bya0IkSZ6_2),.dout(w_dff_B_WAHDLpkr5_2),.clk(gclk));
	jdff dff_B_oJq5gcAZ4_2(.din(w_dff_B_WAHDLpkr5_2),.dout(w_dff_B_oJq5gcAZ4_2),.clk(gclk));
	jdff dff_B_GdhzBQ3w5_2(.din(w_dff_B_oJq5gcAZ4_2),.dout(w_dff_B_GdhzBQ3w5_2),.clk(gclk));
	jdff dff_B_PvTZaMme2_2(.din(w_dff_B_GdhzBQ3w5_2),.dout(w_dff_B_PvTZaMme2_2),.clk(gclk));
	jdff dff_B_qkbJ1AV54_2(.din(w_dff_B_PvTZaMme2_2),.dout(w_dff_B_qkbJ1AV54_2),.clk(gclk));
	jdff dff_B_3EWBsshh3_2(.din(w_dff_B_qkbJ1AV54_2),.dout(w_dff_B_3EWBsshh3_2),.clk(gclk));
	jdff dff_B_mmDfA33w9_2(.din(w_dff_B_3EWBsshh3_2),.dout(w_dff_B_mmDfA33w9_2),.clk(gclk));
	jdff dff_B_EIMOwjdg0_2(.din(w_dff_B_mmDfA33w9_2),.dout(w_dff_B_EIMOwjdg0_2),.clk(gclk));
	jdff dff_B_8Hfq9vft5_2(.din(w_dff_B_EIMOwjdg0_2),.dout(w_dff_B_8Hfq9vft5_2),.clk(gclk));
	jdff dff_B_zXPFMKne4_2(.din(w_dff_B_8Hfq9vft5_2),.dout(w_dff_B_zXPFMKne4_2),.clk(gclk));
	jdff dff_B_4L7NdiLb8_2(.din(w_dff_B_zXPFMKne4_2),.dout(w_dff_B_4L7NdiLb8_2),.clk(gclk));
	jdff dff_B_KeuXjNNN3_2(.din(w_dff_B_4L7NdiLb8_2),.dout(w_dff_B_KeuXjNNN3_2),.clk(gclk));
	jdff dff_B_85JFOAv87_2(.din(w_dff_B_KeuXjNNN3_2),.dout(w_dff_B_85JFOAv87_2),.clk(gclk));
	jdff dff_B_MMZQH4u04_2(.din(w_dff_B_85JFOAv87_2),.dout(w_dff_B_MMZQH4u04_2),.clk(gclk));
	jdff dff_B_ohZ8VlNI6_2(.din(w_dff_B_MMZQH4u04_2),.dout(w_dff_B_ohZ8VlNI6_2),.clk(gclk));
	jdff dff_B_hcpIuflp3_2(.din(w_dff_B_ohZ8VlNI6_2),.dout(w_dff_B_hcpIuflp3_2),.clk(gclk));
	jdff dff_B_jLzE5Uwv9_2(.din(w_dff_B_hcpIuflp3_2),.dout(w_dff_B_jLzE5Uwv9_2),.clk(gclk));
	jdff dff_B_AN0KKKPE5_2(.din(w_dff_B_jLzE5Uwv9_2),.dout(w_dff_B_AN0KKKPE5_2),.clk(gclk));
	jdff dff_B_plw1eKCA3_2(.din(w_dff_B_AN0KKKPE5_2),.dout(w_dff_B_plw1eKCA3_2),.clk(gclk));
	jdff dff_B_WbgLpl9P7_0(.din(n1303),.dout(w_dff_B_WbgLpl9P7_0),.clk(gclk));
	jdff dff_A_o830kju60_1(.dout(w_n1291_0[1]),.din(w_dff_A_o830kju60_1),.clk(gclk));
	jdff dff_B_I4hnYSxQ2_1(.din(n1218),.dout(w_dff_B_I4hnYSxQ2_1),.clk(gclk));
	jdff dff_B_jkJaKtAo0_2(.din(n1126),.dout(w_dff_B_jkJaKtAo0_2),.clk(gclk));
	jdff dff_B_4ItMHm427_2(.din(w_dff_B_jkJaKtAo0_2),.dout(w_dff_B_4ItMHm427_2),.clk(gclk));
	jdff dff_B_nbYo9Rx48_2(.din(w_dff_B_4ItMHm427_2),.dout(w_dff_B_nbYo9Rx48_2),.clk(gclk));
	jdff dff_B_OwOa3Pot5_2(.din(w_dff_B_nbYo9Rx48_2),.dout(w_dff_B_OwOa3Pot5_2),.clk(gclk));
	jdff dff_B_f6MlyqXb1_2(.din(w_dff_B_OwOa3Pot5_2),.dout(w_dff_B_f6MlyqXb1_2),.clk(gclk));
	jdff dff_B_pzHWvknQ4_2(.din(w_dff_B_f6MlyqXb1_2),.dout(w_dff_B_pzHWvknQ4_2),.clk(gclk));
	jdff dff_B_AYkK0VcL3_2(.din(w_dff_B_pzHWvknQ4_2),.dout(w_dff_B_AYkK0VcL3_2),.clk(gclk));
	jdff dff_B_f7hrnO3D2_2(.din(w_dff_B_AYkK0VcL3_2),.dout(w_dff_B_f7hrnO3D2_2),.clk(gclk));
	jdff dff_B_4daHqpxM2_2(.din(w_dff_B_f7hrnO3D2_2),.dout(w_dff_B_4daHqpxM2_2),.clk(gclk));
	jdff dff_B_ltOzQgEJ4_2(.din(w_dff_B_4daHqpxM2_2),.dout(w_dff_B_ltOzQgEJ4_2),.clk(gclk));
	jdff dff_B_vjG45HXm3_2(.din(w_dff_B_ltOzQgEJ4_2),.dout(w_dff_B_vjG45HXm3_2),.clk(gclk));
	jdff dff_B_m2FoSgTj2_2(.din(w_dff_B_vjG45HXm3_2),.dout(w_dff_B_m2FoSgTj2_2),.clk(gclk));
	jdff dff_B_GEVloQc47_2(.din(w_dff_B_m2FoSgTj2_2),.dout(w_dff_B_GEVloQc47_2),.clk(gclk));
	jdff dff_B_B1ngRcMq1_2(.din(w_dff_B_GEVloQc47_2),.dout(w_dff_B_B1ngRcMq1_2),.clk(gclk));
	jdff dff_B_Zqxf87DJ3_2(.din(w_dff_B_B1ngRcMq1_2),.dout(w_dff_B_Zqxf87DJ3_2),.clk(gclk));
	jdff dff_B_qey6le2O2_2(.din(w_dff_B_Zqxf87DJ3_2),.dout(w_dff_B_qey6le2O2_2),.clk(gclk));
	jdff dff_B_8zS87Lyn8_2(.din(w_dff_B_qey6le2O2_2),.dout(w_dff_B_8zS87Lyn8_2),.clk(gclk));
	jdff dff_B_pbCY08Ci3_2(.din(w_dff_B_8zS87Lyn8_2),.dout(w_dff_B_pbCY08Ci3_2),.clk(gclk));
	jdff dff_B_vCleocnw7_2(.din(w_dff_B_pbCY08Ci3_2),.dout(w_dff_B_vCleocnw7_2),.clk(gclk));
	jdff dff_B_kgVGb8NU2_2(.din(w_dff_B_vCleocnw7_2),.dout(w_dff_B_kgVGb8NU2_2),.clk(gclk));
	jdff dff_B_Nh1Yluc92_2(.din(w_dff_B_kgVGb8NU2_2),.dout(w_dff_B_Nh1Yluc92_2),.clk(gclk));
	jdff dff_B_XidOhPvE0_2(.din(w_dff_B_Nh1Yluc92_2),.dout(w_dff_B_XidOhPvE0_2),.clk(gclk));
	jdff dff_B_roFGmJYq1_2(.din(w_dff_B_XidOhPvE0_2),.dout(w_dff_B_roFGmJYq1_2),.clk(gclk));
	jdff dff_B_oR6ruBum6_2(.din(w_dff_B_roFGmJYq1_2),.dout(w_dff_B_oR6ruBum6_2),.clk(gclk));
	jdff dff_B_mnmNpu8t1_2(.din(w_dff_B_oR6ruBum6_2),.dout(w_dff_B_mnmNpu8t1_2),.clk(gclk));
	jdff dff_B_OO6yCJeh7_2(.din(w_dff_B_mnmNpu8t1_2),.dout(w_dff_B_OO6yCJeh7_2),.clk(gclk));
	jdff dff_B_I1ZZlWbr4_2(.din(w_dff_B_OO6yCJeh7_2),.dout(w_dff_B_I1ZZlWbr4_2),.clk(gclk));
	jdff dff_B_OOZZYZsv6_2(.din(w_dff_B_I1ZZlWbr4_2),.dout(w_dff_B_OOZZYZsv6_2),.clk(gclk));
	jdff dff_B_JnnT4mFj7_2(.din(w_dff_B_OOZZYZsv6_2),.dout(w_dff_B_JnnT4mFj7_2),.clk(gclk));
	jdff dff_B_NjwGDvfe4_2(.din(w_dff_B_JnnT4mFj7_2),.dout(w_dff_B_NjwGDvfe4_2),.clk(gclk));
	jdff dff_B_IvMc5iTh9_2(.din(w_dff_B_NjwGDvfe4_2),.dout(w_dff_B_IvMc5iTh9_2),.clk(gclk));
	jdff dff_B_90Vlik5A7_2(.din(w_dff_B_IvMc5iTh9_2),.dout(w_dff_B_90Vlik5A7_2),.clk(gclk));
	jdff dff_B_zj6kbofr7_2(.din(w_dff_B_90Vlik5A7_2),.dout(w_dff_B_zj6kbofr7_2),.clk(gclk));
	jdff dff_B_yPn4o7ol5_2(.din(w_dff_B_zj6kbofr7_2),.dout(w_dff_B_yPn4o7ol5_2),.clk(gclk));
	jdff dff_B_Bk4DPF6d4_2(.din(w_dff_B_yPn4o7ol5_2),.dout(w_dff_B_Bk4DPF6d4_2),.clk(gclk));
	jdff dff_B_QuiMGWJ42_2(.din(w_dff_B_Bk4DPF6d4_2),.dout(w_dff_B_QuiMGWJ42_2),.clk(gclk));
	jdff dff_B_pqmtBimK2_2(.din(w_dff_B_QuiMGWJ42_2),.dout(w_dff_B_pqmtBimK2_2),.clk(gclk));
	jdff dff_B_YHPlKlE47_2(.din(w_dff_B_pqmtBimK2_2),.dout(w_dff_B_YHPlKlE47_2),.clk(gclk));
	jdff dff_B_CofvUyBV3_2(.din(w_dff_B_YHPlKlE47_2),.dout(w_dff_B_CofvUyBV3_2),.clk(gclk));
	jdff dff_B_aV33VNxI7_2(.din(n1200),.dout(w_dff_B_aV33VNxI7_2),.clk(gclk));
	jdff dff_B_Y31JGknQ3_1(.din(n1127),.dout(w_dff_B_Y31JGknQ3_1),.clk(gclk));
	jdff dff_B_acpUoPty5_2(.din(n1028),.dout(w_dff_B_acpUoPty5_2),.clk(gclk));
	jdff dff_B_96J8h7BX2_2(.din(w_dff_B_acpUoPty5_2),.dout(w_dff_B_96J8h7BX2_2),.clk(gclk));
	jdff dff_B_QTJ77WGC4_2(.din(w_dff_B_96J8h7BX2_2),.dout(w_dff_B_QTJ77WGC4_2),.clk(gclk));
	jdff dff_B_ZnDgHNso0_2(.din(w_dff_B_QTJ77WGC4_2),.dout(w_dff_B_ZnDgHNso0_2),.clk(gclk));
	jdff dff_B_AqUB1R5v8_2(.din(w_dff_B_ZnDgHNso0_2),.dout(w_dff_B_AqUB1R5v8_2),.clk(gclk));
	jdff dff_B_wMyLZpig5_2(.din(w_dff_B_AqUB1R5v8_2),.dout(w_dff_B_wMyLZpig5_2),.clk(gclk));
	jdff dff_B_TBntwDWV4_2(.din(w_dff_B_wMyLZpig5_2),.dout(w_dff_B_TBntwDWV4_2),.clk(gclk));
	jdff dff_B_1WpHUZwh8_2(.din(w_dff_B_TBntwDWV4_2),.dout(w_dff_B_1WpHUZwh8_2),.clk(gclk));
	jdff dff_B_DpheNZBm7_2(.din(w_dff_B_1WpHUZwh8_2),.dout(w_dff_B_DpheNZBm7_2),.clk(gclk));
	jdff dff_B_iIcWVjQf7_2(.din(w_dff_B_DpheNZBm7_2),.dout(w_dff_B_iIcWVjQf7_2),.clk(gclk));
	jdff dff_B_uiRjDFcL5_2(.din(w_dff_B_iIcWVjQf7_2),.dout(w_dff_B_uiRjDFcL5_2),.clk(gclk));
	jdff dff_B_DL4b7u6b4_2(.din(w_dff_B_uiRjDFcL5_2),.dout(w_dff_B_DL4b7u6b4_2),.clk(gclk));
	jdff dff_B_AE5YTbSh3_2(.din(w_dff_B_DL4b7u6b4_2),.dout(w_dff_B_AE5YTbSh3_2),.clk(gclk));
	jdff dff_B_o0WHDeI58_2(.din(w_dff_B_AE5YTbSh3_2),.dout(w_dff_B_o0WHDeI58_2),.clk(gclk));
	jdff dff_B_GTZxZd5X6_2(.din(w_dff_B_o0WHDeI58_2),.dout(w_dff_B_GTZxZd5X6_2),.clk(gclk));
	jdff dff_B_NMJEzIe59_2(.din(w_dff_B_GTZxZd5X6_2),.dout(w_dff_B_NMJEzIe59_2),.clk(gclk));
	jdff dff_B_1QPbR1Ov9_2(.din(w_dff_B_NMJEzIe59_2),.dout(w_dff_B_1QPbR1Ov9_2),.clk(gclk));
	jdff dff_B_ztOrIbZr8_2(.din(w_dff_B_1QPbR1Ov9_2),.dout(w_dff_B_ztOrIbZr8_2),.clk(gclk));
	jdff dff_B_xrd6LqJy1_2(.din(w_dff_B_ztOrIbZr8_2),.dout(w_dff_B_xrd6LqJy1_2),.clk(gclk));
	jdff dff_B_dqkQ0NaF9_2(.din(w_dff_B_xrd6LqJy1_2),.dout(w_dff_B_dqkQ0NaF9_2),.clk(gclk));
	jdff dff_B_w7AlJqd71_2(.din(w_dff_B_dqkQ0NaF9_2),.dout(w_dff_B_w7AlJqd71_2),.clk(gclk));
	jdff dff_B_dhmztLHM5_2(.din(w_dff_B_w7AlJqd71_2),.dout(w_dff_B_dhmztLHM5_2),.clk(gclk));
	jdff dff_B_itzEVHu35_2(.din(w_dff_B_dhmztLHM5_2),.dout(w_dff_B_itzEVHu35_2),.clk(gclk));
	jdff dff_B_La0OAicv8_2(.din(w_dff_B_itzEVHu35_2),.dout(w_dff_B_La0OAicv8_2),.clk(gclk));
	jdff dff_B_VaBO4oAj2_2(.din(w_dff_B_La0OAicv8_2),.dout(w_dff_B_VaBO4oAj2_2),.clk(gclk));
	jdff dff_B_wYfqkKbE4_2(.din(w_dff_B_VaBO4oAj2_2),.dout(w_dff_B_wYfqkKbE4_2),.clk(gclk));
	jdff dff_B_6UegZdvZ1_2(.din(w_dff_B_wYfqkKbE4_2),.dout(w_dff_B_6UegZdvZ1_2),.clk(gclk));
	jdff dff_B_a1QEd8z56_2(.din(w_dff_B_6UegZdvZ1_2),.dout(w_dff_B_a1QEd8z56_2),.clk(gclk));
	jdff dff_B_93QEYQGl0_2(.din(w_dff_B_a1QEd8z56_2),.dout(w_dff_B_93QEYQGl0_2),.clk(gclk));
	jdff dff_B_gbaybP8j8_2(.din(w_dff_B_93QEYQGl0_2),.dout(w_dff_B_gbaybP8j8_2),.clk(gclk));
	jdff dff_B_60rFZjMu3_2(.din(w_dff_B_gbaybP8j8_2),.dout(w_dff_B_60rFZjMu3_2),.clk(gclk));
	jdff dff_B_BtUXjWQK2_2(.din(w_dff_B_60rFZjMu3_2),.dout(w_dff_B_BtUXjWQK2_2),.clk(gclk));
	jdff dff_B_hxDe64Qy8_2(.din(w_dff_B_BtUXjWQK2_2),.dout(w_dff_B_hxDe64Qy8_2),.clk(gclk));
	jdff dff_B_4nKzpZvV9_2(.din(w_dff_B_hxDe64Qy8_2),.dout(w_dff_B_4nKzpZvV9_2),.clk(gclk));
	jdff dff_B_oO3i39ic0_2(.din(w_dff_B_4nKzpZvV9_2),.dout(w_dff_B_oO3i39ic0_2),.clk(gclk));
	jdff dff_B_yCfDalDw2_2(.din(w_dff_B_oO3i39ic0_2),.dout(w_dff_B_yCfDalDw2_2),.clk(gclk));
	jdff dff_B_bXXrmGpH8_2(.din(n1101),.dout(w_dff_B_bXXrmGpH8_2),.clk(gclk));
	jdff dff_B_ldSAnnHy2_1(.din(n1029),.dout(w_dff_B_ldSAnnHy2_1),.clk(gclk));
	jdff dff_B_EilGpvvI0_2(.din(n929),.dout(w_dff_B_EilGpvvI0_2),.clk(gclk));
	jdff dff_B_1IqsQON04_2(.din(w_dff_B_EilGpvvI0_2),.dout(w_dff_B_1IqsQON04_2),.clk(gclk));
	jdff dff_B_PiDytZrV8_2(.din(w_dff_B_1IqsQON04_2),.dout(w_dff_B_PiDytZrV8_2),.clk(gclk));
	jdff dff_B_Vz7i4SA42_2(.din(w_dff_B_PiDytZrV8_2),.dout(w_dff_B_Vz7i4SA42_2),.clk(gclk));
	jdff dff_B_bKIarbmF4_2(.din(w_dff_B_Vz7i4SA42_2),.dout(w_dff_B_bKIarbmF4_2),.clk(gclk));
	jdff dff_B_6feI2gmN2_2(.din(w_dff_B_bKIarbmF4_2),.dout(w_dff_B_6feI2gmN2_2),.clk(gclk));
	jdff dff_B_K6i8BFwL1_2(.din(w_dff_B_6feI2gmN2_2),.dout(w_dff_B_K6i8BFwL1_2),.clk(gclk));
	jdff dff_B_lIX68ivf3_2(.din(w_dff_B_K6i8BFwL1_2),.dout(w_dff_B_lIX68ivf3_2),.clk(gclk));
	jdff dff_B_IN3iCCek4_2(.din(w_dff_B_lIX68ivf3_2),.dout(w_dff_B_IN3iCCek4_2),.clk(gclk));
	jdff dff_B_GEDQd7rQ3_2(.din(w_dff_B_IN3iCCek4_2),.dout(w_dff_B_GEDQd7rQ3_2),.clk(gclk));
	jdff dff_B_xiuvo8em2_2(.din(w_dff_B_GEDQd7rQ3_2),.dout(w_dff_B_xiuvo8em2_2),.clk(gclk));
	jdff dff_B_N615QvB30_2(.din(w_dff_B_xiuvo8em2_2),.dout(w_dff_B_N615QvB30_2),.clk(gclk));
	jdff dff_B_lLhgY6Ha1_2(.din(w_dff_B_N615QvB30_2),.dout(w_dff_B_lLhgY6Ha1_2),.clk(gclk));
	jdff dff_B_9lCWDov90_2(.din(w_dff_B_lLhgY6Ha1_2),.dout(w_dff_B_9lCWDov90_2),.clk(gclk));
	jdff dff_B_lyH64LUT2_2(.din(w_dff_B_9lCWDov90_2),.dout(w_dff_B_lyH64LUT2_2),.clk(gclk));
	jdff dff_B_Dos7dgYF2_2(.din(w_dff_B_lyH64LUT2_2),.dout(w_dff_B_Dos7dgYF2_2),.clk(gclk));
	jdff dff_B_HMlrJCcl6_2(.din(w_dff_B_Dos7dgYF2_2),.dout(w_dff_B_HMlrJCcl6_2),.clk(gclk));
	jdff dff_B_3pc51oFf7_2(.din(w_dff_B_HMlrJCcl6_2),.dout(w_dff_B_3pc51oFf7_2),.clk(gclk));
	jdff dff_B_HGvxUgeN8_2(.din(w_dff_B_3pc51oFf7_2),.dout(w_dff_B_HGvxUgeN8_2),.clk(gclk));
	jdff dff_B_sLTAmdti4_2(.din(w_dff_B_HGvxUgeN8_2),.dout(w_dff_B_sLTAmdti4_2),.clk(gclk));
	jdff dff_B_KNDHTW5v0_2(.din(w_dff_B_sLTAmdti4_2),.dout(w_dff_B_KNDHTW5v0_2),.clk(gclk));
	jdff dff_B_SdOVWn6m8_2(.din(w_dff_B_KNDHTW5v0_2),.dout(w_dff_B_SdOVWn6m8_2),.clk(gclk));
	jdff dff_B_x18VzERf0_2(.din(w_dff_B_SdOVWn6m8_2),.dout(w_dff_B_x18VzERf0_2),.clk(gclk));
	jdff dff_B_Z8oWQsmm0_2(.din(w_dff_B_x18VzERf0_2),.dout(w_dff_B_Z8oWQsmm0_2),.clk(gclk));
	jdff dff_B_YIvHtBNZ3_2(.din(w_dff_B_Z8oWQsmm0_2),.dout(w_dff_B_YIvHtBNZ3_2),.clk(gclk));
	jdff dff_B_CQnVwUjY2_2(.din(w_dff_B_YIvHtBNZ3_2),.dout(w_dff_B_CQnVwUjY2_2),.clk(gclk));
	jdff dff_B_p0BB09JE1_2(.din(w_dff_B_CQnVwUjY2_2),.dout(w_dff_B_p0BB09JE1_2),.clk(gclk));
	jdff dff_B_BU6hNa6v8_2(.din(w_dff_B_p0BB09JE1_2),.dout(w_dff_B_BU6hNa6v8_2),.clk(gclk));
	jdff dff_B_JIHRhzCk2_2(.din(w_dff_B_BU6hNa6v8_2),.dout(w_dff_B_JIHRhzCk2_2),.clk(gclk));
	jdff dff_B_Gru3oGwW4_2(.din(w_dff_B_JIHRhzCk2_2),.dout(w_dff_B_Gru3oGwW4_2),.clk(gclk));
	jdff dff_B_Oe2IoQmu2_2(.din(w_dff_B_Gru3oGwW4_2),.dout(w_dff_B_Oe2IoQmu2_2),.clk(gclk));
	jdff dff_B_QdykN0272_2(.din(w_dff_B_Oe2IoQmu2_2),.dout(w_dff_B_QdykN0272_2),.clk(gclk));
	jdff dff_B_XIQ0wdDi2_2(.din(w_dff_B_QdykN0272_2),.dout(w_dff_B_XIQ0wdDi2_2),.clk(gclk));
	jdff dff_B_hPP1DsNg0_2(.din(n1002),.dout(w_dff_B_hPP1DsNg0_2),.clk(gclk));
	jdff dff_B_E7UF84ec7_1(.din(n930),.dout(w_dff_B_E7UF84ec7_1),.clk(gclk));
	jdff dff_B_JJUTEcV79_2(.din(n827),.dout(w_dff_B_JJUTEcV79_2),.clk(gclk));
	jdff dff_B_wb95uZfJ7_2(.din(w_dff_B_JJUTEcV79_2),.dout(w_dff_B_wb95uZfJ7_2),.clk(gclk));
	jdff dff_B_LJKsoh0a8_2(.din(w_dff_B_wb95uZfJ7_2),.dout(w_dff_B_LJKsoh0a8_2),.clk(gclk));
	jdff dff_B_WQ639usY2_2(.din(w_dff_B_LJKsoh0a8_2),.dout(w_dff_B_WQ639usY2_2),.clk(gclk));
	jdff dff_B_khqkRhgq6_2(.din(w_dff_B_WQ639usY2_2),.dout(w_dff_B_khqkRhgq6_2),.clk(gclk));
	jdff dff_B_N4a7jGat6_2(.din(w_dff_B_khqkRhgq6_2),.dout(w_dff_B_N4a7jGat6_2),.clk(gclk));
	jdff dff_B_9SDLVzEy2_2(.din(w_dff_B_N4a7jGat6_2),.dout(w_dff_B_9SDLVzEy2_2),.clk(gclk));
	jdff dff_B_UlAGNrpR5_2(.din(w_dff_B_9SDLVzEy2_2),.dout(w_dff_B_UlAGNrpR5_2),.clk(gclk));
	jdff dff_B_m6luanHx8_2(.din(w_dff_B_UlAGNrpR5_2),.dout(w_dff_B_m6luanHx8_2),.clk(gclk));
	jdff dff_B_3KTBzRWX9_2(.din(w_dff_B_m6luanHx8_2),.dout(w_dff_B_3KTBzRWX9_2),.clk(gclk));
	jdff dff_B_00DuwbEL3_2(.din(w_dff_B_3KTBzRWX9_2),.dout(w_dff_B_00DuwbEL3_2),.clk(gclk));
	jdff dff_B_oNuoyF3A7_2(.din(w_dff_B_00DuwbEL3_2),.dout(w_dff_B_oNuoyF3A7_2),.clk(gclk));
	jdff dff_B_vPfTaCxx6_2(.din(w_dff_B_oNuoyF3A7_2),.dout(w_dff_B_vPfTaCxx6_2),.clk(gclk));
	jdff dff_B_eD3nbWwU9_2(.din(w_dff_B_vPfTaCxx6_2),.dout(w_dff_B_eD3nbWwU9_2),.clk(gclk));
	jdff dff_B_pBTxQ5713_2(.din(w_dff_B_eD3nbWwU9_2),.dout(w_dff_B_pBTxQ5713_2),.clk(gclk));
	jdff dff_B_9ZZIiemO0_2(.din(w_dff_B_pBTxQ5713_2),.dout(w_dff_B_9ZZIiemO0_2),.clk(gclk));
	jdff dff_B_9LB6HFc85_2(.din(w_dff_B_9ZZIiemO0_2),.dout(w_dff_B_9LB6HFc85_2),.clk(gclk));
	jdff dff_B_7FaVvQxr1_2(.din(w_dff_B_9LB6HFc85_2),.dout(w_dff_B_7FaVvQxr1_2),.clk(gclk));
	jdff dff_B_ycYhuZb70_2(.din(w_dff_B_7FaVvQxr1_2),.dout(w_dff_B_ycYhuZb70_2),.clk(gclk));
	jdff dff_B_VqRdzQjE5_2(.din(w_dff_B_ycYhuZb70_2),.dout(w_dff_B_VqRdzQjE5_2),.clk(gclk));
	jdff dff_B_hWqJidKw5_2(.din(w_dff_B_VqRdzQjE5_2),.dout(w_dff_B_hWqJidKw5_2),.clk(gclk));
	jdff dff_B_iCB3jWab0_2(.din(w_dff_B_hWqJidKw5_2),.dout(w_dff_B_iCB3jWab0_2),.clk(gclk));
	jdff dff_B_m2v3M6pB1_2(.din(w_dff_B_iCB3jWab0_2),.dout(w_dff_B_m2v3M6pB1_2),.clk(gclk));
	jdff dff_B_zD1LSr9q4_2(.din(w_dff_B_m2v3M6pB1_2),.dout(w_dff_B_zD1LSr9q4_2),.clk(gclk));
	jdff dff_B_LsO0OAbH8_2(.din(w_dff_B_zD1LSr9q4_2),.dout(w_dff_B_LsO0OAbH8_2),.clk(gclk));
	jdff dff_B_KUvefpuO2_2(.din(w_dff_B_LsO0OAbH8_2),.dout(w_dff_B_KUvefpuO2_2),.clk(gclk));
	jdff dff_B_wQDQTwAC4_2(.din(w_dff_B_KUvefpuO2_2),.dout(w_dff_B_wQDQTwAC4_2),.clk(gclk));
	jdff dff_B_RjcT4uXL9_2(.din(w_dff_B_wQDQTwAC4_2),.dout(w_dff_B_RjcT4uXL9_2),.clk(gclk));
	jdff dff_B_dhFdcFz57_2(.din(w_dff_B_RjcT4uXL9_2),.dout(w_dff_B_dhFdcFz57_2),.clk(gclk));
	jdff dff_B_GT7w1IgP9_2(.din(w_dff_B_dhFdcFz57_2),.dout(w_dff_B_GT7w1IgP9_2),.clk(gclk));
	jdff dff_B_3oDfo5a12_2(.din(n896),.dout(w_dff_B_3oDfo5a12_2),.clk(gclk));
	jdff dff_B_xSfesVRc9_1(.din(n828),.dout(w_dff_B_xSfesVRc9_1),.clk(gclk));
	jdff dff_B_ACgzCzzy6_2(.din(n729),.dout(w_dff_B_ACgzCzzy6_2),.clk(gclk));
	jdff dff_B_EpwGLWxt6_2(.din(w_dff_B_ACgzCzzy6_2),.dout(w_dff_B_EpwGLWxt6_2),.clk(gclk));
	jdff dff_B_0KCCAmmT6_2(.din(w_dff_B_EpwGLWxt6_2),.dout(w_dff_B_0KCCAmmT6_2),.clk(gclk));
	jdff dff_B_IaUUJVzR6_2(.din(w_dff_B_0KCCAmmT6_2),.dout(w_dff_B_IaUUJVzR6_2),.clk(gclk));
	jdff dff_B_p7n522pN3_2(.din(w_dff_B_IaUUJVzR6_2),.dout(w_dff_B_p7n522pN3_2),.clk(gclk));
	jdff dff_B_RemrzikY3_2(.din(w_dff_B_p7n522pN3_2),.dout(w_dff_B_RemrzikY3_2),.clk(gclk));
	jdff dff_B_noqfPgHG4_2(.din(w_dff_B_RemrzikY3_2),.dout(w_dff_B_noqfPgHG4_2),.clk(gclk));
	jdff dff_B_ozmbDJWM2_2(.din(w_dff_B_noqfPgHG4_2),.dout(w_dff_B_ozmbDJWM2_2),.clk(gclk));
	jdff dff_B_CxxdRRVv4_2(.din(w_dff_B_ozmbDJWM2_2),.dout(w_dff_B_CxxdRRVv4_2),.clk(gclk));
	jdff dff_B_wy24JjPb2_2(.din(w_dff_B_CxxdRRVv4_2),.dout(w_dff_B_wy24JjPb2_2),.clk(gclk));
	jdff dff_B_3rOkTWP09_2(.din(w_dff_B_wy24JjPb2_2),.dout(w_dff_B_3rOkTWP09_2),.clk(gclk));
	jdff dff_B_brsTDgjn3_2(.din(w_dff_B_3rOkTWP09_2),.dout(w_dff_B_brsTDgjn3_2),.clk(gclk));
	jdff dff_B_JDBlXzAt8_2(.din(w_dff_B_brsTDgjn3_2),.dout(w_dff_B_JDBlXzAt8_2),.clk(gclk));
	jdff dff_B_3QS68Yb67_2(.din(w_dff_B_JDBlXzAt8_2),.dout(w_dff_B_3QS68Yb67_2),.clk(gclk));
	jdff dff_B_10428VuR9_2(.din(w_dff_B_3QS68Yb67_2),.dout(w_dff_B_10428VuR9_2),.clk(gclk));
	jdff dff_B_RUxOQRP63_2(.din(w_dff_B_10428VuR9_2),.dout(w_dff_B_RUxOQRP63_2),.clk(gclk));
	jdff dff_B_hhPxUJtY2_2(.din(w_dff_B_RUxOQRP63_2),.dout(w_dff_B_hhPxUJtY2_2),.clk(gclk));
	jdff dff_B_9z4zqIHn4_2(.din(w_dff_B_hhPxUJtY2_2),.dout(w_dff_B_9z4zqIHn4_2),.clk(gclk));
	jdff dff_B_ZM71frwi0_2(.din(w_dff_B_9z4zqIHn4_2),.dout(w_dff_B_ZM71frwi0_2),.clk(gclk));
	jdff dff_B_GANWOPY97_2(.din(w_dff_B_ZM71frwi0_2),.dout(w_dff_B_GANWOPY97_2),.clk(gclk));
	jdff dff_B_EaXsR5ef7_2(.din(w_dff_B_GANWOPY97_2),.dout(w_dff_B_EaXsR5ef7_2),.clk(gclk));
	jdff dff_B_zBL5uHAf6_2(.din(w_dff_B_EaXsR5ef7_2),.dout(w_dff_B_zBL5uHAf6_2),.clk(gclk));
	jdff dff_B_lNTWVNJh3_2(.din(w_dff_B_zBL5uHAf6_2),.dout(w_dff_B_lNTWVNJh3_2),.clk(gclk));
	jdff dff_B_gvQiDGAg4_2(.din(w_dff_B_lNTWVNJh3_2),.dout(w_dff_B_gvQiDGAg4_2),.clk(gclk));
	jdff dff_B_jHwY5K0R5_2(.din(w_dff_B_gvQiDGAg4_2),.dout(w_dff_B_jHwY5K0R5_2),.clk(gclk));
	jdff dff_B_mXWLbgXM9_2(.din(w_dff_B_jHwY5K0R5_2),.dout(w_dff_B_mXWLbgXM9_2),.clk(gclk));
	jdff dff_B_FhOXP8Hs1_2(.din(w_dff_B_mXWLbgXM9_2),.dout(w_dff_B_FhOXP8Hs1_2),.clk(gclk));
	jdff dff_B_hscgPvLM9_2(.din(n793),.dout(w_dff_B_hscgPvLM9_2),.clk(gclk));
	jdff dff_B_mrmko7236_1(.din(n730),.dout(w_dff_B_mrmko7236_1),.clk(gclk));
	jdff dff_B_ocB1jjbI3_2(.din(n637),.dout(w_dff_B_ocB1jjbI3_2),.clk(gclk));
	jdff dff_B_AUp4NN9Q9_2(.din(w_dff_B_ocB1jjbI3_2),.dout(w_dff_B_AUp4NN9Q9_2),.clk(gclk));
	jdff dff_B_g3W2f0T00_2(.din(w_dff_B_AUp4NN9Q9_2),.dout(w_dff_B_g3W2f0T00_2),.clk(gclk));
	jdff dff_B_oFVbP1AG1_2(.din(w_dff_B_g3W2f0T00_2),.dout(w_dff_B_oFVbP1AG1_2),.clk(gclk));
	jdff dff_B_XRTOGGnO0_2(.din(w_dff_B_oFVbP1AG1_2),.dout(w_dff_B_XRTOGGnO0_2),.clk(gclk));
	jdff dff_B_83PCAdnc1_2(.din(w_dff_B_XRTOGGnO0_2),.dout(w_dff_B_83PCAdnc1_2),.clk(gclk));
	jdff dff_B_EAlun3y03_2(.din(w_dff_B_83PCAdnc1_2),.dout(w_dff_B_EAlun3y03_2),.clk(gclk));
	jdff dff_B_C4Sp9jHK7_2(.din(w_dff_B_EAlun3y03_2),.dout(w_dff_B_C4Sp9jHK7_2),.clk(gclk));
	jdff dff_B_wY7y3MAm8_2(.din(w_dff_B_C4Sp9jHK7_2),.dout(w_dff_B_wY7y3MAm8_2),.clk(gclk));
	jdff dff_B_GNL0tK2o3_2(.din(w_dff_B_wY7y3MAm8_2),.dout(w_dff_B_GNL0tK2o3_2),.clk(gclk));
	jdff dff_B_BlglAkr03_2(.din(w_dff_B_GNL0tK2o3_2),.dout(w_dff_B_BlglAkr03_2),.clk(gclk));
	jdff dff_B_EN5gKSgN7_2(.din(w_dff_B_BlglAkr03_2),.dout(w_dff_B_EN5gKSgN7_2),.clk(gclk));
	jdff dff_B_JhTLyd5I4_2(.din(w_dff_B_EN5gKSgN7_2),.dout(w_dff_B_JhTLyd5I4_2),.clk(gclk));
	jdff dff_B_uqytermL2_2(.din(w_dff_B_JhTLyd5I4_2),.dout(w_dff_B_uqytermL2_2),.clk(gclk));
	jdff dff_B_tm252inI4_2(.din(w_dff_B_uqytermL2_2),.dout(w_dff_B_tm252inI4_2),.clk(gclk));
	jdff dff_B_Z5Qox28V8_2(.din(w_dff_B_tm252inI4_2),.dout(w_dff_B_Z5Qox28V8_2),.clk(gclk));
	jdff dff_B_wsCNFRPd8_2(.din(w_dff_B_Z5Qox28V8_2),.dout(w_dff_B_wsCNFRPd8_2),.clk(gclk));
	jdff dff_B_n0qtncWA4_2(.din(w_dff_B_wsCNFRPd8_2),.dout(w_dff_B_n0qtncWA4_2),.clk(gclk));
	jdff dff_B_2LhLO1I82_2(.din(w_dff_B_n0qtncWA4_2),.dout(w_dff_B_2LhLO1I82_2),.clk(gclk));
	jdff dff_B_UJcDkIRb8_2(.din(w_dff_B_2LhLO1I82_2),.dout(w_dff_B_UJcDkIRb8_2),.clk(gclk));
	jdff dff_B_HaJrmOX11_2(.din(w_dff_B_UJcDkIRb8_2),.dout(w_dff_B_HaJrmOX11_2),.clk(gclk));
	jdff dff_B_fWLJ4b7X5_2(.din(w_dff_B_HaJrmOX11_2),.dout(w_dff_B_fWLJ4b7X5_2),.clk(gclk));
	jdff dff_B_w3HzIOnA0_2(.din(w_dff_B_fWLJ4b7X5_2),.dout(w_dff_B_w3HzIOnA0_2),.clk(gclk));
	jdff dff_B_7cQ7JSZV7_2(.din(w_dff_B_w3HzIOnA0_2),.dout(w_dff_B_7cQ7JSZV7_2),.clk(gclk));
	jdff dff_B_esxJIrZt0_2(.din(n694),.dout(w_dff_B_esxJIrZt0_2),.clk(gclk));
	jdff dff_B_01Q6TyWu5_1(.din(n638),.dout(w_dff_B_01Q6TyWu5_1),.clk(gclk));
	jdff dff_B_Q0Vv8isl2_2(.din(n552),.dout(w_dff_B_Q0Vv8isl2_2),.clk(gclk));
	jdff dff_B_qkTA4ZCi5_2(.din(w_dff_B_Q0Vv8isl2_2),.dout(w_dff_B_qkTA4ZCi5_2),.clk(gclk));
	jdff dff_B_YPgcGRzk3_2(.din(w_dff_B_qkTA4ZCi5_2),.dout(w_dff_B_YPgcGRzk3_2),.clk(gclk));
	jdff dff_B_Fue7o7j42_2(.din(w_dff_B_YPgcGRzk3_2),.dout(w_dff_B_Fue7o7j42_2),.clk(gclk));
	jdff dff_B_oMGLSwF08_2(.din(w_dff_B_Fue7o7j42_2),.dout(w_dff_B_oMGLSwF08_2),.clk(gclk));
	jdff dff_B_vw7MKNHx7_2(.din(w_dff_B_oMGLSwF08_2),.dout(w_dff_B_vw7MKNHx7_2),.clk(gclk));
	jdff dff_B_OfZUjcP04_2(.din(w_dff_B_vw7MKNHx7_2),.dout(w_dff_B_OfZUjcP04_2),.clk(gclk));
	jdff dff_B_QF3Mb0R18_2(.din(w_dff_B_OfZUjcP04_2),.dout(w_dff_B_QF3Mb0R18_2),.clk(gclk));
	jdff dff_B_rRPojT5y0_2(.din(w_dff_B_QF3Mb0R18_2),.dout(w_dff_B_rRPojT5y0_2),.clk(gclk));
	jdff dff_B_BqiFcAqp9_2(.din(w_dff_B_rRPojT5y0_2),.dout(w_dff_B_BqiFcAqp9_2),.clk(gclk));
	jdff dff_B_262lAmYn2_2(.din(w_dff_B_BqiFcAqp9_2),.dout(w_dff_B_262lAmYn2_2),.clk(gclk));
	jdff dff_B_fj7uJlEA1_2(.din(w_dff_B_262lAmYn2_2),.dout(w_dff_B_fj7uJlEA1_2),.clk(gclk));
	jdff dff_B_vch0NsBX7_2(.din(w_dff_B_fj7uJlEA1_2),.dout(w_dff_B_vch0NsBX7_2),.clk(gclk));
	jdff dff_B_Z1sKEGzN0_2(.din(w_dff_B_vch0NsBX7_2),.dout(w_dff_B_Z1sKEGzN0_2),.clk(gclk));
	jdff dff_B_2j8NJV3h3_2(.din(w_dff_B_Z1sKEGzN0_2),.dout(w_dff_B_2j8NJV3h3_2),.clk(gclk));
	jdff dff_B_TjX9jPaj6_2(.din(w_dff_B_2j8NJV3h3_2),.dout(w_dff_B_TjX9jPaj6_2),.clk(gclk));
	jdff dff_B_X7LZ0EPa1_2(.din(w_dff_B_TjX9jPaj6_2),.dout(w_dff_B_X7LZ0EPa1_2),.clk(gclk));
	jdff dff_B_rka0hyLL2_2(.din(w_dff_B_X7LZ0EPa1_2),.dout(w_dff_B_rka0hyLL2_2),.clk(gclk));
	jdff dff_B_1xmgAlz88_2(.din(w_dff_B_rka0hyLL2_2),.dout(w_dff_B_1xmgAlz88_2),.clk(gclk));
	jdff dff_B_26vWPJ9F8_2(.din(w_dff_B_1xmgAlz88_2),.dout(w_dff_B_26vWPJ9F8_2),.clk(gclk));
	jdff dff_B_5X81MMu62_2(.din(w_dff_B_26vWPJ9F8_2),.dout(w_dff_B_5X81MMu62_2),.clk(gclk));
	jdff dff_B_BwJipq5t9_2(.din(n602),.dout(w_dff_B_BwJipq5t9_2),.clk(gclk));
	jdff dff_B_bbmwRxcR6_1(.din(n553),.dout(w_dff_B_bbmwRxcR6_1),.clk(gclk));
	jdff dff_B_fq4m4c2V8_2(.din(n474),.dout(w_dff_B_fq4m4c2V8_2),.clk(gclk));
	jdff dff_B_ATKUlGrj4_2(.din(w_dff_B_fq4m4c2V8_2),.dout(w_dff_B_ATKUlGrj4_2),.clk(gclk));
	jdff dff_B_LuBiSRHd1_2(.din(w_dff_B_ATKUlGrj4_2),.dout(w_dff_B_LuBiSRHd1_2),.clk(gclk));
	jdff dff_B_jDPZHoBB1_2(.din(w_dff_B_LuBiSRHd1_2),.dout(w_dff_B_jDPZHoBB1_2),.clk(gclk));
	jdff dff_B_xiCAkGiy1_2(.din(w_dff_B_jDPZHoBB1_2),.dout(w_dff_B_xiCAkGiy1_2),.clk(gclk));
	jdff dff_B_01LedSxX2_2(.din(w_dff_B_xiCAkGiy1_2),.dout(w_dff_B_01LedSxX2_2),.clk(gclk));
	jdff dff_B_oBWK4tDx8_2(.din(w_dff_B_01LedSxX2_2),.dout(w_dff_B_oBWK4tDx8_2),.clk(gclk));
	jdff dff_B_1kqkdgZz1_2(.din(w_dff_B_oBWK4tDx8_2),.dout(w_dff_B_1kqkdgZz1_2),.clk(gclk));
	jdff dff_B_t5liWeGQ6_2(.din(w_dff_B_1kqkdgZz1_2),.dout(w_dff_B_t5liWeGQ6_2),.clk(gclk));
	jdff dff_B_93lIZMmJ3_2(.din(w_dff_B_t5liWeGQ6_2),.dout(w_dff_B_93lIZMmJ3_2),.clk(gclk));
	jdff dff_B_jeUgHtb47_2(.din(w_dff_B_93lIZMmJ3_2),.dout(w_dff_B_jeUgHtb47_2),.clk(gclk));
	jdff dff_B_AgUTF43S0_2(.din(w_dff_B_jeUgHtb47_2),.dout(w_dff_B_AgUTF43S0_2),.clk(gclk));
	jdff dff_B_Hc59ebKa1_2(.din(w_dff_B_AgUTF43S0_2),.dout(w_dff_B_Hc59ebKa1_2),.clk(gclk));
	jdff dff_B_tG8c4KYd0_2(.din(w_dff_B_Hc59ebKa1_2),.dout(w_dff_B_tG8c4KYd0_2),.clk(gclk));
	jdff dff_B_rIh6nSeB1_2(.din(w_dff_B_tG8c4KYd0_2),.dout(w_dff_B_rIh6nSeB1_2),.clk(gclk));
	jdff dff_B_yWq0szcb9_2(.din(w_dff_B_rIh6nSeB1_2),.dout(w_dff_B_yWq0szcb9_2),.clk(gclk));
	jdff dff_B_qhsSym3h7_2(.din(w_dff_B_yWq0szcb9_2),.dout(w_dff_B_qhsSym3h7_2),.clk(gclk));
	jdff dff_B_mnwGxLnu0_2(.din(w_dff_B_qhsSym3h7_2),.dout(w_dff_B_mnwGxLnu0_2),.clk(gclk));
	jdff dff_B_zuvg0Oqv6_2(.din(n517),.dout(w_dff_B_zuvg0Oqv6_2),.clk(gclk));
	jdff dff_B_wgPc0zdc6_1(.din(n475),.dout(w_dff_B_wgPc0zdc6_1),.clk(gclk));
	jdff dff_B_VcL1Bh4P4_2(.din(n403),.dout(w_dff_B_VcL1Bh4P4_2),.clk(gclk));
	jdff dff_B_ScNKj7PP7_2(.din(w_dff_B_VcL1Bh4P4_2),.dout(w_dff_B_ScNKj7PP7_2),.clk(gclk));
	jdff dff_B_bROEBImR9_2(.din(w_dff_B_ScNKj7PP7_2),.dout(w_dff_B_bROEBImR9_2),.clk(gclk));
	jdff dff_B_SIamB0yQ1_2(.din(w_dff_B_bROEBImR9_2),.dout(w_dff_B_SIamB0yQ1_2),.clk(gclk));
	jdff dff_B_Xo46XUiJ2_2(.din(w_dff_B_SIamB0yQ1_2),.dout(w_dff_B_Xo46XUiJ2_2),.clk(gclk));
	jdff dff_B_5YmWazk57_2(.din(w_dff_B_Xo46XUiJ2_2),.dout(w_dff_B_5YmWazk57_2),.clk(gclk));
	jdff dff_B_NtzlXOCR4_2(.din(w_dff_B_5YmWazk57_2),.dout(w_dff_B_NtzlXOCR4_2),.clk(gclk));
	jdff dff_B_wuTxWuA16_2(.din(w_dff_B_NtzlXOCR4_2),.dout(w_dff_B_wuTxWuA16_2),.clk(gclk));
	jdff dff_B_NQoEgRUb7_2(.din(w_dff_B_wuTxWuA16_2),.dout(w_dff_B_NQoEgRUb7_2),.clk(gclk));
	jdff dff_B_UfutkyBZ8_2(.din(w_dff_B_NQoEgRUb7_2),.dout(w_dff_B_UfutkyBZ8_2),.clk(gclk));
	jdff dff_B_3DJ74Piq1_2(.din(w_dff_B_UfutkyBZ8_2),.dout(w_dff_B_3DJ74Piq1_2),.clk(gclk));
	jdff dff_B_9pP8DoTt6_2(.din(w_dff_B_3DJ74Piq1_2),.dout(w_dff_B_9pP8DoTt6_2),.clk(gclk));
	jdff dff_B_Zdifc1bG5_2(.din(w_dff_B_9pP8DoTt6_2),.dout(w_dff_B_Zdifc1bG5_2),.clk(gclk));
	jdff dff_B_Houm7mY63_2(.din(w_dff_B_Zdifc1bG5_2),.dout(w_dff_B_Houm7mY63_2),.clk(gclk));
	jdff dff_B_546d4bqi9_2(.din(w_dff_B_Houm7mY63_2),.dout(w_dff_B_546d4bqi9_2),.clk(gclk));
	jdff dff_B_1pHowUne4_2(.din(n439),.dout(w_dff_B_1pHowUne4_2),.clk(gclk));
	jdff dff_B_V1BaO2AM1_1(.din(n404),.dout(w_dff_B_V1BaO2AM1_1),.clk(gclk));
	jdff dff_B_6n5rAh3B4_2(.din(n340),.dout(w_dff_B_6n5rAh3B4_2),.clk(gclk));
	jdff dff_B_kmyotDWx4_2(.din(w_dff_B_6n5rAh3B4_2),.dout(w_dff_B_kmyotDWx4_2),.clk(gclk));
	jdff dff_B_nNOGxE3k7_2(.din(w_dff_B_kmyotDWx4_2),.dout(w_dff_B_nNOGxE3k7_2),.clk(gclk));
	jdff dff_B_ktjlnF2F2_2(.din(w_dff_B_nNOGxE3k7_2),.dout(w_dff_B_ktjlnF2F2_2),.clk(gclk));
	jdff dff_B_IojyvBFz0_2(.din(w_dff_B_ktjlnF2F2_2),.dout(w_dff_B_IojyvBFz0_2),.clk(gclk));
	jdff dff_B_KcR8J3On6_2(.din(w_dff_B_IojyvBFz0_2),.dout(w_dff_B_KcR8J3On6_2),.clk(gclk));
	jdff dff_B_iZgEhadp4_2(.din(w_dff_B_KcR8J3On6_2),.dout(w_dff_B_iZgEhadp4_2),.clk(gclk));
	jdff dff_B_s7ibFKrE6_2(.din(w_dff_B_iZgEhadp4_2),.dout(w_dff_B_s7ibFKrE6_2),.clk(gclk));
	jdff dff_B_l1Ufrj157_2(.din(w_dff_B_s7ibFKrE6_2),.dout(w_dff_B_l1Ufrj157_2),.clk(gclk));
	jdff dff_B_4HYz8xk52_2(.din(w_dff_B_l1Ufrj157_2),.dout(w_dff_B_4HYz8xk52_2),.clk(gclk));
	jdff dff_B_MbPTzIlK1_2(.din(w_dff_B_4HYz8xk52_2),.dout(w_dff_B_MbPTzIlK1_2),.clk(gclk));
	jdff dff_B_980k4pLA3_2(.din(w_dff_B_MbPTzIlK1_2),.dout(w_dff_B_980k4pLA3_2),.clk(gclk));
	jdff dff_B_AhFWDYpV0_2(.din(n368),.dout(w_dff_B_AhFWDYpV0_2),.clk(gclk));
	jdff dff_B_P4zG5qW56_1(.din(n341),.dout(w_dff_B_P4zG5qW56_1),.clk(gclk));
	jdff dff_B_fEJ6gtzE9_2(.din(n284),.dout(w_dff_B_fEJ6gtzE9_2),.clk(gclk));
	jdff dff_B_6uPCicR67_2(.din(w_dff_B_fEJ6gtzE9_2),.dout(w_dff_B_6uPCicR67_2),.clk(gclk));
	jdff dff_B_Iu4Tv95D1_2(.din(w_dff_B_6uPCicR67_2),.dout(w_dff_B_Iu4Tv95D1_2),.clk(gclk));
	jdff dff_B_wxtrgoak2_2(.din(w_dff_B_Iu4Tv95D1_2),.dout(w_dff_B_wxtrgoak2_2),.clk(gclk));
	jdff dff_B_ytWLxDEr9_2(.din(w_dff_B_wxtrgoak2_2),.dout(w_dff_B_ytWLxDEr9_2),.clk(gclk));
	jdff dff_B_J9cF7xaz9_2(.din(w_dff_B_ytWLxDEr9_2),.dout(w_dff_B_J9cF7xaz9_2),.clk(gclk));
	jdff dff_B_EK5ZLz1L6_2(.din(w_dff_B_J9cF7xaz9_2),.dout(w_dff_B_EK5ZLz1L6_2),.clk(gclk));
	jdff dff_B_ZY0becf17_2(.din(w_dff_B_EK5ZLz1L6_2),.dout(w_dff_B_ZY0becf17_2),.clk(gclk));
	jdff dff_B_KI3bghAP8_2(.din(w_dff_B_ZY0becf17_2),.dout(w_dff_B_KI3bghAP8_2),.clk(gclk));
	jdff dff_B_SUc5WIUE5_2(.din(n305),.dout(w_dff_B_SUc5WIUE5_2),.clk(gclk));
	jdff dff_B_9qhXiizZ6_1(.din(n285),.dout(w_dff_B_9qhXiizZ6_1),.clk(gclk));
	jdff dff_B_4R52ri585_2(.din(n235),.dout(w_dff_B_4R52ri585_2),.clk(gclk));
	jdff dff_B_wwb2ZWi00_2(.din(w_dff_B_4R52ri585_2),.dout(w_dff_B_wwb2ZWi00_2),.clk(gclk));
	jdff dff_B_qVa0tE9x1_2(.din(w_dff_B_wwb2ZWi00_2),.dout(w_dff_B_qVa0tE9x1_2),.clk(gclk));
	jdff dff_B_GlxKCXPs3_2(.din(w_dff_B_qVa0tE9x1_2),.dout(w_dff_B_GlxKCXPs3_2),.clk(gclk));
	jdff dff_B_iPgtyqG65_2(.din(w_dff_B_GlxKCXPs3_2),.dout(w_dff_B_iPgtyqG65_2),.clk(gclk));
	jdff dff_B_r5l3dFb60_2(.din(w_dff_B_iPgtyqG65_2),.dout(w_dff_B_r5l3dFb60_2),.clk(gclk));
	jdff dff_B_F4vWvT7A0_2(.din(n249),.dout(w_dff_B_F4vWvT7A0_2),.clk(gclk));
	jdff dff_B_eTtxAsyR5_2(.din(n194),.dout(w_dff_B_eTtxAsyR5_2),.clk(gclk));
	jdff dff_B_qcV5ZJDx2_2(.din(w_dff_B_eTtxAsyR5_2),.dout(w_dff_B_qcV5ZJDx2_2),.clk(gclk));
	jdff dff_B_HzLkcPRY1_2(.din(w_dff_B_qcV5ZJDx2_2),.dout(w_dff_B_HzLkcPRY1_2),.clk(gclk));
	jdff dff_B_2jpNeUUR3_0(.din(n199),.dout(w_dff_B_2jpNeUUR3_0),.clk(gclk));
	jdff dff_A_71loFDDj1_0(.dout(w_n157_0[0]),.din(w_dff_A_71loFDDj1_0),.clk(gclk));
	jdff dff_A_e5uR1iD21_0(.dout(w_dff_A_71loFDDj1_0),.din(w_dff_A_e5uR1iD21_0),.clk(gclk));
	jdff dff_A_cW8jRnKE1_0(.dout(w_n156_0[0]),.din(w_dff_A_cW8jRnKE1_0),.clk(gclk));
	jdff dff_A_DABRaDyw5_0(.dout(w_dff_A_cW8jRnKE1_0),.din(w_dff_A_DABRaDyw5_0),.clk(gclk));
	jdff dff_B_63aFH6jf5_2(.din(n1389),.dout(w_dff_B_63aFH6jf5_2),.clk(gclk));
	jdff dff_B_NXjw3b0q3_1(.din(n1387),.dout(w_dff_B_NXjw3b0q3_1),.clk(gclk));
	jdff dff_B_WvNCcHnA0_2(.din(n1307),.dout(w_dff_B_WvNCcHnA0_2),.clk(gclk));
	jdff dff_B_f8kbonY97_2(.din(w_dff_B_WvNCcHnA0_2),.dout(w_dff_B_f8kbonY97_2),.clk(gclk));
	jdff dff_B_8NfIgwtA4_2(.din(w_dff_B_f8kbonY97_2),.dout(w_dff_B_8NfIgwtA4_2),.clk(gclk));
	jdff dff_B_2ZksKw4p4_2(.din(w_dff_B_8NfIgwtA4_2),.dout(w_dff_B_2ZksKw4p4_2),.clk(gclk));
	jdff dff_B_uJlInG0K5_2(.din(w_dff_B_2ZksKw4p4_2),.dout(w_dff_B_uJlInG0K5_2),.clk(gclk));
	jdff dff_B_fBEpW50U9_2(.din(w_dff_B_uJlInG0K5_2),.dout(w_dff_B_fBEpW50U9_2),.clk(gclk));
	jdff dff_B_XYP0Xn6a7_2(.din(w_dff_B_fBEpW50U9_2),.dout(w_dff_B_XYP0Xn6a7_2),.clk(gclk));
	jdff dff_B_ZmOH45Qj1_2(.din(w_dff_B_XYP0Xn6a7_2),.dout(w_dff_B_ZmOH45Qj1_2),.clk(gclk));
	jdff dff_B_1xEWzVFg6_2(.din(w_dff_B_ZmOH45Qj1_2),.dout(w_dff_B_1xEWzVFg6_2),.clk(gclk));
	jdff dff_B_IopllFTi0_2(.din(w_dff_B_1xEWzVFg6_2),.dout(w_dff_B_IopllFTi0_2),.clk(gclk));
	jdff dff_B_DNcvq4FG5_2(.din(w_dff_B_IopllFTi0_2),.dout(w_dff_B_DNcvq4FG5_2),.clk(gclk));
	jdff dff_B_vBptDxCp8_2(.din(w_dff_B_DNcvq4FG5_2),.dout(w_dff_B_vBptDxCp8_2),.clk(gclk));
	jdff dff_B_JAgECIsB1_2(.din(w_dff_B_vBptDxCp8_2),.dout(w_dff_B_JAgECIsB1_2),.clk(gclk));
	jdff dff_B_iXRYG9OM9_2(.din(w_dff_B_JAgECIsB1_2),.dout(w_dff_B_iXRYG9OM9_2),.clk(gclk));
	jdff dff_B_zigsYATG0_2(.din(w_dff_B_iXRYG9OM9_2),.dout(w_dff_B_zigsYATG0_2),.clk(gclk));
	jdff dff_B_BvKVLXxp5_2(.din(w_dff_B_zigsYATG0_2),.dout(w_dff_B_BvKVLXxp5_2),.clk(gclk));
	jdff dff_B_NlOVZJQk9_2(.din(w_dff_B_BvKVLXxp5_2),.dout(w_dff_B_NlOVZJQk9_2),.clk(gclk));
	jdff dff_B_jZSMzs900_2(.din(w_dff_B_NlOVZJQk9_2),.dout(w_dff_B_jZSMzs900_2),.clk(gclk));
	jdff dff_B_xae5irdm1_2(.din(w_dff_B_jZSMzs900_2),.dout(w_dff_B_xae5irdm1_2),.clk(gclk));
	jdff dff_B_pBanHuaK9_2(.din(w_dff_B_xae5irdm1_2),.dout(w_dff_B_pBanHuaK9_2),.clk(gclk));
	jdff dff_B_tytTMAzz5_2(.din(w_dff_B_pBanHuaK9_2),.dout(w_dff_B_tytTMAzz5_2),.clk(gclk));
	jdff dff_B_2G6giiJ93_2(.din(w_dff_B_tytTMAzz5_2),.dout(w_dff_B_2G6giiJ93_2),.clk(gclk));
	jdff dff_B_pSwy0n4h3_2(.din(w_dff_B_2G6giiJ93_2),.dout(w_dff_B_pSwy0n4h3_2),.clk(gclk));
	jdff dff_B_FQH5nr1b5_2(.din(w_dff_B_pSwy0n4h3_2),.dout(w_dff_B_FQH5nr1b5_2),.clk(gclk));
	jdff dff_B_AnmhUVRA9_2(.din(w_dff_B_FQH5nr1b5_2),.dout(w_dff_B_AnmhUVRA9_2),.clk(gclk));
	jdff dff_B_F2cpkg8H8_2(.din(w_dff_B_AnmhUVRA9_2),.dout(w_dff_B_F2cpkg8H8_2),.clk(gclk));
	jdff dff_B_pitjU4zR9_2(.din(w_dff_B_F2cpkg8H8_2),.dout(w_dff_B_pitjU4zR9_2),.clk(gclk));
	jdff dff_B_uBkY3qeW1_2(.din(w_dff_B_pitjU4zR9_2),.dout(w_dff_B_uBkY3qeW1_2),.clk(gclk));
	jdff dff_B_R2GrY3aD8_2(.din(w_dff_B_uBkY3qeW1_2),.dout(w_dff_B_R2GrY3aD8_2),.clk(gclk));
	jdff dff_B_Jl7i3bOb1_2(.din(w_dff_B_R2GrY3aD8_2),.dout(w_dff_B_Jl7i3bOb1_2),.clk(gclk));
	jdff dff_B_zaYUQXuh4_2(.din(w_dff_B_Jl7i3bOb1_2),.dout(w_dff_B_zaYUQXuh4_2),.clk(gclk));
	jdff dff_B_ubN5tJLJ2_2(.din(w_dff_B_zaYUQXuh4_2),.dout(w_dff_B_ubN5tJLJ2_2),.clk(gclk));
	jdff dff_B_M092GrGo9_2(.din(w_dff_B_ubN5tJLJ2_2),.dout(w_dff_B_M092GrGo9_2),.clk(gclk));
	jdff dff_B_WNO4BPVO5_2(.din(w_dff_B_M092GrGo9_2),.dout(w_dff_B_WNO4BPVO5_2),.clk(gclk));
	jdff dff_B_OmOUMwOM4_2(.din(w_dff_B_WNO4BPVO5_2),.dout(w_dff_B_OmOUMwOM4_2),.clk(gclk));
	jdff dff_B_kaNslhL44_2(.din(w_dff_B_OmOUMwOM4_2),.dout(w_dff_B_kaNslhL44_2),.clk(gclk));
	jdff dff_B_cqXn2RsE7_2(.din(w_dff_B_kaNslhL44_2),.dout(w_dff_B_cqXn2RsE7_2),.clk(gclk));
	jdff dff_B_1bs89Hry2_2(.din(w_dff_B_cqXn2RsE7_2),.dout(w_dff_B_1bs89Hry2_2),.clk(gclk));
	jdff dff_B_kbo3ePki4_2(.din(w_dff_B_1bs89Hry2_2),.dout(w_dff_B_kbo3ePki4_2),.clk(gclk));
	jdff dff_B_g9IC65jP2_2(.din(w_dff_B_kbo3ePki4_2),.dout(w_dff_B_g9IC65jP2_2),.clk(gclk));
	jdff dff_B_vaMCqxmS3_2(.din(w_dff_B_g9IC65jP2_2),.dout(w_dff_B_vaMCqxmS3_2),.clk(gclk));
	jdff dff_B_mYVREC2A6_2(.din(w_dff_B_vaMCqxmS3_2),.dout(w_dff_B_mYVREC2A6_2),.clk(gclk));
	jdff dff_B_0x579tDP8_2(.din(w_dff_B_mYVREC2A6_2),.dout(w_dff_B_0x579tDP8_2),.clk(gclk));
	jdff dff_B_bG0rai9o5_2(.din(w_dff_B_0x579tDP8_2),.dout(w_dff_B_bG0rai9o5_2),.clk(gclk));
	jdff dff_B_IZi3Ndf67_1(.din(n1308),.dout(w_dff_B_IZi3Ndf67_1),.clk(gclk));
	jdff dff_B_s0RBPDHg1_2(.din(n1222),.dout(w_dff_B_s0RBPDHg1_2),.clk(gclk));
	jdff dff_B_HanLoImk7_2(.din(w_dff_B_s0RBPDHg1_2),.dout(w_dff_B_HanLoImk7_2),.clk(gclk));
	jdff dff_B_i0pgx0Z16_2(.din(w_dff_B_HanLoImk7_2),.dout(w_dff_B_i0pgx0Z16_2),.clk(gclk));
	jdff dff_B_iBy4ifVi2_2(.din(w_dff_B_i0pgx0Z16_2),.dout(w_dff_B_iBy4ifVi2_2),.clk(gclk));
	jdff dff_B_vvZ4gUhA0_2(.din(w_dff_B_iBy4ifVi2_2),.dout(w_dff_B_vvZ4gUhA0_2),.clk(gclk));
	jdff dff_B_BJx4rVKg0_2(.din(w_dff_B_vvZ4gUhA0_2),.dout(w_dff_B_BJx4rVKg0_2),.clk(gclk));
	jdff dff_B_qlJRZGE67_2(.din(w_dff_B_BJx4rVKg0_2),.dout(w_dff_B_qlJRZGE67_2),.clk(gclk));
	jdff dff_B_G7W6kMJl5_2(.din(w_dff_B_qlJRZGE67_2),.dout(w_dff_B_G7W6kMJl5_2),.clk(gclk));
	jdff dff_B_5MNwe50O3_2(.din(w_dff_B_G7W6kMJl5_2),.dout(w_dff_B_5MNwe50O3_2),.clk(gclk));
	jdff dff_B_FTIZ3PTc0_2(.din(w_dff_B_5MNwe50O3_2),.dout(w_dff_B_FTIZ3PTc0_2),.clk(gclk));
	jdff dff_B_iJTd623c1_2(.din(w_dff_B_FTIZ3PTc0_2),.dout(w_dff_B_iJTd623c1_2),.clk(gclk));
	jdff dff_B_wkqF6ASz4_2(.din(w_dff_B_iJTd623c1_2),.dout(w_dff_B_wkqF6ASz4_2),.clk(gclk));
	jdff dff_B_Lu7EvZan6_2(.din(w_dff_B_wkqF6ASz4_2),.dout(w_dff_B_Lu7EvZan6_2),.clk(gclk));
	jdff dff_B_mKMRxdbQ6_2(.din(w_dff_B_Lu7EvZan6_2),.dout(w_dff_B_mKMRxdbQ6_2),.clk(gclk));
	jdff dff_B_d4f1OTzO1_2(.din(w_dff_B_mKMRxdbQ6_2),.dout(w_dff_B_d4f1OTzO1_2),.clk(gclk));
	jdff dff_B_wkEdgNyA8_2(.din(w_dff_B_d4f1OTzO1_2),.dout(w_dff_B_wkEdgNyA8_2),.clk(gclk));
	jdff dff_B_qTliLYmf8_2(.din(w_dff_B_wkEdgNyA8_2),.dout(w_dff_B_qTliLYmf8_2),.clk(gclk));
	jdff dff_B_bmAX0loh9_2(.din(w_dff_B_qTliLYmf8_2),.dout(w_dff_B_bmAX0loh9_2),.clk(gclk));
	jdff dff_B_I5evKUXl8_2(.din(w_dff_B_bmAX0loh9_2),.dout(w_dff_B_I5evKUXl8_2),.clk(gclk));
	jdff dff_B_cAl4t5yr7_2(.din(w_dff_B_I5evKUXl8_2),.dout(w_dff_B_cAl4t5yr7_2),.clk(gclk));
	jdff dff_B_MAC51qts6_2(.din(w_dff_B_cAl4t5yr7_2),.dout(w_dff_B_MAC51qts6_2),.clk(gclk));
	jdff dff_B_L9WLI6E84_2(.din(w_dff_B_MAC51qts6_2),.dout(w_dff_B_L9WLI6E84_2),.clk(gclk));
	jdff dff_B_e1YpAWm89_2(.din(w_dff_B_L9WLI6E84_2),.dout(w_dff_B_e1YpAWm89_2),.clk(gclk));
	jdff dff_B_fmkLYH6Y3_2(.din(w_dff_B_e1YpAWm89_2),.dout(w_dff_B_fmkLYH6Y3_2),.clk(gclk));
	jdff dff_B_f7nwM4HE0_2(.din(w_dff_B_fmkLYH6Y3_2),.dout(w_dff_B_f7nwM4HE0_2),.clk(gclk));
	jdff dff_B_3DklKBKb4_2(.din(w_dff_B_f7nwM4HE0_2),.dout(w_dff_B_3DklKBKb4_2),.clk(gclk));
	jdff dff_B_m7nhDawH8_2(.din(w_dff_B_3DklKBKb4_2),.dout(w_dff_B_m7nhDawH8_2),.clk(gclk));
	jdff dff_B_twoavS7N1_2(.din(w_dff_B_m7nhDawH8_2),.dout(w_dff_B_twoavS7N1_2),.clk(gclk));
	jdff dff_B_1EZMyTPq3_2(.din(w_dff_B_twoavS7N1_2),.dout(w_dff_B_1EZMyTPq3_2),.clk(gclk));
	jdff dff_B_K3pDCnNB2_2(.din(w_dff_B_1EZMyTPq3_2),.dout(w_dff_B_K3pDCnNB2_2),.clk(gclk));
	jdff dff_B_YsxVunNc3_2(.din(w_dff_B_K3pDCnNB2_2),.dout(w_dff_B_YsxVunNc3_2),.clk(gclk));
	jdff dff_B_TrjhvAcA3_2(.din(w_dff_B_YsxVunNc3_2),.dout(w_dff_B_TrjhvAcA3_2),.clk(gclk));
	jdff dff_B_5o002yxn8_2(.din(w_dff_B_TrjhvAcA3_2),.dout(w_dff_B_5o002yxn8_2),.clk(gclk));
	jdff dff_B_0elspNfO9_2(.din(w_dff_B_5o002yxn8_2),.dout(w_dff_B_0elspNfO9_2),.clk(gclk));
	jdff dff_B_8DFGrMkU5_2(.din(w_dff_B_0elspNfO9_2),.dout(w_dff_B_8DFGrMkU5_2),.clk(gclk));
	jdff dff_B_rUGFPC6f3_2(.din(w_dff_B_8DFGrMkU5_2),.dout(w_dff_B_rUGFPC6f3_2),.clk(gclk));
	jdff dff_B_ex0Bfp8v6_2(.din(w_dff_B_rUGFPC6f3_2),.dout(w_dff_B_ex0Bfp8v6_2),.clk(gclk));
	jdff dff_B_0Mw3Lr6J3_2(.din(w_dff_B_ex0Bfp8v6_2),.dout(w_dff_B_0Mw3Lr6J3_2),.clk(gclk));
	jdff dff_B_xDLoDmzC7_2(.din(w_dff_B_0Mw3Lr6J3_2),.dout(w_dff_B_xDLoDmzC7_2),.clk(gclk));
	jdff dff_B_5a7iCyKw7_1(.din(n1223),.dout(w_dff_B_5a7iCyKw7_1),.clk(gclk));
	jdff dff_B_xWuhoX1X7_2(.din(n1131),.dout(w_dff_B_xWuhoX1X7_2),.clk(gclk));
	jdff dff_B_h95ajs822_2(.din(w_dff_B_xWuhoX1X7_2),.dout(w_dff_B_h95ajs822_2),.clk(gclk));
	jdff dff_B_uMhWJFrQ3_2(.din(w_dff_B_h95ajs822_2),.dout(w_dff_B_uMhWJFrQ3_2),.clk(gclk));
	jdff dff_B_W4LQSCaJ2_2(.din(w_dff_B_uMhWJFrQ3_2),.dout(w_dff_B_W4LQSCaJ2_2),.clk(gclk));
	jdff dff_B_LM7e9pCe9_2(.din(w_dff_B_W4LQSCaJ2_2),.dout(w_dff_B_LM7e9pCe9_2),.clk(gclk));
	jdff dff_B_pQb67gyp1_2(.din(w_dff_B_LM7e9pCe9_2),.dout(w_dff_B_pQb67gyp1_2),.clk(gclk));
	jdff dff_B_nfUE4tXR6_2(.din(w_dff_B_pQb67gyp1_2),.dout(w_dff_B_nfUE4tXR6_2),.clk(gclk));
	jdff dff_B_pUNhOJ6l1_2(.din(w_dff_B_nfUE4tXR6_2),.dout(w_dff_B_pUNhOJ6l1_2),.clk(gclk));
	jdff dff_B_zbVRkb4F0_2(.din(w_dff_B_pUNhOJ6l1_2),.dout(w_dff_B_zbVRkb4F0_2),.clk(gclk));
	jdff dff_B_olFUxNMp8_2(.din(w_dff_B_zbVRkb4F0_2),.dout(w_dff_B_olFUxNMp8_2),.clk(gclk));
	jdff dff_B_BojOT41K0_2(.din(w_dff_B_olFUxNMp8_2),.dout(w_dff_B_BojOT41K0_2),.clk(gclk));
	jdff dff_B_m0Q8sLYB5_2(.din(w_dff_B_BojOT41K0_2),.dout(w_dff_B_m0Q8sLYB5_2),.clk(gclk));
	jdff dff_B_r7Mjqsdp4_2(.din(w_dff_B_m0Q8sLYB5_2),.dout(w_dff_B_r7Mjqsdp4_2),.clk(gclk));
	jdff dff_B_O6O25vXp3_2(.din(w_dff_B_r7Mjqsdp4_2),.dout(w_dff_B_O6O25vXp3_2),.clk(gclk));
	jdff dff_B_AoYe3P4t7_2(.din(w_dff_B_O6O25vXp3_2),.dout(w_dff_B_AoYe3P4t7_2),.clk(gclk));
	jdff dff_B_EHDWu3SD6_2(.din(w_dff_B_AoYe3P4t7_2),.dout(w_dff_B_EHDWu3SD6_2),.clk(gclk));
	jdff dff_B_ZVfuvzi73_2(.din(w_dff_B_EHDWu3SD6_2),.dout(w_dff_B_ZVfuvzi73_2),.clk(gclk));
	jdff dff_B_9C29qdIr1_2(.din(w_dff_B_ZVfuvzi73_2),.dout(w_dff_B_9C29qdIr1_2),.clk(gclk));
	jdff dff_B_X5MY2tUt9_2(.din(w_dff_B_9C29qdIr1_2),.dout(w_dff_B_X5MY2tUt9_2),.clk(gclk));
	jdff dff_B_Ogz8plhk6_2(.din(w_dff_B_X5MY2tUt9_2),.dout(w_dff_B_Ogz8plhk6_2),.clk(gclk));
	jdff dff_B_UPlVshC21_2(.din(w_dff_B_Ogz8plhk6_2),.dout(w_dff_B_UPlVshC21_2),.clk(gclk));
	jdff dff_B_mvvDJxYs1_2(.din(w_dff_B_UPlVshC21_2),.dout(w_dff_B_mvvDJxYs1_2),.clk(gclk));
	jdff dff_B_oMYsIgpL8_2(.din(w_dff_B_mvvDJxYs1_2),.dout(w_dff_B_oMYsIgpL8_2),.clk(gclk));
	jdff dff_B_PreNpc8t8_2(.din(w_dff_B_oMYsIgpL8_2),.dout(w_dff_B_PreNpc8t8_2),.clk(gclk));
	jdff dff_B_oG5d7WuC0_2(.din(w_dff_B_PreNpc8t8_2),.dout(w_dff_B_oG5d7WuC0_2),.clk(gclk));
	jdff dff_B_vg6e87IX2_2(.din(w_dff_B_oG5d7WuC0_2),.dout(w_dff_B_vg6e87IX2_2),.clk(gclk));
	jdff dff_B_RKLdNgBi0_2(.din(w_dff_B_vg6e87IX2_2),.dout(w_dff_B_RKLdNgBi0_2),.clk(gclk));
	jdff dff_B_lofPN2A51_2(.din(w_dff_B_RKLdNgBi0_2),.dout(w_dff_B_lofPN2A51_2),.clk(gclk));
	jdff dff_B_iypVaiuf5_2(.din(w_dff_B_lofPN2A51_2),.dout(w_dff_B_iypVaiuf5_2),.clk(gclk));
	jdff dff_B_sDLTB4A11_2(.din(w_dff_B_iypVaiuf5_2),.dout(w_dff_B_sDLTB4A11_2),.clk(gclk));
	jdff dff_B_OiK8AIAa3_2(.din(w_dff_B_sDLTB4A11_2),.dout(w_dff_B_OiK8AIAa3_2),.clk(gclk));
	jdff dff_B_LzUwFY2H5_2(.din(w_dff_B_OiK8AIAa3_2),.dout(w_dff_B_LzUwFY2H5_2),.clk(gclk));
	jdff dff_B_k0tfvsBB0_2(.din(w_dff_B_LzUwFY2H5_2),.dout(w_dff_B_k0tfvsBB0_2),.clk(gclk));
	jdff dff_B_PzPgs8xv5_2(.din(w_dff_B_k0tfvsBB0_2),.dout(w_dff_B_PzPgs8xv5_2),.clk(gclk));
	jdff dff_B_NBnXsbqy3_2(.din(w_dff_B_PzPgs8xv5_2),.dout(w_dff_B_NBnXsbqy3_2),.clk(gclk));
	jdff dff_B_3asv6Oq43_2(.din(w_dff_B_NBnXsbqy3_2),.dout(w_dff_B_3asv6Oq43_2),.clk(gclk));
	jdff dff_B_68zJrRQn6_1(.din(n1132),.dout(w_dff_B_68zJrRQn6_1),.clk(gclk));
	jdff dff_B_5OwEFkNk1_2(.din(n1033),.dout(w_dff_B_5OwEFkNk1_2),.clk(gclk));
	jdff dff_B_6AfpDX0Q5_2(.din(w_dff_B_5OwEFkNk1_2),.dout(w_dff_B_6AfpDX0Q5_2),.clk(gclk));
	jdff dff_B_26Pxisgh1_2(.din(w_dff_B_6AfpDX0Q5_2),.dout(w_dff_B_26Pxisgh1_2),.clk(gclk));
	jdff dff_B_JWMmyMSp1_2(.din(w_dff_B_26Pxisgh1_2),.dout(w_dff_B_JWMmyMSp1_2),.clk(gclk));
	jdff dff_B_KLbaXe9X5_2(.din(w_dff_B_JWMmyMSp1_2),.dout(w_dff_B_KLbaXe9X5_2),.clk(gclk));
	jdff dff_B_zdqxO4HL0_2(.din(w_dff_B_KLbaXe9X5_2),.dout(w_dff_B_zdqxO4HL0_2),.clk(gclk));
	jdff dff_B_93Oe04y36_2(.din(w_dff_B_zdqxO4HL0_2),.dout(w_dff_B_93Oe04y36_2),.clk(gclk));
	jdff dff_B_jos6fRZi3_2(.din(w_dff_B_93Oe04y36_2),.dout(w_dff_B_jos6fRZi3_2),.clk(gclk));
	jdff dff_B_6te7F88y9_2(.din(w_dff_B_jos6fRZi3_2),.dout(w_dff_B_6te7F88y9_2),.clk(gclk));
	jdff dff_B_lsfY90UX1_2(.din(w_dff_B_6te7F88y9_2),.dout(w_dff_B_lsfY90UX1_2),.clk(gclk));
	jdff dff_B_gLAVDZFi7_2(.din(w_dff_B_lsfY90UX1_2),.dout(w_dff_B_gLAVDZFi7_2),.clk(gclk));
	jdff dff_B_h9r6XC8H2_2(.din(w_dff_B_gLAVDZFi7_2),.dout(w_dff_B_h9r6XC8H2_2),.clk(gclk));
	jdff dff_B_37yEnHBD8_2(.din(w_dff_B_h9r6XC8H2_2),.dout(w_dff_B_37yEnHBD8_2),.clk(gclk));
	jdff dff_B_XQBSTqUz2_2(.din(w_dff_B_37yEnHBD8_2),.dout(w_dff_B_XQBSTqUz2_2),.clk(gclk));
	jdff dff_B_xFo5YbXJ5_2(.din(w_dff_B_XQBSTqUz2_2),.dout(w_dff_B_xFo5YbXJ5_2),.clk(gclk));
	jdff dff_B_eR3Rib7Z5_2(.din(w_dff_B_xFo5YbXJ5_2),.dout(w_dff_B_eR3Rib7Z5_2),.clk(gclk));
	jdff dff_B_VJN6Tcim2_2(.din(w_dff_B_eR3Rib7Z5_2),.dout(w_dff_B_VJN6Tcim2_2),.clk(gclk));
	jdff dff_B_vJZdUpQX3_2(.din(w_dff_B_VJN6Tcim2_2),.dout(w_dff_B_vJZdUpQX3_2),.clk(gclk));
	jdff dff_B_V586TrTw1_2(.din(w_dff_B_vJZdUpQX3_2),.dout(w_dff_B_V586TrTw1_2),.clk(gclk));
	jdff dff_B_P5tkvkhM7_2(.din(w_dff_B_V586TrTw1_2),.dout(w_dff_B_P5tkvkhM7_2),.clk(gclk));
	jdff dff_B_BRKgUOf11_2(.din(w_dff_B_P5tkvkhM7_2),.dout(w_dff_B_BRKgUOf11_2),.clk(gclk));
	jdff dff_B_yPMyfZje9_2(.din(w_dff_B_BRKgUOf11_2),.dout(w_dff_B_yPMyfZje9_2),.clk(gclk));
	jdff dff_B_ZIjmV4ZI3_2(.din(w_dff_B_yPMyfZje9_2),.dout(w_dff_B_ZIjmV4ZI3_2),.clk(gclk));
	jdff dff_B_BoQb4wAr7_2(.din(w_dff_B_ZIjmV4ZI3_2),.dout(w_dff_B_BoQb4wAr7_2),.clk(gclk));
	jdff dff_B_j6wsByxZ4_2(.din(w_dff_B_BoQb4wAr7_2),.dout(w_dff_B_j6wsByxZ4_2),.clk(gclk));
	jdff dff_B_VjWvqrvv0_2(.din(w_dff_B_j6wsByxZ4_2),.dout(w_dff_B_VjWvqrvv0_2),.clk(gclk));
	jdff dff_B_GuVVIFjE3_2(.din(w_dff_B_VjWvqrvv0_2),.dout(w_dff_B_GuVVIFjE3_2),.clk(gclk));
	jdff dff_B_HFFPNWWF1_2(.din(w_dff_B_GuVVIFjE3_2),.dout(w_dff_B_HFFPNWWF1_2),.clk(gclk));
	jdff dff_B_N2o7P2Iu6_2(.din(w_dff_B_HFFPNWWF1_2),.dout(w_dff_B_N2o7P2Iu6_2),.clk(gclk));
	jdff dff_B_JkOHAxqH1_2(.din(w_dff_B_N2o7P2Iu6_2),.dout(w_dff_B_JkOHAxqH1_2),.clk(gclk));
	jdff dff_B_Vx0eqJSd2_2(.din(w_dff_B_JkOHAxqH1_2),.dout(w_dff_B_Vx0eqJSd2_2),.clk(gclk));
	jdff dff_B_7SaKbanj4_2(.din(w_dff_B_Vx0eqJSd2_2),.dout(w_dff_B_7SaKbanj4_2),.clk(gclk));
	jdff dff_B_JxLDU3Sf6_2(.din(w_dff_B_7SaKbanj4_2),.dout(w_dff_B_JxLDU3Sf6_2),.clk(gclk));
	jdff dff_B_Nkz8yQSe9_1(.din(n1034),.dout(w_dff_B_Nkz8yQSe9_1),.clk(gclk));
	jdff dff_B_oPWwfmOW2_2(.din(n934),.dout(w_dff_B_oPWwfmOW2_2),.clk(gclk));
	jdff dff_B_PDRDQaFX9_2(.din(w_dff_B_oPWwfmOW2_2),.dout(w_dff_B_PDRDQaFX9_2),.clk(gclk));
	jdff dff_B_jHHJ8PDx1_2(.din(w_dff_B_PDRDQaFX9_2),.dout(w_dff_B_jHHJ8PDx1_2),.clk(gclk));
	jdff dff_B_7Xo00ENa2_2(.din(w_dff_B_jHHJ8PDx1_2),.dout(w_dff_B_7Xo00ENa2_2),.clk(gclk));
	jdff dff_B_i6tYNkW57_2(.din(w_dff_B_7Xo00ENa2_2),.dout(w_dff_B_i6tYNkW57_2),.clk(gclk));
	jdff dff_B_4qVXhN027_2(.din(w_dff_B_i6tYNkW57_2),.dout(w_dff_B_4qVXhN027_2),.clk(gclk));
	jdff dff_B_HLzOduDW4_2(.din(w_dff_B_4qVXhN027_2),.dout(w_dff_B_HLzOduDW4_2),.clk(gclk));
	jdff dff_B_91Bkjm9r1_2(.din(w_dff_B_HLzOduDW4_2),.dout(w_dff_B_91Bkjm9r1_2),.clk(gclk));
	jdff dff_B_pUeuR6Vw4_2(.din(w_dff_B_91Bkjm9r1_2),.dout(w_dff_B_pUeuR6Vw4_2),.clk(gclk));
	jdff dff_B_44gx8QK28_2(.din(w_dff_B_pUeuR6Vw4_2),.dout(w_dff_B_44gx8QK28_2),.clk(gclk));
	jdff dff_B_IBDQiS018_2(.din(w_dff_B_44gx8QK28_2),.dout(w_dff_B_IBDQiS018_2),.clk(gclk));
	jdff dff_B_ZBibaqdY2_2(.din(w_dff_B_IBDQiS018_2),.dout(w_dff_B_ZBibaqdY2_2),.clk(gclk));
	jdff dff_B_wSjEQpSB5_2(.din(w_dff_B_ZBibaqdY2_2),.dout(w_dff_B_wSjEQpSB5_2),.clk(gclk));
	jdff dff_B_Uzxdb5j56_2(.din(w_dff_B_wSjEQpSB5_2),.dout(w_dff_B_Uzxdb5j56_2),.clk(gclk));
	jdff dff_B_EIawDFfw6_2(.din(w_dff_B_Uzxdb5j56_2),.dout(w_dff_B_EIawDFfw6_2),.clk(gclk));
	jdff dff_B_nrWNiFgD4_2(.din(w_dff_B_EIawDFfw6_2),.dout(w_dff_B_nrWNiFgD4_2),.clk(gclk));
	jdff dff_B_Z87vWLnY3_2(.din(w_dff_B_nrWNiFgD4_2),.dout(w_dff_B_Z87vWLnY3_2),.clk(gclk));
	jdff dff_B_uUyHDpO56_2(.din(w_dff_B_Z87vWLnY3_2),.dout(w_dff_B_uUyHDpO56_2),.clk(gclk));
	jdff dff_B_d5fzpVRe0_2(.din(w_dff_B_uUyHDpO56_2),.dout(w_dff_B_d5fzpVRe0_2),.clk(gclk));
	jdff dff_B_rkYMmdb34_2(.din(w_dff_B_d5fzpVRe0_2),.dout(w_dff_B_rkYMmdb34_2),.clk(gclk));
	jdff dff_B_Gnv8Uims4_2(.din(w_dff_B_rkYMmdb34_2),.dout(w_dff_B_Gnv8Uims4_2),.clk(gclk));
	jdff dff_B_sds1cPBn4_2(.din(w_dff_B_Gnv8Uims4_2),.dout(w_dff_B_sds1cPBn4_2),.clk(gclk));
	jdff dff_B_0CgY84cr6_2(.din(w_dff_B_sds1cPBn4_2),.dout(w_dff_B_0CgY84cr6_2),.clk(gclk));
	jdff dff_B_KFEh2fMa6_2(.din(w_dff_B_0CgY84cr6_2),.dout(w_dff_B_KFEh2fMa6_2),.clk(gclk));
	jdff dff_B_KXruVjqQ3_2(.din(w_dff_B_KFEh2fMa6_2),.dout(w_dff_B_KXruVjqQ3_2),.clk(gclk));
	jdff dff_B_rXhW6QRZ7_2(.din(w_dff_B_KXruVjqQ3_2),.dout(w_dff_B_rXhW6QRZ7_2),.clk(gclk));
	jdff dff_B_7d3MHg1i2_2(.din(w_dff_B_rXhW6QRZ7_2),.dout(w_dff_B_7d3MHg1i2_2),.clk(gclk));
	jdff dff_B_5rJqiBB32_2(.din(w_dff_B_7d3MHg1i2_2),.dout(w_dff_B_5rJqiBB32_2),.clk(gclk));
	jdff dff_B_mTaS2yNp5_2(.din(w_dff_B_5rJqiBB32_2),.dout(w_dff_B_mTaS2yNp5_2),.clk(gclk));
	jdff dff_B_GETyUF4i3_2(.din(w_dff_B_mTaS2yNp5_2),.dout(w_dff_B_GETyUF4i3_2),.clk(gclk));
	jdff dff_B_3xx9tJ5y5_1(.din(n935),.dout(w_dff_B_3xx9tJ5y5_1),.clk(gclk));
	jdff dff_B_XQYEf3Bs7_2(.din(n832),.dout(w_dff_B_XQYEf3Bs7_2),.clk(gclk));
	jdff dff_B_w2dm33815_2(.din(w_dff_B_XQYEf3Bs7_2),.dout(w_dff_B_w2dm33815_2),.clk(gclk));
	jdff dff_B_wnBR6JA50_2(.din(w_dff_B_w2dm33815_2),.dout(w_dff_B_wnBR6JA50_2),.clk(gclk));
	jdff dff_B_D8xKpJzf6_2(.din(w_dff_B_wnBR6JA50_2),.dout(w_dff_B_D8xKpJzf6_2),.clk(gclk));
	jdff dff_B_XMZRe6bd6_2(.din(w_dff_B_D8xKpJzf6_2),.dout(w_dff_B_XMZRe6bd6_2),.clk(gclk));
	jdff dff_B_xMHIbwiF4_2(.din(w_dff_B_XMZRe6bd6_2),.dout(w_dff_B_xMHIbwiF4_2),.clk(gclk));
	jdff dff_B_x1pnD8RP4_2(.din(w_dff_B_xMHIbwiF4_2),.dout(w_dff_B_x1pnD8RP4_2),.clk(gclk));
	jdff dff_B_WQk8WZbI9_2(.din(w_dff_B_x1pnD8RP4_2),.dout(w_dff_B_WQk8WZbI9_2),.clk(gclk));
	jdff dff_B_9Z23VAxT0_2(.din(w_dff_B_WQk8WZbI9_2),.dout(w_dff_B_9Z23VAxT0_2),.clk(gclk));
	jdff dff_B_SDqwmYCU9_2(.din(w_dff_B_9Z23VAxT0_2),.dout(w_dff_B_SDqwmYCU9_2),.clk(gclk));
	jdff dff_B_pY0hJPWK9_2(.din(w_dff_B_SDqwmYCU9_2),.dout(w_dff_B_pY0hJPWK9_2),.clk(gclk));
	jdff dff_B_LTdyYCPM6_2(.din(w_dff_B_pY0hJPWK9_2),.dout(w_dff_B_LTdyYCPM6_2),.clk(gclk));
	jdff dff_B_HdBg7PPq7_2(.din(w_dff_B_LTdyYCPM6_2),.dout(w_dff_B_HdBg7PPq7_2),.clk(gclk));
	jdff dff_B_9byKDIrc7_2(.din(w_dff_B_HdBg7PPq7_2),.dout(w_dff_B_9byKDIrc7_2),.clk(gclk));
	jdff dff_B_AHT48S058_2(.din(w_dff_B_9byKDIrc7_2),.dout(w_dff_B_AHT48S058_2),.clk(gclk));
	jdff dff_B_cB4Q6WJd3_2(.din(w_dff_B_AHT48S058_2),.dout(w_dff_B_cB4Q6WJd3_2),.clk(gclk));
	jdff dff_B_Z6V9HleY5_2(.din(w_dff_B_cB4Q6WJd3_2),.dout(w_dff_B_Z6V9HleY5_2),.clk(gclk));
	jdff dff_B_xtNDmmBm2_2(.din(w_dff_B_Z6V9HleY5_2),.dout(w_dff_B_xtNDmmBm2_2),.clk(gclk));
	jdff dff_B_nrsyw6Nw7_2(.din(w_dff_B_xtNDmmBm2_2),.dout(w_dff_B_nrsyw6Nw7_2),.clk(gclk));
	jdff dff_B_Frc572ea5_2(.din(w_dff_B_nrsyw6Nw7_2),.dout(w_dff_B_Frc572ea5_2),.clk(gclk));
	jdff dff_B_1htllQC45_2(.din(w_dff_B_Frc572ea5_2),.dout(w_dff_B_1htllQC45_2),.clk(gclk));
	jdff dff_B_XrFlQZ0f1_2(.din(w_dff_B_1htllQC45_2),.dout(w_dff_B_XrFlQZ0f1_2),.clk(gclk));
	jdff dff_B_CsaZPo1K9_2(.din(w_dff_B_XrFlQZ0f1_2),.dout(w_dff_B_CsaZPo1K9_2),.clk(gclk));
	jdff dff_B_9mMRclRs6_2(.din(w_dff_B_CsaZPo1K9_2),.dout(w_dff_B_9mMRclRs6_2),.clk(gclk));
	jdff dff_B_L1plQ7BJ1_2(.din(w_dff_B_9mMRclRs6_2),.dout(w_dff_B_L1plQ7BJ1_2),.clk(gclk));
	jdff dff_B_2ZzMFQ423_2(.din(w_dff_B_L1plQ7BJ1_2),.dout(w_dff_B_2ZzMFQ423_2),.clk(gclk));
	jdff dff_B_1e5eJ58E4_2(.din(w_dff_B_2ZzMFQ423_2),.dout(w_dff_B_1e5eJ58E4_2),.clk(gclk));
	jdff dff_B_b0QFyRaJ4_1(.din(n833),.dout(w_dff_B_b0QFyRaJ4_1),.clk(gclk));
	jdff dff_B_wH2FGRmR6_2(.din(n734),.dout(w_dff_B_wH2FGRmR6_2),.clk(gclk));
	jdff dff_B_7UsRrJa37_2(.din(w_dff_B_wH2FGRmR6_2),.dout(w_dff_B_7UsRrJa37_2),.clk(gclk));
	jdff dff_B_qEwEU1VK5_2(.din(w_dff_B_7UsRrJa37_2),.dout(w_dff_B_qEwEU1VK5_2),.clk(gclk));
	jdff dff_B_KrWbVi1o5_2(.din(w_dff_B_qEwEU1VK5_2),.dout(w_dff_B_KrWbVi1o5_2),.clk(gclk));
	jdff dff_B_OFj3II7e4_2(.din(w_dff_B_KrWbVi1o5_2),.dout(w_dff_B_OFj3II7e4_2),.clk(gclk));
	jdff dff_B_wQuKQmho0_2(.din(w_dff_B_OFj3II7e4_2),.dout(w_dff_B_wQuKQmho0_2),.clk(gclk));
	jdff dff_B_rFM4KIgO3_2(.din(w_dff_B_wQuKQmho0_2),.dout(w_dff_B_rFM4KIgO3_2),.clk(gclk));
	jdff dff_B_KwweXWJv6_2(.din(w_dff_B_rFM4KIgO3_2),.dout(w_dff_B_KwweXWJv6_2),.clk(gclk));
	jdff dff_B_84x0jNk58_2(.din(w_dff_B_KwweXWJv6_2),.dout(w_dff_B_84x0jNk58_2),.clk(gclk));
	jdff dff_B_wmXsjXrg8_2(.din(w_dff_B_84x0jNk58_2),.dout(w_dff_B_wmXsjXrg8_2),.clk(gclk));
	jdff dff_B_zpwBuqvP2_2(.din(w_dff_B_wmXsjXrg8_2),.dout(w_dff_B_zpwBuqvP2_2),.clk(gclk));
	jdff dff_B_sAQQOZ1Q3_2(.din(w_dff_B_zpwBuqvP2_2),.dout(w_dff_B_sAQQOZ1Q3_2),.clk(gclk));
	jdff dff_B_Dl3O1mtC9_2(.din(w_dff_B_sAQQOZ1Q3_2),.dout(w_dff_B_Dl3O1mtC9_2),.clk(gclk));
	jdff dff_B_Yc9nggDa1_2(.din(w_dff_B_Dl3O1mtC9_2),.dout(w_dff_B_Yc9nggDa1_2),.clk(gclk));
	jdff dff_B_4OP5NqJ49_2(.din(w_dff_B_Yc9nggDa1_2),.dout(w_dff_B_4OP5NqJ49_2),.clk(gclk));
	jdff dff_B_k4bqxa922_2(.din(w_dff_B_4OP5NqJ49_2),.dout(w_dff_B_k4bqxa922_2),.clk(gclk));
	jdff dff_B_daLnpbxA3_2(.din(w_dff_B_k4bqxa922_2),.dout(w_dff_B_daLnpbxA3_2),.clk(gclk));
	jdff dff_B_S6m8QAh92_2(.din(w_dff_B_daLnpbxA3_2),.dout(w_dff_B_S6m8QAh92_2),.clk(gclk));
	jdff dff_B_MwqVd59X2_2(.din(w_dff_B_S6m8QAh92_2),.dout(w_dff_B_MwqVd59X2_2),.clk(gclk));
	jdff dff_B_2HiMGl5j1_2(.din(w_dff_B_MwqVd59X2_2),.dout(w_dff_B_2HiMGl5j1_2),.clk(gclk));
	jdff dff_B_yemd9cAo9_2(.din(w_dff_B_2HiMGl5j1_2),.dout(w_dff_B_yemd9cAo9_2),.clk(gclk));
	jdff dff_B_KrDsOy8L9_2(.din(w_dff_B_yemd9cAo9_2),.dout(w_dff_B_KrDsOy8L9_2),.clk(gclk));
	jdff dff_B_6UDR1fBH9_2(.din(w_dff_B_KrDsOy8L9_2),.dout(w_dff_B_6UDR1fBH9_2),.clk(gclk));
	jdff dff_B_bTlMXmHN0_2(.din(w_dff_B_6UDR1fBH9_2),.dout(w_dff_B_bTlMXmHN0_2),.clk(gclk));
	jdff dff_B_a5hMvIXr4_1(.din(n735),.dout(w_dff_B_a5hMvIXr4_1),.clk(gclk));
	jdff dff_B_95TFH98x2_2(.din(n642),.dout(w_dff_B_95TFH98x2_2),.clk(gclk));
	jdff dff_B_FDB44I3s9_2(.din(w_dff_B_95TFH98x2_2),.dout(w_dff_B_FDB44I3s9_2),.clk(gclk));
	jdff dff_B_ZRB8TWo86_2(.din(w_dff_B_FDB44I3s9_2),.dout(w_dff_B_ZRB8TWo86_2),.clk(gclk));
	jdff dff_B_HuVF1xcf4_2(.din(w_dff_B_ZRB8TWo86_2),.dout(w_dff_B_HuVF1xcf4_2),.clk(gclk));
	jdff dff_B_5FPRP90C4_2(.din(w_dff_B_HuVF1xcf4_2),.dout(w_dff_B_5FPRP90C4_2),.clk(gclk));
	jdff dff_B_qSveOskZ7_2(.din(w_dff_B_5FPRP90C4_2),.dout(w_dff_B_qSveOskZ7_2),.clk(gclk));
	jdff dff_B_IRLLnjOa4_2(.din(w_dff_B_qSveOskZ7_2),.dout(w_dff_B_IRLLnjOa4_2),.clk(gclk));
	jdff dff_B_YxIoEKj84_2(.din(w_dff_B_IRLLnjOa4_2),.dout(w_dff_B_YxIoEKj84_2),.clk(gclk));
	jdff dff_B_G6eUWOPl2_2(.din(w_dff_B_YxIoEKj84_2),.dout(w_dff_B_G6eUWOPl2_2),.clk(gclk));
	jdff dff_B_RJY2uDu19_2(.din(w_dff_B_G6eUWOPl2_2),.dout(w_dff_B_RJY2uDu19_2),.clk(gclk));
	jdff dff_B_mQhis6j15_2(.din(w_dff_B_RJY2uDu19_2),.dout(w_dff_B_mQhis6j15_2),.clk(gclk));
	jdff dff_B_vk9FTMO82_2(.din(w_dff_B_mQhis6j15_2),.dout(w_dff_B_vk9FTMO82_2),.clk(gclk));
	jdff dff_B_lLkldlYr8_2(.din(w_dff_B_vk9FTMO82_2),.dout(w_dff_B_lLkldlYr8_2),.clk(gclk));
	jdff dff_B_KmsgppnI8_2(.din(w_dff_B_lLkldlYr8_2),.dout(w_dff_B_KmsgppnI8_2),.clk(gclk));
	jdff dff_B_CVt3WYV58_2(.din(w_dff_B_KmsgppnI8_2),.dout(w_dff_B_CVt3WYV58_2),.clk(gclk));
	jdff dff_B_d5Ww78tP8_2(.din(w_dff_B_CVt3WYV58_2),.dout(w_dff_B_d5Ww78tP8_2),.clk(gclk));
	jdff dff_B_51b1fma64_2(.din(w_dff_B_d5Ww78tP8_2),.dout(w_dff_B_51b1fma64_2),.clk(gclk));
	jdff dff_B_m3qBvm096_2(.din(w_dff_B_51b1fma64_2),.dout(w_dff_B_m3qBvm096_2),.clk(gclk));
	jdff dff_B_gWGqX1cA0_2(.din(w_dff_B_m3qBvm096_2),.dout(w_dff_B_gWGqX1cA0_2),.clk(gclk));
	jdff dff_B_9bJyjAPO7_2(.din(w_dff_B_gWGqX1cA0_2),.dout(w_dff_B_9bJyjAPO7_2),.clk(gclk));
	jdff dff_B_2KqAnSEU2_2(.din(w_dff_B_9bJyjAPO7_2),.dout(w_dff_B_2KqAnSEU2_2),.clk(gclk));
	jdff dff_B_SSFrj5Nk1_1(.din(n643),.dout(w_dff_B_SSFrj5Nk1_1),.clk(gclk));
	jdff dff_B_qFoG6pek1_2(.din(n557),.dout(w_dff_B_qFoG6pek1_2),.clk(gclk));
	jdff dff_B_BC4DsAIz2_2(.din(w_dff_B_qFoG6pek1_2),.dout(w_dff_B_BC4DsAIz2_2),.clk(gclk));
	jdff dff_B_dyvud0fw6_2(.din(w_dff_B_BC4DsAIz2_2),.dout(w_dff_B_dyvud0fw6_2),.clk(gclk));
	jdff dff_B_Z3gK0SMQ1_2(.din(w_dff_B_dyvud0fw6_2),.dout(w_dff_B_Z3gK0SMQ1_2),.clk(gclk));
	jdff dff_B_8zz5iqBf0_2(.din(w_dff_B_Z3gK0SMQ1_2),.dout(w_dff_B_8zz5iqBf0_2),.clk(gclk));
	jdff dff_B_mCLqynJs3_2(.din(w_dff_B_8zz5iqBf0_2),.dout(w_dff_B_mCLqynJs3_2),.clk(gclk));
	jdff dff_B_FBFMEVqD8_2(.din(w_dff_B_mCLqynJs3_2),.dout(w_dff_B_FBFMEVqD8_2),.clk(gclk));
	jdff dff_B_SfHG0bQ89_2(.din(w_dff_B_FBFMEVqD8_2),.dout(w_dff_B_SfHG0bQ89_2),.clk(gclk));
	jdff dff_B_lzBz9qpK8_2(.din(w_dff_B_SfHG0bQ89_2),.dout(w_dff_B_lzBz9qpK8_2),.clk(gclk));
	jdff dff_B_zufUWRD91_2(.din(w_dff_B_lzBz9qpK8_2),.dout(w_dff_B_zufUWRD91_2),.clk(gclk));
	jdff dff_B_wLEgturd6_2(.din(w_dff_B_zufUWRD91_2),.dout(w_dff_B_wLEgturd6_2),.clk(gclk));
	jdff dff_B_orYTpMRz5_2(.din(w_dff_B_wLEgturd6_2),.dout(w_dff_B_orYTpMRz5_2),.clk(gclk));
	jdff dff_B_n0Cmn7y92_2(.din(w_dff_B_orYTpMRz5_2),.dout(w_dff_B_n0Cmn7y92_2),.clk(gclk));
	jdff dff_B_Y6FP9So05_2(.din(w_dff_B_n0Cmn7y92_2),.dout(w_dff_B_Y6FP9So05_2),.clk(gclk));
	jdff dff_B_e38GIF168_2(.din(w_dff_B_Y6FP9So05_2),.dout(w_dff_B_e38GIF168_2),.clk(gclk));
	jdff dff_B_8W6mVw9a0_2(.din(w_dff_B_e38GIF168_2),.dout(w_dff_B_8W6mVw9a0_2),.clk(gclk));
	jdff dff_B_lp1IivzI1_2(.din(w_dff_B_8W6mVw9a0_2),.dout(w_dff_B_lp1IivzI1_2),.clk(gclk));
	jdff dff_B_PIUi5LCX0_2(.din(w_dff_B_lp1IivzI1_2),.dout(w_dff_B_PIUi5LCX0_2),.clk(gclk));
	jdff dff_B_b6JibRo52_1(.din(n558),.dout(w_dff_B_b6JibRo52_1),.clk(gclk));
	jdff dff_B_uDq8J1XC0_2(.din(n479),.dout(w_dff_B_uDq8J1XC0_2),.clk(gclk));
	jdff dff_B_q9b7ZXoW7_2(.din(w_dff_B_uDq8J1XC0_2),.dout(w_dff_B_q9b7ZXoW7_2),.clk(gclk));
	jdff dff_B_guXcKO6u4_2(.din(w_dff_B_q9b7ZXoW7_2),.dout(w_dff_B_guXcKO6u4_2),.clk(gclk));
	jdff dff_B_Jhv0cexv3_2(.din(w_dff_B_guXcKO6u4_2),.dout(w_dff_B_Jhv0cexv3_2),.clk(gclk));
	jdff dff_B_SWTulCdI1_2(.din(w_dff_B_Jhv0cexv3_2),.dout(w_dff_B_SWTulCdI1_2),.clk(gclk));
	jdff dff_B_V5JIIkF60_2(.din(w_dff_B_SWTulCdI1_2),.dout(w_dff_B_V5JIIkF60_2),.clk(gclk));
	jdff dff_B_P7aYFYCH8_2(.din(w_dff_B_V5JIIkF60_2),.dout(w_dff_B_P7aYFYCH8_2),.clk(gclk));
	jdff dff_B_ETEoCqUj7_2(.din(w_dff_B_P7aYFYCH8_2),.dout(w_dff_B_ETEoCqUj7_2),.clk(gclk));
	jdff dff_B_9p4VykO81_2(.din(w_dff_B_ETEoCqUj7_2),.dout(w_dff_B_9p4VykO81_2),.clk(gclk));
	jdff dff_B_Nkvt1q1B3_2(.din(w_dff_B_9p4VykO81_2),.dout(w_dff_B_Nkvt1q1B3_2),.clk(gclk));
	jdff dff_B_gVJ1WyDN5_2(.din(w_dff_B_Nkvt1q1B3_2),.dout(w_dff_B_gVJ1WyDN5_2),.clk(gclk));
	jdff dff_B_kNjXTNPM3_2(.din(w_dff_B_gVJ1WyDN5_2),.dout(w_dff_B_kNjXTNPM3_2),.clk(gclk));
	jdff dff_B_17tYhwAN7_2(.din(w_dff_B_kNjXTNPM3_2),.dout(w_dff_B_17tYhwAN7_2),.clk(gclk));
	jdff dff_B_sIc9ZKYP3_2(.din(w_dff_B_17tYhwAN7_2),.dout(w_dff_B_sIc9ZKYP3_2),.clk(gclk));
	jdff dff_B_74u6g0wf4_2(.din(w_dff_B_sIc9ZKYP3_2),.dout(w_dff_B_74u6g0wf4_2),.clk(gclk));
	jdff dff_B_HyF84s1z6_1(.din(n480),.dout(w_dff_B_HyF84s1z6_1),.clk(gclk));
	jdff dff_B_QJgOlO5S3_2(.din(n408),.dout(w_dff_B_QJgOlO5S3_2),.clk(gclk));
	jdff dff_B_VC5AI2cE2_2(.din(w_dff_B_QJgOlO5S3_2),.dout(w_dff_B_VC5AI2cE2_2),.clk(gclk));
	jdff dff_B_6jvrfecC2_2(.din(w_dff_B_VC5AI2cE2_2),.dout(w_dff_B_6jvrfecC2_2),.clk(gclk));
	jdff dff_B_LHqolNIR7_2(.din(w_dff_B_6jvrfecC2_2),.dout(w_dff_B_LHqolNIR7_2),.clk(gclk));
	jdff dff_B_Lc13rufq5_2(.din(w_dff_B_LHqolNIR7_2),.dout(w_dff_B_Lc13rufq5_2),.clk(gclk));
	jdff dff_B_0iV3cD4D1_2(.din(w_dff_B_Lc13rufq5_2),.dout(w_dff_B_0iV3cD4D1_2),.clk(gclk));
	jdff dff_B_eslJJmNt6_2(.din(w_dff_B_0iV3cD4D1_2),.dout(w_dff_B_eslJJmNt6_2),.clk(gclk));
	jdff dff_B_5Mytq3hu9_2(.din(w_dff_B_eslJJmNt6_2),.dout(w_dff_B_5Mytq3hu9_2),.clk(gclk));
	jdff dff_B_15wlhsPs1_2(.din(w_dff_B_5Mytq3hu9_2),.dout(w_dff_B_15wlhsPs1_2),.clk(gclk));
	jdff dff_B_ZadxiPV94_2(.din(w_dff_B_15wlhsPs1_2),.dout(w_dff_B_ZadxiPV94_2),.clk(gclk));
	jdff dff_B_kbKgaLLY7_2(.din(w_dff_B_ZadxiPV94_2),.dout(w_dff_B_kbKgaLLY7_2),.clk(gclk));
	jdff dff_B_h9fjyNnY5_2(.din(w_dff_B_kbKgaLLY7_2),.dout(w_dff_B_h9fjyNnY5_2),.clk(gclk));
	jdff dff_B_MeQzjXfG9_1(.din(n409),.dout(w_dff_B_MeQzjXfG9_1),.clk(gclk));
	jdff dff_B_ZejeJu0H2_2(.din(n345),.dout(w_dff_B_ZejeJu0H2_2),.clk(gclk));
	jdff dff_B_9ommu0Cu8_2(.din(w_dff_B_ZejeJu0H2_2),.dout(w_dff_B_9ommu0Cu8_2),.clk(gclk));
	jdff dff_B_aXbMf3v88_2(.din(w_dff_B_9ommu0Cu8_2),.dout(w_dff_B_aXbMf3v88_2),.clk(gclk));
	jdff dff_B_hRxqR5J26_2(.din(w_dff_B_aXbMf3v88_2),.dout(w_dff_B_hRxqR5J26_2),.clk(gclk));
	jdff dff_B_3wDR3Q5p8_2(.din(w_dff_B_hRxqR5J26_2),.dout(w_dff_B_3wDR3Q5p8_2),.clk(gclk));
	jdff dff_B_AhWySDnr8_2(.din(w_dff_B_3wDR3Q5p8_2),.dout(w_dff_B_AhWySDnr8_2),.clk(gclk));
	jdff dff_B_MHIfGEIW1_2(.din(w_dff_B_AhWySDnr8_2),.dout(w_dff_B_MHIfGEIW1_2),.clk(gclk));
	jdff dff_B_TIHxiZXZ5_2(.din(w_dff_B_MHIfGEIW1_2),.dout(w_dff_B_TIHxiZXZ5_2),.clk(gclk));
	jdff dff_B_UKDO5yzq0_2(.din(w_dff_B_TIHxiZXZ5_2),.dout(w_dff_B_UKDO5yzq0_2),.clk(gclk));
	jdff dff_B_o71vjIz19_2(.din(n366),.dout(w_dff_B_o71vjIz19_2),.clk(gclk));
	jdff dff_B_d4C0Djht4_1(.din(n346),.dout(w_dff_B_d4C0Djht4_1),.clk(gclk));
	jdff dff_B_QLmmHdBd3_2(.din(n289),.dout(w_dff_B_QLmmHdBd3_2),.clk(gclk));
	jdff dff_B_AD6FBGMr9_2(.din(w_dff_B_QLmmHdBd3_2),.dout(w_dff_B_AD6FBGMr9_2),.clk(gclk));
	jdff dff_B_yU97FjGZ8_2(.din(w_dff_B_AD6FBGMr9_2),.dout(w_dff_B_yU97FjGZ8_2),.clk(gclk));
	jdff dff_B_nQ8IACQD3_2(.din(w_dff_B_yU97FjGZ8_2),.dout(w_dff_B_nQ8IACQD3_2),.clk(gclk));
	jdff dff_B_aOg66IsC9_2(.din(w_dff_B_nQ8IACQD3_2),.dout(w_dff_B_aOg66IsC9_2),.clk(gclk));
	jdff dff_B_nzEs7aAK5_2(.din(w_dff_B_aOg66IsC9_2),.dout(w_dff_B_nzEs7aAK5_2),.clk(gclk));
	jdff dff_B_9ig1YyJM9_2(.din(n303),.dout(w_dff_B_9ig1YyJM9_2),.clk(gclk));
	jdff dff_B_PO4Y0hsc6_2(.din(n241),.dout(w_dff_B_PO4Y0hsc6_2),.clk(gclk));
	jdff dff_B_PDaul29w4_2(.din(w_dff_B_PO4Y0hsc6_2),.dout(w_dff_B_PDaul29w4_2),.clk(gclk));
	jdff dff_B_moe5ArhA2_2(.din(w_dff_B_PDaul29w4_2),.dout(w_dff_B_moe5ArhA2_2),.clk(gclk));
	jdff dff_B_R06sGySs5_0(.din(n246),.dout(w_dff_B_R06sGySs5_0),.clk(gclk));
	jdff dff_A_avPaiqt82_0(.dout(w_n196_0[0]),.din(w_dff_A_avPaiqt82_0),.clk(gclk));
	jdff dff_A_d0yTcVi09_0(.dout(w_dff_A_avPaiqt82_0),.din(w_dff_A_d0yTcVi09_0),.clk(gclk));
	jdff dff_A_lmAUvAnN9_1(.dout(w_n196_0[1]),.din(w_dff_A_lmAUvAnN9_1),.clk(gclk));
	jdff dff_A_Pm0Nd7zt9_1(.dout(w_dff_A_lmAUvAnN9_1),.din(w_dff_A_Pm0Nd7zt9_1),.clk(gclk));
	jdff dff_B_7IYrndFR5_2(.din(n1465),.dout(w_dff_B_7IYrndFR5_2),.clk(gclk));
	jdff dff_B_fcHIml3A7_1(.din(n1463),.dout(w_dff_B_fcHIml3A7_1),.clk(gclk));
	jdff dff_B_VByecPze9_2(.din(n1390),.dout(w_dff_B_VByecPze9_2),.clk(gclk));
	jdff dff_B_bnwwtrCn4_2(.din(w_dff_B_VByecPze9_2),.dout(w_dff_B_bnwwtrCn4_2),.clk(gclk));
	jdff dff_B_qT3ZAFbp1_2(.din(w_dff_B_bnwwtrCn4_2),.dout(w_dff_B_qT3ZAFbp1_2),.clk(gclk));
	jdff dff_B_uhMyfmmT5_2(.din(w_dff_B_qT3ZAFbp1_2),.dout(w_dff_B_uhMyfmmT5_2),.clk(gclk));
	jdff dff_B_QEK7rfsY1_2(.din(w_dff_B_uhMyfmmT5_2),.dout(w_dff_B_QEK7rfsY1_2),.clk(gclk));
	jdff dff_B_9vpFs3On0_2(.din(w_dff_B_QEK7rfsY1_2),.dout(w_dff_B_9vpFs3On0_2),.clk(gclk));
	jdff dff_B_YATb2Jj04_2(.din(w_dff_B_9vpFs3On0_2),.dout(w_dff_B_YATb2Jj04_2),.clk(gclk));
	jdff dff_B_EUSs6NCu4_2(.din(w_dff_B_YATb2Jj04_2),.dout(w_dff_B_EUSs6NCu4_2),.clk(gclk));
	jdff dff_B_HoK8i75Z1_2(.din(w_dff_B_EUSs6NCu4_2),.dout(w_dff_B_HoK8i75Z1_2),.clk(gclk));
	jdff dff_B_QlNHCHsO0_2(.din(w_dff_B_HoK8i75Z1_2),.dout(w_dff_B_QlNHCHsO0_2),.clk(gclk));
	jdff dff_B_lzz0N8Uc5_2(.din(w_dff_B_QlNHCHsO0_2),.dout(w_dff_B_lzz0N8Uc5_2),.clk(gclk));
	jdff dff_B_pPBQNrSV0_2(.din(w_dff_B_lzz0N8Uc5_2),.dout(w_dff_B_pPBQNrSV0_2),.clk(gclk));
	jdff dff_B_Bs8SAgra7_2(.din(w_dff_B_pPBQNrSV0_2),.dout(w_dff_B_Bs8SAgra7_2),.clk(gclk));
	jdff dff_B_Q2eQFoDZ2_2(.din(w_dff_B_Bs8SAgra7_2),.dout(w_dff_B_Q2eQFoDZ2_2),.clk(gclk));
	jdff dff_B_4e4g0vIF9_2(.din(w_dff_B_Q2eQFoDZ2_2),.dout(w_dff_B_4e4g0vIF9_2),.clk(gclk));
	jdff dff_B_NIctntP14_2(.din(w_dff_B_4e4g0vIF9_2),.dout(w_dff_B_NIctntP14_2),.clk(gclk));
	jdff dff_B_DPkKJCks4_2(.din(w_dff_B_NIctntP14_2),.dout(w_dff_B_DPkKJCks4_2),.clk(gclk));
	jdff dff_B_Sg6DnKlH5_2(.din(w_dff_B_DPkKJCks4_2),.dout(w_dff_B_Sg6DnKlH5_2),.clk(gclk));
	jdff dff_B_m6rfshPa9_2(.din(w_dff_B_Sg6DnKlH5_2),.dout(w_dff_B_m6rfshPa9_2),.clk(gclk));
	jdff dff_B_kv0gVde97_2(.din(w_dff_B_m6rfshPa9_2),.dout(w_dff_B_kv0gVde97_2),.clk(gclk));
	jdff dff_B_LYAK9hG93_2(.din(w_dff_B_kv0gVde97_2),.dout(w_dff_B_LYAK9hG93_2),.clk(gclk));
	jdff dff_B_3nU1rMaH3_2(.din(w_dff_B_LYAK9hG93_2),.dout(w_dff_B_3nU1rMaH3_2),.clk(gclk));
	jdff dff_B_Yvk8M88Y8_2(.din(w_dff_B_3nU1rMaH3_2),.dout(w_dff_B_Yvk8M88Y8_2),.clk(gclk));
	jdff dff_B_qow4P8zI1_2(.din(w_dff_B_Yvk8M88Y8_2),.dout(w_dff_B_qow4P8zI1_2),.clk(gclk));
	jdff dff_B_zy8II2T83_2(.din(w_dff_B_qow4P8zI1_2),.dout(w_dff_B_zy8II2T83_2),.clk(gclk));
	jdff dff_B_hXMnjQfh8_2(.din(w_dff_B_zy8II2T83_2),.dout(w_dff_B_hXMnjQfh8_2),.clk(gclk));
	jdff dff_B_QkH2Hj617_2(.din(w_dff_B_hXMnjQfh8_2),.dout(w_dff_B_QkH2Hj617_2),.clk(gclk));
	jdff dff_B_aBGDm4q65_2(.din(w_dff_B_QkH2Hj617_2),.dout(w_dff_B_aBGDm4q65_2),.clk(gclk));
	jdff dff_B_9YmMe76O7_2(.din(w_dff_B_aBGDm4q65_2),.dout(w_dff_B_9YmMe76O7_2),.clk(gclk));
	jdff dff_B_gtvk1xKi7_2(.din(w_dff_B_9YmMe76O7_2),.dout(w_dff_B_gtvk1xKi7_2),.clk(gclk));
	jdff dff_B_SPqnErfz3_2(.din(w_dff_B_gtvk1xKi7_2),.dout(w_dff_B_SPqnErfz3_2),.clk(gclk));
	jdff dff_B_iVZ44Ixp2_2(.din(w_dff_B_SPqnErfz3_2),.dout(w_dff_B_iVZ44Ixp2_2),.clk(gclk));
	jdff dff_B_a4Cj5tGN0_2(.din(w_dff_B_iVZ44Ixp2_2),.dout(w_dff_B_a4Cj5tGN0_2),.clk(gclk));
	jdff dff_B_gdkYer2Z1_2(.din(w_dff_B_a4Cj5tGN0_2),.dout(w_dff_B_gdkYer2Z1_2),.clk(gclk));
	jdff dff_B_zJSwEd6f6_2(.din(w_dff_B_gdkYer2Z1_2),.dout(w_dff_B_zJSwEd6f6_2),.clk(gclk));
	jdff dff_B_OQ9pBsmO5_2(.din(w_dff_B_zJSwEd6f6_2),.dout(w_dff_B_OQ9pBsmO5_2),.clk(gclk));
	jdff dff_B_vfvCQtii6_2(.din(w_dff_B_OQ9pBsmO5_2),.dout(w_dff_B_vfvCQtii6_2),.clk(gclk));
	jdff dff_B_N5nte4gK0_2(.din(w_dff_B_vfvCQtii6_2),.dout(w_dff_B_N5nte4gK0_2),.clk(gclk));
	jdff dff_B_vaU8AVxB7_2(.din(w_dff_B_N5nte4gK0_2),.dout(w_dff_B_vaU8AVxB7_2),.clk(gclk));
	jdff dff_B_drAzDmhn5_2(.din(w_dff_B_vaU8AVxB7_2),.dout(w_dff_B_drAzDmhn5_2),.clk(gclk));
	jdff dff_B_3tOTKcic8_2(.din(w_dff_B_drAzDmhn5_2),.dout(w_dff_B_3tOTKcic8_2),.clk(gclk));
	jdff dff_B_GSLVi2KG7_2(.din(w_dff_B_3tOTKcic8_2),.dout(w_dff_B_GSLVi2KG7_2),.clk(gclk));
	jdff dff_B_0bc0jAd24_2(.din(w_dff_B_GSLVi2KG7_2),.dout(w_dff_B_0bc0jAd24_2),.clk(gclk));
	jdff dff_B_fZkY1zIB6_2(.din(w_dff_B_0bc0jAd24_2),.dout(w_dff_B_fZkY1zIB6_2),.clk(gclk));
	jdff dff_B_Pd21kpZx1_2(.din(w_dff_B_fZkY1zIB6_2),.dout(w_dff_B_Pd21kpZx1_2),.clk(gclk));
	jdff dff_B_xAz4mD5f3_1(.din(n1391),.dout(w_dff_B_xAz4mD5f3_1),.clk(gclk));
	jdff dff_B_q6BFgqL85_2(.din(n1312),.dout(w_dff_B_q6BFgqL85_2),.clk(gclk));
	jdff dff_B_jigvGq0e2_2(.din(w_dff_B_q6BFgqL85_2),.dout(w_dff_B_jigvGq0e2_2),.clk(gclk));
	jdff dff_B_dVV9qFXZ5_2(.din(w_dff_B_jigvGq0e2_2),.dout(w_dff_B_dVV9qFXZ5_2),.clk(gclk));
	jdff dff_B_qssjqL4Q9_2(.din(w_dff_B_dVV9qFXZ5_2),.dout(w_dff_B_qssjqL4Q9_2),.clk(gclk));
	jdff dff_B_sQ7DaFdy4_2(.din(w_dff_B_qssjqL4Q9_2),.dout(w_dff_B_sQ7DaFdy4_2),.clk(gclk));
	jdff dff_B_6MDUZfcK1_2(.din(w_dff_B_sQ7DaFdy4_2),.dout(w_dff_B_6MDUZfcK1_2),.clk(gclk));
	jdff dff_B_UruRfHuH3_2(.din(w_dff_B_6MDUZfcK1_2),.dout(w_dff_B_UruRfHuH3_2),.clk(gclk));
	jdff dff_B_44iIadLG0_2(.din(w_dff_B_UruRfHuH3_2),.dout(w_dff_B_44iIadLG0_2),.clk(gclk));
	jdff dff_B_pFGvHN1P6_2(.din(w_dff_B_44iIadLG0_2),.dout(w_dff_B_pFGvHN1P6_2),.clk(gclk));
	jdff dff_B_Jwm96ixk5_2(.din(w_dff_B_pFGvHN1P6_2),.dout(w_dff_B_Jwm96ixk5_2),.clk(gclk));
	jdff dff_B_MVuqNFAQ4_2(.din(w_dff_B_Jwm96ixk5_2),.dout(w_dff_B_MVuqNFAQ4_2),.clk(gclk));
	jdff dff_B_LJ5MIyFT5_2(.din(w_dff_B_MVuqNFAQ4_2),.dout(w_dff_B_LJ5MIyFT5_2),.clk(gclk));
	jdff dff_B_olNavd7w7_2(.din(w_dff_B_LJ5MIyFT5_2),.dout(w_dff_B_olNavd7w7_2),.clk(gclk));
	jdff dff_B_hnMyeiQQ8_2(.din(w_dff_B_olNavd7w7_2),.dout(w_dff_B_hnMyeiQQ8_2),.clk(gclk));
	jdff dff_B_zB8CuPwy5_2(.din(w_dff_B_hnMyeiQQ8_2),.dout(w_dff_B_zB8CuPwy5_2),.clk(gclk));
	jdff dff_B_DnGTPm9q1_2(.din(w_dff_B_zB8CuPwy5_2),.dout(w_dff_B_DnGTPm9q1_2),.clk(gclk));
	jdff dff_B_qWJRcS0Q2_2(.din(w_dff_B_DnGTPm9q1_2),.dout(w_dff_B_qWJRcS0Q2_2),.clk(gclk));
	jdff dff_B_iqPujPyG7_2(.din(w_dff_B_qWJRcS0Q2_2),.dout(w_dff_B_iqPujPyG7_2),.clk(gclk));
	jdff dff_B_jAzmZZl82_2(.din(w_dff_B_iqPujPyG7_2),.dout(w_dff_B_jAzmZZl82_2),.clk(gclk));
	jdff dff_B_O6SonGJW2_2(.din(w_dff_B_jAzmZZl82_2),.dout(w_dff_B_O6SonGJW2_2),.clk(gclk));
	jdff dff_B_RPAuD1L04_2(.din(w_dff_B_O6SonGJW2_2),.dout(w_dff_B_RPAuD1L04_2),.clk(gclk));
	jdff dff_B_imRTaY8j3_2(.din(w_dff_B_RPAuD1L04_2),.dout(w_dff_B_imRTaY8j3_2),.clk(gclk));
	jdff dff_B_9Fyvj60o4_2(.din(w_dff_B_imRTaY8j3_2),.dout(w_dff_B_9Fyvj60o4_2),.clk(gclk));
	jdff dff_B_aqEN59Os0_2(.din(w_dff_B_9Fyvj60o4_2),.dout(w_dff_B_aqEN59Os0_2),.clk(gclk));
	jdff dff_B_2UUaVsUM1_2(.din(w_dff_B_aqEN59Os0_2),.dout(w_dff_B_2UUaVsUM1_2),.clk(gclk));
	jdff dff_B_kfFmmocH7_2(.din(w_dff_B_2UUaVsUM1_2),.dout(w_dff_B_kfFmmocH7_2),.clk(gclk));
	jdff dff_B_zFGf6PEK0_2(.din(w_dff_B_kfFmmocH7_2),.dout(w_dff_B_zFGf6PEK0_2),.clk(gclk));
	jdff dff_B_YEw0aEIl7_2(.din(w_dff_B_zFGf6PEK0_2),.dout(w_dff_B_YEw0aEIl7_2),.clk(gclk));
	jdff dff_B_yIvWOSUj2_2(.din(w_dff_B_YEw0aEIl7_2),.dout(w_dff_B_yIvWOSUj2_2),.clk(gclk));
	jdff dff_B_Kplq0gJX7_2(.din(w_dff_B_yIvWOSUj2_2),.dout(w_dff_B_Kplq0gJX7_2),.clk(gclk));
	jdff dff_B_nkLYM3ov8_2(.din(w_dff_B_Kplq0gJX7_2),.dout(w_dff_B_nkLYM3ov8_2),.clk(gclk));
	jdff dff_B_Gwh5F2ak5_2(.din(w_dff_B_nkLYM3ov8_2),.dout(w_dff_B_Gwh5F2ak5_2),.clk(gclk));
	jdff dff_B_mZJnrehT5_2(.din(w_dff_B_Gwh5F2ak5_2),.dout(w_dff_B_mZJnrehT5_2),.clk(gclk));
	jdff dff_B_WTzdh0vQ9_2(.din(w_dff_B_mZJnrehT5_2),.dout(w_dff_B_WTzdh0vQ9_2),.clk(gclk));
	jdff dff_B_oyip6Zpf3_2(.din(w_dff_B_WTzdh0vQ9_2),.dout(w_dff_B_oyip6Zpf3_2),.clk(gclk));
	jdff dff_B_unzYtWQN5_2(.din(w_dff_B_oyip6Zpf3_2),.dout(w_dff_B_unzYtWQN5_2),.clk(gclk));
	jdff dff_B_cvWtVvmy8_2(.din(w_dff_B_unzYtWQN5_2),.dout(w_dff_B_cvWtVvmy8_2),.clk(gclk));
	jdff dff_B_RSoabqlo7_2(.din(w_dff_B_cvWtVvmy8_2),.dout(w_dff_B_RSoabqlo7_2),.clk(gclk));
	jdff dff_B_SN2A4cA76_2(.din(w_dff_B_RSoabqlo7_2),.dout(w_dff_B_SN2A4cA76_2),.clk(gclk));
	jdff dff_B_tgvlIUag2_2(.din(w_dff_B_SN2A4cA76_2),.dout(w_dff_B_tgvlIUag2_2),.clk(gclk));
	jdff dff_B_p1ySQhIb4_1(.din(n1313),.dout(w_dff_B_p1ySQhIb4_1),.clk(gclk));
	jdff dff_B_0jZhwfd52_2(.din(n1227),.dout(w_dff_B_0jZhwfd52_2),.clk(gclk));
	jdff dff_B_bwv6OI9X1_2(.din(w_dff_B_0jZhwfd52_2),.dout(w_dff_B_bwv6OI9X1_2),.clk(gclk));
	jdff dff_B_w2r9OyeU9_2(.din(w_dff_B_bwv6OI9X1_2),.dout(w_dff_B_w2r9OyeU9_2),.clk(gclk));
	jdff dff_B_uJ3TkUiB6_2(.din(w_dff_B_w2r9OyeU9_2),.dout(w_dff_B_uJ3TkUiB6_2),.clk(gclk));
	jdff dff_B_iQ6HjADO4_2(.din(w_dff_B_uJ3TkUiB6_2),.dout(w_dff_B_iQ6HjADO4_2),.clk(gclk));
	jdff dff_B_oSJSHojw6_2(.din(w_dff_B_iQ6HjADO4_2),.dout(w_dff_B_oSJSHojw6_2),.clk(gclk));
	jdff dff_B_8GMGOIep7_2(.din(w_dff_B_oSJSHojw6_2),.dout(w_dff_B_8GMGOIep7_2),.clk(gclk));
	jdff dff_B_WlWy4VaC6_2(.din(w_dff_B_8GMGOIep7_2),.dout(w_dff_B_WlWy4VaC6_2),.clk(gclk));
	jdff dff_B_heGH44ag4_2(.din(w_dff_B_WlWy4VaC6_2),.dout(w_dff_B_heGH44ag4_2),.clk(gclk));
	jdff dff_B_4PqX7Zab3_2(.din(w_dff_B_heGH44ag4_2),.dout(w_dff_B_4PqX7Zab3_2),.clk(gclk));
	jdff dff_B_lpC4r68j0_2(.din(w_dff_B_4PqX7Zab3_2),.dout(w_dff_B_lpC4r68j0_2),.clk(gclk));
	jdff dff_B_LXd1zZoD3_2(.din(w_dff_B_lpC4r68j0_2),.dout(w_dff_B_LXd1zZoD3_2),.clk(gclk));
	jdff dff_B_BiXd18tC1_2(.din(w_dff_B_LXd1zZoD3_2),.dout(w_dff_B_BiXd18tC1_2),.clk(gclk));
	jdff dff_B_CawyenJ93_2(.din(w_dff_B_BiXd18tC1_2),.dout(w_dff_B_CawyenJ93_2),.clk(gclk));
	jdff dff_B_CFu21fDh7_2(.din(w_dff_B_CawyenJ93_2),.dout(w_dff_B_CFu21fDh7_2),.clk(gclk));
	jdff dff_B_omETCELq1_2(.din(w_dff_B_CFu21fDh7_2),.dout(w_dff_B_omETCELq1_2),.clk(gclk));
	jdff dff_B_iUBFLVxG4_2(.din(w_dff_B_omETCELq1_2),.dout(w_dff_B_iUBFLVxG4_2),.clk(gclk));
	jdff dff_B_IEFrqQnV0_2(.din(w_dff_B_iUBFLVxG4_2),.dout(w_dff_B_IEFrqQnV0_2),.clk(gclk));
	jdff dff_B_CdsExHPx0_2(.din(w_dff_B_IEFrqQnV0_2),.dout(w_dff_B_CdsExHPx0_2),.clk(gclk));
	jdff dff_B_W8nbYeAN8_2(.din(w_dff_B_CdsExHPx0_2),.dout(w_dff_B_W8nbYeAN8_2),.clk(gclk));
	jdff dff_B_Rwq1Dclc9_2(.din(w_dff_B_W8nbYeAN8_2),.dout(w_dff_B_Rwq1Dclc9_2),.clk(gclk));
	jdff dff_B_Ja0QR4Ji5_2(.din(w_dff_B_Rwq1Dclc9_2),.dout(w_dff_B_Ja0QR4Ji5_2),.clk(gclk));
	jdff dff_B_97D0QIxU7_2(.din(w_dff_B_Ja0QR4Ji5_2),.dout(w_dff_B_97D0QIxU7_2),.clk(gclk));
	jdff dff_B_gqzqYgfg4_2(.din(w_dff_B_97D0QIxU7_2),.dout(w_dff_B_gqzqYgfg4_2),.clk(gclk));
	jdff dff_B_Fx2RNUbk9_2(.din(w_dff_B_gqzqYgfg4_2),.dout(w_dff_B_Fx2RNUbk9_2),.clk(gclk));
	jdff dff_B_XxquX4TF3_2(.din(w_dff_B_Fx2RNUbk9_2),.dout(w_dff_B_XxquX4TF3_2),.clk(gclk));
	jdff dff_B_DsH4y2Yt3_2(.din(w_dff_B_XxquX4TF3_2),.dout(w_dff_B_DsH4y2Yt3_2),.clk(gclk));
	jdff dff_B_UMuBHyn88_2(.din(w_dff_B_DsH4y2Yt3_2),.dout(w_dff_B_UMuBHyn88_2),.clk(gclk));
	jdff dff_B_erApfxOA6_2(.din(w_dff_B_UMuBHyn88_2),.dout(w_dff_B_erApfxOA6_2),.clk(gclk));
	jdff dff_B_u2xWP5EJ2_2(.din(w_dff_B_erApfxOA6_2),.dout(w_dff_B_u2xWP5EJ2_2),.clk(gclk));
	jdff dff_B_OvQo1C3o7_2(.din(w_dff_B_u2xWP5EJ2_2),.dout(w_dff_B_OvQo1C3o7_2),.clk(gclk));
	jdff dff_B_Ogqofr107_2(.din(w_dff_B_OvQo1C3o7_2),.dout(w_dff_B_Ogqofr107_2),.clk(gclk));
	jdff dff_B_2nNPAo0D7_2(.din(w_dff_B_Ogqofr107_2),.dout(w_dff_B_2nNPAo0D7_2),.clk(gclk));
	jdff dff_B_Jd6l7w2P9_2(.din(w_dff_B_2nNPAo0D7_2),.dout(w_dff_B_Jd6l7w2P9_2),.clk(gclk));
	jdff dff_B_qUd31gLq9_2(.din(w_dff_B_Jd6l7w2P9_2),.dout(w_dff_B_qUd31gLq9_2),.clk(gclk));
	jdff dff_B_gwwqRqOS0_2(.din(w_dff_B_qUd31gLq9_2),.dout(w_dff_B_gwwqRqOS0_2),.clk(gclk));
	jdff dff_B_2TijpYi78_2(.din(w_dff_B_gwwqRqOS0_2),.dout(w_dff_B_2TijpYi78_2),.clk(gclk));
	jdff dff_B_Ncrix9Co4_1(.din(n1228),.dout(w_dff_B_Ncrix9Co4_1),.clk(gclk));
	jdff dff_B_Y8wFsNR74_2(.din(n1136),.dout(w_dff_B_Y8wFsNR74_2),.clk(gclk));
	jdff dff_B_Vg88ocSZ6_2(.din(w_dff_B_Y8wFsNR74_2),.dout(w_dff_B_Vg88ocSZ6_2),.clk(gclk));
	jdff dff_B_zV0LuOs57_2(.din(w_dff_B_Vg88ocSZ6_2),.dout(w_dff_B_zV0LuOs57_2),.clk(gclk));
	jdff dff_B_hMxudX500_2(.din(w_dff_B_zV0LuOs57_2),.dout(w_dff_B_hMxudX500_2),.clk(gclk));
	jdff dff_B_s8ceWCYO4_2(.din(w_dff_B_hMxudX500_2),.dout(w_dff_B_s8ceWCYO4_2),.clk(gclk));
	jdff dff_B_oyf71azQ6_2(.din(w_dff_B_s8ceWCYO4_2),.dout(w_dff_B_oyf71azQ6_2),.clk(gclk));
	jdff dff_B_Hap07XHV0_2(.din(w_dff_B_oyf71azQ6_2),.dout(w_dff_B_Hap07XHV0_2),.clk(gclk));
	jdff dff_B_XAircJLx3_2(.din(w_dff_B_Hap07XHV0_2),.dout(w_dff_B_XAircJLx3_2),.clk(gclk));
	jdff dff_B_2FoMNE2y9_2(.din(w_dff_B_XAircJLx3_2),.dout(w_dff_B_2FoMNE2y9_2),.clk(gclk));
	jdff dff_B_pY9HX9700_2(.din(w_dff_B_2FoMNE2y9_2),.dout(w_dff_B_pY9HX9700_2),.clk(gclk));
	jdff dff_B_7ZG8p6cb1_2(.din(w_dff_B_pY9HX9700_2),.dout(w_dff_B_7ZG8p6cb1_2),.clk(gclk));
	jdff dff_B_txF6M97S4_2(.din(w_dff_B_7ZG8p6cb1_2),.dout(w_dff_B_txF6M97S4_2),.clk(gclk));
	jdff dff_B_onCvetXI5_2(.din(w_dff_B_txF6M97S4_2),.dout(w_dff_B_onCvetXI5_2),.clk(gclk));
	jdff dff_B_DRd4W0KS2_2(.din(w_dff_B_onCvetXI5_2),.dout(w_dff_B_DRd4W0KS2_2),.clk(gclk));
	jdff dff_B_wHqNAGMY0_2(.din(w_dff_B_DRd4W0KS2_2),.dout(w_dff_B_wHqNAGMY0_2),.clk(gclk));
	jdff dff_B_opYE9eWC2_2(.din(w_dff_B_wHqNAGMY0_2),.dout(w_dff_B_opYE9eWC2_2),.clk(gclk));
	jdff dff_B_sgkrrRGD7_2(.din(w_dff_B_opYE9eWC2_2),.dout(w_dff_B_sgkrrRGD7_2),.clk(gclk));
	jdff dff_B_IVCPit3L1_2(.din(w_dff_B_sgkrrRGD7_2),.dout(w_dff_B_IVCPit3L1_2),.clk(gclk));
	jdff dff_B_5KKygy3C9_2(.din(w_dff_B_IVCPit3L1_2),.dout(w_dff_B_5KKygy3C9_2),.clk(gclk));
	jdff dff_B_T2X5e5yQ8_2(.din(w_dff_B_5KKygy3C9_2),.dout(w_dff_B_T2X5e5yQ8_2),.clk(gclk));
	jdff dff_B_zKuZnUrH6_2(.din(w_dff_B_T2X5e5yQ8_2),.dout(w_dff_B_zKuZnUrH6_2),.clk(gclk));
	jdff dff_B_Ef1DAYzs8_2(.din(w_dff_B_zKuZnUrH6_2),.dout(w_dff_B_Ef1DAYzs8_2),.clk(gclk));
	jdff dff_B_Kpk2ZwEA6_2(.din(w_dff_B_Ef1DAYzs8_2),.dout(w_dff_B_Kpk2ZwEA6_2),.clk(gclk));
	jdff dff_B_h7zqUyKf9_2(.din(w_dff_B_Kpk2ZwEA6_2),.dout(w_dff_B_h7zqUyKf9_2),.clk(gclk));
	jdff dff_B_FEBK82sH3_2(.din(w_dff_B_h7zqUyKf9_2),.dout(w_dff_B_FEBK82sH3_2),.clk(gclk));
	jdff dff_B_K0zobonR7_2(.din(w_dff_B_FEBK82sH3_2),.dout(w_dff_B_K0zobonR7_2),.clk(gclk));
	jdff dff_B_BEqFulR19_2(.din(w_dff_B_K0zobonR7_2),.dout(w_dff_B_BEqFulR19_2),.clk(gclk));
	jdff dff_B_C0fQjyRv5_2(.din(w_dff_B_BEqFulR19_2),.dout(w_dff_B_C0fQjyRv5_2),.clk(gclk));
	jdff dff_B_bVOlXeOK6_2(.din(w_dff_B_C0fQjyRv5_2),.dout(w_dff_B_bVOlXeOK6_2),.clk(gclk));
	jdff dff_B_2aCrStZ59_2(.din(w_dff_B_bVOlXeOK6_2),.dout(w_dff_B_2aCrStZ59_2),.clk(gclk));
	jdff dff_B_VvNG1HuI7_2(.din(w_dff_B_2aCrStZ59_2),.dout(w_dff_B_VvNG1HuI7_2),.clk(gclk));
	jdff dff_B_5EEBvNvP7_2(.din(w_dff_B_VvNG1HuI7_2),.dout(w_dff_B_5EEBvNvP7_2),.clk(gclk));
	jdff dff_B_lgYGEJcS8_2(.din(w_dff_B_5EEBvNvP7_2),.dout(w_dff_B_lgYGEJcS8_2),.clk(gclk));
	jdff dff_B_O7NpO5ou1_2(.din(w_dff_B_lgYGEJcS8_2),.dout(w_dff_B_O7NpO5ou1_2),.clk(gclk));
	jdff dff_B_mSgxvJiU9_1(.din(n1137),.dout(w_dff_B_mSgxvJiU9_1),.clk(gclk));
	jdff dff_B_U1c0qcFe6_2(.din(n1038),.dout(w_dff_B_U1c0qcFe6_2),.clk(gclk));
	jdff dff_B_dspjIlW31_2(.din(w_dff_B_U1c0qcFe6_2),.dout(w_dff_B_dspjIlW31_2),.clk(gclk));
	jdff dff_B_yqWxRizk1_2(.din(w_dff_B_dspjIlW31_2),.dout(w_dff_B_yqWxRizk1_2),.clk(gclk));
	jdff dff_B_iAoyfUpp6_2(.din(w_dff_B_yqWxRizk1_2),.dout(w_dff_B_iAoyfUpp6_2),.clk(gclk));
	jdff dff_B_71slUsZz2_2(.din(w_dff_B_iAoyfUpp6_2),.dout(w_dff_B_71slUsZz2_2),.clk(gclk));
	jdff dff_B_srbUcKaG7_2(.din(w_dff_B_71slUsZz2_2),.dout(w_dff_B_srbUcKaG7_2),.clk(gclk));
	jdff dff_B_RBHC6Fcb4_2(.din(w_dff_B_srbUcKaG7_2),.dout(w_dff_B_RBHC6Fcb4_2),.clk(gclk));
	jdff dff_B_4J1vW2Yx1_2(.din(w_dff_B_RBHC6Fcb4_2),.dout(w_dff_B_4J1vW2Yx1_2),.clk(gclk));
	jdff dff_B_9kO19CQ53_2(.din(w_dff_B_4J1vW2Yx1_2),.dout(w_dff_B_9kO19CQ53_2),.clk(gclk));
	jdff dff_B_AdGsBN6o7_2(.din(w_dff_B_9kO19CQ53_2),.dout(w_dff_B_AdGsBN6o7_2),.clk(gclk));
	jdff dff_B_A4wK2cUz5_2(.din(w_dff_B_AdGsBN6o7_2),.dout(w_dff_B_A4wK2cUz5_2),.clk(gclk));
	jdff dff_B_mY7vJ0G82_2(.din(w_dff_B_A4wK2cUz5_2),.dout(w_dff_B_mY7vJ0G82_2),.clk(gclk));
	jdff dff_B_WIL0UxPW3_2(.din(w_dff_B_mY7vJ0G82_2),.dout(w_dff_B_WIL0UxPW3_2),.clk(gclk));
	jdff dff_B_IV2gujoy4_2(.din(w_dff_B_WIL0UxPW3_2),.dout(w_dff_B_IV2gujoy4_2),.clk(gclk));
	jdff dff_B_tMXdvZbI5_2(.din(w_dff_B_IV2gujoy4_2),.dout(w_dff_B_tMXdvZbI5_2),.clk(gclk));
	jdff dff_B_nYp4JGmM8_2(.din(w_dff_B_tMXdvZbI5_2),.dout(w_dff_B_nYp4JGmM8_2),.clk(gclk));
	jdff dff_B_CHaodq9V6_2(.din(w_dff_B_nYp4JGmM8_2),.dout(w_dff_B_CHaodq9V6_2),.clk(gclk));
	jdff dff_B_yJIvjSgk6_2(.din(w_dff_B_CHaodq9V6_2),.dout(w_dff_B_yJIvjSgk6_2),.clk(gclk));
	jdff dff_B_6pcU0j1Q8_2(.din(w_dff_B_yJIvjSgk6_2),.dout(w_dff_B_6pcU0j1Q8_2),.clk(gclk));
	jdff dff_B_sMRXcpsK7_2(.din(w_dff_B_6pcU0j1Q8_2),.dout(w_dff_B_sMRXcpsK7_2),.clk(gclk));
	jdff dff_B_vtP9k1hW9_2(.din(w_dff_B_sMRXcpsK7_2),.dout(w_dff_B_vtP9k1hW9_2),.clk(gclk));
	jdff dff_B_cid6UOIn7_2(.din(w_dff_B_vtP9k1hW9_2),.dout(w_dff_B_cid6UOIn7_2),.clk(gclk));
	jdff dff_B_UeWIvyM95_2(.din(w_dff_B_cid6UOIn7_2),.dout(w_dff_B_UeWIvyM95_2),.clk(gclk));
	jdff dff_B_Y5dPiKLC6_2(.din(w_dff_B_UeWIvyM95_2),.dout(w_dff_B_Y5dPiKLC6_2),.clk(gclk));
	jdff dff_B_Ue23enFQ0_2(.din(w_dff_B_Y5dPiKLC6_2),.dout(w_dff_B_Ue23enFQ0_2),.clk(gclk));
	jdff dff_B_givJpf8v0_2(.din(w_dff_B_Ue23enFQ0_2),.dout(w_dff_B_givJpf8v0_2),.clk(gclk));
	jdff dff_B_hHa1j1AN3_2(.din(w_dff_B_givJpf8v0_2),.dout(w_dff_B_hHa1j1AN3_2),.clk(gclk));
	jdff dff_B_S5y9SNT34_2(.din(w_dff_B_hHa1j1AN3_2),.dout(w_dff_B_S5y9SNT34_2),.clk(gclk));
	jdff dff_B_y6vpjOxy1_2(.din(w_dff_B_S5y9SNT34_2),.dout(w_dff_B_y6vpjOxy1_2),.clk(gclk));
	jdff dff_B_xQciGphy7_2(.din(w_dff_B_y6vpjOxy1_2),.dout(w_dff_B_xQciGphy7_2),.clk(gclk));
	jdff dff_B_x2SPxzy90_2(.din(w_dff_B_xQciGphy7_2),.dout(w_dff_B_x2SPxzy90_2),.clk(gclk));
	jdff dff_B_cqPJn0w51_1(.din(n1039),.dout(w_dff_B_cqPJn0w51_1),.clk(gclk));
	jdff dff_B_fq1BFHsr5_2(.din(n939),.dout(w_dff_B_fq1BFHsr5_2),.clk(gclk));
	jdff dff_B_cSzjWdue0_2(.din(w_dff_B_fq1BFHsr5_2),.dout(w_dff_B_cSzjWdue0_2),.clk(gclk));
	jdff dff_B_JBEwOUys6_2(.din(w_dff_B_cSzjWdue0_2),.dout(w_dff_B_JBEwOUys6_2),.clk(gclk));
	jdff dff_B_mtfWq1CC7_2(.din(w_dff_B_JBEwOUys6_2),.dout(w_dff_B_mtfWq1CC7_2),.clk(gclk));
	jdff dff_B_JQQkmHbq4_2(.din(w_dff_B_mtfWq1CC7_2),.dout(w_dff_B_JQQkmHbq4_2),.clk(gclk));
	jdff dff_B_4wTDaToZ7_2(.din(w_dff_B_JQQkmHbq4_2),.dout(w_dff_B_4wTDaToZ7_2),.clk(gclk));
	jdff dff_B_NmSPOJLx6_2(.din(w_dff_B_4wTDaToZ7_2),.dout(w_dff_B_NmSPOJLx6_2),.clk(gclk));
	jdff dff_B_eaefrATz8_2(.din(w_dff_B_NmSPOJLx6_2),.dout(w_dff_B_eaefrATz8_2),.clk(gclk));
	jdff dff_B_mtJULdaF2_2(.din(w_dff_B_eaefrATz8_2),.dout(w_dff_B_mtJULdaF2_2),.clk(gclk));
	jdff dff_B_RiUjBtlv3_2(.din(w_dff_B_mtJULdaF2_2),.dout(w_dff_B_RiUjBtlv3_2),.clk(gclk));
	jdff dff_B_CAOi4r8W1_2(.din(w_dff_B_RiUjBtlv3_2),.dout(w_dff_B_CAOi4r8W1_2),.clk(gclk));
	jdff dff_B_osF680Ms8_2(.din(w_dff_B_CAOi4r8W1_2),.dout(w_dff_B_osF680Ms8_2),.clk(gclk));
	jdff dff_B_uqs5i3tY6_2(.din(w_dff_B_osF680Ms8_2),.dout(w_dff_B_uqs5i3tY6_2),.clk(gclk));
	jdff dff_B_y8oaetqd4_2(.din(w_dff_B_uqs5i3tY6_2),.dout(w_dff_B_y8oaetqd4_2),.clk(gclk));
	jdff dff_B_rQGcMrEs9_2(.din(w_dff_B_y8oaetqd4_2),.dout(w_dff_B_rQGcMrEs9_2),.clk(gclk));
	jdff dff_B_BRNtNuXT4_2(.din(w_dff_B_rQGcMrEs9_2),.dout(w_dff_B_BRNtNuXT4_2),.clk(gclk));
	jdff dff_B_4Sx2gh6V7_2(.din(w_dff_B_BRNtNuXT4_2),.dout(w_dff_B_4Sx2gh6V7_2),.clk(gclk));
	jdff dff_B_sBLIjZ9m4_2(.din(w_dff_B_4Sx2gh6V7_2),.dout(w_dff_B_sBLIjZ9m4_2),.clk(gclk));
	jdff dff_B_X4ong0Kj4_2(.din(w_dff_B_sBLIjZ9m4_2),.dout(w_dff_B_X4ong0Kj4_2),.clk(gclk));
	jdff dff_B_rHnL7PN81_2(.din(w_dff_B_X4ong0Kj4_2),.dout(w_dff_B_rHnL7PN81_2),.clk(gclk));
	jdff dff_B_uKCbPCPY7_2(.din(w_dff_B_rHnL7PN81_2),.dout(w_dff_B_uKCbPCPY7_2),.clk(gclk));
	jdff dff_B_S02Bfd0r7_2(.din(w_dff_B_uKCbPCPY7_2),.dout(w_dff_B_S02Bfd0r7_2),.clk(gclk));
	jdff dff_B_nP7Fmwkm2_2(.din(w_dff_B_S02Bfd0r7_2),.dout(w_dff_B_nP7Fmwkm2_2),.clk(gclk));
	jdff dff_B_dVGylOsn2_2(.din(w_dff_B_nP7Fmwkm2_2),.dout(w_dff_B_dVGylOsn2_2),.clk(gclk));
	jdff dff_B_hPuH5TjQ2_2(.din(w_dff_B_dVGylOsn2_2),.dout(w_dff_B_hPuH5TjQ2_2),.clk(gclk));
	jdff dff_B_5qNVlcW28_2(.din(w_dff_B_hPuH5TjQ2_2),.dout(w_dff_B_5qNVlcW28_2),.clk(gclk));
	jdff dff_B_1jpj3San1_2(.din(w_dff_B_5qNVlcW28_2),.dout(w_dff_B_1jpj3San1_2),.clk(gclk));
	jdff dff_B_APlCJvM38_2(.din(w_dff_B_1jpj3San1_2),.dout(w_dff_B_APlCJvM38_2),.clk(gclk));
	jdff dff_B_oHrmig9b8_1(.din(n940),.dout(w_dff_B_oHrmig9b8_1),.clk(gclk));
	jdff dff_B_rkfsy30s1_2(.din(n837),.dout(w_dff_B_rkfsy30s1_2),.clk(gclk));
	jdff dff_B_Mxo3yYls4_2(.din(w_dff_B_rkfsy30s1_2),.dout(w_dff_B_Mxo3yYls4_2),.clk(gclk));
	jdff dff_B_FqyUuTVD5_2(.din(w_dff_B_Mxo3yYls4_2),.dout(w_dff_B_FqyUuTVD5_2),.clk(gclk));
	jdff dff_B_SMxuUzVq0_2(.din(w_dff_B_FqyUuTVD5_2),.dout(w_dff_B_SMxuUzVq0_2),.clk(gclk));
	jdff dff_B_5dsBJsfb2_2(.din(w_dff_B_SMxuUzVq0_2),.dout(w_dff_B_5dsBJsfb2_2),.clk(gclk));
	jdff dff_B_Ty9VgCsB4_2(.din(w_dff_B_5dsBJsfb2_2),.dout(w_dff_B_Ty9VgCsB4_2),.clk(gclk));
	jdff dff_B_F2dQohVp4_2(.din(w_dff_B_Ty9VgCsB4_2),.dout(w_dff_B_F2dQohVp4_2),.clk(gclk));
	jdff dff_B_DradSCFZ6_2(.din(w_dff_B_F2dQohVp4_2),.dout(w_dff_B_DradSCFZ6_2),.clk(gclk));
	jdff dff_B_jMoggx2e1_2(.din(w_dff_B_DradSCFZ6_2),.dout(w_dff_B_jMoggx2e1_2),.clk(gclk));
	jdff dff_B_BUhoAFux1_2(.din(w_dff_B_jMoggx2e1_2),.dout(w_dff_B_BUhoAFux1_2),.clk(gclk));
	jdff dff_B_m0OZvkKe2_2(.din(w_dff_B_BUhoAFux1_2),.dout(w_dff_B_m0OZvkKe2_2),.clk(gclk));
	jdff dff_B_4t4LIWnU8_2(.din(w_dff_B_m0OZvkKe2_2),.dout(w_dff_B_4t4LIWnU8_2),.clk(gclk));
	jdff dff_B_48IWPnwM2_2(.din(w_dff_B_4t4LIWnU8_2),.dout(w_dff_B_48IWPnwM2_2),.clk(gclk));
	jdff dff_B_LSjNWVPQ1_2(.din(w_dff_B_48IWPnwM2_2),.dout(w_dff_B_LSjNWVPQ1_2),.clk(gclk));
	jdff dff_B_fu1ZQUaY3_2(.din(w_dff_B_LSjNWVPQ1_2),.dout(w_dff_B_fu1ZQUaY3_2),.clk(gclk));
	jdff dff_B_yJfrJwUh2_2(.din(w_dff_B_fu1ZQUaY3_2),.dout(w_dff_B_yJfrJwUh2_2),.clk(gclk));
	jdff dff_B_75uPTHOI5_2(.din(w_dff_B_yJfrJwUh2_2),.dout(w_dff_B_75uPTHOI5_2),.clk(gclk));
	jdff dff_B_oZ2MO2l11_2(.din(w_dff_B_75uPTHOI5_2),.dout(w_dff_B_oZ2MO2l11_2),.clk(gclk));
	jdff dff_B_hfvKoMDr7_2(.din(w_dff_B_oZ2MO2l11_2),.dout(w_dff_B_hfvKoMDr7_2),.clk(gclk));
	jdff dff_B_wyR6zR8Z8_2(.din(w_dff_B_hfvKoMDr7_2),.dout(w_dff_B_wyR6zR8Z8_2),.clk(gclk));
	jdff dff_B_u2l2OQMG6_2(.din(w_dff_B_wyR6zR8Z8_2),.dout(w_dff_B_u2l2OQMG6_2),.clk(gclk));
	jdff dff_B_BpOj8OnA6_2(.din(w_dff_B_u2l2OQMG6_2),.dout(w_dff_B_BpOj8OnA6_2),.clk(gclk));
	jdff dff_B_RaYknB3l7_2(.din(w_dff_B_BpOj8OnA6_2),.dout(w_dff_B_RaYknB3l7_2),.clk(gclk));
	jdff dff_B_SunJ3O1y4_2(.din(w_dff_B_RaYknB3l7_2),.dout(w_dff_B_SunJ3O1y4_2),.clk(gclk));
	jdff dff_B_UyzY5MlU4_2(.din(w_dff_B_SunJ3O1y4_2),.dout(w_dff_B_UyzY5MlU4_2),.clk(gclk));
	jdff dff_B_Ev4CQdpk0_1(.din(n838),.dout(w_dff_B_Ev4CQdpk0_1),.clk(gclk));
	jdff dff_B_0pM1aYEb6_2(.din(n739),.dout(w_dff_B_0pM1aYEb6_2),.clk(gclk));
	jdff dff_B_3GWtVEYO3_2(.din(w_dff_B_0pM1aYEb6_2),.dout(w_dff_B_3GWtVEYO3_2),.clk(gclk));
	jdff dff_B_IX4X35ka6_2(.din(w_dff_B_3GWtVEYO3_2),.dout(w_dff_B_IX4X35ka6_2),.clk(gclk));
	jdff dff_B_DVDEdXfi1_2(.din(w_dff_B_IX4X35ka6_2),.dout(w_dff_B_DVDEdXfi1_2),.clk(gclk));
	jdff dff_B_kebgbYYS2_2(.din(w_dff_B_DVDEdXfi1_2),.dout(w_dff_B_kebgbYYS2_2),.clk(gclk));
	jdff dff_B_s0jgHSUe3_2(.din(w_dff_B_kebgbYYS2_2),.dout(w_dff_B_s0jgHSUe3_2),.clk(gclk));
	jdff dff_B_5M9CLjh65_2(.din(w_dff_B_s0jgHSUe3_2),.dout(w_dff_B_5M9CLjh65_2),.clk(gclk));
	jdff dff_B_Uas4CeUS6_2(.din(w_dff_B_5M9CLjh65_2),.dout(w_dff_B_Uas4CeUS6_2),.clk(gclk));
	jdff dff_B_Znvr1vFd2_2(.din(w_dff_B_Uas4CeUS6_2),.dout(w_dff_B_Znvr1vFd2_2),.clk(gclk));
	jdff dff_B_eKXQWiGV8_2(.din(w_dff_B_Znvr1vFd2_2),.dout(w_dff_B_eKXQWiGV8_2),.clk(gclk));
	jdff dff_B_NsFZQH9p6_2(.din(w_dff_B_eKXQWiGV8_2),.dout(w_dff_B_NsFZQH9p6_2),.clk(gclk));
	jdff dff_B_6E1N0qgj9_2(.din(w_dff_B_NsFZQH9p6_2),.dout(w_dff_B_6E1N0qgj9_2),.clk(gclk));
	jdff dff_B_ctiY2GBW2_2(.din(w_dff_B_6E1N0qgj9_2),.dout(w_dff_B_ctiY2GBW2_2),.clk(gclk));
	jdff dff_B_FSOn4wq39_2(.din(w_dff_B_ctiY2GBW2_2),.dout(w_dff_B_FSOn4wq39_2),.clk(gclk));
	jdff dff_B_03w5wrtF0_2(.din(w_dff_B_FSOn4wq39_2),.dout(w_dff_B_03w5wrtF0_2),.clk(gclk));
	jdff dff_B_BXDoiOag6_2(.din(w_dff_B_03w5wrtF0_2),.dout(w_dff_B_BXDoiOag6_2),.clk(gclk));
	jdff dff_B_KujAZ5lW0_2(.din(w_dff_B_BXDoiOag6_2),.dout(w_dff_B_KujAZ5lW0_2),.clk(gclk));
	jdff dff_B_SCiVOBJu5_2(.din(w_dff_B_KujAZ5lW0_2),.dout(w_dff_B_SCiVOBJu5_2),.clk(gclk));
	jdff dff_B_CjUmJcZb7_2(.din(w_dff_B_SCiVOBJu5_2),.dout(w_dff_B_CjUmJcZb7_2),.clk(gclk));
	jdff dff_B_dozsRspm0_2(.din(w_dff_B_CjUmJcZb7_2),.dout(w_dff_B_dozsRspm0_2),.clk(gclk));
	jdff dff_B_FD27LYtI0_2(.din(w_dff_B_dozsRspm0_2),.dout(w_dff_B_FD27LYtI0_2),.clk(gclk));
	jdff dff_B_DgxOZg6R1_2(.din(w_dff_B_FD27LYtI0_2),.dout(w_dff_B_DgxOZg6R1_2),.clk(gclk));
	jdff dff_B_uh9KG59w7_1(.din(n740),.dout(w_dff_B_uh9KG59w7_1),.clk(gclk));
	jdff dff_B_khBAQAxY9_2(.din(n647),.dout(w_dff_B_khBAQAxY9_2),.clk(gclk));
	jdff dff_B_1a3P04YC0_2(.din(w_dff_B_khBAQAxY9_2),.dout(w_dff_B_1a3P04YC0_2),.clk(gclk));
	jdff dff_B_1eVCw3IS4_2(.din(w_dff_B_1a3P04YC0_2),.dout(w_dff_B_1eVCw3IS4_2),.clk(gclk));
	jdff dff_B_cXspYIdS7_2(.din(w_dff_B_1eVCw3IS4_2),.dout(w_dff_B_cXspYIdS7_2),.clk(gclk));
	jdff dff_B_yOndADZW7_2(.din(w_dff_B_cXspYIdS7_2),.dout(w_dff_B_yOndADZW7_2),.clk(gclk));
	jdff dff_B_aId95FVP0_2(.din(w_dff_B_yOndADZW7_2),.dout(w_dff_B_aId95FVP0_2),.clk(gclk));
	jdff dff_B_Zp74O74J9_2(.din(w_dff_B_aId95FVP0_2),.dout(w_dff_B_Zp74O74J9_2),.clk(gclk));
	jdff dff_B_R2N939fv4_2(.din(w_dff_B_Zp74O74J9_2),.dout(w_dff_B_R2N939fv4_2),.clk(gclk));
	jdff dff_B_m0DtOOQ88_2(.din(w_dff_B_R2N939fv4_2),.dout(w_dff_B_m0DtOOQ88_2),.clk(gclk));
	jdff dff_B_OKb7n73E7_2(.din(w_dff_B_m0DtOOQ88_2),.dout(w_dff_B_OKb7n73E7_2),.clk(gclk));
	jdff dff_B_Knb5uX1Z5_2(.din(w_dff_B_OKb7n73E7_2),.dout(w_dff_B_Knb5uX1Z5_2),.clk(gclk));
	jdff dff_B_KGi53uo27_2(.din(w_dff_B_Knb5uX1Z5_2),.dout(w_dff_B_KGi53uo27_2),.clk(gclk));
	jdff dff_B_hziZrZsd5_2(.din(w_dff_B_KGi53uo27_2),.dout(w_dff_B_hziZrZsd5_2),.clk(gclk));
	jdff dff_B_bIXaZiWu4_2(.din(w_dff_B_hziZrZsd5_2),.dout(w_dff_B_bIXaZiWu4_2),.clk(gclk));
	jdff dff_B_qscKhjSK6_2(.din(w_dff_B_bIXaZiWu4_2),.dout(w_dff_B_qscKhjSK6_2),.clk(gclk));
	jdff dff_B_1grgBQC35_2(.din(w_dff_B_qscKhjSK6_2),.dout(w_dff_B_1grgBQC35_2),.clk(gclk));
	jdff dff_B_mkGiDRUD8_2(.din(w_dff_B_1grgBQC35_2),.dout(w_dff_B_mkGiDRUD8_2),.clk(gclk));
	jdff dff_B_wVmiFhGN1_2(.din(w_dff_B_mkGiDRUD8_2),.dout(w_dff_B_wVmiFhGN1_2),.clk(gclk));
	jdff dff_B_cbKJmi6f7_2(.din(w_dff_B_wVmiFhGN1_2),.dout(w_dff_B_cbKJmi6f7_2),.clk(gclk));
	jdff dff_B_bPimEsZa9_1(.din(n648),.dout(w_dff_B_bPimEsZa9_1),.clk(gclk));
	jdff dff_B_rWJETwad5_2(.din(n562),.dout(w_dff_B_rWJETwad5_2),.clk(gclk));
	jdff dff_B_RnOIm7mA1_2(.din(w_dff_B_rWJETwad5_2),.dout(w_dff_B_RnOIm7mA1_2),.clk(gclk));
	jdff dff_B_2XDlsdfZ8_2(.din(w_dff_B_RnOIm7mA1_2),.dout(w_dff_B_2XDlsdfZ8_2),.clk(gclk));
	jdff dff_B_7hHJbMH16_2(.din(w_dff_B_2XDlsdfZ8_2),.dout(w_dff_B_7hHJbMH16_2),.clk(gclk));
	jdff dff_B_YL4rz5Oc4_2(.din(w_dff_B_7hHJbMH16_2),.dout(w_dff_B_YL4rz5Oc4_2),.clk(gclk));
	jdff dff_B_BBAL9Mm45_2(.din(w_dff_B_YL4rz5Oc4_2),.dout(w_dff_B_BBAL9Mm45_2),.clk(gclk));
	jdff dff_B_4W6g83Ap5_2(.din(w_dff_B_BBAL9Mm45_2),.dout(w_dff_B_4W6g83Ap5_2),.clk(gclk));
	jdff dff_B_kbnzJNs73_2(.din(w_dff_B_4W6g83Ap5_2),.dout(w_dff_B_kbnzJNs73_2),.clk(gclk));
	jdff dff_B_uiGck9g12_2(.din(w_dff_B_kbnzJNs73_2),.dout(w_dff_B_uiGck9g12_2),.clk(gclk));
	jdff dff_B_w9vMPKL08_2(.din(w_dff_B_uiGck9g12_2),.dout(w_dff_B_w9vMPKL08_2),.clk(gclk));
	jdff dff_B_NSeJwMri3_2(.din(w_dff_B_w9vMPKL08_2),.dout(w_dff_B_NSeJwMri3_2),.clk(gclk));
	jdff dff_B_TcPTESMx8_2(.din(w_dff_B_NSeJwMri3_2),.dout(w_dff_B_TcPTESMx8_2),.clk(gclk));
	jdff dff_B_T8WafdQk1_2(.din(w_dff_B_TcPTESMx8_2),.dout(w_dff_B_T8WafdQk1_2),.clk(gclk));
	jdff dff_B_8LVRvV5P4_2(.din(w_dff_B_T8WafdQk1_2),.dout(w_dff_B_8LVRvV5P4_2),.clk(gclk));
	jdff dff_B_USbybAmP6_2(.din(w_dff_B_8LVRvV5P4_2),.dout(w_dff_B_USbybAmP6_2),.clk(gclk));
	jdff dff_B_NAIXv9WN7_2(.din(w_dff_B_USbybAmP6_2),.dout(w_dff_B_NAIXv9WN7_2),.clk(gclk));
	jdff dff_B_Op82aIIH5_1(.din(n563),.dout(w_dff_B_Op82aIIH5_1),.clk(gclk));
	jdff dff_B_5fzhd01t4_2(.din(n484),.dout(w_dff_B_5fzhd01t4_2),.clk(gclk));
	jdff dff_B_Q1EulNwY6_2(.din(w_dff_B_5fzhd01t4_2),.dout(w_dff_B_Q1EulNwY6_2),.clk(gclk));
	jdff dff_B_AECID8ag8_2(.din(w_dff_B_Q1EulNwY6_2),.dout(w_dff_B_AECID8ag8_2),.clk(gclk));
	jdff dff_B_Chug2rJ45_2(.din(w_dff_B_AECID8ag8_2),.dout(w_dff_B_Chug2rJ45_2),.clk(gclk));
	jdff dff_B_ZAKizlQK3_2(.din(w_dff_B_Chug2rJ45_2),.dout(w_dff_B_ZAKizlQK3_2),.clk(gclk));
	jdff dff_B_K433J3Fj6_2(.din(w_dff_B_ZAKizlQK3_2),.dout(w_dff_B_K433J3Fj6_2),.clk(gclk));
	jdff dff_B_iZsWPgul7_2(.din(w_dff_B_K433J3Fj6_2),.dout(w_dff_B_iZsWPgul7_2),.clk(gclk));
	jdff dff_B_fjdZW6g19_2(.din(w_dff_B_iZsWPgul7_2),.dout(w_dff_B_fjdZW6g19_2),.clk(gclk));
	jdff dff_B_enosXykL2_2(.din(w_dff_B_fjdZW6g19_2),.dout(w_dff_B_enosXykL2_2),.clk(gclk));
	jdff dff_B_sZrhq1Gf8_2(.din(w_dff_B_enosXykL2_2),.dout(w_dff_B_sZrhq1Gf8_2),.clk(gclk));
	jdff dff_B_z31PjNrX4_2(.din(w_dff_B_sZrhq1Gf8_2),.dout(w_dff_B_z31PjNrX4_2),.clk(gclk));
	jdff dff_B_ipLRqzef3_2(.din(w_dff_B_z31PjNrX4_2),.dout(w_dff_B_ipLRqzef3_2),.clk(gclk));
	jdff dff_B_hnVkheOv4_2(.din(w_dff_B_ipLRqzef3_2),.dout(w_dff_B_hnVkheOv4_2),.clk(gclk));
	jdff dff_B_vOu5VeOi2_1(.din(n485),.dout(w_dff_B_vOu5VeOi2_1),.clk(gclk));
	jdff dff_B_l59LYDJ84_2(.din(n413),.dout(w_dff_B_l59LYDJ84_2),.clk(gclk));
	jdff dff_B_y8rb9ITS0_2(.din(w_dff_B_l59LYDJ84_2),.dout(w_dff_B_y8rb9ITS0_2),.clk(gclk));
	jdff dff_B_SqeNrBCI9_2(.din(w_dff_B_y8rb9ITS0_2),.dout(w_dff_B_SqeNrBCI9_2),.clk(gclk));
	jdff dff_B_uOME5WZa9_2(.din(w_dff_B_SqeNrBCI9_2),.dout(w_dff_B_uOME5WZa9_2),.clk(gclk));
	jdff dff_B_582O5wJe8_2(.din(w_dff_B_uOME5WZa9_2),.dout(w_dff_B_582O5wJe8_2),.clk(gclk));
	jdff dff_B_9T145DRs4_2(.din(w_dff_B_582O5wJe8_2),.dout(w_dff_B_9T145DRs4_2),.clk(gclk));
	jdff dff_B_0O3cDWAy8_2(.din(w_dff_B_9T145DRs4_2),.dout(w_dff_B_0O3cDWAy8_2),.clk(gclk));
	jdff dff_B_m4MiRyCc2_2(.din(w_dff_B_0O3cDWAy8_2),.dout(w_dff_B_m4MiRyCc2_2),.clk(gclk));
	jdff dff_B_dH3500ym3_2(.din(w_dff_B_m4MiRyCc2_2),.dout(w_dff_B_dH3500ym3_2),.clk(gclk));
	jdff dff_B_jOYZKkVE5_2(.din(w_dff_B_dH3500ym3_2),.dout(w_dff_B_jOYZKkVE5_2),.clk(gclk));
	jdff dff_B_WbZgNx2W0_2(.din(n416),.dout(w_dff_B_WbZgNx2W0_2),.clk(gclk));
	jdff dff_B_HLZqCbhz3_1(.din(n414),.dout(w_dff_B_HLZqCbhz3_1),.clk(gclk));
	jdff dff_B_vdT1MCRY4_2(.din(n350),.dout(w_dff_B_vdT1MCRY4_2),.clk(gclk));
	jdff dff_B_n0IvnRvw2_2(.din(w_dff_B_vdT1MCRY4_2),.dout(w_dff_B_n0IvnRvw2_2),.clk(gclk));
	jdff dff_B_UhWQDQaU0_2(.din(w_dff_B_n0IvnRvw2_2),.dout(w_dff_B_UhWQDQaU0_2),.clk(gclk));
	jdff dff_B_cHuZeCJF9_2(.din(w_dff_B_UhWQDQaU0_2),.dout(w_dff_B_cHuZeCJF9_2),.clk(gclk));
	jdff dff_B_JiTexVVI6_2(.din(w_dff_B_cHuZeCJF9_2),.dout(w_dff_B_JiTexVVI6_2),.clk(gclk));
	jdff dff_B_pKLuxngU2_2(.din(w_dff_B_JiTexVVI6_2),.dout(w_dff_B_pKLuxngU2_2),.clk(gclk));
	jdff dff_B_v1WaF1H94_2(.din(n364),.dout(w_dff_B_v1WaF1H94_2),.clk(gclk));
	jdff dff_B_equHhrx92_2(.din(n295),.dout(w_dff_B_equHhrx92_2),.clk(gclk));
	jdff dff_B_mP9gkpxo4_2(.din(w_dff_B_equHhrx92_2),.dout(w_dff_B_mP9gkpxo4_2),.clk(gclk));
	jdff dff_B_xGVVmCvC2_2(.din(w_dff_B_mP9gkpxo4_2),.dout(w_dff_B_xGVVmCvC2_2),.clk(gclk));
	jdff dff_B_Nlus2vSY4_0(.din(n300),.dout(w_dff_B_Nlus2vSY4_0),.clk(gclk));
	jdff dff_A_UtJmcRHB7_0(.dout(w_n243_0[0]),.din(w_dff_A_UtJmcRHB7_0),.clk(gclk));
	jdff dff_A_wPraWFFy9_0(.dout(w_dff_A_UtJmcRHB7_0),.din(w_dff_A_wPraWFFy9_0),.clk(gclk));
	jdff dff_A_6eIcQALi3_1(.dout(w_n243_0[1]),.din(w_dff_A_6eIcQALi3_1),.clk(gclk));
	jdff dff_A_VyoFlOGM9_1(.dout(w_dff_A_6eIcQALi3_1),.din(w_dff_A_VyoFlOGM9_1),.clk(gclk));
	jdff dff_B_Jk58wg5I9_1(.din(n1532),.dout(w_dff_B_Jk58wg5I9_1),.clk(gclk));
	jdff dff_B_VswOaHDp8_2(.din(n1466),.dout(w_dff_B_VswOaHDp8_2),.clk(gclk));
	jdff dff_B_gyQuQIR00_2(.din(w_dff_B_VswOaHDp8_2),.dout(w_dff_B_gyQuQIR00_2),.clk(gclk));
	jdff dff_B_PWuIdnru6_2(.din(w_dff_B_gyQuQIR00_2),.dout(w_dff_B_PWuIdnru6_2),.clk(gclk));
	jdff dff_B_rrAS1YKE4_2(.din(w_dff_B_PWuIdnru6_2),.dout(w_dff_B_rrAS1YKE4_2),.clk(gclk));
	jdff dff_B_jDGzIUPu7_2(.din(w_dff_B_rrAS1YKE4_2),.dout(w_dff_B_jDGzIUPu7_2),.clk(gclk));
	jdff dff_B_qAueXGVO4_2(.din(w_dff_B_jDGzIUPu7_2),.dout(w_dff_B_qAueXGVO4_2),.clk(gclk));
	jdff dff_B_1wm2OyUI1_2(.din(w_dff_B_qAueXGVO4_2),.dout(w_dff_B_1wm2OyUI1_2),.clk(gclk));
	jdff dff_B_otHU9EIX4_2(.din(w_dff_B_1wm2OyUI1_2),.dout(w_dff_B_otHU9EIX4_2),.clk(gclk));
	jdff dff_B_i0R3tGtH7_2(.din(w_dff_B_otHU9EIX4_2),.dout(w_dff_B_i0R3tGtH7_2),.clk(gclk));
	jdff dff_B_ysPxCx4m1_2(.din(w_dff_B_i0R3tGtH7_2),.dout(w_dff_B_ysPxCx4m1_2),.clk(gclk));
	jdff dff_B_JHLSWOjB5_2(.din(w_dff_B_ysPxCx4m1_2),.dout(w_dff_B_JHLSWOjB5_2),.clk(gclk));
	jdff dff_B_GHJNnxQR7_2(.din(w_dff_B_JHLSWOjB5_2),.dout(w_dff_B_GHJNnxQR7_2),.clk(gclk));
	jdff dff_B_Jb9rvoFV0_2(.din(w_dff_B_GHJNnxQR7_2),.dout(w_dff_B_Jb9rvoFV0_2),.clk(gclk));
	jdff dff_B_wYKYUiNB6_2(.din(w_dff_B_Jb9rvoFV0_2),.dout(w_dff_B_wYKYUiNB6_2),.clk(gclk));
	jdff dff_B_ijcB46EL8_2(.din(w_dff_B_wYKYUiNB6_2),.dout(w_dff_B_ijcB46EL8_2),.clk(gclk));
	jdff dff_B_94t7fViY5_2(.din(w_dff_B_ijcB46EL8_2),.dout(w_dff_B_94t7fViY5_2),.clk(gclk));
	jdff dff_B_jtTjHHDr1_2(.din(w_dff_B_94t7fViY5_2),.dout(w_dff_B_jtTjHHDr1_2),.clk(gclk));
	jdff dff_B_fjn5SRUZ0_2(.din(w_dff_B_jtTjHHDr1_2),.dout(w_dff_B_fjn5SRUZ0_2),.clk(gclk));
	jdff dff_B_WSmMpNTo0_2(.din(w_dff_B_fjn5SRUZ0_2),.dout(w_dff_B_WSmMpNTo0_2),.clk(gclk));
	jdff dff_B_9siyY3d93_2(.din(w_dff_B_WSmMpNTo0_2),.dout(w_dff_B_9siyY3d93_2),.clk(gclk));
	jdff dff_B_B2PypJQY7_2(.din(w_dff_B_9siyY3d93_2),.dout(w_dff_B_B2PypJQY7_2),.clk(gclk));
	jdff dff_B_3CmrlFIu6_2(.din(w_dff_B_B2PypJQY7_2),.dout(w_dff_B_3CmrlFIu6_2),.clk(gclk));
	jdff dff_B_fcglWAlY8_2(.din(w_dff_B_3CmrlFIu6_2),.dout(w_dff_B_fcglWAlY8_2),.clk(gclk));
	jdff dff_B_aWnC45ll6_2(.din(w_dff_B_fcglWAlY8_2),.dout(w_dff_B_aWnC45ll6_2),.clk(gclk));
	jdff dff_B_KUFfFuAc8_2(.din(w_dff_B_aWnC45ll6_2),.dout(w_dff_B_KUFfFuAc8_2),.clk(gclk));
	jdff dff_B_Mqyjql5n2_2(.din(w_dff_B_KUFfFuAc8_2),.dout(w_dff_B_Mqyjql5n2_2),.clk(gclk));
	jdff dff_B_MEQp75cg1_2(.din(w_dff_B_Mqyjql5n2_2),.dout(w_dff_B_MEQp75cg1_2),.clk(gclk));
	jdff dff_B_5ligMp879_2(.din(w_dff_B_MEQp75cg1_2),.dout(w_dff_B_5ligMp879_2),.clk(gclk));
	jdff dff_B_mnZcbAnD2_2(.din(w_dff_B_5ligMp879_2),.dout(w_dff_B_mnZcbAnD2_2),.clk(gclk));
	jdff dff_B_roI7RvcF0_2(.din(w_dff_B_mnZcbAnD2_2),.dout(w_dff_B_roI7RvcF0_2),.clk(gclk));
	jdff dff_B_SFQP6Lyz8_2(.din(w_dff_B_roI7RvcF0_2),.dout(w_dff_B_SFQP6Lyz8_2),.clk(gclk));
	jdff dff_B_4Ba7yUbC7_2(.din(w_dff_B_SFQP6Lyz8_2),.dout(w_dff_B_4Ba7yUbC7_2),.clk(gclk));
	jdff dff_B_gdbDDKO17_2(.din(w_dff_B_4Ba7yUbC7_2),.dout(w_dff_B_gdbDDKO17_2),.clk(gclk));
	jdff dff_B_xDY6n8gT4_2(.din(w_dff_B_gdbDDKO17_2),.dout(w_dff_B_xDY6n8gT4_2),.clk(gclk));
	jdff dff_B_kAAMWXrC9_2(.din(w_dff_B_xDY6n8gT4_2),.dout(w_dff_B_kAAMWXrC9_2),.clk(gclk));
	jdff dff_B_fe0Sx0cY3_2(.din(w_dff_B_kAAMWXrC9_2),.dout(w_dff_B_fe0Sx0cY3_2),.clk(gclk));
	jdff dff_B_vVmjT4eL4_2(.din(w_dff_B_fe0Sx0cY3_2),.dout(w_dff_B_vVmjT4eL4_2),.clk(gclk));
	jdff dff_B_UgcHleqv1_2(.din(w_dff_B_vVmjT4eL4_2),.dout(w_dff_B_UgcHleqv1_2),.clk(gclk));
	jdff dff_B_4yxHmEsr7_2(.din(w_dff_B_UgcHleqv1_2),.dout(w_dff_B_4yxHmEsr7_2),.clk(gclk));
	jdff dff_B_MO9xv4sd5_2(.din(w_dff_B_4yxHmEsr7_2),.dout(w_dff_B_MO9xv4sd5_2),.clk(gclk));
	jdff dff_B_FdfsJ2bu9_2(.din(w_dff_B_MO9xv4sd5_2),.dout(w_dff_B_FdfsJ2bu9_2),.clk(gclk));
	jdff dff_B_KJgi9yBS9_2(.din(w_dff_B_FdfsJ2bu9_2),.dout(w_dff_B_KJgi9yBS9_2),.clk(gclk));
	jdff dff_B_MmSVDjU50_2(.din(w_dff_B_KJgi9yBS9_2),.dout(w_dff_B_MmSVDjU50_2),.clk(gclk));
	jdff dff_B_M7PjRRpN6_2(.din(w_dff_B_MmSVDjU50_2),.dout(w_dff_B_M7PjRRpN6_2),.clk(gclk));
	jdff dff_B_2x6iD6hl6_2(.din(w_dff_B_M7PjRRpN6_2),.dout(w_dff_B_2x6iD6hl6_2),.clk(gclk));
	jdff dff_B_p3ZNSoEw1_2(.din(w_dff_B_2x6iD6hl6_2),.dout(w_dff_B_p3ZNSoEw1_2),.clk(gclk));
	jdff dff_B_1ax3ECta3_0(.din(n1531),.dout(w_dff_B_1ax3ECta3_0),.clk(gclk));
	jdff dff_A_PxH1NRvU1_1(.dout(w_n1519_0[1]),.din(w_dff_A_PxH1NRvU1_1),.clk(gclk));
	jdff dff_B_1aMAG6Sh9_1(.din(n1467),.dout(w_dff_B_1aMAG6Sh9_1),.clk(gclk));
	jdff dff_B_inRuTdfA4_2(.din(n1395),.dout(w_dff_B_inRuTdfA4_2),.clk(gclk));
	jdff dff_B_AlyN7p6I0_2(.din(w_dff_B_inRuTdfA4_2),.dout(w_dff_B_AlyN7p6I0_2),.clk(gclk));
	jdff dff_B_zAGxqyxT5_2(.din(w_dff_B_AlyN7p6I0_2),.dout(w_dff_B_zAGxqyxT5_2),.clk(gclk));
	jdff dff_B_wFlugMFi4_2(.din(w_dff_B_zAGxqyxT5_2),.dout(w_dff_B_wFlugMFi4_2),.clk(gclk));
	jdff dff_B_TxlXRj5I9_2(.din(w_dff_B_wFlugMFi4_2),.dout(w_dff_B_TxlXRj5I9_2),.clk(gclk));
	jdff dff_B_icdHhhTo6_2(.din(w_dff_B_TxlXRj5I9_2),.dout(w_dff_B_icdHhhTo6_2),.clk(gclk));
	jdff dff_B_xi53Znlx0_2(.din(w_dff_B_icdHhhTo6_2),.dout(w_dff_B_xi53Znlx0_2),.clk(gclk));
	jdff dff_B_f7way87Z8_2(.din(w_dff_B_xi53Znlx0_2),.dout(w_dff_B_f7way87Z8_2),.clk(gclk));
	jdff dff_B_WbFIrWsJ2_2(.din(w_dff_B_f7way87Z8_2),.dout(w_dff_B_WbFIrWsJ2_2),.clk(gclk));
	jdff dff_B_A8ztJC4t9_2(.din(w_dff_B_WbFIrWsJ2_2),.dout(w_dff_B_A8ztJC4t9_2),.clk(gclk));
	jdff dff_B_OyhKT9HT2_2(.din(w_dff_B_A8ztJC4t9_2),.dout(w_dff_B_OyhKT9HT2_2),.clk(gclk));
	jdff dff_B_MGtDrr1s5_2(.din(w_dff_B_OyhKT9HT2_2),.dout(w_dff_B_MGtDrr1s5_2),.clk(gclk));
	jdff dff_B_3YmYvg2T6_2(.din(w_dff_B_MGtDrr1s5_2),.dout(w_dff_B_3YmYvg2T6_2),.clk(gclk));
	jdff dff_B_fbiqLisC1_2(.din(w_dff_B_3YmYvg2T6_2),.dout(w_dff_B_fbiqLisC1_2),.clk(gclk));
	jdff dff_B_6uFlHUwT1_2(.din(w_dff_B_fbiqLisC1_2),.dout(w_dff_B_6uFlHUwT1_2),.clk(gclk));
	jdff dff_B_fwn4TuNY9_2(.din(w_dff_B_6uFlHUwT1_2),.dout(w_dff_B_fwn4TuNY9_2),.clk(gclk));
	jdff dff_B_d3Nai7tk8_2(.din(w_dff_B_fwn4TuNY9_2),.dout(w_dff_B_d3Nai7tk8_2),.clk(gclk));
	jdff dff_B_UJVtCxeN7_2(.din(w_dff_B_d3Nai7tk8_2),.dout(w_dff_B_UJVtCxeN7_2),.clk(gclk));
	jdff dff_B_FcJZjd6i2_2(.din(w_dff_B_UJVtCxeN7_2),.dout(w_dff_B_FcJZjd6i2_2),.clk(gclk));
	jdff dff_B_nMCAX8wY4_2(.din(w_dff_B_FcJZjd6i2_2),.dout(w_dff_B_nMCAX8wY4_2),.clk(gclk));
	jdff dff_B_tAKjTtwH1_2(.din(w_dff_B_nMCAX8wY4_2),.dout(w_dff_B_tAKjTtwH1_2),.clk(gclk));
	jdff dff_B_oAtIciFs5_2(.din(w_dff_B_tAKjTtwH1_2),.dout(w_dff_B_oAtIciFs5_2),.clk(gclk));
	jdff dff_B_mmY24BI05_2(.din(w_dff_B_oAtIciFs5_2),.dout(w_dff_B_mmY24BI05_2),.clk(gclk));
	jdff dff_B_GzKuMRKi2_2(.din(w_dff_B_mmY24BI05_2),.dout(w_dff_B_GzKuMRKi2_2),.clk(gclk));
	jdff dff_B_X82b9LiP9_2(.din(w_dff_B_GzKuMRKi2_2),.dout(w_dff_B_X82b9LiP9_2),.clk(gclk));
	jdff dff_B_7bkMfmwt4_2(.din(w_dff_B_X82b9LiP9_2),.dout(w_dff_B_7bkMfmwt4_2),.clk(gclk));
	jdff dff_B_qnyTeGld3_2(.din(w_dff_B_7bkMfmwt4_2),.dout(w_dff_B_qnyTeGld3_2),.clk(gclk));
	jdff dff_B_qGC9KhU82_2(.din(w_dff_B_qnyTeGld3_2),.dout(w_dff_B_qGC9KhU82_2),.clk(gclk));
	jdff dff_B_ZvnobH0V6_2(.din(w_dff_B_qGC9KhU82_2),.dout(w_dff_B_ZvnobH0V6_2),.clk(gclk));
	jdff dff_B_zZ9onDR59_2(.din(w_dff_B_ZvnobH0V6_2),.dout(w_dff_B_zZ9onDR59_2),.clk(gclk));
	jdff dff_B_2Elc3VTP4_2(.din(w_dff_B_zZ9onDR59_2),.dout(w_dff_B_2Elc3VTP4_2),.clk(gclk));
	jdff dff_B_xTZTmmn96_2(.din(w_dff_B_2Elc3VTP4_2),.dout(w_dff_B_xTZTmmn96_2),.clk(gclk));
	jdff dff_B_v4KQNg9H3_2(.din(w_dff_B_xTZTmmn96_2),.dout(w_dff_B_v4KQNg9H3_2),.clk(gclk));
	jdff dff_B_315ukMqs3_2(.din(w_dff_B_v4KQNg9H3_2),.dout(w_dff_B_315ukMqs3_2),.clk(gclk));
	jdff dff_B_I3NbLvJY0_2(.din(w_dff_B_315ukMqs3_2),.dout(w_dff_B_I3NbLvJY0_2),.clk(gclk));
	jdff dff_B_5QTuLfKd5_2(.din(w_dff_B_I3NbLvJY0_2),.dout(w_dff_B_5QTuLfKd5_2),.clk(gclk));
	jdff dff_B_r9hSc30U2_2(.din(w_dff_B_5QTuLfKd5_2),.dout(w_dff_B_r9hSc30U2_2),.clk(gclk));
	jdff dff_B_y4IGddwb1_2(.din(w_dff_B_r9hSc30U2_2),.dout(w_dff_B_y4IGddwb1_2),.clk(gclk));
	jdff dff_B_ElXZYIa20_2(.din(w_dff_B_y4IGddwb1_2),.dout(w_dff_B_ElXZYIa20_2),.clk(gclk));
	jdff dff_B_M3LK1xzU2_2(.din(w_dff_B_ElXZYIa20_2),.dout(w_dff_B_M3LK1xzU2_2),.clk(gclk));
	jdff dff_B_IbvucGwe3_2(.din(w_dff_B_M3LK1xzU2_2),.dout(w_dff_B_IbvucGwe3_2),.clk(gclk));
	jdff dff_B_9qHtF55P1_2(.din(n1448),.dout(w_dff_B_9qHtF55P1_2),.clk(gclk));
	jdff dff_B_lZcZVzdw3_1(.din(n1396),.dout(w_dff_B_lZcZVzdw3_1),.clk(gclk));
	jdff dff_B_XPhmulcQ5_2(.din(n1317),.dout(w_dff_B_XPhmulcQ5_2),.clk(gclk));
	jdff dff_B_ODZG99Yp7_2(.din(w_dff_B_XPhmulcQ5_2),.dout(w_dff_B_ODZG99Yp7_2),.clk(gclk));
	jdff dff_B_bf3OVSsi8_2(.din(w_dff_B_ODZG99Yp7_2),.dout(w_dff_B_bf3OVSsi8_2),.clk(gclk));
	jdff dff_B_iqTgUew23_2(.din(w_dff_B_bf3OVSsi8_2),.dout(w_dff_B_iqTgUew23_2),.clk(gclk));
	jdff dff_B_m4v3d7Kv1_2(.din(w_dff_B_iqTgUew23_2),.dout(w_dff_B_m4v3d7Kv1_2),.clk(gclk));
	jdff dff_B_neuP4lQ52_2(.din(w_dff_B_m4v3d7Kv1_2),.dout(w_dff_B_neuP4lQ52_2),.clk(gclk));
	jdff dff_B_TSUrgaKt8_2(.din(w_dff_B_neuP4lQ52_2),.dout(w_dff_B_TSUrgaKt8_2),.clk(gclk));
	jdff dff_B_wD8Zr9vW6_2(.din(w_dff_B_TSUrgaKt8_2),.dout(w_dff_B_wD8Zr9vW6_2),.clk(gclk));
	jdff dff_B_7Yfwf9aZ7_2(.din(w_dff_B_wD8Zr9vW6_2),.dout(w_dff_B_7Yfwf9aZ7_2),.clk(gclk));
	jdff dff_B_RsgfZ2uu3_2(.din(w_dff_B_7Yfwf9aZ7_2),.dout(w_dff_B_RsgfZ2uu3_2),.clk(gclk));
	jdff dff_B_K1KFsQ2u2_2(.din(w_dff_B_RsgfZ2uu3_2),.dout(w_dff_B_K1KFsQ2u2_2),.clk(gclk));
	jdff dff_B_i2KxM8Re5_2(.din(w_dff_B_K1KFsQ2u2_2),.dout(w_dff_B_i2KxM8Re5_2),.clk(gclk));
	jdff dff_B_OlTIx4ce8_2(.din(w_dff_B_i2KxM8Re5_2),.dout(w_dff_B_OlTIx4ce8_2),.clk(gclk));
	jdff dff_B_mlj6Hy8p2_2(.din(w_dff_B_OlTIx4ce8_2),.dout(w_dff_B_mlj6Hy8p2_2),.clk(gclk));
	jdff dff_B_OgCIYfPB8_2(.din(w_dff_B_mlj6Hy8p2_2),.dout(w_dff_B_OgCIYfPB8_2),.clk(gclk));
	jdff dff_B_SnhMdyTp7_2(.din(w_dff_B_OgCIYfPB8_2),.dout(w_dff_B_SnhMdyTp7_2),.clk(gclk));
	jdff dff_B_cwGQd2xI4_2(.din(w_dff_B_SnhMdyTp7_2),.dout(w_dff_B_cwGQd2xI4_2),.clk(gclk));
	jdff dff_B_A9IIPvHv3_2(.din(w_dff_B_cwGQd2xI4_2),.dout(w_dff_B_A9IIPvHv3_2),.clk(gclk));
	jdff dff_B_4kjnqb1K6_2(.din(w_dff_B_A9IIPvHv3_2),.dout(w_dff_B_4kjnqb1K6_2),.clk(gclk));
	jdff dff_B_YZT9ddvX4_2(.din(w_dff_B_4kjnqb1K6_2),.dout(w_dff_B_YZT9ddvX4_2),.clk(gclk));
	jdff dff_B_JwZKP0fX2_2(.din(w_dff_B_YZT9ddvX4_2),.dout(w_dff_B_JwZKP0fX2_2),.clk(gclk));
	jdff dff_B_1CIVLKIj4_2(.din(w_dff_B_JwZKP0fX2_2),.dout(w_dff_B_1CIVLKIj4_2),.clk(gclk));
	jdff dff_B_Ld4rCjnd4_2(.din(w_dff_B_1CIVLKIj4_2),.dout(w_dff_B_Ld4rCjnd4_2),.clk(gclk));
	jdff dff_B_kRSEWkmn0_2(.din(w_dff_B_Ld4rCjnd4_2),.dout(w_dff_B_kRSEWkmn0_2),.clk(gclk));
	jdff dff_B_pepnupah9_2(.din(w_dff_B_kRSEWkmn0_2),.dout(w_dff_B_pepnupah9_2),.clk(gclk));
	jdff dff_B_FOHMAXDs5_2(.din(w_dff_B_pepnupah9_2),.dout(w_dff_B_FOHMAXDs5_2),.clk(gclk));
	jdff dff_B_Z74a6RK19_2(.din(w_dff_B_FOHMAXDs5_2),.dout(w_dff_B_Z74a6RK19_2),.clk(gclk));
	jdff dff_B_J5YehL8a8_2(.din(w_dff_B_Z74a6RK19_2),.dout(w_dff_B_J5YehL8a8_2),.clk(gclk));
	jdff dff_B_yUuoIbTx8_2(.din(w_dff_B_J5YehL8a8_2),.dout(w_dff_B_yUuoIbTx8_2),.clk(gclk));
	jdff dff_B_EvBpFlVv7_2(.din(w_dff_B_yUuoIbTx8_2),.dout(w_dff_B_EvBpFlVv7_2),.clk(gclk));
	jdff dff_B_JP0xAU0r3_2(.din(w_dff_B_EvBpFlVv7_2),.dout(w_dff_B_JP0xAU0r3_2),.clk(gclk));
	jdff dff_B_3FVv3jQY6_2(.din(w_dff_B_JP0xAU0r3_2),.dout(w_dff_B_3FVv3jQY6_2),.clk(gclk));
	jdff dff_B_pExHhlD19_2(.din(w_dff_B_3FVv3jQY6_2),.dout(w_dff_B_pExHhlD19_2),.clk(gclk));
	jdff dff_B_YVSvoF7J7_2(.din(w_dff_B_pExHhlD19_2),.dout(w_dff_B_YVSvoF7J7_2),.clk(gclk));
	jdff dff_B_WQ1WoQPh9_2(.din(w_dff_B_YVSvoF7J7_2),.dout(w_dff_B_WQ1WoQPh9_2),.clk(gclk));
	jdff dff_B_0fI18B7O1_2(.din(w_dff_B_WQ1WoQPh9_2),.dout(w_dff_B_0fI18B7O1_2),.clk(gclk));
	jdff dff_B_GKDcWaz37_2(.din(w_dff_B_0fI18B7O1_2),.dout(w_dff_B_GKDcWaz37_2),.clk(gclk));
	jdff dff_B_Rp3ucYYc1_2(.din(w_dff_B_GKDcWaz37_2),.dout(w_dff_B_Rp3ucYYc1_2),.clk(gclk));
	jdff dff_B_MCd6ORrO0_2(.din(n1370),.dout(w_dff_B_MCd6ORrO0_2),.clk(gclk));
	jdff dff_B_htxOHOD62_1(.din(n1318),.dout(w_dff_B_htxOHOD62_1),.clk(gclk));
	jdff dff_B_1kv8LCsj3_2(.din(n1232),.dout(w_dff_B_1kv8LCsj3_2),.clk(gclk));
	jdff dff_B_JcQK66OL1_2(.din(w_dff_B_1kv8LCsj3_2),.dout(w_dff_B_JcQK66OL1_2),.clk(gclk));
	jdff dff_B_uaUhpf4s7_2(.din(w_dff_B_JcQK66OL1_2),.dout(w_dff_B_uaUhpf4s7_2),.clk(gclk));
	jdff dff_B_G47l6X8V8_2(.din(w_dff_B_uaUhpf4s7_2),.dout(w_dff_B_G47l6X8V8_2),.clk(gclk));
	jdff dff_B_Ro9KydpO7_2(.din(w_dff_B_G47l6X8V8_2),.dout(w_dff_B_Ro9KydpO7_2),.clk(gclk));
	jdff dff_B_9SuPu77z6_2(.din(w_dff_B_Ro9KydpO7_2),.dout(w_dff_B_9SuPu77z6_2),.clk(gclk));
	jdff dff_B_WrNEXcKN9_2(.din(w_dff_B_9SuPu77z6_2),.dout(w_dff_B_WrNEXcKN9_2),.clk(gclk));
	jdff dff_B_43XMRe7j9_2(.din(w_dff_B_WrNEXcKN9_2),.dout(w_dff_B_43XMRe7j9_2),.clk(gclk));
	jdff dff_B_s2cgr2AW3_2(.din(w_dff_B_43XMRe7j9_2),.dout(w_dff_B_s2cgr2AW3_2),.clk(gclk));
	jdff dff_B_Ozkoba9W8_2(.din(w_dff_B_s2cgr2AW3_2),.dout(w_dff_B_Ozkoba9W8_2),.clk(gclk));
	jdff dff_B_yXxqEg2W1_2(.din(w_dff_B_Ozkoba9W8_2),.dout(w_dff_B_yXxqEg2W1_2),.clk(gclk));
	jdff dff_B_OAtSuQRO1_2(.din(w_dff_B_yXxqEg2W1_2),.dout(w_dff_B_OAtSuQRO1_2),.clk(gclk));
	jdff dff_B_mcp0dSs15_2(.din(w_dff_B_OAtSuQRO1_2),.dout(w_dff_B_mcp0dSs15_2),.clk(gclk));
	jdff dff_B_6A6qlhvf4_2(.din(w_dff_B_mcp0dSs15_2),.dout(w_dff_B_6A6qlhvf4_2),.clk(gclk));
	jdff dff_B_TnKfDes99_2(.din(w_dff_B_6A6qlhvf4_2),.dout(w_dff_B_TnKfDes99_2),.clk(gclk));
	jdff dff_B_cKDrpWUJ7_2(.din(w_dff_B_TnKfDes99_2),.dout(w_dff_B_cKDrpWUJ7_2),.clk(gclk));
	jdff dff_B_vrDEH52I1_2(.din(w_dff_B_cKDrpWUJ7_2),.dout(w_dff_B_vrDEH52I1_2),.clk(gclk));
	jdff dff_B_0xICeWWk8_2(.din(w_dff_B_vrDEH52I1_2),.dout(w_dff_B_0xICeWWk8_2),.clk(gclk));
	jdff dff_B_2q53ClOO1_2(.din(w_dff_B_0xICeWWk8_2),.dout(w_dff_B_2q53ClOO1_2),.clk(gclk));
	jdff dff_B_Yk0RwQoZ2_2(.din(w_dff_B_2q53ClOO1_2),.dout(w_dff_B_Yk0RwQoZ2_2),.clk(gclk));
	jdff dff_B_7HWmukWz4_2(.din(w_dff_B_Yk0RwQoZ2_2),.dout(w_dff_B_7HWmukWz4_2),.clk(gclk));
	jdff dff_B_vskxeJnm5_2(.din(w_dff_B_7HWmukWz4_2),.dout(w_dff_B_vskxeJnm5_2),.clk(gclk));
	jdff dff_B_GliYpxA19_2(.din(w_dff_B_vskxeJnm5_2),.dout(w_dff_B_GliYpxA19_2),.clk(gclk));
	jdff dff_B_ZcvSGS8T6_2(.din(w_dff_B_GliYpxA19_2),.dout(w_dff_B_ZcvSGS8T6_2),.clk(gclk));
	jdff dff_B_mzHnQgh06_2(.din(w_dff_B_ZcvSGS8T6_2),.dout(w_dff_B_mzHnQgh06_2),.clk(gclk));
	jdff dff_B_iFYc1Zr22_2(.din(w_dff_B_mzHnQgh06_2),.dout(w_dff_B_iFYc1Zr22_2),.clk(gclk));
	jdff dff_B_lFIs85bo3_2(.din(w_dff_B_iFYc1Zr22_2),.dout(w_dff_B_lFIs85bo3_2),.clk(gclk));
	jdff dff_B_vRhkfnEJ5_2(.din(w_dff_B_lFIs85bo3_2),.dout(w_dff_B_vRhkfnEJ5_2),.clk(gclk));
	jdff dff_B_wle64HD04_2(.din(w_dff_B_vRhkfnEJ5_2),.dout(w_dff_B_wle64HD04_2),.clk(gclk));
	jdff dff_B_LybolC2y0_2(.din(w_dff_B_wle64HD04_2),.dout(w_dff_B_LybolC2y0_2),.clk(gclk));
	jdff dff_B_Efvx2P9U3_2(.din(w_dff_B_LybolC2y0_2),.dout(w_dff_B_Efvx2P9U3_2),.clk(gclk));
	jdff dff_B_7J8XEpEw9_2(.din(w_dff_B_Efvx2P9U3_2),.dout(w_dff_B_7J8XEpEw9_2),.clk(gclk));
	jdff dff_B_cl5b4eIb2_2(.din(w_dff_B_7J8XEpEw9_2),.dout(w_dff_B_cl5b4eIb2_2),.clk(gclk));
	jdff dff_B_UnKdesTB9_2(.din(w_dff_B_cl5b4eIb2_2),.dout(w_dff_B_UnKdesTB9_2),.clk(gclk));
	jdff dff_B_PCF5qNEU6_2(.din(w_dff_B_UnKdesTB9_2),.dout(w_dff_B_PCF5qNEU6_2),.clk(gclk));
	jdff dff_B_JVkXs9h96_2(.din(n1285),.dout(w_dff_B_JVkXs9h96_2),.clk(gclk));
	jdff dff_B_rlehoPlh3_1(.din(n1233),.dout(w_dff_B_rlehoPlh3_1),.clk(gclk));
	jdff dff_B_qnRqOOAO4_2(.din(n1141),.dout(w_dff_B_qnRqOOAO4_2),.clk(gclk));
	jdff dff_B_ZqoxD9Vg7_2(.din(w_dff_B_qnRqOOAO4_2),.dout(w_dff_B_ZqoxD9Vg7_2),.clk(gclk));
	jdff dff_B_xDle3Ej36_2(.din(w_dff_B_ZqoxD9Vg7_2),.dout(w_dff_B_xDle3Ej36_2),.clk(gclk));
	jdff dff_B_AKAHyaMk5_2(.din(w_dff_B_xDle3Ej36_2),.dout(w_dff_B_AKAHyaMk5_2),.clk(gclk));
	jdff dff_B_2mk9SXaj9_2(.din(w_dff_B_AKAHyaMk5_2),.dout(w_dff_B_2mk9SXaj9_2),.clk(gclk));
	jdff dff_B_Oa14ZuAL2_2(.din(w_dff_B_2mk9SXaj9_2),.dout(w_dff_B_Oa14ZuAL2_2),.clk(gclk));
	jdff dff_B_r7CK5K8f0_2(.din(w_dff_B_Oa14ZuAL2_2),.dout(w_dff_B_r7CK5K8f0_2),.clk(gclk));
	jdff dff_B_TP682LfF3_2(.din(w_dff_B_r7CK5K8f0_2),.dout(w_dff_B_TP682LfF3_2),.clk(gclk));
	jdff dff_B_t5S7MITs9_2(.din(w_dff_B_TP682LfF3_2),.dout(w_dff_B_t5S7MITs9_2),.clk(gclk));
	jdff dff_B_8nU81K8n7_2(.din(w_dff_B_t5S7MITs9_2),.dout(w_dff_B_8nU81K8n7_2),.clk(gclk));
	jdff dff_B_T3GpPOQY2_2(.din(w_dff_B_8nU81K8n7_2),.dout(w_dff_B_T3GpPOQY2_2),.clk(gclk));
	jdff dff_B_eF3Gpsp35_2(.din(w_dff_B_T3GpPOQY2_2),.dout(w_dff_B_eF3Gpsp35_2),.clk(gclk));
	jdff dff_B_ddrW5dNN3_2(.din(w_dff_B_eF3Gpsp35_2),.dout(w_dff_B_ddrW5dNN3_2),.clk(gclk));
	jdff dff_B_w4xr85qT5_2(.din(w_dff_B_ddrW5dNN3_2),.dout(w_dff_B_w4xr85qT5_2),.clk(gclk));
	jdff dff_B_8pU5VBtd7_2(.din(w_dff_B_w4xr85qT5_2),.dout(w_dff_B_8pU5VBtd7_2),.clk(gclk));
	jdff dff_B_GH8vwDxA0_2(.din(w_dff_B_8pU5VBtd7_2),.dout(w_dff_B_GH8vwDxA0_2),.clk(gclk));
	jdff dff_B_eKVAcyeV2_2(.din(w_dff_B_GH8vwDxA0_2),.dout(w_dff_B_eKVAcyeV2_2),.clk(gclk));
	jdff dff_B_mB3RxjI36_2(.din(w_dff_B_eKVAcyeV2_2),.dout(w_dff_B_mB3RxjI36_2),.clk(gclk));
	jdff dff_B_CkRzwcqN2_2(.din(w_dff_B_mB3RxjI36_2),.dout(w_dff_B_CkRzwcqN2_2),.clk(gclk));
	jdff dff_B_Pbp7yQOZ7_2(.din(w_dff_B_CkRzwcqN2_2),.dout(w_dff_B_Pbp7yQOZ7_2),.clk(gclk));
	jdff dff_B_NyT20UKI5_2(.din(w_dff_B_Pbp7yQOZ7_2),.dout(w_dff_B_NyT20UKI5_2),.clk(gclk));
	jdff dff_B_3gwCqjJ39_2(.din(w_dff_B_NyT20UKI5_2),.dout(w_dff_B_3gwCqjJ39_2),.clk(gclk));
	jdff dff_B_glm0SnPP8_2(.din(w_dff_B_3gwCqjJ39_2),.dout(w_dff_B_glm0SnPP8_2),.clk(gclk));
	jdff dff_B_pti3UzU40_2(.din(w_dff_B_glm0SnPP8_2),.dout(w_dff_B_pti3UzU40_2),.clk(gclk));
	jdff dff_B_FoFBl5Dz0_2(.din(w_dff_B_pti3UzU40_2),.dout(w_dff_B_FoFBl5Dz0_2),.clk(gclk));
	jdff dff_B_yWvJUjzJ6_2(.din(w_dff_B_FoFBl5Dz0_2),.dout(w_dff_B_yWvJUjzJ6_2),.clk(gclk));
	jdff dff_B_SZlvdsNo7_2(.din(w_dff_B_yWvJUjzJ6_2),.dout(w_dff_B_SZlvdsNo7_2),.clk(gclk));
	jdff dff_B_oDJxQXXZ3_2(.din(w_dff_B_SZlvdsNo7_2),.dout(w_dff_B_oDJxQXXZ3_2),.clk(gclk));
	jdff dff_B_2lamB7ID9_2(.din(w_dff_B_oDJxQXXZ3_2),.dout(w_dff_B_2lamB7ID9_2),.clk(gclk));
	jdff dff_B_aggaVBfl3_2(.din(w_dff_B_2lamB7ID9_2),.dout(w_dff_B_aggaVBfl3_2),.clk(gclk));
	jdff dff_B_0vKqDatN5_2(.din(w_dff_B_aggaVBfl3_2),.dout(w_dff_B_0vKqDatN5_2),.clk(gclk));
	jdff dff_B_kuIpC0Vp4_2(.din(w_dff_B_0vKqDatN5_2),.dout(w_dff_B_kuIpC0Vp4_2),.clk(gclk));
	jdff dff_B_D3YZD5D76_2(.din(n1194),.dout(w_dff_B_D3YZD5D76_2),.clk(gclk));
	jdff dff_B_gg2FB3My6_1(.din(n1142),.dout(w_dff_B_gg2FB3My6_1),.clk(gclk));
	jdff dff_B_AnYtJzmb0_2(.din(n1043),.dout(w_dff_B_AnYtJzmb0_2),.clk(gclk));
	jdff dff_B_CnCUs4fP3_2(.din(w_dff_B_AnYtJzmb0_2),.dout(w_dff_B_CnCUs4fP3_2),.clk(gclk));
	jdff dff_B_OE7PKV5v8_2(.din(w_dff_B_CnCUs4fP3_2),.dout(w_dff_B_OE7PKV5v8_2),.clk(gclk));
	jdff dff_B_boDm4h6Q6_2(.din(w_dff_B_OE7PKV5v8_2),.dout(w_dff_B_boDm4h6Q6_2),.clk(gclk));
	jdff dff_B_Cu9evJKv3_2(.din(w_dff_B_boDm4h6Q6_2),.dout(w_dff_B_Cu9evJKv3_2),.clk(gclk));
	jdff dff_B_KAXUlKk72_2(.din(w_dff_B_Cu9evJKv3_2),.dout(w_dff_B_KAXUlKk72_2),.clk(gclk));
	jdff dff_B_SSStPbcG2_2(.din(w_dff_B_KAXUlKk72_2),.dout(w_dff_B_SSStPbcG2_2),.clk(gclk));
	jdff dff_B_H4pIjNWc0_2(.din(w_dff_B_SSStPbcG2_2),.dout(w_dff_B_H4pIjNWc0_2),.clk(gclk));
	jdff dff_B_qtWiRgLX7_2(.din(w_dff_B_H4pIjNWc0_2),.dout(w_dff_B_qtWiRgLX7_2),.clk(gclk));
	jdff dff_B_tpxzfHba9_2(.din(w_dff_B_qtWiRgLX7_2),.dout(w_dff_B_tpxzfHba9_2),.clk(gclk));
	jdff dff_B_LAEe8wqC0_2(.din(w_dff_B_tpxzfHba9_2),.dout(w_dff_B_LAEe8wqC0_2),.clk(gclk));
	jdff dff_B_330shDWv3_2(.din(w_dff_B_LAEe8wqC0_2),.dout(w_dff_B_330shDWv3_2),.clk(gclk));
	jdff dff_B_9DurIZci1_2(.din(w_dff_B_330shDWv3_2),.dout(w_dff_B_9DurIZci1_2),.clk(gclk));
	jdff dff_B_BvuxMaUr8_2(.din(w_dff_B_9DurIZci1_2),.dout(w_dff_B_BvuxMaUr8_2),.clk(gclk));
	jdff dff_B_UrosZfpO2_2(.din(w_dff_B_BvuxMaUr8_2),.dout(w_dff_B_UrosZfpO2_2),.clk(gclk));
	jdff dff_B_UKZvIUwg3_2(.din(w_dff_B_UrosZfpO2_2),.dout(w_dff_B_UKZvIUwg3_2),.clk(gclk));
	jdff dff_B_wJxyiGT27_2(.din(w_dff_B_UKZvIUwg3_2),.dout(w_dff_B_wJxyiGT27_2),.clk(gclk));
	jdff dff_B_5BjBczeA7_2(.din(w_dff_B_wJxyiGT27_2),.dout(w_dff_B_5BjBczeA7_2),.clk(gclk));
	jdff dff_B_5CNKYy1E9_2(.din(w_dff_B_5BjBczeA7_2),.dout(w_dff_B_5CNKYy1E9_2),.clk(gclk));
	jdff dff_B_8b3QJ5jh9_2(.din(w_dff_B_5CNKYy1E9_2),.dout(w_dff_B_8b3QJ5jh9_2),.clk(gclk));
	jdff dff_B_QckKYNf06_2(.din(w_dff_B_8b3QJ5jh9_2),.dout(w_dff_B_QckKYNf06_2),.clk(gclk));
	jdff dff_B_cwz65iGh5_2(.din(w_dff_B_QckKYNf06_2),.dout(w_dff_B_cwz65iGh5_2),.clk(gclk));
	jdff dff_B_wY0IsHG82_2(.din(w_dff_B_cwz65iGh5_2),.dout(w_dff_B_wY0IsHG82_2),.clk(gclk));
	jdff dff_B_klWKGcQv2_2(.din(w_dff_B_wY0IsHG82_2),.dout(w_dff_B_klWKGcQv2_2),.clk(gclk));
	jdff dff_B_3IaUNx172_2(.din(w_dff_B_klWKGcQv2_2),.dout(w_dff_B_3IaUNx172_2),.clk(gclk));
	jdff dff_B_lEHS7Zak6_2(.din(w_dff_B_3IaUNx172_2),.dout(w_dff_B_lEHS7Zak6_2),.clk(gclk));
	jdff dff_B_K6D321cK1_2(.din(w_dff_B_lEHS7Zak6_2),.dout(w_dff_B_K6D321cK1_2),.clk(gclk));
	jdff dff_B_tYEhZjTJ3_2(.din(w_dff_B_K6D321cK1_2),.dout(w_dff_B_tYEhZjTJ3_2),.clk(gclk));
	jdff dff_B_0et19v5d5_2(.din(w_dff_B_tYEhZjTJ3_2),.dout(w_dff_B_0et19v5d5_2),.clk(gclk));
	jdff dff_B_SmpoGJ4N8_2(.din(n1095),.dout(w_dff_B_SmpoGJ4N8_2),.clk(gclk));
	jdff dff_B_7bnw41xC0_1(.din(n1044),.dout(w_dff_B_7bnw41xC0_1),.clk(gclk));
	jdff dff_B_p5YvcBGO7_2(.din(n944),.dout(w_dff_B_p5YvcBGO7_2),.clk(gclk));
	jdff dff_B_wSOusyKg6_2(.din(w_dff_B_p5YvcBGO7_2),.dout(w_dff_B_wSOusyKg6_2),.clk(gclk));
	jdff dff_B_3vt0DaiS8_2(.din(w_dff_B_wSOusyKg6_2),.dout(w_dff_B_3vt0DaiS8_2),.clk(gclk));
	jdff dff_B_wEcy0GZO6_2(.din(w_dff_B_3vt0DaiS8_2),.dout(w_dff_B_wEcy0GZO6_2),.clk(gclk));
	jdff dff_B_z4G4z7R83_2(.din(w_dff_B_wEcy0GZO6_2),.dout(w_dff_B_z4G4z7R83_2),.clk(gclk));
	jdff dff_B_uUr8EfHm2_2(.din(w_dff_B_z4G4z7R83_2),.dout(w_dff_B_uUr8EfHm2_2),.clk(gclk));
	jdff dff_B_TbXRX6eS1_2(.din(w_dff_B_uUr8EfHm2_2),.dout(w_dff_B_TbXRX6eS1_2),.clk(gclk));
	jdff dff_B_YmavrFzT1_2(.din(w_dff_B_TbXRX6eS1_2),.dout(w_dff_B_YmavrFzT1_2),.clk(gclk));
	jdff dff_B_4bn01ozy2_2(.din(w_dff_B_YmavrFzT1_2),.dout(w_dff_B_4bn01ozy2_2),.clk(gclk));
	jdff dff_B_Ge5Cc4Kl6_2(.din(w_dff_B_4bn01ozy2_2),.dout(w_dff_B_Ge5Cc4Kl6_2),.clk(gclk));
	jdff dff_B_PimQafJy6_2(.din(w_dff_B_Ge5Cc4Kl6_2),.dout(w_dff_B_PimQafJy6_2),.clk(gclk));
	jdff dff_B_ZEMII0Zt4_2(.din(w_dff_B_PimQafJy6_2),.dout(w_dff_B_ZEMII0Zt4_2),.clk(gclk));
	jdff dff_B_DWDa9spu8_2(.din(w_dff_B_ZEMII0Zt4_2),.dout(w_dff_B_DWDa9spu8_2),.clk(gclk));
	jdff dff_B_voH1uFbB5_2(.din(w_dff_B_DWDa9spu8_2),.dout(w_dff_B_voH1uFbB5_2),.clk(gclk));
	jdff dff_B_d1tQvrDw6_2(.din(w_dff_B_voH1uFbB5_2),.dout(w_dff_B_d1tQvrDw6_2),.clk(gclk));
	jdff dff_B_R0ygIqUD6_2(.din(w_dff_B_d1tQvrDw6_2),.dout(w_dff_B_R0ygIqUD6_2),.clk(gclk));
	jdff dff_B_U1dqrdTD5_2(.din(w_dff_B_R0ygIqUD6_2),.dout(w_dff_B_U1dqrdTD5_2),.clk(gclk));
	jdff dff_B_CKkttcAN6_2(.din(w_dff_B_U1dqrdTD5_2),.dout(w_dff_B_CKkttcAN6_2),.clk(gclk));
	jdff dff_B_KGLorfy53_2(.din(w_dff_B_CKkttcAN6_2),.dout(w_dff_B_KGLorfy53_2),.clk(gclk));
	jdff dff_B_RBtOME0j2_2(.din(w_dff_B_KGLorfy53_2),.dout(w_dff_B_RBtOME0j2_2),.clk(gclk));
	jdff dff_B_TL7zEP7a7_2(.din(w_dff_B_RBtOME0j2_2),.dout(w_dff_B_TL7zEP7a7_2),.clk(gclk));
	jdff dff_B_pzJHSiQL5_2(.din(w_dff_B_TL7zEP7a7_2),.dout(w_dff_B_pzJHSiQL5_2),.clk(gclk));
	jdff dff_B_gWArFEau1_2(.din(w_dff_B_pzJHSiQL5_2),.dout(w_dff_B_gWArFEau1_2),.clk(gclk));
	jdff dff_B_QtAs6B3W4_2(.din(w_dff_B_gWArFEau1_2),.dout(w_dff_B_QtAs6B3W4_2),.clk(gclk));
	jdff dff_B_PGbTllZq5_2(.din(w_dff_B_QtAs6B3W4_2),.dout(w_dff_B_PGbTllZq5_2),.clk(gclk));
	jdff dff_B_ZaSiZtFw1_2(.din(w_dff_B_PGbTllZq5_2),.dout(w_dff_B_ZaSiZtFw1_2),.clk(gclk));
	jdff dff_B_hYJzon4O3_2(.din(n996),.dout(w_dff_B_hYJzon4O3_2),.clk(gclk));
	jdff dff_B_OnoqUXsn8_1(.din(n945),.dout(w_dff_B_OnoqUXsn8_1),.clk(gclk));
	jdff dff_B_KefcasIe6_2(.din(n842),.dout(w_dff_B_KefcasIe6_2),.clk(gclk));
	jdff dff_B_HzG04r9G3_2(.din(w_dff_B_KefcasIe6_2),.dout(w_dff_B_HzG04r9G3_2),.clk(gclk));
	jdff dff_B_fHjGnlhj5_2(.din(w_dff_B_HzG04r9G3_2),.dout(w_dff_B_fHjGnlhj5_2),.clk(gclk));
	jdff dff_B_s6yqWXg95_2(.din(w_dff_B_fHjGnlhj5_2),.dout(w_dff_B_s6yqWXg95_2),.clk(gclk));
	jdff dff_B_n1zXIAZP7_2(.din(w_dff_B_s6yqWXg95_2),.dout(w_dff_B_n1zXIAZP7_2),.clk(gclk));
	jdff dff_B_yV6xjVtf5_2(.din(w_dff_B_n1zXIAZP7_2),.dout(w_dff_B_yV6xjVtf5_2),.clk(gclk));
	jdff dff_B_B7lOt4jv7_2(.din(w_dff_B_yV6xjVtf5_2),.dout(w_dff_B_B7lOt4jv7_2),.clk(gclk));
	jdff dff_B_htayxL4J3_2(.din(w_dff_B_B7lOt4jv7_2),.dout(w_dff_B_htayxL4J3_2),.clk(gclk));
	jdff dff_B_UpNnZp7M1_2(.din(w_dff_B_htayxL4J3_2),.dout(w_dff_B_UpNnZp7M1_2),.clk(gclk));
	jdff dff_B_hRxavixN3_2(.din(w_dff_B_UpNnZp7M1_2),.dout(w_dff_B_hRxavixN3_2),.clk(gclk));
	jdff dff_B_8VSF4nkX0_2(.din(w_dff_B_hRxavixN3_2),.dout(w_dff_B_8VSF4nkX0_2),.clk(gclk));
	jdff dff_B_Y3A3szwY8_2(.din(w_dff_B_8VSF4nkX0_2),.dout(w_dff_B_Y3A3szwY8_2),.clk(gclk));
	jdff dff_B_NRvHbfiu7_2(.din(w_dff_B_Y3A3szwY8_2),.dout(w_dff_B_NRvHbfiu7_2),.clk(gclk));
	jdff dff_B_Yp43ncj11_2(.din(w_dff_B_NRvHbfiu7_2),.dout(w_dff_B_Yp43ncj11_2),.clk(gclk));
	jdff dff_B_mOXjGl9Q4_2(.din(w_dff_B_Yp43ncj11_2),.dout(w_dff_B_mOXjGl9Q4_2),.clk(gclk));
	jdff dff_B_Ik7mrRdj5_2(.din(w_dff_B_mOXjGl9Q4_2),.dout(w_dff_B_Ik7mrRdj5_2),.clk(gclk));
	jdff dff_B_yO9TkDke5_2(.din(w_dff_B_Ik7mrRdj5_2),.dout(w_dff_B_yO9TkDke5_2),.clk(gclk));
	jdff dff_B_MvEKXKAS1_2(.din(w_dff_B_yO9TkDke5_2),.dout(w_dff_B_MvEKXKAS1_2),.clk(gclk));
	jdff dff_B_gYJCljrR4_2(.din(w_dff_B_MvEKXKAS1_2),.dout(w_dff_B_gYJCljrR4_2),.clk(gclk));
	jdff dff_B_za8iUesw8_2(.din(w_dff_B_gYJCljrR4_2),.dout(w_dff_B_za8iUesw8_2),.clk(gclk));
	jdff dff_B_u2NwlTMH0_2(.din(w_dff_B_za8iUesw8_2),.dout(w_dff_B_u2NwlTMH0_2),.clk(gclk));
	jdff dff_B_6Ah8I60j5_2(.din(w_dff_B_u2NwlTMH0_2),.dout(w_dff_B_6Ah8I60j5_2),.clk(gclk));
	jdff dff_B_cKWKrVXj8_2(.din(w_dff_B_6Ah8I60j5_2),.dout(w_dff_B_cKWKrVXj8_2),.clk(gclk));
	jdff dff_B_V85fjSlv9_2(.din(n890),.dout(w_dff_B_V85fjSlv9_2),.clk(gclk));
	jdff dff_B_rB1nKRZA0_1(.din(n843),.dout(w_dff_B_rB1nKRZA0_1),.clk(gclk));
	jdff dff_B_B7KRyNZu6_2(.din(n744),.dout(w_dff_B_B7KRyNZu6_2),.clk(gclk));
	jdff dff_B_HMuKd9D11_2(.din(w_dff_B_B7KRyNZu6_2),.dout(w_dff_B_HMuKd9D11_2),.clk(gclk));
	jdff dff_B_miT1FUoR1_2(.din(w_dff_B_HMuKd9D11_2),.dout(w_dff_B_miT1FUoR1_2),.clk(gclk));
	jdff dff_B_yMvNDoDM5_2(.din(w_dff_B_miT1FUoR1_2),.dout(w_dff_B_yMvNDoDM5_2),.clk(gclk));
	jdff dff_B_sbJNVXe81_2(.din(w_dff_B_yMvNDoDM5_2),.dout(w_dff_B_sbJNVXe81_2),.clk(gclk));
	jdff dff_B_eI9W4oGE3_2(.din(w_dff_B_sbJNVXe81_2),.dout(w_dff_B_eI9W4oGE3_2),.clk(gclk));
	jdff dff_B_B8ee8iVP2_2(.din(w_dff_B_eI9W4oGE3_2),.dout(w_dff_B_B8ee8iVP2_2),.clk(gclk));
	jdff dff_B_PevLuJYF7_2(.din(w_dff_B_B8ee8iVP2_2),.dout(w_dff_B_PevLuJYF7_2),.clk(gclk));
	jdff dff_B_5w3Av6GE3_2(.din(w_dff_B_PevLuJYF7_2),.dout(w_dff_B_5w3Av6GE3_2),.clk(gclk));
	jdff dff_B_p0PG2wGQ8_2(.din(w_dff_B_5w3Av6GE3_2),.dout(w_dff_B_p0PG2wGQ8_2),.clk(gclk));
	jdff dff_B_M8nokPFC0_2(.din(w_dff_B_p0PG2wGQ8_2),.dout(w_dff_B_M8nokPFC0_2),.clk(gclk));
	jdff dff_B_WZnKADMq0_2(.din(w_dff_B_M8nokPFC0_2),.dout(w_dff_B_WZnKADMq0_2),.clk(gclk));
	jdff dff_B_AZvMrFNO5_2(.din(w_dff_B_WZnKADMq0_2),.dout(w_dff_B_AZvMrFNO5_2),.clk(gclk));
	jdff dff_B_xy8eEO6j9_2(.din(w_dff_B_AZvMrFNO5_2),.dout(w_dff_B_xy8eEO6j9_2),.clk(gclk));
	jdff dff_B_bMmjzMxZ7_2(.din(w_dff_B_xy8eEO6j9_2),.dout(w_dff_B_bMmjzMxZ7_2),.clk(gclk));
	jdff dff_B_OerqAZ2r4_2(.din(w_dff_B_bMmjzMxZ7_2),.dout(w_dff_B_OerqAZ2r4_2),.clk(gclk));
	jdff dff_B_jPKYSNFo1_2(.din(w_dff_B_OerqAZ2r4_2),.dout(w_dff_B_jPKYSNFo1_2),.clk(gclk));
	jdff dff_B_388w2Zga0_2(.din(w_dff_B_jPKYSNFo1_2),.dout(w_dff_B_388w2Zga0_2),.clk(gclk));
	jdff dff_B_kpIfSQFC1_2(.din(w_dff_B_388w2Zga0_2),.dout(w_dff_B_kpIfSQFC1_2),.clk(gclk));
	jdff dff_B_VA0c2Vd83_2(.din(w_dff_B_kpIfSQFC1_2),.dout(w_dff_B_VA0c2Vd83_2),.clk(gclk));
	jdff dff_B_iedO2Yhv8_2(.din(n787),.dout(w_dff_B_iedO2Yhv8_2),.clk(gclk));
	jdff dff_B_SLuxqxfn3_1(.din(n745),.dout(w_dff_B_SLuxqxfn3_1),.clk(gclk));
	jdff dff_B_3TAhVC4f7_2(.din(n652),.dout(w_dff_B_3TAhVC4f7_2),.clk(gclk));
	jdff dff_B_w3Yl70fm8_2(.din(w_dff_B_3TAhVC4f7_2),.dout(w_dff_B_w3Yl70fm8_2),.clk(gclk));
	jdff dff_B_L8n5hhGj3_2(.din(w_dff_B_w3Yl70fm8_2),.dout(w_dff_B_L8n5hhGj3_2),.clk(gclk));
	jdff dff_B_huCo1aGm2_2(.din(w_dff_B_L8n5hhGj3_2),.dout(w_dff_B_huCo1aGm2_2),.clk(gclk));
	jdff dff_B_eoxFidYA3_2(.din(w_dff_B_huCo1aGm2_2),.dout(w_dff_B_eoxFidYA3_2),.clk(gclk));
	jdff dff_B_UZxZduZX0_2(.din(w_dff_B_eoxFidYA3_2),.dout(w_dff_B_UZxZduZX0_2),.clk(gclk));
	jdff dff_B_kOKqo6Ms2_2(.din(w_dff_B_UZxZduZX0_2),.dout(w_dff_B_kOKqo6Ms2_2),.clk(gclk));
	jdff dff_B_Rz7r1ZiV0_2(.din(w_dff_B_kOKqo6Ms2_2),.dout(w_dff_B_Rz7r1ZiV0_2),.clk(gclk));
	jdff dff_B_xoXXaG8G1_2(.din(w_dff_B_Rz7r1ZiV0_2),.dout(w_dff_B_xoXXaG8G1_2),.clk(gclk));
	jdff dff_B_okcYbJYB4_2(.din(w_dff_B_xoXXaG8G1_2),.dout(w_dff_B_okcYbJYB4_2),.clk(gclk));
	jdff dff_B_fsoFwImI9_2(.din(w_dff_B_okcYbJYB4_2),.dout(w_dff_B_fsoFwImI9_2),.clk(gclk));
	jdff dff_B_bYvR40qM9_2(.din(w_dff_B_fsoFwImI9_2),.dout(w_dff_B_bYvR40qM9_2),.clk(gclk));
	jdff dff_B_IjvRux7i0_2(.din(w_dff_B_bYvR40qM9_2),.dout(w_dff_B_IjvRux7i0_2),.clk(gclk));
	jdff dff_B_rBo1blwq5_2(.din(w_dff_B_IjvRux7i0_2),.dout(w_dff_B_rBo1blwq5_2),.clk(gclk));
	jdff dff_B_d9KG1JPN5_2(.din(w_dff_B_rBo1blwq5_2),.dout(w_dff_B_d9KG1JPN5_2),.clk(gclk));
	jdff dff_B_lRAeVbAg5_2(.din(w_dff_B_d9KG1JPN5_2),.dout(w_dff_B_lRAeVbAg5_2),.clk(gclk));
	jdff dff_B_1d86I5RD5_2(.din(w_dff_B_lRAeVbAg5_2),.dout(w_dff_B_1d86I5RD5_2),.clk(gclk));
	jdff dff_B_1w0Q7Pzv5_2(.din(n688),.dout(w_dff_B_1w0Q7Pzv5_2),.clk(gclk));
	jdff dff_B_9p2hFyFV9_1(.din(n653),.dout(w_dff_B_9p2hFyFV9_1),.clk(gclk));
	jdff dff_B_YSEJDdHr8_2(.din(n567),.dout(w_dff_B_YSEJDdHr8_2),.clk(gclk));
	jdff dff_B_7QtlJNFC1_2(.din(w_dff_B_YSEJDdHr8_2),.dout(w_dff_B_7QtlJNFC1_2),.clk(gclk));
	jdff dff_B_fecmAZju2_2(.din(w_dff_B_7QtlJNFC1_2),.dout(w_dff_B_fecmAZju2_2),.clk(gclk));
	jdff dff_B_T8h6c7c27_2(.din(w_dff_B_fecmAZju2_2),.dout(w_dff_B_T8h6c7c27_2),.clk(gclk));
	jdff dff_B_o93ULIuq9_2(.din(w_dff_B_T8h6c7c27_2),.dout(w_dff_B_o93ULIuq9_2),.clk(gclk));
	jdff dff_B_ZTAuuj942_2(.din(w_dff_B_o93ULIuq9_2),.dout(w_dff_B_ZTAuuj942_2),.clk(gclk));
	jdff dff_B_ZR2rgU1e0_2(.din(w_dff_B_ZTAuuj942_2),.dout(w_dff_B_ZR2rgU1e0_2),.clk(gclk));
	jdff dff_B_wXvfAy4a7_2(.din(w_dff_B_ZR2rgU1e0_2),.dout(w_dff_B_wXvfAy4a7_2),.clk(gclk));
	jdff dff_B_lkhQmSBd0_2(.din(w_dff_B_wXvfAy4a7_2),.dout(w_dff_B_lkhQmSBd0_2),.clk(gclk));
	jdff dff_B_E9KrE9Jw9_2(.din(w_dff_B_lkhQmSBd0_2),.dout(w_dff_B_E9KrE9Jw9_2),.clk(gclk));
	jdff dff_B_T3444ETd4_2(.din(w_dff_B_E9KrE9Jw9_2),.dout(w_dff_B_T3444ETd4_2),.clk(gclk));
	jdff dff_B_FMTujS1d9_2(.din(w_dff_B_T3444ETd4_2),.dout(w_dff_B_FMTujS1d9_2),.clk(gclk));
	jdff dff_B_P8mzXKyo4_2(.din(w_dff_B_FMTujS1d9_2),.dout(w_dff_B_P8mzXKyo4_2),.clk(gclk));
	jdff dff_B_yETXfUWg6_2(.din(w_dff_B_P8mzXKyo4_2),.dout(w_dff_B_yETXfUWg6_2),.clk(gclk));
	jdff dff_B_Kuevk1gs9_2(.din(n596),.dout(w_dff_B_Kuevk1gs9_2),.clk(gclk));
	jdff dff_B_IdxXSTVP0_1(.din(n568),.dout(w_dff_B_IdxXSTVP0_1),.clk(gclk));
	jdff dff_B_Jdk1nkM12_2(.din(n489),.dout(w_dff_B_Jdk1nkM12_2),.clk(gclk));
	jdff dff_B_9bO056u13_2(.din(w_dff_B_Jdk1nkM12_2),.dout(w_dff_B_9bO056u13_2),.clk(gclk));
	jdff dff_B_bmpZvaVQ5_2(.din(w_dff_B_9bO056u13_2),.dout(w_dff_B_bmpZvaVQ5_2),.clk(gclk));
	jdff dff_B_5yISK2Gy2_2(.din(w_dff_B_bmpZvaVQ5_2),.dout(w_dff_B_5yISK2Gy2_2),.clk(gclk));
	jdff dff_B_REIWgtRT8_2(.din(w_dff_B_5yISK2Gy2_2),.dout(w_dff_B_REIWgtRT8_2),.clk(gclk));
	jdff dff_B_NjLmuidY2_2(.din(w_dff_B_REIWgtRT8_2),.dout(w_dff_B_NjLmuidY2_2),.clk(gclk));
	jdff dff_B_IBGigjUL9_2(.din(w_dff_B_NjLmuidY2_2),.dout(w_dff_B_IBGigjUL9_2),.clk(gclk));
	jdff dff_B_2KEe7e9F6_2(.din(w_dff_B_IBGigjUL9_2),.dout(w_dff_B_2KEe7e9F6_2),.clk(gclk));
	jdff dff_B_ELg0OH7J0_2(.din(w_dff_B_2KEe7e9F6_2),.dout(w_dff_B_ELg0OH7J0_2),.clk(gclk));
	jdff dff_B_qVefu5aa2_2(.din(w_dff_B_ELg0OH7J0_2),.dout(w_dff_B_qVefu5aa2_2),.clk(gclk));
	jdff dff_B_dTMigAAZ6_2(.din(w_dff_B_qVefu5aa2_2),.dout(w_dff_B_dTMigAAZ6_2),.clk(gclk));
	jdff dff_B_p2ZwLPy27_2(.din(n511),.dout(w_dff_B_p2ZwLPy27_2),.clk(gclk));
	jdff dff_B_4uHK7tHT0_1(.din(n490),.dout(w_dff_B_4uHK7tHT0_1),.clk(gclk));
	jdff dff_B_6jM7pCO53_2(.din(n418),.dout(w_dff_B_6jM7pCO53_2),.clk(gclk));
	jdff dff_B_29AIBOeG6_2(.din(w_dff_B_6jM7pCO53_2),.dout(w_dff_B_29AIBOeG6_2),.clk(gclk));
	jdff dff_B_8jVsIgq90_2(.din(w_dff_B_29AIBOeG6_2),.dout(w_dff_B_8jVsIgq90_2),.clk(gclk));
	jdff dff_B_79Va2LeQ9_2(.din(w_dff_B_8jVsIgq90_2),.dout(w_dff_B_79Va2LeQ9_2),.clk(gclk));
	jdff dff_B_4Jefg1ts2_2(.din(w_dff_B_79Va2LeQ9_2),.dout(w_dff_B_4Jefg1ts2_2),.clk(gclk));
	jdff dff_B_f97bKrLE2_2(.din(w_dff_B_4Jefg1ts2_2),.dout(w_dff_B_f97bKrLE2_2),.clk(gclk));
	jdff dff_B_UNGCasGX6_2(.din(w_dff_B_f97bKrLE2_2),.dout(w_dff_B_UNGCasGX6_2),.clk(gclk));
	jdff dff_B_CuSaWmlk0_2(.din(w_dff_B_UNGCasGX6_2),.dout(w_dff_B_CuSaWmlk0_2),.clk(gclk));
	jdff dff_B_KCgyCyz10_2(.din(n433),.dout(w_dff_B_KCgyCyz10_2),.clk(gclk));
	jdff dff_B_4ORAqMPa0_2(.din(w_dff_B_KCgyCyz10_2),.dout(w_dff_B_4ORAqMPa0_2),.clk(gclk));
	jdff dff_B_zrQ40S7o4_2(.din(w_dff_B_4ORAqMPa0_2),.dout(w_dff_B_zrQ40S7o4_2),.clk(gclk));
	jdff dff_B_XEg0eNsw0_1(.din(n419),.dout(w_dff_B_XEg0eNsw0_1),.clk(gclk));
	jdff dff_B_7jFsosD90_1(.din(w_dff_B_XEg0eNsw0_1),.dout(w_dff_B_7jFsosD90_1),.clk(gclk));
	jdff dff_B_APjeyntA5_2(.din(n356),.dout(w_dff_B_APjeyntA5_2),.clk(gclk));
	jdff dff_B_VzrCsoqi0_2(.din(w_dff_B_APjeyntA5_2),.dout(w_dff_B_VzrCsoqi0_2),.clk(gclk));
	jdff dff_B_a8u7jpK85_2(.din(w_dff_B_VzrCsoqi0_2),.dout(w_dff_B_a8u7jpK85_2),.clk(gclk));
	jdff dff_B_PJsyqXJB2_0(.din(n361),.dout(w_dff_B_PJsyqXJB2_0),.clk(gclk));
	jdff dff_A_4mp05Umi5_0(.dout(w_n297_0[0]),.din(w_dff_A_4mp05Umi5_0),.clk(gclk));
	jdff dff_A_ErpNfXoR8_0(.dout(w_dff_A_4mp05Umi5_0),.din(w_dff_A_ErpNfXoR8_0),.clk(gclk));
	jdff dff_A_4pv54OEY1_1(.dout(w_n297_0[1]),.din(w_dff_A_4pv54OEY1_1),.clk(gclk));
	jdff dff_A_dAKuKW9I4_1(.dout(w_dff_A_4pv54OEY1_1),.din(w_dff_A_dAKuKW9I4_1),.clk(gclk));
	jdff dff_B_oYhPHKjl4_1(.din(n1594),.dout(w_dff_B_oYhPHKjl4_1),.clk(gclk));
	jdff dff_B_2iX1qkJR9_2(.din(n1535),.dout(w_dff_B_2iX1qkJR9_2),.clk(gclk));
	jdff dff_B_iPUBaDTI8_2(.din(w_dff_B_2iX1qkJR9_2),.dout(w_dff_B_iPUBaDTI8_2),.clk(gclk));
	jdff dff_B_kvLTVt0Z9_2(.din(w_dff_B_iPUBaDTI8_2),.dout(w_dff_B_kvLTVt0Z9_2),.clk(gclk));
	jdff dff_B_4htIGfre7_2(.din(w_dff_B_kvLTVt0Z9_2),.dout(w_dff_B_4htIGfre7_2),.clk(gclk));
	jdff dff_B_nd5vT7jX8_2(.din(w_dff_B_4htIGfre7_2),.dout(w_dff_B_nd5vT7jX8_2),.clk(gclk));
	jdff dff_B_rXjVEhCa5_2(.din(w_dff_B_nd5vT7jX8_2),.dout(w_dff_B_rXjVEhCa5_2),.clk(gclk));
	jdff dff_B_DkGFepT26_2(.din(w_dff_B_rXjVEhCa5_2),.dout(w_dff_B_DkGFepT26_2),.clk(gclk));
	jdff dff_B_BfvZLibs9_2(.din(w_dff_B_DkGFepT26_2),.dout(w_dff_B_BfvZLibs9_2),.clk(gclk));
	jdff dff_B_zoPKMN4e8_2(.din(w_dff_B_BfvZLibs9_2),.dout(w_dff_B_zoPKMN4e8_2),.clk(gclk));
	jdff dff_B_lJY29jr69_2(.din(w_dff_B_zoPKMN4e8_2),.dout(w_dff_B_lJY29jr69_2),.clk(gclk));
	jdff dff_B_ZYqT0wRN2_2(.din(w_dff_B_lJY29jr69_2),.dout(w_dff_B_ZYqT0wRN2_2),.clk(gclk));
	jdff dff_B_n4tp6VBk4_2(.din(w_dff_B_ZYqT0wRN2_2),.dout(w_dff_B_n4tp6VBk4_2),.clk(gclk));
	jdff dff_B_AAZ0HZk78_2(.din(w_dff_B_n4tp6VBk4_2),.dout(w_dff_B_AAZ0HZk78_2),.clk(gclk));
	jdff dff_B_jUZyEqdB8_2(.din(w_dff_B_AAZ0HZk78_2),.dout(w_dff_B_jUZyEqdB8_2),.clk(gclk));
	jdff dff_B_th0klIpv7_2(.din(w_dff_B_jUZyEqdB8_2),.dout(w_dff_B_th0klIpv7_2),.clk(gclk));
	jdff dff_B_76Gh53Sf5_2(.din(w_dff_B_th0klIpv7_2),.dout(w_dff_B_76Gh53Sf5_2),.clk(gclk));
	jdff dff_B_Z2dBzG2a3_2(.din(w_dff_B_76Gh53Sf5_2),.dout(w_dff_B_Z2dBzG2a3_2),.clk(gclk));
	jdff dff_B_0qQCfqbM7_2(.din(w_dff_B_Z2dBzG2a3_2),.dout(w_dff_B_0qQCfqbM7_2),.clk(gclk));
	jdff dff_B_3FCms8IU6_2(.din(w_dff_B_0qQCfqbM7_2),.dout(w_dff_B_3FCms8IU6_2),.clk(gclk));
	jdff dff_B_ddgBhsn63_2(.din(w_dff_B_3FCms8IU6_2),.dout(w_dff_B_ddgBhsn63_2),.clk(gclk));
	jdff dff_B_Wn0haHJ42_2(.din(w_dff_B_ddgBhsn63_2),.dout(w_dff_B_Wn0haHJ42_2),.clk(gclk));
	jdff dff_B_Qu2HyoT23_2(.din(w_dff_B_Wn0haHJ42_2),.dout(w_dff_B_Qu2HyoT23_2),.clk(gclk));
	jdff dff_B_kSgfh2fp8_2(.din(w_dff_B_Qu2HyoT23_2),.dout(w_dff_B_kSgfh2fp8_2),.clk(gclk));
	jdff dff_B_PSZTaUdt7_2(.din(w_dff_B_kSgfh2fp8_2),.dout(w_dff_B_PSZTaUdt7_2),.clk(gclk));
	jdff dff_B_nGPZtgZs5_2(.din(w_dff_B_PSZTaUdt7_2),.dout(w_dff_B_nGPZtgZs5_2),.clk(gclk));
	jdff dff_B_RZYqVgc03_2(.din(w_dff_B_nGPZtgZs5_2),.dout(w_dff_B_RZYqVgc03_2),.clk(gclk));
	jdff dff_B_3MKWqkmm5_2(.din(w_dff_B_RZYqVgc03_2),.dout(w_dff_B_3MKWqkmm5_2),.clk(gclk));
	jdff dff_B_Q3Z7tuAa4_2(.din(w_dff_B_3MKWqkmm5_2),.dout(w_dff_B_Q3Z7tuAa4_2),.clk(gclk));
	jdff dff_B_qRBu20oN3_2(.din(w_dff_B_Q3Z7tuAa4_2),.dout(w_dff_B_qRBu20oN3_2),.clk(gclk));
	jdff dff_B_F6YZlYos5_2(.din(w_dff_B_qRBu20oN3_2),.dout(w_dff_B_F6YZlYos5_2),.clk(gclk));
	jdff dff_B_7MbxxquT9_2(.din(w_dff_B_F6YZlYos5_2),.dout(w_dff_B_7MbxxquT9_2),.clk(gclk));
	jdff dff_B_b2tvfak68_2(.din(w_dff_B_7MbxxquT9_2),.dout(w_dff_B_b2tvfak68_2),.clk(gclk));
	jdff dff_B_2rWbq4s89_2(.din(w_dff_B_b2tvfak68_2),.dout(w_dff_B_2rWbq4s89_2),.clk(gclk));
	jdff dff_B_aQIXke7N9_2(.din(w_dff_B_2rWbq4s89_2),.dout(w_dff_B_aQIXke7N9_2),.clk(gclk));
	jdff dff_B_isxosnJW5_2(.din(w_dff_B_aQIXke7N9_2),.dout(w_dff_B_isxosnJW5_2),.clk(gclk));
	jdff dff_B_mnqzB8ou4_2(.din(w_dff_B_isxosnJW5_2),.dout(w_dff_B_mnqzB8ou4_2),.clk(gclk));
	jdff dff_B_aWtXyjR17_2(.din(w_dff_B_mnqzB8ou4_2),.dout(w_dff_B_aWtXyjR17_2),.clk(gclk));
	jdff dff_B_2U4AEvCd8_2(.din(w_dff_B_aWtXyjR17_2),.dout(w_dff_B_2U4AEvCd8_2),.clk(gclk));
	jdff dff_B_py8EmL695_2(.din(w_dff_B_2U4AEvCd8_2),.dout(w_dff_B_py8EmL695_2),.clk(gclk));
	jdff dff_B_gHiaeyQm2_2(.din(w_dff_B_py8EmL695_2),.dout(w_dff_B_gHiaeyQm2_2),.clk(gclk));
	jdff dff_B_r96ggMCF1_2(.din(w_dff_B_gHiaeyQm2_2),.dout(w_dff_B_r96ggMCF1_2),.clk(gclk));
	jdff dff_B_bdbI5LpD7_2(.din(w_dff_B_r96ggMCF1_2),.dout(w_dff_B_bdbI5LpD7_2),.clk(gclk));
	jdff dff_B_o10tMNDT3_2(.din(w_dff_B_bdbI5LpD7_2),.dout(w_dff_B_o10tMNDT3_2),.clk(gclk));
	jdff dff_B_8FEdDFRe5_2(.din(w_dff_B_o10tMNDT3_2),.dout(w_dff_B_8FEdDFRe5_2),.clk(gclk));
	jdff dff_B_XM4ocCmk3_2(.din(w_dff_B_8FEdDFRe5_2),.dout(w_dff_B_XM4ocCmk3_2),.clk(gclk));
	jdff dff_B_jZxX9Yif1_2(.din(w_dff_B_XM4ocCmk3_2),.dout(w_dff_B_jZxX9Yif1_2),.clk(gclk));
	jdff dff_B_BVI7x5lT3_0(.din(n1593),.dout(w_dff_B_BVI7x5lT3_0),.clk(gclk));
	jdff dff_A_ZZHp1yH95_1(.dout(w_n1581_0[1]),.din(w_dff_A_ZZHp1yH95_1),.clk(gclk));
	jdff dff_B_zsNagZtx2_1(.din(n1536),.dout(w_dff_B_zsNagZtx2_1),.clk(gclk));
	jdff dff_B_KQN9dBK23_2(.din(n1471),.dout(w_dff_B_KQN9dBK23_2),.clk(gclk));
	jdff dff_B_eURYiopo0_2(.din(w_dff_B_KQN9dBK23_2),.dout(w_dff_B_eURYiopo0_2),.clk(gclk));
	jdff dff_B_ccThDRwu2_2(.din(w_dff_B_eURYiopo0_2),.dout(w_dff_B_ccThDRwu2_2),.clk(gclk));
	jdff dff_B_MA36lqUx7_2(.din(w_dff_B_ccThDRwu2_2),.dout(w_dff_B_MA36lqUx7_2),.clk(gclk));
	jdff dff_B_Oqy4fChH6_2(.din(w_dff_B_MA36lqUx7_2),.dout(w_dff_B_Oqy4fChH6_2),.clk(gclk));
	jdff dff_B_ipOgdIF81_2(.din(w_dff_B_Oqy4fChH6_2),.dout(w_dff_B_ipOgdIF81_2),.clk(gclk));
	jdff dff_B_HonmLwBS7_2(.din(w_dff_B_ipOgdIF81_2),.dout(w_dff_B_HonmLwBS7_2),.clk(gclk));
	jdff dff_B_KCJ4womP2_2(.din(w_dff_B_HonmLwBS7_2),.dout(w_dff_B_KCJ4womP2_2),.clk(gclk));
	jdff dff_B_tjDW81ES4_2(.din(w_dff_B_KCJ4womP2_2),.dout(w_dff_B_tjDW81ES4_2),.clk(gclk));
	jdff dff_B_7wyXYK1F8_2(.din(w_dff_B_tjDW81ES4_2),.dout(w_dff_B_7wyXYK1F8_2),.clk(gclk));
	jdff dff_B_EMR9cLy91_2(.din(w_dff_B_7wyXYK1F8_2),.dout(w_dff_B_EMR9cLy91_2),.clk(gclk));
	jdff dff_B_h9sf2DD17_2(.din(w_dff_B_EMR9cLy91_2),.dout(w_dff_B_h9sf2DD17_2),.clk(gclk));
	jdff dff_B_1QPeJpFK7_2(.din(w_dff_B_h9sf2DD17_2),.dout(w_dff_B_1QPeJpFK7_2),.clk(gclk));
	jdff dff_B_HRpebVMQ4_2(.din(w_dff_B_1QPeJpFK7_2),.dout(w_dff_B_HRpebVMQ4_2),.clk(gclk));
	jdff dff_B_Vjz80nv38_2(.din(w_dff_B_HRpebVMQ4_2),.dout(w_dff_B_Vjz80nv38_2),.clk(gclk));
	jdff dff_B_VwtcjlgE8_2(.din(w_dff_B_Vjz80nv38_2),.dout(w_dff_B_VwtcjlgE8_2),.clk(gclk));
	jdff dff_B_8p9TZ9WH7_2(.din(w_dff_B_VwtcjlgE8_2),.dout(w_dff_B_8p9TZ9WH7_2),.clk(gclk));
	jdff dff_B_GUQdrqMZ4_2(.din(w_dff_B_8p9TZ9WH7_2),.dout(w_dff_B_GUQdrqMZ4_2),.clk(gclk));
	jdff dff_B_dRuvbDyk6_2(.din(w_dff_B_GUQdrqMZ4_2),.dout(w_dff_B_dRuvbDyk6_2),.clk(gclk));
	jdff dff_B_8izDSxvv1_2(.din(w_dff_B_dRuvbDyk6_2),.dout(w_dff_B_8izDSxvv1_2),.clk(gclk));
	jdff dff_B_vW27K4gl9_2(.din(w_dff_B_8izDSxvv1_2),.dout(w_dff_B_vW27K4gl9_2),.clk(gclk));
	jdff dff_B_c8f8wfBy5_2(.din(w_dff_B_vW27K4gl9_2),.dout(w_dff_B_c8f8wfBy5_2),.clk(gclk));
	jdff dff_B_akFMc7ZY1_2(.din(w_dff_B_c8f8wfBy5_2),.dout(w_dff_B_akFMc7ZY1_2),.clk(gclk));
	jdff dff_B_nVeiDsEe8_2(.din(w_dff_B_akFMc7ZY1_2),.dout(w_dff_B_nVeiDsEe8_2),.clk(gclk));
	jdff dff_B_SBu6N85x7_2(.din(w_dff_B_nVeiDsEe8_2),.dout(w_dff_B_SBu6N85x7_2),.clk(gclk));
	jdff dff_B_BRxuSeMW6_2(.din(w_dff_B_SBu6N85x7_2),.dout(w_dff_B_BRxuSeMW6_2),.clk(gclk));
	jdff dff_B_V2KEJ7W12_2(.din(w_dff_B_BRxuSeMW6_2),.dout(w_dff_B_V2KEJ7W12_2),.clk(gclk));
	jdff dff_B_7tv8BPpL8_2(.din(w_dff_B_V2KEJ7W12_2),.dout(w_dff_B_7tv8BPpL8_2),.clk(gclk));
	jdff dff_B_2WkUKoCC5_2(.din(w_dff_B_7tv8BPpL8_2),.dout(w_dff_B_2WkUKoCC5_2),.clk(gclk));
	jdff dff_B_kNuoio7N7_2(.din(w_dff_B_2WkUKoCC5_2),.dout(w_dff_B_kNuoio7N7_2),.clk(gclk));
	jdff dff_B_PRzlvdY87_2(.din(w_dff_B_kNuoio7N7_2),.dout(w_dff_B_PRzlvdY87_2),.clk(gclk));
	jdff dff_B_SVSYuJBJ3_2(.din(w_dff_B_PRzlvdY87_2),.dout(w_dff_B_SVSYuJBJ3_2),.clk(gclk));
	jdff dff_B_jKfmhyGq3_2(.din(w_dff_B_SVSYuJBJ3_2),.dout(w_dff_B_jKfmhyGq3_2),.clk(gclk));
	jdff dff_B_7itRnMKc8_2(.din(w_dff_B_jKfmhyGq3_2),.dout(w_dff_B_7itRnMKc8_2),.clk(gclk));
	jdff dff_B_ZMHvjRCv7_2(.din(w_dff_B_7itRnMKc8_2),.dout(w_dff_B_ZMHvjRCv7_2),.clk(gclk));
	jdff dff_B_PcpCVi0w7_2(.din(w_dff_B_ZMHvjRCv7_2),.dout(w_dff_B_PcpCVi0w7_2),.clk(gclk));
	jdff dff_B_XF04V13S3_2(.din(w_dff_B_PcpCVi0w7_2),.dout(w_dff_B_XF04V13S3_2),.clk(gclk));
	jdff dff_B_fQ5bDZ6e1_2(.din(w_dff_B_XF04V13S3_2),.dout(w_dff_B_fQ5bDZ6e1_2),.clk(gclk));
	jdff dff_B_MWkULhKK5_2(.din(w_dff_B_fQ5bDZ6e1_2),.dout(w_dff_B_MWkULhKK5_2),.clk(gclk));
	jdff dff_B_yDVmqgXH7_2(.din(w_dff_B_MWkULhKK5_2),.dout(w_dff_B_yDVmqgXH7_2),.clk(gclk));
	jdff dff_B_qRHni46W2_2(.din(w_dff_B_yDVmqgXH7_2),.dout(w_dff_B_qRHni46W2_2),.clk(gclk));
	jdff dff_B_FLkG0m4S9_2(.din(n1517),.dout(w_dff_B_FLkG0m4S9_2),.clk(gclk));
	jdff dff_B_jJuYpWOA2_1(.din(n1472),.dout(w_dff_B_jJuYpWOA2_1),.clk(gclk));
	jdff dff_B_5MebQy4y3_2(.din(n1400),.dout(w_dff_B_5MebQy4y3_2),.clk(gclk));
	jdff dff_B_tyil62C34_2(.din(w_dff_B_5MebQy4y3_2),.dout(w_dff_B_tyil62C34_2),.clk(gclk));
	jdff dff_B_wgyVInjP7_2(.din(w_dff_B_tyil62C34_2),.dout(w_dff_B_wgyVInjP7_2),.clk(gclk));
	jdff dff_B_EI2UErS63_2(.din(w_dff_B_wgyVInjP7_2),.dout(w_dff_B_EI2UErS63_2),.clk(gclk));
	jdff dff_B_GaCBY2Zp1_2(.din(w_dff_B_EI2UErS63_2),.dout(w_dff_B_GaCBY2Zp1_2),.clk(gclk));
	jdff dff_B_JShO2dtC3_2(.din(w_dff_B_GaCBY2Zp1_2),.dout(w_dff_B_JShO2dtC3_2),.clk(gclk));
	jdff dff_B_19s6xN4c4_2(.din(w_dff_B_JShO2dtC3_2),.dout(w_dff_B_19s6xN4c4_2),.clk(gclk));
	jdff dff_B_Tcm7HXuR9_2(.din(w_dff_B_19s6xN4c4_2),.dout(w_dff_B_Tcm7HXuR9_2),.clk(gclk));
	jdff dff_B_gfMISfdO3_2(.din(w_dff_B_Tcm7HXuR9_2),.dout(w_dff_B_gfMISfdO3_2),.clk(gclk));
	jdff dff_B_8DVVGD8C6_2(.din(w_dff_B_gfMISfdO3_2),.dout(w_dff_B_8DVVGD8C6_2),.clk(gclk));
	jdff dff_B_Ff1yS4UM3_2(.din(w_dff_B_8DVVGD8C6_2),.dout(w_dff_B_Ff1yS4UM3_2),.clk(gclk));
	jdff dff_B_wUmCV5oz1_2(.din(w_dff_B_Ff1yS4UM3_2),.dout(w_dff_B_wUmCV5oz1_2),.clk(gclk));
	jdff dff_B_uLafZMRB4_2(.din(w_dff_B_wUmCV5oz1_2),.dout(w_dff_B_uLafZMRB4_2),.clk(gclk));
	jdff dff_B_yo6FGxEx2_2(.din(w_dff_B_uLafZMRB4_2),.dout(w_dff_B_yo6FGxEx2_2),.clk(gclk));
	jdff dff_B_utpluYEb2_2(.din(w_dff_B_yo6FGxEx2_2),.dout(w_dff_B_utpluYEb2_2),.clk(gclk));
	jdff dff_B_2qKwkANa9_2(.din(w_dff_B_utpluYEb2_2),.dout(w_dff_B_2qKwkANa9_2),.clk(gclk));
	jdff dff_B_3YeARK4s5_2(.din(w_dff_B_2qKwkANa9_2),.dout(w_dff_B_3YeARK4s5_2),.clk(gclk));
	jdff dff_B_rxn99gtp8_2(.din(w_dff_B_3YeARK4s5_2),.dout(w_dff_B_rxn99gtp8_2),.clk(gclk));
	jdff dff_B_I15Z2ViY3_2(.din(w_dff_B_rxn99gtp8_2),.dout(w_dff_B_I15Z2ViY3_2),.clk(gclk));
	jdff dff_B_yJylDi858_2(.din(w_dff_B_I15Z2ViY3_2),.dout(w_dff_B_yJylDi858_2),.clk(gclk));
	jdff dff_B_3nJajgoy7_2(.din(w_dff_B_yJylDi858_2),.dout(w_dff_B_3nJajgoy7_2),.clk(gclk));
	jdff dff_B_bqEsBQLj2_2(.din(w_dff_B_3nJajgoy7_2),.dout(w_dff_B_bqEsBQLj2_2),.clk(gclk));
	jdff dff_B_WdLbnMT72_2(.din(w_dff_B_bqEsBQLj2_2),.dout(w_dff_B_WdLbnMT72_2),.clk(gclk));
	jdff dff_B_vPDYpPKz5_2(.din(w_dff_B_WdLbnMT72_2),.dout(w_dff_B_vPDYpPKz5_2),.clk(gclk));
	jdff dff_B_R5vCPNJl1_2(.din(w_dff_B_vPDYpPKz5_2),.dout(w_dff_B_R5vCPNJl1_2),.clk(gclk));
	jdff dff_B_Mh8hxsIz2_2(.din(w_dff_B_R5vCPNJl1_2),.dout(w_dff_B_Mh8hxsIz2_2),.clk(gclk));
	jdff dff_B_RhJvNJP53_2(.din(w_dff_B_Mh8hxsIz2_2),.dout(w_dff_B_RhJvNJP53_2),.clk(gclk));
	jdff dff_B_HDt627Dx1_2(.din(w_dff_B_RhJvNJP53_2),.dout(w_dff_B_HDt627Dx1_2),.clk(gclk));
	jdff dff_B_qHekgAvu2_2(.din(w_dff_B_HDt627Dx1_2),.dout(w_dff_B_qHekgAvu2_2),.clk(gclk));
	jdff dff_B_0CAk07Ti4_2(.din(w_dff_B_qHekgAvu2_2),.dout(w_dff_B_0CAk07Ti4_2),.clk(gclk));
	jdff dff_B_t0QCoj4S8_2(.din(w_dff_B_0CAk07Ti4_2),.dout(w_dff_B_t0QCoj4S8_2),.clk(gclk));
	jdff dff_B_rdBYLdR77_2(.din(w_dff_B_t0QCoj4S8_2),.dout(w_dff_B_rdBYLdR77_2),.clk(gclk));
	jdff dff_B_hASYa8Ly5_2(.din(w_dff_B_rdBYLdR77_2),.dout(w_dff_B_hASYa8Ly5_2),.clk(gclk));
	jdff dff_B_fthatEhs0_2(.din(w_dff_B_hASYa8Ly5_2),.dout(w_dff_B_fthatEhs0_2),.clk(gclk));
	jdff dff_B_YcsuVGtl3_2(.din(w_dff_B_fthatEhs0_2),.dout(w_dff_B_YcsuVGtl3_2),.clk(gclk));
	jdff dff_B_c7dTpPDR9_2(.din(w_dff_B_YcsuVGtl3_2),.dout(w_dff_B_c7dTpPDR9_2),.clk(gclk));
	jdff dff_B_GZUGlUZm7_2(.din(w_dff_B_c7dTpPDR9_2),.dout(w_dff_B_GZUGlUZm7_2),.clk(gclk));
	jdff dff_B_o7k5VhFC6_2(.din(w_dff_B_GZUGlUZm7_2),.dout(w_dff_B_o7k5VhFC6_2),.clk(gclk));
	jdff dff_B_3LZA2KGF3_2(.din(n1446),.dout(w_dff_B_3LZA2KGF3_2),.clk(gclk));
	jdff dff_B_mI1SzJPV7_1(.din(n1401),.dout(w_dff_B_mI1SzJPV7_1),.clk(gclk));
	jdff dff_B_MS5RgPOK3_2(.din(n1322),.dout(w_dff_B_MS5RgPOK3_2),.clk(gclk));
	jdff dff_B_qvjMcSCF3_2(.din(w_dff_B_MS5RgPOK3_2),.dout(w_dff_B_qvjMcSCF3_2),.clk(gclk));
	jdff dff_B_pAfmfhW22_2(.din(w_dff_B_qvjMcSCF3_2),.dout(w_dff_B_pAfmfhW22_2),.clk(gclk));
	jdff dff_B_3ArIR8xx7_2(.din(w_dff_B_pAfmfhW22_2),.dout(w_dff_B_3ArIR8xx7_2),.clk(gclk));
	jdff dff_B_4jukcp5a0_2(.din(w_dff_B_3ArIR8xx7_2),.dout(w_dff_B_4jukcp5a0_2),.clk(gclk));
	jdff dff_B_xkjF5DsQ3_2(.din(w_dff_B_4jukcp5a0_2),.dout(w_dff_B_xkjF5DsQ3_2),.clk(gclk));
	jdff dff_B_nmFDYMGB6_2(.din(w_dff_B_xkjF5DsQ3_2),.dout(w_dff_B_nmFDYMGB6_2),.clk(gclk));
	jdff dff_B_kdyF9wor8_2(.din(w_dff_B_nmFDYMGB6_2),.dout(w_dff_B_kdyF9wor8_2),.clk(gclk));
	jdff dff_B_IjgkynGZ4_2(.din(w_dff_B_kdyF9wor8_2),.dout(w_dff_B_IjgkynGZ4_2),.clk(gclk));
	jdff dff_B_ThGcIjRc9_2(.din(w_dff_B_IjgkynGZ4_2),.dout(w_dff_B_ThGcIjRc9_2),.clk(gclk));
	jdff dff_B_BjQXxbml7_2(.din(w_dff_B_ThGcIjRc9_2),.dout(w_dff_B_BjQXxbml7_2),.clk(gclk));
	jdff dff_B_fN3cWTD72_2(.din(w_dff_B_BjQXxbml7_2),.dout(w_dff_B_fN3cWTD72_2),.clk(gclk));
	jdff dff_B_GlbVVF2m8_2(.din(w_dff_B_fN3cWTD72_2),.dout(w_dff_B_GlbVVF2m8_2),.clk(gclk));
	jdff dff_B_KJzueAyN5_2(.din(w_dff_B_GlbVVF2m8_2),.dout(w_dff_B_KJzueAyN5_2),.clk(gclk));
	jdff dff_B_UI78CJEv9_2(.din(w_dff_B_KJzueAyN5_2),.dout(w_dff_B_UI78CJEv9_2),.clk(gclk));
	jdff dff_B_XE56vBG73_2(.din(w_dff_B_UI78CJEv9_2),.dout(w_dff_B_XE56vBG73_2),.clk(gclk));
	jdff dff_B_mDgqSqOO8_2(.din(w_dff_B_XE56vBG73_2),.dout(w_dff_B_mDgqSqOO8_2),.clk(gclk));
	jdff dff_B_bivT0ACb9_2(.din(w_dff_B_mDgqSqOO8_2),.dout(w_dff_B_bivT0ACb9_2),.clk(gclk));
	jdff dff_B_ETGiKMWk9_2(.din(w_dff_B_bivT0ACb9_2),.dout(w_dff_B_ETGiKMWk9_2),.clk(gclk));
	jdff dff_B_IgeJkEo30_2(.din(w_dff_B_ETGiKMWk9_2),.dout(w_dff_B_IgeJkEo30_2),.clk(gclk));
	jdff dff_B_XEYGXgFd2_2(.din(w_dff_B_IgeJkEo30_2),.dout(w_dff_B_XEYGXgFd2_2),.clk(gclk));
	jdff dff_B_0qo0iBGN2_2(.din(w_dff_B_XEYGXgFd2_2),.dout(w_dff_B_0qo0iBGN2_2),.clk(gclk));
	jdff dff_B_VbUsVrxV3_2(.din(w_dff_B_0qo0iBGN2_2),.dout(w_dff_B_VbUsVrxV3_2),.clk(gclk));
	jdff dff_B_00pExPWt1_2(.din(w_dff_B_VbUsVrxV3_2),.dout(w_dff_B_00pExPWt1_2),.clk(gclk));
	jdff dff_B_6cjjXCw71_2(.din(w_dff_B_00pExPWt1_2),.dout(w_dff_B_6cjjXCw71_2),.clk(gclk));
	jdff dff_B_ZLEaQRx80_2(.din(w_dff_B_6cjjXCw71_2),.dout(w_dff_B_ZLEaQRx80_2),.clk(gclk));
	jdff dff_B_VSx8nG8j7_2(.din(w_dff_B_ZLEaQRx80_2),.dout(w_dff_B_VSx8nG8j7_2),.clk(gclk));
	jdff dff_B_K4o352yn0_2(.din(w_dff_B_VSx8nG8j7_2),.dout(w_dff_B_K4o352yn0_2),.clk(gclk));
	jdff dff_B_4Bk24P1w5_2(.din(w_dff_B_K4o352yn0_2),.dout(w_dff_B_4Bk24P1w5_2),.clk(gclk));
	jdff dff_B_5awZzLdr3_2(.din(w_dff_B_4Bk24P1w5_2),.dout(w_dff_B_5awZzLdr3_2),.clk(gclk));
	jdff dff_B_Bb8W7eVh7_2(.din(w_dff_B_5awZzLdr3_2),.dout(w_dff_B_Bb8W7eVh7_2),.clk(gclk));
	jdff dff_B_hDCKSB4k2_2(.din(w_dff_B_Bb8W7eVh7_2),.dout(w_dff_B_hDCKSB4k2_2),.clk(gclk));
	jdff dff_B_GIw7g1rw3_2(.din(w_dff_B_hDCKSB4k2_2),.dout(w_dff_B_GIw7g1rw3_2),.clk(gclk));
	jdff dff_B_6q6Jk2e22_2(.din(w_dff_B_GIw7g1rw3_2),.dout(w_dff_B_6q6Jk2e22_2),.clk(gclk));
	jdff dff_B_l85Ij3Ye7_2(.din(w_dff_B_6q6Jk2e22_2),.dout(w_dff_B_l85Ij3Ye7_2),.clk(gclk));
	jdff dff_B_Js1sOPgh7_2(.din(n1368),.dout(w_dff_B_Js1sOPgh7_2),.clk(gclk));
	jdff dff_B_LbZi72ql7_1(.din(n1323),.dout(w_dff_B_LbZi72ql7_1),.clk(gclk));
	jdff dff_B_YD1atmkx4_2(.din(n1237),.dout(w_dff_B_YD1atmkx4_2),.clk(gclk));
	jdff dff_B_L9fRZkbE5_2(.din(w_dff_B_YD1atmkx4_2),.dout(w_dff_B_L9fRZkbE5_2),.clk(gclk));
	jdff dff_B_IJfShoji8_2(.din(w_dff_B_L9fRZkbE5_2),.dout(w_dff_B_IJfShoji8_2),.clk(gclk));
	jdff dff_B_udOBCeIp6_2(.din(w_dff_B_IJfShoji8_2),.dout(w_dff_B_udOBCeIp6_2),.clk(gclk));
	jdff dff_B_3A8ESZVg6_2(.din(w_dff_B_udOBCeIp6_2),.dout(w_dff_B_3A8ESZVg6_2),.clk(gclk));
	jdff dff_B_fJ7DtA105_2(.din(w_dff_B_3A8ESZVg6_2),.dout(w_dff_B_fJ7DtA105_2),.clk(gclk));
	jdff dff_B_5ZboEowH5_2(.din(w_dff_B_fJ7DtA105_2),.dout(w_dff_B_5ZboEowH5_2),.clk(gclk));
	jdff dff_B_zZyq1RD10_2(.din(w_dff_B_5ZboEowH5_2),.dout(w_dff_B_zZyq1RD10_2),.clk(gclk));
	jdff dff_B_QTtbc1qE5_2(.din(w_dff_B_zZyq1RD10_2),.dout(w_dff_B_QTtbc1qE5_2),.clk(gclk));
	jdff dff_B_iBCncV6B3_2(.din(w_dff_B_QTtbc1qE5_2),.dout(w_dff_B_iBCncV6B3_2),.clk(gclk));
	jdff dff_B_zYn8Ogo56_2(.din(w_dff_B_iBCncV6B3_2),.dout(w_dff_B_zYn8Ogo56_2),.clk(gclk));
	jdff dff_B_wAP5mkC67_2(.din(w_dff_B_zYn8Ogo56_2),.dout(w_dff_B_wAP5mkC67_2),.clk(gclk));
	jdff dff_B_4N4eDkzd6_2(.din(w_dff_B_wAP5mkC67_2),.dout(w_dff_B_4N4eDkzd6_2),.clk(gclk));
	jdff dff_B_gy8SRj9I6_2(.din(w_dff_B_4N4eDkzd6_2),.dout(w_dff_B_gy8SRj9I6_2),.clk(gclk));
	jdff dff_B_hAVVkfDr8_2(.din(w_dff_B_gy8SRj9I6_2),.dout(w_dff_B_hAVVkfDr8_2),.clk(gclk));
	jdff dff_B_ZMha1dJU1_2(.din(w_dff_B_hAVVkfDr8_2),.dout(w_dff_B_ZMha1dJU1_2),.clk(gclk));
	jdff dff_B_n4xlXqnW0_2(.din(w_dff_B_ZMha1dJU1_2),.dout(w_dff_B_n4xlXqnW0_2),.clk(gclk));
	jdff dff_B_ozvO78aK6_2(.din(w_dff_B_n4xlXqnW0_2),.dout(w_dff_B_ozvO78aK6_2),.clk(gclk));
	jdff dff_B_Z3pIL7yF1_2(.din(w_dff_B_ozvO78aK6_2),.dout(w_dff_B_Z3pIL7yF1_2),.clk(gclk));
	jdff dff_B_ncMAgAVV0_2(.din(w_dff_B_Z3pIL7yF1_2),.dout(w_dff_B_ncMAgAVV0_2),.clk(gclk));
	jdff dff_B_GK5mYZBb3_2(.din(w_dff_B_ncMAgAVV0_2),.dout(w_dff_B_GK5mYZBb3_2),.clk(gclk));
	jdff dff_B_9L7cTObu3_2(.din(w_dff_B_GK5mYZBb3_2),.dout(w_dff_B_9L7cTObu3_2),.clk(gclk));
	jdff dff_B_3ufLWbKX6_2(.din(w_dff_B_9L7cTObu3_2),.dout(w_dff_B_3ufLWbKX6_2),.clk(gclk));
	jdff dff_B_uEG9OSjB3_2(.din(w_dff_B_3ufLWbKX6_2),.dout(w_dff_B_uEG9OSjB3_2),.clk(gclk));
	jdff dff_B_cRTjQz4a7_2(.din(w_dff_B_uEG9OSjB3_2),.dout(w_dff_B_cRTjQz4a7_2),.clk(gclk));
	jdff dff_B_SKMJ9imk3_2(.din(w_dff_B_cRTjQz4a7_2),.dout(w_dff_B_SKMJ9imk3_2),.clk(gclk));
	jdff dff_B_JJQPVFb56_2(.din(w_dff_B_SKMJ9imk3_2),.dout(w_dff_B_JJQPVFb56_2),.clk(gclk));
	jdff dff_B_FGseNpCy1_2(.din(w_dff_B_JJQPVFb56_2),.dout(w_dff_B_FGseNpCy1_2),.clk(gclk));
	jdff dff_B_kVwVwxbL3_2(.din(w_dff_B_FGseNpCy1_2),.dout(w_dff_B_kVwVwxbL3_2),.clk(gclk));
	jdff dff_B_I1W31Ccg7_2(.din(w_dff_B_kVwVwxbL3_2),.dout(w_dff_B_I1W31Ccg7_2),.clk(gclk));
	jdff dff_B_7q09bgBt4_2(.din(w_dff_B_I1W31Ccg7_2),.dout(w_dff_B_7q09bgBt4_2),.clk(gclk));
	jdff dff_B_okKF1GY07_2(.din(w_dff_B_7q09bgBt4_2),.dout(w_dff_B_okKF1GY07_2),.clk(gclk));
	jdff dff_B_6HhSHxWD4_2(.din(n1283),.dout(w_dff_B_6HhSHxWD4_2),.clk(gclk));
	jdff dff_B_zIUS8s871_1(.din(n1238),.dout(w_dff_B_zIUS8s871_1),.clk(gclk));
	jdff dff_B_NGDpqiWM6_2(.din(n1146),.dout(w_dff_B_NGDpqiWM6_2),.clk(gclk));
	jdff dff_B_bJa4WDH61_2(.din(w_dff_B_NGDpqiWM6_2),.dout(w_dff_B_bJa4WDH61_2),.clk(gclk));
	jdff dff_B_qaCn5nbH5_2(.din(w_dff_B_bJa4WDH61_2),.dout(w_dff_B_qaCn5nbH5_2),.clk(gclk));
	jdff dff_B_HlsJiCPB2_2(.din(w_dff_B_qaCn5nbH5_2),.dout(w_dff_B_HlsJiCPB2_2),.clk(gclk));
	jdff dff_B_lY9gyQlw8_2(.din(w_dff_B_HlsJiCPB2_2),.dout(w_dff_B_lY9gyQlw8_2),.clk(gclk));
	jdff dff_B_8bHfZIRA7_2(.din(w_dff_B_lY9gyQlw8_2),.dout(w_dff_B_8bHfZIRA7_2),.clk(gclk));
	jdff dff_B_qanxPJZu4_2(.din(w_dff_B_8bHfZIRA7_2),.dout(w_dff_B_qanxPJZu4_2),.clk(gclk));
	jdff dff_B_VG7ja1FN1_2(.din(w_dff_B_qanxPJZu4_2),.dout(w_dff_B_VG7ja1FN1_2),.clk(gclk));
	jdff dff_B_krFEi6Am1_2(.din(w_dff_B_VG7ja1FN1_2),.dout(w_dff_B_krFEi6Am1_2),.clk(gclk));
	jdff dff_B_yKbQhQDw4_2(.din(w_dff_B_krFEi6Am1_2),.dout(w_dff_B_yKbQhQDw4_2),.clk(gclk));
	jdff dff_B_Hqvy0AWD3_2(.din(w_dff_B_yKbQhQDw4_2),.dout(w_dff_B_Hqvy0AWD3_2),.clk(gclk));
	jdff dff_B_frCnMz7W3_2(.din(w_dff_B_Hqvy0AWD3_2),.dout(w_dff_B_frCnMz7W3_2),.clk(gclk));
	jdff dff_B_4iLs0C436_2(.din(w_dff_B_frCnMz7W3_2),.dout(w_dff_B_4iLs0C436_2),.clk(gclk));
	jdff dff_B_CA29PapU9_2(.din(w_dff_B_4iLs0C436_2),.dout(w_dff_B_CA29PapU9_2),.clk(gclk));
	jdff dff_B_nNKIWlm17_2(.din(w_dff_B_CA29PapU9_2),.dout(w_dff_B_nNKIWlm17_2),.clk(gclk));
	jdff dff_B_VkPwFpIc6_2(.din(w_dff_B_nNKIWlm17_2),.dout(w_dff_B_VkPwFpIc6_2),.clk(gclk));
	jdff dff_B_ODiWUEgl9_2(.din(w_dff_B_VkPwFpIc6_2),.dout(w_dff_B_ODiWUEgl9_2),.clk(gclk));
	jdff dff_B_1ZayYYam8_2(.din(w_dff_B_ODiWUEgl9_2),.dout(w_dff_B_1ZayYYam8_2),.clk(gclk));
	jdff dff_B_ftGECzqr9_2(.din(w_dff_B_1ZayYYam8_2),.dout(w_dff_B_ftGECzqr9_2),.clk(gclk));
	jdff dff_B_cuXEpZpm1_2(.din(w_dff_B_ftGECzqr9_2),.dout(w_dff_B_cuXEpZpm1_2),.clk(gclk));
	jdff dff_B_XvSGN2c00_2(.din(w_dff_B_cuXEpZpm1_2),.dout(w_dff_B_XvSGN2c00_2),.clk(gclk));
	jdff dff_B_jTdHultr4_2(.din(w_dff_B_XvSGN2c00_2),.dout(w_dff_B_jTdHultr4_2),.clk(gclk));
	jdff dff_B_0ACKFj0z7_2(.din(w_dff_B_jTdHultr4_2),.dout(w_dff_B_0ACKFj0z7_2),.clk(gclk));
	jdff dff_B_hyn5HOFb7_2(.din(w_dff_B_0ACKFj0z7_2),.dout(w_dff_B_hyn5HOFb7_2),.clk(gclk));
	jdff dff_B_LIatZtMR5_2(.din(w_dff_B_hyn5HOFb7_2),.dout(w_dff_B_LIatZtMR5_2),.clk(gclk));
	jdff dff_B_HSx2JnHT2_2(.din(w_dff_B_LIatZtMR5_2),.dout(w_dff_B_HSx2JnHT2_2),.clk(gclk));
	jdff dff_B_6HZ8KgQp6_2(.din(w_dff_B_HSx2JnHT2_2),.dout(w_dff_B_6HZ8KgQp6_2),.clk(gclk));
	jdff dff_B_DXGNdAQd6_2(.din(w_dff_B_6HZ8KgQp6_2),.dout(w_dff_B_DXGNdAQd6_2),.clk(gclk));
	jdff dff_B_WHme5axn2_2(.din(w_dff_B_DXGNdAQd6_2),.dout(w_dff_B_WHme5axn2_2),.clk(gclk));
	jdff dff_B_8UoqdxrN9_2(.din(n1192),.dout(w_dff_B_8UoqdxrN9_2),.clk(gclk));
	jdff dff_B_qGgjE1Rn5_1(.din(n1147),.dout(w_dff_B_qGgjE1Rn5_1),.clk(gclk));
	jdff dff_B_J6vRyHIx5_2(.din(n1048),.dout(w_dff_B_J6vRyHIx5_2),.clk(gclk));
	jdff dff_B_LeAaHmsT5_2(.din(w_dff_B_J6vRyHIx5_2),.dout(w_dff_B_LeAaHmsT5_2),.clk(gclk));
	jdff dff_B_9ANxlNdu9_2(.din(w_dff_B_LeAaHmsT5_2),.dout(w_dff_B_9ANxlNdu9_2),.clk(gclk));
	jdff dff_B_OhayqCGm0_2(.din(w_dff_B_9ANxlNdu9_2),.dout(w_dff_B_OhayqCGm0_2),.clk(gclk));
	jdff dff_B_WbQT8W073_2(.din(w_dff_B_OhayqCGm0_2),.dout(w_dff_B_WbQT8W073_2),.clk(gclk));
	jdff dff_B_Kcb3axph0_2(.din(w_dff_B_WbQT8W073_2),.dout(w_dff_B_Kcb3axph0_2),.clk(gclk));
	jdff dff_B_vEinAjQ44_2(.din(w_dff_B_Kcb3axph0_2),.dout(w_dff_B_vEinAjQ44_2),.clk(gclk));
	jdff dff_B_sNcA8fvc9_2(.din(w_dff_B_vEinAjQ44_2),.dout(w_dff_B_sNcA8fvc9_2),.clk(gclk));
	jdff dff_B_G1W2vT0s2_2(.din(w_dff_B_sNcA8fvc9_2),.dout(w_dff_B_G1W2vT0s2_2),.clk(gclk));
	jdff dff_B_IYklaDxc3_2(.din(w_dff_B_G1W2vT0s2_2),.dout(w_dff_B_IYklaDxc3_2),.clk(gclk));
	jdff dff_B_ySVQXHtq3_2(.din(w_dff_B_IYklaDxc3_2),.dout(w_dff_B_ySVQXHtq3_2),.clk(gclk));
	jdff dff_B_edYN6leQ4_2(.din(w_dff_B_ySVQXHtq3_2),.dout(w_dff_B_edYN6leQ4_2),.clk(gclk));
	jdff dff_B_zlpNHW0z1_2(.din(w_dff_B_edYN6leQ4_2),.dout(w_dff_B_zlpNHW0z1_2),.clk(gclk));
	jdff dff_B_e1nUaIqS3_2(.din(w_dff_B_zlpNHW0z1_2),.dout(w_dff_B_e1nUaIqS3_2),.clk(gclk));
	jdff dff_B_cWzcx7Zj3_2(.din(w_dff_B_e1nUaIqS3_2),.dout(w_dff_B_cWzcx7Zj3_2),.clk(gclk));
	jdff dff_B_o5Ssbzgm4_2(.din(w_dff_B_cWzcx7Zj3_2),.dout(w_dff_B_o5Ssbzgm4_2),.clk(gclk));
	jdff dff_B_ccHIVRvk7_2(.din(w_dff_B_o5Ssbzgm4_2),.dout(w_dff_B_ccHIVRvk7_2),.clk(gclk));
	jdff dff_B_zsCqAjJ61_2(.din(w_dff_B_ccHIVRvk7_2),.dout(w_dff_B_zsCqAjJ61_2),.clk(gclk));
	jdff dff_B_1wUjJCab7_2(.din(w_dff_B_zsCqAjJ61_2),.dout(w_dff_B_1wUjJCab7_2),.clk(gclk));
	jdff dff_B_ZoewvTH74_2(.din(w_dff_B_1wUjJCab7_2),.dout(w_dff_B_ZoewvTH74_2),.clk(gclk));
	jdff dff_B_6kQtoUCL0_2(.din(w_dff_B_ZoewvTH74_2),.dout(w_dff_B_6kQtoUCL0_2),.clk(gclk));
	jdff dff_B_sswBTdAv5_2(.din(w_dff_B_6kQtoUCL0_2),.dout(w_dff_B_sswBTdAv5_2),.clk(gclk));
	jdff dff_B_RijX5t8b1_2(.din(w_dff_B_sswBTdAv5_2),.dout(w_dff_B_RijX5t8b1_2),.clk(gclk));
	jdff dff_B_htjO9n1L6_2(.din(w_dff_B_RijX5t8b1_2),.dout(w_dff_B_htjO9n1L6_2),.clk(gclk));
	jdff dff_B_rPKIXgGq9_2(.din(w_dff_B_htjO9n1L6_2),.dout(w_dff_B_rPKIXgGq9_2),.clk(gclk));
	jdff dff_B_CSNfWwZN2_2(.din(w_dff_B_rPKIXgGq9_2),.dout(w_dff_B_CSNfWwZN2_2),.clk(gclk));
	jdff dff_B_pravOeJa6_2(.din(n1093),.dout(w_dff_B_pravOeJa6_2),.clk(gclk));
	jdff dff_B_NUJAPVTH1_1(.din(n1049),.dout(w_dff_B_NUJAPVTH1_1),.clk(gclk));
	jdff dff_B_zRSG50vb3_2(.din(n949),.dout(w_dff_B_zRSG50vb3_2),.clk(gclk));
	jdff dff_B_LdNbmbpL6_2(.din(w_dff_B_zRSG50vb3_2),.dout(w_dff_B_LdNbmbpL6_2),.clk(gclk));
	jdff dff_B_eyJX0G1q9_2(.din(w_dff_B_LdNbmbpL6_2),.dout(w_dff_B_eyJX0G1q9_2),.clk(gclk));
	jdff dff_B_gSZYEKnZ8_2(.din(w_dff_B_eyJX0G1q9_2),.dout(w_dff_B_gSZYEKnZ8_2),.clk(gclk));
	jdff dff_B_rtbX6WwV7_2(.din(w_dff_B_gSZYEKnZ8_2),.dout(w_dff_B_rtbX6WwV7_2),.clk(gclk));
	jdff dff_B_G8fcrtJZ6_2(.din(w_dff_B_rtbX6WwV7_2),.dout(w_dff_B_G8fcrtJZ6_2),.clk(gclk));
	jdff dff_B_kel6czC82_2(.din(w_dff_B_G8fcrtJZ6_2),.dout(w_dff_B_kel6czC82_2),.clk(gclk));
	jdff dff_B_wiPHTbKD7_2(.din(w_dff_B_kel6czC82_2),.dout(w_dff_B_wiPHTbKD7_2),.clk(gclk));
	jdff dff_B_kWIfkf4A4_2(.din(w_dff_B_wiPHTbKD7_2),.dout(w_dff_B_kWIfkf4A4_2),.clk(gclk));
	jdff dff_B_QOdgpeCl9_2(.din(w_dff_B_kWIfkf4A4_2),.dout(w_dff_B_QOdgpeCl9_2),.clk(gclk));
	jdff dff_B_Z1pTSHl80_2(.din(w_dff_B_QOdgpeCl9_2),.dout(w_dff_B_Z1pTSHl80_2),.clk(gclk));
	jdff dff_B_M6u4jiNH0_2(.din(w_dff_B_Z1pTSHl80_2),.dout(w_dff_B_M6u4jiNH0_2),.clk(gclk));
	jdff dff_B_Uokl5F1z8_2(.din(w_dff_B_M6u4jiNH0_2),.dout(w_dff_B_Uokl5F1z8_2),.clk(gclk));
	jdff dff_B_DCjcOa3G1_2(.din(w_dff_B_Uokl5F1z8_2),.dout(w_dff_B_DCjcOa3G1_2),.clk(gclk));
	jdff dff_B_CmtaG9eP2_2(.din(w_dff_B_DCjcOa3G1_2),.dout(w_dff_B_CmtaG9eP2_2),.clk(gclk));
	jdff dff_B_R6a7cuxy8_2(.din(w_dff_B_CmtaG9eP2_2),.dout(w_dff_B_R6a7cuxy8_2),.clk(gclk));
	jdff dff_B_2dLhHX765_2(.din(w_dff_B_R6a7cuxy8_2),.dout(w_dff_B_2dLhHX765_2),.clk(gclk));
	jdff dff_B_M9dEtoLm5_2(.din(w_dff_B_2dLhHX765_2),.dout(w_dff_B_M9dEtoLm5_2),.clk(gclk));
	jdff dff_B_6vzcQcFf2_2(.din(w_dff_B_M9dEtoLm5_2),.dout(w_dff_B_6vzcQcFf2_2),.clk(gclk));
	jdff dff_B_nIqNbTDI6_2(.din(w_dff_B_6vzcQcFf2_2),.dout(w_dff_B_nIqNbTDI6_2),.clk(gclk));
	jdff dff_B_6gGDwck35_2(.din(w_dff_B_nIqNbTDI6_2),.dout(w_dff_B_6gGDwck35_2),.clk(gclk));
	jdff dff_B_iCMIOgkW8_2(.din(w_dff_B_6gGDwck35_2),.dout(w_dff_B_iCMIOgkW8_2),.clk(gclk));
	jdff dff_B_2WUixItf6_2(.din(w_dff_B_iCMIOgkW8_2),.dout(w_dff_B_2WUixItf6_2),.clk(gclk));
	jdff dff_B_EqvHgSLD6_2(.din(n994),.dout(w_dff_B_EqvHgSLD6_2),.clk(gclk));
	jdff dff_B_SY1dVtdg4_1(.din(n950),.dout(w_dff_B_SY1dVtdg4_1),.clk(gclk));
	jdff dff_B_fdLQXVQC8_2(.din(n847),.dout(w_dff_B_fdLQXVQC8_2),.clk(gclk));
	jdff dff_B_750sclDP4_2(.din(w_dff_B_fdLQXVQC8_2),.dout(w_dff_B_750sclDP4_2),.clk(gclk));
	jdff dff_B_HYuka2wO9_2(.din(w_dff_B_750sclDP4_2),.dout(w_dff_B_HYuka2wO9_2),.clk(gclk));
	jdff dff_B_X6yIsHbD5_2(.din(w_dff_B_HYuka2wO9_2),.dout(w_dff_B_X6yIsHbD5_2),.clk(gclk));
	jdff dff_B_19xtU5IV1_2(.din(w_dff_B_X6yIsHbD5_2),.dout(w_dff_B_19xtU5IV1_2),.clk(gclk));
	jdff dff_B_KgMNJRlv7_2(.din(w_dff_B_19xtU5IV1_2),.dout(w_dff_B_KgMNJRlv7_2),.clk(gclk));
	jdff dff_B_EXM3HdVp7_2(.din(w_dff_B_KgMNJRlv7_2),.dout(w_dff_B_EXM3HdVp7_2),.clk(gclk));
	jdff dff_B_QALLJNme5_2(.din(w_dff_B_EXM3HdVp7_2),.dout(w_dff_B_QALLJNme5_2),.clk(gclk));
	jdff dff_B_gNGT0SeE9_2(.din(w_dff_B_QALLJNme5_2),.dout(w_dff_B_gNGT0SeE9_2),.clk(gclk));
	jdff dff_B_lxa6Uaao8_2(.din(w_dff_B_gNGT0SeE9_2),.dout(w_dff_B_lxa6Uaao8_2),.clk(gclk));
	jdff dff_B_DoJYQiuo5_2(.din(w_dff_B_lxa6Uaao8_2),.dout(w_dff_B_DoJYQiuo5_2),.clk(gclk));
	jdff dff_B_4jkqOUvD3_2(.din(w_dff_B_DoJYQiuo5_2),.dout(w_dff_B_4jkqOUvD3_2),.clk(gclk));
	jdff dff_B_Y2u2Mk3D1_2(.din(w_dff_B_4jkqOUvD3_2),.dout(w_dff_B_Y2u2Mk3D1_2),.clk(gclk));
	jdff dff_B_xiZ4gCn92_2(.din(w_dff_B_Y2u2Mk3D1_2),.dout(w_dff_B_xiZ4gCn92_2),.clk(gclk));
	jdff dff_B_5q2KSaA64_2(.din(w_dff_B_xiZ4gCn92_2),.dout(w_dff_B_5q2KSaA64_2),.clk(gclk));
	jdff dff_B_Uk2waCTi9_2(.din(w_dff_B_5q2KSaA64_2),.dout(w_dff_B_Uk2waCTi9_2),.clk(gclk));
	jdff dff_B_YuRtDOMr4_2(.din(w_dff_B_Uk2waCTi9_2),.dout(w_dff_B_YuRtDOMr4_2),.clk(gclk));
	jdff dff_B_2FmEnAqX6_2(.din(w_dff_B_YuRtDOMr4_2),.dout(w_dff_B_2FmEnAqX6_2),.clk(gclk));
	jdff dff_B_qKnUK94u4_2(.din(w_dff_B_2FmEnAqX6_2),.dout(w_dff_B_qKnUK94u4_2),.clk(gclk));
	jdff dff_B_xWjgITBo3_2(.din(w_dff_B_qKnUK94u4_2),.dout(w_dff_B_xWjgITBo3_2),.clk(gclk));
	jdff dff_B_YkoF4SCv4_2(.din(n888),.dout(w_dff_B_YkoF4SCv4_2),.clk(gclk));
	jdff dff_B_2GiWZanX5_1(.din(n848),.dout(w_dff_B_2GiWZanX5_1),.clk(gclk));
	jdff dff_B_72qZHXs54_2(.din(n749),.dout(w_dff_B_72qZHXs54_2),.clk(gclk));
	jdff dff_B_aRivU5J29_2(.din(w_dff_B_72qZHXs54_2),.dout(w_dff_B_aRivU5J29_2),.clk(gclk));
	jdff dff_B_NfatX3m43_2(.din(w_dff_B_aRivU5J29_2),.dout(w_dff_B_NfatX3m43_2),.clk(gclk));
	jdff dff_B_aYOv1SLd6_2(.din(w_dff_B_NfatX3m43_2),.dout(w_dff_B_aYOv1SLd6_2),.clk(gclk));
	jdff dff_B_8aJc6ERt4_2(.din(w_dff_B_aYOv1SLd6_2),.dout(w_dff_B_8aJc6ERt4_2),.clk(gclk));
	jdff dff_B_7O0Zkyjx4_2(.din(w_dff_B_8aJc6ERt4_2),.dout(w_dff_B_7O0Zkyjx4_2),.clk(gclk));
	jdff dff_B_Azy82fwj0_2(.din(w_dff_B_7O0Zkyjx4_2),.dout(w_dff_B_Azy82fwj0_2),.clk(gclk));
	jdff dff_B_gAWDaJPw5_2(.din(w_dff_B_Azy82fwj0_2),.dout(w_dff_B_gAWDaJPw5_2),.clk(gclk));
	jdff dff_B_DXuin0ol9_2(.din(w_dff_B_gAWDaJPw5_2),.dout(w_dff_B_DXuin0ol9_2),.clk(gclk));
	jdff dff_B_JZwvDQVf1_2(.din(w_dff_B_DXuin0ol9_2),.dout(w_dff_B_JZwvDQVf1_2),.clk(gclk));
	jdff dff_B_TnlsbTit6_2(.din(w_dff_B_JZwvDQVf1_2),.dout(w_dff_B_TnlsbTit6_2),.clk(gclk));
	jdff dff_B_57tzlzMX0_2(.din(w_dff_B_TnlsbTit6_2),.dout(w_dff_B_57tzlzMX0_2),.clk(gclk));
	jdff dff_B_Lvy2Z4Vx3_2(.din(w_dff_B_57tzlzMX0_2),.dout(w_dff_B_Lvy2Z4Vx3_2),.clk(gclk));
	jdff dff_B_LnA1wPUW8_2(.din(w_dff_B_Lvy2Z4Vx3_2),.dout(w_dff_B_LnA1wPUW8_2),.clk(gclk));
	jdff dff_B_SbImryn38_2(.din(w_dff_B_LnA1wPUW8_2),.dout(w_dff_B_SbImryn38_2),.clk(gclk));
	jdff dff_B_la7O5Nqs2_2(.din(w_dff_B_SbImryn38_2),.dout(w_dff_B_la7O5Nqs2_2),.clk(gclk));
	jdff dff_B_28pqL9by1_2(.din(w_dff_B_la7O5Nqs2_2),.dout(w_dff_B_28pqL9by1_2),.clk(gclk));
	jdff dff_B_cF7Ixm6x1_2(.din(n785),.dout(w_dff_B_cF7Ixm6x1_2),.clk(gclk));
	jdff dff_B_r9B0w8l35_1(.din(n750),.dout(w_dff_B_r9B0w8l35_1),.clk(gclk));
	jdff dff_B_ZEwr4JXt5_2(.din(n657),.dout(w_dff_B_ZEwr4JXt5_2),.clk(gclk));
	jdff dff_B_MesALP467_2(.din(w_dff_B_ZEwr4JXt5_2),.dout(w_dff_B_MesALP467_2),.clk(gclk));
	jdff dff_B_UifpdZWV3_2(.din(w_dff_B_MesALP467_2),.dout(w_dff_B_UifpdZWV3_2),.clk(gclk));
	jdff dff_B_M8txeVwG6_2(.din(w_dff_B_UifpdZWV3_2),.dout(w_dff_B_M8txeVwG6_2),.clk(gclk));
	jdff dff_B_oSMyBzXP0_2(.din(w_dff_B_M8txeVwG6_2),.dout(w_dff_B_oSMyBzXP0_2),.clk(gclk));
	jdff dff_B_XBkNE5nj7_2(.din(w_dff_B_oSMyBzXP0_2),.dout(w_dff_B_XBkNE5nj7_2),.clk(gclk));
	jdff dff_B_mnpElBUh1_2(.din(w_dff_B_XBkNE5nj7_2),.dout(w_dff_B_mnpElBUh1_2),.clk(gclk));
	jdff dff_B_7xLQkOa40_2(.din(w_dff_B_mnpElBUh1_2),.dout(w_dff_B_7xLQkOa40_2),.clk(gclk));
	jdff dff_B_fiMxtoMP6_2(.din(w_dff_B_7xLQkOa40_2),.dout(w_dff_B_fiMxtoMP6_2),.clk(gclk));
	jdff dff_B_pCmurpbL1_2(.din(w_dff_B_fiMxtoMP6_2),.dout(w_dff_B_pCmurpbL1_2),.clk(gclk));
	jdff dff_B_rYaauK352_2(.din(w_dff_B_pCmurpbL1_2),.dout(w_dff_B_rYaauK352_2),.clk(gclk));
	jdff dff_B_L9SLDhoh9_2(.din(w_dff_B_rYaauK352_2),.dout(w_dff_B_L9SLDhoh9_2),.clk(gclk));
	jdff dff_B_u9nCgL5q5_2(.din(w_dff_B_L9SLDhoh9_2),.dout(w_dff_B_u9nCgL5q5_2),.clk(gclk));
	jdff dff_B_yuiA1Rrp4_2(.din(w_dff_B_u9nCgL5q5_2),.dout(w_dff_B_yuiA1Rrp4_2),.clk(gclk));
	jdff dff_B_d8eQmLZH6_2(.din(n686),.dout(w_dff_B_d8eQmLZH6_2),.clk(gclk));
	jdff dff_B_m2Jk00NH5_1(.din(n658),.dout(w_dff_B_m2Jk00NH5_1),.clk(gclk));
	jdff dff_B_1epBzvRe8_2(.din(n572),.dout(w_dff_B_1epBzvRe8_2),.clk(gclk));
	jdff dff_B_0rgXNger8_2(.din(w_dff_B_1epBzvRe8_2),.dout(w_dff_B_0rgXNger8_2),.clk(gclk));
	jdff dff_B_sivrI2256_2(.din(w_dff_B_0rgXNger8_2),.dout(w_dff_B_sivrI2256_2),.clk(gclk));
	jdff dff_B_hRnZjd0z4_2(.din(w_dff_B_sivrI2256_2),.dout(w_dff_B_hRnZjd0z4_2),.clk(gclk));
	jdff dff_B_7J0qZQea2_2(.din(w_dff_B_hRnZjd0z4_2),.dout(w_dff_B_7J0qZQea2_2),.clk(gclk));
	jdff dff_B_7CdF4jer7_2(.din(w_dff_B_7J0qZQea2_2),.dout(w_dff_B_7CdF4jer7_2),.clk(gclk));
	jdff dff_B_XObOW2hW1_2(.din(w_dff_B_7CdF4jer7_2),.dout(w_dff_B_XObOW2hW1_2),.clk(gclk));
	jdff dff_B_jBAZemRm5_2(.din(w_dff_B_XObOW2hW1_2),.dout(w_dff_B_jBAZemRm5_2),.clk(gclk));
	jdff dff_B_dINjm7Ft0_2(.din(w_dff_B_jBAZemRm5_2),.dout(w_dff_B_dINjm7Ft0_2),.clk(gclk));
	jdff dff_B_JCuDsFxD7_2(.din(w_dff_B_dINjm7Ft0_2),.dout(w_dff_B_JCuDsFxD7_2),.clk(gclk));
	jdff dff_B_Bw3OsVie8_2(.din(w_dff_B_JCuDsFxD7_2),.dout(w_dff_B_Bw3OsVie8_2),.clk(gclk));
	jdff dff_B_iknV8gPt0_2(.din(n594),.dout(w_dff_B_iknV8gPt0_2),.clk(gclk));
	jdff dff_B_akOY61NU1_1(.din(n573),.dout(w_dff_B_akOY61NU1_1),.clk(gclk));
	jdff dff_B_HtscdnlW7_2(.din(n494),.dout(w_dff_B_HtscdnlW7_2),.clk(gclk));
	jdff dff_B_dVFGlK9i2_2(.din(w_dff_B_HtscdnlW7_2),.dout(w_dff_B_dVFGlK9i2_2),.clk(gclk));
	jdff dff_B_a6qujakw4_2(.din(w_dff_B_dVFGlK9i2_2),.dout(w_dff_B_a6qujakw4_2),.clk(gclk));
	jdff dff_B_kb1pdHTW2_2(.din(w_dff_B_a6qujakw4_2),.dout(w_dff_B_kb1pdHTW2_2),.clk(gclk));
	jdff dff_B_5YBzyBpb5_2(.din(w_dff_B_kb1pdHTW2_2),.dout(w_dff_B_5YBzyBpb5_2),.clk(gclk));
	jdff dff_B_HonZBjHB0_2(.din(w_dff_B_5YBzyBpb5_2),.dout(w_dff_B_HonZBjHB0_2),.clk(gclk));
	jdff dff_B_a37YOQbf1_2(.din(w_dff_B_HonZBjHB0_2),.dout(w_dff_B_a37YOQbf1_2),.clk(gclk));
	jdff dff_B_sW1vra5Q7_2(.din(w_dff_B_a37YOQbf1_2),.dout(w_dff_B_sW1vra5Q7_2),.clk(gclk));
	jdff dff_B_ct0g8B0Q6_2(.din(n509),.dout(w_dff_B_ct0g8B0Q6_2),.clk(gclk));
	jdff dff_B_7EClZ9OK6_2(.din(w_dff_B_ct0g8B0Q6_2),.dout(w_dff_B_7EClZ9OK6_2),.clk(gclk));
	jdff dff_B_bSzKJyA47_2(.din(w_dff_B_7EClZ9OK6_2),.dout(w_dff_B_bSzKJyA47_2),.clk(gclk));
	jdff dff_B_IxrNAbwX9_1(.din(n495),.dout(w_dff_B_IxrNAbwX9_1),.clk(gclk));
	jdff dff_B_9kJ7FV726_1(.din(w_dff_B_IxrNAbwX9_1),.dout(w_dff_B_9kJ7FV726_1),.clk(gclk));
	jdff dff_B_MIJfWOow1_2(.din(n425),.dout(w_dff_B_MIJfWOow1_2),.clk(gclk));
	jdff dff_B_UcTY9fRj4_2(.din(w_dff_B_MIJfWOow1_2),.dout(w_dff_B_UcTY9fRj4_2),.clk(gclk));
	jdff dff_B_QGJTPq0i6_2(.din(w_dff_B_UcTY9fRj4_2),.dout(w_dff_B_QGJTPq0i6_2),.clk(gclk));
	jdff dff_B_CBpFB20e9_0(.din(n430),.dout(w_dff_B_CBpFB20e9_0),.clk(gclk));
	jdff dff_A_CigddwwK4_0(.dout(w_n358_0[0]),.din(w_dff_A_CigddwwK4_0),.clk(gclk));
	jdff dff_A_PN5thRrM1_0(.dout(w_dff_A_CigddwwK4_0),.din(w_dff_A_PN5thRrM1_0),.clk(gclk));
	jdff dff_A_dB2hOinj9_1(.dout(w_n358_0[1]),.din(w_dff_A_dB2hOinj9_1),.clk(gclk));
	jdff dff_A_iBKlWHFh0_1(.dout(w_dff_A_dB2hOinj9_1),.din(w_dff_A_iBKlWHFh0_1),.clk(gclk));
	jdff dff_B_PRuDwE9Y3_2(.din(n1651),.dout(w_dff_B_PRuDwE9Y3_2),.clk(gclk));
	jdff dff_B_fQdaedm32_1(.din(n1649),.dout(w_dff_B_fQdaedm32_1),.clk(gclk));
	jdff dff_B_To1rGYVT8_2(.din(n1597),.dout(w_dff_B_To1rGYVT8_2),.clk(gclk));
	jdff dff_B_gOnr7dGR8_2(.din(w_dff_B_To1rGYVT8_2),.dout(w_dff_B_gOnr7dGR8_2),.clk(gclk));
	jdff dff_B_rPV06Wdr9_2(.din(w_dff_B_gOnr7dGR8_2),.dout(w_dff_B_rPV06Wdr9_2),.clk(gclk));
	jdff dff_B_4yiI2Aek3_2(.din(w_dff_B_rPV06Wdr9_2),.dout(w_dff_B_4yiI2Aek3_2),.clk(gclk));
	jdff dff_B_gRBa6ZD10_2(.din(w_dff_B_4yiI2Aek3_2),.dout(w_dff_B_gRBa6ZD10_2),.clk(gclk));
	jdff dff_B_2FswoSkg0_2(.din(w_dff_B_gRBa6ZD10_2),.dout(w_dff_B_2FswoSkg0_2),.clk(gclk));
	jdff dff_B_bBDIiziW4_2(.din(w_dff_B_2FswoSkg0_2),.dout(w_dff_B_bBDIiziW4_2),.clk(gclk));
	jdff dff_B_mb1cISqR2_2(.din(w_dff_B_bBDIiziW4_2),.dout(w_dff_B_mb1cISqR2_2),.clk(gclk));
	jdff dff_B_wJjhnMvt3_2(.din(w_dff_B_mb1cISqR2_2),.dout(w_dff_B_wJjhnMvt3_2),.clk(gclk));
	jdff dff_B_93Fd7zLP2_2(.din(w_dff_B_wJjhnMvt3_2),.dout(w_dff_B_93Fd7zLP2_2),.clk(gclk));
	jdff dff_B_Wt3wfxyq9_2(.din(w_dff_B_93Fd7zLP2_2),.dout(w_dff_B_Wt3wfxyq9_2),.clk(gclk));
	jdff dff_B_eG1fY8XZ7_2(.din(w_dff_B_Wt3wfxyq9_2),.dout(w_dff_B_eG1fY8XZ7_2),.clk(gclk));
	jdff dff_B_pMYxWNMv7_2(.din(w_dff_B_eG1fY8XZ7_2),.dout(w_dff_B_pMYxWNMv7_2),.clk(gclk));
	jdff dff_B_aktjuSIn8_2(.din(w_dff_B_pMYxWNMv7_2),.dout(w_dff_B_aktjuSIn8_2),.clk(gclk));
	jdff dff_B_0QUl3x8T0_2(.din(w_dff_B_aktjuSIn8_2),.dout(w_dff_B_0QUl3x8T0_2),.clk(gclk));
	jdff dff_B_xN17xPVe2_2(.din(w_dff_B_0QUl3x8T0_2),.dout(w_dff_B_xN17xPVe2_2),.clk(gclk));
	jdff dff_B_oI0bT2ii7_2(.din(w_dff_B_xN17xPVe2_2),.dout(w_dff_B_oI0bT2ii7_2),.clk(gclk));
	jdff dff_B_3Jg0OAzJ5_2(.din(w_dff_B_oI0bT2ii7_2),.dout(w_dff_B_3Jg0OAzJ5_2),.clk(gclk));
	jdff dff_B_sVdn2fhy7_2(.din(w_dff_B_3Jg0OAzJ5_2),.dout(w_dff_B_sVdn2fhy7_2),.clk(gclk));
	jdff dff_B_fVGi4qnx7_2(.din(w_dff_B_sVdn2fhy7_2),.dout(w_dff_B_fVGi4qnx7_2),.clk(gclk));
	jdff dff_B_AMkpMV9r8_2(.din(w_dff_B_fVGi4qnx7_2),.dout(w_dff_B_AMkpMV9r8_2),.clk(gclk));
	jdff dff_B_K4u83C0p8_2(.din(w_dff_B_AMkpMV9r8_2),.dout(w_dff_B_K4u83C0p8_2),.clk(gclk));
	jdff dff_B_ltjsJ0Mk8_2(.din(w_dff_B_K4u83C0p8_2),.dout(w_dff_B_ltjsJ0Mk8_2),.clk(gclk));
	jdff dff_B_9sfKQkEq8_2(.din(w_dff_B_ltjsJ0Mk8_2),.dout(w_dff_B_9sfKQkEq8_2),.clk(gclk));
	jdff dff_B_8vH6OZhe0_2(.din(w_dff_B_9sfKQkEq8_2),.dout(w_dff_B_8vH6OZhe0_2),.clk(gclk));
	jdff dff_B_utd7gkqZ0_2(.din(w_dff_B_8vH6OZhe0_2),.dout(w_dff_B_utd7gkqZ0_2),.clk(gclk));
	jdff dff_B_wtuzRUED7_2(.din(w_dff_B_utd7gkqZ0_2),.dout(w_dff_B_wtuzRUED7_2),.clk(gclk));
	jdff dff_B_2Seqvs3J0_2(.din(w_dff_B_wtuzRUED7_2),.dout(w_dff_B_2Seqvs3J0_2),.clk(gclk));
	jdff dff_B_vFSIWNtd6_2(.din(w_dff_B_2Seqvs3J0_2),.dout(w_dff_B_vFSIWNtd6_2),.clk(gclk));
	jdff dff_B_qB5EOR3P9_2(.din(w_dff_B_vFSIWNtd6_2),.dout(w_dff_B_qB5EOR3P9_2),.clk(gclk));
	jdff dff_B_2C8aICjN2_2(.din(w_dff_B_qB5EOR3P9_2),.dout(w_dff_B_2C8aICjN2_2),.clk(gclk));
	jdff dff_B_3JP1qNqk0_2(.din(w_dff_B_2C8aICjN2_2),.dout(w_dff_B_3JP1qNqk0_2),.clk(gclk));
	jdff dff_B_9mcI6qZF7_2(.din(w_dff_B_3JP1qNqk0_2),.dout(w_dff_B_9mcI6qZF7_2),.clk(gclk));
	jdff dff_B_ikMCDLfs7_2(.din(w_dff_B_9mcI6qZF7_2),.dout(w_dff_B_ikMCDLfs7_2),.clk(gclk));
	jdff dff_B_vHHCFOAW5_2(.din(w_dff_B_ikMCDLfs7_2),.dout(w_dff_B_vHHCFOAW5_2),.clk(gclk));
	jdff dff_B_c2TpOike2_2(.din(w_dff_B_vHHCFOAW5_2),.dout(w_dff_B_c2TpOike2_2),.clk(gclk));
	jdff dff_B_IjOpXgSA9_2(.din(w_dff_B_c2TpOike2_2),.dout(w_dff_B_IjOpXgSA9_2),.clk(gclk));
	jdff dff_B_CsWSkPJk0_2(.din(w_dff_B_IjOpXgSA9_2),.dout(w_dff_B_CsWSkPJk0_2),.clk(gclk));
	jdff dff_B_bkPas9l87_2(.din(w_dff_B_CsWSkPJk0_2),.dout(w_dff_B_bkPas9l87_2),.clk(gclk));
	jdff dff_B_N84NUNze8_2(.din(w_dff_B_bkPas9l87_2),.dout(w_dff_B_N84NUNze8_2),.clk(gclk));
	jdff dff_B_5oPFgi4G2_2(.din(w_dff_B_N84NUNze8_2),.dout(w_dff_B_5oPFgi4G2_2),.clk(gclk));
	jdff dff_B_SbvijqDi9_2(.din(w_dff_B_5oPFgi4G2_2),.dout(w_dff_B_SbvijqDi9_2),.clk(gclk));
	jdff dff_B_L5qjy5tn6_2(.din(w_dff_B_SbvijqDi9_2),.dout(w_dff_B_L5qjy5tn6_2),.clk(gclk));
	jdff dff_B_6U8373391_2(.din(w_dff_B_L5qjy5tn6_2),.dout(w_dff_B_6U8373391_2),.clk(gclk));
	jdff dff_B_RZlwdoMm0_2(.din(w_dff_B_6U8373391_2),.dout(w_dff_B_RZlwdoMm0_2),.clk(gclk));
	jdff dff_B_vPvA7ghK4_2(.din(w_dff_B_RZlwdoMm0_2),.dout(w_dff_B_vPvA7ghK4_2),.clk(gclk));
	jdff dff_B_7wdXn7xq8_1(.din(n1598),.dout(w_dff_B_7wdXn7xq8_1),.clk(gclk));
	jdff dff_B_MBaxzcXn6_2(.din(n1540),.dout(w_dff_B_MBaxzcXn6_2),.clk(gclk));
	jdff dff_B_ffOzgL0A6_2(.din(w_dff_B_MBaxzcXn6_2),.dout(w_dff_B_ffOzgL0A6_2),.clk(gclk));
	jdff dff_B_DcaIJKdj8_2(.din(w_dff_B_ffOzgL0A6_2),.dout(w_dff_B_DcaIJKdj8_2),.clk(gclk));
	jdff dff_B_aKsbO9YB1_2(.din(w_dff_B_DcaIJKdj8_2),.dout(w_dff_B_aKsbO9YB1_2),.clk(gclk));
	jdff dff_B_vPkuSM7D9_2(.din(w_dff_B_aKsbO9YB1_2),.dout(w_dff_B_vPkuSM7D9_2),.clk(gclk));
	jdff dff_B_ri8K1K2j6_2(.din(w_dff_B_vPkuSM7D9_2),.dout(w_dff_B_ri8K1K2j6_2),.clk(gclk));
	jdff dff_B_NpVHOysA0_2(.din(w_dff_B_ri8K1K2j6_2),.dout(w_dff_B_NpVHOysA0_2),.clk(gclk));
	jdff dff_B_rEtLTi0k3_2(.din(w_dff_B_NpVHOysA0_2),.dout(w_dff_B_rEtLTi0k3_2),.clk(gclk));
	jdff dff_B_vZWYy1ZJ9_2(.din(w_dff_B_rEtLTi0k3_2),.dout(w_dff_B_vZWYy1ZJ9_2),.clk(gclk));
	jdff dff_B_TYm4E5dt4_2(.din(w_dff_B_vZWYy1ZJ9_2),.dout(w_dff_B_TYm4E5dt4_2),.clk(gclk));
	jdff dff_B_IITNda7D9_2(.din(w_dff_B_TYm4E5dt4_2),.dout(w_dff_B_IITNda7D9_2),.clk(gclk));
	jdff dff_B_aM3CxAwF5_2(.din(w_dff_B_IITNda7D9_2),.dout(w_dff_B_aM3CxAwF5_2),.clk(gclk));
	jdff dff_B_O6XAyyGO9_2(.din(w_dff_B_aM3CxAwF5_2),.dout(w_dff_B_O6XAyyGO9_2),.clk(gclk));
	jdff dff_B_yE6j8YpU0_2(.din(w_dff_B_O6XAyyGO9_2),.dout(w_dff_B_yE6j8YpU0_2),.clk(gclk));
	jdff dff_B_pmHyXNkc7_2(.din(w_dff_B_yE6j8YpU0_2),.dout(w_dff_B_pmHyXNkc7_2),.clk(gclk));
	jdff dff_B_jlVxlsF33_2(.din(w_dff_B_pmHyXNkc7_2),.dout(w_dff_B_jlVxlsF33_2),.clk(gclk));
	jdff dff_B_Pd09L2yh1_2(.din(w_dff_B_jlVxlsF33_2),.dout(w_dff_B_Pd09L2yh1_2),.clk(gclk));
	jdff dff_B_OPMTPTxp3_2(.din(w_dff_B_Pd09L2yh1_2),.dout(w_dff_B_OPMTPTxp3_2),.clk(gclk));
	jdff dff_B_IPZr3kO27_2(.din(w_dff_B_OPMTPTxp3_2),.dout(w_dff_B_IPZr3kO27_2),.clk(gclk));
	jdff dff_B_Yf6Wlj752_2(.din(w_dff_B_IPZr3kO27_2),.dout(w_dff_B_Yf6Wlj752_2),.clk(gclk));
	jdff dff_B_gdHjwZcI1_2(.din(w_dff_B_Yf6Wlj752_2),.dout(w_dff_B_gdHjwZcI1_2),.clk(gclk));
	jdff dff_B_2Vg8P0ca2_2(.din(w_dff_B_gdHjwZcI1_2),.dout(w_dff_B_2Vg8P0ca2_2),.clk(gclk));
	jdff dff_B_cI4J6ngt3_2(.din(w_dff_B_2Vg8P0ca2_2),.dout(w_dff_B_cI4J6ngt3_2),.clk(gclk));
	jdff dff_B_RNepMO3g6_2(.din(w_dff_B_cI4J6ngt3_2),.dout(w_dff_B_RNepMO3g6_2),.clk(gclk));
	jdff dff_B_qnbjfDLL2_2(.din(w_dff_B_RNepMO3g6_2),.dout(w_dff_B_qnbjfDLL2_2),.clk(gclk));
	jdff dff_B_vxXFrN1R4_2(.din(w_dff_B_qnbjfDLL2_2),.dout(w_dff_B_vxXFrN1R4_2),.clk(gclk));
	jdff dff_B_qGy1li6f4_2(.din(w_dff_B_vxXFrN1R4_2),.dout(w_dff_B_qGy1li6f4_2),.clk(gclk));
	jdff dff_B_ZD39w16C8_2(.din(w_dff_B_qGy1li6f4_2),.dout(w_dff_B_ZD39w16C8_2),.clk(gclk));
	jdff dff_B_1dRbeTai0_2(.din(w_dff_B_ZD39w16C8_2),.dout(w_dff_B_1dRbeTai0_2),.clk(gclk));
	jdff dff_B_sS4TXpeF5_2(.din(w_dff_B_1dRbeTai0_2),.dout(w_dff_B_sS4TXpeF5_2),.clk(gclk));
	jdff dff_B_w4QzL81w7_2(.din(w_dff_B_sS4TXpeF5_2),.dout(w_dff_B_w4QzL81w7_2),.clk(gclk));
	jdff dff_B_8mFOqBu00_2(.din(w_dff_B_w4QzL81w7_2),.dout(w_dff_B_8mFOqBu00_2),.clk(gclk));
	jdff dff_B_PEGDJIF03_2(.din(w_dff_B_8mFOqBu00_2),.dout(w_dff_B_PEGDJIF03_2),.clk(gclk));
	jdff dff_B_hzKbM6lj2_2(.din(w_dff_B_PEGDJIF03_2),.dout(w_dff_B_hzKbM6lj2_2),.clk(gclk));
	jdff dff_B_RKk958mT8_2(.din(w_dff_B_hzKbM6lj2_2),.dout(w_dff_B_RKk958mT8_2),.clk(gclk));
	jdff dff_B_cSgU2YQR8_2(.din(w_dff_B_RKk958mT8_2),.dout(w_dff_B_cSgU2YQR8_2),.clk(gclk));
	jdff dff_B_k67nTlFJ0_2(.din(w_dff_B_cSgU2YQR8_2),.dout(w_dff_B_k67nTlFJ0_2),.clk(gclk));
	jdff dff_B_j5ssqJ709_2(.din(w_dff_B_k67nTlFJ0_2),.dout(w_dff_B_j5ssqJ709_2),.clk(gclk));
	jdff dff_B_KBP1Yr8X1_2(.din(w_dff_B_j5ssqJ709_2),.dout(w_dff_B_KBP1Yr8X1_2),.clk(gclk));
	jdff dff_B_10j4VEk86_2(.din(w_dff_B_KBP1Yr8X1_2),.dout(w_dff_B_10j4VEk86_2),.clk(gclk));
	jdff dff_B_HCrwfOX29_2(.din(w_dff_B_10j4VEk86_2),.dout(w_dff_B_HCrwfOX29_2),.clk(gclk));
	jdff dff_B_W50Qyrbw6_2(.din(n1579),.dout(w_dff_B_W50Qyrbw6_2),.clk(gclk));
	jdff dff_B_rlviRy9l5_1(.din(n1541),.dout(w_dff_B_rlviRy9l5_1),.clk(gclk));
	jdff dff_B_tt85ceTp2_2(.din(n1476),.dout(w_dff_B_tt85ceTp2_2),.clk(gclk));
	jdff dff_B_YB6HQslk7_2(.din(w_dff_B_tt85ceTp2_2),.dout(w_dff_B_YB6HQslk7_2),.clk(gclk));
	jdff dff_B_UgTW4v2B1_2(.din(w_dff_B_YB6HQslk7_2),.dout(w_dff_B_UgTW4v2B1_2),.clk(gclk));
	jdff dff_B_9UWUFGRU4_2(.din(w_dff_B_UgTW4v2B1_2),.dout(w_dff_B_9UWUFGRU4_2),.clk(gclk));
	jdff dff_B_SP0FId8K8_2(.din(w_dff_B_9UWUFGRU4_2),.dout(w_dff_B_SP0FId8K8_2),.clk(gclk));
	jdff dff_B_ECITgqmX1_2(.din(w_dff_B_SP0FId8K8_2),.dout(w_dff_B_ECITgqmX1_2),.clk(gclk));
	jdff dff_B_pcVGBoLR6_2(.din(w_dff_B_ECITgqmX1_2),.dout(w_dff_B_pcVGBoLR6_2),.clk(gclk));
	jdff dff_B_T3niKc1M2_2(.din(w_dff_B_pcVGBoLR6_2),.dout(w_dff_B_T3niKc1M2_2),.clk(gclk));
	jdff dff_B_jX6oBj0i5_2(.din(w_dff_B_T3niKc1M2_2),.dout(w_dff_B_jX6oBj0i5_2),.clk(gclk));
	jdff dff_B_MvHgLRx49_2(.din(w_dff_B_jX6oBj0i5_2),.dout(w_dff_B_MvHgLRx49_2),.clk(gclk));
	jdff dff_B_VjrxxHLG7_2(.din(w_dff_B_MvHgLRx49_2),.dout(w_dff_B_VjrxxHLG7_2),.clk(gclk));
	jdff dff_B_b6P5lV8Y8_2(.din(w_dff_B_VjrxxHLG7_2),.dout(w_dff_B_b6P5lV8Y8_2),.clk(gclk));
	jdff dff_B_lo1Jo8NM4_2(.din(w_dff_B_b6P5lV8Y8_2),.dout(w_dff_B_lo1Jo8NM4_2),.clk(gclk));
	jdff dff_B_C7ztNqX31_2(.din(w_dff_B_lo1Jo8NM4_2),.dout(w_dff_B_C7ztNqX31_2),.clk(gclk));
	jdff dff_B_clW06KAT5_2(.din(w_dff_B_C7ztNqX31_2),.dout(w_dff_B_clW06KAT5_2),.clk(gclk));
	jdff dff_B_NCBxeYwQ8_2(.din(w_dff_B_clW06KAT5_2),.dout(w_dff_B_NCBxeYwQ8_2),.clk(gclk));
	jdff dff_B_PIUXLQ7r0_2(.din(w_dff_B_NCBxeYwQ8_2),.dout(w_dff_B_PIUXLQ7r0_2),.clk(gclk));
	jdff dff_B_c9Oqtcda7_2(.din(w_dff_B_PIUXLQ7r0_2),.dout(w_dff_B_c9Oqtcda7_2),.clk(gclk));
	jdff dff_B_fOv2905U6_2(.din(w_dff_B_c9Oqtcda7_2),.dout(w_dff_B_fOv2905U6_2),.clk(gclk));
	jdff dff_B_BWvCBIQi6_2(.din(w_dff_B_fOv2905U6_2),.dout(w_dff_B_BWvCBIQi6_2),.clk(gclk));
	jdff dff_B_uhwLdBhe2_2(.din(w_dff_B_BWvCBIQi6_2),.dout(w_dff_B_uhwLdBhe2_2),.clk(gclk));
	jdff dff_B_eQQ9BNKv2_2(.din(w_dff_B_uhwLdBhe2_2),.dout(w_dff_B_eQQ9BNKv2_2),.clk(gclk));
	jdff dff_B_HjkYvuQO4_2(.din(w_dff_B_eQQ9BNKv2_2),.dout(w_dff_B_HjkYvuQO4_2),.clk(gclk));
	jdff dff_B_TMtBTEPy5_2(.din(w_dff_B_HjkYvuQO4_2),.dout(w_dff_B_TMtBTEPy5_2),.clk(gclk));
	jdff dff_B_jZRa4nPc3_2(.din(w_dff_B_TMtBTEPy5_2),.dout(w_dff_B_jZRa4nPc3_2),.clk(gclk));
	jdff dff_B_ASirHnKY8_2(.din(w_dff_B_jZRa4nPc3_2),.dout(w_dff_B_ASirHnKY8_2),.clk(gclk));
	jdff dff_B_6SjSxr2G1_2(.din(w_dff_B_ASirHnKY8_2),.dout(w_dff_B_6SjSxr2G1_2),.clk(gclk));
	jdff dff_B_COsSvsm94_2(.din(w_dff_B_6SjSxr2G1_2),.dout(w_dff_B_COsSvsm94_2),.clk(gclk));
	jdff dff_B_AJBXZuQz9_2(.din(w_dff_B_COsSvsm94_2),.dout(w_dff_B_AJBXZuQz9_2),.clk(gclk));
	jdff dff_B_qQGAcyMx7_2(.din(w_dff_B_AJBXZuQz9_2),.dout(w_dff_B_qQGAcyMx7_2),.clk(gclk));
	jdff dff_B_v2AbIQqE3_2(.din(w_dff_B_qQGAcyMx7_2),.dout(w_dff_B_v2AbIQqE3_2),.clk(gclk));
	jdff dff_B_Ldk91WU46_2(.din(w_dff_B_v2AbIQqE3_2),.dout(w_dff_B_Ldk91WU46_2),.clk(gclk));
	jdff dff_B_A7d9UWtF9_2(.din(w_dff_B_Ldk91WU46_2),.dout(w_dff_B_A7d9UWtF9_2),.clk(gclk));
	jdff dff_B_rzsEWZXU3_2(.din(w_dff_B_A7d9UWtF9_2),.dout(w_dff_B_rzsEWZXU3_2),.clk(gclk));
	jdff dff_B_M07pNaUx9_2(.din(w_dff_B_rzsEWZXU3_2),.dout(w_dff_B_M07pNaUx9_2),.clk(gclk));
	jdff dff_B_nkLIFtgr7_2(.din(w_dff_B_M07pNaUx9_2),.dout(w_dff_B_nkLIFtgr7_2),.clk(gclk));
	jdff dff_B_jAmeWmgd8_2(.din(w_dff_B_nkLIFtgr7_2),.dout(w_dff_B_jAmeWmgd8_2),.clk(gclk));
	jdff dff_B_SlMs5Ypt1_2(.din(w_dff_B_jAmeWmgd8_2),.dout(w_dff_B_SlMs5Ypt1_2),.clk(gclk));
	jdff dff_B_EbZ9Y5HW1_2(.din(n1515),.dout(w_dff_B_EbZ9Y5HW1_2),.clk(gclk));
	jdff dff_B_O45oxs1m1_1(.din(n1477),.dout(w_dff_B_O45oxs1m1_1),.clk(gclk));
	jdff dff_B_GIt6yQGw5_2(.din(n1405),.dout(w_dff_B_GIt6yQGw5_2),.clk(gclk));
	jdff dff_B_uBdElKpA7_2(.din(w_dff_B_GIt6yQGw5_2),.dout(w_dff_B_uBdElKpA7_2),.clk(gclk));
	jdff dff_B_jglgimgk5_2(.din(w_dff_B_uBdElKpA7_2),.dout(w_dff_B_jglgimgk5_2),.clk(gclk));
	jdff dff_B_HNNBXJ0e3_2(.din(w_dff_B_jglgimgk5_2),.dout(w_dff_B_HNNBXJ0e3_2),.clk(gclk));
	jdff dff_B_EUv7Pd5x5_2(.din(w_dff_B_HNNBXJ0e3_2),.dout(w_dff_B_EUv7Pd5x5_2),.clk(gclk));
	jdff dff_B_atYAZREb3_2(.din(w_dff_B_EUv7Pd5x5_2),.dout(w_dff_B_atYAZREb3_2),.clk(gclk));
	jdff dff_B_OklQO3ti5_2(.din(w_dff_B_atYAZREb3_2),.dout(w_dff_B_OklQO3ti5_2),.clk(gclk));
	jdff dff_B_51586D049_2(.din(w_dff_B_OklQO3ti5_2),.dout(w_dff_B_51586D049_2),.clk(gclk));
	jdff dff_B_RX6Unpp46_2(.din(w_dff_B_51586D049_2),.dout(w_dff_B_RX6Unpp46_2),.clk(gclk));
	jdff dff_B_L6jxg9U82_2(.din(w_dff_B_RX6Unpp46_2),.dout(w_dff_B_L6jxg9U82_2),.clk(gclk));
	jdff dff_B_ZqpAp6zJ1_2(.din(w_dff_B_L6jxg9U82_2),.dout(w_dff_B_ZqpAp6zJ1_2),.clk(gclk));
	jdff dff_B_1YWDwpIV6_2(.din(w_dff_B_ZqpAp6zJ1_2),.dout(w_dff_B_1YWDwpIV6_2),.clk(gclk));
	jdff dff_B_zc2ww7O23_2(.din(w_dff_B_1YWDwpIV6_2),.dout(w_dff_B_zc2ww7O23_2),.clk(gclk));
	jdff dff_B_sf3Z0jfs3_2(.din(w_dff_B_zc2ww7O23_2),.dout(w_dff_B_sf3Z0jfs3_2),.clk(gclk));
	jdff dff_B_og8ipIzG0_2(.din(w_dff_B_sf3Z0jfs3_2),.dout(w_dff_B_og8ipIzG0_2),.clk(gclk));
	jdff dff_B_pbacs4S92_2(.din(w_dff_B_og8ipIzG0_2),.dout(w_dff_B_pbacs4S92_2),.clk(gclk));
	jdff dff_B_eQsyoHpB9_2(.din(w_dff_B_pbacs4S92_2),.dout(w_dff_B_eQsyoHpB9_2),.clk(gclk));
	jdff dff_B_copNBME19_2(.din(w_dff_B_eQsyoHpB9_2),.dout(w_dff_B_copNBME19_2),.clk(gclk));
	jdff dff_B_0U5qMBne2_2(.din(w_dff_B_copNBME19_2),.dout(w_dff_B_0U5qMBne2_2),.clk(gclk));
	jdff dff_B_hhX7s2Gr4_2(.din(w_dff_B_0U5qMBne2_2),.dout(w_dff_B_hhX7s2Gr4_2),.clk(gclk));
	jdff dff_B_dlyx0Y127_2(.din(w_dff_B_hhX7s2Gr4_2),.dout(w_dff_B_dlyx0Y127_2),.clk(gclk));
	jdff dff_B_Wh8mMQl34_2(.din(w_dff_B_dlyx0Y127_2),.dout(w_dff_B_Wh8mMQl34_2),.clk(gclk));
	jdff dff_B_pXcWmqzX7_2(.din(w_dff_B_Wh8mMQl34_2),.dout(w_dff_B_pXcWmqzX7_2),.clk(gclk));
	jdff dff_B_gj9jYQON2_2(.din(w_dff_B_pXcWmqzX7_2),.dout(w_dff_B_gj9jYQON2_2),.clk(gclk));
	jdff dff_B_MdM0X7Ni8_2(.din(w_dff_B_gj9jYQON2_2),.dout(w_dff_B_MdM0X7Ni8_2),.clk(gclk));
	jdff dff_B_xD3kKjUQ0_2(.din(w_dff_B_MdM0X7Ni8_2),.dout(w_dff_B_xD3kKjUQ0_2),.clk(gclk));
	jdff dff_B_8bU7kZIR7_2(.din(w_dff_B_xD3kKjUQ0_2),.dout(w_dff_B_8bU7kZIR7_2),.clk(gclk));
	jdff dff_B_B9dGR5wu0_2(.din(w_dff_B_8bU7kZIR7_2),.dout(w_dff_B_B9dGR5wu0_2),.clk(gclk));
	jdff dff_B_YVsFPeV26_2(.din(w_dff_B_B9dGR5wu0_2),.dout(w_dff_B_YVsFPeV26_2),.clk(gclk));
	jdff dff_B_BrYF22Up2_2(.din(w_dff_B_YVsFPeV26_2),.dout(w_dff_B_BrYF22Up2_2),.clk(gclk));
	jdff dff_B_s7WC25b94_2(.din(w_dff_B_BrYF22Up2_2),.dout(w_dff_B_s7WC25b94_2),.clk(gclk));
	jdff dff_B_1jKFPvBD8_2(.din(w_dff_B_s7WC25b94_2),.dout(w_dff_B_1jKFPvBD8_2),.clk(gclk));
	jdff dff_B_q5B90cfv0_2(.din(w_dff_B_1jKFPvBD8_2),.dout(w_dff_B_q5B90cfv0_2),.clk(gclk));
	jdff dff_B_WhphCp273_2(.din(w_dff_B_q5B90cfv0_2),.dout(w_dff_B_WhphCp273_2),.clk(gclk));
	jdff dff_B_aWErp4ZT3_2(.din(w_dff_B_WhphCp273_2),.dout(w_dff_B_aWErp4ZT3_2),.clk(gclk));
	jdff dff_B_T1ZHVrvU9_2(.din(n1444),.dout(w_dff_B_T1ZHVrvU9_2),.clk(gclk));
	jdff dff_B_Q0KMD2eo2_1(.din(n1406),.dout(w_dff_B_Q0KMD2eo2_1),.clk(gclk));
	jdff dff_B_3LotTdUk0_2(.din(n1327),.dout(w_dff_B_3LotTdUk0_2),.clk(gclk));
	jdff dff_B_9WChpInF5_2(.din(w_dff_B_3LotTdUk0_2),.dout(w_dff_B_9WChpInF5_2),.clk(gclk));
	jdff dff_B_Av3Ax3GG9_2(.din(w_dff_B_9WChpInF5_2),.dout(w_dff_B_Av3Ax3GG9_2),.clk(gclk));
	jdff dff_B_lAVYpExO7_2(.din(w_dff_B_Av3Ax3GG9_2),.dout(w_dff_B_lAVYpExO7_2),.clk(gclk));
	jdff dff_B_Skuahs6X6_2(.din(w_dff_B_lAVYpExO7_2),.dout(w_dff_B_Skuahs6X6_2),.clk(gclk));
	jdff dff_B_Kr0RdxBu4_2(.din(w_dff_B_Skuahs6X6_2),.dout(w_dff_B_Kr0RdxBu4_2),.clk(gclk));
	jdff dff_B_gRaHvrKl6_2(.din(w_dff_B_Kr0RdxBu4_2),.dout(w_dff_B_gRaHvrKl6_2),.clk(gclk));
	jdff dff_B_w5jyNEoj4_2(.din(w_dff_B_gRaHvrKl6_2),.dout(w_dff_B_w5jyNEoj4_2),.clk(gclk));
	jdff dff_B_zbx9B9IZ0_2(.din(w_dff_B_w5jyNEoj4_2),.dout(w_dff_B_zbx9B9IZ0_2),.clk(gclk));
	jdff dff_B_4iozQe248_2(.din(w_dff_B_zbx9B9IZ0_2),.dout(w_dff_B_4iozQe248_2),.clk(gclk));
	jdff dff_B_vAVO0Wtk5_2(.din(w_dff_B_4iozQe248_2),.dout(w_dff_B_vAVO0Wtk5_2),.clk(gclk));
	jdff dff_B_3VpJpqqL7_2(.din(w_dff_B_vAVO0Wtk5_2),.dout(w_dff_B_3VpJpqqL7_2),.clk(gclk));
	jdff dff_B_pqCD6kKb8_2(.din(w_dff_B_3VpJpqqL7_2),.dout(w_dff_B_pqCD6kKb8_2),.clk(gclk));
	jdff dff_B_Ovd3VDzZ0_2(.din(w_dff_B_pqCD6kKb8_2),.dout(w_dff_B_Ovd3VDzZ0_2),.clk(gclk));
	jdff dff_B_R7Vb8WBB4_2(.din(w_dff_B_Ovd3VDzZ0_2),.dout(w_dff_B_R7Vb8WBB4_2),.clk(gclk));
	jdff dff_B_Ui3t7buT2_2(.din(w_dff_B_R7Vb8WBB4_2),.dout(w_dff_B_Ui3t7buT2_2),.clk(gclk));
	jdff dff_B_CEydjoAt0_2(.din(w_dff_B_Ui3t7buT2_2),.dout(w_dff_B_CEydjoAt0_2),.clk(gclk));
	jdff dff_B_uAcEd9QB0_2(.din(w_dff_B_CEydjoAt0_2),.dout(w_dff_B_uAcEd9QB0_2),.clk(gclk));
	jdff dff_B_3Q7Hm6xA9_2(.din(w_dff_B_uAcEd9QB0_2),.dout(w_dff_B_3Q7Hm6xA9_2),.clk(gclk));
	jdff dff_B_P0KwbxrD7_2(.din(w_dff_B_3Q7Hm6xA9_2),.dout(w_dff_B_P0KwbxrD7_2),.clk(gclk));
	jdff dff_B_3dwfZuv69_2(.din(w_dff_B_P0KwbxrD7_2),.dout(w_dff_B_3dwfZuv69_2),.clk(gclk));
	jdff dff_B_KpchTjCI8_2(.din(w_dff_B_3dwfZuv69_2),.dout(w_dff_B_KpchTjCI8_2),.clk(gclk));
	jdff dff_B_zFYTX8CP8_2(.din(w_dff_B_KpchTjCI8_2),.dout(w_dff_B_zFYTX8CP8_2),.clk(gclk));
	jdff dff_B_vXMzPBv28_2(.din(w_dff_B_zFYTX8CP8_2),.dout(w_dff_B_vXMzPBv28_2),.clk(gclk));
	jdff dff_B_5DjJHNL86_2(.din(w_dff_B_vXMzPBv28_2),.dout(w_dff_B_5DjJHNL86_2),.clk(gclk));
	jdff dff_B_G2YbobsN1_2(.din(w_dff_B_5DjJHNL86_2),.dout(w_dff_B_G2YbobsN1_2),.clk(gclk));
	jdff dff_B_k7A2pZSS8_2(.din(w_dff_B_G2YbobsN1_2),.dout(w_dff_B_k7A2pZSS8_2),.clk(gclk));
	jdff dff_B_h7gOn26C1_2(.din(w_dff_B_k7A2pZSS8_2),.dout(w_dff_B_h7gOn26C1_2),.clk(gclk));
	jdff dff_B_5IOrGMpb5_2(.din(w_dff_B_h7gOn26C1_2),.dout(w_dff_B_5IOrGMpb5_2),.clk(gclk));
	jdff dff_B_mJyNMxgk5_2(.din(w_dff_B_5IOrGMpb5_2),.dout(w_dff_B_mJyNMxgk5_2),.clk(gclk));
	jdff dff_B_9E7EO7PV7_2(.din(w_dff_B_mJyNMxgk5_2),.dout(w_dff_B_9E7EO7PV7_2),.clk(gclk));
	jdff dff_B_zoqa3g5I7_2(.din(w_dff_B_9E7EO7PV7_2),.dout(w_dff_B_zoqa3g5I7_2),.clk(gclk));
	jdff dff_B_LXPE0yOq1_2(.din(n1366),.dout(w_dff_B_LXPE0yOq1_2),.clk(gclk));
	jdff dff_B_XsKObT771_1(.din(n1328),.dout(w_dff_B_XsKObT771_1),.clk(gclk));
	jdff dff_B_3FDkFYgy2_2(.din(n1242),.dout(w_dff_B_3FDkFYgy2_2),.clk(gclk));
	jdff dff_B_DfyloW6U1_2(.din(w_dff_B_3FDkFYgy2_2),.dout(w_dff_B_DfyloW6U1_2),.clk(gclk));
	jdff dff_B_WpmeYibs2_2(.din(w_dff_B_DfyloW6U1_2),.dout(w_dff_B_WpmeYibs2_2),.clk(gclk));
	jdff dff_B_ismQLkxc5_2(.din(w_dff_B_WpmeYibs2_2),.dout(w_dff_B_ismQLkxc5_2),.clk(gclk));
	jdff dff_B_f1dVwbxx3_2(.din(w_dff_B_ismQLkxc5_2),.dout(w_dff_B_f1dVwbxx3_2),.clk(gclk));
	jdff dff_B_riePBStL7_2(.din(w_dff_B_f1dVwbxx3_2),.dout(w_dff_B_riePBStL7_2),.clk(gclk));
	jdff dff_B_nOoUmHIE0_2(.din(w_dff_B_riePBStL7_2),.dout(w_dff_B_nOoUmHIE0_2),.clk(gclk));
	jdff dff_B_VIEZRoua3_2(.din(w_dff_B_nOoUmHIE0_2),.dout(w_dff_B_VIEZRoua3_2),.clk(gclk));
	jdff dff_B_A6ZGEqzY7_2(.din(w_dff_B_VIEZRoua3_2),.dout(w_dff_B_A6ZGEqzY7_2),.clk(gclk));
	jdff dff_B_lsQDhDfG6_2(.din(w_dff_B_A6ZGEqzY7_2),.dout(w_dff_B_lsQDhDfG6_2),.clk(gclk));
	jdff dff_B_QPmYOZp32_2(.din(w_dff_B_lsQDhDfG6_2),.dout(w_dff_B_QPmYOZp32_2),.clk(gclk));
	jdff dff_B_dfgWMsG67_2(.din(w_dff_B_QPmYOZp32_2),.dout(w_dff_B_dfgWMsG67_2),.clk(gclk));
	jdff dff_B_Oze0BHgY1_2(.din(w_dff_B_dfgWMsG67_2),.dout(w_dff_B_Oze0BHgY1_2),.clk(gclk));
	jdff dff_B_sf5P6DNl2_2(.din(w_dff_B_Oze0BHgY1_2),.dout(w_dff_B_sf5P6DNl2_2),.clk(gclk));
	jdff dff_B_mjhS1ujV9_2(.din(w_dff_B_sf5P6DNl2_2),.dout(w_dff_B_mjhS1ujV9_2),.clk(gclk));
	jdff dff_B_Tz9mdE135_2(.din(w_dff_B_mjhS1ujV9_2),.dout(w_dff_B_Tz9mdE135_2),.clk(gclk));
	jdff dff_B_qKmbLJQm9_2(.din(w_dff_B_Tz9mdE135_2),.dout(w_dff_B_qKmbLJQm9_2),.clk(gclk));
	jdff dff_B_17SqajER6_2(.din(w_dff_B_qKmbLJQm9_2),.dout(w_dff_B_17SqajER6_2),.clk(gclk));
	jdff dff_B_zTJ0d35B7_2(.din(w_dff_B_17SqajER6_2),.dout(w_dff_B_zTJ0d35B7_2),.clk(gclk));
	jdff dff_B_tIJncfAq5_2(.din(w_dff_B_zTJ0d35B7_2),.dout(w_dff_B_tIJncfAq5_2),.clk(gclk));
	jdff dff_B_9bg9qoa78_2(.din(w_dff_B_tIJncfAq5_2),.dout(w_dff_B_9bg9qoa78_2),.clk(gclk));
	jdff dff_B_qjZ2xRDk3_2(.din(w_dff_B_9bg9qoa78_2),.dout(w_dff_B_qjZ2xRDk3_2),.clk(gclk));
	jdff dff_B_T2f1wlHB5_2(.din(w_dff_B_qjZ2xRDk3_2),.dout(w_dff_B_T2f1wlHB5_2),.clk(gclk));
	jdff dff_B_TQ6uh5ey7_2(.din(w_dff_B_T2f1wlHB5_2),.dout(w_dff_B_TQ6uh5ey7_2),.clk(gclk));
	jdff dff_B_e7uPHoos3_2(.din(w_dff_B_TQ6uh5ey7_2),.dout(w_dff_B_e7uPHoos3_2),.clk(gclk));
	jdff dff_B_JB68xpvG4_2(.din(w_dff_B_e7uPHoos3_2),.dout(w_dff_B_JB68xpvG4_2),.clk(gclk));
	jdff dff_B_kH36B8Jr4_2(.din(w_dff_B_JB68xpvG4_2),.dout(w_dff_B_kH36B8Jr4_2),.clk(gclk));
	jdff dff_B_cb5Lomwy8_2(.din(w_dff_B_kH36B8Jr4_2),.dout(w_dff_B_cb5Lomwy8_2),.clk(gclk));
	jdff dff_B_IVyUdDth9_2(.din(w_dff_B_cb5Lomwy8_2),.dout(w_dff_B_IVyUdDth9_2),.clk(gclk));
	jdff dff_B_4unbKKyv2_2(.din(n1281),.dout(w_dff_B_4unbKKyv2_2),.clk(gclk));
	jdff dff_B_NTV0JpaY7_1(.din(n1243),.dout(w_dff_B_NTV0JpaY7_1),.clk(gclk));
	jdff dff_B_M6MPbOP08_2(.din(n1151),.dout(w_dff_B_M6MPbOP08_2),.clk(gclk));
	jdff dff_B_HWIc7Vvh2_2(.din(w_dff_B_M6MPbOP08_2),.dout(w_dff_B_HWIc7Vvh2_2),.clk(gclk));
	jdff dff_B_X7ICUWdi5_2(.din(w_dff_B_HWIc7Vvh2_2),.dout(w_dff_B_X7ICUWdi5_2),.clk(gclk));
	jdff dff_B_Us4ZMLs32_2(.din(w_dff_B_X7ICUWdi5_2),.dout(w_dff_B_Us4ZMLs32_2),.clk(gclk));
	jdff dff_B_EcnpEkef0_2(.din(w_dff_B_Us4ZMLs32_2),.dout(w_dff_B_EcnpEkef0_2),.clk(gclk));
	jdff dff_B_usBG6r4L1_2(.din(w_dff_B_EcnpEkef0_2),.dout(w_dff_B_usBG6r4L1_2),.clk(gclk));
	jdff dff_B_qNQGmkJw9_2(.din(w_dff_B_usBG6r4L1_2),.dout(w_dff_B_qNQGmkJw9_2),.clk(gclk));
	jdff dff_B_9E3q66NZ5_2(.din(w_dff_B_qNQGmkJw9_2),.dout(w_dff_B_9E3q66NZ5_2),.clk(gclk));
	jdff dff_B_wcSI2O9w3_2(.din(w_dff_B_9E3q66NZ5_2),.dout(w_dff_B_wcSI2O9w3_2),.clk(gclk));
	jdff dff_B_GBrbiIcZ4_2(.din(w_dff_B_wcSI2O9w3_2),.dout(w_dff_B_GBrbiIcZ4_2),.clk(gclk));
	jdff dff_B_8UoTzZZQ5_2(.din(w_dff_B_GBrbiIcZ4_2),.dout(w_dff_B_8UoTzZZQ5_2),.clk(gclk));
	jdff dff_B_lng2jslR6_2(.din(w_dff_B_8UoTzZZQ5_2),.dout(w_dff_B_lng2jslR6_2),.clk(gclk));
	jdff dff_B_ohyiPMzs1_2(.din(w_dff_B_lng2jslR6_2),.dout(w_dff_B_ohyiPMzs1_2),.clk(gclk));
	jdff dff_B_GcfzvsZZ4_2(.din(w_dff_B_ohyiPMzs1_2),.dout(w_dff_B_GcfzvsZZ4_2),.clk(gclk));
	jdff dff_B_qyo95S2A8_2(.din(w_dff_B_GcfzvsZZ4_2),.dout(w_dff_B_qyo95S2A8_2),.clk(gclk));
	jdff dff_B_xWGnhoyp6_2(.din(w_dff_B_qyo95S2A8_2),.dout(w_dff_B_xWGnhoyp6_2),.clk(gclk));
	jdff dff_B_xLVuIwOM2_2(.din(w_dff_B_xWGnhoyp6_2),.dout(w_dff_B_xLVuIwOM2_2),.clk(gclk));
	jdff dff_B_ABRvO3Gm6_2(.din(w_dff_B_xLVuIwOM2_2),.dout(w_dff_B_ABRvO3Gm6_2),.clk(gclk));
	jdff dff_B_f2NoFdnG4_2(.din(w_dff_B_ABRvO3Gm6_2),.dout(w_dff_B_f2NoFdnG4_2),.clk(gclk));
	jdff dff_B_F5XSCjvi4_2(.din(w_dff_B_f2NoFdnG4_2),.dout(w_dff_B_F5XSCjvi4_2),.clk(gclk));
	jdff dff_B_r5HJCcq01_2(.din(w_dff_B_F5XSCjvi4_2),.dout(w_dff_B_r5HJCcq01_2),.clk(gclk));
	jdff dff_B_bR87hDVs3_2(.din(w_dff_B_r5HJCcq01_2),.dout(w_dff_B_bR87hDVs3_2),.clk(gclk));
	jdff dff_B_PdAB4Kf17_2(.din(w_dff_B_bR87hDVs3_2),.dout(w_dff_B_PdAB4Kf17_2),.clk(gclk));
	jdff dff_B_5vVkkgl53_2(.din(w_dff_B_PdAB4Kf17_2),.dout(w_dff_B_5vVkkgl53_2),.clk(gclk));
	jdff dff_B_PKyCj2292_2(.din(w_dff_B_5vVkkgl53_2),.dout(w_dff_B_PKyCj2292_2),.clk(gclk));
	jdff dff_B_DANe89Pc6_2(.din(w_dff_B_PKyCj2292_2),.dout(w_dff_B_DANe89Pc6_2),.clk(gclk));
	jdff dff_B_LVaaCOzx9_2(.din(n1190),.dout(w_dff_B_LVaaCOzx9_2),.clk(gclk));
	jdff dff_B_6LIhDnGg7_1(.din(n1152),.dout(w_dff_B_6LIhDnGg7_1),.clk(gclk));
	jdff dff_B_WoIHbr2B5_2(.din(n1053),.dout(w_dff_B_WoIHbr2B5_2),.clk(gclk));
	jdff dff_B_AAN7k6AH0_2(.din(w_dff_B_WoIHbr2B5_2),.dout(w_dff_B_AAN7k6AH0_2),.clk(gclk));
	jdff dff_B_V6xVXnqP7_2(.din(w_dff_B_AAN7k6AH0_2),.dout(w_dff_B_V6xVXnqP7_2),.clk(gclk));
	jdff dff_B_IIkvho6D4_2(.din(w_dff_B_V6xVXnqP7_2),.dout(w_dff_B_IIkvho6D4_2),.clk(gclk));
	jdff dff_B_Z9Z0fINg8_2(.din(w_dff_B_IIkvho6D4_2),.dout(w_dff_B_Z9Z0fINg8_2),.clk(gclk));
	jdff dff_B_1l5vlHV07_2(.din(w_dff_B_Z9Z0fINg8_2),.dout(w_dff_B_1l5vlHV07_2),.clk(gclk));
	jdff dff_B_4waNQHrE1_2(.din(w_dff_B_1l5vlHV07_2),.dout(w_dff_B_4waNQHrE1_2),.clk(gclk));
	jdff dff_B_xdniJO7t6_2(.din(w_dff_B_4waNQHrE1_2),.dout(w_dff_B_xdniJO7t6_2),.clk(gclk));
	jdff dff_B_N6wYs5GC1_2(.din(w_dff_B_xdniJO7t6_2),.dout(w_dff_B_N6wYs5GC1_2),.clk(gclk));
	jdff dff_B_GStbbVmn4_2(.din(w_dff_B_N6wYs5GC1_2),.dout(w_dff_B_GStbbVmn4_2),.clk(gclk));
	jdff dff_B_0nNUjlrC5_2(.din(w_dff_B_GStbbVmn4_2),.dout(w_dff_B_0nNUjlrC5_2),.clk(gclk));
	jdff dff_B_uPr6GIUR6_2(.din(w_dff_B_0nNUjlrC5_2),.dout(w_dff_B_uPr6GIUR6_2),.clk(gclk));
	jdff dff_B_6q25G7C74_2(.din(w_dff_B_uPr6GIUR6_2),.dout(w_dff_B_6q25G7C74_2),.clk(gclk));
	jdff dff_B_ukJulgJa1_2(.din(w_dff_B_6q25G7C74_2),.dout(w_dff_B_ukJulgJa1_2),.clk(gclk));
	jdff dff_B_yjmTH8IW6_2(.din(w_dff_B_ukJulgJa1_2),.dout(w_dff_B_yjmTH8IW6_2),.clk(gclk));
	jdff dff_B_PQGRwwi04_2(.din(w_dff_B_yjmTH8IW6_2),.dout(w_dff_B_PQGRwwi04_2),.clk(gclk));
	jdff dff_B_4rcKrpCa9_2(.din(w_dff_B_PQGRwwi04_2),.dout(w_dff_B_4rcKrpCa9_2),.clk(gclk));
	jdff dff_B_GT3BDYVb2_2(.din(w_dff_B_4rcKrpCa9_2),.dout(w_dff_B_GT3BDYVb2_2),.clk(gclk));
	jdff dff_B_S6rGuAbY3_2(.din(w_dff_B_GT3BDYVb2_2),.dout(w_dff_B_S6rGuAbY3_2),.clk(gclk));
	jdff dff_B_GahVn0W57_2(.din(w_dff_B_S6rGuAbY3_2),.dout(w_dff_B_GahVn0W57_2),.clk(gclk));
	jdff dff_B_ln64X7KU1_2(.din(w_dff_B_GahVn0W57_2),.dout(w_dff_B_ln64X7KU1_2),.clk(gclk));
	jdff dff_B_sMPMIBpe6_2(.din(w_dff_B_ln64X7KU1_2),.dout(w_dff_B_sMPMIBpe6_2),.clk(gclk));
	jdff dff_B_M6F2BNcO5_2(.din(w_dff_B_sMPMIBpe6_2),.dout(w_dff_B_M6F2BNcO5_2),.clk(gclk));
	jdff dff_B_oht5QqZp1_2(.din(n1091),.dout(w_dff_B_oht5QqZp1_2),.clk(gclk));
	jdff dff_B_pX2KoYxw6_1(.din(n1054),.dout(w_dff_B_pX2KoYxw6_1),.clk(gclk));
	jdff dff_B_0uFWQ1TT9_2(.din(n954),.dout(w_dff_B_0uFWQ1TT9_2),.clk(gclk));
	jdff dff_B_jYMCYAoZ6_2(.din(w_dff_B_0uFWQ1TT9_2),.dout(w_dff_B_jYMCYAoZ6_2),.clk(gclk));
	jdff dff_B_lYYjqGL49_2(.din(w_dff_B_jYMCYAoZ6_2),.dout(w_dff_B_lYYjqGL49_2),.clk(gclk));
	jdff dff_B_Xoy6NoAW4_2(.din(w_dff_B_lYYjqGL49_2),.dout(w_dff_B_Xoy6NoAW4_2),.clk(gclk));
	jdff dff_B_IglZLohJ1_2(.din(w_dff_B_Xoy6NoAW4_2),.dout(w_dff_B_IglZLohJ1_2),.clk(gclk));
	jdff dff_B_6k9HpCEw6_2(.din(w_dff_B_IglZLohJ1_2),.dout(w_dff_B_6k9HpCEw6_2),.clk(gclk));
	jdff dff_B_nw8Ev4eU7_2(.din(w_dff_B_6k9HpCEw6_2),.dout(w_dff_B_nw8Ev4eU7_2),.clk(gclk));
	jdff dff_B_SlTpcpa97_2(.din(w_dff_B_nw8Ev4eU7_2),.dout(w_dff_B_SlTpcpa97_2),.clk(gclk));
	jdff dff_B_ZVNo4dll0_2(.din(w_dff_B_SlTpcpa97_2),.dout(w_dff_B_ZVNo4dll0_2),.clk(gclk));
	jdff dff_B_K7ZoG8473_2(.din(w_dff_B_ZVNo4dll0_2),.dout(w_dff_B_K7ZoG8473_2),.clk(gclk));
	jdff dff_B_bPzABTjK8_2(.din(w_dff_B_K7ZoG8473_2),.dout(w_dff_B_bPzABTjK8_2),.clk(gclk));
	jdff dff_B_ElpGkCPY9_2(.din(w_dff_B_bPzABTjK8_2),.dout(w_dff_B_ElpGkCPY9_2),.clk(gclk));
	jdff dff_B_GK7pGRUK9_2(.din(w_dff_B_ElpGkCPY9_2),.dout(w_dff_B_GK7pGRUK9_2),.clk(gclk));
	jdff dff_B_LzD6n1ah9_2(.din(w_dff_B_GK7pGRUK9_2),.dout(w_dff_B_LzD6n1ah9_2),.clk(gclk));
	jdff dff_B_ue5rVFnc3_2(.din(w_dff_B_LzD6n1ah9_2),.dout(w_dff_B_ue5rVFnc3_2),.clk(gclk));
	jdff dff_B_D36rVPAI6_2(.din(w_dff_B_ue5rVFnc3_2),.dout(w_dff_B_D36rVPAI6_2),.clk(gclk));
	jdff dff_B_b9G913cz9_2(.din(w_dff_B_D36rVPAI6_2),.dout(w_dff_B_b9G913cz9_2),.clk(gclk));
	jdff dff_B_G7vm2dvU1_2(.din(w_dff_B_b9G913cz9_2),.dout(w_dff_B_G7vm2dvU1_2),.clk(gclk));
	jdff dff_B_Fl7mkeel8_2(.din(w_dff_B_G7vm2dvU1_2),.dout(w_dff_B_Fl7mkeel8_2),.clk(gclk));
	jdff dff_B_rYhzUowM4_2(.din(w_dff_B_Fl7mkeel8_2),.dout(w_dff_B_rYhzUowM4_2),.clk(gclk));
	jdff dff_B_yMyjy5lP9_2(.din(n992),.dout(w_dff_B_yMyjy5lP9_2),.clk(gclk));
	jdff dff_B_TQIgVv3D2_1(.din(n955),.dout(w_dff_B_TQIgVv3D2_1),.clk(gclk));
	jdff dff_B_xKUoSrrP4_2(.din(n852),.dout(w_dff_B_xKUoSrrP4_2),.clk(gclk));
	jdff dff_B_nD9pGQkj7_2(.din(w_dff_B_xKUoSrrP4_2),.dout(w_dff_B_nD9pGQkj7_2),.clk(gclk));
	jdff dff_B_9DyghPPn3_2(.din(w_dff_B_nD9pGQkj7_2),.dout(w_dff_B_9DyghPPn3_2),.clk(gclk));
	jdff dff_B_72R75wz33_2(.din(w_dff_B_9DyghPPn3_2),.dout(w_dff_B_72R75wz33_2),.clk(gclk));
	jdff dff_B_LQfYXBSY0_2(.din(w_dff_B_72R75wz33_2),.dout(w_dff_B_LQfYXBSY0_2),.clk(gclk));
	jdff dff_B_LbFfgrF16_2(.din(w_dff_B_LQfYXBSY0_2),.dout(w_dff_B_LbFfgrF16_2),.clk(gclk));
	jdff dff_B_rLCUsHLf5_2(.din(w_dff_B_LbFfgrF16_2),.dout(w_dff_B_rLCUsHLf5_2),.clk(gclk));
	jdff dff_B_qyl61W6T4_2(.din(w_dff_B_rLCUsHLf5_2),.dout(w_dff_B_qyl61W6T4_2),.clk(gclk));
	jdff dff_B_sFZEMTdJ3_2(.din(w_dff_B_qyl61W6T4_2),.dout(w_dff_B_sFZEMTdJ3_2),.clk(gclk));
	jdff dff_B_cZmosjrc7_2(.din(w_dff_B_sFZEMTdJ3_2),.dout(w_dff_B_cZmosjrc7_2),.clk(gclk));
	jdff dff_B_ROpFQ6wA0_2(.din(w_dff_B_cZmosjrc7_2),.dout(w_dff_B_ROpFQ6wA0_2),.clk(gclk));
	jdff dff_B_pF6zIYni9_2(.din(w_dff_B_ROpFQ6wA0_2),.dout(w_dff_B_pF6zIYni9_2),.clk(gclk));
	jdff dff_B_nnhxoa7W2_2(.din(w_dff_B_pF6zIYni9_2),.dout(w_dff_B_nnhxoa7W2_2),.clk(gclk));
	jdff dff_B_AyeUgQ4M0_2(.din(w_dff_B_nnhxoa7W2_2),.dout(w_dff_B_AyeUgQ4M0_2),.clk(gclk));
	jdff dff_B_SFfitdX00_2(.din(w_dff_B_AyeUgQ4M0_2),.dout(w_dff_B_SFfitdX00_2),.clk(gclk));
	jdff dff_B_OOSPB0R73_2(.din(w_dff_B_SFfitdX00_2),.dout(w_dff_B_OOSPB0R73_2),.clk(gclk));
	jdff dff_B_lOI0ErTq6_2(.din(w_dff_B_OOSPB0R73_2),.dout(w_dff_B_lOI0ErTq6_2),.clk(gclk));
	jdff dff_B_e8521bL50_2(.din(n886),.dout(w_dff_B_e8521bL50_2),.clk(gclk));
	jdff dff_B_CqXK098R2_1(.din(n853),.dout(w_dff_B_CqXK098R2_1),.clk(gclk));
	jdff dff_B_CPKbHixs6_2(.din(n754),.dout(w_dff_B_CPKbHixs6_2),.clk(gclk));
	jdff dff_B_KODDDt5q0_2(.din(w_dff_B_CPKbHixs6_2),.dout(w_dff_B_KODDDt5q0_2),.clk(gclk));
	jdff dff_B_6PvG91yQ0_2(.din(w_dff_B_KODDDt5q0_2),.dout(w_dff_B_6PvG91yQ0_2),.clk(gclk));
	jdff dff_B_woOb5ry74_2(.din(w_dff_B_6PvG91yQ0_2),.dout(w_dff_B_woOb5ry74_2),.clk(gclk));
	jdff dff_B_XY5MEbzx4_2(.din(w_dff_B_woOb5ry74_2),.dout(w_dff_B_XY5MEbzx4_2),.clk(gclk));
	jdff dff_B_2fCRdRov6_2(.din(w_dff_B_XY5MEbzx4_2),.dout(w_dff_B_2fCRdRov6_2),.clk(gclk));
	jdff dff_B_Eg2j2r7n0_2(.din(w_dff_B_2fCRdRov6_2),.dout(w_dff_B_Eg2j2r7n0_2),.clk(gclk));
	jdff dff_B_J39YEIGX9_2(.din(w_dff_B_Eg2j2r7n0_2),.dout(w_dff_B_J39YEIGX9_2),.clk(gclk));
	jdff dff_B_AiEjmKEm2_2(.din(w_dff_B_J39YEIGX9_2),.dout(w_dff_B_AiEjmKEm2_2),.clk(gclk));
	jdff dff_B_NGJH8CNT2_2(.din(w_dff_B_AiEjmKEm2_2),.dout(w_dff_B_NGJH8CNT2_2),.clk(gclk));
	jdff dff_B_aY6f32F14_2(.din(w_dff_B_NGJH8CNT2_2),.dout(w_dff_B_aY6f32F14_2),.clk(gclk));
	jdff dff_B_WTtcbrbp0_2(.din(w_dff_B_aY6f32F14_2),.dout(w_dff_B_WTtcbrbp0_2),.clk(gclk));
	jdff dff_B_Xto36zXd3_2(.din(w_dff_B_WTtcbrbp0_2),.dout(w_dff_B_Xto36zXd3_2),.clk(gclk));
	jdff dff_B_6HXXvmvm1_2(.din(w_dff_B_Xto36zXd3_2),.dout(w_dff_B_6HXXvmvm1_2),.clk(gclk));
	jdff dff_B_v1rhBZ8R9_2(.din(n783),.dout(w_dff_B_v1rhBZ8R9_2),.clk(gclk));
	jdff dff_B_5jrER1x16_1(.din(n755),.dout(w_dff_B_5jrER1x16_1),.clk(gclk));
	jdff dff_B_2AYq0Bwy9_2(.din(n662),.dout(w_dff_B_2AYq0Bwy9_2),.clk(gclk));
	jdff dff_B_H6BudrGj4_2(.din(w_dff_B_2AYq0Bwy9_2),.dout(w_dff_B_H6BudrGj4_2),.clk(gclk));
	jdff dff_B_3e6kCOJq3_2(.din(w_dff_B_H6BudrGj4_2),.dout(w_dff_B_3e6kCOJq3_2),.clk(gclk));
	jdff dff_B_LUx15ufz7_2(.din(w_dff_B_3e6kCOJq3_2),.dout(w_dff_B_LUx15ufz7_2),.clk(gclk));
	jdff dff_B_crrRVYAr6_2(.din(w_dff_B_LUx15ufz7_2),.dout(w_dff_B_crrRVYAr6_2),.clk(gclk));
	jdff dff_B_Y6t5K9Je2_2(.din(w_dff_B_crrRVYAr6_2),.dout(w_dff_B_Y6t5K9Je2_2),.clk(gclk));
	jdff dff_B_trGqSKB23_2(.din(w_dff_B_Y6t5K9Je2_2),.dout(w_dff_B_trGqSKB23_2),.clk(gclk));
	jdff dff_B_9YpyBDd83_2(.din(w_dff_B_trGqSKB23_2),.dout(w_dff_B_9YpyBDd83_2),.clk(gclk));
	jdff dff_B_uzlyiqiE0_2(.din(w_dff_B_9YpyBDd83_2),.dout(w_dff_B_uzlyiqiE0_2),.clk(gclk));
	jdff dff_B_g63P4pV44_2(.din(w_dff_B_uzlyiqiE0_2),.dout(w_dff_B_g63P4pV44_2),.clk(gclk));
	jdff dff_B_yvjjMG5t8_2(.din(w_dff_B_g63P4pV44_2),.dout(w_dff_B_yvjjMG5t8_2),.clk(gclk));
	jdff dff_B_ntkPcTrO9_2(.din(n684),.dout(w_dff_B_ntkPcTrO9_2),.clk(gclk));
	jdff dff_B_TtpsuMRV5_1(.din(n663),.dout(w_dff_B_TtpsuMRV5_1),.clk(gclk));
	jdff dff_B_gRzaeMXP6_2(.din(n577),.dout(w_dff_B_gRzaeMXP6_2),.clk(gclk));
	jdff dff_B_Jytmd6hd1_2(.din(w_dff_B_gRzaeMXP6_2),.dout(w_dff_B_Jytmd6hd1_2),.clk(gclk));
	jdff dff_B_wgGQbVtJ3_2(.din(w_dff_B_Jytmd6hd1_2),.dout(w_dff_B_wgGQbVtJ3_2),.clk(gclk));
	jdff dff_B_hwJsTtd18_2(.din(w_dff_B_wgGQbVtJ3_2),.dout(w_dff_B_hwJsTtd18_2),.clk(gclk));
	jdff dff_B_B9F1MYl50_2(.din(w_dff_B_hwJsTtd18_2),.dout(w_dff_B_B9F1MYl50_2),.clk(gclk));
	jdff dff_B_rdo5XgCz3_2(.din(w_dff_B_B9F1MYl50_2),.dout(w_dff_B_rdo5XgCz3_2),.clk(gclk));
	jdff dff_B_IVmnjhSB0_2(.din(w_dff_B_rdo5XgCz3_2),.dout(w_dff_B_IVmnjhSB0_2),.clk(gclk));
	jdff dff_B_okQQNJjO8_2(.din(w_dff_B_IVmnjhSB0_2),.dout(w_dff_B_okQQNJjO8_2),.clk(gclk));
	jdff dff_B_XyMDSPbS9_2(.din(n592),.dout(w_dff_B_XyMDSPbS9_2),.clk(gclk));
	jdff dff_B_Hm4uXY3R1_2(.din(w_dff_B_XyMDSPbS9_2),.dout(w_dff_B_Hm4uXY3R1_2),.clk(gclk));
	jdff dff_B_rD2axpKL5_2(.din(w_dff_B_Hm4uXY3R1_2),.dout(w_dff_B_rD2axpKL5_2),.clk(gclk));
	jdff dff_B_xfeIIpLG8_1(.din(n578),.dout(w_dff_B_xfeIIpLG8_1),.clk(gclk));
	jdff dff_B_vue9wlNq3_1(.din(w_dff_B_xfeIIpLG8_1),.dout(w_dff_B_vue9wlNq3_1),.clk(gclk));
	jdff dff_B_8Z4UK4ht2_2(.din(n501),.dout(w_dff_B_8Z4UK4ht2_2),.clk(gclk));
	jdff dff_B_o3kYMXiw6_2(.din(w_dff_B_8Z4UK4ht2_2),.dout(w_dff_B_o3kYMXiw6_2),.clk(gclk));
	jdff dff_B_a9yMZg6v9_2(.din(w_dff_B_o3kYMXiw6_2),.dout(w_dff_B_a9yMZg6v9_2),.clk(gclk));
	jdff dff_B_bGahM8op0_0(.din(n506),.dout(w_dff_B_bGahM8op0_0),.clk(gclk));
	jdff dff_A_dA4xiOw58_0(.dout(w_n427_0[0]),.din(w_dff_A_dA4xiOw58_0),.clk(gclk));
	jdff dff_A_pOvWQzFu1_0(.dout(w_dff_A_dA4xiOw58_0),.din(w_dff_A_pOvWQzFu1_0),.clk(gclk));
	jdff dff_A_2yDzPjus9_1(.dout(w_n427_0[1]),.din(w_dff_A_2yDzPjus9_1),.clk(gclk));
	jdff dff_A_KrIQk1Yq0_1(.dout(w_dff_A_2yDzPjus9_1),.din(w_dff_A_KrIQk1Yq0_1),.clk(gclk));
	jdff dff_B_21KCN8U59_1(.din(n1729),.dout(w_dff_B_21KCN8U59_1),.clk(gclk));
	jdff dff_A_FN7R7Wuv2_1(.dout(w_n1697_0[1]),.din(w_dff_A_FN7R7Wuv2_1),.clk(gclk));
	jdff dff_B_l9V517vC0_1(.din(n1695),.dout(w_dff_B_l9V517vC0_1),.clk(gclk));
	jdff dff_B_kDMst8ru0_2(.din(n1653),.dout(w_dff_B_kDMst8ru0_2),.clk(gclk));
	jdff dff_B_IswEgwWA0_2(.din(w_dff_B_kDMst8ru0_2),.dout(w_dff_B_IswEgwWA0_2),.clk(gclk));
	jdff dff_B_O5n8xANB5_2(.din(w_dff_B_IswEgwWA0_2),.dout(w_dff_B_O5n8xANB5_2),.clk(gclk));
	jdff dff_B_r5E6ob3k8_2(.din(w_dff_B_O5n8xANB5_2),.dout(w_dff_B_r5E6ob3k8_2),.clk(gclk));
	jdff dff_B_Ra1N4xg39_2(.din(w_dff_B_r5E6ob3k8_2),.dout(w_dff_B_Ra1N4xg39_2),.clk(gclk));
	jdff dff_B_GVEJimHn8_2(.din(w_dff_B_Ra1N4xg39_2),.dout(w_dff_B_GVEJimHn8_2),.clk(gclk));
	jdff dff_B_vIy9m4ZJ4_2(.din(w_dff_B_GVEJimHn8_2),.dout(w_dff_B_vIy9m4ZJ4_2),.clk(gclk));
	jdff dff_B_bLhTxWf84_2(.din(w_dff_B_vIy9m4ZJ4_2),.dout(w_dff_B_bLhTxWf84_2),.clk(gclk));
	jdff dff_B_TSGgaxC88_2(.din(w_dff_B_bLhTxWf84_2),.dout(w_dff_B_TSGgaxC88_2),.clk(gclk));
	jdff dff_B_O6AoPGDW7_2(.din(w_dff_B_TSGgaxC88_2),.dout(w_dff_B_O6AoPGDW7_2),.clk(gclk));
	jdff dff_B_CyTUg9zY4_2(.din(w_dff_B_O6AoPGDW7_2),.dout(w_dff_B_CyTUg9zY4_2),.clk(gclk));
	jdff dff_B_R9hX5szf3_2(.din(w_dff_B_CyTUg9zY4_2),.dout(w_dff_B_R9hX5szf3_2),.clk(gclk));
	jdff dff_B_4NvmlHSU1_2(.din(w_dff_B_R9hX5szf3_2),.dout(w_dff_B_4NvmlHSU1_2),.clk(gclk));
	jdff dff_B_zLOVYjFV0_2(.din(w_dff_B_4NvmlHSU1_2),.dout(w_dff_B_zLOVYjFV0_2),.clk(gclk));
	jdff dff_B_Qw0EP8G27_2(.din(w_dff_B_zLOVYjFV0_2),.dout(w_dff_B_Qw0EP8G27_2),.clk(gclk));
	jdff dff_B_pG6bqBe88_2(.din(w_dff_B_Qw0EP8G27_2),.dout(w_dff_B_pG6bqBe88_2),.clk(gclk));
	jdff dff_B_wHzXodWt3_2(.din(w_dff_B_pG6bqBe88_2),.dout(w_dff_B_wHzXodWt3_2),.clk(gclk));
	jdff dff_B_ZcHLUDGF3_2(.din(w_dff_B_wHzXodWt3_2),.dout(w_dff_B_ZcHLUDGF3_2),.clk(gclk));
	jdff dff_B_TPGh4hOh5_2(.din(w_dff_B_ZcHLUDGF3_2),.dout(w_dff_B_TPGh4hOh5_2),.clk(gclk));
	jdff dff_B_2dfuuemb4_2(.din(w_dff_B_TPGh4hOh5_2),.dout(w_dff_B_2dfuuemb4_2),.clk(gclk));
	jdff dff_B_srbJV4312_2(.din(w_dff_B_2dfuuemb4_2),.dout(w_dff_B_srbJV4312_2),.clk(gclk));
	jdff dff_B_v0HKAo3k6_2(.din(w_dff_B_srbJV4312_2),.dout(w_dff_B_v0HKAo3k6_2),.clk(gclk));
	jdff dff_B_bWpJJRTS9_2(.din(w_dff_B_v0HKAo3k6_2),.dout(w_dff_B_bWpJJRTS9_2),.clk(gclk));
	jdff dff_B_1Z2HTE6W6_2(.din(w_dff_B_bWpJJRTS9_2),.dout(w_dff_B_1Z2HTE6W6_2),.clk(gclk));
	jdff dff_B_MX2almsg4_2(.din(w_dff_B_1Z2HTE6W6_2),.dout(w_dff_B_MX2almsg4_2),.clk(gclk));
	jdff dff_B_JtIv3EAd1_2(.din(w_dff_B_MX2almsg4_2),.dout(w_dff_B_JtIv3EAd1_2),.clk(gclk));
	jdff dff_B_XJXSJ4NN7_2(.din(w_dff_B_JtIv3EAd1_2),.dout(w_dff_B_XJXSJ4NN7_2),.clk(gclk));
	jdff dff_B_obN1Fa2Y3_2(.din(w_dff_B_XJXSJ4NN7_2),.dout(w_dff_B_obN1Fa2Y3_2),.clk(gclk));
	jdff dff_B_zXAbX5OI6_2(.din(w_dff_B_obN1Fa2Y3_2),.dout(w_dff_B_zXAbX5OI6_2),.clk(gclk));
	jdff dff_B_HWSRoIsS3_2(.din(w_dff_B_zXAbX5OI6_2),.dout(w_dff_B_HWSRoIsS3_2),.clk(gclk));
	jdff dff_B_U7LQDixK0_2(.din(w_dff_B_HWSRoIsS3_2),.dout(w_dff_B_U7LQDixK0_2),.clk(gclk));
	jdff dff_B_U1gigY8K5_2(.din(w_dff_B_U7LQDixK0_2),.dout(w_dff_B_U1gigY8K5_2),.clk(gclk));
	jdff dff_B_Wk5qA5Vz4_2(.din(w_dff_B_U1gigY8K5_2),.dout(w_dff_B_Wk5qA5Vz4_2),.clk(gclk));
	jdff dff_B_IjAhIE5b4_2(.din(w_dff_B_Wk5qA5Vz4_2),.dout(w_dff_B_IjAhIE5b4_2),.clk(gclk));
	jdff dff_B_uIwFxCoJ9_2(.din(w_dff_B_IjAhIE5b4_2),.dout(w_dff_B_uIwFxCoJ9_2),.clk(gclk));
	jdff dff_B_vUmxW7Al8_2(.din(w_dff_B_uIwFxCoJ9_2),.dout(w_dff_B_vUmxW7Al8_2),.clk(gclk));
	jdff dff_B_JF9L3uyX1_2(.din(w_dff_B_vUmxW7Al8_2),.dout(w_dff_B_JF9L3uyX1_2),.clk(gclk));
	jdff dff_B_9ma0up9x1_2(.din(w_dff_B_JF9L3uyX1_2),.dout(w_dff_B_9ma0up9x1_2),.clk(gclk));
	jdff dff_B_oxLHPdvN3_2(.din(w_dff_B_9ma0up9x1_2),.dout(w_dff_B_oxLHPdvN3_2),.clk(gclk));
	jdff dff_B_TdmzmMNp9_2(.din(w_dff_B_oxLHPdvN3_2),.dout(w_dff_B_TdmzmMNp9_2),.clk(gclk));
	jdff dff_B_P3OCRb2K7_2(.din(w_dff_B_TdmzmMNp9_2),.dout(w_dff_B_P3OCRb2K7_2),.clk(gclk));
	jdff dff_B_J1YjMSLR6_2(.din(w_dff_B_P3OCRb2K7_2),.dout(w_dff_B_J1YjMSLR6_2),.clk(gclk));
	jdff dff_B_FBIuk3mv6_2(.din(w_dff_B_J1YjMSLR6_2),.dout(w_dff_B_FBIuk3mv6_2),.clk(gclk));
	jdff dff_B_xfZV3ANG5_2(.din(w_dff_B_FBIuk3mv6_2),.dout(w_dff_B_xfZV3ANG5_2),.clk(gclk));
	jdff dff_B_tOaXRmgC1_2(.din(w_dff_B_xfZV3ANG5_2),.dout(w_dff_B_tOaXRmgC1_2),.clk(gclk));
	jdff dff_B_9eCQOicP7_2(.din(w_dff_B_tOaXRmgC1_2),.dout(w_dff_B_9eCQOicP7_2),.clk(gclk));
	jdff dff_B_WrJ6V0nm5_2(.din(n1656),.dout(w_dff_B_WrJ6V0nm5_2),.clk(gclk));
	jdff dff_B_t9D5uTt80_1(.din(n1654),.dout(w_dff_B_t9D5uTt80_1),.clk(gclk));
	jdff dff_B_pNYOjhVC9_2(.din(n1602),.dout(w_dff_B_pNYOjhVC9_2),.clk(gclk));
	jdff dff_B_5W9X6wvi3_2(.din(w_dff_B_pNYOjhVC9_2),.dout(w_dff_B_5W9X6wvi3_2),.clk(gclk));
	jdff dff_B_KHjqwb790_2(.din(w_dff_B_5W9X6wvi3_2),.dout(w_dff_B_KHjqwb790_2),.clk(gclk));
	jdff dff_B_dbEq4qeh2_2(.din(w_dff_B_KHjqwb790_2),.dout(w_dff_B_dbEq4qeh2_2),.clk(gclk));
	jdff dff_B_0hyjp00i9_2(.din(w_dff_B_dbEq4qeh2_2),.dout(w_dff_B_0hyjp00i9_2),.clk(gclk));
	jdff dff_B_vZ2J4v7S5_2(.din(w_dff_B_0hyjp00i9_2),.dout(w_dff_B_vZ2J4v7S5_2),.clk(gclk));
	jdff dff_B_XUycLhxH7_2(.din(w_dff_B_vZ2J4v7S5_2),.dout(w_dff_B_XUycLhxH7_2),.clk(gclk));
	jdff dff_B_tCZoC5kF9_2(.din(w_dff_B_XUycLhxH7_2),.dout(w_dff_B_tCZoC5kF9_2),.clk(gclk));
	jdff dff_B_wjaIMfrg1_2(.din(w_dff_B_tCZoC5kF9_2),.dout(w_dff_B_wjaIMfrg1_2),.clk(gclk));
	jdff dff_B_d6EuFWhm9_2(.din(w_dff_B_wjaIMfrg1_2),.dout(w_dff_B_d6EuFWhm9_2),.clk(gclk));
	jdff dff_B_SPKceGUe2_2(.din(w_dff_B_d6EuFWhm9_2),.dout(w_dff_B_SPKceGUe2_2),.clk(gclk));
	jdff dff_B_YCDekAtL9_2(.din(w_dff_B_SPKceGUe2_2),.dout(w_dff_B_YCDekAtL9_2),.clk(gclk));
	jdff dff_B_JlT7ObC32_2(.din(w_dff_B_YCDekAtL9_2),.dout(w_dff_B_JlT7ObC32_2),.clk(gclk));
	jdff dff_B_S8NFVUaB2_2(.din(w_dff_B_JlT7ObC32_2),.dout(w_dff_B_S8NFVUaB2_2),.clk(gclk));
	jdff dff_B_6X0kgRPa3_2(.din(w_dff_B_S8NFVUaB2_2),.dout(w_dff_B_6X0kgRPa3_2),.clk(gclk));
	jdff dff_B_mgBeuNHh3_2(.din(w_dff_B_6X0kgRPa3_2),.dout(w_dff_B_mgBeuNHh3_2),.clk(gclk));
	jdff dff_B_msd059e11_2(.din(w_dff_B_mgBeuNHh3_2),.dout(w_dff_B_msd059e11_2),.clk(gclk));
	jdff dff_B_HulELTYO0_2(.din(w_dff_B_msd059e11_2),.dout(w_dff_B_HulELTYO0_2),.clk(gclk));
	jdff dff_B_W0i79Icr6_2(.din(w_dff_B_HulELTYO0_2),.dout(w_dff_B_W0i79Icr6_2),.clk(gclk));
	jdff dff_B_22ltXU1U5_2(.din(w_dff_B_W0i79Icr6_2),.dout(w_dff_B_22ltXU1U5_2),.clk(gclk));
	jdff dff_B_tY3PL4BS3_2(.din(w_dff_B_22ltXU1U5_2),.dout(w_dff_B_tY3PL4BS3_2),.clk(gclk));
	jdff dff_B_glmeXJvf3_2(.din(w_dff_B_tY3PL4BS3_2),.dout(w_dff_B_glmeXJvf3_2),.clk(gclk));
	jdff dff_B_BTCRbjOH4_2(.din(w_dff_B_glmeXJvf3_2),.dout(w_dff_B_BTCRbjOH4_2),.clk(gclk));
	jdff dff_B_N1EjSTc73_2(.din(w_dff_B_BTCRbjOH4_2),.dout(w_dff_B_N1EjSTc73_2),.clk(gclk));
	jdff dff_B_IGIG1Wu73_2(.din(w_dff_B_N1EjSTc73_2),.dout(w_dff_B_IGIG1Wu73_2),.clk(gclk));
	jdff dff_B_874iPqy03_2(.din(w_dff_B_IGIG1Wu73_2),.dout(w_dff_B_874iPqy03_2),.clk(gclk));
	jdff dff_B_DPySylyg0_2(.din(w_dff_B_874iPqy03_2),.dout(w_dff_B_DPySylyg0_2),.clk(gclk));
	jdff dff_B_K6RHEaGa7_2(.din(w_dff_B_DPySylyg0_2),.dout(w_dff_B_K6RHEaGa7_2),.clk(gclk));
	jdff dff_B_IwEq0MXj4_2(.din(w_dff_B_K6RHEaGa7_2),.dout(w_dff_B_IwEq0MXj4_2),.clk(gclk));
	jdff dff_B_Ghr6fiuS3_2(.din(w_dff_B_IwEq0MXj4_2),.dout(w_dff_B_Ghr6fiuS3_2),.clk(gclk));
	jdff dff_B_ybiFY6b38_2(.din(w_dff_B_Ghr6fiuS3_2),.dout(w_dff_B_ybiFY6b38_2),.clk(gclk));
	jdff dff_B_uZLDrLUz0_2(.din(w_dff_B_ybiFY6b38_2),.dout(w_dff_B_uZLDrLUz0_2),.clk(gclk));
	jdff dff_B_ahSFkCHz7_2(.din(w_dff_B_uZLDrLUz0_2),.dout(w_dff_B_ahSFkCHz7_2),.clk(gclk));
	jdff dff_B_8QPG6n0H4_2(.din(w_dff_B_ahSFkCHz7_2),.dout(w_dff_B_8QPG6n0H4_2),.clk(gclk));
	jdff dff_B_sVk5CXUM7_2(.din(w_dff_B_8QPG6n0H4_2),.dout(w_dff_B_sVk5CXUM7_2),.clk(gclk));
	jdff dff_B_5L8wzYpj0_2(.din(w_dff_B_sVk5CXUM7_2),.dout(w_dff_B_5L8wzYpj0_2),.clk(gclk));
	jdff dff_B_5HqwWtqK8_2(.din(w_dff_B_5L8wzYpj0_2),.dout(w_dff_B_5HqwWtqK8_2),.clk(gclk));
	jdff dff_B_viTqWzlJ5_2(.din(w_dff_B_5HqwWtqK8_2),.dout(w_dff_B_viTqWzlJ5_2),.clk(gclk));
	jdff dff_B_5yoD2A4C2_2(.din(w_dff_B_viTqWzlJ5_2),.dout(w_dff_B_5yoD2A4C2_2),.clk(gclk));
	jdff dff_B_1xWcrS0v9_2(.din(w_dff_B_5yoD2A4C2_2),.dout(w_dff_B_1xWcrS0v9_2),.clk(gclk));
	jdff dff_B_2m7wddaq1_2(.din(w_dff_B_1xWcrS0v9_2),.dout(w_dff_B_2m7wddaq1_2),.clk(gclk));
	jdff dff_B_o9zY27mx9_2(.din(w_dff_B_2m7wddaq1_2),.dout(w_dff_B_o9zY27mx9_2),.clk(gclk));
	jdff dff_B_0qTTQ4Ah9_2(.din(n1605),.dout(w_dff_B_0qTTQ4Ah9_2),.clk(gclk));
	jdff dff_B_XFmAsQRz6_1(.din(n1603),.dout(w_dff_B_XFmAsQRz6_1),.clk(gclk));
	jdff dff_B_fvwodyaw1_2(.din(n1545),.dout(w_dff_B_fvwodyaw1_2),.clk(gclk));
	jdff dff_B_gNgMs2UZ8_2(.din(w_dff_B_fvwodyaw1_2),.dout(w_dff_B_gNgMs2UZ8_2),.clk(gclk));
	jdff dff_B_syuvkTXI7_2(.din(w_dff_B_gNgMs2UZ8_2),.dout(w_dff_B_syuvkTXI7_2),.clk(gclk));
	jdff dff_B_A2vbns6u9_2(.din(w_dff_B_syuvkTXI7_2),.dout(w_dff_B_A2vbns6u9_2),.clk(gclk));
	jdff dff_B_WJ7efmps6_2(.din(w_dff_B_A2vbns6u9_2),.dout(w_dff_B_WJ7efmps6_2),.clk(gclk));
	jdff dff_B_C16YQgUm8_2(.din(w_dff_B_WJ7efmps6_2),.dout(w_dff_B_C16YQgUm8_2),.clk(gclk));
	jdff dff_B_t52tujzu6_2(.din(w_dff_B_C16YQgUm8_2),.dout(w_dff_B_t52tujzu6_2),.clk(gclk));
	jdff dff_B_IkwsdRSm2_2(.din(w_dff_B_t52tujzu6_2),.dout(w_dff_B_IkwsdRSm2_2),.clk(gclk));
	jdff dff_B_JNrRfv6T2_2(.din(w_dff_B_IkwsdRSm2_2),.dout(w_dff_B_JNrRfv6T2_2),.clk(gclk));
	jdff dff_B_QzRvDUp34_2(.din(w_dff_B_JNrRfv6T2_2),.dout(w_dff_B_QzRvDUp34_2),.clk(gclk));
	jdff dff_B_san3x6Xe1_2(.din(w_dff_B_QzRvDUp34_2),.dout(w_dff_B_san3x6Xe1_2),.clk(gclk));
	jdff dff_B_TiZUP3T61_2(.din(w_dff_B_san3x6Xe1_2),.dout(w_dff_B_TiZUP3T61_2),.clk(gclk));
	jdff dff_B_KYWjDAKY4_2(.din(w_dff_B_TiZUP3T61_2),.dout(w_dff_B_KYWjDAKY4_2),.clk(gclk));
	jdff dff_B_hh3gpvA19_2(.din(w_dff_B_KYWjDAKY4_2),.dout(w_dff_B_hh3gpvA19_2),.clk(gclk));
	jdff dff_B_EDB4rhT63_2(.din(w_dff_B_hh3gpvA19_2),.dout(w_dff_B_EDB4rhT63_2),.clk(gclk));
	jdff dff_B_ZdiTDCdE8_2(.din(w_dff_B_EDB4rhT63_2),.dout(w_dff_B_ZdiTDCdE8_2),.clk(gclk));
	jdff dff_B_6zdidnU93_2(.din(w_dff_B_ZdiTDCdE8_2),.dout(w_dff_B_6zdidnU93_2),.clk(gclk));
	jdff dff_B_Pu5UpHsa0_2(.din(w_dff_B_6zdidnU93_2),.dout(w_dff_B_Pu5UpHsa0_2),.clk(gclk));
	jdff dff_B_GTM5hGc03_2(.din(w_dff_B_Pu5UpHsa0_2),.dout(w_dff_B_GTM5hGc03_2),.clk(gclk));
	jdff dff_B_9jsokTcW3_2(.din(w_dff_B_GTM5hGc03_2),.dout(w_dff_B_9jsokTcW3_2),.clk(gclk));
	jdff dff_B_7cCbKGA89_2(.din(w_dff_B_9jsokTcW3_2),.dout(w_dff_B_7cCbKGA89_2),.clk(gclk));
	jdff dff_B_6XVx36N21_2(.din(w_dff_B_7cCbKGA89_2),.dout(w_dff_B_6XVx36N21_2),.clk(gclk));
	jdff dff_B_0FfbOxez7_2(.din(w_dff_B_6XVx36N21_2),.dout(w_dff_B_0FfbOxez7_2),.clk(gclk));
	jdff dff_B_4uYe4nTv3_2(.din(w_dff_B_0FfbOxez7_2),.dout(w_dff_B_4uYe4nTv3_2),.clk(gclk));
	jdff dff_B_uhKaDYun1_2(.din(w_dff_B_4uYe4nTv3_2),.dout(w_dff_B_uhKaDYun1_2),.clk(gclk));
	jdff dff_B_4kvG4O9I4_2(.din(w_dff_B_uhKaDYun1_2),.dout(w_dff_B_4kvG4O9I4_2),.clk(gclk));
	jdff dff_B_zwY4jpUB0_2(.din(w_dff_B_4kvG4O9I4_2),.dout(w_dff_B_zwY4jpUB0_2),.clk(gclk));
	jdff dff_B_CRa0TBPZ1_2(.din(w_dff_B_zwY4jpUB0_2),.dout(w_dff_B_CRa0TBPZ1_2),.clk(gclk));
	jdff dff_B_exNDzymW9_2(.din(w_dff_B_CRa0TBPZ1_2),.dout(w_dff_B_exNDzymW9_2),.clk(gclk));
	jdff dff_B_lTc3NPak9_2(.din(w_dff_B_exNDzymW9_2),.dout(w_dff_B_lTc3NPak9_2),.clk(gclk));
	jdff dff_B_c9qIiq8j2_2(.din(w_dff_B_lTc3NPak9_2),.dout(w_dff_B_c9qIiq8j2_2),.clk(gclk));
	jdff dff_B_py3cDcPl0_2(.din(w_dff_B_c9qIiq8j2_2),.dout(w_dff_B_py3cDcPl0_2),.clk(gclk));
	jdff dff_B_TcBjEos55_2(.din(w_dff_B_py3cDcPl0_2),.dout(w_dff_B_TcBjEos55_2),.clk(gclk));
	jdff dff_B_FrGPuZe21_2(.din(w_dff_B_TcBjEos55_2),.dout(w_dff_B_FrGPuZe21_2),.clk(gclk));
	jdff dff_B_6F0HSgVC7_2(.din(w_dff_B_FrGPuZe21_2),.dout(w_dff_B_6F0HSgVC7_2),.clk(gclk));
	jdff dff_B_e4mtod7U1_2(.din(w_dff_B_6F0HSgVC7_2),.dout(w_dff_B_e4mtod7U1_2),.clk(gclk));
	jdff dff_B_kAtuO9bV5_2(.din(w_dff_B_e4mtod7U1_2),.dout(w_dff_B_kAtuO9bV5_2),.clk(gclk));
	jdff dff_B_PcSwCouR6_2(.din(w_dff_B_kAtuO9bV5_2),.dout(w_dff_B_PcSwCouR6_2),.clk(gclk));
	jdff dff_B_16aT5zsN1_1(.din(n1546),.dout(w_dff_B_16aT5zsN1_1),.clk(gclk));
	jdff dff_B_3pLSN5CG3_2(.din(n1481),.dout(w_dff_B_3pLSN5CG3_2),.clk(gclk));
	jdff dff_B_CazexgUy6_2(.din(w_dff_B_3pLSN5CG3_2),.dout(w_dff_B_CazexgUy6_2),.clk(gclk));
	jdff dff_B_8vyIbKAw5_2(.din(w_dff_B_CazexgUy6_2),.dout(w_dff_B_8vyIbKAw5_2),.clk(gclk));
	jdff dff_B_YnRnSAN96_2(.din(w_dff_B_8vyIbKAw5_2),.dout(w_dff_B_YnRnSAN96_2),.clk(gclk));
	jdff dff_B_IveJ91e54_2(.din(w_dff_B_YnRnSAN96_2),.dout(w_dff_B_IveJ91e54_2),.clk(gclk));
	jdff dff_B_OA9vheDX3_2(.din(w_dff_B_IveJ91e54_2),.dout(w_dff_B_OA9vheDX3_2),.clk(gclk));
	jdff dff_B_w0gPgVsl0_2(.din(w_dff_B_OA9vheDX3_2),.dout(w_dff_B_w0gPgVsl0_2),.clk(gclk));
	jdff dff_B_EnltlGRM5_2(.din(w_dff_B_w0gPgVsl0_2),.dout(w_dff_B_EnltlGRM5_2),.clk(gclk));
	jdff dff_B_NtXKQfB58_2(.din(w_dff_B_EnltlGRM5_2),.dout(w_dff_B_NtXKQfB58_2),.clk(gclk));
	jdff dff_B_2E9D7a5M1_2(.din(w_dff_B_NtXKQfB58_2),.dout(w_dff_B_2E9D7a5M1_2),.clk(gclk));
	jdff dff_B_uRJ3iyoj2_2(.din(w_dff_B_2E9D7a5M1_2),.dout(w_dff_B_uRJ3iyoj2_2),.clk(gclk));
	jdff dff_B_ef8N4YWm2_2(.din(w_dff_B_uRJ3iyoj2_2),.dout(w_dff_B_ef8N4YWm2_2),.clk(gclk));
	jdff dff_B_0dFP5lOF9_2(.din(w_dff_B_ef8N4YWm2_2),.dout(w_dff_B_0dFP5lOF9_2),.clk(gclk));
	jdff dff_B_6CkqVLE86_2(.din(w_dff_B_0dFP5lOF9_2),.dout(w_dff_B_6CkqVLE86_2),.clk(gclk));
	jdff dff_B_jMVzD7GU2_2(.din(w_dff_B_6CkqVLE86_2),.dout(w_dff_B_jMVzD7GU2_2),.clk(gclk));
	jdff dff_B_EzqaJBGg4_2(.din(w_dff_B_jMVzD7GU2_2),.dout(w_dff_B_EzqaJBGg4_2),.clk(gclk));
	jdff dff_B_HHpoGZCe5_2(.din(w_dff_B_EzqaJBGg4_2),.dout(w_dff_B_HHpoGZCe5_2),.clk(gclk));
	jdff dff_B_FyVQqYve0_2(.din(w_dff_B_HHpoGZCe5_2),.dout(w_dff_B_FyVQqYve0_2),.clk(gclk));
	jdff dff_B_3MahnG3q5_2(.din(w_dff_B_FyVQqYve0_2),.dout(w_dff_B_3MahnG3q5_2),.clk(gclk));
	jdff dff_B_uGnD9CkP2_2(.din(w_dff_B_3MahnG3q5_2),.dout(w_dff_B_uGnD9CkP2_2),.clk(gclk));
	jdff dff_B_AqOa60tT2_2(.din(w_dff_B_uGnD9CkP2_2),.dout(w_dff_B_AqOa60tT2_2),.clk(gclk));
	jdff dff_B_SBy6zCVB8_2(.din(w_dff_B_AqOa60tT2_2),.dout(w_dff_B_SBy6zCVB8_2),.clk(gclk));
	jdff dff_B_uhaj9Mai1_2(.din(w_dff_B_SBy6zCVB8_2),.dout(w_dff_B_uhaj9Mai1_2),.clk(gclk));
	jdff dff_B_uSF582VV1_2(.din(w_dff_B_uhaj9Mai1_2),.dout(w_dff_B_uSF582VV1_2),.clk(gclk));
	jdff dff_B_Z62PFuGl9_2(.din(w_dff_B_uSF582VV1_2),.dout(w_dff_B_Z62PFuGl9_2),.clk(gclk));
	jdff dff_B_Q8k6Skgy8_2(.din(w_dff_B_Z62PFuGl9_2),.dout(w_dff_B_Q8k6Skgy8_2),.clk(gclk));
	jdff dff_B_7cNMhV7X9_2(.din(w_dff_B_Q8k6Skgy8_2),.dout(w_dff_B_7cNMhV7X9_2),.clk(gclk));
	jdff dff_B_tHSvPa6A3_2(.din(w_dff_B_7cNMhV7X9_2),.dout(w_dff_B_tHSvPa6A3_2),.clk(gclk));
	jdff dff_B_V0Mg8WqM5_2(.din(w_dff_B_tHSvPa6A3_2),.dout(w_dff_B_V0Mg8WqM5_2),.clk(gclk));
	jdff dff_B_gIZeW8nP4_2(.din(w_dff_B_V0Mg8WqM5_2),.dout(w_dff_B_gIZeW8nP4_2),.clk(gclk));
	jdff dff_B_6bj8HGa52_2(.din(w_dff_B_gIZeW8nP4_2),.dout(w_dff_B_6bj8HGa52_2),.clk(gclk));
	jdff dff_B_Qpys5LsV2_2(.din(w_dff_B_6bj8HGa52_2),.dout(w_dff_B_Qpys5LsV2_2),.clk(gclk));
	jdff dff_B_Wd5rhdrX9_2(.din(w_dff_B_Qpys5LsV2_2),.dout(w_dff_B_Wd5rhdrX9_2),.clk(gclk));
	jdff dff_B_3v7FLQP13_2(.din(w_dff_B_Wd5rhdrX9_2),.dout(w_dff_B_3v7FLQP13_2),.clk(gclk));
	jdff dff_B_5wq6JhJu8_2(.din(w_dff_B_3v7FLQP13_2),.dout(w_dff_B_5wq6JhJu8_2),.clk(gclk));
	jdff dff_B_wnhFjLNo7_2(.din(n1513),.dout(w_dff_B_wnhFjLNo7_2),.clk(gclk));
	jdff dff_B_1GGwFMXf4_1(.din(n1482),.dout(w_dff_B_1GGwFMXf4_1),.clk(gclk));
	jdff dff_B_KVsQxj5R5_2(.din(n1410),.dout(w_dff_B_KVsQxj5R5_2),.clk(gclk));
	jdff dff_B_avIcZMrb1_2(.din(w_dff_B_KVsQxj5R5_2),.dout(w_dff_B_avIcZMrb1_2),.clk(gclk));
	jdff dff_B_iEXG9xPY9_2(.din(w_dff_B_avIcZMrb1_2),.dout(w_dff_B_iEXG9xPY9_2),.clk(gclk));
	jdff dff_B_WkLhh7J52_2(.din(w_dff_B_iEXG9xPY9_2),.dout(w_dff_B_WkLhh7J52_2),.clk(gclk));
	jdff dff_B_frBDfW6X0_2(.din(w_dff_B_WkLhh7J52_2),.dout(w_dff_B_frBDfW6X0_2),.clk(gclk));
	jdff dff_B_sLa1qN8a2_2(.din(w_dff_B_frBDfW6X0_2),.dout(w_dff_B_sLa1qN8a2_2),.clk(gclk));
	jdff dff_B_pRjce0Ks8_2(.din(w_dff_B_sLa1qN8a2_2),.dout(w_dff_B_pRjce0Ks8_2),.clk(gclk));
	jdff dff_B_ytoBCoOm1_2(.din(w_dff_B_pRjce0Ks8_2),.dout(w_dff_B_ytoBCoOm1_2),.clk(gclk));
	jdff dff_B_sEyaELGB1_2(.din(w_dff_B_ytoBCoOm1_2),.dout(w_dff_B_sEyaELGB1_2),.clk(gclk));
	jdff dff_B_i4n86loG1_2(.din(w_dff_B_sEyaELGB1_2),.dout(w_dff_B_i4n86loG1_2),.clk(gclk));
	jdff dff_B_MH75h9N42_2(.din(w_dff_B_i4n86loG1_2),.dout(w_dff_B_MH75h9N42_2),.clk(gclk));
	jdff dff_B_ccx6fG382_2(.din(w_dff_B_MH75h9N42_2),.dout(w_dff_B_ccx6fG382_2),.clk(gclk));
	jdff dff_B_qErzRpsU7_2(.din(w_dff_B_ccx6fG382_2),.dout(w_dff_B_qErzRpsU7_2),.clk(gclk));
	jdff dff_B_KnTHTJ6V6_2(.din(w_dff_B_qErzRpsU7_2),.dout(w_dff_B_KnTHTJ6V6_2),.clk(gclk));
	jdff dff_B_92WceIax7_2(.din(w_dff_B_KnTHTJ6V6_2),.dout(w_dff_B_92WceIax7_2),.clk(gclk));
	jdff dff_B_qgo46wpE7_2(.din(w_dff_B_92WceIax7_2),.dout(w_dff_B_qgo46wpE7_2),.clk(gclk));
	jdff dff_B_fXnTDbjO6_2(.din(w_dff_B_qgo46wpE7_2),.dout(w_dff_B_fXnTDbjO6_2),.clk(gclk));
	jdff dff_B_eUYFIQY90_2(.din(w_dff_B_fXnTDbjO6_2),.dout(w_dff_B_eUYFIQY90_2),.clk(gclk));
	jdff dff_B_NssLkWHN1_2(.din(w_dff_B_eUYFIQY90_2),.dout(w_dff_B_NssLkWHN1_2),.clk(gclk));
	jdff dff_B_zFHoNNH77_2(.din(w_dff_B_NssLkWHN1_2),.dout(w_dff_B_zFHoNNH77_2),.clk(gclk));
	jdff dff_B_V4VrACSw7_2(.din(w_dff_B_zFHoNNH77_2),.dout(w_dff_B_V4VrACSw7_2),.clk(gclk));
	jdff dff_B_GoZvDL4v5_2(.din(w_dff_B_V4VrACSw7_2),.dout(w_dff_B_GoZvDL4v5_2),.clk(gclk));
	jdff dff_B_s9opWJOP0_2(.din(w_dff_B_GoZvDL4v5_2),.dout(w_dff_B_s9opWJOP0_2),.clk(gclk));
	jdff dff_B_FW0RCixr1_2(.din(w_dff_B_s9opWJOP0_2),.dout(w_dff_B_FW0RCixr1_2),.clk(gclk));
	jdff dff_B_6uEMwGVI0_2(.din(w_dff_B_FW0RCixr1_2),.dout(w_dff_B_6uEMwGVI0_2),.clk(gclk));
	jdff dff_B_7aWfhsmM8_2(.din(w_dff_B_6uEMwGVI0_2),.dout(w_dff_B_7aWfhsmM8_2),.clk(gclk));
	jdff dff_B_l7O45QNP2_2(.din(w_dff_B_7aWfhsmM8_2),.dout(w_dff_B_l7O45QNP2_2),.clk(gclk));
	jdff dff_B_rswdLXD06_2(.din(w_dff_B_l7O45QNP2_2),.dout(w_dff_B_rswdLXD06_2),.clk(gclk));
	jdff dff_B_R8TsZpYj4_2(.din(w_dff_B_rswdLXD06_2),.dout(w_dff_B_R8TsZpYj4_2),.clk(gclk));
	jdff dff_B_8gPLJpK13_2(.din(w_dff_B_R8TsZpYj4_2),.dout(w_dff_B_8gPLJpK13_2),.clk(gclk));
	jdff dff_B_icy7nypp6_2(.din(w_dff_B_8gPLJpK13_2),.dout(w_dff_B_icy7nypp6_2),.clk(gclk));
	jdff dff_B_kL36koVf8_2(.din(w_dff_B_icy7nypp6_2),.dout(w_dff_B_kL36koVf8_2),.clk(gclk));
	jdff dff_B_QSdI15m68_2(.din(n1442),.dout(w_dff_B_QSdI15m68_2),.clk(gclk));
	jdff dff_B_03C4d0Nz5_1(.din(n1411),.dout(w_dff_B_03C4d0Nz5_1),.clk(gclk));
	jdff dff_B_ZTRAGPzd5_2(.din(n1332),.dout(w_dff_B_ZTRAGPzd5_2),.clk(gclk));
	jdff dff_B_9mUIdDGm1_2(.din(w_dff_B_ZTRAGPzd5_2),.dout(w_dff_B_9mUIdDGm1_2),.clk(gclk));
	jdff dff_B_sRiNvewp2_2(.din(w_dff_B_9mUIdDGm1_2),.dout(w_dff_B_sRiNvewp2_2),.clk(gclk));
	jdff dff_B_SCk0ElQf8_2(.din(w_dff_B_sRiNvewp2_2),.dout(w_dff_B_SCk0ElQf8_2),.clk(gclk));
	jdff dff_B_6Qw9lyRy7_2(.din(w_dff_B_SCk0ElQf8_2),.dout(w_dff_B_6Qw9lyRy7_2),.clk(gclk));
	jdff dff_B_HcrkmSGr1_2(.din(w_dff_B_6Qw9lyRy7_2),.dout(w_dff_B_HcrkmSGr1_2),.clk(gclk));
	jdff dff_B_PcIRYYr12_2(.din(w_dff_B_HcrkmSGr1_2),.dout(w_dff_B_PcIRYYr12_2),.clk(gclk));
	jdff dff_B_IuBtgw9k2_2(.din(w_dff_B_PcIRYYr12_2),.dout(w_dff_B_IuBtgw9k2_2),.clk(gclk));
	jdff dff_B_cCjUmUSv2_2(.din(w_dff_B_IuBtgw9k2_2),.dout(w_dff_B_cCjUmUSv2_2),.clk(gclk));
	jdff dff_B_mCgLaQyL4_2(.din(w_dff_B_cCjUmUSv2_2),.dout(w_dff_B_mCgLaQyL4_2),.clk(gclk));
	jdff dff_B_SvrCyC528_2(.din(w_dff_B_mCgLaQyL4_2),.dout(w_dff_B_SvrCyC528_2),.clk(gclk));
	jdff dff_B_LVEWAfhX3_2(.din(w_dff_B_SvrCyC528_2),.dout(w_dff_B_LVEWAfhX3_2),.clk(gclk));
	jdff dff_B_rfA7ybRF7_2(.din(w_dff_B_LVEWAfhX3_2),.dout(w_dff_B_rfA7ybRF7_2),.clk(gclk));
	jdff dff_B_6RdFhHoK9_2(.din(w_dff_B_rfA7ybRF7_2),.dout(w_dff_B_6RdFhHoK9_2),.clk(gclk));
	jdff dff_B_IMN8IZXh3_2(.din(w_dff_B_6RdFhHoK9_2),.dout(w_dff_B_IMN8IZXh3_2),.clk(gclk));
	jdff dff_B_i5BBpHps1_2(.din(w_dff_B_IMN8IZXh3_2),.dout(w_dff_B_i5BBpHps1_2),.clk(gclk));
	jdff dff_B_EDWDpFGB3_2(.din(w_dff_B_i5BBpHps1_2),.dout(w_dff_B_EDWDpFGB3_2),.clk(gclk));
	jdff dff_B_LG7Q3p3Z0_2(.din(w_dff_B_EDWDpFGB3_2),.dout(w_dff_B_LG7Q3p3Z0_2),.clk(gclk));
	jdff dff_B_ZIM0uiyb7_2(.din(w_dff_B_LG7Q3p3Z0_2),.dout(w_dff_B_ZIM0uiyb7_2),.clk(gclk));
	jdff dff_B_NRyVUIUT4_2(.din(w_dff_B_ZIM0uiyb7_2),.dout(w_dff_B_NRyVUIUT4_2),.clk(gclk));
	jdff dff_B_3bFWeXvq1_2(.din(w_dff_B_NRyVUIUT4_2),.dout(w_dff_B_3bFWeXvq1_2),.clk(gclk));
	jdff dff_B_fCgLx2Ab8_2(.din(w_dff_B_3bFWeXvq1_2),.dout(w_dff_B_fCgLx2Ab8_2),.clk(gclk));
	jdff dff_B_Qy1bWVMt1_2(.din(w_dff_B_fCgLx2Ab8_2),.dout(w_dff_B_Qy1bWVMt1_2),.clk(gclk));
	jdff dff_B_TOdpPG1v6_2(.din(w_dff_B_Qy1bWVMt1_2),.dout(w_dff_B_TOdpPG1v6_2),.clk(gclk));
	jdff dff_B_S0umS0Q60_2(.din(w_dff_B_TOdpPG1v6_2),.dout(w_dff_B_S0umS0Q60_2),.clk(gclk));
	jdff dff_B_89mD8GuJ6_2(.din(w_dff_B_S0umS0Q60_2),.dout(w_dff_B_89mD8GuJ6_2),.clk(gclk));
	jdff dff_B_vSKpSpCu6_2(.din(w_dff_B_89mD8GuJ6_2),.dout(w_dff_B_vSKpSpCu6_2),.clk(gclk));
	jdff dff_B_2AvGAdzv3_2(.din(w_dff_B_vSKpSpCu6_2),.dout(w_dff_B_2AvGAdzv3_2),.clk(gclk));
	jdff dff_B_B4idFpAm8_2(.din(w_dff_B_2AvGAdzv3_2),.dout(w_dff_B_B4idFpAm8_2),.clk(gclk));
	jdff dff_B_FMdovfI97_2(.din(n1364),.dout(w_dff_B_FMdovfI97_2),.clk(gclk));
	jdff dff_B_3YJs9FYL7_1(.din(n1333),.dout(w_dff_B_3YJs9FYL7_1),.clk(gclk));
	jdff dff_B_O909kjOB6_2(.din(n1247),.dout(w_dff_B_O909kjOB6_2),.clk(gclk));
	jdff dff_B_9cjHc9BA0_2(.din(w_dff_B_O909kjOB6_2),.dout(w_dff_B_9cjHc9BA0_2),.clk(gclk));
	jdff dff_B_MVX68V2I7_2(.din(w_dff_B_9cjHc9BA0_2),.dout(w_dff_B_MVX68V2I7_2),.clk(gclk));
	jdff dff_B_JKNQFBoV8_2(.din(w_dff_B_MVX68V2I7_2),.dout(w_dff_B_JKNQFBoV8_2),.clk(gclk));
	jdff dff_B_uKLSG0b28_2(.din(w_dff_B_JKNQFBoV8_2),.dout(w_dff_B_uKLSG0b28_2),.clk(gclk));
	jdff dff_B_H9Dp2Wn96_2(.din(w_dff_B_uKLSG0b28_2),.dout(w_dff_B_H9Dp2Wn96_2),.clk(gclk));
	jdff dff_B_dFG8EpLY0_2(.din(w_dff_B_H9Dp2Wn96_2),.dout(w_dff_B_dFG8EpLY0_2),.clk(gclk));
	jdff dff_B_kp039gr16_2(.din(w_dff_B_dFG8EpLY0_2),.dout(w_dff_B_kp039gr16_2),.clk(gclk));
	jdff dff_B_3DKnH1Yz6_2(.din(w_dff_B_kp039gr16_2),.dout(w_dff_B_3DKnH1Yz6_2),.clk(gclk));
	jdff dff_B_YPKdWiKd3_2(.din(w_dff_B_3DKnH1Yz6_2),.dout(w_dff_B_YPKdWiKd3_2),.clk(gclk));
	jdff dff_B_gwKTBcxk1_2(.din(w_dff_B_YPKdWiKd3_2),.dout(w_dff_B_gwKTBcxk1_2),.clk(gclk));
	jdff dff_B_VMQBcAm46_2(.din(w_dff_B_gwKTBcxk1_2),.dout(w_dff_B_VMQBcAm46_2),.clk(gclk));
	jdff dff_B_hYocLxTP7_2(.din(w_dff_B_VMQBcAm46_2),.dout(w_dff_B_hYocLxTP7_2),.clk(gclk));
	jdff dff_B_dou3UOQX5_2(.din(w_dff_B_hYocLxTP7_2),.dout(w_dff_B_dou3UOQX5_2),.clk(gclk));
	jdff dff_B_OSju6Gw70_2(.din(w_dff_B_dou3UOQX5_2),.dout(w_dff_B_OSju6Gw70_2),.clk(gclk));
	jdff dff_B_PzPFNVaN8_2(.din(w_dff_B_OSju6Gw70_2),.dout(w_dff_B_PzPFNVaN8_2),.clk(gclk));
	jdff dff_B_wdwGwaL93_2(.din(w_dff_B_PzPFNVaN8_2),.dout(w_dff_B_wdwGwaL93_2),.clk(gclk));
	jdff dff_B_MeVbMxQn0_2(.din(w_dff_B_wdwGwaL93_2),.dout(w_dff_B_MeVbMxQn0_2),.clk(gclk));
	jdff dff_B_XnuWoWXB9_2(.din(w_dff_B_MeVbMxQn0_2),.dout(w_dff_B_XnuWoWXB9_2),.clk(gclk));
	jdff dff_B_iLwZvHKa8_2(.din(w_dff_B_XnuWoWXB9_2),.dout(w_dff_B_iLwZvHKa8_2),.clk(gclk));
	jdff dff_B_R6KMT4Hv1_2(.din(w_dff_B_iLwZvHKa8_2),.dout(w_dff_B_R6KMT4Hv1_2),.clk(gclk));
	jdff dff_B_wkF0Ap7w4_2(.din(w_dff_B_R6KMT4Hv1_2),.dout(w_dff_B_wkF0Ap7w4_2),.clk(gclk));
	jdff dff_B_VHx9nbKy2_2(.din(w_dff_B_wkF0Ap7w4_2),.dout(w_dff_B_VHx9nbKy2_2),.clk(gclk));
	jdff dff_B_syeGgtK06_2(.din(w_dff_B_VHx9nbKy2_2),.dout(w_dff_B_syeGgtK06_2),.clk(gclk));
	jdff dff_B_8f5t40EH4_2(.din(w_dff_B_syeGgtK06_2),.dout(w_dff_B_8f5t40EH4_2),.clk(gclk));
	jdff dff_B_vPZYQ9446_2(.din(w_dff_B_8f5t40EH4_2),.dout(w_dff_B_vPZYQ9446_2),.clk(gclk));
	jdff dff_B_Lm9mW8yr3_2(.din(n1279),.dout(w_dff_B_Lm9mW8yr3_2),.clk(gclk));
	jdff dff_B_r1b8WR3B7_1(.din(n1248),.dout(w_dff_B_r1b8WR3B7_1),.clk(gclk));
	jdff dff_B_x3mFtPrJ8_2(.din(n1156),.dout(w_dff_B_x3mFtPrJ8_2),.clk(gclk));
	jdff dff_B_liXXXrSw7_2(.din(w_dff_B_x3mFtPrJ8_2),.dout(w_dff_B_liXXXrSw7_2),.clk(gclk));
	jdff dff_B_EUqn5DNy8_2(.din(w_dff_B_liXXXrSw7_2),.dout(w_dff_B_EUqn5DNy8_2),.clk(gclk));
	jdff dff_B_L8DOvECq1_2(.din(w_dff_B_EUqn5DNy8_2),.dout(w_dff_B_L8DOvECq1_2),.clk(gclk));
	jdff dff_B_GZwLpp811_2(.din(w_dff_B_L8DOvECq1_2),.dout(w_dff_B_GZwLpp811_2),.clk(gclk));
	jdff dff_B_i7kLmSo80_2(.din(w_dff_B_GZwLpp811_2),.dout(w_dff_B_i7kLmSo80_2),.clk(gclk));
	jdff dff_B_ziWRDt3A1_2(.din(w_dff_B_i7kLmSo80_2),.dout(w_dff_B_ziWRDt3A1_2),.clk(gclk));
	jdff dff_B_zxyjUr9d6_2(.din(w_dff_B_ziWRDt3A1_2),.dout(w_dff_B_zxyjUr9d6_2),.clk(gclk));
	jdff dff_B_Iil3oNRz3_2(.din(w_dff_B_zxyjUr9d6_2),.dout(w_dff_B_Iil3oNRz3_2),.clk(gclk));
	jdff dff_B_9GIOokJC5_2(.din(w_dff_B_Iil3oNRz3_2),.dout(w_dff_B_9GIOokJC5_2),.clk(gclk));
	jdff dff_B_SgO2pyAa9_2(.din(w_dff_B_9GIOokJC5_2),.dout(w_dff_B_SgO2pyAa9_2),.clk(gclk));
	jdff dff_B_k6iOAHRL2_2(.din(w_dff_B_SgO2pyAa9_2),.dout(w_dff_B_k6iOAHRL2_2),.clk(gclk));
	jdff dff_B_qk8FC8x47_2(.din(w_dff_B_k6iOAHRL2_2),.dout(w_dff_B_qk8FC8x47_2),.clk(gclk));
	jdff dff_B_wb14hT8h8_2(.din(w_dff_B_qk8FC8x47_2),.dout(w_dff_B_wb14hT8h8_2),.clk(gclk));
	jdff dff_B_PDZxi2Ag9_2(.din(w_dff_B_wb14hT8h8_2),.dout(w_dff_B_PDZxi2Ag9_2),.clk(gclk));
	jdff dff_B_IGOaujNL1_2(.din(w_dff_B_PDZxi2Ag9_2),.dout(w_dff_B_IGOaujNL1_2),.clk(gclk));
	jdff dff_B_91cugucc0_2(.din(w_dff_B_IGOaujNL1_2),.dout(w_dff_B_91cugucc0_2),.clk(gclk));
	jdff dff_B_PMNHLCSo4_2(.din(w_dff_B_91cugucc0_2),.dout(w_dff_B_PMNHLCSo4_2),.clk(gclk));
	jdff dff_B_Nu2s07Qw3_2(.din(w_dff_B_PMNHLCSo4_2),.dout(w_dff_B_Nu2s07Qw3_2),.clk(gclk));
	jdff dff_B_lIQmthI84_2(.din(w_dff_B_Nu2s07Qw3_2),.dout(w_dff_B_lIQmthI84_2),.clk(gclk));
	jdff dff_B_osVDgbw17_2(.din(w_dff_B_lIQmthI84_2),.dout(w_dff_B_osVDgbw17_2),.clk(gclk));
	jdff dff_B_Z6oTmj7y9_2(.din(w_dff_B_osVDgbw17_2),.dout(w_dff_B_Z6oTmj7y9_2),.clk(gclk));
	jdff dff_B_04xkvR896_2(.din(w_dff_B_Z6oTmj7y9_2),.dout(w_dff_B_04xkvR896_2),.clk(gclk));
	jdff dff_B_y33tYOu80_2(.din(n1188),.dout(w_dff_B_y33tYOu80_2),.clk(gclk));
	jdff dff_B_dFvhUsMM4_1(.din(n1157),.dout(w_dff_B_dFvhUsMM4_1),.clk(gclk));
	jdff dff_B_51y7hsma4_2(.din(n1058),.dout(w_dff_B_51y7hsma4_2),.clk(gclk));
	jdff dff_B_f1KX6mMl1_2(.din(w_dff_B_51y7hsma4_2),.dout(w_dff_B_f1KX6mMl1_2),.clk(gclk));
	jdff dff_B_bIDddtaF4_2(.din(w_dff_B_f1KX6mMl1_2),.dout(w_dff_B_bIDddtaF4_2),.clk(gclk));
	jdff dff_B_GwOFstOW2_2(.din(w_dff_B_bIDddtaF4_2),.dout(w_dff_B_GwOFstOW2_2),.clk(gclk));
	jdff dff_B_TmlORck29_2(.din(w_dff_B_GwOFstOW2_2),.dout(w_dff_B_TmlORck29_2),.clk(gclk));
	jdff dff_B_hbDt7uwv2_2(.din(w_dff_B_TmlORck29_2),.dout(w_dff_B_hbDt7uwv2_2),.clk(gclk));
	jdff dff_B_fAU1TFqW5_2(.din(w_dff_B_hbDt7uwv2_2),.dout(w_dff_B_fAU1TFqW5_2),.clk(gclk));
	jdff dff_B_vnrKLf7b2_2(.din(w_dff_B_fAU1TFqW5_2),.dout(w_dff_B_vnrKLf7b2_2),.clk(gclk));
	jdff dff_B_pAnLs9fe8_2(.din(w_dff_B_vnrKLf7b2_2),.dout(w_dff_B_pAnLs9fe8_2),.clk(gclk));
	jdff dff_B_5eKEgA4p4_2(.din(w_dff_B_pAnLs9fe8_2),.dout(w_dff_B_5eKEgA4p4_2),.clk(gclk));
	jdff dff_B_Y3Aqfz2K4_2(.din(w_dff_B_5eKEgA4p4_2),.dout(w_dff_B_Y3Aqfz2K4_2),.clk(gclk));
	jdff dff_B_pcHUbSNj9_2(.din(w_dff_B_Y3Aqfz2K4_2),.dout(w_dff_B_pcHUbSNj9_2),.clk(gclk));
	jdff dff_B_Wf9ylcjt6_2(.din(w_dff_B_pcHUbSNj9_2),.dout(w_dff_B_Wf9ylcjt6_2),.clk(gclk));
	jdff dff_B_KvGUxGQp0_2(.din(w_dff_B_Wf9ylcjt6_2),.dout(w_dff_B_KvGUxGQp0_2),.clk(gclk));
	jdff dff_B_BeL5p8Pj2_2(.din(w_dff_B_KvGUxGQp0_2),.dout(w_dff_B_BeL5p8Pj2_2),.clk(gclk));
	jdff dff_B_6Iu4fln07_2(.din(w_dff_B_BeL5p8Pj2_2),.dout(w_dff_B_6Iu4fln07_2),.clk(gclk));
	jdff dff_B_YvpQtGn88_2(.din(w_dff_B_6Iu4fln07_2),.dout(w_dff_B_YvpQtGn88_2),.clk(gclk));
	jdff dff_B_Qn9R1tgg8_2(.din(w_dff_B_YvpQtGn88_2),.dout(w_dff_B_Qn9R1tgg8_2),.clk(gclk));
	jdff dff_B_WTLmxP1M8_2(.din(w_dff_B_Qn9R1tgg8_2),.dout(w_dff_B_WTLmxP1M8_2),.clk(gclk));
	jdff dff_B_7FGqqgOK4_2(.din(w_dff_B_WTLmxP1M8_2),.dout(w_dff_B_7FGqqgOK4_2),.clk(gclk));
	jdff dff_B_MV1nrUwB4_2(.din(n1089),.dout(w_dff_B_MV1nrUwB4_2),.clk(gclk));
	jdff dff_B_cexRrHv16_1(.din(n1059),.dout(w_dff_B_cexRrHv16_1),.clk(gclk));
	jdff dff_B_KWlvKiXB7_2(.din(n959),.dout(w_dff_B_KWlvKiXB7_2),.clk(gclk));
	jdff dff_B_oqHToH5b6_2(.din(w_dff_B_KWlvKiXB7_2),.dout(w_dff_B_oqHToH5b6_2),.clk(gclk));
	jdff dff_B_sHph7eFO0_2(.din(w_dff_B_oqHToH5b6_2),.dout(w_dff_B_sHph7eFO0_2),.clk(gclk));
	jdff dff_B_tFYH2YVv9_2(.din(w_dff_B_sHph7eFO0_2),.dout(w_dff_B_tFYH2YVv9_2),.clk(gclk));
	jdff dff_B_8WGE9fUd9_2(.din(w_dff_B_tFYH2YVv9_2),.dout(w_dff_B_8WGE9fUd9_2),.clk(gclk));
	jdff dff_B_iBJUXVJm7_2(.din(w_dff_B_8WGE9fUd9_2),.dout(w_dff_B_iBJUXVJm7_2),.clk(gclk));
	jdff dff_B_1e6Oejm25_2(.din(w_dff_B_iBJUXVJm7_2),.dout(w_dff_B_1e6Oejm25_2),.clk(gclk));
	jdff dff_B_Tyy0JRCP1_2(.din(w_dff_B_1e6Oejm25_2),.dout(w_dff_B_Tyy0JRCP1_2),.clk(gclk));
	jdff dff_B_MD93t9ql0_2(.din(w_dff_B_Tyy0JRCP1_2),.dout(w_dff_B_MD93t9ql0_2),.clk(gclk));
	jdff dff_B_NYJavSmY3_2(.din(w_dff_B_MD93t9ql0_2),.dout(w_dff_B_NYJavSmY3_2),.clk(gclk));
	jdff dff_B_jQGM1Ts92_2(.din(w_dff_B_NYJavSmY3_2),.dout(w_dff_B_jQGM1Ts92_2),.clk(gclk));
	jdff dff_B_hYmhH8Wz1_2(.din(w_dff_B_jQGM1Ts92_2),.dout(w_dff_B_hYmhH8Wz1_2),.clk(gclk));
	jdff dff_B_0zZ2AAQo3_2(.din(w_dff_B_hYmhH8Wz1_2),.dout(w_dff_B_0zZ2AAQo3_2),.clk(gclk));
	jdff dff_B_Cxmen5VL8_2(.din(w_dff_B_0zZ2AAQo3_2),.dout(w_dff_B_Cxmen5VL8_2),.clk(gclk));
	jdff dff_B_JzCAXZbT5_2(.din(w_dff_B_Cxmen5VL8_2),.dout(w_dff_B_JzCAXZbT5_2),.clk(gclk));
	jdff dff_B_z7HxxPCg7_2(.din(w_dff_B_JzCAXZbT5_2),.dout(w_dff_B_z7HxxPCg7_2),.clk(gclk));
	jdff dff_B_7uNOedha2_2(.din(w_dff_B_z7HxxPCg7_2),.dout(w_dff_B_7uNOedha2_2),.clk(gclk));
	jdff dff_B_UZquPyqL3_2(.din(n990),.dout(w_dff_B_UZquPyqL3_2),.clk(gclk));
	jdff dff_B_RcaNpk1T7_1(.din(n960),.dout(w_dff_B_RcaNpk1T7_1),.clk(gclk));
	jdff dff_B_jyD9jlPS1_2(.din(n857),.dout(w_dff_B_jyD9jlPS1_2),.clk(gclk));
	jdff dff_B_M1MrszxR0_2(.din(w_dff_B_jyD9jlPS1_2),.dout(w_dff_B_M1MrszxR0_2),.clk(gclk));
	jdff dff_B_be2rJyGh9_2(.din(w_dff_B_M1MrszxR0_2),.dout(w_dff_B_be2rJyGh9_2),.clk(gclk));
	jdff dff_B_l1sSRFEA6_2(.din(w_dff_B_be2rJyGh9_2),.dout(w_dff_B_l1sSRFEA6_2),.clk(gclk));
	jdff dff_B_obOo6bfF4_2(.din(w_dff_B_l1sSRFEA6_2),.dout(w_dff_B_obOo6bfF4_2),.clk(gclk));
	jdff dff_B_Auk0EMZ11_2(.din(w_dff_B_obOo6bfF4_2),.dout(w_dff_B_Auk0EMZ11_2),.clk(gclk));
	jdff dff_B_pjGDfKvY6_2(.din(w_dff_B_Auk0EMZ11_2),.dout(w_dff_B_pjGDfKvY6_2),.clk(gclk));
	jdff dff_B_a3WcKyJ41_2(.din(w_dff_B_pjGDfKvY6_2),.dout(w_dff_B_a3WcKyJ41_2),.clk(gclk));
	jdff dff_B_6guXQXpl8_2(.din(w_dff_B_a3WcKyJ41_2),.dout(w_dff_B_6guXQXpl8_2),.clk(gclk));
	jdff dff_B_iDqmTMMw8_2(.din(w_dff_B_6guXQXpl8_2),.dout(w_dff_B_iDqmTMMw8_2),.clk(gclk));
	jdff dff_B_obKF3JNN7_2(.din(w_dff_B_iDqmTMMw8_2),.dout(w_dff_B_obKF3JNN7_2),.clk(gclk));
	jdff dff_B_c7kGDYuK5_2(.din(w_dff_B_obKF3JNN7_2),.dout(w_dff_B_c7kGDYuK5_2),.clk(gclk));
	jdff dff_B_2a9Kgfqe3_2(.din(w_dff_B_c7kGDYuK5_2),.dout(w_dff_B_2a9Kgfqe3_2),.clk(gclk));
	jdff dff_B_6GItylHC3_2(.din(w_dff_B_2a9Kgfqe3_2),.dout(w_dff_B_6GItylHC3_2),.clk(gclk));
	jdff dff_B_Wvs81bCN0_2(.din(n884),.dout(w_dff_B_Wvs81bCN0_2),.clk(gclk));
	jdff dff_B_3kdNpIDS2_1(.din(n858),.dout(w_dff_B_3kdNpIDS2_1),.clk(gclk));
	jdff dff_B_4UDEevnT5_2(.din(n759),.dout(w_dff_B_4UDEevnT5_2),.clk(gclk));
	jdff dff_B_uz8Ib7D22_2(.din(w_dff_B_4UDEevnT5_2),.dout(w_dff_B_uz8Ib7D22_2),.clk(gclk));
	jdff dff_B_qwaZHtGz0_2(.din(w_dff_B_uz8Ib7D22_2),.dout(w_dff_B_qwaZHtGz0_2),.clk(gclk));
	jdff dff_B_W3BAzdNv3_2(.din(w_dff_B_qwaZHtGz0_2),.dout(w_dff_B_W3BAzdNv3_2),.clk(gclk));
	jdff dff_B_ioPUdqXo0_2(.din(w_dff_B_W3BAzdNv3_2),.dout(w_dff_B_ioPUdqXo0_2),.clk(gclk));
	jdff dff_B_qJavXmVr2_2(.din(w_dff_B_ioPUdqXo0_2),.dout(w_dff_B_qJavXmVr2_2),.clk(gclk));
	jdff dff_B_6MfAlA2I6_2(.din(w_dff_B_qJavXmVr2_2),.dout(w_dff_B_6MfAlA2I6_2),.clk(gclk));
	jdff dff_B_pZG3zAAN2_2(.din(w_dff_B_6MfAlA2I6_2),.dout(w_dff_B_pZG3zAAN2_2),.clk(gclk));
	jdff dff_B_n3oivF5S0_2(.din(w_dff_B_pZG3zAAN2_2),.dout(w_dff_B_n3oivF5S0_2),.clk(gclk));
	jdff dff_B_RjfTGN7b6_2(.din(w_dff_B_n3oivF5S0_2),.dout(w_dff_B_RjfTGN7b6_2),.clk(gclk));
	jdff dff_B_XovSSTRy2_2(.din(w_dff_B_RjfTGN7b6_2),.dout(w_dff_B_XovSSTRy2_2),.clk(gclk));
	jdff dff_B_1s3Leg2W0_2(.din(n781),.dout(w_dff_B_1s3Leg2W0_2),.clk(gclk));
	jdff dff_B_58V6RV5c9_1(.din(n760),.dout(w_dff_B_58V6RV5c9_1),.clk(gclk));
	jdff dff_B_1DtK8UZq9_2(.din(n667),.dout(w_dff_B_1DtK8UZq9_2),.clk(gclk));
	jdff dff_B_hv0zbFXF1_2(.din(w_dff_B_1DtK8UZq9_2),.dout(w_dff_B_hv0zbFXF1_2),.clk(gclk));
	jdff dff_B_k0T8pjKR3_2(.din(w_dff_B_hv0zbFXF1_2),.dout(w_dff_B_k0T8pjKR3_2),.clk(gclk));
	jdff dff_B_JnbiRzxM6_2(.din(w_dff_B_k0T8pjKR3_2),.dout(w_dff_B_JnbiRzxM6_2),.clk(gclk));
	jdff dff_B_yve8NB3J4_2(.din(w_dff_B_JnbiRzxM6_2),.dout(w_dff_B_yve8NB3J4_2),.clk(gclk));
	jdff dff_B_eJDvWjLt3_2(.din(w_dff_B_yve8NB3J4_2),.dout(w_dff_B_eJDvWjLt3_2),.clk(gclk));
	jdff dff_B_aFnSAuSM5_2(.din(w_dff_B_eJDvWjLt3_2),.dout(w_dff_B_aFnSAuSM5_2),.clk(gclk));
	jdff dff_B_NcfWduB29_2(.din(w_dff_B_aFnSAuSM5_2),.dout(w_dff_B_NcfWduB29_2),.clk(gclk));
	jdff dff_B_uaazYh8H4_2(.din(n682),.dout(w_dff_B_uaazYh8H4_2),.clk(gclk));
	jdff dff_B_FR9pN9Gn5_2(.din(w_dff_B_uaazYh8H4_2),.dout(w_dff_B_FR9pN9Gn5_2),.clk(gclk));
	jdff dff_B_NnRZQt6k9_2(.din(w_dff_B_FR9pN9Gn5_2),.dout(w_dff_B_NnRZQt6k9_2),.clk(gclk));
	jdff dff_B_lctd7zUT2_1(.din(n668),.dout(w_dff_B_lctd7zUT2_1),.clk(gclk));
	jdff dff_B_sNSkNFS63_1(.din(w_dff_B_lctd7zUT2_1),.dout(w_dff_B_sNSkNFS63_1),.clk(gclk));
	jdff dff_B_OxJMzRfB7_2(.din(n584),.dout(w_dff_B_OxJMzRfB7_2),.clk(gclk));
	jdff dff_B_Ms7VltmA1_2(.din(w_dff_B_OxJMzRfB7_2),.dout(w_dff_B_Ms7VltmA1_2),.clk(gclk));
	jdff dff_B_t8ZJcDmB0_2(.din(w_dff_B_Ms7VltmA1_2),.dout(w_dff_B_t8ZJcDmB0_2),.clk(gclk));
	jdff dff_B_wGRbh8jc5_0(.din(n589),.dout(w_dff_B_wGRbh8jc5_0),.clk(gclk));
	jdff dff_A_io4gw1MZ2_0(.dout(w_n503_0[0]),.din(w_dff_A_io4gw1MZ2_0),.clk(gclk));
	jdff dff_A_t6iX48tA8_0(.dout(w_dff_A_io4gw1MZ2_0),.din(w_dff_A_t6iX48tA8_0),.clk(gclk));
	jdff dff_A_YF2EYJSt0_1(.dout(w_n503_0[1]),.din(w_dff_A_YF2EYJSt0_1),.clk(gclk));
	jdff dff_A_qZksD9iJ4_1(.dout(w_dff_A_YF2EYJSt0_1),.din(w_dff_A_qZksD9iJ4_1),.clk(gclk));
	jdff dff_B_BKablcen2_1(.din(n1762),.dout(w_dff_B_BKablcen2_1),.clk(gclk));
	jdff dff_A_bsSlG3hO7_1(.dout(w_n1737_0[1]),.din(w_dff_A_bsSlG3hO7_1),.clk(gclk));
	jdff dff_B_FcTF5d0h3_1(.din(n1735),.dout(w_dff_B_FcTF5d0h3_1),.clk(gclk));
	jdff dff_B_OUBhC1NO7_2(.din(n1699),.dout(w_dff_B_OUBhC1NO7_2),.clk(gclk));
	jdff dff_B_fmJtwFIt2_2(.din(w_dff_B_OUBhC1NO7_2),.dout(w_dff_B_fmJtwFIt2_2),.clk(gclk));
	jdff dff_B_ItwRgNHp0_2(.din(w_dff_B_fmJtwFIt2_2),.dout(w_dff_B_ItwRgNHp0_2),.clk(gclk));
	jdff dff_B_Pw74HCmk5_2(.din(w_dff_B_ItwRgNHp0_2),.dout(w_dff_B_Pw74HCmk5_2),.clk(gclk));
	jdff dff_B_whysWFLh7_2(.din(w_dff_B_Pw74HCmk5_2),.dout(w_dff_B_whysWFLh7_2),.clk(gclk));
	jdff dff_B_vFHUHe1I6_2(.din(w_dff_B_whysWFLh7_2),.dout(w_dff_B_vFHUHe1I6_2),.clk(gclk));
	jdff dff_B_dNBzMi9l1_2(.din(w_dff_B_vFHUHe1I6_2),.dout(w_dff_B_dNBzMi9l1_2),.clk(gclk));
	jdff dff_B_t4aK7ddr9_2(.din(w_dff_B_dNBzMi9l1_2),.dout(w_dff_B_t4aK7ddr9_2),.clk(gclk));
	jdff dff_B_VRfdxMMV1_2(.din(w_dff_B_t4aK7ddr9_2),.dout(w_dff_B_VRfdxMMV1_2),.clk(gclk));
	jdff dff_B_PANLaeBs9_2(.din(w_dff_B_VRfdxMMV1_2),.dout(w_dff_B_PANLaeBs9_2),.clk(gclk));
	jdff dff_B_lPWXXIzo8_2(.din(w_dff_B_PANLaeBs9_2),.dout(w_dff_B_lPWXXIzo8_2),.clk(gclk));
	jdff dff_B_M36Y5qE90_2(.din(w_dff_B_lPWXXIzo8_2),.dout(w_dff_B_M36Y5qE90_2),.clk(gclk));
	jdff dff_B_KfefUwkb1_2(.din(w_dff_B_M36Y5qE90_2),.dout(w_dff_B_KfefUwkb1_2),.clk(gclk));
	jdff dff_B_d71AzNVT2_2(.din(w_dff_B_KfefUwkb1_2),.dout(w_dff_B_d71AzNVT2_2),.clk(gclk));
	jdff dff_B_MMHvZwqM3_2(.din(w_dff_B_d71AzNVT2_2),.dout(w_dff_B_MMHvZwqM3_2),.clk(gclk));
	jdff dff_B_0mPgEUwx9_2(.din(w_dff_B_MMHvZwqM3_2),.dout(w_dff_B_0mPgEUwx9_2),.clk(gclk));
	jdff dff_B_5VK78K6H1_2(.din(w_dff_B_0mPgEUwx9_2),.dout(w_dff_B_5VK78K6H1_2),.clk(gclk));
	jdff dff_B_TP73D6c32_2(.din(w_dff_B_5VK78K6H1_2),.dout(w_dff_B_TP73D6c32_2),.clk(gclk));
	jdff dff_B_lBaP8azp5_2(.din(w_dff_B_TP73D6c32_2),.dout(w_dff_B_lBaP8azp5_2),.clk(gclk));
	jdff dff_B_Uvkgl5ZA7_2(.din(w_dff_B_lBaP8azp5_2),.dout(w_dff_B_Uvkgl5ZA7_2),.clk(gclk));
	jdff dff_B_n4ysy3ao2_2(.din(w_dff_B_Uvkgl5ZA7_2),.dout(w_dff_B_n4ysy3ao2_2),.clk(gclk));
	jdff dff_B_g4XX9DeR3_2(.din(w_dff_B_n4ysy3ao2_2),.dout(w_dff_B_g4XX9DeR3_2),.clk(gclk));
	jdff dff_B_Ov3UanVv7_2(.din(w_dff_B_g4XX9DeR3_2),.dout(w_dff_B_Ov3UanVv7_2),.clk(gclk));
	jdff dff_B_FD0NL8Vi5_2(.din(w_dff_B_Ov3UanVv7_2),.dout(w_dff_B_FD0NL8Vi5_2),.clk(gclk));
	jdff dff_B_VwtkVktY9_2(.din(w_dff_B_FD0NL8Vi5_2),.dout(w_dff_B_VwtkVktY9_2),.clk(gclk));
	jdff dff_B_ZRWJtusi2_2(.din(w_dff_B_VwtkVktY9_2),.dout(w_dff_B_ZRWJtusi2_2),.clk(gclk));
	jdff dff_B_ipL11gTl0_2(.din(w_dff_B_ZRWJtusi2_2),.dout(w_dff_B_ipL11gTl0_2),.clk(gclk));
	jdff dff_B_YJxHvJrQ8_2(.din(w_dff_B_ipL11gTl0_2),.dout(w_dff_B_YJxHvJrQ8_2),.clk(gclk));
	jdff dff_B_sFVwPFI35_2(.din(w_dff_B_YJxHvJrQ8_2),.dout(w_dff_B_sFVwPFI35_2),.clk(gclk));
	jdff dff_B_ZQKVMXdx0_2(.din(w_dff_B_sFVwPFI35_2),.dout(w_dff_B_ZQKVMXdx0_2),.clk(gclk));
	jdff dff_B_EAc4G7fo3_2(.din(w_dff_B_ZQKVMXdx0_2),.dout(w_dff_B_EAc4G7fo3_2),.clk(gclk));
	jdff dff_B_QM6cG2iy0_2(.din(w_dff_B_EAc4G7fo3_2),.dout(w_dff_B_QM6cG2iy0_2),.clk(gclk));
	jdff dff_B_UkqzuT5k3_2(.din(w_dff_B_QM6cG2iy0_2),.dout(w_dff_B_UkqzuT5k3_2),.clk(gclk));
	jdff dff_B_J0lgCcYt9_2(.din(w_dff_B_UkqzuT5k3_2),.dout(w_dff_B_J0lgCcYt9_2),.clk(gclk));
	jdff dff_B_hQQo2If56_2(.din(w_dff_B_J0lgCcYt9_2),.dout(w_dff_B_hQQo2If56_2),.clk(gclk));
	jdff dff_B_2mlZENjF0_2(.din(w_dff_B_hQQo2If56_2),.dout(w_dff_B_2mlZENjF0_2),.clk(gclk));
	jdff dff_B_khVW1U4E7_2(.din(w_dff_B_2mlZENjF0_2),.dout(w_dff_B_khVW1U4E7_2),.clk(gclk));
	jdff dff_B_26yFExap6_2(.din(w_dff_B_khVW1U4E7_2),.dout(w_dff_B_26yFExap6_2),.clk(gclk));
	jdff dff_B_gxIDlyg10_2(.din(w_dff_B_26yFExap6_2),.dout(w_dff_B_gxIDlyg10_2),.clk(gclk));
	jdff dff_B_HfKV2YGx6_2(.din(w_dff_B_gxIDlyg10_2),.dout(w_dff_B_HfKV2YGx6_2),.clk(gclk));
	jdff dff_B_F85Oe1U58_2(.din(w_dff_B_HfKV2YGx6_2),.dout(w_dff_B_F85Oe1U58_2),.clk(gclk));
	jdff dff_B_Dq8tn5gX4_2(.din(w_dff_B_F85Oe1U58_2),.dout(w_dff_B_Dq8tn5gX4_2),.clk(gclk));
	jdff dff_B_ude87cpT0_2(.din(w_dff_B_Dq8tn5gX4_2),.dout(w_dff_B_ude87cpT0_2),.clk(gclk));
	jdff dff_B_T19x75My6_2(.din(w_dff_B_ude87cpT0_2),.dout(w_dff_B_T19x75My6_2),.clk(gclk));
	jdff dff_B_QhLcJXdJ5_2(.din(w_dff_B_T19x75My6_2),.dout(w_dff_B_QhLcJXdJ5_2),.clk(gclk));
	jdff dff_B_VYjkvQDf1_2(.din(w_dff_B_QhLcJXdJ5_2),.dout(w_dff_B_VYjkvQDf1_2),.clk(gclk));
	jdff dff_B_UTmKQY3Q3_2(.din(w_dff_B_VYjkvQDf1_2),.dout(w_dff_B_UTmKQY3Q3_2),.clk(gclk));
	jdff dff_B_a2Kjpush8_2(.din(w_dff_B_UTmKQY3Q3_2),.dout(w_dff_B_a2Kjpush8_2),.clk(gclk));
	jdff dff_B_YwNIF9Vn6_2(.din(n1702),.dout(w_dff_B_YwNIF9Vn6_2),.clk(gclk));
	jdff dff_B_jjFo3b7d1_1(.din(n1700),.dout(w_dff_B_jjFo3b7d1_1),.clk(gclk));
	jdff dff_B_eHB6nEBG0_2(.din(n1658),.dout(w_dff_B_eHB6nEBG0_2),.clk(gclk));
	jdff dff_B_CHEiYN1l4_2(.din(w_dff_B_eHB6nEBG0_2),.dout(w_dff_B_CHEiYN1l4_2),.clk(gclk));
	jdff dff_B_72yhTXIg5_2(.din(w_dff_B_CHEiYN1l4_2),.dout(w_dff_B_72yhTXIg5_2),.clk(gclk));
	jdff dff_B_4La54H0s1_2(.din(w_dff_B_72yhTXIg5_2),.dout(w_dff_B_4La54H0s1_2),.clk(gclk));
	jdff dff_B_RtkH3Ulv6_2(.din(w_dff_B_4La54H0s1_2),.dout(w_dff_B_RtkH3Ulv6_2),.clk(gclk));
	jdff dff_B_6Yrhcs9R7_2(.din(w_dff_B_RtkH3Ulv6_2),.dout(w_dff_B_6Yrhcs9R7_2),.clk(gclk));
	jdff dff_B_Sq5xUdzH9_2(.din(w_dff_B_6Yrhcs9R7_2),.dout(w_dff_B_Sq5xUdzH9_2),.clk(gclk));
	jdff dff_B_uMw4oF765_2(.din(w_dff_B_Sq5xUdzH9_2),.dout(w_dff_B_uMw4oF765_2),.clk(gclk));
	jdff dff_B_kNMwuPsa4_2(.din(w_dff_B_uMw4oF765_2),.dout(w_dff_B_kNMwuPsa4_2),.clk(gclk));
	jdff dff_B_UHhjEkkI4_2(.din(w_dff_B_kNMwuPsa4_2),.dout(w_dff_B_UHhjEkkI4_2),.clk(gclk));
	jdff dff_B_9d4qtsyr5_2(.din(w_dff_B_UHhjEkkI4_2),.dout(w_dff_B_9d4qtsyr5_2),.clk(gclk));
	jdff dff_B_z06po0zU3_2(.din(w_dff_B_9d4qtsyr5_2),.dout(w_dff_B_z06po0zU3_2),.clk(gclk));
	jdff dff_B_VaWOY6TC8_2(.din(w_dff_B_z06po0zU3_2),.dout(w_dff_B_VaWOY6TC8_2),.clk(gclk));
	jdff dff_B_mwnjfS311_2(.din(w_dff_B_VaWOY6TC8_2),.dout(w_dff_B_mwnjfS311_2),.clk(gclk));
	jdff dff_B_ImxED3zz2_2(.din(w_dff_B_mwnjfS311_2),.dout(w_dff_B_ImxED3zz2_2),.clk(gclk));
	jdff dff_B_UEAyJW5l1_2(.din(w_dff_B_ImxED3zz2_2),.dout(w_dff_B_UEAyJW5l1_2),.clk(gclk));
	jdff dff_B_guwLKsvS8_2(.din(w_dff_B_UEAyJW5l1_2),.dout(w_dff_B_guwLKsvS8_2),.clk(gclk));
	jdff dff_B_sHHvjsPS6_2(.din(w_dff_B_guwLKsvS8_2),.dout(w_dff_B_sHHvjsPS6_2),.clk(gclk));
	jdff dff_B_qzHT2KNb3_2(.din(w_dff_B_sHHvjsPS6_2),.dout(w_dff_B_qzHT2KNb3_2),.clk(gclk));
	jdff dff_B_ocGRKwGS9_2(.din(w_dff_B_qzHT2KNb3_2),.dout(w_dff_B_ocGRKwGS9_2),.clk(gclk));
	jdff dff_B_rnd3yGtu5_2(.din(w_dff_B_ocGRKwGS9_2),.dout(w_dff_B_rnd3yGtu5_2),.clk(gclk));
	jdff dff_B_t7kK7vpJ3_2(.din(w_dff_B_rnd3yGtu5_2),.dout(w_dff_B_t7kK7vpJ3_2),.clk(gclk));
	jdff dff_B_khTexeY66_2(.din(w_dff_B_t7kK7vpJ3_2),.dout(w_dff_B_khTexeY66_2),.clk(gclk));
	jdff dff_B_AP9FniQL4_2(.din(w_dff_B_khTexeY66_2),.dout(w_dff_B_AP9FniQL4_2),.clk(gclk));
	jdff dff_B_2CZ094Zn5_2(.din(w_dff_B_AP9FniQL4_2),.dout(w_dff_B_2CZ094Zn5_2),.clk(gclk));
	jdff dff_B_g0ETjYvw9_2(.din(w_dff_B_2CZ094Zn5_2),.dout(w_dff_B_g0ETjYvw9_2),.clk(gclk));
	jdff dff_B_wGwYkgyp5_2(.din(w_dff_B_g0ETjYvw9_2),.dout(w_dff_B_wGwYkgyp5_2),.clk(gclk));
	jdff dff_B_TXFvDDTV0_2(.din(w_dff_B_wGwYkgyp5_2),.dout(w_dff_B_TXFvDDTV0_2),.clk(gclk));
	jdff dff_B_gnDsqmLA8_2(.din(w_dff_B_TXFvDDTV0_2),.dout(w_dff_B_gnDsqmLA8_2),.clk(gclk));
	jdff dff_B_lxBOVhXB5_2(.din(w_dff_B_gnDsqmLA8_2),.dout(w_dff_B_lxBOVhXB5_2),.clk(gclk));
	jdff dff_B_WrAUXnFC0_2(.din(w_dff_B_lxBOVhXB5_2),.dout(w_dff_B_WrAUXnFC0_2),.clk(gclk));
	jdff dff_B_E27KxMi70_2(.din(w_dff_B_WrAUXnFC0_2),.dout(w_dff_B_E27KxMi70_2),.clk(gclk));
	jdff dff_B_7zabKwqo9_2(.din(w_dff_B_E27KxMi70_2),.dout(w_dff_B_7zabKwqo9_2),.clk(gclk));
	jdff dff_B_HeJAS2282_2(.din(w_dff_B_7zabKwqo9_2),.dout(w_dff_B_HeJAS2282_2),.clk(gclk));
	jdff dff_B_7tKD9LPK4_2(.din(w_dff_B_HeJAS2282_2),.dout(w_dff_B_7tKD9LPK4_2),.clk(gclk));
	jdff dff_B_W9udXep88_2(.din(w_dff_B_7tKD9LPK4_2),.dout(w_dff_B_W9udXep88_2),.clk(gclk));
	jdff dff_B_iMWVDoie5_2(.din(w_dff_B_W9udXep88_2),.dout(w_dff_B_iMWVDoie5_2),.clk(gclk));
	jdff dff_B_Gi4ooOp19_2(.din(w_dff_B_iMWVDoie5_2),.dout(w_dff_B_Gi4ooOp19_2),.clk(gclk));
	jdff dff_B_UP7BAiTN3_2(.din(w_dff_B_Gi4ooOp19_2),.dout(w_dff_B_UP7BAiTN3_2),.clk(gclk));
	jdff dff_B_H4cSGW3E7_2(.din(w_dff_B_UP7BAiTN3_2),.dout(w_dff_B_H4cSGW3E7_2),.clk(gclk));
	jdff dff_B_46d62AYL0_2(.din(w_dff_B_H4cSGW3E7_2),.dout(w_dff_B_46d62AYL0_2),.clk(gclk));
	jdff dff_B_PL5uDZ9L5_2(.din(w_dff_B_46d62AYL0_2),.dout(w_dff_B_PL5uDZ9L5_2),.clk(gclk));
	jdff dff_B_v7fAg0fD1_2(.din(w_dff_B_PL5uDZ9L5_2),.dout(w_dff_B_v7fAg0fD1_2),.clk(gclk));
	jdff dff_B_9Pq9g6YL3_2(.din(w_dff_B_v7fAg0fD1_2),.dout(w_dff_B_9Pq9g6YL3_2),.clk(gclk));
	jdff dff_B_mPJtTvrl4_2(.din(n1661),.dout(w_dff_B_mPJtTvrl4_2),.clk(gclk));
	jdff dff_B_J1dXw1Si3_1(.din(n1659),.dout(w_dff_B_J1dXw1Si3_1),.clk(gclk));
	jdff dff_B_DEXGpvSM7_2(.din(n1607),.dout(w_dff_B_DEXGpvSM7_2),.clk(gclk));
	jdff dff_B_eFLJveyf3_2(.din(w_dff_B_DEXGpvSM7_2),.dout(w_dff_B_eFLJveyf3_2),.clk(gclk));
	jdff dff_B_bOCPJfyW8_2(.din(w_dff_B_eFLJveyf3_2),.dout(w_dff_B_bOCPJfyW8_2),.clk(gclk));
	jdff dff_B_36b6XdMD6_2(.din(w_dff_B_bOCPJfyW8_2),.dout(w_dff_B_36b6XdMD6_2),.clk(gclk));
	jdff dff_B_pdwZLhvl3_2(.din(w_dff_B_36b6XdMD6_2),.dout(w_dff_B_pdwZLhvl3_2),.clk(gclk));
	jdff dff_B_odG7Wl2P6_2(.din(w_dff_B_pdwZLhvl3_2),.dout(w_dff_B_odG7Wl2P6_2),.clk(gclk));
	jdff dff_B_2sxTNxK93_2(.din(w_dff_B_odG7Wl2P6_2),.dout(w_dff_B_2sxTNxK93_2),.clk(gclk));
	jdff dff_B_5HARTNgB6_2(.din(w_dff_B_2sxTNxK93_2),.dout(w_dff_B_5HARTNgB6_2),.clk(gclk));
	jdff dff_B_YqYrLMvF8_2(.din(w_dff_B_5HARTNgB6_2),.dout(w_dff_B_YqYrLMvF8_2),.clk(gclk));
	jdff dff_B_G9TyQWZW5_2(.din(w_dff_B_YqYrLMvF8_2),.dout(w_dff_B_G9TyQWZW5_2),.clk(gclk));
	jdff dff_B_JSaBwnQg6_2(.din(w_dff_B_G9TyQWZW5_2),.dout(w_dff_B_JSaBwnQg6_2),.clk(gclk));
	jdff dff_B_DbpJXVVX7_2(.din(w_dff_B_JSaBwnQg6_2),.dout(w_dff_B_DbpJXVVX7_2),.clk(gclk));
	jdff dff_B_fHojTLNq4_2(.din(w_dff_B_DbpJXVVX7_2),.dout(w_dff_B_fHojTLNq4_2),.clk(gclk));
	jdff dff_B_5jDJJQiJ9_2(.din(w_dff_B_fHojTLNq4_2),.dout(w_dff_B_5jDJJQiJ9_2),.clk(gclk));
	jdff dff_B_N384otp13_2(.din(w_dff_B_5jDJJQiJ9_2),.dout(w_dff_B_N384otp13_2),.clk(gclk));
	jdff dff_B_zWavUoES0_2(.din(w_dff_B_N384otp13_2),.dout(w_dff_B_zWavUoES0_2),.clk(gclk));
	jdff dff_B_eku0LzPZ7_2(.din(w_dff_B_zWavUoES0_2),.dout(w_dff_B_eku0LzPZ7_2),.clk(gclk));
	jdff dff_B_VFJ0Nj5D8_2(.din(w_dff_B_eku0LzPZ7_2),.dout(w_dff_B_VFJ0Nj5D8_2),.clk(gclk));
	jdff dff_B_lYXCGiOs8_2(.din(w_dff_B_VFJ0Nj5D8_2),.dout(w_dff_B_lYXCGiOs8_2),.clk(gclk));
	jdff dff_B_6ZsLZ4wK5_2(.din(w_dff_B_lYXCGiOs8_2),.dout(w_dff_B_6ZsLZ4wK5_2),.clk(gclk));
	jdff dff_B_LVfbHczP4_2(.din(w_dff_B_6ZsLZ4wK5_2),.dout(w_dff_B_LVfbHczP4_2),.clk(gclk));
	jdff dff_B_0uX0iXsO9_2(.din(w_dff_B_LVfbHczP4_2),.dout(w_dff_B_0uX0iXsO9_2),.clk(gclk));
	jdff dff_B_hNUFNmTL6_2(.din(w_dff_B_0uX0iXsO9_2),.dout(w_dff_B_hNUFNmTL6_2),.clk(gclk));
	jdff dff_B_nVotZP695_2(.din(w_dff_B_hNUFNmTL6_2),.dout(w_dff_B_nVotZP695_2),.clk(gclk));
	jdff dff_B_p8pibRlP1_2(.din(w_dff_B_nVotZP695_2),.dout(w_dff_B_p8pibRlP1_2),.clk(gclk));
	jdff dff_B_5gPiEYGt8_2(.din(w_dff_B_p8pibRlP1_2),.dout(w_dff_B_5gPiEYGt8_2),.clk(gclk));
	jdff dff_B_xHWM1olY6_2(.din(w_dff_B_5gPiEYGt8_2),.dout(w_dff_B_xHWM1olY6_2),.clk(gclk));
	jdff dff_B_Si4HnNJr4_2(.din(w_dff_B_xHWM1olY6_2),.dout(w_dff_B_Si4HnNJr4_2),.clk(gclk));
	jdff dff_B_vsiNTbZV0_2(.din(w_dff_B_Si4HnNJr4_2),.dout(w_dff_B_vsiNTbZV0_2),.clk(gclk));
	jdff dff_B_2mmrACs66_2(.din(w_dff_B_vsiNTbZV0_2),.dout(w_dff_B_2mmrACs66_2),.clk(gclk));
	jdff dff_B_Yd0GGByz4_2(.din(w_dff_B_2mmrACs66_2),.dout(w_dff_B_Yd0GGByz4_2),.clk(gclk));
	jdff dff_B_Lcm8LdNh2_2(.din(w_dff_B_Yd0GGByz4_2),.dout(w_dff_B_Lcm8LdNh2_2),.clk(gclk));
	jdff dff_B_SAlxpB8D1_2(.din(w_dff_B_Lcm8LdNh2_2),.dout(w_dff_B_SAlxpB8D1_2),.clk(gclk));
	jdff dff_B_x34HdRjl9_2(.din(w_dff_B_SAlxpB8D1_2),.dout(w_dff_B_x34HdRjl9_2),.clk(gclk));
	jdff dff_B_XrvjAUW74_2(.din(w_dff_B_x34HdRjl9_2),.dout(w_dff_B_XrvjAUW74_2),.clk(gclk));
	jdff dff_B_fxaBQXP27_2(.din(w_dff_B_XrvjAUW74_2),.dout(w_dff_B_fxaBQXP27_2),.clk(gclk));
	jdff dff_B_MHLn6Nhr9_2(.din(w_dff_B_fxaBQXP27_2),.dout(w_dff_B_MHLn6Nhr9_2),.clk(gclk));
	jdff dff_B_pKNsPfbR9_2(.din(w_dff_B_MHLn6Nhr9_2),.dout(w_dff_B_pKNsPfbR9_2),.clk(gclk));
	jdff dff_B_J5dSF4jh3_2(.din(w_dff_B_pKNsPfbR9_2),.dout(w_dff_B_J5dSF4jh3_2),.clk(gclk));
	jdff dff_B_NWclf5rq6_2(.din(w_dff_B_J5dSF4jh3_2),.dout(w_dff_B_NWclf5rq6_2),.clk(gclk));
	jdff dff_B_s48Z0v4b3_2(.din(n1610),.dout(w_dff_B_s48Z0v4b3_2),.clk(gclk));
	jdff dff_B_NToFGzAQ7_1(.din(n1608),.dout(w_dff_B_NToFGzAQ7_1),.clk(gclk));
	jdff dff_B_vJXJgwPJ0_2(.din(n1550),.dout(w_dff_B_vJXJgwPJ0_2),.clk(gclk));
	jdff dff_B_CVcrzpfv7_2(.din(w_dff_B_vJXJgwPJ0_2),.dout(w_dff_B_CVcrzpfv7_2),.clk(gclk));
	jdff dff_B_nQi6u14K6_2(.din(w_dff_B_CVcrzpfv7_2),.dout(w_dff_B_nQi6u14K6_2),.clk(gclk));
	jdff dff_B_x120Z6yC1_2(.din(w_dff_B_nQi6u14K6_2),.dout(w_dff_B_x120Z6yC1_2),.clk(gclk));
	jdff dff_B_NM3kxtf45_2(.din(w_dff_B_x120Z6yC1_2),.dout(w_dff_B_NM3kxtf45_2),.clk(gclk));
	jdff dff_B_ATZybB8C1_2(.din(w_dff_B_NM3kxtf45_2),.dout(w_dff_B_ATZybB8C1_2),.clk(gclk));
	jdff dff_B_iIPdcsum9_2(.din(w_dff_B_ATZybB8C1_2),.dout(w_dff_B_iIPdcsum9_2),.clk(gclk));
	jdff dff_B_B2ObvuDJ1_2(.din(w_dff_B_iIPdcsum9_2),.dout(w_dff_B_B2ObvuDJ1_2),.clk(gclk));
	jdff dff_B_mB0evKK29_2(.din(w_dff_B_B2ObvuDJ1_2),.dout(w_dff_B_mB0evKK29_2),.clk(gclk));
	jdff dff_B_z25aOPCP0_2(.din(w_dff_B_mB0evKK29_2),.dout(w_dff_B_z25aOPCP0_2),.clk(gclk));
	jdff dff_B_mCc2ME7p8_2(.din(w_dff_B_z25aOPCP0_2),.dout(w_dff_B_mCc2ME7p8_2),.clk(gclk));
	jdff dff_B_1UZJbKRA5_2(.din(w_dff_B_mCc2ME7p8_2),.dout(w_dff_B_1UZJbKRA5_2),.clk(gclk));
	jdff dff_B_4kijFdoW6_2(.din(w_dff_B_1UZJbKRA5_2),.dout(w_dff_B_4kijFdoW6_2),.clk(gclk));
	jdff dff_B_l6Z6BXob2_2(.din(w_dff_B_4kijFdoW6_2),.dout(w_dff_B_l6Z6BXob2_2),.clk(gclk));
	jdff dff_B_CZOEVuH90_2(.din(w_dff_B_l6Z6BXob2_2),.dout(w_dff_B_CZOEVuH90_2),.clk(gclk));
	jdff dff_B_TY7LN03v8_2(.din(w_dff_B_CZOEVuH90_2),.dout(w_dff_B_TY7LN03v8_2),.clk(gclk));
	jdff dff_B_CYochupi6_2(.din(w_dff_B_TY7LN03v8_2),.dout(w_dff_B_CYochupi6_2),.clk(gclk));
	jdff dff_B_F2Boja8F4_2(.din(w_dff_B_CYochupi6_2),.dout(w_dff_B_F2Boja8F4_2),.clk(gclk));
	jdff dff_B_ssP6s4HK2_2(.din(w_dff_B_F2Boja8F4_2),.dout(w_dff_B_ssP6s4HK2_2),.clk(gclk));
	jdff dff_B_t20TExDa2_2(.din(w_dff_B_ssP6s4HK2_2),.dout(w_dff_B_t20TExDa2_2),.clk(gclk));
	jdff dff_B_ClGlmacp8_2(.din(w_dff_B_t20TExDa2_2),.dout(w_dff_B_ClGlmacp8_2),.clk(gclk));
	jdff dff_B_94sdIFXV0_2(.din(w_dff_B_ClGlmacp8_2),.dout(w_dff_B_94sdIFXV0_2),.clk(gclk));
	jdff dff_B_StdHmQqc6_2(.din(w_dff_B_94sdIFXV0_2),.dout(w_dff_B_StdHmQqc6_2),.clk(gclk));
	jdff dff_B_5yjgYhqu5_2(.din(w_dff_B_StdHmQqc6_2),.dout(w_dff_B_5yjgYhqu5_2),.clk(gclk));
	jdff dff_B_fca5CBu10_2(.din(w_dff_B_5yjgYhqu5_2),.dout(w_dff_B_fca5CBu10_2),.clk(gclk));
	jdff dff_B_p3NBk60j6_2(.din(w_dff_B_fca5CBu10_2),.dout(w_dff_B_p3NBk60j6_2),.clk(gclk));
	jdff dff_B_0ToTjtN56_2(.din(w_dff_B_p3NBk60j6_2),.dout(w_dff_B_0ToTjtN56_2),.clk(gclk));
	jdff dff_B_wn77oDMg1_2(.din(w_dff_B_0ToTjtN56_2),.dout(w_dff_B_wn77oDMg1_2),.clk(gclk));
	jdff dff_B_OwSITP280_2(.din(w_dff_B_wn77oDMg1_2),.dout(w_dff_B_OwSITP280_2),.clk(gclk));
	jdff dff_B_sjpAV16v1_2(.din(w_dff_B_OwSITP280_2),.dout(w_dff_B_sjpAV16v1_2),.clk(gclk));
	jdff dff_B_AfNT8kK71_2(.din(w_dff_B_sjpAV16v1_2),.dout(w_dff_B_AfNT8kK71_2),.clk(gclk));
	jdff dff_B_6h4ar9Ku6_2(.din(w_dff_B_AfNT8kK71_2),.dout(w_dff_B_6h4ar9Ku6_2),.clk(gclk));
	jdff dff_B_iJiDvakS7_2(.din(w_dff_B_6h4ar9Ku6_2),.dout(w_dff_B_iJiDvakS7_2),.clk(gclk));
	jdff dff_B_ZebamhUt0_2(.din(w_dff_B_iJiDvakS7_2),.dout(w_dff_B_ZebamhUt0_2),.clk(gclk));
	jdff dff_B_qgPNeUjA1_2(.din(w_dff_B_ZebamhUt0_2),.dout(w_dff_B_qgPNeUjA1_2),.clk(gclk));
	jdff dff_B_7fjS4I5R0_2(.din(w_dff_B_qgPNeUjA1_2),.dout(w_dff_B_7fjS4I5R0_2),.clk(gclk));
	jdff dff_B_t8ZmUGWO1_2(.din(n1553),.dout(w_dff_B_t8ZmUGWO1_2),.clk(gclk));
	jdff dff_B_Q7YT2tXl2_1(.din(n1551),.dout(w_dff_B_Q7YT2tXl2_1),.clk(gclk));
	jdff dff_B_WYVJMJUn5_2(.din(n1486),.dout(w_dff_B_WYVJMJUn5_2),.clk(gclk));
	jdff dff_B_ScVhj7am9_2(.din(w_dff_B_WYVJMJUn5_2),.dout(w_dff_B_ScVhj7am9_2),.clk(gclk));
	jdff dff_B_ViNS0e246_2(.din(w_dff_B_ScVhj7am9_2),.dout(w_dff_B_ViNS0e246_2),.clk(gclk));
	jdff dff_B_plE4owDJ0_2(.din(w_dff_B_ViNS0e246_2),.dout(w_dff_B_plE4owDJ0_2),.clk(gclk));
	jdff dff_B_hfQVAflm3_2(.din(w_dff_B_plE4owDJ0_2),.dout(w_dff_B_hfQVAflm3_2),.clk(gclk));
	jdff dff_B_BhI42FS42_2(.din(w_dff_B_hfQVAflm3_2),.dout(w_dff_B_BhI42FS42_2),.clk(gclk));
	jdff dff_B_npJAnwln5_2(.din(w_dff_B_BhI42FS42_2),.dout(w_dff_B_npJAnwln5_2),.clk(gclk));
	jdff dff_B_iRAuH4e56_2(.din(w_dff_B_npJAnwln5_2),.dout(w_dff_B_iRAuH4e56_2),.clk(gclk));
	jdff dff_B_Y0uNT97w2_2(.din(w_dff_B_iRAuH4e56_2),.dout(w_dff_B_Y0uNT97w2_2),.clk(gclk));
	jdff dff_B_c0z3FUhU2_2(.din(w_dff_B_Y0uNT97w2_2),.dout(w_dff_B_c0z3FUhU2_2),.clk(gclk));
	jdff dff_B_uNIK081t0_2(.din(w_dff_B_c0z3FUhU2_2),.dout(w_dff_B_uNIK081t0_2),.clk(gclk));
	jdff dff_B_6LMh9R2C2_2(.din(w_dff_B_uNIK081t0_2),.dout(w_dff_B_6LMh9R2C2_2),.clk(gclk));
	jdff dff_B_ZuJihfnl6_2(.din(w_dff_B_6LMh9R2C2_2),.dout(w_dff_B_ZuJihfnl6_2),.clk(gclk));
	jdff dff_B_yWFHp9fQ3_2(.din(w_dff_B_ZuJihfnl6_2),.dout(w_dff_B_yWFHp9fQ3_2),.clk(gclk));
	jdff dff_B_vLvjLSms5_2(.din(w_dff_B_yWFHp9fQ3_2),.dout(w_dff_B_vLvjLSms5_2),.clk(gclk));
	jdff dff_B_iUJ8DrRb0_2(.din(w_dff_B_vLvjLSms5_2),.dout(w_dff_B_iUJ8DrRb0_2),.clk(gclk));
	jdff dff_B_cCIonvuG0_2(.din(w_dff_B_iUJ8DrRb0_2),.dout(w_dff_B_cCIonvuG0_2),.clk(gclk));
	jdff dff_B_EoGS1bbT2_2(.din(w_dff_B_cCIonvuG0_2),.dout(w_dff_B_EoGS1bbT2_2),.clk(gclk));
	jdff dff_B_qRhLGgjD0_2(.din(w_dff_B_EoGS1bbT2_2),.dout(w_dff_B_qRhLGgjD0_2),.clk(gclk));
	jdff dff_B_BjXSP8lL4_2(.din(w_dff_B_qRhLGgjD0_2),.dout(w_dff_B_BjXSP8lL4_2),.clk(gclk));
	jdff dff_B_eA1aXsB79_2(.din(w_dff_B_BjXSP8lL4_2),.dout(w_dff_B_eA1aXsB79_2),.clk(gclk));
	jdff dff_B_DnIDgaQK8_2(.din(w_dff_B_eA1aXsB79_2),.dout(w_dff_B_DnIDgaQK8_2),.clk(gclk));
	jdff dff_B_2kSrcUO43_2(.din(w_dff_B_DnIDgaQK8_2),.dout(w_dff_B_2kSrcUO43_2),.clk(gclk));
	jdff dff_B_E8yQ1OjJ7_2(.din(w_dff_B_2kSrcUO43_2),.dout(w_dff_B_E8yQ1OjJ7_2),.clk(gclk));
	jdff dff_B_bSLruTOz6_2(.din(w_dff_B_E8yQ1OjJ7_2),.dout(w_dff_B_bSLruTOz6_2),.clk(gclk));
	jdff dff_B_OJt0hsBe1_2(.din(w_dff_B_bSLruTOz6_2),.dout(w_dff_B_OJt0hsBe1_2),.clk(gclk));
	jdff dff_B_eJJuzPRJ5_2(.din(w_dff_B_OJt0hsBe1_2),.dout(w_dff_B_eJJuzPRJ5_2),.clk(gclk));
	jdff dff_B_CpjqXGqa7_2(.din(w_dff_B_eJJuzPRJ5_2),.dout(w_dff_B_CpjqXGqa7_2),.clk(gclk));
	jdff dff_B_FhCzXo9Y4_2(.din(w_dff_B_CpjqXGqa7_2),.dout(w_dff_B_FhCzXo9Y4_2),.clk(gclk));
	jdff dff_B_oCKEaP5c6_2(.din(w_dff_B_FhCzXo9Y4_2),.dout(w_dff_B_oCKEaP5c6_2),.clk(gclk));
	jdff dff_B_FbhpoCpu2_2(.din(w_dff_B_oCKEaP5c6_2),.dout(w_dff_B_FbhpoCpu2_2),.clk(gclk));
	jdff dff_B_JzzDAZy18_2(.din(w_dff_B_FbhpoCpu2_2),.dout(w_dff_B_JzzDAZy18_2),.clk(gclk));
	jdff dff_B_KqDwvtXB8_1(.din(n1487),.dout(w_dff_B_KqDwvtXB8_1),.clk(gclk));
	jdff dff_B_4MW1dy5I3_2(.din(n1415),.dout(w_dff_B_4MW1dy5I3_2),.clk(gclk));
	jdff dff_B_xBzRkKfh2_2(.din(w_dff_B_4MW1dy5I3_2),.dout(w_dff_B_xBzRkKfh2_2),.clk(gclk));
	jdff dff_B_tOcnGwwS4_2(.din(w_dff_B_xBzRkKfh2_2),.dout(w_dff_B_tOcnGwwS4_2),.clk(gclk));
	jdff dff_B_CuP3tzkD3_2(.din(w_dff_B_tOcnGwwS4_2),.dout(w_dff_B_CuP3tzkD3_2),.clk(gclk));
	jdff dff_B_ePe6b4s39_2(.din(w_dff_B_CuP3tzkD3_2),.dout(w_dff_B_ePe6b4s39_2),.clk(gclk));
	jdff dff_B_KCEdPDOJ8_2(.din(w_dff_B_ePe6b4s39_2),.dout(w_dff_B_KCEdPDOJ8_2),.clk(gclk));
	jdff dff_B_kjyESEy86_2(.din(w_dff_B_KCEdPDOJ8_2),.dout(w_dff_B_kjyESEy86_2),.clk(gclk));
	jdff dff_B_Cwx4TogP5_2(.din(w_dff_B_kjyESEy86_2),.dout(w_dff_B_Cwx4TogP5_2),.clk(gclk));
	jdff dff_B_XOyxlPop0_2(.din(w_dff_B_Cwx4TogP5_2),.dout(w_dff_B_XOyxlPop0_2),.clk(gclk));
	jdff dff_B_SUnJpseU0_2(.din(w_dff_B_XOyxlPop0_2),.dout(w_dff_B_SUnJpseU0_2),.clk(gclk));
	jdff dff_B_Ad940SHD2_2(.din(w_dff_B_SUnJpseU0_2),.dout(w_dff_B_Ad940SHD2_2),.clk(gclk));
	jdff dff_B_sDMmGItq3_2(.din(w_dff_B_Ad940SHD2_2),.dout(w_dff_B_sDMmGItq3_2),.clk(gclk));
	jdff dff_B_xQwMSEmP7_2(.din(w_dff_B_sDMmGItq3_2),.dout(w_dff_B_xQwMSEmP7_2),.clk(gclk));
	jdff dff_B_TZq1nyMg9_2(.din(w_dff_B_xQwMSEmP7_2),.dout(w_dff_B_TZq1nyMg9_2),.clk(gclk));
	jdff dff_B_GoF85LcZ0_2(.din(w_dff_B_TZq1nyMg9_2),.dout(w_dff_B_GoF85LcZ0_2),.clk(gclk));
	jdff dff_B_ArDhKMWe6_2(.din(w_dff_B_GoF85LcZ0_2),.dout(w_dff_B_ArDhKMWe6_2),.clk(gclk));
	jdff dff_B_FZWaVXJO4_2(.din(w_dff_B_ArDhKMWe6_2),.dout(w_dff_B_FZWaVXJO4_2),.clk(gclk));
	jdff dff_B_ldOADhiu5_2(.din(w_dff_B_FZWaVXJO4_2),.dout(w_dff_B_ldOADhiu5_2),.clk(gclk));
	jdff dff_B_oaREJ4IR5_2(.din(w_dff_B_ldOADhiu5_2),.dout(w_dff_B_oaREJ4IR5_2),.clk(gclk));
	jdff dff_B_8z27Dhzj8_2(.din(w_dff_B_oaREJ4IR5_2),.dout(w_dff_B_8z27Dhzj8_2),.clk(gclk));
	jdff dff_B_N2xtKETd9_2(.din(w_dff_B_8z27Dhzj8_2),.dout(w_dff_B_N2xtKETd9_2),.clk(gclk));
	jdff dff_B_hbCXoDJi4_2(.din(w_dff_B_N2xtKETd9_2),.dout(w_dff_B_hbCXoDJi4_2),.clk(gclk));
	jdff dff_B_tw11y9qt5_2(.din(w_dff_B_hbCXoDJi4_2),.dout(w_dff_B_tw11y9qt5_2),.clk(gclk));
	jdff dff_B_F5wxppnt0_2(.din(w_dff_B_tw11y9qt5_2),.dout(w_dff_B_F5wxppnt0_2),.clk(gclk));
	jdff dff_B_m94nor1V1_2(.din(w_dff_B_F5wxppnt0_2),.dout(w_dff_B_m94nor1V1_2),.clk(gclk));
	jdff dff_B_W4ymwp633_2(.din(w_dff_B_m94nor1V1_2),.dout(w_dff_B_W4ymwp633_2),.clk(gclk));
	jdff dff_B_axL7CF5E3_2(.din(w_dff_B_W4ymwp633_2),.dout(w_dff_B_axL7CF5E3_2),.clk(gclk));
	jdff dff_B_ji4cfoxE8_2(.din(w_dff_B_axL7CF5E3_2),.dout(w_dff_B_ji4cfoxE8_2),.clk(gclk));
	jdff dff_B_XU9zNzmb9_2(.din(w_dff_B_ji4cfoxE8_2),.dout(w_dff_B_XU9zNzmb9_2),.clk(gclk));
	jdff dff_B_7AmvrWmr2_2(.din(n1440),.dout(w_dff_B_7AmvrWmr2_2),.clk(gclk));
	jdff dff_B_fhgkpsz11_1(.din(n1416),.dout(w_dff_B_fhgkpsz11_1),.clk(gclk));
	jdff dff_B_J0m5tXEJ0_2(.din(n1337),.dout(w_dff_B_J0m5tXEJ0_2),.clk(gclk));
	jdff dff_B_M7zkUsJD9_2(.din(w_dff_B_J0m5tXEJ0_2),.dout(w_dff_B_M7zkUsJD9_2),.clk(gclk));
	jdff dff_B_0PW2za2H2_2(.din(w_dff_B_M7zkUsJD9_2),.dout(w_dff_B_0PW2za2H2_2),.clk(gclk));
	jdff dff_B_sBefOyIN1_2(.din(w_dff_B_0PW2za2H2_2),.dout(w_dff_B_sBefOyIN1_2),.clk(gclk));
	jdff dff_B_WOqdT7zu6_2(.din(w_dff_B_sBefOyIN1_2),.dout(w_dff_B_WOqdT7zu6_2),.clk(gclk));
	jdff dff_B_FYe3N1UV9_2(.din(w_dff_B_WOqdT7zu6_2),.dout(w_dff_B_FYe3N1UV9_2),.clk(gclk));
	jdff dff_B_u7h2gh5a1_2(.din(w_dff_B_FYe3N1UV9_2),.dout(w_dff_B_u7h2gh5a1_2),.clk(gclk));
	jdff dff_B_rL7bf5Xe0_2(.din(w_dff_B_u7h2gh5a1_2),.dout(w_dff_B_rL7bf5Xe0_2),.clk(gclk));
	jdff dff_B_6e4h2Ofw5_2(.din(w_dff_B_rL7bf5Xe0_2),.dout(w_dff_B_6e4h2Ofw5_2),.clk(gclk));
	jdff dff_B_yyxgltEE0_2(.din(w_dff_B_6e4h2Ofw5_2),.dout(w_dff_B_yyxgltEE0_2),.clk(gclk));
	jdff dff_B_7iH8rB9v4_2(.din(w_dff_B_yyxgltEE0_2),.dout(w_dff_B_7iH8rB9v4_2),.clk(gclk));
	jdff dff_B_KzE6huZh7_2(.din(w_dff_B_7iH8rB9v4_2),.dout(w_dff_B_KzE6huZh7_2),.clk(gclk));
	jdff dff_B_mQY3A42h5_2(.din(w_dff_B_KzE6huZh7_2),.dout(w_dff_B_mQY3A42h5_2),.clk(gclk));
	jdff dff_B_kn0q0M0M4_2(.din(w_dff_B_mQY3A42h5_2),.dout(w_dff_B_kn0q0M0M4_2),.clk(gclk));
	jdff dff_B_qzmXuNxB3_2(.din(w_dff_B_kn0q0M0M4_2),.dout(w_dff_B_qzmXuNxB3_2),.clk(gclk));
	jdff dff_B_LGULOmy35_2(.din(w_dff_B_qzmXuNxB3_2),.dout(w_dff_B_LGULOmy35_2),.clk(gclk));
	jdff dff_B_WYg5GW4C8_2(.din(w_dff_B_LGULOmy35_2),.dout(w_dff_B_WYg5GW4C8_2),.clk(gclk));
	jdff dff_B_9OEULCYx5_2(.din(w_dff_B_WYg5GW4C8_2),.dout(w_dff_B_9OEULCYx5_2),.clk(gclk));
	jdff dff_B_qbHmGXhI1_2(.din(w_dff_B_9OEULCYx5_2),.dout(w_dff_B_qbHmGXhI1_2),.clk(gclk));
	jdff dff_B_wOTDmG5X4_2(.din(w_dff_B_qbHmGXhI1_2),.dout(w_dff_B_wOTDmG5X4_2),.clk(gclk));
	jdff dff_B_IcJzz89m2_2(.din(w_dff_B_wOTDmG5X4_2),.dout(w_dff_B_IcJzz89m2_2),.clk(gclk));
	jdff dff_B_9SsYb6J03_2(.din(w_dff_B_IcJzz89m2_2),.dout(w_dff_B_9SsYb6J03_2),.clk(gclk));
	jdff dff_B_VNRioU9r3_2(.din(w_dff_B_9SsYb6J03_2),.dout(w_dff_B_VNRioU9r3_2),.clk(gclk));
	jdff dff_B_ApGWT2H27_2(.din(w_dff_B_VNRioU9r3_2),.dout(w_dff_B_ApGWT2H27_2),.clk(gclk));
	jdff dff_B_PemKooQa6_2(.din(w_dff_B_ApGWT2H27_2),.dout(w_dff_B_PemKooQa6_2),.clk(gclk));
	jdff dff_B_LDWxq2Tz1_2(.din(w_dff_B_PemKooQa6_2),.dout(w_dff_B_LDWxq2Tz1_2),.clk(gclk));
	jdff dff_B_oXKCQvLj0_2(.din(n1362),.dout(w_dff_B_oXKCQvLj0_2),.clk(gclk));
	jdff dff_B_RCvdprrW0_1(.din(n1338),.dout(w_dff_B_RCvdprrW0_1),.clk(gclk));
	jdff dff_B_K6oej78G5_2(.din(n1252),.dout(w_dff_B_K6oej78G5_2),.clk(gclk));
	jdff dff_B_mbWKxVcy1_2(.din(w_dff_B_K6oej78G5_2),.dout(w_dff_B_mbWKxVcy1_2),.clk(gclk));
	jdff dff_B_UO3mjFJ69_2(.din(w_dff_B_mbWKxVcy1_2),.dout(w_dff_B_UO3mjFJ69_2),.clk(gclk));
	jdff dff_B_WtkGxZ4T0_2(.din(w_dff_B_UO3mjFJ69_2),.dout(w_dff_B_WtkGxZ4T0_2),.clk(gclk));
	jdff dff_B_yQXfnlFn1_2(.din(w_dff_B_WtkGxZ4T0_2),.dout(w_dff_B_yQXfnlFn1_2),.clk(gclk));
	jdff dff_B_AylUQdnU8_2(.din(w_dff_B_yQXfnlFn1_2),.dout(w_dff_B_AylUQdnU8_2),.clk(gclk));
	jdff dff_B_RhSjcLl70_2(.din(w_dff_B_AylUQdnU8_2),.dout(w_dff_B_RhSjcLl70_2),.clk(gclk));
	jdff dff_B_UxqJJMzN7_2(.din(w_dff_B_RhSjcLl70_2),.dout(w_dff_B_UxqJJMzN7_2),.clk(gclk));
	jdff dff_B_vwIjTXup1_2(.din(w_dff_B_UxqJJMzN7_2),.dout(w_dff_B_vwIjTXup1_2),.clk(gclk));
	jdff dff_B_7Pjut8BE2_2(.din(w_dff_B_vwIjTXup1_2),.dout(w_dff_B_7Pjut8BE2_2),.clk(gclk));
	jdff dff_B_0tfE0Zod5_2(.din(w_dff_B_7Pjut8BE2_2),.dout(w_dff_B_0tfE0Zod5_2),.clk(gclk));
	jdff dff_B_gzXi3Ktd1_2(.din(w_dff_B_0tfE0Zod5_2),.dout(w_dff_B_gzXi3Ktd1_2),.clk(gclk));
	jdff dff_B_oVi7Px857_2(.din(w_dff_B_gzXi3Ktd1_2),.dout(w_dff_B_oVi7Px857_2),.clk(gclk));
	jdff dff_B_IwYVabqU5_2(.din(w_dff_B_oVi7Px857_2),.dout(w_dff_B_IwYVabqU5_2),.clk(gclk));
	jdff dff_B_t2pHHfU22_2(.din(w_dff_B_IwYVabqU5_2),.dout(w_dff_B_t2pHHfU22_2),.clk(gclk));
	jdff dff_B_AkPOQ7AW2_2(.din(w_dff_B_t2pHHfU22_2),.dout(w_dff_B_AkPOQ7AW2_2),.clk(gclk));
	jdff dff_B_ZTAd8W0A4_2(.din(w_dff_B_AkPOQ7AW2_2),.dout(w_dff_B_ZTAd8W0A4_2),.clk(gclk));
	jdff dff_B_JX6xhG9F6_2(.din(w_dff_B_ZTAd8W0A4_2),.dout(w_dff_B_JX6xhG9F6_2),.clk(gclk));
	jdff dff_B_hhOQQPkJ8_2(.din(w_dff_B_JX6xhG9F6_2),.dout(w_dff_B_hhOQQPkJ8_2),.clk(gclk));
	jdff dff_B_6uh1CL0c9_2(.din(w_dff_B_hhOQQPkJ8_2),.dout(w_dff_B_6uh1CL0c9_2),.clk(gclk));
	jdff dff_B_07sf7OJa5_2(.din(w_dff_B_6uh1CL0c9_2),.dout(w_dff_B_07sf7OJa5_2),.clk(gclk));
	jdff dff_B_Mg0dzEFw8_2(.din(w_dff_B_07sf7OJa5_2),.dout(w_dff_B_Mg0dzEFw8_2),.clk(gclk));
	jdff dff_B_rWoV4dyW9_2(.din(w_dff_B_Mg0dzEFw8_2),.dout(w_dff_B_rWoV4dyW9_2),.clk(gclk));
	jdff dff_B_XFi4CKxd4_2(.din(n1277),.dout(w_dff_B_XFi4CKxd4_2),.clk(gclk));
	jdff dff_B_XA6EwYAF0_1(.din(n1253),.dout(w_dff_B_XA6EwYAF0_1),.clk(gclk));
	jdff dff_B_ZgFSeLE93_2(.din(n1161),.dout(w_dff_B_ZgFSeLE93_2),.clk(gclk));
	jdff dff_B_4kXPqXZx7_2(.din(w_dff_B_ZgFSeLE93_2),.dout(w_dff_B_4kXPqXZx7_2),.clk(gclk));
	jdff dff_B_preJuuKJ6_2(.din(w_dff_B_4kXPqXZx7_2),.dout(w_dff_B_preJuuKJ6_2),.clk(gclk));
	jdff dff_B_6JMv849W1_2(.din(w_dff_B_preJuuKJ6_2),.dout(w_dff_B_6JMv849W1_2),.clk(gclk));
	jdff dff_B_nGeIk8gy3_2(.din(w_dff_B_6JMv849W1_2),.dout(w_dff_B_nGeIk8gy3_2),.clk(gclk));
	jdff dff_B_fsE8v4dZ8_2(.din(w_dff_B_nGeIk8gy3_2),.dout(w_dff_B_fsE8v4dZ8_2),.clk(gclk));
	jdff dff_B_z9VJK7IZ7_2(.din(w_dff_B_fsE8v4dZ8_2),.dout(w_dff_B_z9VJK7IZ7_2),.clk(gclk));
	jdff dff_B_kQ3OXmrY2_2(.din(w_dff_B_z9VJK7IZ7_2),.dout(w_dff_B_kQ3OXmrY2_2),.clk(gclk));
	jdff dff_B_d14JP68W0_2(.din(w_dff_B_kQ3OXmrY2_2),.dout(w_dff_B_d14JP68W0_2),.clk(gclk));
	jdff dff_B_sEJTVhfV8_2(.din(w_dff_B_d14JP68W0_2),.dout(w_dff_B_sEJTVhfV8_2),.clk(gclk));
	jdff dff_B_q7VaESVD2_2(.din(w_dff_B_sEJTVhfV8_2),.dout(w_dff_B_q7VaESVD2_2),.clk(gclk));
	jdff dff_B_z3LdGgzA6_2(.din(w_dff_B_q7VaESVD2_2),.dout(w_dff_B_z3LdGgzA6_2),.clk(gclk));
	jdff dff_B_s6Uw1iiy0_2(.din(w_dff_B_z3LdGgzA6_2),.dout(w_dff_B_s6Uw1iiy0_2),.clk(gclk));
	jdff dff_B_AWaUS11O1_2(.din(w_dff_B_s6Uw1iiy0_2),.dout(w_dff_B_AWaUS11O1_2),.clk(gclk));
	jdff dff_B_UHC1K1kB7_2(.din(w_dff_B_AWaUS11O1_2),.dout(w_dff_B_UHC1K1kB7_2),.clk(gclk));
	jdff dff_B_C3mduFv11_2(.din(w_dff_B_UHC1K1kB7_2),.dout(w_dff_B_C3mduFv11_2),.clk(gclk));
	jdff dff_B_NKA4irhU5_2(.din(w_dff_B_C3mduFv11_2),.dout(w_dff_B_NKA4irhU5_2),.clk(gclk));
	jdff dff_B_aLmtdjwg7_2(.din(w_dff_B_NKA4irhU5_2),.dout(w_dff_B_aLmtdjwg7_2),.clk(gclk));
	jdff dff_B_nV1wXi2P0_2(.din(w_dff_B_aLmtdjwg7_2),.dout(w_dff_B_nV1wXi2P0_2),.clk(gclk));
	jdff dff_B_2uCsVlcn6_2(.din(w_dff_B_nV1wXi2P0_2),.dout(w_dff_B_2uCsVlcn6_2),.clk(gclk));
	jdff dff_B_p4KQoNjV9_2(.din(n1186),.dout(w_dff_B_p4KQoNjV9_2),.clk(gclk));
	jdff dff_B_Klmu89BJ8_1(.din(n1162),.dout(w_dff_B_Klmu89BJ8_1),.clk(gclk));
	jdff dff_B_VhtQ0F8U1_2(.din(n1063),.dout(w_dff_B_VhtQ0F8U1_2),.clk(gclk));
	jdff dff_B_S41vNDXG9_2(.din(w_dff_B_VhtQ0F8U1_2),.dout(w_dff_B_S41vNDXG9_2),.clk(gclk));
	jdff dff_B_5FkHNdIs9_2(.din(w_dff_B_S41vNDXG9_2),.dout(w_dff_B_5FkHNdIs9_2),.clk(gclk));
	jdff dff_B_DHaLOYlK7_2(.din(w_dff_B_5FkHNdIs9_2),.dout(w_dff_B_DHaLOYlK7_2),.clk(gclk));
	jdff dff_B_D0p5I5LU2_2(.din(w_dff_B_DHaLOYlK7_2),.dout(w_dff_B_D0p5I5LU2_2),.clk(gclk));
	jdff dff_B_s1sw8CgJ1_2(.din(w_dff_B_D0p5I5LU2_2),.dout(w_dff_B_s1sw8CgJ1_2),.clk(gclk));
	jdff dff_B_Imy5NynV1_2(.din(w_dff_B_s1sw8CgJ1_2),.dout(w_dff_B_Imy5NynV1_2),.clk(gclk));
	jdff dff_B_nrLixpA81_2(.din(w_dff_B_Imy5NynV1_2),.dout(w_dff_B_nrLixpA81_2),.clk(gclk));
	jdff dff_B_4yLsAD8X9_2(.din(w_dff_B_nrLixpA81_2),.dout(w_dff_B_4yLsAD8X9_2),.clk(gclk));
	jdff dff_B_ilrJxCb46_2(.din(w_dff_B_4yLsAD8X9_2),.dout(w_dff_B_ilrJxCb46_2),.clk(gclk));
	jdff dff_B_ws29kss34_2(.din(w_dff_B_ilrJxCb46_2),.dout(w_dff_B_ws29kss34_2),.clk(gclk));
	jdff dff_B_3RbpLpql2_2(.din(w_dff_B_ws29kss34_2),.dout(w_dff_B_3RbpLpql2_2),.clk(gclk));
	jdff dff_B_bO280q4X1_2(.din(w_dff_B_3RbpLpql2_2),.dout(w_dff_B_bO280q4X1_2),.clk(gclk));
	jdff dff_B_O3ciAwDl7_2(.din(w_dff_B_bO280q4X1_2),.dout(w_dff_B_O3ciAwDl7_2),.clk(gclk));
	jdff dff_B_XgTjRMOj1_2(.din(w_dff_B_O3ciAwDl7_2),.dout(w_dff_B_XgTjRMOj1_2),.clk(gclk));
	jdff dff_B_z8K4H9mD3_2(.din(w_dff_B_XgTjRMOj1_2),.dout(w_dff_B_z8K4H9mD3_2),.clk(gclk));
	jdff dff_B_UBQUdD8G3_2(.din(w_dff_B_z8K4H9mD3_2),.dout(w_dff_B_UBQUdD8G3_2),.clk(gclk));
	jdff dff_B_9dj6N0cZ0_2(.din(n1087),.dout(w_dff_B_9dj6N0cZ0_2),.clk(gclk));
	jdff dff_B_lElzpUqB8_1(.din(n1064),.dout(w_dff_B_lElzpUqB8_1),.clk(gclk));
	jdff dff_B_I99xRRJk7_2(.din(n964),.dout(w_dff_B_I99xRRJk7_2),.clk(gclk));
	jdff dff_B_bRlAjyl20_2(.din(w_dff_B_I99xRRJk7_2),.dout(w_dff_B_bRlAjyl20_2),.clk(gclk));
	jdff dff_B_ihixATLA1_2(.din(w_dff_B_bRlAjyl20_2),.dout(w_dff_B_ihixATLA1_2),.clk(gclk));
	jdff dff_B_hC0M6Dok5_2(.din(w_dff_B_ihixATLA1_2),.dout(w_dff_B_hC0M6Dok5_2),.clk(gclk));
	jdff dff_B_hq3ZFMDV9_2(.din(w_dff_B_hC0M6Dok5_2),.dout(w_dff_B_hq3ZFMDV9_2),.clk(gclk));
	jdff dff_B_HD64EQci4_2(.din(w_dff_B_hq3ZFMDV9_2),.dout(w_dff_B_HD64EQci4_2),.clk(gclk));
	jdff dff_B_xMu8lGfQ9_2(.din(w_dff_B_HD64EQci4_2),.dout(w_dff_B_xMu8lGfQ9_2),.clk(gclk));
	jdff dff_B_aXNFyKXY9_2(.din(w_dff_B_xMu8lGfQ9_2),.dout(w_dff_B_aXNFyKXY9_2),.clk(gclk));
	jdff dff_B_dXW1jjuC2_2(.din(w_dff_B_aXNFyKXY9_2),.dout(w_dff_B_dXW1jjuC2_2),.clk(gclk));
	jdff dff_B_9TMbwzxA3_2(.din(w_dff_B_dXW1jjuC2_2),.dout(w_dff_B_9TMbwzxA3_2),.clk(gclk));
	jdff dff_B_YY3jv06z6_2(.din(w_dff_B_9TMbwzxA3_2),.dout(w_dff_B_YY3jv06z6_2),.clk(gclk));
	jdff dff_B_j0QtQlh04_2(.din(w_dff_B_YY3jv06z6_2),.dout(w_dff_B_j0QtQlh04_2),.clk(gclk));
	jdff dff_B_92GYoN5c6_2(.din(w_dff_B_j0QtQlh04_2),.dout(w_dff_B_92GYoN5c6_2),.clk(gclk));
	jdff dff_B_GpUGpCoU0_2(.din(w_dff_B_92GYoN5c6_2),.dout(w_dff_B_GpUGpCoU0_2),.clk(gclk));
	jdff dff_B_FFyMfjKa9_2(.din(n988),.dout(w_dff_B_FFyMfjKa9_2),.clk(gclk));
	jdff dff_B_AEG78ezj7_1(.din(n965),.dout(w_dff_B_AEG78ezj7_1),.clk(gclk));
	jdff dff_B_3pGNk0yz0_2(.din(n862),.dout(w_dff_B_3pGNk0yz0_2),.clk(gclk));
	jdff dff_B_FooUfOxn0_2(.din(w_dff_B_3pGNk0yz0_2),.dout(w_dff_B_FooUfOxn0_2),.clk(gclk));
	jdff dff_B_pMR0IVFP0_2(.din(w_dff_B_FooUfOxn0_2),.dout(w_dff_B_pMR0IVFP0_2),.clk(gclk));
	jdff dff_B_rRswQRFe0_2(.din(w_dff_B_pMR0IVFP0_2),.dout(w_dff_B_rRswQRFe0_2),.clk(gclk));
	jdff dff_B_dzeX0QTt6_2(.din(w_dff_B_rRswQRFe0_2),.dout(w_dff_B_dzeX0QTt6_2),.clk(gclk));
	jdff dff_B_YfGZtyco7_2(.din(w_dff_B_dzeX0QTt6_2),.dout(w_dff_B_YfGZtyco7_2),.clk(gclk));
	jdff dff_B_yC0Dj2CN2_2(.din(w_dff_B_YfGZtyco7_2),.dout(w_dff_B_yC0Dj2CN2_2),.clk(gclk));
	jdff dff_B_YecMjM0H4_2(.din(w_dff_B_yC0Dj2CN2_2),.dout(w_dff_B_YecMjM0H4_2),.clk(gclk));
	jdff dff_B_SsgKgUyf4_2(.din(w_dff_B_YecMjM0H4_2),.dout(w_dff_B_SsgKgUyf4_2),.clk(gclk));
	jdff dff_B_bIphNa268_2(.din(w_dff_B_SsgKgUyf4_2),.dout(w_dff_B_bIphNa268_2),.clk(gclk));
	jdff dff_B_wSkPVZ5H8_2(.din(w_dff_B_bIphNa268_2),.dout(w_dff_B_wSkPVZ5H8_2),.clk(gclk));
	jdff dff_B_R921Ezfz5_2(.din(n882),.dout(w_dff_B_R921Ezfz5_2),.clk(gclk));
	jdff dff_B_mHlV8etn5_1(.din(n863),.dout(w_dff_B_mHlV8etn5_1),.clk(gclk));
	jdff dff_B_ybLsXfET3_2(.din(n764),.dout(w_dff_B_ybLsXfET3_2),.clk(gclk));
	jdff dff_B_i7KImOju7_2(.din(w_dff_B_ybLsXfET3_2),.dout(w_dff_B_i7KImOju7_2),.clk(gclk));
	jdff dff_B_P8FnVOW29_2(.din(w_dff_B_i7KImOju7_2),.dout(w_dff_B_P8FnVOW29_2),.clk(gclk));
	jdff dff_B_cYHompDw4_2(.din(w_dff_B_P8FnVOW29_2),.dout(w_dff_B_cYHompDw4_2),.clk(gclk));
	jdff dff_B_a0jShjwR1_2(.din(w_dff_B_cYHompDw4_2),.dout(w_dff_B_a0jShjwR1_2),.clk(gclk));
	jdff dff_B_cSQmYooW7_2(.din(w_dff_B_a0jShjwR1_2),.dout(w_dff_B_cSQmYooW7_2),.clk(gclk));
	jdff dff_B_JQI5isGO9_2(.din(w_dff_B_cSQmYooW7_2),.dout(w_dff_B_JQI5isGO9_2),.clk(gclk));
	jdff dff_B_EXRxjeOL2_2(.din(w_dff_B_JQI5isGO9_2),.dout(w_dff_B_EXRxjeOL2_2),.clk(gclk));
	jdff dff_B_pEsvVSsL5_2(.din(n779),.dout(w_dff_B_pEsvVSsL5_2),.clk(gclk));
	jdff dff_B_28L4XTPF9_2(.din(w_dff_B_pEsvVSsL5_2),.dout(w_dff_B_28L4XTPF9_2),.clk(gclk));
	jdff dff_B_px5urLfF6_2(.din(w_dff_B_28L4XTPF9_2),.dout(w_dff_B_px5urLfF6_2),.clk(gclk));
	jdff dff_B_ndMJxwyC9_1(.din(n765),.dout(w_dff_B_ndMJxwyC9_1),.clk(gclk));
	jdff dff_B_ny94K4xr4_1(.din(w_dff_B_ndMJxwyC9_1),.dout(w_dff_B_ny94K4xr4_1),.clk(gclk));
	jdff dff_B_6OKlmBQJ6_2(.din(n674),.dout(w_dff_B_6OKlmBQJ6_2),.clk(gclk));
	jdff dff_B_QDOksBRU7_2(.din(w_dff_B_6OKlmBQJ6_2),.dout(w_dff_B_QDOksBRU7_2),.clk(gclk));
	jdff dff_B_ymoeGeBM1_2(.din(w_dff_B_QDOksBRU7_2),.dout(w_dff_B_ymoeGeBM1_2),.clk(gclk));
	jdff dff_B_2G8Dmrc76_0(.din(n679),.dout(w_dff_B_2G8Dmrc76_0),.clk(gclk));
	jdff dff_A_5u9AfVKa4_0(.dout(w_n586_0[0]),.din(w_dff_A_5u9AfVKa4_0),.clk(gclk));
	jdff dff_A_lI9Tl6Ax2_0(.dout(w_dff_A_5u9AfVKa4_0),.din(w_dff_A_lI9Tl6Ax2_0),.clk(gclk));
	jdff dff_A_toJ3qaRi7_1(.dout(w_n586_0[1]),.din(w_dff_A_toJ3qaRi7_1),.clk(gclk));
	jdff dff_A_SA268giF4_1(.dout(w_dff_A_toJ3qaRi7_1),.din(w_dff_A_SA268giF4_1),.clk(gclk));
	jdff dff_B_gTft9evD3_1(.din(n1788),.dout(w_dff_B_gTft9evD3_1),.clk(gclk));
	jdff dff_A_qYRAclYB1_1(.dout(w_n1770_0[1]),.din(w_dff_A_qYRAclYB1_1),.clk(gclk));
	jdff dff_B_OVSklzkW6_1(.din(n1768),.dout(w_dff_B_OVSklzkW6_1),.clk(gclk));
	jdff dff_B_CBTpJeBU1_2(.din(n1739),.dout(w_dff_B_CBTpJeBU1_2),.clk(gclk));
	jdff dff_B_cWF9zexF1_2(.din(w_dff_B_CBTpJeBU1_2),.dout(w_dff_B_cWF9zexF1_2),.clk(gclk));
	jdff dff_B_LhDtNopF9_2(.din(w_dff_B_cWF9zexF1_2),.dout(w_dff_B_LhDtNopF9_2),.clk(gclk));
	jdff dff_B_e1VZUiPv8_2(.din(w_dff_B_LhDtNopF9_2),.dout(w_dff_B_e1VZUiPv8_2),.clk(gclk));
	jdff dff_B_wE7C7L9t3_2(.din(w_dff_B_e1VZUiPv8_2),.dout(w_dff_B_wE7C7L9t3_2),.clk(gclk));
	jdff dff_B_CJ7gv1az3_2(.din(w_dff_B_wE7C7L9t3_2),.dout(w_dff_B_CJ7gv1az3_2),.clk(gclk));
	jdff dff_B_CybqY79d8_2(.din(w_dff_B_CJ7gv1az3_2),.dout(w_dff_B_CybqY79d8_2),.clk(gclk));
	jdff dff_B_NMnYLpWk7_2(.din(w_dff_B_CybqY79d8_2),.dout(w_dff_B_NMnYLpWk7_2),.clk(gclk));
	jdff dff_B_x8EaEdZO8_2(.din(w_dff_B_NMnYLpWk7_2),.dout(w_dff_B_x8EaEdZO8_2),.clk(gclk));
	jdff dff_B_VVrmtqHx5_2(.din(w_dff_B_x8EaEdZO8_2),.dout(w_dff_B_VVrmtqHx5_2),.clk(gclk));
	jdff dff_B_flKJsC0X0_2(.din(w_dff_B_VVrmtqHx5_2),.dout(w_dff_B_flKJsC0X0_2),.clk(gclk));
	jdff dff_B_zJwt8dYs8_2(.din(w_dff_B_flKJsC0X0_2),.dout(w_dff_B_zJwt8dYs8_2),.clk(gclk));
	jdff dff_B_czGG51lP5_2(.din(w_dff_B_zJwt8dYs8_2),.dout(w_dff_B_czGG51lP5_2),.clk(gclk));
	jdff dff_B_fT49r7xT1_2(.din(w_dff_B_czGG51lP5_2),.dout(w_dff_B_fT49r7xT1_2),.clk(gclk));
	jdff dff_B_xxup8haT6_2(.din(w_dff_B_fT49r7xT1_2),.dout(w_dff_B_xxup8haT6_2),.clk(gclk));
	jdff dff_B_ABDIfSrK3_2(.din(w_dff_B_xxup8haT6_2),.dout(w_dff_B_ABDIfSrK3_2),.clk(gclk));
	jdff dff_B_THITAzdv3_2(.din(w_dff_B_ABDIfSrK3_2),.dout(w_dff_B_THITAzdv3_2),.clk(gclk));
	jdff dff_B_6StuxNoU3_2(.din(w_dff_B_THITAzdv3_2),.dout(w_dff_B_6StuxNoU3_2),.clk(gclk));
	jdff dff_B_hSJDsKhL3_2(.din(w_dff_B_6StuxNoU3_2),.dout(w_dff_B_hSJDsKhL3_2),.clk(gclk));
	jdff dff_B_MqvlbyyA9_2(.din(w_dff_B_hSJDsKhL3_2),.dout(w_dff_B_MqvlbyyA9_2),.clk(gclk));
	jdff dff_B_5GRkqyut1_2(.din(w_dff_B_MqvlbyyA9_2),.dout(w_dff_B_5GRkqyut1_2),.clk(gclk));
	jdff dff_B_z2AAoVie6_2(.din(w_dff_B_5GRkqyut1_2),.dout(w_dff_B_z2AAoVie6_2),.clk(gclk));
	jdff dff_B_xFmRr5hD8_2(.din(w_dff_B_z2AAoVie6_2),.dout(w_dff_B_xFmRr5hD8_2),.clk(gclk));
	jdff dff_B_1EI6BfdN1_2(.din(w_dff_B_xFmRr5hD8_2),.dout(w_dff_B_1EI6BfdN1_2),.clk(gclk));
	jdff dff_B_rwsV5ITJ7_2(.din(w_dff_B_1EI6BfdN1_2),.dout(w_dff_B_rwsV5ITJ7_2),.clk(gclk));
	jdff dff_B_i6TtNGgf4_2(.din(w_dff_B_rwsV5ITJ7_2),.dout(w_dff_B_i6TtNGgf4_2),.clk(gclk));
	jdff dff_B_LVa7GPqN8_2(.din(w_dff_B_i6TtNGgf4_2),.dout(w_dff_B_LVa7GPqN8_2),.clk(gclk));
	jdff dff_B_S92yJVOM2_2(.din(w_dff_B_LVa7GPqN8_2),.dout(w_dff_B_S92yJVOM2_2),.clk(gclk));
	jdff dff_B_BbrlAjXw0_2(.din(w_dff_B_S92yJVOM2_2),.dout(w_dff_B_BbrlAjXw0_2),.clk(gclk));
	jdff dff_B_XmjbQ9ms5_2(.din(w_dff_B_BbrlAjXw0_2),.dout(w_dff_B_XmjbQ9ms5_2),.clk(gclk));
	jdff dff_B_04cfFUiZ1_2(.din(w_dff_B_XmjbQ9ms5_2),.dout(w_dff_B_04cfFUiZ1_2),.clk(gclk));
	jdff dff_B_dvjIDWEU1_2(.din(w_dff_B_04cfFUiZ1_2),.dout(w_dff_B_dvjIDWEU1_2),.clk(gclk));
	jdff dff_B_K3vfERUE5_2(.din(w_dff_B_dvjIDWEU1_2),.dout(w_dff_B_K3vfERUE5_2),.clk(gclk));
	jdff dff_B_9P0P5iPE6_2(.din(w_dff_B_K3vfERUE5_2),.dout(w_dff_B_9P0P5iPE6_2),.clk(gclk));
	jdff dff_B_g0v9ARu22_2(.din(w_dff_B_9P0P5iPE6_2),.dout(w_dff_B_g0v9ARu22_2),.clk(gclk));
	jdff dff_B_79ohoplp4_2(.din(w_dff_B_g0v9ARu22_2),.dout(w_dff_B_79ohoplp4_2),.clk(gclk));
	jdff dff_B_7kBKBRLV9_2(.din(w_dff_B_79ohoplp4_2),.dout(w_dff_B_7kBKBRLV9_2),.clk(gclk));
	jdff dff_B_3FU7fnm00_2(.din(w_dff_B_7kBKBRLV9_2),.dout(w_dff_B_3FU7fnm00_2),.clk(gclk));
	jdff dff_B_JKUv5p9S3_2(.din(w_dff_B_3FU7fnm00_2),.dout(w_dff_B_JKUv5p9S3_2),.clk(gclk));
	jdff dff_B_mNSbcnuv1_2(.din(w_dff_B_JKUv5p9S3_2),.dout(w_dff_B_mNSbcnuv1_2),.clk(gclk));
	jdff dff_B_PA4h3NaM5_2(.din(w_dff_B_mNSbcnuv1_2),.dout(w_dff_B_PA4h3NaM5_2),.clk(gclk));
	jdff dff_B_689Pt4u27_2(.din(w_dff_B_PA4h3NaM5_2),.dout(w_dff_B_689Pt4u27_2),.clk(gclk));
	jdff dff_B_aXoTpu649_2(.din(w_dff_B_689Pt4u27_2),.dout(w_dff_B_aXoTpu649_2),.clk(gclk));
	jdff dff_B_Pmw4J4Ih7_2(.din(w_dff_B_aXoTpu649_2),.dout(w_dff_B_Pmw4J4Ih7_2),.clk(gclk));
	jdff dff_B_krbNcL2i3_2(.din(w_dff_B_Pmw4J4Ih7_2),.dout(w_dff_B_krbNcL2i3_2),.clk(gclk));
	jdff dff_B_8Dxmp4ON5_2(.din(w_dff_B_krbNcL2i3_2),.dout(w_dff_B_8Dxmp4ON5_2),.clk(gclk));
	jdff dff_B_B97tuTB35_2(.din(w_dff_B_8Dxmp4ON5_2),.dout(w_dff_B_B97tuTB35_2),.clk(gclk));
	jdff dff_B_p5pi7sEK0_2(.din(w_dff_B_B97tuTB35_2),.dout(w_dff_B_p5pi7sEK0_2),.clk(gclk));
	jdff dff_B_7lIgAyzM7_2(.din(w_dff_B_p5pi7sEK0_2),.dout(w_dff_B_7lIgAyzM7_2),.clk(gclk));
	jdff dff_B_5eC0TGI62_2(.din(w_dff_B_7lIgAyzM7_2),.dout(w_dff_B_5eC0TGI62_2),.clk(gclk));
	jdff dff_B_M75QlrxF7_2(.din(n1742),.dout(w_dff_B_M75QlrxF7_2),.clk(gclk));
	jdff dff_B_IJm0KGB21_1(.din(n1740),.dout(w_dff_B_IJm0KGB21_1),.clk(gclk));
	jdff dff_B_ewmSuU8E4_2(.din(n1704),.dout(w_dff_B_ewmSuU8E4_2),.clk(gclk));
	jdff dff_B_se2OTqVx4_2(.din(w_dff_B_ewmSuU8E4_2),.dout(w_dff_B_se2OTqVx4_2),.clk(gclk));
	jdff dff_B_xpCqhpgU5_2(.din(w_dff_B_se2OTqVx4_2),.dout(w_dff_B_xpCqhpgU5_2),.clk(gclk));
	jdff dff_B_IOrp231l9_2(.din(w_dff_B_xpCqhpgU5_2),.dout(w_dff_B_IOrp231l9_2),.clk(gclk));
	jdff dff_B_z3XbKRlS4_2(.din(w_dff_B_IOrp231l9_2),.dout(w_dff_B_z3XbKRlS4_2),.clk(gclk));
	jdff dff_B_DfeeHPYi6_2(.din(w_dff_B_z3XbKRlS4_2),.dout(w_dff_B_DfeeHPYi6_2),.clk(gclk));
	jdff dff_B_tUQStImV2_2(.din(w_dff_B_DfeeHPYi6_2),.dout(w_dff_B_tUQStImV2_2),.clk(gclk));
	jdff dff_B_MuUMjhc89_2(.din(w_dff_B_tUQStImV2_2),.dout(w_dff_B_MuUMjhc89_2),.clk(gclk));
	jdff dff_B_kFPuXkXY5_2(.din(w_dff_B_MuUMjhc89_2),.dout(w_dff_B_kFPuXkXY5_2),.clk(gclk));
	jdff dff_B_KIpOZCrK4_2(.din(w_dff_B_kFPuXkXY5_2),.dout(w_dff_B_KIpOZCrK4_2),.clk(gclk));
	jdff dff_B_psENIpg98_2(.din(w_dff_B_KIpOZCrK4_2),.dout(w_dff_B_psENIpg98_2),.clk(gclk));
	jdff dff_B_yzVsX0nW7_2(.din(w_dff_B_psENIpg98_2),.dout(w_dff_B_yzVsX0nW7_2),.clk(gclk));
	jdff dff_B_Z50GMZMd8_2(.din(w_dff_B_yzVsX0nW7_2),.dout(w_dff_B_Z50GMZMd8_2),.clk(gclk));
	jdff dff_B_s2X1SFth1_2(.din(w_dff_B_Z50GMZMd8_2),.dout(w_dff_B_s2X1SFth1_2),.clk(gclk));
	jdff dff_B_IPKxiNFC4_2(.din(w_dff_B_s2X1SFth1_2),.dout(w_dff_B_IPKxiNFC4_2),.clk(gclk));
	jdff dff_B_pQXUsDfd1_2(.din(w_dff_B_IPKxiNFC4_2),.dout(w_dff_B_pQXUsDfd1_2),.clk(gclk));
	jdff dff_B_cukDzmpN0_2(.din(w_dff_B_pQXUsDfd1_2),.dout(w_dff_B_cukDzmpN0_2),.clk(gclk));
	jdff dff_B_aX7gAgJ73_2(.din(w_dff_B_cukDzmpN0_2),.dout(w_dff_B_aX7gAgJ73_2),.clk(gclk));
	jdff dff_B_iS20eu445_2(.din(w_dff_B_aX7gAgJ73_2),.dout(w_dff_B_iS20eu445_2),.clk(gclk));
	jdff dff_B_4kMd7Gqp5_2(.din(w_dff_B_iS20eu445_2),.dout(w_dff_B_4kMd7Gqp5_2),.clk(gclk));
	jdff dff_B_V5lSAUpo3_2(.din(w_dff_B_4kMd7Gqp5_2),.dout(w_dff_B_V5lSAUpo3_2),.clk(gclk));
	jdff dff_B_qIBPcK4C0_2(.din(w_dff_B_V5lSAUpo3_2),.dout(w_dff_B_qIBPcK4C0_2),.clk(gclk));
	jdff dff_B_BBE16eG26_2(.din(w_dff_B_qIBPcK4C0_2),.dout(w_dff_B_BBE16eG26_2),.clk(gclk));
	jdff dff_B_y9eYEcky2_2(.din(w_dff_B_BBE16eG26_2),.dout(w_dff_B_y9eYEcky2_2),.clk(gclk));
	jdff dff_B_0roA5NhG1_2(.din(w_dff_B_y9eYEcky2_2),.dout(w_dff_B_0roA5NhG1_2),.clk(gclk));
	jdff dff_B_t4qJS2Tn9_2(.din(w_dff_B_0roA5NhG1_2),.dout(w_dff_B_t4qJS2Tn9_2),.clk(gclk));
	jdff dff_B_t34YdNge6_2(.din(w_dff_B_t4qJS2Tn9_2),.dout(w_dff_B_t34YdNge6_2),.clk(gclk));
	jdff dff_B_XWIUAX9k0_2(.din(w_dff_B_t34YdNge6_2),.dout(w_dff_B_XWIUAX9k0_2),.clk(gclk));
	jdff dff_B_pKQkGmkS1_2(.din(w_dff_B_XWIUAX9k0_2),.dout(w_dff_B_pKQkGmkS1_2),.clk(gclk));
	jdff dff_B_I15EsNas6_2(.din(w_dff_B_pKQkGmkS1_2),.dout(w_dff_B_I15EsNas6_2),.clk(gclk));
	jdff dff_B_GenIUEX24_2(.din(w_dff_B_I15EsNas6_2),.dout(w_dff_B_GenIUEX24_2),.clk(gclk));
	jdff dff_B_rbVrT2E62_2(.din(w_dff_B_GenIUEX24_2),.dout(w_dff_B_rbVrT2E62_2),.clk(gclk));
	jdff dff_B_KqmLfOlG6_2(.din(w_dff_B_rbVrT2E62_2),.dout(w_dff_B_KqmLfOlG6_2),.clk(gclk));
	jdff dff_B_8aEYebXt9_2(.din(w_dff_B_KqmLfOlG6_2),.dout(w_dff_B_8aEYebXt9_2),.clk(gclk));
	jdff dff_B_wc1wAwBc7_2(.din(w_dff_B_8aEYebXt9_2),.dout(w_dff_B_wc1wAwBc7_2),.clk(gclk));
	jdff dff_B_lEmWHFXi5_2(.din(w_dff_B_wc1wAwBc7_2),.dout(w_dff_B_lEmWHFXi5_2),.clk(gclk));
	jdff dff_B_qCGAblvd4_2(.din(w_dff_B_lEmWHFXi5_2),.dout(w_dff_B_qCGAblvd4_2),.clk(gclk));
	jdff dff_B_fmOeRQYn1_2(.din(w_dff_B_qCGAblvd4_2),.dout(w_dff_B_fmOeRQYn1_2),.clk(gclk));
	jdff dff_B_m4o2AZ9N0_2(.din(w_dff_B_fmOeRQYn1_2),.dout(w_dff_B_m4o2AZ9N0_2),.clk(gclk));
	jdff dff_B_fSG9SH0t3_2(.din(w_dff_B_m4o2AZ9N0_2),.dout(w_dff_B_fSG9SH0t3_2),.clk(gclk));
	jdff dff_B_BZGSdULB3_2(.din(w_dff_B_fSG9SH0t3_2),.dout(w_dff_B_BZGSdULB3_2),.clk(gclk));
	jdff dff_B_FSimbVGz8_2(.din(w_dff_B_BZGSdULB3_2),.dout(w_dff_B_FSimbVGz8_2),.clk(gclk));
	jdff dff_B_4TCVkJQQ4_2(.din(w_dff_B_FSimbVGz8_2),.dout(w_dff_B_4TCVkJQQ4_2),.clk(gclk));
	jdff dff_B_dywIAmWK6_2(.din(w_dff_B_4TCVkJQQ4_2),.dout(w_dff_B_dywIAmWK6_2),.clk(gclk));
	jdff dff_B_p4sLLeAm1_2(.din(w_dff_B_dywIAmWK6_2),.dout(w_dff_B_p4sLLeAm1_2),.clk(gclk));
	jdff dff_B_oclFPpvi7_2(.din(w_dff_B_p4sLLeAm1_2),.dout(w_dff_B_oclFPpvi7_2),.clk(gclk));
	jdff dff_B_RnJwT5Ck2_2(.din(n1707),.dout(w_dff_B_RnJwT5Ck2_2),.clk(gclk));
	jdff dff_B_xUhWQ7P78_1(.din(n1705),.dout(w_dff_B_xUhWQ7P78_1),.clk(gclk));
	jdff dff_B_ZnUvd0pB6_2(.din(n1663),.dout(w_dff_B_ZnUvd0pB6_2),.clk(gclk));
	jdff dff_B_R1LkGii23_2(.din(w_dff_B_ZnUvd0pB6_2),.dout(w_dff_B_R1LkGii23_2),.clk(gclk));
	jdff dff_B_ue6fJH8d2_2(.din(w_dff_B_R1LkGii23_2),.dout(w_dff_B_ue6fJH8d2_2),.clk(gclk));
	jdff dff_B_uaUI1tya2_2(.din(w_dff_B_ue6fJH8d2_2),.dout(w_dff_B_uaUI1tya2_2),.clk(gclk));
	jdff dff_B_e0osTeAk0_2(.din(w_dff_B_uaUI1tya2_2),.dout(w_dff_B_e0osTeAk0_2),.clk(gclk));
	jdff dff_B_veltr0Mk4_2(.din(w_dff_B_e0osTeAk0_2),.dout(w_dff_B_veltr0Mk4_2),.clk(gclk));
	jdff dff_B_8I8ntM0i4_2(.din(w_dff_B_veltr0Mk4_2),.dout(w_dff_B_8I8ntM0i4_2),.clk(gclk));
	jdff dff_B_H8gDoiJq2_2(.din(w_dff_B_8I8ntM0i4_2),.dout(w_dff_B_H8gDoiJq2_2),.clk(gclk));
	jdff dff_B_1ZXJWgzi7_2(.din(w_dff_B_H8gDoiJq2_2),.dout(w_dff_B_1ZXJWgzi7_2),.clk(gclk));
	jdff dff_B_broJSCKl3_2(.din(w_dff_B_1ZXJWgzi7_2),.dout(w_dff_B_broJSCKl3_2),.clk(gclk));
	jdff dff_B_AF3h5rwq0_2(.din(w_dff_B_broJSCKl3_2),.dout(w_dff_B_AF3h5rwq0_2),.clk(gclk));
	jdff dff_B_NnnaeN9S3_2(.din(w_dff_B_AF3h5rwq0_2),.dout(w_dff_B_NnnaeN9S3_2),.clk(gclk));
	jdff dff_B_jJnSiXcb6_2(.din(w_dff_B_NnnaeN9S3_2),.dout(w_dff_B_jJnSiXcb6_2),.clk(gclk));
	jdff dff_B_0a4Am7YK2_2(.din(w_dff_B_jJnSiXcb6_2),.dout(w_dff_B_0a4Am7YK2_2),.clk(gclk));
	jdff dff_B_8cipSeC47_2(.din(w_dff_B_0a4Am7YK2_2),.dout(w_dff_B_8cipSeC47_2),.clk(gclk));
	jdff dff_B_54lBBl5N7_2(.din(w_dff_B_8cipSeC47_2),.dout(w_dff_B_54lBBl5N7_2),.clk(gclk));
	jdff dff_B_Ky4Z5DvP9_2(.din(w_dff_B_54lBBl5N7_2),.dout(w_dff_B_Ky4Z5DvP9_2),.clk(gclk));
	jdff dff_B_2ATFLZSG5_2(.din(w_dff_B_Ky4Z5DvP9_2),.dout(w_dff_B_2ATFLZSG5_2),.clk(gclk));
	jdff dff_B_Ge13u8Ls4_2(.din(w_dff_B_2ATFLZSG5_2),.dout(w_dff_B_Ge13u8Ls4_2),.clk(gclk));
	jdff dff_B_f1glNoIf6_2(.din(w_dff_B_Ge13u8Ls4_2),.dout(w_dff_B_f1glNoIf6_2),.clk(gclk));
	jdff dff_B_1NVNZibn5_2(.din(w_dff_B_f1glNoIf6_2),.dout(w_dff_B_1NVNZibn5_2),.clk(gclk));
	jdff dff_B_U5N9KqAq8_2(.din(w_dff_B_1NVNZibn5_2),.dout(w_dff_B_U5N9KqAq8_2),.clk(gclk));
	jdff dff_B_0ukPKVr16_2(.din(w_dff_B_U5N9KqAq8_2),.dout(w_dff_B_0ukPKVr16_2),.clk(gclk));
	jdff dff_B_Kk345oQU3_2(.din(w_dff_B_0ukPKVr16_2),.dout(w_dff_B_Kk345oQU3_2),.clk(gclk));
	jdff dff_B_6Y6NhmMw6_2(.din(w_dff_B_Kk345oQU3_2),.dout(w_dff_B_6Y6NhmMw6_2),.clk(gclk));
	jdff dff_B_wVowZGc66_2(.din(w_dff_B_6Y6NhmMw6_2),.dout(w_dff_B_wVowZGc66_2),.clk(gclk));
	jdff dff_B_g9yUQ3sO8_2(.din(w_dff_B_wVowZGc66_2),.dout(w_dff_B_g9yUQ3sO8_2),.clk(gclk));
	jdff dff_B_GZN7ssAe4_2(.din(w_dff_B_g9yUQ3sO8_2),.dout(w_dff_B_GZN7ssAe4_2),.clk(gclk));
	jdff dff_B_GyvGxgWo0_2(.din(w_dff_B_GZN7ssAe4_2),.dout(w_dff_B_GyvGxgWo0_2),.clk(gclk));
	jdff dff_B_TO8no1gk0_2(.din(w_dff_B_GyvGxgWo0_2),.dout(w_dff_B_TO8no1gk0_2),.clk(gclk));
	jdff dff_B_bzHPAJfm7_2(.din(w_dff_B_TO8no1gk0_2),.dout(w_dff_B_bzHPAJfm7_2),.clk(gclk));
	jdff dff_B_kZDfj2IH8_2(.din(w_dff_B_bzHPAJfm7_2),.dout(w_dff_B_kZDfj2IH8_2),.clk(gclk));
	jdff dff_B_ZKZeaSGl1_2(.din(w_dff_B_kZDfj2IH8_2),.dout(w_dff_B_ZKZeaSGl1_2),.clk(gclk));
	jdff dff_B_jWmgzRKY9_2(.din(w_dff_B_ZKZeaSGl1_2),.dout(w_dff_B_jWmgzRKY9_2),.clk(gclk));
	jdff dff_B_9yQ7bBTg6_2(.din(w_dff_B_jWmgzRKY9_2),.dout(w_dff_B_9yQ7bBTg6_2),.clk(gclk));
	jdff dff_B_0laUZmpq8_2(.din(w_dff_B_9yQ7bBTg6_2),.dout(w_dff_B_0laUZmpq8_2),.clk(gclk));
	jdff dff_B_VS1icB471_2(.din(w_dff_B_0laUZmpq8_2),.dout(w_dff_B_VS1icB471_2),.clk(gclk));
	jdff dff_B_7YdJci8z9_2(.din(w_dff_B_VS1icB471_2),.dout(w_dff_B_7YdJci8z9_2),.clk(gclk));
	jdff dff_B_VyMs4l4N2_2(.din(w_dff_B_7YdJci8z9_2),.dout(w_dff_B_VyMs4l4N2_2),.clk(gclk));
	jdff dff_B_NJPxzKL28_2(.din(w_dff_B_VyMs4l4N2_2),.dout(w_dff_B_NJPxzKL28_2),.clk(gclk));
	jdff dff_B_RVp14ZLk4_2(.din(w_dff_B_NJPxzKL28_2),.dout(w_dff_B_RVp14ZLk4_2),.clk(gclk));
	jdff dff_B_LZLyJm3j4_2(.din(w_dff_B_RVp14ZLk4_2),.dout(w_dff_B_LZLyJm3j4_2),.clk(gclk));
	jdff dff_B_ja0mBXim9_2(.din(n1666),.dout(w_dff_B_ja0mBXim9_2),.clk(gclk));
	jdff dff_B_Z3kybcKC3_1(.din(n1664),.dout(w_dff_B_Z3kybcKC3_1),.clk(gclk));
	jdff dff_B_OPVb36m03_2(.din(n1612),.dout(w_dff_B_OPVb36m03_2),.clk(gclk));
	jdff dff_B_9kUpg01B3_2(.din(w_dff_B_OPVb36m03_2),.dout(w_dff_B_9kUpg01B3_2),.clk(gclk));
	jdff dff_B_7YnxLA981_2(.din(w_dff_B_9kUpg01B3_2),.dout(w_dff_B_7YnxLA981_2),.clk(gclk));
	jdff dff_B_32w9rWTP6_2(.din(w_dff_B_7YnxLA981_2),.dout(w_dff_B_32w9rWTP6_2),.clk(gclk));
	jdff dff_B_MyQzIQD49_2(.din(w_dff_B_32w9rWTP6_2),.dout(w_dff_B_MyQzIQD49_2),.clk(gclk));
	jdff dff_B_3O83F5zh5_2(.din(w_dff_B_MyQzIQD49_2),.dout(w_dff_B_3O83F5zh5_2),.clk(gclk));
	jdff dff_B_086scwRj8_2(.din(w_dff_B_3O83F5zh5_2),.dout(w_dff_B_086scwRj8_2),.clk(gclk));
	jdff dff_B_zs3gKa1G6_2(.din(w_dff_B_086scwRj8_2),.dout(w_dff_B_zs3gKa1G6_2),.clk(gclk));
	jdff dff_B_0Elg8Dxi0_2(.din(w_dff_B_zs3gKa1G6_2),.dout(w_dff_B_0Elg8Dxi0_2),.clk(gclk));
	jdff dff_B_hBFSUMLP1_2(.din(w_dff_B_0Elg8Dxi0_2),.dout(w_dff_B_hBFSUMLP1_2),.clk(gclk));
	jdff dff_B_qr1wgGro3_2(.din(w_dff_B_hBFSUMLP1_2),.dout(w_dff_B_qr1wgGro3_2),.clk(gclk));
	jdff dff_B_R0e5yC4e2_2(.din(w_dff_B_qr1wgGro3_2),.dout(w_dff_B_R0e5yC4e2_2),.clk(gclk));
	jdff dff_B_QIYXvTD87_2(.din(w_dff_B_R0e5yC4e2_2),.dout(w_dff_B_QIYXvTD87_2),.clk(gclk));
	jdff dff_B_tjnddSiO0_2(.din(w_dff_B_QIYXvTD87_2),.dout(w_dff_B_tjnddSiO0_2),.clk(gclk));
	jdff dff_B_Cy7Xh06B4_2(.din(w_dff_B_tjnddSiO0_2),.dout(w_dff_B_Cy7Xh06B4_2),.clk(gclk));
	jdff dff_B_nEAQQnVQ1_2(.din(w_dff_B_Cy7Xh06B4_2),.dout(w_dff_B_nEAQQnVQ1_2),.clk(gclk));
	jdff dff_B_UwGJbpqU0_2(.din(w_dff_B_nEAQQnVQ1_2),.dout(w_dff_B_UwGJbpqU0_2),.clk(gclk));
	jdff dff_B_KIZ64XxM0_2(.din(w_dff_B_UwGJbpqU0_2),.dout(w_dff_B_KIZ64XxM0_2),.clk(gclk));
	jdff dff_B_nAeiZhqK3_2(.din(w_dff_B_KIZ64XxM0_2),.dout(w_dff_B_nAeiZhqK3_2),.clk(gclk));
	jdff dff_B_5hnQ81NF1_2(.din(w_dff_B_nAeiZhqK3_2),.dout(w_dff_B_5hnQ81NF1_2),.clk(gclk));
	jdff dff_B_ddA0HavY3_2(.din(w_dff_B_5hnQ81NF1_2),.dout(w_dff_B_ddA0HavY3_2),.clk(gclk));
	jdff dff_B_cChozTUg5_2(.din(w_dff_B_ddA0HavY3_2),.dout(w_dff_B_cChozTUg5_2),.clk(gclk));
	jdff dff_B_nL861Zk87_2(.din(w_dff_B_cChozTUg5_2),.dout(w_dff_B_nL861Zk87_2),.clk(gclk));
	jdff dff_B_54Vr9SM96_2(.din(w_dff_B_nL861Zk87_2),.dout(w_dff_B_54Vr9SM96_2),.clk(gclk));
	jdff dff_B_gKcCL3Xl1_2(.din(w_dff_B_54Vr9SM96_2),.dout(w_dff_B_gKcCL3Xl1_2),.clk(gclk));
	jdff dff_B_zIRcDqcF0_2(.din(w_dff_B_gKcCL3Xl1_2),.dout(w_dff_B_zIRcDqcF0_2),.clk(gclk));
	jdff dff_B_ZWSCqcPd2_2(.din(w_dff_B_zIRcDqcF0_2),.dout(w_dff_B_ZWSCqcPd2_2),.clk(gclk));
	jdff dff_B_ydOqIiGX8_2(.din(w_dff_B_ZWSCqcPd2_2),.dout(w_dff_B_ydOqIiGX8_2),.clk(gclk));
	jdff dff_B_tqmGzePz4_2(.din(w_dff_B_ydOqIiGX8_2),.dout(w_dff_B_tqmGzePz4_2),.clk(gclk));
	jdff dff_B_00CjC6pd0_2(.din(w_dff_B_tqmGzePz4_2),.dout(w_dff_B_00CjC6pd0_2),.clk(gclk));
	jdff dff_B_zNqGBlgz3_2(.din(w_dff_B_00CjC6pd0_2),.dout(w_dff_B_zNqGBlgz3_2),.clk(gclk));
	jdff dff_B_mBDjjgkK8_2(.din(w_dff_B_zNqGBlgz3_2),.dout(w_dff_B_mBDjjgkK8_2),.clk(gclk));
	jdff dff_B_gLRzJdOx1_2(.din(w_dff_B_mBDjjgkK8_2),.dout(w_dff_B_gLRzJdOx1_2),.clk(gclk));
	jdff dff_B_5oC21Aiy7_2(.din(w_dff_B_gLRzJdOx1_2),.dout(w_dff_B_5oC21Aiy7_2),.clk(gclk));
	jdff dff_B_iGR8yivS8_2(.din(w_dff_B_5oC21Aiy7_2),.dout(w_dff_B_iGR8yivS8_2),.clk(gclk));
	jdff dff_B_xOLGpIMd0_2(.din(w_dff_B_iGR8yivS8_2),.dout(w_dff_B_xOLGpIMd0_2),.clk(gclk));
	jdff dff_B_JrgDec5g1_2(.din(w_dff_B_xOLGpIMd0_2),.dout(w_dff_B_JrgDec5g1_2),.clk(gclk));
	jdff dff_B_xoIVA3GF0_2(.din(w_dff_B_JrgDec5g1_2),.dout(w_dff_B_xoIVA3GF0_2),.clk(gclk));
	jdff dff_B_91rMqHuE3_2(.din(n1615),.dout(w_dff_B_91rMqHuE3_2),.clk(gclk));
	jdff dff_B_WCqwlkD57_1(.din(n1613),.dout(w_dff_B_WCqwlkD57_1),.clk(gclk));
	jdff dff_B_fPiuv2cm9_2(.din(n1555),.dout(w_dff_B_fPiuv2cm9_2),.clk(gclk));
	jdff dff_B_RcopoAdc6_2(.din(w_dff_B_fPiuv2cm9_2),.dout(w_dff_B_RcopoAdc6_2),.clk(gclk));
	jdff dff_B_AZlF2ya14_2(.din(w_dff_B_RcopoAdc6_2),.dout(w_dff_B_AZlF2ya14_2),.clk(gclk));
	jdff dff_B_fW15ihs65_2(.din(w_dff_B_AZlF2ya14_2),.dout(w_dff_B_fW15ihs65_2),.clk(gclk));
	jdff dff_B_zn8AjPi58_2(.din(w_dff_B_fW15ihs65_2),.dout(w_dff_B_zn8AjPi58_2),.clk(gclk));
	jdff dff_B_NRHqG14d8_2(.din(w_dff_B_zn8AjPi58_2),.dout(w_dff_B_NRHqG14d8_2),.clk(gclk));
	jdff dff_B_6WgsknMI6_2(.din(w_dff_B_NRHqG14d8_2),.dout(w_dff_B_6WgsknMI6_2),.clk(gclk));
	jdff dff_B_8sMMocFp3_2(.din(w_dff_B_6WgsknMI6_2),.dout(w_dff_B_8sMMocFp3_2),.clk(gclk));
	jdff dff_B_yktOetWv2_2(.din(w_dff_B_8sMMocFp3_2),.dout(w_dff_B_yktOetWv2_2),.clk(gclk));
	jdff dff_B_bvoWQD3B5_2(.din(w_dff_B_yktOetWv2_2),.dout(w_dff_B_bvoWQD3B5_2),.clk(gclk));
	jdff dff_B_XFc5KKgL0_2(.din(w_dff_B_bvoWQD3B5_2),.dout(w_dff_B_XFc5KKgL0_2),.clk(gclk));
	jdff dff_B_rt4W2dJk9_2(.din(w_dff_B_XFc5KKgL0_2),.dout(w_dff_B_rt4W2dJk9_2),.clk(gclk));
	jdff dff_B_fY2z0SjK8_2(.din(w_dff_B_rt4W2dJk9_2),.dout(w_dff_B_fY2z0SjK8_2),.clk(gclk));
	jdff dff_B_P7Q2Tp9n5_2(.din(w_dff_B_fY2z0SjK8_2),.dout(w_dff_B_P7Q2Tp9n5_2),.clk(gclk));
	jdff dff_B_TdWZf15q6_2(.din(w_dff_B_P7Q2Tp9n5_2),.dout(w_dff_B_TdWZf15q6_2),.clk(gclk));
	jdff dff_B_mpEPL3kk2_2(.din(w_dff_B_TdWZf15q6_2),.dout(w_dff_B_mpEPL3kk2_2),.clk(gclk));
	jdff dff_B_4drblbfP0_2(.din(w_dff_B_mpEPL3kk2_2),.dout(w_dff_B_4drblbfP0_2),.clk(gclk));
	jdff dff_B_sIZefvHT4_2(.din(w_dff_B_4drblbfP0_2),.dout(w_dff_B_sIZefvHT4_2),.clk(gclk));
	jdff dff_B_OsScXjat3_2(.din(w_dff_B_sIZefvHT4_2),.dout(w_dff_B_OsScXjat3_2),.clk(gclk));
	jdff dff_B_gWnmwcgo4_2(.din(w_dff_B_OsScXjat3_2),.dout(w_dff_B_gWnmwcgo4_2),.clk(gclk));
	jdff dff_B_9TslwpQo4_2(.din(w_dff_B_gWnmwcgo4_2),.dout(w_dff_B_9TslwpQo4_2),.clk(gclk));
	jdff dff_B_aOYXxL9T3_2(.din(w_dff_B_9TslwpQo4_2),.dout(w_dff_B_aOYXxL9T3_2),.clk(gclk));
	jdff dff_B_aThpX9yG3_2(.din(w_dff_B_aOYXxL9T3_2),.dout(w_dff_B_aThpX9yG3_2),.clk(gclk));
	jdff dff_B_2tr2JhNf2_2(.din(w_dff_B_aThpX9yG3_2),.dout(w_dff_B_2tr2JhNf2_2),.clk(gclk));
	jdff dff_B_xdjcD8ek1_2(.din(w_dff_B_2tr2JhNf2_2),.dout(w_dff_B_xdjcD8ek1_2),.clk(gclk));
	jdff dff_B_ZUBg0cdR5_2(.din(w_dff_B_xdjcD8ek1_2),.dout(w_dff_B_ZUBg0cdR5_2),.clk(gclk));
	jdff dff_B_enfe3FSn1_2(.din(w_dff_B_ZUBg0cdR5_2),.dout(w_dff_B_enfe3FSn1_2),.clk(gclk));
	jdff dff_B_lWoPGZ4f7_2(.din(w_dff_B_enfe3FSn1_2),.dout(w_dff_B_lWoPGZ4f7_2),.clk(gclk));
	jdff dff_B_yOe9LVJR5_2(.din(w_dff_B_lWoPGZ4f7_2),.dout(w_dff_B_yOe9LVJR5_2),.clk(gclk));
	jdff dff_B_LIjf5T790_2(.din(w_dff_B_yOe9LVJR5_2),.dout(w_dff_B_LIjf5T790_2),.clk(gclk));
	jdff dff_B_lBz3PMqb0_2(.din(w_dff_B_LIjf5T790_2),.dout(w_dff_B_lBz3PMqb0_2),.clk(gclk));
	jdff dff_B_r7CUCfbe3_2(.din(w_dff_B_lBz3PMqb0_2),.dout(w_dff_B_r7CUCfbe3_2),.clk(gclk));
	jdff dff_B_TBk6PQ0Z0_2(.din(w_dff_B_r7CUCfbe3_2),.dout(w_dff_B_TBk6PQ0Z0_2),.clk(gclk));
	jdff dff_B_RkwElSTr3_2(.din(w_dff_B_TBk6PQ0Z0_2),.dout(w_dff_B_RkwElSTr3_2),.clk(gclk));
	jdff dff_B_gP79HKPg5_2(.din(n1558),.dout(w_dff_B_gP79HKPg5_2),.clk(gclk));
	jdff dff_B_C2oGLTtB5_1(.din(n1556),.dout(w_dff_B_C2oGLTtB5_1),.clk(gclk));
	jdff dff_B_av488jlZ9_2(.din(n1491),.dout(w_dff_B_av488jlZ9_2),.clk(gclk));
	jdff dff_B_qXkxlrXA3_2(.din(w_dff_B_av488jlZ9_2),.dout(w_dff_B_qXkxlrXA3_2),.clk(gclk));
	jdff dff_B_zknPNhha5_2(.din(w_dff_B_qXkxlrXA3_2),.dout(w_dff_B_zknPNhha5_2),.clk(gclk));
	jdff dff_B_d1irbzPu0_2(.din(w_dff_B_zknPNhha5_2),.dout(w_dff_B_d1irbzPu0_2),.clk(gclk));
	jdff dff_B_lRuSyQre1_2(.din(w_dff_B_d1irbzPu0_2),.dout(w_dff_B_lRuSyQre1_2),.clk(gclk));
	jdff dff_B_w5oOZ97R7_2(.din(w_dff_B_lRuSyQre1_2),.dout(w_dff_B_w5oOZ97R7_2),.clk(gclk));
	jdff dff_B_Dgu7PPXC1_2(.din(w_dff_B_w5oOZ97R7_2),.dout(w_dff_B_Dgu7PPXC1_2),.clk(gclk));
	jdff dff_B_uyoNLxOB3_2(.din(w_dff_B_Dgu7PPXC1_2),.dout(w_dff_B_uyoNLxOB3_2),.clk(gclk));
	jdff dff_B_zzqO8dRf2_2(.din(w_dff_B_uyoNLxOB3_2),.dout(w_dff_B_zzqO8dRf2_2),.clk(gclk));
	jdff dff_B_R4IDc1Fl4_2(.din(w_dff_B_zzqO8dRf2_2),.dout(w_dff_B_R4IDc1Fl4_2),.clk(gclk));
	jdff dff_B_9Q1NfQnx7_2(.din(w_dff_B_R4IDc1Fl4_2),.dout(w_dff_B_9Q1NfQnx7_2),.clk(gclk));
	jdff dff_B_XUEJ55j08_2(.din(w_dff_B_9Q1NfQnx7_2),.dout(w_dff_B_XUEJ55j08_2),.clk(gclk));
	jdff dff_B_IyDbQTbd1_2(.din(w_dff_B_XUEJ55j08_2),.dout(w_dff_B_IyDbQTbd1_2),.clk(gclk));
	jdff dff_B_IhbNuhZ40_2(.din(w_dff_B_IyDbQTbd1_2),.dout(w_dff_B_IhbNuhZ40_2),.clk(gclk));
	jdff dff_B_LJ65Cxe72_2(.din(w_dff_B_IhbNuhZ40_2),.dout(w_dff_B_LJ65Cxe72_2),.clk(gclk));
	jdff dff_B_EsacYrXN3_2(.din(w_dff_B_LJ65Cxe72_2),.dout(w_dff_B_EsacYrXN3_2),.clk(gclk));
	jdff dff_B_ScNGK3SD7_2(.din(w_dff_B_EsacYrXN3_2),.dout(w_dff_B_ScNGK3SD7_2),.clk(gclk));
	jdff dff_B_lk13Ztqe3_2(.din(w_dff_B_ScNGK3SD7_2),.dout(w_dff_B_lk13Ztqe3_2),.clk(gclk));
	jdff dff_B_9GJa4h0v1_2(.din(w_dff_B_lk13Ztqe3_2),.dout(w_dff_B_9GJa4h0v1_2),.clk(gclk));
	jdff dff_B_VnAcH8bm7_2(.din(w_dff_B_9GJa4h0v1_2),.dout(w_dff_B_VnAcH8bm7_2),.clk(gclk));
	jdff dff_B_gxnA3I7a1_2(.din(w_dff_B_VnAcH8bm7_2),.dout(w_dff_B_gxnA3I7a1_2),.clk(gclk));
	jdff dff_B_jfJLPkd41_2(.din(w_dff_B_gxnA3I7a1_2),.dout(w_dff_B_jfJLPkd41_2),.clk(gclk));
	jdff dff_B_FqDvi7Zh3_2(.din(w_dff_B_jfJLPkd41_2),.dout(w_dff_B_FqDvi7Zh3_2),.clk(gclk));
	jdff dff_B_AWigrkcm2_2(.din(w_dff_B_FqDvi7Zh3_2),.dout(w_dff_B_AWigrkcm2_2),.clk(gclk));
	jdff dff_B_49wzTS1w4_2(.din(w_dff_B_AWigrkcm2_2),.dout(w_dff_B_49wzTS1w4_2),.clk(gclk));
	jdff dff_B_3fSRVEIg5_2(.din(w_dff_B_49wzTS1w4_2),.dout(w_dff_B_3fSRVEIg5_2),.clk(gclk));
	jdff dff_B_3WbzAvAo2_2(.din(w_dff_B_3fSRVEIg5_2),.dout(w_dff_B_3WbzAvAo2_2),.clk(gclk));
	jdff dff_B_ct5dX4hf7_2(.din(w_dff_B_3WbzAvAo2_2),.dout(w_dff_B_ct5dX4hf7_2),.clk(gclk));
	jdff dff_B_XnLifrND1_2(.din(w_dff_B_ct5dX4hf7_2),.dout(w_dff_B_XnLifrND1_2),.clk(gclk));
	jdff dff_B_88iN42Kq8_2(.din(w_dff_B_XnLifrND1_2),.dout(w_dff_B_88iN42Kq8_2),.clk(gclk));
	jdff dff_B_cP8Rbmyk5_2(.din(n1494),.dout(w_dff_B_cP8Rbmyk5_2),.clk(gclk));
	jdff dff_B_I86KhtRw2_1(.din(n1492),.dout(w_dff_B_I86KhtRw2_1),.clk(gclk));
	jdff dff_B_ju7W2gGp6_2(.din(n1420),.dout(w_dff_B_ju7W2gGp6_2),.clk(gclk));
	jdff dff_B_yIS7eXoJ0_2(.din(w_dff_B_ju7W2gGp6_2),.dout(w_dff_B_yIS7eXoJ0_2),.clk(gclk));
	jdff dff_B_seK5TP5Z9_2(.din(w_dff_B_yIS7eXoJ0_2),.dout(w_dff_B_seK5TP5Z9_2),.clk(gclk));
	jdff dff_B_GMiotzNZ0_2(.din(w_dff_B_seK5TP5Z9_2),.dout(w_dff_B_GMiotzNZ0_2),.clk(gclk));
	jdff dff_B_HxEAuNNN4_2(.din(w_dff_B_GMiotzNZ0_2),.dout(w_dff_B_HxEAuNNN4_2),.clk(gclk));
	jdff dff_B_D41Uv9zD2_2(.din(w_dff_B_HxEAuNNN4_2),.dout(w_dff_B_D41Uv9zD2_2),.clk(gclk));
	jdff dff_B_yO5d1ktJ2_2(.din(w_dff_B_D41Uv9zD2_2),.dout(w_dff_B_yO5d1ktJ2_2),.clk(gclk));
	jdff dff_B_fGhgf1iw8_2(.din(w_dff_B_yO5d1ktJ2_2),.dout(w_dff_B_fGhgf1iw8_2),.clk(gclk));
	jdff dff_B_8la4JtVp2_2(.din(w_dff_B_fGhgf1iw8_2),.dout(w_dff_B_8la4JtVp2_2),.clk(gclk));
	jdff dff_B_jE1vvOdw8_2(.din(w_dff_B_8la4JtVp2_2),.dout(w_dff_B_jE1vvOdw8_2),.clk(gclk));
	jdff dff_B_U47nJWp36_2(.din(w_dff_B_jE1vvOdw8_2),.dout(w_dff_B_U47nJWp36_2),.clk(gclk));
	jdff dff_B_pHgLMOTn8_2(.din(w_dff_B_U47nJWp36_2),.dout(w_dff_B_pHgLMOTn8_2),.clk(gclk));
	jdff dff_B_H8y7XJcP4_2(.din(w_dff_B_pHgLMOTn8_2),.dout(w_dff_B_H8y7XJcP4_2),.clk(gclk));
	jdff dff_B_yWJydMai0_2(.din(w_dff_B_H8y7XJcP4_2),.dout(w_dff_B_yWJydMai0_2),.clk(gclk));
	jdff dff_B_QtzlR6zi2_2(.din(w_dff_B_yWJydMai0_2),.dout(w_dff_B_QtzlR6zi2_2),.clk(gclk));
	jdff dff_B_OHufHraA4_2(.din(w_dff_B_QtzlR6zi2_2),.dout(w_dff_B_OHufHraA4_2),.clk(gclk));
	jdff dff_B_qfwGkaqB7_2(.din(w_dff_B_OHufHraA4_2),.dout(w_dff_B_qfwGkaqB7_2),.clk(gclk));
	jdff dff_B_noSn6UwS4_2(.din(w_dff_B_qfwGkaqB7_2),.dout(w_dff_B_noSn6UwS4_2),.clk(gclk));
	jdff dff_B_8lQtiQRp3_2(.din(w_dff_B_noSn6UwS4_2),.dout(w_dff_B_8lQtiQRp3_2),.clk(gclk));
	jdff dff_B_0wOwqwwg6_2(.din(w_dff_B_8lQtiQRp3_2),.dout(w_dff_B_0wOwqwwg6_2),.clk(gclk));
	jdff dff_B_ZsPoO47b0_2(.din(w_dff_B_0wOwqwwg6_2),.dout(w_dff_B_ZsPoO47b0_2),.clk(gclk));
	jdff dff_B_tlnucIfU0_2(.din(w_dff_B_ZsPoO47b0_2),.dout(w_dff_B_tlnucIfU0_2),.clk(gclk));
	jdff dff_B_q8hU2th87_2(.din(w_dff_B_tlnucIfU0_2),.dout(w_dff_B_q8hU2th87_2),.clk(gclk));
	jdff dff_B_lFseBrOB9_2(.din(w_dff_B_q8hU2th87_2),.dout(w_dff_B_lFseBrOB9_2),.clk(gclk));
	jdff dff_B_UbOE9IND1_2(.din(w_dff_B_lFseBrOB9_2),.dout(w_dff_B_UbOE9IND1_2),.clk(gclk));
	jdff dff_B_3uQSKymP1_2(.din(w_dff_B_UbOE9IND1_2),.dout(w_dff_B_3uQSKymP1_2),.clk(gclk));
	jdff dff_B_LJDxjFoi4_1(.din(n1421),.dout(w_dff_B_LJDxjFoi4_1),.clk(gclk));
	jdff dff_B_08VVXDkH0_2(.din(n1342),.dout(w_dff_B_08VVXDkH0_2),.clk(gclk));
	jdff dff_B_O4F29F054_2(.din(w_dff_B_08VVXDkH0_2),.dout(w_dff_B_O4F29F054_2),.clk(gclk));
	jdff dff_B_Dmc46R6q7_2(.din(w_dff_B_O4F29F054_2),.dout(w_dff_B_Dmc46R6q7_2),.clk(gclk));
	jdff dff_B_S7GON89R7_2(.din(w_dff_B_Dmc46R6q7_2),.dout(w_dff_B_S7GON89R7_2),.clk(gclk));
	jdff dff_B_zSLUxsei5_2(.din(w_dff_B_S7GON89R7_2),.dout(w_dff_B_zSLUxsei5_2),.clk(gclk));
	jdff dff_B_YDt6z6cg9_2(.din(w_dff_B_zSLUxsei5_2),.dout(w_dff_B_YDt6z6cg9_2),.clk(gclk));
	jdff dff_B_M1yvTjJl5_2(.din(w_dff_B_YDt6z6cg9_2),.dout(w_dff_B_M1yvTjJl5_2),.clk(gclk));
	jdff dff_B_az8E3v9g6_2(.din(w_dff_B_M1yvTjJl5_2),.dout(w_dff_B_az8E3v9g6_2),.clk(gclk));
	jdff dff_B_tAq2IbZl3_2(.din(w_dff_B_az8E3v9g6_2),.dout(w_dff_B_tAq2IbZl3_2),.clk(gclk));
	jdff dff_B_J5e5KFVe2_2(.din(w_dff_B_tAq2IbZl3_2),.dout(w_dff_B_J5e5KFVe2_2),.clk(gclk));
	jdff dff_B_lTrmwefs6_2(.din(w_dff_B_J5e5KFVe2_2),.dout(w_dff_B_lTrmwefs6_2),.clk(gclk));
	jdff dff_B_7AByAONw9_2(.din(w_dff_B_lTrmwefs6_2),.dout(w_dff_B_7AByAONw9_2),.clk(gclk));
	jdff dff_B_ILkibUJj7_2(.din(w_dff_B_7AByAONw9_2),.dout(w_dff_B_ILkibUJj7_2),.clk(gclk));
	jdff dff_B_WtOB8IT22_2(.din(w_dff_B_ILkibUJj7_2),.dout(w_dff_B_WtOB8IT22_2),.clk(gclk));
	jdff dff_B_ZzF7ou968_2(.din(w_dff_B_WtOB8IT22_2),.dout(w_dff_B_ZzF7ou968_2),.clk(gclk));
	jdff dff_B_V6qDCgDl4_2(.din(w_dff_B_ZzF7ou968_2),.dout(w_dff_B_V6qDCgDl4_2),.clk(gclk));
	jdff dff_B_IoDUvnMM0_2(.din(w_dff_B_V6qDCgDl4_2),.dout(w_dff_B_IoDUvnMM0_2),.clk(gclk));
	jdff dff_B_CdBOnoWr5_2(.din(w_dff_B_IoDUvnMM0_2),.dout(w_dff_B_CdBOnoWr5_2),.clk(gclk));
	jdff dff_B_HA0nb6ci8_2(.din(w_dff_B_CdBOnoWr5_2),.dout(w_dff_B_HA0nb6ci8_2),.clk(gclk));
	jdff dff_B_rvlZNm1Z6_2(.din(w_dff_B_HA0nb6ci8_2),.dout(w_dff_B_rvlZNm1Z6_2),.clk(gclk));
	jdff dff_B_K72b4cU16_2(.din(w_dff_B_rvlZNm1Z6_2),.dout(w_dff_B_K72b4cU16_2),.clk(gclk));
	jdff dff_B_qNrSSy3u2_2(.din(w_dff_B_K72b4cU16_2),.dout(w_dff_B_qNrSSy3u2_2),.clk(gclk));
	jdff dff_B_QUpBqD0A6_2(.din(w_dff_B_qNrSSy3u2_2),.dout(w_dff_B_QUpBqD0A6_2),.clk(gclk));
	jdff dff_B_72tu2LAE3_2(.din(n1360),.dout(w_dff_B_72tu2LAE3_2),.clk(gclk));
	jdff dff_B_5mHjtuOZ5_1(.din(n1343),.dout(w_dff_B_5mHjtuOZ5_1),.clk(gclk));
	jdff dff_B_73sBYgZK7_2(.din(n1257),.dout(w_dff_B_73sBYgZK7_2),.clk(gclk));
	jdff dff_B_HXBvKebs7_2(.din(w_dff_B_73sBYgZK7_2),.dout(w_dff_B_HXBvKebs7_2),.clk(gclk));
	jdff dff_B_NmKTxOY83_2(.din(w_dff_B_HXBvKebs7_2),.dout(w_dff_B_NmKTxOY83_2),.clk(gclk));
	jdff dff_B_ZqNRnkbi7_2(.din(w_dff_B_NmKTxOY83_2),.dout(w_dff_B_ZqNRnkbi7_2),.clk(gclk));
	jdff dff_B_cBfevwWd8_2(.din(w_dff_B_ZqNRnkbi7_2),.dout(w_dff_B_cBfevwWd8_2),.clk(gclk));
	jdff dff_B_QR1ydtWC1_2(.din(w_dff_B_cBfevwWd8_2),.dout(w_dff_B_QR1ydtWC1_2),.clk(gclk));
	jdff dff_B_eO9swGgq0_2(.din(w_dff_B_QR1ydtWC1_2),.dout(w_dff_B_eO9swGgq0_2),.clk(gclk));
	jdff dff_B_2iXHiTP31_2(.din(w_dff_B_eO9swGgq0_2),.dout(w_dff_B_2iXHiTP31_2),.clk(gclk));
	jdff dff_B_VXM7YLfv8_2(.din(w_dff_B_2iXHiTP31_2),.dout(w_dff_B_VXM7YLfv8_2),.clk(gclk));
	jdff dff_B_ythenOWD3_2(.din(w_dff_B_VXM7YLfv8_2),.dout(w_dff_B_ythenOWD3_2),.clk(gclk));
	jdff dff_B_Pdn9LChg6_2(.din(w_dff_B_ythenOWD3_2),.dout(w_dff_B_Pdn9LChg6_2),.clk(gclk));
	jdff dff_B_m4jRz59K9_2(.din(w_dff_B_Pdn9LChg6_2),.dout(w_dff_B_m4jRz59K9_2),.clk(gclk));
	jdff dff_B_EAkevS0z0_2(.din(w_dff_B_m4jRz59K9_2),.dout(w_dff_B_EAkevS0z0_2),.clk(gclk));
	jdff dff_B_2kJUwQqd0_2(.din(w_dff_B_EAkevS0z0_2),.dout(w_dff_B_2kJUwQqd0_2),.clk(gclk));
	jdff dff_B_NJbB9n1W7_2(.din(w_dff_B_2kJUwQqd0_2),.dout(w_dff_B_NJbB9n1W7_2),.clk(gclk));
	jdff dff_B_iSHyyvDm5_2(.din(w_dff_B_NJbB9n1W7_2),.dout(w_dff_B_iSHyyvDm5_2),.clk(gclk));
	jdff dff_B_8wbRfNYU4_2(.din(w_dff_B_iSHyyvDm5_2),.dout(w_dff_B_8wbRfNYU4_2),.clk(gclk));
	jdff dff_B_YVpeK3cy7_2(.din(w_dff_B_8wbRfNYU4_2),.dout(w_dff_B_YVpeK3cy7_2),.clk(gclk));
	jdff dff_B_h00hxkZJ6_2(.din(w_dff_B_YVpeK3cy7_2),.dout(w_dff_B_h00hxkZJ6_2),.clk(gclk));
	jdff dff_B_wQxdIANl7_2(.din(w_dff_B_h00hxkZJ6_2),.dout(w_dff_B_wQxdIANl7_2),.clk(gclk));
	jdff dff_B_bXuZ2R9U2_2(.din(n1275),.dout(w_dff_B_bXuZ2R9U2_2),.clk(gclk));
	jdff dff_B_QNM7Qz8B1_1(.din(n1258),.dout(w_dff_B_QNM7Qz8B1_1),.clk(gclk));
	jdff dff_B_DxcT5UY99_2(.din(n1166),.dout(w_dff_B_DxcT5UY99_2),.clk(gclk));
	jdff dff_B_BTaoT8Xu8_2(.din(w_dff_B_DxcT5UY99_2),.dout(w_dff_B_BTaoT8Xu8_2),.clk(gclk));
	jdff dff_B_fGl5cl8s6_2(.din(w_dff_B_BTaoT8Xu8_2),.dout(w_dff_B_fGl5cl8s6_2),.clk(gclk));
	jdff dff_B_7ppeqsrN5_2(.din(w_dff_B_fGl5cl8s6_2),.dout(w_dff_B_7ppeqsrN5_2),.clk(gclk));
	jdff dff_B_vj44D1I42_2(.din(w_dff_B_7ppeqsrN5_2),.dout(w_dff_B_vj44D1I42_2),.clk(gclk));
	jdff dff_B_0G1sA9Pt8_2(.din(w_dff_B_vj44D1I42_2),.dout(w_dff_B_0G1sA9Pt8_2),.clk(gclk));
	jdff dff_B_DLbnZe7g7_2(.din(w_dff_B_0G1sA9Pt8_2),.dout(w_dff_B_DLbnZe7g7_2),.clk(gclk));
	jdff dff_B_8VQDqMGD3_2(.din(w_dff_B_DLbnZe7g7_2),.dout(w_dff_B_8VQDqMGD3_2),.clk(gclk));
	jdff dff_B_tgA1Zv524_2(.din(w_dff_B_8VQDqMGD3_2),.dout(w_dff_B_tgA1Zv524_2),.clk(gclk));
	jdff dff_B_bS3Fn67k7_2(.din(w_dff_B_tgA1Zv524_2),.dout(w_dff_B_bS3Fn67k7_2),.clk(gclk));
	jdff dff_B_7gA6ZETQ1_2(.din(w_dff_B_bS3Fn67k7_2),.dout(w_dff_B_7gA6ZETQ1_2),.clk(gclk));
	jdff dff_B_khCf8RYj8_2(.din(w_dff_B_7gA6ZETQ1_2),.dout(w_dff_B_khCf8RYj8_2),.clk(gclk));
	jdff dff_B_c0iKoziR7_2(.din(w_dff_B_khCf8RYj8_2),.dout(w_dff_B_c0iKoziR7_2),.clk(gclk));
	jdff dff_B_ZghivQ114_2(.din(w_dff_B_c0iKoziR7_2),.dout(w_dff_B_ZghivQ114_2),.clk(gclk));
	jdff dff_B_5Z0tHiZu1_2(.din(w_dff_B_ZghivQ114_2),.dout(w_dff_B_5Z0tHiZu1_2),.clk(gclk));
	jdff dff_B_iPUyH3sg7_2(.din(w_dff_B_5Z0tHiZu1_2),.dout(w_dff_B_iPUyH3sg7_2),.clk(gclk));
	jdff dff_B_0fgYsl7M7_2(.din(w_dff_B_iPUyH3sg7_2),.dout(w_dff_B_0fgYsl7M7_2),.clk(gclk));
	jdff dff_B_FbDURwN55_2(.din(n1184),.dout(w_dff_B_FbDURwN55_2),.clk(gclk));
	jdff dff_B_w6HJXtga9_1(.din(n1167),.dout(w_dff_B_w6HJXtga9_1),.clk(gclk));
	jdff dff_B_vtMewbRc0_2(.din(n1068),.dout(w_dff_B_vtMewbRc0_2),.clk(gclk));
	jdff dff_B_cX7EzFbw1_2(.din(w_dff_B_vtMewbRc0_2),.dout(w_dff_B_cX7EzFbw1_2),.clk(gclk));
	jdff dff_B_oG3RKuPe3_2(.din(w_dff_B_cX7EzFbw1_2),.dout(w_dff_B_oG3RKuPe3_2),.clk(gclk));
	jdff dff_B_Uy5KFX1F9_2(.din(w_dff_B_oG3RKuPe3_2),.dout(w_dff_B_Uy5KFX1F9_2),.clk(gclk));
	jdff dff_B_S6rwYapD8_2(.din(w_dff_B_Uy5KFX1F9_2),.dout(w_dff_B_S6rwYapD8_2),.clk(gclk));
	jdff dff_B_kzjhLKBF6_2(.din(w_dff_B_S6rwYapD8_2),.dout(w_dff_B_kzjhLKBF6_2),.clk(gclk));
	jdff dff_B_92IMJ7ZM2_2(.din(w_dff_B_kzjhLKBF6_2),.dout(w_dff_B_92IMJ7ZM2_2),.clk(gclk));
	jdff dff_B_iUbH7IrW8_2(.din(w_dff_B_92IMJ7ZM2_2),.dout(w_dff_B_iUbH7IrW8_2),.clk(gclk));
	jdff dff_B_FvDLb4XM7_2(.din(w_dff_B_iUbH7IrW8_2),.dout(w_dff_B_FvDLb4XM7_2),.clk(gclk));
	jdff dff_B_qWN1ySMt7_2(.din(w_dff_B_FvDLb4XM7_2),.dout(w_dff_B_qWN1ySMt7_2),.clk(gclk));
	jdff dff_B_I145K9kq6_2(.din(w_dff_B_qWN1ySMt7_2),.dout(w_dff_B_I145K9kq6_2),.clk(gclk));
	jdff dff_B_2XSfBDqh9_2(.din(w_dff_B_I145K9kq6_2),.dout(w_dff_B_2XSfBDqh9_2),.clk(gclk));
	jdff dff_B_7BEK49uK1_2(.din(w_dff_B_2XSfBDqh9_2),.dout(w_dff_B_7BEK49uK1_2),.clk(gclk));
	jdff dff_B_VfNDgjQa5_2(.din(w_dff_B_7BEK49uK1_2),.dout(w_dff_B_VfNDgjQa5_2),.clk(gclk));
	jdff dff_B_bFThtfdB8_2(.din(n1085),.dout(w_dff_B_bFThtfdB8_2),.clk(gclk));
	jdff dff_B_zz5olJJm3_1(.din(n1069),.dout(w_dff_B_zz5olJJm3_1),.clk(gclk));
	jdff dff_B_mOWuvJG62_2(.din(n969),.dout(w_dff_B_mOWuvJG62_2),.clk(gclk));
	jdff dff_B_WieyFUj92_2(.din(w_dff_B_mOWuvJG62_2),.dout(w_dff_B_WieyFUj92_2),.clk(gclk));
	jdff dff_B_oJvtDd4k6_2(.din(w_dff_B_WieyFUj92_2),.dout(w_dff_B_oJvtDd4k6_2),.clk(gclk));
	jdff dff_B_VEVvxzre2_2(.din(w_dff_B_oJvtDd4k6_2),.dout(w_dff_B_VEVvxzre2_2),.clk(gclk));
	jdff dff_B_IOgruZrP8_2(.din(w_dff_B_VEVvxzre2_2),.dout(w_dff_B_IOgruZrP8_2),.clk(gclk));
	jdff dff_B_cwBUrJLP2_2(.din(w_dff_B_IOgruZrP8_2),.dout(w_dff_B_cwBUrJLP2_2),.clk(gclk));
	jdff dff_B_BERuTnDO0_2(.din(w_dff_B_cwBUrJLP2_2),.dout(w_dff_B_BERuTnDO0_2),.clk(gclk));
	jdff dff_B_9RCoXGYh5_2(.din(w_dff_B_BERuTnDO0_2),.dout(w_dff_B_9RCoXGYh5_2),.clk(gclk));
	jdff dff_B_cGp6XCah9_2(.din(w_dff_B_9RCoXGYh5_2),.dout(w_dff_B_cGp6XCah9_2),.clk(gclk));
	jdff dff_B_dS5O7xwN9_2(.din(w_dff_B_cGp6XCah9_2),.dout(w_dff_B_dS5O7xwN9_2),.clk(gclk));
	jdff dff_B_4ShqpVAq3_2(.din(w_dff_B_dS5O7xwN9_2),.dout(w_dff_B_4ShqpVAq3_2),.clk(gclk));
	jdff dff_B_5E2IGDSn9_2(.din(n986),.dout(w_dff_B_5E2IGDSn9_2),.clk(gclk));
	jdff dff_B_KaaAk79D5_1(.din(n970),.dout(w_dff_B_KaaAk79D5_1),.clk(gclk));
	jdff dff_B_yF3ObJhE0_2(.din(n867),.dout(w_dff_B_yF3ObJhE0_2),.clk(gclk));
	jdff dff_B_BjUNqUy12_2(.din(w_dff_B_yF3ObJhE0_2),.dout(w_dff_B_BjUNqUy12_2),.clk(gclk));
	jdff dff_B_NzqfFX740_2(.din(w_dff_B_BjUNqUy12_2),.dout(w_dff_B_NzqfFX740_2),.clk(gclk));
	jdff dff_B_vte77m381_2(.din(w_dff_B_NzqfFX740_2),.dout(w_dff_B_vte77m381_2),.clk(gclk));
	jdff dff_B_HohZjWKK4_2(.din(w_dff_B_vte77m381_2),.dout(w_dff_B_HohZjWKK4_2),.clk(gclk));
	jdff dff_B_7HnIj5zW7_2(.din(w_dff_B_HohZjWKK4_2),.dout(w_dff_B_7HnIj5zW7_2),.clk(gclk));
	jdff dff_B_hQK9vWSi7_2(.din(w_dff_B_7HnIj5zW7_2),.dout(w_dff_B_hQK9vWSi7_2),.clk(gclk));
	jdff dff_B_AxdmzWHQ1_2(.din(w_dff_B_hQK9vWSi7_2),.dout(w_dff_B_AxdmzWHQ1_2),.clk(gclk));
	jdff dff_B_iCsp48My5_2(.din(n880),.dout(w_dff_B_iCsp48My5_2),.clk(gclk));
	jdff dff_B_HA8qc1Lm5_2(.din(w_dff_B_iCsp48My5_2),.dout(w_dff_B_HA8qc1Lm5_2),.clk(gclk));
	jdff dff_B_P00s8lh91_2(.din(w_dff_B_HA8qc1Lm5_2),.dout(w_dff_B_P00s8lh91_2),.clk(gclk));
	jdff dff_B_dwgyX0h69_1(.din(n868),.dout(w_dff_B_dwgyX0h69_1),.clk(gclk));
	jdff dff_B_B7jVbXwV8_1(.din(w_dff_B_dwgyX0h69_1),.dout(w_dff_B_B7jVbXwV8_1),.clk(gclk));
	jdff dff_B_MJ3UurQN6_2(.din(n771),.dout(w_dff_B_MJ3UurQN6_2),.clk(gclk));
	jdff dff_B_OZfCZq0z4_2(.din(w_dff_B_MJ3UurQN6_2),.dout(w_dff_B_OZfCZq0z4_2),.clk(gclk));
	jdff dff_B_x2wZXyLI6_2(.din(w_dff_B_OZfCZq0z4_2),.dout(w_dff_B_x2wZXyLI6_2),.clk(gclk));
	jdff dff_B_CPt8EioO4_0(.din(n776),.dout(w_dff_B_CPt8EioO4_0),.clk(gclk));
	jdff dff_A_WpIMPUUK4_0(.dout(w_n676_0[0]),.din(w_dff_A_WpIMPUUK4_0),.clk(gclk));
	jdff dff_A_ddDRVV2g5_0(.dout(w_dff_A_WpIMPUUK4_0),.din(w_dff_A_ddDRVV2g5_0),.clk(gclk));
	jdff dff_A_Cvr6BZlL8_1(.dout(w_n676_0[1]),.din(w_dff_A_Cvr6BZlL8_1),.clk(gclk));
	jdff dff_A_u7HtRnIt1_1(.dout(w_dff_A_Cvr6BZlL8_1),.din(w_dff_A_u7HtRnIt1_1),.clk(gclk));
	jdff dff_B_rnOokL9a0_1(.din(n1812),.dout(w_dff_B_rnOokL9a0_1),.clk(gclk));
	jdff dff_B_eemYFfZE1_1(.din(n1799),.dout(w_dff_B_eemYFfZE1_1),.clk(gclk));
	jdff dff_B_qoKI2Mw54_1(.din(w_dff_B_eemYFfZE1_1),.dout(w_dff_B_qoKI2Mw54_1),.clk(gclk));
	jdff dff_B_fekuKRv69_2(.din(n1798),.dout(w_dff_B_fekuKRv69_2),.clk(gclk));
	jdff dff_B_6o46UZoJ2_2(.din(w_dff_B_fekuKRv69_2),.dout(w_dff_B_6o46UZoJ2_2),.clk(gclk));
	jdff dff_B_ScWcUdbH1_2(.din(w_dff_B_6o46UZoJ2_2),.dout(w_dff_B_ScWcUdbH1_2),.clk(gclk));
	jdff dff_B_Fza23mTq3_2(.din(w_dff_B_ScWcUdbH1_2),.dout(w_dff_B_Fza23mTq3_2),.clk(gclk));
	jdff dff_B_FKB9wtSE6_2(.din(w_dff_B_Fza23mTq3_2),.dout(w_dff_B_FKB9wtSE6_2),.clk(gclk));
	jdff dff_B_pwQQ3Vxg0_2(.din(w_dff_B_FKB9wtSE6_2),.dout(w_dff_B_pwQQ3Vxg0_2),.clk(gclk));
	jdff dff_B_OSw2XQzE6_2(.din(w_dff_B_pwQQ3Vxg0_2),.dout(w_dff_B_OSw2XQzE6_2),.clk(gclk));
	jdff dff_B_8h2JOS4D1_2(.din(w_dff_B_OSw2XQzE6_2),.dout(w_dff_B_8h2JOS4D1_2),.clk(gclk));
	jdff dff_B_iSK38hw75_2(.din(w_dff_B_8h2JOS4D1_2),.dout(w_dff_B_iSK38hw75_2),.clk(gclk));
	jdff dff_B_SuNKY6o98_2(.din(w_dff_B_iSK38hw75_2),.dout(w_dff_B_SuNKY6o98_2),.clk(gclk));
	jdff dff_B_WfFvJ3ds6_2(.din(w_dff_B_SuNKY6o98_2),.dout(w_dff_B_WfFvJ3ds6_2),.clk(gclk));
	jdff dff_B_YYfaUxtK7_2(.din(w_dff_B_WfFvJ3ds6_2),.dout(w_dff_B_YYfaUxtK7_2),.clk(gclk));
	jdff dff_B_dYkhZAQ05_2(.din(w_dff_B_YYfaUxtK7_2),.dout(w_dff_B_dYkhZAQ05_2),.clk(gclk));
	jdff dff_B_UhWBAowR8_2(.din(w_dff_B_dYkhZAQ05_2),.dout(w_dff_B_UhWBAowR8_2),.clk(gclk));
	jdff dff_B_3ogD9THR8_2(.din(w_dff_B_UhWBAowR8_2),.dout(w_dff_B_3ogD9THR8_2),.clk(gclk));
	jdff dff_B_1iM6xSUK3_2(.din(w_dff_B_3ogD9THR8_2),.dout(w_dff_B_1iM6xSUK3_2),.clk(gclk));
	jdff dff_B_LbN90txj0_2(.din(w_dff_B_1iM6xSUK3_2),.dout(w_dff_B_LbN90txj0_2),.clk(gclk));
	jdff dff_B_HHx7ipqQ8_2(.din(w_dff_B_LbN90txj0_2),.dout(w_dff_B_HHx7ipqQ8_2),.clk(gclk));
	jdff dff_B_V540786e0_2(.din(w_dff_B_HHx7ipqQ8_2),.dout(w_dff_B_V540786e0_2),.clk(gclk));
	jdff dff_B_ylMcfni99_2(.din(w_dff_B_V540786e0_2),.dout(w_dff_B_ylMcfni99_2),.clk(gclk));
	jdff dff_B_cfL4g4H03_2(.din(w_dff_B_ylMcfni99_2),.dout(w_dff_B_cfL4g4H03_2),.clk(gclk));
	jdff dff_B_waiXJdWJ2_2(.din(w_dff_B_cfL4g4H03_2),.dout(w_dff_B_waiXJdWJ2_2),.clk(gclk));
	jdff dff_B_VjQ6fMhN5_2(.din(w_dff_B_waiXJdWJ2_2),.dout(w_dff_B_VjQ6fMhN5_2),.clk(gclk));
	jdff dff_B_tpLpNfts2_2(.din(w_dff_B_VjQ6fMhN5_2),.dout(w_dff_B_tpLpNfts2_2),.clk(gclk));
	jdff dff_B_Et7EwVPd9_2(.din(w_dff_B_tpLpNfts2_2),.dout(w_dff_B_Et7EwVPd9_2),.clk(gclk));
	jdff dff_B_UJCaMQ2l8_2(.din(w_dff_B_Et7EwVPd9_2),.dout(w_dff_B_UJCaMQ2l8_2),.clk(gclk));
	jdff dff_B_54nb5RJS4_2(.din(w_dff_B_UJCaMQ2l8_2),.dout(w_dff_B_54nb5RJS4_2),.clk(gclk));
	jdff dff_B_ncsG6zO35_2(.din(w_dff_B_54nb5RJS4_2),.dout(w_dff_B_ncsG6zO35_2),.clk(gclk));
	jdff dff_B_AgJoGb7q0_2(.din(w_dff_B_ncsG6zO35_2),.dout(w_dff_B_AgJoGb7q0_2),.clk(gclk));
	jdff dff_B_Dheq6hcl7_2(.din(w_dff_B_AgJoGb7q0_2),.dout(w_dff_B_Dheq6hcl7_2),.clk(gclk));
	jdff dff_B_EC1RA1He8_2(.din(w_dff_B_Dheq6hcl7_2),.dout(w_dff_B_EC1RA1He8_2),.clk(gclk));
	jdff dff_B_i06ei0xs0_2(.din(w_dff_B_EC1RA1He8_2),.dout(w_dff_B_i06ei0xs0_2),.clk(gclk));
	jdff dff_B_32qNexT32_2(.din(w_dff_B_i06ei0xs0_2),.dout(w_dff_B_32qNexT32_2),.clk(gclk));
	jdff dff_B_A61xT71d8_2(.din(w_dff_B_32qNexT32_2),.dout(w_dff_B_A61xT71d8_2),.clk(gclk));
	jdff dff_B_iepEY6QA4_2(.din(w_dff_B_A61xT71d8_2),.dout(w_dff_B_iepEY6QA4_2),.clk(gclk));
	jdff dff_B_bfsOVy8W7_2(.din(w_dff_B_iepEY6QA4_2),.dout(w_dff_B_bfsOVy8W7_2),.clk(gclk));
	jdff dff_B_F1O6xQX38_2(.din(w_dff_B_bfsOVy8W7_2),.dout(w_dff_B_F1O6xQX38_2),.clk(gclk));
	jdff dff_B_XafBI5KU8_2(.din(w_dff_B_F1O6xQX38_2),.dout(w_dff_B_XafBI5KU8_2),.clk(gclk));
	jdff dff_B_V5ZrDsEz6_2(.din(w_dff_B_XafBI5KU8_2),.dout(w_dff_B_V5ZrDsEz6_2),.clk(gclk));
	jdff dff_B_fygMFRAS3_2(.din(w_dff_B_V5ZrDsEz6_2),.dout(w_dff_B_fygMFRAS3_2),.clk(gclk));
	jdff dff_B_BoMWUDut6_2(.din(w_dff_B_fygMFRAS3_2),.dout(w_dff_B_BoMWUDut6_2),.clk(gclk));
	jdff dff_B_VskeT8Gn3_2(.din(w_dff_B_BoMWUDut6_2),.dout(w_dff_B_VskeT8Gn3_2),.clk(gclk));
	jdff dff_B_mfIE8pPi6_2(.din(w_dff_B_VskeT8Gn3_2),.dout(w_dff_B_mfIE8pPi6_2),.clk(gclk));
	jdff dff_B_oQAX6XgK2_2(.din(w_dff_B_mfIE8pPi6_2),.dout(w_dff_B_oQAX6XgK2_2),.clk(gclk));
	jdff dff_B_1tYcAu7d7_2(.din(w_dff_B_oQAX6XgK2_2),.dout(w_dff_B_1tYcAu7d7_2),.clk(gclk));
	jdff dff_B_iS8DQAJU4_2(.din(w_dff_B_1tYcAu7d7_2),.dout(w_dff_B_iS8DQAJU4_2),.clk(gclk));
	jdff dff_B_LD8x03BM6_2(.din(w_dff_B_iS8DQAJU4_2),.dout(w_dff_B_LD8x03BM6_2),.clk(gclk));
	jdff dff_B_eiY4043F5_2(.din(w_dff_B_LD8x03BM6_2),.dout(w_dff_B_eiY4043F5_2),.clk(gclk));
	jdff dff_B_yqGLUhTl0_2(.din(w_dff_B_eiY4043F5_2),.dout(w_dff_B_yqGLUhTl0_2),.clk(gclk));
	jdff dff_B_XsNfQcA90_2(.din(w_dff_B_yqGLUhTl0_2),.dout(w_dff_B_XsNfQcA90_2),.clk(gclk));
	jdff dff_B_kHmAAaLS5_2(.din(w_dff_B_XsNfQcA90_2),.dout(w_dff_B_kHmAAaLS5_2),.clk(gclk));
	jdff dff_B_GzkyVSpP2_2(.din(w_dff_B_kHmAAaLS5_2),.dout(w_dff_B_GzkyVSpP2_2),.clk(gclk));
	jdff dff_B_qbkifT6e7_2(.din(w_dff_B_GzkyVSpP2_2),.dout(w_dff_B_qbkifT6e7_2),.clk(gclk));
	jdff dff_B_wHex4ErG5_2(.din(n1797),.dout(w_dff_B_wHex4ErG5_2),.clk(gclk));
	jdff dff_B_NRorvn3D1_2(.din(w_dff_B_wHex4ErG5_2),.dout(w_dff_B_NRorvn3D1_2),.clk(gclk));
	jdff dff_B_dnrhKfRz2_2(.din(w_dff_B_NRorvn3D1_2),.dout(w_dff_B_dnrhKfRz2_2),.clk(gclk));
	jdff dff_B_iKSGlt2k2_2(.din(w_dff_B_dnrhKfRz2_2),.dout(w_dff_B_iKSGlt2k2_2),.clk(gclk));
	jdff dff_B_6KZtI9BN5_2(.din(w_dff_B_iKSGlt2k2_2),.dout(w_dff_B_6KZtI9BN5_2),.clk(gclk));
	jdff dff_B_BxohSfVY3_2(.din(w_dff_B_6KZtI9BN5_2),.dout(w_dff_B_BxohSfVY3_2),.clk(gclk));
	jdff dff_B_hUDzoFWI9_2(.din(w_dff_B_BxohSfVY3_2),.dout(w_dff_B_hUDzoFWI9_2),.clk(gclk));
	jdff dff_B_ISFZ6qAj6_2(.din(w_dff_B_hUDzoFWI9_2),.dout(w_dff_B_ISFZ6qAj6_2),.clk(gclk));
	jdff dff_B_bZoKpMmg6_2(.din(w_dff_B_ISFZ6qAj6_2),.dout(w_dff_B_bZoKpMmg6_2),.clk(gclk));
	jdff dff_B_ikxFmEcE1_2(.din(w_dff_B_bZoKpMmg6_2),.dout(w_dff_B_ikxFmEcE1_2),.clk(gclk));
	jdff dff_B_FcWayhaS9_2(.din(w_dff_B_ikxFmEcE1_2),.dout(w_dff_B_FcWayhaS9_2),.clk(gclk));
	jdff dff_B_vQ8lOx3G1_2(.din(w_dff_B_FcWayhaS9_2),.dout(w_dff_B_vQ8lOx3G1_2),.clk(gclk));
	jdff dff_B_0dp8mov36_2(.din(w_dff_B_vQ8lOx3G1_2),.dout(w_dff_B_0dp8mov36_2),.clk(gclk));
	jdff dff_B_sFdmXqkX9_2(.din(w_dff_B_0dp8mov36_2),.dout(w_dff_B_sFdmXqkX9_2),.clk(gclk));
	jdff dff_B_WF8y5fMJ1_2(.din(w_dff_B_sFdmXqkX9_2),.dout(w_dff_B_WF8y5fMJ1_2),.clk(gclk));
	jdff dff_B_qq8b4wp45_2(.din(w_dff_B_WF8y5fMJ1_2),.dout(w_dff_B_qq8b4wp45_2),.clk(gclk));
	jdff dff_B_KQBaWEgq6_2(.din(w_dff_B_qq8b4wp45_2),.dout(w_dff_B_KQBaWEgq6_2),.clk(gclk));
	jdff dff_B_euyVptgE5_2(.din(w_dff_B_KQBaWEgq6_2),.dout(w_dff_B_euyVptgE5_2),.clk(gclk));
	jdff dff_B_7pfLpn5v1_2(.din(w_dff_B_euyVptgE5_2),.dout(w_dff_B_7pfLpn5v1_2),.clk(gclk));
	jdff dff_B_fOGfCDcD5_2(.din(w_dff_B_7pfLpn5v1_2),.dout(w_dff_B_fOGfCDcD5_2),.clk(gclk));
	jdff dff_B_8hIqXpWi8_2(.din(w_dff_B_fOGfCDcD5_2),.dout(w_dff_B_8hIqXpWi8_2),.clk(gclk));
	jdff dff_B_9P8HEvje1_2(.din(w_dff_B_8hIqXpWi8_2),.dout(w_dff_B_9P8HEvje1_2),.clk(gclk));
	jdff dff_B_HJ92Qrpr8_2(.din(w_dff_B_9P8HEvje1_2),.dout(w_dff_B_HJ92Qrpr8_2),.clk(gclk));
	jdff dff_B_e6rj65kD3_2(.din(w_dff_B_HJ92Qrpr8_2),.dout(w_dff_B_e6rj65kD3_2),.clk(gclk));
	jdff dff_B_4TqLvPoB2_2(.din(w_dff_B_e6rj65kD3_2),.dout(w_dff_B_4TqLvPoB2_2),.clk(gclk));
	jdff dff_B_mXqIyH7B0_2(.din(w_dff_B_4TqLvPoB2_2),.dout(w_dff_B_mXqIyH7B0_2),.clk(gclk));
	jdff dff_B_rCTg4omV4_2(.din(w_dff_B_mXqIyH7B0_2),.dout(w_dff_B_rCTg4omV4_2),.clk(gclk));
	jdff dff_B_6CKiChEE0_2(.din(w_dff_B_rCTg4omV4_2),.dout(w_dff_B_6CKiChEE0_2),.clk(gclk));
	jdff dff_B_J3iEX8oP7_2(.din(w_dff_B_6CKiChEE0_2),.dout(w_dff_B_J3iEX8oP7_2),.clk(gclk));
	jdff dff_B_x11pYp299_2(.din(w_dff_B_J3iEX8oP7_2),.dout(w_dff_B_x11pYp299_2),.clk(gclk));
	jdff dff_B_fqSX8xtR7_2(.din(w_dff_B_x11pYp299_2),.dout(w_dff_B_fqSX8xtR7_2),.clk(gclk));
	jdff dff_B_aoLxrmVu7_2(.din(w_dff_B_fqSX8xtR7_2),.dout(w_dff_B_aoLxrmVu7_2),.clk(gclk));
	jdff dff_B_l2MwQBq36_2(.din(w_dff_B_aoLxrmVu7_2),.dout(w_dff_B_l2MwQBq36_2),.clk(gclk));
	jdff dff_B_yWm41cbh2_2(.din(w_dff_B_l2MwQBq36_2),.dout(w_dff_B_yWm41cbh2_2),.clk(gclk));
	jdff dff_B_4ft1bbLm8_2(.din(w_dff_B_yWm41cbh2_2),.dout(w_dff_B_4ft1bbLm8_2),.clk(gclk));
	jdff dff_B_SlnWQCht9_2(.din(w_dff_B_4ft1bbLm8_2),.dout(w_dff_B_SlnWQCht9_2),.clk(gclk));
	jdff dff_B_aMCSR9bf3_2(.din(w_dff_B_SlnWQCht9_2),.dout(w_dff_B_aMCSR9bf3_2),.clk(gclk));
	jdff dff_B_8GYIJnRQ1_2(.din(w_dff_B_aMCSR9bf3_2),.dout(w_dff_B_8GYIJnRQ1_2),.clk(gclk));
	jdff dff_B_TJeub2rC8_2(.din(w_dff_B_8GYIJnRQ1_2),.dout(w_dff_B_TJeub2rC8_2),.clk(gclk));
	jdff dff_B_LlKDU5qL8_2(.din(w_dff_B_TJeub2rC8_2),.dout(w_dff_B_LlKDU5qL8_2),.clk(gclk));
	jdff dff_B_3EcdPy3h2_2(.din(w_dff_B_LlKDU5qL8_2),.dout(w_dff_B_3EcdPy3h2_2),.clk(gclk));
	jdff dff_B_2MbxBxlc8_2(.din(w_dff_B_3EcdPy3h2_2),.dout(w_dff_B_2MbxBxlc8_2),.clk(gclk));
	jdff dff_B_47rlAOQB2_2(.din(w_dff_B_2MbxBxlc8_2),.dout(w_dff_B_47rlAOQB2_2),.clk(gclk));
	jdff dff_B_oG65F0kM0_2(.din(w_dff_B_47rlAOQB2_2),.dout(w_dff_B_oG65F0kM0_2),.clk(gclk));
	jdff dff_B_PydkgQ309_2(.din(w_dff_B_oG65F0kM0_2),.dout(w_dff_B_PydkgQ309_2),.clk(gclk));
	jdff dff_B_R0FdWsCi9_2(.din(w_dff_B_PydkgQ309_2),.dout(w_dff_B_R0FdWsCi9_2),.clk(gclk));
	jdff dff_B_PPUprleU2_2(.din(w_dff_B_R0FdWsCi9_2),.dout(w_dff_B_PPUprleU2_2),.clk(gclk));
	jdff dff_B_wCvOxZcE8_2(.din(w_dff_B_PPUprleU2_2),.dout(w_dff_B_wCvOxZcE8_2),.clk(gclk));
	jdff dff_B_qlLGs09n3_2(.din(w_dff_B_wCvOxZcE8_2),.dout(w_dff_B_qlLGs09n3_2),.clk(gclk));
	jdff dff_B_J06WYYku7_2(.din(w_dff_B_qlLGs09n3_2),.dout(w_dff_B_J06WYYku7_2),.clk(gclk));
	jdff dff_B_LYMiaIjV0_2(.din(w_dff_B_J06WYYku7_2),.dout(w_dff_B_LYMiaIjV0_2),.clk(gclk));
	jdff dff_B_3BcFTCck0_2(.din(w_dff_B_LYMiaIjV0_2),.dout(w_dff_B_3BcFTCck0_2),.clk(gclk));
	jdff dff_B_24wYAHYp0_2(.din(w_dff_B_3BcFTCck0_2),.dout(w_dff_B_24wYAHYp0_2),.clk(gclk));
	jdff dff_B_w5zeJbcK1_2(.din(w_dff_B_24wYAHYp0_2),.dout(w_dff_B_w5zeJbcK1_2),.clk(gclk));
	jdff dff_B_h5KCZ1I58_2(.din(w_dff_B_w5zeJbcK1_2),.dout(w_dff_B_h5KCZ1I58_2),.clk(gclk));
	jdff dff_A_AC3zetFj0_1(.dout(w_n1796_0[1]),.din(w_dff_A_AC3zetFj0_1),.clk(gclk));
	jdff dff_B_85yW5gdO3_1(.din(n1794),.dout(w_dff_B_85yW5gdO3_1),.clk(gclk));
	jdff dff_B_8WF4KYqn5_2(.din(n1772),.dout(w_dff_B_8WF4KYqn5_2),.clk(gclk));
	jdff dff_B_Jqn8uaQ92_2(.din(w_dff_B_8WF4KYqn5_2),.dout(w_dff_B_Jqn8uaQ92_2),.clk(gclk));
	jdff dff_B_jy7C6HWf9_2(.din(w_dff_B_Jqn8uaQ92_2),.dout(w_dff_B_jy7C6HWf9_2),.clk(gclk));
	jdff dff_B_Cy9GJQgW8_2(.din(w_dff_B_jy7C6HWf9_2),.dout(w_dff_B_Cy9GJQgW8_2),.clk(gclk));
	jdff dff_B_CCiXw2dm0_2(.din(w_dff_B_Cy9GJQgW8_2),.dout(w_dff_B_CCiXw2dm0_2),.clk(gclk));
	jdff dff_B_QMlT8fwp8_2(.din(w_dff_B_CCiXw2dm0_2),.dout(w_dff_B_QMlT8fwp8_2),.clk(gclk));
	jdff dff_B_UUOvCZ546_2(.din(w_dff_B_QMlT8fwp8_2),.dout(w_dff_B_UUOvCZ546_2),.clk(gclk));
	jdff dff_B_uDvz2kqa7_2(.din(w_dff_B_UUOvCZ546_2),.dout(w_dff_B_uDvz2kqa7_2),.clk(gclk));
	jdff dff_B_SsU40btC3_2(.din(w_dff_B_uDvz2kqa7_2),.dout(w_dff_B_SsU40btC3_2),.clk(gclk));
	jdff dff_B_a9aTANtB6_2(.din(w_dff_B_SsU40btC3_2),.dout(w_dff_B_a9aTANtB6_2),.clk(gclk));
	jdff dff_B_vcyrLHtu7_2(.din(w_dff_B_a9aTANtB6_2),.dout(w_dff_B_vcyrLHtu7_2),.clk(gclk));
	jdff dff_B_h5Efwqro5_2(.din(w_dff_B_vcyrLHtu7_2),.dout(w_dff_B_h5Efwqro5_2),.clk(gclk));
	jdff dff_B_orAWzWoQ9_2(.din(w_dff_B_h5Efwqro5_2),.dout(w_dff_B_orAWzWoQ9_2),.clk(gclk));
	jdff dff_B_CRQ6lrv31_2(.din(w_dff_B_orAWzWoQ9_2),.dout(w_dff_B_CRQ6lrv31_2),.clk(gclk));
	jdff dff_B_cDd7MEgJ8_2(.din(w_dff_B_CRQ6lrv31_2),.dout(w_dff_B_cDd7MEgJ8_2),.clk(gclk));
	jdff dff_B_3HYPkTbX3_2(.din(w_dff_B_cDd7MEgJ8_2),.dout(w_dff_B_3HYPkTbX3_2),.clk(gclk));
	jdff dff_B_BwZAt3Ko7_2(.din(w_dff_B_3HYPkTbX3_2),.dout(w_dff_B_BwZAt3Ko7_2),.clk(gclk));
	jdff dff_B_ufmYqBUq7_2(.din(w_dff_B_BwZAt3Ko7_2),.dout(w_dff_B_ufmYqBUq7_2),.clk(gclk));
	jdff dff_B_71L3SUDj8_2(.din(w_dff_B_ufmYqBUq7_2),.dout(w_dff_B_71L3SUDj8_2),.clk(gclk));
	jdff dff_B_iAicqo8d6_2(.din(w_dff_B_71L3SUDj8_2),.dout(w_dff_B_iAicqo8d6_2),.clk(gclk));
	jdff dff_B_AM2GkTIl7_2(.din(w_dff_B_iAicqo8d6_2),.dout(w_dff_B_AM2GkTIl7_2),.clk(gclk));
	jdff dff_B_zo6ENjUE4_2(.din(w_dff_B_AM2GkTIl7_2),.dout(w_dff_B_zo6ENjUE4_2),.clk(gclk));
	jdff dff_B_PD0ftZX28_2(.din(w_dff_B_zo6ENjUE4_2),.dout(w_dff_B_PD0ftZX28_2),.clk(gclk));
	jdff dff_B_AUJz5OWt4_2(.din(w_dff_B_PD0ftZX28_2),.dout(w_dff_B_AUJz5OWt4_2),.clk(gclk));
	jdff dff_B_VTBdWyW88_2(.din(w_dff_B_AUJz5OWt4_2),.dout(w_dff_B_VTBdWyW88_2),.clk(gclk));
	jdff dff_B_nMBamYQy4_2(.din(w_dff_B_VTBdWyW88_2),.dout(w_dff_B_nMBamYQy4_2),.clk(gclk));
	jdff dff_B_9CqUlWIl8_2(.din(w_dff_B_nMBamYQy4_2),.dout(w_dff_B_9CqUlWIl8_2),.clk(gclk));
	jdff dff_B_FM4MBQ361_2(.din(w_dff_B_9CqUlWIl8_2),.dout(w_dff_B_FM4MBQ361_2),.clk(gclk));
	jdff dff_B_QoMGX0Ri1_2(.din(w_dff_B_FM4MBQ361_2),.dout(w_dff_B_QoMGX0Ri1_2),.clk(gclk));
	jdff dff_B_OJdxKCF99_2(.din(w_dff_B_QoMGX0Ri1_2),.dout(w_dff_B_OJdxKCF99_2),.clk(gclk));
	jdff dff_B_wS5SBU8a9_2(.din(w_dff_B_OJdxKCF99_2),.dout(w_dff_B_wS5SBU8a9_2),.clk(gclk));
	jdff dff_B_Bs5Fozd86_2(.din(w_dff_B_wS5SBU8a9_2),.dout(w_dff_B_Bs5Fozd86_2),.clk(gclk));
	jdff dff_B_Gn2uyNUh3_2(.din(w_dff_B_Bs5Fozd86_2),.dout(w_dff_B_Gn2uyNUh3_2),.clk(gclk));
	jdff dff_B_VQ9xYquK1_2(.din(w_dff_B_Gn2uyNUh3_2),.dout(w_dff_B_VQ9xYquK1_2),.clk(gclk));
	jdff dff_B_lPksMeCS9_2(.din(w_dff_B_VQ9xYquK1_2),.dout(w_dff_B_lPksMeCS9_2),.clk(gclk));
	jdff dff_B_MbFSliPR3_2(.din(w_dff_B_lPksMeCS9_2),.dout(w_dff_B_MbFSliPR3_2),.clk(gclk));
	jdff dff_B_yTXCb2XC6_2(.din(w_dff_B_MbFSliPR3_2),.dout(w_dff_B_yTXCb2XC6_2),.clk(gclk));
	jdff dff_B_3ln4MD2j3_2(.din(w_dff_B_yTXCb2XC6_2),.dout(w_dff_B_3ln4MD2j3_2),.clk(gclk));
	jdff dff_B_57X8Wt5L5_2(.din(w_dff_B_3ln4MD2j3_2),.dout(w_dff_B_57X8Wt5L5_2),.clk(gclk));
	jdff dff_B_TBi551Nz5_2(.din(w_dff_B_57X8Wt5L5_2),.dout(w_dff_B_TBi551Nz5_2),.clk(gclk));
	jdff dff_B_lHpg4irN2_2(.din(w_dff_B_TBi551Nz5_2),.dout(w_dff_B_lHpg4irN2_2),.clk(gclk));
	jdff dff_B_Eg0KSJP98_2(.din(w_dff_B_lHpg4irN2_2),.dout(w_dff_B_Eg0KSJP98_2),.clk(gclk));
	jdff dff_B_2Jy3gg3s6_2(.din(w_dff_B_Eg0KSJP98_2),.dout(w_dff_B_2Jy3gg3s6_2),.clk(gclk));
	jdff dff_B_o7E4ISy59_2(.din(w_dff_B_2Jy3gg3s6_2),.dout(w_dff_B_o7E4ISy59_2),.clk(gclk));
	jdff dff_B_ltad0Hjn0_2(.din(w_dff_B_o7E4ISy59_2),.dout(w_dff_B_ltad0Hjn0_2),.clk(gclk));
	jdff dff_B_uJO1sXxd1_2(.din(w_dff_B_ltad0Hjn0_2),.dout(w_dff_B_uJO1sXxd1_2),.clk(gclk));
	jdff dff_B_T5uxMaiV8_2(.din(w_dff_B_uJO1sXxd1_2),.dout(w_dff_B_T5uxMaiV8_2),.clk(gclk));
	jdff dff_B_033E9Cvb2_2(.din(w_dff_B_T5uxMaiV8_2),.dout(w_dff_B_033E9Cvb2_2),.clk(gclk));
	jdff dff_B_OHakaALJ9_2(.din(w_dff_B_033E9Cvb2_2),.dout(w_dff_B_OHakaALJ9_2),.clk(gclk));
	jdff dff_B_8vHTzRsX1_2(.din(w_dff_B_OHakaALJ9_2),.dout(w_dff_B_8vHTzRsX1_2),.clk(gclk));
	jdff dff_B_gRltySca3_2(.din(w_dff_B_8vHTzRsX1_2),.dout(w_dff_B_gRltySca3_2),.clk(gclk));
	jdff dff_B_2CXTIugB1_2(.din(w_dff_B_gRltySca3_2),.dout(w_dff_B_2CXTIugB1_2),.clk(gclk));
	jdff dff_B_HQF7bk0e2_1(.din(n1778),.dout(w_dff_B_HQF7bk0e2_1),.clk(gclk));
	jdff dff_B_RPpjFPI81_1(.din(w_dff_B_HQF7bk0e2_1),.dout(w_dff_B_RPpjFPI81_1),.clk(gclk));
	jdff dff_B_z32vzuen8_2(.din(n1777),.dout(w_dff_B_z32vzuen8_2),.clk(gclk));
	jdff dff_B_2TxosvpK4_2(.din(w_dff_B_z32vzuen8_2),.dout(w_dff_B_2TxosvpK4_2),.clk(gclk));
	jdff dff_B_2zP9rxji0_2(.din(w_dff_B_2TxosvpK4_2),.dout(w_dff_B_2zP9rxji0_2),.clk(gclk));
	jdff dff_B_tWO7PmSc9_2(.din(w_dff_B_2zP9rxji0_2),.dout(w_dff_B_tWO7PmSc9_2),.clk(gclk));
	jdff dff_B_WlMbHSGw4_2(.din(w_dff_B_tWO7PmSc9_2),.dout(w_dff_B_WlMbHSGw4_2),.clk(gclk));
	jdff dff_B_FpxiYoBb8_2(.din(w_dff_B_WlMbHSGw4_2),.dout(w_dff_B_FpxiYoBb8_2),.clk(gclk));
	jdff dff_B_Dbvpant06_2(.din(w_dff_B_FpxiYoBb8_2),.dout(w_dff_B_Dbvpant06_2),.clk(gclk));
	jdff dff_B_0FjwZUAB1_2(.din(w_dff_B_Dbvpant06_2),.dout(w_dff_B_0FjwZUAB1_2),.clk(gclk));
	jdff dff_B_2ULonY1o0_2(.din(w_dff_B_0FjwZUAB1_2),.dout(w_dff_B_2ULonY1o0_2),.clk(gclk));
	jdff dff_B_G8sLIlY88_2(.din(w_dff_B_2ULonY1o0_2),.dout(w_dff_B_G8sLIlY88_2),.clk(gclk));
	jdff dff_B_fcjllQOJ1_2(.din(w_dff_B_G8sLIlY88_2),.dout(w_dff_B_fcjllQOJ1_2),.clk(gclk));
	jdff dff_B_yEW0P7HF4_2(.din(w_dff_B_fcjllQOJ1_2),.dout(w_dff_B_yEW0P7HF4_2),.clk(gclk));
	jdff dff_B_s8ylfpqX8_2(.din(w_dff_B_yEW0P7HF4_2),.dout(w_dff_B_s8ylfpqX8_2),.clk(gclk));
	jdff dff_B_MV29CfLk2_2(.din(w_dff_B_s8ylfpqX8_2),.dout(w_dff_B_MV29CfLk2_2),.clk(gclk));
	jdff dff_B_DX3fr6qb6_2(.din(w_dff_B_MV29CfLk2_2),.dout(w_dff_B_DX3fr6qb6_2),.clk(gclk));
	jdff dff_B_tlRlAHoH7_2(.din(w_dff_B_DX3fr6qb6_2),.dout(w_dff_B_tlRlAHoH7_2),.clk(gclk));
	jdff dff_B_9L95tK7M0_2(.din(w_dff_B_tlRlAHoH7_2),.dout(w_dff_B_9L95tK7M0_2),.clk(gclk));
	jdff dff_B_QYeBX5YM1_2(.din(w_dff_B_9L95tK7M0_2),.dout(w_dff_B_QYeBX5YM1_2),.clk(gclk));
	jdff dff_B_TCHWB0M38_2(.din(w_dff_B_QYeBX5YM1_2),.dout(w_dff_B_TCHWB0M38_2),.clk(gclk));
	jdff dff_B_aVZyOHo32_2(.din(w_dff_B_TCHWB0M38_2),.dout(w_dff_B_aVZyOHo32_2),.clk(gclk));
	jdff dff_B_X8OHSapp3_2(.din(w_dff_B_aVZyOHo32_2),.dout(w_dff_B_X8OHSapp3_2),.clk(gclk));
	jdff dff_B_PYYePxEZ2_2(.din(w_dff_B_X8OHSapp3_2),.dout(w_dff_B_PYYePxEZ2_2),.clk(gclk));
	jdff dff_B_0Zw2sFuo4_2(.din(w_dff_B_PYYePxEZ2_2),.dout(w_dff_B_0Zw2sFuo4_2),.clk(gclk));
	jdff dff_B_hzZt9EVf5_2(.din(w_dff_B_0Zw2sFuo4_2),.dout(w_dff_B_hzZt9EVf5_2),.clk(gclk));
	jdff dff_B_JvyXTsTy1_2(.din(w_dff_B_hzZt9EVf5_2),.dout(w_dff_B_JvyXTsTy1_2),.clk(gclk));
	jdff dff_B_5darSBRX8_2(.din(w_dff_B_JvyXTsTy1_2),.dout(w_dff_B_5darSBRX8_2),.clk(gclk));
	jdff dff_B_1GVf5QKc6_2(.din(w_dff_B_5darSBRX8_2),.dout(w_dff_B_1GVf5QKc6_2),.clk(gclk));
	jdff dff_B_5D241waB4_2(.din(w_dff_B_1GVf5QKc6_2),.dout(w_dff_B_5D241waB4_2),.clk(gclk));
	jdff dff_B_cWtCDbYR5_2(.din(w_dff_B_5D241waB4_2),.dout(w_dff_B_cWtCDbYR5_2),.clk(gclk));
	jdff dff_B_veMo1N1j1_2(.din(w_dff_B_cWtCDbYR5_2),.dout(w_dff_B_veMo1N1j1_2),.clk(gclk));
	jdff dff_B_0iGAMoMH3_2(.din(w_dff_B_veMo1N1j1_2),.dout(w_dff_B_0iGAMoMH3_2),.clk(gclk));
	jdff dff_B_OlQFWA1y7_2(.din(w_dff_B_0iGAMoMH3_2),.dout(w_dff_B_OlQFWA1y7_2),.clk(gclk));
	jdff dff_B_dkUO5tex3_2(.din(w_dff_B_OlQFWA1y7_2),.dout(w_dff_B_dkUO5tex3_2),.clk(gclk));
	jdff dff_B_KHPZNq1z4_2(.din(w_dff_B_dkUO5tex3_2),.dout(w_dff_B_KHPZNq1z4_2),.clk(gclk));
	jdff dff_B_uVHk9e7I4_2(.din(w_dff_B_KHPZNq1z4_2),.dout(w_dff_B_uVHk9e7I4_2),.clk(gclk));
	jdff dff_B_FFAQXH8y8_2(.din(w_dff_B_uVHk9e7I4_2),.dout(w_dff_B_FFAQXH8y8_2),.clk(gclk));
	jdff dff_B_HkgoVjKt2_2(.din(w_dff_B_FFAQXH8y8_2),.dout(w_dff_B_HkgoVjKt2_2),.clk(gclk));
	jdff dff_B_MS9o8qbU7_2(.din(w_dff_B_HkgoVjKt2_2),.dout(w_dff_B_MS9o8qbU7_2),.clk(gclk));
	jdff dff_B_rXqxLoeU5_2(.din(w_dff_B_MS9o8qbU7_2),.dout(w_dff_B_rXqxLoeU5_2),.clk(gclk));
	jdff dff_B_KHyzEeXE7_2(.din(w_dff_B_rXqxLoeU5_2),.dout(w_dff_B_KHyzEeXE7_2),.clk(gclk));
	jdff dff_B_k6RKacYf8_2(.din(w_dff_B_KHyzEeXE7_2),.dout(w_dff_B_k6RKacYf8_2),.clk(gclk));
	jdff dff_B_kwa01AcH7_2(.din(w_dff_B_k6RKacYf8_2),.dout(w_dff_B_kwa01AcH7_2),.clk(gclk));
	jdff dff_B_iAwdxS9e9_2(.din(w_dff_B_kwa01AcH7_2),.dout(w_dff_B_iAwdxS9e9_2),.clk(gclk));
	jdff dff_B_rWMhrAY43_2(.din(w_dff_B_iAwdxS9e9_2),.dout(w_dff_B_rWMhrAY43_2),.clk(gclk));
	jdff dff_B_WDx2Oece0_2(.din(w_dff_B_rWMhrAY43_2),.dout(w_dff_B_WDx2Oece0_2),.clk(gclk));
	jdff dff_B_LHhYusnr3_2(.din(w_dff_B_WDx2Oece0_2),.dout(w_dff_B_LHhYusnr3_2),.clk(gclk));
	jdff dff_B_mG0hsKCn9_2(.din(w_dff_B_LHhYusnr3_2),.dout(w_dff_B_mG0hsKCn9_2),.clk(gclk));
	jdff dff_B_1ULdHyqg5_2(.din(w_dff_B_mG0hsKCn9_2),.dout(w_dff_B_1ULdHyqg5_2),.clk(gclk));
	jdff dff_B_shCeCe4X9_2(.din(w_dff_B_1ULdHyqg5_2),.dout(w_dff_B_shCeCe4X9_2),.clk(gclk));
	jdff dff_B_38XHFW1a0_2(.din(n1776),.dout(w_dff_B_38XHFW1a0_2),.clk(gclk));
	jdff dff_B_6l6LmxGh8_2(.din(w_dff_B_38XHFW1a0_2),.dout(w_dff_B_6l6LmxGh8_2),.clk(gclk));
	jdff dff_B_pBxWMLd88_2(.din(w_dff_B_6l6LmxGh8_2),.dout(w_dff_B_pBxWMLd88_2),.clk(gclk));
	jdff dff_B_VXmyVpwX6_2(.din(w_dff_B_pBxWMLd88_2),.dout(w_dff_B_VXmyVpwX6_2),.clk(gclk));
	jdff dff_B_IdiO4bbN6_2(.din(w_dff_B_VXmyVpwX6_2),.dout(w_dff_B_IdiO4bbN6_2),.clk(gclk));
	jdff dff_B_NmtiALd18_2(.din(w_dff_B_IdiO4bbN6_2),.dout(w_dff_B_NmtiALd18_2),.clk(gclk));
	jdff dff_B_ao1mXhxw2_2(.din(w_dff_B_NmtiALd18_2),.dout(w_dff_B_ao1mXhxw2_2),.clk(gclk));
	jdff dff_B_ZbBMZt8j7_2(.din(w_dff_B_ao1mXhxw2_2),.dout(w_dff_B_ZbBMZt8j7_2),.clk(gclk));
	jdff dff_B_kk0Uvfm58_2(.din(w_dff_B_ZbBMZt8j7_2),.dout(w_dff_B_kk0Uvfm58_2),.clk(gclk));
	jdff dff_B_lZPcH5UB8_2(.din(w_dff_B_kk0Uvfm58_2),.dout(w_dff_B_lZPcH5UB8_2),.clk(gclk));
	jdff dff_B_ArcWtZyl0_2(.din(w_dff_B_lZPcH5UB8_2),.dout(w_dff_B_ArcWtZyl0_2),.clk(gclk));
	jdff dff_B_Ei18dZBy1_2(.din(w_dff_B_ArcWtZyl0_2),.dout(w_dff_B_Ei18dZBy1_2),.clk(gclk));
	jdff dff_B_mNppE8HK5_2(.din(w_dff_B_Ei18dZBy1_2),.dout(w_dff_B_mNppE8HK5_2),.clk(gclk));
	jdff dff_B_1cqeLFF82_2(.din(w_dff_B_mNppE8HK5_2),.dout(w_dff_B_1cqeLFF82_2),.clk(gclk));
	jdff dff_B_gjrizHwI6_2(.din(w_dff_B_1cqeLFF82_2),.dout(w_dff_B_gjrizHwI6_2),.clk(gclk));
	jdff dff_B_Nr7qpHFG9_2(.din(w_dff_B_gjrizHwI6_2),.dout(w_dff_B_Nr7qpHFG9_2),.clk(gclk));
	jdff dff_B_Tp75y8Qm0_2(.din(w_dff_B_Nr7qpHFG9_2),.dout(w_dff_B_Tp75y8Qm0_2),.clk(gclk));
	jdff dff_B_uulUz8c12_2(.din(w_dff_B_Tp75y8Qm0_2),.dout(w_dff_B_uulUz8c12_2),.clk(gclk));
	jdff dff_B_xBauWA2G6_2(.din(w_dff_B_uulUz8c12_2),.dout(w_dff_B_xBauWA2G6_2),.clk(gclk));
	jdff dff_B_ueKq4WmA4_2(.din(w_dff_B_xBauWA2G6_2),.dout(w_dff_B_ueKq4WmA4_2),.clk(gclk));
	jdff dff_B_nLC5pjLh4_2(.din(w_dff_B_ueKq4WmA4_2),.dout(w_dff_B_nLC5pjLh4_2),.clk(gclk));
	jdff dff_B_fNwM23435_2(.din(w_dff_B_nLC5pjLh4_2),.dout(w_dff_B_fNwM23435_2),.clk(gclk));
	jdff dff_B_UoJcFxZb4_2(.din(w_dff_B_fNwM23435_2),.dout(w_dff_B_UoJcFxZb4_2),.clk(gclk));
	jdff dff_B_hHUbooTL0_2(.din(w_dff_B_UoJcFxZb4_2),.dout(w_dff_B_hHUbooTL0_2),.clk(gclk));
	jdff dff_B_t6v06zX06_2(.din(w_dff_B_hHUbooTL0_2),.dout(w_dff_B_t6v06zX06_2),.clk(gclk));
	jdff dff_B_m4yMbSoz3_2(.din(w_dff_B_t6v06zX06_2),.dout(w_dff_B_m4yMbSoz3_2),.clk(gclk));
	jdff dff_B_p9bNeZhd7_2(.din(w_dff_B_m4yMbSoz3_2),.dout(w_dff_B_p9bNeZhd7_2),.clk(gclk));
	jdff dff_B_xDLC4G8i6_2(.din(w_dff_B_p9bNeZhd7_2),.dout(w_dff_B_xDLC4G8i6_2),.clk(gclk));
	jdff dff_B_Acwt59K28_2(.din(w_dff_B_xDLC4G8i6_2),.dout(w_dff_B_Acwt59K28_2),.clk(gclk));
	jdff dff_B_QQ75cPNx1_2(.din(w_dff_B_Acwt59K28_2),.dout(w_dff_B_QQ75cPNx1_2),.clk(gclk));
	jdff dff_B_BOTMtTsc3_2(.din(w_dff_B_QQ75cPNx1_2),.dout(w_dff_B_BOTMtTsc3_2),.clk(gclk));
	jdff dff_B_JwATBW8Q0_2(.din(w_dff_B_BOTMtTsc3_2),.dout(w_dff_B_JwATBW8Q0_2),.clk(gclk));
	jdff dff_B_l4CR5KVy8_2(.din(w_dff_B_JwATBW8Q0_2),.dout(w_dff_B_l4CR5KVy8_2),.clk(gclk));
	jdff dff_B_PVYLwQFE2_2(.din(w_dff_B_l4CR5KVy8_2),.dout(w_dff_B_PVYLwQFE2_2),.clk(gclk));
	jdff dff_B_1Epdjbom5_2(.din(w_dff_B_PVYLwQFE2_2),.dout(w_dff_B_1Epdjbom5_2),.clk(gclk));
	jdff dff_B_L93FNHMi3_2(.din(w_dff_B_1Epdjbom5_2),.dout(w_dff_B_L93FNHMi3_2),.clk(gclk));
	jdff dff_B_EZ7VocIB0_2(.din(w_dff_B_L93FNHMi3_2),.dout(w_dff_B_EZ7VocIB0_2),.clk(gclk));
	jdff dff_B_puR35NMM1_2(.din(w_dff_B_EZ7VocIB0_2),.dout(w_dff_B_puR35NMM1_2),.clk(gclk));
	jdff dff_B_5ePNdsAh0_2(.din(w_dff_B_puR35NMM1_2),.dout(w_dff_B_5ePNdsAh0_2),.clk(gclk));
	jdff dff_B_d7n0X0my4_2(.din(w_dff_B_5ePNdsAh0_2),.dout(w_dff_B_d7n0X0my4_2),.clk(gclk));
	jdff dff_B_jWC2VfwL4_2(.din(w_dff_B_d7n0X0my4_2),.dout(w_dff_B_jWC2VfwL4_2),.clk(gclk));
	jdff dff_B_HZj48SdY2_2(.din(w_dff_B_jWC2VfwL4_2),.dout(w_dff_B_HZj48SdY2_2),.clk(gclk));
	jdff dff_B_49podTqW6_2(.din(w_dff_B_HZj48SdY2_2),.dout(w_dff_B_49podTqW6_2),.clk(gclk));
	jdff dff_B_XmgPat7m5_2(.din(w_dff_B_49podTqW6_2),.dout(w_dff_B_XmgPat7m5_2),.clk(gclk));
	jdff dff_B_uokwtuQD7_2(.din(w_dff_B_XmgPat7m5_2),.dout(w_dff_B_uokwtuQD7_2),.clk(gclk));
	jdff dff_B_OsJdbdGz5_2(.din(w_dff_B_uokwtuQD7_2),.dout(w_dff_B_OsJdbdGz5_2),.clk(gclk));
	jdff dff_B_VPkaGOVS6_2(.din(w_dff_B_OsJdbdGz5_2),.dout(w_dff_B_VPkaGOVS6_2),.clk(gclk));
	jdff dff_B_deH8Th2h3_2(.din(w_dff_B_VPkaGOVS6_2),.dout(w_dff_B_deH8Th2h3_2),.clk(gclk));
	jdff dff_B_UGOBmCau4_2(.din(w_dff_B_deH8Th2h3_2),.dout(w_dff_B_UGOBmCau4_2),.clk(gclk));
	jdff dff_B_7d4n6SbI0_2(.din(w_dff_B_UGOBmCau4_2),.dout(w_dff_B_7d4n6SbI0_2),.clk(gclk));
	jdff dff_B_3OSCaDKz1_2(.din(w_dff_B_7d4n6SbI0_2),.dout(w_dff_B_3OSCaDKz1_2),.clk(gclk));
	jdff dff_B_8KA5KVCB4_2(.din(n1775),.dout(w_dff_B_8KA5KVCB4_2),.clk(gclk));
	jdff dff_B_qWUxsDRZ7_1(.din(n1773),.dout(w_dff_B_qWUxsDRZ7_1),.clk(gclk));
	jdff dff_B_xD076iXe6_2(.din(n1744),.dout(w_dff_B_xD076iXe6_2),.clk(gclk));
	jdff dff_B_kyesZ4rs8_2(.din(w_dff_B_xD076iXe6_2),.dout(w_dff_B_kyesZ4rs8_2),.clk(gclk));
	jdff dff_B_oik7KltN4_2(.din(w_dff_B_kyesZ4rs8_2),.dout(w_dff_B_oik7KltN4_2),.clk(gclk));
	jdff dff_B_e5tzgqE57_2(.din(w_dff_B_oik7KltN4_2),.dout(w_dff_B_e5tzgqE57_2),.clk(gclk));
	jdff dff_B_oKcMerhe6_2(.din(w_dff_B_e5tzgqE57_2),.dout(w_dff_B_oKcMerhe6_2),.clk(gclk));
	jdff dff_B_Vryh36YB6_2(.din(w_dff_B_oKcMerhe6_2),.dout(w_dff_B_Vryh36YB6_2),.clk(gclk));
	jdff dff_B_6xBYqasI9_2(.din(w_dff_B_Vryh36YB6_2),.dout(w_dff_B_6xBYqasI9_2),.clk(gclk));
	jdff dff_B_19wc5L0r5_2(.din(w_dff_B_6xBYqasI9_2),.dout(w_dff_B_19wc5L0r5_2),.clk(gclk));
	jdff dff_B_aEX32HKi5_2(.din(w_dff_B_19wc5L0r5_2),.dout(w_dff_B_aEX32HKi5_2),.clk(gclk));
	jdff dff_B_sqvRMQzC6_2(.din(w_dff_B_aEX32HKi5_2),.dout(w_dff_B_sqvRMQzC6_2),.clk(gclk));
	jdff dff_B_RSfjmcyd9_2(.din(w_dff_B_sqvRMQzC6_2),.dout(w_dff_B_RSfjmcyd9_2),.clk(gclk));
	jdff dff_B_gqbnx4fx0_2(.din(w_dff_B_RSfjmcyd9_2),.dout(w_dff_B_gqbnx4fx0_2),.clk(gclk));
	jdff dff_B_qJCpyv0l2_2(.din(w_dff_B_gqbnx4fx0_2),.dout(w_dff_B_qJCpyv0l2_2),.clk(gclk));
	jdff dff_B_M9aDvJwx7_2(.din(w_dff_B_qJCpyv0l2_2),.dout(w_dff_B_M9aDvJwx7_2),.clk(gclk));
	jdff dff_B_Y1ZmAn6a6_2(.din(w_dff_B_M9aDvJwx7_2),.dout(w_dff_B_Y1ZmAn6a6_2),.clk(gclk));
	jdff dff_B_9fo6GBzZ7_2(.din(w_dff_B_Y1ZmAn6a6_2),.dout(w_dff_B_9fo6GBzZ7_2),.clk(gclk));
	jdff dff_B_82v8wYhk2_2(.din(w_dff_B_9fo6GBzZ7_2),.dout(w_dff_B_82v8wYhk2_2),.clk(gclk));
	jdff dff_B_um04Y1dA1_2(.din(w_dff_B_82v8wYhk2_2),.dout(w_dff_B_um04Y1dA1_2),.clk(gclk));
	jdff dff_B_fd7C7USc6_2(.din(w_dff_B_um04Y1dA1_2),.dout(w_dff_B_fd7C7USc6_2),.clk(gclk));
	jdff dff_B_G3UktORU8_2(.din(w_dff_B_fd7C7USc6_2),.dout(w_dff_B_G3UktORU8_2),.clk(gclk));
	jdff dff_B_fH7pNbZu5_2(.din(w_dff_B_G3UktORU8_2),.dout(w_dff_B_fH7pNbZu5_2),.clk(gclk));
	jdff dff_B_WKNN1m8k1_2(.din(w_dff_B_fH7pNbZu5_2),.dout(w_dff_B_WKNN1m8k1_2),.clk(gclk));
	jdff dff_B_p3qWDmPL3_2(.din(w_dff_B_WKNN1m8k1_2),.dout(w_dff_B_p3qWDmPL3_2),.clk(gclk));
	jdff dff_B_lCPAivWe7_2(.din(w_dff_B_p3qWDmPL3_2),.dout(w_dff_B_lCPAivWe7_2),.clk(gclk));
	jdff dff_B_DhRAhByB2_2(.din(w_dff_B_lCPAivWe7_2),.dout(w_dff_B_DhRAhByB2_2),.clk(gclk));
	jdff dff_B_VIdwCA4l9_2(.din(w_dff_B_DhRAhByB2_2),.dout(w_dff_B_VIdwCA4l9_2),.clk(gclk));
	jdff dff_B_6MPY2VgM1_2(.din(w_dff_B_VIdwCA4l9_2),.dout(w_dff_B_6MPY2VgM1_2),.clk(gclk));
	jdff dff_B_zNWNzSBz5_2(.din(w_dff_B_6MPY2VgM1_2),.dout(w_dff_B_zNWNzSBz5_2),.clk(gclk));
	jdff dff_B_j9BTXpGQ8_2(.din(w_dff_B_zNWNzSBz5_2),.dout(w_dff_B_j9BTXpGQ8_2),.clk(gclk));
	jdff dff_B_59sPQ6fC3_2(.din(w_dff_B_j9BTXpGQ8_2),.dout(w_dff_B_59sPQ6fC3_2),.clk(gclk));
	jdff dff_B_GBHLQwtx8_2(.din(w_dff_B_59sPQ6fC3_2),.dout(w_dff_B_GBHLQwtx8_2),.clk(gclk));
	jdff dff_B_InKxkVFR3_2(.din(w_dff_B_GBHLQwtx8_2),.dout(w_dff_B_InKxkVFR3_2),.clk(gclk));
	jdff dff_B_ow5G3P7x5_2(.din(w_dff_B_InKxkVFR3_2),.dout(w_dff_B_ow5G3P7x5_2),.clk(gclk));
	jdff dff_B_XL2a7IEz7_2(.din(w_dff_B_ow5G3P7x5_2),.dout(w_dff_B_XL2a7IEz7_2),.clk(gclk));
	jdff dff_B_NGDDQFOp9_2(.din(w_dff_B_XL2a7IEz7_2),.dout(w_dff_B_NGDDQFOp9_2),.clk(gclk));
	jdff dff_B_sRVDEl1N3_2(.din(w_dff_B_NGDDQFOp9_2),.dout(w_dff_B_sRVDEl1N3_2),.clk(gclk));
	jdff dff_B_xrPVKBRL4_2(.din(w_dff_B_sRVDEl1N3_2),.dout(w_dff_B_xrPVKBRL4_2),.clk(gclk));
	jdff dff_B_qIUimjEC6_2(.din(w_dff_B_xrPVKBRL4_2),.dout(w_dff_B_qIUimjEC6_2),.clk(gclk));
	jdff dff_B_LowstA8A8_2(.din(w_dff_B_qIUimjEC6_2),.dout(w_dff_B_LowstA8A8_2),.clk(gclk));
	jdff dff_B_sC89UURm6_2(.din(w_dff_B_LowstA8A8_2),.dout(w_dff_B_sC89UURm6_2),.clk(gclk));
	jdff dff_B_yoHj2H7U8_2(.din(w_dff_B_sC89UURm6_2),.dout(w_dff_B_yoHj2H7U8_2),.clk(gclk));
	jdff dff_B_adlzWLRy3_2(.din(w_dff_B_yoHj2H7U8_2),.dout(w_dff_B_adlzWLRy3_2),.clk(gclk));
	jdff dff_B_epf9saWp2_2(.din(w_dff_B_adlzWLRy3_2),.dout(w_dff_B_epf9saWp2_2),.clk(gclk));
	jdff dff_B_Weh4jPJS0_2(.din(w_dff_B_epf9saWp2_2),.dout(w_dff_B_Weh4jPJS0_2),.clk(gclk));
	jdff dff_B_gRug1Bad9_2(.din(w_dff_B_Weh4jPJS0_2),.dout(w_dff_B_gRug1Bad9_2),.clk(gclk));
	jdff dff_B_I6IYIYEb0_2(.din(w_dff_B_gRug1Bad9_2),.dout(w_dff_B_I6IYIYEb0_2),.clk(gclk));
	jdff dff_B_DevLermn5_2(.din(w_dff_B_I6IYIYEb0_2),.dout(w_dff_B_DevLermn5_2),.clk(gclk));
	jdff dff_B_12hr5EGl3_2(.din(w_dff_B_DevLermn5_2),.dout(w_dff_B_12hr5EGl3_2),.clk(gclk));
	jdff dff_B_CWGCbJ0w0_1(.din(n1750),.dout(w_dff_B_CWGCbJ0w0_1),.clk(gclk));
	jdff dff_B_d4ZAE1QM3_1(.din(w_dff_B_CWGCbJ0w0_1),.dout(w_dff_B_d4ZAE1QM3_1),.clk(gclk));
	jdff dff_B_faJ9xdeC4_2(.din(n1749),.dout(w_dff_B_faJ9xdeC4_2),.clk(gclk));
	jdff dff_B_nF5ANBtQ5_2(.din(w_dff_B_faJ9xdeC4_2),.dout(w_dff_B_nF5ANBtQ5_2),.clk(gclk));
	jdff dff_B_C0XUzrGO1_2(.din(w_dff_B_nF5ANBtQ5_2),.dout(w_dff_B_C0XUzrGO1_2),.clk(gclk));
	jdff dff_B_yM3dHu371_2(.din(w_dff_B_C0XUzrGO1_2),.dout(w_dff_B_yM3dHu371_2),.clk(gclk));
	jdff dff_B_qsKw82EM9_2(.din(w_dff_B_yM3dHu371_2),.dout(w_dff_B_qsKw82EM9_2),.clk(gclk));
	jdff dff_B_qY83BAly6_2(.din(w_dff_B_qsKw82EM9_2),.dout(w_dff_B_qY83BAly6_2),.clk(gclk));
	jdff dff_B_Jwc7aw7h2_2(.din(w_dff_B_qY83BAly6_2),.dout(w_dff_B_Jwc7aw7h2_2),.clk(gclk));
	jdff dff_B_8t6SukKM3_2(.din(w_dff_B_Jwc7aw7h2_2),.dout(w_dff_B_8t6SukKM3_2),.clk(gclk));
	jdff dff_B_lZXZY2CY6_2(.din(w_dff_B_8t6SukKM3_2),.dout(w_dff_B_lZXZY2CY6_2),.clk(gclk));
	jdff dff_B_E6XZIp867_2(.din(w_dff_B_lZXZY2CY6_2),.dout(w_dff_B_E6XZIp867_2),.clk(gclk));
	jdff dff_B_ivekI5sQ4_2(.din(w_dff_B_E6XZIp867_2),.dout(w_dff_B_ivekI5sQ4_2),.clk(gclk));
	jdff dff_B_cqHO71de8_2(.din(w_dff_B_ivekI5sQ4_2),.dout(w_dff_B_cqHO71de8_2),.clk(gclk));
	jdff dff_B_QD0UR4Vz9_2(.din(w_dff_B_cqHO71de8_2),.dout(w_dff_B_QD0UR4Vz9_2),.clk(gclk));
	jdff dff_B_RV1zZGpt4_2(.din(w_dff_B_QD0UR4Vz9_2),.dout(w_dff_B_RV1zZGpt4_2),.clk(gclk));
	jdff dff_B_s7RlcEsX7_2(.din(w_dff_B_RV1zZGpt4_2),.dout(w_dff_B_s7RlcEsX7_2),.clk(gclk));
	jdff dff_B_J44t7Nwn4_2(.din(w_dff_B_s7RlcEsX7_2),.dout(w_dff_B_J44t7Nwn4_2),.clk(gclk));
	jdff dff_B_Y3jwTgdq1_2(.din(w_dff_B_J44t7Nwn4_2),.dout(w_dff_B_Y3jwTgdq1_2),.clk(gclk));
	jdff dff_B_sbN9BVqF3_2(.din(w_dff_B_Y3jwTgdq1_2),.dout(w_dff_B_sbN9BVqF3_2),.clk(gclk));
	jdff dff_B_hWWuQbSl0_2(.din(w_dff_B_sbN9BVqF3_2),.dout(w_dff_B_hWWuQbSl0_2),.clk(gclk));
	jdff dff_B_AphpyBUy8_2(.din(w_dff_B_hWWuQbSl0_2),.dout(w_dff_B_AphpyBUy8_2),.clk(gclk));
	jdff dff_B_j50asqdf6_2(.din(w_dff_B_AphpyBUy8_2),.dout(w_dff_B_j50asqdf6_2),.clk(gclk));
	jdff dff_B_HjQi7iLm1_2(.din(w_dff_B_j50asqdf6_2),.dout(w_dff_B_HjQi7iLm1_2),.clk(gclk));
	jdff dff_B_FGXlemH91_2(.din(w_dff_B_HjQi7iLm1_2),.dout(w_dff_B_FGXlemH91_2),.clk(gclk));
	jdff dff_B_Eb0oQOHA8_2(.din(w_dff_B_FGXlemH91_2),.dout(w_dff_B_Eb0oQOHA8_2),.clk(gclk));
	jdff dff_B_abzWY0ir1_2(.din(w_dff_B_Eb0oQOHA8_2),.dout(w_dff_B_abzWY0ir1_2),.clk(gclk));
	jdff dff_B_hat5Xztu7_2(.din(w_dff_B_abzWY0ir1_2),.dout(w_dff_B_hat5Xztu7_2),.clk(gclk));
	jdff dff_B_NoUV1BRL3_2(.din(w_dff_B_hat5Xztu7_2),.dout(w_dff_B_NoUV1BRL3_2),.clk(gclk));
	jdff dff_B_W50ncMDH3_2(.din(w_dff_B_NoUV1BRL3_2),.dout(w_dff_B_W50ncMDH3_2),.clk(gclk));
	jdff dff_B_st73XXd01_2(.din(w_dff_B_W50ncMDH3_2),.dout(w_dff_B_st73XXd01_2),.clk(gclk));
	jdff dff_B_36MSZ6Yb8_2(.din(w_dff_B_st73XXd01_2),.dout(w_dff_B_36MSZ6Yb8_2),.clk(gclk));
	jdff dff_B_zVlBygQ15_2(.din(w_dff_B_36MSZ6Yb8_2),.dout(w_dff_B_zVlBygQ15_2),.clk(gclk));
	jdff dff_B_wFXBDUk77_2(.din(w_dff_B_zVlBygQ15_2),.dout(w_dff_B_wFXBDUk77_2),.clk(gclk));
	jdff dff_B_3R4mOfJH5_2(.din(w_dff_B_wFXBDUk77_2),.dout(w_dff_B_3R4mOfJH5_2),.clk(gclk));
	jdff dff_B_wO8axMbp6_2(.din(w_dff_B_3R4mOfJH5_2),.dout(w_dff_B_wO8axMbp6_2),.clk(gclk));
	jdff dff_B_MSlP7h3A3_2(.din(w_dff_B_wO8axMbp6_2),.dout(w_dff_B_MSlP7h3A3_2),.clk(gclk));
	jdff dff_B_m21HxMrG0_2(.din(w_dff_B_MSlP7h3A3_2),.dout(w_dff_B_m21HxMrG0_2),.clk(gclk));
	jdff dff_B_VhroFn5w0_2(.din(w_dff_B_m21HxMrG0_2),.dout(w_dff_B_VhroFn5w0_2),.clk(gclk));
	jdff dff_B_oBLqhJkX1_2(.din(w_dff_B_VhroFn5w0_2),.dout(w_dff_B_oBLqhJkX1_2),.clk(gclk));
	jdff dff_B_HUoWclQQ1_2(.din(w_dff_B_oBLqhJkX1_2),.dout(w_dff_B_HUoWclQQ1_2),.clk(gclk));
	jdff dff_B_rrvRyZfs8_2(.din(w_dff_B_HUoWclQQ1_2),.dout(w_dff_B_rrvRyZfs8_2),.clk(gclk));
	jdff dff_B_cHFib2jT1_2(.din(w_dff_B_rrvRyZfs8_2),.dout(w_dff_B_cHFib2jT1_2),.clk(gclk));
	jdff dff_B_C1kslyPO6_2(.din(w_dff_B_cHFib2jT1_2),.dout(w_dff_B_C1kslyPO6_2),.clk(gclk));
	jdff dff_B_mgDUfXp27_2(.din(w_dff_B_C1kslyPO6_2),.dout(w_dff_B_mgDUfXp27_2),.clk(gclk));
	jdff dff_B_fGsuuLXw7_2(.din(w_dff_B_mgDUfXp27_2),.dout(w_dff_B_fGsuuLXw7_2),.clk(gclk));
	jdff dff_B_chfeBSJ11_2(.din(w_dff_B_fGsuuLXw7_2),.dout(w_dff_B_chfeBSJ11_2),.clk(gclk));
	jdff dff_B_2EAVDkLl7_2(.din(n1748),.dout(w_dff_B_2EAVDkLl7_2),.clk(gclk));
	jdff dff_B_ngLYd4XY5_2(.din(w_dff_B_2EAVDkLl7_2),.dout(w_dff_B_ngLYd4XY5_2),.clk(gclk));
	jdff dff_B_gzg6flQI8_2(.din(w_dff_B_ngLYd4XY5_2),.dout(w_dff_B_gzg6flQI8_2),.clk(gclk));
	jdff dff_B_R4yFSMeE1_2(.din(w_dff_B_gzg6flQI8_2),.dout(w_dff_B_R4yFSMeE1_2),.clk(gclk));
	jdff dff_B_YdBBbARr4_2(.din(w_dff_B_R4yFSMeE1_2),.dout(w_dff_B_YdBBbARr4_2),.clk(gclk));
	jdff dff_B_avlYpuqv7_2(.din(w_dff_B_YdBBbARr4_2),.dout(w_dff_B_avlYpuqv7_2),.clk(gclk));
	jdff dff_B_bGdUGE8j5_2(.din(w_dff_B_avlYpuqv7_2),.dout(w_dff_B_bGdUGE8j5_2),.clk(gclk));
	jdff dff_B_umVXL3Dw4_2(.din(w_dff_B_bGdUGE8j5_2),.dout(w_dff_B_umVXL3Dw4_2),.clk(gclk));
	jdff dff_B_jI5YRURc6_2(.din(w_dff_B_umVXL3Dw4_2),.dout(w_dff_B_jI5YRURc6_2),.clk(gclk));
	jdff dff_B_7XKxpy8r3_2(.din(w_dff_B_jI5YRURc6_2),.dout(w_dff_B_7XKxpy8r3_2),.clk(gclk));
	jdff dff_B_jKJ5sE8T3_2(.din(w_dff_B_7XKxpy8r3_2),.dout(w_dff_B_jKJ5sE8T3_2),.clk(gclk));
	jdff dff_B_Hk7b3xWK1_2(.din(w_dff_B_jKJ5sE8T3_2),.dout(w_dff_B_Hk7b3xWK1_2),.clk(gclk));
	jdff dff_B_ew6PZ2WT2_2(.din(w_dff_B_Hk7b3xWK1_2),.dout(w_dff_B_ew6PZ2WT2_2),.clk(gclk));
	jdff dff_B_4eQudNhd7_2(.din(w_dff_B_ew6PZ2WT2_2),.dout(w_dff_B_4eQudNhd7_2),.clk(gclk));
	jdff dff_B_VrgPTmQO6_2(.din(w_dff_B_4eQudNhd7_2),.dout(w_dff_B_VrgPTmQO6_2),.clk(gclk));
	jdff dff_B_GQEYkhqY1_2(.din(w_dff_B_VrgPTmQO6_2),.dout(w_dff_B_GQEYkhqY1_2),.clk(gclk));
	jdff dff_B_cVhU0I1q0_2(.din(w_dff_B_GQEYkhqY1_2),.dout(w_dff_B_cVhU0I1q0_2),.clk(gclk));
	jdff dff_B_ymzaI4fb8_2(.din(w_dff_B_cVhU0I1q0_2),.dout(w_dff_B_ymzaI4fb8_2),.clk(gclk));
	jdff dff_B_7iL8PC3L6_2(.din(w_dff_B_ymzaI4fb8_2),.dout(w_dff_B_7iL8PC3L6_2),.clk(gclk));
	jdff dff_B_OhBTwph58_2(.din(w_dff_B_7iL8PC3L6_2),.dout(w_dff_B_OhBTwph58_2),.clk(gclk));
	jdff dff_B_MIx31jh04_2(.din(w_dff_B_OhBTwph58_2),.dout(w_dff_B_MIx31jh04_2),.clk(gclk));
	jdff dff_B_9Qko8Pqy1_2(.din(w_dff_B_MIx31jh04_2),.dout(w_dff_B_9Qko8Pqy1_2),.clk(gclk));
	jdff dff_B_IrmeGxQh5_2(.din(w_dff_B_9Qko8Pqy1_2),.dout(w_dff_B_IrmeGxQh5_2),.clk(gclk));
	jdff dff_B_10HN8qt34_2(.din(w_dff_B_IrmeGxQh5_2),.dout(w_dff_B_10HN8qt34_2),.clk(gclk));
	jdff dff_B_FPoNjL1f0_2(.din(w_dff_B_10HN8qt34_2),.dout(w_dff_B_FPoNjL1f0_2),.clk(gclk));
	jdff dff_B_Ql9V8Nh02_2(.din(w_dff_B_FPoNjL1f0_2),.dout(w_dff_B_Ql9V8Nh02_2),.clk(gclk));
	jdff dff_B_eZlUtsJ09_2(.din(w_dff_B_Ql9V8Nh02_2),.dout(w_dff_B_eZlUtsJ09_2),.clk(gclk));
	jdff dff_B_GUQEn7xA6_2(.din(w_dff_B_eZlUtsJ09_2),.dout(w_dff_B_GUQEn7xA6_2),.clk(gclk));
	jdff dff_B_fWE6NGUT7_2(.din(w_dff_B_GUQEn7xA6_2),.dout(w_dff_B_fWE6NGUT7_2),.clk(gclk));
	jdff dff_B_7TruB4oG3_2(.din(w_dff_B_fWE6NGUT7_2),.dout(w_dff_B_7TruB4oG3_2),.clk(gclk));
	jdff dff_B_0kioKlY41_2(.din(w_dff_B_7TruB4oG3_2),.dout(w_dff_B_0kioKlY41_2),.clk(gclk));
	jdff dff_B_tJtqcomJ2_2(.din(w_dff_B_0kioKlY41_2),.dout(w_dff_B_tJtqcomJ2_2),.clk(gclk));
	jdff dff_B_0hdK8N0n6_2(.din(w_dff_B_tJtqcomJ2_2),.dout(w_dff_B_0hdK8N0n6_2),.clk(gclk));
	jdff dff_B_kuez1BPk2_2(.din(w_dff_B_0hdK8N0n6_2),.dout(w_dff_B_kuez1BPk2_2),.clk(gclk));
	jdff dff_B_egoPkZ047_2(.din(w_dff_B_kuez1BPk2_2),.dout(w_dff_B_egoPkZ047_2),.clk(gclk));
	jdff dff_B_e3ktsPK58_2(.din(w_dff_B_egoPkZ047_2),.dout(w_dff_B_e3ktsPK58_2),.clk(gclk));
	jdff dff_B_yGNuGTbC4_2(.din(w_dff_B_e3ktsPK58_2),.dout(w_dff_B_yGNuGTbC4_2),.clk(gclk));
	jdff dff_B_RO0r7OBj8_2(.din(w_dff_B_yGNuGTbC4_2),.dout(w_dff_B_RO0r7OBj8_2),.clk(gclk));
	jdff dff_B_1Z4GYRlm9_2(.din(w_dff_B_RO0r7OBj8_2),.dout(w_dff_B_1Z4GYRlm9_2),.clk(gclk));
	jdff dff_B_apBpyLGa3_2(.din(w_dff_B_1Z4GYRlm9_2),.dout(w_dff_B_apBpyLGa3_2),.clk(gclk));
	jdff dff_B_1Kk16XHi5_2(.din(w_dff_B_apBpyLGa3_2),.dout(w_dff_B_1Kk16XHi5_2),.clk(gclk));
	jdff dff_B_n1TXBwYX3_2(.din(w_dff_B_1Kk16XHi5_2),.dout(w_dff_B_n1TXBwYX3_2),.clk(gclk));
	jdff dff_B_LrNu2tmv7_2(.din(w_dff_B_n1TXBwYX3_2),.dout(w_dff_B_LrNu2tmv7_2),.clk(gclk));
	jdff dff_B_gvhiwkz56_2(.din(w_dff_B_LrNu2tmv7_2),.dout(w_dff_B_gvhiwkz56_2),.clk(gclk));
	jdff dff_B_mJ3gr90N8_2(.din(w_dff_B_gvhiwkz56_2),.dout(w_dff_B_mJ3gr90N8_2),.clk(gclk));
	jdff dff_B_srHe9ezn4_2(.din(w_dff_B_mJ3gr90N8_2),.dout(w_dff_B_srHe9ezn4_2),.clk(gclk));
	jdff dff_B_t3UUnhQ63_2(.din(w_dff_B_srHe9ezn4_2),.dout(w_dff_B_t3UUnhQ63_2),.clk(gclk));
	jdff dff_B_j4DIVSxT5_2(.din(n1747),.dout(w_dff_B_j4DIVSxT5_2),.clk(gclk));
	jdff dff_B_1cUf0YGg3_1(.din(n1745),.dout(w_dff_B_1cUf0YGg3_1),.clk(gclk));
	jdff dff_B_fYLZYovA4_2(.din(n1709),.dout(w_dff_B_fYLZYovA4_2),.clk(gclk));
	jdff dff_B_vSbmGcqz5_2(.din(w_dff_B_fYLZYovA4_2),.dout(w_dff_B_vSbmGcqz5_2),.clk(gclk));
	jdff dff_B_jQbvSLKP1_2(.din(w_dff_B_vSbmGcqz5_2),.dout(w_dff_B_jQbvSLKP1_2),.clk(gclk));
	jdff dff_B_gszgBOQm4_2(.din(w_dff_B_jQbvSLKP1_2),.dout(w_dff_B_gszgBOQm4_2),.clk(gclk));
	jdff dff_B_RuqD6PyM5_2(.din(w_dff_B_gszgBOQm4_2),.dout(w_dff_B_RuqD6PyM5_2),.clk(gclk));
	jdff dff_B_52HjBxyi4_2(.din(w_dff_B_RuqD6PyM5_2),.dout(w_dff_B_52HjBxyi4_2),.clk(gclk));
	jdff dff_B_NRd8nkEE1_2(.din(w_dff_B_52HjBxyi4_2),.dout(w_dff_B_NRd8nkEE1_2),.clk(gclk));
	jdff dff_B_sN5CeOlZ1_2(.din(w_dff_B_NRd8nkEE1_2),.dout(w_dff_B_sN5CeOlZ1_2),.clk(gclk));
	jdff dff_B_PIYKBRiq6_2(.din(w_dff_B_sN5CeOlZ1_2),.dout(w_dff_B_PIYKBRiq6_2),.clk(gclk));
	jdff dff_B_VfWB5LxK4_2(.din(w_dff_B_PIYKBRiq6_2),.dout(w_dff_B_VfWB5LxK4_2),.clk(gclk));
	jdff dff_B_sKybOTp39_2(.din(w_dff_B_VfWB5LxK4_2),.dout(w_dff_B_sKybOTp39_2),.clk(gclk));
	jdff dff_B_ApqATlrs4_2(.din(w_dff_B_sKybOTp39_2),.dout(w_dff_B_ApqATlrs4_2),.clk(gclk));
	jdff dff_B_mr0OaWUT2_2(.din(w_dff_B_ApqATlrs4_2),.dout(w_dff_B_mr0OaWUT2_2),.clk(gclk));
	jdff dff_B_ARTueBT24_2(.din(w_dff_B_mr0OaWUT2_2),.dout(w_dff_B_ARTueBT24_2),.clk(gclk));
	jdff dff_B_6KuKY68J7_2(.din(w_dff_B_ARTueBT24_2),.dout(w_dff_B_6KuKY68J7_2),.clk(gclk));
	jdff dff_B_hk87IMgY3_2(.din(w_dff_B_6KuKY68J7_2),.dout(w_dff_B_hk87IMgY3_2),.clk(gclk));
	jdff dff_B_887I8Jxa2_2(.din(w_dff_B_hk87IMgY3_2),.dout(w_dff_B_887I8Jxa2_2),.clk(gclk));
	jdff dff_B_yZjRqMe42_2(.din(w_dff_B_887I8Jxa2_2),.dout(w_dff_B_yZjRqMe42_2),.clk(gclk));
	jdff dff_B_NM0Y1hWn2_2(.din(w_dff_B_yZjRqMe42_2),.dout(w_dff_B_NM0Y1hWn2_2),.clk(gclk));
	jdff dff_B_CGQvG3yf8_2(.din(w_dff_B_NM0Y1hWn2_2),.dout(w_dff_B_CGQvG3yf8_2),.clk(gclk));
	jdff dff_B_FBwPxAJx6_2(.din(w_dff_B_CGQvG3yf8_2),.dout(w_dff_B_FBwPxAJx6_2),.clk(gclk));
	jdff dff_B_Cd4ay4Wa8_2(.din(w_dff_B_FBwPxAJx6_2),.dout(w_dff_B_Cd4ay4Wa8_2),.clk(gclk));
	jdff dff_B_q8ta6jqp4_2(.din(w_dff_B_Cd4ay4Wa8_2),.dout(w_dff_B_q8ta6jqp4_2),.clk(gclk));
	jdff dff_B_iU8oq5SF4_2(.din(w_dff_B_q8ta6jqp4_2),.dout(w_dff_B_iU8oq5SF4_2),.clk(gclk));
	jdff dff_B_WcSJHpsH8_2(.din(w_dff_B_iU8oq5SF4_2),.dout(w_dff_B_WcSJHpsH8_2),.clk(gclk));
	jdff dff_B_sqHZn5su3_2(.din(w_dff_B_WcSJHpsH8_2),.dout(w_dff_B_sqHZn5su3_2),.clk(gclk));
	jdff dff_B_6UbglX4O2_2(.din(w_dff_B_sqHZn5su3_2),.dout(w_dff_B_6UbglX4O2_2),.clk(gclk));
	jdff dff_B_UxQgDpqq2_2(.din(w_dff_B_6UbglX4O2_2),.dout(w_dff_B_UxQgDpqq2_2),.clk(gclk));
	jdff dff_B_TYNlJLSn7_2(.din(w_dff_B_UxQgDpqq2_2),.dout(w_dff_B_TYNlJLSn7_2),.clk(gclk));
	jdff dff_B_HhpQE4kW9_2(.din(w_dff_B_TYNlJLSn7_2),.dout(w_dff_B_HhpQE4kW9_2),.clk(gclk));
	jdff dff_B_VVfQdY1B5_2(.din(w_dff_B_HhpQE4kW9_2),.dout(w_dff_B_VVfQdY1B5_2),.clk(gclk));
	jdff dff_B_Mf1IWDy81_2(.din(w_dff_B_VVfQdY1B5_2),.dout(w_dff_B_Mf1IWDy81_2),.clk(gclk));
	jdff dff_B_ZzQJFCZZ6_2(.din(w_dff_B_Mf1IWDy81_2),.dout(w_dff_B_ZzQJFCZZ6_2),.clk(gclk));
	jdff dff_B_UQ776D743_2(.din(w_dff_B_ZzQJFCZZ6_2),.dout(w_dff_B_UQ776D743_2),.clk(gclk));
	jdff dff_B_VMc7Faea5_2(.din(w_dff_B_UQ776D743_2),.dout(w_dff_B_VMc7Faea5_2),.clk(gclk));
	jdff dff_B_xB2zWgPK7_2(.din(w_dff_B_VMc7Faea5_2),.dout(w_dff_B_xB2zWgPK7_2),.clk(gclk));
	jdff dff_B_KjwqDgQE0_2(.din(w_dff_B_xB2zWgPK7_2),.dout(w_dff_B_KjwqDgQE0_2),.clk(gclk));
	jdff dff_B_UaOu27yt3_2(.din(w_dff_B_KjwqDgQE0_2),.dout(w_dff_B_UaOu27yt3_2),.clk(gclk));
	jdff dff_B_E0t5ECdE0_2(.din(w_dff_B_UaOu27yt3_2),.dout(w_dff_B_E0t5ECdE0_2),.clk(gclk));
	jdff dff_B_E1e5RC7n4_2(.din(w_dff_B_E0t5ECdE0_2),.dout(w_dff_B_E1e5RC7n4_2),.clk(gclk));
	jdff dff_B_B1p262JB2_2(.din(w_dff_B_E1e5RC7n4_2),.dout(w_dff_B_B1p262JB2_2),.clk(gclk));
	jdff dff_B_a4Ke2SEk4_2(.din(w_dff_B_B1p262JB2_2),.dout(w_dff_B_a4Ke2SEk4_2),.clk(gclk));
	jdff dff_B_lRuyGLG24_2(.din(w_dff_B_a4Ke2SEk4_2),.dout(w_dff_B_lRuyGLG24_2),.clk(gclk));
	jdff dff_B_CBStuMlU2_2(.din(w_dff_B_lRuyGLG24_2),.dout(w_dff_B_CBStuMlU2_2),.clk(gclk));
	jdff dff_B_MOifhJCc8_1(.din(n1715),.dout(w_dff_B_MOifhJCc8_1),.clk(gclk));
	jdff dff_B_lVWo6LPI0_1(.din(w_dff_B_MOifhJCc8_1),.dout(w_dff_B_lVWo6LPI0_1),.clk(gclk));
	jdff dff_B_W1fImlgg1_2(.din(n1714),.dout(w_dff_B_W1fImlgg1_2),.clk(gclk));
	jdff dff_B_gy0E2syy4_2(.din(w_dff_B_W1fImlgg1_2),.dout(w_dff_B_gy0E2syy4_2),.clk(gclk));
	jdff dff_B_8ILM1cof0_2(.din(w_dff_B_gy0E2syy4_2),.dout(w_dff_B_8ILM1cof0_2),.clk(gclk));
	jdff dff_B_XUi5sFrJ6_2(.din(w_dff_B_8ILM1cof0_2),.dout(w_dff_B_XUi5sFrJ6_2),.clk(gclk));
	jdff dff_B_kpE5Vyk67_2(.din(w_dff_B_XUi5sFrJ6_2),.dout(w_dff_B_kpE5Vyk67_2),.clk(gclk));
	jdff dff_B_5qnMg1bU9_2(.din(w_dff_B_kpE5Vyk67_2),.dout(w_dff_B_5qnMg1bU9_2),.clk(gclk));
	jdff dff_B_ziY8UmGG3_2(.din(w_dff_B_5qnMg1bU9_2),.dout(w_dff_B_ziY8UmGG3_2),.clk(gclk));
	jdff dff_B_jXk44IW77_2(.din(w_dff_B_ziY8UmGG3_2),.dout(w_dff_B_jXk44IW77_2),.clk(gclk));
	jdff dff_B_xBNwlM3J6_2(.din(w_dff_B_jXk44IW77_2),.dout(w_dff_B_xBNwlM3J6_2),.clk(gclk));
	jdff dff_B_xhbjBwyY2_2(.din(w_dff_B_xBNwlM3J6_2),.dout(w_dff_B_xhbjBwyY2_2),.clk(gclk));
	jdff dff_B_QOnKBiC72_2(.din(w_dff_B_xhbjBwyY2_2),.dout(w_dff_B_QOnKBiC72_2),.clk(gclk));
	jdff dff_B_GiLeXQaB9_2(.din(w_dff_B_QOnKBiC72_2),.dout(w_dff_B_GiLeXQaB9_2),.clk(gclk));
	jdff dff_B_CbburaLq0_2(.din(w_dff_B_GiLeXQaB9_2),.dout(w_dff_B_CbburaLq0_2),.clk(gclk));
	jdff dff_B_7c29jQdE0_2(.din(w_dff_B_CbburaLq0_2),.dout(w_dff_B_7c29jQdE0_2),.clk(gclk));
	jdff dff_B_KssGcenL7_2(.din(w_dff_B_7c29jQdE0_2),.dout(w_dff_B_KssGcenL7_2),.clk(gclk));
	jdff dff_B_ujDKBUXA5_2(.din(w_dff_B_KssGcenL7_2),.dout(w_dff_B_ujDKBUXA5_2),.clk(gclk));
	jdff dff_B_Xq3z0dH93_2(.din(w_dff_B_ujDKBUXA5_2),.dout(w_dff_B_Xq3z0dH93_2),.clk(gclk));
	jdff dff_B_vWFAv8EE2_2(.din(w_dff_B_Xq3z0dH93_2),.dout(w_dff_B_vWFAv8EE2_2),.clk(gclk));
	jdff dff_B_D5Uwx2WR9_2(.din(w_dff_B_vWFAv8EE2_2),.dout(w_dff_B_D5Uwx2WR9_2),.clk(gclk));
	jdff dff_B_7MqjbenK8_2(.din(w_dff_B_D5Uwx2WR9_2),.dout(w_dff_B_7MqjbenK8_2),.clk(gclk));
	jdff dff_B_cdfS37n29_2(.din(w_dff_B_7MqjbenK8_2),.dout(w_dff_B_cdfS37n29_2),.clk(gclk));
	jdff dff_B_LH8nCjx98_2(.din(w_dff_B_cdfS37n29_2),.dout(w_dff_B_LH8nCjx98_2),.clk(gclk));
	jdff dff_B_BA4Bn5JB6_2(.din(w_dff_B_LH8nCjx98_2),.dout(w_dff_B_BA4Bn5JB6_2),.clk(gclk));
	jdff dff_B_y1TIZDIi7_2(.din(w_dff_B_BA4Bn5JB6_2),.dout(w_dff_B_y1TIZDIi7_2),.clk(gclk));
	jdff dff_B_hjIWMQYH1_2(.din(w_dff_B_y1TIZDIi7_2),.dout(w_dff_B_hjIWMQYH1_2),.clk(gclk));
	jdff dff_B_enC1StP34_2(.din(w_dff_B_hjIWMQYH1_2),.dout(w_dff_B_enC1StP34_2),.clk(gclk));
	jdff dff_B_cVEEZnhd5_2(.din(w_dff_B_enC1StP34_2),.dout(w_dff_B_cVEEZnhd5_2),.clk(gclk));
	jdff dff_B_6aTtpjm30_2(.din(w_dff_B_cVEEZnhd5_2),.dout(w_dff_B_6aTtpjm30_2),.clk(gclk));
	jdff dff_B_59GPI1Sd1_2(.din(w_dff_B_6aTtpjm30_2),.dout(w_dff_B_59GPI1Sd1_2),.clk(gclk));
	jdff dff_B_hhpnrpPS4_2(.din(w_dff_B_59GPI1Sd1_2),.dout(w_dff_B_hhpnrpPS4_2),.clk(gclk));
	jdff dff_B_HOyvwsa40_2(.din(w_dff_B_hhpnrpPS4_2),.dout(w_dff_B_HOyvwsa40_2),.clk(gclk));
	jdff dff_B_9gvnNtA70_2(.din(w_dff_B_HOyvwsa40_2),.dout(w_dff_B_9gvnNtA70_2),.clk(gclk));
	jdff dff_B_2S7GHZ3H9_2(.din(w_dff_B_9gvnNtA70_2),.dout(w_dff_B_2S7GHZ3H9_2),.clk(gclk));
	jdff dff_B_owyP0Yx30_2(.din(w_dff_B_2S7GHZ3H9_2),.dout(w_dff_B_owyP0Yx30_2),.clk(gclk));
	jdff dff_B_tCP1VM0J5_2(.din(w_dff_B_owyP0Yx30_2),.dout(w_dff_B_tCP1VM0J5_2),.clk(gclk));
	jdff dff_B_1gNVAssC9_2(.din(w_dff_B_tCP1VM0J5_2),.dout(w_dff_B_1gNVAssC9_2),.clk(gclk));
	jdff dff_B_rZ9LUbfm1_2(.din(w_dff_B_1gNVAssC9_2),.dout(w_dff_B_rZ9LUbfm1_2),.clk(gclk));
	jdff dff_B_bELAnydM6_2(.din(w_dff_B_rZ9LUbfm1_2),.dout(w_dff_B_bELAnydM6_2),.clk(gclk));
	jdff dff_B_kyT5jDZT2_2(.din(w_dff_B_bELAnydM6_2),.dout(w_dff_B_kyT5jDZT2_2),.clk(gclk));
	jdff dff_B_mWxr1naH6_2(.din(w_dff_B_kyT5jDZT2_2),.dout(w_dff_B_mWxr1naH6_2),.clk(gclk));
	jdff dff_B_Cy9xGHOQ5_2(.din(w_dff_B_mWxr1naH6_2),.dout(w_dff_B_Cy9xGHOQ5_2),.clk(gclk));
	jdff dff_B_NDQiaCOP5_2(.din(n1713),.dout(w_dff_B_NDQiaCOP5_2),.clk(gclk));
	jdff dff_B_zte6Kcty8_2(.din(w_dff_B_NDQiaCOP5_2),.dout(w_dff_B_zte6Kcty8_2),.clk(gclk));
	jdff dff_B_pLwJsyDp8_2(.din(w_dff_B_zte6Kcty8_2),.dout(w_dff_B_pLwJsyDp8_2),.clk(gclk));
	jdff dff_B_n1SXt6eE9_2(.din(w_dff_B_pLwJsyDp8_2),.dout(w_dff_B_n1SXt6eE9_2),.clk(gclk));
	jdff dff_B_PYuac0zV5_2(.din(w_dff_B_n1SXt6eE9_2),.dout(w_dff_B_PYuac0zV5_2),.clk(gclk));
	jdff dff_B_G83IlmWl6_2(.din(w_dff_B_PYuac0zV5_2),.dout(w_dff_B_G83IlmWl6_2),.clk(gclk));
	jdff dff_B_EHe0aV8Q0_2(.din(w_dff_B_G83IlmWl6_2),.dout(w_dff_B_EHe0aV8Q0_2),.clk(gclk));
	jdff dff_B_3IGIPZVt7_2(.din(w_dff_B_EHe0aV8Q0_2),.dout(w_dff_B_3IGIPZVt7_2),.clk(gclk));
	jdff dff_B_jucUOgts6_2(.din(w_dff_B_3IGIPZVt7_2),.dout(w_dff_B_jucUOgts6_2),.clk(gclk));
	jdff dff_B_OxboZAsz4_2(.din(w_dff_B_jucUOgts6_2),.dout(w_dff_B_OxboZAsz4_2),.clk(gclk));
	jdff dff_B_tUqE9xah2_2(.din(w_dff_B_OxboZAsz4_2),.dout(w_dff_B_tUqE9xah2_2),.clk(gclk));
	jdff dff_B_GyA2b7Tc5_2(.din(w_dff_B_tUqE9xah2_2),.dout(w_dff_B_GyA2b7Tc5_2),.clk(gclk));
	jdff dff_B_cogp0iZV3_2(.din(w_dff_B_GyA2b7Tc5_2),.dout(w_dff_B_cogp0iZV3_2),.clk(gclk));
	jdff dff_B_dfHMjl051_2(.din(w_dff_B_cogp0iZV3_2),.dout(w_dff_B_dfHMjl051_2),.clk(gclk));
	jdff dff_B_N8NCNmHB5_2(.din(w_dff_B_dfHMjl051_2),.dout(w_dff_B_N8NCNmHB5_2),.clk(gclk));
	jdff dff_B_F6Vzk1BR9_2(.din(w_dff_B_N8NCNmHB5_2),.dout(w_dff_B_F6Vzk1BR9_2),.clk(gclk));
	jdff dff_B_0aaFObD03_2(.din(w_dff_B_F6Vzk1BR9_2),.dout(w_dff_B_0aaFObD03_2),.clk(gclk));
	jdff dff_B_ezSLIK7a4_2(.din(w_dff_B_0aaFObD03_2),.dout(w_dff_B_ezSLIK7a4_2),.clk(gclk));
	jdff dff_B_7MPW1RIy8_2(.din(w_dff_B_ezSLIK7a4_2),.dout(w_dff_B_7MPW1RIy8_2),.clk(gclk));
	jdff dff_B_k6dWuvBb1_2(.din(w_dff_B_7MPW1RIy8_2),.dout(w_dff_B_k6dWuvBb1_2),.clk(gclk));
	jdff dff_B_rI2td8W11_2(.din(w_dff_B_k6dWuvBb1_2),.dout(w_dff_B_rI2td8W11_2),.clk(gclk));
	jdff dff_B_NeLpJ9J22_2(.din(w_dff_B_rI2td8W11_2),.dout(w_dff_B_NeLpJ9J22_2),.clk(gclk));
	jdff dff_B_5i5q6OnL2_2(.din(w_dff_B_NeLpJ9J22_2),.dout(w_dff_B_5i5q6OnL2_2),.clk(gclk));
	jdff dff_B_Zc8aYGpA9_2(.din(w_dff_B_5i5q6OnL2_2),.dout(w_dff_B_Zc8aYGpA9_2),.clk(gclk));
	jdff dff_B_lLdbZKoH9_2(.din(w_dff_B_Zc8aYGpA9_2),.dout(w_dff_B_lLdbZKoH9_2),.clk(gclk));
	jdff dff_B_3eWry5JS6_2(.din(w_dff_B_lLdbZKoH9_2),.dout(w_dff_B_3eWry5JS6_2),.clk(gclk));
	jdff dff_B_FLlRzHmu3_2(.din(w_dff_B_3eWry5JS6_2),.dout(w_dff_B_FLlRzHmu3_2),.clk(gclk));
	jdff dff_B_EDf6ugCK0_2(.din(w_dff_B_FLlRzHmu3_2),.dout(w_dff_B_EDf6ugCK0_2),.clk(gclk));
	jdff dff_B_9wvPUEAv1_2(.din(w_dff_B_EDf6ugCK0_2),.dout(w_dff_B_9wvPUEAv1_2),.clk(gclk));
	jdff dff_B_yFTwmcv21_2(.din(w_dff_B_9wvPUEAv1_2),.dout(w_dff_B_yFTwmcv21_2),.clk(gclk));
	jdff dff_B_anBSeP584_2(.din(w_dff_B_yFTwmcv21_2),.dout(w_dff_B_anBSeP584_2),.clk(gclk));
	jdff dff_B_PjVOV9nZ7_2(.din(w_dff_B_anBSeP584_2),.dout(w_dff_B_PjVOV9nZ7_2),.clk(gclk));
	jdff dff_B_6Ldbww9W2_2(.din(w_dff_B_PjVOV9nZ7_2),.dout(w_dff_B_6Ldbww9W2_2),.clk(gclk));
	jdff dff_B_riiEll2j1_2(.din(w_dff_B_6Ldbww9W2_2),.dout(w_dff_B_riiEll2j1_2),.clk(gclk));
	jdff dff_B_mppRzF617_2(.din(w_dff_B_riiEll2j1_2),.dout(w_dff_B_mppRzF617_2),.clk(gclk));
	jdff dff_B_Qseosek06_2(.din(w_dff_B_mppRzF617_2),.dout(w_dff_B_Qseosek06_2),.clk(gclk));
	jdff dff_B_J2fetmqx3_2(.din(w_dff_B_Qseosek06_2),.dout(w_dff_B_J2fetmqx3_2),.clk(gclk));
	jdff dff_B_S6MH5rPa7_2(.din(w_dff_B_J2fetmqx3_2),.dout(w_dff_B_S6MH5rPa7_2),.clk(gclk));
	jdff dff_B_j7uGJMBe1_2(.din(w_dff_B_S6MH5rPa7_2),.dout(w_dff_B_j7uGJMBe1_2),.clk(gclk));
	jdff dff_B_MloNm4do6_2(.din(w_dff_B_j7uGJMBe1_2),.dout(w_dff_B_MloNm4do6_2),.clk(gclk));
	jdff dff_B_9KOoqiZj9_2(.din(w_dff_B_MloNm4do6_2),.dout(w_dff_B_9KOoqiZj9_2),.clk(gclk));
	jdff dff_B_rkl99rgz3_2(.din(w_dff_B_9KOoqiZj9_2),.dout(w_dff_B_rkl99rgz3_2),.clk(gclk));
	jdff dff_B_hmcBy8Y75_2(.din(w_dff_B_rkl99rgz3_2),.dout(w_dff_B_hmcBy8Y75_2),.clk(gclk));
	jdff dff_B_rttDH4w78_2(.din(n1712),.dout(w_dff_B_rttDH4w78_2),.clk(gclk));
	jdff dff_B_SN63Z6ww0_1(.din(n1710),.dout(w_dff_B_SN63Z6ww0_1),.clk(gclk));
	jdff dff_B_2w8MVoH53_2(.din(n1668),.dout(w_dff_B_2w8MVoH53_2),.clk(gclk));
	jdff dff_B_e46VTKop9_2(.din(w_dff_B_2w8MVoH53_2),.dout(w_dff_B_e46VTKop9_2),.clk(gclk));
	jdff dff_B_LSisNa268_2(.din(w_dff_B_e46VTKop9_2),.dout(w_dff_B_LSisNa268_2),.clk(gclk));
	jdff dff_B_oFCdudBJ2_2(.din(w_dff_B_LSisNa268_2),.dout(w_dff_B_oFCdudBJ2_2),.clk(gclk));
	jdff dff_B_2DjnVYRp1_2(.din(w_dff_B_oFCdudBJ2_2),.dout(w_dff_B_2DjnVYRp1_2),.clk(gclk));
	jdff dff_B_ssWz4MEp5_2(.din(w_dff_B_2DjnVYRp1_2),.dout(w_dff_B_ssWz4MEp5_2),.clk(gclk));
	jdff dff_B_of32stQY3_2(.din(w_dff_B_ssWz4MEp5_2),.dout(w_dff_B_of32stQY3_2),.clk(gclk));
	jdff dff_B_XHpujecB2_2(.din(w_dff_B_of32stQY3_2),.dout(w_dff_B_XHpujecB2_2),.clk(gclk));
	jdff dff_B_zWPvtu2x9_2(.din(w_dff_B_XHpujecB2_2),.dout(w_dff_B_zWPvtu2x9_2),.clk(gclk));
	jdff dff_B_W2e9vhvR8_2(.din(w_dff_B_zWPvtu2x9_2),.dout(w_dff_B_W2e9vhvR8_2),.clk(gclk));
	jdff dff_B_8gKzIHv56_2(.din(w_dff_B_W2e9vhvR8_2),.dout(w_dff_B_8gKzIHv56_2),.clk(gclk));
	jdff dff_B_ZFsO7iqZ2_2(.din(w_dff_B_8gKzIHv56_2),.dout(w_dff_B_ZFsO7iqZ2_2),.clk(gclk));
	jdff dff_B_YON7aJgk8_2(.din(w_dff_B_ZFsO7iqZ2_2),.dout(w_dff_B_YON7aJgk8_2),.clk(gclk));
	jdff dff_B_wC2KjiuU5_2(.din(w_dff_B_YON7aJgk8_2),.dout(w_dff_B_wC2KjiuU5_2),.clk(gclk));
	jdff dff_B_b7JHQl2A4_2(.din(w_dff_B_wC2KjiuU5_2),.dout(w_dff_B_b7JHQl2A4_2),.clk(gclk));
	jdff dff_B_2kGRweaU6_2(.din(w_dff_B_b7JHQl2A4_2),.dout(w_dff_B_2kGRweaU6_2),.clk(gclk));
	jdff dff_B_42bTzYJ90_2(.din(w_dff_B_2kGRweaU6_2),.dout(w_dff_B_42bTzYJ90_2),.clk(gclk));
	jdff dff_B_FxxJ7s439_2(.din(w_dff_B_42bTzYJ90_2),.dout(w_dff_B_FxxJ7s439_2),.clk(gclk));
	jdff dff_B_VGKt2nH15_2(.din(w_dff_B_FxxJ7s439_2),.dout(w_dff_B_VGKt2nH15_2),.clk(gclk));
	jdff dff_B_eWXal43W1_2(.din(w_dff_B_VGKt2nH15_2),.dout(w_dff_B_eWXal43W1_2),.clk(gclk));
	jdff dff_B_czxxPufb9_2(.din(w_dff_B_eWXal43W1_2),.dout(w_dff_B_czxxPufb9_2),.clk(gclk));
	jdff dff_B_LQTbmUYy2_2(.din(w_dff_B_czxxPufb9_2),.dout(w_dff_B_LQTbmUYy2_2),.clk(gclk));
	jdff dff_B_nIXyuSJv5_2(.din(w_dff_B_LQTbmUYy2_2),.dout(w_dff_B_nIXyuSJv5_2),.clk(gclk));
	jdff dff_B_1Vojf63D9_2(.din(w_dff_B_nIXyuSJv5_2),.dout(w_dff_B_1Vojf63D9_2),.clk(gclk));
	jdff dff_B_2z0zJWmN0_2(.din(w_dff_B_1Vojf63D9_2),.dout(w_dff_B_2z0zJWmN0_2),.clk(gclk));
	jdff dff_B_1q4wkFhO8_2(.din(w_dff_B_2z0zJWmN0_2),.dout(w_dff_B_1q4wkFhO8_2),.clk(gclk));
	jdff dff_B_fm9r7YsV2_2(.din(w_dff_B_1q4wkFhO8_2),.dout(w_dff_B_fm9r7YsV2_2),.clk(gclk));
	jdff dff_B_BYvTr5Qp6_2(.din(w_dff_B_fm9r7YsV2_2),.dout(w_dff_B_BYvTr5Qp6_2),.clk(gclk));
	jdff dff_B_WNFPVwXA5_2(.din(w_dff_B_BYvTr5Qp6_2),.dout(w_dff_B_WNFPVwXA5_2),.clk(gclk));
	jdff dff_B_sUnW1Sx40_2(.din(w_dff_B_WNFPVwXA5_2),.dout(w_dff_B_sUnW1Sx40_2),.clk(gclk));
	jdff dff_B_kgzbo2OC7_2(.din(w_dff_B_sUnW1Sx40_2),.dout(w_dff_B_kgzbo2OC7_2),.clk(gclk));
	jdff dff_B_VZgp7J896_2(.din(w_dff_B_kgzbo2OC7_2),.dout(w_dff_B_VZgp7J896_2),.clk(gclk));
	jdff dff_B_cIbOwcwU2_2(.din(w_dff_B_VZgp7J896_2),.dout(w_dff_B_cIbOwcwU2_2),.clk(gclk));
	jdff dff_B_bKuJ5P6R3_2(.din(w_dff_B_cIbOwcwU2_2),.dout(w_dff_B_bKuJ5P6R3_2),.clk(gclk));
	jdff dff_B_f1dZ6x8c1_2(.din(w_dff_B_bKuJ5P6R3_2),.dout(w_dff_B_f1dZ6x8c1_2),.clk(gclk));
	jdff dff_B_1DOe9Pgg1_2(.din(w_dff_B_f1dZ6x8c1_2),.dout(w_dff_B_1DOe9Pgg1_2),.clk(gclk));
	jdff dff_B_U28oDTfI7_2(.din(w_dff_B_1DOe9Pgg1_2),.dout(w_dff_B_U28oDTfI7_2),.clk(gclk));
	jdff dff_B_qBi4lIwq1_2(.din(w_dff_B_U28oDTfI7_2),.dout(w_dff_B_qBi4lIwq1_2),.clk(gclk));
	jdff dff_B_ZjWGrG8E2_2(.din(w_dff_B_qBi4lIwq1_2),.dout(w_dff_B_ZjWGrG8E2_2),.clk(gclk));
	jdff dff_B_hWflD2Rx4_2(.din(w_dff_B_ZjWGrG8E2_2),.dout(w_dff_B_hWflD2Rx4_2),.clk(gclk));
	jdff dff_B_dQiY6pmy6_1(.din(n1674),.dout(w_dff_B_dQiY6pmy6_1),.clk(gclk));
	jdff dff_B_O32QGbkt5_1(.din(w_dff_B_dQiY6pmy6_1),.dout(w_dff_B_O32QGbkt5_1),.clk(gclk));
	jdff dff_B_RClOnliE9_2(.din(n1673),.dout(w_dff_B_RClOnliE9_2),.clk(gclk));
	jdff dff_B_cz818Th53_2(.din(w_dff_B_RClOnliE9_2),.dout(w_dff_B_cz818Th53_2),.clk(gclk));
	jdff dff_B_AgdktrfV4_2(.din(w_dff_B_cz818Th53_2),.dout(w_dff_B_AgdktrfV4_2),.clk(gclk));
	jdff dff_B_SyU2s1Sj8_2(.din(w_dff_B_AgdktrfV4_2),.dout(w_dff_B_SyU2s1Sj8_2),.clk(gclk));
	jdff dff_B_TmYQ4m1W4_2(.din(w_dff_B_SyU2s1Sj8_2),.dout(w_dff_B_TmYQ4m1W4_2),.clk(gclk));
	jdff dff_B_uVMWVjQb0_2(.din(w_dff_B_TmYQ4m1W4_2),.dout(w_dff_B_uVMWVjQb0_2),.clk(gclk));
	jdff dff_B_uagxMc4J3_2(.din(w_dff_B_uVMWVjQb0_2),.dout(w_dff_B_uagxMc4J3_2),.clk(gclk));
	jdff dff_B_nedMcWL41_2(.din(w_dff_B_uagxMc4J3_2),.dout(w_dff_B_nedMcWL41_2),.clk(gclk));
	jdff dff_B_EJ602wVC7_2(.din(w_dff_B_nedMcWL41_2),.dout(w_dff_B_EJ602wVC7_2),.clk(gclk));
	jdff dff_B_zNRMbOVC5_2(.din(w_dff_B_EJ602wVC7_2),.dout(w_dff_B_zNRMbOVC5_2),.clk(gclk));
	jdff dff_B_O0XDEz0J2_2(.din(w_dff_B_zNRMbOVC5_2),.dout(w_dff_B_O0XDEz0J2_2),.clk(gclk));
	jdff dff_B_tMbhbP9K9_2(.din(w_dff_B_O0XDEz0J2_2),.dout(w_dff_B_tMbhbP9K9_2),.clk(gclk));
	jdff dff_B_GtMLA1TE7_2(.din(w_dff_B_tMbhbP9K9_2),.dout(w_dff_B_GtMLA1TE7_2),.clk(gclk));
	jdff dff_B_CfVVt80c6_2(.din(w_dff_B_GtMLA1TE7_2),.dout(w_dff_B_CfVVt80c6_2),.clk(gclk));
	jdff dff_B_PNLk8pWd3_2(.din(w_dff_B_CfVVt80c6_2),.dout(w_dff_B_PNLk8pWd3_2),.clk(gclk));
	jdff dff_B_amDPAmdF1_2(.din(w_dff_B_PNLk8pWd3_2),.dout(w_dff_B_amDPAmdF1_2),.clk(gclk));
	jdff dff_B_zqrndod36_2(.din(w_dff_B_amDPAmdF1_2),.dout(w_dff_B_zqrndod36_2),.clk(gclk));
	jdff dff_B_fT7OgN7M8_2(.din(w_dff_B_zqrndod36_2),.dout(w_dff_B_fT7OgN7M8_2),.clk(gclk));
	jdff dff_B_CG8ZfgVv1_2(.din(w_dff_B_fT7OgN7M8_2),.dout(w_dff_B_CG8ZfgVv1_2),.clk(gclk));
	jdff dff_B_druNSZnM0_2(.din(w_dff_B_CG8ZfgVv1_2),.dout(w_dff_B_druNSZnM0_2),.clk(gclk));
	jdff dff_B_wDy28X018_2(.din(w_dff_B_druNSZnM0_2),.dout(w_dff_B_wDy28X018_2),.clk(gclk));
	jdff dff_B_VvoJFzTR3_2(.din(w_dff_B_wDy28X018_2),.dout(w_dff_B_VvoJFzTR3_2),.clk(gclk));
	jdff dff_B_EB4uBugq0_2(.din(w_dff_B_VvoJFzTR3_2),.dout(w_dff_B_EB4uBugq0_2),.clk(gclk));
	jdff dff_B_2T1XdtDl1_2(.din(w_dff_B_EB4uBugq0_2),.dout(w_dff_B_2T1XdtDl1_2),.clk(gclk));
	jdff dff_B_BbgYCdJ65_2(.din(w_dff_B_2T1XdtDl1_2),.dout(w_dff_B_BbgYCdJ65_2),.clk(gclk));
	jdff dff_B_Kz6osrUH9_2(.din(w_dff_B_BbgYCdJ65_2),.dout(w_dff_B_Kz6osrUH9_2),.clk(gclk));
	jdff dff_B_J4nBOsCP7_2(.din(w_dff_B_Kz6osrUH9_2),.dout(w_dff_B_J4nBOsCP7_2),.clk(gclk));
	jdff dff_B_IQTdUg0M8_2(.din(w_dff_B_J4nBOsCP7_2),.dout(w_dff_B_IQTdUg0M8_2),.clk(gclk));
	jdff dff_B_vqVDl74n0_2(.din(w_dff_B_IQTdUg0M8_2),.dout(w_dff_B_vqVDl74n0_2),.clk(gclk));
	jdff dff_B_s38a6tfY1_2(.din(w_dff_B_vqVDl74n0_2),.dout(w_dff_B_s38a6tfY1_2),.clk(gclk));
	jdff dff_B_HFPoG2LJ8_2(.din(w_dff_B_s38a6tfY1_2),.dout(w_dff_B_HFPoG2LJ8_2),.clk(gclk));
	jdff dff_B_nYTioUsq0_2(.din(w_dff_B_HFPoG2LJ8_2),.dout(w_dff_B_nYTioUsq0_2),.clk(gclk));
	jdff dff_B_gwJqSQnA4_2(.din(w_dff_B_nYTioUsq0_2),.dout(w_dff_B_gwJqSQnA4_2),.clk(gclk));
	jdff dff_B_lBSLs1DI8_2(.din(w_dff_B_gwJqSQnA4_2),.dout(w_dff_B_lBSLs1DI8_2),.clk(gclk));
	jdff dff_B_NN8zJ1x25_2(.din(w_dff_B_lBSLs1DI8_2),.dout(w_dff_B_NN8zJ1x25_2),.clk(gclk));
	jdff dff_B_OZfqgxWB4_2(.din(w_dff_B_NN8zJ1x25_2),.dout(w_dff_B_OZfqgxWB4_2),.clk(gclk));
	jdff dff_B_6Y8cJT6S0_2(.din(w_dff_B_OZfqgxWB4_2),.dout(w_dff_B_6Y8cJT6S0_2),.clk(gclk));
	jdff dff_B_gsjuqBPn0_2(.din(n1672),.dout(w_dff_B_gsjuqBPn0_2),.clk(gclk));
	jdff dff_B_l7Sj046f1_2(.din(w_dff_B_gsjuqBPn0_2),.dout(w_dff_B_l7Sj046f1_2),.clk(gclk));
	jdff dff_B_RZB5afjY7_2(.din(w_dff_B_l7Sj046f1_2),.dout(w_dff_B_RZB5afjY7_2),.clk(gclk));
	jdff dff_B_imRLAERZ0_2(.din(w_dff_B_RZB5afjY7_2),.dout(w_dff_B_imRLAERZ0_2),.clk(gclk));
	jdff dff_B_t5lxNJun8_2(.din(w_dff_B_imRLAERZ0_2),.dout(w_dff_B_t5lxNJun8_2),.clk(gclk));
	jdff dff_B_Z0BtaOVv9_2(.din(w_dff_B_t5lxNJun8_2),.dout(w_dff_B_Z0BtaOVv9_2),.clk(gclk));
	jdff dff_B_7ftk6shM5_2(.din(w_dff_B_Z0BtaOVv9_2),.dout(w_dff_B_7ftk6shM5_2),.clk(gclk));
	jdff dff_B_SJYor4cu9_2(.din(w_dff_B_7ftk6shM5_2),.dout(w_dff_B_SJYor4cu9_2),.clk(gclk));
	jdff dff_B_PYdspwWx5_2(.din(w_dff_B_SJYor4cu9_2),.dout(w_dff_B_PYdspwWx5_2),.clk(gclk));
	jdff dff_B_TdwCeMJV4_2(.din(w_dff_B_PYdspwWx5_2),.dout(w_dff_B_TdwCeMJV4_2),.clk(gclk));
	jdff dff_B_r2JSgjXJ2_2(.din(w_dff_B_TdwCeMJV4_2),.dout(w_dff_B_r2JSgjXJ2_2),.clk(gclk));
	jdff dff_B_vNvxmP1U6_2(.din(w_dff_B_r2JSgjXJ2_2),.dout(w_dff_B_vNvxmP1U6_2),.clk(gclk));
	jdff dff_B_EJ1Pm7es9_2(.din(w_dff_B_vNvxmP1U6_2),.dout(w_dff_B_EJ1Pm7es9_2),.clk(gclk));
	jdff dff_B_rQDUj1Vr9_2(.din(w_dff_B_EJ1Pm7es9_2),.dout(w_dff_B_rQDUj1Vr9_2),.clk(gclk));
	jdff dff_B_GNSPR3aJ4_2(.din(w_dff_B_rQDUj1Vr9_2),.dout(w_dff_B_GNSPR3aJ4_2),.clk(gclk));
	jdff dff_B_JI6uYzf38_2(.din(w_dff_B_GNSPR3aJ4_2),.dout(w_dff_B_JI6uYzf38_2),.clk(gclk));
	jdff dff_B_9C6Rr72o8_2(.din(w_dff_B_JI6uYzf38_2),.dout(w_dff_B_9C6Rr72o8_2),.clk(gclk));
	jdff dff_B_aLlZACOc9_2(.din(w_dff_B_9C6Rr72o8_2),.dout(w_dff_B_aLlZACOc9_2),.clk(gclk));
	jdff dff_B_RULpIXsq8_2(.din(w_dff_B_aLlZACOc9_2),.dout(w_dff_B_RULpIXsq8_2),.clk(gclk));
	jdff dff_B_Zsy0vRJv1_2(.din(w_dff_B_RULpIXsq8_2),.dout(w_dff_B_Zsy0vRJv1_2),.clk(gclk));
	jdff dff_B_IXMaCWHe2_2(.din(w_dff_B_Zsy0vRJv1_2),.dout(w_dff_B_IXMaCWHe2_2),.clk(gclk));
	jdff dff_B_GA5bSx567_2(.din(w_dff_B_IXMaCWHe2_2),.dout(w_dff_B_GA5bSx567_2),.clk(gclk));
	jdff dff_B_8ZFvWMEG0_2(.din(w_dff_B_GA5bSx567_2),.dout(w_dff_B_8ZFvWMEG0_2),.clk(gclk));
	jdff dff_B_2rgNDfTq6_2(.din(w_dff_B_8ZFvWMEG0_2),.dout(w_dff_B_2rgNDfTq6_2),.clk(gclk));
	jdff dff_B_2Sgye0nx5_2(.din(w_dff_B_2rgNDfTq6_2),.dout(w_dff_B_2Sgye0nx5_2),.clk(gclk));
	jdff dff_B_CGz959fP4_2(.din(w_dff_B_2Sgye0nx5_2),.dout(w_dff_B_CGz959fP4_2),.clk(gclk));
	jdff dff_B_UMDIFo0e1_2(.din(w_dff_B_CGz959fP4_2),.dout(w_dff_B_UMDIFo0e1_2),.clk(gclk));
	jdff dff_B_YXTPGBjk7_2(.din(w_dff_B_UMDIFo0e1_2),.dout(w_dff_B_YXTPGBjk7_2),.clk(gclk));
	jdff dff_B_HdXbFFF26_2(.din(w_dff_B_YXTPGBjk7_2),.dout(w_dff_B_HdXbFFF26_2),.clk(gclk));
	jdff dff_B_JAJzgZW73_2(.din(w_dff_B_HdXbFFF26_2),.dout(w_dff_B_JAJzgZW73_2),.clk(gclk));
	jdff dff_B_SlyuKEI28_2(.din(w_dff_B_JAJzgZW73_2),.dout(w_dff_B_SlyuKEI28_2),.clk(gclk));
	jdff dff_B_7gktJ1yw4_2(.din(w_dff_B_SlyuKEI28_2),.dout(w_dff_B_7gktJ1yw4_2),.clk(gclk));
	jdff dff_B_Jns0gf7Z7_2(.din(w_dff_B_7gktJ1yw4_2),.dout(w_dff_B_Jns0gf7Z7_2),.clk(gclk));
	jdff dff_B_Oky6VBgY6_2(.din(w_dff_B_Jns0gf7Z7_2),.dout(w_dff_B_Oky6VBgY6_2),.clk(gclk));
	jdff dff_B_AZEJgdk93_2(.din(w_dff_B_Oky6VBgY6_2),.dout(w_dff_B_AZEJgdk93_2),.clk(gclk));
	jdff dff_B_XYX6scPp4_2(.din(w_dff_B_AZEJgdk93_2),.dout(w_dff_B_XYX6scPp4_2),.clk(gclk));
	jdff dff_B_XK6G5zYL8_2(.din(w_dff_B_XYX6scPp4_2),.dout(w_dff_B_XK6G5zYL8_2),.clk(gclk));
	jdff dff_B_cHEqulFX0_2(.din(w_dff_B_XK6G5zYL8_2),.dout(w_dff_B_cHEqulFX0_2),.clk(gclk));
	jdff dff_B_kJbWkHSd9_2(.din(w_dff_B_cHEqulFX0_2),.dout(w_dff_B_kJbWkHSd9_2),.clk(gclk));
	jdff dff_B_Gi5MsAd61_2(.din(n1671),.dout(w_dff_B_Gi5MsAd61_2),.clk(gclk));
	jdff dff_B_df8nTyr38_1(.din(n1669),.dout(w_dff_B_df8nTyr38_1),.clk(gclk));
	jdff dff_B_Kc3JxjFy3_2(.din(n1617),.dout(w_dff_B_Kc3JxjFy3_2),.clk(gclk));
	jdff dff_B_ab32jLiY5_2(.din(w_dff_B_Kc3JxjFy3_2),.dout(w_dff_B_ab32jLiY5_2),.clk(gclk));
	jdff dff_B_OdUybZNN6_2(.din(w_dff_B_ab32jLiY5_2),.dout(w_dff_B_OdUybZNN6_2),.clk(gclk));
	jdff dff_B_MahVShMK0_2(.din(w_dff_B_OdUybZNN6_2),.dout(w_dff_B_MahVShMK0_2),.clk(gclk));
	jdff dff_B_WpV9de4t7_2(.din(w_dff_B_MahVShMK0_2),.dout(w_dff_B_WpV9de4t7_2),.clk(gclk));
	jdff dff_B_neJ2wEdv6_2(.din(w_dff_B_WpV9de4t7_2),.dout(w_dff_B_neJ2wEdv6_2),.clk(gclk));
	jdff dff_B_8bp1GZPb0_2(.din(w_dff_B_neJ2wEdv6_2),.dout(w_dff_B_8bp1GZPb0_2),.clk(gclk));
	jdff dff_B_bhOwstdk1_2(.din(w_dff_B_8bp1GZPb0_2),.dout(w_dff_B_bhOwstdk1_2),.clk(gclk));
	jdff dff_B_HROPr6sp4_2(.din(w_dff_B_bhOwstdk1_2),.dout(w_dff_B_HROPr6sp4_2),.clk(gclk));
	jdff dff_B_udesApIZ9_2(.din(w_dff_B_HROPr6sp4_2),.dout(w_dff_B_udesApIZ9_2),.clk(gclk));
	jdff dff_B_LDMCuwR39_2(.din(w_dff_B_udesApIZ9_2),.dout(w_dff_B_LDMCuwR39_2),.clk(gclk));
	jdff dff_B_jFyLK0dc0_2(.din(w_dff_B_LDMCuwR39_2),.dout(w_dff_B_jFyLK0dc0_2),.clk(gclk));
	jdff dff_B_uimemobK6_2(.din(w_dff_B_jFyLK0dc0_2),.dout(w_dff_B_uimemobK6_2),.clk(gclk));
	jdff dff_B_vPCTWK6K1_2(.din(w_dff_B_uimemobK6_2),.dout(w_dff_B_vPCTWK6K1_2),.clk(gclk));
	jdff dff_B_PGVuK9349_2(.din(w_dff_B_vPCTWK6K1_2),.dout(w_dff_B_PGVuK9349_2),.clk(gclk));
	jdff dff_B_9Ii5kWkm0_2(.din(w_dff_B_PGVuK9349_2),.dout(w_dff_B_9Ii5kWkm0_2),.clk(gclk));
	jdff dff_B_3TsY9hxj0_2(.din(w_dff_B_9Ii5kWkm0_2),.dout(w_dff_B_3TsY9hxj0_2),.clk(gclk));
	jdff dff_B_YSVlqAD68_2(.din(w_dff_B_3TsY9hxj0_2),.dout(w_dff_B_YSVlqAD68_2),.clk(gclk));
	jdff dff_B_UI7fXv842_2(.din(w_dff_B_YSVlqAD68_2),.dout(w_dff_B_UI7fXv842_2),.clk(gclk));
	jdff dff_B_ZvBh2sIL5_2(.din(w_dff_B_UI7fXv842_2),.dout(w_dff_B_ZvBh2sIL5_2),.clk(gclk));
	jdff dff_B_dVzk8pWh9_2(.din(w_dff_B_ZvBh2sIL5_2),.dout(w_dff_B_dVzk8pWh9_2),.clk(gclk));
	jdff dff_B_hgfIgNlB0_2(.din(w_dff_B_dVzk8pWh9_2),.dout(w_dff_B_hgfIgNlB0_2),.clk(gclk));
	jdff dff_B_GBdlN8tU1_2(.din(w_dff_B_hgfIgNlB0_2),.dout(w_dff_B_GBdlN8tU1_2),.clk(gclk));
	jdff dff_B_RryZuItE0_2(.din(w_dff_B_GBdlN8tU1_2),.dout(w_dff_B_RryZuItE0_2),.clk(gclk));
	jdff dff_B_yvTMCjiP7_2(.din(w_dff_B_RryZuItE0_2),.dout(w_dff_B_yvTMCjiP7_2),.clk(gclk));
	jdff dff_B_RkzM8Yi26_2(.din(w_dff_B_yvTMCjiP7_2),.dout(w_dff_B_RkzM8Yi26_2),.clk(gclk));
	jdff dff_B_NTPSMIke1_2(.din(w_dff_B_RkzM8Yi26_2),.dout(w_dff_B_NTPSMIke1_2),.clk(gclk));
	jdff dff_B_eUYmdRU37_2(.din(w_dff_B_NTPSMIke1_2),.dout(w_dff_B_eUYmdRU37_2),.clk(gclk));
	jdff dff_B_MhSWmCHF2_2(.din(w_dff_B_eUYmdRU37_2),.dout(w_dff_B_MhSWmCHF2_2),.clk(gclk));
	jdff dff_B_wqkcv9TC5_2(.din(w_dff_B_MhSWmCHF2_2),.dout(w_dff_B_wqkcv9TC5_2),.clk(gclk));
	jdff dff_B_doWquLHD6_2(.din(w_dff_B_wqkcv9TC5_2),.dout(w_dff_B_doWquLHD6_2),.clk(gclk));
	jdff dff_B_pA8vGTAg6_2(.din(w_dff_B_doWquLHD6_2),.dout(w_dff_B_pA8vGTAg6_2),.clk(gclk));
	jdff dff_B_0m6J8dqN9_2(.din(w_dff_B_pA8vGTAg6_2),.dout(w_dff_B_0m6J8dqN9_2),.clk(gclk));
	jdff dff_B_4MiELK345_2(.din(w_dff_B_0m6J8dqN9_2),.dout(w_dff_B_4MiELK345_2),.clk(gclk));
	jdff dff_B_47ewNo307_2(.din(w_dff_B_4MiELK345_2),.dout(w_dff_B_47ewNo307_2),.clk(gclk));
	jdff dff_B_wjKxITkK3_2(.din(w_dff_B_47ewNo307_2),.dout(w_dff_B_wjKxITkK3_2),.clk(gclk));
	jdff dff_B_WJYGTsHj0_1(.din(n1623),.dout(w_dff_B_WJYGTsHj0_1),.clk(gclk));
	jdff dff_B_Hip9cB0c0_1(.din(w_dff_B_WJYGTsHj0_1),.dout(w_dff_B_Hip9cB0c0_1),.clk(gclk));
	jdff dff_B_fqZYClF17_2(.din(n1622),.dout(w_dff_B_fqZYClF17_2),.clk(gclk));
	jdff dff_B_XBTvMr9v1_2(.din(w_dff_B_fqZYClF17_2),.dout(w_dff_B_XBTvMr9v1_2),.clk(gclk));
	jdff dff_B_ghMS6MsN1_2(.din(w_dff_B_XBTvMr9v1_2),.dout(w_dff_B_ghMS6MsN1_2),.clk(gclk));
	jdff dff_B_59i6FpCy2_2(.din(w_dff_B_ghMS6MsN1_2),.dout(w_dff_B_59i6FpCy2_2),.clk(gclk));
	jdff dff_B_moRsaybu7_2(.din(w_dff_B_59i6FpCy2_2),.dout(w_dff_B_moRsaybu7_2),.clk(gclk));
	jdff dff_B_rcFslrCy7_2(.din(w_dff_B_moRsaybu7_2),.dout(w_dff_B_rcFslrCy7_2),.clk(gclk));
	jdff dff_B_hSELKlPW8_2(.din(w_dff_B_rcFslrCy7_2),.dout(w_dff_B_hSELKlPW8_2),.clk(gclk));
	jdff dff_B_UG3916dJ5_2(.din(w_dff_B_hSELKlPW8_2),.dout(w_dff_B_UG3916dJ5_2),.clk(gclk));
	jdff dff_B_dZRTrxZB6_2(.din(w_dff_B_UG3916dJ5_2),.dout(w_dff_B_dZRTrxZB6_2),.clk(gclk));
	jdff dff_B_b1N6H1r40_2(.din(w_dff_B_dZRTrxZB6_2),.dout(w_dff_B_b1N6H1r40_2),.clk(gclk));
	jdff dff_B_5IbtYzTC1_2(.din(w_dff_B_b1N6H1r40_2),.dout(w_dff_B_5IbtYzTC1_2),.clk(gclk));
	jdff dff_B_OCzzEgDC8_2(.din(w_dff_B_5IbtYzTC1_2),.dout(w_dff_B_OCzzEgDC8_2),.clk(gclk));
	jdff dff_B_ipgcKSCe3_2(.din(w_dff_B_OCzzEgDC8_2),.dout(w_dff_B_ipgcKSCe3_2),.clk(gclk));
	jdff dff_B_R4VJ3Sr68_2(.din(w_dff_B_ipgcKSCe3_2),.dout(w_dff_B_R4VJ3Sr68_2),.clk(gclk));
	jdff dff_B_2wY2V7gg0_2(.din(w_dff_B_R4VJ3Sr68_2),.dout(w_dff_B_2wY2V7gg0_2),.clk(gclk));
	jdff dff_B_1evDCg2j8_2(.din(w_dff_B_2wY2V7gg0_2),.dout(w_dff_B_1evDCg2j8_2),.clk(gclk));
	jdff dff_B_t4L0GnZx2_2(.din(w_dff_B_1evDCg2j8_2),.dout(w_dff_B_t4L0GnZx2_2),.clk(gclk));
	jdff dff_B_zFJza9Af3_2(.din(w_dff_B_t4L0GnZx2_2),.dout(w_dff_B_zFJza9Af3_2),.clk(gclk));
	jdff dff_B_AZzzrBBw1_2(.din(w_dff_B_zFJza9Af3_2),.dout(w_dff_B_AZzzrBBw1_2),.clk(gclk));
	jdff dff_B_VXIVymVf9_2(.din(w_dff_B_AZzzrBBw1_2),.dout(w_dff_B_VXIVymVf9_2),.clk(gclk));
	jdff dff_B_uVoM8roE6_2(.din(w_dff_B_VXIVymVf9_2),.dout(w_dff_B_uVoM8roE6_2),.clk(gclk));
	jdff dff_B_ZhdP4AXv9_2(.din(w_dff_B_uVoM8roE6_2),.dout(w_dff_B_ZhdP4AXv9_2),.clk(gclk));
	jdff dff_B_3XsMJqFg2_2(.din(w_dff_B_ZhdP4AXv9_2),.dout(w_dff_B_3XsMJqFg2_2),.clk(gclk));
	jdff dff_B_w0xk2gsv6_2(.din(w_dff_B_3XsMJqFg2_2),.dout(w_dff_B_w0xk2gsv6_2),.clk(gclk));
	jdff dff_B_93wGTiVo5_2(.din(w_dff_B_w0xk2gsv6_2),.dout(w_dff_B_93wGTiVo5_2),.clk(gclk));
	jdff dff_B_V89d4gDM0_2(.din(w_dff_B_93wGTiVo5_2),.dout(w_dff_B_V89d4gDM0_2),.clk(gclk));
	jdff dff_B_ng2Se3Qv8_2(.din(w_dff_B_V89d4gDM0_2),.dout(w_dff_B_ng2Se3Qv8_2),.clk(gclk));
	jdff dff_B_7RSODiMM0_2(.din(w_dff_B_ng2Se3Qv8_2),.dout(w_dff_B_7RSODiMM0_2),.clk(gclk));
	jdff dff_B_xEekS89M6_2(.din(w_dff_B_7RSODiMM0_2),.dout(w_dff_B_xEekS89M6_2),.clk(gclk));
	jdff dff_B_zJbCZklX8_2(.din(w_dff_B_xEekS89M6_2),.dout(w_dff_B_zJbCZklX8_2),.clk(gclk));
	jdff dff_B_ipcv16086_2(.din(w_dff_B_zJbCZklX8_2),.dout(w_dff_B_ipcv16086_2),.clk(gclk));
	jdff dff_B_TTARY8Rj9_2(.din(w_dff_B_ipcv16086_2),.dout(w_dff_B_TTARY8Rj9_2),.clk(gclk));
	jdff dff_B_a3zElpLN1_2(.din(w_dff_B_TTARY8Rj9_2),.dout(w_dff_B_a3zElpLN1_2),.clk(gclk));
	jdff dff_B_KWKAVASx4_2(.din(n1621),.dout(w_dff_B_KWKAVASx4_2),.clk(gclk));
	jdff dff_B_P1kuuF9V8_2(.din(w_dff_B_KWKAVASx4_2),.dout(w_dff_B_P1kuuF9V8_2),.clk(gclk));
	jdff dff_B_RGR5oJBC5_2(.din(w_dff_B_P1kuuF9V8_2),.dout(w_dff_B_RGR5oJBC5_2),.clk(gclk));
	jdff dff_B_Zd3O4XIk4_2(.din(w_dff_B_RGR5oJBC5_2),.dout(w_dff_B_Zd3O4XIk4_2),.clk(gclk));
	jdff dff_B_xRXXHCDU5_2(.din(w_dff_B_Zd3O4XIk4_2),.dout(w_dff_B_xRXXHCDU5_2),.clk(gclk));
	jdff dff_B_zNHXZvMf2_2(.din(w_dff_B_xRXXHCDU5_2),.dout(w_dff_B_zNHXZvMf2_2),.clk(gclk));
	jdff dff_B_BCyv68xR5_2(.din(w_dff_B_zNHXZvMf2_2),.dout(w_dff_B_BCyv68xR5_2),.clk(gclk));
	jdff dff_B_znL5EFci3_2(.din(w_dff_B_BCyv68xR5_2),.dout(w_dff_B_znL5EFci3_2),.clk(gclk));
	jdff dff_B_VZoOeUAS0_2(.din(w_dff_B_znL5EFci3_2),.dout(w_dff_B_VZoOeUAS0_2),.clk(gclk));
	jdff dff_B_su47rQAO5_2(.din(w_dff_B_VZoOeUAS0_2),.dout(w_dff_B_su47rQAO5_2),.clk(gclk));
	jdff dff_B_Vh8qAGoS0_2(.din(w_dff_B_su47rQAO5_2),.dout(w_dff_B_Vh8qAGoS0_2),.clk(gclk));
	jdff dff_B_TDBdd1qY1_2(.din(w_dff_B_Vh8qAGoS0_2),.dout(w_dff_B_TDBdd1qY1_2),.clk(gclk));
	jdff dff_B_3764zBtX5_2(.din(w_dff_B_TDBdd1qY1_2),.dout(w_dff_B_3764zBtX5_2),.clk(gclk));
	jdff dff_B_NnQj9aBl4_2(.din(w_dff_B_3764zBtX5_2),.dout(w_dff_B_NnQj9aBl4_2),.clk(gclk));
	jdff dff_B_nBeaxeVp2_2(.din(w_dff_B_NnQj9aBl4_2),.dout(w_dff_B_nBeaxeVp2_2),.clk(gclk));
	jdff dff_B_hWjvjyXJ5_2(.din(w_dff_B_nBeaxeVp2_2),.dout(w_dff_B_hWjvjyXJ5_2),.clk(gclk));
	jdff dff_B_w6Yd3EN50_2(.din(w_dff_B_hWjvjyXJ5_2),.dout(w_dff_B_w6Yd3EN50_2),.clk(gclk));
	jdff dff_B_uwE98vtO7_2(.din(w_dff_B_w6Yd3EN50_2),.dout(w_dff_B_uwE98vtO7_2),.clk(gclk));
	jdff dff_B_dIrjrwRw6_2(.din(w_dff_B_uwE98vtO7_2),.dout(w_dff_B_dIrjrwRw6_2),.clk(gclk));
	jdff dff_B_vlMeF1YR0_2(.din(w_dff_B_dIrjrwRw6_2),.dout(w_dff_B_vlMeF1YR0_2),.clk(gclk));
	jdff dff_B_GkYapuNh0_2(.din(w_dff_B_vlMeF1YR0_2),.dout(w_dff_B_GkYapuNh0_2),.clk(gclk));
	jdff dff_B_Djwi7hZv2_2(.din(w_dff_B_GkYapuNh0_2),.dout(w_dff_B_Djwi7hZv2_2),.clk(gclk));
	jdff dff_B_dlcXEriD3_2(.din(w_dff_B_Djwi7hZv2_2),.dout(w_dff_B_dlcXEriD3_2),.clk(gclk));
	jdff dff_B_p1SbDHGp7_2(.din(w_dff_B_dlcXEriD3_2),.dout(w_dff_B_p1SbDHGp7_2),.clk(gclk));
	jdff dff_B_YEAecKDB7_2(.din(w_dff_B_p1SbDHGp7_2),.dout(w_dff_B_YEAecKDB7_2),.clk(gclk));
	jdff dff_B_agpdSzXV4_2(.din(w_dff_B_YEAecKDB7_2),.dout(w_dff_B_agpdSzXV4_2),.clk(gclk));
	jdff dff_B_7c1YjoS18_2(.din(w_dff_B_agpdSzXV4_2),.dout(w_dff_B_7c1YjoS18_2),.clk(gclk));
	jdff dff_B_Uyo0hUlD6_2(.din(w_dff_B_7c1YjoS18_2),.dout(w_dff_B_Uyo0hUlD6_2),.clk(gclk));
	jdff dff_B_lhHaqCbk2_2(.din(w_dff_B_Uyo0hUlD6_2),.dout(w_dff_B_lhHaqCbk2_2),.clk(gclk));
	jdff dff_B_Jg0HP3nZ6_2(.din(w_dff_B_lhHaqCbk2_2),.dout(w_dff_B_Jg0HP3nZ6_2),.clk(gclk));
	jdff dff_B_r2J4KLyT0_2(.din(w_dff_B_Jg0HP3nZ6_2),.dout(w_dff_B_r2J4KLyT0_2),.clk(gclk));
	jdff dff_B_Q5bAYjee7_2(.din(w_dff_B_r2J4KLyT0_2),.dout(w_dff_B_Q5bAYjee7_2),.clk(gclk));
	jdff dff_B_APvONUqZ7_2(.din(w_dff_B_Q5bAYjee7_2),.dout(w_dff_B_APvONUqZ7_2),.clk(gclk));
	jdff dff_B_5BiHwCAM0_2(.din(w_dff_B_APvONUqZ7_2),.dout(w_dff_B_5BiHwCAM0_2),.clk(gclk));
	jdff dff_B_6V8zst9C7_2(.din(w_dff_B_5BiHwCAM0_2),.dout(w_dff_B_6V8zst9C7_2),.clk(gclk));
	jdff dff_B_jQ8wPSVW4_2(.din(n1620),.dout(w_dff_B_jQ8wPSVW4_2),.clk(gclk));
	jdff dff_B_LwpMB43I2_1(.din(n1618),.dout(w_dff_B_LwpMB43I2_1),.clk(gclk));
	jdff dff_B_GugcLrnm6_2(.din(n1560),.dout(w_dff_B_GugcLrnm6_2),.clk(gclk));
	jdff dff_B_AbZlQYC56_2(.din(w_dff_B_GugcLrnm6_2),.dout(w_dff_B_AbZlQYC56_2),.clk(gclk));
	jdff dff_B_TZ8AIovi4_2(.din(w_dff_B_AbZlQYC56_2),.dout(w_dff_B_TZ8AIovi4_2),.clk(gclk));
	jdff dff_B_RHITzt4v1_2(.din(w_dff_B_TZ8AIovi4_2),.dout(w_dff_B_RHITzt4v1_2),.clk(gclk));
	jdff dff_B_NoDuwryF8_2(.din(w_dff_B_RHITzt4v1_2),.dout(w_dff_B_NoDuwryF8_2),.clk(gclk));
	jdff dff_B_wyoowKMJ2_2(.din(w_dff_B_NoDuwryF8_2),.dout(w_dff_B_wyoowKMJ2_2),.clk(gclk));
	jdff dff_B_DjjCQl1h6_2(.din(w_dff_B_wyoowKMJ2_2),.dout(w_dff_B_DjjCQl1h6_2),.clk(gclk));
	jdff dff_B_OnTXUDJC7_2(.din(w_dff_B_DjjCQl1h6_2),.dout(w_dff_B_OnTXUDJC7_2),.clk(gclk));
	jdff dff_B_mWvhFxjm4_2(.din(w_dff_B_OnTXUDJC7_2),.dout(w_dff_B_mWvhFxjm4_2),.clk(gclk));
	jdff dff_B_j91NeEOV8_2(.din(w_dff_B_mWvhFxjm4_2),.dout(w_dff_B_j91NeEOV8_2),.clk(gclk));
	jdff dff_B_ba1GqPRL1_2(.din(w_dff_B_j91NeEOV8_2),.dout(w_dff_B_ba1GqPRL1_2),.clk(gclk));
	jdff dff_B_COn85NbT6_2(.din(w_dff_B_ba1GqPRL1_2),.dout(w_dff_B_COn85NbT6_2),.clk(gclk));
	jdff dff_B_F1bmglqz6_2(.din(w_dff_B_COn85NbT6_2),.dout(w_dff_B_F1bmglqz6_2),.clk(gclk));
	jdff dff_B_rusZJjk15_2(.din(w_dff_B_F1bmglqz6_2),.dout(w_dff_B_rusZJjk15_2),.clk(gclk));
	jdff dff_B_rjQ0MfK38_2(.din(w_dff_B_rusZJjk15_2),.dout(w_dff_B_rjQ0MfK38_2),.clk(gclk));
	jdff dff_B_uPzjkIAx0_2(.din(w_dff_B_rjQ0MfK38_2),.dout(w_dff_B_uPzjkIAx0_2),.clk(gclk));
	jdff dff_B_GVjPtiHJ5_2(.din(w_dff_B_uPzjkIAx0_2),.dout(w_dff_B_GVjPtiHJ5_2),.clk(gclk));
	jdff dff_B_EWDpgouP8_2(.din(w_dff_B_GVjPtiHJ5_2),.dout(w_dff_B_EWDpgouP8_2),.clk(gclk));
	jdff dff_B_EYyV6B744_2(.din(w_dff_B_EWDpgouP8_2),.dout(w_dff_B_EYyV6B744_2),.clk(gclk));
	jdff dff_B_SIrYyk2z7_2(.din(w_dff_B_EYyV6B744_2),.dout(w_dff_B_SIrYyk2z7_2),.clk(gclk));
	jdff dff_B_fXrWZS0D5_2(.din(w_dff_B_SIrYyk2z7_2),.dout(w_dff_B_fXrWZS0D5_2),.clk(gclk));
	jdff dff_B_SCO1RFWY4_2(.din(w_dff_B_fXrWZS0D5_2),.dout(w_dff_B_SCO1RFWY4_2),.clk(gclk));
	jdff dff_B_whHMKccd6_2(.din(w_dff_B_SCO1RFWY4_2),.dout(w_dff_B_whHMKccd6_2),.clk(gclk));
	jdff dff_B_qWG4D4Zx9_2(.din(w_dff_B_whHMKccd6_2),.dout(w_dff_B_qWG4D4Zx9_2),.clk(gclk));
	jdff dff_B_uD3e3aUz3_2(.din(w_dff_B_qWG4D4Zx9_2),.dout(w_dff_B_uD3e3aUz3_2),.clk(gclk));
	jdff dff_B_n9LNErZ02_2(.din(w_dff_B_uD3e3aUz3_2),.dout(w_dff_B_n9LNErZ02_2),.clk(gclk));
	jdff dff_B_oQp4IJEg0_2(.din(w_dff_B_n9LNErZ02_2),.dout(w_dff_B_oQp4IJEg0_2),.clk(gclk));
	jdff dff_B_2kZfCFYy1_2(.din(w_dff_B_oQp4IJEg0_2),.dout(w_dff_B_2kZfCFYy1_2),.clk(gclk));
	jdff dff_B_PUckGBek7_2(.din(w_dff_B_2kZfCFYy1_2),.dout(w_dff_B_PUckGBek7_2),.clk(gclk));
	jdff dff_B_63oH4BDt9_2(.din(w_dff_B_PUckGBek7_2),.dout(w_dff_B_63oH4BDt9_2),.clk(gclk));
	jdff dff_B_7oxKpmbY9_2(.din(w_dff_B_63oH4BDt9_2),.dout(w_dff_B_7oxKpmbY9_2),.clk(gclk));
	jdff dff_B_baoqdbM52_2(.din(w_dff_B_7oxKpmbY9_2),.dout(w_dff_B_baoqdbM52_2),.clk(gclk));
	jdff dff_B_c2yjbTwH0_1(.din(n1566),.dout(w_dff_B_c2yjbTwH0_1),.clk(gclk));
	jdff dff_B_SlEBjpw15_1(.din(w_dff_B_c2yjbTwH0_1),.dout(w_dff_B_SlEBjpw15_1),.clk(gclk));
	jdff dff_B_x7ZnNhe53_2(.din(n1565),.dout(w_dff_B_x7ZnNhe53_2),.clk(gclk));
	jdff dff_B_8DnKZYTP2_2(.din(w_dff_B_x7ZnNhe53_2),.dout(w_dff_B_8DnKZYTP2_2),.clk(gclk));
	jdff dff_B_YkQjSEPa4_2(.din(w_dff_B_8DnKZYTP2_2),.dout(w_dff_B_YkQjSEPa4_2),.clk(gclk));
	jdff dff_B_SzWCiNbT8_2(.din(w_dff_B_YkQjSEPa4_2),.dout(w_dff_B_SzWCiNbT8_2),.clk(gclk));
	jdff dff_B_fN38XyAa7_2(.din(w_dff_B_SzWCiNbT8_2),.dout(w_dff_B_fN38XyAa7_2),.clk(gclk));
	jdff dff_B_q4503rNP6_2(.din(w_dff_B_fN38XyAa7_2),.dout(w_dff_B_q4503rNP6_2),.clk(gclk));
	jdff dff_B_gDkx0rSA9_2(.din(w_dff_B_q4503rNP6_2),.dout(w_dff_B_gDkx0rSA9_2),.clk(gclk));
	jdff dff_B_lsTORZFR4_2(.din(w_dff_B_gDkx0rSA9_2),.dout(w_dff_B_lsTORZFR4_2),.clk(gclk));
	jdff dff_B_eMvivkk69_2(.din(w_dff_B_lsTORZFR4_2),.dout(w_dff_B_eMvivkk69_2),.clk(gclk));
	jdff dff_B_2dOYPNCN6_2(.din(w_dff_B_eMvivkk69_2),.dout(w_dff_B_2dOYPNCN6_2),.clk(gclk));
	jdff dff_B_4lEFZheb6_2(.din(w_dff_B_2dOYPNCN6_2),.dout(w_dff_B_4lEFZheb6_2),.clk(gclk));
	jdff dff_B_z5VFRaH92_2(.din(w_dff_B_4lEFZheb6_2),.dout(w_dff_B_z5VFRaH92_2),.clk(gclk));
	jdff dff_B_Bhhd5Y0G9_2(.din(w_dff_B_z5VFRaH92_2),.dout(w_dff_B_Bhhd5Y0G9_2),.clk(gclk));
	jdff dff_B_pG3vB1Ii5_2(.din(w_dff_B_Bhhd5Y0G9_2),.dout(w_dff_B_pG3vB1Ii5_2),.clk(gclk));
	jdff dff_B_FqJ8Xvwo0_2(.din(w_dff_B_pG3vB1Ii5_2),.dout(w_dff_B_FqJ8Xvwo0_2),.clk(gclk));
	jdff dff_B_h1yJEpBM9_2(.din(w_dff_B_FqJ8Xvwo0_2),.dout(w_dff_B_h1yJEpBM9_2),.clk(gclk));
	jdff dff_B_A8eIH1ei6_2(.din(w_dff_B_h1yJEpBM9_2),.dout(w_dff_B_A8eIH1ei6_2),.clk(gclk));
	jdff dff_B_68fSbukW8_2(.din(w_dff_B_A8eIH1ei6_2),.dout(w_dff_B_68fSbukW8_2),.clk(gclk));
	jdff dff_B_gNwX56j45_2(.din(w_dff_B_68fSbukW8_2),.dout(w_dff_B_gNwX56j45_2),.clk(gclk));
	jdff dff_B_UNdv8N1s5_2(.din(w_dff_B_gNwX56j45_2),.dout(w_dff_B_UNdv8N1s5_2),.clk(gclk));
	jdff dff_B_ZI6kZ0CH1_2(.din(w_dff_B_UNdv8N1s5_2),.dout(w_dff_B_ZI6kZ0CH1_2),.clk(gclk));
	jdff dff_B_Xj80AD3f2_2(.din(w_dff_B_ZI6kZ0CH1_2),.dout(w_dff_B_Xj80AD3f2_2),.clk(gclk));
	jdff dff_B_ItotBtzo2_2(.din(w_dff_B_Xj80AD3f2_2),.dout(w_dff_B_ItotBtzo2_2),.clk(gclk));
	jdff dff_B_zeBcSGFn5_2(.din(w_dff_B_ItotBtzo2_2),.dout(w_dff_B_zeBcSGFn5_2),.clk(gclk));
	jdff dff_B_M96nUBHJ0_2(.din(w_dff_B_zeBcSGFn5_2),.dout(w_dff_B_M96nUBHJ0_2),.clk(gclk));
	jdff dff_B_aggZNkns5_2(.din(w_dff_B_M96nUBHJ0_2),.dout(w_dff_B_aggZNkns5_2),.clk(gclk));
	jdff dff_B_CwnYIZsQ2_2(.din(w_dff_B_aggZNkns5_2),.dout(w_dff_B_CwnYIZsQ2_2),.clk(gclk));
	jdff dff_B_cKmGXSGE9_2(.din(w_dff_B_CwnYIZsQ2_2),.dout(w_dff_B_cKmGXSGE9_2),.clk(gclk));
	jdff dff_B_BxO64W1V2_2(.din(w_dff_B_cKmGXSGE9_2),.dout(w_dff_B_BxO64W1V2_2),.clk(gclk));
	jdff dff_B_vtUutOwt3_2(.din(n1564),.dout(w_dff_B_vtUutOwt3_2),.clk(gclk));
	jdff dff_B_7sTMXM465_2(.din(w_dff_B_vtUutOwt3_2),.dout(w_dff_B_7sTMXM465_2),.clk(gclk));
	jdff dff_B_KKyuNzo66_2(.din(w_dff_B_7sTMXM465_2),.dout(w_dff_B_KKyuNzo66_2),.clk(gclk));
	jdff dff_B_DDkdSG1i2_2(.din(w_dff_B_KKyuNzo66_2),.dout(w_dff_B_DDkdSG1i2_2),.clk(gclk));
	jdff dff_B_mBhy0BFq7_2(.din(w_dff_B_DDkdSG1i2_2),.dout(w_dff_B_mBhy0BFq7_2),.clk(gclk));
	jdff dff_B_l7L0FhuG2_2(.din(w_dff_B_mBhy0BFq7_2),.dout(w_dff_B_l7L0FhuG2_2),.clk(gclk));
	jdff dff_B_u28Jy0qd1_2(.din(w_dff_B_l7L0FhuG2_2),.dout(w_dff_B_u28Jy0qd1_2),.clk(gclk));
	jdff dff_B_DRJyE8b40_2(.din(w_dff_B_u28Jy0qd1_2),.dout(w_dff_B_DRJyE8b40_2),.clk(gclk));
	jdff dff_B_JiYLPRuo6_2(.din(w_dff_B_DRJyE8b40_2),.dout(w_dff_B_JiYLPRuo6_2),.clk(gclk));
	jdff dff_B_5vuPtkq32_2(.din(w_dff_B_JiYLPRuo6_2),.dout(w_dff_B_5vuPtkq32_2),.clk(gclk));
	jdff dff_B_UdjggULq0_2(.din(w_dff_B_5vuPtkq32_2),.dout(w_dff_B_UdjggULq0_2),.clk(gclk));
	jdff dff_B_DNFsz12B0_2(.din(w_dff_B_UdjggULq0_2),.dout(w_dff_B_DNFsz12B0_2),.clk(gclk));
	jdff dff_B_ny3lv2Jd9_2(.din(w_dff_B_DNFsz12B0_2),.dout(w_dff_B_ny3lv2Jd9_2),.clk(gclk));
	jdff dff_B_hhnvwzLR4_2(.din(w_dff_B_ny3lv2Jd9_2),.dout(w_dff_B_hhnvwzLR4_2),.clk(gclk));
	jdff dff_B_gnsUch1D4_2(.din(w_dff_B_hhnvwzLR4_2),.dout(w_dff_B_gnsUch1D4_2),.clk(gclk));
	jdff dff_B_0f9njkGx2_2(.din(w_dff_B_gnsUch1D4_2),.dout(w_dff_B_0f9njkGx2_2),.clk(gclk));
	jdff dff_B_fDmKdxwM5_2(.din(w_dff_B_0f9njkGx2_2),.dout(w_dff_B_fDmKdxwM5_2),.clk(gclk));
	jdff dff_B_ELoFqzoL2_2(.din(w_dff_B_fDmKdxwM5_2),.dout(w_dff_B_ELoFqzoL2_2),.clk(gclk));
	jdff dff_B_hYN2DRpR5_2(.din(w_dff_B_ELoFqzoL2_2),.dout(w_dff_B_hYN2DRpR5_2),.clk(gclk));
	jdff dff_B_fEbKfBrj6_2(.din(w_dff_B_hYN2DRpR5_2),.dout(w_dff_B_fEbKfBrj6_2),.clk(gclk));
	jdff dff_B_98wTQw1G1_2(.din(w_dff_B_fEbKfBrj6_2),.dout(w_dff_B_98wTQw1G1_2),.clk(gclk));
	jdff dff_B_GBiiiZej1_2(.din(w_dff_B_98wTQw1G1_2),.dout(w_dff_B_GBiiiZej1_2),.clk(gclk));
	jdff dff_B_lnUtt5NM5_2(.din(w_dff_B_GBiiiZej1_2),.dout(w_dff_B_lnUtt5NM5_2),.clk(gclk));
	jdff dff_B_YNTsZpgP4_2(.din(w_dff_B_lnUtt5NM5_2),.dout(w_dff_B_YNTsZpgP4_2),.clk(gclk));
	jdff dff_B_UwOKQZCP9_2(.din(w_dff_B_YNTsZpgP4_2),.dout(w_dff_B_UwOKQZCP9_2),.clk(gclk));
	jdff dff_B_z27gR8kK1_2(.din(w_dff_B_UwOKQZCP9_2),.dout(w_dff_B_z27gR8kK1_2),.clk(gclk));
	jdff dff_B_LMPaQdI47_2(.din(w_dff_B_z27gR8kK1_2),.dout(w_dff_B_LMPaQdI47_2),.clk(gclk));
	jdff dff_B_tXTTbGDF2_2(.din(w_dff_B_LMPaQdI47_2),.dout(w_dff_B_tXTTbGDF2_2),.clk(gclk));
	jdff dff_B_YSqoSBQi6_2(.din(w_dff_B_tXTTbGDF2_2),.dout(w_dff_B_YSqoSBQi6_2),.clk(gclk));
	jdff dff_B_5TA3ku9h4_2(.din(w_dff_B_YSqoSBQi6_2),.dout(w_dff_B_5TA3ku9h4_2),.clk(gclk));
	jdff dff_B_oAJS2gxH9_2(.din(w_dff_B_5TA3ku9h4_2),.dout(w_dff_B_oAJS2gxH9_2),.clk(gclk));
	jdff dff_B_p4XeoJmg1_2(.din(n1563),.dout(w_dff_B_p4XeoJmg1_2),.clk(gclk));
	jdff dff_B_eAljtyPM9_1(.din(n1561),.dout(w_dff_B_eAljtyPM9_1),.clk(gclk));
	jdff dff_B_dcRyaz0x3_2(.din(n1496),.dout(w_dff_B_dcRyaz0x3_2),.clk(gclk));
	jdff dff_B_VfX6BxUF7_2(.din(w_dff_B_dcRyaz0x3_2),.dout(w_dff_B_VfX6BxUF7_2),.clk(gclk));
	jdff dff_B_innOVUcS8_2(.din(w_dff_B_VfX6BxUF7_2),.dout(w_dff_B_innOVUcS8_2),.clk(gclk));
	jdff dff_B_FaLf88IZ5_2(.din(w_dff_B_innOVUcS8_2),.dout(w_dff_B_FaLf88IZ5_2),.clk(gclk));
	jdff dff_B_edtbpbmp0_2(.din(w_dff_B_FaLf88IZ5_2),.dout(w_dff_B_edtbpbmp0_2),.clk(gclk));
	jdff dff_B_H6OjrtMF1_2(.din(w_dff_B_edtbpbmp0_2),.dout(w_dff_B_H6OjrtMF1_2),.clk(gclk));
	jdff dff_B_iTrgwVPV5_2(.din(w_dff_B_H6OjrtMF1_2),.dout(w_dff_B_iTrgwVPV5_2),.clk(gclk));
	jdff dff_B_S1rTYZ5R5_2(.din(w_dff_B_iTrgwVPV5_2),.dout(w_dff_B_S1rTYZ5R5_2),.clk(gclk));
	jdff dff_B_GqmIozHi6_2(.din(w_dff_B_S1rTYZ5R5_2),.dout(w_dff_B_GqmIozHi6_2),.clk(gclk));
	jdff dff_B_PICjZBWz6_2(.din(w_dff_B_GqmIozHi6_2),.dout(w_dff_B_PICjZBWz6_2),.clk(gclk));
	jdff dff_B_FlKleEVC8_2(.din(w_dff_B_PICjZBWz6_2),.dout(w_dff_B_FlKleEVC8_2),.clk(gclk));
	jdff dff_B_hDozs50r1_2(.din(w_dff_B_FlKleEVC8_2),.dout(w_dff_B_hDozs50r1_2),.clk(gclk));
	jdff dff_B_CNEgWOUT6_2(.din(w_dff_B_hDozs50r1_2),.dout(w_dff_B_CNEgWOUT6_2),.clk(gclk));
	jdff dff_B_Bn6sZ6mb0_2(.din(w_dff_B_CNEgWOUT6_2),.dout(w_dff_B_Bn6sZ6mb0_2),.clk(gclk));
	jdff dff_B_LYJCQMxE4_2(.din(w_dff_B_Bn6sZ6mb0_2),.dout(w_dff_B_LYJCQMxE4_2),.clk(gclk));
	jdff dff_B_wXJDgVuo0_2(.din(w_dff_B_LYJCQMxE4_2),.dout(w_dff_B_wXJDgVuo0_2),.clk(gclk));
	jdff dff_B_DZ0VPlyn8_2(.din(w_dff_B_wXJDgVuo0_2),.dout(w_dff_B_DZ0VPlyn8_2),.clk(gclk));
	jdff dff_B_FegmY1Od9_2(.din(w_dff_B_DZ0VPlyn8_2),.dout(w_dff_B_FegmY1Od9_2),.clk(gclk));
	jdff dff_B_qTyaly0q4_2(.din(w_dff_B_FegmY1Od9_2),.dout(w_dff_B_qTyaly0q4_2),.clk(gclk));
	jdff dff_B_cQKEC7547_2(.din(w_dff_B_qTyaly0q4_2),.dout(w_dff_B_cQKEC7547_2),.clk(gclk));
	jdff dff_B_uz5NnPzy5_2(.din(w_dff_B_cQKEC7547_2),.dout(w_dff_B_uz5NnPzy5_2),.clk(gclk));
	jdff dff_B_duFxJ8s00_2(.din(w_dff_B_uz5NnPzy5_2),.dout(w_dff_B_duFxJ8s00_2),.clk(gclk));
	jdff dff_B_SC7R0snO2_2(.din(w_dff_B_duFxJ8s00_2),.dout(w_dff_B_SC7R0snO2_2),.clk(gclk));
	jdff dff_B_91KWYDUn6_2(.din(w_dff_B_SC7R0snO2_2),.dout(w_dff_B_91KWYDUn6_2),.clk(gclk));
	jdff dff_B_lCxN2mNQ5_2(.din(w_dff_B_91KWYDUn6_2),.dout(w_dff_B_lCxN2mNQ5_2),.clk(gclk));
	jdff dff_B_AuWPTUae7_2(.din(w_dff_B_lCxN2mNQ5_2),.dout(w_dff_B_AuWPTUae7_2),.clk(gclk));
	jdff dff_B_77y9GENH0_2(.din(w_dff_B_AuWPTUae7_2),.dout(w_dff_B_77y9GENH0_2),.clk(gclk));
	jdff dff_B_3aHAWKT57_2(.din(w_dff_B_77y9GENH0_2),.dout(w_dff_B_3aHAWKT57_2),.clk(gclk));
	jdff dff_B_c3bULSld1_1(.din(n1502),.dout(w_dff_B_c3bULSld1_1),.clk(gclk));
	jdff dff_B_jkG7Gnh21_1(.din(w_dff_B_c3bULSld1_1),.dout(w_dff_B_jkG7Gnh21_1),.clk(gclk));
	jdff dff_B_3lm5RqDx4_2(.din(n1501),.dout(w_dff_B_3lm5RqDx4_2),.clk(gclk));
	jdff dff_B_ZmTez0jb0_2(.din(w_dff_B_3lm5RqDx4_2),.dout(w_dff_B_ZmTez0jb0_2),.clk(gclk));
	jdff dff_B_QHzUqkc97_2(.din(w_dff_B_ZmTez0jb0_2),.dout(w_dff_B_QHzUqkc97_2),.clk(gclk));
	jdff dff_B_6IBFZh2k8_2(.din(w_dff_B_QHzUqkc97_2),.dout(w_dff_B_6IBFZh2k8_2),.clk(gclk));
	jdff dff_B_AuJfrlsY4_2(.din(w_dff_B_6IBFZh2k8_2),.dout(w_dff_B_AuJfrlsY4_2),.clk(gclk));
	jdff dff_B_8mW2OEhD4_2(.din(w_dff_B_AuJfrlsY4_2),.dout(w_dff_B_8mW2OEhD4_2),.clk(gclk));
	jdff dff_B_DfMVywnC4_2(.din(w_dff_B_8mW2OEhD4_2),.dout(w_dff_B_DfMVywnC4_2),.clk(gclk));
	jdff dff_B_aOvUAm1s6_2(.din(w_dff_B_DfMVywnC4_2),.dout(w_dff_B_aOvUAm1s6_2),.clk(gclk));
	jdff dff_B_ekBohHdc3_2(.din(w_dff_B_aOvUAm1s6_2),.dout(w_dff_B_ekBohHdc3_2),.clk(gclk));
	jdff dff_B_M87LqWdH1_2(.din(w_dff_B_ekBohHdc3_2),.dout(w_dff_B_M87LqWdH1_2),.clk(gclk));
	jdff dff_B_JT8HwOxL6_2(.din(w_dff_B_M87LqWdH1_2),.dout(w_dff_B_JT8HwOxL6_2),.clk(gclk));
	jdff dff_B_A3UkykDj6_2(.din(w_dff_B_JT8HwOxL6_2),.dout(w_dff_B_A3UkykDj6_2),.clk(gclk));
	jdff dff_B_uNVEeAel7_2(.din(w_dff_B_A3UkykDj6_2),.dout(w_dff_B_uNVEeAel7_2),.clk(gclk));
	jdff dff_B_Phg1ej875_2(.din(w_dff_B_uNVEeAel7_2),.dout(w_dff_B_Phg1ej875_2),.clk(gclk));
	jdff dff_B_bkF9Tx1m0_2(.din(w_dff_B_Phg1ej875_2),.dout(w_dff_B_bkF9Tx1m0_2),.clk(gclk));
	jdff dff_B_FRuFpevk2_2(.din(w_dff_B_bkF9Tx1m0_2),.dout(w_dff_B_FRuFpevk2_2),.clk(gclk));
	jdff dff_B_9drKR0pB5_2(.din(w_dff_B_FRuFpevk2_2),.dout(w_dff_B_9drKR0pB5_2),.clk(gclk));
	jdff dff_B_OyvTpN4s8_2(.din(w_dff_B_9drKR0pB5_2),.dout(w_dff_B_OyvTpN4s8_2),.clk(gclk));
	jdff dff_B_AycQ6MKX1_2(.din(w_dff_B_OyvTpN4s8_2),.dout(w_dff_B_AycQ6MKX1_2),.clk(gclk));
	jdff dff_B_cR2o2IGY3_2(.din(w_dff_B_AycQ6MKX1_2),.dout(w_dff_B_cR2o2IGY3_2),.clk(gclk));
	jdff dff_B_pfK1Zg7E2_2(.din(w_dff_B_cR2o2IGY3_2),.dout(w_dff_B_pfK1Zg7E2_2),.clk(gclk));
	jdff dff_B_yFKj9PKM2_2(.din(w_dff_B_pfK1Zg7E2_2),.dout(w_dff_B_yFKj9PKM2_2),.clk(gclk));
	jdff dff_B_SHUOJgeh1_2(.din(w_dff_B_yFKj9PKM2_2),.dout(w_dff_B_SHUOJgeh1_2),.clk(gclk));
	jdff dff_B_CC0YeSiT7_2(.din(w_dff_B_SHUOJgeh1_2),.dout(w_dff_B_CC0YeSiT7_2),.clk(gclk));
	jdff dff_B_0ytc6keY6_2(.din(w_dff_B_CC0YeSiT7_2),.dout(w_dff_B_0ytc6keY6_2),.clk(gclk));
	jdff dff_B_kGcpJOVY7_2(.din(n1500),.dout(w_dff_B_kGcpJOVY7_2),.clk(gclk));
	jdff dff_B_J4JWlldT8_2(.din(w_dff_B_kGcpJOVY7_2),.dout(w_dff_B_J4JWlldT8_2),.clk(gclk));
	jdff dff_B_kObFjjDR0_2(.din(w_dff_B_J4JWlldT8_2),.dout(w_dff_B_kObFjjDR0_2),.clk(gclk));
	jdff dff_B_iED7qo193_2(.din(w_dff_B_kObFjjDR0_2),.dout(w_dff_B_iED7qo193_2),.clk(gclk));
	jdff dff_B_E8JasFAi5_2(.din(w_dff_B_iED7qo193_2),.dout(w_dff_B_E8JasFAi5_2),.clk(gclk));
	jdff dff_B_AvWwjkFq5_2(.din(w_dff_B_E8JasFAi5_2),.dout(w_dff_B_AvWwjkFq5_2),.clk(gclk));
	jdff dff_B_M2709WEX8_2(.din(w_dff_B_AvWwjkFq5_2),.dout(w_dff_B_M2709WEX8_2),.clk(gclk));
	jdff dff_B_BgXFYNdH3_2(.din(w_dff_B_M2709WEX8_2),.dout(w_dff_B_BgXFYNdH3_2),.clk(gclk));
	jdff dff_B_Op3T7d9G6_2(.din(w_dff_B_BgXFYNdH3_2),.dout(w_dff_B_Op3T7d9G6_2),.clk(gclk));
	jdff dff_B_GGjH24kH3_2(.din(w_dff_B_Op3T7d9G6_2),.dout(w_dff_B_GGjH24kH3_2),.clk(gclk));
	jdff dff_B_AJOeFvkt2_2(.din(w_dff_B_GGjH24kH3_2),.dout(w_dff_B_AJOeFvkt2_2),.clk(gclk));
	jdff dff_B_JDPIXf858_2(.din(w_dff_B_AJOeFvkt2_2),.dout(w_dff_B_JDPIXf858_2),.clk(gclk));
	jdff dff_B_RcXo07651_2(.din(w_dff_B_JDPIXf858_2),.dout(w_dff_B_RcXo07651_2),.clk(gclk));
	jdff dff_B_gasTXOml2_2(.din(w_dff_B_RcXo07651_2),.dout(w_dff_B_gasTXOml2_2),.clk(gclk));
	jdff dff_B_FMzdovn09_2(.din(w_dff_B_gasTXOml2_2),.dout(w_dff_B_FMzdovn09_2),.clk(gclk));
	jdff dff_B_7kEQqkeJ4_2(.din(w_dff_B_FMzdovn09_2),.dout(w_dff_B_7kEQqkeJ4_2),.clk(gclk));
	jdff dff_B_7Y8VCaGV4_2(.din(w_dff_B_7kEQqkeJ4_2),.dout(w_dff_B_7Y8VCaGV4_2),.clk(gclk));
	jdff dff_B_uZOvTSdZ3_2(.din(w_dff_B_7Y8VCaGV4_2),.dout(w_dff_B_uZOvTSdZ3_2),.clk(gclk));
	jdff dff_B_Q0GSHaYs1_2(.din(w_dff_B_uZOvTSdZ3_2),.dout(w_dff_B_Q0GSHaYs1_2),.clk(gclk));
	jdff dff_B_XAHFpnQC3_2(.din(w_dff_B_Q0GSHaYs1_2),.dout(w_dff_B_XAHFpnQC3_2),.clk(gclk));
	jdff dff_B_ROfSh6Eo9_2(.din(w_dff_B_XAHFpnQC3_2),.dout(w_dff_B_ROfSh6Eo9_2),.clk(gclk));
	jdff dff_B_HgsUEgEm5_2(.din(w_dff_B_ROfSh6Eo9_2),.dout(w_dff_B_HgsUEgEm5_2),.clk(gclk));
	jdff dff_B_DQXPQeFA6_2(.din(w_dff_B_HgsUEgEm5_2),.dout(w_dff_B_DQXPQeFA6_2),.clk(gclk));
	jdff dff_B_GZgteWl33_2(.din(w_dff_B_DQXPQeFA6_2),.dout(w_dff_B_GZgteWl33_2),.clk(gclk));
	jdff dff_B_MkF20I2O9_2(.din(w_dff_B_GZgteWl33_2),.dout(w_dff_B_MkF20I2O9_2),.clk(gclk));
	jdff dff_B_oDtEooSa4_2(.din(w_dff_B_MkF20I2O9_2),.dout(w_dff_B_oDtEooSa4_2),.clk(gclk));
	jdff dff_B_w3yWoLIG5_2(.din(w_dff_B_oDtEooSa4_2),.dout(w_dff_B_w3yWoLIG5_2),.clk(gclk));
	jdff dff_B_1ZVbO9WY8_2(.din(n1499),.dout(w_dff_B_1ZVbO9WY8_2),.clk(gclk));
	jdff dff_B_Qgbz1cZp2_1(.din(n1497),.dout(w_dff_B_Qgbz1cZp2_1),.clk(gclk));
	jdff dff_B_piQY7FD69_2(.din(n1425),.dout(w_dff_B_piQY7FD69_2),.clk(gclk));
	jdff dff_B_MjDz38Rb0_2(.din(w_dff_B_piQY7FD69_2),.dout(w_dff_B_MjDz38Rb0_2),.clk(gclk));
	jdff dff_B_NkNoymbq0_2(.din(w_dff_B_MjDz38Rb0_2),.dout(w_dff_B_NkNoymbq0_2),.clk(gclk));
	jdff dff_B_kbq4Q1ix0_2(.din(w_dff_B_NkNoymbq0_2),.dout(w_dff_B_kbq4Q1ix0_2),.clk(gclk));
	jdff dff_B_GsCu1Mc82_2(.din(w_dff_B_kbq4Q1ix0_2),.dout(w_dff_B_GsCu1Mc82_2),.clk(gclk));
	jdff dff_B_gsBRj3eu6_2(.din(w_dff_B_GsCu1Mc82_2),.dout(w_dff_B_gsBRj3eu6_2),.clk(gclk));
	jdff dff_B_GiL44ctW6_2(.din(w_dff_B_gsBRj3eu6_2),.dout(w_dff_B_GiL44ctW6_2),.clk(gclk));
	jdff dff_B_t4jjJZ4n9_2(.din(w_dff_B_GiL44ctW6_2),.dout(w_dff_B_t4jjJZ4n9_2),.clk(gclk));
	jdff dff_B_8AMbdcLi9_2(.din(w_dff_B_t4jjJZ4n9_2),.dout(w_dff_B_8AMbdcLi9_2),.clk(gclk));
	jdff dff_B_zuHQfkPo9_2(.din(w_dff_B_8AMbdcLi9_2),.dout(w_dff_B_zuHQfkPo9_2),.clk(gclk));
	jdff dff_B_2qWfIzGz7_2(.din(w_dff_B_zuHQfkPo9_2),.dout(w_dff_B_2qWfIzGz7_2),.clk(gclk));
	jdff dff_B_CdpdPQOS9_2(.din(w_dff_B_2qWfIzGz7_2),.dout(w_dff_B_CdpdPQOS9_2),.clk(gclk));
	jdff dff_B_2LbnHy5O1_2(.din(w_dff_B_CdpdPQOS9_2),.dout(w_dff_B_2LbnHy5O1_2),.clk(gclk));
	jdff dff_B_KejJAvHh6_2(.din(w_dff_B_2LbnHy5O1_2),.dout(w_dff_B_KejJAvHh6_2),.clk(gclk));
	jdff dff_B_SV2YQmhc9_2(.din(w_dff_B_KejJAvHh6_2),.dout(w_dff_B_SV2YQmhc9_2),.clk(gclk));
	jdff dff_B_N24Ub3J52_2(.din(w_dff_B_SV2YQmhc9_2),.dout(w_dff_B_N24Ub3J52_2),.clk(gclk));
	jdff dff_B_zVqUjW0n6_2(.din(w_dff_B_N24Ub3J52_2),.dout(w_dff_B_zVqUjW0n6_2),.clk(gclk));
	jdff dff_B_J71eQzl57_2(.din(w_dff_B_zVqUjW0n6_2),.dout(w_dff_B_J71eQzl57_2),.clk(gclk));
	jdff dff_B_HZDIJFTy6_2(.din(w_dff_B_J71eQzl57_2),.dout(w_dff_B_HZDIJFTy6_2),.clk(gclk));
	jdff dff_B_po3Xfo5O2_2(.din(w_dff_B_HZDIJFTy6_2),.dout(w_dff_B_po3Xfo5O2_2),.clk(gclk));
	jdff dff_B_um4wzFQ99_2(.din(w_dff_B_po3Xfo5O2_2),.dout(w_dff_B_um4wzFQ99_2),.clk(gclk));
	jdff dff_B_CWHlLOav1_2(.din(w_dff_B_um4wzFQ99_2),.dout(w_dff_B_CWHlLOav1_2),.clk(gclk));
	jdff dff_B_95dXR3pb1_2(.din(w_dff_B_CWHlLOav1_2),.dout(w_dff_B_95dXR3pb1_2),.clk(gclk));
	jdff dff_B_EzliOta12_2(.din(w_dff_B_95dXR3pb1_2),.dout(w_dff_B_EzliOta12_2),.clk(gclk));
	jdff dff_B_OiPdZfzd9_1(.din(n1431),.dout(w_dff_B_OiPdZfzd9_1),.clk(gclk));
	jdff dff_B_WWR6ioqC4_1(.din(w_dff_B_OiPdZfzd9_1),.dout(w_dff_B_WWR6ioqC4_1),.clk(gclk));
	jdff dff_B_doWhhhXj9_2(.din(n1430),.dout(w_dff_B_doWhhhXj9_2),.clk(gclk));
	jdff dff_B_NymjAeOs9_2(.din(w_dff_B_doWhhhXj9_2),.dout(w_dff_B_NymjAeOs9_2),.clk(gclk));
	jdff dff_B_lXDpwh3A1_2(.din(w_dff_B_NymjAeOs9_2),.dout(w_dff_B_lXDpwh3A1_2),.clk(gclk));
	jdff dff_B_ER9wpk1s2_2(.din(w_dff_B_lXDpwh3A1_2),.dout(w_dff_B_ER9wpk1s2_2),.clk(gclk));
	jdff dff_B_580gmNBR1_2(.din(w_dff_B_ER9wpk1s2_2),.dout(w_dff_B_580gmNBR1_2),.clk(gclk));
	jdff dff_B_5XsftpV22_2(.din(w_dff_B_580gmNBR1_2),.dout(w_dff_B_5XsftpV22_2),.clk(gclk));
	jdff dff_B_DqEmxztK3_2(.din(w_dff_B_5XsftpV22_2),.dout(w_dff_B_DqEmxztK3_2),.clk(gclk));
	jdff dff_B_fiR0a2pm3_2(.din(w_dff_B_DqEmxztK3_2),.dout(w_dff_B_fiR0a2pm3_2),.clk(gclk));
	jdff dff_B_EGmb7ZUH8_2(.din(w_dff_B_fiR0a2pm3_2),.dout(w_dff_B_EGmb7ZUH8_2),.clk(gclk));
	jdff dff_B_qKlxcxXJ3_2(.din(w_dff_B_EGmb7ZUH8_2),.dout(w_dff_B_qKlxcxXJ3_2),.clk(gclk));
	jdff dff_B_ArxJjXMQ5_2(.din(w_dff_B_qKlxcxXJ3_2),.dout(w_dff_B_ArxJjXMQ5_2),.clk(gclk));
	jdff dff_B_ZjEzips51_2(.din(w_dff_B_ArxJjXMQ5_2),.dout(w_dff_B_ZjEzips51_2),.clk(gclk));
	jdff dff_B_pwy0Ktlq6_2(.din(w_dff_B_ZjEzips51_2),.dout(w_dff_B_pwy0Ktlq6_2),.clk(gclk));
	jdff dff_B_gzqJSMd32_2(.din(w_dff_B_pwy0Ktlq6_2),.dout(w_dff_B_gzqJSMd32_2),.clk(gclk));
	jdff dff_B_gipH3PPL1_2(.din(w_dff_B_gzqJSMd32_2),.dout(w_dff_B_gipH3PPL1_2),.clk(gclk));
	jdff dff_B_hogzUncN2_2(.din(w_dff_B_gipH3PPL1_2),.dout(w_dff_B_hogzUncN2_2),.clk(gclk));
	jdff dff_B_42pL21Zb0_2(.din(w_dff_B_hogzUncN2_2),.dout(w_dff_B_42pL21Zb0_2),.clk(gclk));
	jdff dff_B_utlxdGBp8_2(.din(w_dff_B_42pL21Zb0_2),.dout(w_dff_B_utlxdGBp8_2),.clk(gclk));
	jdff dff_B_ONUyUNkJ2_2(.din(w_dff_B_utlxdGBp8_2),.dout(w_dff_B_ONUyUNkJ2_2),.clk(gclk));
	jdff dff_B_hE1OpSM45_2(.din(w_dff_B_ONUyUNkJ2_2),.dout(w_dff_B_hE1OpSM45_2),.clk(gclk));
	jdff dff_B_S3RGNprc3_2(.din(w_dff_B_hE1OpSM45_2),.dout(w_dff_B_S3RGNprc3_2),.clk(gclk));
	jdff dff_B_8v4kmHIr0_2(.din(n1429),.dout(w_dff_B_8v4kmHIr0_2),.clk(gclk));
	jdff dff_B_oNAkpXc45_2(.din(w_dff_B_8v4kmHIr0_2),.dout(w_dff_B_oNAkpXc45_2),.clk(gclk));
	jdff dff_B_J3Fv31er0_2(.din(w_dff_B_oNAkpXc45_2),.dout(w_dff_B_J3Fv31er0_2),.clk(gclk));
	jdff dff_B_sy6vPOu41_2(.din(w_dff_B_J3Fv31er0_2),.dout(w_dff_B_sy6vPOu41_2),.clk(gclk));
	jdff dff_B_pexyw1il9_2(.din(w_dff_B_sy6vPOu41_2),.dout(w_dff_B_pexyw1il9_2),.clk(gclk));
	jdff dff_B_cQqQwQ7A9_2(.din(w_dff_B_pexyw1il9_2),.dout(w_dff_B_cQqQwQ7A9_2),.clk(gclk));
	jdff dff_B_fKPmDFBN9_2(.din(w_dff_B_cQqQwQ7A9_2),.dout(w_dff_B_fKPmDFBN9_2),.clk(gclk));
	jdff dff_B_UuNmlEi89_2(.din(w_dff_B_fKPmDFBN9_2),.dout(w_dff_B_UuNmlEi89_2),.clk(gclk));
	jdff dff_B_GWOzs5ni6_2(.din(w_dff_B_UuNmlEi89_2),.dout(w_dff_B_GWOzs5ni6_2),.clk(gclk));
	jdff dff_B_piPFD9aN1_2(.din(w_dff_B_GWOzs5ni6_2),.dout(w_dff_B_piPFD9aN1_2),.clk(gclk));
	jdff dff_B_1Ph9KQoK7_2(.din(w_dff_B_piPFD9aN1_2),.dout(w_dff_B_1Ph9KQoK7_2),.clk(gclk));
	jdff dff_B_3nFcw1C58_2(.din(w_dff_B_1Ph9KQoK7_2),.dout(w_dff_B_3nFcw1C58_2),.clk(gclk));
	jdff dff_B_1t08g69X5_2(.din(w_dff_B_3nFcw1C58_2),.dout(w_dff_B_1t08g69X5_2),.clk(gclk));
	jdff dff_B_ncdylhJS9_2(.din(w_dff_B_1t08g69X5_2),.dout(w_dff_B_ncdylhJS9_2),.clk(gclk));
	jdff dff_B_VgY1Hdjs5_2(.din(w_dff_B_ncdylhJS9_2),.dout(w_dff_B_VgY1Hdjs5_2),.clk(gclk));
	jdff dff_B_rPA5s7yn8_2(.din(w_dff_B_VgY1Hdjs5_2),.dout(w_dff_B_rPA5s7yn8_2),.clk(gclk));
	jdff dff_B_VjpRjuk45_2(.din(w_dff_B_rPA5s7yn8_2),.dout(w_dff_B_VjpRjuk45_2),.clk(gclk));
	jdff dff_B_xasKGlYQ8_2(.din(w_dff_B_VjpRjuk45_2),.dout(w_dff_B_xasKGlYQ8_2),.clk(gclk));
	jdff dff_B_felqBjNZ5_2(.din(w_dff_B_xasKGlYQ8_2),.dout(w_dff_B_felqBjNZ5_2),.clk(gclk));
	jdff dff_B_ZPYw7DlJ2_2(.din(w_dff_B_felqBjNZ5_2),.dout(w_dff_B_ZPYw7DlJ2_2),.clk(gclk));
	jdff dff_B_UV0Eixpq8_2(.din(w_dff_B_ZPYw7DlJ2_2),.dout(w_dff_B_UV0Eixpq8_2),.clk(gclk));
	jdff dff_B_HPnERQSg0_2(.din(w_dff_B_UV0Eixpq8_2),.dout(w_dff_B_HPnERQSg0_2),.clk(gclk));
	jdff dff_B_P5aKcMzV6_2(.din(w_dff_B_HPnERQSg0_2),.dout(w_dff_B_P5aKcMzV6_2),.clk(gclk));
	jdff dff_B_obud84Fq6_2(.din(n1428),.dout(w_dff_B_obud84Fq6_2),.clk(gclk));
	jdff dff_B_xvrIb0mS9_1(.din(n1426),.dout(w_dff_B_xvrIb0mS9_1),.clk(gclk));
	jdff dff_B_UZP12VuM1_2(.din(n1347),.dout(w_dff_B_UZP12VuM1_2),.clk(gclk));
	jdff dff_B_X46FJYec7_2(.din(w_dff_B_UZP12VuM1_2),.dout(w_dff_B_X46FJYec7_2),.clk(gclk));
	jdff dff_B_hpqdlP1B8_2(.din(w_dff_B_X46FJYec7_2),.dout(w_dff_B_hpqdlP1B8_2),.clk(gclk));
	jdff dff_B_8oI7eOp77_2(.din(w_dff_B_hpqdlP1B8_2),.dout(w_dff_B_8oI7eOp77_2),.clk(gclk));
	jdff dff_B_o6bquFzt8_2(.din(w_dff_B_8oI7eOp77_2),.dout(w_dff_B_o6bquFzt8_2),.clk(gclk));
	jdff dff_B_ckWZdXUX0_2(.din(w_dff_B_o6bquFzt8_2),.dout(w_dff_B_ckWZdXUX0_2),.clk(gclk));
	jdff dff_B_5azc3tdZ1_2(.din(w_dff_B_ckWZdXUX0_2),.dout(w_dff_B_5azc3tdZ1_2),.clk(gclk));
	jdff dff_B_Dq587cjY0_2(.din(w_dff_B_5azc3tdZ1_2),.dout(w_dff_B_Dq587cjY0_2),.clk(gclk));
	jdff dff_B_WYhCNK918_2(.din(w_dff_B_Dq587cjY0_2),.dout(w_dff_B_WYhCNK918_2),.clk(gclk));
	jdff dff_B_OCoodkJc4_2(.din(w_dff_B_WYhCNK918_2),.dout(w_dff_B_OCoodkJc4_2),.clk(gclk));
	jdff dff_B_UI7bWbGz9_2(.din(w_dff_B_OCoodkJc4_2),.dout(w_dff_B_UI7bWbGz9_2),.clk(gclk));
	jdff dff_B_bGvhDLWC7_2(.din(w_dff_B_UI7bWbGz9_2),.dout(w_dff_B_bGvhDLWC7_2),.clk(gclk));
	jdff dff_B_RhCtjxKE0_2(.din(w_dff_B_bGvhDLWC7_2),.dout(w_dff_B_RhCtjxKE0_2),.clk(gclk));
	jdff dff_B_KvpPmaY98_2(.din(w_dff_B_RhCtjxKE0_2),.dout(w_dff_B_KvpPmaY98_2),.clk(gclk));
	jdff dff_B_wof6xHnK4_2(.din(w_dff_B_KvpPmaY98_2),.dout(w_dff_B_wof6xHnK4_2),.clk(gclk));
	jdff dff_B_LKRcOnkX0_2(.din(w_dff_B_wof6xHnK4_2),.dout(w_dff_B_LKRcOnkX0_2),.clk(gclk));
	jdff dff_B_op1iX8rY0_2(.din(w_dff_B_LKRcOnkX0_2),.dout(w_dff_B_op1iX8rY0_2),.clk(gclk));
	jdff dff_B_OW6n44te8_2(.din(w_dff_B_op1iX8rY0_2),.dout(w_dff_B_OW6n44te8_2),.clk(gclk));
	jdff dff_B_rpq5eHw38_2(.din(w_dff_B_OW6n44te8_2),.dout(w_dff_B_rpq5eHw38_2),.clk(gclk));
	jdff dff_B_sIGu0EXt3_2(.din(w_dff_B_rpq5eHw38_2),.dout(w_dff_B_sIGu0EXt3_2),.clk(gclk));
	jdff dff_B_Rauj33Hx7_1(.din(n1353),.dout(w_dff_B_Rauj33Hx7_1),.clk(gclk));
	jdff dff_B_qLfpP2yC6_1(.din(w_dff_B_Rauj33Hx7_1),.dout(w_dff_B_qLfpP2yC6_1),.clk(gclk));
	jdff dff_B_ieZrxodV4_2(.din(n1352),.dout(w_dff_B_ieZrxodV4_2),.clk(gclk));
	jdff dff_B_h12KJgud2_2(.din(w_dff_B_ieZrxodV4_2),.dout(w_dff_B_h12KJgud2_2),.clk(gclk));
	jdff dff_B_c8XFa7nk8_2(.din(w_dff_B_h12KJgud2_2),.dout(w_dff_B_c8XFa7nk8_2),.clk(gclk));
	jdff dff_B_DCEYz4Lr7_2(.din(w_dff_B_c8XFa7nk8_2),.dout(w_dff_B_DCEYz4Lr7_2),.clk(gclk));
	jdff dff_B_BtuclDl46_2(.din(w_dff_B_DCEYz4Lr7_2),.dout(w_dff_B_BtuclDl46_2),.clk(gclk));
	jdff dff_B_NOJpTwrO2_2(.din(w_dff_B_BtuclDl46_2),.dout(w_dff_B_NOJpTwrO2_2),.clk(gclk));
	jdff dff_B_Fe9Tkhlu7_2(.din(w_dff_B_NOJpTwrO2_2),.dout(w_dff_B_Fe9Tkhlu7_2),.clk(gclk));
	jdff dff_B_o8BBL3m74_2(.din(w_dff_B_Fe9Tkhlu7_2),.dout(w_dff_B_o8BBL3m74_2),.clk(gclk));
	jdff dff_B_FFEWbkTz0_2(.din(w_dff_B_o8BBL3m74_2),.dout(w_dff_B_FFEWbkTz0_2),.clk(gclk));
	jdff dff_B_FNwXay5i3_2(.din(w_dff_B_FFEWbkTz0_2),.dout(w_dff_B_FNwXay5i3_2),.clk(gclk));
	jdff dff_B_Tt7NSMvs7_2(.din(w_dff_B_FNwXay5i3_2),.dout(w_dff_B_Tt7NSMvs7_2),.clk(gclk));
	jdff dff_B_snCwN42f3_2(.din(w_dff_B_Tt7NSMvs7_2),.dout(w_dff_B_snCwN42f3_2),.clk(gclk));
	jdff dff_B_FZ8SdgGh0_2(.din(w_dff_B_snCwN42f3_2),.dout(w_dff_B_FZ8SdgGh0_2),.clk(gclk));
	jdff dff_B_APAPQfSQ3_2(.din(w_dff_B_FZ8SdgGh0_2),.dout(w_dff_B_APAPQfSQ3_2),.clk(gclk));
	jdff dff_B_3QZVNOAL8_2(.din(w_dff_B_APAPQfSQ3_2),.dout(w_dff_B_3QZVNOAL8_2),.clk(gclk));
	jdff dff_B_2JQWDic04_2(.din(w_dff_B_3QZVNOAL8_2),.dout(w_dff_B_2JQWDic04_2),.clk(gclk));
	jdff dff_B_FySL7aDB0_2(.din(w_dff_B_2JQWDic04_2),.dout(w_dff_B_FySL7aDB0_2),.clk(gclk));
	jdff dff_B_Z8bmcoua3_2(.din(n1351),.dout(w_dff_B_Z8bmcoua3_2),.clk(gclk));
	jdff dff_B_81FDSwIW1_2(.din(w_dff_B_Z8bmcoua3_2),.dout(w_dff_B_81FDSwIW1_2),.clk(gclk));
	jdff dff_B_lWxB88oV9_2(.din(w_dff_B_81FDSwIW1_2),.dout(w_dff_B_lWxB88oV9_2),.clk(gclk));
	jdff dff_B_WGblt9En9_2(.din(w_dff_B_lWxB88oV9_2),.dout(w_dff_B_WGblt9En9_2),.clk(gclk));
	jdff dff_B_xPNbKXED9_2(.din(w_dff_B_WGblt9En9_2),.dout(w_dff_B_xPNbKXED9_2),.clk(gclk));
	jdff dff_B_lLgwbKra1_2(.din(w_dff_B_xPNbKXED9_2),.dout(w_dff_B_lLgwbKra1_2),.clk(gclk));
	jdff dff_B_CkXWAS8q2_2(.din(w_dff_B_lLgwbKra1_2),.dout(w_dff_B_CkXWAS8q2_2),.clk(gclk));
	jdff dff_B_PywBbwpA8_2(.din(w_dff_B_CkXWAS8q2_2),.dout(w_dff_B_PywBbwpA8_2),.clk(gclk));
	jdff dff_B_b4YVCQlx5_2(.din(w_dff_B_PywBbwpA8_2),.dout(w_dff_B_b4YVCQlx5_2),.clk(gclk));
	jdff dff_B_QhXkmSDI0_2(.din(w_dff_B_b4YVCQlx5_2),.dout(w_dff_B_QhXkmSDI0_2),.clk(gclk));
	jdff dff_B_siap2Erl7_2(.din(w_dff_B_QhXkmSDI0_2),.dout(w_dff_B_siap2Erl7_2),.clk(gclk));
	jdff dff_B_ZDgohWOT2_2(.din(w_dff_B_siap2Erl7_2),.dout(w_dff_B_ZDgohWOT2_2),.clk(gclk));
	jdff dff_B_7DeUiXoB2_2(.din(w_dff_B_ZDgohWOT2_2),.dout(w_dff_B_7DeUiXoB2_2),.clk(gclk));
	jdff dff_B_kIZfLlmz3_2(.din(w_dff_B_7DeUiXoB2_2),.dout(w_dff_B_kIZfLlmz3_2),.clk(gclk));
	jdff dff_B_imIW2sWm4_2(.din(w_dff_B_kIZfLlmz3_2),.dout(w_dff_B_imIW2sWm4_2),.clk(gclk));
	jdff dff_B_MFs6FmlM3_2(.din(w_dff_B_imIW2sWm4_2),.dout(w_dff_B_MFs6FmlM3_2),.clk(gclk));
	jdff dff_B_X1CLj5ET8_2(.din(w_dff_B_MFs6FmlM3_2),.dout(w_dff_B_X1CLj5ET8_2),.clk(gclk));
	jdff dff_B_sOSGaqFI5_2(.din(w_dff_B_X1CLj5ET8_2),.dout(w_dff_B_sOSGaqFI5_2),.clk(gclk));
	jdff dff_B_4OFR99W31_2(.din(w_dff_B_sOSGaqFI5_2),.dout(w_dff_B_4OFR99W31_2),.clk(gclk));
	jdff dff_B_fF22xHZ72_1(.din(n1348),.dout(w_dff_B_fF22xHZ72_1),.clk(gclk));
	jdff dff_B_LpHrC3td5_2(.din(n1262),.dout(w_dff_B_LpHrC3td5_2),.clk(gclk));
	jdff dff_B_3bRU1I8S0_2(.din(w_dff_B_LpHrC3td5_2),.dout(w_dff_B_3bRU1I8S0_2),.clk(gclk));
	jdff dff_B_mHldo0tM9_2(.din(w_dff_B_3bRU1I8S0_2),.dout(w_dff_B_mHldo0tM9_2),.clk(gclk));
	jdff dff_B_OT2uoaZ40_2(.din(w_dff_B_mHldo0tM9_2),.dout(w_dff_B_OT2uoaZ40_2),.clk(gclk));
	jdff dff_B_doxB9s1K8_2(.din(w_dff_B_OT2uoaZ40_2),.dout(w_dff_B_doxB9s1K8_2),.clk(gclk));
	jdff dff_B_Oalguq2R5_2(.din(w_dff_B_doxB9s1K8_2),.dout(w_dff_B_Oalguq2R5_2),.clk(gclk));
	jdff dff_B_rsqeRcUk3_2(.din(w_dff_B_Oalguq2R5_2),.dout(w_dff_B_rsqeRcUk3_2),.clk(gclk));
	jdff dff_B_WcySLL2d2_2(.din(w_dff_B_rsqeRcUk3_2),.dout(w_dff_B_WcySLL2d2_2),.clk(gclk));
	jdff dff_B_rRChLAt44_2(.din(w_dff_B_WcySLL2d2_2),.dout(w_dff_B_rRChLAt44_2),.clk(gclk));
	jdff dff_B_5oOxccy72_2(.din(w_dff_B_rRChLAt44_2),.dout(w_dff_B_5oOxccy72_2),.clk(gclk));
	jdff dff_B_A6Q4mzqB0_2(.din(w_dff_B_5oOxccy72_2),.dout(w_dff_B_A6Q4mzqB0_2),.clk(gclk));
	jdff dff_B_qLh1rJOC9_2(.din(w_dff_B_A6Q4mzqB0_2),.dout(w_dff_B_qLh1rJOC9_2),.clk(gclk));
	jdff dff_B_5TeLkKGR2_2(.din(w_dff_B_qLh1rJOC9_2),.dout(w_dff_B_5TeLkKGR2_2),.clk(gclk));
	jdff dff_B_EMvmhfn53_2(.din(w_dff_B_5TeLkKGR2_2),.dout(w_dff_B_EMvmhfn53_2),.clk(gclk));
	jdff dff_B_h8AWiYyk6_2(.din(w_dff_B_EMvmhfn53_2),.dout(w_dff_B_h8AWiYyk6_2),.clk(gclk));
	jdff dff_B_5D5Qzu784_2(.din(w_dff_B_h8AWiYyk6_2),.dout(w_dff_B_5D5Qzu784_2),.clk(gclk));
	jdff dff_B_mp4WhI0R0_2(.din(w_dff_B_5D5Qzu784_2),.dout(w_dff_B_mp4WhI0R0_2),.clk(gclk));
	jdff dff_B_4RzogzYx1_2(.din(n1273),.dout(w_dff_B_4RzogzYx1_2),.clk(gclk));
	jdff dff_B_YfxulAEM9_1(.din(n1268),.dout(w_dff_B_YfxulAEM9_1),.clk(gclk));
	jdff dff_B_DY66GdNE4_1(.din(w_dff_B_YfxulAEM9_1),.dout(w_dff_B_DY66GdNE4_1),.clk(gclk));
	jdff dff_B_6YIX5qiW0_2(.din(n1267),.dout(w_dff_B_6YIX5qiW0_2),.clk(gclk));
	jdff dff_B_cFZ7vhnJ3_2(.din(w_dff_B_6YIX5qiW0_2),.dout(w_dff_B_cFZ7vhnJ3_2),.clk(gclk));
	jdff dff_B_LvMbsXMz4_2(.din(w_dff_B_cFZ7vhnJ3_2),.dout(w_dff_B_LvMbsXMz4_2),.clk(gclk));
	jdff dff_B_0afRMXRA5_2(.din(w_dff_B_LvMbsXMz4_2),.dout(w_dff_B_0afRMXRA5_2),.clk(gclk));
	jdff dff_B_YbhA4pNj6_2(.din(w_dff_B_0afRMXRA5_2),.dout(w_dff_B_YbhA4pNj6_2),.clk(gclk));
	jdff dff_B_PkWTiQfA4_2(.din(w_dff_B_YbhA4pNj6_2),.dout(w_dff_B_PkWTiQfA4_2),.clk(gclk));
	jdff dff_B_xOupLYoq8_2(.din(w_dff_B_PkWTiQfA4_2),.dout(w_dff_B_xOupLYoq8_2),.clk(gclk));
	jdff dff_B_uKeiKftv8_2(.din(w_dff_B_xOupLYoq8_2),.dout(w_dff_B_uKeiKftv8_2),.clk(gclk));
	jdff dff_B_9vJRf5FY2_2(.din(w_dff_B_uKeiKftv8_2),.dout(w_dff_B_9vJRf5FY2_2),.clk(gclk));
	jdff dff_B_HXqP3gBQ3_2(.din(w_dff_B_9vJRf5FY2_2),.dout(w_dff_B_HXqP3gBQ3_2),.clk(gclk));
	jdff dff_B_EorAVzXZ9_2(.din(w_dff_B_HXqP3gBQ3_2),.dout(w_dff_B_EorAVzXZ9_2),.clk(gclk));
	jdff dff_B_oivbJ5lx0_2(.din(w_dff_B_EorAVzXZ9_2),.dout(w_dff_B_oivbJ5lx0_2),.clk(gclk));
	jdff dff_B_1tzjXXiY8_2(.din(w_dff_B_oivbJ5lx0_2),.dout(w_dff_B_1tzjXXiY8_2),.clk(gclk));
	jdff dff_B_IIVSuTXM6_2(.din(n1266),.dout(w_dff_B_IIVSuTXM6_2),.clk(gclk));
	jdff dff_B_qzKKlDqP2_2(.din(w_dff_B_IIVSuTXM6_2),.dout(w_dff_B_qzKKlDqP2_2),.clk(gclk));
	jdff dff_B_Qh1da2da3_2(.din(w_dff_B_qzKKlDqP2_2),.dout(w_dff_B_Qh1da2da3_2),.clk(gclk));
	jdff dff_B_6e6bukUb7_2(.din(w_dff_B_Qh1da2da3_2),.dout(w_dff_B_6e6bukUb7_2),.clk(gclk));
	jdff dff_B_JzfdNGzG1_2(.din(w_dff_B_6e6bukUb7_2),.dout(w_dff_B_JzfdNGzG1_2),.clk(gclk));
	jdff dff_B_XUaFS7bj0_2(.din(w_dff_B_JzfdNGzG1_2),.dout(w_dff_B_XUaFS7bj0_2),.clk(gclk));
	jdff dff_B_v4Nt48gh8_2(.din(w_dff_B_XUaFS7bj0_2),.dout(w_dff_B_v4Nt48gh8_2),.clk(gclk));
	jdff dff_B_jd1pvwFq1_2(.din(w_dff_B_v4Nt48gh8_2),.dout(w_dff_B_jd1pvwFq1_2),.clk(gclk));
	jdff dff_B_jHy9EOol7_2(.din(w_dff_B_jd1pvwFq1_2),.dout(w_dff_B_jHy9EOol7_2),.clk(gclk));
	jdff dff_B_gH8pRmX97_2(.din(w_dff_B_jHy9EOol7_2),.dout(w_dff_B_gH8pRmX97_2),.clk(gclk));
	jdff dff_B_LfQ2JeJl7_2(.din(w_dff_B_gH8pRmX97_2),.dout(w_dff_B_LfQ2JeJl7_2),.clk(gclk));
	jdff dff_B_x8VQxSHb2_2(.din(w_dff_B_LfQ2JeJl7_2),.dout(w_dff_B_x8VQxSHb2_2),.clk(gclk));
	jdff dff_B_8uHJxpYY7_2(.din(w_dff_B_x8VQxSHb2_2),.dout(w_dff_B_8uHJxpYY7_2),.clk(gclk));
	jdff dff_B_5YJDHX9f4_2(.din(w_dff_B_8uHJxpYY7_2),.dout(w_dff_B_5YJDHX9f4_2),.clk(gclk));
	jdff dff_B_wCNWPAxc6_2(.din(w_dff_B_5YJDHX9f4_2),.dout(w_dff_B_wCNWPAxc6_2),.clk(gclk));
	jdff dff_B_rMz0XjOQ0_1(.din(n1263),.dout(w_dff_B_rMz0XjOQ0_1),.clk(gclk));
	jdff dff_B_yh3oE8w74_2(.din(n1171),.dout(w_dff_B_yh3oE8w74_2),.clk(gclk));
	jdff dff_B_Kt4m0qyQ8_2(.din(w_dff_B_yh3oE8w74_2),.dout(w_dff_B_Kt4m0qyQ8_2),.clk(gclk));
	jdff dff_B_0tysaLwm9_2(.din(w_dff_B_Kt4m0qyQ8_2),.dout(w_dff_B_0tysaLwm9_2),.clk(gclk));
	jdff dff_B_soh2w2Vt2_2(.din(w_dff_B_0tysaLwm9_2),.dout(w_dff_B_soh2w2Vt2_2),.clk(gclk));
	jdff dff_B_vHZeM2a86_2(.din(w_dff_B_soh2w2Vt2_2),.dout(w_dff_B_vHZeM2a86_2),.clk(gclk));
	jdff dff_B_ZIxMueCJ2_2(.din(w_dff_B_vHZeM2a86_2),.dout(w_dff_B_ZIxMueCJ2_2),.clk(gclk));
	jdff dff_B_QHf1iKAe8_2(.din(w_dff_B_ZIxMueCJ2_2),.dout(w_dff_B_QHf1iKAe8_2),.clk(gclk));
	jdff dff_B_L6B3r8fA2_2(.din(w_dff_B_QHf1iKAe8_2),.dout(w_dff_B_L6B3r8fA2_2),.clk(gclk));
	jdff dff_B_7UNYeD0A0_2(.din(w_dff_B_L6B3r8fA2_2),.dout(w_dff_B_7UNYeD0A0_2),.clk(gclk));
	jdff dff_B_JiOSGKO16_2(.din(w_dff_B_7UNYeD0A0_2),.dout(w_dff_B_JiOSGKO16_2),.clk(gclk));
	jdff dff_B_n2uwMoUY0_2(.din(w_dff_B_JiOSGKO16_2),.dout(w_dff_B_n2uwMoUY0_2),.clk(gclk));
	jdff dff_B_tlkm3Xnl4_2(.din(w_dff_B_n2uwMoUY0_2),.dout(w_dff_B_tlkm3Xnl4_2),.clk(gclk));
	jdff dff_B_nXIyRATt2_2(.din(w_dff_B_tlkm3Xnl4_2),.dout(w_dff_B_nXIyRATt2_2),.clk(gclk));
	jdff dff_B_gsC6wqNH0_2(.din(w_dff_B_nXIyRATt2_2),.dout(w_dff_B_gsC6wqNH0_2),.clk(gclk));
	jdff dff_B_LUhwgJYf1_2(.din(n1182),.dout(w_dff_B_LUhwgJYf1_2),.clk(gclk));
	jdff dff_B_l1BIsj2K7_2(.din(w_dff_B_LUhwgJYf1_2),.dout(w_dff_B_l1BIsj2K7_2),.clk(gclk));
	jdff dff_B_FMMA80sR8_1(.din(n1177),.dout(w_dff_B_FMMA80sR8_1),.clk(gclk));
	jdff dff_B_T8VZlarh2_1(.din(w_dff_B_FMMA80sR8_1),.dout(w_dff_B_T8VZlarh2_1),.clk(gclk));
	jdff dff_B_sqZW4AaN1_2(.din(n1176),.dout(w_dff_B_sqZW4AaN1_2),.clk(gclk));
	jdff dff_B_mB61WCyw8_2(.din(w_dff_B_sqZW4AaN1_2),.dout(w_dff_B_mB61WCyw8_2),.clk(gclk));
	jdff dff_B_yG5hC4mr5_2(.din(w_dff_B_mB61WCyw8_2),.dout(w_dff_B_yG5hC4mr5_2),.clk(gclk));
	jdff dff_B_rAP4h9PY5_2(.din(w_dff_B_yG5hC4mr5_2),.dout(w_dff_B_rAP4h9PY5_2),.clk(gclk));
	jdff dff_B_iYdgua2v5_2(.din(w_dff_B_rAP4h9PY5_2),.dout(w_dff_B_iYdgua2v5_2),.clk(gclk));
	jdff dff_B_CHRacBht2_2(.din(w_dff_B_iYdgua2v5_2),.dout(w_dff_B_CHRacBht2_2),.clk(gclk));
	jdff dff_B_tcyb7Ah26_2(.din(w_dff_B_CHRacBht2_2),.dout(w_dff_B_tcyb7Ah26_2),.clk(gclk));
	jdff dff_B_NqSMCDDU1_2(.din(w_dff_B_tcyb7Ah26_2),.dout(w_dff_B_NqSMCDDU1_2),.clk(gclk));
	jdff dff_B_bHlhii1X8_2(.din(w_dff_B_NqSMCDDU1_2),.dout(w_dff_B_bHlhii1X8_2),.clk(gclk));
	jdff dff_B_tNYKdjia8_2(.din(n1175),.dout(w_dff_B_tNYKdjia8_2),.clk(gclk));
	jdff dff_B_lE9E1rrc1_2(.din(w_dff_B_tNYKdjia8_2),.dout(w_dff_B_lE9E1rrc1_2),.clk(gclk));
	jdff dff_B_40Gezdqh1_2(.din(w_dff_B_lE9E1rrc1_2),.dout(w_dff_B_40Gezdqh1_2),.clk(gclk));
	jdff dff_B_9Xzy9A743_2(.din(w_dff_B_40Gezdqh1_2),.dout(w_dff_B_9Xzy9A743_2),.clk(gclk));
	jdff dff_B_4Pdrrfuv6_2(.din(w_dff_B_9Xzy9A743_2),.dout(w_dff_B_4Pdrrfuv6_2),.clk(gclk));
	jdff dff_B_nKYygaBl3_2(.din(w_dff_B_4Pdrrfuv6_2),.dout(w_dff_B_nKYygaBl3_2),.clk(gclk));
	jdff dff_B_VgjF3Ddo0_2(.din(w_dff_B_nKYygaBl3_2),.dout(w_dff_B_VgjF3Ddo0_2),.clk(gclk));
	jdff dff_B_eNnSARLR1_2(.din(w_dff_B_VgjF3Ddo0_2),.dout(w_dff_B_eNnSARLR1_2),.clk(gclk));
	jdff dff_B_6JUHd4Uy0_2(.din(w_dff_B_eNnSARLR1_2),.dout(w_dff_B_6JUHd4Uy0_2),.clk(gclk));
	jdff dff_B_6EwDfvpH1_2(.din(w_dff_B_6JUHd4Uy0_2),.dout(w_dff_B_6EwDfvpH1_2),.clk(gclk));
	jdff dff_B_3iHvH29H0_2(.din(w_dff_B_6EwDfvpH1_2),.dout(w_dff_B_3iHvH29H0_2),.clk(gclk));
	jdff dff_B_EaFpkXqV1_1(.din(n1172),.dout(w_dff_B_EaFpkXqV1_1),.clk(gclk));
	jdff dff_B_Y00VNV5P6_2(.din(n1073),.dout(w_dff_B_Y00VNV5P6_2),.clk(gclk));
	jdff dff_B_tz2glaSP3_2(.din(w_dff_B_Y00VNV5P6_2),.dout(w_dff_B_tz2glaSP3_2),.clk(gclk));
	jdff dff_B_OljZJaSS9_2(.din(w_dff_B_tz2glaSP3_2),.dout(w_dff_B_OljZJaSS9_2),.clk(gclk));
	jdff dff_B_IbXrYaYB1_2(.din(w_dff_B_OljZJaSS9_2),.dout(w_dff_B_IbXrYaYB1_2),.clk(gclk));
	jdff dff_B_GWQHjMTX7_2(.din(w_dff_B_IbXrYaYB1_2),.dout(w_dff_B_GWQHjMTX7_2),.clk(gclk));
	jdff dff_B_hyat70PT0_2(.din(w_dff_B_GWQHjMTX7_2),.dout(w_dff_B_hyat70PT0_2),.clk(gclk));
	jdff dff_B_CSDHSm5r4_2(.din(w_dff_B_hyat70PT0_2),.dout(w_dff_B_CSDHSm5r4_2),.clk(gclk));
	jdff dff_B_ydb2yCIh5_2(.din(w_dff_B_CSDHSm5r4_2),.dout(w_dff_B_ydb2yCIh5_2),.clk(gclk));
	jdff dff_B_q3BEP2P83_2(.din(w_dff_B_ydb2yCIh5_2),.dout(w_dff_B_q3BEP2P83_2),.clk(gclk));
	jdff dff_B_ScIGnvEV2_2(.din(w_dff_B_q3BEP2P83_2),.dout(w_dff_B_ScIGnvEV2_2),.clk(gclk));
	jdff dff_B_vR19TmIW5_2(.din(w_dff_B_ScIGnvEV2_2),.dout(w_dff_B_vR19TmIW5_2),.clk(gclk));
	jdff dff_B_iLqcGY7d8_2(.din(n1083),.dout(w_dff_B_iLqcGY7d8_2),.clk(gclk));
	jdff dff_B_vTgByL8q6_2(.din(w_dff_B_iLqcGY7d8_2),.dout(w_dff_B_vTgByL8q6_2),.clk(gclk));
	jdff dff_B_QBuWzmQu0_2(.din(w_dff_B_vTgByL8q6_2),.dout(w_dff_B_QBuWzmQu0_2),.clk(gclk));
	jdff dff_B_NavRGwX05_2(.din(n1078),.dout(w_dff_B_NavRGwX05_2),.clk(gclk));
	jdff dff_B_4rgkupxz3_2(.din(w_dff_B_NavRGwX05_2),.dout(w_dff_B_4rgkupxz3_2),.clk(gclk));
	jdff dff_B_AgB7gdh96_2(.din(w_dff_B_4rgkupxz3_2),.dout(w_dff_B_AgB7gdh96_2),.clk(gclk));
	jdff dff_B_D0Rwz3jX7_2(.din(w_dff_B_AgB7gdh96_2),.dout(w_dff_B_D0Rwz3jX7_2),.clk(gclk));
	jdff dff_B_s8ukJ44q7_2(.din(w_dff_B_D0Rwz3jX7_2),.dout(w_dff_B_s8ukJ44q7_2),.clk(gclk));
	jdff dff_B_t1JgZ43E2_2(.din(n1077),.dout(w_dff_B_t1JgZ43E2_2),.clk(gclk));
	jdff dff_B_CGtPIEal5_2(.din(w_dff_B_t1JgZ43E2_2),.dout(w_dff_B_CGtPIEal5_2),.clk(gclk));
	jdff dff_B_zMlyabps6_2(.din(w_dff_B_CGtPIEal5_2),.dout(w_dff_B_zMlyabps6_2),.clk(gclk));
	jdff dff_B_YgOjHMXK5_2(.din(w_dff_B_zMlyabps6_2),.dout(w_dff_B_YgOjHMXK5_2),.clk(gclk));
	jdff dff_B_uAvbnW1L3_2(.din(w_dff_B_YgOjHMXK5_2),.dout(w_dff_B_uAvbnW1L3_2),.clk(gclk));
	jdff dff_B_9asOxlze8_2(.din(w_dff_B_uAvbnW1L3_2),.dout(w_dff_B_9asOxlze8_2),.clk(gclk));
	jdff dff_B_x50Fva0C5_2(.din(w_dff_B_9asOxlze8_2),.dout(w_dff_B_x50Fva0C5_2),.clk(gclk));
	jdff dff_B_U2eEKYyt1_1(.din(n1074),.dout(w_dff_B_U2eEKYyt1_1),.clk(gclk));
	jdff dff_B_B786o5QK3_2(.din(n974),.dout(w_dff_B_B786o5QK3_2),.clk(gclk));
	jdff dff_B_PnWj6IOu5_2(.din(w_dff_B_B786o5QK3_2),.dout(w_dff_B_PnWj6IOu5_2),.clk(gclk));
	jdff dff_B_y1XSpmK04_2(.din(w_dff_B_PnWj6IOu5_2),.dout(w_dff_B_y1XSpmK04_2),.clk(gclk));
	jdff dff_B_enB6kYnQ0_2(.din(w_dff_B_y1XSpmK04_2),.dout(w_dff_B_enB6kYnQ0_2),.clk(gclk));
	jdff dff_B_XIqwfjWb0_2(.din(w_dff_B_enB6kYnQ0_2),.dout(w_dff_B_XIqwfjWb0_2),.clk(gclk));
	jdff dff_B_RgoM6Jzc8_2(.din(w_dff_B_XIqwfjWb0_2),.dout(w_dff_B_RgoM6Jzc8_2),.clk(gclk));
	jdff dff_B_6UsLvbar2_2(.din(w_dff_B_RgoM6Jzc8_2),.dout(w_dff_B_6UsLvbar2_2),.clk(gclk));
	jdff dff_B_c4z6oQvR5_2(.din(w_dff_B_6UsLvbar2_2),.dout(w_dff_B_c4z6oQvR5_2),.clk(gclk));
	jdff dff_B_1XvQhRLC2_2(.din(n984),.dout(w_dff_B_1XvQhRLC2_2),.clk(gclk));
	jdff dff_B_HnC3DcPT0_2(.din(w_dff_B_1XvQhRLC2_2),.dout(w_dff_B_HnC3DcPT0_2),.clk(gclk));
	jdff dff_B_P6yanSA50_2(.din(w_dff_B_HnC3DcPT0_2),.dout(w_dff_B_P6yanSA50_2),.clk(gclk));
	jdff dff_B_1PruDQuf8_2(.din(w_dff_B_P6yanSA50_2),.dout(w_dff_B_1PruDQuf8_2),.clk(gclk));
	jdff dff_B_lgtWnk074_2(.din(n983),.dout(w_dff_B_lgtWnk074_2),.clk(gclk));
	jdff dff_B_1aKC89GH2_2(.din(w_dff_B_lgtWnk074_2),.dout(w_dff_B_1aKC89GH2_2),.clk(gclk));
	jdff dff_B_gu26uhNi2_2(.din(w_dff_B_1aKC89GH2_2),.dout(w_dff_B_gu26uhNi2_2),.clk(gclk));
	jdff dff_A_hWGiBTey5_0(.dout(w_n980_0[0]),.din(w_dff_A_hWGiBTey5_0),.clk(gclk));
	jdff dff_A_j2iJF3dD4_0(.dout(w_dff_A_hWGiBTey5_0),.din(w_dff_A_j2iJF3dD4_0),.clk(gclk));
	jdff dff_A_cTYpb9Uc5_0(.dout(w_dff_A_j2iJF3dD4_0),.din(w_dff_A_cTYpb9Uc5_0),.clk(gclk));
	jdff dff_B_0eI2STGI0_2(.din(n980),.dout(w_dff_B_0eI2STGI0_2),.clk(gclk));
	jdff dff_A_Tj1mn60e8_0(.dout(w_n877_0[0]),.din(w_dff_A_Tj1mn60e8_0),.clk(gclk));
	jdff dff_A_CHYnw0Mb4_0(.dout(w_dff_A_Tj1mn60e8_0),.din(w_dff_A_CHYnw0Mb4_0),.clk(gclk));
	jdff dff_A_nVhSQM5i0_0(.dout(w_dff_A_CHYnw0Mb4_0),.din(w_dff_A_nVhSQM5i0_0),.clk(gclk));
	jdff dff_B_91FhsFt05_2(.din(n877),.dout(w_dff_B_91FhsFt05_2),.clk(gclk));
	jdff dff_A_GSJ5BpHw4_0(.dout(w_n875_0[0]),.din(w_dff_A_GSJ5BpHw4_0),.clk(gclk));
	jdff dff_A_U3lV2lY70_0(.dout(w_dff_A_GSJ5BpHw4_0),.din(w_dff_A_U3lV2lY70_0),.clk(gclk));
	jdff dff_B_yVRLDYHI0_2(.din(n874),.dout(w_dff_B_yVRLDYHI0_2),.clk(gclk));
	jdff dff_B_wglqkA0O8_2(.din(w_dff_B_yVRLDYHI0_2),.dout(w_dff_B_wglqkA0O8_2),.clk(gclk));
	jdff dff_B_sHzh34fk5_2(.din(w_dff_B_wglqkA0O8_2),.dout(w_dff_B_sHzh34fk5_2),.clk(gclk));
	jdff dff_A_Fe3KFXMD4_1(.dout(w_dff_A_spfPBIUn3_0),.din(w_dff_A_Fe3KFXMD4_1),.clk(gclk));
	jdff dff_A_spfPBIUn3_0(.dout(w_dff_A_95A7I1Kf9_0),.din(w_dff_A_spfPBIUn3_0),.clk(gclk));
	jdff dff_A_95A7I1Kf9_0(.dout(w_dff_A_EqG0Wzs46_0),.din(w_dff_A_95A7I1Kf9_0),.clk(gclk));
	jdff dff_A_EqG0Wzs46_0(.dout(w_dff_A_uPVtwYRJ4_0),.din(w_dff_A_EqG0Wzs46_0),.clk(gclk));
	jdff dff_A_uPVtwYRJ4_0(.dout(w_dff_A_C4CjRsh24_0),.din(w_dff_A_uPVtwYRJ4_0),.clk(gclk));
	jdff dff_A_C4CjRsh24_0(.dout(w_dff_A_V0en8nbW3_0),.din(w_dff_A_C4CjRsh24_0),.clk(gclk));
	jdff dff_A_V0en8nbW3_0(.dout(w_dff_A_ZjhSb9Oq4_0),.din(w_dff_A_V0en8nbW3_0),.clk(gclk));
	jdff dff_A_ZjhSb9Oq4_0(.dout(w_dff_A_EvJcgQzi7_0),.din(w_dff_A_ZjhSb9Oq4_0),.clk(gclk));
	jdff dff_A_EvJcgQzi7_0(.dout(w_dff_A_6HaGyRM36_0),.din(w_dff_A_EvJcgQzi7_0),.clk(gclk));
	jdff dff_A_6HaGyRM36_0(.dout(w_dff_A_gNoPZlNg0_0),.din(w_dff_A_6HaGyRM36_0),.clk(gclk));
	jdff dff_A_gNoPZlNg0_0(.dout(w_dff_A_cfH63hYN2_0),.din(w_dff_A_gNoPZlNg0_0),.clk(gclk));
	jdff dff_A_cfH63hYN2_0(.dout(w_dff_A_6D3v2Ycd2_0),.din(w_dff_A_cfH63hYN2_0),.clk(gclk));
	jdff dff_A_6D3v2Ycd2_0(.dout(w_dff_A_kgko3x4Q8_0),.din(w_dff_A_6D3v2Ycd2_0),.clk(gclk));
	jdff dff_A_kgko3x4Q8_0(.dout(w_dff_A_jDHW5v3Q0_0),.din(w_dff_A_kgko3x4Q8_0),.clk(gclk));
	jdff dff_A_jDHW5v3Q0_0(.dout(w_dff_A_L86RYP2Y6_0),.din(w_dff_A_jDHW5v3Q0_0),.clk(gclk));
	jdff dff_A_L86RYP2Y6_0(.dout(w_dff_A_Bhzq0YMv5_0),.din(w_dff_A_L86RYP2Y6_0),.clk(gclk));
	jdff dff_A_Bhzq0YMv5_0(.dout(w_dff_A_TbH3fasC7_0),.din(w_dff_A_Bhzq0YMv5_0),.clk(gclk));
	jdff dff_A_TbH3fasC7_0(.dout(w_dff_A_3gq02Vfb6_0),.din(w_dff_A_TbH3fasC7_0),.clk(gclk));
	jdff dff_A_3gq02Vfb6_0(.dout(w_dff_A_hZKeKtNB7_0),.din(w_dff_A_3gq02Vfb6_0),.clk(gclk));
	jdff dff_A_hZKeKtNB7_0(.dout(w_dff_A_80GCqJf52_0),.din(w_dff_A_hZKeKtNB7_0),.clk(gclk));
	jdff dff_A_80GCqJf52_0(.dout(w_dff_A_AP83QNGI4_0),.din(w_dff_A_80GCqJf52_0),.clk(gclk));
	jdff dff_A_AP83QNGI4_0(.dout(w_dff_A_46Jazfvb7_0),.din(w_dff_A_AP83QNGI4_0),.clk(gclk));
	jdff dff_A_46Jazfvb7_0(.dout(w_dff_A_8JMTCC4G7_0),.din(w_dff_A_46Jazfvb7_0),.clk(gclk));
	jdff dff_A_8JMTCC4G7_0(.dout(w_dff_A_igBzCly85_0),.din(w_dff_A_8JMTCC4G7_0),.clk(gclk));
	jdff dff_A_igBzCly85_0(.dout(w_dff_A_67uThCbv0_0),.din(w_dff_A_igBzCly85_0),.clk(gclk));
	jdff dff_A_67uThCbv0_0(.dout(w_dff_A_BMfnBHBV9_0),.din(w_dff_A_67uThCbv0_0),.clk(gclk));
	jdff dff_A_BMfnBHBV9_0(.dout(w_dff_A_KH7iVs1y8_0),.din(w_dff_A_BMfnBHBV9_0),.clk(gclk));
	jdff dff_A_KH7iVs1y8_0(.dout(w_dff_A_5sBtDR4h7_0),.din(w_dff_A_KH7iVs1y8_0),.clk(gclk));
	jdff dff_A_5sBtDR4h7_0(.dout(w_dff_A_3TARjgSY8_0),.din(w_dff_A_5sBtDR4h7_0),.clk(gclk));
	jdff dff_A_3TARjgSY8_0(.dout(w_dff_A_PXQYzuSd2_0),.din(w_dff_A_3TARjgSY8_0),.clk(gclk));
	jdff dff_A_PXQYzuSd2_0(.dout(w_dff_A_A5UXe75s6_0),.din(w_dff_A_PXQYzuSd2_0),.clk(gclk));
	jdff dff_A_A5UXe75s6_0(.dout(w_dff_A_VPlY73v35_0),.din(w_dff_A_A5UXe75s6_0),.clk(gclk));
	jdff dff_A_VPlY73v35_0(.dout(w_dff_A_9wkwbeZy1_0),.din(w_dff_A_VPlY73v35_0),.clk(gclk));
	jdff dff_A_9wkwbeZy1_0(.dout(w_dff_A_4k9ggX7N0_0),.din(w_dff_A_9wkwbeZy1_0),.clk(gclk));
	jdff dff_A_4k9ggX7N0_0(.dout(w_dff_A_IJrmdSH98_0),.din(w_dff_A_4k9ggX7N0_0),.clk(gclk));
	jdff dff_A_IJrmdSH98_0(.dout(w_dff_A_s9CQY1F47_0),.din(w_dff_A_IJrmdSH98_0),.clk(gclk));
	jdff dff_A_s9CQY1F47_0(.dout(w_dff_A_L4l8MKV24_0),.din(w_dff_A_s9CQY1F47_0),.clk(gclk));
	jdff dff_A_L4l8MKV24_0(.dout(w_dff_A_ep9F4Npv2_0),.din(w_dff_A_L4l8MKV24_0),.clk(gclk));
	jdff dff_A_ep9F4Npv2_0(.dout(w_dff_A_s7o1HIsz7_0),.din(w_dff_A_ep9F4Npv2_0),.clk(gclk));
	jdff dff_A_s7o1HIsz7_0(.dout(w_dff_A_Ot1OUzNt5_0),.din(w_dff_A_s7o1HIsz7_0),.clk(gclk));
	jdff dff_A_Ot1OUzNt5_0(.dout(w_dff_A_5OqTouOM2_0),.din(w_dff_A_Ot1OUzNt5_0),.clk(gclk));
	jdff dff_A_5OqTouOM2_0(.dout(w_dff_A_yjgt2cjq9_0),.din(w_dff_A_5OqTouOM2_0),.clk(gclk));
	jdff dff_A_yjgt2cjq9_0(.dout(w_dff_A_FCyEI8Ij2_0),.din(w_dff_A_yjgt2cjq9_0),.clk(gclk));
	jdff dff_A_FCyEI8Ij2_0(.dout(w_dff_A_XwTCm0QV6_0),.din(w_dff_A_FCyEI8Ij2_0),.clk(gclk));
	jdff dff_A_XwTCm0QV6_0(.dout(w_dff_A_ib8Pv4T83_0),.din(w_dff_A_XwTCm0QV6_0),.clk(gclk));
	jdff dff_A_ib8Pv4T83_0(.dout(w_dff_A_IoObJSrG4_0),.din(w_dff_A_ib8Pv4T83_0),.clk(gclk));
	jdff dff_A_IoObJSrG4_0(.dout(w_dff_A_i9lHLVO34_0),.din(w_dff_A_IoObJSrG4_0),.clk(gclk));
	jdff dff_A_i9lHLVO34_0(.dout(w_dff_A_8NAOYYnA8_0),.din(w_dff_A_i9lHLVO34_0),.clk(gclk));
	jdff dff_A_8NAOYYnA8_0(.dout(w_dff_A_0yLf0eDj1_0),.din(w_dff_A_8NAOYYnA8_0),.clk(gclk));
	jdff dff_A_0yLf0eDj1_0(.dout(w_dff_A_eAGRm9zi7_0),.din(w_dff_A_0yLf0eDj1_0),.clk(gclk));
	jdff dff_A_eAGRm9zi7_0(.dout(w_dff_A_Yabd95VT8_0),.din(w_dff_A_eAGRm9zi7_0),.clk(gclk));
	jdff dff_A_Yabd95VT8_0(.dout(w_dff_A_e21pVVJK5_0),.din(w_dff_A_Yabd95VT8_0),.clk(gclk));
	jdff dff_A_e21pVVJK5_0(.dout(w_dff_A_bCnAN8eK6_0),.din(w_dff_A_e21pVVJK5_0),.clk(gclk));
	jdff dff_A_bCnAN8eK6_0(.dout(w_dff_A_jEjHb6RW0_0),.din(w_dff_A_bCnAN8eK6_0),.clk(gclk));
	jdff dff_A_jEjHb6RW0_0(.dout(w_dff_A_OTF0tl1Z2_0),.din(w_dff_A_jEjHb6RW0_0),.clk(gclk));
	jdff dff_A_OTF0tl1Z2_0(.dout(w_dff_A_aA7Uiq1F0_0),.din(w_dff_A_OTF0tl1Z2_0),.clk(gclk));
	jdff dff_A_aA7Uiq1F0_0(.dout(w_dff_A_vqsK2C1f4_0),.din(w_dff_A_aA7Uiq1F0_0),.clk(gclk));
	jdff dff_A_vqsK2C1f4_0(.dout(w_dff_A_14hF01UT8_0),.din(w_dff_A_vqsK2C1f4_0),.clk(gclk));
	jdff dff_A_14hF01UT8_0(.dout(w_dff_A_mFl9UivU7_0),.din(w_dff_A_14hF01UT8_0),.clk(gclk));
	jdff dff_A_mFl9UivU7_0(.dout(w_dff_A_kOkCmNTa2_0),.din(w_dff_A_mFl9UivU7_0),.clk(gclk));
	jdff dff_A_kOkCmNTa2_0(.dout(w_dff_A_BlFefluR4_0),.din(w_dff_A_kOkCmNTa2_0),.clk(gclk));
	jdff dff_A_BlFefluR4_0(.dout(w_dff_A_4TduGLqi5_0),.din(w_dff_A_BlFefluR4_0),.clk(gclk));
	jdff dff_A_4TduGLqi5_0(.dout(w_dff_A_798Pic9G4_0),.din(w_dff_A_4TduGLqi5_0),.clk(gclk));
	jdff dff_A_798Pic9G4_0(.dout(w_dff_A_90x6earD2_0),.din(w_dff_A_798Pic9G4_0),.clk(gclk));
	jdff dff_A_90x6earD2_0(.dout(w_dff_A_EDcuu3vf3_0),.din(w_dff_A_90x6earD2_0),.clk(gclk));
	jdff dff_A_EDcuu3vf3_0(.dout(w_dff_A_gTxKXYil8_0),.din(w_dff_A_EDcuu3vf3_0),.clk(gclk));
	jdff dff_A_gTxKXYil8_0(.dout(w_dff_A_XQeKpwe45_0),.din(w_dff_A_gTxKXYil8_0),.clk(gclk));
	jdff dff_A_XQeKpwe45_0(.dout(w_dff_A_AlFKrb5A8_0),.din(w_dff_A_XQeKpwe45_0),.clk(gclk));
	jdff dff_A_AlFKrb5A8_0(.dout(w_dff_A_l3ffOSui7_0),.din(w_dff_A_AlFKrb5A8_0),.clk(gclk));
	jdff dff_A_l3ffOSui7_0(.dout(w_dff_A_K8tqUTVv5_0),.din(w_dff_A_l3ffOSui7_0),.clk(gclk));
	jdff dff_A_K8tqUTVv5_0(.dout(w_dff_A_HNGQKIgh5_0),.din(w_dff_A_K8tqUTVv5_0),.clk(gclk));
	jdff dff_A_HNGQKIgh5_0(.dout(w_dff_A_sBFbWx9O6_0),.din(w_dff_A_HNGQKIgh5_0),.clk(gclk));
	jdff dff_A_sBFbWx9O6_0(.dout(w_dff_A_WB9YxVfw4_0),.din(w_dff_A_sBFbWx9O6_0),.clk(gclk));
	jdff dff_A_WB9YxVfw4_0(.dout(G545gat),.din(w_dff_A_WB9YxVfw4_0),.clk(gclk));
	jdff dff_A_NslXWg0x3_2(.dout(w_dff_A_I5WThFvY9_0),.din(w_dff_A_NslXWg0x3_2),.clk(gclk));
	jdff dff_A_I5WThFvY9_0(.dout(w_dff_A_5rbu215e2_0),.din(w_dff_A_I5WThFvY9_0),.clk(gclk));
	jdff dff_A_5rbu215e2_0(.dout(w_dff_A_LPvp6EMm3_0),.din(w_dff_A_5rbu215e2_0),.clk(gclk));
	jdff dff_A_LPvp6EMm3_0(.dout(w_dff_A_pGhZ6fo68_0),.din(w_dff_A_LPvp6EMm3_0),.clk(gclk));
	jdff dff_A_pGhZ6fo68_0(.dout(w_dff_A_vFbWPHOG9_0),.din(w_dff_A_pGhZ6fo68_0),.clk(gclk));
	jdff dff_A_vFbWPHOG9_0(.dout(w_dff_A_Mr0aDnxi3_0),.din(w_dff_A_vFbWPHOG9_0),.clk(gclk));
	jdff dff_A_Mr0aDnxi3_0(.dout(w_dff_A_jhmVoLMs2_0),.din(w_dff_A_Mr0aDnxi3_0),.clk(gclk));
	jdff dff_A_jhmVoLMs2_0(.dout(w_dff_A_euC441m84_0),.din(w_dff_A_jhmVoLMs2_0),.clk(gclk));
	jdff dff_A_euC441m84_0(.dout(w_dff_A_F4hX5uHX8_0),.din(w_dff_A_euC441m84_0),.clk(gclk));
	jdff dff_A_F4hX5uHX8_0(.dout(w_dff_A_AI2F0nfn2_0),.din(w_dff_A_F4hX5uHX8_0),.clk(gclk));
	jdff dff_A_AI2F0nfn2_0(.dout(w_dff_A_f3mjBQUq4_0),.din(w_dff_A_AI2F0nfn2_0),.clk(gclk));
	jdff dff_A_f3mjBQUq4_0(.dout(w_dff_A_0WOiSrou4_0),.din(w_dff_A_f3mjBQUq4_0),.clk(gclk));
	jdff dff_A_0WOiSrou4_0(.dout(w_dff_A_cYLQHQBX9_0),.din(w_dff_A_0WOiSrou4_0),.clk(gclk));
	jdff dff_A_cYLQHQBX9_0(.dout(w_dff_A_eonTJ2wl7_0),.din(w_dff_A_cYLQHQBX9_0),.clk(gclk));
	jdff dff_A_eonTJ2wl7_0(.dout(w_dff_A_XeqP43tG6_0),.din(w_dff_A_eonTJ2wl7_0),.clk(gclk));
	jdff dff_A_XeqP43tG6_0(.dout(w_dff_A_UOwWTtj39_0),.din(w_dff_A_XeqP43tG6_0),.clk(gclk));
	jdff dff_A_UOwWTtj39_0(.dout(w_dff_A_fIalWi3U6_0),.din(w_dff_A_UOwWTtj39_0),.clk(gclk));
	jdff dff_A_fIalWi3U6_0(.dout(w_dff_A_8wTPooyb8_0),.din(w_dff_A_fIalWi3U6_0),.clk(gclk));
	jdff dff_A_8wTPooyb8_0(.dout(w_dff_A_aZ5rjZAr3_0),.din(w_dff_A_8wTPooyb8_0),.clk(gclk));
	jdff dff_A_aZ5rjZAr3_0(.dout(w_dff_A_UPEs4K000_0),.din(w_dff_A_aZ5rjZAr3_0),.clk(gclk));
	jdff dff_A_UPEs4K000_0(.dout(w_dff_A_axL163r37_0),.din(w_dff_A_UPEs4K000_0),.clk(gclk));
	jdff dff_A_axL163r37_0(.dout(w_dff_A_Jj1EUh8x7_0),.din(w_dff_A_axL163r37_0),.clk(gclk));
	jdff dff_A_Jj1EUh8x7_0(.dout(w_dff_A_rh3nVGxM1_0),.din(w_dff_A_Jj1EUh8x7_0),.clk(gclk));
	jdff dff_A_rh3nVGxM1_0(.dout(w_dff_A_eVuzDtIV0_0),.din(w_dff_A_rh3nVGxM1_0),.clk(gclk));
	jdff dff_A_eVuzDtIV0_0(.dout(w_dff_A_MzRNPNfU3_0),.din(w_dff_A_eVuzDtIV0_0),.clk(gclk));
	jdff dff_A_MzRNPNfU3_0(.dout(w_dff_A_YXKRck8f6_0),.din(w_dff_A_MzRNPNfU3_0),.clk(gclk));
	jdff dff_A_YXKRck8f6_0(.dout(w_dff_A_88pVLx314_0),.din(w_dff_A_YXKRck8f6_0),.clk(gclk));
	jdff dff_A_88pVLx314_0(.dout(w_dff_A_3EdiyTJZ3_0),.din(w_dff_A_88pVLx314_0),.clk(gclk));
	jdff dff_A_3EdiyTJZ3_0(.dout(w_dff_A_qwSl4dj92_0),.din(w_dff_A_3EdiyTJZ3_0),.clk(gclk));
	jdff dff_A_qwSl4dj92_0(.dout(w_dff_A_lBMi7rQc6_0),.din(w_dff_A_qwSl4dj92_0),.clk(gclk));
	jdff dff_A_lBMi7rQc6_0(.dout(w_dff_A_tPeRy6r72_0),.din(w_dff_A_lBMi7rQc6_0),.clk(gclk));
	jdff dff_A_tPeRy6r72_0(.dout(w_dff_A_HR5LP9AX2_0),.din(w_dff_A_tPeRy6r72_0),.clk(gclk));
	jdff dff_A_HR5LP9AX2_0(.dout(w_dff_A_7eglWOl51_0),.din(w_dff_A_HR5LP9AX2_0),.clk(gclk));
	jdff dff_A_7eglWOl51_0(.dout(w_dff_A_56AO8c590_0),.din(w_dff_A_7eglWOl51_0),.clk(gclk));
	jdff dff_A_56AO8c590_0(.dout(w_dff_A_eVUbKRmL7_0),.din(w_dff_A_56AO8c590_0),.clk(gclk));
	jdff dff_A_eVUbKRmL7_0(.dout(w_dff_A_QDLcDh6t8_0),.din(w_dff_A_eVUbKRmL7_0),.clk(gclk));
	jdff dff_A_QDLcDh6t8_0(.dout(w_dff_A_yPHr171L6_0),.din(w_dff_A_QDLcDh6t8_0),.clk(gclk));
	jdff dff_A_yPHr171L6_0(.dout(w_dff_A_ZZ4hvhWL9_0),.din(w_dff_A_yPHr171L6_0),.clk(gclk));
	jdff dff_A_ZZ4hvhWL9_0(.dout(w_dff_A_XvX4plDk1_0),.din(w_dff_A_ZZ4hvhWL9_0),.clk(gclk));
	jdff dff_A_XvX4plDk1_0(.dout(w_dff_A_1a3VfOzx3_0),.din(w_dff_A_XvX4plDk1_0),.clk(gclk));
	jdff dff_A_1a3VfOzx3_0(.dout(w_dff_A_75n9HyO70_0),.din(w_dff_A_1a3VfOzx3_0),.clk(gclk));
	jdff dff_A_75n9HyO70_0(.dout(w_dff_A_wQMs33ol9_0),.din(w_dff_A_75n9HyO70_0),.clk(gclk));
	jdff dff_A_wQMs33ol9_0(.dout(w_dff_A_d51U9rm39_0),.din(w_dff_A_wQMs33ol9_0),.clk(gclk));
	jdff dff_A_d51U9rm39_0(.dout(w_dff_A_xomWgcyQ5_0),.din(w_dff_A_d51U9rm39_0),.clk(gclk));
	jdff dff_A_xomWgcyQ5_0(.dout(w_dff_A_eutneaXU6_0),.din(w_dff_A_xomWgcyQ5_0),.clk(gclk));
	jdff dff_A_eutneaXU6_0(.dout(w_dff_A_9fKHYyrl0_0),.din(w_dff_A_eutneaXU6_0),.clk(gclk));
	jdff dff_A_9fKHYyrl0_0(.dout(w_dff_A_fyhr0Jde6_0),.din(w_dff_A_9fKHYyrl0_0),.clk(gclk));
	jdff dff_A_fyhr0Jde6_0(.dout(w_dff_A_tEs4guOG1_0),.din(w_dff_A_fyhr0Jde6_0),.clk(gclk));
	jdff dff_A_tEs4guOG1_0(.dout(w_dff_A_dp3mvErr8_0),.din(w_dff_A_tEs4guOG1_0),.clk(gclk));
	jdff dff_A_dp3mvErr8_0(.dout(w_dff_A_wynkwt1E3_0),.din(w_dff_A_dp3mvErr8_0),.clk(gclk));
	jdff dff_A_wynkwt1E3_0(.dout(w_dff_A_y2v0RrB84_0),.din(w_dff_A_wynkwt1E3_0),.clk(gclk));
	jdff dff_A_y2v0RrB84_0(.dout(w_dff_A_eYPdsBSX3_0),.din(w_dff_A_y2v0RrB84_0),.clk(gclk));
	jdff dff_A_eYPdsBSX3_0(.dout(w_dff_A_yV8RrRx57_0),.din(w_dff_A_eYPdsBSX3_0),.clk(gclk));
	jdff dff_A_yV8RrRx57_0(.dout(w_dff_A_Q9puzdqY5_0),.din(w_dff_A_yV8RrRx57_0),.clk(gclk));
	jdff dff_A_Q9puzdqY5_0(.dout(w_dff_A_05HWikCa1_0),.din(w_dff_A_Q9puzdqY5_0),.clk(gclk));
	jdff dff_A_05HWikCa1_0(.dout(w_dff_A_SuWjL1B27_0),.din(w_dff_A_05HWikCa1_0),.clk(gclk));
	jdff dff_A_SuWjL1B27_0(.dout(w_dff_A_9KudURsQ1_0),.din(w_dff_A_SuWjL1B27_0),.clk(gclk));
	jdff dff_A_9KudURsQ1_0(.dout(w_dff_A_v5nks1rE4_0),.din(w_dff_A_9KudURsQ1_0),.clk(gclk));
	jdff dff_A_v5nks1rE4_0(.dout(w_dff_A_umQly1M49_0),.din(w_dff_A_v5nks1rE4_0),.clk(gclk));
	jdff dff_A_umQly1M49_0(.dout(w_dff_A_sk2oOwGJ4_0),.din(w_dff_A_umQly1M49_0),.clk(gclk));
	jdff dff_A_sk2oOwGJ4_0(.dout(w_dff_A_T6E2pNcF1_0),.din(w_dff_A_sk2oOwGJ4_0),.clk(gclk));
	jdff dff_A_T6E2pNcF1_0(.dout(w_dff_A_uwSLX6KQ6_0),.din(w_dff_A_T6E2pNcF1_0),.clk(gclk));
	jdff dff_A_uwSLX6KQ6_0(.dout(w_dff_A_6CYW7BgD0_0),.din(w_dff_A_uwSLX6KQ6_0),.clk(gclk));
	jdff dff_A_6CYW7BgD0_0(.dout(w_dff_A_VrJxdA0N5_0),.din(w_dff_A_6CYW7BgD0_0),.clk(gclk));
	jdff dff_A_VrJxdA0N5_0(.dout(w_dff_A_mQuFLoBo3_0),.din(w_dff_A_VrJxdA0N5_0),.clk(gclk));
	jdff dff_A_mQuFLoBo3_0(.dout(w_dff_A_ypOMHuoY4_0),.din(w_dff_A_mQuFLoBo3_0),.clk(gclk));
	jdff dff_A_ypOMHuoY4_0(.dout(w_dff_A_ef3ofoF17_0),.din(w_dff_A_ypOMHuoY4_0),.clk(gclk));
	jdff dff_A_ef3ofoF17_0(.dout(w_dff_A_CGlm3Azc7_0),.din(w_dff_A_ef3ofoF17_0),.clk(gclk));
	jdff dff_A_CGlm3Azc7_0(.dout(w_dff_A_0EJiQWms3_0),.din(w_dff_A_CGlm3Azc7_0),.clk(gclk));
	jdff dff_A_0EJiQWms3_0(.dout(G1581gat),.din(w_dff_A_0EJiQWms3_0),.clk(gclk));
	jdff dff_A_aqNNkNcQ8_2(.dout(w_dff_A_Bcadps6G9_0),.din(w_dff_A_aqNNkNcQ8_2),.clk(gclk));
	jdff dff_A_Bcadps6G9_0(.dout(w_dff_A_JngHxxGD0_0),.din(w_dff_A_Bcadps6G9_0),.clk(gclk));
	jdff dff_A_JngHxxGD0_0(.dout(w_dff_A_qnXymM9S5_0),.din(w_dff_A_JngHxxGD0_0),.clk(gclk));
	jdff dff_A_qnXymM9S5_0(.dout(w_dff_A_XFGSbv049_0),.din(w_dff_A_qnXymM9S5_0),.clk(gclk));
	jdff dff_A_XFGSbv049_0(.dout(w_dff_A_iAPNqVDe6_0),.din(w_dff_A_XFGSbv049_0),.clk(gclk));
	jdff dff_A_iAPNqVDe6_0(.dout(w_dff_A_7JWiMhIr6_0),.din(w_dff_A_iAPNqVDe6_0),.clk(gclk));
	jdff dff_A_7JWiMhIr6_0(.dout(w_dff_A_DIApHEs70_0),.din(w_dff_A_7JWiMhIr6_0),.clk(gclk));
	jdff dff_A_DIApHEs70_0(.dout(w_dff_A_uqToj7HG0_0),.din(w_dff_A_DIApHEs70_0),.clk(gclk));
	jdff dff_A_uqToj7HG0_0(.dout(w_dff_A_iRIcnbg91_0),.din(w_dff_A_uqToj7HG0_0),.clk(gclk));
	jdff dff_A_iRIcnbg91_0(.dout(w_dff_A_lXmb7PkR3_0),.din(w_dff_A_iRIcnbg91_0),.clk(gclk));
	jdff dff_A_lXmb7PkR3_0(.dout(w_dff_A_ykG41ovV2_0),.din(w_dff_A_lXmb7PkR3_0),.clk(gclk));
	jdff dff_A_ykG41ovV2_0(.dout(w_dff_A_0OoSYOW68_0),.din(w_dff_A_ykG41ovV2_0),.clk(gclk));
	jdff dff_A_0OoSYOW68_0(.dout(w_dff_A_p11g2EET9_0),.din(w_dff_A_0OoSYOW68_0),.clk(gclk));
	jdff dff_A_p11g2EET9_0(.dout(w_dff_A_wR0RbipV7_0),.din(w_dff_A_p11g2EET9_0),.clk(gclk));
	jdff dff_A_wR0RbipV7_0(.dout(w_dff_A_CuuGmkAA3_0),.din(w_dff_A_wR0RbipV7_0),.clk(gclk));
	jdff dff_A_CuuGmkAA3_0(.dout(w_dff_A_x21qsiKw8_0),.din(w_dff_A_CuuGmkAA3_0),.clk(gclk));
	jdff dff_A_x21qsiKw8_0(.dout(w_dff_A_U19Zw9DS5_0),.din(w_dff_A_x21qsiKw8_0),.clk(gclk));
	jdff dff_A_U19Zw9DS5_0(.dout(w_dff_A_wTBy4Y314_0),.din(w_dff_A_U19Zw9DS5_0),.clk(gclk));
	jdff dff_A_wTBy4Y314_0(.dout(w_dff_A_3ZPyqDpN0_0),.din(w_dff_A_wTBy4Y314_0),.clk(gclk));
	jdff dff_A_3ZPyqDpN0_0(.dout(w_dff_A_emNpalZw6_0),.din(w_dff_A_3ZPyqDpN0_0),.clk(gclk));
	jdff dff_A_emNpalZw6_0(.dout(w_dff_A_JgSWAHOr3_0),.din(w_dff_A_emNpalZw6_0),.clk(gclk));
	jdff dff_A_JgSWAHOr3_0(.dout(w_dff_A_iENyi0Ou2_0),.din(w_dff_A_JgSWAHOr3_0),.clk(gclk));
	jdff dff_A_iENyi0Ou2_0(.dout(w_dff_A_l8YRJB5X1_0),.din(w_dff_A_iENyi0Ou2_0),.clk(gclk));
	jdff dff_A_l8YRJB5X1_0(.dout(w_dff_A_ngCzv0wq8_0),.din(w_dff_A_l8YRJB5X1_0),.clk(gclk));
	jdff dff_A_ngCzv0wq8_0(.dout(w_dff_A_7jrJ0Wn38_0),.din(w_dff_A_ngCzv0wq8_0),.clk(gclk));
	jdff dff_A_7jrJ0Wn38_0(.dout(w_dff_A_vhVA9I2D5_0),.din(w_dff_A_7jrJ0Wn38_0),.clk(gclk));
	jdff dff_A_vhVA9I2D5_0(.dout(w_dff_A_nGdAGcDr6_0),.din(w_dff_A_vhVA9I2D5_0),.clk(gclk));
	jdff dff_A_nGdAGcDr6_0(.dout(w_dff_A_MvXObyMj3_0),.din(w_dff_A_nGdAGcDr6_0),.clk(gclk));
	jdff dff_A_MvXObyMj3_0(.dout(w_dff_A_Ge9b69P73_0),.din(w_dff_A_MvXObyMj3_0),.clk(gclk));
	jdff dff_A_Ge9b69P73_0(.dout(w_dff_A_ioWSYgyo1_0),.din(w_dff_A_Ge9b69P73_0),.clk(gclk));
	jdff dff_A_ioWSYgyo1_0(.dout(w_dff_A_rDyev51K2_0),.din(w_dff_A_ioWSYgyo1_0),.clk(gclk));
	jdff dff_A_rDyev51K2_0(.dout(w_dff_A_KuPz8kQQ4_0),.din(w_dff_A_rDyev51K2_0),.clk(gclk));
	jdff dff_A_KuPz8kQQ4_0(.dout(w_dff_A_086ab7BX0_0),.din(w_dff_A_KuPz8kQQ4_0),.clk(gclk));
	jdff dff_A_086ab7BX0_0(.dout(w_dff_A_8d3JbXYl3_0),.din(w_dff_A_086ab7BX0_0),.clk(gclk));
	jdff dff_A_8d3JbXYl3_0(.dout(w_dff_A_XIdSLnhK1_0),.din(w_dff_A_8d3JbXYl3_0),.clk(gclk));
	jdff dff_A_XIdSLnhK1_0(.dout(w_dff_A_4C0Rxurq5_0),.din(w_dff_A_XIdSLnhK1_0),.clk(gclk));
	jdff dff_A_4C0Rxurq5_0(.dout(w_dff_A_YiMzQWIM0_0),.din(w_dff_A_4C0Rxurq5_0),.clk(gclk));
	jdff dff_A_YiMzQWIM0_0(.dout(w_dff_A_sBLe3Nxr3_0),.din(w_dff_A_YiMzQWIM0_0),.clk(gclk));
	jdff dff_A_sBLe3Nxr3_0(.dout(w_dff_A_sK0OXaTN4_0),.din(w_dff_A_sBLe3Nxr3_0),.clk(gclk));
	jdff dff_A_sK0OXaTN4_0(.dout(w_dff_A_kHePytj39_0),.din(w_dff_A_sK0OXaTN4_0),.clk(gclk));
	jdff dff_A_kHePytj39_0(.dout(w_dff_A_XkN0OuQz6_0),.din(w_dff_A_kHePytj39_0),.clk(gclk));
	jdff dff_A_XkN0OuQz6_0(.dout(w_dff_A_9CQ9uvkB1_0),.din(w_dff_A_XkN0OuQz6_0),.clk(gclk));
	jdff dff_A_9CQ9uvkB1_0(.dout(w_dff_A_xFxhVMVn4_0),.din(w_dff_A_9CQ9uvkB1_0),.clk(gclk));
	jdff dff_A_xFxhVMVn4_0(.dout(w_dff_A_p9jxaPIf0_0),.din(w_dff_A_xFxhVMVn4_0),.clk(gclk));
	jdff dff_A_p9jxaPIf0_0(.dout(w_dff_A_HMnq1jw19_0),.din(w_dff_A_p9jxaPIf0_0),.clk(gclk));
	jdff dff_A_HMnq1jw19_0(.dout(w_dff_A_UdjTtzgm6_0),.din(w_dff_A_HMnq1jw19_0),.clk(gclk));
	jdff dff_A_UdjTtzgm6_0(.dout(w_dff_A_mmcb6lT62_0),.din(w_dff_A_UdjTtzgm6_0),.clk(gclk));
	jdff dff_A_mmcb6lT62_0(.dout(w_dff_A_sZBaC4AJ7_0),.din(w_dff_A_mmcb6lT62_0),.clk(gclk));
	jdff dff_A_sZBaC4AJ7_0(.dout(w_dff_A_6OPiAxXu3_0),.din(w_dff_A_sZBaC4AJ7_0),.clk(gclk));
	jdff dff_A_6OPiAxXu3_0(.dout(w_dff_A_IgyQ1NGe8_0),.din(w_dff_A_6OPiAxXu3_0),.clk(gclk));
	jdff dff_A_IgyQ1NGe8_0(.dout(w_dff_A_lHISZ7A64_0),.din(w_dff_A_IgyQ1NGe8_0),.clk(gclk));
	jdff dff_A_lHISZ7A64_0(.dout(w_dff_A_zV21c5Ja7_0),.din(w_dff_A_lHISZ7A64_0),.clk(gclk));
	jdff dff_A_zV21c5Ja7_0(.dout(w_dff_A_QhYHca3w4_0),.din(w_dff_A_zV21c5Ja7_0),.clk(gclk));
	jdff dff_A_QhYHca3w4_0(.dout(w_dff_A_dvsVWLrZ3_0),.din(w_dff_A_QhYHca3w4_0),.clk(gclk));
	jdff dff_A_dvsVWLrZ3_0(.dout(w_dff_A_MQ6t6Fq74_0),.din(w_dff_A_dvsVWLrZ3_0),.clk(gclk));
	jdff dff_A_MQ6t6Fq74_0(.dout(w_dff_A_rTDSSZh00_0),.din(w_dff_A_MQ6t6Fq74_0),.clk(gclk));
	jdff dff_A_rTDSSZh00_0(.dout(w_dff_A_ku56SRiv8_0),.din(w_dff_A_rTDSSZh00_0),.clk(gclk));
	jdff dff_A_ku56SRiv8_0(.dout(w_dff_A_Ui8RXGmf2_0),.din(w_dff_A_ku56SRiv8_0),.clk(gclk));
	jdff dff_A_Ui8RXGmf2_0(.dout(w_dff_A_jo8J4tIO0_0),.din(w_dff_A_Ui8RXGmf2_0),.clk(gclk));
	jdff dff_A_jo8J4tIO0_0(.dout(w_dff_A_lhCUuOAq9_0),.din(w_dff_A_jo8J4tIO0_0),.clk(gclk));
	jdff dff_A_lhCUuOAq9_0(.dout(w_dff_A_9dS3Pf2z3_0),.din(w_dff_A_lhCUuOAq9_0),.clk(gclk));
	jdff dff_A_9dS3Pf2z3_0(.dout(w_dff_A_D4LRZqVc4_0),.din(w_dff_A_9dS3Pf2z3_0),.clk(gclk));
	jdff dff_A_D4LRZqVc4_0(.dout(w_dff_A_cG1P65du0_0),.din(w_dff_A_D4LRZqVc4_0),.clk(gclk));
	jdff dff_A_cG1P65du0_0(.dout(w_dff_A_jo7a9cxF6_0),.din(w_dff_A_cG1P65du0_0),.clk(gclk));
	jdff dff_A_jo7a9cxF6_0(.dout(w_dff_A_8AhaQ92M4_0),.din(w_dff_A_jo7a9cxF6_0),.clk(gclk));
	jdff dff_A_8AhaQ92M4_0(.dout(w_dff_A_2aFfJTxd9_0),.din(w_dff_A_8AhaQ92M4_0),.clk(gclk));
	jdff dff_A_2aFfJTxd9_0(.dout(w_dff_A_uyEcTvc40_0),.din(w_dff_A_2aFfJTxd9_0),.clk(gclk));
	jdff dff_A_uyEcTvc40_0(.dout(w_dff_A_OdNAlUUY1_0),.din(w_dff_A_uyEcTvc40_0),.clk(gclk));
	jdff dff_A_OdNAlUUY1_0(.dout(G1901gat),.din(w_dff_A_OdNAlUUY1_0),.clk(gclk));
	jdff dff_A_ia5znL6j8_2(.dout(w_dff_A_Sil0NLgq3_0),.din(w_dff_A_ia5znL6j8_2),.clk(gclk));
	jdff dff_A_Sil0NLgq3_0(.dout(w_dff_A_VT5zNKAv4_0),.din(w_dff_A_Sil0NLgq3_0),.clk(gclk));
	jdff dff_A_VT5zNKAv4_0(.dout(w_dff_A_ir5PzM1t9_0),.din(w_dff_A_VT5zNKAv4_0),.clk(gclk));
	jdff dff_A_ir5PzM1t9_0(.dout(w_dff_A_1WKU4g5p9_0),.din(w_dff_A_ir5PzM1t9_0),.clk(gclk));
	jdff dff_A_1WKU4g5p9_0(.dout(w_dff_A_1onpxYXY2_0),.din(w_dff_A_1WKU4g5p9_0),.clk(gclk));
	jdff dff_A_1onpxYXY2_0(.dout(w_dff_A_1zanhRZy4_0),.din(w_dff_A_1onpxYXY2_0),.clk(gclk));
	jdff dff_A_1zanhRZy4_0(.dout(w_dff_A_3e91Gvn39_0),.din(w_dff_A_1zanhRZy4_0),.clk(gclk));
	jdff dff_A_3e91Gvn39_0(.dout(w_dff_A_006MIS991_0),.din(w_dff_A_3e91Gvn39_0),.clk(gclk));
	jdff dff_A_006MIS991_0(.dout(w_dff_A_12b4hOkc4_0),.din(w_dff_A_006MIS991_0),.clk(gclk));
	jdff dff_A_12b4hOkc4_0(.dout(w_dff_A_RaRIIDE68_0),.din(w_dff_A_12b4hOkc4_0),.clk(gclk));
	jdff dff_A_RaRIIDE68_0(.dout(w_dff_A_yaWVbUjb0_0),.din(w_dff_A_RaRIIDE68_0),.clk(gclk));
	jdff dff_A_yaWVbUjb0_0(.dout(w_dff_A_kKb2a76c1_0),.din(w_dff_A_yaWVbUjb0_0),.clk(gclk));
	jdff dff_A_kKb2a76c1_0(.dout(w_dff_A_a9hHyqNs9_0),.din(w_dff_A_kKb2a76c1_0),.clk(gclk));
	jdff dff_A_a9hHyqNs9_0(.dout(w_dff_A_52yL5Oir8_0),.din(w_dff_A_a9hHyqNs9_0),.clk(gclk));
	jdff dff_A_52yL5Oir8_0(.dout(w_dff_A_kMpLpclI6_0),.din(w_dff_A_52yL5Oir8_0),.clk(gclk));
	jdff dff_A_kMpLpclI6_0(.dout(w_dff_A_oucS8qp29_0),.din(w_dff_A_kMpLpclI6_0),.clk(gclk));
	jdff dff_A_oucS8qp29_0(.dout(w_dff_A_ZYdeFAQq7_0),.din(w_dff_A_oucS8qp29_0),.clk(gclk));
	jdff dff_A_ZYdeFAQq7_0(.dout(w_dff_A_sv5qDQit8_0),.din(w_dff_A_ZYdeFAQq7_0),.clk(gclk));
	jdff dff_A_sv5qDQit8_0(.dout(w_dff_A_cHT48gSs5_0),.din(w_dff_A_sv5qDQit8_0),.clk(gclk));
	jdff dff_A_cHT48gSs5_0(.dout(w_dff_A_Gzjyp4tK6_0),.din(w_dff_A_cHT48gSs5_0),.clk(gclk));
	jdff dff_A_Gzjyp4tK6_0(.dout(w_dff_A_8H9vCOIc4_0),.din(w_dff_A_Gzjyp4tK6_0),.clk(gclk));
	jdff dff_A_8H9vCOIc4_0(.dout(w_dff_A_62FQUY7e9_0),.din(w_dff_A_8H9vCOIc4_0),.clk(gclk));
	jdff dff_A_62FQUY7e9_0(.dout(w_dff_A_hrELfqsW8_0),.din(w_dff_A_62FQUY7e9_0),.clk(gclk));
	jdff dff_A_hrELfqsW8_0(.dout(w_dff_A_KDBF3E607_0),.din(w_dff_A_hrELfqsW8_0),.clk(gclk));
	jdff dff_A_KDBF3E607_0(.dout(w_dff_A_ohHlkvwA4_0),.din(w_dff_A_KDBF3E607_0),.clk(gclk));
	jdff dff_A_ohHlkvwA4_0(.dout(w_dff_A_lVYVVi217_0),.din(w_dff_A_ohHlkvwA4_0),.clk(gclk));
	jdff dff_A_lVYVVi217_0(.dout(w_dff_A_ojj653AN2_0),.din(w_dff_A_lVYVVi217_0),.clk(gclk));
	jdff dff_A_ojj653AN2_0(.dout(w_dff_A_PzchLUhG1_0),.din(w_dff_A_ojj653AN2_0),.clk(gclk));
	jdff dff_A_PzchLUhG1_0(.dout(w_dff_A_304jaEvm3_0),.din(w_dff_A_PzchLUhG1_0),.clk(gclk));
	jdff dff_A_304jaEvm3_0(.dout(w_dff_A_8SnIt23R3_0),.din(w_dff_A_304jaEvm3_0),.clk(gclk));
	jdff dff_A_8SnIt23R3_0(.dout(w_dff_A_2dkQMxX12_0),.din(w_dff_A_8SnIt23R3_0),.clk(gclk));
	jdff dff_A_2dkQMxX12_0(.dout(w_dff_A_sTkaVVIg9_0),.din(w_dff_A_2dkQMxX12_0),.clk(gclk));
	jdff dff_A_sTkaVVIg9_0(.dout(w_dff_A_cQXSYRbY8_0),.din(w_dff_A_sTkaVVIg9_0),.clk(gclk));
	jdff dff_A_cQXSYRbY8_0(.dout(w_dff_A_zSo2aDVP3_0),.din(w_dff_A_cQXSYRbY8_0),.clk(gclk));
	jdff dff_A_zSo2aDVP3_0(.dout(w_dff_A_HPhFy2ab9_0),.din(w_dff_A_zSo2aDVP3_0),.clk(gclk));
	jdff dff_A_HPhFy2ab9_0(.dout(w_dff_A_3tdAzL8v3_0),.din(w_dff_A_HPhFy2ab9_0),.clk(gclk));
	jdff dff_A_3tdAzL8v3_0(.dout(w_dff_A_5FcrTReg5_0),.din(w_dff_A_3tdAzL8v3_0),.clk(gclk));
	jdff dff_A_5FcrTReg5_0(.dout(w_dff_A_6eUgR59u9_0),.din(w_dff_A_5FcrTReg5_0),.clk(gclk));
	jdff dff_A_6eUgR59u9_0(.dout(w_dff_A_8CUDCYJB8_0),.din(w_dff_A_6eUgR59u9_0),.clk(gclk));
	jdff dff_A_8CUDCYJB8_0(.dout(w_dff_A_nDsTolMs8_0),.din(w_dff_A_8CUDCYJB8_0),.clk(gclk));
	jdff dff_A_nDsTolMs8_0(.dout(w_dff_A_R7vr0vRE3_0),.din(w_dff_A_nDsTolMs8_0),.clk(gclk));
	jdff dff_A_R7vr0vRE3_0(.dout(w_dff_A_kgUuWbe53_0),.din(w_dff_A_R7vr0vRE3_0),.clk(gclk));
	jdff dff_A_kgUuWbe53_0(.dout(w_dff_A_7NRKMlg45_0),.din(w_dff_A_kgUuWbe53_0),.clk(gclk));
	jdff dff_A_7NRKMlg45_0(.dout(w_dff_A_Y8H8L4Mh7_0),.din(w_dff_A_7NRKMlg45_0),.clk(gclk));
	jdff dff_A_Y8H8L4Mh7_0(.dout(w_dff_A_9uTIdewM4_0),.din(w_dff_A_Y8H8L4Mh7_0),.clk(gclk));
	jdff dff_A_9uTIdewM4_0(.dout(w_dff_A_5cH6oclo9_0),.din(w_dff_A_9uTIdewM4_0),.clk(gclk));
	jdff dff_A_5cH6oclo9_0(.dout(w_dff_A_VmwPEXiV7_0),.din(w_dff_A_5cH6oclo9_0),.clk(gclk));
	jdff dff_A_VmwPEXiV7_0(.dout(w_dff_A_FmS0ciSa2_0),.din(w_dff_A_VmwPEXiV7_0),.clk(gclk));
	jdff dff_A_FmS0ciSa2_0(.dout(w_dff_A_RVgKvPYQ5_0),.din(w_dff_A_FmS0ciSa2_0),.clk(gclk));
	jdff dff_A_RVgKvPYQ5_0(.dout(w_dff_A_1PDFdbZK4_0),.din(w_dff_A_RVgKvPYQ5_0),.clk(gclk));
	jdff dff_A_1PDFdbZK4_0(.dout(w_dff_A_VMHJ3NcX1_0),.din(w_dff_A_1PDFdbZK4_0),.clk(gclk));
	jdff dff_A_VMHJ3NcX1_0(.dout(w_dff_A_s5vgirpi1_0),.din(w_dff_A_VMHJ3NcX1_0),.clk(gclk));
	jdff dff_A_s5vgirpi1_0(.dout(w_dff_A_KozlldQB5_0),.din(w_dff_A_s5vgirpi1_0),.clk(gclk));
	jdff dff_A_KozlldQB5_0(.dout(w_dff_A_fuQVxD3L5_0),.din(w_dff_A_KozlldQB5_0),.clk(gclk));
	jdff dff_A_fuQVxD3L5_0(.dout(w_dff_A_aO651zeA7_0),.din(w_dff_A_fuQVxD3L5_0),.clk(gclk));
	jdff dff_A_aO651zeA7_0(.dout(w_dff_A_mpVyZMfs2_0),.din(w_dff_A_aO651zeA7_0),.clk(gclk));
	jdff dff_A_mpVyZMfs2_0(.dout(w_dff_A_TjdUyd1m3_0),.din(w_dff_A_mpVyZMfs2_0),.clk(gclk));
	jdff dff_A_TjdUyd1m3_0(.dout(w_dff_A_hmaBXeqC7_0),.din(w_dff_A_TjdUyd1m3_0),.clk(gclk));
	jdff dff_A_hmaBXeqC7_0(.dout(w_dff_A_JhClA7XN6_0),.din(w_dff_A_hmaBXeqC7_0),.clk(gclk));
	jdff dff_A_JhClA7XN6_0(.dout(w_dff_A_d1D5AJHx9_0),.din(w_dff_A_JhClA7XN6_0),.clk(gclk));
	jdff dff_A_d1D5AJHx9_0(.dout(w_dff_A_R2OefjDr9_0),.din(w_dff_A_d1D5AJHx9_0),.clk(gclk));
	jdff dff_A_R2OefjDr9_0(.dout(w_dff_A_2F0U9oUi3_0),.din(w_dff_A_R2OefjDr9_0),.clk(gclk));
	jdff dff_A_2F0U9oUi3_0(.dout(w_dff_A_bCQyzGeO1_0),.din(w_dff_A_2F0U9oUi3_0),.clk(gclk));
	jdff dff_A_bCQyzGeO1_0(.dout(w_dff_A_EtvmkPLL6_0),.din(w_dff_A_bCQyzGeO1_0),.clk(gclk));
	jdff dff_A_EtvmkPLL6_0(.dout(w_dff_A_fnBrgqSm5_0),.din(w_dff_A_EtvmkPLL6_0),.clk(gclk));
	jdff dff_A_fnBrgqSm5_0(.dout(G2223gat),.din(w_dff_A_fnBrgqSm5_0),.clk(gclk));
	jdff dff_A_aLbf6XPK1_2(.dout(w_dff_A_QaP3D5ZU3_0),.din(w_dff_A_aLbf6XPK1_2),.clk(gclk));
	jdff dff_A_QaP3D5ZU3_0(.dout(w_dff_A_LjmKnrxD5_0),.din(w_dff_A_QaP3D5ZU3_0),.clk(gclk));
	jdff dff_A_LjmKnrxD5_0(.dout(w_dff_A_ENeHB0fV4_0),.din(w_dff_A_LjmKnrxD5_0),.clk(gclk));
	jdff dff_A_ENeHB0fV4_0(.dout(w_dff_A_R54V7n3i8_0),.din(w_dff_A_ENeHB0fV4_0),.clk(gclk));
	jdff dff_A_R54V7n3i8_0(.dout(w_dff_A_o52T4KMF8_0),.din(w_dff_A_R54V7n3i8_0),.clk(gclk));
	jdff dff_A_o52T4KMF8_0(.dout(w_dff_A_CvZlUgDk0_0),.din(w_dff_A_o52T4KMF8_0),.clk(gclk));
	jdff dff_A_CvZlUgDk0_0(.dout(w_dff_A_GvQDGDh67_0),.din(w_dff_A_CvZlUgDk0_0),.clk(gclk));
	jdff dff_A_GvQDGDh67_0(.dout(w_dff_A_bh2APSLp6_0),.din(w_dff_A_GvQDGDh67_0),.clk(gclk));
	jdff dff_A_bh2APSLp6_0(.dout(w_dff_A_DGYHpj5P7_0),.din(w_dff_A_bh2APSLp6_0),.clk(gclk));
	jdff dff_A_DGYHpj5P7_0(.dout(w_dff_A_8TK6d1gG5_0),.din(w_dff_A_DGYHpj5P7_0),.clk(gclk));
	jdff dff_A_8TK6d1gG5_0(.dout(w_dff_A_sHry7NyT4_0),.din(w_dff_A_8TK6d1gG5_0),.clk(gclk));
	jdff dff_A_sHry7NyT4_0(.dout(w_dff_A_IeOFZFFC1_0),.din(w_dff_A_sHry7NyT4_0),.clk(gclk));
	jdff dff_A_IeOFZFFC1_0(.dout(w_dff_A_4eZgLYV21_0),.din(w_dff_A_IeOFZFFC1_0),.clk(gclk));
	jdff dff_A_4eZgLYV21_0(.dout(w_dff_A_HXmEf8aN3_0),.din(w_dff_A_4eZgLYV21_0),.clk(gclk));
	jdff dff_A_HXmEf8aN3_0(.dout(w_dff_A_KNF8iGyM1_0),.din(w_dff_A_HXmEf8aN3_0),.clk(gclk));
	jdff dff_A_KNF8iGyM1_0(.dout(w_dff_A_pPliMtAK0_0),.din(w_dff_A_KNF8iGyM1_0),.clk(gclk));
	jdff dff_A_pPliMtAK0_0(.dout(w_dff_A_qSsHN3Ix4_0),.din(w_dff_A_pPliMtAK0_0),.clk(gclk));
	jdff dff_A_qSsHN3Ix4_0(.dout(w_dff_A_Ed2k6v438_0),.din(w_dff_A_qSsHN3Ix4_0),.clk(gclk));
	jdff dff_A_Ed2k6v438_0(.dout(w_dff_A_8rgolz4m2_0),.din(w_dff_A_Ed2k6v438_0),.clk(gclk));
	jdff dff_A_8rgolz4m2_0(.dout(w_dff_A_tLr9nbjR6_0),.din(w_dff_A_8rgolz4m2_0),.clk(gclk));
	jdff dff_A_tLr9nbjR6_0(.dout(w_dff_A_x3AzODmj5_0),.din(w_dff_A_tLr9nbjR6_0),.clk(gclk));
	jdff dff_A_x3AzODmj5_0(.dout(w_dff_A_QfUUn8bN6_0),.din(w_dff_A_x3AzODmj5_0),.clk(gclk));
	jdff dff_A_QfUUn8bN6_0(.dout(w_dff_A_4HLVI9dQ5_0),.din(w_dff_A_QfUUn8bN6_0),.clk(gclk));
	jdff dff_A_4HLVI9dQ5_0(.dout(w_dff_A_4s8PTElj1_0),.din(w_dff_A_4HLVI9dQ5_0),.clk(gclk));
	jdff dff_A_4s8PTElj1_0(.dout(w_dff_A_IAgpnSlD3_0),.din(w_dff_A_4s8PTElj1_0),.clk(gclk));
	jdff dff_A_IAgpnSlD3_0(.dout(w_dff_A_yUAUJ1wR1_0),.din(w_dff_A_IAgpnSlD3_0),.clk(gclk));
	jdff dff_A_yUAUJ1wR1_0(.dout(w_dff_A_xSNHOa6j7_0),.din(w_dff_A_yUAUJ1wR1_0),.clk(gclk));
	jdff dff_A_xSNHOa6j7_0(.dout(w_dff_A_29fDN8L70_0),.din(w_dff_A_xSNHOa6j7_0),.clk(gclk));
	jdff dff_A_29fDN8L70_0(.dout(w_dff_A_tIPN73wT6_0),.din(w_dff_A_29fDN8L70_0),.clk(gclk));
	jdff dff_A_tIPN73wT6_0(.dout(w_dff_A_Efcch7jW2_0),.din(w_dff_A_tIPN73wT6_0),.clk(gclk));
	jdff dff_A_Efcch7jW2_0(.dout(w_dff_A_xkCiVbQh7_0),.din(w_dff_A_Efcch7jW2_0),.clk(gclk));
	jdff dff_A_xkCiVbQh7_0(.dout(w_dff_A_y6ohbpy86_0),.din(w_dff_A_xkCiVbQh7_0),.clk(gclk));
	jdff dff_A_y6ohbpy86_0(.dout(w_dff_A_jQkCx8Dp7_0),.din(w_dff_A_y6ohbpy86_0),.clk(gclk));
	jdff dff_A_jQkCx8Dp7_0(.dout(w_dff_A_O4CF5uWf1_0),.din(w_dff_A_jQkCx8Dp7_0),.clk(gclk));
	jdff dff_A_O4CF5uWf1_0(.dout(w_dff_A_yb2Ku54r4_0),.din(w_dff_A_O4CF5uWf1_0),.clk(gclk));
	jdff dff_A_yb2Ku54r4_0(.dout(w_dff_A_kEJvZqUP9_0),.din(w_dff_A_yb2Ku54r4_0),.clk(gclk));
	jdff dff_A_kEJvZqUP9_0(.dout(w_dff_A_YxJMjaIZ1_0),.din(w_dff_A_kEJvZqUP9_0),.clk(gclk));
	jdff dff_A_YxJMjaIZ1_0(.dout(w_dff_A_JXwZ7n5C8_0),.din(w_dff_A_YxJMjaIZ1_0),.clk(gclk));
	jdff dff_A_JXwZ7n5C8_0(.dout(w_dff_A_GQ0A3ISV9_0),.din(w_dff_A_JXwZ7n5C8_0),.clk(gclk));
	jdff dff_A_GQ0A3ISV9_0(.dout(w_dff_A_PKYKLMPJ9_0),.din(w_dff_A_GQ0A3ISV9_0),.clk(gclk));
	jdff dff_A_PKYKLMPJ9_0(.dout(w_dff_A_w2qDXOxp3_0),.din(w_dff_A_PKYKLMPJ9_0),.clk(gclk));
	jdff dff_A_w2qDXOxp3_0(.dout(w_dff_A_rhiqZhER5_0),.din(w_dff_A_w2qDXOxp3_0),.clk(gclk));
	jdff dff_A_rhiqZhER5_0(.dout(w_dff_A_OaFrd7Qy4_0),.din(w_dff_A_rhiqZhER5_0),.clk(gclk));
	jdff dff_A_OaFrd7Qy4_0(.dout(w_dff_A_MB4GHscJ8_0),.din(w_dff_A_OaFrd7Qy4_0),.clk(gclk));
	jdff dff_A_MB4GHscJ8_0(.dout(w_dff_A_RzZ07c8e1_0),.din(w_dff_A_MB4GHscJ8_0),.clk(gclk));
	jdff dff_A_RzZ07c8e1_0(.dout(w_dff_A_5Fx9KCuE9_0),.din(w_dff_A_RzZ07c8e1_0),.clk(gclk));
	jdff dff_A_5Fx9KCuE9_0(.dout(w_dff_A_D37uXOCo7_0),.din(w_dff_A_5Fx9KCuE9_0),.clk(gclk));
	jdff dff_A_D37uXOCo7_0(.dout(w_dff_A_1nID5NdP6_0),.din(w_dff_A_D37uXOCo7_0),.clk(gclk));
	jdff dff_A_1nID5NdP6_0(.dout(w_dff_A_OoY8hnye1_0),.din(w_dff_A_1nID5NdP6_0),.clk(gclk));
	jdff dff_A_OoY8hnye1_0(.dout(w_dff_A_XUsa8Kup5_0),.din(w_dff_A_OoY8hnye1_0),.clk(gclk));
	jdff dff_A_XUsa8Kup5_0(.dout(w_dff_A_DWsRDCbR6_0),.din(w_dff_A_XUsa8Kup5_0),.clk(gclk));
	jdff dff_A_DWsRDCbR6_0(.dout(w_dff_A_9gCRsJK16_0),.din(w_dff_A_DWsRDCbR6_0),.clk(gclk));
	jdff dff_A_9gCRsJK16_0(.dout(w_dff_A_PzUR5csb4_0),.din(w_dff_A_9gCRsJK16_0),.clk(gclk));
	jdff dff_A_PzUR5csb4_0(.dout(w_dff_A_Qvmd2M0y3_0),.din(w_dff_A_PzUR5csb4_0),.clk(gclk));
	jdff dff_A_Qvmd2M0y3_0(.dout(w_dff_A_vBQUKRdX7_0),.din(w_dff_A_Qvmd2M0y3_0),.clk(gclk));
	jdff dff_A_vBQUKRdX7_0(.dout(w_dff_A_cu0Bw0H98_0),.din(w_dff_A_vBQUKRdX7_0),.clk(gclk));
	jdff dff_A_cu0Bw0H98_0(.dout(w_dff_A_5IdgGGfG5_0),.din(w_dff_A_cu0Bw0H98_0),.clk(gclk));
	jdff dff_A_5IdgGGfG5_0(.dout(w_dff_A_8GlWDUqT0_0),.din(w_dff_A_5IdgGGfG5_0),.clk(gclk));
	jdff dff_A_8GlWDUqT0_0(.dout(w_dff_A_x1Lz4r392_0),.din(w_dff_A_8GlWDUqT0_0),.clk(gclk));
	jdff dff_A_x1Lz4r392_0(.dout(w_dff_A_sjG6wrnR9_0),.din(w_dff_A_x1Lz4r392_0),.clk(gclk));
	jdff dff_A_sjG6wrnR9_0(.dout(w_dff_A_K1mxTCAS4_0),.din(w_dff_A_sjG6wrnR9_0),.clk(gclk));
	jdff dff_A_K1mxTCAS4_0(.dout(w_dff_A_FNChFH696_0),.din(w_dff_A_K1mxTCAS4_0),.clk(gclk));
	jdff dff_A_FNChFH696_0(.dout(G2548gat),.din(w_dff_A_FNChFH696_0),.clk(gclk));
	jdff dff_A_vopQHw7W8_2(.dout(w_dff_A_mFoBwehz9_0),.din(w_dff_A_vopQHw7W8_2),.clk(gclk));
	jdff dff_A_mFoBwehz9_0(.dout(w_dff_A_lpEAnQPX0_0),.din(w_dff_A_mFoBwehz9_0),.clk(gclk));
	jdff dff_A_lpEAnQPX0_0(.dout(w_dff_A_k1XBAUvs0_0),.din(w_dff_A_lpEAnQPX0_0),.clk(gclk));
	jdff dff_A_k1XBAUvs0_0(.dout(w_dff_A_aDnyrkFj7_0),.din(w_dff_A_k1XBAUvs0_0),.clk(gclk));
	jdff dff_A_aDnyrkFj7_0(.dout(w_dff_A_8aONQoL34_0),.din(w_dff_A_aDnyrkFj7_0),.clk(gclk));
	jdff dff_A_8aONQoL34_0(.dout(w_dff_A_I6kKjmlw7_0),.din(w_dff_A_8aONQoL34_0),.clk(gclk));
	jdff dff_A_I6kKjmlw7_0(.dout(w_dff_A_9ddu3VGz6_0),.din(w_dff_A_I6kKjmlw7_0),.clk(gclk));
	jdff dff_A_9ddu3VGz6_0(.dout(w_dff_A_uFeY0ZwY9_0),.din(w_dff_A_9ddu3VGz6_0),.clk(gclk));
	jdff dff_A_uFeY0ZwY9_0(.dout(w_dff_A_vrqJFr1D4_0),.din(w_dff_A_uFeY0ZwY9_0),.clk(gclk));
	jdff dff_A_vrqJFr1D4_0(.dout(w_dff_A_mj9nnrBL8_0),.din(w_dff_A_vrqJFr1D4_0),.clk(gclk));
	jdff dff_A_mj9nnrBL8_0(.dout(w_dff_A_nAKHURSR4_0),.din(w_dff_A_mj9nnrBL8_0),.clk(gclk));
	jdff dff_A_nAKHURSR4_0(.dout(w_dff_A_WAmUxhqR9_0),.din(w_dff_A_nAKHURSR4_0),.clk(gclk));
	jdff dff_A_WAmUxhqR9_0(.dout(w_dff_A_iy2miqlv3_0),.din(w_dff_A_WAmUxhqR9_0),.clk(gclk));
	jdff dff_A_iy2miqlv3_0(.dout(w_dff_A_31IDM0L67_0),.din(w_dff_A_iy2miqlv3_0),.clk(gclk));
	jdff dff_A_31IDM0L67_0(.dout(w_dff_A_uUYaAqXH4_0),.din(w_dff_A_31IDM0L67_0),.clk(gclk));
	jdff dff_A_uUYaAqXH4_0(.dout(w_dff_A_yRdRrBuj7_0),.din(w_dff_A_uUYaAqXH4_0),.clk(gclk));
	jdff dff_A_yRdRrBuj7_0(.dout(w_dff_A_pWk8ihPO5_0),.din(w_dff_A_yRdRrBuj7_0),.clk(gclk));
	jdff dff_A_pWk8ihPO5_0(.dout(w_dff_A_SrPpZCxu8_0),.din(w_dff_A_pWk8ihPO5_0),.clk(gclk));
	jdff dff_A_SrPpZCxu8_0(.dout(w_dff_A_YxRUQL8A5_0),.din(w_dff_A_SrPpZCxu8_0),.clk(gclk));
	jdff dff_A_YxRUQL8A5_0(.dout(w_dff_A_xFDMzeuG3_0),.din(w_dff_A_YxRUQL8A5_0),.clk(gclk));
	jdff dff_A_xFDMzeuG3_0(.dout(w_dff_A_Wss4OJSK2_0),.din(w_dff_A_xFDMzeuG3_0),.clk(gclk));
	jdff dff_A_Wss4OJSK2_0(.dout(w_dff_A_tbOMpMK81_0),.din(w_dff_A_Wss4OJSK2_0),.clk(gclk));
	jdff dff_A_tbOMpMK81_0(.dout(w_dff_A_dkf8Q8G94_0),.din(w_dff_A_tbOMpMK81_0),.clk(gclk));
	jdff dff_A_dkf8Q8G94_0(.dout(w_dff_A_tKwFEqj33_0),.din(w_dff_A_dkf8Q8G94_0),.clk(gclk));
	jdff dff_A_tKwFEqj33_0(.dout(w_dff_A_aDsSbgmo4_0),.din(w_dff_A_tKwFEqj33_0),.clk(gclk));
	jdff dff_A_aDsSbgmo4_0(.dout(w_dff_A_EgsBPe6D2_0),.din(w_dff_A_aDsSbgmo4_0),.clk(gclk));
	jdff dff_A_EgsBPe6D2_0(.dout(w_dff_A_SZ00c0SZ2_0),.din(w_dff_A_EgsBPe6D2_0),.clk(gclk));
	jdff dff_A_SZ00c0SZ2_0(.dout(w_dff_A_TwVRXF2y6_0),.din(w_dff_A_SZ00c0SZ2_0),.clk(gclk));
	jdff dff_A_TwVRXF2y6_0(.dout(w_dff_A_jGUshw0S7_0),.din(w_dff_A_TwVRXF2y6_0),.clk(gclk));
	jdff dff_A_jGUshw0S7_0(.dout(w_dff_A_BXzfYPKT0_0),.din(w_dff_A_jGUshw0S7_0),.clk(gclk));
	jdff dff_A_BXzfYPKT0_0(.dout(w_dff_A_6M4fPLVj7_0),.din(w_dff_A_BXzfYPKT0_0),.clk(gclk));
	jdff dff_A_6M4fPLVj7_0(.dout(w_dff_A_DnJ8TZiW0_0),.din(w_dff_A_6M4fPLVj7_0),.clk(gclk));
	jdff dff_A_DnJ8TZiW0_0(.dout(w_dff_A_iOdFmewz0_0),.din(w_dff_A_DnJ8TZiW0_0),.clk(gclk));
	jdff dff_A_iOdFmewz0_0(.dout(w_dff_A_OzQ2Ebdd0_0),.din(w_dff_A_iOdFmewz0_0),.clk(gclk));
	jdff dff_A_OzQ2Ebdd0_0(.dout(w_dff_A_WOJr8laE8_0),.din(w_dff_A_OzQ2Ebdd0_0),.clk(gclk));
	jdff dff_A_WOJr8laE8_0(.dout(w_dff_A_8AFyvlss7_0),.din(w_dff_A_WOJr8laE8_0),.clk(gclk));
	jdff dff_A_8AFyvlss7_0(.dout(w_dff_A_IpUk4VZL0_0),.din(w_dff_A_8AFyvlss7_0),.clk(gclk));
	jdff dff_A_IpUk4VZL0_0(.dout(w_dff_A_z5vgm3J21_0),.din(w_dff_A_IpUk4VZL0_0),.clk(gclk));
	jdff dff_A_z5vgm3J21_0(.dout(w_dff_A_jOe6T4Zy3_0),.din(w_dff_A_z5vgm3J21_0),.clk(gclk));
	jdff dff_A_jOe6T4Zy3_0(.dout(w_dff_A_uMbOQooM9_0),.din(w_dff_A_jOe6T4Zy3_0),.clk(gclk));
	jdff dff_A_uMbOQooM9_0(.dout(w_dff_A_6y1SwXfO1_0),.din(w_dff_A_uMbOQooM9_0),.clk(gclk));
	jdff dff_A_6y1SwXfO1_0(.dout(w_dff_A_kI8w5MOE7_0),.din(w_dff_A_6y1SwXfO1_0),.clk(gclk));
	jdff dff_A_kI8w5MOE7_0(.dout(w_dff_A_b4Nm84XW8_0),.din(w_dff_A_kI8w5MOE7_0),.clk(gclk));
	jdff dff_A_b4Nm84XW8_0(.dout(w_dff_A_zRsSBkzh1_0),.din(w_dff_A_b4Nm84XW8_0),.clk(gclk));
	jdff dff_A_zRsSBkzh1_0(.dout(w_dff_A_Mg9D5fXL3_0),.din(w_dff_A_zRsSBkzh1_0),.clk(gclk));
	jdff dff_A_Mg9D5fXL3_0(.dout(w_dff_A_kjm8Wqfw8_0),.din(w_dff_A_Mg9D5fXL3_0),.clk(gclk));
	jdff dff_A_kjm8Wqfw8_0(.dout(w_dff_A_b0En7ZcL2_0),.din(w_dff_A_kjm8Wqfw8_0),.clk(gclk));
	jdff dff_A_b0En7ZcL2_0(.dout(w_dff_A_9vZ9g4sh5_0),.din(w_dff_A_b0En7ZcL2_0),.clk(gclk));
	jdff dff_A_9vZ9g4sh5_0(.dout(w_dff_A_UFs2y91Z8_0),.din(w_dff_A_9vZ9g4sh5_0),.clk(gclk));
	jdff dff_A_UFs2y91Z8_0(.dout(w_dff_A_4OtmtBbg9_0),.din(w_dff_A_UFs2y91Z8_0),.clk(gclk));
	jdff dff_A_4OtmtBbg9_0(.dout(w_dff_A_SGeC2zRk4_0),.din(w_dff_A_4OtmtBbg9_0),.clk(gclk));
	jdff dff_A_SGeC2zRk4_0(.dout(w_dff_A_Lo1pvlvF9_0),.din(w_dff_A_SGeC2zRk4_0),.clk(gclk));
	jdff dff_A_Lo1pvlvF9_0(.dout(w_dff_A_jmE8YK7I1_0),.din(w_dff_A_Lo1pvlvF9_0),.clk(gclk));
	jdff dff_A_jmE8YK7I1_0(.dout(w_dff_A_cPWEKegT1_0),.din(w_dff_A_jmE8YK7I1_0),.clk(gclk));
	jdff dff_A_cPWEKegT1_0(.dout(w_dff_A_iWmkvgPp6_0),.din(w_dff_A_cPWEKegT1_0),.clk(gclk));
	jdff dff_A_iWmkvgPp6_0(.dout(w_dff_A_0zhb5H5M3_0),.din(w_dff_A_iWmkvgPp6_0),.clk(gclk));
	jdff dff_A_0zhb5H5M3_0(.dout(w_dff_A_cfY3Mtns9_0),.din(w_dff_A_0zhb5H5M3_0),.clk(gclk));
	jdff dff_A_cfY3Mtns9_0(.dout(w_dff_A_9MDZ3hWf6_0),.din(w_dff_A_cfY3Mtns9_0),.clk(gclk));
	jdff dff_A_9MDZ3hWf6_0(.dout(w_dff_A_6RkZudg36_0),.din(w_dff_A_9MDZ3hWf6_0),.clk(gclk));
	jdff dff_A_6RkZudg36_0(.dout(G2877gat),.din(w_dff_A_6RkZudg36_0),.clk(gclk));
	jdff dff_A_xPsKA8QQ4_2(.dout(w_dff_A_VtaktCyZ6_0),.din(w_dff_A_xPsKA8QQ4_2),.clk(gclk));
	jdff dff_A_VtaktCyZ6_0(.dout(w_dff_A_TpZoPvat8_0),.din(w_dff_A_VtaktCyZ6_0),.clk(gclk));
	jdff dff_A_TpZoPvat8_0(.dout(w_dff_A_tNbZIGhQ7_0),.din(w_dff_A_TpZoPvat8_0),.clk(gclk));
	jdff dff_A_tNbZIGhQ7_0(.dout(w_dff_A_HRd7yJal4_0),.din(w_dff_A_tNbZIGhQ7_0),.clk(gclk));
	jdff dff_A_HRd7yJal4_0(.dout(w_dff_A_zIfZ8yh84_0),.din(w_dff_A_HRd7yJal4_0),.clk(gclk));
	jdff dff_A_zIfZ8yh84_0(.dout(w_dff_A_mHBE1IYC9_0),.din(w_dff_A_zIfZ8yh84_0),.clk(gclk));
	jdff dff_A_mHBE1IYC9_0(.dout(w_dff_A_IrB2qO3r4_0),.din(w_dff_A_mHBE1IYC9_0),.clk(gclk));
	jdff dff_A_IrB2qO3r4_0(.dout(w_dff_A_eJ66f0YT0_0),.din(w_dff_A_IrB2qO3r4_0),.clk(gclk));
	jdff dff_A_eJ66f0YT0_0(.dout(w_dff_A_nhzZEO2k6_0),.din(w_dff_A_eJ66f0YT0_0),.clk(gclk));
	jdff dff_A_nhzZEO2k6_0(.dout(w_dff_A_ddUKiAET7_0),.din(w_dff_A_nhzZEO2k6_0),.clk(gclk));
	jdff dff_A_ddUKiAET7_0(.dout(w_dff_A_ZvWBmQti6_0),.din(w_dff_A_ddUKiAET7_0),.clk(gclk));
	jdff dff_A_ZvWBmQti6_0(.dout(w_dff_A_0tMGJ2us5_0),.din(w_dff_A_ZvWBmQti6_0),.clk(gclk));
	jdff dff_A_0tMGJ2us5_0(.dout(w_dff_A_uuxNTB2n0_0),.din(w_dff_A_0tMGJ2us5_0),.clk(gclk));
	jdff dff_A_uuxNTB2n0_0(.dout(w_dff_A_dSX1gFKq9_0),.din(w_dff_A_uuxNTB2n0_0),.clk(gclk));
	jdff dff_A_dSX1gFKq9_0(.dout(w_dff_A_L4P54gpI0_0),.din(w_dff_A_dSX1gFKq9_0),.clk(gclk));
	jdff dff_A_L4P54gpI0_0(.dout(w_dff_A_9uzdJkUP9_0),.din(w_dff_A_L4P54gpI0_0),.clk(gclk));
	jdff dff_A_9uzdJkUP9_0(.dout(w_dff_A_yiuPU3LY2_0),.din(w_dff_A_9uzdJkUP9_0),.clk(gclk));
	jdff dff_A_yiuPU3LY2_0(.dout(w_dff_A_LQfmxIMN5_0),.din(w_dff_A_yiuPU3LY2_0),.clk(gclk));
	jdff dff_A_LQfmxIMN5_0(.dout(w_dff_A_1QeAzK8O0_0),.din(w_dff_A_LQfmxIMN5_0),.clk(gclk));
	jdff dff_A_1QeAzK8O0_0(.dout(w_dff_A_ZirUxbJy9_0),.din(w_dff_A_1QeAzK8O0_0),.clk(gclk));
	jdff dff_A_ZirUxbJy9_0(.dout(w_dff_A_a9z1lfKH1_0),.din(w_dff_A_ZirUxbJy9_0),.clk(gclk));
	jdff dff_A_a9z1lfKH1_0(.dout(w_dff_A_BCRZdo1t0_0),.din(w_dff_A_a9z1lfKH1_0),.clk(gclk));
	jdff dff_A_BCRZdo1t0_0(.dout(w_dff_A_y5odsYue8_0),.din(w_dff_A_BCRZdo1t0_0),.clk(gclk));
	jdff dff_A_y5odsYue8_0(.dout(w_dff_A_etjNtSsz3_0),.din(w_dff_A_y5odsYue8_0),.clk(gclk));
	jdff dff_A_etjNtSsz3_0(.dout(w_dff_A_fsiO41dQ7_0),.din(w_dff_A_etjNtSsz3_0),.clk(gclk));
	jdff dff_A_fsiO41dQ7_0(.dout(w_dff_A_SxwruHad3_0),.din(w_dff_A_fsiO41dQ7_0),.clk(gclk));
	jdff dff_A_SxwruHad3_0(.dout(w_dff_A_NLAVcwWt9_0),.din(w_dff_A_SxwruHad3_0),.clk(gclk));
	jdff dff_A_NLAVcwWt9_0(.dout(w_dff_A_21jvGW8Y0_0),.din(w_dff_A_NLAVcwWt9_0),.clk(gclk));
	jdff dff_A_21jvGW8Y0_0(.dout(w_dff_A_BjOUEZux0_0),.din(w_dff_A_21jvGW8Y0_0),.clk(gclk));
	jdff dff_A_BjOUEZux0_0(.dout(w_dff_A_0euBjbWc6_0),.din(w_dff_A_BjOUEZux0_0),.clk(gclk));
	jdff dff_A_0euBjbWc6_0(.dout(w_dff_A_EKGJ3hDJ1_0),.din(w_dff_A_0euBjbWc6_0),.clk(gclk));
	jdff dff_A_EKGJ3hDJ1_0(.dout(w_dff_A_WpFJcSxo9_0),.din(w_dff_A_EKGJ3hDJ1_0),.clk(gclk));
	jdff dff_A_WpFJcSxo9_0(.dout(w_dff_A_0DEEoLFt8_0),.din(w_dff_A_WpFJcSxo9_0),.clk(gclk));
	jdff dff_A_0DEEoLFt8_0(.dout(w_dff_A_3CxfT8b73_0),.din(w_dff_A_0DEEoLFt8_0),.clk(gclk));
	jdff dff_A_3CxfT8b73_0(.dout(w_dff_A_fOrt9ejS3_0),.din(w_dff_A_3CxfT8b73_0),.clk(gclk));
	jdff dff_A_fOrt9ejS3_0(.dout(w_dff_A_I3sMw07c3_0),.din(w_dff_A_fOrt9ejS3_0),.clk(gclk));
	jdff dff_A_I3sMw07c3_0(.dout(w_dff_A_3yLcQN5i9_0),.din(w_dff_A_I3sMw07c3_0),.clk(gclk));
	jdff dff_A_3yLcQN5i9_0(.dout(w_dff_A_goBP1uOm8_0),.din(w_dff_A_3yLcQN5i9_0),.clk(gclk));
	jdff dff_A_goBP1uOm8_0(.dout(w_dff_A_9HQ5FCA44_0),.din(w_dff_A_goBP1uOm8_0),.clk(gclk));
	jdff dff_A_9HQ5FCA44_0(.dout(w_dff_A_oqiLpstc0_0),.din(w_dff_A_9HQ5FCA44_0),.clk(gclk));
	jdff dff_A_oqiLpstc0_0(.dout(w_dff_A_CxWcVPBl4_0),.din(w_dff_A_oqiLpstc0_0),.clk(gclk));
	jdff dff_A_CxWcVPBl4_0(.dout(w_dff_A_SJkGpVdc0_0),.din(w_dff_A_CxWcVPBl4_0),.clk(gclk));
	jdff dff_A_SJkGpVdc0_0(.dout(w_dff_A_jmZeOd3P8_0),.din(w_dff_A_SJkGpVdc0_0),.clk(gclk));
	jdff dff_A_jmZeOd3P8_0(.dout(w_dff_A_PxTx5HK61_0),.din(w_dff_A_jmZeOd3P8_0),.clk(gclk));
	jdff dff_A_PxTx5HK61_0(.dout(w_dff_A_aqfX5RqX1_0),.din(w_dff_A_PxTx5HK61_0),.clk(gclk));
	jdff dff_A_aqfX5RqX1_0(.dout(w_dff_A_Ulav9pLt5_0),.din(w_dff_A_aqfX5RqX1_0),.clk(gclk));
	jdff dff_A_Ulav9pLt5_0(.dout(w_dff_A_UKs76Q702_0),.din(w_dff_A_Ulav9pLt5_0),.clk(gclk));
	jdff dff_A_UKs76Q702_0(.dout(w_dff_A_KQWdSDpY3_0),.din(w_dff_A_UKs76Q702_0),.clk(gclk));
	jdff dff_A_KQWdSDpY3_0(.dout(w_dff_A_RQzzZAYD7_0),.din(w_dff_A_KQWdSDpY3_0),.clk(gclk));
	jdff dff_A_RQzzZAYD7_0(.dout(w_dff_A_a41ksy7G6_0),.din(w_dff_A_RQzzZAYD7_0),.clk(gclk));
	jdff dff_A_a41ksy7G6_0(.dout(w_dff_A_fn4jRplA1_0),.din(w_dff_A_a41ksy7G6_0),.clk(gclk));
	jdff dff_A_fn4jRplA1_0(.dout(w_dff_A_FChtwYNV6_0),.din(w_dff_A_fn4jRplA1_0),.clk(gclk));
	jdff dff_A_FChtwYNV6_0(.dout(w_dff_A_Km7j8Yhc0_0),.din(w_dff_A_FChtwYNV6_0),.clk(gclk));
	jdff dff_A_Km7j8Yhc0_0(.dout(w_dff_A_wF9lnkhh2_0),.din(w_dff_A_Km7j8Yhc0_0),.clk(gclk));
	jdff dff_A_wF9lnkhh2_0(.dout(w_dff_A_hyne3PJx7_0),.din(w_dff_A_wF9lnkhh2_0),.clk(gclk));
	jdff dff_A_hyne3PJx7_0(.dout(w_dff_A_r2P9juUz5_0),.din(w_dff_A_hyne3PJx7_0),.clk(gclk));
	jdff dff_A_r2P9juUz5_0(.dout(G3211gat),.din(w_dff_A_r2P9juUz5_0),.clk(gclk));
	jdff dff_A_ByNtDrk64_2(.dout(w_dff_A_MOy45Gta4_0),.din(w_dff_A_ByNtDrk64_2),.clk(gclk));
	jdff dff_A_MOy45Gta4_0(.dout(w_dff_A_5Tx3mpaO2_0),.din(w_dff_A_MOy45Gta4_0),.clk(gclk));
	jdff dff_A_5Tx3mpaO2_0(.dout(w_dff_A_8TC1SORo5_0),.din(w_dff_A_5Tx3mpaO2_0),.clk(gclk));
	jdff dff_A_8TC1SORo5_0(.dout(w_dff_A_onfZaWLE0_0),.din(w_dff_A_8TC1SORo5_0),.clk(gclk));
	jdff dff_A_onfZaWLE0_0(.dout(w_dff_A_aVugbHoH2_0),.din(w_dff_A_onfZaWLE0_0),.clk(gclk));
	jdff dff_A_aVugbHoH2_0(.dout(w_dff_A_ghdKFs9E3_0),.din(w_dff_A_aVugbHoH2_0),.clk(gclk));
	jdff dff_A_ghdKFs9E3_0(.dout(w_dff_A_cOxkFxM15_0),.din(w_dff_A_ghdKFs9E3_0),.clk(gclk));
	jdff dff_A_cOxkFxM15_0(.dout(w_dff_A_s1VdefxO8_0),.din(w_dff_A_cOxkFxM15_0),.clk(gclk));
	jdff dff_A_s1VdefxO8_0(.dout(w_dff_A_GqlkSCUu6_0),.din(w_dff_A_s1VdefxO8_0),.clk(gclk));
	jdff dff_A_GqlkSCUu6_0(.dout(w_dff_A_y6rU666g2_0),.din(w_dff_A_GqlkSCUu6_0),.clk(gclk));
	jdff dff_A_y6rU666g2_0(.dout(w_dff_A_KqlqJ8e55_0),.din(w_dff_A_y6rU666g2_0),.clk(gclk));
	jdff dff_A_KqlqJ8e55_0(.dout(w_dff_A_BjBnoNwL7_0),.din(w_dff_A_KqlqJ8e55_0),.clk(gclk));
	jdff dff_A_BjBnoNwL7_0(.dout(w_dff_A_h9whmFh97_0),.din(w_dff_A_BjBnoNwL7_0),.clk(gclk));
	jdff dff_A_h9whmFh97_0(.dout(w_dff_A_pxFwMPUY1_0),.din(w_dff_A_h9whmFh97_0),.clk(gclk));
	jdff dff_A_pxFwMPUY1_0(.dout(w_dff_A_qeH9taZC0_0),.din(w_dff_A_pxFwMPUY1_0),.clk(gclk));
	jdff dff_A_qeH9taZC0_0(.dout(w_dff_A_vmW6vxdh5_0),.din(w_dff_A_qeH9taZC0_0),.clk(gclk));
	jdff dff_A_vmW6vxdh5_0(.dout(w_dff_A_Ayckzlpl6_0),.din(w_dff_A_vmW6vxdh5_0),.clk(gclk));
	jdff dff_A_Ayckzlpl6_0(.dout(w_dff_A_pIwsWaUa8_0),.din(w_dff_A_Ayckzlpl6_0),.clk(gclk));
	jdff dff_A_pIwsWaUa8_0(.dout(w_dff_A_O8hG4fWQ0_0),.din(w_dff_A_pIwsWaUa8_0),.clk(gclk));
	jdff dff_A_O8hG4fWQ0_0(.dout(w_dff_A_Q5jClSu92_0),.din(w_dff_A_O8hG4fWQ0_0),.clk(gclk));
	jdff dff_A_Q5jClSu92_0(.dout(w_dff_A_Lns7Ijju7_0),.din(w_dff_A_Q5jClSu92_0),.clk(gclk));
	jdff dff_A_Lns7Ijju7_0(.dout(w_dff_A_uWQ2yjvK6_0),.din(w_dff_A_Lns7Ijju7_0),.clk(gclk));
	jdff dff_A_uWQ2yjvK6_0(.dout(w_dff_A_KMyGcg4b7_0),.din(w_dff_A_uWQ2yjvK6_0),.clk(gclk));
	jdff dff_A_KMyGcg4b7_0(.dout(w_dff_A_G45DwoiU0_0),.din(w_dff_A_KMyGcg4b7_0),.clk(gclk));
	jdff dff_A_G45DwoiU0_0(.dout(w_dff_A_9qtxAklF2_0),.din(w_dff_A_G45DwoiU0_0),.clk(gclk));
	jdff dff_A_9qtxAklF2_0(.dout(w_dff_A_qnEAhHQt3_0),.din(w_dff_A_9qtxAklF2_0),.clk(gclk));
	jdff dff_A_qnEAhHQt3_0(.dout(w_dff_A_pIaS6yfF6_0),.din(w_dff_A_qnEAhHQt3_0),.clk(gclk));
	jdff dff_A_pIaS6yfF6_0(.dout(w_dff_A_y4X44ksk0_0),.din(w_dff_A_pIaS6yfF6_0),.clk(gclk));
	jdff dff_A_y4X44ksk0_0(.dout(w_dff_A_RwLuFJSC5_0),.din(w_dff_A_y4X44ksk0_0),.clk(gclk));
	jdff dff_A_RwLuFJSC5_0(.dout(w_dff_A_2PPGMt3j5_0),.din(w_dff_A_RwLuFJSC5_0),.clk(gclk));
	jdff dff_A_2PPGMt3j5_0(.dout(w_dff_A_FFA0ajUg8_0),.din(w_dff_A_2PPGMt3j5_0),.clk(gclk));
	jdff dff_A_FFA0ajUg8_0(.dout(w_dff_A_r9hNANWG7_0),.din(w_dff_A_FFA0ajUg8_0),.clk(gclk));
	jdff dff_A_r9hNANWG7_0(.dout(w_dff_A_yB5jntl06_0),.din(w_dff_A_r9hNANWG7_0),.clk(gclk));
	jdff dff_A_yB5jntl06_0(.dout(w_dff_A_vSW29hvO5_0),.din(w_dff_A_yB5jntl06_0),.clk(gclk));
	jdff dff_A_vSW29hvO5_0(.dout(w_dff_A_ghCvYGAd8_0),.din(w_dff_A_vSW29hvO5_0),.clk(gclk));
	jdff dff_A_ghCvYGAd8_0(.dout(w_dff_A_GbNOzueq6_0),.din(w_dff_A_ghCvYGAd8_0),.clk(gclk));
	jdff dff_A_GbNOzueq6_0(.dout(w_dff_A_QJRJU3N02_0),.din(w_dff_A_GbNOzueq6_0),.clk(gclk));
	jdff dff_A_QJRJU3N02_0(.dout(w_dff_A_yXVuvWgT5_0),.din(w_dff_A_QJRJU3N02_0),.clk(gclk));
	jdff dff_A_yXVuvWgT5_0(.dout(w_dff_A_9Qz7LQBP5_0),.din(w_dff_A_yXVuvWgT5_0),.clk(gclk));
	jdff dff_A_9Qz7LQBP5_0(.dout(w_dff_A_TmM8lxpT3_0),.din(w_dff_A_9Qz7LQBP5_0),.clk(gclk));
	jdff dff_A_TmM8lxpT3_0(.dout(w_dff_A_qLkWJwRB1_0),.din(w_dff_A_TmM8lxpT3_0),.clk(gclk));
	jdff dff_A_qLkWJwRB1_0(.dout(w_dff_A_krxee2Uc9_0),.din(w_dff_A_qLkWJwRB1_0),.clk(gclk));
	jdff dff_A_krxee2Uc9_0(.dout(w_dff_A_UfKtTvOK1_0),.din(w_dff_A_krxee2Uc9_0),.clk(gclk));
	jdff dff_A_UfKtTvOK1_0(.dout(w_dff_A_AWGoDzqR1_0),.din(w_dff_A_UfKtTvOK1_0),.clk(gclk));
	jdff dff_A_AWGoDzqR1_0(.dout(w_dff_A_vxcXAnTc6_0),.din(w_dff_A_AWGoDzqR1_0),.clk(gclk));
	jdff dff_A_vxcXAnTc6_0(.dout(w_dff_A_6902Kq5q3_0),.din(w_dff_A_vxcXAnTc6_0),.clk(gclk));
	jdff dff_A_6902Kq5q3_0(.dout(w_dff_A_0zMcmGsi4_0),.din(w_dff_A_6902Kq5q3_0),.clk(gclk));
	jdff dff_A_0zMcmGsi4_0(.dout(w_dff_A_mTmxVBjj2_0),.din(w_dff_A_0zMcmGsi4_0),.clk(gclk));
	jdff dff_A_mTmxVBjj2_0(.dout(w_dff_A_J4dk22Yl9_0),.din(w_dff_A_mTmxVBjj2_0),.clk(gclk));
	jdff dff_A_J4dk22Yl9_0(.dout(w_dff_A_4CdmSuGL9_0),.din(w_dff_A_J4dk22Yl9_0),.clk(gclk));
	jdff dff_A_4CdmSuGL9_0(.dout(w_dff_A_nHWK10bh2_0),.din(w_dff_A_4CdmSuGL9_0),.clk(gclk));
	jdff dff_A_nHWK10bh2_0(.dout(w_dff_A_8VRwnKMI3_0),.din(w_dff_A_nHWK10bh2_0),.clk(gclk));
	jdff dff_A_8VRwnKMI3_0(.dout(w_dff_A_MQl52QAR1_0),.din(w_dff_A_8VRwnKMI3_0),.clk(gclk));
	jdff dff_A_MQl52QAR1_0(.dout(G3552gat),.din(w_dff_A_MQl52QAR1_0),.clk(gclk));
	jdff dff_A_nMXYqaCW1_2(.dout(w_dff_A_YYpgINDy3_0),.din(w_dff_A_nMXYqaCW1_2),.clk(gclk));
	jdff dff_A_YYpgINDy3_0(.dout(w_dff_A_lwrrrB3p7_0),.din(w_dff_A_YYpgINDy3_0),.clk(gclk));
	jdff dff_A_lwrrrB3p7_0(.dout(w_dff_A_B8fJ0ntx2_0),.din(w_dff_A_lwrrrB3p7_0),.clk(gclk));
	jdff dff_A_B8fJ0ntx2_0(.dout(w_dff_A_YjvteGTd2_0),.din(w_dff_A_B8fJ0ntx2_0),.clk(gclk));
	jdff dff_A_YjvteGTd2_0(.dout(w_dff_A_yaTgu2VO1_0),.din(w_dff_A_YjvteGTd2_0),.clk(gclk));
	jdff dff_A_yaTgu2VO1_0(.dout(w_dff_A_SEcWP5OR6_0),.din(w_dff_A_yaTgu2VO1_0),.clk(gclk));
	jdff dff_A_SEcWP5OR6_0(.dout(w_dff_A_D1OXEpw21_0),.din(w_dff_A_SEcWP5OR6_0),.clk(gclk));
	jdff dff_A_D1OXEpw21_0(.dout(w_dff_A_v8GX5eHi7_0),.din(w_dff_A_D1OXEpw21_0),.clk(gclk));
	jdff dff_A_v8GX5eHi7_0(.dout(w_dff_A_ZUHgF6Eb5_0),.din(w_dff_A_v8GX5eHi7_0),.clk(gclk));
	jdff dff_A_ZUHgF6Eb5_0(.dout(w_dff_A_u6QIqdzu5_0),.din(w_dff_A_ZUHgF6Eb5_0),.clk(gclk));
	jdff dff_A_u6QIqdzu5_0(.dout(w_dff_A_o5NFb3Ii8_0),.din(w_dff_A_u6QIqdzu5_0),.clk(gclk));
	jdff dff_A_o5NFb3Ii8_0(.dout(w_dff_A_35zqimbM6_0),.din(w_dff_A_o5NFb3Ii8_0),.clk(gclk));
	jdff dff_A_35zqimbM6_0(.dout(w_dff_A_kusZDYTx2_0),.din(w_dff_A_35zqimbM6_0),.clk(gclk));
	jdff dff_A_kusZDYTx2_0(.dout(w_dff_A_cgnjCkye7_0),.din(w_dff_A_kusZDYTx2_0),.clk(gclk));
	jdff dff_A_cgnjCkye7_0(.dout(w_dff_A_Y0bRhwzn5_0),.din(w_dff_A_cgnjCkye7_0),.clk(gclk));
	jdff dff_A_Y0bRhwzn5_0(.dout(w_dff_A_JdIDhnLx5_0),.din(w_dff_A_Y0bRhwzn5_0),.clk(gclk));
	jdff dff_A_JdIDhnLx5_0(.dout(w_dff_A_jsWGIM580_0),.din(w_dff_A_JdIDhnLx5_0),.clk(gclk));
	jdff dff_A_jsWGIM580_0(.dout(w_dff_A_Z9J2BnBh3_0),.din(w_dff_A_jsWGIM580_0),.clk(gclk));
	jdff dff_A_Z9J2BnBh3_0(.dout(w_dff_A_izzOODcx7_0),.din(w_dff_A_Z9J2BnBh3_0),.clk(gclk));
	jdff dff_A_izzOODcx7_0(.dout(w_dff_A_vyoYzxX94_0),.din(w_dff_A_izzOODcx7_0),.clk(gclk));
	jdff dff_A_vyoYzxX94_0(.dout(w_dff_A_r4KHrzwQ1_0),.din(w_dff_A_vyoYzxX94_0),.clk(gclk));
	jdff dff_A_r4KHrzwQ1_0(.dout(w_dff_A_JrmBbtdJ8_0),.din(w_dff_A_r4KHrzwQ1_0),.clk(gclk));
	jdff dff_A_JrmBbtdJ8_0(.dout(w_dff_A_M6jBHEeD8_0),.din(w_dff_A_JrmBbtdJ8_0),.clk(gclk));
	jdff dff_A_M6jBHEeD8_0(.dout(w_dff_A_y10g4YGS6_0),.din(w_dff_A_M6jBHEeD8_0),.clk(gclk));
	jdff dff_A_y10g4YGS6_0(.dout(w_dff_A_nHcE0DUg9_0),.din(w_dff_A_y10g4YGS6_0),.clk(gclk));
	jdff dff_A_nHcE0DUg9_0(.dout(w_dff_A_0BhYfPlQ7_0),.din(w_dff_A_nHcE0DUg9_0),.clk(gclk));
	jdff dff_A_0BhYfPlQ7_0(.dout(w_dff_A_ywoydGKi4_0),.din(w_dff_A_0BhYfPlQ7_0),.clk(gclk));
	jdff dff_A_ywoydGKi4_0(.dout(w_dff_A_FeWTgB8k8_0),.din(w_dff_A_ywoydGKi4_0),.clk(gclk));
	jdff dff_A_FeWTgB8k8_0(.dout(w_dff_A_yNnk6Uvw5_0),.din(w_dff_A_FeWTgB8k8_0),.clk(gclk));
	jdff dff_A_yNnk6Uvw5_0(.dout(w_dff_A_9QLcHwXy2_0),.din(w_dff_A_yNnk6Uvw5_0),.clk(gclk));
	jdff dff_A_9QLcHwXy2_0(.dout(w_dff_A_96No0DOe8_0),.din(w_dff_A_9QLcHwXy2_0),.clk(gclk));
	jdff dff_A_96No0DOe8_0(.dout(w_dff_A_TbQglCN53_0),.din(w_dff_A_96No0DOe8_0),.clk(gclk));
	jdff dff_A_TbQglCN53_0(.dout(w_dff_A_pI0ROOVO7_0),.din(w_dff_A_TbQglCN53_0),.clk(gclk));
	jdff dff_A_pI0ROOVO7_0(.dout(w_dff_A_19zbZyDP2_0),.din(w_dff_A_pI0ROOVO7_0),.clk(gclk));
	jdff dff_A_19zbZyDP2_0(.dout(w_dff_A_wtQSMymi6_0),.din(w_dff_A_19zbZyDP2_0),.clk(gclk));
	jdff dff_A_wtQSMymi6_0(.dout(w_dff_A_pNM5oZap1_0),.din(w_dff_A_wtQSMymi6_0),.clk(gclk));
	jdff dff_A_pNM5oZap1_0(.dout(w_dff_A_OZvvVaKl1_0),.din(w_dff_A_pNM5oZap1_0),.clk(gclk));
	jdff dff_A_OZvvVaKl1_0(.dout(w_dff_A_PzCWopPt7_0),.din(w_dff_A_OZvvVaKl1_0),.clk(gclk));
	jdff dff_A_PzCWopPt7_0(.dout(w_dff_A_9S4vkzzc3_0),.din(w_dff_A_PzCWopPt7_0),.clk(gclk));
	jdff dff_A_9S4vkzzc3_0(.dout(w_dff_A_Qi5Sacb09_0),.din(w_dff_A_9S4vkzzc3_0),.clk(gclk));
	jdff dff_A_Qi5Sacb09_0(.dout(w_dff_A_LLzdCRSK6_0),.din(w_dff_A_Qi5Sacb09_0),.clk(gclk));
	jdff dff_A_LLzdCRSK6_0(.dout(w_dff_A_8C7GdqWL1_0),.din(w_dff_A_LLzdCRSK6_0),.clk(gclk));
	jdff dff_A_8C7GdqWL1_0(.dout(w_dff_A_fcA96LoP8_0),.din(w_dff_A_8C7GdqWL1_0),.clk(gclk));
	jdff dff_A_fcA96LoP8_0(.dout(w_dff_A_dTCWqSlQ2_0),.din(w_dff_A_fcA96LoP8_0),.clk(gclk));
	jdff dff_A_dTCWqSlQ2_0(.dout(w_dff_A_R0aARRQc7_0),.din(w_dff_A_dTCWqSlQ2_0),.clk(gclk));
	jdff dff_A_R0aARRQc7_0(.dout(w_dff_A_5Mm8Y8dt2_0),.din(w_dff_A_R0aARRQc7_0),.clk(gclk));
	jdff dff_A_5Mm8Y8dt2_0(.dout(w_dff_A_Idj8UVp15_0),.din(w_dff_A_5Mm8Y8dt2_0),.clk(gclk));
	jdff dff_A_Idj8UVp15_0(.dout(w_dff_A_Rdzpgkfa3_0),.din(w_dff_A_Idj8UVp15_0),.clk(gclk));
	jdff dff_A_Rdzpgkfa3_0(.dout(w_dff_A_ykGrHtUK1_0),.din(w_dff_A_Rdzpgkfa3_0),.clk(gclk));
	jdff dff_A_ykGrHtUK1_0(.dout(w_dff_A_Er4tz4if6_0),.din(w_dff_A_ykGrHtUK1_0),.clk(gclk));
	jdff dff_A_Er4tz4if6_0(.dout(G3895gat),.din(w_dff_A_Er4tz4if6_0),.clk(gclk));
	jdff dff_A_jS7LkhAz1_2(.dout(w_dff_A_rYdq5y3o6_0),.din(w_dff_A_jS7LkhAz1_2),.clk(gclk));
	jdff dff_A_rYdq5y3o6_0(.dout(w_dff_A_aNacdnhV0_0),.din(w_dff_A_rYdq5y3o6_0),.clk(gclk));
	jdff dff_A_aNacdnhV0_0(.dout(w_dff_A_YpzLEucd6_0),.din(w_dff_A_aNacdnhV0_0),.clk(gclk));
	jdff dff_A_YpzLEucd6_0(.dout(w_dff_A_hGThfReO3_0),.din(w_dff_A_YpzLEucd6_0),.clk(gclk));
	jdff dff_A_hGThfReO3_0(.dout(w_dff_A_qRNHv9At6_0),.din(w_dff_A_hGThfReO3_0),.clk(gclk));
	jdff dff_A_qRNHv9At6_0(.dout(w_dff_A_11EZkWzy2_0),.din(w_dff_A_qRNHv9At6_0),.clk(gclk));
	jdff dff_A_11EZkWzy2_0(.dout(w_dff_A_95CyLDFD7_0),.din(w_dff_A_11EZkWzy2_0),.clk(gclk));
	jdff dff_A_95CyLDFD7_0(.dout(w_dff_A_L1mesjpJ0_0),.din(w_dff_A_95CyLDFD7_0),.clk(gclk));
	jdff dff_A_L1mesjpJ0_0(.dout(w_dff_A_YbnuNaDi3_0),.din(w_dff_A_L1mesjpJ0_0),.clk(gclk));
	jdff dff_A_YbnuNaDi3_0(.dout(w_dff_A_D9Wqwrpl1_0),.din(w_dff_A_YbnuNaDi3_0),.clk(gclk));
	jdff dff_A_D9Wqwrpl1_0(.dout(w_dff_A_Dmrc0wNa9_0),.din(w_dff_A_D9Wqwrpl1_0),.clk(gclk));
	jdff dff_A_Dmrc0wNa9_0(.dout(w_dff_A_9Vst5bMJ3_0),.din(w_dff_A_Dmrc0wNa9_0),.clk(gclk));
	jdff dff_A_9Vst5bMJ3_0(.dout(w_dff_A_btsBmhzI6_0),.din(w_dff_A_9Vst5bMJ3_0),.clk(gclk));
	jdff dff_A_btsBmhzI6_0(.dout(w_dff_A_P8hvuDZx6_0),.din(w_dff_A_btsBmhzI6_0),.clk(gclk));
	jdff dff_A_P8hvuDZx6_0(.dout(w_dff_A_fpSGDsJV3_0),.din(w_dff_A_P8hvuDZx6_0),.clk(gclk));
	jdff dff_A_fpSGDsJV3_0(.dout(w_dff_A_JPcHcMZo9_0),.din(w_dff_A_fpSGDsJV3_0),.clk(gclk));
	jdff dff_A_JPcHcMZo9_0(.dout(w_dff_A_AHEyVeYx6_0),.din(w_dff_A_JPcHcMZo9_0),.clk(gclk));
	jdff dff_A_AHEyVeYx6_0(.dout(w_dff_A_CaUtmfT38_0),.din(w_dff_A_AHEyVeYx6_0),.clk(gclk));
	jdff dff_A_CaUtmfT38_0(.dout(w_dff_A_OTz6aHL36_0),.din(w_dff_A_CaUtmfT38_0),.clk(gclk));
	jdff dff_A_OTz6aHL36_0(.dout(w_dff_A_7E1PTGuK9_0),.din(w_dff_A_OTz6aHL36_0),.clk(gclk));
	jdff dff_A_7E1PTGuK9_0(.dout(w_dff_A_JxfX8zAx4_0),.din(w_dff_A_7E1PTGuK9_0),.clk(gclk));
	jdff dff_A_JxfX8zAx4_0(.dout(w_dff_A_4ogO21bK2_0),.din(w_dff_A_JxfX8zAx4_0),.clk(gclk));
	jdff dff_A_4ogO21bK2_0(.dout(w_dff_A_mrEdarCm7_0),.din(w_dff_A_4ogO21bK2_0),.clk(gclk));
	jdff dff_A_mrEdarCm7_0(.dout(w_dff_A_e1XVe4sA1_0),.din(w_dff_A_mrEdarCm7_0),.clk(gclk));
	jdff dff_A_e1XVe4sA1_0(.dout(w_dff_A_tH9kGI2s0_0),.din(w_dff_A_e1XVe4sA1_0),.clk(gclk));
	jdff dff_A_tH9kGI2s0_0(.dout(w_dff_A_L5zbAgZ49_0),.din(w_dff_A_tH9kGI2s0_0),.clk(gclk));
	jdff dff_A_L5zbAgZ49_0(.dout(w_dff_A_UbOOOFqZ1_0),.din(w_dff_A_L5zbAgZ49_0),.clk(gclk));
	jdff dff_A_UbOOOFqZ1_0(.dout(w_dff_A_FKG7jUTr7_0),.din(w_dff_A_UbOOOFqZ1_0),.clk(gclk));
	jdff dff_A_FKG7jUTr7_0(.dout(w_dff_A_fhSc2Xbt9_0),.din(w_dff_A_FKG7jUTr7_0),.clk(gclk));
	jdff dff_A_fhSc2Xbt9_0(.dout(w_dff_A_bYyJYapF5_0),.din(w_dff_A_fhSc2Xbt9_0),.clk(gclk));
	jdff dff_A_bYyJYapF5_0(.dout(w_dff_A_bMoVnqGV3_0),.din(w_dff_A_bYyJYapF5_0),.clk(gclk));
	jdff dff_A_bMoVnqGV3_0(.dout(w_dff_A_3fh4P4QS4_0),.din(w_dff_A_bMoVnqGV3_0),.clk(gclk));
	jdff dff_A_3fh4P4QS4_0(.dout(w_dff_A_aWvbuDCF3_0),.din(w_dff_A_3fh4P4QS4_0),.clk(gclk));
	jdff dff_A_aWvbuDCF3_0(.dout(w_dff_A_PFEd0Xos4_0),.din(w_dff_A_aWvbuDCF3_0),.clk(gclk));
	jdff dff_A_PFEd0Xos4_0(.dout(w_dff_A_e6iNcabG9_0),.din(w_dff_A_PFEd0Xos4_0),.clk(gclk));
	jdff dff_A_e6iNcabG9_0(.dout(w_dff_A_eUgayTAz1_0),.din(w_dff_A_e6iNcabG9_0),.clk(gclk));
	jdff dff_A_eUgayTAz1_0(.dout(w_dff_A_FHm4QNY21_0),.din(w_dff_A_eUgayTAz1_0),.clk(gclk));
	jdff dff_A_FHm4QNY21_0(.dout(w_dff_A_0q13euX98_0),.din(w_dff_A_FHm4QNY21_0),.clk(gclk));
	jdff dff_A_0q13euX98_0(.dout(w_dff_A_IR2pIF1V0_0),.din(w_dff_A_0q13euX98_0),.clk(gclk));
	jdff dff_A_IR2pIF1V0_0(.dout(w_dff_A_BPW7a3Os3_0),.din(w_dff_A_IR2pIF1V0_0),.clk(gclk));
	jdff dff_A_BPW7a3Os3_0(.dout(w_dff_A_dyBO7idN3_0),.din(w_dff_A_BPW7a3Os3_0),.clk(gclk));
	jdff dff_A_dyBO7idN3_0(.dout(w_dff_A_fHtNZdYZ2_0),.din(w_dff_A_dyBO7idN3_0),.clk(gclk));
	jdff dff_A_fHtNZdYZ2_0(.dout(w_dff_A_x2JstJLm6_0),.din(w_dff_A_fHtNZdYZ2_0),.clk(gclk));
	jdff dff_A_x2JstJLm6_0(.dout(w_dff_A_KfmLhOCS4_0),.din(w_dff_A_x2JstJLm6_0),.clk(gclk));
	jdff dff_A_KfmLhOCS4_0(.dout(w_dff_A_RqhStVCN8_0),.din(w_dff_A_KfmLhOCS4_0),.clk(gclk));
	jdff dff_A_RqhStVCN8_0(.dout(w_dff_A_rfkhjkw56_0),.din(w_dff_A_RqhStVCN8_0),.clk(gclk));
	jdff dff_A_rfkhjkw56_0(.dout(w_dff_A_TsEFZypi0_0),.din(w_dff_A_rfkhjkw56_0),.clk(gclk));
	jdff dff_A_TsEFZypi0_0(.dout(G4241gat),.din(w_dff_A_TsEFZypi0_0),.clk(gclk));
	jdff dff_A_jXnwwKqc6_2(.dout(w_dff_A_EyhkW8kI9_0),.din(w_dff_A_jXnwwKqc6_2),.clk(gclk));
	jdff dff_A_EyhkW8kI9_0(.dout(w_dff_A_HHYTkiHh7_0),.din(w_dff_A_EyhkW8kI9_0),.clk(gclk));
	jdff dff_A_HHYTkiHh7_0(.dout(w_dff_A_pr4g7m6B6_0),.din(w_dff_A_HHYTkiHh7_0),.clk(gclk));
	jdff dff_A_pr4g7m6B6_0(.dout(w_dff_A_2sMFBNzG1_0),.din(w_dff_A_pr4g7m6B6_0),.clk(gclk));
	jdff dff_A_2sMFBNzG1_0(.dout(w_dff_A_YFyweRcv5_0),.din(w_dff_A_2sMFBNzG1_0),.clk(gclk));
	jdff dff_A_YFyweRcv5_0(.dout(w_dff_A_3KCa8cg62_0),.din(w_dff_A_YFyweRcv5_0),.clk(gclk));
	jdff dff_A_3KCa8cg62_0(.dout(w_dff_A_dBclAjSs5_0),.din(w_dff_A_3KCa8cg62_0),.clk(gclk));
	jdff dff_A_dBclAjSs5_0(.dout(w_dff_A_OGYqzOkd6_0),.din(w_dff_A_dBclAjSs5_0),.clk(gclk));
	jdff dff_A_OGYqzOkd6_0(.dout(w_dff_A_DlFXrXBO9_0),.din(w_dff_A_OGYqzOkd6_0),.clk(gclk));
	jdff dff_A_DlFXrXBO9_0(.dout(w_dff_A_lz2DAHkv1_0),.din(w_dff_A_DlFXrXBO9_0),.clk(gclk));
	jdff dff_A_lz2DAHkv1_0(.dout(w_dff_A_foRu15oU4_0),.din(w_dff_A_lz2DAHkv1_0),.clk(gclk));
	jdff dff_A_foRu15oU4_0(.dout(w_dff_A_N6AyBItT9_0),.din(w_dff_A_foRu15oU4_0),.clk(gclk));
	jdff dff_A_N6AyBItT9_0(.dout(w_dff_A_jDlaZ5oN0_0),.din(w_dff_A_N6AyBItT9_0),.clk(gclk));
	jdff dff_A_jDlaZ5oN0_0(.dout(w_dff_A_4k5Arbv01_0),.din(w_dff_A_jDlaZ5oN0_0),.clk(gclk));
	jdff dff_A_4k5Arbv01_0(.dout(w_dff_A_wrJKIFmZ3_0),.din(w_dff_A_4k5Arbv01_0),.clk(gclk));
	jdff dff_A_wrJKIFmZ3_0(.dout(w_dff_A_eOHTfR564_0),.din(w_dff_A_wrJKIFmZ3_0),.clk(gclk));
	jdff dff_A_eOHTfR564_0(.dout(w_dff_A_dpkBOj0d6_0),.din(w_dff_A_eOHTfR564_0),.clk(gclk));
	jdff dff_A_dpkBOj0d6_0(.dout(w_dff_A_zeFohYIq0_0),.din(w_dff_A_dpkBOj0d6_0),.clk(gclk));
	jdff dff_A_zeFohYIq0_0(.dout(w_dff_A_m1RaIO4f8_0),.din(w_dff_A_zeFohYIq0_0),.clk(gclk));
	jdff dff_A_m1RaIO4f8_0(.dout(w_dff_A_4sTr0x073_0),.din(w_dff_A_m1RaIO4f8_0),.clk(gclk));
	jdff dff_A_4sTr0x073_0(.dout(w_dff_A_lhDRANhY5_0),.din(w_dff_A_4sTr0x073_0),.clk(gclk));
	jdff dff_A_lhDRANhY5_0(.dout(w_dff_A_U97lU8Df2_0),.din(w_dff_A_lhDRANhY5_0),.clk(gclk));
	jdff dff_A_U97lU8Df2_0(.dout(w_dff_A_cTpNyUj90_0),.din(w_dff_A_U97lU8Df2_0),.clk(gclk));
	jdff dff_A_cTpNyUj90_0(.dout(w_dff_A_85YsmSJS4_0),.din(w_dff_A_cTpNyUj90_0),.clk(gclk));
	jdff dff_A_85YsmSJS4_0(.dout(w_dff_A_Wi2L1H9b2_0),.din(w_dff_A_85YsmSJS4_0),.clk(gclk));
	jdff dff_A_Wi2L1H9b2_0(.dout(w_dff_A_32JurMhH5_0),.din(w_dff_A_Wi2L1H9b2_0),.clk(gclk));
	jdff dff_A_32JurMhH5_0(.dout(w_dff_A_q6kNwUVp2_0),.din(w_dff_A_32JurMhH5_0),.clk(gclk));
	jdff dff_A_q6kNwUVp2_0(.dout(w_dff_A_VKwdWK2t8_0),.din(w_dff_A_q6kNwUVp2_0),.clk(gclk));
	jdff dff_A_VKwdWK2t8_0(.dout(w_dff_A_YCY0nPRx8_0),.din(w_dff_A_VKwdWK2t8_0),.clk(gclk));
	jdff dff_A_YCY0nPRx8_0(.dout(w_dff_A_DeD0Xxjt4_0),.din(w_dff_A_YCY0nPRx8_0),.clk(gclk));
	jdff dff_A_DeD0Xxjt4_0(.dout(w_dff_A_aTOxYAW03_0),.din(w_dff_A_DeD0Xxjt4_0),.clk(gclk));
	jdff dff_A_aTOxYAW03_0(.dout(w_dff_A_5iGNlgD84_0),.din(w_dff_A_aTOxYAW03_0),.clk(gclk));
	jdff dff_A_5iGNlgD84_0(.dout(w_dff_A_LOCMHPqz1_0),.din(w_dff_A_5iGNlgD84_0),.clk(gclk));
	jdff dff_A_LOCMHPqz1_0(.dout(w_dff_A_fuEUCixC4_0),.din(w_dff_A_LOCMHPqz1_0),.clk(gclk));
	jdff dff_A_fuEUCixC4_0(.dout(w_dff_A_YcGhvpYK5_0),.din(w_dff_A_fuEUCixC4_0),.clk(gclk));
	jdff dff_A_YcGhvpYK5_0(.dout(w_dff_A_Kq8QgNPy8_0),.din(w_dff_A_YcGhvpYK5_0),.clk(gclk));
	jdff dff_A_Kq8QgNPy8_0(.dout(w_dff_A_IDge9Oud0_0),.din(w_dff_A_Kq8QgNPy8_0),.clk(gclk));
	jdff dff_A_IDge9Oud0_0(.dout(w_dff_A_NafXWdyD9_0),.din(w_dff_A_IDge9Oud0_0),.clk(gclk));
	jdff dff_A_NafXWdyD9_0(.dout(w_dff_A_moFZvKrK4_0),.din(w_dff_A_NafXWdyD9_0),.clk(gclk));
	jdff dff_A_moFZvKrK4_0(.dout(w_dff_A_jlJU8G6u5_0),.din(w_dff_A_moFZvKrK4_0),.clk(gclk));
	jdff dff_A_jlJU8G6u5_0(.dout(w_dff_A_XEIVmxyX6_0),.din(w_dff_A_jlJU8G6u5_0),.clk(gclk));
	jdff dff_A_XEIVmxyX6_0(.dout(w_dff_A_J2NaBzCs1_0),.din(w_dff_A_XEIVmxyX6_0),.clk(gclk));
	jdff dff_A_J2NaBzCs1_0(.dout(w_dff_A_eYorYIE99_0),.din(w_dff_A_J2NaBzCs1_0),.clk(gclk));
	jdff dff_A_eYorYIE99_0(.dout(w_dff_A_0P7PXjZ73_0),.din(w_dff_A_eYorYIE99_0),.clk(gclk));
	jdff dff_A_0P7PXjZ73_0(.dout(G4591gat),.din(w_dff_A_0P7PXjZ73_0),.clk(gclk));
	jdff dff_A_InJoAco86_2(.dout(w_dff_A_8tFjG5Nu4_0),.din(w_dff_A_InJoAco86_2),.clk(gclk));
	jdff dff_A_8tFjG5Nu4_0(.dout(w_dff_A_adZFhVWt3_0),.din(w_dff_A_8tFjG5Nu4_0),.clk(gclk));
	jdff dff_A_adZFhVWt3_0(.dout(w_dff_A_khQeFtbi2_0),.din(w_dff_A_adZFhVWt3_0),.clk(gclk));
	jdff dff_A_khQeFtbi2_0(.dout(w_dff_A_pawRfK1G2_0),.din(w_dff_A_khQeFtbi2_0),.clk(gclk));
	jdff dff_A_pawRfK1G2_0(.dout(w_dff_A_lHQnDnJv7_0),.din(w_dff_A_pawRfK1G2_0),.clk(gclk));
	jdff dff_A_lHQnDnJv7_0(.dout(w_dff_A_kiy4hM7B1_0),.din(w_dff_A_lHQnDnJv7_0),.clk(gclk));
	jdff dff_A_kiy4hM7B1_0(.dout(w_dff_A_WZQwmKDJ9_0),.din(w_dff_A_kiy4hM7B1_0),.clk(gclk));
	jdff dff_A_WZQwmKDJ9_0(.dout(w_dff_A_oeFFh1Qd8_0),.din(w_dff_A_WZQwmKDJ9_0),.clk(gclk));
	jdff dff_A_oeFFh1Qd8_0(.dout(w_dff_A_KNo4ep9N4_0),.din(w_dff_A_oeFFh1Qd8_0),.clk(gclk));
	jdff dff_A_KNo4ep9N4_0(.dout(w_dff_A_LFG5QP5K3_0),.din(w_dff_A_KNo4ep9N4_0),.clk(gclk));
	jdff dff_A_LFG5QP5K3_0(.dout(w_dff_A_4wOkTt5C8_0),.din(w_dff_A_LFG5QP5K3_0),.clk(gclk));
	jdff dff_A_4wOkTt5C8_0(.dout(w_dff_A_7VtlChLr7_0),.din(w_dff_A_4wOkTt5C8_0),.clk(gclk));
	jdff dff_A_7VtlChLr7_0(.dout(w_dff_A_VteV8FS84_0),.din(w_dff_A_7VtlChLr7_0),.clk(gclk));
	jdff dff_A_VteV8FS84_0(.dout(w_dff_A_tlx0rhtQ9_0),.din(w_dff_A_VteV8FS84_0),.clk(gclk));
	jdff dff_A_tlx0rhtQ9_0(.dout(w_dff_A_92ta0ssu8_0),.din(w_dff_A_tlx0rhtQ9_0),.clk(gclk));
	jdff dff_A_92ta0ssu8_0(.dout(w_dff_A_AEKKLIYV7_0),.din(w_dff_A_92ta0ssu8_0),.clk(gclk));
	jdff dff_A_AEKKLIYV7_0(.dout(w_dff_A_0ixeKnDn9_0),.din(w_dff_A_AEKKLIYV7_0),.clk(gclk));
	jdff dff_A_0ixeKnDn9_0(.dout(w_dff_A_PqXnSlV98_0),.din(w_dff_A_0ixeKnDn9_0),.clk(gclk));
	jdff dff_A_PqXnSlV98_0(.dout(w_dff_A_lgn9l7ch1_0),.din(w_dff_A_PqXnSlV98_0),.clk(gclk));
	jdff dff_A_lgn9l7ch1_0(.dout(w_dff_A_KpNFLpMX4_0),.din(w_dff_A_lgn9l7ch1_0),.clk(gclk));
	jdff dff_A_KpNFLpMX4_0(.dout(w_dff_A_aWKhFH2m5_0),.din(w_dff_A_KpNFLpMX4_0),.clk(gclk));
	jdff dff_A_aWKhFH2m5_0(.dout(w_dff_A_VZdekvL53_0),.din(w_dff_A_aWKhFH2m5_0),.clk(gclk));
	jdff dff_A_VZdekvL53_0(.dout(w_dff_A_tAEldFgU2_0),.din(w_dff_A_VZdekvL53_0),.clk(gclk));
	jdff dff_A_tAEldFgU2_0(.dout(w_dff_A_GUwmpE9s6_0),.din(w_dff_A_tAEldFgU2_0),.clk(gclk));
	jdff dff_A_GUwmpE9s6_0(.dout(w_dff_A_AdUBg0mg6_0),.din(w_dff_A_GUwmpE9s6_0),.clk(gclk));
	jdff dff_A_AdUBg0mg6_0(.dout(w_dff_A_rP6G0iiV7_0),.din(w_dff_A_AdUBg0mg6_0),.clk(gclk));
	jdff dff_A_rP6G0iiV7_0(.dout(w_dff_A_kRm8IWAG9_0),.din(w_dff_A_rP6G0iiV7_0),.clk(gclk));
	jdff dff_A_kRm8IWAG9_0(.dout(w_dff_A_zknHFImh4_0),.din(w_dff_A_kRm8IWAG9_0),.clk(gclk));
	jdff dff_A_zknHFImh4_0(.dout(w_dff_A_bjuChTcd4_0),.din(w_dff_A_zknHFImh4_0),.clk(gclk));
	jdff dff_A_bjuChTcd4_0(.dout(w_dff_A_Py5PRoml6_0),.din(w_dff_A_bjuChTcd4_0),.clk(gclk));
	jdff dff_A_Py5PRoml6_0(.dout(w_dff_A_XYMOkY597_0),.din(w_dff_A_Py5PRoml6_0),.clk(gclk));
	jdff dff_A_XYMOkY597_0(.dout(w_dff_A_pgIJinxr2_0),.din(w_dff_A_XYMOkY597_0),.clk(gclk));
	jdff dff_A_pgIJinxr2_0(.dout(w_dff_A_gR9x8sir8_0),.din(w_dff_A_pgIJinxr2_0),.clk(gclk));
	jdff dff_A_gR9x8sir8_0(.dout(w_dff_A_mTznjd3V1_0),.din(w_dff_A_gR9x8sir8_0),.clk(gclk));
	jdff dff_A_mTznjd3V1_0(.dout(w_dff_A_po6byZm51_0),.din(w_dff_A_mTznjd3V1_0),.clk(gclk));
	jdff dff_A_po6byZm51_0(.dout(w_dff_A_NkEXzxnV6_0),.din(w_dff_A_po6byZm51_0),.clk(gclk));
	jdff dff_A_NkEXzxnV6_0(.dout(w_dff_A_bRrItFUZ7_0),.din(w_dff_A_NkEXzxnV6_0),.clk(gclk));
	jdff dff_A_bRrItFUZ7_0(.dout(w_dff_A_Z4r2umF19_0),.din(w_dff_A_bRrItFUZ7_0),.clk(gclk));
	jdff dff_A_Z4r2umF19_0(.dout(w_dff_A_w9Y5PU9q1_0),.din(w_dff_A_Z4r2umF19_0),.clk(gclk));
	jdff dff_A_w9Y5PU9q1_0(.dout(w_dff_A_53xL7dgN4_0),.din(w_dff_A_w9Y5PU9q1_0),.clk(gclk));
	jdff dff_A_53xL7dgN4_0(.dout(w_dff_A_mocf161Y5_0),.din(w_dff_A_53xL7dgN4_0),.clk(gclk));
	jdff dff_A_mocf161Y5_0(.dout(G4946gat),.din(w_dff_A_mocf161Y5_0),.clk(gclk));
	jdff dff_A_XOoOUeVN7_2(.dout(w_dff_A_2XzYw5Sx7_0),.din(w_dff_A_XOoOUeVN7_2),.clk(gclk));
	jdff dff_A_2XzYw5Sx7_0(.dout(w_dff_A_54or12fq0_0),.din(w_dff_A_2XzYw5Sx7_0),.clk(gclk));
	jdff dff_A_54or12fq0_0(.dout(w_dff_A_OWIeZrdq8_0),.din(w_dff_A_54or12fq0_0),.clk(gclk));
	jdff dff_A_OWIeZrdq8_0(.dout(w_dff_A_3RK770oa1_0),.din(w_dff_A_OWIeZrdq8_0),.clk(gclk));
	jdff dff_A_3RK770oa1_0(.dout(w_dff_A_vMMXiNqg9_0),.din(w_dff_A_3RK770oa1_0),.clk(gclk));
	jdff dff_A_vMMXiNqg9_0(.dout(w_dff_A_ELqyL6p15_0),.din(w_dff_A_vMMXiNqg9_0),.clk(gclk));
	jdff dff_A_ELqyL6p15_0(.dout(w_dff_A_ubsyBGdE0_0),.din(w_dff_A_ELqyL6p15_0),.clk(gclk));
	jdff dff_A_ubsyBGdE0_0(.dout(w_dff_A_pHQzrwBN7_0),.din(w_dff_A_ubsyBGdE0_0),.clk(gclk));
	jdff dff_A_pHQzrwBN7_0(.dout(w_dff_A_X9yQ8z6n0_0),.din(w_dff_A_pHQzrwBN7_0),.clk(gclk));
	jdff dff_A_X9yQ8z6n0_0(.dout(w_dff_A_xTgPQv3V5_0),.din(w_dff_A_X9yQ8z6n0_0),.clk(gclk));
	jdff dff_A_xTgPQv3V5_0(.dout(w_dff_A_37HwXmjE4_0),.din(w_dff_A_xTgPQv3V5_0),.clk(gclk));
	jdff dff_A_37HwXmjE4_0(.dout(w_dff_A_aNyO50tc7_0),.din(w_dff_A_37HwXmjE4_0),.clk(gclk));
	jdff dff_A_aNyO50tc7_0(.dout(w_dff_A_dRVfjY9J9_0),.din(w_dff_A_aNyO50tc7_0),.clk(gclk));
	jdff dff_A_dRVfjY9J9_0(.dout(w_dff_A_OURD4cKj9_0),.din(w_dff_A_dRVfjY9J9_0),.clk(gclk));
	jdff dff_A_OURD4cKj9_0(.dout(w_dff_A_tD30K2Zm8_0),.din(w_dff_A_OURD4cKj9_0),.clk(gclk));
	jdff dff_A_tD30K2Zm8_0(.dout(w_dff_A_86Ws02WH4_0),.din(w_dff_A_tD30K2Zm8_0),.clk(gclk));
	jdff dff_A_86Ws02WH4_0(.dout(w_dff_A_BWIjOuxE1_0),.din(w_dff_A_86Ws02WH4_0),.clk(gclk));
	jdff dff_A_BWIjOuxE1_0(.dout(w_dff_A_GJAHJOxT4_0),.din(w_dff_A_BWIjOuxE1_0),.clk(gclk));
	jdff dff_A_GJAHJOxT4_0(.dout(w_dff_A_dyiAxvMi1_0),.din(w_dff_A_GJAHJOxT4_0),.clk(gclk));
	jdff dff_A_dyiAxvMi1_0(.dout(w_dff_A_cXVsAY8B3_0),.din(w_dff_A_dyiAxvMi1_0),.clk(gclk));
	jdff dff_A_cXVsAY8B3_0(.dout(w_dff_A_m1o9RK7j9_0),.din(w_dff_A_cXVsAY8B3_0),.clk(gclk));
	jdff dff_A_m1o9RK7j9_0(.dout(w_dff_A_G0pxffjw2_0),.din(w_dff_A_m1o9RK7j9_0),.clk(gclk));
	jdff dff_A_G0pxffjw2_0(.dout(w_dff_A_vnjbYvWV6_0),.din(w_dff_A_G0pxffjw2_0),.clk(gclk));
	jdff dff_A_vnjbYvWV6_0(.dout(w_dff_A_MSSxBnnR7_0),.din(w_dff_A_vnjbYvWV6_0),.clk(gclk));
	jdff dff_A_MSSxBnnR7_0(.dout(w_dff_A_u6Pp6xdQ7_0),.din(w_dff_A_MSSxBnnR7_0),.clk(gclk));
	jdff dff_A_u6Pp6xdQ7_0(.dout(w_dff_A_jFP94YyL3_0),.din(w_dff_A_u6Pp6xdQ7_0),.clk(gclk));
	jdff dff_A_jFP94YyL3_0(.dout(w_dff_A_IrK5KcnO6_0),.din(w_dff_A_jFP94YyL3_0),.clk(gclk));
	jdff dff_A_IrK5KcnO6_0(.dout(w_dff_A_0URgGxv48_0),.din(w_dff_A_IrK5KcnO6_0),.clk(gclk));
	jdff dff_A_0URgGxv48_0(.dout(w_dff_A_WCz3bCSs5_0),.din(w_dff_A_0URgGxv48_0),.clk(gclk));
	jdff dff_A_WCz3bCSs5_0(.dout(w_dff_A_Is2VsdUM2_0),.din(w_dff_A_WCz3bCSs5_0),.clk(gclk));
	jdff dff_A_Is2VsdUM2_0(.dout(w_dff_A_K1iWiehT4_0),.din(w_dff_A_Is2VsdUM2_0),.clk(gclk));
	jdff dff_A_K1iWiehT4_0(.dout(w_dff_A_zA4Jzm3R2_0),.din(w_dff_A_K1iWiehT4_0),.clk(gclk));
	jdff dff_A_zA4Jzm3R2_0(.dout(w_dff_A_9AqNdbqI6_0),.din(w_dff_A_zA4Jzm3R2_0),.clk(gclk));
	jdff dff_A_9AqNdbqI6_0(.dout(w_dff_A_ds57DFHj0_0),.din(w_dff_A_9AqNdbqI6_0),.clk(gclk));
	jdff dff_A_ds57DFHj0_0(.dout(w_dff_A_AbnSA8Wv8_0),.din(w_dff_A_ds57DFHj0_0),.clk(gclk));
	jdff dff_A_AbnSA8Wv8_0(.dout(w_dff_A_fGrLnsBi1_0),.din(w_dff_A_AbnSA8Wv8_0),.clk(gclk));
	jdff dff_A_fGrLnsBi1_0(.dout(w_dff_A_QCqrNgOf5_0),.din(w_dff_A_fGrLnsBi1_0),.clk(gclk));
	jdff dff_A_QCqrNgOf5_0(.dout(w_dff_A_DXzQ8kFL2_0),.din(w_dff_A_QCqrNgOf5_0),.clk(gclk));
	jdff dff_A_DXzQ8kFL2_0(.dout(G5308gat),.din(w_dff_A_DXzQ8kFL2_0),.clk(gclk));
	jdff dff_A_2eploXL89_2(.dout(w_dff_A_UdC9gNAX3_0),.din(w_dff_A_2eploXL89_2),.clk(gclk));
	jdff dff_A_UdC9gNAX3_0(.dout(w_dff_A_5FU17UXK0_0),.din(w_dff_A_UdC9gNAX3_0),.clk(gclk));
	jdff dff_A_5FU17UXK0_0(.dout(w_dff_A_rXGbqFUD2_0),.din(w_dff_A_5FU17UXK0_0),.clk(gclk));
	jdff dff_A_rXGbqFUD2_0(.dout(w_dff_A_JKUfwg6E9_0),.din(w_dff_A_rXGbqFUD2_0),.clk(gclk));
	jdff dff_A_JKUfwg6E9_0(.dout(w_dff_A_zJDzzZVk4_0),.din(w_dff_A_JKUfwg6E9_0),.clk(gclk));
	jdff dff_A_zJDzzZVk4_0(.dout(w_dff_A_raXzRdUI4_0),.din(w_dff_A_zJDzzZVk4_0),.clk(gclk));
	jdff dff_A_raXzRdUI4_0(.dout(w_dff_A_P1LIRME81_0),.din(w_dff_A_raXzRdUI4_0),.clk(gclk));
	jdff dff_A_P1LIRME81_0(.dout(w_dff_A_12yhYJn96_0),.din(w_dff_A_P1LIRME81_0),.clk(gclk));
	jdff dff_A_12yhYJn96_0(.dout(w_dff_A_R5faY6Ud2_0),.din(w_dff_A_12yhYJn96_0),.clk(gclk));
	jdff dff_A_R5faY6Ud2_0(.dout(w_dff_A_PzJMzCiL0_0),.din(w_dff_A_R5faY6Ud2_0),.clk(gclk));
	jdff dff_A_PzJMzCiL0_0(.dout(w_dff_A_8SeXCYUG5_0),.din(w_dff_A_PzJMzCiL0_0),.clk(gclk));
	jdff dff_A_8SeXCYUG5_0(.dout(w_dff_A_L3rDwbIB9_0),.din(w_dff_A_8SeXCYUG5_0),.clk(gclk));
	jdff dff_A_L3rDwbIB9_0(.dout(w_dff_A_VIsmJmRc0_0),.din(w_dff_A_L3rDwbIB9_0),.clk(gclk));
	jdff dff_A_VIsmJmRc0_0(.dout(w_dff_A_0qff5Z2H6_0),.din(w_dff_A_VIsmJmRc0_0),.clk(gclk));
	jdff dff_A_0qff5Z2H6_0(.dout(w_dff_A_mCB9qQjo0_0),.din(w_dff_A_0qff5Z2H6_0),.clk(gclk));
	jdff dff_A_mCB9qQjo0_0(.dout(w_dff_A_XSjJk7rX7_0),.din(w_dff_A_mCB9qQjo0_0),.clk(gclk));
	jdff dff_A_XSjJk7rX7_0(.dout(w_dff_A_1CRZe30o4_0),.din(w_dff_A_XSjJk7rX7_0),.clk(gclk));
	jdff dff_A_1CRZe30o4_0(.dout(w_dff_A_QsA7PpOn5_0),.din(w_dff_A_1CRZe30o4_0),.clk(gclk));
	jdff dff_A_QsA7PpOn5_0(.dout(w_dff_A_5UOx81rq2_0),.din(w_dff_A_QsA7PpOn5_0),.clk(gclk));
	jdff dff_A_5UOx81rq2_0(.dout(w_dff_A_8Se1HEYT5_0),.din(w_dff_A_5UOx81rq2_0),.clk(gclk));
	jdff dff_A_8Se1HEYT5_0(.dout(w_dff_A_BYiFPuHT0_0),.din(w_dff_A_8Se1HEYT5_0),.clk(gclk));
	jdff dff_A_BYiFPuHT0_0(.dout(w_dff_A_vEpqnFMt4_0),.din(w_dff_A_BYiFPuHT0_0),.clk(gclk));
	jdff dff_A_vEpqnFMt4_0(.dout(w_dff_A_vCxMsaqY4_0),.din(w_dff_A_vEpqnFMt4_0),.clk(gclk));
	jdff dff_A_vCxMsaqY4_0(.dout(w_dff_A_832snTKX6_0),.din(w_dff_A_vCxMsaqY4_0),.clk(gclk));
	jdff dff_A_832snTKX6_0(.dout(w_dff_A_slnmOMLo7_0),.din(w_dff_A_832snTKX6_0),.clk(gclk));
	jdff dff_A_slnmOMLo7_0(.dout(w_dff_A_FxSLtNzd0_0),.din(w_dff_A_slnmOMLo7_0),.clk(gclk));
	jdff dff_A_FxSLtNzd0_0(.dout(w_dff_A_y1ewrchc5_0),.din(w_dff_A_FxSLtNzd0_0),.clk(gclk));
	jdff dff_A_y1ewrchc5_0(.dout(w_dff_A_wWB6wqIg1_0),.din(w_dff_A_y1ewrchc5_0),.clk(gclk));
	jdff dff_A_wWB6wqIg1_0(.dout(w_dff_A_iTNRMvBc4_0),.din(w_dff_A_wWB6wqIg1_0),.clk(gclk));
	jdff dff_A_iTNRMvBc4_0(.dout(w_dff_A_U1rrjxAt8_0),.din(w_dff_A_iTNRMvBc4_0),.clk(gclk));
	jdff dff_A_U1rrjxAt8_0(.dout(w_dff_A_5AQSyvdS8_0),.din(w_dff_A_U1rrjxAt8_0),.clk(gclk));
	jdff dff_A_5AQSyvdS8_0(.dout(w_dff_A_wCpHk9zz9_0),.din(w_dff_A_5AQSyvdS8_0),.clk(gclk));
	jdff dff_A_wCpHk9zz9_0(.dout(w_dff_A_7g3GfLQ00_0),.din(w_dff_A_wCpHk9zz9_0),.clk(gclk));
	jdff dff_A_7g3GfLQ00_0(.dout(w_dff_A_LFKCZbbW1_0),.din(w_dff_A_7g3GfLQ00_0),.clk(gclk));
	jdff dff_A_LFKCZbbW1_0(.dout(w_dff_A_FbP4X9Z62_0),.din(w_dff_A_LFKCZbbW1_0),.clk(gclk));
	jdff dff_A_FbP4X9Z62_0(.dout(G5672gat),.din(w_dff_A_FbP4X9Z62_0),.clk(gclk));
	jdff dff_A_Y7aiHoy19_2(.dout(w_dff_A_HJm9H9L25_0),.din(w_dff_A_Y7aiHoy19_2),.clk(gclk));
	jdff dff_A_HJm9H9L25_0(.dout(w_dff_A_Xkr3vQ0J9_0),.din(w_dff_A_HJm9H9L25_0),.clk(gclk));
	jdff dff_A_Xkr3vQ0J9_0(.dout(w_dff_A_L028gl8T8_0),.din(w_dff_A_Xkr3vQ0J9_0),.clk(gclk));
	jdff dff_A_L028gl8T8_0(.dout(w_dff_A_dfwW0gsq6_0),.din(w_dff_A_L028gl8T8_0),.clk(gclk));
	jdff dff_A_dfwW0gsq6_0(.dout(w_dff_A_Lv2BQzXU1_0),.din(w_dff_A_dfwW0gsq6_0),.clk(gclk));
	jdff dff_A_Lv2BQzXU1_0(.dout(w_dff_A_6ZHXvjvc4_0),.din(w_dff_A_Lv2BQzXU1_0),.clk(gclk));
	jdff dff_A_6ZHXvjvc4_0(.dout(w_dff_A_auGLRn7K2_0),.din(w_dff_A_6ZHXvjvc4_0),.clk(gclk));
	jdff dff_A_auGLRn7K2_0(.dout(w_dff_A_R7GgadRq3_0),.din(w_dff_A_auGLRn7K2_0),.clk(gclk));
	jdff dff_A_R7GgadRq3_0(.dout(w_dff_A_9H7xgTXh8_0),.din(w_dff_A_R7GgadRq3_0),.clk(gclk));
	jdff dff_A_9H7xgTXh8_0(.dout(w_dff_A_Z5YGKIa88_0),.din(w_dff_A_9H7xgTXh8_0),.clk(gclk));
	jdff dff_A_Z5YGKIa88_0(.dout(w_dff_A_7aUXMkwn7_0),.din(w_dff_A_Z5YGKIa88_0),.clk(gclk));
	jdff dff_A_7aUXMkwn7_0(.dout(w_dff_A_QGce68b84_0),.din(w_dff_A_7aUXMkwn7_0),.clk(gclk));
	jdff dff_A_QGce68b84_0(.dout(w_dff_A_OVGBUYaL5_0),.din(w_dff_A_QGce68b84_0),.clk(gclk));
	jdff dff_A_OVGBUYaL5_0(.dout(w_dff_A_9gXgKaXw0_0),.din(w_dff_A_OVGBUYaL5_0),.clk(gclk));
	jdff dff_A_9gXgKaXw0_0(.dout(w_dff_A_Ejheg2bu0_0),.din(w_dff_A_9gXgKaXw0_0),.clk(gclk));
	jdff dff_A_Ejheg2bu0_0(.dout(w_dff_A_NCiURC5E0_0),.din(w_dff_A_Ejheg2bu0_0),.clk(gclk));
	jdff dff_A_NCiURC5E0_0(.dout(w_dff_A_BjBWmdEn8_0),.din(w_dff_A_NCiURC5E0_0),.clk(gclk));
	jdff dff_A_BjBWmdEn8_0(.dout(w_dff_A_uPUZ9dsM6_0),.din(w_dff_A_BjBWmdEn8_0),.clk(gclk));
	jdff dff_A_uPUZ9dsM6_0(.dout(w_dff_A_aYyvOcxe5_0),.din(w_dff_A_uPUZ9dsM6_0),.clk(gclk));
	jdff dff_A_aYyvOcxe5_0(.dout(w_dff_A_Nct9yvsP4_0),.din(w_dff_A_aYyvOcxe5_0),.clk(gclk));
	jdff dff_A_Nct9yvsP4_0(.dout(w_dff_A_XGldcTk53_0),.din(w_dff_A_Nct9yvsP4_0),.clk(gclk));
	jdff dff_A_XGldcTk53_0(.dout(w_dff_A_jiqcNkw18_0),.din(w_dff_A_XGldcTk53_0),.clk(gclk));
	jdff dff_A_jiqcNkw18_0(.dout(w_dff_A_VpvSj5dJ7_0),.din(w_dff_A_jiqcNkw18_0),.clk(gclk));
	jdff dff_A_VpvSj5dJ7_0(.dout(w_dff_A_ZtyUiTBv8_0),.din(w_dff_A_VpvSj5dJ7_0),.clk(gclk));
	jdff dff_A_ZtyUiTBv8_0(.dout(w_dff_A_cOrt3WrE8_0),.din(w_dff_A_ZtyUiTBv8_0),.clk(gclk));
	jdff dff_A_cOrt3WrE8_0(.dout(w_dff_A_2ZSKEUyj8_0),.din(w_dff_A_cOrt3WrE8_0),.clk(gclk));
	jdff dff_A_2ZSKEUyj8_0(.dout(w_dff_A_RqyyAWIx9_0),.din(w_dff_A_2ZSKEUyj8_0),.clk(gclk));
	jdff dff_A_RqyyAWIx9_0(.dout(w_dff_A_wErVqJat2_0),.din(w_dff_A_RqyyAWIx9_0),.clk(gclk));
	jdff dff_A_wErVqJat2_0(.dout(w_dff_A_gPzvwB2F7_0),.din(w_dff_A_wErVqJat2_0),.clk(gclk));
	jdff dff_A_gPzvwB2F7_0(.dout(w_dff_A_zVweBWe90_0),.din(w_dff_A_gPzvwB2F7_0),.clk(gclk));
	jdff dff_A_zVweBWe90_0(.dout(w_dff_A_tqURTRsT5_0),.din(w_dff_A_zVweBWe90_0),.clk(gclk));
	jdff dff_A_tqURTRsT5_0(.dout(w_dff_A_UyeQsIq00_0),.din(w_dff_A_tqURTRsT5_0),.clk(gclk));
	jdff dff_A_UyeQsIq00_0(.dout(G5971gat),.din(w_dff_A_UyeQsIq00_0),.clk(gclk));
	jdff dff_A_wIpjPOmp5_2(.dout(w_dff_A_AtNUbuPZ6_0),.din(w_dff_A_wIpjPOmp5_2),.clk(gclk));
	jdff dff_A_AtNUbuPZ6_0(.dout(w_dff_A_BJinPbYE0_0),.din(w_dff_A_AtNUbuPZ6_0),.clk(gclk));
	jdff dff_A_BJinPbYE0_0(.dout(w_dff_A_m8BbU3kq9_0),.din(w_dff_A_BJinPbYE0_0),.clk(gclk));
	jdff dff_A_m8BbU3kq9_0(.dout(w_dff_A_gYrjFtuP1_0),.din(w_dff_A_m8BbU3kq9_0),.clk(gclk));
	jdff dff_A_gYrjFtuP1_0(.dout(w_dff_A_qYnAGmuk8_0),.din(w_dff_A_gYrjFtuP1_0),.clk(gclk));
	jdff dff_A_qYnAGmuk8_0(.dout(w_dff_A_SjvbUbv44_0),.din(w_dff_A_qYnAGmuk8_0),.clk(gclk));
	jdff dff_A_SjvbUbv44_0(.dout(w_dff_A_4HVpanFh3_0),.din(w_dff_A_SjvbUbv44_0),.clk(gclk));
	jdff dff_A_4HVpanFh3_0(.dout(w_dff_A_dOzpNVyM5_0),.din(w_dff_A_4HVpanFh3_0),.clk(gclk));
	jdff dff_A_dOzpNVyM5_0(.dout(w_dff_A_oKk0otOe0_0),.din(w_dff_A_dOzpNVyM5_0),.clk(gclk));
	jdff dff_A_oKk0otOe0_0(.dout(w_dff_A_z7oGsaG63_0),.din(w_dff_A_oKk0otOe0_0),.clk(gclk));
	jdff dff_A_z7oGsaG63_0(.dout(w_dff_A_S6k56uct6_0),.din(w_dff_A_z7oGsaG63_0),.clk(gclk));
	jdff dff_A_S6k56uct6_0(.dout(w_dff_A_aazInrlM5_0),.din(w_dff_A_S6k56uct6_0),.clk(gclk));
	jdff dff_A_aazInrlM5_0(.dout(w_dff_A_GAW4iidl0_0),.din(w_dff_A_aazInrlM5_0),.clk(gclk));
	jdff dff_A_GAW4iidl0_0(.dout(w_dff_A_dyvtR10S5_0),.din(w_dff_A_GAW4iidl0_0),.clk(gclk));
	jdff dff_A_dyvtR10S5_0(.dout(w_dff_A_S4sEj3uH1_0),.din(w_dff_A_dyvtR10S5_0),.clk(gclk));
	jdff dff_A_S4sEj3uH1_0(.dout(w_dff_A_44n3h7Zq3_0),.din(w_dff_A_S4sEj3uH1_0),.clk(gclk));
	jdff dff_A_44n3h7Zq3_0(.dout(w_dff_A_i5zczjgk3_0),.din(w_dff_A_44n3h7Zq3_0),.clk(gclk));
	jdff dff_A_i5zczjgk3_0(.dout(w_dff_A_YffjuMFx5_0),.din(w_dff_A_i5zczjgk3_0),.clk(gclk));
	jdff dff_A_YffjuMFx5_0(.dout(w_dff_A_LOi9yVsM4_0),.din(w_dff_A_YffjuMFx5_0),.clk(gclk));
	jdff dff_A_LOi9yVsM4_0(.dout(w_dff_A_To8wRyRH4_0),.din(w_dff_A_LOi9yVsM4_0),.clk(gclk));
	jdff dff_A_To8wRyRH4_0(.dout(w_dff_A_Raho7Dv51_0),.din(w_dff_A_To8wRyRH4_0),.clk(gclk));
	jdff dff_A_Raho7Dv51_0(.dout(w_dff_A_TgRyoHRk7_0),.din(w_dff_A_Raho7Dv51_0),.clk(gclk));
	jdff dff_A_TgRyoHRk7_0(.dout(w_dff_A_xcMEHyMM7_0),.din(w_dff_A_TgRyoHRk7_0),.clk(gclk));
	jdff dff_A_xcMEHyMM7_0(.dout(w_dff_A_LR86UzAt5_0),.din(w_dff_A_xcMEHyMM7_0),.clk(gclk));
	jdff dff_A_LR86UzAt5_0(.dout(w_dff_A_uLTMz8aG0_0),.din(w_dff_A_LR86UzAt5_0),.clk(gclk));
	jdff dff_A_uLTMz8aG0_0(.dout(w_dff_A_9MW6V2Xb8_0),.din(w_dff_A_uLTMz8aG0_0),.clk(gclk));
	jdff dff_A_9MW6V2Xb8_0(.dout(w_dff_A_DSmQh9sG8_0),.din(w_dff_A_9MW6V2Xb8_0),.clk(gclk));
	jdff dff_A_DSmQh9sG8_0(.dout(w_dff_A_aRvqhXWD3_0),.din(w_dff_A_DSmQh9sG8_0),.clk(gclk));
	jdff dff_A_aRvqhXWD3_0(.dout(w_dff_A_ds6SS5sf0_0),.din(w_dff_A_aRvqhXWD3_0),.clk(gclk));
	jdff dff_A_ds6SS5sf0_0(.dout(G6123gat),.din(w_dff_A_ds6SS5sf0_0),.clk(gclk));
	jdff dff_A_UloyOVAB2_2(.dout(w_dff_A_Ibwud07n3_0),.din(w_dff_A_UloyOVAB2_2),.clk(gclk));
	jdff dff_A_Ibwud07n3_0(.dout(w_dff_A_o2tDNQ8L1_0),.din(w_dff_A_Ibwud07n3_0),.clk(gclk));
	jdff dff_A_o2tDNQ8L1_0(.dout(w_dff_A_cYTGn0w85_0),.din(w_dff_A_o2tDNQ8L1_0),.clk(gclk));
	jdff dff_A_cYTGn0w85_0(.dout(w_dff_A_UFDwGYHv6_0),.din(w_dff_A_cYTGn0w85_0),.clk(gclk));
	jdff dff_A_UFDwGYHv6_0(.dout(w_dff_A_hHgul19L0_0),.din(w_dff_A_UFDwGYHv6_0),.clk(gclk));
	jdff dff_A_hHgul19L0_0(.dout(w_dff_A_LxKvx0D30_0),.din(w_dff_A_hHgul19L0_0),.clk(gclk));
	jdff dff_A_LxKvx0D30_0(.dout(w_dff_A_cVgx0giF9_0),.din(w_dff_A_LxKvx0D30_0),.clk(gclk));
	jdff dff_A_cVgx0giF9_0(.dout(w_dff_A_GJ77rgCE8_0),.din(w_dff_A_cVgx0giF9_0),.clk(gclk));
	jdff dff_A_GJ77rgCE8_0(.dout(w_dff_A_qWSMzihb6_0),.din(w_dff_A_GJ77rgCE8_0),.clk(gclk));
	jdff dff_A_qWSMzihb6_0(.dout(w_dff_A_gCAghKsR7_0),.din(w_dff_A_qWSMzihb6_0),.clk(gclk));
	jdff dff_A_gCAghKsR7_0(.dout(w_dff_A_fOl9z5zx4_0),.din(w_dff_A_gCAghKsR7_0),.clk(gclk));
	jdff dff_A_fOl9z5zx4_0(.dout(w_dff_A_TsmY1Nzz1_0),.din(w_dff_A_fOl9z5zx4_0),.clk(gclk));
	jdff dff_A_TsmY1Nzz1_0(.dout(w_dff_A_2FglyBmi3_0),.din(w_dff_A_TsmY1Nzz1_0),.clk(gclk));
	jdff dff_A_2FglyBmi3_0(.dout(w_dff_A_DREhNRDh2_0),.din(w_dff_A_2FglyBmi3_0),.clk(gclk));
	jdff dff_A_DREhNRDh2_0(.dout(w_dff_A_bE73Pfdf2_0),.din(w_dff_A_DREhNRDh2_0),.clk(gclk));
	jdff dff_A_bE73Pfdf2_0(.dout(w_dff_A_jcKUJfu46_0),.din(w_dff_A_bE73Pfdf2_0),.clk(gclk));
	jdff dff_A_jcKUJfu46_0(.dout(w_dff_A_GeOOR1Kw8_0),.din(w_dff_A_jcKUJfu46_0),.clk(gclk));
	jdff dff_A_GeOOR1Kw8_0(.dout(w_dff_A_lcIhxg9N3_0),.din(w_dff_A_GeOOR1Kw8_0),.clk(gclk));
	jdff dff_A_lcIhxg9N3_0(.dout(w_dff_A_ElhITZKE8_0),.din(w_dff_A_lcIhxg9N3_0),.clk(gclk));
	jdff dff_A_ElhITZKE8_0(.dout(w_dff_A_o2wrKTho2_0),.din(w_dff_A_ElhITZKE8_0),.clk(gclk));
	jdff dff_A_o2wrKTho2_0(.dout(w_dff_A_xOGH776w5_0),.din(w_dff_A_o2wrKTho2_0),.clk(gclk));
	jdff dff_A_xOGH776w5_0(.dout(w_dff_A_9WEhy4VH4_0),.din(w_dff_A_xOGH776w5_0),.clk(gclk));
	jdff dff_A_9WEhy4VH4_0(.dout(w_dff_A_Ds88u79W7_0),.din(w_dff_A_9WEhy4VH4_0),.clk(gclk));
	jdff dff_A_Ds88u79W7_0(.dout(w_dff_A_AJXQP84v1_0),.din(w_dff_A_Ds88u79W7_0),.clk(gclk));
	jdff dff_A_AJXQP84v1_0(.dout(w_dff_A_GTAKWQ9M5_0),.din(w_dff_A_AJXQP84v1_0),.clk(gclk));
	jdff dff_A_GTAKWQ9M5_0(.dout(w_dff_A_tWXmNiTj5_0),.din(w_dff_A_GTAKWQ9M5_0),.clk(gclk));
	jdff dff_A_tWXmNiTj5_0(.dout(w_dff_A_NsXp71H74_0),.din(w_dff_A_tWXmNiTj5_0),.clk(gclk));
	jdff dff_A_NsXp71H74_0(.dout(G6150gat),.din(w_dff_A_NsXp71H74_0),.clk(gclk));
	jdff dff_A_JVdXQdwf8_2(.dout(w_dff_A_1zH06zMy1_0),.din(w_dff_A_JVdXQdwf8_2),.clk(gclk));
	jdff dff_A_1zH06zMy1_0(.dout(w_dff_A_x3873p1D6_0),.din(w_dff_A_1zH06zMy1_0),.clk(gclk));
	jdff dff_A_x3873p1D6_0(.dout(w_dff_A_kmw9SK7V6_0),.din(w_dff_A_x3873p1D6_0),.clk(gclk));
	jdff dff_A_kmw9SK7V6_0(.dout(w_dff_A_PRf3HOJn2_0),.din(w_dff_A_kmw9SK7V6_0),.clk(gclk));
	jdff dff_A_PRf3HOJn2_0(.dout(w_dff_A_2KmzX7Ao7_0),.din(w_dff_A_PRf3HOJn2_0),.clk(gclk));
	jdff dff_A_2KmzX7Ao7_0(.dout(w_dff_A_HmgcqW901_0),.din(w_dff_A_2KmzX7Ao7_0),.clk(gclk));
	jdff dff_A_HmgcqW901_0(.dout(w_dff_A_gOZAnXRZ1_0),.din(w_dff_A_HmgcqW901_0),.clk(gclk));
	jdff dff_A_gOZAnXRZ1_0(.dout(w_dff_A_wGEJkh7A6_0),.din(w_dff_A_gOZAnXRZ1_0),.clk(gclk));
	jdff dff_A_wGEJkh7A6_0(.dout(w_dff_A_b388iv6w3_0),.din(w_dff_A_wGEJkh7A6_0),.clk(gclk));
	jdff dff_A_b388iv6w3_0(.dout(w_dff_A_GDfxKoOG2_0),.din(w_dff_A_b388iv6w3_0),.clk(gclk));
	jdff dff_A_GDfxKoOG2_0(.dout(w_dff_A_0yI39X0Y7_0),.din(w_dff_A_GDfxKoOG2_0),.clk(gclk));
	jdff dff_A_0yI39X0Y7_0(.dout(w_dff_A_T2NoHBtC4_0),.din(w_dff_A_0yI39X0Y7_0),.clk(gclk));
	jdff dff_A_T2NoHBtC4_0(.dout(w_dff_A_f2cnQIQF6_0),.din(w_dff_A_T2NoHBtC4_0),.clk(gclk));
	jdff dff_A_f2cnQIQF6_0(.dout(w_dff_A_NutVUu4T7_0),.din(w_dff_A_f2cnQIQF6_0),.clk(gclk));
	jdff dff_A_NutVUu4T7_0(.dout(w_dff_A_1JVCAbvN6_0),.din(w_dff_A_NutVUu4T7_0),.clk(gclk));
	jdff dff_A_1JVCAbvN6_0(.dout(w_dff_A_vlOyO0CB5_0),.din(w_dff_A_1JVCAbvN6_0),.clk(gclk));
	jdff dff_A_vlOyO0CB5_0(.dout(w_dff_A_UflzVYxz0_0),.din(w_dff_A_vlOyO0CB5_0),.clk(gclk));
	jdff dff_A_UflzVYxz0_0(.dout(w_dff_A_H3lqwzVH4_0),.din(w_dff_A_UflzVYxz0_0),.clk(gclk));
	jdff dff_A_H3lqwzVH4_0(.dout(w_dff_A_3NCNoKhF9_0),.din(w_dff_A_H3lqwzVH4_0),.clk(gclk));
	jdff dff_A_3NCNoKhF9_0(.dout(w_dff_A_kKO7wThK9_0),.din(w_dff_A_3NCNoKhF9_0),.clk(gclk));
	jdff dff_A_kKO7wThK9_0(.dout(w_dff_A_7RolqyXH1_0),.din(w_dff_A_kKO7wThK9_0),.clk(gclk));
	jdff dff_A_7RolqyXH1_0(.dout(w_dff_A_2liRurwf0_0),.din(w_dff_A_7RolqyXH1_0),.clk(gclk));
	jdff dff_A_2liRurwf0_0(.dout(w_dff_A_kvydyW6B5_0),.din(w_dff_A_2liRurwf0_0),.clk(gclk));
	jdff dff_A_kvydyW6B5_0(.dout(w_dff_A_mEJGlNto5_0),.din(w_dff_A_kvydyW6B5_0),.clk(gclk));
	jdff dff_A_mEJGlNto5_0(.dout(w_dff_A_bu2MqwBY3_0),.din(w_dff_A_mEJGlNto5_0),.clk(gclk));
	jdff dff_A_bu2MqwBY3_0(.dout(G6160gat),.din(w_dff_A_bu2MqwBY3_0),.clk(gclk));
	jdff dff_A_CyfQuo9O5_2(.dout(w_dff_A_6QsmgJCT4_0),.din(w_dff_A_CyfQuo9O5_2),.clk(gclk));
	jdff dff_A_6QsmgJCT4_0(.dout(w_dff_A_QLgpwxGr1_0),.din(w_dff_A_6QsmgJCT4_0),.clk(gclk));
	jdff dff_A_QLgpwxGr1_0(.dout(w_dff_A_OhEcXmMH6_0),.din(w_dff_A_QLgpwxGr1_0),.clk(gclk));
	jdff dff_A_OhEcXmMH6_0(.dout(w_dff_A_f0sM1qhK3_0),.din(w_dff_A_OhEcXmMH6_0),.clk(gclk));
	jdff dff_A_f0sM1qhK3_0(.dout(w_dff_A_bKDVYeOx0_0),.din(w_dff_A_f0sM1qhK3_0),.clk(gclk));
	jdff dff_A_bKDVYeOx0_0(.dout(w_dff_A_7fgkbALf7_0),.din(w_dff_A_bKDVYeOx0_0),.clk(gclk));
	jdff dff_A_7fgkbALf7_0(.dout(w_dff_A_TzUaa2e52_0),.din(w_dff_A_7fgkbALf7_0),.clk(gclk));
	jdff dff_A_TzUaa2e52_0(.dout(w_dff_A_pumQyfY82_0),.din(w_dff_A_TzUaa2e52_0),.clk(gclk));
	jdff dff_A_pumQyfY82_0(.dout(w_dff_A_KTleP3A94_0),.din(w_dff_A_pumQyfY82_0),.clk(gclk));
	jdff dff_A_KTleP3A94_0(.dout(w_dff_A_67r9RmrV8_0),.din(w_dff_A_KTleP3A94_0),.clk(gclk));
	jdff dff_A_67r9RmrV8_0(.dout(w_dff_A_LWKSoOGR7_0),.din(w_dff_A_67r9RmrV8_0),.clk(gclk));
	jdff dff_A_LWKSoOGR7_0(.dout(w_dff_A_gzmOcQbw7_0),.din(w_dff_A_LWKSoOGR7_0),.clk(gclk));
	jdff dff_A_gzmOcQbw7_0(.dout(w_dff_A_o5JiHedi3_0),.din(w_dff_A_gzmOcQbw7_0),.clk(gclk));
	jdff dff_A_o5JiHedi3_0(.dout(w_dff_A_F6Qgon7N7_0),.din(w_dff_A_o5JiHedi3_0),.clk(gclk));
	jdff dff_A_F6Qgon7N7_0(.dout(w_dff_A_AKaExpA45_0),.din(w_dff_A_F6Qgon7N7_0),.clk(gclk));
	jdff dff_A_AKaExpA45_0(.dout(w_dff_A_rSedN8Au7_0),.din(w_dff_A_AKaExpA45_0),.clk(gclk));
	jdff dff_A_rSedN8Au7_0(.dout(w_dff_A_c36Gp4Km5_0),.din(w_dff_A_rSedN8Au7_0),.clk(gclk));
	jdff dff_A_c36Gp4Km5_0(.dout(w_dff_A_lSJDeB477_0),.din(w_dff_A_c36Gp4Km5_0),.clk(gclk));
	jdff dff_A_lSJDeB477_0(.dout(w_dff_A_Kahl07kv5_0),.din(w_dff_A_lSJDeB477_0),.clk(gclk));
	jdff dff_A_Kahl07kv5_0(.dout(w_dff_A_w7zOwIuP6_0),.din(w_dff_A_Kahl07kv5_0),.clk(gclk));
	jdff dff_A_w7zOwIuP6_0(.dout(w_dff_A_FM5DeNXp3_0),.din(w_dff_A_w7zOwIuP6_0),.clk(gclk));
	jdff dff_A_FM5DeNXp3_0(.dout(w_dff_A_2KiYTUpU1_0),.din(w_dff_A_FM5DeNXp3_0),.clk(gclk));
	jdff dff_A_2KiYTUpU1_0(.dout(w_dff_A_sD0cSjtY8_0),.din(w_dff_A_2KiYTUpU1_0),.clk(gclk));
	jdff dff_A_sD0cSjtY8_0(.dout(w_dff_A_PzmSJC3Q3_0),.din(w_dff_A_sD0cSjtY8_0),.clk(gclk));
	jdff dff_A_PzmSJC3Q3_0(.dout(G6170gat),.din(w_dff_A_PzmSJC3Q3_0),.clk(gclk));
	jdff dff_A_MLPL8Tm53_2(.dout(w_dff_A_1cUE5gY61_0),.din(w_dff_A_MLPL8Tm53_2),.clk(gclk));
	jdff dff_A_1cUE5gY61_0(.dout(w_dff_A_Nx2zFIdU0_0),.din(w_dff_A_1cUE5gY61_0),.clk(gclk));
	jdff dff_A_Nx2zFIdU0_0(.dout(w_dff_A_YbuSdF7k1_0),.din(w_dff_A_Nx2zFIdU0_0),.clk(gclk));
	jdff dff_A_YbuSdF7k1_0(.dout(w_dff_A_PliTLY538_0),.din(w_dff_A_YbuSdF7k1_0),.clk(gclk));
	jdff dff_A_PliTLY538_0(.dout(w_dff_A_IGbAi8d80_0),.din(w_dff_A_PliTLY538_0),.clk(gclk));
	jdff dff_A_IGbAi8d80_0(.dout(w_dff_A_g2HGkiKj8_0),.din(w_dff_A_IGbAi8d80_0),.clk(gclk));
	jdff dff_A_g2HGkiKj8_0(.dout(w_dff_A_5tgjmMIm3_0),.din(w_dff_A_g2HGkiKj8_0),.clk(gclk));
	jdff dff_A_5tgjmMIm3_0(.dout(w_dff_A_SHFAsCLF7_0),.din(w_dff_A_5tgjmMIm3_0),.clk(gclk));
	jdff dff_A_SHFAsCLF7_0(.dout(w_dff_A_hGGFY9fF8_0),.din(w_dff_A_SHFAsCLF7_0),.clk(gclk));
	jdff dff_A_hGGFY9fF8_0(.dout(w_dff_A_R0UyvXsu2_0),.din(w_dff_A_hGGFY9fF8_0),.clk(gclk));
	jdff dff_A_R0UyvXsu2_0(.dout(w_dff_A_Dczdn4nl2_0),.din(w_dff_A_R0UyvXsu2_0),.clk(gclk));
	jdff dff_A_Dczdn4nl2_0(.dout(w_dff_A_QhXh7hU81_0),.din(w_dff_A_Dczdn4nl2_0),.clk(gclk));
	jdff dff_A_QhXh7hU81_0(.dout(w_dff_A_Gv9ZysSp0_0),.din(w_dff_A_QhXh7hU81_0),.clk(gclk));
	jdff dff_A_Gv9ZysSp0_0(.dout(w_dff_A_gDevGOR13_0),.din(w_dff_A_Gv9ZysSp0_0),.clk(gclk));
	jdff dff_A_gDevGOR13_0(.dout(w_dff_A_p0BmH3YN4_0),.din(w_dff_A_gDevGOR13_0),.clk(gclk));
	jdff dff_A_p0BmH3YN4_0(.dout(w_dff_A_VATKnVjT6_0),.din(w_dff_A_p0BmH3YN4_0),.clk(gclk));
	jdff dff_A_VATKnVjT6_0(.dout(w_dff_A_h0gD6GjZ9_0),.din(w_dff_A_VATKnVjT6_0),.clk(gclk));
	jdff dff_A_h0gD6GjZ9_0(.dout(w_dff_A_vziCFJVO1_0),.din(w_dff_A_h0gD6GjZ9_0),.clk(gclk));
	jdff dff_A_vziCFJVO1_0(.dout(w_dff_A_Zy7WuMtb2_0),.din(w_dff_A_vziCFJVO1_0),.clk(gclk));
	jdff dff_A_Zy7WuMtb2_0(.dout(w_dff_A_aUNKkEc46_0),.din(w_dff_A_Zy7WuMtb2_0),.clk(gclk));
	jdff dff_A_aUNKkEc46_0(.dout(w_dff_A_PLHlw61x0_0),.din(w_dff_A_aUNKkEc46_0),.clk(gclk));
	jdff dff_A_PLHlw61x0_0(.dout(w_dff_A_OOLKuQoX2_0),.din(w_dff_A_PLHlw61x0_0),.clk(gclk));
	jdff dff_A_OOLKuQoX2_0(.dout(G6180gat),.din(w_dff_A_OOLKuQoX2_0),.clk(gclk));
	jdff dff_A_n713uqzH6_2(.dout(w_dff_A_1zyePD0k0_0),.din(w_dff_A_n713uqzH6_2),.clk(gclk));
	jdff dff_A_1zyePD0k0_0(.dout(w_dff_A_8EkLrFWD9_0),.din(w_dff_A_1zyePD0k0_0),.clk(gclk));
	jdff dff_A_8EkLrFWD9_0(.dout(w_dff_A_mkIIKsEY7_0),.din(w_dff_A_8EkLrFWD9_0),.clk(gclk));
	jdff dff_A_mkIIKsEY7_0(.dout(w_dff_A_VsZYpE2W6_0),.din(w_dff_A_mkIIKsEY7_0),.clk(gclk));
	jdff dff_A_VsZYpE2W6_0(.dout(w_dff_A_uG58UR1Y7_0),.din(w_dff_A_VsZYpE2W6_0),.clk(gclk));
	jdff dff_A_uG58UR1Y7_0(.dout(w_dff_A_37vdwpRh7_0),.din(w_dff_A_uG58UR1Y7_0),.clk(gclk));
	jdff dff_A_37vdwpRh7_0(.dout(w_dff_A_2VlvsQ2N5_0),.din(w_dff_A_37vdwpRh7_0),.clk(gclk));
	jdff dff_A_2VlvsQ2N5_0(.dout(w_dff_A_G4rarnNb2_0),.din(w_dff_A_2VlvsQ2N5_0),.clk(gclk));
	jdff dff_A_G4rarnNb2_0(.dout(w_dff_A_bFGW1Aob9_0),.din(w_dff_A_G4rarnNb2_0),.clk(gclk));
	jdff dff_A_bFGW1Aob9_0(.dout(w_dff_A_n1RWEHcT4_0),.din(w_dff_A_bFGW1Aob9_0),.clk(gclk));
	jdff dff_A_n1RWEHcT4_0(.dout(w_dff_A_Q1Hj46AI5_0),.din(w_dff_A_n1RWEHcT4_0),.clk(gclk));
	jdff dff_A_Q1Hj46AI5_0(.dout(w_dff_A_2r7e5l4a2_0),.din(w_dff_A_Q1Hj46AI5_0),.clk(gclk));
	jdff dff_A_2r7e5l4a2_0(.dout(w_dff_A_XKnSYu4M6_0),.din(w_dff_A_2r7e5l4a2_0),.clk(gclk));
	jdff dff_A_XKnSYu4M6_0(.dout(w_dff_A_K1QTPPHV9_0),.din(w_dff_A_XKnSYu4M6_0),.clk(gclk));
	jdff dff_A_K1QTPPHV9_0(.dout(w_dff_A_RRmvn2mA0_0),.din(w_dff_A_K1QTPPHV9_0),.clk(gclk));
	jdff dff_A_RRmvn2mA0_0(.dout(w_dff_A_Qp7kegdR0_0),.din(w_dff_A_RRmvn2mA0_0),.clk(gclk));
	jdff dff_A_Qp7kegdR0_0(.dout(w_dff_A_SxJHOqFh5_0),.din(w_dff_A_Qp7kegdR0_0),.clk(gclk));
	jdff dff_A_SxJHOqFh5_0(.dout(w_dff_A_7GqKYvYY1_0),.din(w_dff_A_SxJHOqFh5_0),.clk(gclk));
	jdff dff_A_7GqKYvYY1_0(.dout(w_dff_A_yCy4gWd84_0),.din(w_dff_A_7GqKYvYY1_0),.clk(gclk));
	jdff dff_A_yCy4gWd84_0(.dout(w_dff_A_IR1hYRdO8_0),.din(w_dff_A_yCy4gWd84_0),.clk(gclk));
	jdff dff_A_IR1hYRdO8_0(.dout(G6190gat),.din(w_dff_A_IR1hYRdO8_0),.clk(gclk));
	jdff dff_A_uHImcr829_2(.dout(w_dff_A_PuntIyzd3_0),.din(w_dff_A_uHImcr829_2),.clk(gclk));
	jdff dff_A_PuntIyzd3_0(.dout(w_dff_A_9hC8YyDW0_0),.din(w_dff_A_PuntIyzd3_0),.clk(gclk));
	jdff dff_A_9hC8YyDW0_0(.dout(w_dff_A_MAVKxQfy9_0),.din(w_dff_A_9hC8YyDW0_0),.clk(gclk));
	jdff dff_A_MAVKxQfy9_0(.dout(w_dff_A_OU1juCpu3_0),.din(w_dff_A_MAVKxQfy9_0),.clk(gclk));
	jdff dff_A_OU1juCpu3_0(.dout(w_dff_A_vQsYsFQ84_0),.din(w_dff_A_OU1juCpu3_0),.clk(gclk));
	jdff dff_A_vQsYsFQ84_0(.dout(w_dff_A_6JaZ3H5x0_0),.din(w_dff_A_vQsYsFQ84_0),.clk(gclk));
	jdff dff_A_6JaZ3H5x0_0(.dout(w_dff_A_L0aAgzoy5_0),.din(w_dff_A_6JaZ3H5x0_0),.clk(gclk));
	jdff dff_A_L0aAgzoy5_0(.dout(w_dff_A_YqFbGUtE6_0),.din(w_dff_A_L0aAgzoy5_0),.clk(gclk));
	jdff dff_A_YqFbGUtE6_0(.dout(w_dff_A_3chAuc6C7_0),.din(w_dff_A_YqFbGUtE6_0),.clk(gclk));
	jdff dff_A_3chAuc6C7_0(.dout(w_dff_A_gJqYnwRf4_0),.din(w_dff_A_3chAuc6C7_0),.clk(gclk));
	jdff dff_A_gJqYnwRf4_0(.dout(w_dff_A_HyR4pv8i8_0),.din(w_dff_A_gJqYnwRf4_0),.clk(gclk));
	jdff dff_A_HyR4pv8i8_0(.dout(w_dff_A_H31sQU3z4_0),.din(w_dff_A_HyR4pv8i8_0),.clk(gclk));
	jdff dff_A_H31sQU3z4_0(.dout(w_dff_A_VXuuPWYE1_0),.din(w_dff_A_H31sQU3z4_0),.clk(gclk));
	jdff dff_A_VXuuPWYE1_0(.dout(w_dff_A_cEQ7hE1d9_0),.din(w_dff_A_VXuuPWYE1_0),.clk(gclk));
	jdff dff_A_cEQ7hE1d9_0(.dout(w_dff_A_fWBN7M7R5_0),.din(w_dff_A_cEQ7hE1d9_0),.clk(gclk));
	jdff dff_A_fWBN7M7R5_0(.dout(w_dff_A_3IpZdmmt8_0),.din(w_dff_A_fWBN7M7R5_0),.clk(gclk));
	jdff dff_A_3IpZdmmt8_0(.dout(w_dff_A_fsnear8F0_0),.din(w_dff_A_3IpZdmmt8_0),.clk(gclk));
	jdff dff_A_fsnear8F0_0(.dout(w_dff_A_peG6gmsc2_0),.din(w_dff_A_fsnear8F0_0),.clk(gclk));
	jdff dff_A_peG6gmsc2_0(.dout(G6200gat),.din(w_dff_A_peG6gmsc2_0),.clk(gclk));
	jdff dff_A_IVpIwNKv9_2(.dout(w_dff_A_6hil7dpQ8_0),.din(w_dff_A_IVpIwNKv9_2),.clk(gclk));
	jdff dff_A_6hil7dpQ8_0(.dout(w_dff_A_z9BO7XGP7_0),.din(w_dff_A_6hil7dpQ8_0),.clk(gclk));
	jdff dff_A_z9BO7XGP7_0(.dout(w_dff_A_iC1YrsCy7_0),.din(w_dff_A_z9BO7XGP7_0),.clk(gclk));
	jdff dff_A_iC1YrsCy7_0(.dout(w_dff_A_DvFndVcE9_0),.din(w_dff_A_iC1YrsCy7_0),.clk(gclk));
	jdff dff_A_DvFndVcE9_0(.dout(w_dff_A_ODlpoHVs5_0),.din(w_dff_A_DvFndVcE9_0),.clk(gclk));
	jdff dff_A_ODlpoHVs5_0(.dout(w_dff_A_XfuX7JNC6_0),.din(w_dff_A_ODlpoHVs5_0),.clk(gclk));
	jdff dff_A_XfuX7JNC6_0(.dout(w_dff_A_xbvxqzN21_0),.din(w_dff_A_XfuX7JNC6_0),.clk(gclk));
	jdff dff_A_xbvxqzN21_0(.dout(w_dff_A_HqOzHMBf3_0),.din(w_dff_A_xbvxqzN21_0),.clk(gclk));
	jdff dff_A_HqOzHMBf3_0(.dout(w_dff_A_qWw2ImB81_0),.din(w_dff_A_HqOzHMBf3_0),.clk(gclk));
	jdff dff_A_qWw2ImB81_0(.dout(w_dff_A_MTKcdpiO3_0),.din(w_dff_A_qWw2ImB81_0),.clk(gclk));
	jdff dff_A_MTKcdpiO3_0(.dout(w_dff_A_ybVgRRSY6_0),.din(w_dff_A_MTKcdpiO3_0),.clk(gclk));
	jdff dff_A_ybVgRRSY6_0(.dout(w_dff_A_iGfZIBto7_0),.din(w_dff_A_ybVgRRSY6_0),.clk(gclk));
	jdff dff_A_iGfZIBto7_0(.dout(w_dff_A_EKf6nyf00_0),.din(w_dff_A_iGfZIBto7_0),.clk(gclk));
	jdff dff_A_EKf6nyf00_0(.dout(w_dff_A_3bgR5Esy3_0),.din(w_dff_A_EKf6nyf00_0),.clk(gclk));
	jdff dff_A_3bgR5Esy3_0(.dout(w_dff_A_HgzcCpoD4_0),.din(w_dff_A_3bgR5Esy3_0),.clk(gclk));
	jdff dff_A_HgzcCpoD4_0(.dout(w_dff_A_qEnI3H503_0),.din(w_dff_A_HgzcCpoD4_0),.clk(gclk));
	jdff dff_A_qEnI3H503_0(.dout(G6210gat),.din(w_dff_A_qEnI3H503_0),.clk(gclk));
	jdff dff_A_J9KkTH2x8_2(.dout(w_dff_A_3TFql5wV6_0),.din(w_dff_A_J9KkTH2x8_2),.clk(gclk));
	jdff dff_A_3TFql5wV6_0(.dout(w_dff_A_Cg14zy3H6_0),.din(w_dff_A_3TFql5wV6_0),.clk(gclk));
	jdff dff_A_Cg14zy3H6_0(.dout(w_dff_A_TKmPl4h12_0),.din(w_dff_A_Cg14zy3H6_0),.clk(gclk));
	jdff dff_A_TKmPl4h12_0(.dout(w_dff_A_BMz3zrYF4_0),.din(w_dff_A_TKmPl4h12_0),.clk(gclk));
	jdff dff_A_BMz3zrYF4_0(.dout(w_dff_A_xjsRzz3e0_0),.din(w_dff_A_BMz3zrYF4_0),.clk(gclk));
	jdff dff_A_xjsRzz3e0_0(.dout(w_dff_A_HPuBL4Zj8_0),.din(w_dff_A_xjsRzz3e0_0),.clk(gclk));
	jdff dff_A_HPuBL4Zj8_0(.dout(w_dff_A_rAePVV5H4_0),.din(w_dff_A_HPuBL4Zj8_0),.clk(gclk));
	jdff dff_A_rAePVV5H4_0(.dout(w_dff_A_GC3C7Ipp8_0),.din(w_dff_A_rAePVV5H4_0),.clk(gclk));
	jdff dff_A_GC3C7Ipp8_0(.dout(w_dff_A_XICinNMW7_0),.din(w_dff_A_GC3C7Ipp8_0),.clk(gclk));
	jdff dff_A_XICinNMW7_0(.dout(w_dff_A_jWnHqDMP3_0),.din(w_dff_A_XICinNMW7_0),.clk(gclk));
	jdff dff_A_jWnHqDMP3_0(.dout(w_dff_A_7YPS7KFr9_0),.din(w_dff_A_jWnHqDMP3_0),.clk(gclk));
	jdff dff_A_7YPS7KFr9_0(.dout(w_dff_A_vqTTAhJa6_0),.din(w_dff_A_7YPS7KFr9_0),.clk(gclk));
	jdff dff_A_vqTTAhJa6_0(.dout(w_dff_A_TI6FyUpQ0_0),.din(w_dff_A_vqTTAhJa6_0),.clk(gclk));
	jdff dff_A_TI6FyUpQ0_0(.dout(w_dff_A_MzFxhQaF3_0),.din(w_dff_A_TI6FyUpQ0_0),.clk(gclk));
	jdff dff_A_MzFxhQaF3_0(.dout(G6220gat),.din(w_dff_A_MzFxhQaF3_0),.clk(gclk));
	jdff dff_A_SiAvJkIH2_2(.dout(w_dff_A_DMQvcXa57_0),.din(w_dff_A_SiAvJkIH2_2),.clk(gclk));
	jdff dff_A_DMQvcXa57_0(.dout(w_dff_A_iaGQDlki6_0),.din(w_dff_A_DMQvcXa57_0),.clk(gclk));
	jdff dff_A_iaGQDlki6_0(.dout(w_dff_A_C5FUBbPf2_0),.din(w_dff_A_iaGQDlki6_0),.clk(gclk));
	jdff dff_A_C5FUBbPf2_0(.dout(w_dff_A_Jirr21g67_0),.din(w_dff_A_C5FUBbPf2_0),.clk(gclk));
	jdff dff_A_Jirr21g67_0(.dout(w_dff_A_5cSz67HW5_0),.din(w_dff_A_Jirr21g67_0),.clk(gclk));
	jdff dff_A_5cSz67HW5_0(.dout(w_dff_A_pVwqnoch6_0),.din(w_dff_A_5cSz67HW5_0),.clk(gclk));
	jdff dff_A_pVwqnoch6_0(.dout(w_dff_A_jPJSMjq68_0),.din(w_dff_A_pVwqnoch6_0),.clk(gclk));
	jdff dff_A_jPJSMjq68_0(.dout(w_dff_A_CzVrvDbH0_0),.din(w_dff_A_jPJSMjq68_0),.clk(gclk));
	jdff dff_A_CzVrvDbH0_0(.dout(w_dff_A_sNlDG9Kl8_0),.din(w_dff_A_CzVrvDbH0_0),.clk(gclk));
	jdff dff_A_sNlDG9Kl8_0(.dout(w_dff_A_CKVihfhb3_0),.din(w_dff_A_sNlDG9Kl8_0),.clk(gclk));
	jdff dff_A_CKVihfhb3_0(.dout(w_dff_A_OxoA2Dmw7_0),.din(w_dff_A_CKVihfhb3_0),.clk(gclk));
	jdff dff_A_OxoA2Dmw7_0(.dout(w_dff_A_MJmxjNUa6_0),.din(w_dff_A_OxoA2Dmw7_0),.clk(gclk));
	jdff dff_A_MJmxjNUa6_0(.dout(G6230gat),.din(w_dff_A_MJmxjNUa6_0),.clk(gclk));
	jdff dff_A_iPOTMMlN8_2(.dout(w_dff_A_Mcel7Ici0_0),.din(w_dff_A_iPOTMMlN8_2),.clk(gclk));
	jdff dff_A_Mcel7Ici0_0(.dout(w_dff_A_mLuGV0qZ8_0),.din(w_dff_A_Mcel7Ici0_0),.clk(gclk));
	jdff dff_A_mLuGV0qZ8_0(.dout(w_dff_A_RTLILm7e3_0),.din(w_dff_A_mLuGV0qZ8_0),.clk(gclk));
	jdff dff_A_RTLILm7e3_0(.dout(w_dff_A_PguZKwg88_0),.din(w_dff_A_RTLILm7e3_0),.clk(gclk));
	jdff dff_A_PguZKwg88_0(.dout(w_dff_A_NUqmzJqp4_0),.din(w_dff_A_PguZKwg88_0),.clk(gclk));
	jdff dff_A_NUqmzJqp4_0(.dout(w_dff_A_q8EXGjNW0_0),.din(w_dff_A_NUqmzJqp4_0),.clk(gclk));
	jdff dff_A_q8EXGjNW0_0(.dout(w_dff_A_z8DsJDDU7_0),.din(w_dff_A_q8EXGjNW0_0),.clk(gclk));
	jdff dff_A_z8DsJDDU7_0(.dout(w_dff_A_1SYlCHVO7_0),.din(w_dff_A_z8DsJDDU7_0),.clk(gclk));
	jdff dff_A_1SYlCHVO7_0(.dout(w_dff_A_KvCKM18V3_0),.din(w_dff_A_1SYlCHVO7_0),.clk(gclk));
	jdff dff_A_KvCKM18V3_0(.dout(w_dff_A_HmcJ3q5s3_0),.din(w_dff_A_KvCKM18V3_0),.clk(gclk));
	jdff dff_A_HmcJ3q5s3_0(.dout(G6240gat),.din(w_dff_A_HmcJ3q5s3_0),.clk(gclk));
	jdff dff_A_ZynMqCJa0_2(.dout(w_dff_A_EfzsPbLb3_0),.din(w_dff_A_ZynMqCJa0_2),.clk(gclk));
	jdff dff_A_EfzsPbLb3_0(.dout(w_dff_A_lzkEW5DO4_0),.din(w_dff_A_EfzsPbLb3_0),.clk(gclk));
	jdff dff_A_lzkEW5DO4_0(.dout(w_dff_A_T3BcHT3C2_0),.din(w_dff_A_lzkEW5DO4_0),.clk(gclk));
	jdff dff_A_T3BcHT3C2_0(.dout(w_dff_A_hHw8iqDQ9_0),.din(w_dff_A_T3BcHT3C2_0),.clk(gclk));
	jdff dff_A_hHw8iqDQ9_0(.dout(w_dff_A_LH6lzpir2_0),.din(w_dff_A_hHw8iqDQ9_0),.clk(gclk));
	jdff dff_A_LH6lzpir2_0(.dout(w_dff_A_Wl1wMhsX8_0),.din(w_dff_A_LH6lzpir2_0),.clk(gclk));
	jdff dff_A_Wl1wMhsX8_0(.dout(w_dff_A_O7PPRNrY9_0),.din(w_dff_A_Wl1wMhsX8_0),.clk(gclk));
	jdff dff_A_O7PPRNrY9_0(.dout(w_dff_A_aqTIs5RT3_0),.din(w_dff_A_O7PPRNrY9_0),.clk(gclk));
	jdff dff_A_aqTIs5RT3_0(.dout(G6250gat),.din(w_dff_A_aqTIs5RT3_0),.clk(gclk));
	jdff dff_A_DQBFPbwp8_2(.dout(w_dff_A_7Eum09t90_0),.din(w_dff_A_DQBFPbwp8_2),.clk(gclk));
	jdff dff_A_7Eum09t90_0(.dout(w_dff_A_1DK9Zo400_0),.din(w_dff_A_7Eum09t90_0),.clk(gclk));
	jdff dff_A_1DK9Zo400_0(.dout(w_dff_A_u1PNOSYe3_0),.din(w_dff_A_1DK9Zo400_0),.clk(gclk));
	jdff dff_A_u1PNOSYe3_0(.dout(w_dff_A_brfkCIms5_0),.din(w_dff_A_u1PNOSYe3_0),.clk(gclk));
	jdff dff_A_brfkCIms5_0(.dout(w_dff_A_GclQeXAU6_0),.din(w_dff_A_brfkCIms5_0),.clk(gclk));
	jdff dff_A_GclQeXAU6_0(.dout(w_dff_A_Tyc7mDF21_0),.din(w_dff_A_GclQeXAU6_0),.clk(gclk));
	jdff dff_A_Tyc7mDF21_0(.dout(G6260gat),.din(w_dff_A_Tyc7mDF21_0),.clk(gclk));
	jdff dff_A_6HD4c7010_2(.dout(w_dff_A_H101jjJm2_0),.din(w_dff_A_6HD4c7010_2),.clk(gclk));
	jdff dff_A_H101jjJm2_0(.dout(w_dff_A_iCKC4Clq9_0),.din(w_dff_A_H101jjJm2_0),.clk(gclk));
	jdff dff_A_iCKC4Clq9_0(.dout(w_dff_A_NHm2bFxY2_0),.din(w_dff_A_iCKC4Clq9_0),.clk(gclk));
	jdff dff_A_NHm2bFxY2_0(.dout(w_dff_A_equOPP612_0),.din(w_dff_A_NHm2bFxY2_0),.clk(gclk));
	jdff dff_A_equOPP612_0(.dout(G6270gat),.din(w_dff_A_equOPP612_0),.clk(gclk));
	jdff dff_A_onIovUsr0_2(.dout(w_dff_A_ghfVfWMO9_0),.din(w_dff_A_onIovUsr0_2),.clk(gclk));
	jdff dff_A_ghfVfWMO9_0(.dout(w_dff_A_SMJRn6R92_0),.din(w_dff_A_ghfVfWMO9_0),.clk(gclk));
	jdff dff_A_SMJRn6R92_0(.dout(G6280gat),.din(w_dff_A_SMJRn6R92_0),.clk(gclk));
	jdff dff_A_mVaqxWQK4_2(.dout(G6288gat),.din(w_dff_A_mVaqxWQK4_2),.clk(gclk));
endmodule

