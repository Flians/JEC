// Benchmark "c3540" written by ABC on Sun May 24 21:27:50 2020

module c3540 ( 
    G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
    G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200,
    G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274,
    G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698,
    G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107,
    G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
    G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270,
    G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire n72, n73, n74, n75, n76, n77, n79, n80, n81, n82, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n124, n125, n126,
    n127, n128, n129, n130, n132, n133, n134, n135, n136, n137, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n517, n518, n519, n520, n521, n522, n523, n524, n525,
    n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
    n575, n576, n577, n578, n579, n580, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n610, n611, n612,
    n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
    n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
    n795, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
    n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1170, n1171, n1172, n1173, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186;
  jnot g0000(.din(G77), .dout(n72));
  jnot g0001(.din(G50), .dout(n73));
  jnot g0002(.din(G58), .dout(n74));
  jnot g0003(.din(G68), .dout(n75));
  jand g0004(.dina(n75), .dinb(n74), .dout(n76));
  jand g0005(.dina(n76), .dinb(n73), .dout(n77));
  jand g0006(.dina(n77), .dinb(n72), .dout(G353));
  jnot g0007(.din(G87), .dout(n79));
  jnot g0008(.din(G97), .dout(n80));
  jnot g0009(.din(G107), .dout(n81));
  jand g0010(.dina(n81), .dinb(n80), .dout(n82));
  jor  g0011(.dina(n82), .dinb(n79), .dout(G355));
  jnot g0012(.din(G250), .dout(n84));
  jnot g0013(.din(G257), .dout(n85));
  jnot g0014(.din(G264), .dout(n86));
  jand g0015(.dina(n86), .dinb(n85), .dout(n87));
  jor  g0016(.dina(n87), .dinb(n84), .dout(n88));
  jnot g0017(.din(G13), .dout(n89));
  jand g0018(.dina(n89), .dinb(G1), .dout(n90));
  jand g0019(.dina(n90), .dinb(G20), .dout(n91));
  jand g0020(.dina(n91), .dinb(n88), .dout(n92));
  jor  g0021(.dina(n85), .dinb(n80), .dout(n93));
  jnot g0022(.din(G244), .dout(n94));
  jor  g0023(.dina(n94), .dinb(n72), .dout(n95));
  jnot g0024(.din(G238), .dout(n96));
  jor  g0025(.dina(n96), .dinb(n75), .dout(n97));
  jand g0026(.dina(n97), .dinb(n95), .dout(n98));
  jnot g0027(.din(G226), .dout(n99));
  jor  g0028(.dina(n99), .dinb(n73), .dout(n100));
  jand g0029(.dina(n100), .dinb(n98), .dout(n101));
  jand g0030(.dina(n101), .dinb(n93), .dout(n102));
  jnot g0031(.din(G232), .dout(n103));
  jor  g0032(.dina(n103), .dinb(n74), .dout(n104));
  jnot g0033(.din(G116), .dout(n105));
  jnot g0034(.din(G270), .dout(n106));
  jor  g0035(.dina(n106), .dinb(n105), .dout(n107));
  jand g0036(.dina(n107), .dinb(n104), .dout(n108));
  jor  g0037(.dina(n86), .dinb(n81), .dout(n109));
  jand g0038(.dina(n109), .dinb(n108), .dout(n110));
  jand g0039(.dina(G20), .dinb(G1), .dout(n111));
  jnot g0040(.din(n111), .dout(n112));
  jor  g0041(.dina(n84), .dinb(n79), .dout(n113));
  jand g0042(.dina(n113), .dinb(n112), .dout(n114));
  jand g0043(.dina(n114), .dinb(n110), .dout(n115));
  jand g0044(.dina(n115), .dinb(n102), .dout(n116));
  jnot g0045(.din(n76), .dout(n117));
  jand g0046(.dina(n117), .dinb(G50), .dout(n118));
  jnot g0047(.din(n118), .dout(n119));
  jand g0048(.dina(n111), .dinb(G13), .dout(n120));
  jand g0049(.dina(n120), .dinb(n119), .dout(n121));
  jor  g0050(.dina(n121), .dinb(n116), .dout(n122));
  jor  g0051(.dina(n122), .dinb(n92), .dout(G361));
  jxor g0052(.dina(G270), .dinb(n86), .dout(n124));
  jxor g0053(.dina(G257), .dinb(G250), .dout(n125));
  jxor g0054(.dina(n125), .dinb(n124), .dout(n126));
  jnot g0055(.din(n126), .dout(n127));
  jxor g0056(.dina(G244), .dinb(n96), .dout(n128));
  jxor g0057(.dina(G232), .dinb(G226), .dout(n129));
  jxor g0058(.dina(n129), .dinb(n128), .dout(n130));
  jxor g0059(.dina(n130), .dinb(n127), .dout(G358));
  jxor g0060(.dina(G58), .dinb(G50), .dout(n132));
  jxor g0061(.dina(G77), .dinb(G68), .dout(n133));
  jxor g0062(.dina(n133), .dinb(n132), .dout(n134));
  jxor g0063(.dina(G116), .dinb(n81), .dout(n135));
  jxor g0064(.dina(G97), .dinb(G87), .dout(n136));
  jxor g0065(.dina(n136), .dinb(n135), .dout(n137));
  jxor g0066(.dina(n137), .dinb(n134), .dout(G351));
  jand g0067(.dina(G13), .dinb(G1), .dout(n139));
  jand g0068(.dina(n111), .dinb(G33), .dout(n140));
  jor  g0069(.dina(n140), .dinb(n139), .dout(n141));
  jnot g0070(.din(G1), .dout(n142));
  jand g0071(.dina(G13), .dinb(n142), .dout(n143));
  jand g0072(.dina(n143), .dinb(G20), .dout(n144));
  jor  g0073(.dina(n144), .dinb(n141), .dout(n145));
  jand g0074(.dina(G33), .dinb(n142), .dout(n146));
  jor  g0075(.dina(n146), .dinb(n145), .dout(n147));
  jnot g0076(.din(n147), .dout(n148));
  jand g0077(.dina(n148), .dinb(G116), .dout(n149));
  jand g0078(.dina(G116), .dinb(G20), .dout(n150));
  jnot g0079(.din(G20), .dout(n151));
  jand g0080(.dina(G283), .dinb(G33), .dout(n152));
  jnot g0081(.din(G33), .dout(n153));
  jand g0082(.dina(G97), .dinb(n153), .dout(n154));
  jor  g0083(.dina(n154), .dinb(n152), .dout(n155));
  jand g0084(.dina(n155), .dinb(n151), .dout(n156));
  jor  g0085(.dina(n156), .dinb(n150), .dout(n157));
  jand g0086(.dina(n157), .dinb(n141), .dout(n158));
  jand g0087(.dina(n144), .dinb(n105), .dout(n159));
  jor  g0088(.dina(n159), .dinb(n158), .dout(n160));
  jor  g0089(.dina(n160), .dinb(n149), .dout(n161));
  jnot g0090(.din(n161), .dout(n162));
  jnot g0091(.din(G41), .dout(n163));
  jand g0092(.dina(G45), .dinb(n142), .dout(n164));
  jand g0093(.dina(n164), .dinb(n163), .dout(n165));
  jnot g0094(.din(n139), .dout(n166));
  jand g0095(.dina(G41), .dinb(G33), .dout(n167));
  jor  g0096(.dina(n167), .dinb(n166), .dout(n168));
  jand g0097(.dina(n168), .dinb(G274), .dout(n169));
  jand g0098(.dina(n169), .dinb(n165), .dout(n170));
  jnot g0099(.din(n167), .dout(n171));
  jand g0100(.dina(n171), .dinb(n139), .dout(n172));
  jand g0101(.dina(G1698), .dinb(n153), .dout(n173));
  jand g0102(.dina(n173), .dinb(G264), .dout(n174));
  jand g0103(.dina(G303), .dinb(G33), .dout(n175));
  jnot g0104(.din(G1698), .dout(n176));
  jand g0105(.dina(n176), .dinb(n153), .dout(n177));
  jand g0106(.dina(n177), .dinb(G257), .dout(n178));
  jor  g0107(.dina(n178), .dinb(n175), .dout(n179));
  jor  g0108(.dina(n179), .dinb(n174), .dout(n180));
  jand g0109(.dina(n180), .dinb(n172), .dout(n181));
  jnot g0110(.din(n165), .dout(n182));
  jand g0111(.dina(n168), .dinb(G270), .dout(n183));
  jand g0112(.dina(n183), .dinb(n182), .dout(n184));
  jor  g0113(.dina(n184), .dinb(n181), .dout(n185));
  jor  g0114(.dina(n185), .dinb(n170), .dout(n186));
  jand g0115(.dina(n186), .dinb(G169), .dout(n187));
  jnot g0116(.din(n187), .dout(n188));
  jnot g0117(.din(G179), .dout(n189));
  jor  g0118(.dina(n186), .dinb(n189), .dout(n190));
  jand g0119(.dina(n190), .dinb(n188), .dout(n191));
  jor  g0120(.dina(n191), .dinb(n162), .dout(n192));
  jand g0121(.dina(n186), .dinb(G200), .dout(n193));
  jnot g0122(.din(n186), .dout(n194));
  jand g0123(.dina(n194), .dinb(G190), .dout(n195));
  jor  g0124(.dina(n195), .dinb(n161), .dout(n196));
  jor  g0125(.dina(n196), .dinb(n193), .dout(n197));
  jand g0126(.dina(n197), .dinb(n192), .dout(n198));
  jnot g0127(.din(G169), .dout(n199));
  jand g0128(.dina(n168), .dinb(G264), .dout(n200));
  jand g0129(.dina(n200), .dinb(n182), .dout(n201));
  jand g0130(.dina(n173), .dinb(G257), .dout(n202));
  jand g0131(.dina(G294), .dinb(G33), .dout(n203));
  jnot g0132(.din(n203), .dout(n204));
  jor  g0133(.dina(G1698), .dinb(G33), .dout(n205));
  jor  g0134(.dina(n205), .dinb(n84), .dout(n206));
  jand g0135(.dina(n206), .dinb(n204), .dout(n207));
  jnot g0136(.din(n207), .dout(n208));
  jor  g0137(.dina(n208), .dinb(n202), .dout(n209));
  jand g0138(.dina(n209), .dinb(n172), .dout(n210));
  jor  g0139(.dina(n210), .dinb(n170), .dout(n211));
  jor  g0140(.dina(n211), .dinb(n201), .dout(n212));
  jand g0141(.dina(n212), .dinb(n199), .dout(n213));
  jand g0142(.dina(n148), .dinb(G107), .dout(n214));
  jor  g0143(.dina(n140), .dinb(G13), .dout(n215));
  jand g0144(.dina(n81), .dinb(G20), .dout(n216));
  jand g0145(.dina(n216), .dinb(n215), .dout(n217));
  jand g0146(.dina(G116), .dinb(G33), .dout(n218));
  jand g0147(.dina(G87), .dinb(n153), .dout(n219));
  jor  g0148(.dina(n219), .dinb(n218), .dout(n220));
  jand g0149(.dina(n220), .dinb(n141), .dout(n221));
  jand g0150(.dina(n221), .dinb(n151), .dout(n222));
  jor  g0151(.dina(n222), .dinb(n217), .dout(n223));
  jor  g0152(.dina(n223), .dinb(n214), .dout(n224));
  jnot g0153(.din(n224), .dout(n225));
  jnot g0154(.din(n201), .dout(n226));
  jnot g0155(.din(G274), .dout(n227));
  jor  g0156(.dina(n172), .dinb(n227), .dout(n228));
  jor  g0157(.dina(n228), .dinb(n182), .dout(n229));
  jnot g0158(.din(n202), .dout(n230));
  jand g0159(.dina(n207), .dinb(n230), .dout(n231));
  jor  g0160(.dina(n231), .dinb(n168), .dout(n232));
  jand g0161(.dina(n232), .dinb(n229), .dout(n233));
  jand g0162(.dina(n233), .dinb(n226), .dout(n234));
  jand g0163(.dina(n234), .dinb(n189), .dout(n235));
  jor  g0164(.dina(n235), .dinb(n225), .dout(n236));
  jor  g0165(.dina(n236), .dinb(n213), .dout(n237));
  jand g0166(.dina(n234), .dinb(G190), .dout(n238));
  jand g0167(.dina(n212), .dinb(G200), .dout(n239));
  jor  g0168(.dina(n239), .dinb(n224), .dout(n240));
  jor  g0169(.dina(n240), .dinb(n238), .dout(n241));
  jand g0170(.dina(n241), .dinb(n237), .dout(n242));
  jand g0171(.dina(n173), .dinb(G244), .dout(n243));
  jnot g0172(.din(n243), .dout(n244));
  jnot g0173(.din(n218), .dout(n245));
  jor  g0174(.dina(n205), .dinb(n96), .dout(n246));
  jand g0175(.dina(n246), .dinb(n245), .dout(n247));
  jand g0176(.dina(n247), .dinb(n244), .dout(n248));
  jand g0177(.dina(n248), .dinb(n172), .dout(n249));
  jor  g0178(.dina(n164), .dinb(n84), .dout(n250));
  jand g0179(.dina(n164), .dinb(G274), .dout(n251));
  jnot g0180(.din(n251), .dout(n252));
  jand g0181(.dina(n252), .dinb(n250), .dout(n253));
  jand g0182(.dina(n253), .dinb(n168), .dout(n254));
  jor  g0183(.dina(n254), .dinb(n249), .dout(n255));
  jand g0184(.dina(n255), .dinb(n189), .dout(n256));
  jor  g0185(.dina(n147), .dinb(n79), .dout(n257));
  jand g0186(.dina(n80), .dinb(n79), .dout(n258));
  jand g0187(.dina(n258), .dinb(n81), .dout(n259));
  jand g0188(.dina(n259), .dinb(G20), .dout(n260));
  jnot g0189(.din(n141), .dout(n261));
  jand g0190(.dina(G97), .dinb(G33), .dout(n262));
  jnot g0191(.din(n262), .dout(n263));
  jor  g0192(.dina(n75), .dinb(G33), .dout(n264));
  jand g0193(.dina(n264), .dinb(n151), .dout(n265));
  jand g0194(.dina(n265), .dinb(n263), .dout(n266));
  jor  g0195(.dina(n266), .dinb(n261), .dout(n267));
  jor  g0196(.dina(n267), .dinb(n260), .dout(n268));
  jand g0197(.dina(n144), .dinb(n79), .dout(n269));
  jnot g0198(.din(n269), .dout(n270));
  jand g0199(.dina(n270), .dinb(n268), .dout(n271));
  jand g0200(.dina(n271), .dinb(n257), .dout(n272));
  jnot g0201(.din(n247), .dout(n273));
  jor  g0202(.dina(n273), .dinb(n243), .dout(n274));
  jor  g0203(.dina(n274), .dinb(n168), .dout(n275));
  jnot g0204(.din(n250), .dout(n276));
  jor  g0205(.dina(n251), .dinb(n276), .dout(n277));
  jor  g0206(.dina(n277), .dinb(n172), .dout(n278));
  jand g0207(.dina(n278), .dinb(n275), .dout(n279));
  jand g0208(.dina(n279), .dinb(n199), .dout(n280));
  jor  g0209(.dina(n280), .dinb(n272), .dout(n281));
  jor  g0210(.dina(n281), .dinb(n256), .dout(n282));
  jand g0211(.dina(n279), .dinb(G200), .dout(n283));
  jnot g0212(.din(n257), .dout(n284));
  jnot g0213(.din(n260), .dout(n285));
  jand g0214(.dina(G68), .dinb(n153), .dout(n286));
  jor  g0215(.dina(n286), .dinb(G20), .dout(n287));
  jor  g0216(.dina(n287), .dinb(n262), .dout(n288));
  jand g0217(.dina(n288), .dinb(n141), .dout(n289));
  jand g0218(.dina(n289), .dinb(n285), .dout(n290));
  jor  g0219(.dina(n269), .dinb(n290), .dout(n291));
  jor  g0220(.dina(n291), .dinb(n284), .dout(n292));
  jand g0221(.dina(n255), .dinb(G190), .dout(n293));
  jor  g0222(.dina(n293), .dinb(n292), .dout(n294));
  jor  g0223(.dina(n294), .dinb(n283), .dout(n295));
  jand g0224(.dina(n295), .dinb(n282), .dout(n296));
  jand g0225(.dina(n168), .dinb(G257), .dout(n297));
  jand g0226(.dina(n297), .dinb(n182), .dout(n298));
  jnot g0227(.din(n298), .dout(n299));
  jor  g0228(.dina(n176), .dinb(G33), .dout(n300));
  jor  g0229(.dina(n300), .dinb(n84), .dout(n301));
  jnot g0230(.din(n152), .dout(n302));
  jor  g0231(.dina(n205), .dinb(n94), .dout(n303));
  jand g0232(.dina(n303), .dinb(n302), .dout(n304));
  jand g0233(.dina(n304), .dinb(n301), .dout(n305));
  jor  g0234(.dina(n305), .dinb(n168), .dout(n306));
  jand g0235(.dina(n306), .dinb(n229), .dout(n307));
  jand g0236(.dina(n307), .dinb(n299), .dout(n308));
  jand g0237(.dina(n308), .dinb(G190), .dout(n309));
  jor  g0238(.dina(n147), .dinb(n80), .dout(n310));
  jnot g0239(.din(n310), .dout(n311));
  jxor g0240(.dina(G107), .dinb(G97), .dout(n312));
  jand g0241(.dina(n312), .dinb(G20), .dout(n313));
  jnot g0242(.din(n313), .dout(n314));
  jand g0243(.dina(G107), .dinb(G33), .dout(n315));
  jand g0244(.dina(G77), .dinb(n153), .dout(n316));
  jor  g0245(.dina(n316), .dinb(G20), .dout(n317));
  jor  g0246(.dina(n317), .dinb(n315), .dout(n318));
  jand g0247(.dina(n318), .dinb(n141), .dout(n319));
  jand g0248(.dina(n319), .dinb(n314), .dout(n320));
  jand g0249(.dina(n144), .dinb(n80), .dout(n321));
  jor  g0250(.dina(n321), .dinb(n320), .dout(n322));
  jor  g0251(.dina(n322), .dinb(n311), .dout(n323));
  jand g0252(.dina(n173), .dinb(G250), .dout(n324));
  jand g0253(.dina(n177), .dinb(G244), .dout(n325));
  jor  g0254(.dina(n325), .dinb(n152), .dout(n326));
  jor  g0255(.dina(n326), .dinb(n324), .dout(n327));
  jand g0256(.dina(n327), .dinb(n172), .dout(n328));
  jor  g0257(.dina(n328), .dinb(n170), .dout(n329));
  jor  g0258(.dina(n329), .dinb(n298), .dout(n330));
  jand g0259(.dina(n330), .dinb(G200), .dout(n331));
  jor  g0260(.dina(n331), .dinb(n323), .dout(n332));
  jor  g0261(.dina(n332), .dinb(n309), .dout(n333));
  jor  g0262(.dina(n308), .dinb(G169), .dout(n334));
  jnot g0263(.din(n334), .dout(n335));
  jnot g0264(.din(n315), .dout(n336));
  jor  g0265(.dina(n72), .dinb(G33), .dout(n337));
  jand g0266(.dina(n337), .dinb(n151), .dout(n338));
  jand g0267(.dina(n338), .dinb(n336), .dout(n339));
  jor  g0268(.dina(n339), .dinb(n261), .dout(n340));
  jor  g0269(.dina(n340), .dinb(n313), .dout(n341));
  jnot g0270(.din(n321), .dout(n342));
  jand g0271(.dina(n342), .dinb(n341), .dout(n343));
  jand g0272(.dina(n343), .dinb(n310), .dout(n344));
  jand g0273(.dina(n308), .dinb(n189), .dout(n345));
  jor  g0274(.dina(n345), .dinb(n344), .dout(n346));
  jor  g0275(.dina(n346), .dinb(n335), .dout(n347));
  jand g0276(.dina(n347), .dinb(n333), .dout(n348));
  jand g0277(.dina(n348), .dinb(n296), .dout(n349));
  jand g0278(.dina(n349), .dinb(n242), .dout(n350));
  jand g0279(.dina(n350), .dinb(n198), .dout(n351));
  jnot g0280(.din(G45), .dout(n352));
  jand g0281(.dina(n352), .dinb(n163), .dout(n353));
  jor  g0282(.dina(n353), .dinb(G1), .dout(n354));
  jnot g0283(.din(n354), .dout(n355));
  jand g0284(.dina(n355), .dinb(n169), .dout(n356));
  jnot g0285(.din(n356), .dout(n357));
  jand g0286(.dina(n173), .dinb(G238), .dout(n358));
  jand g0287(.dina(n177), .dinb(G232), .dout(n359));
  jor  g0288(.dina(n359), .dinb(n315), .dout(n360));
  jor  g0289(.dina(n360), .dinb(n358), .dout(n361));
  jand g0290(.dina(n361), .dinb(n172), .dout(n362));
  jnot g0291(.din(n362), .dout(n363));
  jor  g0292(.dina(n355), .dinb(n94), .dout(n364));
  jor  g0293(.dina(n364), .dinb(n172), .dout(n365));
  jand g0294(.dina(n365), .dinb(n363), .dout(n366));
  jand g0295(.dina(n366), .dinb(n357), .dout(n367));
  jnot g0296(.din(n367), .dout(n368));
  jand g0297(.dina(n368), .dinb(n199), .dout(n369));
  jand g0298(.dina(G87), .dinb(G33), .dout(n370));
  jand g0299(.dina(G58), .dinb(n153), .dout(n371));
  jor  g0300(.dina(n371), .dinb(n370), .dout(n372));
  jand g0301(.dina(n372), .dinb(n151), .dout(n373));
  jand g0302(.dina(n373), .dinb(n141), .dout(n374));
  jand g0303(.dina(n139), .dinb(n151), .dout(n375));
  jnot g0304(.din(n375), .dout(n376));
  jand g0305(.dina(G20), .dinb(n142), .dout(n377));
  jnot g0306(.din(n377), .dout(n378));
  jand g0307(.dina(n378), .dinb(G77), .dout(n379));
  jand g0308(.dina(n379), .dinb(n376), .dout(n380));
  jand g0309(.dina(n144), .dinb(n72), .dout(n381));
  jor  g0310(.dina(n381), .dinb(n380), .dout(n382));
  jor  g0311(.dina(n382), .dinb(n374), .dout(n383));
  jnot g0312(.din(n383), .dout(n384));
  jand g0313(.dina(n367), .dinb(n189), .dout(n385));
  jor  g0314(.dina(n385), .dinb(n384), .dout(n386));
  jor  g0315(.dina(n386), .dinb(n369), .dout(n387));
  jnot g0316(.din(G200), .dout(n388));
  jor  g0317(.dina(n367), .dinb(n388), .dout(n389));
  jnot g0318(.din(n389), .dout(n390));
  jand g0319(.dina(n367), .dinb(G190), .dout(n391));
  jor  g0320(.dina(n391), .dinb(n383), .dout(n392));
  jor  g0321(.dina(n392), .dinb(n390), .dout(n393));
  jand g0322(.dina(n393), .dinb(n387), .dout(n394));
  jnot g0323(.din(n394), .dout(n395));
  jand g0324(.dina(n168), .dinb(G238), .dout(n396));
  jand g0325(.dina(n396), .dinb(n354), .dout(n397));
  jand g0326(.dina(n173), .dinb(G232), .dout(n398));
  jand g0327(.dina(n177), .dinb(G226), .dout(n399));
  jor  g0328(.dina(n399), .dinb(n262), .dout(n400));
  jor  g0329(.dina(n400), .dinb(n398), .dout(n401));
  jand g0330(.dina(n401), .dinb(n172), .dout(n402));
  jor  g0331(.dina(n402), .dinb(n356), .dout(n403));
  jor  g0332(.dina(n403), .dinb(n397), .dout(n404));
  jnot g0333(.din(n404), .dout(n405));
  jor  g0334(.dina(n405), .dinb(G169), .dout(n406));
  jand g0335(.dina(G77), .dinb(G33), .dout(n407));
  jand g0336(.dina(G50), .dinb(n153), .dout(n408));
  jor  g0337(.dina(n408), .dinb(n407), .dout(n409));
  jand g0338(.dina(n409), .dinb(n141), .dout(n410));
  jand g0339(.dina(n410), .dinb(n151), .dout(n411));
  jand g0340(.dina(n75), .dinb(G20), .dout(n412));
  jand g0341(.dina(n412), .dinb(n215), .dout(n413));
  jand g0342(.dina(n378), .dinb(n261), .dout(n414));
  jand g0343(.dina(n414), .dinb(G68), .dout(n415));
  jor  g0344(.dina(n415), .dinb(n413), .dout(n416));
  jor  g0345(.dina(n416), .dinb(n411), .dout(n417));
  jor  g0346(.dina(n404), .dinb(G179), .dout(n418));
  jand g0347(.dina(n418), .dinb(n417), .dout(n419));
  jand g0348(.dina(n419), .dinb(n406), .dout(n420));
  jand g0349(.dina(n405), .dinb(G190), .dout(n421));
  jand g0350(.dina(n404), .dinb(G200), .dout(n422));
  jor  g0351(.dina(n422), .dinb(n417), .dout(n423));
  jor  g0352(.dina(n423), .dinb(n421), .dout(n424));
  jnot g0353(.din(n424), .dout(n425));
  jor  g0354(.dina(n425), .dinb(n420), .dout(n426));
  jand g0355(.dina(n168), .dinb(G226), .dout(n427));
  jand g0356(.dina(n427), .dinb(n354), .dout(n428));
  jnot g0357(.din(n428), .dout(n429));
  jand g0358(.dina(n173), .dinb(G223), .dout(n430));
  jnot g0359(.din(n430), .dout(n431));
  jnot g0360(.din(n407), .dout(n432));
  jnot g0361(.din(G222), .dout(n433));
  jor  g0362(.dina(n205), .dinb(n433), .dout(n434));
  jand g0363(.dina(n434), .dinb(n432), .dout(n435));
  jand g0364(.dina(n435), .dinb(n431), .dout(n436));
  jor  g0365(.dina(n436), .dinb(n168), .dout(n437));
  jand g0366(.dina(n437), .dinb(n357), .dout(n438));
  jand g0367(.dina(n438), .dinb(n429), .dout(n439));
  jor  g0368(.dina(n439), .dinb(G169), .dout(n440));
  jand g0369(.dina(G33), .dinb(n151), .dout(n441));
  jand g0370(.dina(n441), .dinb(G58), .dout(n442));
  jnot g0371(.din(n442), .dout(n443));
  jor  g0372(.dina(n77), .dinb(n151), .dout(n444));
  jand g0373(.dina(n153), .dinb(n151), .dout(n445));
  jand g0374(.dina(n445), .dinb(G150), .dout(n446));
  jnot g0375(.din(n446), .dout(n447));
  jand g0376(.dina(n447), .dinb(n444), .dout(n448));
  jand g0377(.dina(n448), .dinb(n443), .dout(n449));
  jor  g0378(.dina(n449), .dinb(n261), .dout(n450));
  jnot g0379(.din(n450), .dout(n451));
  jnot g0380(.din(n144), .dout(n452));
  jand g0381(.dina(n452), .dinb(n73), .dout(n453));
  jnot g0382(.din(n453), .dout(n454));
  jor  g0383(.dina(n414), .dinb(n73), .dout(n455));
  jand g0384(.dina(n455), .dinb(n454), .dout(n456));
  jor  g0385(.dina(n456), .dinb(n451), .dout(n457));
  jnot g0386(.din(n435), .dout(n458));
  jor  g0387(.dina(n458), .dinb(n430), .dout(n459));
  jand g0388(.dina(n459), .dinb(n172), .dout(n460));
  jor  g0389(.dina(n460), .dinb(n356), .dout(n461));
  jor  g0390(.dina(n461), .dinb(n428), .dout(n462));
  jor  g0391(.dina(n462), .dinb(G179), .dout(n463));
  jand g0392(.dina(n463), .dinb(n457), .dout(n464));
  jand g0393(.dina(n464), .dinb(n440), .dout(n465));
  jand g0394(.dina(n439), .dinb(G190), .dout(n466));
  jnot g0395(.din(n466), .dout(n467));
  jnot g0396(.din(n456), .dout(n468));
  jand g0397(.dina(n468), .dinb(n450), .dout(n469));
  jor  g0398(.dina(n439), .dinb(n388), .dout(n470));
  jand g0399(.dina(n470), .dinb(n469), .dout(n471));
  jand g0400(.dina(n471), .dinb(n467), .dout(n472));
  jor  g0401(.dina(n472), .dinb(n465), .dout(n473));
  jand g0402(.dina(n168), .dinb(G232), .dout(n474));
  jand g0403(.dina(n474), .dinb(n354), .dout(n475));
  jand g0404(.dina(n173), .dinb(G226), .dout(n476));
  jand g0405(.dina(n177), .dinb(G223), .dout(n477));
  jor  g0406(.dina(n477), .dinb(n370), .dout(n478));
  jor  g0407(.dina(n478), .dinb(n476), .dout(n479));
  jand g0408(.dina(n479), .dinb(n172), .dout(n480));
  jor  g0409(.dina(n480), .dinb(n356), .dout(n481));
  jor  g0410(.dina(n481), .dinb(n475), .dout(n482));
  jnot g0411(.din(n482), .dout(n483));
  jor  g0412(.dina(n483), .dinb(G169), .dout(n484));
  jnot g0413(.din(G159), .dout(n485));
  jnot g0414(.din(n445), .dout(n486));
  jor  g0415(.dina(n486), .dinb(n485), .dout(n487));
  jxor g0416(.dina(G68), .dinb(G58), .dout(n488));
  jor  g0417(.dina(n488), .dinb(n151), .dout(n489));
  jand g0418(.dina(n441), .dinb(G68), .dout(n490));
  jnot g0419(.din(n490), .dout(n491));
  jand g0420(.dina(n491), .dinb(n489), .dout(n492));
  jand g0421(.dina(n492), .dinb(n487), .dout(n493));
  jor  g0422(.dina(n493), .dinb(n261), .dout(n494));
  jnot g0423(.din(n494), .dout(n495));
  jand g0424(.dina(n452), .dinb(n74), .dout(n496));
  jnot g0425(.din(n496), .dout(n497));
  jor  g0426(.dina(n414), .dinb(n74), .dout(n498));
  jand g0427(.dina(n498), .dinb(n497), .dout(n499));
  jor  g0428(.dina(n499), .dinb(n495), .dout(n500));
  jor  g0429(.dina(n482), .dinb(G179), .dout(n501));
  jand g0430(.dina(n501), .dinb(n500), .dout(n502));
  jand g0431(.dina(n502), .dinb(n484), .dout(n503));
  jor  g0432(.dina(n483), .dinb(n388), .dout(n504));
  jnot g0433(.din(n499), .dout(n505));
  jand g0434(.dina(n505), .dinb(n494), .dout(n506));
  jnot g0435(.din(G190), .dout(n507));
  jor  g0436(.dina(n482), .dinb(n507), .dout(n508));
  jand g0437(.dina(n508), .dinb(n506), .dout(n509));
  jand g0438(.dina(n509), .dinb(n504), .dout(n510));
  jor  g0439(.dina(n510), .dinb(n503), .dout(n511));
  jor  g0440(.dina(n511), .dinb(n473), .dout(n512));
  jor  g0441(.dina(n512), .dinb(n426), .dout(n513));
  jor  g0442(.dina(n513), .dinb(n395), .dout(n514));
  jnot g0443(.din(n514), .dout(n515));
  jand g0444(.dina(n515), .dinb(n351), .dout(G372));
  jnot g0445(.din(n213), .dout(n517));
  jor  g0446(.dina(n212), .dinb(G179), .dout(n518));
  jand g0447(.dina(n518), .dinb(n224), .dout(n519));
  jand g0448(.dina(n519), .dinb(n517), .dout(n520));
  jnot g0449(.din(n238), .dout(n521));
  jor  g0450(.dina(n234), .dinb(n388), .dout(n522));
  jand g0451(.dina(n522), .dinb(n225), .dout(n523));
  jand g0452(.dina(n523), .dinb(n521), .dout(n524));
  jor  g0453(.dina(n524), .dinb(n520), .dout(n525));
  jnot g0454(.din(n256), .dout(n526));
  jor  g0455(.dina(n255), .dinb(G169), .dout(n527));
  jand g0456(.dina(n527), .dinb(n292), .dout(n528));
  jand g0457(.dina(n528), .dinb(n526), .dout(n529));
  jnot g0458(.din(n283), .dout(n530));
  jor  g0459(.dina(n279), .dinb(n507), .dout(n531));
  jand g0460(.dina(n531), .dinb(n272), .dout(n532));
  jand g0461(.dina(n532), .dinb(n530), .dout(n533));
  jor  g0462(.dina(n533), .dinb(n529), .dout(n534));
  jnot g0463(.din(n309), .dout(n535));
  jor  g0464(.dina(n308), .dinb(n388), .dout(n536));
  jand g0465(.dina(n536), .dinb(n344), .dout(n537));
  jand g0466(.dina(n537), .dinb(n535), .dout(n538));
  jor  g0467(.dina(n330), .dinb(G179), .dout(n539));
  jand g0468(.dina(n539), .dinb(n323), .dout(n540));
  jand g0469(.dina(n540), .dinb(n334), .dout(n541));
  jor  g0470(.dina(n541), .dinb(n538), .dout(n542));
  jor  g0471(.dina(n542), .dinb(n534), .dout(n543));
  jor  g0472(.dina(n543), .dinb(n525), .dout(n544));
  jor  g0473(.dina(n544), .dinb(n192), .dout(n545));
  jor  g0474(.dina(n543), .dinb(n237), .dout(n546));
  jor  g0475(.dina(n347), .dinb(n533), .dout(n547));
  jand g0476(.dina(n547), .dinb(n282), .dout(n548));
  jand g0477(.dina(n548), .dinb(n546), .dout(n549));
  jand g0478(.dina(n549), .dinb(n545), .dout(n550));
  jor  g0479(.dina(n550), .dinb(n514), .dout(n551));
  jnot g0480(.din(n551), .dout(n552));
  jnot g0481(.din(n472), .dout(n553));
  jand g0482(.dina(n503), .dinb(n553), .dout(n554));
  jnot g0483(.din(n554), .dout(n555));
  jnot g0484(.din(n465), .dout(n556));
  jnot g0485(.din(n420), .dout(n557));
  jor  g0486(.dina(n425), .dinb(n387), .dout(n558));
  jand g0487(.dina(n558), .dinb(n557), .dout(n559));
  jor  g0488(.dina(n559), .dinb(n512), .dout(n560));
  jand g0489(.dina(n560), .dinb(n556), .dout(n561));
  jand g0490(.dina(n561), .dinb(n555), .dout(n562));
  jnot g0491(.din(n562), .dout(n563));
  jor  g0492(.dina(n563), .dinb(n552), .dout(G369));
  jand g0493(.dina(n143), .dinb(G213), .dout(n565));
  jand g0494(.dina(n565), .dinb(n151), .dout(n566));
  jand g0495(.dina(n566), .dinb(G343), .dout(n567));
  jor  g0496(.dina(n567), .dinb(n237), .dout(n568));
  jnot g0497(.din(n568), .dout(n569));
  jnot g0498(.din(n192), .dout(n570));
  jnot g0499(.din(n567), .dout(n571));
  jand g0500(.dina(n571), .dinb(n570), .dout(n572));
  jand g0501(.dina(n572), .dinb(n242), .dout(n573));
  jor  g0502(.dina(n573), .dinb(n569), .dout(n574));
  jand g0503(.dina(n567), .dinb(n161), .dout(n575));
  jxor g0504(.dina(n575), .dinb(n198), .dout(n576));
  jand g0505(.dina(n576), .dinb(G330), .dout(n577));
  jand g0506(.dina(n567), .dinb(n224), .dout(n578));
  jxor g0507(.dina(n578), .dinb(n242), .dout(n579));
  jand g0508(.dina(n579), .dinb(n577), .dout(n580));
  jor  g0509(.dina(n580), .dinb(n574), .dout(G399));
  jand g0510(.dina(n91), .dinb(n163), .dout(n582));
  jand g0511(.dina(n582), .dinb(n118), .dout(n583));
  jor  g0512(.dina(n567), .dinb(n550), .dout(n584));
  jnot g0513(.din(n198), .dout(n585));
  jor  g0514(.dina(n544), .dinb(n585), .dout(n586));
  jand g0515(.dina(n571), .dinb(n586), .dout(n587));
  jnot g0516(.din(n190), .dout(n588));
  jand g0517(.dina(n308), .dinb(n255), .dout(n589));
  jand g0518(.dina(n589), .dinb(n588), .dout(n590));
  jand g0519(.dina(n590), .dinb(n234), .dout(n591));
  jand g0520(.dina(n279), .dinb(n189), .dout(n592));
  jand g0521(.dina(n592), .dinb(n330), .dout(n593));
  jand g0522(.dina(n593), .dinb(n186), .dout(n594));
  jand g0523(.dina(n594), .dinb(n212), .dout(n595));
  jor  g0524(.dina(n595), .dinb(n571), .dout(n596));
  jor  g0525(.dina(n596), .dinb(n591), .dout(n597));
  jand g0526(.dina(n597), .dinb(G330), .dout(n598));
  jnot g0527(.din(n598), .dout(n599));
  jor  g0528(.dina(n599), .dinb(n587), .dout(n600));
  jand g0529(.dina(n600), .dinb(n584), .dout(n601));
  jnot g0530(.din(n601), .dout(n602));
  jand g0531(.dina(n602), .dinb(n142), .dout(n603));
  jnot g0532(.din(n582), .dout(n604));
  jand g0533(.dina(n259), .dinb(n105), .dout(n605));
  jand g0534(.dina(n605), .dinb(G1), .dout(n606));
  jand g0535(.dina(n606), .dinb(n604), .dout(n607));
  jor  g0536(.dina(n607), .dinb(n603), .dout(n608));
  jor  g0537(.dina(n608), .dinb(n583), .dout(G364));
  jand g0538(.dina(G45), .dinb(G13), .dout(n610));
  jand g0539(.dina(n610), .dinb(n151), .dout(n611));
  jor  g0540(.dina(n611), .dinb(n142), .dout(n612));
  jnot g0541(.din(n612), .dout(n613));
  jand g0542(.dina(n613), .dinb(n604), .dout(n614));
  jnot g0543(.din(n614), .dout(n615));
  jxor g0544(.dina(n576), .dinb(G330), .dout(n616));
  jand g0545(.dina(n616), .dinb(n615), .dout(n617));
  jand g0546(.dina(n153), .dinb(n89), .dout(n618));
  jand g0547(.dina(n618), .dinb(n151), .dout(n619));
  jnot g0548(.din(n619), .dout(n620));
  jor  g0549(.dina(n620), .dinb(n576), .dout(n621));
  jand g0550(.dina(n507), .dinb(G20), .dout(n622));
  jnot g0551(.din(n622), .dout(n623));
  jand g0552(.dina(G200), .dinb(G20), .dout(n624));
  jnot g0553(.din(n624), .dout(n625));
  jand g0554(.dina(G179), .dinb(G20), .dout(n626));
  jnot g0555(.din(n626), .dout(n627));
  jand g0556(.dina(n627), .dinb(n625), .dout(n628));
  jand g0557(.dina(n628), .dinb(n623), .dout(n629));
  jand g0558(.dina(n629), .dinb(G97), .dout(n630));
  jnot g0559(.din(n630), .dout(n631));
  jand g0560(.dina(n624), .dinb(n189), .dout(n632));
  jand g0561(.dina(n632), .dinb(G190), .dout(n633));
  jand g0562(.dina(n633), .dinb(G87), .dout(n634));
  jnot g0563(.din(n634), .dout(n635));
  jand g0564(.dina(n635), .dinb(n631), .dout(n636));
  jand g0565(.dina(n626), .dinb(n388), .dout(n637));
  jand g0566(.dina(n637), .dinb(n507), .dout(n638));
  jand g0567(.dina(n638), .dinb(G77), .dout(n639));
  jand g0568(.dina(n628), .dinb(n622), .dout(n640));
  jand g0569(.dina(n640), .dinb(G159), .dout(n641));
  jor  g0570(.dina(n641), .dinb(n639), .dout(n642));
  jor  g0571(.dina(n642), .dinb(G33), .dout(n643));
  jnot g0572(.din(n643), .dout(n644));
  jand g0573(.dina(n644), .dinb(n636), .dout(n645));
  jand g0574(.dina(n637), .dinb(G190), .dout(n646));
  jand g0575(.dina(n646), .dinb(G58), .dout(n647));
  jand g0576(.dina(n632), .dinb(n507), .dout(n648));
  jand g0577(.dina(n648), .dinb(G107), .dout(n649));
  jand g0578(.dina(n626), .dinb(G200), .dout(n650));
  jand g0579(.dina(n650), .dinb(G190), .dout(n651));
  jand g0580(.dina(n651), .dinb(G50), .dout(n652));
  jand g0581(.dina(n650), .dinb(n507), .dout(n653));
  jand g0582(.dina(n653), .dinb(G68), .dout(n654));
  jor  g0583(.dina(n654), .dinb(n652), .dout(n655));
  jor  g0584(.dina(n655), .dinb(n649), .dout(n656));
  jor  g0585(.dina(n656), .dinb(n647), .dout(n657));
  jnot g0586(.din(n657), .dout(n658));
  jand g0587(.dina(n658), .dinb(n645), .dout(n659));
  jnot g0588(.din(n659), .dout(n660));
  jand g0589(.dina(n646), .dinb(G322), .dout(n661));
  jand g0590(.dina(n633), .dinb(G303), .dout(n662));
  jand g0591(.dina(n629), .dinb(G294), .dout(n663));
  jor  g0592(.dina(n663), .dinb(n662), .dout(n664));
  jand g0593(.dina(n651), .dinb(G326), .dout(n665));
  jor  g0594(.dina(n665), .dinb(n664), .dout(n666));
  jand g0595(.dina(n640), .dinb(G329), .dout(n667));
  jor  g0596(.dina(n667), .dinb(n153), .dout(n668));
  jand g0597(.dina(n638), .dinb(G311), .dout(n669));
  jand g0598(.dina(n653), .dinb(G317), .dout(n670));
  jor  g0599(.dina(n670), .dinb(n669), .dout(n671));
  jand g0600(.dina(n648), .dinb(G283), .dout(n672));
  jor  g0601(.dina(n672), .dinb(n671), .dout(n673));
  jor  g0602(.dina(n673), .dinb(n668), .dout(n674));
  jor  g0603(.dina(n674), .dinb(n666), .dout(n675));
  jor  g0604(.dina(n675), .dinb(n661), .dout(n676));
  jand g0605(.dina(n676), .dinb(n660), .dout(n677));
  jand g0606(.dina(n139), .dinb(G169), .dout(n678));
  jor  g0607(.dina(n678), .dinb(n375), .dout(n679));
  jnot g0608(.din(n679), .dout(n680));
  jor  g0609(.dina(n680), .dinb(n677), .dout(n681));
  jand g0610(.dina(n680), .dinb(n620), .dout(n682));
  jor  g0611(.dina(n134), .dinb(n352), .dout(n683));
  jand g0612(.dina(n91), .dinb(G33), .dout(n684));
  jnot g0613(.din(n684), .dout(n685));
  jand g0614(.dina(n118), .dinb(n352), .dout(n686));
  jor  g0615(.dina(n686), .dinb(n685), .dout(n687));
  jnot g0616(.din(n687), .dout(n688));
  jand g0617(.dina(n688), .dinb(n683), .dout(n689));
  jnot g0618(.din(n91), .dout(n690));
  jand g0619(.dina(n690), .dinb(n105), .dout(n691));
  jand g0620(.dina(n91), .dinb(n153), .dout(n692));
  jand g0621(.dina(n692), .dinb(G355), .dout(n693));
  jor  g0622(.dina(n693), .dinb(n691), .dout(n694));
  jor  g0623(.dina(n694), .dinb(n689), .dout(n695));
  jand g0624(.dina(n695), .dinb(n682), .dout(n696));
  jnot g0625(.din(n696), .dout(n697));
  jand g0626(.dina(n697), .dinb(n681), .dout(n698));
  jand g0627(.dina(n698), .dinb(n621), .dout(n699));
  jand g0628(.dina(n699), .dinb(n614), .dout(n700));
  jor  g0629(.dina(n700), .dinb(n617), .dout(G396));
  jand g0630(.dina(n567), .dinb(n383), .dout(n702));
  jxor g0631(.dina(n702), .dinb(n394), .dout(n703));
  jnot g0632(.din(n703), .dout(n704));
  jand g0633(.dina(n704), .dinb(n618), .dout(n705));
  jnot g0634(.din(n705), .dout(n706));
  jand g0635(.dina(n653), .dinb(G150), .dout(n707));
  jand g0636(.dina(n651), .dinb(G137), .dout(n708));
  jand g0637(.dina(n633), .dinb(G50), .dout(n709));
  jor  g0638(.dina(n709), .dinb(n708), .dout(n710));
  jand g0639(.dina(n646), .dinb(G143), .dout(n711));
  jor  g0640(.dina(n711), .dinb(n710), .dout(n712));
  jor  g0641(.dina(n712), .dinb(n707), .dout(n713));
  jand g0642(.dina(n638), .dinb(G159), .dout(n714));
  jand g0643(.dina(n640), .dinb(G132), .dout(n715));
  jor  g0644(.dina(n715), .dinb(n714), .dout(n716));
  jand g0645(.dina(n629), .dinb(G58), .dout(n717));
  jand g0646(.dina(n648), .dinb(G68), .dout(n718));
  jor  g0647(.dina(n718), .dinb(n717), .dout(n719));
  jor  g0648(.dina(n719), .dinb(G33), .dout(n720));
  jor  g0649(.dina(n720), .dinb(n716), .dout(n721));
  jor  g0650(.dina(n721), .dinb(n713), .dout(n722));
  jand g0651(.dina(n653), .dinb(G283), .dout(n723));
  jand g0652(.dina(n640), .dinb(G311), .dout(n724));
  jor  g0653(.dina(n724), .dinb(n723), .dout(n725));
  jand g0654(.dina(n633), .dinb(G107), .dout(n726));
  jor  g0655(.dina(n726), .dinb(n630), .dout(n727));
  jor  g0656(.dina(n727), .dinb(n725), .dout(n728));
  jand g0657(.dina(n646), .dinb(G294), .dout(n729));
  jand g0658(.dina(n638), .dinb(G116), .dout(n730));
  jor  g0659(.dina(n730), .dinb(n729), .dout(n731));
  jand g0660(.dina(n651), .dinb(G303), .dout(n732));
  jand g0661(.dina(n648), .dinb(G87), .dout(n733));
  jor  g0662(.dina(n733), .dinb(n732), .dout(n734));
  jor  g0663(.dina(n734), .dinb(n731), .dout(n735));
  jor  g0664(.dina(n735), .dinb(n728), .dout(n736));
  jor  g0665(.dina(n736), .dinb(n153), .dout(n737));
  jand g0666(.dina(n737), .dinb(n722), .dout(n738));
  jor  g0667(.dina(n738), .dinb(n680), .dout(n739));
  jnot g0668(.din(n618), .dout(n740));
  jand g0669(.dina(n680), .dinb(n740), .dout(n741));
  jand g0670(.dina(n741), .dinb(n72), .dout(n742));
  jnot g0671(.din(n742), .dout(n743));
  jand g0672(.dina(n743), .dinb(n739), .dout(n744));
  jand g0673(.dina(n744), .dinb(n614), .dout(n745));
  jand g0674(.dina(n745), .dinb(n706), .dout(n746));
  jnot g0675(.din(n746), .dout(n747));
  jor  g0676(.dina(n584), .dinb(n395), .dout(n748));
  jand g0677(.dina(n350), .dinb(n570), .dout(n749));
  jand g0678(.dina(n349), .dinb(n520), .dout(n750));
  jnot g0679(.din(n548), .dout(n751));
  jor  g0680(.dina(n751), .dinb(n750), .dout(n752));
  jor  g0681(.dina(n752), .dinb(n749), .dout(n753));
  jand g0682(.dina(n571), .dinb(n753), .dout(n754));
  jor  g0683(.dina(n703), .dinb(n754), .dout(n755));
  jand g0684(.dina(n755), .dinb(n748), .dout(n756));
  jxor g0685(.dina(n756), .dinb(n600), .dout(n757));
  jor  g0686(.dina(n757), .dinb(n614), .dout(n758));
  jand g0687(.dina(n758), .dinb(n747), .dout(n759));
  jnot g0688(.din(n759), .dout(G384));
  jnot g0689(.din(n90), .dout(n761));
  jand g0690(.dina(n112), .dinb(n761), .dout(n762));
  jnot g0691(.din(n566), .dout(n763));
  jand g0692(.dina(n763), .dinb(n503), .dout(n764));
  jand g0693(.dina(n566), .dinb(n500), .dout(n765));
  jxor g0694(.dina(n765), .dinb(n511), .dout(n766));
  jnot g0695(.din(n766), .dout(n767));
  jor  g0696(.dina(n567), .dinb(n559), .dout(n768));
  jnot g0697(.din(n768), .dout(n769));
  jand g0698(.dina(n567), .dinb(n417), .dout(n770));
  jxor g0699(.dina(n770), .dinb(n426), .dout(n771));
  jnot g0700(.din(n771), .dout(n772));
  jand g0701(.dina(n772), .dinb(n703), .dout(n773));
  jand g0702(.dina(n773), .dinb(n754), .dout(n774));
  jor  g0703(.dina(n774), .dinb(n769), .dout(n775));
  jand g0704(.dina(n775), .dinb(n767), .dout(n776));
  jor  g0705(.dina(n776), .dinb(n764), .dout(n777));
  jand g0706(.dina(n773), .dinb(n767), .dout(n778));
  jxor g0707(.dina(n778), .dinb(n514), .dout(n779));
  jor  g0708(.dina(n779), .dinb(n600), .dout(n780));
  jor  g0709(.dina(n567), .dinb(n551), .dout(n781));
  jand g0710(.dina(n781), .dinb(n562), .dout(n782));
  jxor g0711(.dina(n782), .dinb(n780), .dout(n783));
  jxor g0712(.dina(n783), .dinb(n777), .dout(n784));
  jand g0713(.dina(n784), .dinb(n762), .dout(n785));
  jor  g0714(.dina(n75), .dinb(n74), .dout(n786));
  jand g0715(.dina(n786), .dinb(G77), .dout(n787));
  jor  g0716(.dina(n787), .dinb(n73), .dout(n788));
  jand g0717(.dina(G58), .dinb(G50), .dout(n789));
  jor  g0718(.dina(n789), .dinb(G68), .dout(n790));
  jand g0719(.dina(n790), .dinb(n90), .dout(n791));
  jand g0720(.dina(n791), .dinb(n788), .dout(n792));
  jand g0721(.dina(n312), .dinb(n120), .dout(n793));
  jand g0722(.dina(n793), .dinb(G116), .dout(n794));
  jor  g0723(.dina(n794), .dinb(n792), .dout(n795));
  jor  g0724(.dina(n795), .dinb(n785), .dout(G367));
  jand g0725(.dina(n567), .dinb(n292), .dout(n797));
  jxor g0726(.dina(n797), .dinb(n534), .dout(n798));
  jand g0727(.dina(n798), .dinb(n619), .dout(n799));
  jnot g0728(.din(n799), .dout(n800));
  jand g0729(.dina(n684), .dinb(n126), .dout(n801));
  jnot g0730(.din(n682), .dout(n802));
  jand g0731(.dina(n690), .dinb(G87), .dout(n803));
  jor  g0732(.dina(n803), .dinb(n802), .dout(n804));
  jor  g0733(.dina(n804), .dinb(n801), .dout(n805));
  jand g0734(.dina(n805), .dinb(n614), .dout(n806));
  jand g0735(.dina(n646), .dinb(G303), .dout(n807));
  jand g0736(.dina(n638), .dinb(G283), .dout(n808));
  jor  g0737(.dina(n808), .dinb(n807), .dout(n809));
  jand g0738(.dina(n651), .dinb(G311), .dout(n810));
  jand g0739(.dina(n633), .dinb(G116), .dout(n811));
  jor  g0740(.dina(n811), .dinb(n810), .dout(n812));
  jand g0741(.dina(n653), .dinb(G294), .dout(n813));
  jand g0742(.dina(n640), .dinb(G317), .dout(n814));
  jor  g0743(.dina(n814), .dinb(n813), .dout(n815));
  jand g0744(.dina(n629), .dinb(G107), .dout(n816));
  jand g0745(.dina(n648), .dinb(G97), .dout(n817));
  jor  g0746(.dina(n817), .dinb(n816), .dout(n818));
  jor  g0747(.dina(n818), .dinb(n815), .dout(n819));
  jor  g0748(.dina(n819), .dinb(n812), .dout(n820));
  jor  g0749(.dina(n820), .dinb(n809), .dout(n821));
  jand g0750(.dina(n821), .dinb(G33), .dout(n822));
  jand g0751(.dina(n638), .dinb(G50), .dout(n823));
  jand g0752(.dina(n640), .dinb(G137), .dout(n824));
  jor  g0753(.dina(n824), .dinb(n823), .dout(n825));
  jand g0754(.dina(n651), .dinb(G143), .dout(n826));
  jand g0755(.dina(n653), .dinb(G159), .dout(n827));
  jor  g0756(.dina(n827), .dinb(n826), .dout(n828));
  jand g0757(.dina(n633), .dinb(G58), .dout(n829));
  jand g0758(.dina(n629), .dinb(G68), .dout(n830));
  jor  g0759(.dina(n830), .dinb(n829), .dout(n831));
  jand g0760(.dina(n646), .dinb(G150), .dout(n832));
  jand g0761(.dina(n648), .dinb(G77), .dout(n833));
  jor  g0762(.dina(n833), .dinb(n832), .dout(n834));
  jor  g0763(.dina(n834), .dinb(n831), .dout(n835));
  jor  g0764(.dina(n835), .dinb(n828), .dout(n836));
  jor  g0765(.dina(n836), .dinb(n825), .dout(n837));
  jand g0766(.dina(n837), .dinb(n153), .dout(n838));
  jor  g0767(.dina(n838), .dinb(n822), .dout(n839));
  jor  g0768(.dina(n839), .dinb(n680), .dout(n840));
  jand g0769(.dina(n840), .dinb(n806), .dout(n841));
  jand g0770(.dina(n841), .dinb(n800), .dout(n842));
  jnot g0771(.din(n842), .dout(n843));
  jand g0772(.dina(n567), .dinb(n323), .dout(n844));
  jxor g0773(.dina(n844), .dinb(n542), .dout(n845));
  jnot g0774(.din(n845), .dout(n846));
  jand g0775(.dina(n846), .dinb(n580), .dout(n847));
  jand g0776(.dina(n571), .dinb(n541), .dout(n848));
  jand g0777(.dina(n579), .dinb(n348), .dout(n849));
  jand g0778(.dina(n849), .dinb(n572), .dout(n850));
  jand g0779(.dina(n569), .dinb(n333), .dout(n851));
  jor  g0780(.dina(n851), .dinb(n850), .dout(n852));
  jor  g0781(.dina(n852), .dinb(n848), .dout(n853));
  jxor g0782(.dina(n853), .dinb(n798), .dout(n854));
  jxor g0783(.dina(n854), .dinb(n847), .dout(n855));
  jor  g0784(.dina(n855), .dinb(n613), .dout(n856));
  jnot g0785(.din(n573), .dout(n857));
  jor  g0786(.dina(n579), .dinb(n572), .dout(n858));
  jand g0787(.dina(n858), .dinb(n857), .dout(n859));
  jxor g0788(.dina(n859), .dinb(n577), .dout(n860));
  jnot g0789(.din(n860), .dout(n861));
  jxor g0790(.dina(n580), .dinb(n574), .dout(n862));
  jxor g0791(.dina(n862), .dinb(n845), .dout(n863));
  jor  g0792(.dina(n863), .dinb(n861), .dout(n864));
  jand g0793(.dina(n864), .dinb(n601), .dout(n865));
  jor  g0794(.dina(n855), .dinb(n604), .dout(n866));
  jor  g0795(.dina(n866), .dinb(n865), .dout(n867));
  jand g0796(.dina(n867), .dinb(n856), .dout(n868));
  jand g0797(.dina(n868), .dinb(n843), .dout(n869));
  jnot g0798(.din(n869), .dout(G387));
  jor  g0799(.dina(n602), .dinb(n604), .dout(n871));
  jand g0800(.dina(n871), .dinb(n861), .dout(n872));
  jand g0801(.dina(n860), .dinb(n601), .dout(n873));
  jand g0802(.dina(n873), .dinb(n613), .dout(n874));
  jor  g0803(.dina(n874), .dinb(n614), .dout(n875));
  jor  g0804(.dina(n875), .dinb(n872), .dout(n876));
  jor  g0805(.dina(n620), .dinb(n579), .dout(n877));
  jand g0806(.dina(n653), .dinb(G58), .dout(n878));
  jand g0807(.dina(n638), .dinb(G68), .dout(n879));
  jor  g0808(.dina(n879), .dinb(n817), .dout(n880));
  jor  g0809(.dina(n880), .dinb(G33), .dout(n881));
  jor  g0810(.dina(n881), .dinb(n878), .dout(n882));
  jnot g0811(.din(n882), .dout(n883));
  jand g0812(.dina(n629), .dinb(G87), .dout(n884));
  jnot g0813(.din(n884), .dout(n885));
  jand g0814(.dina(n633), .dinb(G77), .dout(n886));
  jnot g0815(.din(n886), .dout(n887));
  jand g0816(.dina(n887), .dinb(n885), .dout(n888));
  jand g0817(.dina(n646), .dinb(G50), .dout(n889));
  jand g0818(.dina(n640), .dinb(G150), .dout(n890));
  jor  g0819(.dina(n890), .dinb(n889), .dout(n891));
  jand g0820(.dina(n651), .dinb(G159), .dout(n892));
  jor  g0821(.dina(n892), .dinb(n891), .dout(n893));
  jnot g0822(.din(n893), .dout(n894));
  jand g0823(.dina(n894), .dinb(n888), .dout(n895));
  jand g0824(.dina(n895), .dinb(n883), .dout(n896));
  jnot g0825(.din(n896), .dout(n897));
  jand g0826(.dina(n653), .dinb(G311), .dout(n898));
  jand g0827(.dina(n633), .dinb(G294), .dout(n899));
  jand g0828(.dina(n629), .dinb(G283), .dout(n900));
  jor  g0829(.dina(n900), .dinb(n899), .dout(n901));
  jand g0830(.dina(n651), .dinb(G322), .dout(n902));
  jand g0831(.dina(n640), .dinb(G326), .dout(n903));
  jor  g0832(.dina(n903), .dinb(n902), .dout(n904));
  jor  g0833(.dina(n904), .dinb(n901), .dout(n905));
  jand g0834(.dina(n638), .dinb(G303), .dout(n906));
  jand g0835(.dina(n648), .dinb(G116), .dout(n907));
  jor  g0836(.dina(n907), .dinb(n906), .dout(n908));
  jand g0837(.dina(n646), .dinb(G317), .dout(n909));
  jor  g0838(.dina(n909), .dinb(n908), .dout(n910));
  jor  g0839(.dina(n910), .dinb(n153), .dout(n911));
  jor  g0840(.dina(n911), .dinb(n905), .dout(n912));
  jor  g0841(.dina(n912), .dinb(n898), .dout(n913));
  jand g0842(.dina(n913), .dinb(n897), .dout(n914));
  jor  g0843(.dina(n914), .dinb(n680), .dout(n915));
  jand g0844(.dina(n690), .dinb(n81), .dout(n916));
  jnot g0845(.din(n916), .dout(n917));
  jnot g0846(.din(n605), .dout(n918));
  jand g0847(.dina(n692), .dinb(n918), .dout(n919));
  jnot g0848(.din(n919), .dout(n920));
  jand g0849(.dina(n130), .dinb(G45), .dout(n921));
  jor  g0850(.dina(n921), .dinb(n685), .dout(n922));
  jand g0851(.dina(n922), .dinb(n920), .dout(n923));
  jand g0852(.dina(G77), .dinb(G68), .dout(n924));
  jnot g0853(.din(n924), .dout(n925));
  jand g0854(.dina(G58), .dinb(n73), .dout(n926));
  jand g0855(.dina(n926), .dinb(n925), .dout(n927));
  jand g0856(.dina(n927), .dinb(n605), .dout(n928));
  jand g0857(.dina(n928), .dinb(n352), .dout(n929));
  jor  g0858(.dina(n929), .dinb(n923), .dout(n930));
  jand g0859(.dina(n930), .dinb(n917), .dout(n931));
  jor  g0860(.dina(n931), .dinb(n802), .dout(n932));
  jand g0861(.dina(n932), .dinb(n915), .dout(n933));
  jand g0862(.dina(n933), .dinb(n877), .dout(n934));
  jand g0863(.dina(n934), .dinb(n614), .dout(n935));
  jnot g0864(.din(n935), .dout(n936));
  jand g0865(.dina(n936), .dinb(n876), .dout(n937));
  jnot g0866(.din(n937), .dout(G393));
  jnot g0867(.din(n863), .dout(n939));
  jnot g0868(.din(n873), .dout(n940));
  jor  g0869(.dina(n940), .dinb(n939), .dout(n941));
  jor  g0870(.dina(n941), .dinb(n604), .dout(n942));
  jor  g0871(.dina(n875), .dinb(n863), .dout(n943));
  jand g0872(.dina(n845), .dinb(n619), .dout(n944));
  jnot g0873(.din(n944), .dout(n945));
  jand g0874(.dina(n690), .dinb(G97), .dout(n946));
  jand g0875(.dina(n684), .dinb(n137), .dout(n947));
  jor  g0876(.dina(n947), .dinb(n802), .dout(n948));
  jor  g0877(.dina(n948), .dinb(n946), .dout(n949));
  jand g0878(.dina(n653), .dinb(G50), .dout(n950));
  jand g0879(.dina(n638), .dinb(G58), .dout(n951));
  jor  g0880(.dina(n951), .dinb(n950), .dout(n952));
  jand g0881(.dina(n646), .dinb(G159), .dout(n953));
  jand g0882(.dina(n633), .dinb(G68), .dout(n954));
  jor  g0883(.dina(n954), .dinb(n953), .dout(n955));
  jand g0884(.dina(n651), .dinb(G150), .dout(n956));
  jor  g0885(.dina(n956), .dinb(n733), .dout(n957));
  jand g0886(.dina(n640), .dinb(G143), .dout(n958));
  jand g0887(.dina(n629), .dinb(G77), .dout(n959));
  jor  g0888(.dina(n959), .dinb(n958), .dout(n960));
  jor  g0889(.dina(n960), .dinb(n957), .dout(n961));
  jor  g0890(.dina(n961), .dinb(n955), .dout(n962));
  jor  g0891(.dina(n962), .dinb(n952), .dout(n963));
  jand g0892(.dina(n963), .dinb(n153), .dout(n964));
  jand g0893(.dina(n638), .dinb(G294), .dout(n965));
  jand g0894(.dina(n640), .dinb(G322), .dout(n966));
  jor  g0895(.dina(n966), .dinb(n965), .dout(n967));
  jand g0896(.dina(n646), .dinb(G311), .dout(n968));
  jand g0897(.dina(n651), .dinb(G317), .dout(n969));
  jor  g0898(.dina(n969), .dinb(n968), .dout(n970));
  jand g0899(.dina(n653), .dinb(G303), .dout(n971));
  jor  g0900(.dina(n971), .dinb(n649), .dout(n972));
  jor  g0901(.dina(n972), .dinb(n970), .dout(n973));
  jand g0902(.dina(n633), .dinb(G283), .dout(n974));
  jand g0903(.dina(n629), .dinb(G116), .dout(n975));
  jor  g0904(.dina(n975), .dinb(n974), .dout(n976));
  jor  g0905(.dina(n976), .dinb(n973), .dout(n977));
  jor  g0906(.dina(n977), .dinb(n967), .dout(n978));
  jand g0907(.dina(n978), .dinb(G33), .dout(n979));
  jor  g0908(.dina(n979), .dinb(n680), .dout(n980));
  jor  g0909(.dina(n980), .dinb(n964), .dout(n981));
  jand g0910(.dina(n981), .dinb(n614), .dout(n982));
  jand g0911(.dina(n982), .dinb(n949), .dout(n983));
  jand g0912(.dina(n983), .dinb(n945), .dout(n984));
  jnot g0913(.din(n984), .dout(n985));
  jand g0914(.dina(n985), .dinb(n943), .dout(n986));
  jand g0915(.dina(n986), .dinb(n942), .dout(n987));
  jnot g0916(.din(n987), .dout(G390));
  jand g0917(.dina(n766), .dinb(n618), .dout(n989));
  jnot g0918(.din(n989), .dout(n990));
  jand g0919(.dina(n651), .dinb(G128), .dout(n991));
  jand g0920(.dina(n640), .dinb(G125), .dout(n992));
  jor  g0921(.dina(n992), .dinb(n991), .dout(n993));
  jand g0922(.dina(n648), .dinb(G50), .dout(n994));
  jand g0923(.dina(n653), .dinb(G137), .dout(n995));
  jor  g0924(.dina(n995), .dinb(n994), .dout(n996));
  jor  g0925(.dina(n996), .dinb(G33), .dout(n997));
  jor  g0926(.dina(n997), .dinb(n993), .dout(n998));
  jand g0927(.dina(n638), .dinb(G143), .dout(n999));
  jand g0928(.dina(n633), .dinb(G150), .dout(n1000));
  jand g0929(.dina(n629), .dinb(G159), .dout(n1001));
  jand g0930(.dina(n646), .dinb(G132), .dout(n1002));
  jor  g0931(.dina(n1002), .dinb(n1001), .dout(n1003));
  jor  g0932(.dina(n1003), .dinb(n1000), .dout(n1004));
  jor  g0933(.dina(n1004), .dinb(n999), .dout(n1005));
  jor  g0934(.dina(n1005), .dinb(n998), .dout(n1006));
  jand g0935(.dina(n651), .dinb(G283), .dout(n1007));
  jand g0936(.dina(n638), .dinb(G97), .dout(n1008));
  jor  g0937(.dina(n1008), .dinb(n153), .dout(n1009));
  jor  g0938(.dina(n1009), .dinb(n1007), .dout(n1010));
  jand g0939(.dina(n646), .dinb(G116), .dout(n1011));
  jand g0940(.dina(n640), .dinb(G294), .dout(n1012));
  jor  g0941(.dina(n1012), .dinb(n1011), .dout(n1013));
  jand g0942(.dina(n653), .dinb(G107), .dout(n1014));
  jor  g0943(.dina(n1014), .dinb(n634), .dout(n1015));
  jor  g0944(.dina(n1015), .dinb(n1013), .dout(n1016));
  jor  g0945(.dina(n1016), .dinb(n1010), .dout(n1017));
  jor  g0946(.dina(n1017), .dinb(n959), .dout(n1018));
  jor  g0947(.dina(n1018), .dinb(n718), .dout(n1019));
  jand g0948(.dina(n1019), .dinb(n1006), .dout(n1020));
  jor  g0949(.dina(n1020), .dinb(n680), .dout(n1021));
  jand g0950(.dina(n741), .dinb(n74), .dout(n1022));
  jnot g0951(.din(n1022), .dout(n1023));
  jand g0952(.dina(n1023), .dinb(n1021), .dout(n1024));
  jand g0953(.dina(n1024), .dinb(n614), .dout(n1025));
  jand g0954(.dina(n1025), .dinb(n990), .dout(n1026));
  jnot g0955(.din(n1026), .dout(n1027));
  jor  g0956(.dina(n600), .dinb(n514), .dout(n1028));
  jand g0957(.dina(n1028), .dinb(n782), .dout(n1029));
  jnot g0958(.din(n387), .dout(n1030));
  jand g0959(.dina(n571), .dinb(n1030), .dout(n1031));
  jnot g0960(.din(n1031), .dout(n1032));
  jand g0961(.dina(n1032), .dinb(n748), .dout(n1033));
  jor  g0962(.dina(n567), .dinb(n351), .dout(n1034));
  jand g0963(.dina(n598), .dinb(n1034), .dout(n1035));
  jand g0964(.dina(n703), .dinb(n1035), .dout(n1036));
  jxor g0965(.dina(n1036), .dinb(n771), .dout(n1037));
  jxor g0966(.dina(n1037), .dinb(n1033), .dout(n1038));
  jand g0967(.dina(n1038), .dinb(n1029), .dout(n1039));
  jor  g0968(.dina(n1039), .dinb(n604), .dout(n1040));
  jand g0969(.dina(n1040), .dinb(n613), .dout(n1041));
  jor  g0970(.dina(n704), .dinb(n600), .dout(n1042));
  jor  g0971(.dina(n1042), .dinb(n771), .dout(n1043));
  jxor g0972(.dina(n775), .dinb(n767), .dout(n1044));
  jxor g0973(.dina(n1044), .dinb(n1043), .dout(n1045));
  jor  g0974(.dina(n1045), .dinb(n1041), .dout(n1046));
  jnot g0975(.din(n1039), .dout(n1047));
  jnot g0976(.din(n1043), .dout(n1048));
  jxor g0977(.dina(n1044), .dinb(n1048), .dout(n1049));
  jor  g0978(.dina(n1049), .dinb(n604), .dout(n1050));
  jor  g0979(.dina(n1050), .dinb(n1047), .dout(n1051));
  jand g0980(.dina(n1051), .dinb(n1046), .dout(n1052));
  jand g0981(.dina(n1052), .dinb(n1027), .dout(n1053));
  jnot g0982(.din(n1053), .dout(G378));
  jxor g0983(.dina(n1036), .dinb(n772), .dout(n1055));
  jxor g0984(.dina(n1055), .dinb(n1033), .dout(n1056));
  jor  g0985(.dina(n1045), .dinb(n1056), .dout(n1057));
  jand g0986(.dina(n1029), .dinb(n613), .dout(n1058));
  jand g0987(.dina(n1058), .dinb(n1057), .dout(n1059));
  jand g0988(.dina(n1048), .dinb(n767), .dout(n1060));
  jand g0989(.dina(n566), .dinb(n457), .dout(n1061));
  jxor g0990(.dina(n1061), .dinb(n473), .dout(n1062));
  jxor g0991(.dina(n1062), .dinb(n777), .dout(n1063));
  jxor g0992(.dina(n1063), .dinb(n1060), .dout(n1064));
  jor  g0993(.dina(n1064), .dinb(n1059), .dout(n1065));
  jor  g0994(.dina(n1065), .dinb(n614), .dout(n1066));
  jand g0995(.dina(n1062), .dinb(n618), .dout(n1067));
  jnot g0996(.din(n1067), .dout(n1068));
  jand g0997(.dina(G50), .dinb(G41), .dout(n1069));
  jor  g0998(.dina(n1069), .dinb(n680), .dout(n1070));
  jand g0999(.dina(n638), .dinb(G137), .dout(n1071));
  jand g1000(.dina(n633), .dinb(G143), .dout(n1072));
  jand g1001(.dina(n651), .dinb(G125), .dout(n1073));
  jor  g1002(.dina(n1073), .dinb(n1072), .dout(n1074));
  jor  g1003(.dina(n1074), .dinb(n1071), .dout(n1075));
  jand g1004(.dina(n640), .dinb(G124), .dout(n1076));
  jand g1005(.dina(n629), .dinb(G150), .dout(n1077));
  jand g1006(.dina(n646), .dinb(G128), .dout(n1078));
  jor  g1007(.dina(n1078), .dinb(n1077), .dout(n1079));
  jor  g1008(.dina(n1079), .dinb(n1076), .dout(n1080));
  jand g1009(.dina(n648), .dinb(G159), .dout(n1081));
  jand g1010(.dina(n653), .dinb(G132), .dout(n1082));
  jor  g1011(.dina(n1082), .dinb(n1081), .dout(n1083));
  jor  g1012(.dina(n1083), .dinb(G33), .dout(n1084));
  jor  g1013(.dina(n1084), .dinb(n1080), .dout(n1085));
  jor  g1014(.dina(n1085), .dinb(n1075), .dout(n1086));
  jand g1015(.dina(n653), .dinb(G97), .dout(n1087));
  jand g1016(.dina(n646), .dinb(G107), .dout(n1088));
  jor  g1017(.dina(n1088), .dinb(n1087), .dout(n1089));
  jnot g1018(.din(n1089), .dout(n1090));
  jand g1019(.dina(n648), .dinb(G58), .dout(n1091));
  jnot g1020(.din(n1091), .dout(n1092));
  jand g1021(.dina(n1092), .dinb(n887), .dout(n1093));
  jand g1022(.dina(n1093), .dinb(n1090), .dout(n1094));
  jand g1023(.dina(n640), .dinb(G283), .dout(n1095));
  jor  g1024(.dina(n1095), .dinb(n830), .dout(n1096));
  jand g1025(.dina(n651), .dinb(G116), .dout(n1097));
  jand g1026(.dina(n638), .dinb(G87), .dout(n1098));
  jor  g1027(.dina(n1098), .dinb(n1097), .dout(n1099));
  jor  g1028(.dina(n1099), .dinb(n1096), .dout(n1100));
  jnot g1029(.din(n1100), .dout(n1101));
  jand g1030(.dina(n1101), .dinb(n1094), .dout(n1102));
  jand g1031(.dina(n1102), .dinb(G33), .dout(n1103));
  jnot g1032(.din(n1103), .dout(n1104));
  jand g1033(.dina(n1104), .dinb(n1086), .dout(n1105));
  jand g1034(.dina(n1105), .dinb(n163), .dout(n1106));
  jor  g1035(.dina(n1106), .dinb(n1070), .dout(n1107));
  jand g1036(.dina(n741), .dinb(n73), .dout(n1108));
  jnot g1037(.din(n1108), .dout(n1109));
  jand g1038(.dina(n1109), .dinb(n1107), .dout(n1110));
  jand g1039(.dina(n1110), .dinb(n1068), .dout(n1111));
  jand g1040(.dina(n1111), .dinb(n614), .dout(n1112));
  jnot g1041(.din(n1112), .dout(n1113));
  jand g1042(.dina(n1113), .dinb(n1066), .dout(n1114));
  jnot g1043(.din(n1114), .dout(G375));
  jand g1044(.dina(n771), .dinb(n618), .dout(n1116));
  jnot g1045(.din(n1116), .dout(n1117));
  jand g1046(.dina(n646), .dinb(G283), .dout(n1118));
  jand g1047(.dina(n633), .dinb(G97), .dout(n1119));
  jand g1048(.dina(n653), .dinb(G116), .dout(n1120));
  jor  g1049(.dina(n1120), .dinb(n1119), .dout(n1121));
  jand g1050(.dina(n640), .dinb(G303), .dout(n1122));
  jor  g1051(.dina(n1122), .dinb(n1121), .dout(n1123));
  jor  g1052(.dina(n1123), .dinb(n1118), .dout(n1124));
  jor  g1053(.dina(n884), .dinb(n833), .dout(n1125));
  jand g1054(.dina(n651), .dinb(G294), .dout(n1126));
  jand g1055(.dina(n638), .dinb(G107), .dout(n1127));
  jor  g1056(.dina(n1127), .dinb(n1126), .dout(n1128));
  jor  g1057(.dina(n1128), .dinb(n153), .dout(n1129));
  jor  g1058(.dina(n1129), .dinb(n1125), .dout(n1130));
  jor  g1059(.dina(n1130), .dinb(n1124), .dout(n1131));
  jand g1060(.dina(n646), .dinb(G137), .dout(n1132));
  jand g1061(.dina(n633), .dinb(G159), .dout(n1133));
  jand g1062(.dina(n638), .dinb(G150), .dout(n1134));
  jor  g1063(.dina(n1134), .dinb(n1133), .dout(n1135));
  jand g1064(.dina(n651), .dinb(G132), .dout(n1136));
  jand g1065(.dina(n629), .dinb(G50), .dout(n1137));
  jor  g1066(.dina(n1137), .dinb(n1091), .dout(n1138));
  jor  g1067(.dina(n1138), .dinb(n1136), .dout(n1139));
  jand g1068(.dina(n653), .dinb(G143), .dout(n1140));
  jand g1069(.dina(n640), .dinb(G128), .dout(n1141));
  jor  g1070(.dina(n1141), .dinb(n1140), .dout(n1142));
  jor  g1071(.dina(n1142), .dinb(G33), .dout(n1143));
  jor  g1072(.dina(n1143), .dinb(n1139), .dout(n1144));
  jor  g1073(.dina(n1144), .dinb(n1135), .dout(n1145));
  jor  g1074(.dina(n1145), .dinb(n1132), .dout(n1146));
  jand g1075(.dina(n1146), .dinb(n1131), .dout(n1147));
  jor  g1076(.dina(n1147), .dinb(n680), .dout(n1148));
  jand g1077(.dina(n741), .dinb(n75), .dout(n1149));
  jnot g1078(.din(n1149), .dout(n1150));
  jand g1079(.dina(n1150), .dinb(n1148), .dout(n1151));
  jand g1080(.dina(n1151), .dinb(n1117), .dout(n1152));
  jand g1081(.dina(n1152), .dinb(n614), .dout(n1153));
  jnot g1082(.din(n1153), .dout(n1154));
  jor  g1083(.dina(n1041), .dinb(n1056), .dout(n1155));
  jnot g1084(.din(n1029), .dout(n1156));
  jor  g1085(.dina(n1040), .dinb(n1156), .dout(n1157));
  jand g1086(.dina(n1157), .dinb(n1155), .dout(n1158));
  jand g1087(.dina(n1158), .dinb(n1154), .dout(n1159));
  jnot g1088(.din(n1159), .dout(G381));
  jand g1089(.dina(n1114), .dinb(n1053), .dout(n1161));
  jand g1090(.dina(n1159), .dinb(n759), .dout(n1162));
  jand g1091(.dina(n987), .dinb(n869), .dout(n1163));
  jnot g1092(.din(G396), .dout(n1164));
  jand g1093(.dina(n937), .dinb(n1164), .dout(n1165));
  jand g1094(.dina(n1165), .dinb(n1163), .dout(n1166));
  jand g1095(.dina(n1166), .dinb(n1162), .dout(n1167));
  jand g1096(.dina(n1167), .dinb(n1161), .dout(n1168));
  jnot g1097(.din(n1168), .dout(G407));
  jnot g1098(.din(G343), .dout(n1170));
  jand g1099(.dina(n1161), .dinb(n1170), .dout(n1171));
  jnot g1100(.din(G213), .dout(n1172));
  jor  g1101(.dina(n1168), .dinb(n1172), .dout(n1173));
  jor  g1102(.dina(n1173), .dinb(n1171), .dout(G409));
  jxor g1103(.dina(n937), .dinb(n1164), .dout(n1175));
  jxor g1104(.dina(n987), .dinb(n869), .dout(n1176));
  jxor g1105(.dina(n1176), .dinb(n1175), .dout(n1177));
  jand g1106(.dina(n1170), .dinb(G213), .dout(n1178));
  jxor g1107(.dina(n1159), .dinb(G384), .dout(n1179));
  jxor g1108(.dina(n1179), .dinb(G2897), .dout(n1180));
  jand g1109(.dina(n1180), .dinb(n1178), .dout(n1181));
  jnot g1110(.din(n1178), .dout(n1182));
  jxor g1111(.dina(n1114), .dinb(n1053), .dout(n1183));
  jxor g1112(.dina(n1183), .dinb(n1179), .dout(n1184));
  jand g1113(.dina(n1184), .dinb(n1182), .dout(n1185));
  jor  g1114(.dina(n1185), .dinb(n1181), .dout(n1186));
  jxor g1115(.dina(n1186), .dinb(n1177), .dout(G405));
  jxor g1116(.dina(n1184), .dinb(n1177), .dout(G402));
endmodule


