/*

top:
	jxor: 698
	jspl: 1602
	jspl3: 1627
	jnot: 590
	jdff: 786
	jor: 1333
	jand: 2824

Summary:
	jxor: 698
	jspl: 1602
	jspl3: 1627
	jnot: 590
	jdff: 786
	jor: 1333
	jand: 2824

The maximum logic level gap of any gate:
	top: 145
*/

module gf_sin(gclk, a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, sin0, sin1, sin2, sin3, sin4, sin5, sin6, sin7, sin8, sin9, sin10, sin11, sin12, sin13, sin14, sin15, sin16, sin17, sin18, sin19, sin20, sin21, sin22, sin23, sin24);
	input gclk;
	input a0;
	input a1;
	input a2;
	input a3;
	input a4;
	input a5;
	input a6;
	input a7;
	input a8;
	input a9;
	input a10;
	input a11;
	input a12;
	input a13;
	input a14;
	input a15;
	input a16;
	input a17;
	input a18;
	input a19;
	input a20;
	input a21;
	input a22;
	input a23;
	output sin0;
	output sin1;
	output sin2;
	output sin3;
	output sin4;
	output sin5;
	output sin6;
	output sin7;
	output sin8;
	output sin9;
	output sin10;
	output sin11;
	output sin12;
	output sin13;
	output sin14;
	output sin15;
	output sin16;
	output sin17;
	output sin18;
	output sin19;
	output sin20;
	output sin21;
	output sin22;
	output sin23;
	output sin24;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1837;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire n1852;
	wire n1853;
	wire n1854;
	wire n1855;
	wire n1856;
	wire n1857;
	wire n1858;
	wire n1859;
	wire n1860;
	wire n1861;
	wire n1862;
	wire n1863;
	wire n1864;
	wire n1865;
	wire n1866;
	wire n1867;
	wire n1868;
	wire n1869;
	wire n1870;
	wire n1871;
	wire n1872;
	wire n1873;
	wire n1874;
	wire n1875;
	wire n1876;
	wire n1877;
	wire n1878;
	wire n1879;
	wire n1880;
	wire n1881;
	wire n1882;
	wire n1883;
	wire n1884;
	wire n1885;
	wire n1886;
	wire n1887;
	wire n1888;
	wire n1889;
	wire n1890;
	wire n1891;
	wire n1892;
	wire n1893;
	wire n1894;
	wire n1895;
	wire n1896;
	wire n1897;
	wire n1898;
	wire n1899;
	wire n1900;
	wire n1901;
	wire n1902;
	wire n1903;
	wire n1904;
	wire n1905;
	wire n1906;
	wire n1907;
	wire n1908;
	wire n1909;
	wire n1910;
	wire n1911;
	wire n1912;
	wire n1913;
	wire n1914;
	wire n1915;
	wire n1916;
	wire n1917;
	wire n1918;
	wire n1919;
	wire n1920;
	wire n1921;
	wire n1922;
	wire n1923;
	wire n1924;
	wire n1925;
	wire n1926;
	wire n1927;
	wire n1928;
	wire n1929;
	wire n1930;
	wire n1931;
	wire n1932;
	wire n1933;
	wire n1934;
	wire n1935;
	wire n1936;
	wire n1937;
	wire n1938;
	wire n1939;
	wire n1940;
	wire n1941;
	wire n1942;
	wire n1943;
	wire n1944;
	wire n1945;
	wire n1946;
	wire n1947;
	wire n1948;
	wire n1949;
	wire n1950;
	wire n1951;
	wire n1952;
	wire n1953;
	wire n1954;
	wire n1955;
	wire n1956;
	wire n1957;
	wire n1958;
	wire n1959;
	wire n1960;
	wire n1961;
	wire n1962;
	wire n1963;
	wire n1964;
	wire n1965;
	wire n1966;
	wire n1967;
	wire n1968;
	wire n1969;
	wire n1970;
	wire n1971;
	wire n1972;
	wire n1973;
	wire n1974;
	wire n1975;
	wire n1976;
	wire n1977;
	wire n1978;
	wire n1979;
	wire n1980;
	wire n1981;
	wire n1982;
	wire n1983;
	wire n1984;
	wire n1985;
	wire n1986;
	wire n1987;
	wire n1988;
	wire n1989;
	wire n1990;
	wire n1991;
	wire n1992;
	wire n1993;
	wire n1994;
	wire n1995;
	wire n1996;
	wire n1997;
	wire n1998;
	wire n1999;
	wire n2000;
	wire n2001;
	wire n2002;
	wire n2003;
	wire n2004;
	wire n2005;
	wire n2006;
	wire n2007;
	wire n2008;
	wire n2009;
	wire n2010;
	wire n2011;
	wire n2012;
	wire n2013;
	wire n2014;
	wire n2015;
	wire n2016;
	wire n2017;
	wire n2018;
	wire n2019;
	wire n2020;
	wire n2021;
	wire n2022;
	wire n2023;
	wire n2024;
	wire n2025;
	wire n2026;
	wire n2027;
	wire n2028;
	wire n2029;
	wire n2030;
	wire n2031;
	wire n2032;
	wire n2033;
	wire n2034;
	wire n2035;
	wire n2036;
	wire n2037;
	wire n2038;
	wire n2039;
	wire n2040;
	wire n2041;
	wire n2042;
	wire n2043;
	wire n2044;
	wire n2045;
	wire n2046;
	wire n2047;
	wire n2048;
	wire n2049;
	wire n2050;
	wire n2051;
	wire n2052;
	wire n2053;
	wire n2054;
	wire n2055;
	wire n2056;
	wire n2057;
	wire n2058;
	wire n2059;
	wire n2060;
	wire n2061;
	wire n2062;
	wire n2063;
	wire n2064;
	wire n2065;
	wire n2066;
	wire n2067;
	wire n2068;
	wire n2069;
	wire n2070;
	wire n2071;
	wire n2072;
	wire n2073;
	wire n2074;
	wire n2075;
	wire n2076;
	wire n2077;
	wire n2078;
	wire n2079;
	wire n2080;
	wire n2081;
	wire n2082;
	wire n2083;
	wire n2084;
	wire n2085;
	wire n2086;
	wire n2087;
	wire n2088;
	wire n2089;
	wire n2090;
	wire n2091;
	wire n2092;
	wire n2093;
	wire n2094;
	wire n2095;
	wire n2096;
	wire n2097;
	wire n2098;
	wire n2099;
	wire n2100;
	wire n2101;
	wire n2102;
	wire n2103;
	wire n2104;
	wire n2105;
	wire n2106;
	wire n2107;
	wire n2108;
	wire n2109;
	wire n2110;
	wire n2111;
	wire n2112;
	wire n2113;
	wire n2114;
	wire n2115;
	wire n2116;
	wire n2117;
	wire n2118;
	wire n2119;
	wire n2120;
	wire n2121;
	wire n2122;
	wire n2123;
	wire n2124;
	wire n2125;
	wire n2126;
	wire n2127;
	wire n2128;
	wire n2129;
	wire n2130;
	wire n2131;
	wire n2132;
	wire n2133;
	wire n2134;
	wire n2135;
	wire n2136;
	wire n2137;
	wire n2138;
	wire n2139;
	wire n2140;
	wire n2141;
	wire n2142;
	wire n2143;
	wire n2144;
	wire n2145;
	wire n2146;
	wire n2147;
	wire n2148;
	wire n2149;
	wire n2150;
	wire n2151;
	wire n2152;
	wire n2153;
	wire n2154;
	wire n2155;
	wire n2156;
	wire n2157;
	wire n2158;
	wire n2159;
	wire n2160;
	wire n2161;
	wire n2162;
	wire n2163;
	wire n2164;
	wire n2165;
	wire n2166;
	wire n2167;
	wire n2168;
	wire n2169;
	wire n2170;
	wire n2171;
	wire n2172;
	wire n2173;
	wire n2174;
	wire n2175;
	wire n2176;
	wire n2177;
	wire n2178;
	wire n2179;
	wire n2180;
	wire n2181;
	wire n2182;
	wire n2183;
	wire n2184;
	wire n2185;
	wire n2186;
	wire n2187;
	wire n2188;
	wire n2189;
	wire n2190;
	wire n2191;
	wire n2192;
	wire n2193;
	wire n2194;
	wire n2195;
	wire n2196;
	wire n2197;
	wire n2198;
	wire n2199;
	wire n2200;
	wire n2201;
	wire n2202;
	wire n2203;
	wire n2204;
	wire n2205;
	wire n2206;
	wire n2207;
	wire n2208;
	wire n2209;
	wire n2210;
	wire n2211;
	wire n2212;
	wire n2213;
	wire n2214;
	wire n2215;
	wire n2216;
	wire n2217;
	wire n2218;
	wire n2219;
	wire n2220;
	wire n2221;
	wire n2222;
	wire n2223;
	wire n2224;
	wire n2225;
	wire n2226;
	wire n2227;
	wire n2228;
	wire n2229;
	wire n2230;
	wire n2231;
	wire n2232;
	wire n2233;
	wire n2234;
	wire n2235;
	wire n2236;
	wire n2237;
	wire n2238;
	wire n2239;
	wire n2240;
	wire n2241;
	wire n2242;
	wire n2243;
	wire n2244;
	wire n2245;
	wire n2246;
	wire n2247;
	wire n2248;
	wire n2249;
	wire n2250;
	wire n2251;
	wire n2252;
	wire n2253;
	wire n2254;
	wire n2255;
	wire n2256;
	wire n2257;
	wire n2258;
	wire n2259;
	wire n2260;
	wire n2261;
	wire n2262;
	wire n2263;
	wire n2264;
	wire n2265;
	wire n2266;
	wire n2267;
	wire n2268;
	wire n2269;
	wire n2270;
	wire n2271;
	wire n2272;
	wire n2273;
	wire n2274;
	wire n2275;
	wire n2276;
	wire n2277;
	wire n2278;
	wire n2279;
	wire n2280;
	wire n2281;
	wire n2282;
	wire n2283;
	wire n2284;
	wire n2285;
	wire n2286;
	wire n2287;
	wire n2288;
	wire n2289;
	wire n2290;
	wire n2291;
	wire n2292;
	wire n2293;
	wire n2294;
	wire n2295;
	wire n2296;
	wire n2297;
	wire n2298;
	wire n2299;
	wire n2300;
	wire n2301;
	wire n2302;
	wire n2303;
	wire n2304;
	wire n2305;
	wire n2306;
	wire n2307;
	wire n2308;
	wire n2309;
	wire n2310;
	wire n2311;
	wire n2312;
	wire n2313;
	wire n2314;
	wire n2315;
	wire n2316;
	wire n2317;
	wire n2318;
	wire n2319;
	wire n2320;
	wire n2321;
	wire n2322;
	wire n2323;
	wire n2324;
	wire n2325;
	wire n2326;
	wire n2327;
	wire n2328;
	wire n2329;
	wire n2330;
	wire n2331;
	wire n2332;
	wire n2333;
	wire n2334;
	wire n2335;
	wire n2336;
	wire n2337;
	wire n2338;
	wire n2339;
	wire n2340;
	wire n2341;
	wire n2342;
	wire n2343;
	wire n2344;
	wire n2345;
	wire n2346;
	wire n2347;
	wire n2348;
	wire n2349;
	wire n2350;
	wire n2351;
	wire n2352;
	wire n2353;
	wire n2354;
	wire n2355;
	wire n2356;
	wire n2357;
	wire n2358;
	wire n2359;
	wire n2360;
	wire n2361;
	wire n2362;
	wire n2363;
	wire n2364;
	wire n2365;
	wire n2366;
	wire n2367;
	wire n2368;
	wire n2369;
	wire n2370;
	wire n2371;
	wire n2372;
	wire n2373;
	wire n2374;
	wire n2375;
	wire n2376;
	wire n2377;
	wire n2378;
	wire n2379;
	wire n2380;
	wire n2381;
	wire n2382;
	wire n2383;
	wire n2384;
	wire n2385;
	wire n2386;
	wire n2387;
	wire n2388;
	wire n2389;
	wire n2390;
	wire n2391;
	wire n2392;
	wire n2393;
	wire n2394;
	wire n2395;
	wire n2396;
	wire n2397;
	wire n2398;
	wire n2399;
	wire n2400;
	wire n2401;
	wire n2402;
	wire n2403;
	wire n2404;
	wire n2405;
	wire n2406;
	wire n2407;
	wire n2408;
	wire n2409;
	wire n2410;
	wire n2411;
	wire n2412;
	wire n2413;
	wire n2414;
	wire n2415;
	wire n2416;
	wire n2417;
	wire n2418;
	wire n2419;
	wire n2420;
	wire n2421;
	wire n2422;
	wire n2423;
	wire n2424;
	wire n2425;
	wire n2426;
	wire n2427;
	wire n2428;
	wire n2429;
	wire n2430;
	wire n2431;
	wire n2432;
	wire n2433;
	wire n2434;
	wire n2435;
	wire n2436;
	wire n2437;
	wire n2438;
	wire n2439;
	wire n2440;
	wire n2441;
	wire n2442;
	wire n2443;
	wire n2444;
	wire n2445;
	wire n2446;
	wire n2447;
	wire n2448;
	wire n2449;
	wire n2450;
	wire n2451;
	wire n2452;
	wire n2453;
	wire n2454;
	wire n2455;
	wire n2456;
	wire n2457;
	wire n2458;
	wire n2459;
	wire n2460;
	wire n2461;
	wire n2462;
	wire n2463;
	wire n2464;
	wire n2465;
	wire n2466;
	wire n2467;
	wire n2468;
	wire n2469;
	wire n2470;
	wire n2471;
	wire n2472;
	wire n2473;
	wire n2474;
	wire n2475;
	wire n2476;
	wire n2477;
	wire n2478;
	wire n2479;
	wire n2480;
	wire n2481;
	wire n2482;
	wire n2483;
	wire n2484;
	wire n2485;
	wire n2486;
	wire n2487;
	wire n2488;
	wire n2489;
	wire n2490;
	wire n2491;
	wire n2492;
	wire n2493;
	wire n2494;
	wire n2495;
	wire n2496;
	wire n2497;
	wire n2498;
	wire n2499;
	wire n2500;
	wire n2501;
	wire n2502;
	wire n2503;
	wire n2504;
	wire n2505;
	wire n2506;
	wire n2507;
	wire n2508;
	wire n2509;
	wire n2510;
	wire n2511;
	wire n2512;
	wire n2513;
	wire n2514;
	wire n2515;
	wire n2516;
	wire n2517;
	wire n2518;
	wire n2519;
	wire n2520;
	wire n2521;
	wire n2522;
	wire n2523;
	wire n2524;
	wire n2525;
	wire n2526;
	wire n2527;
	wire n2528;
	wire n2529;
	wire n2530;
	wire n2531;
	wire n2532;
	wire n2533;
	wire n2534;
	wire n2535;
	wire n2536;
	wire n2537;
	wire n2538;
	wire n2539;
	wire n2540;
	wire n2541;
	wire n2542;
	wire n2543;
	wire n2544;
	wire n2545;
	wire n2546;
	wire n2547;
	wire n2548;
	wire n2549;
	wire n2550;
	wire n2551;
	wire n2552;
	wire n2553;
	wire n2554;
	wire n2555;
	wire n2556;
	wire n2557;
	wire n2558;
	wire n2559;
	wire n2560;
	wire n2561;
	wire n2562;
	wire n2563;
	wire n2564;
	wire n2565;
	wire n2566;
	wire n2567;
	wire n2568;
	wire n2569;
	wire n2570;
	wire n2571;
	wire n2572;
	wire n2573;
	wire n2574;
	wire n2575;
	wire n2576;
	wire n2577;
	wire n2578;
	wire n2579;
	wire n2580;
	wire n2581;
	wire n2582;
	wire n2583;
	wire n2584;
	wire n2585;
	wire n2586;
	wire n2587;
	wire n2588;
	wire n2589;
	wire n2590;
	wire n2591;
	wire n2592;
	wire n2593;
	wire n2594;
	wire n2595;
	wire n2596;
	wire n2597;
	wire n2598;
	wire n2599;
	wire n2600;
	wire n2601;
	wire n2602;
	wire n2603;
	wire n2604;
	wire n2605;
	wire n2606;
	wire n2607;
	wire n2608;
	wire n2609;
	wire n2610;
	wire n2611;
	wire n2612;
	wire n2613;
	wire n2614;
	wire n2615;
	wire n2616;
	wire n2617;
	wire n2618;
	wire n2619;
	wire n2620;
	wire n2621;
	wire n2622;
	wire n2623;
	wire n2624;
	wire n2625;
	wire n2626;
	wire n2627;
	wire n2628;
	wire n2629;
	wire n2630;
	wire n2631;
	wire n2632;
	wire n2633;
	wire n2634;
	wire n2635;
	wire n2636;
	wire n2637;
	wire n2638;
	wire n2639;
	wire n2640;
	wire n2641;
	wire n2642;
	wire n2643;
	wire n2644;
	wire n2645;
	wire n2646;
	wire n2647;
	wire n2648;
	wire n2649;
	wire n2650;
	wire n2651;
	wire n2652;
	wire n2653;
	wire n2654;
	wire n2655;
	wire n2656;
	wire n2657;
	wire n2658;
	wire n2659;
	wire n2660;
	wire n2661;
	wire n2662;
	wire n2663;
	wire n2664;
	wire n2665;
	wire n2666;
	wire n2667;
	wire n2668;
	wire n2669;
	wire n2670;
	wire n2671;
	wire n2672;
	wire n2673;
	wire n2674;
	wire n2675;
	wire n2676;
	wire n2677;
	wire n2678;
	wire n2679;
	wire n2680;
	wire n2681;
	wire n2682;
	wire n2683;
	wire n2684;
	wire n2685;
	wire n2686;
	wire n2687;
	wire n2688;
	wire n2689;
	wire n2690;
	wire n2691;
	wire n2692;
	wire n2693;
	wire n2694;
	wire n2695;
	wire n2696;
	wire n2697;
	wire n2698;
	wire n2699;
	wire n2700;
	wire n2701;
	wire n2702;
	wire n2703;
	wire n2704;
	wire n2705;
	wire n2706;
	wire n2707;
	wire n2708;
	wire n2709;
	wire n2710;
	wire n2711;
	wire n2712;
	wire n2713;
	wire n2714;
	wire n2715;
	wire n2716;
	wire n2717;
	wire n2718;
	wire n2719;
	wire n2720;
	wire n2721;
	wire n2722;
	wire n2723;
	wire n2724;
	wire n2725;
	wire n2726;
	wire n2727;
	wire n2728;
	wire n2729;
	wire n2730;
	wire n2731;
	wire n2732;
	wire n2733;
	wire n2734;
	wire n2735;
	wire n2736;
	wire n2737;
	wire n2738;
	wire n2739;
	wire n2740;
	wire n2741;
	wire n2742;
	wire n2743;
	wire n2744;
	wire n2745;
	wire n2746;
	wire n2747;
	wire n2748;
	wire n2749;
	wire n2750;
	wire n2751;
	wire n2752;
	wire n2753;
	wire n2754;
	wire n2755;
	wire n2756;
	wire n2757;
	wire n2758;
	wire n2759;
	wire n2760;
	wire n2761;
	wire n2762;
	wire n2763;
	wire n2764;
	wire n2765;
	wire n2766;
	wire n2767;
	wire n2768;
	wire n2769;
	wire n2770;
	wire n2771;
	wire n2772;
	wire n2773;
	wire n2774;
	wire n2775;
	wire n2776;
	wire n2777;
	wire n2778;
	wire n2779;
	wire n2780;
	wire n2781;
	wire n2782;
	wire n2783;
	wire n2784;
	wire n2785;
	wire n2786;
	wire n2787;
	wire n2788;
	wire n2789;
	wire n2790;
	wire n2791;
	wire n2792;
	wire n2793;
	wire n2794;
	wire n2795;
	wire n2796;
	wire n2797;
	wire n2798;
	wire n2799;
	wire n2800;
	wire n2801;
	wire n2802;
	wire n2803;
	wire n2804;
	wire n2805;
	wire n2806;
	wire n2807;
	wire n2808;
	wire n2809;
	wire n2810;
	wire n2811;
	wire n2812;
	wire n2813;
	wire n2814;
	wire n2815;
	wire n2816;
	wire n2817;
	wire n2818;
	wire n2819;
	wire n2820;
	wire n2821;
	wire n2822;
	wire n2823;
	wire n2824;
	wire n2825;
	wire n2826;
	wire n2827;
	wire n2828;
	wire n2829;
	wire n2830;
	wire n2831;
	wire n2832;
	wire n2833;
	wire n2834;
	wire n2835;
	wire n2836;
	wire n2837;
	wire n2838;
	wire n2839;
	wire n2840;
	wire n2841;
	wire n2842;
	wire n2843;
	wire n2844;
	wire n2845;
	wire n2846;
	wire n2847;
	wire n2848;
	wire n2849;
	wire n2850;
	wire n2851;
	wire n2852;
	wire n2853;
	wire n2854;
	wire n2855;
	wire n2856;
	wire n2857;
	wire n2858;
	wire n2859;
	wire n2860;
	wire n2861;
	wire n2862;
	wire n2863;
	wire n2864;
	wire n2865;
	wire n2866;
	wire n2867;
	wire n2868;
	wire n2869;
	wire n2870;
	wire n2871;
	wire n2872;
	wire n2873;
	wire n2874;
	wire n2875;
	wire n2876;
	wire n2877;
	wire n2878;
	wire n2879;
	wire n2880;
	wire n2881;
	wire n2882;
	wire n2883;
	wire n2884;
	wire n2885;
	wire n2886;
	wire n2887;
	wire n2888;
	wire n2889;
	wire n2890;
	wire n2891;
	wire n2892;
	wire n2893;
	wire n2894;
	wire n2895;
	wire n2896;
	wire n2897;
	wire n2898;
	wire n2899;
	wire n2900;
	wire n2901;
	wire n2902;
	wire n2903;
	wire n2904;
	wire n2905;
	wire n2906;
	wire n2907;
	wire n2908;
	wire n2909;
	wire n2910;
	wire n2911;
	wire n2912;
	wire n2913;
	wire n2914;
	wire n2915;
	wire n2916;
	wire n2917;
	wire n2918;
	wire n2919;
	wire n2920;
	wire n2921;
	wire n2922;
	wire n2923;
	wire n2924;
	wire n2925;
	wire n2926;
	wire n2927;
	wire n2928;
	wire n2929;
	wire n2930;
	wire n2931;
	wire n2932;
	wire n2933;
	wire n2934;
	wire n2935;
	wire n2936;
	wire n2937;
	wire n2938;
	wire n2939;
	wire n2940;
	wire n2941;
	wire n2942;
	wire n2943;
	wire n2944;
	wire n2945;
	wire n2946;
	wire n2947;
	wire n2948;
	wire n2949;
	wire n2950;
	wire n2951;
	wire n2952;
	wire n2953;
	wire n2954;
	wire n2955;
	wire n2956;
	wire n2957;
	wire n2958;
	wire n2959;
	wire n2960;
	wire n2961;
	wire n2962;
	wire n2963;
	wire n2964;
	wire n2965;
	wire n2966;
	wire n2967;
	wire n2968;
	wire n2969;
	wire n2970;
	wire n2971;
	wire n2972;
	wire n2973;
	wire n2974;
	wire n2975;
	wire n2976;
	wire n2977;
	wire n2978;
	wire n2979;
	wire n2980;
	wire n2981;
	wire n2982;
	wire n2983;
	wire n2984;
	wire n2985;
	wire n2986;
	wire n2987;
	wire n2988;
	wire n2989;
	wire n2990;
	wire n2991;
	wire n2992;
	wire n2993;
	wire n2994;
	wire n2995;
	wire n2996;
	wire n2997;
	wire n2998;
	wire n2999;
	wire n3000;
	wire n3001;
	wire n3002;
	wire n3003;
	wire n3004;
	wire n3005;
	wire n3006;
	wire n3007;
	wire n3008;
	wire n3009;
	wire n3010;
	wire n3011;
	wire n3012;
	wire n3013;
	wire n3014;
	wire n3015;
	wire n3016;
	wire n3017;
	wire n3018;
	wire n3019;
	wire n3020;
	wire n3021;
	wire n3022;
	wire n3023;
	wire n3024;
	wire n3025;
	wire n3026;
	wire n3027;
	wire n3028;
	wire n3029;
	wire n3030;
	wire n3031;
	wire n3032;
	wire n3033;
	wire n3034;
	wire n3035;
	wire n3036;
	wire n3037;
	wire n3038;
	wire n3039;
	wire n3040;
	wire n3041;
	wire n3042;
	wire n3043;
	wire n3044;
	wire n3045;
	wire n3046;
	wire n3047;
	wire n3048;
	wire n3049;
	wire n3050;
	wire n3051;
	wire n3052;
	wire n3053;
	wire n3054;
	wire n3055;
	wire n3056;
	wire n3057;
	wire n3058;
	wire n3059;
	wire n3060;
	wire n3061;
	wire n3062;
	wire n3063;
	wire n3064;
	wire n3065;
	wire n3066;
	wire n3067;
	wire n3068;
	wire n3069;
	wire n3070;
	wire n3071;
	wire n3072;
	wire n3073;
	wire n3074;
	wire n3075;
	wire n3076;
	wire n3077;
	wire n3078;
	wire n3079;
	wire n3080;
	wire n3081;
	wire n3082;
	wire n3083;
	wire n3084;
	wire n3085;
	wire n3086;
	wire n3087;
	wire n3088;
	wire n3089;
	wire n3090;
	wire n3091;
	wire n3092;
	wire n3093;
	wire n3094;
	wire n3095;
	wire n3096;
	wire n3097;
	wire n3098;
	wire n3099;
	wire n3100;
	wire n3101;
	wire n3102;
	wire n3103;
	wire n3104;
	wire n3105;
	wire n3106;
	wire n3107;
	wire n3108;
	wire n3109;
	wire n3110;
	wire n3111;
	wire n3112;
	wire n3113;
	wire n3114;
	wire n3115;
	wire n3116;
	wire n3117;
	wire n3118;
	wire n3119;
	wire n3120;
	wire n3121;
	wire n3122;
	wire n3123;
	wire n3124;
	wire n3125;
	wire n3126;
	wire n3128;
	wire n3129;
	wire n3130;
	wire n3131;
	wire n3132;
	wire n3133;
	wire n3134;
	wire n3135;
	wire n3136;
	wire n3137;
	wire n3138;
	wire n3139;
	wire n3140;
	wire n3141;
	wire n3142;
	wire n3143;
	wire n3144;
	wire n3145;
	wire n3146;
	wire n3147;
	wire n3148;
	wire n3149;
	wire n3150;
	wire n3151;
	wire n3152;
	wire n3153;
	wire n3154;
	wire n3155;
	wire n3156;
	wire n3157;
	wire n3158;
	wire n3159;
	wire n3160;
	wire n3161;
	wire n3162;
	wire n3163;
	wire n3164;
	wire n3165;
	wire n3166;
	wire n3167;
	wire n3168;
	wire n3169;
	wire n3170;
	wire n3171;
	wire n3172;
	wire n3173;
	wire n3174;
	wire n3175;
	wire n3176;
	wire n3177;
	wire n3178;
	wire n3179;
	wire n3180;
	wire n3181;
	wire n3182;
	wire n3183;
	wire n3184;
	wire n3185;
	wire n3186;
	wire n3187;
	wire n3188;
	wire n3189;
	wire n3190;
	wire n3191;
	wire n3192;
	wire n3193;
	wire n3194;
	wire n3195;
	wire n3196;
	wire n3197;
	wire n3198;
	wire n3199;
	wire n3200;
	wire n3201;
	wire n3202;
	wire n3203;
	wire n3204;
	wire n3205;
	wire n3206;
	wire n3207;
	wire n3208;
	wire n3209;
	wire n3210;
	wire n3211;
	wire n3212;
	wire n3213;
	wire n3214;
	wire n3215;
	wire n3216;
	wire n3217;
	wire n3218;
	wire n3219;
	wire n3220;
	wire n3221;
	wire n3222;
	wire n3223;
	wire n3224;
	wire n3225;
	wire n3226;
	wire n3227;
	wire n3228;
	wire n3229;
	wire n3230;
	wire n3231;
	wire n3232;
	wire n3233;
	wire n3234;
	wire n3235;
	wire n3236;
	wire n3237;
	wire n3238;
	wire n3239;
	wire n3240;
	wire n3241;
	wire n3242;
	wire n3243;
	wire n3244;
	wire n3245;
	wire n3246;
	wire n3247;
	wire n3248;
	wire n3249;
	wire n3250;
	wire n3251;
	wire n3252;
	wire n3253;
	wire n3254;
	wire n3255;
	wire n3256;
	wire n3257;
	wire n3258;
	wire n3259;
	wire n3260;
	wire n3261;
	wire n3262;
	wire n3263;
	wire n3264;
	wire n3265;
	wire n3266;
	wire n3267;
	wire n3268;
	wire n3269;
	wire n3270;
	wire n3271;
	wire n3272;
	wire n3273;
	wire n3274;
	wire n3275;
	wire n3276;
	wire n3277;
	wire n3278;
	wire n3279;
	wire n3280;
	wire n3281;
	wire n3282;
	wire n3283;
	wire n3284;
	wire n3285;
	wire n3286;
	wire n3287;
	wire n3288;
	wire n3289;
	wire n3290;
	wire n3291;
	wire n3292;
	wire n3293;
	wire n3294;
	wire n3295;
	wire n3296;
	wire n3297;
	wire n3298;
	wire n3299;
	wire n3300;
	wire n3301;
	wire n3302;
	wire n3303;
	wire n3304;
	wire n3305;
	wire n3306;
	wire n3307;
	wire n3308;
	wire n3309;
	wire n3310;
	wire n3311;
	wire n3312;
	wire n3313;
	wire n3314;
	wire n3315;
	wire n3316;
	wire n3317;
	wire n3318;
	wire n3319;
	wire n3320;
	wire n3321;
	wire n3322;
	wire n3323;
	wire n3324;
	wire n3325;
	wire n3326;
	wire n3327;
	wire n3328;
	wire n3329;
	wire n3330;
	wire n3331;
	wire n3332;
	wire n3333;
	wire n3334;
	wire n3335;
	wire n3336;
	wire n3337;
	wire n3338;
	wire n3339;
	wire n3340;
	wire n3341;
	wire n3342;
	wire n3343;
	wire n3344;
	wire n3345;
	wire n3346;
	wire n3347;
	wire n3348;
	wire n3349;
	wire n3350;
	wire n3351;
	wire n3352;
	wire n3353;
	wire n3354;
	wire n3355;
	wire n3356;
	wire n3357;
	wire n3358;
	wire n3359;
	wire n3360;
	wire n3361;
	wire n3362;
	wire n3363;
	wire n3364;
	wire n3365;
	wire n3366;
	wire n3367;
	wire n3368;
	wire n3369;
	wire n3370;
	wire n3371;
	wire n3372;
	wire n3373;
	wire n3374;
	wire n3375;
	wire n3376;
	wire n3377;
	wire n3378;
	wire n3379;
	wire n3380;
	wire n3381;
	wire n3382;
	wire n3383;
	wire n3384;
	wire n3385;
	wire n3386;
	wire n3387;
	wire n3388;
	wire n3389;
	wire n3390;
	wire n3391;
	wire n3392;
	wire n3393;
	wire n3394;
	wire n3395;
	wire n3396;
	wire n3397;
	wire n3398;
	wire n3399;
	wire n3400;
	wire n3401;
	wire n3402;
	wire n3403;
	wire n3404;
	wire n3405;
	wire n3406;
	wire n3407;
	wire n3408;
	wire n3409;
	wire n3410;
	wire n3411;
	wire n3412;
	wire n3413;
	wire n3414;
	wire n3415;
	wire n3416;
	wire n3417;
	wire n3418;
	wire n3419;
	wire n3420;
	wire n3421;
	wire n3422;
	wire n3423;
	wire n3424;
	wire n3425;
	wire n3426;
	wire n3427;
	wire n3428;
	wire n3429;
	wire n3430;
	wire n3431;
	wire n3432;
	wire n3433;
	wire n3434;
	wire n3435;
	wire n3436;
	wire n3437;
	wire n3438;
	wire n3439;
	wire n3440;
	wire n3441;
	wire n3442;
	wire n3443;
	wire n3444;
	wire n3445;
	wire n3446;
	wire n3447;
	wire n3448;
	wire n3449;
	wire n3450;
	wire n3451;
	wire n3452;
	wire n3453;
	wire n3454;
	wire n3455;
	wire n3456;
	wire n3457;
	wire n3458;
	wire n3459;
	wire n3460;
	wire n3461;
	wire n3462;
	wire n3463;
	wire n3464;
	wire n3465;
	wire n3466;
	wire n3467;
	wire n3468;
	wire n3469;
	wire n3470;
	wire n3471;
	wire n3472;
	wire n3473;
	wire n3474;
	wire n3475;
	wire n3476;
	wire n3477;
	wire n3478;
	wire n3479;
	wire n3480;
	wire n3481;
	wire n3482;
	wire n3483;
	wire n3484;
	wire n3485;
	wire n3486;
	wire n3487;
	wire n3488;
	wire n3489;
	wire n3490;
	wire n3491;
	wire n3492;
	wire n3493;
	wire n3494;
	wire n3495;
	wire n3496;
	wire n3497;
	wire n3498;
	wire n3499;
	wire n3500;
	wire n3501;
	wire n3502;
	wire n3503;
	wire n3504;
	wire n3505;
	wire n3506;
	wire n3507;
	wire n3508;
	wire n3509;
	wire n3510;
	wire n3511;
	wire n3512;
	wire n3513;
	wire n3514;
	wire n3515;
	wire n3516;
	wire n3517;
	wire n3518;
	wire n3519;
	wire n3520;
	wire n3521;
	wire n3522;
	wire n3523;
	wire n3524;
	wire n3525;
	wire n3526;
	wire n3527;
	wire n3528;
	wire n3529;
	wire n3530;
	wire n3531;
	wire n3532;
	wire n3533;
	wire n3534;
	wire n3535;
	wire n3536;
	wire n3537;
	wire n3538;
	wire n3539;
	wire n3540;
	wire n3541;
	wire n3542;
	wire n3543;
	wire n3544;
	wire n3545;
	wire n3546;
	wire n3547;
	wire n3548;
	wire n3549;
	wire n3550;
	wire n3551;
	wire n3552;
	wire n3553;
	wire n3554;
	wire n3555;
	wire n3556;
	wire n3557;
	wire n3558;
	wire n3559;
	wire n3560;
	wire n3561;
	wire n3562;
	wire n3563;
	wire n3564;
	wire n3565;
	wire n3566;
	wire n3567;
	wire n3568;
	wire n3569;
	wire n3570;
	wire n3571;
	wire n3572;
	wire n3573;
	wire n3574;
	wire n3575;
	wire n3576;
	wire n3577;
	wire n3578;
	wire n3579;
	wire n3580;
	wire n3581;
	wire n3582;
	wire n3583;
	wire n3584;
	wire n3585;
	wire n3586;
	wire n3587;
	wire n3588;
	wire n3589;
	wire n3590;
	wire n3591;
	wire n3592;
	wire n3593;
	wire n3594;
	wire n3595;
	wire n3596;
	wire n3597;
	wire n3598;
	wire n3599;
	wire n3600;
	wire n3601;
	wire n3602;
	wire n3603;
	wire n3604;
	wire n3605;
	wire n3606;
	wire n3607;
	wire n3608;
	wire n3609;
	wire n3610;
	wire n3611;
	wire n3612;
	wire n3613;
	wire n3614;
	wire n3615;
	wire n3616;
	wire n3617;
	wire n3618;
	wire n3619;
	wire n3620;
	wire n3621;
	wire n3622;
	wire n3623;
	wire n3624;
	wire n3625;
	wire n3626;
	wire n3627;
	wire n3628;
	wire n3629;
	wire n3630;
	wire n3631;
	wire n3632;
	wire n3633;
	wire n3634;
	wire n3635;
	wire n3636;
	wire n3637;
	wire n3638;
	wire n3639;
	wire n3640;
	wire n3641;
	wire n3642;
	wire n3643;
	wire n3644;
	wire n3645;
	wire n3646;
	wire n3647;
	wire n3648;
	wire n3649;
	wire n3650;
	wire n3651;
	wire n3652;
	wire n3653;
	wire n3654;
	wire n3655;
	wire n3656;
	wire n3657;
	wire n3658;
	wire n3659;
	wire n3660;
	wire n3661;
	wire n3662;
	wire n3663;
	wire n3664;
	wire n3665;
	wire n3666;
	wire n3667;
	wire n3668;
	wire n3669;
	wire n3670;
	wire n3671;
	wire n3672;
	wire n3673;
	wire n3674;
	wire n3675;
	wire n3676;
	wire n3677;
	wire n3678;
	wire n3679;
	wire n3680;
	wire n3681;
	wire n3682;
	wire n3683;
	wire n3684;
	wire n3685;
	wire n3686;
	wire n3687;
	wire n3688;
	wire n3689;
	wire n3690;
	wire n3691;
	wire n3692;
	wire n3693;
	wire n3694;
	wire n3695;
	wire n3696;
	wire n3697;
	wire n3698;
	wire n3699;
	wire n3700;
	wire n3701;
	wire n3702;
	wire n3703;
	wire n3704;
	wire n3705;
	wire n3706;
	wire n3707;
	wire n3708;
	wire n3709;
	wire n3710;
	wire n3711;
	wire n3712;
	wire n3713;
	wire n3714;
	wire n3715;
	wire n3716;
	wire n3717;
	wire n3718;
	wire n3719;
	wire n3720;
	wire n3721;
	wire n3722;
	wire n3723;
	wire n3724;
	wire n3725;
	wire n3726;
	wire n3727;
	wire n3728;
	wire n3729;
	wire n3730;
	wire n3731;
	wire n3732;
	wire n3733;
	wire n3734;
	wire n3735;
	wire n3736;
	wire n3737;
	wire n3738;
	wire n3739;
	wire n3740;
	wire n3741;
	wire n3742;
	wire n3743;
	wire n3744;
	wire n3745;
	wire n3746;
	wire n3747;
	wire n3748;
	wire n3749;
	wire n3750;
	wire n3751;
	wire n3752;
	wire n3753;
	wire n3754;
	wire n3755;
	wire n3756;
	wire n3757;
	wire n3758;
	wire n3759;
	wire n3760;
	wire n3761;
	wire n3762;
	wire n3763;
	wire n3764;
	wire n3765;
	wire n3766;
	wire n3767;
	wire n3768;
	wire n3769;
	wire n3770;
	wire n3771;
	wire n3772;
	wire n3773;
	wire n3774;
	wire n3775;
	wire n3779;
	wire n3780;
	wire n3781;
	wire n3782;
	wire n3783;
	wire n3784;
	wire n3785;
	wire n3786;
	wire n3787;
	wire n3788;
	wire n3789;
	wire n3790;
	wire n3791;
	wire n3792;
	wire n3793;
	wire n3794;
	wire n3795;
	wire n3796;
	wire n3797;
	wire n3798;
	wire n3799;
	wire n3800;
	wire n3801;
	wire n3802;
	wire n3803;
	wire n3804;
	wire n3805;
	wire n3806;
	wire n3807;
	wire n3808;
	wire n3809;
	wire n3810;
	wire n3811;
	wire n3812;
	wire n3813;
	wire n3814;
	wire n3815;
	wire n3816;
	wire n3817;
	wire n3818;
	wire n3819;
	wire n3820;
	wire n3821;
	wire n3822;
	wire n3823;
	wire n3824;
	wire n3825;
	wire n3826;
	wire n3827;
	wire n3828;
	wire n3829;
	wire n3830;
	wire n3831;
	wire n3832;
	wire n3833;
	wire n3834;
	wire n3835;
	wire n3836;
	wire n3837;
	wire n3838;
	wire n3839;
	wire n3840;
	wire n3841;
	wire n3842;
	wire n3843;
	wire n3844;
	wire n3845;
	wire n3846;
	wire n3847;
	wire n3848;
	wire n3849;
	wire n3850;
	wire n3851;
	wire n3852;
	wire n3853;
	wire n3854;
	wire n3855;
	wire n3856;
	wire n3857;
	wire n3858;
	wire n3859;
	wire n3860;
	wire n3861;
	wire n3862;
	wire n3863;
	wire n3864;
	wire n3865;
	wire n3866;
	wire n3867;
	wire n3868;
	wire n3869;
	wire n3870;
	wire n3871;
	wire n3872;
	wire n3873;
	wire n3874;
	wire n3875;
	wire n3876;
	wire n3877;
	wire n3878;
	wire n3879;
	wire n3880;
	wire n3881;
	wire n3882;
	wire n3883;
	wire n3884;
	wire n3885;
	wire n3886;
	wire n3887;
	wire n3888;
	wire n3889;
	wire n3890;
	wire n3891;
	wire n3892;
	wire n3893;
	wire n3894;
	wire n3895;
	wire n3896;
	wire n3897;
	wire n3898;
	wire n3899;
	wire n3900;
	wire n3901;
	wire n3902;
	wire n3903;
	wire n3904;
	wire n3905;
	wire n3906;
	wire n3907;
	wire n3908;
	wire n3909;
	wire n3910;
	wire n3911;
	wire n3912;
	wire n3913;
	wire n3914;
	wire n3915;
	wire n3916;
	wire n3917;
	wire n3918;
	wire n3919;
	wire n3920;
	wire n3921;
	wire n3922;
	wire n3923;
	wire n3924;
	wire n3925;
	wire n3926;
	wire n3927;
	wire n3928;
	wire n3929;
	wire n3930;
	wire n3931;
	wire n3932;
	wire n3933;
	wire n3934;
	wire n3935;
	wire n3936;
	wire n3937;
	wire n3938;
	wire n3939;
	wire n3940;
	wire n3941;
	wire n3942;
	wire n3943;
	wire n3944;
	wire n3945;
	wire n3946;
	wire n3947;
	wire n3948;
	wire n3949;
	wire n3950;
	wire n3951;
	wire n3952;
	wire n3953;
	wire n3954;
	wire n3955;
	wire n3956;
	wire n3957;
	wire n3958;
	wire n3959;
	wire n3960;
	wire n3961;
	wire n3962;
	wire n3963;
	wire n3964;
	wire n3965;
	wire n3966;
	wire n3967;
	wire n3968;
	wire n3969;
	wire n3970;
	wire n3971;
	wire n3972;
	wire n3973;
	wire n3974;
	wire n3975;
	wire n3976;
	wire n3977;
	wire n3978;
	wire n3979;
	wire n3980;
	wire n3981;
	wire n3982;
	wire n3983;
	wire n3984;
	wire n3985;
	wire n3986;
	wire n3987;
	wire n3988;
	wire n3989;
	wire n3990;
	wire n3991;
	wire n3992;
	wire n3993;
	wire n3994;
	wire n3995;
	wire n3996;
	wire n3997;
	wire n3998;
	wire n3999;
	wire n4000;
	wire n4001;
	wire n4002;
	wire n4003;
	wire n4004;
	wire n4005;
	wire n4006;
	wire n4007;
	wire n4008;
	wire n4009;
	wire n4010;
	wire n4011;
	wire n4012;
	wire n4013;
	wire n4014;
	wire n4015;
	wire n4016;
	wire n4017;
	wire n4018;
	wire n4019;
	wire n4020;
	wire n4021;
	wire n4022;
	wire n4023;
	wire n4024;
	wire n4025;
	wire n4026;
	wire n4027;
	wire n4028;
	wire n4029;
	wire n4030;
	wire n4031;
	wire n4032;
	wire n4033;
	wire n4034;
	wire n4035;
	wire n4036;
	wire n4037;
	wire n4038;
	wire n4039;
	wire n4040;
	wire n4041;
	wire n4042;
	wire n4043;
	wire n4044;
	wire n4045;
	wire n4046;
	wire n4047;
	wire n4048;
	wire n4049;
	wire n4050;
	wire n4051;
	wire n4052;
	wire n4053;
	wire n4054;
	wire n4055;
	wire n4056;
	wire n4057;
	wire n4058;
	wire n4059;
	wire n4060;
	wire n4061;
	wire n4062;
	wire n4063;
	wire n4064;
	wire n4065;
	wire n4066;
	wire n4067;
	wire n4068;
	wire n4069;
	wire n4070;
	wire n4071;
	wire n4072;
	wire n4073;
	wire n4074;
	wire n4075;
	wire n4076;
	wire n4077;
	wire n4078;
	wire n4079;
	wire n4080;
	wire n4081;
	wire n4082;
	wire n4083;
	wire n4084;
	wire n4085;
	wire n4086;
	wire n4087;
	wire n4088;
	wire n4089;
	wire n4090;
	wire n4091;
	wire n4093;
	wire n4094;
	wire n4095;
	wire n4096;
	wire n4097;
	wire n4098;
	wire n4099;
	wire n4100;
	wire n4101;
	wire n4102;
	wire n4103;
	wire n4104;
	wire n4105;
	wire n4106;
	wire n4107;
	wire n4108;
	wire n4109;
	wire n4110;
	wire n4111;
	wire n4112;
	wire n4113;
	wire n4114;
	wire n4115;
	wire n4116;
	wire n4117;
	wire n4118;
	wire n4119;
	wire n4120;
	wire n4121;
	wire n4122;
	wire n4123;
	wire n4124;
	wire n4125;
	wire n4126;
	wire n4127;
	wire n4128;
	wire n4129;
	wire n4130;
	wire n4131;
	wire n4132;
	wire n4133;
	wire n4134;
	wire n4135;
	wire n4136;
	wire n4137;
	wire n4138;
	wire n4139;
	wire n4140;
	wire n4141;
	wire n4142;
	wire n4143;
	wire n4144;
	wire n4145;
	wire n4146;
	wire n4147;
	wire n4148;
	wire n4149;
	wire n4150;
	wire n4151;
	wire n4152;
	wire n4153;
	wire n4154;
	wire n4155;
	wire n4156;
	wire n4157;
	wire n4158;
	wire n4159;
	wire n4160;
	wire n4161;
	wire n4162;
	wire n4163;
	wire n4164;
	wire n4165;
	wire n4166;
	wire n4167;
	wire n4168;
	wire n4169;
	wire n4170;
	wire n4171;
	wire n4172;
	wire n4173;
	wire n4174;
	wire n4175;
	wire n4176;
	wire n4177;
	wire n4178;
	wire n4179;
	wire n4180;
	wire n4181;
	wire n4182;
	wire n4183;
	wire n4184;
	wire n4185;
	wire n4186;
	wire n4187;
	wire n4188;
	wire n4189;
	wire n4190;
	wire n4191;
	wire n4192;
	wire n4193;
	wire n4194;
	wire n4195;
	wire n4196;
	wire n4197;
	wire n4198;
	wire n4199;
	wire n4200;
	wire n4201;
	wire n4202;
	wire n4203;
	wire n4204;
	wire n4205;
	wire n4206;
	wire n4207;
	wire n4208;
	wire n4209;
	wire n4210;
	wire n4211;
	wire n4212;
	wire n4213;
	wire n4214;
	wire n4215;
	wire n4216;
	wire n4219;
	wire n4220;
	wire n4221;
	wire n4222;
	wire n4223;
	wire n4224;
	wire n4225;
	wire n4226;
	wire n4227;
	wire n4228;
	wire n4229;
	wire n4230;
	wire n4231;
	wire n4232;
	wire n4233;
	wire n4234;
	wire n4235;
	wire n4236;
	wire n4237;
	wire n4238;
	wire n4239;
	wire n4240;
	wire n4241;
	wire n4242;
	wire n4243;
	wire n4244;
	wire n4245;
	wire n4246;
	wire n4247;
	wire n4248;
	wire n4250;
	wire n4251;
	wire n4252;
	wire n4253;
	wire n4254;
	wire n4255;
	wire n4256;
	wire n4257;
	wire n4258;
	wire n4259;
	wire n4260;
	wire n4261;
	wire n4262;
	wire n4263;
	wire n4264;
	wire n4265;
	wire n4266;
	wire n4267;
	wire n4268;
	wire n4269;
	wire n4270;
	wire n4271;
	wire n4272;
	wire n4273;
	wire n4274;
	wire n4275;
	wire n4276;
	wire n4277;
	wire n4278;
	wire n4279;
	wire n4280;
	wire n4281;
	wire n4282;
	wire n4283;
	wire n4284;
	wire n4285;
	wire n4286;
	wire n4287;
	wire n4288;
	wire n4289;
	wire n4290;
	wire n4291;
	wire n4292;
	wire n4293;
	wire n4294;
	wire n4295;
	wire n4296;
	wire n4297;
	wire n4298;
	wire n4299;
	wire n4300;
	wire n4301;
	wire n4302;
	wire n4303;
	wire n4304;
	wire n4305;
	wire n4306;
	wire n4307;
	wire n4308;
	wire n4309;
	wire n4310;
	wire n4311;
	wire n4312;
	wire n4313;
	wire n4314;
	wire n4315;
	wire n4316;
	wire n4317;
	wire n4318;
	wire n4319;
	wire n4320;
	wire n4321;
	wire n4322;
	wire n4323;
	wire n4324;
	wire n4325;
	wire n4326;
	wire n4327;
	wire n4328;
	wire n4329;
	wire n4330;
	wire n4331;
	wire n4332;
	wire n4333;
	wire n4334;
	wire n4335;
	wire n4336;
	wire n4337;
	wire n4338;
	wire n4339;
	wire n4340;
	wire n4341;
	wire n4342;
	wire n4343;
	wire n4344;
	wire n4345;
	wire n4346;
	wire n4347;
	wire n4348;
	wire n4349;
	wire n4350;
	wire n4351;
	wire n4352;
	wire n4353;
	wire n4354;
	wire n4355;
	wire n4356;
	wire n4357;
	wire n4358;
	wire n4359;
	wire n4360;
	wire n4361;
	wire n4362;
	wire n4364;
	wire n4365;
	wire n4366;
	wire n4367;
	wire n4368;
	wire n4369;
	wire n4370;
	wire n4371;
	wire n4372;
	wire n4373;
	wire n4374;
	wire n4375;
	wire n4376;
	wire n4377;
	wire n4378;
	wire n4379;
	wire n4380;
	wire n4381;
	wire n4382;
	wire n4383;
	wire n4384;
	wire n4385;
	wire n4386;
	wire n4387;
	wire n4388;
	wire n4389;
	wire n4390;
	wire n4391;
	wire n4392;
	wire n4393;
	wire n4394;
	wire n4395;
	wire n4396;
	wire n4397;
	wire n4398;
	wire n4399;
	wire n4400;
	wire n4401;
	wire n4402;
	wire n4403;
	wire n4404;
	wire n4405;
	wire n4406;
	wire n4407;
	wire n4408;
	wire n4409;
	wire n4410;
	wire n4411;
	wire n4412;
	wire n4413;
	wire n4414;
	wire n4415;
	wire n4416;
	wire n4417;
	wire n4418;
	wire n4419;
	wire n4420;
	wire n4421;
	wire n4422;
	wire n4423;
	wire n4424;
	wire n4425;
	wire n4426;
	wire n4427;
	wire n4428;
	wire n4429;
	wire n4430;
	wire n4431;
	wire n4432;
	wire n4433;
	wire n4434;
	wire n4435;
	wire n4436;
	wire n4437;
	wire n4438;
	wire n4439;
	wire n4440;
	wire n4441;
	wire n4442;
	wire n4443;
	wire n4444;
	wire n4445;
	wire n4446;
	wire n4447;
	wire n4448;
	wire n4449;
	wire n4450;
	wire n4451;
	wire n4452;
	wire n4453;
	wire n4454;
	wire n4456;
	wire n4457;
	wire n4458;
	wire n4459;
	wire n4460;
	wire n4461;
	wire n4462;
	wire n4463;
	wire n4464;
	wire n4465;
	wire n4466;
	wire n4467;
	wire n4468;
	wire n4469;
	wire n4470;
	wire n4471;
	wire n4472;
	wire n4473;
	wire n4474;
	wire n4475;
	wire n4476;
	wire n4477;
	wire n4478;
	wire n4479;
	wire n4480;
	wire n4481;
	wire n4482;
	wire n4483;
	wire n4484;
	wire n4485;
	wire n4486;
	wire n4487;
	wire n4488;
	wire n4489;
	wire n4490;
	wire n4491;
	wire n4492;
	wire n4493;
	wire n4494;
	wire n4495;
	wire n4496;
	wire n4497;
	wire n4498;
	wire n4499;
	wire n4500;
	wire n4501;
	wire n4502;
	wire n4503;
	wire n4504;
	wire n4505;
	wire n4506;
	wire n4507;
	wire n4508;
	wire n4509;
	wire n4510;
	wire n4511;
	wire n4512;
	wire n4513;
	wire n4514;
	wire n4515;
	wire n4516;
	wire n4517;
	wire n4518;
	wire n4519;
	wire n4520;
	wire n4521;
	wire n4522;
	wire n4523;
	wire n4524;
	wire n4525;
	wire n4526;
	wire n4527;
	wire n4528;
	wire n4529;
	wire n4530;
	wire n4531;
	wire n4532;
	wire n4533;
	wire n4534;
	wire n4535;
	wire n4536;
	wire n4537;
	wire n4538;
	wire n4539;
	wire n4540;
	wire n4541;
	wire n4542;
	wire n4543;
	wire n4544;
	wire n4546;
	wire n4547;
	wire n4548;
	wire n4549;
	wire n4550;
	wire n4551;
	wire n4552;
	wire n4553;
	wire n4554;
	wire n4555;
	wire n4556;
	wire n4557;
	wire n4558;
	wire n4559;
	wire n4560;
	wire n4561;
	wire n4562;
	wire n4563;
	wire n4564;
	wire n4565;
	wire n4566;
	wire n4567;
	wire n4568;
	wire n4569;
	wire n4570;
	wire n4571;
	wire n4572;
	wire n4573;
	wire n4574;
	wire n4575;
	wire n4576;
	wire n4577;
	wire n4578;
	wire n4579;
	wire n4580;
	wire n4581;
	wire n4582;
	wire n4583;
	wire n4584;
	wire n4585;
	wire n4586;
	wire n4587;
	wire n4588;
	wire n4589;
	wire n4590;
	wire n4591;
	wire n4592;
	wire n4593;
	wire n4594;
	wire n4595;
	wire n4596;
	wire n4597;
	wire n4598;
	wire n4599;
	wire n4600;
	wire n4601;
	wire n4602;
	wire n4603;
	wire n4604;
	wire n4605;
	wire n4606;
	wire n4607;
	wire n4608;
	wire n4609;
	wire n4610;
	wire n4611;
	wire n4612;
	wire n4613;
	wire n4614;
	wire n4615;
	wire n4616;
	wire n4617;
	wire n4618;
	wire n4619;
	wire n4620;
	wire n4621;
	wire n4622;
	wire n4623;
	wire n4624;
	wire n4625;
	wire n4626;
	wire n4627;
	wire n4628;
	wire n4629;
	wire n4630;
	wire n4632;
	wire n4633;
	wire n4634;
	wire n4635;
	wire n4636;
	wire n4637;
	wire n4638;
	wire n4639;
	wire n4640;
	wire n4641;
	wire n4642;
	wire n4643;
	wire n4644;
	wire n4645;
	wire n4646;
	wire n4647;
	wire n4648;
	wire n4649;
	wire n4650;
	wire n4651;
	wire n4652;
	wire n4653;
	wire n4654;
	wire n4655;
	wire n4656;
	wire n4657;
	wire n4658;
	wire n4659;
	wire n4660;
	wire n4661;
	wire n4662;
	wire n4663;
	wire n4664;
	wire n4665;
	wire n4666;
	wire n4667;
	wire n4668;
	wire n4669;
	wire n4670;
	wire n4671;
	wire n4672;
	wire n4673;
	wire n4674;
	wire n4675;
	wire n4676;
	wire n4677;
	wire n4678;
	wire n4679;
	wire n4680;
	wire n4681;
	wire n4682;
	wire n4683;
	wire n4684;
	wire n4685;
	wire n4686;
	wire n4687;
	wire n4688;
	wire n4689;
	wire n4690;
	wire n4691;
	wire n4692;
	wire n4693;
	wire n4694;
	wire n4695;
	wire n4696;
	wire n4697;
	wire n4698;
	wire n4699;
	wire n4700;
	wire n4701;
	wire n4702;
	wire n4703;
	wire n4704;
	wire n4705;
	wire n4706;
	wire n4707;
	wire n4708;
	wire n4709;
	wire n4710;
	wire n4711;
	wire n4712;
	wire n4713;
	wire n4714;
	wire n4716;
	wire n4717;
	wire n4718;
	wire n4719;
	wire n4720;
	wire n4721;
	wire n4722;
	wire n4723;
	wire n4724;
	wire n4725;
	wire n4726;
	wire n4727;
	wire n4728;
	wire n4729;
	wire n4730;
	wire n4731;
	wire n4732;
	wire n4733;
	wire n4734;
	wire n4735;
	wire n4736;
	wire n4737;
	wire n4738;
	wire n4739;
	wire n4740;
	wire n4741;
	wire n4742;
	wire n4743;
	wire n4744;
	wire n4745;
	wire n4746;
	wire n4747;
	wire n4748;
	wire n4749;
	wire n4750;
	wire n4751;
	wire n4752;
	wire n4753;
	wire n4754;
	wire n4755;
	wire n4756;
	wire n4757;
	wire n4758;
	wire n4759;
	wire n4760;
	wire n4761;
	wire n4762;
	wire n4763;
	wire n4764;
	wire n4765;
	wire n4766;
	wire n4767;
	wire n4768;
	wire n4769;
	wire n4770;
	wire n4771;
	wire n4772;
	wire n4773;
	wire n4774;
	wire n4775;
	wire n4776;
	wire n4777;
	wire n4778;
	wire n4779;
	wire n4780;
	wire n4781;
	wire n4782;
	wire n4783;
	wire n4784;
	wire n4785;
	wire n4786;
	wire n4787;
	wire n4789;
	wire n4790;
	wire n4791;
	wire n4792;
	wire n4793;
	wire n4794;
	wire n4795;
	wire n4796;
	wire n4797;
	wire n4798;
	wire n4799;
	wire n4800;
	wire n4801;
	wire n4802;
	wire n4803;
	wire n4804;
	wire n4805;
	wire n4806;
	wire n4807;
	wire n4808;
	wire n4809;
	wire n4810;
	wire n4811;
	wire n4812;
	wire n4813;
	wire n4814;
	wire n4815;
	wire n4816;
	wire n4817;
	wire n4818;
	wire n4819;
	wire n4820;
	wire n4821;
	wire n4822;
	wire n4823;
	wire n4824;
	wire n4825;
	wire n4826;
	wire n4827;
	wire n4828;
	wire n4829;
	wire n4830;
	wire n4831;
	wire n4832;
	wire n4833;
	wire n4834;
	wire n4835;
	wire n4836;
	wire n4837;
	wire n4838;
	wire n4839;
	wire n4840;
	wire n4841;
	wire n4842;
	wire n4843;
	wire n4844;
	wire n4845;
	wire n4846;
	wire n4847;
	wire n4848;
	wire n4849;
	wire n4850;
	wire n4851;
	wire n4852;
	wire n4853;
	wire n4854;
	wire n4855;
	wire n4856;
	wire n4857;
	wire n4858;
	wire n4859;
	wire n4860;
	wire n4861;
	wire n4862;
	wire n4863;
	wire n4864;
	wire n4865;
	wire n4866;
	wire n4867;
	wire n4868;
	wire n4869;
	wire n4871;
	wire n4872;
	wire n4873;
	wire n4874;
	wire n4875;
	wire n4876;
	wire n4877;
	wire n4878;
	wire n4879;
	wire n4880;
	wire n4881;
	wire n4882;
	wire n4883;
	wire n4884;
	wire n4885;
	wire n4886;
	wire n4887;
	wire n4888;
	wire n4889;
	wire n4890;
	wire n4891;
	wire n4892;
	wire n4893;
	wire n4894;
	wire n4895;
	wire n4896;
	wire n4897;
	wire n4898;
	wire n4899;
	wire n4900;
	wire n4901;
	wire n4902;
	wire n4903;
	wire n4904;
	wire n4905;
	wire n4906;
	wire n4907;
	wire n4908;
	wire n4909;
	wire n4910;
	wire n4911;
	wire n4912;
	wire n4913;
	wire n4914;
	wire n4915;
	wire n4916;
	wire n4917;
	wire n4918;
	wire n4919;
	wire n4920;
	wire n4921;
	wire n4922;
	wire n4923;
	wire n4924;
	wire n4925;
	wire n4926;
	wire n4927;
	wire n4928;
	wire n4929;
	wire n4930;
	wire n4931;
	wire n4932;
	wire n4933;
	wire n4934;
	wire n4935;
	wire n4937;
	wire n4938;
	wire n4939;
	wire n4940;
	wire n4941;
	wire n4942;
	wire n4943;
	wire n4944;
	wire n4945;
	wire n4946;
	wire n4947;
	wire n4948;
	wire n4949;
	wire n4950;
	wire n4951;
	wire n4952;
	wire n4953;
	wire n4954;
	wire n4955;
	wire n4956;
	wire n4957;
	wire n4958;
	wire n4959;
	wire n4960;
	wire n4961;
	wire n4962;
	wire n4963;
	wire n4964;
	wire n4965;
	wire n4966;
	wire n4967;
	wire n4968;
	wire n4969;
	wire n4970;
	wire n4971;
	wire n4972;
	wire n4973;
	wire n4974;
	wire n4975;
	wire n4976;
	wire n4977;
	wire n4978;
	wire n4979;
	wire n4980;
	wire n4981;
	wire n4982;
	wire n4983;
	wire n4984;
	wire n4985;
	wire n4986;
	wire n4987;
	wire n4988;
	wire n4989;
	wire n4990;
	wire n4991;
	wire n4992;
	wire n4993;
	wire n4994;
	wire n4995;
	wire n4996;
	wire n4997;
	wire n4998;
	wire n4999;
	wire n5000;
	wire n5001;
	wire n5002;
	wire n5003;
	wire n5004;
	wire n5005;
	wire n5007;
	wire n5008;
	wire n5009;
	wire n5010;
	wire n5011;
	wire n5012;
	wire n5013;
	wire n5014;
	wire n5015;
	wire n5016;
	wire n5017;
	wire n5018;
	wire n5019;
	wire n5020;
	wire n5021;
	wire n5022;
	wire n5023;
	wire n5024;
	wire n5025;
	wire n5026;
	wire n5027;
	wire n5028;
	wire n5029;
	wire n5030;
	wire n5031;
	wire n5032;
	wire n5033;
	wire n5034;
	wire n5035;
	wire n5036;
	wire n5037;
	wire n5038;
	wire n5039;
	wire n5040;
	wire n5041;
	wire n5042;
	wire n5043;
	wire n5044;
	wire n5045;
	wire n5046;
	wire n5047;
	wire n5048;
	wire n5049;
	wire n5050;
	wire n5051;
	wire n5052;
	wire n5053;
	wire n5054;
	wire n5055;
	wire n5056;
	wire n5057;
	wire n5058;
	wire n5059;
	wire n5061;
	wire n5062;
	wire n5063;
	wire n5064;
	wire n5065;
	wire n5066;
	wire n5067;
	wire n5068;
	wire n5069;
	wire n5070;
	wire n5071;
	wire n5072;
	wire n5073;
	wire n5074;
	wire n5075;
	wire n5076;
	wire n5077;
	wire n5078;
	wire n5079;
	wire n5080;
	wire n5081;
	wire n5082;
	wire n5083;
	wire n5084;
	wire n5085;
	wire n5086;
	wire n5087;
	wire n5088;
	wire n5089;
	wire n5090;
	wire n5091;
	wire n5092;
	wire n5093;
	wire n5094;
	wire n5095;
	wire n5096;
	wire n5097;
	wire n5098;
	wire n5099;
	wire n5100;
	wire n5101;
	wire n5102;
	wire n5103;
	wire n5104;
	wire n5105;
	wire n5106;
	wire n5107;
	wire n5108;
	wire n5109;
	wire n5110;
	wire n5111;
	wire n5112;
	wire n5113;
	wire n5114;
	wire n5116;
	wire n5117;
	wire n5118;
	wire n5119;
	wire n5120;
	wire n5121;
	wire n5122;
	wire n5123;
	wire n5124;
	wire n5125;
	wire n5126;
	wire n5127;
	wire n5128;
	wire n5129;
	wire n5130;
	wire n5131;
	wire n5132;
	wire n5133;
	wire n5134;
	wire n5135;
	wire n5136;
	wire n5137;
	wire n5138;
	wire n5139;
	wire n5140;
	wire n5141;
	wire n5142;
	wire n5143;
	wire n5144;
	wire n5145;
	wire n5146;
	wire n5147;
	wire n5148;
	wire n5149;
	wire n5150;
	wire n5151;
	wire n5152;
	wire n5153;
	wire n5154;
	wire n5155;
	wire n5156;
	wire n5157;
	wire n5158;
	wire n5159;
	wire n5160;
	wire n5161;
	wire n5162;
	wire n5163;
	wire n5164;
	wire n5165;
	wire n5167;
	wire n5168;
	wire n5169;
	wire n5170;
	wire n5171;
	wire n5172;
	wire n5173;
	wire n5174;
	wire n5175;
	wire n5176;
	wire n5177;
	wire n5178;
	wire n5179;
	wire n5180;
	wire n5181;
	wire n5182;
	wire n5183;
	wire n5184;
	wire n5185;
	wire n5186;
	wire n5187;
	wire n5188;
	wire n5189;
	wire n5190;
	wire n5191;
	wire n5192;
	wire n5193;
	wire n5194;
	wire n5195;
	wire n5196;
	wire n5197;
	wire n5198;
	wire n5199;
	wire n5200;
	wire n5201;
	wire n5202;
	wire n5203;
	wire n5204;
	wire n5205;
	wire n5206;
	wire n5207;
	wire n5208;
	wire n5209;
	wire n5210;
	wire n5211;
	wire n5213;
	wire n5214;
	wire n5215;
	wire n5216;
	wire n5217;
	wire n5218;
	wire n5219;
	wire n5220;
	wire n5221;
	wire n5222;
	wire n5223;
	wire n5224;
	wire n5225;
	wire n5226;
	wire n5227;
	wire n5228;
	wire n5229;
	wire n5230;
	wire n5231;
	wire n5232;
	wire n5233;
	wire n5234;
	wire n5235;
	wire n5236;
	wire n5237;
	wire n5238;
	wire n5239;
	wire n5240;
	wire n5241;
	wire n5242;
	wire n5243;
	wire n5244;
	wire n5245;
	wire n5246;
	wire n5247;
	wire n5248;
	wire n5249;
	wire n5251;
	wire n5252;
	wire n5253;
	wire n5254;
	wire n5255;
	wire n5256;
	wire n5257;
	wire n5258;
	wire n5259;
	wire n5260;
	wire n5261;
	wire n5262;
	wire n5263;
	wire n5264;
	wire n5265;
	wire n5266;
	wire n5267;
	wire n5268;
	wire n5269;
	wire n5270;
	wire n5271;
	wire n5272;
	wire n5273;
	wire n5274;
	wire n5275;
	wire n5276;
	wire n5277;
	wire n5278;
	wire n5279;
	wire n5280;
	wire n5281;
	wire n5282;
	wire n5283;
	wire n5284;
	wire n5285;
	wire n5286;
	wire n5287;
	wire n5288;
	wire n5289;
	wire n5290;
	wire n5291;
	wire n5292;
	wire n5293;
	wire n5294;
	wire n5295;
	wire n5296;
	wire n5297;
	wire n5298;
	wire n5299;
	wire n5300;
	wire n5301;
	wire n5302;
	wire n5303;
	wire n5304;
	wire n5305;
	wire n5306;
	wire n5307;
	wire n5308;
	wire n5309;
	wire n5310;
	wire n5311;
	wire n5312;
	wire n5313;
	wire n5314;
	wire n5315;
	wire n5316;
	wire n5317;
	wire n5318;
	wire n5319;
	wire n5320;
	wire n5321;
	wire n5322;
	wire n5323;
	wire n5324;
	wire n5325;
	wire n5326;
	wire n5327;
	wire n5328;
	wire n5329;
	wire n5330;
	wire n5331;
	wire n5332;
	wire n5333;
	wire n5334;
	wire n5335;
	wire n5336;
	wire n5337;
	wire n5338;
	wire n5339;
	wire n5340;
	wire n5341;
	wire n5342;
	wire n5343;
	wire n5344;
	wire n5345;
	wire n5346;
	wire n5347;
	wire n5348;
	wire n5349;
	wire n5350;
	wire n5351;
	wire n5352;
	wire n5354;
	wire n5355;
	wire n5356;
	wire n5357;
	wire n5358;
	wire n5359;
	wire n5360;
	wire n5361;
	wire n5362;
	wire n5363;
	wire n5364;
	wire n5365;
	wire n5366;
	wire n5367;
	wire n5368;
	wire n5369;
	wire n5370;
	wire n5371;
	wire n5372;
	wire n5373;
	wire n5374;
	wire n5375;
	wire n5376;
	wire n5377;
	wire n5378;
	wire n5379;
	wire n5381;
	wire n5382;
	wire n5383;
	wire n5384;
	wire n5385;
	wire n5386;
	wire n5387;
	wire n5388;
	wire n5389;
	wire n5390;
	wire n5391;
	wire n5392;
	wire n5393;
	wire n5394;
	wire n5395;
	wire n5396;
	wire n5397;
	wire n5398;
	wire n5399;
	wire n5400;
	wire n5401;
	wire n5403;
	wire n5404;
	wire n5405;
	wire n5406;
	wire n5407;
	wire n5408;
	wire n5409;
	wire n5410;
	wire n5411;
	wire n5412;
	wire n5413;
	wire n5414;
	wire n5415;
	wire n5416;
	wire n5417;
	wire n5418;
	wire n5419;
	wire n5421;
	wire n5422;
	wire n5423;
	wire n5424;
	wire n5425;
	wire n5426;
	wire n5427;
	wire n5428;
	wire n5429;
	wire n5430;
	wire n5431;
	wire n5432;
	wire n5433;
	wire n5434;
	wire n5435;
	wire n5436;
	wire n5437;
	wire n5438;
	wire n5439;
	wire n5440;
	wire n5441;
	wire n5442;
	wire n5444;
	wire n5445;
	wire n5446;
	wire n5447;
	wire n5448;
	wire n5449;
	wire n5450;
	wire n5451;
	wire n5452;
	wire n5453;
	wire n5454;
	wire n5455;
	wire n5456;
	wire n5458;
	wire n5459;
	wire n5460;
	wire n5461;
	wire n5462;
	wire n5463;
	wire n5464;
	wire n5465;
	wire n5466;
	wire n5467;
	wire n5468;
	wire n5469;
	wire n5470;
	wire n5471;
	wire n5472;
	wire n5473;
	wire n5474;
	wire n5475;
	wire n5476;
	wire n5478;
	wire n5479;
	wire n5480;
	wire n5481;
	wire n5482;
	wire n5483;
	wire n5484;
	wire n5485;
	wire n5486;
	wire n5487;
	wire n5488;
	wire n5490;
	wire n5491;
	wire n5492;
	wire n5493;
	wire n5494;
	wire n5495;
	wire n5496;
	wire n5497;
	wire n5498;
	wire n5499;
	wire n5500;
	wire n5501;
	wire n5502;
	wire n5503;
	wire[2:0] w_a0_0;
	wire[2:0] w_a1_0;
	wire[1:0] w_a2_0;
	wire[1:0] w_a3_0;
	wire[1:0] w_a4_0;
	wire[1:0] w_a5_0;
	wire[1:0] w_a6_0;
	wire[1:0] w_a7_0;
	wire[1:0] w_a8_0;
	wire[1:0] w_a9_0;
	wire[1:0] w_a10_0;
	wire[1:0] w_a11_0;
	wire[1:0] w_a12_0;
	wire[1:0] w_a13_0;
	wire[1:0] w_a14_0;
	wire[1:0] w_a15_0;
	wire[1:0] w_a16_0;
	wire[1:0] w_a17_0;
	wire[1:0] w_a18_0;
	wire[2:0] w_a19_0;
	wire[2:0] w_a20_0;
	wire[1:0] w_a21_0;
	wire[2:0] w_a22_0;
	wire[1:0] w_sin0_0;
	wire sin0_fa_;
	wire[2:0] w_n49_0;
	wire[2:0] w_n49_1;
	wire[2:0] w_n49_2;
	wire[2:0] w_n49_3;
	wire[2:0] w_n49_4;
	wire[2:0] w_n49_5;
	wire[2:0] w_n49_6;
	wire[2:0] w_n49_7;
	wire[2:0] w_n49_8;
	wire[2:0] w_n49_9;
	wire[2:0] w_n50_0;
	wire[1:0] w_n51_0;
	wire[1:0] w_n52_0;
	wire[1:0] w_n53_0;
	wire[1:0] w_n54_0;
	wire[1:0] w_n55_0;
	wire[1:0] w_n56_0;
	wire[1:0] w_n57_0;
	wire[1:0] w_n58_0;
	wire[1:0] w_n59_0;
	wire[1:0] w_n60_0;
	wire[1:0] w_n61_0;
	wire[1:0] w_n62_0;
	wire[1:0] w_n63_0;
	wire[1:0] w_n64_0;
	wire[1:0] w_n65_0;
	wire[1:0] w_n66_0;
	wire[1:0] w_n67_0;
	wire[1:0] w_n68_0;
	wire[1:0] w_n69_0;
	wire[2:0] w_n70_0;
	wire[1:0] w_n70_1;
	wire[1:0] w_n71_0;
	wire[1:0] w_n72_0;
	wire[1:0] w_n73_0;
	wire[2:0] w_n74_0;
	wire[1:0] w_n74_1;
	wire[2:0] w_n75_0;
	wire[2:0] w_n75_1;
	wire[1:0] w_n75_2;
	wire[2:0] w_n77_0;
	wire[2:0] w_n77_1;
	wire[2:0] w_n77_2;
	wire[2:0] w_n77_3;
	wire[2:0] w_n77_4;
	wire[2:0] w_n77_5;
	wire[2:0] w_n77_6;
	wire[2:0] w_n77_7;
	wire[2:0] w_n77_8;
	wire[2:0] w_n77_9;
	wire[2:0] w_n78_0;
	wire[2:0] w_n78_1;
	wire[2:0] w_n78_2;
	wire[2:0] w_n78_3;
	wire[1:0] w_n80_0;
	wire[2:0] w_n81_0;
	wire[2:0] w_n83_0;
	wire[2:0] w_n84_0;
	wire[2:0] w_n85_0;
	wire[1:0] w_n85_1;
	wire[2:0] w_n87_0;
	wire[1:0] w_n88_0;
	wire[2:0] w_n90_0;
	wire[2:0] w_n91_0;
	wire[1:0] w_n91_1;
	wire[2:0] w_n92_0;
	wire[2:0] w_n92_1;
	wire[2:0] w_n92_2;
	wire[2:0] w_n92_3;
	wire[2:0] w_n93_0;
	wire[2:0] w_n93_1;
	wire[2:0] w_n94_0;
	wire[2:0] w_n94_1;
	wire[2:0] w_n94_2;
	wire[1:0] w_n95_0;
	wire[2:0] w_n96_0;
	wire[1:0] w_n96_1;
	wire[2:0] w_n97_0;
	wire[1:0] w_n97_1;
	wire[2:0] w_n98_0;
	wire[2:0] w_n98_1;
	wire[2:0] w_n98_2;
	wire[2:0] w_n98_3;
	wire[2:0] w_n99_0;
	wire[2:0] w_n99_1;
	wire[2:0] w_n99_2;
	wire[1:0] w_n99_3;
	wire[2:0] w_n100_0;
	wire[2:0] w_n100_1;
	wire[2:0] w_n100_2;
	wire[2:0] w_n100_3;
	wire[2:0] w_n100_4;
	wire[2:0] w_n100_5;
	wire[2:0] w_n100_6;
	wire[2:0] w_n100_7;
	wire[2:0] w_n100_8;
	wire[2:0] w_n101_0;
	wire[2:0] w_n101_1;
	wire[2:0] w_n101_2;
	wire[2:0] w_n101_3;
	wire[2:0] w_n102_0;
	wire[2:0] w_n102_1;
	wire[2:0] w_n102_2;
	wire[1:0] w_n102_3;
	wire[2:0] w_n103_0;
	wire[1:0] w_n103_1;
	wire[2:0] w_n105_0;
	wire[1:0] w_n105_1;
	wire[2:0] w_n106_0;
	wire[1:0] w_n106_1;
	wire[1:0] w_n107_0;
	wire[2:0] w_n108_0;
	wire[2:0] w_n108_1;
	wire[2:0] w_n108_2;
	wire[2:0] w_n108_3;
	wire[2:0] w_n108_4;
	wire[1:0] w_n109_0;
	wire[2:0] w_n110_0;
	wire[2:0] w_n110_1;
	wire[2:0] w_n111_0;
	wire[1:0] w_n111_1;
	wire[2:0] w_n112_0;
	wire[2:0] w_n112_1;
	wire[2:0] w_n112_2;
	wire[2:0] w_n112_3;
	wire[1:0] w_n112_4;
	wire[2:0] w_n113_0;
	wire[2:0] w_n113_1;
	wire[2:0] w_n113_2;
	wire[2:0] w_n114_0;
	wire[2:0] w_n114_1;
	wire[2:0] w_n114_2;
	wire[2:0] w_n114_3;
	wire[2:0] w_n115_0;
	wire[1:0] w_n115_1;
	wire[2:0] w_n116_0;
	wire[2:0] w_n116_1;
	wire[2:0] w_n116_2;
	wire[1:0] w_n116_3;
	wire[2:0] w_n117_0;
	wire[1:0] w_n117_1;
	wire[2:0] w_n118_0;
	wire[2:0] w_n118_1;
	wire[2:0] w_n118_2;
	wire[2:0] w_n118_3;
	wire[2:0] w_n118_4;
	wire[2:0] w_n118_5;
	wire[2:0] w_n118_6;
	wire[1:0] w_n119_0;
	wire[2:0] w_n120_0;
	wire[2:0] w_n120_1;
	wire[2:0] w_n120_2;
	wire[2:0] w_n123_0;
	wire[2:0] w_n123_1;
	wire[1:0] w_n123_2;
	wire[2:0] w_n124_0;
	wire[2:0] w_n124_1;
	wire[2:0] w_n124_2;
	wire[2:0] w_n125_0;
	wire[2:0] w_n125_1;
	wire[2:0] w_n125_2;
	wire[2:0] w_n125_3;
	wire[2:0] w_n125_4;
	wire[1:0] w_n125_5;
	wire[2:0] w_n126_0;
	wire[2:0] w_n126_1;
	wire[2:0] w_n126_2;
	wire[2:0] w_n126_3;
	wire[1:0] w_n126_4;
	wire[2:0] w_n127_0;
	wire[2:0] w_n127_1;
	wire[2:0] w_n127_2;
	wire[1:0] w_n127_3;
	wire[2:0] w_n128_0;
	wire[2:0] w_n128_1;
	wire[2:0] w_n128_2;
	wire[1:0] w_n128_3;
	wire[2:0] w_n129_0;
	wire[2:0] w_n129_1;
	wire[2:0] w_n130_0;
	wire[2:0] w_n130_1;
	wire[2:0] w_n130_2;
	wire[1:0] w_n130_3;
	wire[1:0] w_n131_0;
	wire[2:0] w_n132_0;
	wire[2:0] w_n133_0;
	wire[2:0] w_n133_1;
	wire[1:0] w_n133_2;
	wire[2:0] w_n134_0;
	wire[1:0] w_n134_1;
	wire[2:0] w_n135_0;
	wire[2:0] w_n135_1;
	wire[2:0] w_n135_2;
	wire[2:0] w_n135_3;
	wire[2:0] w_n135_4;
	wire[2:0] w_n136_0;
	wire[2:0] w_n136_1;
	wire[1:0] w_n136_2;
	wire[2:0] w_n137_0;
	wire[2:0] w_n137_1;
	wire[1:0] w_n137_2;
	wire[2:0] w_n138_0;
	wire[2:0] w_n138_1;
	wire[2:0] w_n138_2;
	wire[2:0] w_n138_3;
	wire[1:0] w_n138_4;
	wire[2:0] w_n139_0;
	wire[1:0] w_n139_1;
	wire[2:0] w_n140_0;
	wire[2:0] w_n140_1;
	wire[2:0] w_n140_2;
	wire[1:0] w_n140_3;
	wire[1:0] w_n141_0;
	wire[2:0] w_n142_0;
	wire[2:0] w_n142_1;
	wire[1:0] w_n142_2;
	wire[2:0] w_n143_0;
	wire[1:0] w_n143_1;
	wire[2:0] w_n144_0;
	wire[2:0] w_n144_1;
	wire[2:0] w_n144_2;
	wire[2:0] w_n144_3;
	wire[2:0] w_n144_4;
	wire[2:0] w_n144_5;
	wire[2:0] w_n144_6;
	wire[2:0] w_n145_0;
	wire[2:0] w_n145_1;
	wire[2:0] w_n145_2;
	wire[1:0] w_n145_3;
	wire[1:0] w_n146_0;
	wire[2:0] w_n147_0;
	wire[2:0] w_n147_1;
	wire[1:0] w_n147_2;
	wire[2:0] w_n148_0;
	wire[1:0] w_n148_1;
	wire[1:0] w_n150_0;
	wire[2:0] w_n151_0;
	wire[2:0] w_n151_1;
	wire[2:0] w_n151_2;
	wire[2:0] w_n152_0;
	wire[2:0] w_n152_1;
	wire[2:0] w_n152_2;
	wire[2:0] w_n154_0;
	wire[2:0] w_n154_1;
	wire[2:0] w_n154_2;
	wire[2:0] w_n154_3;
	wire[2:0] w_n154_4;
	wire[2:0] w_n154_5;
	wire[2:0] w_n154_6;
	wire[2:0] w_n155_0;
	wire[2:0] w_n155_1;
	wire[2:0] w_n155_2;
	wire[2:0] w_n155_3;
	wire[2:0] w_n157_0;
	wire[2:0] w_n157_1;
	wire[2:0] w_n157_2;
	wire[1:0] w_n157_3;
	wire[2:0] w_n158_0;
	wire[2:0] w_n158_1;
	wire[2:0] w_n159_0;
	wire[1:0] w_n159_1;
	wire[2:0] w_n160_0;
	wire[2:0] w_n160_1;
	wire[2:0] w_n160_2;
	wire[2:0] w_n161_0;
	wire[2:0] w_n162_0;
	wire[2:0] w_n162_1;
	wire[1:0] w_n162_2;
	wire[2:0] w_n165_0;
	wire[2:0] w_n165_1;
	wire[2:0] w_n165_2;
	wire[2:0] w_n166_0;
	wire[2:0] w_n166_1;
	wire[2:0] w_n166_2;
	wire[2:0] w_n167_0;
	wire[2:0] w_n167_1;
	wire[2:0] w_n167_2;
	wire[2:0] w_n167_3;
	wire[2:0] w_n168_0;
	wire[2:0] w_n168_1;
	wire[1:0] w_n168_2;
	wire[2:0] w_n169_0;
	wire[2:0] w_n169_1;
	wire[1:0] w_n169_2;
	wire[2:0] w_n170_0;
	wire[2:0] w_n170_1;
	wire[2:0] w_n170_2;
	wire[1:0] w_n170_3;
	wire[2:0] w_n171_0;
	wire[2:0] w_n171_1;
	wire[2:0] w_n171_2;
	wire[2:0] w_n171_3;
	wire[1:0] w_n171_4;
	wire[1:0] w_n172_0;
	wire[2:0] w_n173_0;
	wire[2:0] w_n173_1;
	wire[2:0] w_n174_0;
	wire[2:0] w_n174_1;
	wire[2:0] w_n174_2;
	wire[2:0] w_n174_3;
	wire[2:0] w_n174_4;
	wire[2:0] w_n174_5;
	wire[2:0] w_n174_6;
	wire[2:0] w_n176_0;
	wire[2:0] w_n176_1;
	wire[1:0] w_n177_0;
	wire[2:0] w_n180_0;
	wire[1:0] w_n180_1;
	wire[2:0] w_n182_0;
	wire[2:0] w_n182_1;
	wire[2:0] w_n182_2;
	wire[1:0] w_n182_3;
	wire[2:0] w_n183_0;
	wire[2:0] w_n184_0;
	wire[2:0] w_n184_1;
	wire[2:0] w_n184_2;
	wire[2:0] w_n184_3;
	wire[2:0] w_n184_4;
	wire[2:0] w_n184_5;
	wire[2:0] w_n184_6;
	wire[2:0] w_n185_0;
	wire[2:0] w_n185_1;
	wire[2:0] w_n185_2;
	wire[2:0] w_n185_3;
	wire[1:0] w_n186_0;
	wire[2:0] w_n187_0;
	wire[2:0] w_n187_1;
	wire[1:0] w_n187_2;
	wire[2:0] w_n188_0;
	wire[2:0] w_n188_1;
	wire[1:0] w_n188_2;
	wire[1:0] w_n189_0;
	wire[2:0] w_n190_0;
	wire[2:0] w_n190_1;
	wire[2:0] w_n191_0;
	wire[2:0] w_n191_1;
	wire[2:0] w_n191_2;
	wire[2:0] w_n191_3;
	wire[2:0] w_n192_0;
	wire[2:0] w_n192_1;
	wire[2:0] w_n192_2;
	wire[1:0] w_n192_3;
	wire[2:0] w_n193_0;
	wire[2:0] w_n193_1;
	wire[1:0] w_n193_2;
	wire[2:0] w_n194_0;
	wire[2:0] w_n195_0;
	wire[2:0] w_n195_1;
	wire[1:0] w_n195_2;
	wire[2:0] w_n197_0;
	wire[2:0] w_n197_1;
	wire[2:0] w_n197_2;
	wire[1:0] w_n197_3;
	wire[2:0] w_n198_0;
	wire[1:0] w_n198_1;
	wire[2:0] w_n203_0;
	wire[1:0] w_n203_1;
	wire[2:0] w_n204_0;
	wire[2:0] w_n204_1;
	wire[2:0] w_n204_2;
	wire[1:0] w_n205_0;
	wire[2:0] w_n206_0;
	wire[2:0] w_n206_1;
	wire[1:0] w_n206_2;
	wire[2:0] w_n207_0;
	wire[2:0] w_n207_1;
	wire[2:0] w_n207_2;
	wire[1:0] w_n207_3;
	wire[1:0] w_n212_0;
	wire[2:0] w_n213_0;
	wire[2:0] w_n213_1;
	wire[2:0] w_n213_2;
	wire[1:0] w_n213_3;
	wire[1:0] w_n214_0;
	wire[2:0] w_n215_0;
	wire[2:0] w_n215_1;
	wire[2:0] w_n215_2;
	wire[2:0] w_n215_3;
	wire[2:0] w_n216_0;
	wire[2:0] w_n217_0;
	wire[2:0] w_n217_1;
	wire[2:0] w_n217_2;
	wire[2:0] w_n217_3;
	wire[1:0] w_n217_4;
	wire[2:0] w_n218_0;
	wire[2:0] w_n218_1;
	wire[2:0] w_n218_2;
	wire[2:0] w_n218_3;
	wire[2:0] w_n221_0;
	wire[2:0] w_n221_1;
	wire[2:0] w_n221_2;
	wire[2:0] w_n221_3;
	wire[2:0] w_n222_0;
	wire[2:0] w_n222_1;
	wire[2:0] w_n222_2;
	wire[1:0] w_n222_3;
	wire[2:0] w_n223_0;
	wire[2:0] w_n223_1;
	wire[2:0] w_n223_2;
	wire[1:0] w_n223_3;
	wire[2:0] w_n224_0;
	wire[2:0] w_n224_1;
	wire[2:0] w_n224_2;
	wire[2:0] w_n224_3;
	wire[2:0] w_n224_4;
	wire[1:0] w_n224_5;
	wire[2:0] w_n226_0;
	wire[2:0] w_n226_1;
	wire[2:0] w_n226_2;
	wire[1:0] w_n229_0;
	wire[2:0] w_n230_0;
	wire[2:0] w_n230_1;
	wire[2:0] w_n230_2;
	wire[1:0] w_n230_3;
	wire[2:0] w_n231_0;
	wire[1:0] w_n231_1;
	wire[2:0] w_n232_0;
	wire[2:0] w_n232_1;
	wire[2:0] w_n232_2;
	wire[2:0] w_n232_3;
	wire[2:0] w_n232_4;
	wire[2:0] w_n233_0;
	wire[2:0] w_n233_1;
	wire[1:0] w_n233_2;
	wire[2:0] w_n234_0;
	wire[2:0] w_n235_0;
	wire[2:0] w_n235_1;
	wire[1:0] w_n235_2;
	wire[2:0] w_n236_0;
	wire[2:0] w_n236_1;
	wire[2:0] w_n238_0;
	wire[2:0] w_n238_1;
	wire[1:0] w_n238_2;
	wire[1:0] w_n239_0;
	wire[2:0] w_n240_0;
	wire[2:0] w_n240_1;
	wire[1:0] w_n240_2;
	wire[1:0] w_n241_0;
	wire[2:0] w_n244_0;
	wire[2:0] w_n244_1;
	wire[2:0] w_n244_2;
	wire[1:0] w_n244_3;
	wire[2:0] w_n245_0;
	wire[2:0] w_n245_1;
	wire[1:0] w_n245_2;
	wire[2:0] w_n246_0;
	wire[1:0] w_n247_0;
	wire[2:0] w_n248_0;
	wire[2:0] w_n248_1;
	wire[2:0] w_n248_2;
	wire[2:0] w_n248_3;
	wire[2:0] w_n249_0;
	wire[2:0] w_n249_1;
	wire[1:0] w_n249_2;
	wire[2:0] w_n250_0;
	wire[2:0] w_n250_1;
	wire[2:0] w_n250_2;
	wire[2:0] w_n251_0;
	wire[2:0] w_n252_0;
	wire[2:0] w_n252_1;
	wire[2:0] w_n252_2;
	wire[2:0] w_n252_3;
	wire[1:0] w_n252_4;
	wire[2:0] w_n253_0;
	wire[2:0] w_n253_1;
	wire[2:0] w_n253_2;
	wire[2:0] w_n253_3;
	wire[2:0] w_n253_4;
	wire[2:0] w_n253_5;
	wire[2:0] w_n253_6;
	wire[2:0] w_n254_0;
	wire[2:0] w_n255_0;
	wire[2:0] w_n255_1;
	wire[1:0] w_n255_2;
	wire[1:0] w_n260_0;
	wire[2:0] w_n261_0;
	wire[2:0] w_n261_1;
	wire[2:0] w_n261_2;
	wire[2:0] w_n262_0;
	wire[2:0] w_n262_1;
	wire[2:0] w_n262_2;
	wire[2:0] w_n262_3;
	wire[2:0] w_n262_4;
	wire[1:0] w_n262_5;
	wire[2:0] w_n263_0;
	wire[2:0] w_n263_1;
	wire[2:0] w_n263_2;
	wire[2:0] w_n263_3;
	wire[1:0] w_n263_4;
	wire[1:0] w_n264_0;
	wire[2:0] w_n265_0;
	wire[2:0] w_n265_1;
	wire[1:0] w_n265_2;
	wire[2:0] w_n266_0;
	wire[2:0] w_n266_1;
	wire[2:0] w_n267_0;
	wire[2:0] w_n267_1;
	wire[2:0] w_n267_2;
	wire[1:0] w_n267_3;
	wire[2:0] w_n268_0;
	wire[2:0] w_n268_1;
	wire[1:0] w_n268_2;
	wire[2:0] w_n269_0;
	wire[2:0] w_n269_1;
	wire[2:0] w_n269_2;
	wire[1:0] w_n273_0;
	wire[1:0] w_n274_0;
	wire[2:0] w_n275_0;
	wire[2:0] w_n275_1;
	wire[1:0] w_n275_2;
	wire[2:0] w_n276_0;
	wire[2:0] w_n276_1;
	wire[2:0] w_n276_2;
	wire[2:0] w_n276_3;
	wire[1:0] w_n277_0;
	wire[2:0] w_n278_0;
	wire[2:0] w_n278_1;
	wire[2:0] w_n279_0;
	wire[2:0] w_n280_0;
	wire[2:0] w_n280_1;
	wire[2:0] w_n280_2;
	wire[2:0] w_n281_0;
	wire[2:0] w_n282_0;
	wire[2:0] w_n282_1;
	wire[2:0] w_n283_0;
	wire[2:0] w_n283_1;
	wire[1:0] w_n283_2;
	wire[2:0] w_n286_0;
	wire[2:0] w_n286_1;
	wire[2:0] w_n286_2;
	wire[1:0] w_n286_3;
	wire[1:0] w_n287_0;
	wire[2:0] w_n288_0;
	wire[2:0] w_n288_1;
	wire[1:0] w_n288_2;
	wire[2:0] w_n289_0;
	wire[1:0] w_n289_1;
	wire[2:0] w_n290_0;
	wire[2:0] w_n290_1;
	wire[2:0] w_n290_2;
	wire[2:0] w_n290_3;
	wire[1:0] w_n293_0;
	wire[2:0] w_n294_0;
	wire[2:0] w_n294_1;
	wire[2:0] w_n294_2;
	wire[2:0] w_n294_3;
	wire[2:0] w_n295_0;
	wire[1:0] w_n296_0;
	wire[2:0] w_n297_0;
	wire[2:0] w_n297_1;
	wire[1:0] w_n299_0;
	wire[2:0] w_n300_0;
	wire[2:0] w_n300_1;
	wire[2:0] w_n300_2;
	wire[1:0] w_n300_3;
	wire[2:0] w_n301_0;
	wire[1:0] w_n301_1;
	wire[2:0] w_n302_0;
	wire[2:0] w_n303_0;
	wire[2:0] w_n305_0;
	wire[2:0] w_n305_1;
	wire[2:0] w_n305_2;
	wire[1:0] w_n307_0;
	wire[1:0] w_n308_0;
	wire[2:0] w_n309_0;
	wire[2:0] w_n309_1;
	wire[2:0] w_n309_2;
	wire[2:0] w_n310_0;
	wire[2:0] w_n310_1;
	wire[2:0] w_n310_2;
	wire[2:0] w_n311_0;
	wire[2:0] w_n311_1;
	wire[2:0] w_n311_2;
	wire[1:0] w_n312_0;
	wire[2:0] w_n313_0;
	wire[2:0] w_n313_1;
	wire[2:0] w_n314_0;
	wire[2:0] w_n315_0;
	wire[2:0] w_n315_1;
	wire[1:0] w_n315_2;
	wire[2:0] w_n316_0;
	wire[1:0] w_n320_0;
	wire[2:0] w_n321_0;
	wire[2:0] w_n321_1;
	wire[2:0] w_n321_2;
	wire[1:0] w_n321_3;
	wire[1:0] w_n324_0;
	wire[1:0] w_n325_0;
	wire[2:0] w_n327_0;
	wire[2:0] w_n327_1;
	wire[2:0] w_n329_0;
	wire[1:0] w_n329_1;
	wire[2:0] w_n330_0;
	wire[2:0] w_n331_0;
	wire[2:0] w_n331_1;
	wire[2:0] w_n331_2;
	wire[2:0] w_n332_0;
	wire[2:0] w_n332_1;
	wire[2:0] w_n332_2;
	wire[1:0] w_n332_3;
	wire[2:0] w_n333_0;
	wire[2:0] w_n333_1;
	wire[1:0] w_n333_2;
	wire[1:0] w_n334_0;
	wire[2:0] w_n335_0;
	wire[2:0] w_n336_0;
	wire[2:0] w_n336_1;
	wire[2:0] w_n336_2;
	wire[2:0] w_n337_0;
	wire[2:0] w_n337_1;
	wire[2:0] w_n337_2;
	wire[2:0] w_n338_0;
	wire[2:0] w_n339_0;
	wire[2:0] w_n339_1;
	wire[2:0] w_n339_2;
	wire[2:0] w_n339_3;
	wire[1:0] w_n339_4;
	wire[2:0] w_n340_0;
	wire[2:0] w_n340_1;
	wire[2:0] w_n344_0;
	wire[2:0] w_n344_1;
	wire[2:0] w_n344_2;
	wire[1:0] w_n344_3;
	wire[1:0] w_n345_0;
	wire[2:0] w_n346_0;
	wire[2:0] w_n346_1;
	wire[2:0] w_n346_2;
	wire[2:0] w_n347_0;
	wire[2:0] w_n347_1;
	wire[2:0] w_n347_2;
	wire[1:0] w_n350_0;
	wire[2:0] w_n351_0;
	wire[1:0] w_n351_1;
	wire[2:0] w_n352_0;
	wire[1:0] w_n352_1;
	wire[2:0] w_n353_0;
	wire[2:0] w_n353_1;
	wire[2:0] w_n353_2;
	wire[1:0] w_n355_0;
	wire[2:0] w_n359_0;
	wire[2:0] w_n360_0;
	wire[2:0] w_n361_0;
	wire[2:0] w_n361_1;
	wire[2:0] w_n361_2;
	wire[1:0] w_n362_0;
	wire[2:0] w_n366_0;
	wire[2:0] w_n366_1;
	wire[2:0] w_n366_2;
	wire[1:0] w_n366_3;
	wire[2:0] w_n370_0;
	wire[2:0] w_n370_1;
	wire[2:0] w_n370_2;
	wire[1:0] w_n370_3;
	wire[1:0] w_n372_0;
	wire[2:0] w_n373_0;
	wire[2:0] w_n374_0;
	wire[2:0] w_n374_1;
	wire[2:0] w_n374_2;
	wire[1:0] w_n374_3;
	wire[2:0] w_n377_0;
	wire[2:0] w_n377_1;
	wire[2:0] w_n377_2;
	wire[2:0] w_n377_3;
	wire[2:0] w_n378_0;
	wire[2:0] w_n378_1;
	wire[2:0] w_n378_2;
	wire[1:0] w_n378_3;
	wire[1:0] w_n381_0;
	wire[2:0] w_n382_0;
	wire[2:0] w_n382_1;
	wire[1:0] w_n382_2;
	wire[2:0] w_n383_0;
	wire[2:0] w_n383_1;
	wire[2:0] w_n383_2;
	wire[2:0] w_n384_0;
	wire[2:0] w_n384_1;
	wire[2:0] w_n384_2;
	wire[1:0] w_n384_3;
	wire[1:0] w_n385_0;
	wire[1:0] w_n386_0;
	wire[2:0] w_n387_0;
	wire[2:0] w_n387_1;
	wire[2:0] w_n387_2;
	wire[1:0] w_n387_3;
	wire[2:0] w_n388_0;
	wire[1:0] w_n388_1;
	wire[2:0] w_n389_0;
	wire[2:0] w_n389_1;
	wire[2:0] w_n389_2;
	wire[2:0] w_n389_3;
	wire[1:0] w_n394_0;
	wire[2:0] w_n395_0;
	wire[2:0] w_n395_1;
	wire[2:0] w_n395_2;
	wire[1:0] w_n396_0;
	wire[2:0] w_n398_0;
	wire[2:0] w_n399_0;
	wire[2:0] w_n400_0;
	wire[2:0] w_n401_0;
	wire[1:0] w_n402_0;
	wire[2:0] w_n403_0;
	wire[2:0] w_n404_0;
	wire[2:0] w_n404_1;
	wire[1:0] w_n407_0;
	wire[2:0] w_n409_0;
	wire[2:0] w_n409_1;
	wire[2:0] w_n409_2;
	wire[1:0] w_n410_0;
	wire[2:0] w_n411_0;
	wire[2:0] w_n411_1;
	wire[1:0] w_n411_2;
	wire[1:0] w_n413_0;
	wire[2:0] w_n415_0;
	wire[2:0] w_n415_1;
	wire[2:0] w_n415_2;
	wire[2:0] w_n417_0;
	wire[2:0] w_n418_0;
	wire[2:0] w_n418_1;
	wire[1:0] w_n418_2;
	wire[1:0] w_n420_0;
	wire[1:0] w_n425_0;
	wire[2:0] w_n426_0;
	wire[2:0] w_n427_0;
	wire[2:0] w_n427_1;
	wire[2:0] w_n427_2;
	wire[2:0] w_n429_0;
	wire[2:0] w_n429_1;
	wire[2:0] w_n430_0;
	wire[1:0] w_n430_1;
	wire[1:0] w_n433_0;
	wire[2:0] w_n434_0;
	wire[2:0] w_n434_1;
	wire[2:0] w_n434_2;
	wire[2:0] w_n435_0;
	wire[2:0] w_n435_1;
	wire[2:0] w_n435_2;
	wire[2:0] w_n436_0;
	wire[2:0] w_n437_0;
	wire[2:0] w_n437_1;
	wire[2:0] w_n438_0;
	wire[2:0] w_n438_1;
	wire[1:0] w_n438_2;
	wire[2:0] w_n439_0;
	wire[2:0] w_n439_1;
	wire[2:0] w_n439_2;
	wire[2:0] w_n439_3;
	wire[1:0] w_n439_4;
	wire[2:0] w_n443_0;
	wire[1:0] w_n443_1;
	wire[2:0] w_n445_0;
	wire[2:0] w_n445_1;
	wire[2:0] w_n445_2;
	wire[2:0] w_n446_0;
	wire[2:0] w_n446_1;
	wire[1:0] w_n446_2;
	wire[2:0] w_n447_0;
	wire[2:0] w_n448_0;
	wire[2:0] w_n448_1;
	wire[1:0] w_n448_2;
	wire[1:0] w_n452_0;
	wire[1:0] w_n455_0;
	wire[2:0] w_n456_0;
	wire[2:0] w_n457_0;
	wire[2:0] w_n459_0;
	wire[2:0] w_n460_0;
	wire[2:0] w_n460_1;
	wire[2:0] w_n460_2;
	wire[1:0] w_n460_3;
	wire[2:0] w_n461_0;
	wire[2:0] w_n462_0;
	wire[2:0] w_n462_1;
	wire[1:0] w_n462_2;
	wire[2:0] w_n463_0;
	wire[2:0] w_n467_0;
	wire[2:0] w_n467_1;
	wire[2:0] w_n467_2;
	wire[2:0] w_n468_0;
	wire[2:0] w_n470_0;
	wire[1:0] w_n477_0;
	wire[1:0] w_n480_0;
	wire[2:0] w_n481_0;
	wire[1:0] w_n481_1;
	wire[1:0] w_n482_0;
	wire[2:0] w_n486_0;
	wire[2:0] w_n486_1;
	wire[2:0] w_n488_0;
	wire[2:0] w_n488_1;
	wire[2:0] w_n488_2;
	wire[1:0] w_n488_3;
	wire[2:0] w_n489_0;
	wire[2:0] w_n489_1;
	wire[2:0] w_n489_2;
	wire[1:0] w_n489_3;
	wire[1:0] w_n491_0;
	wire[1:0] w_n492_0;
	wire[2:0] w_n495_0;
	wire[1:0] w_n496_0;
	wire[2:0] w_n497_0;
	wire[1:0] w_n497_1;
	wire[1:0] w_n500_0;
	wire[1:0] w_n504_0;
	wire[1:0] w_n505_0;
	wire[2:0] w_n506_0;
	wire[2:0] w_n506_1;
	wire[2:0] w_n506_2;
	wire[1:0] w_n509_0;
	wire[2:0] w_n510_0;
	wire[2:0] w_n510_1;
	wire[2:0] w_n510_2;
	wire[1:0] w_n510_3;
	wire[2:0] w_n513_0;
	wire[1:0] w_n514_0;
	wire[2:0] w_n516_0;
	wire[2:0] w_n517_0;
	wire[2:0] w_n519_0;
	wire[2:0] w_n519_1;
	wire[2:0] w_n519_2;
	wire[2:0] w_n519_3;
	wire[2:0] w_n519_4;
	wire[2:0] w_n519_5;
	wire[1:0] w_n521_0;
	wire[1:0] w_n522_0;
	wire[1:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n525_0;
	wire[1:0] w_n526_0;
	wire[2:0] w_n527_0;
	wire[2:0] w_n527_1;
	wire[2:0] w_n527_2;
	wire[2:0] w_n527_3;
	wire[1:0] w_n528_0;
	wire[1:0] w_n530_0;
	wire[1:0] w_n531_0;
	wire[1:0] w_n532_0;
	wire[2:0] w_n534_0;
	wire[2:0] w_n534_1;
	wire[2:0] w_n534_2;
	wire[2:0] w_n535_0;
	wire[2:0] w_n535_1;
	wire[1:0] w_n535_2;
	wire[1:0] w_n537_0;
	wire[2:0] w_n539_0;
	wire[2:0] w_n539_1;
	wire[2:0] w_n540_0;
	wire[1:0] w_n543_0;
	wire[1:0] w_n544_0;
	wire[2:0] w_n546_0;
	wire[1:0] w_n551_0;
	wire[2:0] w_n552_0;
	wire[1:0] w_n553_0;
	wire[1:0] w_n555_0;
	wire[1:0] w_n557_0;
	wire[1:0] w_n559_0;
	wire[1:0] w_n560_0;
	wire[2:0] w_n561_0;
	wire[1:0] w_n561_1;
	wire[2:0] w_n562_0;
	wire[1:0] w_n562_1;
	wire[1:0] w_n563_0;
	wire[1:0] w_n567_0;
	wire[2:0] w_n568_0;
	wire[2:0] w_n569_0;
	wire[2:0] w_n569_1;
	wire[1:0] w_n569_2;
	wire[2:0] w_n570_0;
	wire[2:0] w_n570_1;
	wire[1:0] w_n570_2;
	wire[1:0] w_n572_0;
	wire[1:0] w_n574_0;
	wire[1:0] w_n575_0;
	wire[1:0] w_n577_0;
	wire[1:0] w_n579_0;
	wire[1:0] w_n582_0;
	wire[1:0] w_n583_0;
	wire[2:0] w_n586_0;
	wire[2:0] w_n587_0;
	wire[2:0] w_n587_1;
	wire[2:0] w_n587_2;
	wire[1:0] w_n587_3;
	wire[2:0] w_n588_0;
	wire[1:0] w_n593_0;
	wire[2:0] w_n594_0;
	wire[1:0] w_n598_0;
	wire[1:0] w_n599_0;
	wire[2:0] w_n600_0;
	wire[2:0] w_n600_1;
	wire[2:0] w_n600_2;
	wire[1:0] w_n601_0;
	wire[1:0] w_n602_0;
	wire[1:0] w_n603_0;
	wire[1:0] w_n604_0;
	wire[2:0] w_n607_0;
	wire[2:0] w_n607_1;
	wire[1:0] w_n607_2;
	wire[1:0] w_n609_0;
	wire[1:0] w_n610_0;
	wire[1:0] w_n612_0;
	wire[1:0] w_n613_0;
	wire[1:0] w_n616_0;
	wire[2:0] w_n617_0;
	wire[1:0] w_n619_0;
	wire[2:0] w_n624_0;
	wire[1:0] w_n625_0;
	wire[1:0] w_n628_0;
	wire[2:0] w_n630_0;
	wire[2:0] w_n634_0;
	wire[1:0] w_n644_0;
	wire[1:0] w_n645_0;
	wire[1:0] w_n646_0;
	wire[1:0] w_n648_0;
	wire[2:0] w_n652_0;
	wire[2:0] w_n654_0;
	wire[1:0] w_n655_0;
	wire[1:0] w_n660_0;
	wire[1:0] w_n661_0;
	wire[1:0] w_n663_0;
	wire[1:0] w_n666_0;
	wire[1:0] w_n667_0;
	wire[1:0] w_n669_0;
	wire[1:0] w_n673_0;
	wire[2:0] w_n676_0;
	wire[2:0] w_n677_0;
	wire[1:0] w_n677_1;
	wire[2:0] w_n684_0;
	wire[1:0] w_n685_0;
	wire[1:0] w_n686_0;
	wire[2:0] w_n689_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n697_0;
	wire[1:0] w_n700_0;
	wire[1:0] w_n702_0;
	wire[2:0] w_n705_0;
	wire[1:0] w_n706_0;
	wire[1:0] w_n708_0;
	wire[2:0] w_n716_0;
	wire[2:0] w_n716_1;
	wire[2:0] w_n716_2;
	wire[2:0] w_n716_3;
	wire[2:0] w_n716_4;
	wire[2:0] w_n716_5;
	wire[2:0] w_n716_6;
	wire[2:0] w_n716_7;
	wire[2:0] w_n716_8;
	wire[2:0] w_n717_0;
	wire[2:0] w_n717_1;
	wire[2:0] w_n717_2;
	wire[1:0] w_n717_3;
	wire[1:0] w_n720_0;
	wire[1:0] w_n723_0;
	wire[1:0] w_n725_0;
	wire[1:0] w_n727_0;
	wire[1:0] w_n744_0;
	wire[1:0] w_n749_0;
	wire[1:0] w_n751_0;
	wire[2:0] w_n752_0;
	wire[1:0] w_n766_0;
	wire[2:0] w_n777_0;
	wire[1:0] w_n785_0;
	wire[1:0] w_n786_0;
	wire[1:0] w_n787_0;
	wire[1:0] w_n788_0;
	wire[1:0] w_n796_0;
	wire[1:0] w_n802_0;
	wire[1:0] w_n803_0;
	wire[1:0] w_n813_0;
	wire[1:0] w_n814_0;
	wire[2:0] w_n815_0;
	wire[1:0] w_n815_1;
	wire[1:0] w_n816_0;
	wire[2:0] w_n817_0;
	wire[2:0] w_n817_1;
	wire[1:0] w_n824_0;
	wire[2:0] w_n825_0;
	wire[2:0] w_n825_1;
	wire[1:0] w_n826_0;
	wire[2:0] w_n827_0;
	wire[1:0] w_n834_0;
	wire[1:0] w_n835_0;
	wire[1:0] w_n841_0;
	wire[1:0] w_n842_0;
	wire[1:0] w_n847_0;
	wire[2:0] w_n849_0;
	wire[2:0] w_n850_0;
	wire[2:0] w_n852_0;
	wire[1:0] w_n852_1;
	wire[2:0] w_n853_0;
	wire[1:0] w_n856_0;
	wire[1:0] w_n858_0;
	wire[1:0] w_n862_0;
	wire[1:0] w_n863_0;
	wire[1:0] w_n866_0;
	wire[1:0] w_n871_0;
	wire[2:0] w_n876_0;
	wire[1:0] w_n876_1;
	wire[2:0] w_n877_0;
	wire[2:0] w_n878_0;
	wire[2:0] w_n878_1;
	wire[2:0] w_n880_0;
	wire[2:0] w_n880_1;
	wire[2:0] w_n880_2;
	wire[2:0] w_n880_3;
	wire[2:0] w_n880_4;
	wire[2:0] w_n880_5;
	wire[1:0] w_n880_6;
	wire[2:0] w_n881_0;
	wire[2:0] w_n881_1;
	wire[2:0] w_n881_2;
	wire[2:0] w_n881_3;
	wire[2:0] w_n881_4;
	wire[2:0] w_n884_0;
	wire[1:0] w_n884_1;
	wire[2:0] w_n886_0;
	wire[1:0] w_n886_1;
	wire[2:0] w_n896_0;
	wire[2:0] w_n897_0;
	wire[2:0] w_n897_1;
	wire[1:0] w_n897_2;
	wire[1:0] w_n903_0;
	wire[2:0] w_n904_0;
	wire[1:0] w_n904_1;
	wire[2:0] w_n912_0;
	wire[2:0] w_n915_0;
	wire[1:0] w_n919_0;
	wire[1:0] w_n921_0;
	wire[2:0] w_n924_0;
	wire[2:0] w_n930_0;
	wire[2:0] w_n930_1;
	wire[1:0] w_n930_2;
	wire[1:0] w_n931_0;
	wire[1:0] w_n965_0;
	wire[1:0] w_n966_0;
	wire[1:0] w_n968_0;
	wire[1:0] w_n974_0;
	wire[1:0] w_n975_0;
	wire[2:0] w_n987_0;
	wire[1:0] w_n987_1;
	wire[2:0] w_n989_0;
	wire[2:0] w_n989_1;
	wire[1:0] w_n989_2;
	wire[2:0] w_n992_0;
	wire[2:0] w_n992_1;
	wire[2:0] w_n992_2;
	wire[2:0] w_n992_3;
	wire[2:0] w_n994_0;
	wire[2:0] w_n994_1;
	wire[2:0] w_n994_2;
	wire[2:0] w_n994_3;
	wire[2:0] w_n994_4;
	wire[2:0] w_n994_5;
	wire[1:0] w_n994_6;
	wire[2:0] w_n996_0;
	wire[2:0] w_n996_1;
	wire[2:0] w_n996_2;
	wire[2:0] w_n996_3;
	wire[2:0] w_n996_4;
	wire[2:0] w_n997_0;
	wire[2:0] w_n997_1;
	wire[2:0] w_n997_2;
	wire[2:0] w_n997_3;
	wire[1:0] w_n997_4;
	wire[1:0] w_n1001_0;
	wire[1:0] w_n1002_0;
	wire[2:0] w_n1005_0;
	wire[2:0] w_n1005_1;
	wire[2:0] w_n1005_2;
	wire[2:0] w_n1005_3;
	wire[1:0] w_n1005_4;
	wire[1:0] w_n1006_0;
	wire[1:0] w_n1009_0;
	wire[1:0] w_n1012_0;
	wire[2:0] w_n1016_0;
	wire[1:0] w_n1016_1;
	wire[1:0] w_n1017_0;
	wire[1:0] w_n1019_0;
	wire[1:0] w_n1021_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1023_0;
	wire[2:0] w_n1024_0;
	wire[2:0] w_n1025_0;
	wire[1:0] w_n1026_0;
	wire[1:0] w_n1030_0;
	wire[1:0] w_n1032_0;
	wire[1:0] w_n1033_0;
	wire[2:0] w_n1035_0;
	wire[2:0] w_n1035_1;
	wire[2:0] w_n1035_2;
	wire[2:0] w_n1039_0;
	wire[1:0] w_n1040_0;
	wire[1:0] w_n1043_0;
	wire[1:0] w_n1045_0;
	wire[1:0] w_n1050_0;
	wire[1:0] w_n1053_0;
	wire[2:0] w_n1055_0;
	wire[2:0] w_n1055_1;
	wire[1:0] w_n1055_2;
	wire[1:0] w_n1056_0;
	wire[1:0] w_n1057_0;
	wire[1:0] w_n1060_0;
	wire[2:0] w_n1064_0;
	wire[1:0] w_n1064_1;
	wire[1:0] w_n1066_0;
	wire[1:0] w_n1069_0;
	wire[1:0] w_n1071_0;
	wire[2:0] w_n1072_0;
	wire[1:0] w_n1072_1;
	wire[2:0] w_n1073_0;
	wire[1:0] w_n1073_1;
	wire[2:0] w_n1074_0;
	wire[2:0] w_n1074_1;
	wire[1:0] w_n1078_0;
	wire[1:0] w_n1079_0;
	wire[1:0] w_n1080_0;
	wire[1:0] w_n1085_0;
	wire[2:0] w_n1087_0;
	wire[1:0] w_n1088_0;
	wire[1:0] w_n1093_0;
	wire[1:0] w_n1094_0;
	wire[2:0] w_n1095_0;
	wire[2:0] w_n1095_1;
	wire[2:0] w_n1095_2;
	wire[2:0] w_n1096_0;
	wire[1:0] w_n1097_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1104_0;
	wire[2:0] w_n1105_0;
	wire[1:0] w_n1109_0;
	wire[2:0] w_n1110_0;
	wire[2:0] w_n1114_0;
	wire[2:0] w_n1115_0;
	wire[1:0] w_n1115_1;
	wire[1:0] w_n1120_0;
	wire[1:0] w_n1122_0;
	wire[1:0] w_n1124_0;
	wire[2:0] w_n1127_0;
	wire[1:0] w_n1130_0;
	wire[1:0] w_n1133_0;
	wire[2:0] w_n1135_0;
	wire[1:0] w_n1135_1;
	wire[1:0] w_n1140_0;
	wire[1:0] w_n1147_0;
	wire[2:0] w_n1149_0;
	wire[2:0] w_n1149_1;
	wire[1:0] w_n1150_0;
	wire[2:0] w_n1151_0;
	wire[2:0] w_n1151_1;
	wire[2:0] w_n1152_0;
	wire[2:0] w_n1152_1;
	wire[1:0] w_n1152_2;
	wire[2:0] w_n1154_0;
	wire[2:0] w_n1154_1;
	wire[2:0] w_n1154_2;
	wire[2:0] w_n1154_3;
	wire[2:0] w_n1154_4;
	wire[2:0] w_n1154_5;
	wire[2:0] w_n1154_6;
	wire[2:0] w_n1154_7;
	wire[2:0] w_n1154_8;
	wire[2:0] w_n1154_9;
	wire[2:0] w_n1154_10;
	wire[2:0] w_n1156_0;
	wire[2:0] w_n1156_1;
	wire[2:0] w_n1156_2;
	wire[2:0] w_n1156_3;
	wire[2:0] w_n1156_4;
	wire[2:0] w_n1156_5;
	wire[2:0] w_n1156_6;
	wire[2:0] w_n1156_7;
	wire[2:0] w_n1156_8;
	wire[2:0] w_n1156_9;
	wire[2:0] w_n1156_10;
	wire[2:0] w_n1156_11;
	wire[1:0] w_n1156_12;
	wire[1:0] w_n1158_0;
	wire[2:0] w_n1160_0;
	wire[2:0] w_n1160_1;
	wire[1:0] w_n1160_2;
	wire[2:0] w_n1163_0;
	wire[2:0] w_n1164_0;
	wire[2:0] w_n1164_1;
	wire[2:0] w_n1164_2;
	wire[2:0] w_n1164_3;
	wire[2:0] w_n1166_0;
	wire[2:0] w_n1166_1;
	wire[2:0] w_n1166_2;
	wire[2:0] w_n1166_3;
	wire[2:0] w_n1166_4;
	wire[2:0] w_n1166_5;
	wire[1:0] w_n1166_6;
	wire[2:0] w_n1168_0;
	wire[2:0] w_n1168_1;
	wire[2:0] w_n1168_2;
	wire[2:0] w_n1168_3;
	wire[2:0] w_n1168_4;
	wire[2:0] w_n1170_0;
	wire[2:0] w_n1170_1;
	wire[2:0] w_n1170_2;
	wire[2:0] w_n1170_3;
	wire[1:0] w_n1170_4;
	wire[1:0] w_n1173_0;
	wire[1:0] w_n1176_0;
	wire[2:0] w_n1178_0;
	wire[1:0] w_n1180_0;
	wire[1:0] w_n1181_0;
	wire[1:0] w_n1185_0;
	wire[1:0] w_n1186_0;
	wire[1:0] w_n1188_0;
	wire[1:0] w_n1189_0;
	wire[1:0] w_n1192_0;
	wire[2:0] w_n1196_0;
	wire[1:0] w_n1196_1;
	wire[1:0] w_n1205_0;
	wire[1:0] w_n1215_0;
	wire[1:0] w_n1226_0;
	wire[2:0] w_n1232_0;
	wire[1:0] w_n1235_0;
	wire[1:0] w_n1243_0;
	wire[1:0] w_n1249_0;
	wire[1:0] w_n1250_0;
	wire[2:0] w_n1252_0;
	wire[1:0] w_n1253_0;
	wire[2:0] w_n1254_0;
	wire[2:0] w_n1254_1;
	wire[1:0] w_n1254_2;
	wire[2:0] w_n1255_0;
	wire[2:0] w_n1255_1;
	wire[1:0] w_n1255_2;
	wire[2:0] w_n1257_0;
	wire[2:0] w_n1257_1;
	wire[2:0] w_n1257_2;
	wire[2:0] w_n1257_3;
	wire[2:0] w_n1257_4;
	wire[2:0] w_n1257_5;
	wire[2:0] w_n1257_6;
	wire[2:0] w_n1257_7;
	wire[2:0] w_n1257_8;
	wire[2:0] w_n1257_9;
	wire[2:0] w_n1257_10;
	wire[2:0] w_n1257_11;
	wire[2:0] w_n1257_12;
	wire[2:0] w_n1257_13;
	wire[2:0] w_n1259_0;
	wire[2:0] w_n1259_1;
	wire[2:0] w_n1259_2;
	wire[2:0] w_n1259_3;
	wire[2:0] w_n1259_4;
	wire[2:0] w_n1259_5;
	wire[2:0] w_n1259_6;
	wire[2:0] w_n1259_7;
	wire[2:0] w_n1259_8;
	wire[1:0] w_n1259_9;
	wire[2:0] w_n1260_0;
	wire[2:0] w_n1261_0;
	wire[2:0] w_n1261_1;
	wire[2:0] w_n1261_2;
	wire[2:0] w_n1266_0;
	wire[2:0] w_n1266_1;
	wire[2:0] w_n1266_2;
	wire[2:0] w_n1266_3;
	wire[2:0] w_n1266_4;
	wire[2:0] w_n1266_5;
	wire[1:0] w_n1266_6;
	wire[1:0] w_n1268_0;
	wire[2:0] w_n1270_0;
	wire[2:0] w_n1270_1;
	wire[2:0] w_n1270_2;
	wire[2:0] w_n1270_3;
	wire[2:0] w_n1272_0;
	wire[2:0] w_n1272_1;
	wire[2:0] w_n1272_2;
	wire[2:0] w_n1272_3;
	wire[2:0] w_n1272_4;
	wire[2:0] w_n1294_0;
	wire[2:0] w_n1295_0;
	wire[2:0] w_n1295_1;
	wire[2:0] w_n1295_2;
	wire[2:0] w_n1295_3;
	wire[1:0] w_n1299_0;
	wire[1:0] w_n1300_0;
	wire[1:0] w_n1302_0;
	wire[1:0] w_n1312_0;
	wire[1:0] w_n1313_0;
	wire[1:0] w_n1319_0;
	wire[2:0] w_n1322_0;
	wire[2:0] w_n1322_1;
	wire[2:0] w_n1331_0;
	wire[1:0] w_n1332_0;
	wire[1:0] w_n1339_0;
	wire[1:0] w_n1343_0;
	wire[2:0] w_n1345_0;
	wire[2:0] w_n1345_1;
	wire[1:0] w_n1346_0;
	wire[2:0] w_n1353_0;
	wire[2:0] w_n1353_1;
	wire[2:0] w_n1353_2;
	wire[2:0] w_n1353_3;
	wire[2:0] w_n1353_4;
	wire[2:0] w_n1353_5;
	wire[2:0] w_n1354_0;
	wire[2:0] w_n1354_1;
	wire[2:0] w_n1354_2;
	wire[2:0] w_n1354_3;
	wire[2:0] w_n1356_0;
	wire[2:0] w_n1356_1;
	wire[2:0] w_n1356_2;
	wire[2:0] w_n1356_3;
	wire[2:0] w_n1356_4;
	wire[2:0] w_n1356_5;
	wire[2:0] w_n1356_6;
	wire[2:0] w_n1356_7;
	wire[2:0] w_n1356_8;
	wire[2:0] w_n1356_9;
	wire[2:0] w_n1356_10;
	wire[2:0] w_n1356_11;
	wire[1:0] w_n1356_12;
	wire[2:0] w_n1360_0;
	wire[2:0] w_n1360_1;
	wire[2:0] w_n1360_2;
	wire[2:0] w_n1360_3;
	wire[2:0] w_n1360_4;
	wire[2:0] w_n1360_5;
	wire[1:0] w_n1360_6;
	wire[1:0] w_n1363_0;
	wire[2:0] w_n1365_0;
	wire[2:0] w_n1366_0;
	wire[1:0] w_n1366_1;
	wire[1:0] w_n1375_0;
	wire[1:0] w_n1378_0;
	wire[1:0] w_n1381_0;
	wire[1:0] w_n1385_0;
	wire[1:0] w_n1387_0;
	wire[1:0] w_n1392_0;
	wire[2:0] w_n1400_0;
	wire[2:0] w_n1402_0;
	wire[2:0] w_n1402_1;
	wire[2:0] w_n1403_0;
	wire[1:0] w_n1403_1;
	wire[2:0] w_n1404_0;
	wire[1:0] w_n1406_0;
	wire[1:0] w_n1407_0;
	wire[1:0] w_n1415_0;
	wire[2:0] w_n1416_0;
	wire[2:0] w_n1416_1;
	wire[1:0] w_n1416_2;
	wire[2:0] w_n1418_0;
	wire[2:0] w_n1418_1;
	wire[2:0] w_n1418_2;
	wire[1:0] w_n1425_0;
	wire[1:0] w_n1426_0;
	wire[1:0] w_n1427_0;
	wire[1:0] w_n1429_0;
	wire[1:0] w_n1432_0;
	wire[2:0] w_n1434_0;
	wire[2:0] w_n1434_1;
	wire[2:0] w_n1434_2;
	wire[2:0] w_n1434_3;
	wire[2:0] w_n1434_4;
	wire[2:0] w_n1434_5;
	wire[2:0] w_n1434_6;
	wire[2:0] w_n1438_0;
	wire[2:0] w_n1438_1;
	wire[2:0] w_n1438_2;
	wire[2:0] w_n1438_3;
	wire[2:0] w_n1438_4;
	wire[2:0] w_n1438_5;
	wire[2:0] w_n1438_6;
	wire[2:0] w_n1438_7;
	wire[2:0] w_n1438_8;
	wire[2:0] w_n1438_9;
	wire[2:0] w_n1438_10;
	wire[2:0] w_n1438_11;
	wire[2:0] w_n1438_12;
	wire[2:0] w_n1438_13;
	wire[2:0] w_n1438_14;
	wire[2:0] w_n1438_15;
	wire[2:0] w_n1438_16;
	wire[2:0] w_n1438_17;
	wire[2:0] w_n1438_18;
	wire[2:0] w_n1438_19;
	wire[2:0] w_n1438_20;
	wire[1:0] w_n1438_21;
	wire[1:0] w_n1441_0;
	wire[1:0] w_n1444_0;
	wire[1:0] w_n1447_0;
	wire[1:0] w_n1448_0;
	wire[1:0] w_n1452_0;
	wire[1:0] w_n1456_0;
	wire[2:0] w_n1459_0;
	wire[2:0] w_n1460_0;
	wire[2:0] w_n1460_1;
	wire[1:0] w_n1467_0;
	wire[1:0] w_n1470_0;
	wire[2:0] w_n1474_0;
	wire[2:0] w_n1474_1;
	wire[2:0] w_n1474_2;
	wire[2:0] w_n1474_3;
	wire[2:0] w_n1474_4;
	wire[2:0] w_n1474_5;
	wire[2:0] w_n1474_6;
	wire[1:0] w_n1474_7;
	wire[1:0] w_n1478_0;
	wire[2:0] w_n1480_0;
	wire[2:0] w_n1480_1;
	wire[2:0] w_n1480_2;
	wire[2:0] w_n1480_3;
	wire[2:0] w_n1480_4;
	wire[2:0] w_n1480_5;
	wire[2:0] w_n1480_6;
	wire[2:0] w_n1480_7;
	wire[2:0] w_n1480_8;
	wire[2:0] w_n1480_9;
	wire[1:0] w_n1480_10;
	wire[2:0] w_n1485_0;
	wire[2:0] w_n1485_1;
	wire[2:0] w_n1485_2;
	wire[2:0] w_n1485_3;
	wire[2:0] w_n1485_4;
	wire[1:0] w_n1489_0;
	wire[2:0] w_n1490_0;
	wire[2:0] w_n1490_1;
	wire[2:0] w_n1490_2;
	wire[2:0] w_n1490_3;
	wire[2:0] w_n1490_4;
	wire[1:0] w_n1490_5;
	wire[1:0] w_n1491_0;
	wire[2:0] w_n1493_0;
	wire[2:0] w_n1493_1;
	wire[2:0] w_n1493_2;
	wire[2:0] w_n1493_3;
	wire[2:0] w_n1493_4;
	wire[1:0] w_n1493_5;
	wire[2:0] w_n1494_0;
	wire[2:0] w_n1494_1;
	wire[2:0] w_n1494_2;
	wire[2:0] w_n1494_3;
	wire[2:0] w_n1494_4;
	wire[2:0] w_n1494_5;
	wire[1:0] w_n1494_6;
	wire[2:0] w_n1499_0;
	wire[2:0] w_n1499_1;
	wire[2:0] w_n1499_2;
	wire[2:0] w_n1499_3;
	wire[2:0] w_n1499_4;
	wire[2:0] w_n1499_5;
	wire[2:0] w_n1500_0;
	wire[2:0] w_n1500_1;
	wire[2:0] w_n1500_2;
	wire[2:0] w_n1500_3;
	wire[2:0] w_n1500_4;
	wire[1:0] w_n1500_5;
	wire[2:0] w_n1504_0;
	wire[2:0] w_n1504_1;
	wire[2:0] w_n1504_2;
	wire[2:0] w_n1504_3;
	wire[2:0] w_n1505_0;
	wire[2:0] w_n1505_1;
	wire[2:0] w_n1505_2;
	wire[2:0] w_n1505_3;
	wire[2:0] w_n1505_4;
	wire[1:0] w_n1508_0;
	wire[1:0] w_n1509_0;
	wire[1:0] w_n1511_0;
	wire[1:0] w_n1513_0;
	wire[2:0] w_n1516_0;
	wire[1:0] w_n1518_0;
	wire[1:0] w_n1520_0;
	wire[1:0] w_n1523_0;
	wire[1:0] w_n1528_0;
	wire[2:0] w_n1529_0;
	wire[1:0] w_n1531_0;
	wire[2:0] w_n1532_0;
	wire[1:0] w_n1533_0;
	wire[2:0] w_n1534_0;
	wire[2:0] w_n1539_0;
	wire[2:0] w_n1539_1;
	wire[2:0] w_n1539_2;
	wire[1:0] w_n1541_0;
	wire[2:0] w_n1542_0;
	wire[2:0] w_n1542_1;
	wire[2:0] w_n1542_2;
	wire[1:0] w_n1545_0;
	wire[1:0] w_n1547_0;
	wire[2:0] w_n1549_0;
	wire[2:0] w_n1549_1;
	wire[2:0] w_n1549_2;
	wire[2:0] w_n1549_3;
	wire[2:0] w_n1549_4;
	wire[2:0] w_n1551_0;
	wire[2:0] w_n1551_1;
	wire[2:0] w_n1551_2;
	wire[2:0] w_n1551_3;
	wire[2:0] w_n1551_4;
	wire[1:0] w_n1555_0;
	wire[1:0] w_n1556_0;
	wire[1:0] w_n1557_0;
	wire[2:0] w_n1558_0;
	wire[2:0] w_n1558_1;
	wire[2:0] w_n1558_2;
	wire[2:0] w_n1558_3;
	wire[1:0] w_n1558_4;
	wire[2:0] w_n1560_0;
	wire[2:0] w_n1560_1;
	wire[2:0] w_n1560_2;
	wire[2:0] w_n1560_3;
	wire[2:0] w_n1560_4;
	wire[1:0] w_n1563_0;
	wire[1:0] w_n1564_0;
	wire[1:0] w_n1566_0;
	wire[1:0] w_n1567_0;
	wire[1:0] w_n1575_0;
	wire[2:0] w_n1576_0;
	wire[1:0] w_n1584_0;
	wire[1:0] w_n1592_0;
	wire[1:0] w_n1593_0;
	wire[1:0] w_n1594_0;
	wire[1:0] w_n1595_0;
	wire[1:0] w_n1598_0;
	wire[1:0] w_n1601_0;
	wire[1:0] w_n1604_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1613_0;
	wire[1:0] w_n1614_0;
	wire[1:0] w_n1615_0;
	wire[1:0] w_n1616_0;
	wire[2:0] w_n1622_0;
	wire[2:0] w_n1622_1;
	wire[2:0] w_n1622_2;
	wire[2:0] w_n1622_3;
	wire[1:0] w_n1622_4;
	wire[1:0] w_n1625_0;
	wire[1:0] w_n1626_0;
	wire[1:0] w_n1629_0;
	wire[1:0] w_n1630_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1632_0;
	wire[1:0] w_n1640_0;
	wire[1:0] w_n1648_0;
	wire[2:0] w_n1649_0;
	wire[2:0] w_n1651_0;
	wire[1:0] w_n1651_1;
	wire[2:0] w_n1656_0;
	wire[2:0] w_n1656_1;
	wire[1:0] w_n1659_0;
	wire[1:0] w_n1660_0;
	wire[1:0] w_n1661_0;
	wire[1:0] w_n1662_0;
	wire[1:0] w_n1663_0;
	wire[2:0] w_n1664_0;
	wire[1:0] w_n1673_0;
	wire[1:0] w_n1674_0;
	wire[1:0] w_n1680_0;
	wire[1:0] w_n1687_0;
	wire[1:0] w_n1696_0;
	wire[1:0] w_n1697_0;
	wire[1:0] w_n1699_0;
	wire[1:0] w_n1700_0;
	wire[1:0] w_n1702_0;
	wire[1:0] w_n1703_0;
	wire[1:0] w_n1705_0;
	wire[1:0] w_n1706_0;
	wire[1:0] w_n1708_0;
	wire[1:0] w_n1709_0;
	wire[1:0] w_n1710_0;
	wire[1:0] w_n1718_0;
	wire[1:0] w_n1725_0;
	wire[1:0] w_n1733_0;
	wire[1:0] w_n1734_0;
	wire[1:0] w_n1736_0;
	wire[1:0] w_n1737_0;
	wire[1:0] w_n1743_0;
	wire[2:0] w_n1744_0;
	wire[1:0] w_n1746_0;
	wire[1:0] w_n1747_0;
	wire[1:0] w_n1754_0;
	wire[1:0] w_n1755_0;
	wire[1:0] w_n1756_0;
	wire[1:0] w_n1757_0;
	wire[1:0] w_n1759_0;
	wire[1:0] w_n1763_0;
	wire[1:0] w_n1764_0;
	wire[1:0] w_n1765_0;
	wire[1:0] w_n1766_0;
	wire[2:0] w_n1767_0;
	wire[1:0] w_n1768_0;
	wire[1:0] w_n1770_0;
	wire[1:0] w_n1778_0;
	wire[1:0] w_n1783_0;
	wire[1:0] w_n1793_0;
	wire[1:0] w_n1794_0;
	wire[1:0] w_n1796_0;
	wire[1:0] w_n1799_0;
	wire[1:0] w_n1800_0;
	wire[1:0] w_n1802_0;
	wire[1:0] w_n1804_0;
	wire[1:0] w_n1806_0;
	wire[1:0] w_n1811_0;
	wire[1:0] w_n1812_0;
	wire[2:0] w_n1813_0;
	wire[1:0] w_n1813_1;
	wire[1:0] w_n1814_0;
	wire[1:0] w_n1815_0;
	wire[1:0] w_n1823_0;
	wire[1:0] w_n1830_0;
	wire[1:0] w_n1832_0;
	wire[1:0] w_n1833_0;
	wire[1:0] w_n1835_0;
	wire[1:0] w_n1836_0;
	wire[1:0] w_n1838_0;
	wire[1:0] w_n1839_0;
	wire[1:0] w_n1840_0;
	wire[1:0] w_n1842_0;
	wire[1:0] w_n1843_0;
	wire[1:0] w_n1844_0;
	wire[1:0] w_n1846_0;
	wire[1:0] w_n1850_0;
	wire[1:0] w_n1860_0;
	wire[1:0] w_n1865_0;
	wire[1:0] w_n1867_0;
	wire[2:0] w_n1868_0;
	wire[1:0] w_n1873_0;
	wire[1:0] w_n1885_0;
	wire[1:0] w_n1886_0;
	wire[1:0] w_n1888_0;
	wire[2:0] w_n1890_0;
	wire[2:0] w_n1895_0;
	wire[2:0] w_n1902_0;
	wire[1:0] w_n1903_0;
	wire[1:0] w_n1904_0;
	wire[2:0] w_n1908_0;
	wire[1:0] w_n1910_0;
	wire[1:0] w_n1921_0;
	wire[1:0] w_n1922_0;
	wire[1:0] w_n1930_0;
	wire[1:0] w_n1933_0;
	wire[1:0] w_n1938_0;
	wire[1:0] w_n1939_0;
	wire[1:0] w_n1940_0;
	wire[1:0] w_n1950_0;
	wire[1:0] w_n1953_0;
	wire[1:0] w_n1954_0;
	wire[2:0] w_n1955_0;
	wire[2:0] w_n1956_0;
	wire[2:0] w_n1956_1;
	wire[2:0] w_n1956_2;
	wire[2:0] w_n1956_3;
	wire[2:0] w_n1956_4;
	wire[2:0] w_n1956_5;
	wire[2:0] w_n1956_6;
	wire[1:0] w_n1956_7;
	wire[2:0] w_n1957_0;
	wire[2:0] w_n1958_0;
	wire[1:0] w_n1958_1;
	wire[2:0] w_n1959_0;
	wire[2:0] w_n1960_0;
	wire[2:0] w_n1961_0;
	wire[1:0] w_n1962_0;
	wire[1:0] w_n1965_0;
	wire[1:0] w_n1970_0;
	wire[1:0] w_n1974_0;
	wire[1:0] w_n1979_0;
	wire[1:0] w_n1984_0;
	wire[2:0] w_n1987_0;
	wire[2:0] w_n1993_0;
	wire[1:0] w_n1994_0;
	wire[1:0] w_n1996_0;
	wire[1:0] w_n1999_0;
	wire[1:0] w_n2002_0;
	wire[1:0] w_n2014_0;
	wire[1:0] w_n2023_0;
	wire[1:0] w_n2026_0;
	wire[1:0] w_n2029_0;
	wire[1:0] w_n2037_0;
	wire[1:0] w_n2040_0;
	wire[1:0] w_n2041_0;
	wire[1:0] w_n2044_0;
	wire[1:0] w_n2045_0;
	wire[1:0] w_n2046_0;
	wire[1:0] w_n2049_0;
	wire[2:0] w_n2051_0;
	wire[2:0] w_n2051_1;
	wire[2:0] w_n2051_2;
	wire[2:0] w_n2051_3;
	wire[2:0] w_n2051_4;
	wire[2:0] w_n2051_5;
	wire[2:0] w_n2051_6;
	wire[2:0] w_n2051_7;
	wire[1:0] w_n2051_8;
	wire[1:0] w_n2058_0;
	wire[1:0] w_n2059_0;
	wire[1:0] w_n2060_0;
	wire[1:0] w_n2061_0;
	wire[1:0] w_n2062_0;
	wire[1:0] w_n2070_0;
	wire[1:0] w_n2078_0;
	wire[1:0] w_n2086_0;
	wire[1:0] w_n2087_0;
	wire[1:0] w_n2088_0;
	wire[1:0] w_n2089_0;
	wire[1:0] w_n2090_0;
	wire[2:0] w_n2091_0;
	wire[1:0] w_n2091_1;
	wire[2:0] w_n2092_0;
	wire[1:0] w_n2093_0;
	wire[2:0] w_n2094_0;
	wire[2:0] w_n2094_1;
	wire[2:0] w_n2094_2;
	wire[2:0] w_n2094_3;
	wire[2:0] w_n2094_4;
	wire[2:0] w_n2094_5;
	wire[2:0] w_n2094_6;
	wire[1:0] w_n2095_0;
	wire[2:0] w_n2096_0;
	wire[1:0] w_n2096_1;
	wire[2:0] w_n2097_0;
	wire[2:0] w_n2098_0;
	wire[1:0] w_n2099_0;
	wire[1:0] w_n2100_0;
	wire[2:0] w_n2101_0;
	wire[1:0] w_n2101_1;
	wire[2:0] w_n2103_0;
	wire[1:0] w_n2105_0;
	wire[2:0] w_n2107_0;
	wire[1:0] w_n2110_0;
	wire[2:0] w_n2112_0;
	wire[1:0] w_n2112_1;
	wire[1:0] w_n2115_0;
	wire[2:0] w_n2116_0;
	wire[2:0] w_n2116_1;
	wire[2:0] w_n2116_2;
	wire[1:0] w_n2120_0;
	wire[1:0] w_n2126_0;
	wire[2:0] w_n2127_0;
	wire[1:0] w_n2127_1;
	wire[1:0] w_n2130_0;
	wire[2:0] w_n2134_0;
	wire[2:0] w_n2135_0;
	wire[2:0] w_n2142_0;
	wire[2:0] w_n2146_0;
	wire[1:0] w_n2147_0;
	wire[1:0] w_n2149_0;
	wire[1:0] w_n2154_0;
	wire[2:0] w_n2155_0;
	wire[1:0] w_n2155_1;
	wire[2:0] w_n2166_0;
	wire[1:0] w_n2167_0;
	wire[1:0] w_n2169_0;
	wire[1:0] w_n2172_0;
	wire[1:0] w_n2175_0;
	wire[1:0] w_n2183_0;
	wire[1:0] w_n2186_0;
	wire[1:0] w_n2187_0;
	wire[1:0] w_n2190_0;
	wire[1:0] w_n2191_0;
	wire[1:0] w_n2192_0;
	wire[1:0] w_n2195_0;
	wire[1:0] w_n2203_0;
	wire[1:0] w_n2211_0;
	wire[1:0] w_n2219_0;
	wire[1:0] w_n2220_0;
	wire[1:0] w_n2221_0;
	wire[1:0] w_n2226_0;
	wire[1:0] w_n2227_0;
	wire[1:0] w_n2228_0;
	wire[1:0] w_n2229_0;
	wire[1:0] w_n2230_0;
	wire[1:0] w_n2231_0;
	wire[1:0] w_n2232_0;
	wire[2:0] w_n2233_0;
	wire[1:0] w_n2233_1;
	wire[2:0] w_n2234_0;
	wire[2:0] w_n2235_0;
	wire[2:0] w_n2236_0;
	wire[2:0] w_n2236_1;
	wire[2:0] w_n2236_2;
	wire[2:0] w_n2236_3;
	wire[2:0] w_n2236_4;
	wire[1:0] w_n2236_5;
	wire[2:0] w_n2238_0;
	wire[1:0] w_n2238_1;
	wire[2:0] w_n2244_0;
	wire[1:0] w_n2248_0;
	wire[1:0] w_n2249_0;
	wire[1:0] w_n2251_0;
	wire[2:0] w_n2252_0;
	wire[2:0] w_n2252_1;
	wire[2:0] w_n2252_2;
	wire[2:0] w_n2252_3;
	wire[2:0] w_n2252_4;
	wire[2:0] w_n2252_5;
	wire[2:0] w_n2252_6;
	wire[2:0] w_n2252_7;
	wire[1:0] w_n2255_0;
	wire[2:0] w_n2256_0;
	wire[2:0] w_n2256_1;
	wire[2:0] w_n2256_2;
	wire[2:0] w_n2256_3;
	wire[2:0] w_n2256_4;
	wire[2:0] w_n2256_5;
	wire[1:0] w_n2258_0;
	wire[1:0] w_n2260_0;
	wire[1:0] w_n2263_0;
	wire[2:0] w_n2277_0;
	wire[1:0] w_n2278_0;
	wire[1:0] w_n2280_0;
	wire[1:0] w_n2283_0;
	wire[1:0] w_n2286_0;
	wire[1:0] w_n2289_0;
	wire[1:0] w_n2297_0;
	wire[1:0] w_n2299_0;
	wire[1:0] w_n2301_0;
	wire[1:0] w_n2302_0;
	wire[1:0] w_n2305_0;
	wire[1:0] w_n2306_0;
	wire[1:0] w_n2309_0;
	wire[1:0] w_n2310_0;
	wire[1:0] w_n2311_0;
	wire[1:0] w_n2312_0;
	wire[1:0] w_n2315_0;
	wire[1:0] w_n2318_0;
	wire[1:0] w_n2326_0;
	wire[1:0] w_n2334_0;
	wire[1:0] w_n2342_0;
	wire[1:0] w_n2343_0;
	wire[1:0] w_n2344_0;
	wire[1:0] w_n2345_0;
	wire[1:0] w_n2346_0;
	wire[1:0] w_n2347_0;
	wire[2:0] w_n2348_0;
	wire[1:0] w_n2348_1;
	wire[2:0] w_n2349_0;
	wire[2:0] w_n2350_0;
	wire[2:0] w_n2351_0;
	wire[2:0] w_n2351_1;
	wire[2:0] w_n2351_2;
	wire[2:0] w_n2351_3;
	wire[2:0] w_n2351_4;
	wire[2:0] w_n2351_5;
	wire[2:0] w_n2351_6;
	wire[2:0] w_n2351_7;
	wire[1:0] w_n2351_8;
	wire[2:0] w_n2352_0;
	wire[2:0] w_n2353_0;
	wire[2:0] w_n2353_1;
	wire[2:0] w_n2355_0;
	wire[2:0] w_n2355_1;
	wire[2:0] w_n2355_2;
	wire[2:0] w_n2355_3;
	wire[2:0] w_n2355_4;
	wire[2:0] w_n2355_5;
	wire[2:0] w_n2355_6;
	wire[1:0] w_n2355_7;
	wire[2:0] w_n2357_0;
	wire[2:0] w_n2357_1;
	wire[2:0] w_n2357_2;
	wire[2:0] w_n2357_3;
	wire[2:0] w_n2357_4;
	wire[2:0] w_n2357_5;
	wire[2:0] w_n2357_6;
	wire[2:0] w_n2357_7;
	wire[2:0] w_n2359_0;
	wire[2:0] w_n2359_1;
	wire[2:0] w_n2359_2;
	wire[2:0] w_n2359_3;
	wire[2:0] w_n2359_4;
	wire[2:0] w_n2359_5;
	wire[2:0] w_n2359_6;
	wire[2:0] w_n2359_7;
	wire[1:0] w_n2364_0;
	wire[1:0] w_n2366_0;
	wire[1:0] w_n2370_0;
	wire[1:0] w_n2372_0;
	wire[1:0] w_n2375_0;
	wire[1:0] w_n2377_0;
	wire[1:0] w_n2384_0;
	wire[1:0] w_n2386_0;
	wire[1:0] w_n2394_0;
	wire[2:0] w_n2395_0;
	wire[1:0] w_n2402_0;
	wire[1:0] w_n2409_0;
	wire[2:0] w_n2412_0;
	wire[1:0] w_n2413_0;
	wire[1:0] w_n2415_0;
	wire[1:0] w_n2418_0;
	wire[1:0] w_n2421_0;
	wire[1:0] w_n2424_0;
	wire[1:0] w_n2425_0;
	wire[1:0] w_n2426_0;
	wire[1:0] w_n2434_0;
	wire[1:0] w_n2442_0;
	wire[1:0] w_n2443_0;
	wire[1:0] w_n2444_0;
	wire[1:0] w_n2447_0;
	wire[1:0] w_n2455_0;
	wire[2:0] w_n2456_0;
	wire[1:0] w_n2457_0;
	wire[1:0] w_n2462_0;
	wire[1:0] w_n2463_0;
	wire[1:0] w_n2464_0;
	wire[1:0] w_n2465_0;
	wire[1:0] w_n2466_0;
	wire[1:0] w_n2467_0;
	wire[2:0] w_n2468_0;
	wire[1:0] w_n2468_1;
	wire[2:0] w_n2469_0;
	wire[2:0] w_n2470_0;
	wire[2:0] w_n2471_0;
	wire[2:0] w_n2471_1;
	wire[2:0] w_n2471_2;
	wire[2:0] w_n2471_3;
	wire[2:0] w_n2471_4;
	wire[2:0] w_n2471_5;
	wire[2:0] w_n2471_6;
	wire[1:0] w_n2471_7;
	wire[2:0] w_n2472_0;
	wire[2:0] w_n2473_0;
	wire[1:0] w_n2473_1;
	wire[1:0] w_n2482_0;
	wire[2:0] w_n2483_0;
	wire[1:0] w_n2483_1;
	wire[2:0] w_n2484_0;
	wire[2:0] w_n2484_1;
	wire[1:0] w_n2486_0;
	wire[2:0] w_n2488_0;
	wire[2:0] w_n2488_1;
	wire[2:0] w_n2488_2;
	wire[2:0] w_n2488_3;
	wire[2:0] w_n2491_0;
	wire[2:0] w_n2491_1;
	wire[2:0] w_n2491_2;
	wire[2:0] w_n2491_3;
	wire[1:0] w_n2494_0;
	wire[1:0] w_n2495_0;
	wire[1:0] w_n2497_0;
	wire[1:0] w_n2498_0;
	wire[1:0] w_n2500_0;
	wire[2:0] w_n2501_0;
	wire[2:0] w_n2502_0;
	wire[1:0] w_n2503_0;
	wire[1:0] w_n2504_0;
	wire[2:0] w_n2505_0;
	wire[1:0] w_n2505_1;
	wire[2:0] w_n2506_0;
	wire[2:0] w_n2506_1;
	wire[2:0] w_n2506_2;
	wire[2:0] w_n2506_3;
	wire[2:0] w_n2506_4;
	wire[2:0] w_n2506_5;
	wire[2:0] w_n2506_6;
	wire[2:0] w_n2506_7;
	wire[1:0] w_n2508_0;
	wire[1:0] w_n2510_0;
	wire[2:0] w_n2513_0;
	wire[1:0] w_n2513_1;
	wire[2:0] w_n2519_0;
	wire[1:0] w_n2520_0;
	wire[1:0] w_n2521_0;
	wire[1:0] w_n2528_0;
	wire[1:0] w_n2531_0;
	wire[1:0] w_n2534_0;
	wire[1:0] w_n2537_0;
	wire[1:0] w_n2540_0;
	wire[1:0] w_n2543_0;
	wire[1:0] w_n2551_0;
	wire[1:0] w_n2559_0;
	wire[1:0] w_n2567_0;
	wire[1:0] w_n2568_0;
	wire[1:0] w_n2569_0;
	wire[1:0] w_n2570_0;
	wire[1:0] w_n2573_0;
	wire[1:0] w_n2576_0;
	wire[1:0] w_n2577_0;
	wire[1:0] w_n2578_0;
	wire[1:0] w_n2579_0;
	wire[1:0] w_n2580_0;
	wire[1:0] w_n2581_0;
	wire[1:0] w_n2582_0;
	wire[2:0] w_n2583_0;
	wire[1:0] w_n2583_1;
	wire[1:0] w_n2586_0;
	wire[1:0] w_n2594_0;
	wire[1:0] w_n2596_0;
	wire[1:0] w_n2598_0;
	wire[1:0] w_n2600_0;
	wire[2:0] w_n2601_0;
	wire[2:0] w_n2602_0;
	wire[1:0] w_n2604_0;
	wire[1:0] w_n2606_0;
	wire[1:0] w_n2613_0;
	wire[1:0] w_n2617_0;
	wire[1:0] w_n2618_0;
	wire[2:0] w_n2623_0;
	wire[1:0] w_n2628_0;
	wire[1:0] w_n2631_0;
	wire[2:0] w_n2636_0;
	wire[1:0] w_n2637_0;
	wire[1:0] w_n2639_0;
	wire[1:0] w_n2642_0;
	wire[1:0] w_n2645_0;
	wire[1:0] w_n2653_0;
	wire[2:0] w_n2654_0;
	wire[1:0] w_n2655_0;
	wire[1:0] w_n2659_0;
	wire[1:0] w_n2660_0;
	wire[1:0] w_n2661_0;
	wire[1:0] w_n2662_0;
	wire[1:0] w_n2665_0;
	wire[1:0] w_n2673_0;
	wire[1:0] w_n2676_0;
	wire[1:0] w_n2677_0;
	wire[1:0] w_n2678_0;
	wire[1:0] w_n2679_0;
	wire[2:0] w_n2680_0;
	wire[1:0] w_n2680_1;
	wire[2:0] w_n2681_0;
	wire[2:0] w_n2682_0;
	wire[2:0] w_n2683_0;
	wire[2:0] w_n2683_1;
	wire[1:0] w_n2683_2;
	wire[2:0] w_n2684_0;
	wire[2:0] w_n2684_1;
	wire[2:0] w_n2684_2;
	wire[1:0] w_n2684_3;
	wire[1:0] w_n2685_0;
	wire[2:0] w_n2687_0;
	wire[2:0] w_n2687_1;
	wire[2:0] w_n2687_2;
	wire[1:0] w_n2687_3;
	wire[1:0] w_n2688_0;
	wire[2:0] w_n2690_0;
	wire[2:0] w_n2690_1;
	wire[2:0] w_n2690_2;
	wire[1:0] w_n2691_0;
	wire[1:0] w_n2695_0;
	wire[1:0] w_n2698_0;
	wire[1:0] w_n2703_0;
	wire[1:0] w_n2706_0;
	wire[2:0] w_n2707_0;
	wire[2:0] w_n2707_1;
	wire[2:0] w_n2707_2;
	wire[2:0] w_n2707_3;
	wire[2:0] w_n2707_4;
	wire[2:0] w_n2707_5;
	wire[2:0] w_n2707_6;
	wire[1:0] w_n2707_7;
	wire[1:0] w_n2710_0;
	wire[1:0] w_n2712_0;
	wire[1:0] w_n2715_0;
	wire[2:0] w_n2717_0;
	wire[1:0] w_n2725_0;
	wire[1:0] w_n2729_0;
	wire[1:0] w_n2732_0;
	wire[2:0] w_n2738_0;
	wire[2:0] w_n2743_0;
	wire[1:0] w_n2744_0;
	wire[1:0] w_n2751_0;
	wire[2:0] w_n2759_0;
	wire[1:0] w_n2760_0;
	wire[1:0] w_n2762_0;
	wire[1:0] w_n2765_0;
	wire[1:0] w_n2768_0;
	wire[1:0] w_n2769_0;
	wire[1:0] w_n2770_0;
	wire[1:0] w_n2771_0;
	wire[1:0] w_n2772_0;
	wire[1:0] w_n2773_0;
	wire[1:0] w_n2777_0;
	wire[1:0] w_n2785_0;
	wire[1:0] w_n2793_0;
	wire[1:0] w_n2794_0;
	wire[1:0] w_n2795_0;
	wire[1:0] w_n2796_0;
	wire[2:0] w_n2797_0;
	wire[1:0] w_n2797_1;
	wire[2:0] w_n2798_0;
	wire[2:0] w_n2799_0;
	wire[2:0] w_n2800_0;
	wire[2:0] w_n2800_1;
	wire[2:0] w_n2800_2;
	wire[2:0] w_n2800_3;
	wire[2:0] w_n2800_4;
	wire[2:0] w_n2800_5;
	wire[2:0] w_n2800_6;
	wire[1:0] w_n2800_7;
	wire[1:0] w_n2801_0;
	wire[2:0] w_n2802_0;
	wire[2:0] w_n2802_1;
	wire[1:0] w_n2804_0;
	wire[2:0] w_n2806_0;
	wire[2:0] w_n2807_0;
	wire[2:0] w_n2807_1;
	wire[2:0] w_n2807_2;
	wire[2:0] w_n2807_3;
	wire[2:0] w_n2807_4;
	wire[2:0] w_n2807_5;
	wire[2:0] w_n2807_6;
	wire[2:0] w_n2807_7;
	wire[2:0] w_n2809_0;
	wire[2:0] w_n2810_0;
	wire[2:0] w_n2810_1;
	wire[2:0] w_n2810_2;
	wire[2:0] w_n2810_3;
	wire[2:0] w_n2810_4;
	wire[2:0] w_n2810_5;
	wire[2:0] w_n2810_6;
	wire[1:0] w_n2810_7;
	wire[2:0] w_n2813_0;
	wire[2:0] w_n2813_1;
	wire[2:0] w_n2813_2;
	wire[2:0] w_n2813_3;
	wire[2:0] w_n2813_4;
	wire[2:0] w_n2813_5;
	wire[2:0] w_n2813_6;
	wire[2:0] w_n2815_0;
	wire[2:0] w_n2816_0;
	wire[2:0] w_n2816_1;
	wire[2:0] w_n2816_2;
	wire[2:0] w_n2816_3;
	wire[2:0] w_n2816_4;
	wire[2:0] w_n2816_5;
	wire[2:0] w_n2816_6;
	wire[2:0] w_n2816_7;
	wire[1:0] w_n2820_0;
	wire[1:0] w_n2823_0;
	wire[1:0] w_n2824_0;
	wire[2:0] w_n2825_0;
	wire[2:0] w_n2825_1;
	wire[1:0] w_n2833_0;
	wire[1:0] w_n2835_0;
	wire[2:0] w_n2836_0;
	wire[2:0] w_n2836_1;
	wire[1:0] w_n2845_0;
	wire[1:0] w_n2847_0;
	wire[1:0] w_n2857_0;
	wire[1:0] w_n2859_0;
	wire[1:0] w_n2865_0;
	wire[2:0] w_n2867_0;
	wire[1:0] w_n2867_1;
	wire[1:0] w_n2870_0;
	wire[1:0] w_n2878_0;
	wire[1:0] w_n2879_0;
	wire[1:0] w_n2881_0;
	wire[1:0] w_n2889_0;
	wire[1:0] w_n2891_0;
	wire[1:0] w_n2892_0;
	wire[1:0] w_n2894_0;
	wire[1:0] w_n2895_0;
	wire[1:0] w_n2897_0;
	wire[1:0] w_n2898_0;
	wire[1:0] w_n2902_0;
	wire[1:0] w_n2903_0;
	wire[1:0] w_n2906_0;
	wire[1:0] w_n2909_0;
	wire[1:0] w_n2918_0;
	wire[2:0] w_n2923_0;
	wire[2:0] w_n2923_1;
	wire[2:0] w_n2923_2;
	wire[2:0] w_n2923_3;
	wire[1:0] w_n2927_0;
	wire[1:0] w_n2929_0;
	wire[1:0] w_n2931_0;
	wire[1:0] w_n2932_0;
	wire[1:0] w_n2934_0;
	wire[1:0] w_n2938_0;
	wire[1:0] w_n2942_0;
	wire[2:0] w_n2943_0;
	wire[2:0] w_n2943_1;
	wire[1:0] w_n2943_2;
	wire[1:0] w_n2944_0;
	wire[1:0] w_n2948_0;
	wire[1:0] w_n2950_0;
	wire[1:0] w_n2953_0;
	wire[1:0] w_n2954_0;
	wire[1:0] w_n2964_0;
	wire[1:0] w_n2968_0;
	wire[1:0] w_n2971_0;
	wire[2:0] w_n2973_0;
	wire[1:0] w_n2974_0;
	wire[1:0] w_n2976_0;
	wire[1:0] w_n2979_0;
	wire[1:0] w_n2987_0;
	wire[2:0] w_n2988_0;
	wire[1:0] w_n2990_0;
	wire[1:0] w_n2994_0;
	wire[1:0] w_n2995_0;
	wire[1:0] w_n2996_0;
	wire[1:0] w_n2999_0;
	wire[1:0] w_n3002_0;
	wire[1:0] w_n3003_0;
	wire[1:0] w_n3004_0;
	wire[2:0] w_n3005_0;
	wire[1:0] w_n3005_1;
	wire[2:0] w_n3006_0;
	wire[2:0] w_n3007_0;
	wire[2:0] w_n3008_0;
	wire[2:0] w_n3008_1;
	wire[2:0] w_n3008_2;
	wire[2:0] w_n3008_3;
	wire[2:0] w_n3008_4;
	wire[2:0] w_n3008_5;
	wire[2:0] w_n3008_6;
	wire[2:0] w_n3008_7;
	wire[1:0] w_n3009_0;
	wire[2:0] w_n3010_0;
	wire[2:0] w_n3010_1;
	wire[1:0] w_n3018_0;
	wire[1:0] w_n3019_0;
	wire[1:0] w_n3020_0;
	wire[1:0] w_n3021_0;
	wire[2:0] w_n3023_0;
	wire[2:0] w_n3023_1;
	wire[2:0] w_n3023_2;
	wire[2:0] w_n3023_3;
	wire[2:0] w_n3023_4;
	wire[2:0] w_n3023_5;
	wire[2:0] w_n3023_6;
	wire[2:0] w_n3023_7;
	wire[2:0] w_n3023_8;
	wire[2:0] w_n3023_9;
	wire[2:0] w_n3023_10;
	wire[2:0] w_n3024_0;
	wire[2:0] w_n3025_0;
	wire[1:0] w_n3026_0;
	wire[1:0] w_n3027_0;
	wire[2:0] w_n3028_0;
	wire[1:0] w_n3028_1;
	wire[2:0] w_n3029_0;
	wire[2:0] w_n3029_1;
	wire[2:0] w_n3029_2;
	wire[2:0] w_n3029_3;
	wire[2:0] w_n3029_4;
	wire[2:0] w_n3029_5;
	wire[2:0] w_n3029_6;
	wire[2:0] w_n3029_7;
	wire[2:0] w_n3042_0;
	wire[1:0] w_n3043_0;
	wire[1:0] w_n3044_0;
	wire[1:0] w_n3050_0;
	wire[1:0] w_n3053_0;
	wire[1:0] w_n3059_0;
	wire[1:0] w_n3065_0;
	wire[1:0] w_n3069_0;
	wire[1:0] w_n3070_0;
	wire[1:0] w_n3071_0;
	wire[1:0] w_n3072_0;
	wire[1:0] w_n3073_0;
	wire[1:0] w_n3074_0;
	wire[1:0] w_n3075_0;
	wire[2:0] w_n3076_0;
	wire[1:0] w_n3079_0;
	wire[1:0] w_n3085_0;
	wire[1:0] w_n3087_0;
	wire[1:0] w_n3089_0;
	wire[2:0] w_n3090_0;
	wire[2:0] w_n3091_0;
	wire[1:0] w_n3093_0;
	wire[1:0] w_n3098_0;
	wire[1:0] w_n3106_0;
	wire[2:0] w_n3118_0;
	wire[2:0] w_n3121_0;
	wire[1:0] w_n3126_0;
	wire[1:0] w_n3130_0;
	wire[1:0] w_n3131_0;
	wire[1:0] w_n3132_0;
	wire[1:0] w_n3136_0;
	wire[1:0] w_n3138_0;
	wire[1:0] w_n3139_0;
	wire[2:0] w_n3140_0;
	wire[2:0] w_n3141_0;
	wire[2:0] w_n3142_0;
	wire[2:0] w_n3143_0;
	wire[1:0] w_n3143_1;
	wire[2:0] w_n3144_0;
	wire[2:0] w_n3144_1;
	wire[1:0] w_n3145_0;
	wire[2:0] w_n3147_0;
	wire[2:0] w_n3147_1;
	wire[1:0] w_n3148_0;
	wire[1:0] w_n3150_0;
	wire[1:0] w_n3154_0;
	wire[1:0] w_n3157_0;
	wire[1:0] w_n3162_0;
	wire[1:0] w_n3165_0;
	wire[2:0] w_n3166_0;
	wire[2:0] w_n3166_1;
	wire[2:0] w_n3166_2;
	wire[2:0] w_n3166_3;
	wire[2:0] w_n3166_4;
	wire[2:0] w_n3166_5;
	wire[2:0] w_n3166_6;
	wire[2:0] w_n3166_7;
	wire[2:0] w_n3166_8;
	wire[1:0] w_n3169_0;
	wire[1:0] w_n3171_0;
	wire[1:0] w_n3174_0;
	wire[1:0] w_n3177_0;
	wire[2:0] w_n3179_0;
	wire[1:0] w_n3185_0;
	wire[2:0] w_n3190_0;
	wire[2:0] w_n3191_0;
	wire[1:0] w_n3194_0;
	wire[1:0] w_n3200_0;
	wire[2:0] w_n3201_0;
	wire[1:0] w_n3202_0;
	wire[2:0] w_n3203_0;
	wire[2:0] w_n3203_1;
	wire[2:0] w_n3203_2;
	wire[2:0] w_n3203_3;
	wire[2:0] w_n3203_4;
	wire[2:0] w_n3203_5;
	wire[2:0] w_n3203_6;
	wire[2:0] w_n3203_7;
	wire[1:0] w_n3203_8;
	wire[1:0] w_n3204_0;
	wire[2:0] w_n3205_0;
	wire[2:0] w_n3205_1;
	wire[1:0] w_n3207_0;
	wire[2:0] w_n3209_0;
	wire[2:0] w_n3210_0;
	wire[2:0] w_n3210_1;
	wire[2:0] w_n3210_2;
	wire[2:0] w_n3210_3;
	wire[2:0] w_n3210_4;
	wire[2:0] w_n3210_5;
	wire[2:0] w_n3210_6;
	wire[2:0] w_n3210_7;
	wire[2:0] w_n3212_0;
	wire[2:0] w_n3213_0;
	wire[2:0] w_n3213_1;
	wire[2:0] w_n3213_2;
	wire[2:0] w_n3213_3;
	wire[2:0] w_n3213_4;
	wire[2:0] w_n3213_5;
	wire[2:0] w_n3213_6;
	wire[1:0] w_n3213_7;
	wire[2:0] w_n3216_0;
	wire[2:0] w_n3216_1;
	wire[2:0] w_n3216_2;
	wire[2:0] w_n3216_3;
	wire[2:0] w_n3216_4;
	wire[2:0] w_n3216_5;
	wire[2:0] w_n3216_6;
	wire[2:0] w_n3216_7;
	wire[2:0] w_n3218_0;
	wire[2:0] w_n3219_0;
	wire[2:0] w_n3219_1;
	wire[2:0] w_n3219_2;
	wire[2:0] w_n3219_3;
	wire[2:0] w_n3219_4;
	wire[2:0] w_n3219_5;
	wire[2:0] w_n3219_6;
	wire[2:0] w_n3219_7;
	wire[1:0] w_n3223_0;
	wire[1:0] w_n3227_0;
	wire[1:0] w_n3228_0;
	wire[2:0] w_n3229_0;
	wire[2:0] w_n3229_1;
	wire[1:0] w_n3237_0;
	wire[1:0] w_n3240_0;
	wire[1:0] w_n3241_0;
	wire[2:0] w_n3242_0;
	wire[2:0] w_n3242_1;
	wire[1:0] w_n3250_0;
	wire[1:0] w_n3252_0;
	wire[1:0] w_n3260_0;
	wire[1:0] w_n3262_0;
	wire[1:0] w_n3270_0;
	wire[1:0] w_n3272_0;
	wire[1:0] w_n3280_0;
	wire[1:0] w_n3289_0;
	wire[1:0] w_n3292_0;
	wire[1:0] w_n3301_0;
	wire[1:0] w_n3304_0;
	wire[1:0] w_n3311_0;
	wire[2:0] w_n3312_0;
	wire[1:0] w_n3315_0;
	wire[1:0] w_n3323_0;
	wire[1:0] w_n3324_0;
	wire[1:0] w_n3326_0;
	wire[1:0] w_n3334_0;
	wire[1:0] w_n3337_0;
	wire[1:0] w_n3338_0;
	wire[1:0] w_n3341_0;
	wire[1:0] w_n3343_0;
	wire[1:0] w_n3345_0;
	wire[1:0] w_n3346_0;
	wire[1:0] w_n3348_0;
	wire[1:0] w_n3349_0;
	wire[1:0] w_n3351_0;
	wire[1:0] w_n3352_0;
	wire[1:0] w_n3354_0;
	wire[1:0] w_n3355_0;
	wire[1:0] w_n3357_0;
	wire[1:0] w_n3358_0;
	wire[1:0] w_n3360_0;
	wire[1:0] w_n3361_0;
	wire[1:0] w_n3363_0;
	wire[1:0] w_n3368_0;
	wire[1:0] w_n3371_0;
	wire[1:0] w_n3380_0;
	wire[1:0] w_n3381_0;
	wire[1:0] w_n3382_0;
	wire[2:0] w_n3384_0;
	wire[2:0] w_n3384_1;
	wire[2:0] w_n3384_2;
	wire[2:0] w_n3384_3;
	wire[2:0] w_n3384_4;
	wire[2:0] w_n3384_5;
	wire[2:0] w_n3384_6;
	wire[1:0] w_n3384_7;
	wire[2:0] w_n3386_0;
	wire[2:0] w_n3386_1;
	wire[2:0] w_n3386_2;
	wire[2:0] w_n3386_3;
	wire[1:0] w_n3386_4;
	wire[2:0] w_n3388_0;
	wire[2:0] w_n3388_1;
	wire[2:0] w_n3388_2;
	wire[2:0] w_n3388_3;
	wire[2:0] w_n3388_4;
	wire[2:0] w_n3390_0;
	wire[2:0] w_n3390_1;
	wire[2:0] w_n3390_2;
	wire[2:0] w_n3390_3;
	wire[2:0] w_n3390_4;
	wire[1:0] w_n3395_0;
	wire[1:0] w_n3396_0;
	wire[1:0] w_n3397_0;
	wire[1:0] w_n3399_0;
	wire[1:0] w_n3407_0;
	wire[1:0] w_n3408_0;
	wire[1:0] w_n3409_0;
	wire[1:0] w_n3414_0;
	wire[2:0] w_n3415_0;
	wire[1:0] w_n3415_1;
	wire[1:0] w_n3416_0;
	wire[1:0] w_n3418_0;
	wire[1:0] w_n3420_0;
	wire[1:0] w_n3429_0;
	wire[2:0] w_n3435_0;
	wire[1:0] w_n3440_0;
	wire[2:0] w_n3441_0;
	wire[2:0] w_n3441_1;
	wire[2:0] w_n3441_2;
	wire[2:0] w_n3441_3;
	wire[2:0] w_n3441_4;
	wire[2:0] w_n3441_5;
	wire[2:0] w_n3441_6;
	wire[2:0] w_n3441_7;
	wire[1:0] w_n3442_0;
	wire[2:0] w_n3443_0;
	wire[2:0] w_n3443_1;
	wire[1:0] w_n3451_0;
	wire[1:0] w_n3452_0;
	wire[1:0] w_n3454_0;
	wire[2:0] w_n3455_0;
	wire[2:0] w_n3455_1;
	wire[2:0] w_n3455_2;
	wire[2:0] w_n3455_3;
	wire[2:0] w_n3455_4;
	wire[2:0] w_n3456_0;
	wire[1:0] w_n3459_0;
	wire[2:0] w_n3460_0;
	wire[2:0] w_n3461_0;
	wire[2:0] w_n3461_1;
	wire[2:0] w_n3461_2;
	wire[2:0] w_n3461_3;
	wire[2:0] w_n3461_4;
	wire[2:0] w_n3461_5;
	wire[2:0] w_n3461_6;
	wire[2:0] w_n3461_7;
	wire[2:0] w_n3461_8;
	wire[1:0] w_n3463_0;
	wire[2:0] w_n3468_0;
	wire[2:0] w_n3470_0;
	wire[2:0] w_n3481_0;
	wire[1:0] w_n3488_0;
	wire[1:0] w_n3489_0;
	wire[2:0] w_n3494_0;
	wire[2:0] w_n3495_0;
	wire[2:0] w_n3495_1;
	wire[2:0] w_n3495_2;
	wire[2:0] w_n3495_3;
	wire[2:0] w_n3495_4;
	wire[2:0] w_n3495_5;
	wire[2:0] w_n3495_6;
	wire[2:0] w_n3495_7;
	wire[1:0] w_n3495_8;
	wire[1:0] w_n3496_0;
	wire[2:0] w_n3497_0;
	wire[2:0] w_n3509_0;
	wire[2:0] w_n3510_0;
	wire[2:0] w_n3510_1;
	wire[2:0] w_n3510_2;
	wire[2:0] w_n3510_3;
	wire[2:0] w_n3510_4;
	wire[2:0] w_n3510_5;
	wire[2:0] w_n3510_6;
	wire[2:0] w_n3510_7;
	wire[2:0] w_n3510_8;
	wire[2:0] w_n3511_0;
	wire[1:0] w_n3512_0;
	wire[2:0] w_n3513_0;
	wire[2:0] w_n3513_1;
	wire[1:0] w_n3514_0;
	wire[1:0] w_n3518_0;
	wire[1:0] w_n3519_0;
	wire[2:0] w_n3520_0;
	wire[1:0] w_n3521_0;
	wire[1:0] w_n3522_0;
	wire[1:0] w_n3526_0;
	wire[2:0] w_n3529_0;
	wire[1:0] w_n3532_0;
	wire[2:0] w_n3537_0;
	wire[2:0] w_n3537_1;
	wire[2:0] w_n3543_0;
	wire[1:0] w_n3546_0;
	wire[2:0] w_n3547_0;
	wire[2:0] w_n3547_1;
	wire[2:0] w_n3547_2;
	wire[2:0] w_n3547_3;
	wire[2:0] w_n3547_4;
	wire[2:0] w_n3547_5;
	wire[2:0] w_n3547_6;
	wire[2:0] w_n3547_7;
	wire[2:0] w_n3548_0;
	wire[2:0] w_n3549_0;
	wire[2:0] w_n3550_0;
	wire[2:0] w_n3550_1;
	wire[2:0] w_n3552_0;
	wire[2:0] w_n3552_1;
	wire[2:0] w_n3552_2;
	wire[2:0] w_n3552_3;
	wire[2:0] w_n3552_4;
	wire[2:0] w_n3552_5;
	wire[2:0] w_n3552_6;
	wire[2:0] w_n3552_7;
	wire[2:0] w_n3554_0;
	wire[2:0] w_n3554_1;
	wire[2:0] w_n3554_2;
	wire[2:0] w_n3554_3;
	wire[2:0] w_n3554_4;
	wire[2:0] w_n3554_5;
	wire[2:0] w_n3554_6;
	wire[2:0] w_n3554_7;
	wire[1:0] w_n3554_8;
	wire[2:0] w_n3557_0;
	wire[1:0] w_n3557_1;
	wire[2:0] w_n3558_0;
	wire[2:0] w_n3558_1;
	wire[2:0] w_n3558_2;
	wire[2:0] w_n3558_3;
	wire[2:0] w_n3558_4;
	wire[2:0] w_n3558_5;
	wire[2:0] w_n3558_6;
	wire[1:0] w_n3562_0;
	wire[1:0] w_n3563_0;
	wire[1:0] w_n3565_0;
	wire[2:0] w_n3566_0;
	wire[2:0] w_n3566_1;
	wire[1:0] w_n3574_0;
	wire[1:0] w_n3575_0;
	wire[1:0] w_n3576_0;
	wire[1:0] w_n3577_0;
	wire[1:0] w_n3578_0;
	wire[2:0] w_n3579_0;
	wire[2:0] w_n3579_1;
	wire[1:0] w_n3587_0;
	wire[1:0] w_n3588_0;
	wire[1:0] w_n3589_0;
	wire[1:0] w_n3590_0;
	wire[1:0] w_n3598_0;
	wire[1:0] w_n3599_0;
	wire[1:0] w_n3600_0;
	wire[1:0] w_n3601_0;
	wire[1:0] w_n3609_0;
	wire[1:0] w_n3610_0;
	wire[1:0] w_n3611_0;
	wire[1:0] w_n3612_0;
	wire[1:0] w_n3620_0;
	wire[1:0] w_n3621_0;
	wire[1:0] w_n3622_0;
	wire[1:0] w_n3623_0;
	wire[1:0] w_n3631_0;
	wire[1:0] w_n3632_0;
	wire[1:0] w_n3633_0;
	wire[1:0] w_n3634_0;
	wire[1:0] w_n3642_0;
	wire[1:0] w_n3643_0;
	wire[1:0] w_n3644_0;
	wire[1:0] w_n3645_0;
	wire[1:0] w_n3653_0;
	wire[1:0] w_n3654_0;
	wire[1:0] w_n3655_0;
	wire[1:0] w_n3656_0;
	wire[1:0] w_n3664_0;
	wire[1:0] w_n3665_0;
	wire[1:0] w_n3676_0;
	wire[1:0] w_n3678_0;
	wire[1:0] w_n3681_0;
	wire[1:0] w_n3682_0;
	wire[1:0] w_n3685_0;
	wire[1:0] w_n3686_0;
	wire[1:0] w_n3688_0;
	wire[1:0] w_n3695_0;
	wire[1:0] w_n3698_0;
	wire[1:0] w_n3700_0;
	wire[1:0] w_n3701_0;
	wire[1:0] w_n3702_0;
	wire[1:0] w_n3705_0;
	wire[1:0] w_n3709_0;
	wire[1:0] w_n3713_0;
	wire[1:0] w_n3714_0;
	wire[1:0] w_n3718_0;
	wire[1:0] w_n3720_0;
	wire[1:0] w_n3725_0;
	wire[2:0] w_n3733_0;
	wire[1:0] w_n3734_0;
	wire[1:0] w_n3738_0;
	wire[1:0] w_n3742_0;
	wire[1:0] w_n3760_0;
	wire[2:0] w_n3761_0;
	wire[1:0] w_n3763_0;
	wire[1:0] w_n3766_0;
	wire[1:0] w_n3770_0;
	wire[1:0] w_n3773_0;
	wire[1:0] w_n3780_0;
	wire[1:0] w_n3787_0;
	wire[1:0] w_n3789_0;
	wire[1:0] w_n3790_0;
	wire[1:0] w_n3798_0;
	wire[1:0] w_n3799_0;
	wire[1:0] w_n3801_0;
	wire[1:0] w_n3809_0;
	wire[1:0] w_n3810_0;
	wire[1:0] w_n3811_0;
	wire[1:0] w_n3819_0;
	wire[1:0] w_n3820_0;
	wire[1:0] w_n3821_0;
	wire[1:0] w_n3824_0;
	wire[2:0] w_n3825_0;
	wire[1:0] w_n3826_0;
	wire[2:0] w_n3833_0;
	wire[1:0] w_n3836_0;
	wire[2:0] w_n3837_0;
	wire[2:0] w_n3837_1;
	wire[2:0] w_n3837_2;
	wire[2:0] w_n3837_3;
	wire[2:0] w_n3837_4;
	wire[2:0] w_n3837_5;
	wire[2:0] w_n3837_6;
	wire[2:0] w_n3837_7;
	wire[1:0] w_n3837_8;
	wire[2:0] w_n3838_0;
	wire[1:0] w_n3838_1;
	wire[1:0] w_n3839_0;
	wire[1:0] w_n3840_0;
	wire[2:0] w_n3841_0;
	wire[2:0] w_n3842_0;
	wire[2:0] w_n3842_1;
	wire[1:0] w_n3850_0;
	wire[2:0] w_n3851_0;
	wire[2:0] w_n3852_0;
	wire[1:0] w_n3853_0;
	wire[1:0] w_n3854_0;
	wire[1:0] w_n3868_0;
	wire[1:0] w_n3871_0;
	wire[1:0] w_n3875_0;
	wire[1:0] w_n3881_0;
	wire[1:0] w_n3887_0;
	wire[2:0] w_n3892_0;
	wire[1:0] w_n3895_0;
	wire[1:0] w_n3910_0;
	wire[1:0] w_n3959_0;
	wire[1:0] w_n3961_0;
	wire[1:0] w_n3963_0;
	wire[1:0] w_n3968_0;
	wire[1:0] w_n3969_0;
	wire[1:0] w_n3971_0;
	wire[1:0] w_n3972_0;
	wire[1:0] w_n3982_0;
	wire[1:0] w_n3985_0;
	wire[1:0] w_n3989_0;
	wire[1:0] w_n3992_0;
	wire[1:0] w_n3998_0;
	wire[1:0] w_n4006_0;
	wire[1:0] w_n4008_0;
	wire[1:0] w_n4009_0;
	wire[1:0] w_n4017_0;
	wire[1:0] w_n4018_0;
	wire[1:0] w_n4020_0;
	wire[1:0] w_n4028_0;
	wire[1:0] w_n4029_0;
	wire[1:0] w_n4030_0;
	wire[1:0] w_n4038_0;
	wire[1:0] w_n4039_0;
	wire[1:0] w_n4040_0;
	wire[1:0] w_n4043_0;
	wire[1:0] w_n4051_0;
	wire[2:0] w_n4059_0;
	wire[1:0] w_n4062_0;
	wire[2:0] w_n4063_0;
	wire[2:0] w_n4063_1;
	wire[2:0] w_n4063_2;
	wire[2:0] w_n4063_3;
	wire[2:0] w_n4063_4;
	wire[2:0] w_n4063_5;
	wire[2:0] w_n4063_6;
	wire[2:0] w_n4063_7;
	wire[1:0] w_n4063_8;
	wire[2:0] w_n4064_0;
	wire[2:0] w_n4065_0;
	wire[2:0] w_n4066_0;
	wire[2:0] w_n4066_1;
	wire[1:0] w_n4074_0;
	wire[2:0] w_n4075_0;
	wire[1:0] w_n4075_1;
	wire[1:0] w_n4076_0;
	wire[2:0] w_n4088_0;
	wire[1:0] w_n4089_0;
	wire[1:0] w_n4090_0;
	wire[1:0] w_n4091_0;
	wire[2:0] w_n4093_0;
	wire[2:0] w_n4093_1;
	wire[2:0] w_n4093_2;
	wire[2:0] w_n4093_3;
	wire[2:0] w_n4093_4;
	wire[2:0] w_n4093_5;
	wire[2:0] w_n4093_6;
	wire[2:0] w_n4093_7;
	wire[2:0] w_n4093_8;
	wire[2:0] w_n4093_9;
	wire[2:0] w_n4093_10;
	wire[1:0] w_n4093_11;
	wire[1:0] w_n4094_0;
	wire[1:0] w_n4096_0;
	wire[1:0] w_n4097_0;
	wire[1:0] w_n4100_0;
	wire[1:0] w_n4101_0;
	wire[1:0] w_n4108_0;
	wire[1:0] w_n4112_0;
	wire[1:0] w_n4115_0;
	wire[1:0] w_n4120_0;
	wire[1:0] w_n4128_0;
	wire[1:0] w_n4130_0;
	wire[1:0] w_n4132_0;
	wire[1:0] w_n4140_0;
	wire[1:0] w_n4141_0;
	wire[1:0] w_n4143_0;
	wire[1:0] w_n4151_0;
	wire[1:0] w_n4152_0;
	wire[1:0] w_n4153_0;
	wire[1:0] w_n4161_0;
	wire[1:0] w_n4162_0;
	wire[1:0] w_n4163_0;
	wire[1:0] w_n4194_0;
	wire[1:0] w_n4203_0;
	wire[2:0] w_n4213_0;
	wire[2:0] w_n4213_1;
	wire[2:0] w_n4213_2;
	wire[2:0] w_n4213_3;
	wire[2:0] w_n4213_4;
	wire[2:0] w_n4213_5;
	wire[2:0] w_n4213_6;
	wire[2:0] w_n4214_0;
	wire[2:0] w_n4215_0;
	wire[2:0] w_n4215_1;
	wire[1:0] w_n4225_0;
	wire[2:0] w_n4226_0;
	wire[1:0] w_n4227_0;
	wire[2:0] w_n4237_0;
	wire[2:0] w_n4242_0;
	wire[1:0] w_n4243_0;
	wire[2:0] w_n4244_0;
	wire[1:0] w_n4245_0;
	wire[1:0] w_n4250_0;
	wire[1:0] w_n4251_0;
	wire[1:0] w_n4254_0;
	wire[1:0] w_n4266_0;
	wire[1:0] w_n4270_0;
	wire[1:0] w_n4271_0;
	wire[1:0] w_n4274_0;
	wire[1:0] w_n4276_0;
	wire[1:0] w_n4278_0;
	wire[1:0] w_n4281_0;
	wire[1:0] w_n4285_0;
	wire[1:0] w_n4290_0;
	wire[1:0] w_n4295_0;
	wire[1:0] w_n4303_0;
	wire[1:0] w_n4305_0;
	wire[1:0] w_n4307_0;
	wire[1:0] w_n4315_0;
	wire[1:0] w_n4316_0;
	wire[1:0] w_n4317_0;
	wire[1:0] w_n4325_0;
	wire[1:0] w_n4326_0;
	wire[1:0] w_n4327_0;
	wire[1:0] w_n4335_0;
	wire[1:0] w_n4336_0;
	wire[1:0] w_n4337_0;
	wire[2:0] w_n4338_0;
	wire[2:0] w_n4338_1;
	wire[2:0] w_n4343_0;
	wire[2:0] w_n4343_1;
	wire[1:0] w_n4343_2;
	wire[1:0] w_n4344_0;
	wire[2:0] w_n4349_0;
	wire[2:0] w_n4349_1;
	wire[1:0] w_n4355_0;
	wire[1:0] w_n4356_0;
	wire[2:0] w_n4357_0;
	wire[1:0] w_n4358_0;
	wire[1:0] w_n4359_0;
	wire[1:0] w_n4360_0;
	wire[1:0] w_n4361_0;
	wire[1:0] w_n4364_0;
	wire[1:0] w_n4366_0;
	wire[1:0] w_n4367_0;
	wire[1:0] w_n4369_0;
	wire[1:0] w_n4381_0;
	wire[1:0] w_n4382_0;
	wire[1:0] w_n4385_0;
	wire[1:0] w_n4388_0;
	wire[1:0] w_n4391_0;
	wire[1:0] w_n4396_0;
	wire[1:0] w_n4401_0;
	wire[1:0] w_n4409_0;
	wire[1:0] w_n4411_0;
	wire[1:0] w_n4413_0;
	wire[1:0] w_n4421_0;
	wire[1:0] w_n4422_0;
	wire[1:0] w_n4424_0;
	wire[1:0] w_n4432_0;
	wire[1:0] w_n4433_0;
	wire[1:0] w_n4434_0;
	wire[1:0] w_n4442_0;
	wire[1:0] w_n4443_0;
	wire[1:0] w_n4448_0;
	wire[1:0] w_n4449_0;
	wire[1:0] w_n4450_0;
	wire[2:0] w_n4451_0;
	wire[1:0] w_n4452_0;
	wire[1:0] w_n4453_0;
	wire[1:0] w_n4454_0;
	wire[1:0] w_n4456_0;
	wire[1:0] w_n4457_0;
	wire[1:0] w_n4459_0;
	wire[1:0] w_n4469_0;
	wire[1:0] w_n4470_0;
	wire[1:0] w_n4473_0;
	wire[1:0] w_n4480_0;
	wire[1:0] w_n4484_0;
	wire[1:0] w_n4489_0;
	wire[1:0] w_n4495_0;
	wire[1:0] w_n4496_0;
	wire[1:0] w_n4497_0;
	wire[1:0] w_n4505_0;
	wire[1:0] w_n4506_0;
	wire[1:0] w_n4508_0;
	wire[1:0] w_n4516_0;
	wire[1:0] w_n4517_0;
	wire[1:0] w_n4518_0;
	wire[1:0] w_n4526_0;
	wire[1:0] w_n4527_0;
	wire[1:0] w_n4528_0;
	wire[1:0] w_n4536_0;
	wire[1:0] w_n4537_0;
	wire[1:0] w_n4538_0;
	wire[2:0] w_n4539_0;
	wire[1:0] w_n4540_0;
	wire[1:0] w_n4541_0;
	wire[1:0] w_n4542_0;
	wire[1:0] w_n4543_0;
	wire[1:0] w_n4546_0;
	wire[1:0] w_n4547_0;
	wire[1:0] w_n4549_0;
	wire[1:0] w_n4556_0;
	wire[2:0] w_n4558_0;
	wire[1:0] w_n4563_0;
	wire[1:0] w_n4564_0;
	wire[1:0] w_n4567_0;
	wire[1:0] w_n4572_0;
	wire[1:0] w_n4575_0;
	wire[1:0] w_n4580_0;
	wire[1:0] w_n4583_0;
	wire[1:0] w_n4584_0;
	wire[1:0] w_n4585_0;
	wire[1:0] w_n4586_0;
	wire[1:0] w_n4594_0;
	wire[1:0] w_n4595_0;
	wire[1:0] w_n4603_0;
	wire[1:0] w_n4604_0;
	wire[1:0] w_n4606_0;
	wire[1:0] w_n4614_0;
	wire[1:0] w_n4615_0;
	wire[1:0] w_n4616_0;
	wire[1:0] w_n4622_0;
	wire[1:0] w_n4623_0;
	wire[1:0] w_n4624_0;
	wire[2:0] w_n4625_0;
	wire[1:0] w_n4626_0;
	wire[1:0] w_n4627_0;
	wire[1:0] w_n4628_0;
	wire[1:0] w_n4629_0;
	wire[1:0] w_n4632_0;
	wire[1:0] w_n4633_0;
	wire[1:0] w_n4635_0;
	wire[1:0] w_n4643_0;
	wire[1:0] w_n4652_0;
	wire[1:0] w_n4653_0;
	wire[1:0] w_n4656_0;
	wire[1:0] w_n4659_0;
	wire[1:0] w_n4663_0;
	wire[1:0] w_n4667_0;
	wire[1:0] w_n4668_0;
	wire[1:0] w_n4671_0;
	wire[1:0] w_n4674_0;
	wire[1:0] w_n4675_0;
	wire[1:0] w_n4676_0;
	wire[1:0] w_n4677_0;
	wire[1:0] w_n4685_0;
	wire[1:0] w_n4686_0;
	wire[1:0] w_n4694_0;
	wire[1:0] w_n4695_0;
	wire[1:0] w_n4697_0;
	wire[1:0] w_n4705_0;
	wire[1:0] w_n4706_0;
	wire[1:0] w_n4707_0;
	wire[1:0] w_n4708_0;
	wire[2:0] w_n4709_0;
	wire[1:0] w_n4710_0;
	wire[1:0] w_n4711_0;
	wire[1:0] w_n4712_0;
	wire[1:0] w_n4713_0;
	wire[1:0] w_n4716_0;
	wire[1:0] w_n4717_0;
	wire[1:0] w_n4719_0;
	wire[2:0] w_n4722_0;
	wire[1:0] w_n4727_0;
	wire[1:0] w_n4731_0;
	wire[1:0] w_n4739_0;
	wire[1:0] w_n4740_0;
	wire[1:0] w_n4743_0;
	wire[1:0] w_n4746_0;
	wire[1:0] w_n4747_0;
	wire[1:0] w_n4748_0;
	wire[1:0] w_n4749_0;
	wire[1:0] w_n4757_0;
	wire[1:0] w_n4758_0;
	wire[1:0] w_n4759_0;
	wire[1:0] w_n4767_0;
	wire[1:0] w_n4768_0;
	wire[1:0] w_n4769_0;
	wire[1:0] w_n4770_0;
	wire[2:0] w_n4771_0;
	wire[1:0] w_n4773_0;
	wire[2:0] w_n4782_0;
	wire[1:0] w_n4783_0;
	wire[1:0] w_n4784_0;
	wire[1:0] w_n4785_0;
	wire[1:0] w_n4786_0;
	wire[1:0] w_n4789_0;
	wire[1:0] w_n4790_0;
	wire[1:0] w_n4793_0;
	wire[1:0] w_n4811_0;
	wire[1:0] w_n4813_0;
	wire[1:0] w_n4814_0;
	wire[1:0] w_n4817_0;
	wire[1:0] w_n4822_0;
	wire[1:0] w_n4825_0;
	wire[1:0] w_n4828_0;
	wire[2:0] w_n4829_0;
	wire[1:0] w_n4830_0;
	wire[1:0] w_n4833_0;
	wire[1:0] w_n4834_0;
	wire[1:0] w_n4842_0;
	wire[1:0] w_n4843_0;
	wire[1:0] w_n4845_0;
	wire[1:0] w_n4853_0;
	wire[1:0] w_n4854_0;
	wire[1:0] w_n4855_0;
	wire[1:0] w_n4861_0;
	wire[1:0] w_n4862_0;
	wire[1:0] w_n4863_0;
	wire[2:0] w_n4864_0;
	wire[1:0] w_n4865_0;
	wire[1:0] w_n4866_0;
	wire[1:0] w_n4867_0;
	wire[1:0] w_n4868_0;
	wire[1:0] w_n4871_0;
	wire[1:0] w_n4872_0;
	wire[1:0] w_n4874_0;
	wire[1:0] w_n4886_0;
	wire[1:0] w_n4887_0;
	wire[1:0] w_n4890_0;
	wire[1:0] w_n4893_0;
	wire[1:0] w_n4897_0;
	wire[1:0] w_n4901_0;
	wire[1:0] w_n4902_0;
	wire[1:0] w_n4905_0;
	wire[1:0] w_n4908_0;
	wire[2:0] w_n4914_0;
	wire[1:0] w_n4915_0;
	wire[1:0] w_n4916_0;
	wire[1:0] w_n4918_0;
	wire[1:0] w_n4926_0;
	wire[1:0] w_n4927_0;
	wire[1:0] w_n4928_0;
	wire[1:0] w_n4929_0;
	wire[2:0] w_n4930_0;
	wire[1:0] w_n4931_0;
	wire[1:0] w_n4932_0;
	wire[1:0] w_n4933_0;
	wire[1:0] w_n4934_0;
	wire[1:0] w_n4937_0;
	wire[1:0] w_n4938_0;
	wire[1:0] w_n4940_0;
	wire[1:0] w_n4952_0;
	wire[1:0] w_n4953_0;
	wire[1:0] w_n4956_0;
	wire[1:0] w_n4961_0;
	wire[1:0] w_n4969_0;
	wire[2:0] w_n4970_0;
	wire[1:0] w_n4972_0;
	wire[1:0] w_n4974_0;
	wire[1:0] w_n4982_0;
	wire[1:0] w_n4983_0;
	wire[1:0] w_n4988_0;
	wire[1:0] w_n4996_0;
	wire[1:0] w_n4997_0;
	wire[1:0] w_n4998_0;
	wire[1:0] w_n4999_0;
	wire[2:0] w_n5000_0;
	wire[1:0] w_n5001_0;
	wire[1:0] w_n5002_0;
	wire[1:0] w_n5003_0;
	wire[1:0] w_n5004_0;
	wire[1:0] w_n5007_0;
	wire[1:0] w_n5008_0;
	wire[1:0] w_n5010_0;
	wire[1:0] w_n5016_0;
	wire[1:0] w_n5017_0;
	wire[1:0] w_n5020_0;
	wire[1:0] w_n5023_0;
	wire[1:0] w_n5028_0;
	wire[1:0] w_n5029_0;
	wire[1:0] w_n5030_0;
	wire[1:0] w_n5034_0;
	wire[1:0] w_n5035_0;
	wire[1:0] w_n5043_0;
	wire[1:0] w_n5044_0;
	wire[1:0] w_n5045_0;
	wire[1:0] w_n5051_0;
	wire[1:0] w_n5052_0;
	wire[1:0] w_n5053_0;
	wire[2:0] w_n5054_0;
	wire[1:0] w_n5055_0;
	wire[1:0] w_n5056_0;
	wire[1:0] w_n5057_0;
	wire[1:0] w_n5058_0;
	wire[1:0] w_n5061_0;
	wire[1:0] w_n5062_0;
	wire[1:0] w_n5064_0;
	wire[1:0] w_n5070_0;
	wire[1:0] w_n5076_0;
	wire[1:0] w_n5077_0;
	wire[1:0] w_n5080_0;
	wire[1:0] w_n5083_0;
	wire[1:0] w_n5088_0;
	wire[1:0] w_n5096_0;
	wire[1:0] w_n5097_0;
	wire[1:0] w_n5100_0;
	wire[1:0] w_n5101_0;
	wire[2:0] w_n5102_0;
	wire[1:0] w_n5105_0;
	wire[1:0] w_n5106_0;
	wire[1:0] w_n5107_0;
	wire[1:0] w_n5108_0;
	wire[2:0] w_n5109_0;
	wire[1:0] w_n5110_0;
	wire[1:0] w_n5111_0;
	wire[1:0] w_n5112_0;
	wire[1:0] w_n5113_0;
	wire[1:0] w_n5116_0;
	wire[1:0] w_n5117_0;
	wire[1:0] w_n5119_0;
	wire[1:0] w_n5122_0;
	wire[1:0] w_n5134_0;
	wire[1:0] w_n5135_0;
	wire[1:0] w_n5138_0;
	wire[1:0] w_n5143_0;
	wire[1:0] w_n5145_0;
	wire[1:0] w_n5146_0;
	wire[1:0] w_n5147_0;
	wire[1:0] w_n5148_0;
	wire[1:0] w_n5156_0;
	wire[1:0] w_n5157_0;
	wire[1:0] w_n5158_0;
	wire[1:0] w_n5159_0;
	wire[2:0] w_n5160_0;
	wire[1:0] w_n5161_0;
	wire[1:0] w_n5162_0;
	wire[1:0] w_n5163_0;
	wire[1:0] w_n5164_0;
	wire[1:0] w_n5167_0;
	wire[1:0] w_n5168_0;
	wire[1:0] w_n5170_0;
	wire[1:0] w_n5184_0;
	wire[1:0] w_n5185_0;
	wire[1:0] w_n5188_0;
	wire[1:0] w_n5191_0;
	wire[1:0] w_n5193_0;
	wire[1:0] w_n5196_0;
	wire[1:0] w_n5197_0;
	wire[1:0] w_n5203_0;
	wire[1:0] w_n5204_0;
	wire[1:0] w_n5205_0;
	wire[2:0] w_n5206_0;
	wire[1:0] w_n5207_0;
	wire[1:0] w_n5208_0;
	wire[1:0] w_n5209_0;
	wire[1:0] w_n5210_0;
	wire[1:0] w_n5213_0;
	wire[1:0] w_n5214_0;
	wire[1:0] w_n5216_0;
	wire[1:0] w_n5219_0;
	wire[1:0] w_n5229_0;
	wire[1:0] w_n5230_0;
	wire[1:0] w_n5233_0;
	wire[2:0] w_n5236_0;
	wire[1:0] w_n5238_0;
	wire[1:0] w_n5239_0;
	wire[1:0] w_n5240_0;
	wire[1:0] w_n5243_0;
	wire[2:0] w_n5244_0;
	wire[1:0] w_n5245_0;
	wire[1:0] w_n5246_0;
	wire[1:0] w_n5247_0;
	wire[1:0] w_n5248_0;
	wire[1:0] w_n5252_0;
	wire[1:0] w_n5253_0;
	wire[1:0] w_n5323_0;
	wire[2:0] w_n5332_0;
	wire[1:0] w_n5332_1;
	wire[1:0] w_n5334_0;
	wire[1:0] w_n5346_0;
	wire[2:0] w_n5347_0;
	wire[1:0] w_n5349_0;
	wire[1:0] w_n5350_0;
	wire[1:0] w_n5351_0;
	wire[1:0] w_n5354_0;
	wire[1:0] w_n5356_0;
	wire[1:0] w_n5357_0;
	wire[2:0] w_n5368_0;
	wire[1:0] w_n5369_0;
	wire[1:0] w_n5370_0;
	wire[1:0] w_n5371_0;
	wire[2:0] w_n5377_0;
	wire[1:0] w_n5378_0;
	wire[1:0] w_n5379_0;
	wire[2:0] w_n5390_0;
	wire[1:0] w_n5390_1;
	wire[1:0] w_n5395_0;
	wire[1:0] w_n5397_0;
	wire[1:0] w_n5398_0;
	wire[1:0] w_n5399_0;
	wire[2:0] w_n5400_0;
	wire[2:0] w_n5404_0;
	wire[1:0] w_n5405_0;
	wire[1:0] w_n5406_0;
	wire[2:0] w_n5415_0;
	wire[1:0] w_n5415_1;
	wire[1:0] w_n5416_0;
	wire[2:0] w_n5417_0;
	wire[1:0] w_n5418_0;
	wire[1:0] w_n5421_0;
	wire[2:0] w_n5431_0;
	wire[2:0] w_n5432_0;
	wire[1:0] w_n5435_0;
	wire[1:0] w_n5437_0;
	wire[2:0] w_n5438_0;
	wire[1:0] w_n5440_0;
	wire[1:0] w_n5441_0;
	wire[1:0] w_n5444_0;
	wire[1:0] w_n5446_0;
	wire[1:0] w_n5447_0;
	wire[1:0] w_n5449_0;
	wire[2:0] w_n5452_0;
	wire[1:0] w_n5452_1;
	wire[1:0] w_n5453_0;
	wire[2:0] w_n5454_0;
	wire[1:0] w_n5455_0;
	wire[1:0] w_n5458_0;
	wire[2:0] w_n5459_0;
	wire[1:0] w_n5461_0;
	wire[2:0] w_n5462_0;
	wire[1:0] w_n5463_0;
	wire[1:0] w_n5465_0;
	wire[1:0] w_n5466_0;
	wire[1:0] w_n5470_0;
	wire[1:0] w_n5471_0;
	wire[1:0] w_n5474_0;
	wire[1:0] w_n5476_0;
	wire[1:0] w_n5480_0;
	wire[1:0] w_n5483_0;
	wire[1:0] w_n5484_0;
	wire[1:0] w_n5487_0;
	wire w_dff_A_nhphmE1W6_0;
	wire w_dff_A_aq1r8Nrv9_0;
	wire w_dff_A_BnrGsSKY8_0;
	wire w_dff_A_9OrtdDC35_0;
	wire w_dff_A_GI8REpUn5_0;
	wire w_dff_A_i9IctGI95_0;
	wire w_dff_A_IuwzUmsQ4_0;
	wire w_dff_A_k4Whxaqa7_0;
	wire w_dff_A_H7NfKn0e1_1;
	wire w_dff_A_8u2TGooJ9_1;
	wire w_dff_A_zthfvi4X4_0;
	wire w_dff_A_STnUsJAO6_0;
	wire w_dff_A_MPoSOk006_0;
	wire w_dff_A_AZO8FXmC7_0;
	wire w_dff_A_mfNsh70O0_1;
	wire w_dff_A_wpA3GKq05_1;
	wire w_dff_A_MITM5qKS5_0;
	wire w_dff_A_CfbEZi267_0;
	wire w_dff_A_Ee8k0hks1_0;
	wire w_dff_A_cUDtSJyJ3_0;
	wire w_dff_A_DRpHc2cG9_1;
	wire w_dff_A_BPbGrQYz5_1;
	wire w_dff_A_Dd9u7gyD3_0;
	wire w_dff_A_lq02Zg2a4_0;
	wire w_dff_A_KCQwo8UC3_0;
	wire w_dff_A_xH2PJntQ0_0;
	wire w_dff_A_TJ7EiHcb4_1;
	wire w_dff_A_55rtkZ763_1;
	wire w_dff_A_Bg5Nu4RH8_0;
	wire w_dff_A_pThksnDn4_0;
	wire w_dff_A_yQupp8fW5_0;
	wire w_dff_A_B2o3GbHy5_0;
	wire w_dff_A_ppYAdYzc9_0;
	wire w_dff_A_ygimsAm25_0;
	wire w_dff_A_GkIFZOZv8_0;
	wire w_dff_A_MzbPBSaa5_0;
	wire w_dff_A_xKT4koJY9_0;
	wire w_dff_A_lykm64H75_0;
	wire w_dff_A_rj3wy9UT4_0;
	wire w_dff_A_fbO785X92_0;
	wire w_dff_A_Bppkcx0L3_1;
	wire w_dff_A_bDwv7Pyo2_1;
	wire w_dff_A_EdZtp1rz5_1;
	wire w_dff_A_Yd2y2bpJ5_1;
	wire w_dff_A_TQJu4EWX8_1;
	wire w_dff_A_9NWZDZCv5_1;
	wire w_dff_B_qpX2ZoCZ3_0;
	wire w_dff_A_g1w0aTHP1_0;
	wire w_dff_A_urx9Osvr5_0;
	wire w_dff_A_XhYdEVGP9_0;
	wire w_dff_A_cAl4L0fX0_0;
	wire w_dff_A_8BQJrza76_0;
	wire w_dff_A_uFawYx0e7_1;
	wire w_dff_A_imlgG5NP4_1;
	wire w_dff_A_KitWvW7m5_0;
	wire w_dff_A_EUkGuJ364_0;
	wire w_dff_A_Iu0AqP8D9_0;
	wire w_dff_A_wOYd2JLH5_1;
	wire w_dff_A_suv5RVkp5_1;
	wire w_dff_B_79XZBc8E3_1;
	wire w_dff_B_qjcjo5yK6_1;
	wire w_dff_B_pNwtQMbW3_0;
	wire w_dff_A_wA1LpPh75_1;
	wire w_dff_A_rXux2KXN2_1;
	wire w_dff_A_Ms0ywCUm8_1;
	wire w_dff_B_1F1gfXBh4_2;
	wire w_dff_B_VKoVih2S8_2;
	wire w_dff_B_zipXXgMG7_2;
	wire w_dff_B_3Y7HE1ps2_2;
	wire w_dff_B_r7mfL8Xx3_2;
	wire w_dff_B_2ZCumULd4_2;
	wire w_dff_B_lgQ2CJpm0_2;
	wire w_dff_B_tCtVDcet3_2;
	wire w_dff_B_f8hVMZUo0_2;
	wire w_dff_B_KcdrDF0c4_2;
	wire w_dff_B_TAg8WBza2_2;
	wire w_dff_B_KrYqum444_2;
	wire w_dff_B_QG15WaUo1_2;
	wire w_dff_B_nx4o88U60_2;
	wire w_dff_B_UhS4FA638_2;
	wire w_dff_B_JDNh7iiZ2_2;
	wire w_dff_B_OxKRY7227_2;
	wire w_dff_B_AU3fIqR25_2;
	wire w_dff_B_Kth0DFSO8_2;
	wire w_dff_B_g0gyRwvL0_2;
	wire w_dff_B_sHUH4X1Q0_2;
	wire w_dff_B_DNAmQGUn9_2;
	wire w_dff_B_aV2a0Cps4_2;
	wire w_dff_B_tZeRuOxq7_2;
	wire w_dff_B_3sZmPu2P2_2;
	wire w_dff_B_ZePAYJ262_2;
	wire w_dff_B_T8xTOSvj0_2;
	wire w_dff_B_n7qHaveF2_2;
	wire w_dff_B_zzK0lWC83_2;
	wire w_dff_B_WAsBDibx6_2;
	wire w_dff_B_YtehPBPw5_2;
	wire w_dff_B_ZCj9Sgpe9_2;
	wire w_dff_B_R9p6zXHr1_2;
	wire w_dff_B_rfl1FEMf9_2;
	wire w_dff_B_F7eW0GgV7_2;
	wire w_dff_B_aeFwX27L8_2;
	wire w_dff_B_VRSTJzhP5_2;
	wire w_dff_B_o3Y9g7EF3_2;
	wire w_dff_B_jLQg0u2Q6_2;
	wire w_dff_B_GcjS3Fik0_2;
	wire w_dff_B_gCZ78ql51_2;
	wire w_dff_B_O8Z66YzX5_2;
	wire w_dff_B_SZI9QF5N6_2;
	wire w_dff_B_FX9Tqe2G0_2;
	wire w_dff_B_Vf48OteZ5_2;
	wire w_dff_B_BjWISscr8_2;
	wire w_dff_B_vj2wDx672_2;
	wire w_dff_B_wDPUzVfv3_2;
	wire w_dff_B_qjQmfUAx7_2;
	wire w_dff_B_Azfpz1S68_2;
	wire w_dff_B_hcgaCqcM6_2;
	wire w_dff_B_3UeVQoDM4_2;
	wire w_dff_B_Q4AQdZVD8_2;
	wire w_dff_B_mHlD39nI3_2;
	wire w_dff_B_iEZyaL1c4_2;
	wire w_dff_B_XbZFELvh9_2;
	wire w_dff_B_mPS8lHRW8_2;
	wire w_dff_B_HcZRw80p2_2;
	wire w_dff_B_OmqXnA2Q9_2;
	wire w_dff_B_DYxtLUtm1_2;
	wire w_dff_B_D1Vf5IR67_2;
	wire w_dff_B_YaBbk4dy6_2;
	wire w_dff_B_skCxo6cn5_2;
	wire w_dff_B_oLai4ogo7_2;
	wire w_dff_B_oCqZeK9A2_2;
	wire w_dff_B_t8rZiQpd3_2;
	wire w_dff_B_g8A50B8m5_2;
	wire w_dff_B_dWR5q1Fo9_2;
	wire w_dff_B_pHDyiLtD2_2;
	wire w_dff_B_NMNpQCzb9_2;
	wire w_dff_B_l40YQyJq7_2;
	wire w_dff_B_BT3ftis21_2;
	wire w_dff_B_piv4UxAW4_2;
	wire w_dff_B_YaZOEOUM2_2;
	wire w_dff_B_7yHGmmnQ4_2;
	wire w_dff_B_Eqw1Eoid2_2;
	wire w_dff_B_gxMfK08z8_2;
	wire w_dff_B_wrNl0mPO3_2;
	wire w_dff_B_5wg4ZqNC2_2;
	wire w_dff_B_QZ2jD26B7_2;
	wire w_dff_B_mgLcBMrq0_2;
	wire w_dff_B_oqKx0yJG3_2;
	wire w_dff_B_a5YMA9Xd5_2;
	wire w_dff_B_nj95YJpD7_2;
	wire w_dff_B_ic5w4RTK2_2;
	wire w_dff_B_dXIi2qk55_2;
	wire w_dff_B_esowjK944_2;
	wire w_dff_B_lV2zAyrv2_2;
	wire w_dff_B_wdHBHGlt9_2;
	wire w_dff_B_12H6lgze3_2;
	wire w_dff_B_cfAJE7kt4_2;
	wire w_dff_B_6uoYTNQ31_2;
	wire w_dff_B_T5nNgsKl4_2;
	wire w_dff_B_2an2B9t30_2;
	wire w_dff_B_hHzmKy4M6_2;
	wire w_dff_B_cRoA1fFK0_2;
	wire w_dff_B_hTwIDE0m7_2;
	wire w_dff_B_Guqptcbx6_2;
	wire w_dff_B_VCH2f1942_2;
	wire w_dff_B_IANTEjUk4_2;
	wire w_dff_B_jUUEGEbz3_2;
	wire w_dff_B_5ILDH56V2_2;
	wire w_dff_B_fSqyH1h07_2;
	wire w_dff_B_66DMoCJC3_2;
	wire w_dff_B_0HtgoPMs5_2;
	wire w_dff_B_Vtxq4e4r5_2;
	wire w_dff_B_xGEbT75K7_2;
	wire w_dff_B_vH0bzWc02_2;
	wire w_dff_B_w7n94gEX8_2;
	wire w_dff_B_YFN78Xne8_2;
	wire w_dff_B_G3xf6Y8X5_2;
	wire w_dff_B_WeiAwsGA5_2;
	wire w_dff_B_AJtHLJFq3_2;
	wire w_dff_B_sgIIXb0q8_2;
	wire w_dff_B_rsT1Gty44_2;
	wire w_dff_B_trnnJA641_2;
	wire w_dff_B_uHnlTEZm1_2;
	wire w_dff_B_uipMsoLk5_2;
	wire w_dff_B_cdI1whfO0_2;
	wire w_dff_B_68oxuLKL0_2;
	wire w_dff_B_hdmnGyEV0_2;
	wire w_dff_B_6F56Vpri7_2;
	wire w_dff_B_rKPkvx055_2;
	wire w_dff_A_L0OSZQeM0_0;
	wire w_dff_A_EzVOOBro3_0;
	wire w_dff_A_S76g9eo65_0;
	wire w_dff_A_ym8OQgjx3_0;
	wire w_dff_A_SAnq582t7_0;
	wire w_dff_A_3DhaB3OS0_2;
	wire w_dff_A_kWqmFeRs7_2;
	wire w_dff_A_srR7HyzS7_2;
	wire w_dff_A_OBpDxHwd5_2;
	wire w_dff_A_Dhx2dUCK6_2;
	wire w_dff_A_SBZ1jIyq3_2;
	wire w_dff_A_reKGcl5w9_2;
	wire w_dff_A_3CAYALH19_2;
	wire w_dff_A_3WCqoWx00_2;
	wire w_dff_A_WClAtgeI0_2;
	wire w_dff_A_41HVUZn98_2;
	wire w_dff_A_mLXrjMgu6_2;
	wire w_dff_A_RYsBOHbI4_2;
	wire w_dff_A_dLlsKCHL4_2;
	wire w_dff_A_NX8QHL285_2;
	wire w_dff_A_xRtQnvNO0_2;
	wire w_dff_A_0QscNQfu9_2;
	wire w_dff_A_5TgjVQ6D2_2;
	wire w_dff_A_wdCcFoKc2_2;
	wire w_dff_A_7nV63SFc6_2;
	wire w_dff_A_F9b0VBf80_2;
	wire w_dff_A_D1Do9hXi2_2;
	wire w_dff_A_Wr6rtGAY9_2;
	wire w_dff_A_51A04pXA4_2;
	wire w_dff_A_Hfc4Msnq2_2;
	wire w_dff_A_WbIvKlhB1_2;
	wire w_dff_A_KiShnFwz1_2;
	wire w_dff_A_ON4G458g6_2;
	wire w_dff_A_yEunRhnk7_2;
	wire w_dff_A_S1qxlL0P9_2;
	wire w_dff_A_SdjizuFJ5_2;
	wire w_dff_A_DqhU2h8p0_2;
	wire w_dff_A_6KqLycjQ3_2;
	wire w_dff_A_s366T35O6_2;
	wire w_dff_A_NpGDyYQY8_2;
	wire w_dff_A_bbaWNdBH9_2;
	wire w_dff_A_1rxV4xZO2_2;
	wire w_dff_A_IOp0rUXs9_2;
	wire w_dff_A_YwlGR1es5_2;
	wire w_dff_A_6OZN7T3U7_2;
	wire w_dff_A_qPkaeIQa7_2;
	wire w_dff_A_TbPrP1sW3_2;
	wire w_dff_A_IxICBTvT9_2;
	wire w_dff_A_9fZQPXhh0_0;
	wire w_dff_A_jveqLtSa7_1;
	wire w_dff_A_0wlIeazr9_0;
	wire w_dff_A_xMHNluYy5_0;
	wire w_dff_A_ghwMUcgR8_0;
	wire w_dff_A_ruo15GOT6_0;
	wire w_dff_A_bxvqYTYx4_0;
	wire w_dff_A_zf31BzpE2_0;
	wire w_dff_A_A2xONnuD7_0;
	wire w_dff_A_vrPoZQgf4_0;
	wire w_dff_A_AlQfCFvp1_0;
	wire w_dff_A_c4lpFFo59_0;
	wire w_dff_A_qqLHRbws4_0;
	wire w_dff_A_ws4tWc4i8_0;
	wire w_dff_A_CepdS1678_0;
	wire w_dff_A_kXRcecfy2_0;
	wire w_dff_A_rxmmLz2D9_0;
	wire w_dff_A_y8pPL52h4_0;
	wire w_dff_A_nhCEAzVC8_0;
	wire w_dff_A_4X71YBkO2_0;
	wire w_dff_A_gvfmGipg2_0;
	wire w_dff_A_JzuBWyFX9_1;
	wire w_dff_A_RcIzSiyI2_2;
	wire w_dff_A_e7OvVlbE3_0;
	wire w_dff_A_x8u3rqMD0_0;
	wire w_dff_A_P2fU1v5w1_0;
	wire w_dff_A_3xwklP8D3_0;
	wire w_dff_A_1GEFQsI24_0;
	wire w_dff_A_e2sVsjtH3_0;
	wire w_dff_A_O2BO2SuL6_0;
	wire w_dff_A_ZJQET9YO9_0;
	wire w_dff_A_mc8ahk2U2_0;
	wire w_dff_A_49KuOZhG8_0;
	wire w_dff_A_GCpml2Rb2_0;
	wire w_dff_A_9FdPHtPY2_0;
	wire w_dff_A_mSsyGlbX9_0;
	wire w_dff_A_HLhGPyqR3_0;
	wire w_dff_A_1O6kJoWc7_0;
	wire w_dff_A_w2WYrEui2_0;
	wire w_dff_A_lAXy6uRz5_0;
	wire w_dff_A_AftDaAqX0_0;
	wire w_dff_A_7Fzu6oUl4_0;
	wire w_dff_A_zlRC7fJ27_0;
	wire w_dff_A_eAGqGZV06_0;
	wire w_dff_A_VdNX6NyX9_0;
	wire w_dff_A_MT890JFd0_0;
	wire w_dff_A_11Rao2mE8_0;
	wire w_dff_A_Sb9gVHhB4_0;
	wire w_dff_A_hvUl05Pf1_0;
	wire w_dff_A_9OZLVE5l3_0;
	wire w_dff_A_jtnIGmFe4_0;
	wire w_dff_A_zUG6Bm9Q7_0;
	wire w_dff_A_XxcD9WVy3_0;
	wire w_dff_A_RyqwCY9u2_0;
	wire w_dff_A_FxOhrNQK7_0;
	wire w_dff_A_Qn7JLtK60_0;
	wire w_dff_A_oSQJc16z0_0;
	wire w_dff_A_FKebBWTn9_0;
	wire w_dff_A_Yzu5N13E9_0;
	wire w_dff_A_ckZ4nhGs3_0;
	wire w_dff_A_rRcHmzzS2_0;
	wire w_dff_A_SFMSlVxD8_0;
	wire w_dff_A_cUSIBKFX0_0;
	wire w_dff_A_zCNYNeL25_0;
	wire w_dff_A_d8buYoeM8_0;
	wire w_dff_A_LSNUlBTH4_0;
	wire w_dff_A_UEaQSzRB1_0;
	wire w_dff_A_lqrq3xOV2_0;
	wire w_dff_A_aLvUiHOn0_2;
	wire w_dff_A_36xkr33S4_0;
	wire w_dff_A_o55eBeBQ4_0;
	wire w_dff_A_I44ZRdTT2_0;
	wire w_dff_A_BBmXfpbl4_0;
	wire w_dff_A_0ub60h0U0_0;
	wire w_dff_A_MZFFVovT9_0;
	wire w_dff_A_IHLM9I733_0;
	wire w_dff_A_KLHWcDfI4_0;
	wire w_dff_A_Hd0B8Jnf1_0;
	wire w_dff_A_2vEbmlFC5_0;
	wire w_dff_A_hSQHa8jX8_0;
	wire w_dff_A_3RiqyP598_0;
	wire w_dff_A_m7toEkNz9_0;
	wire w_dff_A_g8OhgRoj8_0;
	wire w_dff_A_nigqpQkF5_0;
	wire w_dff_A_A1jV4zv96_0;
	wire w_dff_A_2I9T2eCA4_0;
	wire w_dff_A_KicReXWK1_0;
	wire w_dff_A_3XaUSEr87_0;
	wire w_dff_A_NkYjzl1y2_0;
	wire w_dff_A_KnkghA6m8_0;
	wire w_dff_A_fIQ9wPgT5_0;
	wire w_dff_A_sYPqM0Ne0_0;
	wire w_dff_A_1dBbuaDt8_0;
	wire w_dff_A_ddmVdl7d3_0;
	wire w_dff_A_MltskOaQ4_0;
	wire w_dff_A_dLbVsA956_0;
	wire w_dff_A_byJOwl0s0_0;
	wire w_dff_A_KwEVwRUv5_0;
	wire w_dff_A_QujEOu9A6_0;
	wire w_dff_A_c53COlZH7_0;
	wire w_dff_A_EkkJoVIu3_0;
	wire w_dff_A_FtCXtbQg9_0;
	wire w_dff_A_vAmYOYGm1_0;
	wire w_dff_A_ZESBphvC5_0;
	wire w_dff_A_uRDFrFV11_0;
	wire w_dff_A_JJxzZPom5_0;
	wire w_dff_A_zLTGmJ074_0;
	wire w_dff_A_6Q65BMSk9_0;
	wire w_dff_A_g2OhW2KO0_0;
	wire w_dff_A_MkI2c3Bi5_0;
	wire w_dff_A_N1eAxMfr7_2;
	wire w_dff_A_Rq5spMDm0_0;
	wire w_dff_A_i9nintPf9_0;
	wire w_dff_A_AblW14053_0;
	wire w_dff_A_6dVfI5uI0_0;
	wire w_dff_A_n8tTywNa8_0;
	wire w_dff_A_UMCcn4bR2_0;
	wire w_dff_A_NUur3pNc7_0;
	wire w_dff_A_p3ALE3In6_0;
	wire w_dff_A_NNjP8ur99_0;
	wire w_dff_A_I6THQCKm2_0;
	wire w_dff_A_oDiZMTry0_0;
	wire w_dff_A_T9qHtUv04_0;
	wire w_dff_A_J261o2Ss1_0;
	wire w_dff_A_gb1thYBX5_0;
	wire w_dff_A_OOVB7UZJ9_0;
	wire w_dff_A_PduTcBVN6_0;
	wire w_dff_A_2Rx7qi8X1_0;
	wire w_dff_A_ibZGM0ph6_0;
	wire w_dff_A_LlfKHEXB0_0;
	wire w_dff_A_dZYeahfo5_0;
	wire w_dff_A_MVwpyAgL3_0;
	wire w_dff_A_Dxjd7JBQ6_0;
	wire w_dff_A_Z7ToR5508_0;
	wire w_dff_A_xr2NpMAe7_0;
	wire w_dff_A_B2LKw6Hh0_0;
	wire w_dff_A_ny4AM0fk2_0;
	wire w_dff_A_jNH3n5Mv4_0;
	wire w_dff_A_B1EZ8cCP3_0;
	wire w_dff_A_gZpOUTGo5_0;
	wire w_dff_A_ns0uvPKF4_0;
	wire w_dff_A_D5etW4Tb0_0;
	wire w_dff_A_TMcxvjUk7_0;
	wire w_dff_A_wuUwQJDP6_0;
	wire w_dff_A_ZnA4sBYo1_0;
	wire w_dff_A_qmQpENUI5_0;
	wire w_dff_A_UmRC19KI8_0;
	wire w_dff_A_UhCzM3vJ9_0;
	wire w_dff_A_9rl593Pk8_0;
	wire w_dff_A_Qcnenz3c3_0;
	wire w_dff_A_GzWX4srB6_0;
	wire w_dff_A_GpXyXXB64_2;
	wire w_dff_A_ALipnorC1_0;
	wire w_dff_A_XhjQDMNB6_0;
	wire w_dff_A_7H1A6hjr8_0;
	wire w_dff_A_84qVARgy6_0;
	wire w_dff_A_cwKIrz4B6_0;
	wire w_dff_A_9YKuMTny4_0;
	wire w_dff_A_kAOXuQAV5_0;
	wire w_dff_A_PeA6fPhU6_0;
	wire w_dff_A_D7FMRUwh7_0;
	wire w_dff_A_miLhcljX0_0;
	wire w_dff_A_fa7iecpj0_0;
	wire w_dff_A_r0qUSK9q1_0;
	wire w_dff_A_7AXVUXh24_0;
	wire w_dff_A_v9AKyfJg1_0;
	wire w_dff_A_h3u6UiJg2_0;
	wire w_dff_A_88rRlTUG7_0;
	wire w_dff_A_UlO6ny3g1_0;
	wire w_dff_A_EW0FfGZY6_0;
	wire w_dff_A_JhvnjQke7_0;
	wire w_dff_A_lGeebp1P5_0;
	wire w_dff_A_DAsj5WNq9_0;
	wire w_dff_A_joayAzx24_0;
	wire w_dff_A_8D4lveQN6_0;
	wire w_dff_A_uVeIlb1G3_0;
	wire w_dff_A_7uCWuWUr2_0;
	wire w_dff_A_Mq2S7sZk4_0;
	wire w_dff_A_nER4U6K48_0;
	wire w_dff_A_IZv0YM7F1_0;
	wire w_dff_A_crm6Esgu7_0;
	wire w_dff_A_OFoQEhMQ7_0;
	wire w_dff_A_T3cjDN794_0;
	wire w_dff_A_70WuzKR46_0;
	wire w_dff_A_17BjVtui6_0;
	wire w_dff_A_A6PQVR7i4_0;
	wire w_dff_A_azR70T864_0;
	wire w_dff_A_6eS7l4G83_0;
	wire w_dff_A_rreE02PC5_0;
	wire w_dff_A_e5QaUZSQ6_0;
	wire w_dff_A_Kjg55Kq01_2;
	wire w_dff_A_exl6Wb7n2_0;
	wire w_dff_A_ClGP5wdM3_0;
	wire w_dff_A_u3xdwEuT4_0;
	wire w_dff_A_iEubiO8B1_0;
	wire w_dff_A_ruNAGpa23_0;
	wire w_dff_A_mCcryNGs9_0;
	wire w_dff_A_NCFpvP1o3_0;
	wire w_dff_A_KIkikeco2_0;
	wire w_dff_A_e1vnGn374_0;
	wire w_dff_A_sMop9cDf7_0;
	wire w_dff_A_r2Fd3AFe4_0;
	wire w_dff_A_z2psqKaj4_0;
	wire w_dff_A_dza0UVxx8_0;
	wire w_dff_A_Xq7W6AMn2_0;
	wire w_dff_A_FY2QkzWg3_0;
	wire w_dff_A_HqbCpj6h4_0;
	wire w_dff_A_FVmRCHvx7_0;
	wire w_dff_A_YeI9e0lF3_0;
	wire w_dff_A_izyZBich0_0;
	wire w_dff_A_8tKQAvOq7_0;
	wire w_dff_A_YXYPFMNK8_0;
	wire w_dff_A_BPX4faWu2_0;
	wire w_dff_A_gAdfh5234_0;
	wire w_dff_A_Af6nxECs9_0;
	wire w_dff_A_3xZjHrmI4_0;
	wire w_dff_A_Oy88hPKX9_0;
	wire w_dff_A_nE3iIpth5_0;
	wire w_dff_A_tMJTaLlv9_0;
	wire w_dff_A_n8Gz5rOt8_0;
	wire w_dff_A_bgY8fUOw5_0;
	wire w_dff_A_S6B5c8LW1_0;
	wire w_dff_A_rGTXUjBc0_0;
	wire w_dff_A_svb5edEV5_0;
	wire w_dff_A_QJRbqGjc5_0;
	wire w_dff_A_TXtnJcIN5_0;
	wire w_dff_A_hqtUx4ZL7_0;
	wire w_dff_A_jawdh4xz8_2;
	wire w_dff_A_9iV3vboV8_0;
	wire w_dff_A_mUGqYtG34_0;
	wire w_dff_A_PHsUUrIT5_0;
	wire w_dff_A_5dj5NOr98_0;
	wire w_dff_A_9epO0p3g9_0;
	wire w_dff_A_JduSHjIT0_0;
	wire w_dff_A_9iJivsOC3_0;
	wire w_dff_A_Ym1Im8Jw5_0;
	wire w_dff_A_S5O0Fwqf6_0;
	wire w_dff_A_R9HyIRHj3_0;
	wire w_dff_A_BiKzDwcT5_0;
	wire w_dff_A_OsQhl5lF6_0;
	wire w_dff_A_pzaFM3mo6_0;
	wire w_dff_A_n0WZ2Xct9_0;
	wire w_dff_A_VqCDgc329_0;
	wire w_dff_A_3Uak3UhB5_0;
	wire w_dff_A_LxsMLQuO6_0;
	wire w_dff_A_5ZFq95xx6_0;
	wire w_dff_A_2cwPZCds0_0;
	wire w_dff_A_zSbL8nS36_0;
	wire w_dff_A_fhU1izvd1_0;
	wire w_dff_A_JmUqeRJK8_0;
	wire w_dff_A_D73D64gy7_0;
	wire w_dff_A_1zth1a1g5_0;
	wire w_dff_A_Qx9kCEGX2_0;
	wire w_dff_A_EpvSigF52_0;
	wire w_dff_A_DtBBIc706_0;
	wire w_dff_A_uGsoqZmV7_0;
	wire w_dff_A_x4HO3zVQ9_0;
	wire w_dff_A_fMOgHJeK9_0;
	wire w_dff_A_B6YdI7do9_0;
	wire w_dff_A_gHKRirfE3_0;
	wire w_dff_A_Cn401hVH9_0;
	wire w_dff_A_D333eUok3_0;
	wire w_dff_A_Pe38P7pN5_2;
	wire w_dff_A_nCtEnPSJ2_0;
	wire w_dff_A_Ma3O3KvU1_0;
	wire w_dff_A_Ep7KrQup3_0;
	wire w_dff_A_e6ZbUdPx9_0;
	wire w_dff_A_msOno7Ka6_0;
	wire w_dff_A_tqzbhEqh8_0;
	wire w_dff_A_fsO3fsos1_0;
	wire w_dff_A_ghzjACQP6_0;
	wire w_dff_A_TDvTJT7n3_0;
	wire w_dff_A_CXJZvFPU5_0;
	wire w_dff_A_uyTcqu9B1_0;
	wire w_dff_A_Q2bnUvrU5_0;
	wire w_dff_A_wbCW6RWZ7_0;
	wire w_dff_A_zU6d6cKq6_0;
	wire w_dff_A_5b9FxAtZ5_0;
	wire w_dff_A_IDaLhTdA5_0;
	wire w_dff_A_VT3BquvT5_0;
	wire w_dff_A_f21aEBkc3_0;
	wire w_dff_A_mMSm4fmZ2_0;
	wire w_dff_A_g14aAOT03_0;
	wire w_dff_A_tAQiefrK0_0;
	wire w_dff_A_XNb9bnLK7_0;
	wire w_dff_A_Z4LR6hMY9_0;
	wire w_dff_A_8XUyS7db8_0;
	wire w_dff_A_jjEQFNqj1_0;
	wire w_dff_A_1troq28w6_0;
	wire w_dff_A_VYoYmtW93_0;
	wire w_dff_A_GPXb8OUm1_0;
	wire w_dff_A_uZYSGDVi8_0;
	wire w_dff_A_2VRka1ES2_0;
	wire w_dff_A_YkMkjnyG3_0;
	wire w_dff_A_gSW324tT4_0;
	wire w_dff_A_64zGTwWk3_2;
	wire w_dff_A_uoBovu303_0;
	wire w_dff_A_lWdZZcdk5_0;
	wire w_dff_A_XBM05sUU2_0;
	wire w_dff_A_DO1RDvC50_0;
	wire w_dff_A_AjYtVRkR7_0;
	wire w_dff_A_bK1kIERF9_0;
	wire w_dff_A_AKHF9kOM8_0;
	wire w_dff_A_KhCy3EHF8_0;
	wire w_dff_A_glSHPEDr3_0;
	wire w_dff_A_hxHpYU7r5_0;
	wire w_dff_A_8GHlr7Q89_0;
	wire w_dff_A_VOejKKPC9_0;
	wire w_dff_A_7pUuxhwX7_0;
	wire w_dff_A_P99XQ2265_0;
	wire w_dff_A_VF9FwnGg7_0;
	wire w_dff_A_DdghD26L5_0;
	wire w_dff_A_BDvvNO2J5_0;
	wire w_dff_A_hCOdVZp18_0;
	wire w_dff_A_4hSfu2Ow5_0;
	wire w_dff_A_DYm5XO3d1_0;
	wire w_dff_A_gpyHIEUg6_0;
	wire w_dff_A_ag1chzb80_0;
	wire w_dff_A_b8ff46Sh1_0;
	wire w_dff_A_5RXLLOWz5_0;
	wire w_dff_A_Q9sgvRmZ2_0;
	wire w_dff_A_GaacqGqW2_0;
	wire w_dff_A_LWnl3p6B3_0;
	wire w_dff_A_wFRmwx9C7_0;
	wire w_dff_A_YDV1FGeX0_0;
	wire w_dff_A_kHcegJFv5_0;
	wire w_dff_A_xitZ0m6h4_2;
	wire w_dff_A_GFtWDc9i0_0;
	wire w_dff_A_yD4fRJtr7_0;
	wire w_dff_A_6U0Wy77e6_0;
	wire w_dff_A_eIl7S7ze6_0;
	wire w_dff_A_33AONRCr6_0;
	wire w_dff_A_rk23tv952_0;
	wire w_dff_A_PDy9BJo49_0;
	wire w_dff_A_IrWmIFaR5_0;
	wire w_dff_A_dkMNYgt21_0;
	wire w_dff_A_oj0DwjpZ0_0;
	wire w_dff_A_PYfLi9Z31_0;
	wire w_dff_A_MPxYtxEM6_0;
	wire w_dff_A_71LUllYi9_0;
	wire w_dff_A_4JHIOQn55_0;
	wire w_dff_A_PBGcaEpT1_0;
	wire w_dff_A_S3P1buBC1_0;
	wire w_dff_A_jaYVMiG42_0;
	wire w_dff_A_aXInF5FS1_0;
	wire w_dff_A_iY0Av4zl2_0;
	wire w_dff_A_baKc940N6_0;
	wire w_dff_A_1w93GRRl7_0;
	wire w_dff_A_bilfhlDs8_0;
	wire w_dff_A_kgM4MgPf9_0;
	wire w_dff_A_W4XVNCal3_0;
	wire w_dff_A_HOYph2ei1_0;
	wire w_dff_A_kkT9ksFJ8_0;
	wire w_dff_A_7wsIWUxq1_0;
	wire w_dff_A_ds9s3jEa9_0;
	wire w_dff_A_8Yxnvs8b7_2;
	wire w_dff_A_SYPWSNcc7_0;
	wire w_dff_A_mFPo1r7P1_0;
	wire w_dff_A_2qRNLAHc7_0;
	wire w_dff_A_0TrraRCu0_0;
	wire w_dff_A_DNxIYxTd3_0;
	wire w_dff_A_o9SgQY2c2_0;
	wire w_dff_A_SdQ2osBz4_0;
	wire w_dff_A_ormlNuEr7_0;
	wire w_dff_A_y88nNxrE7_0;
	wire w_dff_A_bJsBhGGJ6_0;
	wire w_dff_A_gsNmYIGd5_0;
	wire w_dff_A_307EDnhC9_0;
	wire w_dff_A_ruBncPID5_0;
	wire w_dff_A_SuvKsSB52_0;
	wire w_dff_A_dy3ZYaHg3_0;
	wire w_dff_A_h3PoJ9bF4_0;
	wire w_dff_A_moWmkxYx5_0;
	wire w_dff_A_3AYTVXA91_0;
	wire w_dff_A_KQIyPtLu6_0;
	wire w_dff_A_WOFOicfO2_0;
	wire w_dff_A_3FiKsycw7_0;
	wire w_dff_A_2K98D7ug1_0;
	wire w_dff_A_bX9MNSnE5_0;
	wire w_dff_A_Dz8B5NhD2_0;
	wire w_dff_A_yfk4EEVA6_0;
	wire w_dff_A_dWWTNci52_0;
	wire w_dff_A_xTdiVglx2_2;
	wire w_dff_A_iKz2u3Ft2_0;
	wire w_dff_A_Kv10FGAn7_0;
	wire w_dff_A_MdLREMMe9_0;
	wire w_dff_A_ynVVe63h9_0;
	wire w_dff_A_c0lGk08l2_0;
	wire w_dff_A_4VhsE6I25_0;
	wire w_dff_A_bz8fAUZd0_0;
	wire w_dff_A_PXFejuCE3_0;
	wire w_dff_A_LpZgHsik2_0;
	wire w_dff_A_h4NgCVKe9_0;
	wire w_dff_A_oSsmJyKB3_0;
	wire w_dff_A_AOWMjE2N9_0;
	wire w_dff_A_eypCkUHH9_0;
	wire w_dff_A_4tRQtxpw5_0;
	wire w_dff_A_eRIEMAlA4_0;
	wire w_dff_A_k8ncxhei8_0;
	wire w_dff_A_1WFopbwc6_0;
	wire w_dff_A_Urc2OIlf8_0;
	wire w_dff_A_rrE04nif2_0;
	wire w_dff_A_8WsMtF2e0_0;
	wire w_dff_A_dqTM58VY9_0;
	wire w_dff_A_jBCqwqHM5_0;
	wire w_dff_A_p10qzOdw2_0;
	wire w_dff_A_kZdX2cu59_0;
	wire w_dff_A_aayeK3ua3_2;
	wire w_dff_A_VGdSfmU19_0;
	wire w_dff_A_V5ASmAJW4_0;
	wire w_dff_A_G7f3wmJt0_0;
	wire w_dff_A_jtyFGDub8_0;
	wire w_dff_A_f84gTufo3_0;
	wire w_dff_A_75J3istD6_0;
	wire w_dff_A_zZaK0t8K5_0;
	wire w_dff_A_cc09lsfE2_0;
	wire w_dff_A_Cm7P6Bt25_0;
	wire w_dff_A_O2tfOzqU8_0;
	wire w_dff_A_qFyzp0X27_0;
	wire w_dff_A_zoeSuDYo6_0;
	wire w_dff_A_vYCuIY6O1_0;
	wire w_dff_A_qvYGC0N36_0;
	wire w_dff_A_IHTE9jDe2_0;
	wire w_dff_A_HTxnzyPQ0_0;
	wire w_dff_A_eJSGrcMc5_0;
	wire w_dff_A_IlR0jRwe6_0;
	wire w_dff_A_rEIHsrsR0_0;
	wire w_dff_A_SLBpBbuv5_0;
	wire w_dff_A_2Pm6Yf1P8_0;
	wire w_dff_A_iRJl67vO2_0;
	wire w_dff_A_AXUFYtJ77_2;
	wire w_dff_A_5TAVS12D0_0;
	wire w_dff_A_vLnUZfVP7_0;
	wire w_dff_A_Kqhxnf8I0_0;
	wire w_dff_A_uF89uJ3j4_0;
	wire w_dff_A_3bidzuuM6_0;
	wire w_dff_A_Pp8SQXoO2_0;
	wire w_dff_A_MFRpCeGw4_0;
	wire w_dff_A_3IOEKufs7_0;
	wire w_dff_A_R0rBZZB28_0;
	wire w_dff_A_16JrRSM28_0;
	wire w_dff_A_GngooLNm4_0;
	wire w_dff_A_n1YSv8a61_0;
	wire w_dff_A_jdCWc5VP2_0;
	wire w_dff_A_1T4GIvtJ0_0;
	wire w_dff_A_Ti15zLwd1_0;
	wire w_dff_A_RgMAxGqo5_0;
	wire w_dff_A_BEXiJ5Yu3_0;
	wire w_dff_A_7DylCnW46_0;
	wire w_dff_A_ziewSLq43_0;
	wire w_dff_A_eolJeCl28_0;
	wire w_dff_A_i53FbZmW9_2;
	wire w_dff_A_hVj1eVRn2_0;
	wire w_dff_A_czrKWigV5_0;
	wire w_dff_A_OguOl2FX5_0;
	wire w_dff_A_NBsStWDP9_0;
	wire w_dff_A_0NaOZ1y67_0;
	wire w_dff_A_AfnOP99w3_0;
	wire w_dff_A_AwtUWFMI1_0;
	wire w_dff_A_M5tqbj6J2_0;
	wire w_dff_A_GiTQ42wU7_0;
	wire w_dff_A_aW7cCnZQ8_0;
	wire w_dff_A_fVmUA1oC1_0;
	wire w_dff_A_oeUyyrxc7_0;
	wire w_dff_A_ThJfWili0_0;
	wire w_dff_A_S99gi9db1_0;
	wire w_dff_A_HbdVtext7_0;
	wire w_dff_A_XnyY5NX66_0;
	wire w_dff_A_f9nbxHLb0_0;
	wire w_dff_A_9hSL2wJF7_0;
	wire w_dff_A_MRzbRLbX5_2;
	wire w_dff_A_bmcMeNgS4_0;
	wire w_dff_A_wDSIqWH43_0;
	wire w_dff_A_mgBB9fcK0_0;
	wire w_dff_A_CVdXtpmj5_0;
	wire w_dff_A_wkRbPaiG1_0;
	wire w_dff_A_79qiRzi08_0;
	wire w_dff_A_yCs0SDH25_0;
	wire w_dff_A_Tbr0acDy0_0;
	wire w_dff_A_JLox2jbS0_0;
	wire w_dff_A_K8h2N7414_0;
	wire w_dff_A_aOa6z9ue3_0;
	wire w_dff_A_P17RISnR3_0;
	wire w_dff_A_pW5IAoT87_0;
	wire w_dff_A_bBrHfNIo9_0;
	wire w_dff_A_JrSD9GXH9_0;
	wire w_dff_A_lnGqSLfY2_0;
	wire w_dff_A_MetX8NB96_2;
	wire w_dff_A_kFCIRYxd1_0;
	wire w_dff_A_6Y8hv5bq5_0;
	wire w_dff_A_ZQME5H1p6_0;
	wire w_dff_A_qgc6oGFr0_0;
	wire w_dff_A_bPL7G4gV4_0;
	wire w_dff_A_7xpwiQHR9_0;
	wire w_dff_A_5GHgZTa38_0;
	wire w_dff_A_rJ46syzs8_0;
	wire w_dff_A_OTlabvXC5_0;
	wire w_dff_A_1I877Ghn7_0;
	wire w_dff_A_vzSImIZ66_0;
	wire w_dff_A_T2c3bCeS4_0;
	wire w_dff_A_HbkmqjKA8_0;
	wire w_dff_A_XEFqRjOB6_0;
	wire w_dff_A_HU6Y95fG4_2;
	wire w_dff_A_fkSelirA5_0;
	wire w_dff_A_s9XgZCGz4_0;
	wire w_dff_A_ldn8tt7l8_0;
	wire w_dff_A_tooFhoxr9_0;
	wire w_dff_A_dC4MAl1s5_0;
	wire w_dff_A_FmpBvojb2_0;
	wire w_dff_A_UAdGPHSE4_0;
	wire w_dff_A_TKRQg00C4_0;
	wire w_dff_A_tPk8mCWW7_0;
	wire w_dff_A_FeGbU0Yv3_0;
	wire w_dff_A_fhuCuywo1_0;
	wire w_dff_A_GPqiqml02_2;
	wire w_dff_A_yfQkah866_0;
	wire w_dff_A_bUPQneH97_0;
	wire w_dff_A_KFuKxUiF3_0;
	wire w_dff_A_XiktjTX59_0;
	wire w_dff_A_8MC6z9Bx5_0;
	wire w_dff_A_BR5L0SJE6_0;
	wire w_dff_A_RyEZ8Cq11_0;
	wire w_dff_A_VKAVuqlZ6_0;
	wire w_dff_A_MLj3FGzh5_0;
	wire w_dff_A_1nMlhPpu8_2;
	wire w_dff_A_w7E0o7ab6_0;
	wire w_dff_A_V4HYM5qa8_0;
	wire w_dff_A_Zk6ZIW6G3_0;
	wire w_dff_A_Nng9uJFY2_0;
	wire w_dff_A_svTt3Rct3_0;
	wire w_dff_A_6A34fKVP7_0;
	wire w_dff_A_5DqkBfTU6_0;
	wire w_dff_A_AlCqYWkD8_2;
	wire w_dff_A_gNv4B3hs4_0;
	wire w_dff_A_zJu0IT1w5_0;
	wire w_dff_A_M6b6oqqB4_0;
	wire w_dff_A_OJtixmIZ4_0;
	wire w_dff_A_wcSxKrSD1_0;
	wire w_dff_A_QgvCi3b43_2;
	wire w_dff_A_nRfPDqbs5_0;
	wire w_dff_A_vzTX9Gql9_0;
	wire w_dff_A_eEF03FKE6_0;
	wire w_dff_A_S1RJz5WQ3_0;
	wire w_dff_A_khtMLhmf2_2;
	wire w_dff_A_ufMNppQ99_0;
	wire w_dff_A_JKLHkgMy0_0;
	wire w_dff_A_WEvisCtm5_0;
	wire w_dff_A_d1DL4wzM4_2;
	wire w_dff_A_6D1oDIwG4_0;
	wire w_dff_A_xOJ1iUnI3_0;
	jnot g0000(.din(w_a22_0[2]),.dout(n49),.clk(gclk));
	jor g0001(.dina(w_a1_0[2]),.dinb(w_a0_0[2]),.dout(n50),.clk(gclk));
	jor g0002(.dina(w_n50_0[2]),.dinb(w_a2_0[1]),.dout(n51),.clk(gclk));
	jor g0003(.dina(w_n51_0[1]),.dinb(w_a3_0[1]),.dout(n52),.clk(gclk));
	jor g0004(.dina(w_n52_0[1]),.dinb(w_a4_0[1]),.dout(n53),.clk(gclk));
	jor g0005(.dina(w_n53_0[1]),.dinb(w_a5_0[1]),.dout(n54),.clk(gclk));
	jor g0006(.dina(w_n54_0[1]),.dinb(w_a6_0[1]),.dout(n55),.clk(gclk));
	jor g0007(.dina(w_n55_0[1]),.dinb(w_a7_0[1]),.dout(n56),.clk(gclk));
	jor g0008(.dina(w_n56_0[1]),.dinb(w_a8_0[1]),.dout(n57),.clk(gclk));
	jor g0009(.dina(w_n57_0[1]),.dinb(w_a9_0[1]),.dout(n58),.clk(gclk));
	jor g0010(.dina(w_n58_0[1]),.dinb(w_a10_0[1]),.dout(n59),.clk(gclk));
	jor g0011(.dina(w_n59_0[1]),.dinb(w_a11_0[1]),.dout(n60),.clk(gclk));
	jor g0012(.dina(w_n60_0[1]),.dinb(w_a12_0[1]),.dout(n61),.clk(gclk));
	jor g0013(.dina(w_n61_0[1]),.dinb(w_a13_0[1]),.dout(n62),.clk(gclk));
	jor g0014(.dina(w_n62_0[1]),.dinb(w_a14_0[1]),.dout(n63),.clk(gclk));
	jor g0015(.dina(w_n63_0[1]),.dinb(w_a15_0[1]),.dout(n64),.clk(gclk));
	jor g0016(.dina(w_n64_0[1]),.dinb(w_a16_0[1]),.dout(n65),.clk(gclk));
	jor g0017(.dina(w_n65_0[1]),.dinb(w_a17_0[1]),.dout(n66),.clk(gclk));
	jor g0018(.dina(w_n66_0[1]),.dinb(w_a18_0[1]),.dout(n67),.clk(gclk));
	jor g0019(.dina(w_n67_0[1]),.dinb(w_a19_0[2]),.dout(n68),.clk(gclk));
	jand g0020(.dina(w_n68_0[1]),.dinb(w_n49_9[2]),.dout(n69),.clk(gclk));
	jxor g0021(.dina(w_n69_0[1]),.dinb(w_a20_0[2]),.dout(n70),.clk(gclk));
	jnot g0022(.din(w_a21_0[1]),.dout(n71),.clk(gclk));
	jor g0023(.dina(w_n68_0[0]),.dinb(w_a20_0[1]),.dout(n72),.clk(gclk));
	jand g0024(.dina(w_n72_0[1]),.dinb(w_n49_9[1]),.dout(n73),.clk(gclk));
	jxor g0025(.dina(w_n73_0[1]),.dinb(w_n71_0[1]),.dout(n74),.clk(gclk));
	jor g0026(.dina(w_n74_1[1]),.dinb(w_n70_1[1]),.dout(n75),.clk(gclk));
	jand g0027(.dina(w_n63_0[0]),.dinb(w_n49_9[0]),.dout(n76),.clk(gclk));
	jxor g0028(.dina(n76),.dinb(w_a15_0[0]),.dout(n77),.clk(gclk));
	jor g0029(.dina(w_n77_9[2]),.dinb(w_n75_2[1]),.dout(n78),.clk(gclk));
	jnot g0030(.din(w_a19_0[1]),.dout(n79),.clk(gclk));
	jand g0031(.dina(w_n67_0[0]),.dinb(w_n49_8[2]),.dout(n80),.clk(gclk));
	jxor g0032(.dina(w_n80_0[1]),.dinb(n79),.dout(n81),.clk(gclk));
	jand g0033(.dina(w_n66_0[0]),.dinb(w_n49_8[1]),.dout(n82),.clk(gclk));
	jxor g0034(.dina(n82),.dinb(w_a18_0[0]),.dout(n83),.clk(gclk));
	jnot g0035(.din(w_n83_0[2]),.dout(n84),.clk(gclk));
	jand g0036(.dina(w_n84_0[2]),.dinb(w_n81_0[2]),.dout(n85),.clk(gclk));
	jand g0037(.dina(w_n65_0[0]),.dinb(w_n49_8[0]),.dout(n86),.clk(gclk));
	jxor g0038(.dina(n86),.dinb(w_a17_0[0]),.dout(n87),.clk(gclk));
	jnot g0039(.din(w_n87_0[2]),.dout(n88),.clk(gclk));
	jand g0040(.dina(w_n64_0[0]),.dinb(w_n49_7[2]),.dout(n89),.clk(gclk));
	jxor g0041(.dina(n89),.dinb(w_a16_0[0]),.dout(n90),.clk(gclk));
	jand g0042(.dina(w_n90_0[2]),.dinb(w_n88_0[1]),.dout(n91),.clk(gclk));
	jand g0043(.dina(w_n91_1[1]),.dinb(w_n85_1[1]),.dout(n92),.clk(gclk));
	jnot g0044(.din(w_n92_3[2]),.dout(n93),.clk(gclk));
	jor g0045(.dina(w_n93_1[2]),.dinb(w_n78_3[2]),.dout(n94),.clk(gclk));
	jxor g0046(.dina(w_n80_0[0]),.dinb(w_a19_0[0]),.dout(n95),.clk(gclk));
	jand g0047(.dina(w_n83_0[1]),.dinb(w_n95_0[1]),.dout(n96),.clk(gclk));
	jand g0048(.dina(w_n90_0[1]),.dinb(w_n87_0[1]),.dout(n97),.clk(gclk));
	jand g0049(.dina(w_n97_1[1]),.dinb(w_n96_1[1]),.dout(n98),.clk(gclk));
	jnot g0050(.din(w_n98_3[2]),.dout(n99),.clk(gclk));
	jnot g0051(.din(w_n77_9[1]),.dout(n100),.clk(gclk));
	jor g0052(.dina(w_n100_8[2]),.dinb(w_n75_2[0]),.dout(n101),.clk(gclk));
	jor g0053(.dina(w_n101_3[2]),.dinb(w_n99_3[1]),.dout(n102),.clk(gclk));
	jand g0054(.dina(w_n102_3[1]),.dinb(w_n94_2[2]),.dout(n103),.clk(gclk));
	jnot g0055(.din(w_a20_0[0]),.dout(n104),.clk(gclk));
	jxor g0056(.dina(w_n69_0[0]),.dinb(n104),.dout(n105),.clk(gclk));
	jxor g0057(.dina(w_n73_0[0]),.dinb(w_a21_0[0]),.dout(n106),.clk(gclk));
	jor g0058(.dina(w_n106_1[1]),.dinb(w_n105_1[1]),.dout(n107),.clk(gclk));
	jor g0059(.dina(w_n107_0[1]),.dinb(w_n100_8[1]),.dout(n108),.clk(gclk));
	jnot g0060(.din(w_n90_0[0]),.dout(n109),.clk(gclk));
	jand g0061(.dina(w_n109_0[1]),.dinb(w_n88_0[0]),.dout(n110),.clk(gclk));
	jand g0062(.dina(w_n83_0[0]),.dinb(w_n81_0[1]),.dout(n111),.clk(gclk));
	jand g0063(.dina(w_n111_1[1]),.dinb(w_n110_1[2]),.dout(n112),.clk(gclk));
	jnot g0064(.din(w_n112_4[1]),.dout(n113),.clk(gclk));
	jor g0065(.dina(w_n113_2[2]),.dinb(w_n108_4[2]),.dout(n114),.clk(gclk));
	jand g0066(.dina(w_n109_0[0]),.dinb(w_n87_0[0]),.dout(n115),.clk(gclk));
	jand g0067(.dina(w_n115_1[1]),.dinb(w_n96_1[0]),.dout(n116),.clk(gclk));
	jand g0068(.dina(w_n74_1[0]),.dinb(w_n105_1[0]),.dout(n117),.clk(gclk));
	jand g0069(.dina(w_n117_1[1]),.dinb(w_n100_8[0]),.dout(n118),.clk(gclk));
	jand g0070(.dina(w_n118_6[2]),.dinb(w_n116_3[1]),.dout(n119),.clk(gclk));
	jnot g0071(.din(w_n119_0[1]),.dout(n120),.clk(gclk));
	jand g0072(.dina(w_n120_2[2]),.dinb(w_n114_3[2]),.dout(n121),.clk(gclk));
	jand g0073(.dina(n121),.dinb(w_n103_1[1]),.dout(n122),.clk(gclk));
	jnot g0074(.din(w_n116_3[0]),.dout(n123),.clk(gclk));
	jor g0075(.dina(w_n123_2[1]),.dinb(w_n108_4[1]),.dout(n124),.clk(gclk));
	jor g0076(.dina(w_n107_0[0]),.dinb(w_n77_9[0]),.dout(n125),.clk(gclk));
	jand g0077(.dina(w_n111_1[0]),.dinb(w_n91_1[0]),.dout(n126),.clk(gclk));
	jnot g0078(.din(w_n126_4[1]),.dout(n127),.clk(gclk));
	jor g0079(.dina(w_n127_3[1]),.dinb(w_n125_5[1]),.dout(n128),.clk(gclk));
	jand g0080(.dina(w_n128_3[1]),.dinb(w_n124_2[2]),.dout(n129),.clk(gclk));
	jand g0081(.dina(w_n111_0[2]),.dinb(w_n97_1[0]),.dout(n130),.clk(gclk));
	jand g0082(.dina(w_n130_3[1]),.dinb(w_n117_1[0]),.dout(n131),.clk(gclk));
	jand g0083(.dina(w_n131_0[1]),.dinb(w_n77_8[2]),.dout(n132),.clk(gclk));
	jnot g0084(.din(w_n132_0[2]),.dout(n133),.clk(gclk));
	jor g0085(.dina(w_n74_0[2]),.dinb(w_n105_0[2]),.dout(n134),.clk(gclk));
	jor g0086(.dina(w_n134_1[1]),.dinb(w_n100_7[2]),.dout(n135),.clk(gclk));
	jor g0087(.dina(w_n135_4[2]),.dinb(w_n123_2[0]),.dout(n136),.clk(gclk));
	jand g0088(.dina(w_n136_2[1]),.dinb(w_n133_2[1]),.dout(n137),.clk(gclk));
	jor g0089(.dina(w_n134_1[0]),.dinb(w_n77_8[1]),.dout(n138),.clk(gclk));
	jand g0090(.dina(w_n84_0[1]),.dinb(w_n95_0[0]),.dout(n139),.clk(gclk));
	jand g0091(.dina(w_n139_1[1]),.dinb(w_n115_1[0]),.dout(n140),.clk(gclk));
	jnot g0092(.din(w_n140_3[1]),.dout(n141),.clk(gclk));
	jor g0093(.dina(w_n141_0[1]),.dinb(w_n138_4[1]),.dout(n142),.clk(gclk));
	jand g0094(.dina(w_n106_1[0]),.dinb(w_n70_1[0]),.dout(n143),.clk(gclk));
	jand g0095(.dina(w_n143_1[1]),.dinb(w_n100_7[1]),.dout(n144),.clk(gclk));
	jand g0096(.dina(w_n139_1[0]),.dinb(w_n97_0[2]),.dout(n145),.clk(gclk));
	jand g0097(.dina(w_n145_3[1]),.dinb(w_n144_6[2]),.dout(n146),.clk(gclk));
	jnot g0098(.din(w_n146_0[1]),.dout(n147),.clk(gclk));
	jand g0099(.dina(w_n147_2[1]),.dinb(w_n142_2[1]),.dout(n148),.clk(gclk));
	jand g0100(.dina(w_n148_1[1]),.dinb(w_n137_2[1]),.dout(n149),.clk(gclk));
	jand g0101(.dina(n149),.dinb(w_n129_1[2]),.dout(n150),.clk(gclk));
	jnot g0102(.din(w_n130_3[0]),.dout(n151),.clk(gclk));
	jor g0103(.dina(w_n135_4[1]),.dinb(w_n151_2[2]),.dout(n152),.clk(gclk));
	jand g0104(.dina(w_n152_2[2]),.dinb(w_n150_0[1]),.dout(n153),.clk(gclk));
	jand g0105(.dina(w_n143_1[0]),.dinb(w_n77_8[0]),.dout(n154),.clk(gclk));
	jand g0106(.dina(w_n139_0[2]),.dinb(w_n91_0[2]),.dout(n155),.clk(gclk));
	jand g0107(.dina(w_n155_3[2]),.dinb(w_n154_6[2]),.dout(n156),.clk(gclk));
	jnot g0108(.din(n156),.dout(n157),.clk(gclk));
	jor g0109(.dina(w_n125_5[0]),.dinb(w_n123_1[2]),.dout(n158),.clk(gclk));
	jor g0110(.dina(w_n123_1[1]),.dinb(w_n75_1[2]),.dout(n159),.clk(gclk));
	jor g0111(.dina(w_n159_1[1]),.dinb(w_n100_7[0]),.dout(n160),.clk(gclk));
	jand g0112(.dina(w_n160_2[2]),.dinb(w_n158_1[2]),.dout(n161),.clk(gclk));
	jor g0113(.dina(w_n138_4[0]),.dinb(w_n151_2[1]),.dout(n162),.clk(gclk));
	jand g0114(.dina(w_n162_2[1]),.dinb(w_n161_0[2]),.dout(n163),.clk(gclk));
	jand g0115(.dina(n163),.dinb(w_n157_3[1]),.dout(n164),.clk(gclk));
	jnot g0116(.din(w_n155_3[1]),.dout(n165),.clk(gclk));
	jor g0117(.dina(w_n165_2[2]),.dinb(w_n138_3[2]),.dout(n166),.clk(gclk));
	jand g0118(.dina(w_n115_0[2]),.dinb(w_n111_0[1]),.dout(n167),.clk(gclk));
	jnot g0119(.din(w_n167_3[2]),.dout(n168),.clk(gclk));
	jor g0120(.dina(w_n168_2[1]),.dinb(w_n138_3[1]),.dout(n169),.clk(gclk));
	jand g0121(.dina(w_n169_2[1]),.dinb(w_n166_2[2]),.dout(n170),.clk(gclk));
	jand g0122(.dina(w_n96_0[2]),.dinb(w_n91_0[1]),.dout(n171),.clk(gclk));
	jand g0123(.dina(w_n171_4[1]),.dinb(w_n144_6[1]),.dout(n172),.clk(gclk));
	jnot g0124(.din(w_n172_0[1]),.dout(n173),.clk(gclk));
	jand g0125(.dina(w_n117_0[2]),.dinb(w_n77_7[2]),.dout(n174),.clk(gclk));
	jand g0126(.dina(w_n174_6[2]),.dinb(w_n167_3[1]),.dout(n175),.clk(gclk));
	jnot g0127(.din(n175),.dout(n176),.clk(gclk));
	jand g0128(.dina(w_n176_1[2]),.dinb(w_n173_1[2]),.dout(n177),.clk(gclk));
	jand g0129(.dina(w_n177_0[1]),.dinb(w_n170_3[1]),.dout(n178),.clk(gclk));
	jand g0130(.dina(n178),.dinb(n164),.dout(n179),.clk(gclk));
	jand g0131(.dina(n179),.dinb(n153),.dout(n180),.clk(gclk));
	jand g0132(.dina(w_n180_1[1]),.dinb(n122),.dout(n181),.clk(gclk));
	jor g0133(.dina(w_n168_2[0]),.dinb(w_n101_3[1]),.dout(n182),.clk(gclk));
	jand g0134(.dina(w_n74_0[1]),.dinb(w_n70_0[2]),.dout(n183),.clk(gclk));
	jand g0135(.dina(w_n183_0[2]),.dinb(w_n77_7[1]),.dout(n184),.clk(gclk));
	jand g0136(.dina(w_n115_0[1]),.dinb(w_n85_1[0]),.dout(n185),.clk(gclk));
	jand g0137(.dina(w_n185_3[2]),.dinb(w_n184_6[2]),.dout(n186),.clk(gclk));
	jnot g0138(.din(w_n186_0[1]),.dout(n187),.clk(gclk));
	jor g0139(.dina(w_n138_3[0]),.dinb(w_n127_3[0]),.dout(n188),.clk(gclk));
	jand g0140(.dina(w_n188_2[1]),.dinb(w_n187_2[1]),.dout(n189),.clk(gclk));
	jand g0141(.dina(w_n189_0[1]),.dinb(w_n182_3[1]),.dout(n190),.clk(gclk));
	jor g0142(.dina(w_n138_2[2]),.dinb(w_n123_1[0]),.dout(n191),.clk(gclk));
	jand g0143(.dina(w_n139_0[1]),.dinb(w_n110_1[1]),.dout(n192),.clk(gclk));
	jnot g0144(.din(w_n192_3[1]),.dout(n193),.clk(gclk));
	jor g0145(.dina(w_n193_2[1]),.dinb(w_n75_1[1]),.dout(n194),.clk(gclk));
	jor g0146(.dina(w_n194_0[2]),.dinb(w_n77_7[0]),.dout(n195),.clk(gclk));
	jand g0147(.dina(w_n118_6[1]),.dinb(w_n92_3[1]),.dout(n196),.clk(gclk));
	jnot g0148(.din(n196),.dout(n197),.clk(gclk));
	jand g0149(.dina(w_n197_3[1]),.dinb(w_n195_2[1]),.dout(n198),.clk(gclk));
	jand g0150(.dina(w_n198_1[1]),.dinb(w_n191_3[2]),.dout(n199),.clk(gclk));
	jand g0151(.dina(n199),.dinb(w_n190_1[2]),.dout(n200),.clk(gclk));
	jor g0152(.dina(w_n84_0[0]),.dinb(w_n81_0[0]),.dout(n201),.clk(gclk));
	jnot g0153(.din(w_n110_1[0]),.dout(n202),.clk(gclk));
	jor g0154(.dina(n202),.dinb(n201),.dout(n203),.clk(gclk));
	jor g0155(.dina(w_n203_1[1]),.dinb(w_n125_4[2]),.dout(n204),.clk(gclk));
	jand g0156(.dina(w_n140_3[0]),.dinb(w_n154_6[1]),.dout(n205),.clk(gclk));
	jnot g0157(.din(w_n205_0[1]),.dout(n206),.clk(gclk));
	jor g0158(.dina(w_n193_2[0]),.dinb(w_n125_4[1]),.dout(n207),.clk(gclk));
	jand g0159(.dina(w_n207_3[1]),.dinb(w_n206_2[1]),.dout(n208),.clk(gclk));
	jand g0160(.dina(n208),.dinb(w_n204_2[2]),.dout(n209),.clk(gclk));
	jand g0161(.dina(n209),.dinb(n200),.dout(n210),.clk(gclk));
	jand g0162(.dina(n210),.dinb(n181),.dout(n211),.clk(gclk));
	jand g0163(.dina(w_n140_2[2]),.dinb(w_n184_6[1]),.dout(n212),.clk(gclk));
	jnot g0164(.din(w_n212_0[1]),.dout(n213),.clk(gclk));
	jand g0165(.dina(w_n145_3[0]),.dinb(w_n154_6[0]),.dout(n214),.clk(gclk));
	jnot g0166(.din(w_n214_0[1]),.dout(n215),.clk(gclk));
	jor g0167(.dina(w_n106_0[2]),.dinb(w_n70_0[1]),.dout(n216),.clk(gclk));
	jor g0168(.dina(w_n216_0[2]),.dinb(w_n100_6[2]),.dout(n217),.clk(gclk));
	jor g0169(.dina(w_n217_4[1]),.dinb(w_n165_2[1]),.dout(n218),.clk(gclk));
	jand g0170(.dina(w_n218_3[2]),.dinb(w_n215_3[2]),.dout(n219),.clk(gclk));
	jand g0171(.dina(n219),.dinb(w_n213_3[1]),.dout(n220),.clk(gclk));
	jor g0172(.dina(w_n193_1[2]),.dinb(w_n135_4[0]),.dout(n221),.clk(gclk));
	jor g0173(.dina(w_n159_1[0]),.dinb(w_n77_6[2]),.dout(n222),.clk(gclk));
	jand g0174(.dina(w_n106_0[1]),.dinb(w_n105_0[1]),.dout(n223),.clk(gclk));
	jand g0175(.dina(w_n77_6[1]),.dinb(w_n223_3[1]),.dout(n224),.clk(gclk));
	jand g0176(.dina(w_n171_4[0]),.dinb(w_n224_5[1]),.dout(n225),.clk(gclk));
	jnot g0177(.din(n225),.dout(n226),.clk(gclk));
	jand g0178(.dina(w_n226_2[2]),.dinb(w_n222_3[1]),.dout(n227),.clk(gclk));
	jand g0179(.dina(n227),.dinb(w_n221_3[2]),.dout(n228),.clk(gclk));
	jand g0180(.dina(n228),.dinb(n220),.dout(n229),.clk(gclk));
	jand g0181(.dina(w_n97_0[1]),.dinb(w_n85_0[2]),.dout(n230),.clk(gclk));
	jnot g0182(.din(w_n230_3[1]),.dout(n231),.clk(gclk));
	jor g0183(.dina(w_n231_1[1]),.dinb(w_n135_3[2]),.dout(n232),.clk(gclk));
	jor g0184(.dina(w_n138_2[1]),.dinb(w_n93_1[1]),.dout(n233),.clk(gclk));
	jand g0185(.dina(w_n233_2[1]),.dinb(w_n232_4[2]),.dout(n234),.clk(gclk));
	jor g0186(.dina(w_n135_3[1]),.dinb(w_n127_2[2]),.dout(n235),.clk(gclk));
	jor g0187(.dina(w_n168_1[2]),.dinb(w_n135_3[0]),.dout(n236),.clk(gclk));
	jand g0188(.dina(w_n236_1[2]),.dinb(w_n235_2[1]),.dout(n237),.clk(gclk));
	jor g0189(.dina(w_n127_2[1]),.dinb(w_n101_3[0]),.dout(n238),.clk(gclk));
	jand g0190(.dina(w_n174_6[1]),.dinb(w_n112_4[0]),.dout(n239),.clk(gclk));
	jnot g0191(.din(w_n239_0[1]),.dout(n240),.clk(gclk));
	jand g0192(.dina(w_n240_2[1]),.dinb(w_n238_2[1]),.dout(n241),.clk(gclk));
	jand g0193(.dina(w_n241_0[1]),.dinb(n237),.dout(n242),.clk(gclk));
	jand g0194(.dina(n242),.dinb(w_n234_0[2]),.dout(n243),.clk(gclk));
	jor g0195(.dina(w_n231_1[0]),.dinb(w_n108_4[0]),.dout(n244),.clk(gclk));
	jor g0196(.dina(w_n217_4[0]),.dinb(w_n123_0[2]),.dout(n245),.clk(gclk));
	jand g0197(.dina(w_n245_2[1]),.dinb(w_n244_3[1]),.dout(n246),.clk(gclk));
	jand g0198(.dina(w_n230_3[0]),.dinb(w_n174_6[0]),.dout(n247),.clk(gclk));
	jnot g0199(.din(w_n247_0[1]),.dout(n248),.clk(gclk));
	jnot g0200(.din(w_n185_3[1]),.dout(n249),.clk(gclk));
	jor g0201(.dina(w_n249_2[1]),.dinb(w_n217_3[2]),.dout(n250),.clk(gclk));
	jand g0202(.dina(w_n250_2[2]),.dinb(w_n248_3[2]),.dout(n251),.clk(gclk));
	jor g0203(.dina(w_n203_1[0]),.dinb(w_n78_3[1]),.dout(n252),.clk(gclk));
	jand g0204(.dina(w_n183_0[1]),.dinb(w_n100_6[1]),.dout(n253),.clk(gclk));
	jand g0205(.dina(w_n140_2[1]),.dinb(w_n253_6[2]),.dout(n254),.clk(gclk));
	jnot g0206(.din(w_n254_0[2]),.dout(n255),.clk(gclk));
	jand g0207(.dina(w_n255_2[1]),.dinb(w_n252_4[1]),.dout(n256),.clk(gclk));
	jand g0208(.dina(n256),.dinb(w_n251_0[2]),.dout(n257),.clk(gclk));
	jand g0209(.dina(n257),.dinb(w_n246_0[2]),.dout(n258),.clk(gclk));
	jand g0210(.dina(n258),.dinb(n243),.dout(n259),.clk(gclk));
	jand g0211(.dina(n259),.dinb(w_n229_0[1]),.dout(n260),.clk(gclk));
	jor g0212(.dina(w_n217_3[1]),.dinb(w_n127_2[0]),.dout(n261),.clk(gclk));
	jand g0213(.dina(w_n100_6[0]),.dinb(w_n223_3[0]),.dout(n262),.clk(gclk));
	jand g0214(.dina(w_n110_0[2]),.dinb(w_n85_0[1]),.dout(n263),.clk(gclk));
	jand g0215(.dina(w_n263_4[1]),.dinb(w_n262_5[1]),.dout(n264),.clk(gclk));
	jnot g0216(.din(w_n264_0[1]),.dout(n265),.clk(gclk));
	jand g0217(.dina(w_n184_6[0]),.dinb(w_n98_3[1]),.dout(n266),.clk(gclk));
	jnot g0218(.din(w_n266_1[2]),.dout(n267),.clk(gclk));
	jnot g0219(.din(w_n263_4[0]),.dout(n268),.clk(gclk));
	jor g0220(.dina(w_n268_2[1]),.dinb(w_n135_2[2]),.dout(n269),.clk(gclk));
	jand g0221(.dina(w_n269_2[2]),.dinb(w_n267_3[1]),.dout(n270),.clk(gclk));
	jand g0222(.dina(n270),.dinb(w_n265_2[1]),.dout(n271),.clk(gclk));
	jand g0223(.dina(n271),.dinb(w_n261_2[2]),.dout(n272),.clk(gclk));
	jand g0224(.dina(n272),.dinb(w_n260_0[1]),.dout(n273),.clk(gclk));
	jand g0225(.dina(w_n145_2[2]),.dinb(w_n118_6[0]),.dout(n274),.clk(gclk));
	jnot g0226(.din(w_n274_0[1]),.dout(n275),.clk(gclk));
	jor g0227(.dina(w_n165_2[0]),.dinb(w_n108_3[2]),.dout(n276),.clk(gclk));
	jand g0228(.dina(w_n276_3[2]),.dinb(w_n275_2[1]),.dout(n277),.clk(gclk));
	jor g0229(.dina(w_n113_2[1]),.dinb(w_n78_3[0]),.dout(n278),.clk(gclk));
	jor g0230(.dina(w_n203_0[2]),.dinb(w_n134_0[2]),.dout(n279),.clk(gclk));
	jor g0231(.dina(w_n279_0[2]),.dinb(w_n77_6[0]),.dout(n280),.clk(gclk));
	jand g0232(.dina(w_n280_2[2]),.dinb(w_n278_1[2]),.dout(n281),.clk(gclk));
	jand g0233(.dina(w_n145_2[1]),.dinb(w_n262_5[0]),.dout(n282),.clk(gclk));
	jnot g0234(.din(w_n282_1[2]),.dout(n283),.clk(gclk));
	jand g0235(.dina(w_n283_2[1]),.dinb(w_n281_0[2]),.dout(n284),.clk(gclk));
	jand g0236(.dina(n284),.dinb(w_n277_0[1]),.dout(n285),.clk(gclk));
	jor g0237(.dina(w_n279_0[1]),.dinb(w_n100_5[2]),.dout(n286),.clk(gclk));
	jand g0238(.dina(w_n263_3[2]),.dinb(w_n184_5[2]),.dout(n287),.clk(gclk));
	jnot g0239(.din(w_n287_0[1]),.dout(n288),.clk(gclk));
	jnot g0240(.din(w_n171_3[2]),.dout(n289),.clk(gclk));
	jor g0241(.dina(w_n289_1[1]),.dinb(w_n135_2[1]),.dout(n290),.clk(gclk));
	jand g0242(.dina(w_n290_3[2]),.dinb(w_n288_2[1]),.dout(n291),.clk(gclk));
	jand g0243(.dina(n291),.dinb(w_n286_3[1]),.dout(n292),.clk(gclk));
	jand g0244(.dina(n292),.dinb(n285),.dout(n293),.clk(gclk));
	jor g0245(.dina(w_n138_2[0]),.dinb(w_n99_3[0]),.dout(n294),.clk(gclk));
	jand g0246(.dina(w_n140_2[0]),.dinb(w_n223_2[2]),.dout(n295),.clk(gclk));
	jand g0247(.dina(w_n295_0[2]),.dinb(w_n77_5[2]),.dout(n296),.clk(gclk));
	jnot g0248(.din(w_n296_0[1]),.dout(n297),.clk(gclk));
	jand g0249(.dina(w_n297_1[2]),.dinb(w_n294_3[2]),.dout(n298),.clk(gclk));
	jand g0250(.dina(w_n154_5[2]),.dinb(w_n92_3[0]),.dout(n299),.clk(gclk));
	jnot g0251(.din(w_n299_0[1]),.dout(n300),.clk(gclk));
	jand g0252(.dina(w_n145_2[0]),.dinb(w_n183_0[0]),.dout(n301),.clk(gclk));
	jand g0253(.dina(w_n301_1[1]),.dinb(w_n100_5[1]),.dout(n302),.clk(gclk));
	jnot g0254(.din(w_n302_0[2]),.dout(n303),.clk(gclk));
	jand g0255(.dina(w_n303_0[2]),.dinb(w_n300_3[1]),.dout(n304),.clk(gclk));
	jor g0256(.dina(w_n113_2[0]),.dinb(w_n101_2[2]),.dout(n305),.clk(gclk));
	jand g0257(.dina(w_n305_2[2]),.dinb(n304),.dout(n306),.clk(gclk));
	jand g0258(.dina(n306),.dinb(n298),.dout(n307),.clk(gclk));
	jand g0259(.dina(w_n145_1[2]),.dinb(w_n224_5[0]),.dout(n308),.clk(gclk));
	jnot g0260(.din(w_n308_0[1]),.dout(n309),.clk(gclk));
	jor g0261(.dina(w_n289_1[0]),.dinb(w_n125_4[0]),.dout(n310),.clk(gclk));
	jand g0262(.dina(w_n110_0[1]),.dinb(w_n96_0[1]),.dout(n311),.clk(gclk));
	jand g0263(.dina(w_n311_2[2]),.dinb(w_n224_4[2]),.dout(n312),.clk(gclk));
	jnot g0264(.din(w_n312_0[1]),.dout(n313),.clk(gclk));
	jand g0265(.dina(w_n230_2[2]),.dinb(w_n144_6[0]),.dout(n314),.clk(gclk));
	jnot g0266(.din(w_n314_0[2]),.dout(n315),.clk(gclk));
	jand g0267(.dina(w_n315_2[1]),.dinb(w_n313_1[2]),.dout(n316),.clk(gclk));
	jand g0268(.dina(w_n316_0[2]),.dinb(w_n310_2[2]),.dout(n317),.clk(gclk));
	jand g0269(.dina(n317),.dinb(w_n309_2[2]),.dout(n318),.clk(gclk));
	jand g0270(.dina(n318),.dinb(w_n307_0[1]),.dout(n319),.clk(gclk));
	jand g0271(.dina(n319),.dinb(w_n293_0[1]),.dout(n320),.clk(gclk));
	jor g0272(.dina(w_n165_1[2]),.dinb(w_n101_2[1]),.dout(n321),.clk(gclk));
	jand g0273(.dina(w_n321_3[1]),.dinb(w_n320_0[1]),.dout(n322),.clk(gclk));
	jand g0274(.dina(n322),.dinb(w_n273_0[1]),.dout(n323),.clk(gclk));
	jand g0275(.dina(n323),.dinb(n211),.dout(n324),.clk(gclk));
	jnot g0276(.din(w_n324_0[1]),.dout(n325),.clk(gclk));
	jand g0277(.dina(w_n294_3[1]),.dinb(w_n191_3[1]),.dout(n326),.clk(gclk));
	jor g0278(.dina(w_n289_0[2]),.dinb(w_n108_3[1]),.dout(n327),.clk(gclk));
	jand g0279(.dina(w_n327_1[2]),.dinb(w_n280_2[1]),.dout(n328),.clk(gclk));
	jand g0280(.dina(n328),.dinb(n326),.dout(n329),.clk(gclk));
	jand g0281(.dina(w_n253_6[1]),.dinb(w_n92_2[2]),.dout(n330),.clk(gclk));
	jnot g0282(.din(w_n330_0[2]),.dout(n331),.clk(gclk));
	jor g0283(.dina(w_n168_1[1]),.dinb(w_n78_2[2]),.dout(n332),.clk(gclk));
	jor g0284(.dina(w_n108_3[0]),.dinb(w_n93_1[0]),.dout(n333),.clk(gclk));
	jand g0285(.dina(w_n333_2[1]),.dinb(w_n332_3[1]),.dout(n334),.clk(gclk));
	jand g0286(.dina(w_n334_0[1]),.dinb(w_n331_2[2]),.dout(n335),.clk(gclk));
	jor g0287(.dina(w_n216_0[1]),.dinb(w_n77_5[1]),.dout(n336),.clk(gclk));
	jor g0288(.dina(w_n168_1[0]),.dinb(w_n336_2[2]),.dout(n337),.clk(gclk));
	jand g0289(.dina(w_n337_2[2]),.dinb(w_n250_2[1]),.dout(n338),.clk(gclk));
	jor g0290(.dina(w_n193_1[1]),.dinb(w_n108_2[2]),.dout(n339),.clk(gclk));
	jand g0291(.dina(w_n339_4[1]),.dinb(w_n176_1[1]),.dout(n340),.clk(gclk));
	jand g0292(.dina(w_n340_1[2]),.dinb(w_n133_2[0]),.dout(n341),.clk(gclk));
	jand g0293(.dina(n341),.dinb(w_n338_0[2]),.dout(n342),.clk(gclk));
	jand g0294(.dina(n342),.dinb(w_n335_0[2]),.dout(n343),.clk(gclk));
	jor g0295(.dina(w_n203_0[1]),.dinb(w_n108_2[1]),.dout(n344),.clk(gclk));
	jand g0296(.dina(w_n269_2[1]),.dinb(w_n188_2[0]),.dout(n345),.clk(gclk));
	jor g0297(.dina(w_n268_2[0]),.dinb(w_n125_3[2]),.dout(n346),.clk(gclk));
	jor g0298(.dina(w_n268_1[2]),.dinb(w_n138_1[2]),.dout(n347),.clk(gclk));
	jand g0299(.dina(w_n347_2[2]),.dinb(w_n346_2[2]),.dout(n348),.clk(gclk));
	jand g0300(.dina(n348),.dinb(w_n345_0[1]),.dout(n349),.clk(gclk));
	jand g0301(.dina(n349),.dinb(w_n344_3[1]),.dout(n350),.clk(gclk));
	jand g0302(.dina(w_n305_2[1]),.dinb(w_n238_2[0]),.dout(n351),.clk(gclk));
	jand g0303(.dina(w_n351_1[1]),.dinb(w_n288_2[0]),.dout(n352),.clk(gclk));
	jor g0304(.dina(w_n127_1[2]),.dinb(w_n108_2[0]),.dout(n353),.clk(gclk));
	jand g0305(.dina(w_n353_2[2]),.dinb(w_n195_2[0]),.dout(n354),.clk(gclk));
	jand g0306(.dina(n354),.dinb(w_n161_0[1]),.dout(n355),.clk(gclk));
	jand g0307(.dina(w_n355_0[1]),.dinb(w_n352_1[1]),.dout(n356),.clk(gclk));
	jand g0308(.dina(n356),.dinb(w_n350_0[1]),.dout(n357),.clk(gclk));
	jand g0309(.dina(n357),.dinb(n343),.dout(n358),.clk(gclk));
	jand g0310(.dina(n358),.dinb(w_n329_1[1]),.dout(n359),.clk(gclk));
	jand g0311(.dina(w_n171_3[1]),.dinb(w_n262_4[2]),.dout(n360),.clk(gclk));
	jnot g0312(.din(w_n360_0[2]),.dout(n361),.clk(gclk));
	jand g0313(.dina(w_n361_2[2]),.dinb(w_n120_2[1]),.dout(n362),.clk(gclk));
	jand g0314(.dina(w_n117_0[1]),.dinb(w_n112_3[2]),.dout(n363),.clk(gclk));
	jor g0315(.dina(n363),.dinb(w_n302_0[1]),.dout(n364),.clk(gclk));
	jnot g0316(.din(n364),.dout(n365),.clk(gclk));
	jor g0317(.dina(w_n249_2[0]),.dinb(w_n125_3[1]),.dout(n366),.clk(gclk));
	jand g0318(.dina(w_n366_3[1]),.dinb(w_n297_1[1]),.dout(n367),.clk(gclk));
	jand g0319(.dina(n367),.dinb(n365),.dout(n368),.clk(gclk));
	jand g0320(.dina(n368),.dinb(w_n362_0[1]),.dout(n369),.clk(gclk));
	jor g0321(.dina(w_n135_2[0]),.dinb(w_n99_2[2]),.dout(n370),.clk(gclk));
	jand g0322(.dina(w_n215_3[1]),.dinb(w_n206_2[0]),.dout(n371),.clk(gclk));
	jand g0323(.dina(n371),.dinb(w_n370_3[1]),.dout(n372),.clk(gclk));
	jor g0324(.dina(w_n231_0[2]),.dinb(w_n75_1[0]),.dout(n373),.clk(gclk));
	jor g0325(.dina(w_n373_0[2]),.dinb(w_n100_5[0]),.dout(n374),.clk(gclk));
	jand g0326(.dina(w_n374_3[1]),.dinb(w_n207_3[0]),.dout(n375),.clk(gclk));
	jand g0327(.dina(n375),.dinb(w_n372_0[1]),.dout(n376),.clk(gclk));
	jor g0328(.dina(w_n138_1[1]),.dinb(w_n113_1[2]),.dout(n377),.clk(gclk));
	jor g0329(.dina(w_n165_1[1]),.dinb(w_n78_2[1]),.dout(n378),.clk(gclk));
	jand g0330(.dina(w_n378_3[1]),.dinb(w_n377_3[2]),.dout(n379),.clk(gclk));
	jand g0331(.dina(w_n236_1[1]),.dinb(w_n162_2[0]),.dout(n380),.clk(gclk));
	jand g0332(.dina(n380),.dinb(n379),.dout(n381),.clk(gclk));
	jor g0333(.dina(w_n168_0[2]),.dinb(w_n108_1[2]),.dout(n382),.clk(gclk));
	jor g0334(.dina(w_n165_1[0]),.dinb(w_n336_2[1]),.dout(n383),.clk(gclk));
	jor g0335(.dina(w_n151_2[0]),.dinb(w_n101_2[0]),.dout(n384),.clk(gclk));
	jand g0336(.dina(w_n384_3[1]),.dinb(w_n383_2[2]),.dout(n385),.clk(gclk));
	jand g0337(.dina(w_n385_0[1]),.dinb(w_n382_2[1]),.dout(n386),.clk(gclk));
	jor g0338(.dina(w_n268_1[1]),.dinb(w_n101_1[2]),.dout(n387),.clk(gclk));
	jand g0339(.dina(w_n387_3[1]),.dinb(w_n310_2[1]),.dout(n388),.clk(gclk));
	jor g0340(.dina(w_n127_1[1]),.dinb(w_n336_2[0]),.dout(n389),.clk(gclk));
	jand g0341(.dina(w_n389_3[2]),.dinb(w_n218_3[1]),.dout(n390),.clk(gclk));
	jand g0342(.dina(n390),.dinb(w_n388_1[1]),.dout(n391),.clk(gclk));
	jand g0343(.dina(n391),.dinb(w_n386_0[1]),.dout(n392),.clk(gclk));
	jand g0344(.dina(n392),.dinb(w_n381_0[1]),.dout(n393),.clk(gclk));
	jand g0345(.dina(n393),.dinb(n376),.dout(n394),.clk(gclk));
	jor g0346(.dina(w_n217_3[0]),.dinb(w_n93_0[2]),.dout(n395),.clk(gclk));
	jand g0347(.dina(w_n395_2[2]),.dinb(w_n321_3[0]),.dout(n396),.clk(gclk));
	jand g0348(.dina(w_n396_0[1]),.dinb(w_n255_2[0]),.dout(n397),.clk(gclk));
	jand g0349(.dina(n397),.dinb(w_n309_2[1]),.dout(n398),.clk(gclk));
	jand g0350(.dina(w_n311_2[1]),.dinb(w_n118_5[2]),.dout(n399),.clk(gclk));
	jand g0351(.dina(w_n263_3[1]),.dinb(w_n174_5[2]),.dout(n400),.clk(gclk));
	jor g0352(.dina(w_n400_0[2]),.dinb(w_n399_0[2]),.dout(n401),.clk(gclk));
	jnot g0353(.din(w_n401_0[2]),.dout(n402),.clk(gclk));
	jor g0354(.dina(w_n141_0[0]),.dinb(w_n75_0[2]),.dout(n403),.clk(gclk));
	jor g0355(.dina(w_n403_0[2]),.dinb(w_n77_5[0]),.dout(n404),.clk(gclk));
	jand g0356(.dina(w_n404_1[2]),.dinb(w_n233_2[0]),.dout(n405),.clk(gclk));
	jand g0357(.dina(n405),.dinb(w_n283_2[0]),.dout(n406),.clk(gclk));
	jand g0358(.dina(n406),.dinb(w_n402_0[1]),.dout(n407),.clk(gclk));
	jand g0359(.dina(w_n407_0[1]),.dinb(w_n398_0[2]),.dout(n408),.clk(gclk));
	jor g0360(.dina(w_n165_0[2]),.dinb(w_n125_3[0]),.dout(n409),.clk(gclk));
	jand g0361(.dina(w_n171_3[0]),.dinb(w_n118_5[1]),.dout(n410),.clk(gclk));
	jnot g0362(.din(w_n410_0[1]),.dout(n411),.clk(gclk));
	jand g0363(.dina(w_n411_2[1]),.dinb(w_n409_2[2]),.dout(n412),.clk(gclk));
	jand g0364(.dina(w_n230_2[1]),.dinb(w_n223_2[1]),.dout(n413),.clk(gclk));
	jand g0365(.dina(w_n413_0[1]),.dinb(w_n100_4[2]),.dout(n414),.clk(gclk));
	jnot g0366(.din(n414),.dout(n415),.clk(gclk));
	jand g0367(.dina(w_n415_2[2]),.dinb(w_n286_3[0]),.dout(n416),.clk(gclk));
	jand g0368(.dina(n416),.dinb(n412),.dout(n417),.clk(gclk));
	jor g0369(.dina(w_n249_1[2]),.dinb(w_n101_1[1]),.dout(n418),.clk(gclk));
	jand g0370(.dina(w_n226_2[1]),.dinb(w_n94_2[1]),.dout(n419),.clk(gclk));
	jand g0371(.dina(n419),.dinb(w_n418_2[1]),.dout(n420),.clk(gclk));
	jand g0372(.dina(w_n420_0[1]),.dinb(w_n417_0[2]),.dout(n421),.clk(gclk));
	jand g0373(.dina(n421),.dinb(n408),.dout(n422),.clk(gclk));
	jand g0374(.dina(n422),.dinb(w_n394_0[1]),.dout(n423),.clk(gclk));
	jand g0375(.dina(n423),.dinb(n369),.dout(n424),.clk(gclk));
	jand g0376(.dina(n424),.dinb(w_n359_0[2]),.dout(n425),.clk(gclk));
	jand g0377(.dina(w_n140_1[2]),.dinb(w_n118_5[0]),.dout(n426),.clk(gclk));
	jnot g0378(.din(w_n426_0[2]),.dout(n427),.clk(gclk));
	jand g0379(.dina(w_n411_2[0]),.dinb(w_n120_2[0]),.dout(n428),.clk(gclk));
	jor g0380(.dina(w_n127_1[0]),.dinb(w_n78_2[0]),.dout(n429),.clk(gclk));
	jand g0381(.dina(w_n429_1[2]),.dinb(w_n278_1[1]),.dout(n430),.clk(gclk));
	jand g0382(.dina(w_n430_1[1]),.dinb(n428),.dout(n431),.clk(gclk));
	jand g0383(.dina(n431),.dinb(w_n352_1[0]),.dout(n432),.clk(gclk));
	jand g0384(.dina(w_n311_2[0]),.dinb(w_n174_5[1]),.dout(n433),.clk(gclk));
	jnot g0385(.din(w_n433_0[1]),.dout(n434),.clk(gclk));
	jor g0386(.dina(w_n217_2[2]),.dinb(w_n289_0[1]),.dout(n435),.clk(gclk));
	jand g0387(.dina(w_n435_2[2]),.dinb(w_n434_2[2]),.dout(n436),.clk(gclk));
	jand g0388(.dina(w_n346_2[1]),.dinb(w_n245_2[0]),.dout(n437),.clk(gclk));
	jor g0389(.dina(w_n217_2[1]),.dinb(w_n99_2[1]),.dout(n438),.clk(gclk));
	jor g0390(.dina(w_n336_1[2]),.dinb(w_n99_2[0]),.dout(n439),.clk(gclk));
	jand g0391(.dina(w_n439_4[1]),.dinb(w_n438_2[1]),.dout(n440),.clk(gclk));
	jand g0392(.dina(n440),.dinb(w_n437_1[2]),.dout(n441),.clk(gclk));
	jand g0393(.dina(n441),.dinb(w_n436_0[2]),.dout(n442),.clk(gclk));
	jand g0394(.dina(n442),.dinb(n432),.dout(n443),.clk(gclk));
	jnot g0395(.din(w_n145_1[1]),.dout(n444),.clk(gclk));
	jor g0396(.dina(w_n217_2[0]),.dinb(n444),.dout(n445),.clk(gclk));
	jnot g0397(.din(w_n399_0[1]),.dout(n446),.clk(gclk));
	jand g0398(.dina(w_n174_5[0]),.dinb(w_n140_1[1]),.dout(n447),.clk(gclk));
	jnot g0399(.din(w_n447_0[2]),.dout(n448),.clk(gclk));
	jand g0400(.dina(w_n448_2[1]),.dinb(w_n446_2[1]),.dout(n449),.clk(gclk));
	jand g0401(.dina(n449),.dinb(w_n445_2[2]),.dout(n450),.clk(gclk));
	jand g0402(.dina(n450),.dinb(w_n275_2[0]),.dout(n451),.clk(gclk));
	jand g0403(.dina(n451),.dinb(w_n443_1[1]),.dout(n452),.clk(gclk));
	jand g0404(.dina(w_n452_0[1]),.dinb(w_n427_2[2]),.dout(n453),.clk(gclk));
	jnot g0405(.din(n453),.dout(n454),.clk(gclk));
	jand g0406(.dina(w_n344_3[0]),.dinb(w_n327_1[1]),.dout(n455),.clk(gclk));
	jand g0407(.dina(w_n455_0[1]),.dinb(w_n310_2[0]),.dout(n456),.clk(gclk));
	jnot g0408(.din(w_n301_1[0]),.dout(n457),.clk(gclk));
	jand g0409(.dina(w_n457_0[2]),.dinb(w_n124_2[1]),.dout(n458),.clk(gclk));
	jand g0410(.dina(n458),.dinb(w_n456_0[2]),.dout(n459),.clk(gclk));
	jor g0411(.dina(w_n101_1[0]),.dinb(w_n93_0[1]),.dout(n460),.clk(gclk));
	jand g0412(.dina(w_n460_3[1]),.dinb(w_n418_2[0]),.dout(n461),.clk(gclk));
	jor g0413(.dina(w_n249_1[1]),.dinb(w_n78_1[2]),.dout(n462),.clk(gclk));
	jand g0414(.dina(w_n462_2[1]),.dinb(w_n374_3[0]),.dout(n463),.clk(gclk));
	jand g0415(.dina(w_n463_0[2]),.dinb(w_n461_0[2]),.dout(n464),.clk(gclk));
	jand g0416(.dina(n464),.dinb(w_n459_0[2]),.dout(n465),.clk(gclk));
	jnot g0417(.din(n465),.dout(n466),.clk(gclk));
	jor g0418(.dina(w_n125_2[2]),.dinb(w_n99_1[2]),.dout(n467),.clk(gclk));
	jand g0419(.dina(w_n467_2[2]),.dinb(w_n332_3[0]),.dout(n468),.clk(gclk));
	jnot g0420(.din(w_n468_0[2]),.dout(n469),.clk(gclk));
	jand g0421(.dina(w_n311_1[2]),.dinb(w_n253_6[0]),.dout(n470),.clk(gclk));
	jand g0422(.dina(w_n263_3[0]),.dinb(w_n223_2[0]),.dout(n471),.clk(gclk));
	jor g0423(.dina(n471),.dinb(w_n470_0[2]),.dout(n472),.clk(gclk));
	jor g0424(.dina(n472),.dinb(n469),.dout(n473),.clk(gclk));
	jand g0425(.dina(w_n158_1[1]),.dinb(w_n94_2[0]),.dout(n474),.clk(gclk));
	jand g0426(.dina(w_n415_2[1]),.dinb(w_n267_3[0]),.dout(n475),.clk(gclk));
	jand g0427(.dina(n475),.dinb(w_n213_3[0]),.dout(n476),.clk(gclk));
	jand g0428(.dina(n476),.dinb(n474),.dout(n477),.clk(gclk));
	jnot g0429(.din(w_n477_0[1]),.dout(n478),.clk(gclk));
	jor g0430(.dina(n478),.dinb(n473),.dout(n479),.clk(gclk));
	jor g0431(.dina(n479),.dinb(n466),.dout(n480),.clk(gclk));
	jor g0432(.dina(w_n193_1[0]),.dinb(w_n217_1[2]),.dout(n481),.clk(gclk));
	jand g0433(.dina(w_n481_1[1]),.dinb(w_n218_3[0]),.dout(n482),.clk(gclk));
	jand g0434(.dina(w_n482_0[1]),.dinb(w_n383_2[1]),.dout(n483),.clk(gclk));
	jnot g0435(.din(n483),.dout(n484),.clk(gclk));
	jor g0436(.dina(n484),.dinb(w_n480_0[1]),.dout(n485),.clk(gclk));
	jor g0437(.dina(n485),.dinb(n454),.dout(n486),.clk(gclk));
	jand g0438(.dina(w_n167_3[0]),.dinb(w_n253_5[2]),.dout(n487),.clk(gclk));
	jnot g0439(.din(n487),.dout(n488),.clk(gclk));
	jor g0440(.dina(w_n151_1[2]),.dinb(w_n125_2[1]),.dout(n489),.clk(gclk));
	jand g0441(.dina(w_n489_3[1]),.dinb(w_n353_2[1]),.dout(n490),.clk(gclk));
	jand g0442(.dina(n490),.dinb(w_n488_3[1]),.dout(n491),.clk(gclk));
	jand g0443(.dina(w_n409_2[1]),.dinb(w_n207_2[2]),.dout(n492),.clk(gclk));
	jand g0444(.dina(w_n339_4[0]),.dinb(w_n276_3[1]),.dout(n493),.clk(gclk));
	jand g0445(.dina(n493),.dinb(w_n492_0[1]),.dout(n494),.clk(gclk));
	jand g0446(.dina(w_n130_2[2]),.dinb(w_n184_5[1]),.dout(n495),.clk(gclk));
	jor g0447(.dina(w_n495_0[2]),.dinb(w_n254_0[1]),.dout(n496),.clk(gclk));
	jnot g0448(.din(w_n496_0[1]),.dout(n497),.clk(gclk));
	jand g0449(.dina(w_n497_1[1]),.dinb(w_n382_2[0]),.dout(n498),.clk(gclk));
	jand g0450(.dina(n498),.dinb(n494),.dout(n499),.clk(gclk));
	jand g0451(.dina(n499),.dinb(w_n491_0[1]),.dout(n500),.clk(gclk));
	jand g0452(.dina(w_n430_1[0]),.dinb(w_n351_1[0]),.dout(n501),.clk(gclk));
	jand g0453(.dina(n501),.dinb(w_n500_0[1]),.dout(n502),.clk(gclk));
	jnot g0454(.din(n502),.dout(n503),.clk(gclk));
	jor g0455(.dina(n503),.dinb(w_n480_0[0]),.dout(n504),.clk(gclk));
	jand g0456(.dina(w_n366_3[0]),.dinb(w_n331_2[1]),.dout(n505),.clk(gclk));
	jor g0457(.dina(w_n231_0[1]),.dinb(w_n125_2[0]),.dout(n506),.clk(gclk));
	jand g0458(.dina(w_n506_2[2]),.dinb(w_n333_2[0]),.dout(n507),.clk(gclk));
	jand g0459(.dina(n507),.dinb(w_n114_3[1]),.dout(n508),.clk(gclk));
	jand g0460(.dina(n508),.dinb(w_n505_0[1]),.dout(n509),.clk(gclk));
	jor g0461(.dina(w_n125_1[2]),.dinb(w_n113_1[1]),.dout(n510),.clk(gclk));
	jand g0462(.dina(w_n244_3[0]),.dinb(w_n187_2[0]),.dout(n511),.clk(gclk));
	jand g0463(.dina(n511),.dinb(w_n510_3[1]),.dout(n512),.clk(gclk));
	jand g0464(.dina(n512),.dinb(w_n509_0[1]),.dout(n513),.clk(gclk));
	jand g0465(.dina(w_n513_0[2]),.dinb(w_n128_3[0]),.dout(n514),.clk(gclk));
	jnot g0466(.din(w_n514_0[1]),.dout(n515),.clk(gclk));
	jor g0467(.dina(n515),.dinb(w_n504_0[1]),.dout(n516),.clk(gclk));
	jxor g0468(.dina(w_n516_0[2]),.dinb(w_n486_1[2]),.dout(n517),.clk(gclk));
	jand g0469(.dina(w_n51_0[0]),.dinb(w_n49_7[1]),.dout(n518),.clk(gclk));
	jxor g0470(.dina(n518),.dinb(w_a3_0[0]),.dout(n519),.clk(gclk));
	jand g0471(.dina(w_n519_5[2]),.dinb(w_n517_0[2]),.dout(n520),.clk(gclk));
	jnot g0472(.din(n520),.dout(n521),.clk(gclk));
	jand g0473(.dina(w_n388_1[0]),.dinb(w_n250_2[0]),.dout(n522),.clk(gclk));
	jand g0474(.dina(w_n253_5[1]),.dinb(w_n116_2[2]),.dout(n523),.clk(gclk));
	jor g0475(.dina(w_n172_0[0]),.dinb(w_n523_0[1]),.dout(n524),.clk(gclk));
	jnot g0476(.din(w_n524_0[1]),.dout(n525),.clk(gclk));
	jor g0477(.dina(w_n151_1[1]),.dinb(w_n216_0[0]),.dout(n526),.clk(gclk));
	jor g0478(.dina(w_n526_0[1]),.dinb(w_n77_4[2]),.dout(n527),.clk(gclk));
	jand g0479(.dina(w_n527_3[2]),.dinb(w_n445_2[1]),.dout(n528),.clk(gclk));
	jand g0480(.dina(w_n528_0[1]),.dinb(w_n525_0[1]),.dout(n529),.clk(gclk));
	jand g0481(.dina(n529),.dinb(w_n522_0[1]),.dout(n530),.clk(gclk));
	jand g0482(.dina(w_n333_1[2]),.dinb(w_n147_2[0]),.dout(n531),.clk(gclk));
	jand g0483(.dina(w_n531_0[1]),.dinb(w_n294_3[0]),.dout(n532),.clk(gclk));
	jand g0484(.dina(w_n532_0[1]),.dinb(w_n530_0[1]),.dout(n533),.clk(gclk));
	jor g0485(.dina(w_n99_1[1]),.dinb(w_n78_1[1]),.dout(n534),.clk(gclk));
	jor g0486(.dina(w_n249_1[0]),.dinb(w_n135_1[2]),.dout(n535),.clk(gclk));
	jand g0487(.dina(w_n191_3[0]),.dinb(w_n182_3[0]),.dout(n536),.clk(gclk));
	jand g0488(.dina(n536),.dinb(w_n535_2[1]),.dout(n537),.clk(gclk));
	jand g0489(.dina(w_n537_0[1]),.dinb(w_n534_2[2]),.dout(n538),.clk(gclk));
	jand g0490(.dina(w_n384_3[0]),.dinb(w_n235_2[0]),.dout(n539),.clk(gclk));
	jand g0491(.dina(w_n506_2[1]),.dinb(w_n207_2[1]),.dout(n540),.clk(gclk));
	jand g0492(.dina(w_n540_0[2]),.dinb(w_n539_1[2]),.dout(n541),.clk(gclk));
	jand g0493(.dina(n541),.dinb(w_n267_2[2]),.dout(n542),.clk(gclk));
	jand g0494(.dina(n542),.dinb(n538),.dout(n543),.clk(gclk));
	jor g0495(.dina(w_n495_0[1]),.dinb(w_n312_0[0]),.dout(n544),.clk(gclk));
	jnot g0496(.din(w_n544_0[1]),.dout(n545),.clk(gclk));
	jand g0497(.dina(w_n382_1[2]),.dinb(w_n204_2[1]),.dout(n546),.clk(gclk));
	jand g0498(.dina(w_n546_0[2]),.dinb(w_n133_1[2]),.dout(n547),.clk(gclk));
	jand g0499(.dina(n547),.dinb(n545),.dout(n548),.clk(gclk));
	jand g0500(.dina(n548),.dinb(w_n407_0[0]),.dout(n549),.clk(gclk));
	jand g0501(.dina(n549),.dinb(w_n543_0[1]),.dout(n550),.clk(gclk));
	jand g0502(.dina(n550),.dinb(n533),.dout(n551),.clk(gclk));
	jand g0503(.dina(w_n331_2[0]),.dinb(w_n114_3[0]),.dout(n552),.clk(gclk));
	jand g0504(.dina(w_n112_3[1]),.dinb(w_n262_4[1]),.dout(n553),.clk(gclk));
	jor g0505(.dina(w_n433_0[0]),.dinb(w_n553_0[1]),.dout(n554),.clk(gclk));
	jor g0506(.dina(n554),.dinb(w_n296_0[0]),.dout(n555),.clk(gclk));
	jnot g0507(.din(w_n555_0[1]),.dout(n556),.clk(gclk));
	jand g0508(.dina(w_n269_2[0]),.dinb(w_n252_4[0]),.dout(n557),.clk(gclk));
	jand g0509(.dina(w_n395_2[1]),.dinb(w_n160_2[1]),.dout(n558),.clk(gclk));
	jand g0510(.dina(n558),.dinb(w_n557_0[1]),.dout(n559),.clk(gclk));
	jand g0511(.dina(w_n559_0[1]),.dinb(n556),.dout(n560),.clk(gclk));
	jor g0512(.dina(w_n268_1[0]),.dinb(w_n336_1[1]),.dout(n561),.clk(gclk));
	jand g0513(.dina(w_n561_1[1]),.dinb(w_n321_2[2]),.dout(n562),.clk(gclk));
	jand g0514(.dina(w_n562_1[1]),.dinb(w_n197_3[0]),.dout(n563),.clk(gclk));
	jand g0515(.dina(w_n563_0[1]),.dinb(w_n560_0[1]),.dout(n564),.clk(gclk));
	jand g0516(.dina(n564),.dinb(w_n552_0[2]),.dout(n565),.clk(gclk));
	jand g0517(.dina(n565),.dinb(w_n551_0[1]),.dout(n566),.clk(gclk));
	jand g0518(.dina(w_n370_3[0]),.dinb(w_n303_0[1]),.dout(n567),.clk(gclk));
	jand g0519(.dina(w_n567_0[1]),.dinb(w_n245_1[2]),.dout(n568),.clk(gclk));
	jor g0520(.dina(w_n135_1[1]),.dinb(w_n113_1[0]),.dout(n569),.clk(gclk));
	jor g0521(.dina(w_n193_0[2]),.dinb(w_n336_1[0]),.dout(n570),.clk(gclk));
	jand g0522(.dina(w_n570_2[1]),.dinb(w_n569_2[1]),.dout(n571),.clk(gclk));
	jand g0523(.dina(n571),.dinb(w_n136_2[0]),.dout(n572),.clk(gclk));
	jand g0524(.dina(w_n572_0[1]),.dinb(w_n102_3[0]),.dout(n573),.clk(gclk));
	jand g0525(.dina(n573),.dinb(w_n568_0[2]),.dout(n574),.clk(gclk));
	jand g0526(.dina(w_n194_0[1]),.dinb(w_n152_2[1]),.dout(n575),.clk(gclk));
	jnot g0527(.din(w_n575_0[1]),.dout(n576),.clk(gclk));
	jand g0528(.dina(w_n230_2[0]),.dinb(w_n118_4[2]),.dout(n577),.clk(gclk));
	jor g0529(.dina(w_n577_0[1]),.dinb(w_n205_0[0]),.dout(n578),.clk(gclk));
	jand g0530(.dina(w_n118_4[1]),.dinb(w_n98_3[0]),.dout(n579),.clk(gclk));
	jor g0531(.dina(w_n579_0[1]),.dinb(w_n254_0[0]),.dout(n580),.clk(gclk));
	jor g0532(.dina(n580),.dinb(n578),.dout(n581),.clk(gclk));
	jor g0533(.dina(n581),.dinb(n576),.dout(n582),.clk(gclk));
	jnot g0534(.din(w_n582_0[1]),.dout(n583),.clk(gclk));
	jand g0535(.dina(w_n481_1[0]),.dinb(w_n462_2[0]),.dout(n584),.clk(gclk));
	jand g0536(.dina(w_n467_2[1]),.dinb(w_n383_2[0]),.dout(n585),.clk(gclk));
	jand g0537(.dina(n585),.dinb(n584),.dout(n586),.clk(gclk));
	jor g0538(.dina(w_n151_1[0]),.dinb(w_n78_1[0]),.dout(n587),.clk(gclk));
	jand g0539(.dina(w_n587_3[1]),.dinb(w_n166_2[1]),.dout(n588),.clk(gclk));
	jand g0540(.dina(w_n232_4[1]),.dinb(w_n128_2[2]),.dout(n589),.clk(gclk));
	jand g0541(.dina(n589),.dinb(w_n588_0[2]),.dout(n590),.clk(gclk));
	jand g0542(.dina(n590),.dinb(w_n586_0[2]),.dout(n591),.clk(gclk));
	jand g0543(.dina(w_n438_2[0]),.dinb(w_n244_2[2]),.dout(n592),.clk(gclk));
	jand g0544(.dina(n592),.dinb(w_n248_3[1]),.dout(n593),.clk(gclk));
	jand g0545(.dina(w_n409_2[0]),.dinb(w_n290_3[1]),.dout(n594),.clk(gclk));
	jand g0546(.dina(w_n594_0[2]),.dinb(w_n378_3[0]),.dout(n595),.clk(gclk));
	jand g0547(.dina(n595),.dinb(w_n593_0[1]),.dout(n596),.clk(gclk));
	jand g0548(.dina(n596),.dinb(n591),.dout(n597),.clk(gclk));
	jand g0549(.dina(n597),.dinb(w_n583_0[1]),.dout(n598),.clk(gclk));
	jand g0550(.dina(w_n185_3[0]),.dinb(w_n118_4[0]),.dout(n599),.clk(gclk));
	jnot g0551(.din(w_n599_0[1]),.dout(n600),.clk(gclk));
	jand g0552(.dina(w_n600_2[2]),.dinb(w_n418_1[2]),.dout(n601),.clk(gclk));
	jand g0553(.dina(w_n309_2[0]),.dinb(w_n236_1[0]),.dout(n602),.clk(gclk));
	jand g0554(.dina(w_n602_0[1]),.dinb(w_n305_2[0]),.dout(n603),.clk(gclk));
	jand g0555(.dina(w_n603_0[1]),.dinb(w_n601_0[1]),.dout(n604),.clk(gclk));
	jand g0556(.dina(w_n604_0[1]),.dinb(w_n598_0[1]),.dout(n605),.clk(gclk));
	jand g0557(.dina(n605),.dinb(w_n574_0[1]),.dout(n606),.clk(gclk));
	jand g0558(.dina(n606),.dinb(n566),.dout(n607),.clk(gclk));
	jnot g0559(.din(w_n417_0[1]),.dout(n608),.clk(gclk));
	jand g0560(.dina(w_n192_3[0]),.dinb(w_n154_5[1]),.dout(n609),.clk(gclk));
	jand g0561(.dina(w_n154_5[0]),.dinb(w_n98_2[2]),.dout(n610),.clk(gclk));
	jor g0562(.dina(w_n610_0[1]),.dinb(w_n609_0[1]),.dout(n611),.clk(gclk));
	jand g0563(.dina(w_n144_5[2]),.dinb(w_n92_2[1]),.dout(n612),.clk(gclk));
	jand g0564(.dina(w_n144_5[1]),.dinb(w_n112_3[0]),.dout(n613),.clk(gclk));
	jor g0565(.dina(w_n613_0[1]),.dinb(w_n612_0[1]),.dout(n614),.clk(gclk));
	jor g0566(.dina(n614),.dinb(n611),.dout(n615),.clk(gclk));
	jor g0567(.dina(n615),.dinb(w_n360_0[1]),.dout(n616),.clk(gclk));
	jand g0568(.dina(w_n144_5[0]),.dinb(w_n98_2[1]),.dout(n617),.clk(gclk));
	jand g0569(.dina(w_n116_2[1]),.dinb(w_n184_5[0]),.dout(n618),.clk(gclk));
	jand g0570(.dina(w_n126_4[0]),.dinb(w_n253_5[0]),.dout(n619),.clk(gclk));
	jor g0571(.dina(w_n619_0[1]),.dinb(n618),.dout(n620),.clk(gclk));
	jor g0572(.dina(w_n266_1[1]),.dinb(n620),.dout(n621),.clk(gclk));
	jor g0573(.dina(n621),.dinb(w_n617_0[2]),.dout(n622),.clk(gclk));
	jor g0574(.dina(n622),.dinb(w_n616_0[1]),.dout(n623),.clk(gclk));
	jand g0575(.dina(w_n116_2[0]),.dinb(w_n223_1[2]),.dout(n624),.clk(gclk));
	jand g0576(.dina(w_n624_0[2]),.dinb(w_n100_4[1]),.dout(n625),.clk(gclk));
	jand g0577(.dina(w_n263_2[2]),.dinb(w_n224_4[1]),.dout(n626),.clk(gclk));
	jor g0578(.dina(n626),.dinb(w_n625_0[1]),.dout(n627),.clk(gclk));
	jor g0579(.dina(n627),.dinb(w_n599_0[0]),.dout(n628),.clk(gclk));
	jor g0580(.dina(w_n628_0[1]),.dinb(w_n447_0[1]),.dout(n629),.clk(gclk));
	jand g0581(.dina(w_n167_2[2]),.dinb(w_n262_4[0]),.dout(n630),.clk(gclk));
	jand g0582(.dina(w_n184_4[2]),.dinb(w_n92_2[0]),.dout(n631),.clk(gclk));
	jor g0583(.dina(n631),.dinb(w_n630_0[2]),.dout(n632),.clk(gclk));
	jor g0584(.dina(n632),.dinb(w_n330_0[1]),.dout(n633),.clk(gclk));
	jand g0585(.dina(w_n130_2[1]),.dinb(w_n262_3[2]),.dout(n634),.clk(gclk));
	jor g0586(.dina(w_n634_0[2]),.dinb(n633),.dout(n635),.clk(gclk));
	jor g0587(.dina(n635),.dinb(n629),.dout(n636),.clk(gclk));
	jor g0588(.dina(n636),.dinb(n623),.dout(n637),.clk(gclk));
	jor g0589(.dina(n637),.dinb(n608),.dout(n638),.clk(gclk));
	jand g0590(.dina(w_n174_4[2]),.dinb(w_n116_1[2]),.dout(n639),.clk(gclk));
	jand g0591(.dina(w_n112_2[2]),.dinb(w_n184_4[1]),.dout(n640),.clk(gclk));
	jor g0592(.dina(w_n295_0[1]),.dinb(n640),.dout(n641),.clk(gclk));
	jor g0593(.dina(n641),.dinb(n639),.dout(n642),.clk(gclk));
	jor g0594(.dina(n642),.dinb(w_n301_0[2]),.dout(n643),.clk(gclk));
	jor g0595(.dina(n643),.dinb(w_n212_0[0]),.dout(n644),.clk(gclk));
	jand g0596(.dina(w_n413_0[0]),.dinb(w_n77_4[1]),.dout(n645),.clk(gclk));
	jand g0597(.dina(w_n185_2[2]),.dinb(w_n262_3[1]),.dout(n646),.clk(gclk));
	jor g0598(.dina(w_n646_0[1]),.dinb(w_n645_0[1]),.dout(n647),.clk(gclk));
	jand g0599(.dina(w_n185_2[1]),.dinb(w_n253_4[2]),.dout(n648),.clk(gclk));
	jor g0600(.dina(w_n495_0[0]),.dinb(w_n648_0[1]),.dout(n649),.clk(gclk));
	jor g0601(.dina(n649),.dinb(n647),.dout(n650),.clk(gclk));
	jand g0602(.dina(w_n311_1[1]),.dinb(w_n262_3[0]),.dout(n651),.clk(gclk));
	jand g0603(.dina(w_n263_2[1]),.dinb(w_n154_4[2]),.dout(n652),.clk(gclk));
	jor g0604(.dina(w_n652_0[2]),.dinb(n651),.dout(n653),.clk(gclk));
	jand g0605(.dina(w_n171_2[2]),.dinb(w_n154_4[1]),.dout(n654),.clk(gclk));
	jand g0606(.dina(w_n192_2[2]),.dinb(w_n174_4[1]),.dout(n655),.clk(gclk));
	jor g0607(.dina(w_n655_0[1]),.dinb(w_n654_0[2]),.dout(n656),.clk(gclk));
	jor g0608(.dina(n656),.dinb(w_n400_0[1]),.dout(n657),.clk(gclk));
	jor g0609(.dina(n657),.dinb(n653),.dout(n658),.clk(gclk));
	jor g0610(.dina(n658),.dinb(n650),.dout(n659),.clk(gclk));
	jand g0611(.dina(w_n167_2[1]),.dinb(w_n184_4[0]),.dout(n660),.clk(gclk));
	jor g0612(.dina(w_n660_0[1]),.dinb(w_n470_0[1]),.dout(n661),.clk(gclk));
	jand g0613(.dina(w_n174_4[0]),.dinb(w_n126_3[2]),.dout(n662),.clk(gclk));
	jand g0614(.dina(w_n185_2[0]),.dinb(w_n224_4[0]),.dout(n663),.clk(gclk));
	jor g0615(.dina(w_n663_0[1]),.dinb(n662),.dout(n664),.clk(gclk));
	jor g0616(.dina(n664),.dinb(w_n661_0[1]),.dout(n665),.clk(gclk));
	jand g0617(.dina(w_n311_1[0]),.dinb(w_n143_0[2]),.dout(n666),.clk(gclk));
	jand g0618(.dina(w_n666_0[1]),.dinb(w_n100_4[0]),.dout(n667),.clk(gclk));
	jor g0619(.dina(w_n667_0[1]),.dinb(w_n553_0[0]),.dout(n668),.clk(gclk));
	jand g0620(.dina(w_n311_0[2]),.dinb(w_n184_3[2]),.dout(n669),.clk(gclk));
	jor g0621(.dina(w_n669_0[1]),.dinb(n668),.dout(n670),.clk(gclk));
	jor g0622(.dina(n670),.dinb(n665),.dout(n671),.clk(gclk));
	jand g0623(.dina(w_n154_4[0]),.dinb(w_n130_2[0]),.dout(n672),.clk(gclk));
	jand g0624(.dina(w_n174_3[2]),.dinb(w_n145_1[0]),.dout(n673),.clk(gclk));
	jor g0625(.dina(w_n673_0[1]),.dinb(n672),.dout(n674),.clk(gclk));
	jand g0626(.dina(w_n192_2[1]),.dinb(w_n184_3[1]),.dout(n675),.clk(gclk));
	jand g0627(.dina(w_n112_2[1]),.dinb(w_n224_3[2]),.dout(n676),.clk(gclk));
	jand g0628(.dina(w_n155_3[0]),.dinb(w_n262_2[2]),.dout(n677),.clk(gclk));
	jor g0629(.dina(w_n677_1[1]),.dinb(w_n676_0[2]),.dout(n678),.clk(gclk));
	jor g0630(.dina(n678),.dinb(n675),.dout(n679),.clk(gclk));
	jor g0631(.dina(n679),.dinb(n674),.dout(n680),.clk(gclk));
	jor g0632(.dina(n680),.dinb(n671),.dout(n681),.clk(gclk));
	jor g0633(.dina(n681),.dinb(n659),.dout(n682),.clk(gclk));
	jor g0634(.dina(n682),.dinb(w_n644_0[1]),.dout(n683),.clk(gclk));
	jand g0635(.dina(w_n131_0[0]),.dinb(w_n100_3[2]),.dout(n684),.clk(gclk));
	jand g0636(.dina(w_n185_1[2]),.dinb(w_n154_3[2]),.dout(n685),.clk(gclk));
	jand g0637(.dina(w_n154_3[1]),.dinb(w_n112_2[0]),.dout(n686),.clk(gclk));
	jor g0638(.dina(w_n686_0[1]),.dinb(w_n685_0[1]),.dout(n687),.clk(gclk));
	jor g0639(.dina(n687),.dinb(w_n684_0[2]),.dout(n688),.clk(gclk));
	jand g0640(.dina(w_n155_2[2]),.dinb(w_n224_3[1]),.dout(n689),.clk(gclk));
	jand g0641(.dina(w_n263_2[0]),.dinb(w_n118_3[2]),.dout(n690),.clk(gclk));
	jor g0642(.dina(w_n690_0[1]),.dinb(w_n689_0[2]),.dout(n691),.clk(gclk));
	jor g0643(.dina(n691),.dinb(w_n314_0[1]),.dout(n692),.clk(gclk));
	jor g0644(.dina(n692),.dinb(n688),.dout(n693),.clk(gclk));
	jand g0645(.dina(w_n185_1[1]),.dinb(w_n174_3[1]),.dout(n694),.clk(gclk));
	jand g0646(.dina(w_n167_2[0]),.dinb(w_n118_3[1]),.dout(n695),.clk(gclk));
	jor g0647(.dina(n695),.dinb(n694),.dout(n696),.clk(gclk));
	jand g0648(.dina(w_n143_0[1]),.dinb(w_n126_3[1]),.dout(n697),.clk(gclk));
	jor g0649(.dina(w_n697_0[1]),.dinb(w_n579_0[0]),.dout(n698),.clk(gclk));
	jor g0650(.dina(n698),.dinb(n696),.dout(n699),.clk(gclk));
	jand g0651(.dina(w_n174_3[0]),.dinb(w_n155_2[1]),.dout(n700),.clk(gclk));
	jand g0652(.dina(w_n118_3[0]),.dinb(w_n112_1[2]),.dout(n701),.clk(gclk));
	jor g0653(.dina(n701),.dinb(w_n700_0[1]),.dout(n702),.clk(gclk));
	jor g0654(.dina(w_n702_0[1]),.dinb(n699),.dout(n703),.clk(gclk));
	jor g0655(.dina(n703),.dinb(n693),.dout(n704),.clk(gclk));
	jand g0656(.dina(w_n171_2[1]),.dinb(w_n253_4[1]),.dout(n705),.clk(gclk));
	jand g0657(.dina(w_n624_0[1]),.dinb(w_n77_4[0]),.dout(n706),.clk(gclk));
	jand g0658(.dina(w_n167_1[2]),.dinb(w_n144_4[2]),.dout(n707),.clk(gclk));
	jand g0659(.dina(w_n192_2[0]),.dinb(w_n223_1[1]),.dout(n708),.clk(gclk));
	jand g0660(.dina(w_n708_0[1]),.dinb(w_n77_3[2]),.dout(n709),.clk(gclk));
	jor g0661(.dina(n709),.dinb(n707),.dout(n710),.clk(gclk));
	jor g0662(.dina(n710),.dinb(w_n186_0[0]),.dout(n711),.clk(gclk));
	jor g0663(.dina(n711),.dinb(w_n706_0[1]),.dout(n712),.clk(gclk));
	jor g0664(.dina(n712),.dinb(w_n705_0[2]),.dout(n713),.clk(gclk));
	jor g0665(.dina(n713),.dinb(n704),.dout(n714),.clk(gclk));
	jor g0666(.dina(n714),.dinb(n683),.dout(n715),.clk(gclk));
	jor g0667(.dina(n715),.dinb(n638),.dout(n716),.clk(gclk));
	jor g0668(.dina(w_n194_0[0]),.dinb(w_n100_3[1]),.dout(n717),.clk(gclk));
	jand g0669(.dina(w_n171_2[0]),.dinb(w_n223_1[0]),.dout(n718),.clk(gclk));
	jor g0670(.dina(n718),.dinb(w_n673_0[0]),.dout(n719),.clk(gclk));
	jnot g0671(.din(n719),.dout(n720),.clk(gclk));
	jand g0672(.dina(w_n720_0[1]),.dinb(w_n717_3[1]),.dout(n721),.clk(gclk));
	jand g0673(.dina(w_n240_2[0]),.dinb(w_n197_2[2]),.dout(n722),.clk(gclk));
	jand g0674(.dina(n722),.dinb(n721),.dout(n723),.clk(gclk));
	jnot g0675(.din(w_n723_0[1]),.dout(n724),.clk(gclk));
	jor g0676(.dina(w_n399_0[0]),.dinb(w_n282_1[1]),.dout(n725),.clk(gclk));
	jand g0677(.dina(w_n263_1[2]),.dinb(w_n144_4[1]),.dout(n726),.clk(gclk));
	jand g0678(.dina(w_n98_2[0]),.dinb(w_n262_2[1]),.dout(n727),.clk(gclk));
	jor g0679(.dina(w_n727_0[1]),.dinb(n726),.dout(n728),.clk(gclk));
	jand g0680(.dina(w_n174_2[2]),.dinb(w_n92_1[2]),.dout(n729),.clk(gclk));
	jor g0681(.dina(w_n684_0[1]),.dinb(n729),.dout(n730),.clk(gclk));
	jor g0682(.dina(n730),.dinb(n728),.dout(n731),.clk(gclk));
	jor g0683(.dina(n731),.dinb(w_n725_0[1]),.dout(n732),.clk(gclk));
	jor g0684(.dina(w_n630_0[1]),.dinb(w_n652_0[1]),.dout(n733),.clk(gclk));
	jor g0685(.dina(n733),.dinb(w_n299_0[0]),.dout(n734),.clk(gclk));
	jor g0686(.dina(n734),.dinb(w_n677_1[0]),.dout(n735),.clk(gclk));
	jor g0687(.dina(n735),.dinb(n732),.dout(n736),.clk(gclk));
	jand g0688(.dina(w_n708_0[0]),.dinb(w_n100_3[0]),.dout(n737),.clk(gclk));
	jor g0689(.dina(n737),.dinb(w_n706_0[0]),.dout(n738),.clk(gclk));
	jor g0690(.dina(n738),.dinb(w_n426_0[1]),.dout(n739),.clk(gclk));
	jor g0691(.dina(n739),.dinb(w_n400_0[0]),.dout(n740),.clk(gclk));
	jand g0692(.dina(w_n126_3[0]),.dinb(w_n224_3[0]),.dout(n741),.clk(gclk));
	jor g0693(.dina(w_n676_0[1]),.dinb(n741),.dout(n742),.clk(gclk));
	jor g0694(.dina(w_n690_0[0]),.dinb(n742),.dout(n743),.clk(gclk));
	jor g0695(.dina(w_n308_0[0]),.dinb(w_n132_0[1]),.dout(n744),.clk(gclk));
	jor g0696(.dina(w_n744_0[1]),.dinb(n743),.dout(n745),.clk(gclk));
	jor g0697(.dina(n745),.dinb(n740),.dout(n746),.clk(gclk));
	jor g0698(.dina(n746),.dinb(n736),.dout(n747),.clk(gclk));
	jor g0699(.dina(n747),.dinb(n724),.dout(n748),.clk(gclk));
	jand g0700(.dina(w_n154_3[0]),.dinb(w_n126_2[2]),.dout(n749),.clk(gclk));
	jand g0701(.dina(w_n130_1[2]),.dinb(w_n224_2[2]),.dout(n750),.clk(gclk));
	jor g0702(.dina(n750),.dinb(w_n749_0[1]),.dout(n751),.clk(gclk));
	jand g0703(.dina(w_n144_4[0]),.dinb(w_n116_1[1]),.dout(n752),.clk(gclk));
	jand g0704(.dina(w_n126_2[1]),.dinb(w_n118_2[2]),.dout(n753),.clk(gclk));
	jor g0705(.dina(n753),.dinb(w_n752_0[2]),.dout(n754),.clk(gclk));
	jor g0706(.dina(n754),.dinb(w_n617_0[1]),.dout(n755),.clk(gclk));
	jor g0707(.dina(n755),.dinb(w_n751_0[1]),.dout(n756),.clk(gclk));
	jor g0708(.dina(n756),.dinb(w_n264_0[0]),.dout(n757),.clk(gclk));
	jand g0709(.dina(w_n154_2[2]),.dinb(w_n116_1[0]),.dout(n758),.clk(gclk));
	jand g0710(.dina(w_n192_1[2]),.dinb(w_n118_2[1]),.dout(n759),.clk(gclk));
	jor g0711(.dina(n759),.dinb(w_n686_0[0]),.dout(n760),.clk(gclk));
	jor g0712(.dina(n760),.dinb(n758),.dout(n761),.clk(gclk));
	jand g0713(.dina(w_n140_1[0]),.dinb(w_n144_3[2]),.dout(n762),.clk(gclk));
	jand g0714(.dina(w_n155_2[0]),.dinb(w_n184_3[0]),.dout(n763),.clk(gclk));
	jor g0715(.dina(n763),.dinb(n762),.dout(n764),.clk(gclk));
	jor g0716(.dina(n764),.dinb(n761),.dout(n765),.clk(gclk));
	jand g0717(.dina(w_n230_1[2]),.dinb(w_n253_4[0]),.dout(n766),.clk(gclk));
	jand g0718(.dina(w_n174_2[1]),.dinb(w_n171_1[2]),.dout(n767),.clk(gclk));
	jand g0719(.dina(w_n144_3[1]),.dinb(w_n130_1[1]),.dout(n768),.clk(gclk));
	jor g0720(.dina(w_n609_0[0]),.dinb(n768),.dout(n769),.clk(gclk));
	jor g0721(.dina(n769),.dinb(n767),.dout(n770),.clk(gclk));
	jor g0722(.dina(n770),.dinb(w_n766_0[1]),.dout(n771),.clk(gclk));
	jor g0723(.dina(n771),.dinb(n765),.dout(n772),.clk(gclk));
	jor g0724(.dina(n772),.dinb(n757),.dout(n773),.clk(gclk));
	jand g0725(.dina(w_n666_0[0]),.dinb(w_n77_3[1]),.dout(n774),.clk(gclk));
	jor g0726(.dina(w_n689_0[1]),.dinb(n774),.dout(n775),.clk(gclk));
	jor g0727(.dina(n775),.dinb(w_n610_0[0]),.dout(n776),.clk(gclk));
	jand g0728(.dina(w_n167_1[1]),.dinb(w_n154_2[1]),.dout(n777),.clk(gclk));
	jand g0729(.dina(w_n224_2[1]),.dinb(w_n92_1[1]),.dout(n778),.clk(gclk));
	jor g0730(.dina(n778),.dinb(w_n663_0[0]),.dout(n779),.clk(gclk));
	jor g0731(.dina(n779),.dinb(w_n777_0[2]),.dout(n780),.clk(gclk));
	jor g0732(.dina(n780),.dinb(w_n702_0[0]),.dout(n781),.clk(gclk));
	jor g0733(.dina(n781),.dinb(n776),.dout(n782),.clk(gclk));
	jor g0734(.dina(n782),.dinb(w_n644_0[0]),.dout(n783),.clk(gclk));
	jor g0735(.dina(n783),.dinb(n773),.dout(n784),.clk(gclk));
	jor g0736(.dina(w_n410_0[0]),.dinb(w_n266_1[0]),.dout(n785),.clk(gclk));
	jor g0737(.dina(w_n785_0[1]),.dinb(w_n496_0[0]),.dout(n786),.clk(gclk));
	jnot g0738(.din(w_n170_3[0]),.dout(n787),.clk(gclk));
	jand g0739(.dina(w_n171_1[1]),.dinb(w_n184_2[2]),.dout(n788),.clk(gclk));
	jor g0740(.dina(w_n669_0[0]),.dinb(w_n788_0[1]),.dout(n789),.clk(gclk));
	jor g0741(.dina(n789),.dinb(w_n705_0[1]),.dout(n790),.clk(gclk));
	jor g0742(.dina(n790),.dinb(w_n787_0[1]),.dout(n791),.clk(gclk));
	jor g0743(.dina(n791),.dinb(w_n786_0[1]),.dout(n792),.clk(gclk));
	jand g0744(.dina(w_n126_2[0]),.dinb(w_n184_2[1]),.dout(n793),.clk(gclk));
	jor g0745(.dina(w_n645_0[0]),.dinb(n793),.dout(n794),.clk(gclk));
	jand g0746(.dina(w_n130_1[0]),.dinb(w_n253_3[2]),.dout(n795),.clk(gclk));
	jand g0747(.dina(w_n253_3[1]),.dinb(w_n112_1[1]),.dout(n796),.clk(gclk));
	jor g0748(.dina(w_n796_0[1]),.dinb(n795),.dout(n797),.clk(gclk));
	jand g0749(.dina(w_n263_1[1]),.dinb(w_n253_3[0]),.dout(n798),.clk(gclk));
	jor g0750(.dina(w_n648_0[0]),.dinb(n798),.dout(n799),.clk(gclk));
	jor g0751(.dina(n799),.dinb(n797),.dout(n800),.clk(gclk));
	jor g0752(.dina(n800),.dinb(n794),.dout(n801),.clk(gclk));
	jand g0753(.dina(w_n230_1[1]),.dinb(w_n154_2[0]),.dout(n802),.clk(gclk));
	jor g0754(.dina(w_n330_0[0]),.dinb(w_n802_0[1]),.dout(n803),.clk(gclk));
	jor g0755(.dina(w_n803_0[1]),.dinb(n801),.dout(n804),.clk(gclk));
	jor g0756(.dina(w_n613_0[0]),.dinb(w_n470_0[0]),.dout(n805),.clk(gclk));
	jand g0757(.dina(w_n144_3[0]),.dinb(w_n126_1[2]),.dout(n806),.clk(gclk));
	jor g0758(.dina(n806),.dinb(w_n523_0[0]),.dout(n807),.clk(gclk));
	jor g0759(.dina(n807),.dinb(n805),.dout(n808),.clk(gclk));
	jor g0760(.dina(n808),.dinb(w_n146_0[0]),.dout(n809),.clk(gclk));
	jor g0761(.dina(n809),.dinb(n804),.dout(n810),.clk(gclk));
	jor g0762(.dina(n810),.dinb(n792),.dout(n811),.clk(gclk));
	jor g0763(.dina(n811),.dinb(n784),.dout(n812),.clk(gclk));
	jor g0764(.dina(n812),.dinb(n748),.dout(n813),.clk(gclk));
	jand g0765(.dina(w_n813_0[1]),.dinb(w_n716_8[2]),.dout(n814),.clk(gclk));
	jor g0766(.dina(w_n814_0[1]),.dinb(w_n607_2[1]),.dout(n815),.clk(gclk));
	jnot g0767(.din(w_n725_0[0]),.dout(n816),.clk(gclk));
	jand g0768(.dina(w_n534_2[1]),.dinb(w_n347_2[1]),.dout(n817),.clk(gclk));
	jand g0769(.dina(w_n527_3[1]),.dinb(w_n395_2[0]),.dout(n818),.clk(gclk));
	jand g0770(.dina(n818),.dinb(w_n817_1[2]),.dout(n819),.clk(gclk));
	jand g0771(.dina(n819),.dinb(w_n816_0[1]),.dout(n820),.clk(gclk));
	jand g0772(.dina(w_n332_2[2]),.dinb(w_n269_1[2]),.dout(n821),.clk(gclk));
	jand g0773(.dina(n821),.dinb(w_n300_3[0]),.dout(n822),.clk(gclk));
	jand g0774(.dina(n822),.dinb(w_n378_2[2]),.dout(n823),.clk(gclk));
	jand g0775(.dina(n823),.dinb(n820),.dout(n824),.clk(gclk));
	jor g0776(.dina(w_n268_0[2]),.dinb(w_n217_1[1]),.dout(n825),.clk(gclk));
	jand g0777(.dina(w_n195_1[2]),.dinb(w_n160_2[0]),.dout(n826),.clk(gclk));
	jand g0778(.dina(w_n826_0[1]),.dinb(w_n427_2[1]),.dout(n827),.clk(gclk));
	jand g0779(.dina(w_n827_0[2]),.dinb(w_n825_1[2]),.dout(n828),.clk(gclk));
	jand g0780(.dina(w_n561_1[0]),.dinb(w_n351_0[2]),.dout(n829),.clk(gclk));
	jnot g0781(.din(w_n744_0[0]),.dout(n830),.clk(gclk));
	jand g0782(.dina(n830),.dinb(n829),.dout(n831),.clk(gclk));
	jand g0783(.dina(n831),.dinb(n828),.dout(n832),.clk(gclk));
	jand g0784(.dina(n832),.dinb(w_n824_0[1]),.dout(n833),.clk(gclk));
	jand g0785(.dina(n833),.dinb(w_n723_0[0]),.dout(n834),.clk(gclk));
	jand g0786(.dina(w_n389_3[1]),.dinb(w_n191_2[2]),.dout(n835),.clk(gclk));
	jand g0787(.dina(w_n835_0[1]),.dinb(w_n294_2[2]),.dout(n836),.clk(gclk));
	jand g0788(.dina(n836),.dinb(w_n539_1[1]),.dout(n837),.clk(gclk));
	jand g0789(.dina(n837),.dinb(w_n265_2[0]),.dout(n838),.clk(gclk));
	jand g0790(.dina(w_n276_3[0]),.dinb(w_n142_2[0]),.dout(n839),.clk(gclk));
	jand g0791(.dina(n839),.dinb(w_n572_0[0]),.dout(n840),.clk(gclk));
	jand g0792(.dina(w_n221_3[1]),.dinb(w_n162_1[2]),.dout(n841),.clk(gclk));
	jand g0793(.dina(w_n841_0[1]),.dinb(w_n435_2[1]),.dout(n842),.clk(gclk));
	jand g0794(.dina(w_n842_0[1]),.dinb(w_n506_2[0]),.dout(n843),.clk(gclk));
	jand g0795(.dina(n843),.dinb(n840),.dout(n844),.clk(gclk));
	jand g0796(.dina(n844),.dinb(n838),.dout(n845),.clk(gclk));
	jand g0797(.dina(w_n403_0[1]),.dinb(w_n114_2[2]),.dout(n846),.clk(gclk));
	jand g0798(.dina(n846),.dinb(w_n245_1[1]),.dout(n847),.clk(gclk));
	jand g0799(.dina(w_n847_0[1]),.dinb(w_n457_0[1]),.dout(n848),.clk(gclk));
	jand g0800(.dina(n848),.dinb(w_n213_2[2]),.dout(n849),.clk(gclk));
	jand g0801(.dina(w_n321_2[1]),.dinb(w_n286_2[2]),.dout(n850),.clk(gclk));
	jand g0802(.dina(w_n850_0[2]),.dinb(w_n370_2[2]),.dout(n851),.clk(gclk));
	jor g0803(.dina(w_n336_0[2]),.dinb(w_n113_0[2]),.dout(n852),.clk(gclk));
	jand g0804(.dina(w_n852_1[1]),.dinb(w_n218_2[2]),.dout(n853),.clk(gclk));
	jand g0805(.dina(w_n461_0[1]),.dinb(w_n236_0[2]),.dout(n854),.clk(gclk));
	jand g0806(.dina(n854),.dinb(w_n853_0[2]),.dout(n855),.clk(gclk));
	jand g0807(.dina(n855),.dinb(n851),.dout(n856),.clk(gclk));
	jand g0808(.dina(w_n856_0[1]),.dinb(w_n849_0[2]),.dout(n857),.clk(gclk));
	jand g0809(.dina(n857),.dinb(n845),.dout(n858),.clk(gclk));
	jnot g0810(.din(w_n786_0[0]),.dout(n859),.clk(gclk));
	jand g0811(.dina(w_n456_0[1]),.dinb(w_n170_2[2]),.dout(n860),.clk(gclk));
	jand g0812(.dina(n860),.dinb(n859),.dout(n861),.clk(gclk));
	jand g0813(.dina(w_n374_2[2]),.dinb(w_n353_2[0]),.dout(n862),.clk(gclk));
	jand g0814(.dina(w_n510_3[0]),.dinb(w_n489_3[0]),.dout(n863),.clk(gclk));
	jand g0815(.dina(w_n366_2[2]),.dinb(w_n346_2[0]),.dout(n864),.clk(gclk));
	jand g0816(.dina(n864),.dinb(w_n863_0[1]),.dout(n865),.clk(gclk));
	jand g0817(.dina(n865),.dinb(w_n862_0[1]),.dout(n866),.clk(gclk));
	jnot g0818(.din(w_n803_0[0]),.dout(n867),.clk(gclk));
	jand g0819(.dina(n867),.dinb(w_n866_0[1]),.dout(n868),.clk(gclk));
	jand g0820(.dina(w_n377_3[1]),.dinb(w_n204_2[0]),.dout(n869),.clk(gclk));
	jand g0821(.dina(w_n188_1[2]),.dinb(w_n158_1[0]),.dout(n870),.clk(gclk));
	jand g0822(.dina(n870),.dinb(n869),.dout(n871),.clk(gclk));
	jand g0823(.dina(w_n871_0[1]),.dinb(w_n147_1[2]),.dout(n872),.clk(gclk));
	jand g0824(.dina(n872),.dinb(n868),.dout(n873),.clk(gclk));
	jand g0825(.dina(n873),.dinb(n861),.dout(n874),.clk(gclk));
	jand g0826(.dina(n874),.dinb(w_n858_0[1]),.dout(n875),.clk(gclk));
	jand g0827(.dina(n875),.dinb(w_n834_0[1]),.dout(n876),.clk(gclk));
	jxor g0828(.dina(w_n876_1[1]),.dinb(w_n716_8[1]),.dout(n877),.clk(gclk));
	jand g0829(.dina(w_n877_0[2]),.dinb(w_n815_1[1]),.dout(n878),.clk(gclk));
	jand g0830(.dina(w_n57_0[0]),.dinb(w_n49_7[0]),.dout(n879),.clk(gclk));
	jxor g0831(.dina(n879),.dinb(w_a9_0[0]),.dout(n880),.clk(gclk));
	jnot g0832(.din(w_n880_6[1]),.dout(n881),.clk(gclk));
	jand g0833(.dina(w_n881_4[2]),.dinb(w_n878_1[2]),.dout(n882),.clk(gclk));
	jand g0834(.dina(w_n370_2[1]),.dinb(w_n221_3[0]),.dout(n883),.clk(gclk));
	jand g0835(.dina(w_n377_3[0]),.dinb(w_n233_1[2]),.dout(n884),.clk(gclk));
	jand g0836(.dina(w_n884_1[1]),.dinb(n883),.dout(n885),.clk(gclk));
	jand g0837(.dina(n885),.dinb(w_n361_2[1]),.dout(n886),.clk(gclk));
	jand g0838(.dina(w_n267_2[1]),.dinb(w_n129_1[1]),.dout(n887),.clk(gclk));
	jand g0839(.dina(n887),.dinb(w_n294_2[1]),.dout(n888),.clk(gclk));
	jand g0840(.dina(n888),.dinb(w_n886_1[1]),.dout(n889),.clk(gclk));
	jand g0841(.dina(w_n387_3[0]),.dinb(w_n222_3[0]),.dout(n890),.clk(gclk));
	jand g0842(.dina(n890),.dinb(w_n600_2[1]),.dout(n891),.clk(gclk));
	jand g0843(.dina(n891),.dinb(w_n448_2[0]),.dout(n892),.clk(gclk));
	jand g0844(.dina(w_n587_3[0]),.dinb(w_n335_0[1]),.dout(n893),.clk(gclk));
	jand g0845(.dina(n893),.dinb(n892),.dout(n894),.clk(gclk));
	jand g0846(.dina(n894),.dinb(n889),.dout(n895),.clk(gclk));
	jand g0847(.dina(n895),.dinb(w_n417_0[0]),.dout(n896),.clk(gclk));
	jor g0848(.dina(w_n151_0[2]),.dinb(w_n108_1[1]),.dout(n897),.clk(gclk));
	jand g0849(.dina(w_n897_2[1]),.dinb(w_n366_2[1]),.dout(n898),.clk(gclk));
	jand g0850(.dina(n898),.dinb(w_n463_0[1]),.dout(n899),.clk(gclk));
	jand g0851(.dina(w_n481_0[2]),.dinb(w_n290_3[0]),.dout(n900),.clk(gclk));
	jand g0852(.dina(n900),.dinb(w_n825_1[1]),.dout(n901),.clk(gclk));
	jand g0853(.dina(n901),.dinb(w_n557_0[0]),.dout(n902),.clk(gclk));
	jand g0854(.dina(n902),.dinb(n899),.dout(n903),.clk(gclk));
	jand g0855(.dina(w_n418_1[1]),.dinb(w_n261_2[1]),.dout(n904),.clk(gclk));
	jand g0856(.dina(w_n904_1[1]),.dinb(w_n546_0[1]),.dout(n905),.clk(gclk));
	jand g0857(.dina(w_n344_2[2]),.dinb(w_n281_0[1]),.dout(n906),.clk(gclk));
	jand g0858(.dina(n906),.dinb(n905),.dout(n907),.clk(gclk));
	jand g0859(.dina(w_n445_2[0]),.dinb(w_n152_2[0]),.dout(n908),.clk(gclk));
	jand g0860(.dina(w_n378_2[1]),.dinb(w_n305_1[2]),.dout(n909),.clk(gclk));
	jand g0861(.dina(n909),.dinb(w_n339_3[2]),.dout(n910),.clk(gclk));
	jand g0862(.dina(n910),.dinb(n908),.dout(n911),.clk(gclk));
	jand g0863(.dina(n911),.dinb(n907),.dout(n912),.clk(gclk));
	jand g0864(.dina(w_n912_0[2]),.dinb(w_n903_0[1]),.dout(n913),.clk(gclk));
	jand g0865(.dina(n913),.dinb(w_n849_0[1]),.dout(n914),.clk(gclk));
	jand g0866(.dina(w_n569_2[0]),.dinb(w_n535_2[0]),.dout(n915),.clk(gclk));
	jand g0867(.dina(w_n915_0[2]),.dinb(w_n527_3[0]),.dout(n916),.clk(gclk));
	jand g0868(.dina(w_n562_1[0]),.dinb(w_n315_2[0]),.dout(n917),.clk(gclk));
	jand g0869(.dina(n917),.dinb(n916),.dout(n918),.clk(gclk));
	jnot g0870(.din(w_n697_0[0]),.dout(n919),.clk(gclk));
	jand g0871(.dina(w_n919_0[1]),.dinb(w_n439_4[0]),.dout(n920),.clk(gclk));
	jand g0872(.dina(n920),.dinb(w_n338_0[1]),.dout(n921),.clk(gclk));
	jand g0873(.dina(w_n853_0[1]),.dinb(w_n921_0[1]),.dout(n922),.clk(gclk));
	jand g0874(.dina(n922),.dinb(n918),.dout(n923),.clk(gclk));
	jand g0875(.dina(w_n717_3[0]),.dinb(w_n169_2[0]),.dout(n924),.clk(gclk));
	jand g0876(.dina(w_n924_0[2]),.dinb(w_n187_1[2]),.dout(n925),.clk(gclk));
	jand g0877(.dina(n925),.dinb(w_n160_1[2]),.dout(n926),.clk(gclk));
	jand g0878(.dina(n926),.dinb(w_n310_1[2]),.dout(n927),.clk(gclk));
	jand g0879(.dina(n927),.dinb(n923),.dout(n928),.clk(gclk));
	jand g0880(.dina(n928),.dinb(n914),.dout(n929),.clk(gclk));
	jand g0881(.dina(n929),.dinb(w_n896_0[2]),.dout(n930),.clk(gclk));
	jand g0882(.dina(w_n876_1[0]),.dinb(w_n930_2[1]),.dout(n931),.clk(gclk));
	jnot g0883(.din(w_n522_0[0]),.dout(n932),.clk(gclk));
	jnot g0884(.din(w_n528_0[0]),.dout(n933),.clk(gclk));
	jor g0885(.dina(n933),.dinb(w_n524_0[0]),.dout(n934),.clk(gclk));
	jor g0886(.dina(n934),.dinb(n932),.dout(n935),.clk(gclk));
	jnot g0887(.din(w_n532_0[0]),.dout(n936),.clk(gclk));
	jor g0888(.dina(n936),.dinb(n935),.dout(n937),.clk(gclk));
	jand g0889(.dina(w_n167_1[0]),.dinb(w_n224_2[0]),.dout(n938),.clk(gclk));
	jor g0890(.dina(w_n752_0[1]),.dinb(n938),.dout(n939),.clk(gclk));
	jor g0891(.dina(n939),.dinb(w_n685_0[0]),.dout(n940),.clk(gclk));
	jor g0892(.dina(n940),.dinb(w_n727_0[0]),.dout(n941),.clk(gclk));
	jand g0893(.dina(w_n192_1[1]),.dinb(w_n253_2[2]),.dout(n942),.clk(gclk));
	jor g0894(.dina(w_n766_0[0]),.dinb(n942),.dout(n943),.clk(gclk));
	jor g0895(.dina(n943),.dinb(w_n751_0[0]),.dout(n944),.clk(gclk));
	jor g0896(.dina(n944),.dinb(w_n266_0[2]),.dout(n945),.clk(gclk));
	jor g0897(.dina(n945),.dinb(n941),.dout(n946),.clk(gclk));
	jand g0898(.dina(w_n295_0[0]),.dinb(w_n100_2[2]),.dout(n947),.clk(gclk));
	jor g0899(.dina(n947),.dinb(w_n612_0[0]),.dout(n948),.clk(gclk));
	jor g0900(.dina(n948),.dinb(w_n282_1[0]),.dout(n949),.clk(gclk));
	jor g0901(.dina(n949),.dinb(w_n401_0[1]),.dout(n950),.clk(gclk));
	jor g0902(.dina(w_n661_0[0]),.dinb(w_n132_0[0]),.dout(n951),.clk(gclk));
	jor g0903(.dina(n951),.dinb(w_n544_0[0]),.dout(n952),.clk(gclk));
	jor g0904(.dina(n952),.dinb(n950),.dout(n953),.clk(gclk));
	jor g0905(.dina(n953),.dinb(n946),.dout(n954),.clk(gclk));
	jor g0906(.dina(n954),.dinb(n937),.dout(n955),.clk(gclk));
	jnot g0907(.din(w_n552_0[1]),.dout(n956),.clk(gclk));
	jnot g0908(.din(w_n559_0[0]),.dout(n957),.clk(gclk));
	jor g0909(.dina(n957),.dinb(w_n555_0[0]),.dout(n958),.clk(gclk));
	jnot g0910(.din(w_n563_0[0]),.dout(n959),.clk(gclk));
	jor g0911(.dina(n959),.dinb(n958),.dout(n960),.clk(gclk));
	jor g0912(.dina(n960),.dinb(n956),.dout(n961),.clk(gclk));
	jor g0913(.dina(n961),.dinb(n955),.dout(n962),.clk(gclk));
	jnot g0914(.din(w_n574_0[0]),.dout(n963),.clk(gclk));
	jor g0915(.dina(w_n655_0[0]),.dinb(w_n646_0[0]),.dout(n964),.clk(gclk));
	jand g0916(.dina(w_n155_1[2]),.dinb(w_n118_2[0]),.dout(n965),.clk(gclk));
	jand g0917(.dina(w_n253_2[1]),.dinb(w_n98_1[2]),.dout(n966),.clk(gclk));
	jor g0918(.dina(w_n966_0[1]),.dinb(w_n965_0[1]),.dout(n967),.clk(gclk));
	jor g0919(.dina(n967),.dinb(n964),.dout(n968),.clk(gclk));
	jand g0920(.dina(w_n155_1[1]),.dinb(w_n144_2[2]),.dout(n969),.clk(gclk));
	jor g0921(.dina(w_n634_0[1]),.dinb(n969),.dout(n970),.clk(gclk));
	jor g0922(.dina(w_n802_0[0]),.dinb(w_n619_0[0]),.dout(n971),.clk(gclk));
	jor g0923(.dina(n971),.dinb(n970),.dout(n972),.clk(gclk));
	jor g0924(.dina(n972),.dinb(w_n968_0[1]),.dout(n973),.clk(gclk));
	jand g0925(.dina(w_n230_1[0]),.dinb(w_n184_2[0]),.dout(n974),.clk(gclk));
	jand g0926(.dina(w_n174_2[0]),.dinb(w_n98_1[1]),.dout(n975),.clk(gclk));
	jor g0927(.dina(w_n975_0[1]),.dinb(w_n974_0[1]),.dout(n976),.clk(gclk));
	jor g0928(.dina(n976),.dinb(w_n247_0[0]),.dout(n977),.clk(gclk));
	jand g0929(.dina(w_n155_1[0]),.dinb(w_n253_2[0]),.dout(n978),.clk(gclk));
	jor g0930(.dina(n978),.dinb(w_n654_0[1]),.dout(n979),.clk(gclk));
	jor g0931(.dina(n979),.dinb(w_n677_0[2]),.dout(n980),.clk(gclk));
	jor g0932(.dina(n980),.dinb(n977),.dout(n981),.clk(gclk));
	jor g0933(.dina(n981),.dinb(n973),.dout(n982),.clk(gclk));
	jor g0934(.dina(n982),.dinb(w_n582_0[0]),.dout(n983),.clk(gclk));
	jnot g0935(.din(w_n604_0[0]),.dout(n984),.clk(gclk));
	jor g0936(.dina(n984),.dinb(n983),.dout(n985),.clk(gclk));
	jor g0937(.dina(n985),.dinb(n963),.dout(n986),.clk(gclk));
	jor g0938(.dina(n986),.dinb(n962),.dout(n987),.clk(gclk));
	jand g0939(.dina(w_n814_0[0]),.dinb(w_n987_1[1]),.dout(n988),.clk(gclk));
	jor g0940(.dina(n988),.dinb(w_n931_0[1]),.dout(n989),.clk(gclk));
	jand g0941(.dina(w_n989_2[1]),.dinb(w_n880_6[0]),.dout(n990),.clk(gclk));
	jor g0942(.dina(n990),.dinb(n882),.dout(n991),.clk(gclk));
	jor g0943(.dina(w_n931_0[0]),.dinb(w_n815_1[0]),.dout(n992),.clk(gclk));
	jand g0944(.dina(w_n58_0[0]),.dinb(w_n49_6[2]),.dout(n993),.clk(gclk));
	jxor g0945(.dina(n993),.dinb(w_a10_0[0]),.dout(n994),.clk(gclk));
	jand g0946(.dina(w_n994_6[1]),.dinb(w_n992_3[2]),.dout(n995),.clk(gclk));
	jnot g0947(.din(w_n994_6[0]),.dout(n996),.clk(gclk));
	jor g0948(.dina(w_n877_0[1]),.dinb(w_n987_1[0]),.dout(n997),.clk(gclk));
	jand g0949(.dina(w_n997_4[1]),.dinb(w_n996_4[2]),.dout(n998),.clk(gclk));
	jor g0950(.dina(n998),.dinb(n995),.dout(n999),.clk(gclk));
	jnot g0951(.din(n999),.dout(n1000),.clk(gclk));
	jor g0952(.dina(n1000),.dinb(n991),.dout(n1001),.clk(gclk));
	jand g0953(.dina(w_n250_1[2]),.dinb(w_n120_1[2]),.dout(n1002),.clk(gclk));
	jand g0954(.dina(w_n488_3[0]),.dinb(w_n409_1[2]),.dout(n1003),.clk(gclk));
	jand g0955(.dina(w_n192_1[0]),.dinb(w_n144_2[1]),.dout(n1004),.clk(gclk));
	jnot g0956(.din(n1004),.dout(n1005),.clk(gclk));
	jand g0957(.dina(w_n1005_4[1]),.dinb(w_n570_2[0]),.dout(n1006),.clk(gclk));
	jand g0958(.dina(w_n333_1[1]),.dinb(w_n245_1[0]),.dout(n1007),.clk(gclk));
	jand g0959(.dina(n1007),.dinb(w_n1006_0[1]),.dout(n1008),.clk(gclk));
	jand g0960(.dina(n1008),.dinb(n1003),.dout(n1009),.clk(gclk));
	jand g0961(.dina(w_n1009_0[1]),.dinb(w_n352_0[2]),.dout(n1010),.clk(gclk));
	jand g0962(.dina(n1010),.dinb(w_n1002_0[1]),.dout(n1011),.clk(gclk));
	jand g0963(.dina(w_n344_2[1]),.dinb(w_n187_1[1]),.dout(n1012),.clk(gclk));
	jand g0964(.dina(w_n1012_0[1]),.dinb(w_n897_2[0]),.dout(n1013),.clk(gclk));
	jand g0965(.dina(n1013),.dinb(w_n398_0[1]),.dout(n1014),.clk(gclk));
	jand g0966(.dina(n1014),.dinb(w_n166_2[0]),.dout(n1015),.clk(gclk));
	jand g0967(.dina(n1015),.dinb(n1011),.dout(n1016),.clk(gclk));
	jnot g0968(.din(w_n785_0[0]),.dout(n1017),.clk(gclk));
	jand g0969(.dina(w_n332_2[1]),.dinb(w_n128_2[1]),.dout(n1018),.clk(gclk));
	jand g0970(.dina(w_n404_1[1]),.dinb(w_n252_3[2]),.dout(n1019),.clk(gclk));
	jand g0971(.dina(w_n1019_0[1]),.dinb(w_n841_0[0]),.dout(n1020),.clk(gclk));
	jand g0972(.dina(n1020),.dinb(n1018),.dout(n1021),.clk(gclk));
	jand g0973(.dina(w_n1021_0[1]),.dinb(w_n1017_0[1]),.dout(n1022),.clk(gclk));
	jand g0974(.dina(w_n278_1[0]),.dinb(w_n261_2[0]),.dout(n1023),.clk(gclk));
	jand g0975(.dina(w_n1023_0[1]),.dinb(w_n240_1[2]),.dout(n1024),.clk(gclk));
	jand g0976(.dina(w_n195_1[1]),.dinb(w_n158_0[2]),.dout(n1025),.clk(gclk));
	jor g0977(.dina(w_n965_0[0]),.dinb(w_n314_0[0]),.dout(n1026),.clk(gclk));
	jnot g0978(.din(w_n1026_0[1]),.dout(n1027),.clk(gclk));
	jand g0979(.dina(n1027),.dinb(w_n1025_0[2]),.dout(n1028),.clk(gclk));
	jand g0980(.dina(n1028),.dinb(w_n1024_0[2]),.dout(n1029),.clk(gclk));
	jand g0981(.dina(w_n527_2[2]),.dinb(w_n340_1[1]),.dout(n1030),.clk(gclk));
	jand g0982(.dina(w_n1030_0[1]),.dinb(n1029),.dout(n1031),.clk(gclk));
	jand g0983(.dina(n1031),.dinb(w_n1022_0[1]),.dout(n1032),.clk(gclk));
	jand g0984(.dina(w_n275_1[2]),.dinb(w_n152_1[2]),.dout(n1033),.clk(gclk));
	jand g0985(.dina(w_n301_0[1]),.dinb(w_n77_3[0]),.dout(n1034),.clk(gclk));
	jnot g0986(.din(n1034),.dout(n1035),.clk(gclk));
	jand g0987(.dina(w_n1035_2[2]),.dinb(w_n384_2[2]),.dout(n1036),.clk(gclk));
	jand g0988(.dina(w_n506_1[2]),.dinb(w_n438_1[2]),.dout(n1037),.clk(gclk));
	jand g0989(.dina(n1037),.dinb(n1036),.dout(n1038),.clk(gclk));
	jand g0990(.dina(n1038),.dinb(w_n1033_0[1]),.dout(n1039),.clk(gclk));
	jor g0991(.dina(w_n796_0[0]),.dinb(w_n426_0[0]),.dout(n1040),.clk(gclk));
	jnot g0992(.din(w_n1040_0[1]),.dout(n1041),.clk(gclk));
	jand g0993(.dina(n1041),.dinb(w_n234_0[1]),.dout(n1042),.clk(gclk));
	jand g0994(.dina(w_n347_2[0]),.dinb(w_n310_1[1]),.dout(n1043),.clk(gclk));
	jand g0995(.dina(w_n1043_0[1]),.dinb(w_n402_0[0]),.dout(n1044),.clk(gclk));
	jand g0996(.dina(n1044),.dinb(n1042),.dout(n1045),.clk(gclk));
	jand g0997(.dina(w_n1045_0[1]),.dinb(w_n159_0[2]),.dout(n1046),.clk(gclk));
	jand g0998(.dina(n1046),.dinb(w_n1039_0[2]),.dout(n1047),.clk(gclk));
	jand g0999(.dina(n1047),.dinb(w_n1032_0[1]),.dout(n1048),.clk(gclk));
	jand g1000(.dina(w_n569_1[2]),.dinb(w_n382_1[1]),.dout(n1049),.clk(gclk));
	jand g1001(.dina(n1049),.dinb(w_n269_1[1]),.dout(n1050),.clk(gclk));
	jand g1002(.dina(w_n1050_0[1]),.dinb(w_n377_2[2]),.dout(n1051),.clk(gclk));
	jand g1003(.dina(w_n420_0[0]),.dinb(w_n248_3[0]),.dout(n1052),.clk(gclk));
	jand g1004(.dina(n1052),.dinb(n1051),.dout(n1053),.clk(gclk));
	jand g1005(.dina(w_n1053_0[1]),.dinb(n1048),.dout(n1054),.clk(gclk));
	jand g1006(.dina(n1054),.dinb(w_n1016_1[1]),.dout(n1055),.clk(gclk));
	jand g1007(.dina(w_n915_0[1]),.dinb(w_n133_1[1]),.dout(n1056),.clk(gclk));
	jand g1008(.dina(w_n429_1[1]),.dinb(w_n332_2[0]),.dout(n1057),.clk(gclk));
	jand g1009(.dina(w_n1057_0[1]),.dinb(w_n215_3[0]),.dout(n1058),.clk(gclk));
	jand g1010(.dina(n1058),.dinb(w_n437_1[1]),.dout(n1059),.clk(gclk));
	jand g1011(.dina(n1059),.dinb(w_n1056_0[1]),.dout(n1060),.clk(gclk));
	jand g1012(.dina(w_n835_0[0]),.dinb(w_n489_2[2]),.dout(n1061),.clk(gclk));
	jand g1013(.dina(w_n497_1[0]),.dinb(w_n238_1[2]),.dout(n1062),.clk(gclk));
	jand g1014(.dina(n1062),.dinb(n1061),.dout(n1063),.clk(gclk));
	jand g1015(.dina(w_n300_2[2]),.dinb(w_n136_1[2]),.dout(n1064),.clk(gclk));
	jand g1016(.dina(w_n1064_1[1]),.dinb(w_n148_1[0]),.dout(n1065),.clk(gclk));
	jand g1017(.dina(w_n377_2[1]),.dinb(w_n315_1[2]),.dout(n1066),.clk(gclk));
	jand g1018(.dina(w_n1066_0[1]),.dinb(n1065),.dout(n1067),.clk(gclk));
	jand g1019(.dina(n1067),.dinb(n1063),.dout(n1068),.clk(gclk));
	jand g1020(.dina(n1068),.dinb(w_n1060_0[1]),.dout(n1069),.clk(gclk));
	jand g1021(.dina(w_n1069_0[1]),.dinb(w_n570_1[2]),.dout(n1070),.clk(gclk));
	jand g1022(.dina(n1070),.dinb(w_n370_2[0]),.dout(n1071),.clk(gclk));
	jand g1023(.dina(w_n378_2[0]),.dinb(w_n226_2[0]),.dout(n1072),.clk(gclk));
	jnot g1024(.din(w_n577_0[0]),.dout(n1073),.clk(gclk));
	jand g1025(.dina(w_n1073_1[1]),.dinb(w_n460_3[0]),.dout(n1074),.clk(gclk));
	jand g1026(.dina(w_n1074_1[2]),.dinb(w_n197_2[1]),.dout(n1075),.clk(gclk));
	jand g1027(.dina(w_n427_2[0]),.dinb(w_n129_1[0]),.dout(n1076),.clk(gclk));
	jand g1028(.dina(n1076),.dinb(n1075),.dout(n1077),.clk(gclk));
	jand g1029(.dina(n1077),.dinb(w_n904_1[0]),.dout(n1078),.clk(gclk));
	jand g1030(.dina(w_n1078_0[1]),.dinb(w_n1012_0[0]),.dout(n1079),.clk(gclk));
	jand g1031(.dina(w_n445_1[2]),.dinb(w_n395_1[2]),.dout(n1080),.clk(gclk));
	jand g1032(.dina(w_n1080_0[1]),.dinb(w_n850_0[1]),.dout(n1081),.clk(gclk));
	jand g1033(.dina(n1081),.dinb(w_n1079_0[1]),.dout(n1082),.clk(gclk));
	jand g1034(.dina(n1082),.dinb(w_n1072_1[1]),.dout(n1083),.clk(gclk));
	jand g1035(.dina(n1083),.dinb(w_n1071_0[1]),.dout(n1084),.clk(gclk));
	jand g1036(.dina(w_n310_1[0]),.dinb(w_n222_2[2]),.dout(n1085),.clk(gclk));
	jand g1037(.dina(w_n1085_0[1]),.dinb(w_n435_2[0]),.dout(n1086),.clk(gclk));
	jand g1038(.dina(n1086),.dinb(w_n248_2[2]),.dout(n1087),.clk(gclk));
	jand g1039(.dina(w_n294_2[0]),.dinb(w_n114_2[1]),.dout(n1088),.clk(gclk));
	jand g1040(.dina(w_n1088_0[1]),.dinb(w_n366_2[0]),.dout(n1089),.clk(gclk));
	jand g1041(.dina(n1089),.dinb(w_n1087_0[2]),.dout(n1090),.clk(gclk));
	jand g1042(.dina(w_n467_2[0]),.dinb(w_n218_2[1]),.dout(n1091),.clk(gclk));
	jand g1043(.dina(w_n313_1[1]),.dinb(w_n276_2[2]),.dout(n1092),.clk(gclk));
	jand g1044(.dina(n1092),.dinb(n1091),.dout(n1093),.clk(gclk));
	jand g1045(.dina(w_n185_1[0]),.dinb(w_n144_2[0]),.dout(n1094),.clk(gclk));
	jnot g1046(.din(w_n1094_0[1]),.dout(n1095),.clk(gclk));
	jand g1047(.dina(w_n462_1[2]),.dinb(w_n206_1[2]),.dout(n1096),.clk(gclk));
	jand g1048(.dina(w_n1096_0[2]),.dinb(w_n1095_2[2]),.dout(n1097),.clk(gclk));
	jand g1049(.dina(w_n232_4[0]),.dinb(w_n160_1[1]),.dout(n1098),.clk(gclk));
	jand g1050(.dina(n1098),.dinb(w_n1097_0[1]),.dout(n1099),.clk(gclk));
	jand g1051(.dina(n1099),.dinb(w_n1093_0[1]),.dout(n1100),.clk(gclk));
	jand g1052(.dina(w_n290_2[2]),.dinb(w_n204_1[2]),.dout(n1101),.clk(gclk));
	jand g1053(.dina(n1101),.dinb(w_n446_2[0]),.dout(n1102),.clk(gclk));
	jand g1054(.dina(w_n280_2[0]),.dinb(w_n157_3[0]),.dout(n1103),.clk(gclk));
	jand g1055(.dina(n1103),.dinb(w_n267_2[0]),.dout(n1104),.clk(gclk));
	jand g1056(.dina(w_n506_1[1]),.dinb(w_n404_1[0]),.dout(n1105),.clk(gclk));
	jand g1057(.dina(w_n1105_0[2]),.dinb(w_n362_0[0]),.dout(n1106),.clk(gclk));
	jand g1058(.dina(n1106),.dinb(w_n1104_0[1]),.dout(n1107),.clk(gclk));
	jand g1059(.dina(n1107),.dinb(w_n1102_0[1]),.dout(n1108),.clk(gclk));
	jand g1060(.dina(n1108),.dinb(n1100),.dout(n1109),.clk(gclk));
	jand g1061(.dina(w_n717_2[2]),.dinb(w_n173_1[1]),.dout(n1110),.clk(gclk));
	jand g1062(.dina(w_n1110_0[2]),.dinb(w_n288_1[2]),.dout(n1111),.clk(gclk));
	jand g1063(.dina(n1111),.dinb(w_n1109_0[1]),.dout(n1112),.clk(gclk));
	jand g1064(.dina(n1112),.dinb(n1090),.dout(n1113),.clk(gclk));
	jand g1065(.dina(n1113),.dinb(n1084),.dout(n1114),.clk(gclk));
	jxor g1066(.dina(w_n1114_0[2]),.dinb(w_n1055_2[1]),.dout(n1115),.clk(gclk));
	jor g1067(.dina(w_n1114_0[1]),.dinb(w_n1055_2[0]),.dout(n1116),.clk(gclk));
	jand g1068(.dina(w_n1005_4[0]),.dinb(w_n374_2[1]),.dout(n1117),.clk(gclk));
	jand g1069(.dina(w_n446_1[2]),.dinb(w_n267_1[2]),.dout(n1118),.clk(gclk));
	jand g1070(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jand g1071(.dina(n1119),.dinb(w_n603_0[0]),.dout(n1120),.clk(gclk));
	jand g1072(.dina(w_n467_1[2]),.dinb(w_n339_3[1]),.dout(n1121),.clk(gclk));
	jand g1073(.dina(n1121),.dinb(w_n346_1[2]),.dout(n1122),.clk(gclk));
	jand g1074(.dina(w_n1088_0[0]),.dinb(w_n492_0[0]),.dout(n1123),.clk(gclk));
	jand g1075(.dina(n1123),.dinb(w_n448_1[2]),.dout(n1124),.clk(gclk));
	jand g1076(.dina(w_n1124_0[1]),.dinb(w_n1122_0[1]),.dout(n1125),.clk(gclk));
	jand g1077(.dina(n1125),.dinb(w_n1120_0[1]),.dout(n1126),.clk(gclk));
	jand g1078(.dina(w_n1073_1[0]),.dinb(w_n313_1[0]),.dout(n1127),.clk(gclk));
	jand g1079(.dina(w_n415_2[0]),.dinb(w_n327_1[0]),.dout(n1128),.clk(gclk));
	jand g1080(.dina(w_n429_1[0]),.dinb(w_n252_3[1]),.dout(n1129),.clk(gclk));
	jand g1081(.dina(n1129),.dinb(n1128),.dout(n1130),.clk(gclk));
	jand g1082(.dina(w_n1130_0[1]),.dinb(w_n527_2[1]),.dout(n1131),.clk(gclk));
	jand g1083(.dina(w_n570_1[1]),.dinb(w_n297_1[0]),.dout(n1132),.clk(gclk));
	jand g1084(.dina(n1132),.dinb(w_n222_2[1]),.dout(n1133),.clk(gclk));
	jand g1085(.dina(w_n1133_0[1]),.dinb(w_n255_1[2]),.dout(n1134),.clk(gclk));
	jand g1086(.dina(n1134),.dinb(w_n238_1[1]),.dout(n1135),.clk(gclk));
	jand g1087(.dina(w_n1135_1[1]),.dinb(n1131),.dout(n1136),.clk(gclk));
	jand g1088(.dina(n1136),.dinb(w_n1127_0[2]),.dout(n1137),.clk(gclk));
	jand g1089(.dina(n1137),.dinb(n1126),.dout(n1138),.clk(gclk));
	jand g1090(.dina(w_n510_2[2]),.dinb(w_n221_2[2]),.dout(n1139),.clk(gclk));
	jand g1091(.dina(n1139),.dinb(w_n180_1[0]),.dout(n1140),.clk(gclk));
	jand g1092(.dina(w_n720_0[0]),.dinb(w_n332_1[2]),.dout(n1141),.clk(gclk));
	jand g1093(.dina(n1141),.dinb(w_n593_0[0]),.dout(n1142),.clk(gclk));
	jand g1094(.dina(n1142),.dinb(w_n372_0[0]),.dout(n1143),.clk(gclk));
	jand g1095(.dina(n1143),.dinb(w_n600_2[0]),.dout(n1144),.clk(gclk));
	jand g1096(.dina(w_n921_0[0]),.dinb(w_n191_2[1]),.dout(n1145),.clk(gclk));
	jand g1097(.dina(n1145),.dinb(w_n293_0[0]),.dout(n1146),.clk(gclk));
	jand g1098(.dina(n1146),.dinb(n1144),.dout(n1147),.clk(gclk));
	jand g1099(.dina(w_n1147_0[1]),.dinb(w_n1140_0[1]),.dout(n1148),.clk(gclk));
	jand g1100(.dina(n1148),.dinb(n1138),.dout(n1149),.clk(gclk));
	jnot g1101(.din(w_n1149_1[2]),.dout(n1150),.clk(gclk));
	jand g1102(.dina(w_n1150_0[1]),.dinb(n1116),.dout(n1151),.clk(gclk));
	jor g1103(.dina(w_n1151_1[2]),.dinb(w_n1115_1[1]),.dout(n1152),.clk(gclk));
	jand g1104(.dina(w_n53_0[0]),.dinb(w_n49_6[1]),.dout(n1153),.clk(gclk));
	jxor g1105(.dina(n1153),.dinb(w_a5_0[0]),.dout(n1154),.clk(gclk));
	jor g1106(.dina(w_n1154_10[2]),.dinb(w_n1152_2[1]),.dout(n1155),.clk(gclk));
	jnot g1107(.din(w_n1154_10[1]),.dout(n1156),.clk(gclk));
	jand g1108(.dina(w_n1114_0[0]),.dinb(w_n1055_1[2]),.dout(n1157),.clk(gclk));
	jnot g1109(.din(n1157),.dout(n1158),.clk(gclk));
	jand g1110(.dina(w_n1149_1[1]),.dinb(w_n1158_0[1]),.dout(n1159),.clk(gclk));
	jor g1111(.dina(n1159),.dinb(w_n1115_1[0]),.dout(n1160),.clk(gclk));
	jor g1112(.dina(w_n1160_2[1]),.dinb(w_n1156_12[1]),.dout(n1161),.clk(gclk));
	jand g1113(.dina(n1161),.dinb(n1155),.dout(n1162),.clk(gclk));
	jand g1114(.dina(w_n1151_1[1]),.dinb(w_n1158_0[0]),.dout(n1163),.clk(gclk));
	jnot g1115(.din(w_n1163_0[2]),.dout(n1164),.clk(gclk));
	jand g1116(.dina(w_n54_0[0]),.dinb(w_n49_6[0]),.dout(n1165),.clk(gclk));
	jxor g1117(.dina(n1165),.dinb(w_a6_0[0]),.dout(n1166),.clk(gclk));
	jand g1118(.dina(w_n1166_6[1]),.dinb(w_n1164_3[2]),.dout(n1167),.clk(gclk));
	jnot g1119(.din(w_n1166_6[0]),.dout(n1168),.clk(gclk));
	jnot g1120(.din(w_n1115_0[2]),.dout(n1169),.clk(gclk));
	jor g1121(.dina(w_n1150_0[0]),.dinb(n1169),.dout(n1170),.clk(gclk));
	jand g1122(.dina(w_n1170_4[1]),.dinb(w_n1168_4[2]),.dout(n1171),.clk(gclk));
	jor g1123(.dina(n1171),.dinb(n1167),.dout(n1172),.clk(gclk));
	jand g1124(.dina(n1172),.dinb(n1162),.dout(n1173),.clk(gclk));
	jnot g1125(.din(w_n1173_0[1]),.dout(n1174),.clk(gclk));
	jor g1126(.dina(n1174),.dinb(w_n1001_0[1]),.dout(n1175),.clk(gclk));
	jand g1127(.dina(w_n827_0[1]),.dinb(w_n506_1[0]),.dout(n1176),.clk(gclk));
	jnot g1128(.din(w_n1176_0[1]),.dout(n1177),.clk(gclk));
	jand g1129(.dina(w_n387_2[2]),.dinb(w_n173_1[0]),.dout(n1178),.clk(gclk));
	jnot g1130(.din(w_n1178_0[2]),.dout(n1179),.clk(gclk));
	jor g1131(.dina(w_n447_0[0]),.dinb(w_n975_0[0]),.dout(n1180),.clk(gclk));
	jor g1132(.dina(w_n1180_0[1]),.dinb(w_n634_0[0]),.dout(n1181),.clk(gclk));
	jor g1133(.dina(w_n1181_0[1]),.dinb(n1179),.dout(n1182),.clk(gclk));
	jor g1134(.dina(n1182),.dinb(n1177),.dout(n1183),.clk(gclk));
	jor g1135(.dina(n1183),.dinb(w_n787_0[0]),.dout(n1184),.clk(gclk));
	jor g1136(.dina(w_n660_0[0]),.dinb(w_n302_0[0]),.dout(n1185),.clk(gclk));
	jor g1137(.dina(w_n1185_0[1]),.dinb(w_n282_0[2]),.dout(n1186),.clk(gclk));
	jor g1138(.dina(w_n1186_0[1]),.dinb(w_n676_0[0]),.dout(n1187),.clk(gclk));
	jor g1139(.dina(n1187),.dinb(w_n274_0[0]),.dout(n1188),.clk(gclk));
	jor g1140(.dina(w_n1188_0[1]),.dinb(w_n677_0[1]),.dout(n1189),.clk(gclk));
	jor g1141(.dina(w_n1189_0[1]),.dinb(n1184),.dout(n1190),.clk(gclk));
	jand g1142(.dina(w_n374_2[0]),.dinb(w_n276_2[1]),.dout(n1191),.clk(gclk));
	jand g1143(.dina(n1191),.dinb(w_n1035_2[1]),.dout(n1192),.clk(gclk));
	jand g1144(.dina(w_n1192_0[1]),.dinb(w_n136_1[1]),.dout(n1193),.clk(gclk));
	jand g1145(.dina(w_n863_0[0]),.dinb(w_n244_2[1]),.dout(n1194),.clk(gclk));
	jand g1146(.dina(n1194),.dinb(w_n1019_0[0]),.dout(n1195),.clk(gclk));
	jand g1147(.dina(n1195),.dinb(n1193),.dout(n1196),.clk(gclk));
	jnot g1148(.din(w_n1196_1[1]),.dout(n1197),.clk(gclk));
	jnot g1149(.din(w_n1056_0[0]),.dout(n1198),.clk(gclk));
	jnot g1150(.din(w_n437_1[0]),.dout(n1199),.clk(gclk));
	jand g1151(.dina(w_n126_1[1]),.dinb(w_n262_2[0]),.dout(n1200),.clk(gclk));
	jor g1152(.dina(n1200),.dinb(w_n630_0[0]),.dout(n1201),.clk(gclk));
	jor g1153(.dina(n1201),.dinb(w_n214_0[0]),.dout(n1202),.clk(gclk));
	jor g1154(.dina(n1202),.dinb(n1199),.dout(n1203),.clk(gclk));
	jor g1155(.dina(n1203),.dinb(n1198),.dout(n1204),.clk(gclk));
	jand g1156(.dina(w_n439_3[2]),.dinb(w_n409_1[1]),.dout(n1205),.clk(gclk));
	jnot g1157(.din(w_n1205_0[1]),.dout(n1206),.clk(gclk));
	jor g1158(.dina(n1206),.dinb(n1204),.dout(n1207),.clk(gclk));
	jor g1159(.dina(n1207),.dinb(n1197),.dout(n1208),.clk(gclk));
	jor g1160(.dina(w_n617_0[0]),.dinb(w_n752_0[0]),.dout(n1209),.clk(gclk));
	jor g1161(.dina(w_n788_0[0]),.dinb(w_n667_0[0]),.dout(n1210),.clk(gclk));
	jor g1162(.dina(n1210),.dinb(n1209),.dout(n1211),.clk(gclk));
	jor g1163(.dina(w_n705_0[0]),.dinb(w_n625_0[0]),.dout(n1212),.clk(gclk));
	jor g1164(.dina(n1212),.dinb(w_n654_0[0]),.dout(n1213),.clk(gclk));
	jor g1165(.dina(n1213),.dinb(n1211),.dout(n1214),.clk(gclk));
	jor g1166(.dina(w_n287_0[0]),.dinb(w_n777_0[1]),.dout(n1215),.clk(gclk));
	jor g1167(.dina(w_n1215_0[1]),.dinb(w_n968_0[0]),.dout(n1216),.clk(gclk));
	jor g1168(.dina(n1216),.dinb(n1214),.dout(n1217),.clk(gclk));
	jand g1169(.dina(w_n92_1[0]),.dinb(w_n262_1[2]),.dout(n1218),.clk(gclk));
	jand g1170(.dina(w_n224_1[2]),.dinb(w_n98_1[0]),.dout(n1219),.clk(gclk));
	jor g1171(.dina(n1219),.dinb(n1218),.dout(n1220),.clk(gclk));
	jor g1172(.dina(w_n1094_0[0]),.dinb(n1220),.dout(n1221),.clk(gclk));
	jor g1173(.dina(n1221),.dinb(w_n700_0[0]),.dout(n1222),.clk(gclk));
	jor g1174(.dina(n1222),.dinb(w_n616_0[0]),.dout(n1223),.clk(gclk));
	jor g1175(.dina(n1223),.dinb(n1217),.dout(n1224),.clk(gclk));
	jand g1176(.dina(w_n1006_0[0]),.dinb(w_n527_2[0]),.dout(n1225),.clk(gclk));
	jand g1177(.dina(n1225),.dinb(w_n286_2[1]),.dout(n1226),.clk(gclk));
	jnot g1178(.din(w_n1226_0[1]),.dout(n1227),.clk(gclk));
	jor g1179(.dina(n1227),.dinb(n1224),.dout(n1228),.clk(gclk));
	jor g1180(.dina(n1228),.dinb(n1208),.dout(n1229),.clk(gclk));
	jor g1181(.dina(n1229),.dinb(n1190),.dout(n1230),.clk(gclk));
	jand g1182(.dina(n1230),.dinb(w_n987_0[2]),.dout(n1231),.clk(gclk));
	jor g1183(.dina(n1231),.dinb(w_n1055_1[1]),.dout(n1232),.clk(gclk));
	jnot g1184(.din(w_n1181_0[0]),.dout(n1233),.clk(gclk));
	jand g1185(.dina(n1233),.dinb(w_n1178_0[1]),.dout(n1234),.clk(gclk));
	jand g1186(.dina(n1234),.dinb(w_n1176_0[0]),.dout(n1235),.clk(gclk));
	jand g1187(.dina(w_n1235_0[1]),.dinb(w_n170_2[1]),.dout(n1236),.clk(gclk));
	jnot g1188(.din(w_n1189_0[0]),.dout(n1237),.clk(gclk));
	jand g1189(.dina(n1237),.dinb(n1236),.dout(n1238),.clk(gclk));
	jand g1190(.dina(w_n1205_0[0]),.dinb(w_n1060_0[0]),.dout(n1239),.clk(gclk));
	jand g1191(.dina(n1239),.dinb(w_n1196_1[0]),.dout(n1240),.clk(gclk));
	jand g1192(.dina(w_n1085_0[0]),.dinb(w_n290_2[1]),.dout(n1241),.clk(gclk));
	jand g1193(.dina(n1241),.dinb(w_n329_1[0]),.dout(n1242),.clk(gclk));
	jnot g1194(.din(w_n1215_0[0]),.dout(n1243),.clk(gclk));
	jand g1195(.dina(w_n1243_0[1]),.dinb(w_n586_0[1]),.dout(n1244),.clk(gclk));
	jand g1196(.dina(n1244),.dinb(n1242),.dout(n1245),.clk(gclk));
	jand g1197(.dina(w_n1095_2[1]),.dinb(w_n103_1[0]),.dout(n1246),.clk(gclk));
	jand g1198(.dina(n1246),.dinb(w_n218_2[0]),.dout(n1247),.clk(gclk));
	jand g1199(.dina(n1247),.dinb(w_n886_1[0]),.dout(n1248),.clk(gclk));
	jand g1200(.dina(n1248),.dinb(n1245),.dout(n1249),.clk(gclk));
	jand g1201(.dina(w_n1226_0[0]),.dinb(w_n1249_0[1]),.dout(n1250),.clk(gclk));
	jand g1202(.dina(w_n1250_0[1]),.dinb(n1240),.dout(n1251),.clk(gclk));
	jand g1203(.dina(n1251),.dinb(n1238),.dout(n1252),.clk(gclk));
	jand g1204(.dina(w_n1252_0[2]),.dinb(w_n607_2[0]),.dout(n1253),.clk(gclk));
	jor g1205(.dina(w_n1253_0[1]),.dinb(w_n1232_0[2]),.dout(n1254),.clk(gclk));
	jnot g1206(.din(w_n1254_2[1]),.dout(n1255),.clk(gclk));
	jand g1207(.dina(w_n56_0[0]),.dinb(w_n49_5[2]),.dout(n1256),.clk(gclk));
	jxor g1208(.dina(n1256),.dinb(w_a8_0[0]),.dout(n1257),.clk(gclk));
	jand g1209(.dina(w_n1257_13[2]),.dinb(w_n1255_2[1]),.dout(n1258),.clk(gclk));
	jnot g1210(.din(w_n1257_13[1]),.dout(n1259),.clk(gclk));
	jxor g1211(.dina(w_n1252_0[1]),.dinb(w_n607_1[2]),.dout(n1260),.clk(gclk));
	jand g1212(.dina(w_n1260_0[2]),.dinb(w_n1055_1[0]),.dout(n1261),.clk(gclk));
	jand g1213(.dina(w_n1261_2[2]),.dinb(w_n1259_9[1]),.dout(n1262),.clk(gclk));
	jor g1214(.dina(n1262),.dinb(n1258),.dout(n1263),.clk(gclk));
	jnot g1215(.din(n1263),.dout(n1264),.clk(gclk));
	jand g1216(.dina(w_n55_0[0]),.dinb(w_n49_5[1]),.dout(n1265),.clk(gclk));
	jxor g1217(.dina(n1265),.dinb(w_a7_0[0]),.dout(n1266),.clk(gclk));
	jnot g1218(.din(w_n1253_0[0]),.dout(n1267),.clk(gclk));
	jor g1219(.dina(w_n1252_0[0]),.dinb(w_n607_1[1]),.dout(n1268),.clk(gclk));
	jor g1220(.dina(w_n1268_0[1]),.dinb(w_n1055_0[2]),.dout(n1269),.clk(gclk));
	jand g1221(.dina(n1269),.dinb(n1267),.dout(n1270),.clk(gclk));
	jand g1222(.dina(w_n1270_3[2]),.dinb(w_n1266_6[1]),.dout(n1271),.clk(gclk));
	jnot g1223(.din(w_n1266_6[0]),.dout(n1272),.clk(gclk));
	jnot g1224(.din(w_n1016_1[0]),.dout(n1273),.clk(gclk));
	jnot g1225(.din(w_n1022_0[0]),.dout(n1274),.clk(gclk));
	jnot g1226(.din(w_n1024_0[1]),.dout(n1275),.clk(gclk));
	jnot g1227(.din(w_n1025_0[1]),.dout(n1276),.clk(gclk));
	jor g1228(.dina(w_n1026_0[0]),.dinb(n1276),.dout(n1277),.clk(gclk));
	jor g1229(.dina(n1277),.dinb(n1275),.dout(n1278),.clk(gclk));
	jnot g1230(.din(w_n1030_0[0]),.dout(n1279),.clk(gclk));
	jor g1231(.dina(n1279),.dinb(n1278),.dout(n1280),.clk(gclk));
	jor g1232(.dina(n1280),.dinb(n1274),.dout(n1281),.clk(gclk));
	jnot g1233(.din(w_n1039_0[1]),.dout(n1282),.clk(gclk));
	jnot g1234(.din(w_n234_0[0]),.dout(n1283),.clk(gclk));
	jor g1235(.dina(w_n1040_0[0]),.dinb(n1283),.dout(n1284),.clk(gclk));
	jnot g1236(.din(w_n1043_0[0]),.dout(n1285),.clk(gclk));
	jor g1237(.dina(n1285),.dinb(w_n401_0[0]),.dout(n1286),.clk(gclk));
	jor g1238(.dina(n1286),.dinb(n1284),.dout(n1287),.clk(gclk));
	jor g1239(.dina(n1287),.dinb(w_n624_0[0]),.dout(n1288),.clk(gclk));
	jor g1240(.dina(n1288),.dinb(n1282),.dout(n1289),.clk(gclk));
	jor g1241(.dina(n1289),.dinb(n1281),.dout(n1290),.clk(gclk));
	jnot g1242(.din(w_n1053_0[0]),.dout(n1291),.clk(gclk));
	jor g1243(.dina(n1291),.dinb(n1290),.dout(n1292),.clk(gclk));
	jor g1244(.dina(n1292),.dinb(n1273),.dout(n1293),.clk(gclk));
	jand g1245(.dina(w_n1268_0[0]),.dinb(n1293),.dout(n1294),.clk(gclk));
	jor g1246(.dina(w_n1260_0[1]),.dinb(w_n1294_0[2]),.dout(n1295),.clk(gclk));
	jand g1247(.dina(w_n1295_3[2]),.dinb(w_n1272_4[2]),.dout(n1296),.clk(gclk));
	jor g1248(.dina(n1296),.dinb(n1271),.dout(n1297),.clk(gclk));
	jand g1249(.dina(n1297),.dinb(n1264),.dout(n1298),.clk(gclk));
	jnot g1250(.din(n1298),.dout(n1299),.clk(gclk));
	jxor g1251(.dina(w_n1173_0[0]),.dinb(w_n1001_0[0]),.dout(n1300),.clk(gclk));
	jor g1252(.dina(w_n1300_0[1]),.dinb(w_n1299_0[1]),.dout(n1301),.clk(gclk));
	jand g1253(.dina(n1301),.dinb(n1175),.dout(n1302),.clk(gclk));
	jor g1254(.dina(w_n1302_0[1]),.dinb(w_n521_0[1]),.dout(n1303),.clk(gclk));
	jnot g1255(.din(w_n601_0[0]),.dout(n1304),.clk(gclk));
	jor g1256(.dina(w_n684_0[0]),.dinb(w_n966_0[0]),.dout(n1305),.clk(gclk));
	jor g1257(.dina(w_n689_0[0]),.dinb(w_n266_0[1]),.dout(n1306),.clk(gclk));
	jor g1258(.dina(n1306),.dinb(n1305),.dout(n1307),.clk(gclk));
	jnot g1259(.din(w_n1074_1[1]),.dout(n1308),.clk(gclk));
	jor g1260(.dina(w_n282_0[1]),.dinb(w_n749_0[0]),.dout(n1309),.clk(gclk));
	jor g1261(.dina(n1309),.dinb(n1308),.dout(n1310),.clk(gclk));
	jor g1262(.dina(n1310),.dinb(n1307),.dout(n1311),.clk(gclk));
	jor g1263(.dina(n1311),.dinb(n1304),.dout(n1312),.clk(gclk));
	jand g1264(.dina(w_n353_1[2]),.dinb(w_n197_2[0]),.dout(n1313),.clk(gclk));
	jand g1265(.dina(w_n280_1[2]),.dinb(w_n114_2[0]),.dout(n1314),.clk(gclk));
	jand g1266(.dina(n1314),.dinb(w_n1313_0[1]),.dout(n1315),.clk(gclk));
	jnot g1267(.din(n1315),.dout(n1316),.clk(gclk));
	jor g1268(.dina(n1316),.dinb(w_n1312_0[1]),.dout(n1317),.clk(gclk));
	jnot g1269(.din(w_n1105_0[1]),.dout(n1318),.clk(gclk));
	jor g1270(.dina(n1318),.dinb(w_n777_0[0]),.dout(n1319),.clk(gclk));
	jor g1271(.dina(w_n1319_0[1]),.dinb(w_n974_0[0]),.dout(n1320),.clk(gclk));
	jnot g1272(.din(n1320),.dout(n1321),.clk(gclk));
	jand g1273(.dina(w_n411_1[2]),.dinb(w_n265_1[2]),.dout(n1322),.clk(gclk));
	jand g1274(.dina(w_n1005_3[2]),.dinb(w_n439_3[1]),.dout(n1323),.clk(gclk));
	jand g1275(.dina(n1323),.dinb(w_n1322_1[2]),.dout(n1324),.clk(gclk));
	jand g1276(.dina(w_n1064_1[0]),.dinb(w_n826_0[0]),.dout(n1325),.clk(gclk));
	jand g1277(.dina(n1325),.dinb(n1324),.dout(n1326),.clk(gclk));
	jor g1278(.dina(w_n360_0[0]),.dinb(w_n652_0[0]),.dout(n1327),.clk(gclk));
	jnot g1279(.din(n1327),.dout(n1328),.clk(gclk));
	jand g1280(.dina(n1328),.dinb(w_n1130_0[0]),.dout(n1329),.clk(gclk));
	jand g1281(.dina(n1329),.dinb(n1326),.dout(n1330),.clk(gclk));
	jand g1282(.dina(n1330),.dinb(n1321),.dout(n1331),.clk(gclk));
	jand g1283(.dina(w_n409_1[0]),.dinb(w_n346_1[1]),.dout(n1332),.clk(gclk));
	jand g1284(.dina(w_n374_1[2]),.dinb(w_n288_1[1]),.dout(n1333),.clk(gclk));
	jand g1285(.dina(n1333),.dinb(w_n1332_0[1]),.dout(n1334),.clk(gclk));
	jand g1286(.dina(n1334),.dinb(w_n387_2[1]),.dout(n1335),.clk(gclk));
	jand g1287(.dina(w_n434_2[1]),.dinb(w_n255_1[1]),.dout(n1336),.clk(gclk));
	jand g1288(.dina(n1336),.dinb(w_n133_1[0]),.dout(n1337),.clk(gclk));
	jand g1289(.dina(n1337),.dinb(w_n561_0[2]),.dout(n1338),.clk(gclk));
	jand g1290(.dina(n1338),.dinb(n1335),.dout(n1339),.clk(gclk));
	jand g1291(.dina(w_n232_3[2]),.dinb(w_n206_1[1]),.dout(n1340),.clk(gclk));
	jand g1292(.dina(n1340),.dinb(w_n226_1[2]),.dout(n1341),.clk(gclk));
	jand g1293(.dina(w_n316_0[1]),.dinb(w_n148_0[2]),.dout(n1342),.clk(gclk));
	jand g1294(.dina(n1342),.dinb(n1341),.dout(n1343),.clk(gclk));
	jor g1295(.dina(w_n239_0[0]),.dinb(w_n119_0[0]),.dout(n1344),.clk(gclk));
	jnot g1296(.din(n1344),.dout(n1345),.clk(gclk));
	jand g1297(.dina(w_n852_1[0]),.dinb(w_n261_1[2]),.dout(n1346),.clk(gclk));
	jand g1298(.dina(w_n1346_0[1]),.dinb(w_n188_1[1]),.dout(n1347),.clk(gclk));
	jand g1299(.dina(n1347),.dinb(w_n1345_1[2]),.dout(n1348),.clk(gclk));
	jand g1300(.dina(n1348),.dinb(w_n1343_0[1]),.dout(n1349),.clk(gclk));
	jand g1301(.dina(n1349),.dinb(w_n1339_0[1]),.dout(n1350),.clk(gclk));
	jand g1302(.dina(n1350),.dinb(w_n1331_0[2]),.dout(n1351),.clk(gclk));
	jnot g1303(.din(n1351),.dout(n1352),.clk(gclk));
	jor g1304(.dina(n1352),.dinb(n1317),.dout(n1353),.clk(gclk));
	jnot g1305(.din(w_n1353_5[2]),.dout(n1354),.clk(gclk));
	jand g1306(.dina(w_n59_0[0]),.dinb(w_n49_5[0]),.dout(n1355),.clk(gclk));
	jxor g1307(.dina(n1355),.dinb(w_a11_0[0]),.dout(n1356),.clk(gclk));
	jand g1308(.dina(w_n1356_12[1]),.dinb(w_n1354_3[2]),.dout(n1357),.clk(gclk));
	jnot g1309(.din(n1357),.dout(n1358),.clk(gclk));
	jand g1310(.dina(w_n60_0[0]),.dinb(w_n49_4[2]),.dout(n1359),.clk(gclk));
	jxor g1311(.dina(n1359),.dinb(w_a12_0[0]),.dout(n1360),.clk(gclk));
	jand g1312(.dina(w_n1360_6[1]),.dinb(w_n1353_5[1]),.dout(n1361),.clk(gclk));
	jxor g1313(.dina(n1361),.dinb(w_n716_8[0]),.dout(n1362),.clk(gclk));
	jand g1314(.dina(n1362),.dinb(n1358),.dout(n1363),.clk(gclk));
	jand g1315(.dina(w_n1005_3[1]),.dinb(w_n207_2[0]),.dout(n1364),.clk(gclk));
	jand g1316(.dina(n1364),.dinb(w_n233_1[1]),.dout(n1365),.clk(gclk));
	jand g1317(.dina(w_n434_2[0]),.dinb(w_n415_1[2]),.dout(n1366),.clk(gclk));
	jand g1318(.dina(w_n387_2[0]),.dinb(w_n305_1[1]),.dout(n1367),.clk(gclk));
	jand g1319(.dina(n1367),.dinb(w_n1366_1[1]),.dout(n1368),.clk(gclk));
	jand g1320(.dina(n1368),.dinb(w_n1365_0[2]),.dout(n1369),.clk(gclk));
	jand g1321(.dina(w_n1345_1[1]),.dinb(w_n170_2[0]),.dout(n1370),.clk(gclk));
	jand g1322(.dina(n1370),.dinb(w_n1243_0[0]),.dout(n1371),.clk(gclk));
	jand g1323(.dina(w_n339_3[0]),.dinb(w_n157_2[2]),.dout(n1372),.clk(gclk));
	jand g1324(.dina(n1372),.dinb(w_n337_2[1]),.dout(n1373),.clk(gclk));
	jand g1325(.dina(n1373),.dinb(w_n488_2[2]),.dout(n1374),.clk(gclk));
	jand g1326(.dina(n1374),.dinb(n1371),.dout(n1375),.clk(gclk));
	jand g1327(.dina(w_n1375_0[1]),.dinb(w_n1346_0[0]),.dout(n1376),.clk(gclk));
	jand g1328(.dina(w_n345_0[0]),.dinb(w_n152_1[1]),.dout(n1377),.clk(gclk));
	jand g1329(.dina(n1377),.dinb(w_n276_2[0]),.dout(n1378),.clk(gclk));
	jand g1330(.dina(w_n1378_0[1]),.dinb(n1376),.dout(n1379),.clk(gclk));
	jand g1331(.dina(n1379),.dinb(n1369),.dout(n1380),.clk(gclk));
	jand g1332(.dina(n1380),.dinb(w_n1071_0[0]),.dout(n1381),.clk(gclk));
	jand g1333(.dina(w_n177_0[0]),.dinb(w_n103_0[2]),.dout(n1382),.clk(gclk));
	jand g1334(.dina(w_n438_1[1]),.dinb(w_n235_1[2]),.dout(n1383),.clk(gclk));
	jand g1335(.dina(n1383),.dinb(n1382),.dout(n1384),.clk(gclk));
	jand g1336(.dina(n1384),.dinb(w_n1097_0[0]),.dout(n1385),.clk(gclk));
	jand g1337(.dina(w_n1385_0[1]),.dinb(w_n460_2[2]),.dout(n1386),.clk(gclk));
	jand g1338(.dina(n1386),.dinb(w_n232_3[1]),.dout(n1387),.clk(gclk));
	jand g1339(.dina(w_n817_1[1]),.dinb(w_n382_1[0]),.dout(n1388),.clk(gclk));
	jand g1340(.dina(w_n594_0[1]),.dinb(w_n418_1[0]),.dout(n1389),.clk(gclk));
	jand g1341(.dina(w_n294_1[2]),.dinb(w_n286_2[0]),.dout(n1390),.clk(gclk));
	jand g1342(.dina(n1390),.dinb(n1389),.dout(n1391),.clk(gclk));
	jand g1343(.dina(n1391),.dinb(n1388),.dout(n1392),.clk(gclk));
	jand g1344(.dina(w_n1392_0[1]),.dinb(w_n281_0[0]),.dout(n1393),.clk(gclk));
	jand g1345(.dina(w_n862_0[0]),.dinb(w_n527_1[2]),.dout(n1394),.clk(gclk));
	jand g1346(.dina(n1394),.dinb(w_n842_0[0]),.dout(n1395),.clk(gclk));
	jand g1347(.dina(n1395),.dinb(w_n1322_1[1]),.dout(n1396),.clk(gclk));
	jand g1348(.dina(n1396),.dinb(w_n439_3[0]),.dout(n1397),.clk(gclk));
	jand g1349(.dina(n1397),.dinb(n1393),.dout(n1398),.clk(gclk));
	jand g1350(.dina(n1398),.dinb(w_n1387_0[1]),.dout(n1399),.clk(gclk));
	jand g1351(.dina(n1399),.dinb(w_n1381_0[1]),.dout(n1400),.clk(gclk));
	jor g1352(.dina(w_n1400_0[2]),.dinb(w_n1149_1[0]),.dout(n1401),.clk(gclk));
	jand g1353(.dina(n1401),.dinb(w_n486_1[1]),.dout(n1402),.clk(gclk));
	jxor g1354(.dina(w_n1400_0[1]),.dinb(w_n1149_0[2]),.dout(n1403),.clk(gclk));
	jand g1355(.dina(w_n1403_1[1]),.dinb(w_n519_5[1]),.dout(n1404),.clk(gclk));
	jnot g1356(.din(w_n1404_0[2]),.dout(n1405),.clk(gclk));
	jand g1357(.dina(n1405),.dinb(w_n1402_1[2]),.dout(n1406),.clk(gclk));
	jand g1358(.dina(w_n1406_0[1]),.dinb(w_n1363_0[1]),.dout(n1407),.clk(gclk));
	jand g1359(.dina(w_n1255_2[0]),.dinb(w_n880_5[2]),.dout(n1408),.clk(gclk));
	jand g1360(.dina(w_n1261_2[1]),.dinb(w_n881_4[1]),.dout(n1409),.clk(gclk));
	jor g1361(.dina(n1409),.dinb(n1408),.dout(n1410),.clk(gclk));
	jnot g1362(.din(n1410),.dout(n1411),.clk(gclk));
	jand g1363(.dina(w_n1270_3[1]),.dinb(w_n1257_13[0]),.dout(n1412),.clk(gclk));
	jand g1364(.dina(w_n1295_3[1]),.dinb(w_n1259_9[0]),.dout(n1413),.clk(gclk));
	jor g1365(.dina(n1413),.dinb(n1412),.dout(n1414),.clk(gclk));
	jand g1366(.dina(n1414),.dinb(n1411),.dout(n1415),.clk(gclk));
	jnot g1367(.din(w_n1152_2[0]),.dout(n1416),.clk(gclk));
	jand g1368(.dina(w_n1168_4[1]),.dinb(w_n1416_2[1]),.dout(n1417),.clk(gclk));
	jnot g1369(.din(w_n1160_2[0]),.dout(n1418),.clk(gclk));
	jand g1370(.dina(w_n1166_5[2]),.dinb(w_n1418_2[2]),.dout(n1419),.clk(gclk));
	jor g1371(.dina(n1419),.dinb(n1417),.dout(n1420),.clk(gclk));
	jnot g1372(.din(n1420),.dout(n1421),.clk(gclk));
	jand g1373(.dina(w_n1266_5[2]),.dinb(w_n1164_3[1]),.dout(n1422),.clk(gclk));
	jand g1374(.dina(w_n1272_4[1]),.dinb(w_n1170_4[0]),.dout(n1423),.clk(gclk));
	jor g1375(.dina(n1423),.dinb(n1422),.dout(n1424),.clk(gclk));
	jand g1376(.dina(n1424),.dinb(n1421),.dout(n1425),.clk(gclk));
	jxor g1377(.dina(w_n1425_0[1]),.dinb(w_n1415_0[1]),.dout(n1426),.clk(gclk));
	jxor g1378(.dina(w_n1426_0[1]),.dinb(w_n1407_0[1]),.dout(n1427),.clk(gclk));
	jnot g1379(.din(w_n1427_0[1]),.dout(n1428),.clk(gclk));
	jxor g1380(.dina(w_n1302_0[0]),.dinb(w_n521_0[0]),.dout(n1429),.clk(gclk));
	jnot g1381(.din(w_n1429_0[1]),.dout(n1430),.clk(gclk));
	jor g1382(.dina(n1430),.dinb(n1428),.dout(n1431),.clk(gclk));
	jand g1383(.dina(n1431),.dinb(n1303),.dout(n1432),.clk(gclk));
	jand g1384(.dina(w_n61_0[0]),.dinb(w_n49_4[1]),.dout(n1433),.clk(gclk));
	jxor g1385(.dina(n1433),.dinb(w_a13_0[0]),.dout(n1434),.clk(gclk));
	jand g1386(.dina(w_n1434_6[2]),.dinb(w_n1354_3[1]),.dout(n1435),.clk(gclk));
	jnot g1387(.din(n1435),.dout(n1436),.clk(gclk));
	jand g1388(.dina(w_n62_0[0]),.dinb(w_n49_4[0]),.dout(n1437),.clk(gclk));
	jxor g1389(.dina(n1437),.dinb(w_a14_0[0]),.dout(n1438),.clk(gclk));
	jand g1390(.dina(w_n1438_21[1]),.dinb(w_n1353_5[0]),.dout(n1439),.clk(gclk));
	jxor g1391(.dina(n1439),.dinb(w_n716_7[2]),.dout(n1440),.clk(gclk));
	jand g1392(.dina(n1440),.dinb(n1436),.dout(n1441),.clk(gclk));
	jand g1393(.dina(w_n516_0[1]),.dinb(w_n486_1[0]),.dout(n1442),.clk(gclk));
	jand g1394(.dina(w_n1343_0[0]),.dinb(w_n361_2[0]),.dout(n1443),.clk(gclk));
	jand g1395(.dina(n1443),.dinb(w_n252_3[0]),.dout(n1444),.clk(gclk));
	jand g1396(.dina(w_n569_1[1]),.dinb(w_n321_2[0]),.dout(n1445),.clk(gclk));
	jand g1397(.dina(n1445),.dinb(w_n575_0[0]),.dout(n1446),.clk(gclk));
	jand g1398(.dina(n1446),.dinb(w_n381_0[0]),.dout(n1447),.clk(gclk));
	jand g1399(.dina(w_n347_1[2]),.dinb(w_n102_2[2]),.dout(n1448),.clk(gclk));
	jand g1400(.dina(w_n269_1[0]),.dinb(w_n191_2[0]),.dout(n1449),.clk(gclk));
	jand g1401(.dina(n1449),.dinb(w_n173_0[2]),.dout(n1450),.clk(gclk));
	jand g1402(.dina(n1450),.dinb(w_n1448_0[1]),.dout(n1451),.clk(gclk));
	jand g1403(.dina(w_n290_2[0]),.dinb(w_n233_1[0]),.dout(n1452),.clk(gclk));
	jand g1404(.dina(w_n1452_0[1]),.dinb(w_n157_2[1]),.dout(n1453),.clk(gclk));
	jand g1405(.dina(n1453),.dinb(n1451),.dout(n1454),.clk(gclk));
	jand g1406(.dina(n1454),.dinb(w_n1447_0[1]),.dout(n1455),.clk(gclk));
	jand g1407(.dina(n1455),.dinb(w_n1444_0[1]),.dout(n1456),.clk(gclk));
	jand g1408(.dina(w_n249_0[2]),.dinb(w_n99_1[0]),.dout(n1457),.clk(gclk));
	jor g1409(.dina(n1457),.dinb(w_n134_0[1]),.dout(n1458),.clk(gclk));
	jand g1410(.dina(w_n1005_3[0]),.dinb(w_n283_1[2]),.dout(n1459),.clk(gclk));
	jand g1411(.dina(w_n587_2[2]),.dinb(w_n182_2[2]),.dout(n1460),.clk(gclk));
	jand g1412(.dina(w_n309_1[2]),.dinb(w_n403_0[0]),.dout(n1461),.clk(gclk));
	jand g1413(.dina(n1461),.dinb(w_n1460_1[2]),.dout(n1462),.clk(gclk));
	jand g1414(.dina(n1462),.dinb(w_n1459_0[2]),.dout(n1463),.clk(gclk));
	jand g1415(.dina(w_n384_2[1]),.dinb(w_n221_2[1]),.dout(n1464),.clk(gclk));
	jand g1416(.dina(n1464),.dinb(w_n170_1[2]),.dout(n1465),.clk(gclk));
	jand g1417(.dina(n1465),.dinb(w_n919_0[0]),.dout(n1466),.clk(gclk));
	jand g1418(.dina(n1466),.dinb(n1463),.dout(n1467),.clk(gclk));
	jand g1419(.dina(w_n279_0[0]),.dinb(w_n159_0[1]),.dout(n1468),.clk(gclk));
	jand g1420(.dina(n1468),.dinb(w_n534_2[0]),.dout(n1469),.clk(gclk));
	jand g1421(.dina(n1469),.dinb(w_n215_2[2]),.dout(n1470),.clk(gclk));
	jand g1422(.dina(w_n1470_0[1]),.dinb(w_n1064_0[2]),.dout(n1471),.clk(gclk));
	jand g1423(.dina(n1471),.dinb(w_n1467_0[1]),.dout(n1472),.clk(gclk));
	jand g1424(.dina(n1472),.dinb(n1458),.dout(n1473),.clk(gclk));
	jand g1425(.dina(n1473),.dinb(w_n1456_0[1]),.dout(n1474),.clk(gclk));
	jxor g1426(.dina(w_n1494_6[1]),.dinb(w_n1441_0[1]),.dout(n1478),.clk(gclk));
	jnot g1427(.din(w_n1478_0[1]),.dout(n1479),.clk(gclk));
	jnot g1428(.din(w_n1356_12[0]),.dout(n1480),.clk(gclk));
	jand g1429(.dina(w_n1480_10[1]),.dinb(w_n878_1[1]),.dout(n1481),.clk(gclk));
	jand g1430(.dina(w_n1356_11[2]),.dinb(w_n989_2[0]),.dout(n1482),.clk(gclk));
	jor g1431(.dina(n1482),.dinb(n1481),.dout(n1483),.clk(gclk));
	jand g1432(.dina(w_n1360_6[0]),.dinb(w_n992_3[1]),.dout(n1484),.clk(gclk));
	jnot g1433(.din(w_n1360_5[2]),.dout(n1485),.clk(gclk));
	jand g1434(.dina(w_n1485_4[2]),.dinb(w_n997_4[0]),.dout(n1486),.clk(gclk));
	jor g1435(.dina(n1486),.dinb(n1484),.dout(n1487),.clk(gclk));
	jnot g1436(.din(n1487),.dout(n1488),.clk(gclk));
	jor g1437(.dina(n1488),.dinb(n1483),.dout(n1489),.clk(gclk));
	jnot g1438(.din(w_n517_0[1]),.dout(n1490),.clk(gclk));
	jnot g1439(.din(w_n486_0[2]),.dout(n1491),.clk(gclk));
	jnot g1440(.din(w_n516_0[0]),.dout(n1492),.clk(gclk));
	jand g1441(.dina(n1492),.dinb(w_n1491_0[1]),.dout(n1493),.clk(gclk));
	jnot g1442(.din(w_n1474_7[1]),.dout(n1494),.clk(gclk));
	jand g1443(.dina(w_n1493_5[1]),.dinb(w_n519_5[0]),.dout(n1497),.clk(gclk));
	jand g1444(.dina(w_n52_0[0]),.dinb(w_n49_3[2]),.dout(n1498),.clk(gclk));
	jxor g1445(.dina(n1498),.dinb(w_a4_0[0]),.dout(n1499),.clk(gclk));
	jnot g1446(.din(w_n1499_5[2]),.dout(n1500),.clk(gclk));
	jxor g1447(.dina(w_n1500_5[1]),.dinb(w_n1474_7[0]),.dout(n1501),.clk(gclk));
	jor g1448(.dina(n1501),.dinb(w_n1490_5[1]),.dout(n1502),.clk(gclk));
	jnot g1449(.din(n1502),.dout(n1503),.clk(gclk));
	jnot g1450(.din(w_n519_4[2]),.dout(n1504),.clk(gclk));
	jand g1451(.dina(w_n1474_6[2]),.dinb(w_n1490_5[0]),.dout(n1505),.clk(gclk));
	jand g1452(.dina(w_n1505_4[2]),.dinb(w_n1504_3[2]),.dout(n1506),.clk(gclk));
	jor g1453(.dina(n1506),.dinb(n1503),.dout(n1507),.clk(gclk));
	jor g1454(.dina(n1507),.dinb(n1497),.dout(n1508),.clk(gclk));
	jand g1455(.dina(w_n1508_0[1]),.dinb(w_n1489_0[1]),.dout(n1509),.clk(gclk));
	jnot g1456(.din(w_n1509_0[1]),.dout(n1510),.clk(gclk));
	jor g1457(.dina(w_n1508_0[0]),.dinb(w_n1489_0[0]),.dout(n1511),.clk(gclk));
	jand g1458(.dina(w_n1511_0[1]),.dinb(w_n1478_0[0]),.dout(n1512),.clk(gclk));
	jand g1459(.dina(n1512),.dinb(n1510),.dout(n1513),.clk(gclk));
	jor g1460(.dina(w_n1513_0[1]),.dinb(n1479),.dout(n1514),.clk(gclk));
	jnot g1461(.din(w_n1511_0[0]),.dout(n1515),.clk(gclk));
	jor g1462(.dina(w_n1513_0[0]),.dinb(n1515),.dout(n1516),.clk(gclk));
	jor g1463(.dina(w_n1516_0[2]),.dinb(w_n1509_0[0]),.dout(n1517),.clk(gclk));
	jand g1464(.dina(n1517),.dinb(n1514),.dout(n1518),.clk(gclk));
	jor g1465(.dina(w_n1518_0[1]),.dinb(w_n1432_0[1]),.dout(n1519),.clk(gclk));
	jxor g1466(.dina(w_n1518_0[0]),.dinb(w_n1432_0[0]),.dout(n1520),.clk(gclk));
	jand g1467(.dina(w_n1425_0[0]),.dinb(w_n1415_0[0]),.dout(n1521),.clk(gclk));
	jand g1468(.dina(w_n1426_0[0]),.dinb(w_n1407_0[0]),.dout(n1522),.clk(gclk));
	jor g1469(.dina(n1522),.dinb(n1521),.dout(n1523),.clk(gclk));
	jand g1470(.dina(w_n1360_5[1]),.dinb(w_n1354_3[0]),.dout(n1524),.clk(gclk));
	jnot g1471(.din(n1524),.dout(n1525),.clk(gclk));
	jand g1472(.dina(w_n1434_6[1]),.dinb(w_n1353_4[2]),.dout(n1526),.clk(gclk));
	jxor g1473(.dina(n1526),.dinb(w_n716_7[1]),.dout(n1527),.clk(gclk));
	jand g1474(.dina(n1527),.dinb(n1525),.dout(n1528),.clk(gclk));
	jnot g1475(.din(w_n997_3[2]),.dout(n1529),.clk(gclk));
	jand g1476(.dina(w_n1480_10[0]),.dinb(w_n1529_0[2]),.dout(n1530),.clk(gclk));
	jor g1477(.dina(w_n876_0[2]),.dinb(w_n930_2[0]),.dout(n1531),.clk(gclk));
	jand g1478(.dina(w_n1531_0[1]),.dinb(w_n987_0[1]),.dout(n1532),.clk(gclk));
	jor g1479(.dina(w_n813_0[0]),.dinb(w_n716_7[0]),.dout(n1533),.clk(gclk));
	jand g1480(.dina(w_n1533_0[1]),.dinb(w_n1532_0[2]),.dout(n1534),.clk(gclk));
	jand g1481(.dina(w_n1356_11[1]),.dinb(w_n1534_0[2]),.dout(n1535),.clk(gclk));
	jor g1482(.dina(n1535),.dinb(n1530),.dout(n1536),.clk(gclk));
	jnot g1483(.din(n1536),.dout(n1537),.clk(gclk));
	jor g1484(.dina(w_n1531_0[0]),.dinb(w_n607_1[0]),.dout(n1538),.clk(gclk));
	jand g1485(.dina(n1538),.dinb(w_n1533_0[0]),.dout(n1539),.clk(gclk));
	jand g1486(.dina(w_n994_5[2]),.dinb(w_n1539_2[2]),.dout(n1540),.clk(gclk));
	jxor g1487(.dina(w_n876_0[1]),.dinb(w_n930_1[2]),.dout(n1541),.clk(gclk));
	jor g1488(.dina(w_n1541_0[1]),.dinb(w_n1532_0[1]),.dout(n1542),.clk(gclk));
	jand g1489(.dina(w_n996_4[1]),.dinb(w_n1542_2[2]),.dout(n1543),.clk(gclk));
	jor g1490(.dina(n1543),.dinb(n1540),.dout(n1544),.clk(gclk));
	jand g1491(.dina(n1544),.dinb(n1537),.dout(n1545),.clk(gclk));
	jand g1492(.dina(w_n1545_0[1]),.dinb(w_n1528_0[1]),.dout(n1546),.clk(gclk));
	jand g1493(.dina(w_n1400_0[0]),.dinb(w_n1149_0[1]),.dout(n1547),.clk(gclk));
	jnot g1494(.din(w_n1547_0[1]),.dout(n1548),.clk(gclk));
	jand g1495(.dina(n1548),.dinb(w_n1402_1[1]),.dout(n1549),.clk(gclk));
	jand g1496(.dina(w_n1549_4[2]),.dinb(w_n1154_10[0]),.dout(n1550),.clk(gclk));
	jand g1497(.dina(w_n1403_1[0]),.dinb(w_n1491_0[0]),.dout(n1551),.clk(gclk));
	jand g1498(.dina(w_n1551_4[2]),.dinb(w_n1156_12[0]),.dout(n1552),.clk(gclk));
	jor g1499(.dina(n1552),.dinb(n1550),.dout(n1553),.clk(gclk));
	jnot g1500(.din(n1553),.dout(n1554),.clk(gclk));
	jnot g1501(.din(w_n1403_0[2]),.dout(n1555),.clk(gclk));
	jor g1502(.dina(w_n1547_0[0]),.dinb(w_n486_0[1]),.dout(n1556),.clk(gclk));
	jand g1503(.dina(w_n1556_0[1]),.dinb(w_n1555_0[1]),.dout(n1557),.clk(gclk));
	jnot g1504(.din(w_n1557_0[1]),.dout(n1558),.clk(gclk));
	jand g1505(.dina(w_n1558_4[1]),.dinb(w_n1499_5[1]),.dout(n1559),.clk(gclk));
	jor g1506(.dina(w_n1403_0[1]),.dinb(w_n1402_1[0]),.dout(n1560),.clk(gclk));
	jand g1507(.dina(w_n1560_4[2]),.dinb(w_n1500_5[0]),.dout(n1561),.clk(gclk));
	jor g1508(.dina(n1561),.dinb(n1559),.dout(n1562),.clk(gclk));
	jand g1509(.dina(n1562),.dinb(n1554),.dout(n1563),.clk(gclk));
	jxor g1510(.dina(w_n1545_0[0]),.dinb(w_n1528_0[0]),.dout(n1564),.clk(gclk));
	jand g1511(.dina(w_n1564_0[1]),.dinb(w_n1563_0[1]),.dout(n1565),.clk(gclk));
	jor g1512(.dina(n1565),.dinb(n1546),.dout(n1566),.clk(gclk));
	jxor g1513(.dina(w_n1566_0[1]),.dinb(w_n1523_0[1]),.dout(n1567),.clk(gclk));
	jand g1514(.dina(w_n1255_1[2]),.dinb(w_n994_5[1]),.dout(n1568),.clk(gclk));
	jand g1515(.dina(w_n1261_2[0]),.dinb(w_n996_4[0]),.dout(n1569),.clk(gclk));
	jor g1516(.dina(n1569),.dinb(n1568),.dout(n1570),.clk(gclk));
	jnot g1517(.din(n1570),.dout(n1571),.clk(gclk));
	jand g1518(.dina(w_n1270_3[0]),.dinb(w_n880_5[1]),.dout(n1572),.clk(gclk));
	jand g1519(.dina(w_n1295_3[0]),.dinb(w_n881_4[0]),.dout(n1573),.clk(gclk));
	jor g1520(.dina(n1573),.dinb(n1572),.dout(n1574),.clk(gclk));
	jand g1521(.dina(n1574),.dinb(n1571),.dout(n1575),.clk(gclk));
	jnot g1522(.din(w_n1170_3[2]),.dout(n1576),.clk(gclk));
	jand g1523(.dina(w_n1259_8[2]),.dinb(w_n1576_0[2]),.dout(n1577),.clk(gclk));
	jand g1524(.dina(w_n1257_12[2]),.dinb(w_n1163_0[1]),.dout(n1578),.clk(gclk));
	jor g1525(.dina(n1578),.dinb(n1577),.dout(n1579),.clk(gclk));
	jnot g1526(.din(n1579),.dout(n1580),.clk(gclk));
	jand g1527(.dina(w_n1266_5[1]),.dinb(w_n1160_1[2]),.dout(n1581),.clk(gclk));
	jand g1528(.dina(w_n1272_4[0]),.dinb(w_n1152_1[2]),.dout(n1582),.clk(gclk));
	jor g1529(.dina(n1582),.dinb(n1581),.dout(n1583),.clk(gclk));
	jand g1530(.dina(n1583),.dinb(n1580),.dout(n1584),.clk(gclk));
	jand g1531(.dina(w_n1551_4[1]),.dinb(w_n1168_4[0]),.dout(n1585),.clk(gclk));
	jand g1532(.dina(w_n1549_4[1]),.dinb(w_n1166_5[1]),.dout(n1586),.clk(gclk));
	jor g1533(.dina(n1586),.dinb(n1585),.dout(n1587),.clk(gclk));
	jnot g1534(.din(n1587),.dout(n1588),.clk(gclk));
	jand g1535(.dina(w_n1558_4[0]),.dinb(w_n1154_9[2]),.dout(n1589),.clk(gclk));
	jand g1536(.dina(w_n1560_4[1]),.dinb(w_n1156_11[2]),.dout(n1590),.clk(gclk));
	jor g1537(.dina(n1590),.dinb(n1589),.dout(n1591),.clk(gclk));
	jand g1538(.dina(n1591),.dinb(n1588),.dout(n1592),.clk(gclk));
	jxor g1539(.dina(w_n1592_0[1]),.dinb(w_n1584_0[1]),.dout(n1593),.clk(gclk));
	jxor g1540(.dina(w_n1593_0[1]),.dinb(w_n1575_0[1]),.dout(n1594),.clk(gclk));
	jxor g1541(.dina(w_n1594_0[1]),.dinb(w_n1567_0[1]),.dout(n1595),.clk(gclk));
	jand g1542(.dina(w_n1595_0[1]),.dinb(w_n1520_0[1]),.dout(n1596),.clk(gclk));
	jnot g1543(.din(n1596),.dout(n1597),.clk(gclk));
	jand g1544(.dina(n1597),.dinb(n1519),.dout(n1598),.clk(gclk));
	jand g1545(.dina(w_n1566_0[0]),.dinb(w_n1523_0[0]),.dout(n1599),.clk(gclk));
	jand g1546(.dina(w_n1594_0[0]),.dinb(w_n1567_0[0]),.dout(n1600),.clk(gclk));
	jor g1547(.dina(n1600),.dinb(n1599),.dout(n1601),.clk(gclk));
	jand g1548(.dina(w_n1592_0[0]),.dinb(w_n1584_0[0]),.dout(n1602),.clk(gclk));
	jand g1549(.dina(w_n1593_0[0]),.dinb(w_n1575_0[0]),.dout(n1603),.clk(gclk));
	jor g1550(.dina(n1603),.dinb(n1602),.dout(n1604),.clk(gclk));
	jand g1551(.dina(w_n1494_6[0]),.dinb(w_n1441_0[0]),.dout(n1605),.clk(gclk));
	jand g1552(.dina(w_n1499_5[0]),.dinb(w_n1493_5[0]),.dout(n1606),.clk(gclk));
	jnot g1553(.din(n1606),.dout(n1607),.clk(gclk));
	jxor g1554(.dina(w_n1474_6[1]),.dinb(w_n1156_11[1]),.dout(n1608),.clk(gclk));
	jor g1555(.dina(n1608),.dinb(w_n1490_4[2]),.dout(n1609),.clk(gclk));
	jand g1556(.dina(w_n1505_4[1]),.dinb(w_n1500_4[2]),.dout(n1610),.clk(gclk));
	jnot g1557(.din(n1610),.dout(n1611),.clk(gclk));
	jand g1558(.dina(n1611),.dinb(n1609),.dout(n1612),.clk(gclk));
	jand g1559(.dina(n1612),.dinb(n1607),.dout(n1613),.clk(gclk));
	jxor g1560(.dina(w_n1613_0[1]),.dinb(w_n1605_0[1]),.dout(n1614),.clk(gclk));
	jxor g1561(.dina(w_n1614_0[1]),.dinb(w_n1604_0[1]),.dout(n1615),.clk(gclk));
	jxor g1562(.dina(w_n1615_0[1]),.dinb(w_n1601_0[1]),.dout(n1616),.clk(gclk));
	jand g1563(.dina(w_n1485_4[1]),.dinb(w_n878_1[0]),.dout(n1617),.clk(gclk));
	jand g1564(.dina(w_n1360_5[0]),.dinb(w_n989_1[2]),.dout(n1618),.clk(gclk));
	jor g1565(.dina(n1618),.dinb(n1617),.dout(n1619),.clk(gclk));
	jnot g1566(.din(n1619),.dout(n1620),.clk(gclk));
	jand g1567(.dina(w_n1434_6[0]),.dinb(w_n992_3[0]),.dout(n1621),.clk(gclk));
	jnot g1568(.din(w_n1434_5[2]),.dout(n1622),.clk(gclk));
	jand g1569(.dina(w_n1622_4[1]),.dinb(w_n997_3[1]),.dout(n1623),.clk(gclk));
	jor g1570(.dina(n1623),.dinb(n1621),.dout(n1624),.clk(gclk));
	jand g1571(.dina(n1624),.dinb(n1620),.dout(n1625),.clk(gclk));
	jand g1572(.dina(w_n1494_5[2]),.dinb(w_n519_4[1]),.dout(n1626),.clk(gclk));
	jand g1573(.dina(w_n1438_21[0]),.dinb(w_n1354_2[2]),.dout(n1627),.clk(gclk));
	jor g1574(.dina(n1627),.dinb(w_n930_1[1]),.dout(n1628),.clk(gclk));
	jnot g1575(.din(n1628),.dout(n1629),.clk(gclk));
	jxor g1576(.dina(w_n1629_0[1]),.dinb(w_n1626_0[1]),.dout(n1630),.clk(gclk));
	jxor g1577(.dina(w_n1630_0[1]),.dinb(w_n1625_0[1]),.dout(n1631),.clk(gclk));
	jxor g1578(.dina(w_n1631_0[1]),.dinb(w_n1516_0[1]),.dout(n1632),.clk(gclk));
	jand g1579(.dina(w_n1551_4[0]),.dinb(w_n1272_3[2]),.dout(n1633),.clk(gclk));
	jand g1580(.dina(w_n1549_4[0]),.dinb(w_n1266_5[0]),.dout(n1634),.clk(gclk));
	jor g1581(.dina(n1634),.dinb(n1633),.dout(n1635),.clk(gclk));
	jnot g1582(.din(n1635),.dout(n1636),.clk(gclk));
	jand g1583(.dina(w_n1558_3[2]),.dinb(w_n1166_5[0]),.dout(n1637),.clk(gclk));
	jand g1584(.dina(w_n1560_4[0]),.dinb(w_n1168_3[2]),.dout(n1638),.clk(gclk));
	jor g1585(.dina(n1638),.dinb(n1637),.dout(n1639),.clk(gclk));
	jand g1586(.dina(n1639),.dinb(n1636),.dout(n1640),.clk(gclk));
	jand g1587(.dina(w_n1259_8[1]),.dinb(w_n1416_2[0]),.dout(n1641),.clk(gclk));
	jand g1588(.dina(w_n1257_12[1]),.dinb(w_n1418_2[1]),.dout(n1642),.clk(gclk));
	jor g1589(.dina(n1642),.dinb(n1641),.dout(n1643),.clk(gclk));
	jnot g1590(.din(n1643),.dout(n1644),.clk(gclk));
	jand g1591(.dina(w_n1164_3[0]),.dinb(w_n880_5[0]),.dout(n1645),.clk(gclk));
	jand g1592(.dina(w_n1170_3[1]),.dinb(w_n881_3[2]),.dout(n1646),.clk(gclk));
	jor g1593(.dina(n1646),.dinb(n1645),.dout(n1647),.clk(gclk));
	jand g1594(.dina(n1647),.dinb(n1644),.dout(n1648),.clk(gclk));
	jnot g1595(.din(w_n1295_2[2]),.dout(n1649),.clk(gclk));
	jand g1596(.dina(w_n1649_0[2]),.dinb(w_n996_3[2]),.dout(n1650),.clk(gclk));
	jnot g1597(.din(w_n1270_2[2]),.dout(n1651),.clk(gclk));
	jand g1598(.dina(w_n1651_1[1]),.dinb(w_n994_5[0]),.dout(n1652),.clk(gclk));
	jor g1599(.dina(n1652),.dinb(n1650),.dout(n1653),.clk(gclk));
	jnot g1600(.din(n1653),.dout(n1654),.clk(gclk));
	jand g1601(.dina(w_n1356_11[0]),.dinb(w_n1254_2[0]),.dout(n1655),.clk(gclk));
	jnot g1602(.din(w_n1261_1[2]),.dout(n1656),.clk(gclk));
	jand g1603(.dina(w_n1480_9[2]),.dinb(w_n1656_1[2]),.dout(n1657),.clk(gclk));
	jor g1604(.dina(n1657),.dinb(n1655),.dout(n1658),.clk(gclk));
	jand g1605(.dina(n1658),.dinb(n1654),.dout(n1659),.clk(gclk));
	jxor g1606(.dina(w_n1659_0[1]),.dinb(w_n1648_0[1]),.dout(n1660),.clk(gclk));
	jxor g1607(.dina(w_n1660_0[1]),.dinb(w_n1640_0[1]),.dout(n1661),.clk(gclk));
	jxor g1608(.dina(w_n1661_0[1]),.dinb(w_n1632_0[1]),.dout(n1662),.clk(gclk));
	jxor g1609(.dina(w_n1662_0[1]),.dinb(w_n1616_0[1]),.dout(n1663),.clk(gclk));
	jxor g1610(.dina(w_n1663_0[1]),.dinb(w_n1598_0[1]),.dout(n1664),.clk(gclk));
	jand g1611(.dina(w_n1551_3[2]),.dinb(w_n1500_4[1]),.dout(n1665),.clk(gclk));
	jand g1612(.dina(w_n1549_3[2]),.dinb(w_n1499_4[2]),.dout(n1666),.clk(gclk));
	jor g1613(.dina(n1666),.dinb(n1665),.dout(n1667),.clk(gclk));
	jnot g1614(.din(n1667),.dout(n1668),.clk(gclk));
	jor g1615(.dina(w_n1557_0[0]),.dinb(w_n1504_3[1]),.dout(n1669),.clk(gclk));
	jnot g1616(.din(n1669),.dout(n1670),.clk(gclk));
	jand g1617(.dina(w_n1560_3[2]),.dinb(w_n1504_3[0]),.dout(n1671),.clk(gclk));
	jor g1618(.dina(n1671),.dinb(n1670),.dout(n1672),.clk(gclk));
	jand g1619(.dina(n1672),.dinb(n1668),.dout(n1673),.clk(gclk));
	jxor g1620(.dina(w_n1406_0[0]),.dinb(w_n1363_0[0]),.dout(n1674),.clk(gclk));
	jand g1621(.dina(w_n1674_0[1]),.dinb(w_n1673_0[1]),.dout(n1675),.clk(gclk));
	jand g1622(.dina(w_n1354_2[1]),.dinb(w_n994_4[2]),.dout(n1676),.clk(gclk));
	jnot g1623(.din(n1676),.dout(n1677),.clk(gclk));
	jand g1624(.dina(w_n1356_10[2]),.dinb(w_n1353_4[1]),.dout(n1678),.clk(gclk));
	jxor g1625(.dina(n1678),.dinb(w_n716_6[2]),.dout(n1679),.clk(gclk));
	jand g1626(.dina(n1679),.dinb(n1677),.dout(n1680),.clk(gclk));
	jor g1627(.dina(w_n1257_12[0]),.dinb(w_n1542_2[1]),.dout(n1681),.clk(gclk));
	jor g1628(.dina(w_n1259_8[0]),.dinb(w_n1539_2[1]),.dout(n1682),.clk(gclk));
	jand g1629(.dina(n1682),.dinb(n1681),.dout(n1683),.clk(gclk));
	jand g1630(.dina(w_n992_2[2]),.dinb(w_n880_4[2]),.dout(n1684),.clk(gclk));
	jand g1631(.dina(w_n997_3[0]),.dinb(w_n881_3[1]),.dout(n1685),.clk(gclk));
	jor g1632(.dina(n1685),.dinb(n1684),.dout(n1686),.clk(gclk));
	jand g1633(.dina(n1686),.dinb(n1683),.dout(n1687),.clk(gclk));
	jand g1634(.dina(w_n1687_0[1]),.dinb(w_n1680_0[1]),.dout(n1688),.clk(gclk));
	jand g1635(.dina(w_n1266_4[2]),.dinb(w_n1255_1[1]),.dout(n1689),.clk(gclk));
	jand g1636(.dina(w_n1272_3[1]),.dinb(w_n1261_1[1]),.dout(n1690),.clk(gclk));
	jor g1637(.dina(n1690),.dinb(n1689),.dout(n1691),.clk(gclk));
	jnot g1638(.din(n1691),.dout(n1692),.clk(gclk));
	jand g1639(.dina(w_n1270_2[1]),.dinb(w_n1166_4[2]),.dout(n1693),.clk(gclk));
	jand g1640(.dina(w_n1295_2[1]),.dinb(w_n1168_3[1]),.dout(n1694),.clk(gclk));
	jor g1641(.dina(n1694),.dinb(n1693),.dout(n1695),.clk(gclk));
	jand g1642(.dina(n1695),.dinb(n1692),.dout(n1696),.clk(gclk));
	jxor g1643(.dina(w_n1687_0[0]),.dinb(w_n1680_0[0]),.dout(n1697),.clk(gclk));
	jand g1644(.dina(w_n1697_0[1]),.dinb(w_n1696_0[1]),.dout(n1698),.clk(gclk));
	jor g1645(.dina(n1698),.dinb(n1688),.dout(n1699),.clk(gclk));
	jxor g1646(.dina(w_n1674_0[0]),.dinb(w_n1673_0[0]),.dout(n1700),.clk(gclk));
	jand g1647(.dina(w_n1700_0[1]),.dinb(w_n1699_0[1]),.dout(n1701),.clk(gclk));
	jor g1648(.dina(n1701),.dinb(n1675),.dout(n1702),.clk(gclk));
	jxor g1649(.dina(w_n1564_0[0]),.dinb(w_n1563_0[0]),.dout(n1703),.clk(gclk));
	jand g1650(.dina(w_n1703_0[1]),.dinb(w_n1702_0[1]),.dout(n1704),.clk(gclk));
	jxor g1651(.dina(w_n1429_0[0]),.dinb(w_n1427_0[0]),.dout(n1705),.clk(gclk));
	jxor g1652(.dina(w_n1703_0[0]),.dinb(w_n1702_0[0]),.dout(n1706),.clk(gclk));
	jand g1653(.dina(w_n1706_0[1]),.dinb(w_n1705_0[1]),.dout(n1707),.clk(gclk));
	jor g1654(.dina(n1707),.dinb(n1704),.dout(n1708),.clk(gclk));
	jxor g1655(.dina(w_n1595_0[0]),.dinb(w_n1520_0[0]),.dout(n1709),.clk(gclk));
	jand g1656(.dina(w_n1709_0[1]),.dinb(w_n1708_0[1]),.dout(n1710),.clk(gclk));
	jnot g1657(.din(w_n1710_0[1]),.dout(n1711),.clk(gclk));
	jor g1658(.dina(w_n1266_4[1]),.dinb(w_n1542_2[0]),.dout(n1712),.clk(gclk));
	jor g1659(.dina(w_n1272_3[0]),.dinb(w_n1539_2[0]),.dout(n1713),.clk(gclk));
	jand g1660(.dina(n1713),.dinb(n1712),.dout(n1714),.clk(gclk));
	jand g1661(.dina(w_n1257_11[2]),.dinb(w_n992_2[1]),.dout(n1715),.clk(gclk));
	jand g1662(.dina(w_n1259_7[2]),.dinb(w_n997_2[2]),.dout(n1716),.clk(gclk));
	jor g1663(.dina(n1716),.dinb(n1715),.dout(n1717),.clk(gclk));
	jand g1664(.dina(n1717),.dinb(n1714),.dout(n1718),.clk(gclk));
	jor g1665(.dina(w_n1254_1[2]),.dinb(w_n1168_3[0]),.dout(n1719),.clk(gclk));
	jor g1666(.dina(w_n1656_1[1]),.dinb(w_n1166_4[1]),.dout(n1720),.clk(gclk));
	jand g1667(.dina(n1720),.dinb(n1719),.dout(n1721),.clk(gclk));
	jand g1668(.dina(w_n1270_2[0]),.dinb(w_n1154_9[1]),.dout(n1722),.clk(gclk));
	jand g1669(.dina(w_n1295_2[0]),.dinb(w_n1156_11[0]),.dout(n1723),.clk(gclk));
	jor g1670(.dina(n1723),.dinb(n1722),.dout(n1724),.clk(gclk));
	jand g1671(.dina(n1724),.dinb(n1721),.dout(n1725),.clk(gclk));
	jand g1672(.dina(w_n1725_0[1]),.dinb(w_n1718_0[1]),.dout(n1726),.clk(gclk));
	jor g1673(.dina(w_n1499_4[1]),.dinb(w_n1170_3[0]),.dout(n1727),.clk(gclk));
	jor g1674(.dina(w_n1500_4[0]),.dinb(w_n1164_2[2]),.dout(n1728),.clk(gclk));
	jand g1675(.dina(n1728),.dinb(n1727),.dout(n1729),.clk(gclk));
	jand g1676(.dina(w_n1160_1[1]),.dinb(w_n519_4[0]),.dout(n1730),.clk(gclk));
	jand g1677(.dina(w_n1152_1[1]),.dinb(w_n1504_2[2]),.dout(n1731),.clk(gclk));
	jor g1678(.dina(n1731),.dinb(n1730),.dout(n1732),.clk(gclk));
	jand g1679(.dina(n1732),.dinb(n1729),.dout(n1733),.clk(gclk));
	jxor g1680(.dina(w_n1725_0[0]),.dinb(w_n1718_0[0]),.dout(n1734),.clk(gclk));
	jand g1681(.dina(w_n1734_0[1]),.dinb(w_n1733_0[1]),.dout(n1735),.clk(gclk));
	jor g1682(.dina(n1735),.dinb(n1726),.dout(n1736),.clk(gclk));
	jxor g1683(.dina(w_n1697_0[0]),.dinb(w_n1696_0[0]),.dout(n1737),.clk(gclk));
	jand g1684(.dina(w_n1737_0[1]),.dinb(w_n1736_0[1]),.dout(n1738),.clk(gclk));
	jand g1685(.dina(w_n1354_2[0]),.dinb(w_n880_4[1]),.dout(n1739),.clk(gclk));
	jnot g1686(.din(n1739),.dout(n1740),.clk(gclk));
	jand g1687(.dina(w_n1353_4[0]),.dinb(w_n994_4[1]),.dout(n1741),.clk(gclk));
	jxor g1688(.dina(n1741),.dinb(w_n716_6[1]),.dout(n1742),.clk(gclk));
	jand g1689(.dina(n1742),.dinb(n1740),.dout(n1743),.clk(gclk));
	jand g1690(.dina(w_n1115_0[1]),.dinb(w_n519_3[2]),.dout(n1744),.clk(gclk));
	jnot g1691(.din(w_n1744_0[2]),.dout(n1745),.clk(gclk));
	jand g1692(.dina(n1745),.dinb(w_n1151_1[0]),.dout(n1746),.clk(gclk));
	jand g1693(.dina(w_n1746_0[1]),.dinb(w_n1743_0[1]),.dout(n1747),.clk(gclk));
	jor g1694(.dina(w_n1499_4[0]),.dinb(w_n1152_1[0]),.dout(n1748),.clk(gclk));
	jor g1695(.dina(w_n1500_3[2]),.dinb(w_n1160_1[0]),.dout(n1749),.clk(gclk));
	jand g1696(.dina(n1749),.dinb(n1748),.dout(n1750),.clk(gclk));
	jand g1697(.dina(w_n1164_2[1]),.dinb(w_n1154_9[0]),.dout(n1751),.clk(gclk));
	jand g1698(.dina(w_n1170_2[2]),.dinb(w_n1156_10[2]),.dout(n1752),.clk(gclk));
	jor g1699(.dina(n1752),.dinb(n1751),.dout(n1753),.clk(gclk));
	jand g1700(.dina(n1753),.dinb(n1750),.dout(n1754),.clk(gclk));
	jxor g1701(.dina(w_n1754_0[1]),.dinb(w_n1747_0[1]),.dout(n1755),.clk(gclk));
	jxor g1702(.dina(w_n1755_0[1]),.dinb(w_n1404_0[1]),.dout(n1756),.clk(gclk));
	jxor g1703(.dina(w_n1737_0[0]),.dinb(w_n1736_0[0]),.dout(n1757),.clk(gclk));
	jand g1704(.dina(w_n1757_0[1]),.dinb(w_n1756_0[1]),.dout(n1758),.clk(gclk));
	jor g1705(.dina(n1758),.dinb(n1738),.dout(n1759),.clk(gclk));
	jnot g1706(.din(w_n1759_0[1]),.dout(n1760),.clk(gclk));
	jand g1707(.dina(w_n1754_0[0]),.dinb(w_n1747_0[0]),.dout(n1761),.clk(gclk));
	jand g1708(.dina(w_n1755_0[0]),.dinb(w_n1404_0[0]),.dout(n1762),.clk(gclk));
	jor g1709(.dina(n1762),.dinb(n1761),.dout(n1763),.clk(gclk));
	jxor g1710(.dina(w_n1300_0[0]),.dinb(w_n1299_0[0]),.dout(n1764),.clk(gclk));
	jxor g1711(.dina(w_n1764_0[1]),.dinb(w_n1763_0[1]),.dout(n1765),.clk(gclk));
	jxor g1712(.dina(w_n1700_0[0]),.dinb(w_n1699_0[0]),.dout(n1766),.clk(gclk));
	jxor g1713(.dina(w_n1766_0[1]),.dinb(w_n1765_0[1]),.dout(n1767),.clk(gclk));
	jnot g1714(.din(w_n1767_0[2]),.dout(n1768),.clk(gclk));
	jxor g1715(.dina(w_n1746_0[0]),.dinb(w_n1743_0[0]),.dout(n1769),.clk(gclk));
	jnot g1716(.din(n1769),.dout(n1770),.clk(gclk));
	jand g1717(.dina(w_n1168_2[2]),.dinb(w_n878_0[2]),.dout(n1771),.clk(gclk));
	jand g1718(.dina(w_n1166_4[0]),.dinb(w_n989_1[1]),.dout(n1772),.clk(gclk));
	jor g1719(.dina(n1772),.dinb(n1771),.dout(n1773),.clk(gclk));
	jand g1720(.dina(w_n1266_4[0]),.dinb(w_n992_2[0]),.dout(n1774),.clk(gclk));
	jand g1721(.dina(w_n1272_2[2]),.dinb(w_n997_2[1]),.dout(n1775),.clk(gclk));
	jor g1722(.dina(n1775),.dinb(n1774),.dout(n1776),.clk(gclk));
	jnot g1723(.din(n1776),.dout(n1777),.clk(gclk));
	jor g1724(.dina(n1777),.dinb(n1773),.dout(n1778),.clk(gclk));
	jand g1725(.dina(w_n1354_1[2]),.dinb(w_n1257_11[1]),.dout(n1779),.clk(gclk));
	jnot g1726(.din(n1779),.dout(n1780),.clk(gclk));
	jand g1727(.dina(w_n1353_3[2]),.dinb(w_n880_4[0]),.dout(n1781),.clk(gclk));
	jxor g1728(.dina(n1781),.dinb(w_n716_6[0]),.dout(n1782),.clk(gclk));
	jand g1729(.dina(n1782),.dinb(n1780),.dout(n1783),.clk(gclk));
	jnot g1730(.din(w_n1783_0[1]),.dout(n1784),.clk(gclk));
	jor g1731(.dina(n1784),.dinb(w_n1778_0[1]),.dout(n1785),.clk(gclk));
	jand g1732(.dina(w_n1255_1[0]),.dinb(w_n1154_8[2]),.dout(n1786),.clk(gclk));
	jand g1733(.dina(w_n1261_1[0]),.dinb(w_n1156_10[1]),.dout(n1787),.clk(gclk));
	jor g1734(.dina(n1787),.dinb(n1786),.dout(n1788),.clk(gclk));
	jand g1735(.dina(w_n1499_3[2]),.dinb(w_n1270_1[2]),.dout(n1789),.clk(gclk));
	jand g1736(.dina(w_n1500_3[1]),.dinb(w_n1295_1[2]),.dout(n1790),.clk(gclk));
	jor g1737(.dina(n1790),.dinb(n1789),.dout(n1791),.clk(gclk));
	jnot g1738(.din(n1791),.dout(n1792),.clk(gclk));
	jor g1739(.dina(n1792),.dinb(n1788),.dout(n1793),.clk(gclk));
	jxor g1740(.dina(w_n1783_0[0]),.dinb(w_n1778_0[0]),.dout(n1794),.clk(gclk));
	jor g1741(.dina(w_n1794_0[1]),.dinb(w_n1793_0[1]),.dout(n1795),.clk(gclk));
	jand g1742(.dina(n1795),.dinb(n1785),.dout(n1796),.clk(gclk));
	jor g1743(.dina(w_n1796_0[1]),.dinb(w_n1770_0[1]),.dout(n1797),.clk(gclk));
	jnot g1744(.din(n1797),.dout(n1798),.clk(gclk));
	jxor g1745(.dina(w_n1796_0[0]),.dinb(w_n1770_0[0]),.dout(n1799),.clk(gclk));
	jxor g1746(.dina(w_n1734_0[0]),.dinb(w_n1733_0[0]),.dout(n1800),.clk(gclk));
	jand g1747(.dina(w_n1800_0[1]),.dinb(w_n1799_0[1]),.dout(n1801),.clk(gclk));
	jor g1748(.dina(n1801),.dinb(n1798),.dout(n1802),.clk(gclk));
	jnot g1749(.din(w_n1802_0[1]),.dout(n1803),.clk(gclk));
	jxor g1750(.dina(w_n1757_0[0]),.dinb(w_n1756_0[0]),.dout(n1804),.clk(gclk));
	jnot g1751(.din(w_n1804_0[1]),.dout(n1805),.clk(gclk));
	jand g1752(.dina(n1805),.dinb(n1803),.dout(n1806),.clk(gclk));
	jand g1753(.dina(w_n1354_1[1]),.dinb(w_n1266_3[2]),.dout(n1807),.clk(gclk));
	jnot g1754(.din(n1807),.dout(n1808),.clk(gclk));
	jand g1755(.dina(w_n1353_3[1]),.dinb(w_n1257_11[0]),.dout(n1809),.clk(gclk));
	jxor g1756(.dina(n1809),.dinb(w_n716_5[2]),.dout(n1810),.clk(gclk));
	jand g1757(.dina(n1810),.dinb(n1808),.dout(n1811),.clk(gclk));
	jnot g1758(.din(w_n1260_0[0]),.dout(n1812),.clk(gclk));
	jor g1759(.dina(w_n1812_0[1]),.dinb(w_n1504_2[1]),.dout(n1813),.clk(gclk));
	jand g1760(.dina(w_n1813_1[1]),.dinb(w_n1294_0[1]),.dout(n1814),.clk(gclk));
	jand g1761(.dina(w_n1814_0[1]),.dinb(w_n1811_0[1]),.dout(n1815),.clk(gclk));
	jand g1762(.dina(w_n1815_0[1]),.dinb(w_n1744_0[1]),.dout(n1816),.clk(gclk));
	jor g1763(.dina(w_n1168_2[1]),.dinb(w_n992_1[2]),.dout(n1817),.clk(gclk));
	jor g1764(.dina(w_n1166_3[2]),.dinb(w_n997_2[0]),.dout(n1818),.clk(gclk));
	jand g1765(.dina(n1818),.dinb(n1817),.dout(n1819),.clk(gclk));
	jand g1766(.dina(w_n1154_8[1]),.dinb(w_n1539_1[2]),.dout(n1820),.clk(gclk));
	jand g1767(.dina(w_n1156_10[0]),.dinb(w_n1542_1[2]),.dout(n1821),.clk(gclk));
	jor g1768(.dina(n1821),.dinb(n1820),.dout(n1822),.clk(gclk));
	jand g1769(.dina(n1822),.dinb(n1819),.dout(n1823),.clk(gclk));
	jor g1770(.dina(w_n1295_1[1]),.dinb(w_n519_3[1]),.dout(n1824),.clk(gclk));
	jor g1771(.dina(w_n1270_1[1]),.dinb(w_n1504_2[0]),.dout(n1825),.clk(gclk));
	jand g1772(.dina(n1825),.dinb(n1824),.dout(n1826),.clk(gclk));
	jand g1773(.dina(w_n1499_3[1]),.dinb(w_n1254_1[1]),.dout(n1827),.clk(gclk));
	jand g1774(.dina(w_n1500_3[0]),.dinb(w_n1656_1[0]),.dout(n1828),.clk(gclk));
	jor g1775(.dina(n1828),.dinb(n1827),.dout(n1829),.clk(gclk));
	jand g1776(.dina(n1829),.dinb(n1826),.dout(n1830),.clk(gclk));
	jand g1777(.dina(w_n1830_0[1]),.dinb(w_n1823_0[1]),.dout(n1831),.clk(gclk));
	jxor g1778(.dina(w_n1814_0[0]),.dinb(w_n1811_0[0]),.dout(n1832),.clk(gclk));
	jxor g1779(.dina(w_n1830_0[0]),.dinb(w_n1823_0[0]),.dout(n1833),.clk(gclk));
	jand g1780(.dina(w_n1833_0[1]),.dinb(w_n1832_0[1]),.dout(n1834),.clk(gclk));
	jor g1781(.dina(n1834),.dinb(n1831),.dout(n1835),.clk(gclk));
	jxor g1782(.dina(w_n1815_0[0]),.dinb(w_n1744_0[0]),.dout(n1836),.clk(gclk));
	jand g1783(.dina(w_n1836_0[1]),.dinb(w_n1835_0[1]),.dout(n1837),.clk(gclk));
	jor g1784(.dina(n1837),.dinb(n1816),.dout(n1838),.clk(gclk));
	jxor g1785(.dina(w_n1800_0[0]),.dinb(w_n1799_0[0]),.dout(n1839),.clk(gclk));
	jor g1786(.dina(w_n1839_0[1]),.dinb(w_n1838_0[1]),.dout(n1840),.clk(gclk));
	jnot g1787(.din(w_n1840_0[1]),.dout(n1841),.clk(gclk));
	jxor g1788(.dina(w_n1836_0[0]),.dinb(w_n1835_0[0]),.dout(n1842),.clk(gclk));
	jxor g1789(.dina(w_n1794_0[0]),.dinb(w_n1793_0[0]),.dout(n1843),.clk(gclk));
	jand g1790(.dina(w_n1843_0[1]),.dinb(w_n1842_0[1]),.dout(n1844),.clk(gclk));
	jnot g1791(.din(w_n1844_0[1]),.dout(n1845),.clk(gclk));
	jor g1792(.dina(w_n1843_0[0]),.dinb(w_n1842_0[0]),.dout(n1846),.clk(gclk));
	jnot g1793(.din(w_n1846_0[1]),.dout(n1847),.clk(gclk));
	jand g1794(.dina(w_n877_0[0]),.dinb(w_n519_3[0]),.dout(n1848),.clk(gclk));
	jnot g1795(.din(n1848),.dout(n1849),.clk(gclk));
	jand g1796(.dina(w_n1541_0[0]),.dinb(w_n519_2[2]),.dout(n1850),.clk(gclk));
	jand g1797(.dina(w_n1850_0[1]),.dinb(w_n1353_3[0]),.dout(n1851),.clk(gclk));
	jand g1798(.dina(w_n1500_2[2]),.dinb(w_n716_5[1]),.dout(n1852),.clk(gclk));
	jor g1799(.dina(n1852),.dinb(n1851),.dout(n1853),.clk(gclk));
	jand g1800(.dina(w_n1156_9[2]),.dinb(w_n930_1[0]),.dout(n1854),.clk(gclk));
	jand g1801(.dina(w_n1154_8[0]),.dinb(w_n716_5[0]),.dout(n1855),.clk(gclk));
	jand g1802(.dina(n1855),.dinb(w_n1353_2[2]),.dout(n1856),.clk(gclk));
	jor g1803(.dina(n1856),.dinb(n1854),.dout(n1857),.clk(gclk));
	jnot g1804(.din(n1857),.dout(n1858),.clk(gclk));
	jand g1805(.dina(n1858),.dinb(n1853),.dout(n1859),.clk(gclk));
	jand g1806(.dina(n1859),.dinb(n1849),.dout(n1860),.clk(gclk));
	jnot g1807(.din(w_n1860_0[1]),.dout(n1861),.clk(gclk));
	jor g1808(.dina(w_n1353_2[1]),.dinb(w_n1156_9[1]),.dout(n1862),.clk(gclk));
	jand g1809(.dina(w_n1353_2[0]),.dinb(w_n1166_3[1]),.dout(n1863),.clk(gclk));
	jxor g1810(.dina(n1863),.dinb(w_n716_4[2]),.dout(n1864),.clk(gclk));
	jand g1811(.dina(n1864),.dinb(n1862),.dout(n1865),.clk(gclk));
	jor g1812(.dina(w_n1850_0[0]),.dinb(w_n815_0[2]),.dout(n1866),.clk(gclk));
	jnot g1813(.din(n1866),.dout(n1867),.clk(gclk));
	jxor g1814(.dina(w_n1867_0[1]),.dinb(w_n1865_0[1]),.dout(n1868),.clk(gclk));
	jnot g1815(.din(w_n1868_0[2]),.dout(n1869),.clk(gclk));
	jor g1816(.dina(w_n878_0[1]),.dinb(w_n519_2[1]),.dout(n1870),.clk(gclk));
	jor g1817(.dina(w_n989_1[0]),.dinb(w_n1504_1[2]),.dout(n1871),.clk(gclk));
	jand g1818(.dina(n1871),.dinb(n1870),.dout(n1872),.clk(gclk));
	jor g1819(.dina(w_n1499_3[0]),.dinb(w_n997_1[2]),.dout(n1873),.clk(gclk));
	jnot g1820(.din(w_n1873_0[1]),.dout(n1874),.clk(gclk));
	jand g1821(.dina(w_n1499_2[2]),.dinb(w_n1534_0[1]),.dout(n1875),.clk(gclk));
	jor g1822(.dina(n1875),.dinb(n1874),.dout(n1876),.clk(gclk));
	jor g1823(.dina(n1876),.dinb(n1872),.dout(n1877),.clk(gclk));
	jor g1824(.dina(n1877),.dinb(n1869),.dout(n1878),.clk(gclk));
	jand g1825(.dina(n1878),.dinb(n1861),.dout(n1879),.clk(gclk));
	jand g1826(.dina(w_n1542_1[1]),.dinb(w_n1504_1[1]),.dout(n1880),.clk(gclk));
	jand g1827(.dina(w_n1539_1[1]),.dinb(w_n519_2[0]),.dout(n1881),.clk(gclk));
	jor g1828(.dina(n1881),.dinb(n1880),.dout(n1882),.clk(gclk));
	jor g1829(.dina(w_n1500_2[1]),.dinb(w_n992_1[1]),.dout(n1883),.clk(gclk));
	jand g1830(.dina(n1883),.dinb(w_n1873_0[0]),.dout(n1884),.clk(gclk));
	jand g1831(.dina(n1884),.dinb(n1882),.dout(n1885),.clk(gclk));
	jor g1832(.dina(w_n1885_0[1]),.dinb(w_n1868_0[1]),.dout(n1886),.clk(gclk));
	jnot g1833(.din(w_n1886_0[1]),.dout(n1887),.clk(gclk));
	jor g1834(.dina(n1887),.dinb(n1879),.dout(n1888),.clk(gclk));
	jor g1835(.dina(w_n1888_0[1]),.dinb(w_n1813_1[0]),.dout(n1889),.clk(gclk));
	jand g1836(.dina(w_n1867_0[0]),.dinb(w_n1865_0[0]),.dout(n1890),.clk(gclk));
	jand g1837(.dina(w_n1354_1[0]),.dinb(w_n1166_3[0]),.dout(n1891),.clk(gclk));
	jnot g1838(.din(n1891),.dout(n1892),.clk(gclk));
	jand g1839(.dina(w_n1353_1[2]),.dinb(w_n1266_3[1]),.dout(n1893),.clk(gclk));
	jxor g1840(.dina(n1893),.dinb(w_n716_4[1]),.dout(n1894),.clk(gclk));
	jand g1841(.dina(n1894),.dinb(n1892),.dout(n1895),.clk(gclk));
	jor g1842(.dina(w_n1500_2[0]),.dinb(w_n1539_1[0]),.dout(n1896),.clk(gclk));
	jor g1843(.dina(w_n1499_2[1]),.dinb(w_n1542_1[0]),.dout(n1897),.clk(gclk));
	jand g1844(.dina(n1897),.dinb(n1896),.dout(n1898),.clk(gclk));
	jand g1845(.dina(w_n1154_7[2]),.dinb(w_n992_1[0]),.dout(n1899),.clk(gclk));
	jand g1846(.dina(w_n1156_9[0]),.dinb(w_n997_1[1]),.dout(n1900),.clk(gclk));
	jor g1847(.dina(n1900),.dinb(n1899),.dout(n1901),.clk(gclk));
	jand g1848(.dina(n1901),.dinb(n1898),.dout(n1902),.clk(gclk));
	jxor g1849(.dina(w_n1902_0[2]),.dinb(w_n1895_0[2]),.dout(n1903),.clk(gclk));
	jxor g1850(.dina(w_n1903_0[1]),.dinb(w_n1890_0[2]),.dout(n1904),.clk(gclk));
	jnot g1851(.din(w_n1904_0[1]),.dout(n1905),.clk(gclk));
	jand g1852(.dina(n1905),.dinb(n1889),.dout(n1906),.clk(gclk));
	jand g1853(.dina(w_n1888_0[0]),.dinb(w_n1813_0[2]),.dout(n1907),.clk(gclk));
	jxor g1854(.dina(w_n1833_0[0]),.dinb(w_n1832_0[0]),.dout(n1908),.clk(gclk));
	jnot g1855(.din(w_n1908_0[2]),.dout(n1909),.clk(gclk));
	jand g1856(.dina(w_n1902_0[1]),.dinb(w_n1895_0[1]),.dout(n1910),.clk(gclk));
	jnot g1857(.din(w_n1910_0[1]),.dout(n1911),.clk(gclk));
	jnot g1858(.din(w_n1890_0[1]),.dout(n1912),.clk(gclk));
	jnot g1859(.din(w_n1895_0[0]),.dout(n1913),.clk(gclk));
	jxor g1860(.dina(w_n1902_0[0]),.dinb(n1913),.dout(n1914),.clk(gclk));
	jor g1861(.dina(n1914),.dinb(n1912),.dout(n1915),.clk(gclk));
	jand g1862(.dina(n1915),.dinb(n1911),.dout(n1916),.clk(gclk));
	jand g1863(.dina(n1916),.dinb(n1909),.dout(n1917),.clk(gclk));
	jor g1864(.dina(n1917),.dinb(n1907),.dout(n1918),.clk(gclk));
	jor g1865(.dina(n1918),.dinb(n1906),.dout(n1919),.clk(gclk));
	jand g1866(.dina(w_n1903_0[0]),.dinb(w_n1890_0[0]),.dout(n1920),.clk(gclk));
	jor g1867(.dina(n1920),.dinb(w_n1910_0[0]),.dout(n1921),.clk(gclk));
	jand g1868(.dina(w_n1921_0[1]),.dinb(w_n1908_0[1]),.dout(n1922),.clk(gclk));
	jnot g1869(.din(w_n1922_0[1]),.dout(n1923),.clk(gclk));
	jand g1870(.dina(n1923),.dinb(n1919),.dout(n1924),.clk(gclk));
	jor g1871(.dina(n1924),.dinb(n1847),.dout(n1925),.clk(gclk));
	jand g1872(.dina(n1925),.dinb(n1845),.dout(n1926),.clk(gclk));
	jor g1873(.dina(n1926),.dinb(n1841),.dout(n1927),.clk(gclk));
	jand g1874(.dina(w_n1804_0[0]),.dinb(w_n1802_0[0]),.dout(n1928),.clk(gclk));
	jand g1875(.dina(w_n1839_0[0]),.dinb(w_n1838_0[0]),.dout(n1929),.clk(gclk));
	jor g1876(.dina(n1929),.dinb(n1928),.dout(n1930),.clk(gclk));
	jnot g1877(.din(w_n1930_0[1]),.dout(n1931),.clk(gclk));
	jand g1878(.dina(n1931),.dinb(n1927),.dout(n1932),.clk(gclk));
	jor g1879(.dina(n1932),.dinb(w_n1806_0[1]),.dout(n1933),.clk(gclk));
	jand g1880(.dina(w_n1933_0[1]),.dinb(w_n1768_0[1]),.dout(n1934),.clk(gclk));
	jor g1881(.dina(n1934),.dinb(n1760),.dout(n1935),.clk(gclk));
	jand g1882(.dina(w_n1764_0[0]),.dinb(w_n1763_0[0]),.dout(n1936),.clk(gclk));
	jand g1883(.dina(w_n1766_0[0]),.dinb(w_n1765_0[0]),.dout(n1937),.clk(gclk));
	jor g1884(.dina(n1937),.dinb(n1936),.dout(n1938),.clk(gclk));
	jxor g1885(.dina(w_n1706_0[0]),.dinb(w_n1705_0[0]),.dout(n1939),.clk(gclk));
	jand g1886(.dina(w_n1939_0[1]),.dinb(w_n1938_0[1]),.dout(n1940),.clk(gclk));
	jnot g1887(.din(w_n1940_0[1]),.dout(n1941),.clk(gclk));
	jor g1888(.dina(w_n1933_0[0]),.dinb(w_n1768_0[0]),.dout(n1942),.clk(gclk));
	jand g1889(.dina(n1942),.dinb(n1941),.dout(n1943),.clk(gclk));
	jand g1890(.dina(n1943),.dinb(n1935),.dout(n1944),.clk(gclk));
	jnot g1891(.din(w_n1938_0[0]),.dout(n1945),.clk(gclk));
	jnot g1892(.din(w_n1939_0[0]),.dout(n1946),.clk(gclk));
	jand g1893(.dina(n1946),.dinb(n1945),.dout(n1947),.clk(gclk));
	jnot g1894(.din(n1947),.dout(n1948),.clk(gclk));
	jor g1895(.dina(w_n1709_0[0]),.dinb(w_n1708_0[0]),.dout(n1949),.clk(gclk));
	jand g1896(.dina(n1949),.dinb(n1948),.dout(n1950),.clk(gclk));
	jnot g1897(.din(w_n1950_0[1]),.dout(n1951),.clk(gclk));
	jor g1898(.dina(n1951),.dinb(n1944),.dout(n1952),.clk(gclk));
	jand g1899(.dina(n1952),.dinb(n1711),.dout(n1953),.clk(gclk));
	jxor g1900(.dina(w_n1953_0[1]),.dinb(w_n1664_0[2]),.dout(n1954),.clk(gclk));
	jxor g1901(.dina(w_n1954_0[1]),.dinb(w_n425_0[1]),.dout(n1955),.clk(gclk));
	jnot g1902(.din(w_n1955_0[2]),.dout(n1956),.clk(gclk));
	jxor g1903(.dina(w_n1360_4[2]),.dinb(w_n1480_9[1]),.dout(n1957),.clk(gclk));
	jnot g1904(.din(w_n1957_0[2]),.dout(n1958),.clk(gclk));
	jand g1905(.dina(w_n1958_1[1]),.dinb(w_n1956_7[1]),.dout(n1959),.clk(gclk));
	jand g1906(.dina(w_n1954_0[0]),.dinb(w_n425_0[0]),.dout(n1960),.clk(gclk));
	jand g1907(.dina(w_n445_1[1]),.dinb(w_n327_0[2]),.dout(n1961),.clk(gclk));
	jand g1908(.dina(w_n337_2[0]),.dinb(w_n215_2[1]),.dout(n1962),.clk(gclk));
	jand g1909(.dina(w_n467_1[1]),.dinb(w_n147_1[1]),.dout(n1963),.clk(gclk));
	jand g1910(.dina(n1963),.dinb(w_n1962_0[1]),.dout(n1964),.clk(gclk));
	jand g1911(.dina(n1964),.dinb(w_n924_0[1]),.dout(n1965),.clk(gclk));
	jand g1912(.dina(w_n1965_0[1]),.dinb(w_n526_0[0]),.dout(n1966),.clk(gclk));
	jand g1913(.dina(w_n534_1[2]),.dinb(w_n290_1[2]),.dout(n1967),.clk(gclk));
	jand g1914(.dina(w_n462_1[1]),.dinb(w_n176_1[0]),.dout(n1968),.clk(gclk));
	jand g1915(.dina(n1968),.dinb(w_n353_1[1]),.dout(n1969),.clk(gclk));
	jand g1916(.dina(n1969),.dinb(n1967),.dout(n1970),.clk(gclk));
	jand g1917(.dina(w_n510_2[1]),.dinb(w_n415_1[1]),.dout(n1971),.clk(gclk));
	jand g1918(.dina(n1971),.dinb(w_n460_2[1]),.dout(n1972),.clk(gclk));
	jand g1919(.dina(n1972),.dinb(w_n1970_0[1]),.dout(n1973),.clk(gclk));
	jand g1920(.dina(n1973),.dinb(n1966),.dout(n1974),.clk(gclk));
	jand g1921(.dina(w_n1974_0[1]),.dinb(w_n1961_0[2]),.dout(n1975),.clk(gclk));
	jand g1922(.dina(w_n1087_0[1]),.dinb(w_n297_0[2]),.dout(n1976),.clk(gclk));
	jand g1923(.dina(w_n321_1[2]),.dinb(w_n213_2[1]),.dout(n1977),.clk(gclk));
	jand g1924(.dina(n1977),.dinb(w_n1005_2[2]),.dout(n1978),.clk(gclk));
	jand g1925(.dina(w_n188_1[0]),.dinb(w_n157_2[0]),.dout(n1979),.clk(gclk));
	jand g1926(.dina(w_n1979_0[1]),.dinb(n1978),.dout(n1980),.clk(gclk));
	jand g1927(.dina(n1980),.dinb(n1976),.dout(n1981),.clk(gclk));
	jand g1928(.dina(w_n1024_0[0]),.dinb(w_n276_1[2]),.dout(n1982),.clk(gclk));
	jand g1929(.dina(w_n546_0[0]),.dinb(w_n207_1[2]),.dout(n1983),.clk(gclk));
	jand g1930(.dina(w_n448_1[1]),.dinb(w_n389_3[0]),.dout(n1984),.clk(gclk));
	jand g1931(.dina(w_n1984_0[1]),.dinb(w_n588_0[1]),.dout(n1985),.clk(gclk));
	jand g1932(.dina(n1985),.dinb(n1983),.dout(n1986),.clk(gclk));
	jand g1933(.dina(n1986),.dinb(n1982),.dout(n1987),.clk(gclk));
	jand g1934(.dina(w_n437_0[2]),.dinb(w_n103_0[1]),.dout(n1988),.clk(gclk));
	jand g1935(.dina(n1988),.dinb(w_n383_1[2]),.dout(n1989),.clk(gclk));
	jand g1936(.dina(n1989),.dinb(w_n1987_0[2]),.dout(n1990),.clk(gclk));
	jand g1937(.dina(n1990),.dinb(w_n489_2[1]),.dout(n1991),.clk(gclk));
	jand g1938(.dina(n1991),.dinb(n1981),.dout(n1992),.clk(gclk));
	jand g1939(.dina(n1992),.dinb(n1975),.dout(n1993),.clk(gclk));
	jnot g1940(.din(w_n1993_0[2]),.dout(n1994),.clk(gclk));
	jnot g1941(.din(w_n1598_0[0]),.dout(n1995),.clk(gclk));
	jand g1942(.dina(w_n1663_0[0]),.dinb(n1995),.dout(n1996),.clk(gclk));
	jnot g1943(.din(w_n1664_0[1]),.dout(n1997),.clk(gclk));
	jnot g1944(.din(w_n1806_0[0]),.dout(n1998),.clk(gclk));
	jnot g1945(.din(w_n1813_0[1]),.dout(n1999),.clk(gclk));
	jand g1946(.dina(w_n1885_0[0]),.dinb(w_n1868_0[0]),.dout(n2000),.clk(gclk));
	jor g1947(.dina(n2000),.dinb(w_n1860_0[0]),.dout(n2001),.clk(gclk));
	jand g1948(.dina(w_n1886_0[0]),.dinb(n2001),.dout(n2002),.clk(gclk));
	jand g1949(.dina(w_n2002_0[1]),.dinb(w_n1999_0[1]),.dout(n2003),.clk(gclk));
	jor g1950(.dina(w_n1904_0[0]),.dinb(n2003),.dout(n2004),.clk(gclk));
	jor g1951(.dina(w_n2002_0[0]),.dinb(w_n1999_0[0]),.dout(n2005),.clk(gclk));
	jor g1952(.dina(w_n1921_0[0]),.dinb(w_n1908_0[0]),.dout(n2006),.clk(gclk));
	jand g1953(.dina(n2006),.dinb(n2005),.dout(n2007),.clk(gclk));
	jand g1954(.dina(n2007),.dinb(n2004),.dout(n2008),.clk(gclk));
	jor g1955(.dina(w_n1922_0[0]),.dinb(n2008),.dout(n2009),.clk(gclk));
	jand g1956(.dina(n2009),.dinb(w_n1846_0[0]),.dout(n2010),.clk(gclk));
	jor g1957(.dina(n2010),.dinb(w_n1844_0[0]),.dout(n2011),.clk(gclk));
	jand g1958(.dina(n2011),.dinb(w_n1840_0[0]),.dout(n2012),.clk(gclk));
	jor g1959(.dina(w_n1930_0[0]),.dinb(n2012),.dout(n2013),.clk(gclk));
	jand g1960(.dina(n2013),.dinb(n1998),.dout(n2014),.clk(gclk));
	jor g1961(.dina(w_n2014_0[1]),.dinb(w_n1767_0[1]),.dout(n2015),.clk(gclk));
	jand g1962(.dina(n2015),.dinb(w_n1759_0[0]),.dout(n2016),.clk(gclk));
	jand g1963(.dina(w_n2014_0[0]),.dinb(w_n1767_0[0]),.dout(n2017),.clk(gclk));
	jor g1964(.dina(n2017),.dinb(w_n1940_0[0]),.dout(n2018),.clk(gclk));
	jor g1965(.dina(n2018),.dinb(n2016),.dout(n2019),.clk(gclk));
	jand g1966(.dina(w_n1950_0[0]),.dinb(n2019),.dout(n2020),.clk(gclk));
	jor g1967(.dina(n2020),.dinb(w_n1710_0[0]),.dout(n2021),.clk(gclk));
	jand g1968(.dina(n2021),.dinb(n1997),.dout(n2022),.clk(gclk));
	jor g1969(.dina(n2022),.dinb(w_n1996_0[1]),.dout(n2023),.clk(gclk));
	jand g1970(.dina(w_n1615_0[0]),.dinb(w_n1601_0[0]),.dout(n2024),.clk(gclk));
	jand g1971(.dina(w_n1662_0[0]),.dinb(w_n1616_0[0]),.dout(n2025),.clk(gclk));
	jor g1972(.dina(n2025),.dinb(n2024),.dout(n2026),.clk(gclk));
	jand g1973(.dina(w_n1631_0[0]),.dinb(w_n1516_0[0]),.dout(n2027),.clk(gclk));
	jand g1974(.dina(w_n1661_0[0]),.dinb(w_n1632_0[0]),.dout(n2028),.clk(gclk));
	jor g1975(.dina(n2028),.dinb(n2027),.dout(n2029),.clk(gclk));
	jand g1976(.dina(w_n1493_4[2]),.dinb(w_n1154_7[1]),.dout(n2030),.clk(gclk));
	jnot g1977(.din(n2030),.dout(n2031),.clk(gclk));
	jxor g1978(.dina(w_n1474_6[0]),.dinb(w_n1168_2[0]),.dout(n2032),.clk(gclk));
	jor g1979(.dina(n2032),.dinb(w_n1490_4[1]),.dout(n2033),.clk(gclk));
	jand g1980(.dina(w_n1505_4[0]),.dinb(w_n1156_8[2]),.dout(n2034),.clk(gclk));
	jnot g1981(.din(n2034),.dout(n2035),.clk(gclk));
	jand g1982(.dina(n2035),.dinb(n2033),.dout(n2036),.clk(gclk));
	jand g1983(.dina(n2036),.dinb(n2031),.dout(n2037),.clk(gclk));
	jand g1984(.dina(w_n1629_0[0]),.dinb(w_n1626_0[0]),.dout(n2038),.clk(gclk));
	jand g1985(.dina(w_n1630_0[0]),.dinb(w_n1625_0[0]),.dout(n2039),.clk(gclk));
	jor g1986(.dina(n2039),.dinb(n2038),.dout(n2040),.clk(gclk));
	jxor g1987(.dina(w_n2040_0[1]),.dinb(w_n2037_0[1]),.dout(n2041),.clk(gclk));
	jand g1988(.dina(w_n1659_0[0]),.dinb(w_n1648_0[0]),.dout(n2042),.clk(gclk));
	jand g1989(.dina(w_n1660_0[0]),.dinb(w_n1640_0[0]),.dout(n2043),.clk(gclk));
	jor g1990(.dina(n2043),.dinb(n2042),.dout(n2044),.clk(gclk));
	jxor g1991(.dina(w_n2044_0[1]),.dinb(w_n2041_0[1]),.dout(n2045),.clk(gclk));
	jxor g1992(.dina(w_n2045_0[1]),.dinb(w_n2029_0[1]),.dout(n2046),.clk(gclk));
	jand g1993(.dina(w_n1613_0[0]),.dinb(w_n1605_0[0]),.dout(n2047),.clk(gclk));
	jand g1994(.dina(w_n1614_0[0]),.dinb(w_n1604_0[0]),.dout(n2048),.clk(gclk));
	jor g1995(.dina(n2048),.dinb(n2047),.dout(n2049),.clk(gclk));
	jand g1996(.dina(w_n1438_20[2]),.dinb(w_n1534_0[0]),.dout(n2050),.clk(gclk));
	jnot g1997(.din(w_n1438_20[1]),.dout(n2051),.clk(gclk));
	jand g1998(.dina(w_n2051_8[1]),.dinb(w_n1529_0[1]),.dout(n2052),.clk(gclk));
	jor g1999(.dina(n2052),.dinb(n2050),.dout(n2053),.clk(gclk));
	jnot g2000(.din(n2053),.dout(n2054),.clk(gclk));
	jand g2001(.dina(w_n1434_5[1]),.dinb(w_n1539_0[2]),.dout(n2055),.clk(gclk));
	jand g2002(.dina(w_n1622_4[0]),.dinb(w_n1542_0[2]),.dout(n2056),.clk(gclk));
	jor g2003(.dina(n2056),.dinb(n2055),.dout(n2057),.clk(gclk));
	jand g2004(.dina(n2057),.dinb(n2054),.dout(n2058),.clk(gclk));
	jand g2005(.dina(w_n1499_2[0]),.dinb(w_n1494_5[1]),.dout(n2059),.clk(gclk));
	jxor g2006(.dina(w_n2059_0[1]),.dinb(w_n716_4[0]),.dout(n2060),.clk(gclk));
	jxor g2007(.dina(w_n2060_0[1]),.dinb(w_n2058_0[1]),.dout(n2061),.clk(gclk));
	jxor g2008(.dina(w_n2061_0[1]),.dinb(w_n2049_0[1]),.dout(n2062),.clk(gclk));
	jand g2009(.dina(w_n1551_3[1]),.dinb(w_n1259_7[1]),.dout(n2063),.clk(gclk));
	jand g2010(.dina(w_n1549_3[1]),.dinb(w_n1257_10[2]),.dout(n2064),.clk(gclk));
	jor g2011(.dina(n2064),.dinb(n2063),.dout(n2065),.clk(gclk));
	jnot g2012(.din(n2065),.dout(n2066),.clk(gclk));
	jand g2013(.dina(w_n1558_3[1]),.dinb(w_n1266_3[0]),.dout(n2067),.clk(gclk));
	jand g2014(.dina(w_n1560_3[1]),.dinb(w_n1272_2[1]),.dout(n2068),.clk(gclk));
	jor g2015(.dina(n2068),.dinb(n2067),.dout(n2069),.clk(gclk));
	jand g2016(.dina(n2069),.dinb(n2066),.dout(n2070),.clk(gclk));
	jand g2017(.dina(w_n1416_1[2]),.dinb(w_n881_3[0]),.dout(n2071),.clk(gclk));
	jand g2018(.dina(w_n1418_2[0]),.dinb(w_n880_3[2]),.dout(n2072),.clk(gclk));
	jor g2019(.dina(n2072),.dinb(n2071),.dout(n2073),.clk(gclk));
	jnot g2020(.din(n2073),.dout(n2074),.clk(gclk));
	jand g2021(.dina(w_n1164_2[0]),.dinb(w_n994_4[0]),.dout(n2075),.clk(gclk));
	jand g2022(.dina(w_n1170_2[1]),.dinb(w_n996_3[1]),.dout(n2076),.clk(gclk));
	jor g2023(.dina(n2076),.dinb(n2075),.dout(n2077),.clk(gclk));
	jand g2024(.dina(n2077),.dinb(n2074),.dout(n2078),.clk(gclk));
	jand g2025(.dina(w_n1480_9[0]),.dinb(w_n1649_0[1]),.dout(n2079),.clk(gclk));
	jand g2026(.dina(w_n1356_10[1]),.dinb(w_n1651_1[0]),.dout(n2080),.clk(gclk));
	jor g2027(.dina(n2080),.dinb(n2079),.dout(n2081),.clk(gclk));
	jnot g2028(.din(n2081),.dout(n2082),.clk(gclk));
	jand g2029(.dina(w_n1360_4[1]),.dinb(w_n1254_1[0]),.dout(n2083),.clk(gclk));
	jand g2030(.dina(w_n1485_4[0]),.dinb(w_n1656_0[2]),.dout(n2084),.clk(gclk));
	jor g2031(.dina(n2084),.dinb(n2083),.dout(n2085),.clk(gclk));
	jand g2032(.dina(n2085),.dinb(n2082),.dout(n2086),.clk(gclk));
	jxor g2033(.dina(w_n2086_0[1]),.dinb(w_n2078_0[1]),.dout(n2087),.clk(gclk));
	jxor g2034(.dina(w_n2087_0[1]),.dinb(w_n2070_0[1]),.dout(n2088),.clk(gclk));
	jxor g2035(.dina(w_n2088_0[1]),.dinb(w_n2062_0[1]),.dout(n2089),.clk(gclk));
	jxor g2036(.dina(w_n2089_0[1]),.dinb(w_n2046_0[1]),.dout(n2090),.clk(gclk));
	jxor g2037(.dina(w_n2090_0[1]),.dinb(w_n2026_0[1]),.dout(n2091),.clk(gclk));
	jxor g2038(.dina(w_n2091_1[1]),.dinb(w_n2023_0[1]),.dout(n2092),.clk(gclk));
	jxor g2039(.dina(w_n2092_0[2]),.dinb(w_n1994_0[1]),.dout(n2093),.clk(gclk));
	jxor g2040(.dina(w_n2093_0[1]),.dinb(w_n1960_0[2]),.dout(n2094),.clk(gclk));
	jxor g2041(.dina(w_n2094_6[2]),.dinb(w_n1955_0[1]),.dout(n2095),.clk(gclk));
	jnot g2042(.din(w_n2095_0[1]),.dout(n2096),.clk(gclk));
	jxor g2043(.dina(w_n1259_7[0]),.dinb(w_n880_3[1]),.dout(n2097),.clk(gclk));
	jnot g2044(.din(w_n2097_0[2]),.dout(n2098),.clk(gclk));
	jxor g2045(.dina(w_n1356_10[0]),.dinb(w_n996_3[0]),.dout(n2099),.clk(gclk));
	jnot g2046(.din(w_n2099_0[1]),.dout(n2100),.clk(gclk));
	jand g2047(.dina(w_n2100_0[1]),.dinb(w_n2098_0[2]),.dout(n2101),.clk(gclk));
	jand g2048(.dina(w_n2101_1[1]),.dinb(w_n2096_1[1]),.dout(n2102),.clk(gclk));
	jand g2049(.dina(w_n2099_0[0]),.dinb(w_n2098_0[1]),.dout(n2103),.clk(gclk));
	jand g2050(.dina(w_n2103_0[2]),.dinb(w_n2094_6[1]),.dout(n2104),.clk(gclk));
	jxor g2051(.dina(w_n994_3[2]),.dinb(w_n881_2[2]),.dout(n2105),.clk(gclk));
	jnot g2052(.din(w_n2105_0[1]),.dout(n2106),.clk(gclk));
	jand g2053(.dina(n2106),.dinb(w_n2097_0[1]),.dout(n2107),.clk(gclk));
	jand g2054(.dina(w_n2107_0[2]),.dinb(w_n1956_7[0]),.dout(n2108),.clk(gclk));
	jor g2055(.dina(n2108),.dinb(n2104),.dout(n2109),.clk(gclk));
	jor g2056(.dina(n2109),.dinb(n2102),.dout(n2110),.clk(gclk));
	jnot g2057(.din(w_n2110_0[1]),.dout(n2111),.clk(gclk));
	jand g2058(.dina(w_n2098_0[0]),.dinb(w_n1956_6[2]),.dout(n2112),.clk(gclk));
	jnot g2059(.din(w_n2112_1[1]),.dout(n2113),.clk(gclk));
	jand g2060(.dina(n2113),.dinb(w_n1356_9[2]),.dout(n2114),.clk(gclk));
	jand g2061(.dina(n2114),.dinb(n2111),.dout(n2115),.clk(gclk));
	jnot g2062(.din(w_n2094_6[0]),.dout(n2116),.clk(gclk));
	jor g2063(.dina(w_n2116_2[2]),.dinb(w_n1956_6[1]),.dout(n2117),.clk(gclk));
	jnot g2064(.din(w_n1996_0[0]),.dout(n2118),.clk(gclk));
	jor g2065(.dina(w_n1953_0[0]),.dinb(w_n1664_0[0]),.dout(n2119),.clk(gclk));
	jand g2066(.dina(n2119),.dinb(n2118),.dout(n2120),.clk(gclk));
	jxor g2067(.dina(w_n2091_1[0]),.dinb(w_n2120_0[1]),.dout(n2121),.clk(gclk));
	jand g2068(.dina(n2121),.dinb(w_n1994_0[0]),.dout(n2122),.clk(gclk));
	jnot g2069(.din(w_n1960_0[1]),.dout(n2123),.clk(gclk));
	jxor g2070(.dina(w_n2092_0[1]),.dinb(w_n1993_0[1]),.dout(n2124),.clk(gclk));
	jand g2071(.dina(n2124),.dinb(n2123),.dout(n2125),.clk(gclk));
	jor g2072(.dina(n2125),.dinb(n2122),.dout(n2126),.clk(gclk));
	jand g2073(.dina(w_n852_0[2]),.dinb(w_n600_1[2]),.dout(n2127),.clk(gclk));
	jand g2074(.dina(w_n331_1[2]),.dinb(w_n204_1[1]),.dout(n2128),.clk(gclk));
	jand g2075(.dina(n2128),.dinb(w_n435_1[2]),.dout(n2129),.clk(gclk));
	jand g2076(.dina(n2129),.dinb(w_n2127_1[1]),.dout(n2130),.clk(gclk));
	jand g2077(.dina(w_n2130_0[1]),.dinb(w_n1961_0[1]),.dout(n2131),.clk(gclk));
	jand g2078(.dina(w_n395_1[1]),.dinb(w_n265_1[1]),.dout(n2132),.clk(gclk));
	jand g2079(.dina(n2132),.dinb(w_n825_1[0]),.dout(n2133),.clk(gclk));
	jand g2080(.dina(n2133),.dinb(w_n491_0[0]),.dout(n2134),.clk(gclk));
	jnot g2081(.din(w_n1180_0[0]),.dout(n2135),.clk(gclk));
	jand g2082(.dina(w_n1345_1[0]),.dinb(w_n2135_0[2]),.dout(n2136),.clk(gclk));
	jand g2083(.dina(n2136),.dinb(w_n2134_0[2]),.dout(n2137),.clk(gclk));
	jand g2084(.dina(n2137),.dinb(n2131),.dout(n2138),.clk(gclk));
	jand g2085(.dina(w_n366_1[2]),.dinb(w_n218_1[2]),.dout(n2139),.clk(gclk));
	jand g2086(.dina(n2139),.dinb(w_n411_1[1]),.dout(n2140),.clk(gclk));
	jand g2087(.dina(w_n1035_2[0]),.dinb(w_n248_2[1]),.dout(n2141),.clk(gclk));
	jand g2088(.dina(n2141),.dinb(w_n527_1[1]),.dout(n2142),.clk(gclk));
	jand g2089(.dina(w_n2142_0[2]),.dinb(w_n586_0[0]),.dout(n2143),.clk(gclk));
	jand g2090(.dina(n2143),.dinb(w_n510_2[0]),.dout(n2144),.clk(gclk));
	jand g2091(.dina(n2144),.dinb(n2140),.dout(n2145),.clk(gclk));
	jand g2092(.dina(n2145),.dinb(n2138),.dout(n2146),.clk(gclk));
	jand g2093(.dina(w_n562_0[2]),.dinb(w_n543_0[0]),.dout(n2147),.clk(gclk));
	jand g2094(.dina(w_n2147_0[1]),.dinb(w_n2146_0[2]),.dout(n2148),.clk(gclk));
	jand g2095(.dina(w_n114_1[2]),.dinb(w_n102_2[1]),.dout(n2149),.clk(gclk));
	jand g2096(.dina(w_n347_1[1]),.dinb(w_n213_2[0]),.dout(n2150),.clk(gclk));
	jand g2097(.dina(n2150),.dinb(w_n2149_0[1]),.dout(n2151),.clk(gclk));
	jand g2098(.dina(w_n439_2[2]),.dinb(w_n339_2[2]),.dout(n2152),.clk(gclk));
	jand g2099(.dina(n2152),.dinb(w_n430_0[2]),.dout(n2153),.clk(gclk));
	jand g2100(.dina(n2153),.dinb(n2151),.dout(n2154),.clk(gclk));
	jand g2101(.dina(w_n570_1[0]),.dinb(w_n897_1[2]),.dout(n2155),.clk(gclk));
	jand g2102(.dina(w_n374_1[1]),.dinb(w_n250_1[1]),.dout(n2156),.clk(gclk));
	jand g2103(.dina(n2156),.dinb(w_n2155_1[1]),.dout(n2157),.clk(gclk));
	jand g2104(.dina(w_n1459_0[1]),.dinb(w_n1072_1[0]),.dout(n2158),.clk(gclk));
	jand g2105(.dina(n2158),.dinb(n2157),.dout(n2159),.clk(gclk));
	jand g2106(.dina(n2159),.dinb(w_n2154_0[1]),.dout(n2160),.clk(gclk));
	jand g2107(.dina(w_n1095_2[0]),.dinb(w_n886_0[2]),.dout(n2161),.clk(gclk));
	jand g2108(.dina(w_n269_0[2]),.dinb(w_n195_1[0]),.dout(n2162),.clk(gclk));
	jand g2109(.dina(n2162),.dinb(n2161),.dout(n2163),.clk(gclk));
	jand g2110(.dina(n2163),.dinb(n2160),.dout(n2164),.clk(gclk));
	jand g2111(.dina(n2164),.dinb(w_n180_0[2]),.dout(n2165),.clk(gclk));
	jand g2112(.dina(n2165),.dinb(n2148),.dout(n2166),.clk(gclk));
	jand g2113(.dina(w_n2090_0[0]),.dinb(w_n2026_0[0]),.dout(n2167),.clk(gclk));
	jand g2114(.dina(w_n2091_0[2]),.dinb(w_n2023_0[0]),.dout(n2168),.clk(gclk));
	jor g2115(.dina(n2168),.dinb(w_n2167_0[1]),.dout(n2169),.clk(gclk));
	jand g2116(.dina(w_n2045_0[0]),.dinb(w_n2029_0[0]),.dout(n2170),.clk(gclk));
	jand g2117(.dina(w_n2089_0[0]),.dinb(w_n2046_0[0]),.dout(n2171),.clk(gclk));
	jor g2118(.dina(n2171),.dinb(n2170),.dout(n2172),.clk(gclk));
	jand g2119(.dina(w_n2061_0[0]),.dinb(w_n2049_0[0]),.dout(n2173),.clk(gclk));
	jand g2120(.dina(w_n2088_0[0]),.dinb(w_n2062_0[0]),.dout(n2174),.clk(gclk));
	jor g2121(.dina(n2174),.dinb(n2173),.dout(n2175),.clk(gclk));
	jand g2122(.dina(w_n1505_3[2]),.dinb(w_n1168_1[2]),.dout(n2176),.clk(gclk));
	jnot g2123(.din(n2176),.dout(n2177),.clk(gclk));
	jxor g2124(.dina(w_n1474_5[2]),.dinb(w_n1272_2[0]),.dout(n2178),.clk(gclk));
	jor g2125(.dina(n2178),.dinb(w_n1490_4[0]),.dout(n2179),.clk(gclk));
	jand g2126(.dina(w_n1493_4[1]),.dinb(w_n1166_2[2]),.dout(n2180),.clk(gclk));
	jnot g2127(.din(n2180),.dout(n2181),.clk(gclk));
	jand g2128(.dina(n2181),.dinb(n2179),.dout(n2182),.clk(gclk));
	jand g2129(.dina(n2182),.dinb(n2177),.dout(n2183),.clk(gclk));
	jand g2130(.dina(w_n2059_0[0]),.dinb(w_n716_3[2]),.dout(n2184),.clk(gclk));
	jand g2131(.dina(w_n2060_0[0]),.dinb(w_n2058_0[0]),.dout(n2185),.clk(gclk));
	jor g2132(.dina(n2185),.dinb(n2184),.dout(n2186),.clk(gclk));
	jxor g2133(.dina(w_n2186_0[1]),.dinb(w_n2183_0[1]),.dout(n2187),.clk(gclk));
	jand g2134(.dina(w_n2086_0[0]),.dinb(w_n2078_0[0]),.dout(n2188),.clk(gclk));
	jand g2135(.dina(w_n2087_0[0]),.dinb(w_n2070_0[0]),.dout(n2189),.clk(gclk));
	jor g2136(.dina(n2189),.dinb(n2188),.dout(n2190),.clk(gclk));
	jxor g2137(.dina(w_n2190_0[1]),.dinb(w_n2187_0[1]),.dout(n2191),.clk(gclk));
	jxor g2138(.dina(w_n2191_0[1]),.dinb(w_n2175_0[1]),.dout(n2192),.clk(gclk));
	jand g2139(.dina(w_n2040_0[0]),.dinb(w_n2037_0[0]),.dout(n2193),.clk(gclk));
	jand g2140(.dina(w_n2044_0[0]),.dinb(w_n2041_0[0]),.dout(n2194),.clk(gclk));
	jor g2141(.dina(n2194),.dinb(n2193),.dout(n2195),.clk(gclk));
	jand g2142(.dina(w_n1551_3[0]),.dinb(w_n881_2[1]),.dout(n2196),.clk(gclk));
	jand g2143(.dina(w_n1549_3[0]),.dinb(w_n880_3[0]),.dout(n2197),.clk(gclk));
	jor g2144(.dina(n2197),.dinb(n2196),.dout(n2198),.clk(gclk));
	jnot g2145(.din(n2198),.dout(n2199),.clk(gclk));
	jand g2146(.dina(w_n1558_3[0]),.dinb(w_n1257_10[1]),.dout(n2200),.clk(gclk));
	jand g2147(.dina(w_n1560_3[0]),.dinb(w_n1259_6[2]),.dout(n2201),.clk(gclk));
	jor g2148(.dina(n2201),.dinb(n2200),.dout(n2202),.clk(gclk));
	jand g2149(.dina(n2202),.dinb(n2199),.dout(n2203),.clk(gclk));
	jand g2150(.dina(w_n1434_5[0]),.dinb(w_n1255_0[2]),.dout(n2204),.clk(gclk));
	jand g2151(.dina(w_n1622_3[2]),.dinb(w_n1261_0[2]),.dout(n2205),.clk(gclk));
	jor g2152(.dina(n2205),.dinb(n2204),.dout(n2206),.clk(gclk));
	jnot g2153(.din(n2206),.dout(n2207),.clk(gclk));
	jand g2154(.dina(w_n1360_4[0]),.dinb(w_n1270_1[0]),.dout(n2208),.clk(gclk));
	jand g2155(.dina(w_n1485_3[2]),.dinb(w_n1295_1[0]),.dout(n2209),.clk(gclk));
	jor g2156(.dina(n2209),.dinb(n2208),.dout(n2210),.clk(gclk));
	jand g2157(.dina(n2210),.dinb(n2207),.dout(n2211),.clk(gclk));
	jand g2158(.dina(w_n1416_1[1]),.dinb(w_n996_2[2]),.dout(n2212),.clk(gclk));
	jand g2159(.dina(w_n1418_1[2]),.dinb(w_n994_3[1]),.dout(n2213),.clk(gclk));
	jor g2160(.dina(n2213),.dinb(n2212),.dout(n2214),.clk(gclk));
	jnot g2161(.din(n2214),.dout(n2215),.clk(gclk));
	jand g2162(.dina(w_n1356_9[1]),.dinb(w_n1164_1[2]),.dout(n2216),.clk(gclk));
	jand g2163(.dina(w_n1480_8[2]),.dinb(w_n1170_2[0]),.dout(n2217),.clk(gclk));
	jor g2164(.dina(n2217),.dinb(n2216),.dout(n2218),.clk(gclk));
	jand g2165(.dina(n2218),.dinb(n2215),.dout(n2219),.clk(gclk));
	jxor g2166(.dina(w_n2219_0[1]),.dinb(w_n2211_0[1]),.dout(n2220),.clk(gclk));
	jxor g2167(.dina(w_n2220_0[1]),.dinb(w_n2203_0[1]),.dout(n2221),.clk(gclk));
	jand g2168(.dina(w_n2051_8[0]),.dinb(w_n815_0[1]),.dout(n2222),.clk(gclk));
	jand g2169(.dina(w_n1438_20[0]),.dinb(w_n989_0[2]),.dout(n2223),.clk(gclk));
	jor g2170(.dina(n2223),.dinb(w_n1529_0[0]),.dout(n2224),.clk(gclk));
	jor g2171(.dina(n2224),.dinb(n2222),.dout(n2225),.clk(gclk));
	jnot g2172(.din(n2225),.dout(n2226),.clk(gclk));
	jand g2173(.dina(w_n1494_5[0]),.dinb(w_n1154_7[0]),.dout(n2227),.clk(gclk));
	jxor g2174(.dina(w_n2227_0[1]),.dinb(w_n716_3[1]),.dout(n2228),.clk(gclk));
	jxor g2175(.dina(w_n2228_0[1]),.dinb(w_n2226_0[1]),.dout(n2229),.clk(gclk));
	jxor g2176(.dina(w_n2229_0[1]),.dinb(w_n2221_0[1]),.dout(n2230),.clk(gclk));
	jxor g2177(.dina(w_n2230_0[1]),.dinb(w_n2195_0[1]),.dout(n2231),.clk(gclk));
	jxor g2178(.dina(w_n2231_0[1]),.dinb(w_n2192_0[1]),.dout(n2232),.clk(gclk));
	jxor g2179(.dina(w_n2232_0[1]),.dinb(w_n2172_0[1]),.dout(n2233),.clk(gclk));
	jxor g2180(.dina(w_n2233_1[1]),.dinb(w_n2169_0[1]),.dout(n2234),.clk(gclk));
	jxor g2181(.dina(w_n2234_0[2]),.dinb(w_n2166_0[2]),.dout(n2235),.clk(gclk));
	jxor g2182(.dina(w_n2235_0[2]),.dinb(w_n2126_0[1]),.dout(n2236),.clk(gclk));
	jxor g2183(.dina(w_n2236_5[1]),.dinb(n2117),.dout(n2237),.clk(gclk));
	jnot g2184(.din(n2237),.dout(n2238),.clk(gclk));
	jand g2185(.dina(w_n2238_1[1]),.dinb(w_n2101_1[0]),.dout(n2239),.clk(gclk));
	jand g2186(.dina(w_n2107_0[1]),.dinb(w_n2094_5[2]),.dout(n2240),.clk(gclk));
	jand g2187(.dina(w_n2236_5[0]),.dinb(w_n2103_0[1]),.dout(n2241),.clk(gclk));
	jor g2188(.dina(n2241),.dinb(n2240),.dout(n2242),.clk(gclk));
	jand g2189(.dina(w_n2105_0[0]),.dinb(w_n2097_0[0]),.dout(n2243),.clk(gclk));
	jand g2190(.dina(n2243),.dinb(w_n2100_0[0]),.dout(n2244),.clk(gclk));
	jand g2191(.dina(w_n2244_0[2]),.dinb(w_n1956_6[0]),.dout(n2245),.clk(gclk));
	jor g2192(.dina(n2245),.dinb(n2242),.dout(n2246),.clk(gclk));
	jor g2193(.dina(n2246),.dinb(n2239),.dout(n2247),.clk(gclk));
	jnot g2194(.din(n2247),.dout(n2248),.clk(gclk));
	jand g2195(.dina(w_n2248_0[1]),.dinb(w_n2115_0[1]),.dout(n2249),.clk(gclk));
	jand g2196(.dina(w_n2249_0[1]),.dinb(w_n1959_0[2]),.dout(n2250),.clk(gclk));
	jxor g2197(.dina(w_n2249_0[0]),.dinb(w_n1959_0[1]),.dout(n2251),.clk(gclk));
	jnot g2198(.din(w_n2101_0[2]),.dout(n2252),.clk(gclk));
	jor g2199(.dina(w_n2092_0[0]),.dinb(w_n1993_0[0]),.dout(n2253),.clk(gclk));
	jor g2200(.dina(w_n2093_0[0]),.dinb(w_n1960_0[0]),.dout(n2254),.clk(gclk));
	jand g2201(.dina(n2254),.dinb(n2253),.dout(n2255),.clk(gclk));
	jxor g2202(.dina(w_n2235_0[1]),.dinb(w_n2255_0[1]),.dout(n2256),.clk(gclk));
	jand g2203(.dina(w_n2256_5[2]),.dinb(w_n1955_0[0]),.dout(n2257),.clk(gclk));
	jor g2204(.dina(n2257),.dinb(w_n2116_2[1]),.dout(n2258),.clk(gclk));
	jor g2205(.dina(w_n2234_0[1]),.dinb(w_n2166_0[1]),.dout(n2259),.clk(gclk));
	jnot g2206(.din(w_n2166_0[0]),.dout(n2260),.clk(gclk));
	jxor g2207(.dina(w_n2234_0[0]),.dinb(w_n2260_0[1]),.dout(n2261),.clk(gclk));
	jor g2208(.dina(n2261),.dinb(w_n2255_0[0]),.dout(n2262),.clk(gclk));
	jand g2209(.dina(n2262),.dinb(n2259),.dout(n2263),.clk(gclk));
	jand g2210(.dina(w_n1127_0[1]),.dinb(w_n129_0[2]),.dout(n2264),.clk(gclk));
	jand g2211(.dina(n2264),.dinb(w_n445_1[0]),.dout(n2265),.clk(gclk));
	jand g2212(.dina(n2265),.dinb(w_n222_2[0]),.dout(n2266),.clk(gclk));
	jand g2213(.dina(n2266),.dinb(w_n2154_0[0]),.dout(n2267),.clk(gclk));
	jand g2214(.dina(n2267),.dinb(w_n1016_0[2]),.dout(n2268),.clk(gclk));
	jand g2215(.dina(w_n434_1[2]),.dinb(w_n221_2[0]),.dout(n2269),.clk(gclk));
	jand g2216(.dina(n2269),.dinb(w_n244_2[0]),.dout(n2270),.clk(gclk));
	jand g2217(.dina(w_n337_1[2]),.dinb(w_n232_3[0]),.dout(n2271),.clk(gclk));
	jand g2218(.dina(w_n717_2[1]),.dinb(w_n197_1[2]),.dout(n2272),.clk(gclk));
	jand g2219(.dina(n2272),.dinb(n2271),.dout(n2273),.clk(gclk));
	jand g2220(.dina(n2273),.dinb(w_n329_0[2]),.dout(n2274),.clk(gclk));
	jand g2221(.dina(n2274),.dinb(w_n394_0[0]),.dout(n2275),.clk(gclk));
	jand g2222(.dina(n2275),.dinb(n2270),.dout(n2276),.clk(gclk));
	jand g2223(.dina(n2276),.dinb(n2268),.dout(n2277),.clk(gclk));
	jand g2224(.dina(w_n2232_0[0]),.dinb(w_n2172_0[0]),.dout(n2278),.clk(gclk));
	jand g2225(.dina(w_n2233_1[0]),.dinb(w_n2169_0[0]),.dout(n2279),.clk(gclk));
	jor g2226(.dina(n2279),.dinb(w_n2278_0[1]),.dout(n2280),.clk(gclk));
	jand g2227(.dina(w_n2191_0[0]),.dinb(w_n2175_0[0]),.dout(n2281),.clk(gclk));
	jand g2228(.dina(w_n2231_0[0]),.dinb(w_n2192_0[0]),.dout(n2282),.clk(gclk));
	jor g2229(.dina(n2282),.dinb(n2281),.dout(n2283),.clk(gclk));
	jand g2230(.dina(w_n2229_0[0]),.dinb(w_n2221_0[0]),.dout(n2284),.clk(gclk));
	jand g2231(.dina(w_n2230_0[0]),.dinb(w_n2195_0[0]),.dout(n2285),.clk(gclk));
	jor g2232(.dina(n2285),.dinb(n2284),.dout(n2286),.clk(gclk));
	jand g2233(.dina(w_n2227_0[0]),.dinb(w_n716_3[0]),.dout(n2287),.clk(gclk));
	jand g2234(.dina(w_n2228_0[0]),.dinb(w_n2226_0[0]),.dout(n2288),.clk(gclk));
	jor g2235(.dina(n2288),.dinb(n2287),.dout(n2289),.clk(gclk));
	jand g2236(.dina(w_n1485_3[1]),.dinb(w_n1576_0[1]),.dout(n2290),.clk(gclk));
	jand g2237(.dina(w_n1360_3[2]),.dinb(w_n1163_0[0]),.dout(n2291),.clk(gclk));
	jor g2238(.dina(n2291),.dinb(n2290),.dout(n2292),.clk(gclk));
	jnot g2239(.din(n2292),.dout(n2293),.clk(gclk));
	jand g2240(.dina(w_n1356_9[0]),.dinb(w_n1160_0[2]),.dout(n2294),.clk(gclk));
	jand g2241(.dina(w_n1480_8[1]),.dinb(w_n1152_0[2]),.dout(n2295),.clk(gclk));
	jor g2242(.dina(n2295),.dinb(n2294),.dout(n2296),.clk(gclk));
	jand g2243(.dina(n2296),.dinb(n2293),.dout(n2297),.clk(gclk));
	jand g2244(.dina(w_n1532_0[0]),.dinb(w_n716_2[2]),.dout(n2298),.clk(gclk));
	jnot g2245(.din(n2298),.dout(n2299),.clk(gclk));
	jand g2246(.dina(w_n930_0[2]),.dinb(w_n607_0[2]),.dout(n2300),.clk(gclk));
	jnot g2247(.din(n2300),.dout(n2301),.clk(gclk));
	jand g2248(.dina(w_n1494_4[2]),.dinb(w_n1166_2[1]),.dout(n2302),.clk(gclk));
	jand g2249(.dina(w_n2301_0[1]),.dinb(w_n2302_0[1]),.dout(n2303),.clk(gclk));
	jand g2250(.dina(n2303),.dinb(w_n2299_0[1]),.dout(n2304),.clk(gclk));
	jnot g2251(.din(n2304),.dout(n2305),.clk(gclk));
	jand g2252(.dina(w_n2305_0[1]),.dinb(w_n2301_0[0]),.dout(n2306),.clk(gclk));
	jand g2253(.dina(w_n2306_0[1]),.dinb(w_n2299_0[0]),.dout(n2307),.clk(gclk));
	jand g2254(.dina(w_n2305_0[0]),.dinb(w_n2302_0[0]),.dout(n2308),.clk(gclk));
	jor g2255(.dina(n2308),.dinb(n2307),.dout(n2309),.clk(gclk));
	jxor g2256(.dina(w_n2309_0[1]),.dinb(w_n2297_0[1]),.dout(n2310),.clk(gclk));
	jxor g2257(.dina(w_n2310_0[1]),.dinb(w_n2289_0[1]),.dout(n2311),.clk(gclk));
	jxor g2258(.dina(w_n2311_0[1]),.dinb(w_n2286_0[1]),.dout(n2312),.clk(gclk));
	jand g2259(.dina(w_n2186_0[0]),.dinb(w_n2183_0[0]),.dout(n2313),.clk(gclk));
	jand g2260(.dina(w_n2190_0[0]),.dinb(w_n2187_0[0]),.dout(n2314),.clk(gclk));
	jor g2261(.dina(n2314),.dinb(n2313),.dout(n2315),.clk(gclk));
	jand g2262(.dina(w_n2219_0[0]),.dinb(w_n2211_0[0]),.dout(n2316),.clk(gclk));
	jand g2263(.dina(w_n2220_0[0]),.dinb(w_n2203_0[0]),.dout(n2317),.clk(gclk));
	jor g2264(.dina(n2317),.dinb(n2316),.dout(n2318),.clk(gclk));
	jand g2265(.dina(w_n1622_3[1]),.dinb(w_n1649_0[0]),.dout(n2319),.clk(gclk));
	jand g2266(.dina(w_n1434_4[2]),.dinb(w_n1651_0[2]),.dout(n2320),.clk(gclk));
	jor g2267(.dina(n2320),.dinb(n2319),.dout(n2321),.clk(gclk));
	jnot g2268(.din(n2321),.dout(n2322),.clk(gclk));
	jand g2269(.dina(w_n2051_7[2]),.dinb(w_n1656_0[1]),.dout(n2323),.clk(gclk));
	jand g2270(.dina(w_n1438_19[2]),.dinb(w_n1254_0[2]),.dout(n2324),.clk(gclk));
	jor g2271(.dina(n2324),.dinb(n2323),.dout(n2325),.clk(gclk));
	jand g2272(.dina(n2325),.dinb(n2322),.dout(n2326),.clk(gclk));
	jand g2273(.dina(w_n1551_2[2]),.dinb(w_n996_2[1]),.dout(n2327),.clk(gclk));
	jand g2274(.dina(w_n1549_2[2]),.dinb(w_n994_3[0]),.dout(n2328),.clk(gclk));
	jor g2275(.dina(n2328),.dinb(n2327),.dout(n2329),.clk(gclk));
	jnot g2276(.din(n2329),.dout(n2330),.clk(gclk));
	jand g2277(.dina(w_n1558_2[2]),.dinb(w_n880_2[2]),.dout(n2331),.clk(gclk));
	jand g2278(.dina(w_n1560_2[2]),.dinb(w_n881_2[0]),.dout(n2332),.clk(gclk));
	jor g2279(.dina(n2332),.dinb(n2331),.dout(n2333),.clk(gclk));
	jand g2280(.dina(n2333),.dinb(n2330),.dout(n2334),.clk(gclk));
	jand g2281(.dina(w_n1505_3[1]),.dinb(w_n1272_1[2]),.dout(n2335),.clk(gclk));
	jnot g2282(.din(n2335),.dout(n2336),.clk(gclk));
	jxor g2283(.dina(w_n1474_5[1]),.dinb(w_n1259_6[1]),.dout(n2337),.clk(gclk));
	jor g2284(.dina(n2337),.dinb(w_n1490_3[2]),.dout(n2338),.clk(gclk));
	jand g2285(.dina(w_n1493_4[0]),.dinb(w_n1266_2[2]),.dout(n2339),.clk(gclk));
	jnot g2286(.din(n2339),.dout(n2340),.clk(gclk));
	jand g2287(.dina(n2340),.dinb(n2338),.dout(n2341),.clk(gclk));
	jand g2288(.dina(n2341),.dinb(n2336),.dout(n2342),.clk(gclk));
	jxor g2289(.dina(w_n2342_0[1]),.dinb(w_n2334_0[1]),.dout(n2343),.clk(gclk));
	jxor g2290(.dina(w_n2343_0[1]),.dinb(w_n2326_0[1]),.dout(n2344),.clk(gclk));
	jxor g2291(.dina(w_n2344_0[1]),.dinb(w_n2318_0[1]),.dout(n2345),.clk(gclk));
	jxor g2292(.dina(w_n2345_0[1]),.dinb(w_n2315_0[1]),.dout(n2346),.clk(gclk));
	jxor g2293(.dina(w_n2346_0[1]),.dinb(w_n2312_0[1]),.dout(n2347),.clk(gclk));
	jxor g2294(.dina(w_n2347_0[1]),.dinb(w_n2283_0[1]),.dout(n2348),.clk(gclk));
	jxor g2295(.dina(w_n2348_1[1]),.dinb(w_n2280_0[1]),.dout(n2349),.clk(gclk));
	jxor g2296(.dina(w_n2349_0[2]),.dinb(w_n2277_0[2]),.dout(n2350),.clk(gclk));
	jxor g2297(.dina(w_n2350_0[2]),.dinb(w_n2263_0[1]),.dout(n2351),.clk(gclk));
	jxor g2298(.dina(w_n2351_8[1]),.dinb(w_n2256_5[1]),.dout(n2352),.clk(gclk));
	jxor g2299(.dina(w_n2352_0[2]),.dinb(w_n2258_0[1]),.dout(n2353),.clk(gclk));
	jor g2300(.dina(w_n2353_1[2]),.dinb(w_n2252_7[2]),.dout(n2354),.clk(gclk));
	jnot g2301(.din(w_n2103_0[0]),.dout(n2355),.clk(gclk));
	jor g2302(.dina(w_n2351_8[0]),.dinb(w_n2355_7[1]),.dout(n2356),.clk(gclk));
	jnot g2303(.din(w_n2244_0[1]),.dout(n2357),.clk(gclk));
	jor g2304(.dina(w_n2357_7[2]),.dinb(w_n2116_2[0]),.dout(n2358),.clk(gclk));
	jnot g2305(.din(w_n2107_0[0]),.dout(n2359),.clk(gclk));
	jor g2306(.dina(w_n2256_5[0]),.dinb(w_n2359_7[2]),.dout(n2360),.clk(gclk));
	jand g2307(.dina(n2360),.dinb(n2358),.dout(n2361),.clk(gclk));
	jand g2308(.dina(n2361),.dinb(n2356),.dout(n2362),.clk(gclk));
	jand g2309(.dina(n2362),.dinb(n2354),.dout(n2363),.clk(gclk));
	jxor g2310(.dina(n2363),.dinb(w_n1480_8[0]),.dout(n2364),.clk(gclk));
	jand g2311(.dina(w_n2364_0[1]),.dinb(w_n2251_0[1]),.dout(n2365),.clk(gclk));
	jor g2312(.dina(n2365),.dinb(n2250),.dout(n2366),.clk(gclk));
	jor g2313(.dina(w_n2351_7[2]),.dinb(w_n2256_4[2]),.dout(n2367),.clk(gclk));
	jxor g2314(.dina(w_n2351_7[1]),.dinb(w_n2236_4[2]),.dout(n2368),.clk(gclk));
	jor g2315(.dina(n2368),.dinb(w_n2258_0[0]),.dout(n2369),.clk(gclk));
	jand g2316(.dina(n2369),.dinb(n2367),.dout(n2370),.clk(gclk));
	jor g2317(.dina(w_n2349_0[1]),.dinb(w_n2277_0[1]),.dout(n2371),.clk(gclk));
	jnot g2318(.din(w_n2277_0[0]),.dout(n2372),.clk(gclk));
	jxor g2319(.dina(w_n2349_0[0]),.dinb(w_n2372_0[1]),.dout(n2373),.clk(gclk));
	jor g2320(.dina(n2373),.dinb(w_n2263_0[0]),.dout(n2374),.clk(gclk));
	jand g2321(.dina(n2374),.dinb(n2371),.dout(n2375),.clk(gclk));
	jand g2322(.dina(w_n439_2[1]),.dinb(w_n427_1[2]),.dout(n2376),.clk(gclk));
	jand g2323(.dina(n2376),.dinb(w_n1096_0[1]),.dout(n2377),.clk(gclk));
	jand g2324(.dina(w_n2377_0[1]),.dinb(w_n283_1[1]),.dout(n2378),.clk(gclk));
	jand g2325(.dina(n2378),.dinb(w_n866_0[0]),.dout(n2379),.clk(gclk));
	jand g2326(.dina(w_n160_1[0]),.dinb(w_n124_2[0]),.dout(n2380),.clk(gclk));
	jand g2327(.dina(n2380),.dinb(w_n1345_0[2]),.dout(n2381),.clk(gclk));
	jand g2328(.dina(n2381),.dinb(w_n218_1[1]),.dout(n2382),.clk(gclk));
	jand g2329(.dina(n2382),.dinb(w_n1135_1[0]),.dout(n2383),.clk(gclk));
	jand g2330(.dina(n2383),.dinb(n2379),.dout(n2384),.clk(gclk));
	jand g2331(.dina(w_n2384_0[1]),.dinb(w_n137_2[0]),.dout(n2385),.clk(gclk));
	jand g2332(.dina(n2385),.dinb(w_n404_0[2]),.dout(n2386),.clk(gclk));
	jand g2333(.dina(w_n340_1[0]),.dinb(w_n457_0[0]),.dout(n2387),.clk(gclk));
	jand g2334(.dina(n2387),.dinb(w_n411_1[0]),.dout(n2388),.clk(gclk));
	jand g2335(.dina(w_n467_1[0]),.dinb(w_n235_1[1]),.dout(n2389),.clk(gclk));
	jand g2336(.dina(n2389),.dinb(w_n309_1[1]),.dout(n2390),.clk(gclk));
	jand g2337(.dina(n2390),.dinb(w_n294_1[1]),.dout(n2391),.clk(gclk));
	jand g2338(.dina(n2391),.dinb(n2388),.dout(n2392),.clk(gclk));
	jand g2339(.dina(w_n337_1[1]),.dinb(w_n102_2[0]),.dout(n2393),.clk(gclk));
	jand g2340(.dina(n2393),.dinb(w_n327_0[1]),.dout(n2394),.clk(gclk));
	jand g2341(.dina(w_n300_2[1]),.dinb(w_n248_2[0]),.dout(n2395),.clk(gclk));
	jand g2342(.dina(w_n2395_0[2]),.dinb(w_n409_0[2]),.dout(n2396),.clk(gclk));
	jand g2343(.dina(n2396),.dinb(w_n2394_0[1]),.dout(n2397),.clk(gclk));
	jand g2344(.dina(w_n587_2[1]),.dinb(w_n305_1[0]),.dout(n2398),.clk(gclk));
	jand g2345(.dina(n2398),.dinb(w_n1057_0[0]),.dout(n2399),.clk(gclk));
	jand g2346(.dina(n2399),.dinb(w_n315_1[1]),.dout(n2400),.clk(gclk));
	jand g2347(.dina(n2400),.dinb(w_n530_0[0]),.dout(n2401),.clk(gclk));
	jand g2348(.dina(n2401),.dinb(n2397),.dout(n2402),.clk(gclk));
	jand g2349(.dina(w_n2402_0[1]),.dinb(w_n370_1[2]),.dout(n2403),.clk(gclk));
	jand g2350(.dina(w_n534_1[1]),.dinb(w_n245_0[2]),.dout(n2404),.clk(gclk));
	jand g2351(.dina(w_n600_1[1]),.dinb(w_n384_2[0]),.dout(n2405),.clk(gclk));
	jand g2352(.dina(n2405),.dinb(n2404),.dout(n2406),.clk(gclk));
	jand g2353(.dina(w_n361_1[2]),.dinb(w_n213_1[2]),.dout(n2407),.clk(gclk));
	jand g2354(.dina(n2407),.dinb(w_n170_1[1]),.dout(n2408),.clk(gclk));
	jand g2355(.dina(n2408),.dinb(n2406),.dout(n2409),.clk(gclk));
	jand g2356(.dina(w_n2409_0[1]),.dinb(n2403),.dout(n2410),.clk(gclk));
	jand g2357(.dina(n2410),.dinb(n2392),.dout(n2411),.clk(gclk));
	jand g2358(.dina(n2411),.dinb(w_n2386_0[1]),.dout(n2412),.clk(gclk));
	jand g2359(.dina(w_n2347_0[0]),.dinb(w_n2283_0[0]),.dout(n2413),.clk(gclk));
	jand g2360(.dina(w_n2348_1[0]),.dinb(w_n2280_0[0]),.dout(n2414),.clk(gclk));
	jor g2361(.dina(n2414),.dinb(w_n2413_0[1]),.dout(n2415),.clk(gclk));
	jand g2362(.dina(w_n2311_0[0]),.dinb(w_n2286_0[0]),.dout(n2416),.clk(gclk));
	jand g2363(.dina(w_n2346_0[0]),.dinb(w_n2312_0[0]),.dout(n2417),.clk(gclk));
	jor g2364(.dina(n2417),.dinb(n2416),.dout(n2418),.clk(gclk));
	jand g2365(.dina(w_n2309_0[0]),.dinb(w_n2297_0[0]),.dout(n2419),.clk(gclk));
	jand g2366(.dina(w_n2310_0[0]),.dinb(w_n2289_0[0]),.dout(n2420),.clk(gclk));
	jor g2367(.dina(n2420),.dinb(n2419),.dout(n2421),.clk(gclk));
	jand g2368(.dina(w_n2344_0[0]),.dinb(w_n2318_0[0]),.dout(n2422),.clk(gclk));
	jand g2369(.dina(w_n2345_0[0]),.dinb(w_n2315_0[0]),.dout(n2423),.clk(gclk));
	jor g2370(.dina(n2423),.dinb(n2422),.dout(n2424),.clk(gclk));
	jxor g2371(.dina(w_n2424_0[1]),.dinb(w_n2421_0[1]),.dout(n2425),.clk(gclk));
	jnot g2372(.din(w_n2306_0[0]),.dout(n2426),.clk(gclk));
	jand g2373(.dina(w_n1551_2[1]),.dinb(w_n1480_7[2]),.dout(n2427),.clk(gclk));
	jand g2374(.dina(w_n1549_2[1]),.dinb(w_n1356_8[2]),.dout(n2428),.clk(gclk));
	jor g2375(.dina(n2428),.dinb(n2427),.dout(n2429),.clk(gclk));
	jnot g2376(.din(n2429),.dout(n2430),.clk(gclk));
	jand g2377(.dina(w_n1558_2[1]),.dinb(w_n994_2[2]),.dout(n2431),.clk(gclk));
	jand g2378(.dina(w_n1560_2[1]),.dinb(w_n996_2[0]),.dout(n2432),.clk(gclk));
	jor g2379(.dina(n2432),.dinb(n2431),.dout(n2433),.clk(gclk));
	jand g2380(.dina(n2433),.dinb(n2430),.dout(n2434),.clk(gclk));
	jand g2381(.dina(w_n1493_3[2]),.dinb(w_n1257_10[0]),.dout(n2435),.clk(gclk));
	jnot g2382(.din(n2435),.dout(n2436),.clk(gclk));
	jxor g2383(.dina(w_n1474_5[0]),.dinb(w_n881_1[2]),.dout(n2437),.clk(gclk));
	jor g2384(.dina(n2437),.dinb(w_n1490_3[1]),.dout(n2438),.clk(gclk));
	jand g2385(.dina(w_n1505_3[0]),.dinb(w_n1259_6[0]),.dout(n2439),.clk(gclk));
	jnot g2386(.din(n2439),.dout(n2440),.clk(gclk));
	jand g2387(.dina(n2440),.dinb(n2438),.dout(n2441),.clk(gclk));
	jand g2388(.dina(n2441),.dinb(n2436),.dout(n2442),.clk(gclk));
	jxor g2389(.dina(w_n2442_0[1]),.dinb(w_n2434_0[1]),.dout(n2443),.clk(gclk));
	jxor g2390(.dina(w_n2443_0[1]),.dinb(w_n2426_0[1]),.dout(n2444),.clk(gclk));
	jand g2391(.dina(w_n2342_0[0]),.dinb(w_n2334_0[0]),.dout(n2445),.clk(gclk));
	jand g2392(.dina(w_n2343_0[0]),.dinb(w_n2326_0[0]),.dout(n2446),.clk(gclk));
	jor g2393(.dina(n2446),.dinb(n2445),.dout(n2447),.clk(gclk));
	jand g2394(.dina(w_n1485_3[0]),.dinb(w_n1416_1[0]),.dout(n2448),.clk(gclk));
	jand g2395(.dina(w_n1360_3[1]),.dinb(w_n1418_1[1]),.dout(n2449),.clk(gclk));
	jor g2396(.dina(n2449),.dinb(n2448),.dout(n2450),.clk(gclk));
	jnot g2397(.din(n2450),.dout(n2451),.clk(gclk));
	jand g2398(.dina(w_n1434_4[1]),.dinb(w_n1164_1[1]),.dout(n2452),.clk(gclk));
	jand g2399(.dina(w_n1622_3[0]),.dinb(w_n1170_1[2]),.dout(n2453),.clk(gclk));
	jor g2400(.dina(n2453),.dinb(n2452),.dout(n2454),.clk(gclk));
	jand g2401(.dina(n2454),.dinb(n2451),.dout(n2455),.clk(gclk));
	jand g2402(.dina(w_n1494_4[1]),.dinb(w_n1266_2[1]),.dout(n2456),.clk(gclk));
	jnot g2403(.din(w_n2456_0[2]),.dout(n2457),.clk(gclk));
	jand g2404(.dina(w_n1438_19[1]),.dinb(w_n1651_0[1]),.dout(n2458),.clk(gclk));
	jnot g2405(.din(n2458),.dout(n2459),.clk(gclk));
	jand g2406(.dina(w_n1438_19[0]),.dinb(w_n1812_0[0]),.dout(n2460),.clk(gclk));
	jor g2407(.dina(n2460),.dinb(w_n1294_0[0]),.dout(n2461),.clk(gclk));
	jand g2408(.dina(n2461),.dinb(n2459),.dout(n2462),.clk(gclk));
	jxor g2409(.dina(w_n2462_0[1]),.dinb(w_n2457_0[1]),.dout(n2463),.clk(gclk));
	jxor g2410(.dina(w_n2463_0[1]),.dinb(w_n2455_0[1]),.dout(n2464),.clk(gclk));
	jxor g2411(.dina(w_n2464_0[1]),.dinb(w_n2447_0[1]),.dout(n2465),.clk(gclk));
	jxor g2412(.dina(w_n2465_0[1]),.dinb(w_n2444_0[1]),.dout(n2466),.clk(gclk));
	jxor g2413(.dina(w_n2466_0[1]),.dinb(w_n2425_0[1]),.dout(n2467),.clk(gclk));
	jxor g2414(.dina(w_n2467_0[1]),.dinb(w_n2418_0[1]),.dout(n2468),.clk(gclk));
	jxor g2415(.dina(w_n2468_1[1]),.dinb(w_n2415_0[1]),.dout(n2469),.clk(gclk));
	jxor g2416(.dina(w_n2469_0[2]),.dinb(w_n2412_0[2]),.dout(n2470),.clk(gclk));
	jxor g2417(.dina(w_n2470_0[2]),.dinb(w_n2375_0[1]),.dout(n2471),.clk(gclk));
	jxor g2418(.dina(w_n2471_7[1]),.dinb(w_n2351_7[0]),.dout(n2472),.clk(gclk));
	jxor g2419(.dina(w_n2472_0[2]),.dinb(w_n2370_0[1]),.dout(n2473),.clk(gclk));
	jor g2420(.dina(w_n2473_1[1]),.dinb(w_n2252_7[1]),.dout(n2474),.clk(gclk));
	jor g2421(.dina(w_n2351_6[2]),.dinb(w_n2359_7[1]),.dout(n2475),.clk(gclk));
	jor g2422(.dina(w_n2471_7[0]),.dinb(w_n2355_7[0]),.dout(n2476),.clk(gclk));
	jand g2423(.dina(n2476),.dinb(n2475),.dout(n2477),.clk(gclk));
	jor g2424(.dina(w_n2357_7[1]),.dinb(w_n2256_4[1]),.dout(n2478),.clk(gclk));
	jand g2425(.dina(n2478),.dinb(n2477),.dout(n2479),.clk(gclk));
	jand g2426(.dina(n2479),.dinb(n2474),.dout(n2480),.clk(gclk));
	jxor g2427(.dina(n2480),.dinb(w_n1356_8[1]),.dout(n2481),.clk(gclk));
	jnot g2428(.din(n2481),.dout(n2482),.clk(gclk));
	jxor g2429(.dina(w_n1438_18[2]),.dinb(w_n1434_4[0]),.dout(n2483),.clk(gclk));
	jand g2430(.dina(w_n2483_1[1]),.dinb(w_n1958_1[0]),.dout(n2484),.clk(gclk));
	jand g2431(.dina(w_n2484_1[2]),.dinb(w_n2096_1[0]),.dout(n2485),.clk(gclk));
	jxor g2432(.dina(w_n1434_3[2]),.dinb(w_n1485_2[2]),.dout(n2486),.clk(gclk));
	jnot g2433(.din(w_n2486_0[1]),.dout(n2487),.clk(gclk));
	jand g2434(.dina(n2487),.dinb(w_n1957_0[1]),.dout(n2488),.clk(gclk));
	jand g2435(.dina(w_n2488_3[2]),.dinb(w_n1956_5[2]),.dout(n2489),.clk(gclk));
	jnot g2436(.din(w_n2483_1[0]),.dout(n2490),.clk(gclk));
	jand g2437(.dina(n2490),.dinb(w_n1958_0[2]),.dout(n2491),.clk(gclk));
	jand g2438(.dina(w_n2491_3[2]),.dinb(w_n2094_5[1]),.dout(n2492),.clk(gclk));
	jor g2439(.dina(n2492),.dinb(n2489),.dout(n2493),.clk(gclk));
	jor g2440(.dina(n2493),.dinb(n2485),.dout(n2494),.clk(gclk));
	jand g2441(.dina(w_n1956_5[1]),.dinb(w_n1438_18[1]),.dout(n2495),.clk(gclk));
	jand g2442(.dina(w_n2495_0[1]),.dinb(w_n1958_0[1]),.dout(n2496),.clk(gclk));
	jxor g2443(.dina(n2496),.dinb(w_n2494_0[1]),.dout(n2497),.clk(gclk));
	jxor g2444(.dina(w_n2497_0[1]),.dinb(w_n2482_0[1]),.dout(n2498),.clk(gclk));
	jxor g2445(.dina(w_n2498_0[1]),.dinb(w_n2366_0[1]),.dout(n2499),.clk(gclk));
	jnot g2446(.din(n2499),.dout(n2500),.clk(gclk));
	jxor g2447(.dina(w_n1166_2[0]),.dinb(w_n1156_8[1]),.dout(n2501),.clk(gclk));
	jnot g2448(.din(w_n2501_0[2]),.dout(n2502),.clk(gclk));
	jxor g2449(.dina(w_n1272_1[1]),.dinb(w_n1257_9[2]),.dout(n2503),.clk(gclk));
	jnot g2450(.din(w_n2503_0[1]),.dout(n2504),.clk(gclk));
	jand g2451(.dina(w_n2504_0[1]),.dinb(w_n2502_0[2]),.dout(n2505),.clk(gclk));
	jnot g2452(.din(w_n2505_1[1]),.dout(n2506),.clk(gclk));
	jand g2453(.dina(w_n2134_0[1]),.dinb(w_n583_0[0]),.dout(n2507),.clk(gclk));
	jand g2454(.dina(w_n1366_1[0]),.dinb(w_n238_1[0]),.dout(n2508),.clk(gclk));
	jand g2455(.dina(w_n2508_0[1]),.dinb(n2507),.dout(n2509),.clk(gclk));
	jand g2456(.dina(w_n1002_0[0]),.dinb(w_n332_1[1]),.dout(n2510),.clk(gclk));
	jand g2457(.dina(w_n2510_0[1]),.dinb(w_n1987_0[1]),.dout(n2511),.clk(gclk));
	jand g2458(.dina(n2511),.dinb(n2509),.dout(n2512),.clk(gclk));
	jand g2459(.dina(w_n162_1[1]),.dinb(w_n124_1[2]),.dout(n2513),.clk(gclk));
	jand g2460(.dina(w_n2513_1[1]),.dinb(w_n1064_0[1]),.dout(n2514),.clk(gclk));
	jand g2461(.dina(w_n847_0[0]),.dinb(w_n539_1[0]),.dout(n2515),.clk(gclk));
	jand g2462(.dina(n2515),.dinb(n2514),.dout(n2516),.clk(gclk));
	jand g2463(.dina(n2516),.dinb(w_n531_0[0]),.dout(n2517),.clk(gclk));
	jand g2464(.dina(n2517),.dinb(w_n1249_0[0]),.dout(n2518),.clk(gclk));
	jand g2465(.dina(n2518),.dinb(n2512),.dout(n2519),.clk(gclk));
	jnot g2466(.din(w_n2519_0[2]),.dout(n2520),.clk(gclk));
	jand g2467(.dina(w_n2467_0[0]),.dinb(w_n2418_0[0]),.dout(n2521),.clk(gclk));
	jnot g2468(.din(w_n2521_0[1]),.dout(n2522),.clk(gclk));
	jnot g2469(.din(w_n2413_0[0]),.dout(n2523),.clk(gclk));
	jnot g2470(.din(w_n2278_0[0]),.dout(n2524),.clk(gclk));
	jnot g2471(.din(w_n2167_0[0]),.dout(n2525),.clk(gclk));
	jnot g2472(.din(w_n2091_0[1]),.dout(n2526),.clk(gclk));
	jor g2473(.dina(n2526),.dinb(w_n2120_0[0]),.dout(n2527),.clk(gclk));
	jand g2474(.dina(n2527),.dinb(n2525),.dout(n2528),.clk(gclk));
	jnot g2475(.din(w_n2233_0[2]),.dout(n2529),.clk(gclk));
	jor g2476(.dina(n2529),.dinb(w_n2528_0[1]),.dout(n2530),.clk(gclk));
	jand g2477(.dina(n2530),.dinb(n2524),.dout(n2531),.clk(gclk));
	jnot g2478(.din(w_n2348_0[2]),.dout(n2532),.clk(gclk));
	jor g2479(.dina(n2532),.dinb(w_n2531_0[1]),.dout(n2533),.clk(gclk));
	jand g2480(.dina(n2533),.dinb(n2523),.dout(n2534),.clk(gclk));
	jnot g2481(.din(w_n2468_1[0]),.dout(n2535),.clk(gclk));
	jor g2482(.dina(n2535),.dinb(w_n2534_0[1]),.dout(n2536),.clk(gclk));
	jand g2483(.dina(n2536),.dinb(n2522),.dout(n2537),.clk(gclk));
	jand g2484(.dina(w_n2424_0[0]),.dinb(w_n2421_0[0]),.dout(n2538),.clk(gclk));
	jand g2485(.dina(w_n2466_0[0]),.dinb(w_n2425_0[0]),.dout(n2539),.clk(gclk));
	jor g2486(.dina(n2539),.dinb(n2538),.dout(n2540),.clk(gclk));
	jand g2487(.dina(w_n2464_0[0]),.dinb(w_n2447_0[0]),.dout(n2541),.clk(gclk));
	jand g2488(.dina(w_n2465_0[0]),.dinb(w_n2444_0[0]),.dout(n2542),.clk(gclk));
	jor g2489(.dina(n2542),.dinb(n2541),.dout(n2543),.clk(gclk));
	jand g2490(.dina(w_n1505_2[2]),.dinb(w_n881_1[1]),.dout(n2544),.clk(gclk));
	jnot g2491(.din(n2544),.dout(n2545),.clk(gclk));
	jxor g2492(.dina(w_n1474_4[2]),.dinb(w_n996_1[2]),.dout(n2546),.clk(gclk));
	jor g2493(.dina(n2546),.dinb(w_n1490_3[0]),.dout(n2547),.clk(gclk));
	jand g2494(.dina(w_n1493_3[1]),.dinb(w_n880_2[1]),.dout(n2548),.clk(gclk));
	jnot g2495(.din(n2548),.dout(n2549),.clk(gclk));
	jand g2496(.dina(n2549),.dinb(n2547),.dout(n2550),.clk(gclk));
	jand g2497(.dina(n2550),.dinb(n2545),.dout(n2551),.clk(gclk));
	jand g2498(.dina(w_n1434_3[1]),.dinb(w_n1418_1[0]),.dout(n2552),.clk(gclk));
	jand g2499(.dina(w_n1622_2[2]),.dinb(w_n1416_0[2]),.dout(n2553),.clk(gclk));
	jor g2500(.dina(n2553),.dinb(n2552),.dout(n2554),.clk(gclk));
	jnot g2501(.din(n2554),.dout(n2555),.clk(gclk));
	jand g2502(.dina(w_n2051_7[1]),.dinb(w_n1170_1[1]),.dout(n2556),.clk(gclk));
	jand g2503(.dina(w_n1438_18[0]),.dinb(w_n1164_1[0]),.dout(n2557),.clk(gclk));
	jor g2504(.dina(n2557),.dinb(n2556),.dout(n2558),.clk(gclk));
	jand g2505(.dina(n2558),.dinb(n2555),.dout(n2559),.clk(gclk));
	jand g2506(.dina(w_n1551_2[0]),.dinb(w_n1485_2[1]),.dout(n2560),.clk(gclk));
	jand g2507(.dina(w_n1549_2[0]),.dinb(w_n1360_3[0]),.dout(n2561),.clk(gclk));
	jor g2508(.dina(n2561),.dinb(n2560),.dout(n2562),.clk(gclk));
	jnot g2509(.din(n2562),.dout(n2563),.clk(gclk));
	jand g2510(.dina(w_n1558_2[0]),.dinb(w_n1356_8[0]),.dout(n2564),.clk(gclk));
	jand g2511(.dina(w_n1560_2[0]),.dinb(w_n1480_7[1]),.dout(n2565),.clk(gclk));
	jor g2512(.dina(n2565),.dinb(n2564),.dout(n2566),.clk(gclk));
	jand g2513(.dina(n2566),.dinb(n2563),.dout(n2567),.clk(gclk));
	jxor g2514(.dina(w_n2567_0[1]),.dinb(w_n2559_0[1]),.dout(n2568),.clk(gclk));
	jxor g2515(.dina(w_n2568_0[1]),.dinb(w_n2551_0[1]),.dout(n2569),.clk(gclk));
	jxor g2516(.dina(w_n2569_0[1]),.dinb(w_n2543_0[1]),.dout(n2570),.clk(gclk));
	jand g2517(.dina(w_n2442_0[0]),.dinb(w_n2434_0[0]),.dout(n2571),.clk(gclk));
	jand g2518(.dina(w_n2443_0[0]),.dinb(w_n2426_0[0]),.dout(n2572),.clk(gclk));
	jor g2519(.dina(n2572),.dinb(n2571),.dout(n2573),.clk(gclk));
	jand g2520(.dina(w_n2462_0[0]),.dinb(w_n2457_0[0]),.dout(n2574),.clk(gclk));
	jand g2521(.dina(w_n2463_0[0]),.dinb(w_n2455_0[0]),.dout(n2575),.clk(gclk));
	jor g2522(.dina(n2575),.dinb(n2574),.dout(n2576),.clk(gclk));
	jxor g2523(.dina(w_n2576_0[1]),.dinb(w_n2573_0[1]),.dout(n2577),.clk(gclk));
	jand g2524(.dina(w_n1494_4[0]),.dinb(w_n1257_9[1]),.dout(n2578),.clk(gclk));
	jxor g2525(.dina(w_n2456_0[1]),.dinb(w_n1232_0[1]),.dout(n2579),.clk(gclk));
	jxor g2526(.dina(w_n2579_0[1]),.dinb(w_n2578_0[1]),.dout(n2580),.clk(gclk));
	jxor g2527(.dina(w_n2580_0[1]),.dinb(w_n2577_0[1]),.dout(n2581),.clk(gclk));
	jxor g2528(.dina(w_n2581_0[1]),.dinb(w_n2570_0[1]),.dout(n2582),.clk(gclk));
	jxor g2529(.dina(w_n2582_0[1]),.dinb(w_n2540_0[1]),.dout(n2583),.clk(gclk));
	jxor g2530(.dina(w_n2583_1[1]),.dinb(w_n2537_0[1]),.dout(n2584),.clk(gclk));
	jand g2531(.dina(n2584),.dinb(w_n2520_0[1]),.dout(n2585),.clk(gclk));
	jnot g2532(.din(w_n2412_0[1]),.dout(n2586),.clk(gclk));
	jxor g2533(.dina(w_n2468_0[2]),.dinb(w_n2534_0[0]),.dout(n2587),.clk(gclk));
	jand g2534(.dina(n2587),.dinb(w_n2586_0[1]),.dout(n2588),.clk(gclk));
	jxor g2535(.dina(w_n2348_0[1]),.dinb(w_n2531_0[0]),.dout(n2589),.clk(gclk));
	jand g2536(.dina(n2589),.dinb(w_n2372_0[0]),.dout(n2590),.clk(gclk));
	jxor g2537(.dina(w_n2233_0[1]),.dinb(w_n2528_0[0]),.dout(n2591),.clk(gclk));
	jand g2538(.dina(n2591),.dinb(w_n2260_0[0]),.dout(n2592),.clk(gclk));
	jand g2539(.dina(w_n2235_0[0]),.dinb(w_n2126_0[0]),.dout(n2593),.clk(gclk));
	jor g2540(.dina(n2593),.dinb(n2592),.dout(n2594),.clk(gclk));
	jand g2541(.dina(w_n2350_0[1]),.dinb(w_n2594_0[1]),.dout(n2595),.clk(gclk));
	jor g2542(.dina(n2595),.dinb(n2590),.dout(n2596),.clk(gclk));
	jand g2543(.dina(w_n2470_0[1]),.dinb(w_n2596_0[1]),.dout(n2597),.clk(gclk));
	jor g2544(.dina(n2597),.dinb(n2588),.dout(n2598),.clk(gclk));
	jand g2545(.dina(w_n2468_0[1]),.dinb(w_n2415_0[0]),.dout(n2599),.clk(gclk));
	jor g2546(.dina(n2599),.dinb(w_n2521_0[0]),.dout(n2600),.clk(gclk));
	jxor g2547(.dina(w_n2583_1[0]),.dinb(w_n2600_0[1]),.dout(n2601),.clk(gclk));
	jxor g2548(.dina(w_n2601_0[2]),.dinb(w_n2519_0[1]),.dout(n2602),.clk(gclk));
	jand g2549(.dina(w_n2602_0[2]),.dinb(w_n2598_0[1]),.dout(n2603),.clk(gclk));
	jor g2550(.dina(n2603),.dinb(n2585),.dout(n2604),.clk(gclk));
	jand g2551(.dina(w_n389_2[2]),.dinb(w_n120_1[1]),.dout(n2605),.clk(gclk));
	jand g2552(.dina(n2605),.dinb(w_n551_0[0]),.dout(n2606),.clk(gclk));
	jand g2553(.dina(w_n489_2[0]),.dinb(w_n215_2[0]),.dout(n2607),.clk(gclk));
	jand g2554(.dina(w_n244_1[2]),.dinb(w_n162_1[0]),.dout(n2608),.clk(gclk));
	jand g2555(.dina(w_n275_1[1]),.dinb(w_n255_1[0]),.dout(n2609),.clk(gclk));
	jand g2556(.dina(n2609),.dinb(n2608),.dout(n2610),.clk(gclk));
	jand g2557(.dina(w_n321_1[1]),.dinb(w_n288_1[0]),.dout(n2611),.clk(gclk));
	jand g2558(.dina(n2611),.dinb(n2610),.dout(n2612),.clk(gclk));
	jand g2559(.dina(n2612),.dinb(n2607),.dout(n2613),.clk(gclk));
	jand g2560(.dina(w_n448_1[0]),.dinb(w_n238_0[2]),.dout(n2614),.clk(gclk));
	jand g2561(.dina(w_n221_1[2]),.dinb(w_n124_1[1]),.dout(n2615),.clk(gclk));
	jand g2562(.dina(n2615),.dinb(w_n261_1[1]),.dout(n2616),.clk(gclk));
	jand g2563(.dina(n2616),.dinb(n2614),.dout(n2617),.clk(gclk));
	jand g2564(.dina(w_n383_1[1]),.dinb(w_n300_2[0]),.dout(n2618),.clk(gclk));
	jand g2565(.dina(w_n2618_0[1]),.dinb(w_n377_2[0]),.dout(n2619),.clk(gclk));
	jand g2566(.dina(n2619),.dinb(w_n339_2[1]),.dout(n2620),.clk(gclk));
	jand g2567(.dina(n2620),.dinb(w_n2617_0[1]),.dout(n2621),.clk(gclk));
	jand g2568(.dina(n2621),.dinb(w_n2613_0[1]),.dout(n2622),.clk(gclk));
	jand g2569(.dina(w_n427_1[1]),.dinb(w_n206_1[0]),.dout(n2623),.clk(gclk));
	jand g2570(.dina(w_n467_0[2]),.dinb(w_n460_2[0]),.dout(n2624),.clk(gclk));
	jand g2571(.dina(n2624),.dinb(w_n2623_0[2]),.dout(n2625),.clk(gclk));
	jand g2572(.dina(n2625),.dinb(w_n853_0[0]),.dout(n2626),.clk(gclk));
	jand g2573(.dina(w_n1322_1[0]),.dinb(w_n170_1[0]),.dout(n2627),.clk(gclk));
	jand g2574(.dina(w_n1035_1[2]),.dinb(w_n1005_2[1]),.dout(n2628),.clk(gclk));
	jand g2575(.dina(w_n2628_0[1]),.dinb(n2627),.dout(n2629),.clk(gclk));
	jand g2576(.dina(n2629),.dinb(n2626),.dout(n2630),.clk(gclk));
	jand g2577(.dina(n2630),.dinb(w_n560_0[0]),.dout(n2631),.clk(gclk));
	jand g2578(.dina(w_n2631_0[1]),.dinb(w_n455_0[0]),.dout(n2632),.clk(gclk));
	jand g2579(.dina(w_n1095_1[2]),.dinb(w_n232_2[2]),.dout(n2633),.clk(gclk));
	jand g2580(.dina(n2633),.dinb(n2632),.dout(n2634),.clk(gclk));
	jand g2581(.dina(n2634),.dinb(n2622),.dout(n2635),.clk(gclk));
	jand g2582(.dina(n2635),.dinb(w_n2606_0[1]),.dout(n2636),.clk(gclk));
	jand g2583(.dina(w_n2582_0[0]),.dinb(w_n2540_0[0]),.dout(n2637),.clk(gclk));
	jand g2584(.dina(w_n2583_0[2]),.dinb(w_n2600_0[0]),.dout(n2638),.clk(gclk));
	jor g2585(.dina(n2638),.dinb(w_n2637_0[1]),.dout(n2639),.clk(gclk));
	jand g2586(.dina(w_n2569_0[0]),.dinb(w_n2543_0[0]),.dout(n2640),.clk(gclk));
	jand g2587(.dina(w_n2581_0[0]),.dinb(w_n2570_0[0]),.dout(n2641),.clk(gclk));
	jor g2588(.dina(n2641),.dinb(n2640),.dout(n2642),.clk(gclk));
	jand g2589(.dina(w_n2576_0[0]),.dinb(w_n2573_0[0]),.dout(n2643),.clk(gclk));
	jand g2590(.dina(w_n2580_0[0]),.dinb(w_n2577_0[0]),.dout(n2644),.clk(gclk));
	jor g2591(.dina(n2644),.dinb(n2643),.dout(n2645),.clk(gclk));
	jand g2592(.dina(w_n1551_1[2]),.dinb(w_n1622_2[1]),.dout(n2646),.clk(gclk));
	jand g2593(.dina(w_n1549_1[2]),.dinb(w_n1434_3[0]),.dout(n2647),.clk(gclk));
	jor g2594(.dina(n2647),.dinb(n2646),.dout(n2648),.clk(gclk));
	jnot g2595(.din(n2648),.dout(n2649),.clk(gclk));
	jand g2596(.dina(w_n1558_1[2]),.dinb(w_n1360_2[2]),.dout(n2650),.clk(gclk));
	jand g2597(.dina(w_n1560_1[2]),.dinb(w_n1485_2[0]),.dout(n2651),.clk(gclk));
	jor g2598(.dina(n2651),.dinb(n2650),.dout(n2652),.clk(gclk));
	jand g2599(.dina(n2652),.dinb(n2649),.dout(n2653),.clk(gclk));
	jand g2600(.dina(w_n1494_3[2]),.dinb(w_n880_2[0]),.dout(n2654),.clk(gclk));
	jnot g2601(.din(w_n1151_0[2]),.dout(n2655),.clk(gclk));
	jand g2602(.dina(w_n2051_7[0]),.dinb(w_n2655_0[1]),.dout(n2656),.clk(gclk));
	jand g2603(.dina(w_n1438_17[2]),.dinb(w_n1418_0[2]),.dout(n2657),.clk(gclk));
	jor g2604(.dina(n2657),.dinb(w_n1576_0[0]),.dout(n2658),.clk(gclk));
	jor g2605(.dina(n2658),.dinb(n2656),.dout(n2659),.clk(gclk));
	jxor g2606(.dina(w_n2659_0[1]),.dinb(w_n2654_0[2]),.dout(n2660),.clk(gclk));
	jxor g2607(.dina(w_n2660_0[1]),.dinb(w_n2653_0[1]),.dout(n2661),.clk(gclk));
	jxor g2608(.dina(w_n2661_0[1]),.dinb(w_n2645_0[1]),.dout(n2662),.clk(gclk));
	jand g2609(.dina(w_n2567_0[0]),.dinb(w_n2559_0[0]),.dout(n2663),.clk(gclk));
	jand g2610(.dina(w_n2568_0[0]),.dinb(w_n2551_0[0]),.dout(n2664),.clk(gclk));
	jor g2611(.dina(n2664),.dinb(n2663),.dout(n2665),.clk(gclk));
	jand g2612(.dina(w_n1505_2[1]),.dinb(w_n996_1[1]),.dout(n2666),.clk(gclk));
	jnot g2613(.din(n2666),.dout(n2667),.clk(gclk));
	jxor g2614(.dina(w_n1474_4[1]),.dinb(w_n1480_7[0]),.dout(n2668),.clk(gclk));
	jor g2615(.dina(n2668),.dinb(w_n1490_2[2]),.dout(n2669),.clk(gclk));
	jand g2616(.dina(w_n1493_3[0]),.dinb(w_n994_2[1]),.dout(n2670),.clk(gclk));
	jnot g2617(.din(n2670),.dout(n2671),.clk(gclk));
	jand g2618(.dina(n2671),.dinb(n2669),.dout(n2672),.clk(gclk));
	jand g2619(.dina(n2672),.dinb(n2667),.dout(n2673),.clk(gclk));
	jand g2620(.dina(w_n2456_0[0]),.dinb(w_n1232_0[0]),.dout(n2674),.clk(gclk));
	jand g2621(.dina(w_n2579_0[0]),.dinb(w_n2578_0[0]),.dout(n2675),.clk(gclk));
	jor g2622(.dina(n2675),.dinb(n2674),.dout(n2676),.clk(gclk));
	jxor g2623(.dina(w_n2676_0[1]),.dinb(w_n2673_0[1]),.dout(n2677),.clk(gclk));
	jxor g2624(.dina(w_n2677_0[1]),.dinb(w_n2665_0[1]),.dout(n2678),.clk(gclk));
	jxor g2625(.dina(w_n2678_0[1]),.dinb(w_n2662_0[1]),.dout(n2679),.clk(gclk));
	jxor g2626(.dina(w_n2679_0[1]),.dinb(w_n2642_0[1]),.dout(n2680),.clk(gclk));
	jxor g2627(.dina(w_n2680_1[1]),.dinb(w_n2639_0[1]),.dout(n2681),.clk(gclk));
	jxor g2628(.dina(w_n2681_0[2]),.dinb(w_n2636_0[2]),.dout(n2682),.clk(gclk));
	jxor g2629(.dina(w_n2682_0[2]),.dinb(w_n2604_0[1]),.dout(n2683),.clk(gclk));
	jxor g2630(.dina(w_n2602_0[1]),.dinb(w_n2598_0[0]),.dout(n2684),.clk(gclk));
	jand g2631(.dina(w_n2684_3[1]),.dinb(w_n2683_2[1]),.dout(n2685),.clk(gclk));
	jnot g2632(.din(w_n2685_0[1]),.dout(n2686),.clk(gclk));
	jxor g2633(.dina(w_n2470_0[0]),.dinb(w_n2596_0[0]),.dout(n2687),.clk(gclk));
	jand g2634(.dina(w_n2684_3[0]),.dinb(w_n2687_3[1]),.dout(n2688),.clk(gclk));
	jnot g2635(.din(w_n2688_0[1]),.dout(n2689),.clk(gclk));
	jxor g2636(.dina(w_n2350_0[0]),.dinb(w_n2594_0[0]),.dout(n2690),.clk(gclk));
	jand g2637(.dina(w_n2687_3[0]),.dinb(w_n2690_2[2]),.dout(n2691),.clk(gclk));
	jnot g2638(.din(w_n2691_0[1]),.dout(n2692),.clk(gclk));
	jxor g2639(.dina(w_n2687_2[2]),.dinb(w_n2351_6[1]),.dout(n2693),.clk(gclk));
	jor g2640(.dina(n2693),.dinb(w_n2370_0[0]),.dout(n2694),.clk(gclk));
	jand g2641(.dina(n2694),.dinb(n2692),.dout(n2695),.clk(gclk));
	jxor g2642(.dina(w_n2684_2[2]),.dinb(w_n2471_6[2]),.dout(n2696),.clk(gclk));
	jor g2643(.dina(n2696),.dinb(w_n2695_0[1]),.dout(n2697),.clk(gclk));
	jand g2644(.dina(n2697),.dinb(n2689),.dout(n2698),.clk(gclk));
	jor g2645(.dina(w_n2601_0[1]),.dinb(w_n2519_0[0]),.dout(n2699),.clk(gclk));
	jor g2646(.dina(w_n2469_0[1]),.dinb(w_n2412_0[0]),.dout(n2700),.clk(gclk));
	jxor g2647(.dina(w_n2469_0[0]),.dinb(w_n2586_0[0]),.dout(n2701),.clk(gclk));
	jor g2648(.dina(n2701),.dinb(w_n2375_0[0]),.dout(n2702),.clk(gclk));
	jand g2649(.dina(n2702),.dinb(n2700),.dout(n2703),.clk(gclk));
	jxor g2650(.dina(w_n2601_0[0]),.dinb(w_n2520_0[0]),.dout(n2704),.clk(gclk));
	jor g2651(.dina(n2704),.dinb(w_n2703_0[1]),.dout(n2705),.clk(gclk));
	jand g2652(.dina(n2705),.dinb(n2699),.dout(n2706),.clk(gclk));
	jxor g2653(.dina(w_n2682_0[1]),.dinb(w_n2706_0[1]),.dout(n2707),.clk(gclk));
	jxor g2654(.dina(w_n2684_2[1]),.dinb(w_n2707_7[1]),.dout(n2708),.clk(gclk));
	jor g2655(.dina(n2708),.dinb(w_n2698_0[1]),.dout(n2709),.clk(gclk));
	jand g2656(.dina(n2709),.dinb(n2686),.dout(n2710),.clk(gclk));
	jor g2657(.dina(w_n2681_0[1]),.dinb(w_n2636_0[1]),.dout(n2711),.clk(gclk));
	jnot g2658(.din(w_n2636_0[0]),.dout(n2712),.clk(gclk));
	jxor g2659(.dina(w_n2681_0[0]),.dinb(w_n2712_0[1]),.dout(n2713),.clk(gclk));
	jor g2660(.dina(n2713),.dinb(w_n2706_0[0]),.dout(n2714),.clk(gclk));
	jand g2661(.dina(n2714),.dinb(n2711),.dout(n2715),.clk(gclk));
	jand g2662(.dina(w_n232_2[1]),.dinb(w_n157_1[2]),.dout(n2716),.clk(gclk));
	jand g2663(.dina(n2716),.dinb(w_n481_0[1]),.dout(n2717),.clk(gclk));
	jand g2664(.dina(w_n246_0[1]),.dinb(w_n235_1[0]),.dout(n2718),.clk(gclk));
	jand g2665(.dina(n2718),.dinb(w_n2717_0[2]),.dout(n2719),.clk(gclk));
	jand g2666(.dina(w_n817_1[0]),.dinb(w_n904_0[2]),.dout(n2720),.clk(gclk));
	jand g2667(.dina(n2720),.dinb(n2719),.dout(n2721),.clk(gclk));
	jand g2668(.dina(w_n370_1[1]),.dinb(w_n355_0[0]),.dout(n2722),.clk(gclk));
	jand g2669(.dina(w_n226_1[1]),.dinb(w_n187_1[0]),.dout(n2723),.clk(gclk));
	jand g2670(.dina(w_n1095_1[1]),.dinb(w_n102_1[2]),.dout(n2724),.clk(gclk));
	jand g2671(.dina(n2724),.dinb(w_n429_0[2]),.dout(n2725),.clk(gclk));
	jand g2672(.dina(w_n2725_0[1]),.dinb(n2723),.dout(n2726),.clk(gclk));
	jand g2673(.dina(n2726),.dinb(n2722),.dout(n2727),.clk(gclk));
	jand g2674(.dina(n2727),.dinb(w_n1135_0[2]),.dout(n2728),.clk(gclk));
	jand g2675(.dina(n2728),.dinb(n2721),.dout(n2729),.clk(gclk));
	jand g2676(.dina(w_n445_0[2]),.dinb(w_n147_1[0]),.dout(n2730),.clk(gclk));
	jand g2677(.dina(n2730),.dinb(w_n240_1[1]),.dout(n2731),.clk(gclk));
	jand g2678(.dina(n2731),.dinb(w_n2729_0[1]),.dout(n2732),.clk(gclk));
	jand g2679(.dina(w_n460_1[2]),.dinb(w_n169_1[2]),.dout(n2733),.clk(gclk));
	jand g2680(.dina(n2733),.dinb(w_n600_1[0]),.dout(n2734),.clk(gclk));
	jand g2681(.dina(w_n489_1[2]),.dinb(w_n128_2[0]),.dout(n2735),.clk(gclk));
	jand g2682(.dina(n2735),.dinb(w_n378_1[2]),.dout(n2736),.clk(gclk));
	jand g2683(.dina(n2736),.dinb(w_n1093_0[0]),.dout(n2737),.clk(gclk));
	jand g2684(.dina(n2737),.dinb(n2734),.dout(n2738),.clk(gclk));
	jand g2685(.dina(w_n2738_0[2]),.dinb(w_n1105_0[0]),.dout(n2739),.clk(gclk));
	jand g2686(.dina(n2739),.dinb(w_n384_1[2]),.dout(n2740),.clk(gclk));
	jand g2687(.dina(w_n852_0[1]),.dinb(w_n439_2[0]),.dout(n2741),.clk(gclk));
	jand g2688(.dina(w_n488_2[1]),.dinb(w_n438_1[0]),.dout(n2742),.clk(gclk));
	jand g2689(.dina(n2742),.dinb(w_n280_1[1]),.dout(n2743),.clk(gclk));
	jand g2690(.dina(w_n331_1[1]),.dinb(w_n315_1[0]),.dout(n2744),.clk(gclk));
	jand g2691(.dina(w_n510_1[2]),.dinb(w_n166_1[2]),.dout(n2745),.clk(gclk));
	jand g2692(.dina(n2745),.dinb(w_n2744_0[1]),.dout(n2746),.clk(gclk));
	jand g2693(.dina(n2746),.dinb(w_n2743_0[2]),.dout(n2747),.clk(gclk));
	jand g2694(.dina(w_n1459_0[0]),.dinb(w_n191_1[2]),.dout(n2748),.clk(gclk));
	jand g2695(.dina(n2748),.dinb(w_n456_0[0]),.dout(n2749),.clk(gclk));
	jand g2696(.dina(n2749),.dinb(n2747),.dout(n2750),.clk(gclk));
	jand g2697(.dina(n2750),.dinb(n2741),.dout(n2751),.clk(gclk));
	jand g2698(.dina(w_n1452_0[0]),.dinb(w_n373_0[1]),.dout(n2752),.clk(gclk));
	jand g2699(.dina(w_n562_0[1]),.dinb(w_n377_1[2]),.dout(n2753),.clk(gclk));
	jand g2700(.dina(n2753),.dinb(n2752),.dout(n2754),.clk(gclk));
	jand g2701(.dina(w_n2142_0[1]),.dinb(w_n602_0[0]),.dout(n2755),.clk(gclk));
	jand g2702(.dina(n2755),.dinb(n2754),.dout(n2756),.clk(gclk));
	jand g2703(.dina(n2756),.dinb(w_n2751_0[1]),.dout(n2757),.clk(gclk));
	jand g2704(.dina(n2757),.dinb(n2740),.dout(n2758),.clk(gclk));
	jand g2705(.dina(n2758),.dinb(w_n2732_0[1]),.dout(n2759),.clk(gclk));
	jand g2706(.dina(w_n2679_0[0]),.dinb(w_n2642_0[0]),.dout(n2760),.clk(gclk));
	jand g2707(.dina(w_n2680_1[0]),.dinb(w_n2639_0[0]),.dout(n2761),.clk(gclk));
	jor g2708(.dina(n2761),.dinb(w_n2760_0[1]),.dout(n2762),.clk(gclk));
	jand g2709(.dina(w_n2661_0[0]),.dinb(w_n2645_0[0]),.dout(n2763),.clk(gclk));
	jand g2710(.dina(w_n2678_0[0]),.dinb(w_n2662_0[0]),.dout(n2764),.clk(gclk));
	jor g2711(.dina(n2764),.dinb(n2763),.dout(n2765),.clk(gclk));
	jand g2712(.dina(w_n2676_0[0]),.dinb(w_n2673_0[0]),.dout(n2766),.clk(gclk));
	jand g2713(.dina(w_n2677_0[0]),.dinb(w_n2665_0[0]),.dout(n2767),.clk(gclk));
	jor g2714(.dina(n2767),.dinb(n2766),.dout(n2768),.clk(gclk));
	jand g2715(.dina(w_n1494_3[1]),.dinb(w_n994_2[0]),.dout(n2769),.clk(gclk));
	jnot g2716(.din(w_n2654_0[1]),.dout(n2770),.clk(gclk));
	jxor g2717(.dina(w_n2770_0[1]),.dinb(w_n1151_0[1]),.dout(n2771),.clk(gclk));
	jxor g2718(.dina(w_n2771_0[1]),.dinb(w_n2769_0[1]),.dout(n2772),.clk(gclk));
	jxor g2719(.dina(w_n2772_0[1]),.dinb(w_n2768_0[1]),.dout(n2773),.clk(gclk));
	jnot g2720(.din(w_n2659_0[0]),.dout(n2774),.clk(gclk));
	jand g2721(.dina(n2774),.dinb(w_n2770_0[0]),.dout(n2775),.clk(gclk));
	jand g2722(.dina(w_n2660_0[0]),.dinb(w_n2653_0[0]),.dout(n2776),.clk(gclk));
	jor g2723(.dina(n2776),.dinb(n2775),.dout(n2777),.clk(gclk));
	jand g2724(.dina(w_n1549_1[1]),.dinb(w_n1438_17[1]),.dout(n2778),.clk(gclk));
	jand g2725(.dina(w_n1551_1[1]),.dinb(w_n2051_6[2]),.dout(n2779),.clk(gclk));
	jor g2726(.dina(n2779),.dinb(n2778),.dout(n2780),.clk(gclk));
	jnot g2727(.din(n2780),.dout(n2781),.clk(gclk));
	jand g2728(.dina(w_n1558_1[1]),.dinb(w_n1434_2[2]),.dout(n2782),.clk(gclk));
	jand g2729(.dina(w_n1560_1[1]),.dinb(w_n1622_2[0]),.dout(n2783),.clk(gclk));
	jor g2730(.dina(n2783),.dinb(n2782),.dout(n2784),.clk(gclk));
	jand g2731(.dina(n2784),.dinb(n2781),.dout(n2785),.clk(gclk));
	jand g2732(.dina(w_n1493_2[2]),.dinb(w_n1356_7[2]),.dout(n2786),.clk(gclk));
	jnot g2733(.din(n2786),.dout(n2787),.clk(gclk));
	jxor g2734(.dina(w_n1474_4[0]),.dinb(w_n1485_1[2]),.dout(n2788),.clk(gclk));
	jor g2735(.dina(n2788),.dinb(w_n1490_2[1]),.dout(n2789),.clk(gclk));
	jand g2736(.dina(w_n1505_2[0]),.dinb(w_n1480_6[2]),.dout(n2790),.clk(gclk));
	jnot g2737(.din(n2790),.dout(n2791),.clk(gclk));
	jand g2738(.dina(n2791),.dinb(n2789),.dout(n2792),.clk(gclk));
	jand g2739(.dina(n2792),.dinb(n2787),.dout(n2793),.clk(gclk));
	jxor g2740(.dina(w_n2793_0[1]),.dinb(w_n2785_0[1]),.dout(n2794),.clk(gclk));
	jxor g2741(.dina(w_n2794_0[1]),.dinb(w_n2777_0[1]),.dout(n2795),.clk(gclk));
	jxor g2742(.dina(w_n2795_0[1]),.dinb(w_n2773_0[1]),.dout(n2796),.clk(gclk));
	jxor g2743(.dina(w_n2796_0[1]),.dinb(w_n2765_0[1]),.dout(n2797),.clk(gclk));
	jxor g2744(.dina(w_n2797_1[1]),.dinb(w_n2762_0[1]),.dout(n2798),.clk(gclk));
	jxor g2745(.dina(w_n2798_0[2]),.dinb(w_n2759_0[2]),.dout(n2799),.clk(gclk));
	jxor g2746(.dina(w_n2799_0[2]),.dinb(w_n2715_0[1]),.dout(n2800),.clk(gclk));
	jxor g2747(.dina(w_n2800_7[1]),.dinb(w_n2707_7[0]),.dout(n2801),.clk(gclk));
	jxor g2748(.dina(w_n2801_0[1]),.dinb(w_n2710_0[1]),.dout(n2802),.clk(gclk));
	jor g2749(.dina(w_n2802_1[2]),.dinb(w_n2506_7[2]),.dout(n2803),.clk(gclk));
	jxor g2750(.dina(w_n1266_2[0]),.dinb(w_n1168_1[1]),.dout(n2804),.clk(gclk));
	jnot g2751(.din(w_n2804_0[1]),.dout(n2805),.clk(gclk));
	jand g2752(.dina(n2805),.dinb(w_n2501_0[1]),.dout(n2806),.clk(gclk));
	jnot g2753(.din(w_n2806_0[2]),.dout(n2807),.clk(gclk));
	jor g2754(.dina(w_n2807_7[2]),.dinb(w_n2707_6[2]),.dout(n2808),.clk(gclk));
	jand g2755(.dina(w_n2503_0[0]),.dinb(w_n2502_0[1]),.dout(n2809),.clk(gclk));
	jnot g2756(.din(w_n2809_0[2]),.dout(n2810),.clk(gclk));
	jor g2757(.dina(w_n2810_7[1]),.dinb(w_n2800_7[0]),.dout(n2811),.clk(gclk));
	jand g2758(.dina(n2811),.dinb(n2808),.dout(n2812),.clk(gclk));
	jxor g2759(.dina(w_n2602_0[0]),.dinb(w_n2703_0[0]),.dout(n2813),.clk(gclk));
	jand g2760(.dina(w_n2804_0[0]),.dinb(w_n2504_0[0]),.dout(n2814),.clk(gclk));
	jand g2761(.dina(n2814),.dinb(w_n2501_0[0]),.dout(n2815),.clk(gclk));
	jnot g2762(.din(w_n2815_0[2]),.dout(n2816),.clk(gclk));
	jor g2763(.dina(w_n2816_7[2]),.dinb(w_n2813_6[2]),.dout(n2817),.clk(gclk));
	jand g2764(.dina(n2817),.dinb(n2812),.dout(n2818),.clk(gclk));
	jand g2765(.dina(n2818),.dinb(n2803),.dout(n2819),.clk(gclk));
	jxor g2766(.dina(n2819),.dinb(w_n1257_9[0]),.dout(n2820),.clk(gclk));
	jor g2767(.dina(w_n2820_0[1]),.dinb(w_n2500_0[1]),.dout(n2821),.clk(gclk));
	jxor g2768(.dina(w_n2364_0[0]),.dinb(w_n2251_0[0]),.dout(n2822),.clk(gclk));
	jnot g2769(.din(n2822),.dout(n2823),.clk(gclk));
	jxor g2770(.dina(w_n2813_6[1]),.dinb(w_n2707_6[1]),.dout(n2824),.clk(gclk));
	jxor g2771(.dina(w_n2824_0[1]),.dinb(w_n2698_0[0]),.dout(n2825),.clk(gclk));
	jor g2772(.dina(w_n2825_1[2]),.dinb(w_n2506_7[1]),.dout(n2826),.clk(gclk));
	jor g2773(.dina(w_n2810_7[0]),.dinb(w_n2707_6[0]),.dout(n2827),.clk(gclk));
	jor g2774(.dina(w_n2807_7[1]),.dinb(w_n2813_6[0]),.dout(n2828),.clk(gclk));
	jand g2775(.dina(n2828),.dinb(n2827),.dout(n2829),.clk(gclk));
	jor g2776(.dina(w_n2816_7[1]),.dinb(w_n2471_6[1]),.dout(n2830),.clk(gclk));
	jand g2777(.dina(n2830),.dinb(n2829),.dout(n2831),.clk(gclk));
	jand g2778(.dina(n2831),.dinb(n2826),.dout(n2832),.clk(gclk));
	jxor g2779(.dina(n2832),.dinb(w_n1257_8[2]),.dout(n2833),.clk(gclk));
	jor g2780(.dina(w_n2833_0[1]),.dinb(w_n2823_0[1]),.dout(n2834),.clk(gclk));
	jxor g2781(.dina(w_n2813_5[2]),.dinb(w_n2471_6[0]),.dout(n2835),.clk(gclk));
	jxor g2782(.dina(w_n2835_0[1]),.dinb(w_n2695_0[0]),.dout(n2836),.clk(gclk));
	jor g2783(.dina(w_n2836_1[2]),.dinb(w_n2506_7[0]),.dout(n2837),.clk(gclk));
	jor g2784(.dina(w_n2807_7[0]),.dinb(w_n2471_5[2]),.dout(n2838),.clk(gclk));
	jor g2785(.dina(w_n2810_6[2]),.dinb(w_n2813_5[1]),.dout(n2839),.clk(gclk));
	jand g2786(.dina(n2839),.dinb(n2838),.dout(n2840),.clk(gclk));
	jor g2787(.dina(w_n2816_7[0]),.dinb(w_n2351_6[0]),.dout(n2841),.clk(gclk));
	jand g2788(.dina(n2841),.dinb(n2840),.dout(n2842),.clk(gclk));
	jand g2789(.dina(n2842),.dinb(n2837),.dout(n2843),.clk(gclk));
	jxor g2790(.dina(n2843),.dinb(w_n1257_8[1]),.dout(n2844),.clk(gclk));
	jnot g2791(.din(n2844),.dout(n2845),.clk(gclk));
	jor g2792(.dina(w_n2115_0[0]),.dinb(w_n1480_6[1]),.dout(n2846),.clk(gclk));
	jxor g2793(.dina(n2846),.dinb(w_n2248_0[0]),.dout(n2847),.clk(gclk));
	jand g2794(.dina(w_n2847_0[1]),.dinb(w_n2845_0[1]),.dout(n2848),.clk(gclk));
	jor g2795(.dina(w_n2506_6[2]),.dinb(w_n2473_1[0]),.dout(n2849),.clk(gclk));
	jor g2796(.dina(w_n2807_6[2]),.dinb(w_n2351_5[2]),.dout(n2850),.clk(gclk));
	jor g2797(.dina(w_n2810_6[1]),.dinb(w_n2471_5[1]),.dout(n2851),.clk(gclk));
	jand g2798(.dina(n2851),.dinb(n2850),.dout(n2852),.clk(gclk));
	jor g2799(.dina(w_n2816_6[2]),.dinb(w_n2256_4[0]),.dout(n2853),.clk(gclk));
	jand g2800(.dina(n2853),.dinb(n2852),.dout(n2854),.clk(gclk));
	jand g2801(.dina(n2854),.dinb(n2849),.dout(n2855),.clk(gclk));
	jxor g2802(.dina(n2855),.dinb(w_n1257_8[0]),.dout(n2856),.clk(gclk));
	jnot g2803(.din(n2856),.dout(n2857),.clk(gclk));
	jand g2804(.dina(w_n2112_1[0]),.dinb(w_n1356_7[1]),.dout(n2858),.clk(gclk));
	jxor g2805(.dina(n2858),.dinb(w_n2110_0[0]),.dout(n2859),.clk(gclk));
	jand g2806(.dina(w_n2859_0[1]),.dinb(w_n2857_0[1]),.dout(n2860),.clk(gclk));
	jand g2807(.dina(w_n2505_1[0]),.dinb(w_n2096_0[2]),.dout(n2861),.clk(gclk));
	jand g2808(.dina(w_n2806_0[1]),.dinb(w_n1956_5[0]),.dout(n2862),.clk(gclk));
	jand g2809(.dina(w_n2809_0[1]),.dinb(w_n2094_5[0]),.dout(n2863),.clk(gclk));
	jor g2810(.dina(n2863),.dinb(n2862),.dout(n2864),.clk(gclk));
	jor g2811(.dina(n2864),.dinb(n2861),.dout(n2865),.clk(gclk));
	jnot g2812(.din(w_n2865_0[1]),.dout(n2866),.clk(gclk));
	jand g2813(.dina(w_n2502_0[0]),.dinb(w_n1956_4[2]),.dout(n2867),.clk(gclk));
	jnot g2814(.din(w_n2867_1[1]),.dout(n2868),.clk(gclk));
	jand g2815(.dina(n2868),.dinb(w_n1257_7[2]),.dout(n2869),.clk(gclk));
	jand g2816(.dina(n2869),.dinb(n2866),.dout(n2870),.clk(gclk));
	jand g2817(.dina(w_n2505_0[2]),.dinb(w_n2238_1[0]),.dout(n2871),.clk(gclk));
	jand g2818(.dina(w_n2806_0[0]),.dinb(w_n2094_4[2]),.dout(n2872),.clk(gclk));
	jand g2819(.dina(w_n2809_0[0]),.dinb(w_n2236_4[1]),.dout(n2873),.clk(gclk));
	jor g2820(.dina(n2873),.dinb(n2872),.dout(n2874),.clk(gclk));
	jand g2821(.dina(w_n2815_0[1]),.dinb(w_n1956_4[1]),.dout(n2875),.clk(gclk));
	jor g2822(.dina(n2875),.dinb(n2874),.dout(n2876),.clk(gclk));
	jor g2823(.dina(n2876),.dinb(n2871),.dout(n2877),.clk(gclk));
	jnot g2824(.din(n2877),.dout(n2878),.clk(gclk));
	jand g2825(.dina(w_n2878_0[1]),.dinb(w_n2870_0[1]),.dout(n2879),.clk(gclk));
	jand g2826(.dina(w_n2879_0[1]),.dinb(w_n2112_0[2]),.dout(n2880),.clk(gclk));
	jxor g2827(.dina(w_n2879_0[0]),.dinb(w_n2112_0[1]),.dout(n2881),.clk(gclk));
	jor g2828(.dina(w_n2506_6[1]),.dinb(w_n2353_1[1]),.dout(n2882),.clk(gclk));
	jor g2829(.dina(w_n2810_6[0]),.dinb(w_n2351_5[1]),.dout(n2883),.clk(gclk));
	jor g2830(.dina(w_n2816_6[1]),.dinb(w_n2116_1[2]),.dout(n2884),.clk(gclk));
	jor g2831(.dina(w_n2807_6[1]),.dinb(w_n2256_3[2]),.dout(n2885),.clk(gclk));
	jand g2832(.dina(n2885),.dinb(n2884),.dout(n2886),.clk(gclk));
	jand g2833(.dina(n2886),.dinb(n2883),.dout(n2887),.clk(gclk));
	jand g2834(.dina(n2887),.dinb(n2882),.dout(n2888),.clk(gclk));
	jxor g2835(.dina(n2888),.dinb(w_n1259_5[2]),.dout(n2889),.clk(gclk));
	jand g2836(.dina(w_n2889_0[1]),.dinb(w_n2881_0[1]),.dout(n2890),.clk(gclk));
	jor g2837(.dina(n2890),.dinb(n2880),.dout(n2891),.clk(gclk));
	jxor g2838(.dina(w_n2859_0[0]),.dinb(w_n2857_0[0]),.dout(n2892),.clk(gclk));
	jand g2839(.dina(w_n2892_0[1]),.dinb(w_n2891_0[1]),.dout(n2893),.clk(gclk));
	jor g2840(.dina(n2893),.dinb(n2860),.dout(n2894),.clk(gclk));
	jxor g2841(.dina(w_n2847_0[0]),.dinb(w_n2845_0[0]),.dout(n2895),.clk(gclk));
	jand g2842(.dina(w_n2895_0[1]),.dinb(w_n2894_0[1]),.dout(n2896),.clk(gclk));
	jor g2843(.dina(n2896),.dinb(n2848),.dout(n2897),.clk(gclk));
	jxor g2844(.dina(w_n2833_0[0]),.dinb(w_n2823_0[0]),.dout(n2898),.clk(gclk));
	jand g2845(.dina(w_n2898_0[1]),.dinb(w_n2897_0[1]),.dout(n2899),.clk(gclk));
	jnot g2846(.din(n2899),.dout(n2900),.clk(gclk));
	jand g2847(.dina(n2900),.dinb(n2834),.dout(n2901),.clk(gclk));
	jnot g2848(.din(n2901),.dout(n2902),.clk(gclk));
	jxor g2849(.dina(w_n2820_0[0]),.dinb(w_n2500_0[0]),.dout(n2903),.clk(gclk));
	jand g2850(.dina(w_n2903_0[1]),.dinb(w_n2902_0[1]),.dout(n2904),.clk(gclk));
	jnot g2851(.din(n2904),.dout(n2905),.clk(gclk));
	jand g2852(.dina(n2905),.dinb(n2821),.dout(n2906),.clk(gclk));
	jand g2853(.dina(w_n2497_0[0]),.dinb(w_n2482_0[0]),.dout(n2907),.clk(gclk));
	jand g2854(.dina(w_n2498_0[0]),.dinb(w_n2366_0[0]),.dout(n2908),.clk(gclk));
	jor g2855(.dina(n2908),.dinb(n2907),.dout(n2909),.clk(gclk));
	jor g2856(.dina(w_n2836_1[1]),.dinb(w_n2252_7[0]),.dout(n2910),.clk(gclk));
	jor g2857(.dina(w_n2471_5[0]),.dinb(w_n2359_7[0]),.dout(n2911),.clk(gclk));
	jor g2858(.dina(w_n2813_5[0]),.dinb(w_n2355_6[2]),.dout(n2912),.clk(gclk));
	jand g2859(.dina(n2912),.dinb(n2911),.dout(n2913),.clk(gclk));
	jor g2860(.dina(w_n2351_5[0]),.dinb(w_n2357_7[0]),.dout(n2914),.clk(gclk));
	jand g2861(.dina(n2914),.dinb(n2913),.dout(n2915),.clk(gclk));
	jand g2862(.dina(n2915),.dinb(n2910),.dout(n2916),.clk(gclk));
	jxor g2863(.dina(n2916),.dinb(w_n1356_7[0]),.dout(n2917),.clk(gclk));
	jnot g2864(.din(n2917),.dout(n2918),.clk(gclk));
	jand g2865(.dina(w_n2484_1[1]),.dinb(w_n2238_0[2]),.dout(n2919),.clk(gclk));
	jand g2866(.dina(w_n2491_3[1]),.dinb(w_n2236_4[0]),.dout(n2920),.clk(gclk));
	jand g2867(.dina(w_n2488_3[1]),.dinb(w_n2094_4[1]),.dout(n2921),.clk(gclk));
	jand g2868(.dina(w_n2483_0[2]),.dinb(w_n1957_0[0]),.dout(n2922),.clk(gclk));
	jand g2869(.dina(n2922),.dinb(w_n2486_0[0]),.dout(n2923),.clk(gclk));
	jand g2870(.dina(w_n2923_3[2]),.dinb(w_n1956_4[0]),.dout(n2924),.clk(gclk));
	jor g2871(.dina(n2924),.dinb(n2921),.dout(n2925),.clk(gclk));
	jor g2872(.dina(n2925),.dinb(n2920),.dout(n2926),.clk(gclk));
	jor g2873(.dina(n2926),.dinb(n2919),.dout(n2927),.clk(gclk));
	jor g2874(.dina(w_n1959_0[0]),.dinb(w_n2051_6[1]),.dout(n2928),.clk(gclk));
	jor g2875(.dina(n2928),.dinb(w_n2494_0[0]),.dout(n2929),.clk(gclk));
	jand g2876(.dina(w_n2929_0[1]),.dinb(w_n1438_17[0]),.dout(n2930),.clk(gclk));
	jxor g2877(.dina(n2930),.dinb(w_n2927_0[1]),.dout(n2931),.clk(gclk));
	jxor g2878(.dina(w_n2931_0[1]),.dinb(w_n2918_0[1]),.dout(n2932),.clk(gclk));
	jxor g2879(.dina(w_n2932_0[1]),.dinb(w_n2909_0[1]),.dout(n2933),.clk(gclk));
	jnot g2880(.din(n2933),.dout(n2934),.clk(gclk));
	jnot g2881(.din(w_n2637_0[0]),.dout(n2935),.clk(gclk));
	jnot g2882(.din(w_n2583_0[1]),.dout(n2936),.clk(gclk));
	jor g2883(.dina(n2936),.dinb(w_n2537_0[0]),.dout(n2937),.clk(gclk));
	jand g2884(.dina(n2937),.dinb(n2935),.dout(n2938),.clk(gclk));
	jxor g2885(.dina(w_n2680_0[2]),.dinb(w_n2938_0[1]),.dout(n2939),.clk(gclk));
	jand g2886(.dina(n2939),.dinb(w_n2712_0[0]),.dout(n2940),.clk(gclk));
	jand g2887(.dina(w_n2682_0[0]),.dinb(w_n2604_0[0]),.dout(n2941),.clk(gclk));
	jor g2888(.dina(n2941),.dinb(n2940),.dout(n2942),.clk(gclk));
	jxor g2889(.dina(w_n2799_0[1]),.dinb(w_n2942_0[1]),.dout(n2943),.clk(gclk));
	jand g2890(.dina(w_n2943_2[1]),.dinb(w_n2683_2[0]),.dout(n2944),.clk(gclk));
	jnot g2891(.din(w_n2944_0[1]),.dout(n2945),.clk(gclk));
	jxor g2892(.dina(w_n2943_2[0]),.dinb(w_n2707_5[2]),.dout(n2946),.clk(gclk));
	jor g2893(.dina(n2946),.dinb(w_n2710_0[0]),.dout(n2947),.clk(gclk));
	jand g2894(.dina(n2947),.dinb(n2945),.dout(n2948),.clk(gclk));
	jor g2895(.dina(w_n2798_0[1]),.dinb(w_n2759_0[1]),.dout(n2949),.clk(gclk));
	jnot g2896(.din(w_n2759_0[0]),.dout(n2950),.clk(gclk));
	jxor g2897(.dina(w_n2798_0[0]),.dinb(w_n2950_0[1]),.dout(n2951),.clk(gclk));
	jor g2898(.dina(n2951),.dinb(w_n2715_0[0]),.dout(n2952),.clk(gclk));
	jand g2899(.dina(n2952),.dinb(n2949),.dout(n2953),.clk(gclk));
	jand g2900(.dina(w_n535_1[2]),.dinb(w_n337_1[0]),.dout(n2954),.clk(gclk));
	jand g2901(.dina(w_n2954_0[1]),.dinb(w_n1120_0[0]),.dout(n2955),.clk(gclk));
	jand g2902(.dina(n2955),.dinb(w_n2743_0[1]),.dout(n2956),.clk(gclk));
	jand g2903(.dina(n2956),.dinb(w_n436_0[1]),.dout(n2957),.clk(gclk));
	jand g2904(.dina(w_n1322_0[2]),.dinb(w_n137_1[2]),.dout(n2958),.clk(gclk));
	jand g2905(.dina(w_n717_2[0]),.dinb(w_n386_0[0]),.dout(n2959),.clk(gclk));
	jand g2906(.dina(n2959),.dinb(n2958),.dout(n2960),.clk(gclk));
	jand g2907(.dina(n2960),.dinb(n2957),.dout(n2961),.clk(gclk));
	jand g2908(.dina(w_n1124_0[0]),.dinb(w_n396_0[0]),.dout(n2962),.clk(gclk));
	jand g2909(.dina(n2962),.dinb(w_n215_1[2]),.dout(n2963),.clk(gclk));
	jand g2910(.dina(w_n250_1[0]),.dinb(w_n204_1[0]),.dout(n2964),.clk(gclk));
	jand g2911(.dina(w_n2964_0[1]),.dinb(w_n128_1[2]),.dout(n2965),.clk(gclk));
	jand g2912(.dina(w_n1035_1[1]),.dinb(w_n94_1[2]),.dout(n2966),.clk(gclk));
	jand g2913(.dina(n2966),.dinb(w_n388_0[2]),.dout(n2967),.clk(gclk));
	jand g2914(.dina(n2967),.dinb(n2965),.dout(n2968),.clk(gclk));
	jand g2915(.dina(w_n2968_0[1]),.dinb(w_n361_1[1]),.dout(n2969),.clk(gclk));
	jand g2916(.dina(n2969),.dinb(w_n1378_0[0]),.dout(n2970),.clk(gclk));
	jand g2917(.dina(n2970),.dinb(n2963),.dout(n2971),.clk(gclk));
	jand g2918(.dina(w_n2971_0[1]),.dinb(w_n2729_0[0]),.dout(n2972),.clk(gclk));
	jand g2919(.dina(n2972),.dinb(n2961),.dout(n2973),.clk(gclk));
	jand g2920(.dina(w_n2796_0[0]),.dinb(w_n2765_0[0]),.dout(n2974),.clk(gclk));
	jand g2921(.dina(w_n2797_1[0]),.dinb(w_n2762_0[0]),.dout(n2975),.clk(gclk));
	jor g2922(.dina(n2975),.dinb(w_n2974_0[1]),.dout(n2976),.clk(gclk));
	jand g2923(.dina(w_n2772_0[0]),.dinb(w_n2768_0[0]),.dout(n2977),.clk(gclk));
	jand g2924(.dina(w_n2795_0[0]),.dinb(w_n2773_0[0]),.dout(n2978),.clk(gclk));
	jor g2925(.dina(n2978),.dinb(n2977),.dout(n2979),.clk(gclk));
	jand g2926(.dina(w_n1505_1[2]),.dinb(w_n1485_1[1]),.dout(n2980),.clk(gclk));
	jnot g2927(.din(n2980),.dout(n2981),.clk(gclk));
	jxor g2928(.dina(w_n1474_3[2]),.dinb(w_n1622_1[2]),.dout(n2982),.clk(gclk));
	jor g2929(.dina(n2982),.dinb(w_n1490_2[0]),.dout(n2983),.clk(gclk));
	jand g2930(.dina(w_n1493_2[1]),.dinb(w_n1360_2[1]),.dout(n2984),.clk(gclk));
	jnot g2931(.din(n2984),.dout(n2985),.clk(gclk));
	jand g2932(.dina(n2985),.dinb(n2983),.dout(n2986),.clk(gclk));
	jand g2933(.dina(n2986),.dinb(n2981),.dout(n2987),.clk(gclk));
	jand g2934(.dina(w_n1494_3[0]),.dinb(w_n1356_6[2]),.dout(n2988),.clk(gclk));
	jand g2935(.dina(w_n1438_16[2]),.dinb(w_n1555_0[0]),.dout(n2989),.clk(gclk));
	jnot g2936(.din(n2989),.dout(n2990),.clk(gclk));
	jor g2937(.dina(w_n2990_0[1]),.dinb(w_n1556_0[0]),.dout(n2991),.clk(gclk));
	jand g2938(.dina(w_n2990_0[0]),.dinb(w_n1402_0[2]),.dout(n2992),.clk(gclk));
	jnot g2939(.din(n2992),.dout(n2993),.clk(gclk));
	jand g2940(.dina(n2993),.dinb(n2991),.dout(n2994),.clk(gclk));
	jxor g2941(.dina(w_n2994_0[1]),.dinb(w_n2988_0[2]),.dout(n2995),.clk(gclk));
	jxor g2942(.dina(w_n2995_0[1]),.dinb(w_n2987_0[1]),.dout(n2996),.clk(gclk));
	jand g2943(.dina(w_n2654_0[0]),.dinb(w_n2655_0[0]),.dout(n2997),.clk(gclk));
	jand g2944(.dina(w_n2771_0[0]),.dinb(w_n2769_0[0]),.dout(n2998),.clk(gclk));
	jor g2945(.dina(n2998),.dinb(n2997),.dout(n2999),.clk(gclk));
	jand g2946(.dina(w_n2793_0[0]),.dinb(w_n2785_0[0]),.dout(n3000),.clk(gclk));
	jand g2947(.dina(w_n2794_0[0]),.dinb(w_n2777_0[0]),.dout(n3001),.clk(gclk));
	jor g2948(.dina(n3001),.dinb(n3000),.dout(n3002),.clk(gclk));
	jxor g2949(.dina(w_n3002_0[1]),.dinb(w_n2999_0[1]),.dout(n3003),.clk(gclk));
	jxor g2950(.dina(w_n3003_0[1]),.dinb(w_n2996_0[1]),.dout(n3004),.clk(gclk));
	jxor g2951(.dina(w_n3004_0[1]),.dinb(w_n2979_0[1]),.dout(n3005),.clk(gclk));
	jxor g2952(.dina(w_n3005_1[1]),.dinb(w_n2976_0[1]),.dout(n3006),.clk(gclk));
	jxor g2953(.dina(w_n3006_0[2]),.dinb(w_n2973_0[2]),.dout(n3007),.clk(gclk));
	jxor g2954(.dina(w_n3007_0[2]),.dinb(w_n2953_0[1]),.dout(n3008),.clk(gclk));
	jxor g2955(.dina(w_n3008_7[2]),.dinb(w_n2800_6[2]),.dout(n3009),.clk(gclk));
	jxor g2956(.dina(w_n3009_0[1]),.dinb(w_n2948_0[1]),.dout(n3010),.clk(gclk));
	jor g2957(.dina(w_n3010_1[2]),.dinb(w_n2506_6[0]),.dout(n3011),.clk(gclk));
	jor g2958(.dina(w_n3008_7[1]),.dinb(w_n2810_5[2]),.dout(n3012),.clk(gclk));
	jor g2959(.dina(w_n2807_6[0]),.dinb(w_n2800_6[1]),.dout(n3013),.clk(gclk));
	jand g2960(.dina(n3013),.dinb(n3012),.dout(n3014),.clk(gclk));
	jor g2961(.dina(w_n2816_6[0]),.dinb(w_n2707_5[1]),.dout(n3015),.clk(gclk));
	jand g2962(.dina(n3015),.dinb(n3014),.dout(n3016),.clk(gclk));
	jand g2963(.dina(n3016),.dinb(n3011),.dout(n3017),.clk(gclk));
	jxor g2964(.dina(n3017),.dinb(w_n1257_7[1]),.dout(n3018),.clk(gclk));
	jxor g2965(.dina(w_n3018_0[1]),.dinb(w_n2934_0[1]),.dout(n3019),.clk(gclk));
	jxor g2966(.dina(w_n3019_0[1]),.dinb(w_n2906_0[1]),.dout(n3020),.clk(gclk));
	jnot g2967(.din(w_a2_0[0]),.dout(n3021),.clk(gclk));
	jand g2968(.dina(w_n50_0[1]),.dinb(w_n49_3[1]),.dout(n3022),.clk(gclk));
	jxor g2969(.dina(n3022),.dinb(w_n3021_0[1]),.dout(n3023),.clk(gclk));
	jxor g2970(.dina(w_n3023_10[2]),.dinb(w_n519_1[2]),.dout(n3024),.clk(gclk));
	jnot g2971(.din(w_n3024_0[2]),.dout(n3025),.clk(gclk));
	jxor g2972(.dina(w_n1500_1[2]),.dinb(w_n1154_6[2]),.dout(n3026),.clk(gclk));
	jnot g2973(.din(w_n3026_0[1]),.dout(n3027),.clk(gclk));
	jand g2974(.dina(w_n3027_0[1]),.dinb(w_n3025_0[2]),.dout(n3028),.clk(gclk));
	jnot g2975(.din(w_n3028_1[1]),.dout(n3029),.clk(gclk));
	jand g2976(.dina(w_n1102_0[0]),.dinb(w_n275_1[0]),.dout(n3030),.clk(gclk));
	jand g2977(.dina(n3030),.dinb(w_n398_0[0]),.dout(n3031),.clk(gclk));
	jand g2978(.dina(n3031),.dinb(w_n1375_0[0]),.dout(n3032),.clk(gclk));
	jand g2979(.dina(w_n525_0[0]),.dinb(w_n248_1[2]),.dout(n3033),.clk(gclk));
	jand g2980(.dina(n3033),.dinb(w_n437_0[1]),.dout(n3034),.clk(gclk));
	jand g2981(.dina(w_n817_0[2]),.dinb(w_n366_1[1]),.dout(n3035),.clk(gclk));
	jand g2982(.dina(n3035),.dinb(w_n460_1[1]),.dout(n3036),.clk(gclk));
	jand g2983(.dina(n3036),.dinb(n3034),.dout(n3037),.clk(gclk));
	jand g2984(.dina(n3037),.dinb(w_n1196_0[2]),.dout(n3038),.clk(gclk));
	jand g2985(.dina(n3038),.dinb(n3032),.dout(n3039),.clk(gclk));
	jand g2986(.dina(w_n537_0[0]),.dinb(w_n344_2[0]),.dout(n3040),.clk(gclk));
	jand g2987(.dina(n3040),.dinb(n3039),.dout(n3041),.clk(gclk));
	jand g2988(.dina(n3041),.dinb(w_n896_0[1]),.dout(n3042),.clk(gclk));
	jnot g2989(.din(w_n3042_0[2]),.dout(n3043),.clk(gclk));
	jand g2990(.dina(w_n3004_0[0]),.dinb(w_n2979_0[0]),.dout(n3044),.clk(gclk));
	jnot g2991(.din(w_n3044_0[1]),.dout(n3045),.clk(gclk));
	jnot g2992(.din(w_n2974_0[0]),.dout(n3046),.clk(gclk));
	jnot g2993(.din(w_n2760_0[0]),.dout(n3047),.clk(gclk));
	jnot g2994(.din(w_n2680_0[1]),.dout(n3048),.clk(gclk));
	jor g2995(.dina(n3048),.dinb(w_n2938_0[0]),.dout(n3049),.clk(gclk));
	jand g2996(.dina(n3049),.dinb(n3047),.dout(n3050),.clk(gclk));
	jnot g2997(.din(w_n2797_0[2]),.dout(n3051),.clk(gclk));
	jor g2998(.dina(n3051),.dinb(w_n3050_0[1]),.dout(n3052),.clk(gclk));
	jand g2999(.dina(n3052),.dinb(n3046),.dout(n3053),.clk(gclk));
	jnot g3000(.din(w_n3005_1[0]),.dout(n3054),.clk(gclk));
	jor g3001(.dina(n3054),.dinb(w_n3053_0[1]),.dout(n3055),.clk(gclk));
	jand g3002(.dina(n3055),.dinb(n3045),.dout(n3056),.clk(gclk));
	jand g3003(.dina(w_n3002_0[0]),.dinb(w_n2999_0[0]),.dout(n3057),.clk(gclk));
	jand g3004(.dina(w_n3003_0[0]),.dinb(w_n2996_0[0]),.dout(n3058),.clk(gclk));
	jor g3005(.dina(n3058),.dinb(n3057),.dout(n3059),.clk(gclk));
	jand g3006(.dina(w_n1493_2[0]),.dinb(w_n1434_2[1]),.dout(n3060),.clk(gclk));
	jxor g3007(.dina(w_n1474_3[1]),.dinb(w_n1438_16[1]),.dout(n3061),.clk(gclk));
	jand g3008(.dina(n3061),.dinb(w_n517_0[0]),.dout(n3062),.clk(gclk));
	jand g3009(.dina(w_n1505_1[1]),.dinb(w_n1622_1[1]),.dout(n3063),.clk(gclk));
	jor g3010(.dina(n3063),.dinb(n3062),.dout(n3064),.clk(gclk));
	jor g3011(.dina(n3064),.dinb(n3060),.dout(n3065),.clk(gclk));
	jor g3012(.dina(w_n2994_0[0]),.dinb(w_n2988_0[1]),.dout(n3066),.clk(gclk));
	jand g3013(.dina(w_n2995_0[0]),.dinb(w_n2987_0[0]),.dout(n3067),.clk(gclk));
	jnot g3014(.din(n3067),.dout(n3068),.clk(gclk));
	jand g3015(.dina(n3068),.dinb(n3066),.dout(n3069),.clk(gclk));
	jxor g3016(.dina(w_n3069_0[1]),.dinb(w_n3065_0[1]),.dout(n3070),.clk(gclk));
	jand g3017(.dina(w_n1494_2[2]),.dinb(w_n1360_2[0]),.dout(n3071),.clk(gclk));
	jnot g3018(.din(w_n2988_0[0]),.dout(n3072),.clk(gclk));
	jxor g3019(.dina(w_n3072_0[1]),.dinb(w_n1402_0[1]),.dout(n3073),.clk(gclk));
	jxor g3020(.dina(w_n3073_0[1]),.dinb(w_n3071_0[1]),.dout(n3074),.clk(gclk));
	jxor g3021(.dina(w_n3074_0[1]),.dinb(w_n3070_0[1]),.dout(n3075),.clk(gclk));
	jxor g3022(.dina(w_n3075_0[1]),.dinb(w_n3059_0[1]),.dout(n3076),.clk(gclk));
	jxor g3023(.dina(w_n3076_0[2]),.dinb(n3056),.dout(n3077),.clk(gclk));
	jand g3024(.dina(n3077),.dinb(w_n3043_0[1]),.dout(n3078),.clk(gclk));
	jnot g3025(.din(w_n2973_0[1]),.dout(n3079),.clk(gclk));
	jxor g3026(.dina(w_n3005_0[2]),.dinb(w_n3053_0[0]),.dout(n3080),.clk(gclk));
	jand g3027(.dina(n3080),.dinb(w_n3079_0[1]),.dout(n3081),.clk(gclk));
	jxor g3028(.dina(w_n2797_0[1]),.dinb(w_n3050_0[0]),.dout(n3082),.clk(gclk));
	jand g3029(.dina(n3082),.dinb(w_n2950_0[0]),.dout(n3083),.clk(gclk));
	jand g3030(.dina(w_n2799_0[0]),.dinb(w_n2942_0[0]),.dout(n3084),.clk(gclk));
	jor g3031(.dina(n3084),.dinb(n3083),.dout(n3085),.clk(gclk));
	jand g3032(.dina(w_n3007_0[1]),.dinb(w_n3085_0[1]),.dout(n3086),.clk(gclk));
	jor g3033(.dina(n3086),.dinb(n3081),.dout(n3087),.clk(gclk));
	jand g3034(.dina(w_n3005_0[1]),.dinb(w_n2976_0[0]),.dout(n3088),.clk(gclk));
	jor g3035(.dina(n3088),.dinb(w_n3044_0[0]),.dout(n3089),.clk(gclk));
	jxor g3036(.dina(w_n3076_0[1]),.dinb(w_n3089_0[1]),.dout(n3090),.clk(gclk));
	jxor g3037(.dina(w_n3090_0[2]),.dinb(w_n3042_0[1]),.dout(n3091),.clk(gclk));
	jand g3038(.dina(w_n3091_0[2]),.dinb(w_n3087_0[1]),.dout(n3092),.clk(gclk));
	jor g3039(.dina(n3092),.dinb(n3078),.dout(n3093),.clk(gclk));
	jand g3040(.dina(w_n1095_1[0]),.dinb(w_n359_0[1]),.dout(n3094),.clk(gclk));
	jand g3041(.dina(w_n429_0[1]),.dinb(w_n94_1[1]),.dout(n3095),.clk(gclk));
	jand g3042(.dina(w_n434_1[1]),.dinb(w_n366_1[0]),.dout(n3096),.clk(gclk));
	jand g3043(.dina(n3096),.dinb(w_n389_2[1]),.dout(n3097),.clk(gclk));
	jand g3044(.dina(n3097),.dinb(n3095),.dout(n3098),.clk(gclk));
	jand g3045(.dina(w_n252_2[2]),.dinb(w_n187_0[2]),.dout(n3099),.clk(gclk));
	jand g3046(.dina(n3099),.dinb(w_n1017_0[0]),.dout(n3100),.clk(gclk));
	jand g3047(.dina(n3100),.dinb(w_n3098_0[1]),.dout(n3101),.clk(gclk));
	jand g3048(.dina(w_n309_1[0]),.dinb(w_n303_0[0]),.dout(n3102),.clk(gclk));
	jand g3049(.dina(w_n1073_0[2]),.dinb(w_n395_1[0]),.dout(n3103),.clk(gclk));
	jand g3050(.dina(n3103),.dinb(w_n222_1[2]),.dout(n3104),.clk(gclk));
	jand g3051(.dina(n3104),.dinb(n3102),.dout(n3105),.clk(gclk));
	jand g3052(.dina(n3105),.dinb(n3101),.dout(n3106),.clk(gclk));
	jand g3053(.dina(w_n3106_0[1]),.dinb(w_n897_1[1]),.dout(n3107),.clk(gclk));
	jand g3054(.dina(w_n1110_0[1]),.dinb(w_n221_1[1]),.dout(n3108),.clk(gclk));
	jand g3055(.dina(n3108),.dinb(w_n2717_0[1]),.dout(n3109),.clk(gclk));
	jand g3056(.dina(n3109),.dinb(w_n1039_0[0]),.dout(n3110),.clk(gclk));
	jand g3057(.dina(n3110),.dinb(w_n240_1[0]),.dout(n3111),.clk(gclk));
	jand g3058(.dina(n3111),.dinb(n3107),.dout(n3112),.clk(gclk));
	jand g3059(.dina(w_n1460_1[1]),.dinb(w_n148_0[1]),.dout(n3113),.clk(gclk));
	jand g3060(.dina(n3113),.dinb(w_n439_1[2]),.dout(n3114),.clk(gclk));
	jand g3061(.dina(n3114),.dinb(w_n2738_0[1]),.dout(n3115),.clk(gclk));
	jand g3062(.dina(n3115),.dinb(w_n278_0[2]),.dout(n3116),.clk(gclk));
	jand g3063(.dina(n3116),.dinb(n3112),.dout(n3117),.clk(gclk));
	jand g3064(.dina(n3117),.dinb(n3094),.dout(n3118),.clk(gclk));
	jand g3065(.dina(w_n3075_0[0]),.dinb(w_n3059_0[0]),.dout(n3119),.clk(gclk));
	jand g3066(.dina(w_n3076_0[0]),.dinb(w_n3089_0[0]),.dout(n3120),.clk(gclk));
	jor g3067(.dina(n3120),.dinb(n3119),.dout(n3121),.clk(gclk));
	jor g3068(.dina(w_n3069_0[0]),.dinb(w_n3065_0[0]),.dout(n3122),.clk(gclk));
	jand g3069(.dina(w_n3074_0[0]),.dinb(w_n3070_0[0]),.dout(n3123),.clk(gclk));
	jnot g3070(.din(n3123),.dout(n3124),.clk(gclk));
	jand g3071(.dina(n3124),.dinb(n3122),.dout(n3125),.clk(gclk));
	jnot g3072(.din(n3125),.dout(n3126),.clk(gclk));
	jand g3073(.dina(w_n3073_0[0]),.dinb(w_n3071_0[0]),.dout(n3128),.clk(gclk));
	jnot g3074(.din(n3128),.dout(n3129),.clk(gclk));
	jand g3075(.dina(n3129),.dinb(w_n3072_0[0]),.dout(n3130),.clk(gclk));
	jand g3076(.dina(w_n1494_2[1]),.dinb(w_n1434_2[0]),.dout(n3131),.clk(gclk));
	jand g3077(.dina(w_n1438_16[0]),.dinb(w_n1490_1[2]),.dout(n3132),.clk(gclk));
	jnot g3078(.din(w_n3132_0[1]),.dout(n3133),.clk(gclk));
	jor g3079(.dina(n3133),.dinb(w_n1493_1[2]),.dout(n3134),.clk(gclk));
	jor g3080(.dina(w_n3132_0[0]),.dinb(w_n1474_3[0]),.dout(n3135),.clk(gclk));
	jand g3081(.dina(n3135),.dinb(n3134),.dout(n3136),.clk(gclk));
	jxor g3082(.dina(w_n3136_0[1]),.dinb(w_n3131_0[1]),.dout(n3137),.clk(gclk));
	jnot g3083(.din(n3137),.dout(n3138),.clk(gclk));
	jxor g3084(.dina(w_n3138_0[1]),.dinb(w_n3130_0[1]),.dout(n3139),.clk(gclk));
	jxor g3085(.dina(w_n3139_0[1]),.dinb(w_n3126_0[1]),.dout(n3140),.clk(gclk));
	jxor g3086(.dina(w_n3140_0[2]),.dinb(w_n3121_0[2]),.dout(n3141),.clk(gclk));
	jxor g3087(.dina(w_n3141_0[2]),.dinb(w_n3118_0[2]),.dout(n3142),.clk(gclk));
	jxor g3088(.dina(w_n3142_0[2]),.dinb(w_n3093_0[1]),.dout(n3143),.clk(gclk));
	jxor g3089(.dina(w_n3091_0[1]),.dinb(w_n3087_0[0]),.dout(n3144),.clk(gclk));
	jand g3090(.dina(w_n3144_1[2]),.dinb(w_n3143_1[1]),.dout(n3145),.clk(gclk));
	jnot g3091(.din(w_n3145_0[1]),.dout(n3146),.clk(gclk));
	jxor g3092(.dina(w_n3007_0[0]),.dinb(w_n3085_0[0]),.dout(n3147),.clk(gclk));
	jand g3093(.dina(w_n3144_1[1]),.dinb(w_n3147_1[2]),.dout(n3148),.clk(gclk));
	jnot g3094(.din(w_n3148_0[1]),.dout(n3149),.clk(gclk));
	jand g3095(.dina(w_n3147_1[1]),.dinb(w_n2943_1[2]),.dout(n3150),.clk(gclk));
	jnot g3096(.din(w_n3150_0[1]),.dout(n3151),.clk(gclk));
	jxor g3097(.dina(w_n3147_1[0]),.dinb(w_n2800_6[0]),.dout(n3152),.clk(gclk));
	jor g3098(.dina(n3152),.dinb(w_n2948_0[0]),.dout(n3153),.clk(gclk));
	jand g3099(.dina(n3153),.dinb(n3151),.dout(n3154),.clk(gclk));
	jxor g3100(.dina(w_n3144_1[0]),.dinb(w_n3008_7[0]),.dout(n3155),.clk(gclk));
	jor g3101(.dina(n3155),.dinb(w_n3154_0[1]),.dout(n3156),.clk(gclk));
	jand g3102(.dina(n3156),.dinb(n3149),.dout(n3157),.clk(gclk));
	jor g3103(.dina(w_n3090_0[1]),.dinb(w_n3042_0[0]),.dout(n3158),.clk(gclk));
	jor g3104(.dina(w_n3006_0[1]),.dinb(w_n2973_0[0]),.dout(n3159),.clk(gclk));
	jxor g3105(.dina(w_n3006_0[0]),.dinb(w_n3079_0[0]),.dout(n3160),.clk(gclk));
	jor g3106(.dina(n3160),.dinb(w_n2953_0[0]),.dout(n3161),.clk(gclk));
	jand g3107(.dina(n3161),.dinb(n3159),.dout(n3162),.clk(gclk));
	jxor g3108(.dina(w_n3090_0[0]),.dinb(w_n3043_0[0]),.dout(n3163),.clk(gclk));
	jor g3109(.dina(n3163),.dinb(w_n3162_0[1]),.dout(n3164),.clk(gclk));
	jand g3110(.dina(n3164),.dinb(n3158),.dout(n3165),.clk(gclk));
	jxor g3111(.dina(w_n3142_0[1]),.dinb(w_n3165_0[1]),.dout(n3166),.clk(gclk));
	jxor g3112(.dina(w_n3144_0[2]),.dinb(w_n3166_8[2]),.dout(n3167),.clk(gclk));
	jor g3113(.dina(n3167),.dinb(w_n3157_0[1]),.dout(n3168),.clk(gclk));
	jand g3114(.dina(n3168),.dinb(n3146),.dout(n3169),.clk(gclk));
	jor g3115(.dina(w_n3141_0[1]),.dinb(w_n3118_0[1]),.dout(n3170),.clk(gclk));
	jnot g3116(.din(w_n3118_0[0]),.dout(n3171),.clk(gclk));
	jxor g3117(.dina(w_n3141_0[0]),.dinb(w_n3171_0[1]),.dout(n3172),.clk(gclk));
	jor g3118(.dina(n3172),.dinb(w_n3165_0[0]),.dout(n3173),.clk(gclk));
	jand g3119(.dina(n3173),.dinb(n3170),.dout(n3174),.clk(gclk));
	jand g3120(.dina(w_n587_2[0]),.dinb(w_n275_0[2]),.dout(n3175),.clk(gclk));
	jand g3121(.dina(n3175),.dinb(w_n389_2[0]),.dout(n3176),.clk(gclk));
	jand g3122(.dina(n3176),.dinb(w_n2725_0[0]),.dout(n3177),.clk(gclk));
	jand g3123(.dina(w_n3177_0[1]),.dinb(w_n198_1[0]),.dout(n3178),.clk(gclk));
	jand g3124(.dina(w_n825_0[2]),.dinb(w_n142_1[2]),.dout(n3179),.clk(gclk));
	jand g3125(.dina(w_n3179_0[2]),.dinb(w_n1979_0[0]),.dout(n3180),.clk(gclk));
	jand g3126(.dina(n3180),.dinb(n3178),.dout(n3181),.clk(gclk));
	jand g3127(.dina(n3181),.dinb(w_n2147_0[0]),.dout(n3182),.clk(gclk));
	jand g3128(.dina(w_n1005_2[0]),.dinb(w_n717_1[2]),.dout(n3183),.clk(gclk));
	jand g3129(.dina(n3183),.dinb(w_n2744_0[0]),.dout(n3184),.clk(gclk));
	jand g3130(.dina(n3184),.dinb(w_n286_1[2]),.dout(n3185),.clk(gclk));
	jand g3131(.dina(w_n3185_0[1]),.dinb(w_n1366_0[2]),.dout(n3186),.clk(gclk));
	jand g3132(.dina(n3186),.dinb(w_n912_0[1]),.dout(n3187),.clk(gclk));
	jand g3133(.dina(n3187),.dinb(w_n468_0[1]),.dout(n3188),.clk(gclk));
	jand g3134(.dina(n3188),.dinb(n3182),.dout(n3189),.clk(gclk));
	jand g3135(.dina(n3189),.dinb(w_n2386_0[0]),.dout(n3190),.clk(gclk));
	jnot g3136(.din(w_n3190_0[2]),.dout(n3191),.clk(gclk));
	jand g3137(.dina(w_n3139_0[0]),.dinb(w_n3126_0[0]),.dout(n3192),.clk(gclk));
	jand g3138(.dina(w_n3140_0[1]),.dinb(w_n3121_0[1]),.dout(n3193),.clk(gclk));
	jor g3139(.dina(n3193),.dinb(n3192),.dout(n3194),.clk(gclk));
	jxor g3140(.dina(w_n2483_0[1]),.dinb(n1442),.dout(n3195),.clk(gclk));
	jor g3141(.dina(n3195),.dinb(w_n1474_2[2]),.dout(n3196),.clk(gclk));
	jor g3142(.dina(w_n3136_0[0]),.dinb(w_n3131_0[0]),.dout(n3197),.clk(gclk));
	jor g3143(.dina(w_n3138_0[0]),.dinb(w_n3130_0[0]),.dout(n3198),.clk(gclk));
	jand g3144(.dina(n3198),.dinb(n3197),.dout(n3199),.clk(gclk));
	jxor g3145(.dina(n3199),.dinb(n3196),.dout(n3200),.clk(gclk));
	jxor g3146(.dina(w_n3200_0[1]),.dinb(w_n3194_0[1]),.dout(n3201),.clk(gclk));
	jxor g3147(.dina(w_n3201_0[2]),.dinb(w_n3191_0[2]),.dout(n3202),.clk(gclk));
	jxor g3148(.dina(w_n3202_0[1]),.dinb(w_n3174_0[1]),.dout(n3203),.clk(gclk));
	jxor g3149(.dina(w_n3203_8[1]),.dinb(w_n3166_8[1]),.dout(n3204),.clk(gclk));
	jxor g3150(.dina(w_n3204_0[1]),.dinb(w_n3169_0[1]),.dout(n3205),.clk(gclk));
	jor g3151(.dina(w_n3205_1[2]),.dinb(w_n3029_7[2]),.dout(n3206),.clk(gclk));
	jxor g3152(.dina(w_n1499_1[2]),.dinb(w_n1504_1[0]),.dout(n3207),.clk(gclk));
	jnot g3153(.din(w_n3207_0[1]),.dout(n3208),.clk(gclk));
	jand g3154(.dina(n3208),.dinb(w_n3024_0[1]),.dout(n3209),.clk(gclk));
	jnot g3155(.din(w_n3209_0[2]),.dout(n3210),.clk(gclk));
	jor g3156(.dina(w_n3210_7[2]),.dinb(w_n3166_8[0]),.dout(n3211),.clk(gclk));
	jand g3157(.dina(w_n3026_0[0]),.dinb(w_n3025_0[1]),.dout(n3212),.clk(gclk));
	jnot g3158(.din(w_n3212_0[2]),.dout(n3213),.clk(gclk));
	jor g3159(.dina(w_n3213_7[1]),.dinb(w_n3203_8[0]),.dout(n3214),.clk(gclk));
	jand g3160(.dina(n3214),.dinb(n3211),.dout(n3215),.clk(gclk));
	jxor g3161(.dina(w_n3091_0[0]),.dinb(w_n3162_0[0]),.dout(n3216),.clk(gclk));
	jand g3162(.dina(w_n3207_0[0]),.dinb(w_n3024_0[0]),.dout(n3217),.clk(gclk));
	jand g3163(.dina(n3217),.dinb(w_n3027_0[0]),.dout(n3218),.clk(gclk));
	jnot g3164(.din(w_n3218_0[2]),.dout(n3219),.clk(gclk));
	jor g3165(.dina(w_n3219_7[2]),.dinb(w_n3216_7[2]),.dout(n3220),.clk(gclk));
	jand g3166(.dina(n3220),.dinb(n3215),.dout(n3221),.clk(gclk));
	jand g3167(.dina(n3221),.dinb(n3206),.dout(n3222),.clk(gclk));
	jxor g3168(.dina(n3222),.dinb(w_n1154_6[1]),.dout(n3223),.clk(gclk));
	jor g3169(.dina(w_n3223_0[1]),.dinb(w_n3020_0[1]),.dout(n3224),.clk(gclk));
	jnot g3170(.din(n3224),.dout(n3225),.clk(gclk));
	jxor g3171(.dina(w_n2903_0[0]),.dinb(w_n2902_0[0]),.dout(n3226),.clk(gclk));
	jnot g3172(.din(n3226),.dout(n3227),.clk(gclk));
	jxor g3173(.dina(w_n3216_7[1]),.dinb(w_n3166_7[2]),.dout(n3228),.clk(gclk));
	jxor g3174(.dina(w_n3228_0[1]),.dinb(w_n3157_0[0]),.dout(n3229),.clk(gclk));
	jor g3175(.dina(w_n3229_1[2]),.dinb(w_n3029_7[1]),.dout(n3230),.clk(gclk));
	jor g3176(.dina(w_n3213_7[0]),.dinb(w_n3166_7[1]),.dout(n3231),.clk(gclk));
	jor g3177(.dina(w_n3210_7[1]),.dinb(w_n3216_7[0]),.dout(n3232),.clk(gclk));
	jand g3178(.dina(n3232),.dinb(n3231),.dout(n3233),.clk(gclk));
	jor g3179(.dina(w_n3219_7[1]),.dinb(w_n3008_6[2]),.dout(n3234),.clk(gclk));
	jand g3180(.dina(n3234),.dinb(n3233),.dout(n3235),.clk(gclk));
	jand g3181(.dina(n3235),.dinb(n3230),.dout(n3236),.clk(gclk));
	jxor g3182(.dina(n3236),.dinb(w_n1154_6[0]),.dout(n3237),.clk(gclk));
	jor g3183(.dina(w_n3237_0[1]),.dinb(w_n3227_0[1]),.dout(n3238),.clk(gclk));
	jnot g3184(.din(n3238),.dout(n3239),.clk(gclk));
	jxor g3185(.dina(w_n2898_0[0]),.dinb(w_n2897_0[0]),.dout(n3240),.clk(gclk));
	jxor g3186(.dina(w_n3216_6[2]),.dinb(w_n3008_6[1]),.dout(n3241),.clk(gclk));
	jxor g3187(.dina(w_n3241_0[1]),.dinb(w_n3154_0[0]),.dout(n3242),.clk(gclk));
	jor g3188(.dina(w_n3242_1[2]),.dinb(w_n3029_7[0]),.dout(n3243),.clk(gclk));
	jor g3189(.dina(w_n3213_6[2]),.dinb(w_n3216_6[1]),.dout(n3244),.clk(gclk));
	jor g3190(.dina(w_n3210_7[0]),.dinb(w_n3008_6[0]),.dout(n3245),.clk(gclk));
	jor g3191(.dina(w_n3219_7[0]),.dinb(w_n2800_5[2]),.dout(n3246),.clk(gclk));
	jand g3192(.dina(n3246),.dinb(n3245),.dout(n3247),.clk(gclk));
	jand g3193(.dina(n3247),.dinb(n3244),.dout(n3248),.clk(gclk));
	jand g3194(.dina(n3248),.dinb(n3243),.dout(n3249),.clk(gclk));
	jxor g3195(.dina(n3249),.dinb(w_n1156_8[0]),.dout(n3250),.clk(gclk));
	jand g3196(.dina(w_n3250_0[1]),.dinb(w_n3240_0[1]),.dout(n3251),.clk(gclk));
	jxor g3197(.dina(w_n2895_0[0]),.dinb(w_n2894_0[0]),.dout(n3252),.clk(gclk));
	jor g3198(.dina(w_n3029_6[2]),.dinb(w_n3010_1[1]),.dout(n3253),.clk(gclk));
	jor g3199(.dina(w_n3210_6[2]),.dinb(w_n2800_5[1]),.dout(n3254),.clk(gclk));
	jor g3200(.dina(w_n3213_6[1]),.dinb(w_n3008_5[2]),.dout(n3255),.clk(gclk));
	jor g3201(.dina(w_n3219_6[2]),.dinb(w_n2707_5[0]),.dout(n3256),.clk(gclk));
	jand g3202(.dina(n3256),.dinb(n3255),.dout(n3257),.clk(gclk));
	jand g3203(.dina(n3257),.dinb(n3254),.dout(n3258),.clk(gclk));
	jand g3204(.dina(n3258),.dinb(n3253),.dout(n3259),.clk(gclk));
	jxor g3205(.dina(n3259),.dinb(w_n1156_7[2]),.dout(n3260),.clk(gclk));
	jand g3206(.dina(w_n3260_0[1]),.dinb(w_n3252_0[1]),.dout(n3261),.clk(gclk));
	jxor g3207(.dina(w_n2892_0[0]),.dinb(w_n2891_0[0]),.dout(n3262),.clk(gclk));
	jor g3208(.dina(w_n3029_6[1]),.dinb(w_n2802_1[1]),.dout(n3263),.clk(gclk));
	jor g3209(.dina(w_n3213_6[0]),.dinb(w_n2800_5[0]),.dout(n3264),.clk(gclk));
	jor g3210(.dina(w_n3210_6[1]),.dinb(w_n2707_4[2]),.dout(n3265),.clk(gclk));
	jor g3211(.dina(w_n3219_6[1]),.dinb(w_n2813_4[2]),.dout(n3266),.clk(gclk));
	jand g3212(.dina(n3266),.dinb(n3265),.dout(n3267),.clk(gclk));
	jand g3213(.dina(n3267),.dinb(n3264),.dout(n3268),.clk(gclk));
	jand g3214(.dina(n3268),.dinb(n3263),.dout(n3269),.clk(gclk));
	jxor g3215(.dina(n3269),.dinb(w_n1156_7[1]),.dout(n3270),.clk(gclk));
	jand g3216(.dina(w_n3270_0[1]),.dinb(w_n3262_0[1]),.dout(n3271),.clk(gclk));
	jxor g3217(.dina(w_n2889_0[0]),.dinb(w_n2881_0[0]),.dout(n3272),.clk(gclk));
	jor g3218(.dina(w_n3029_6[0]),.dinb(w_n2825_1[1]),.dout(n3273),.clk(gclk));
	jor g3219(.dina(w_n3210_6[0]),.dinb(w_n2813_4[1]),.dout(n3274),.clk(gclk));
	jor g3220(.dina(w_n3213_5[2]),.dinb(w_n2707_4[1]),.dout(n3275),.clk(gclk));
	jor g3221(.dina(w_n3219_6[0]),.dinb(w_n2471_4[2]),.dout(n3276),.clk(gclk));
	jand g3222(.dina(n3276),.dinb(n3275),.dout(n3277),.clk(gclk));
	jand g3223(.dina(n3277),.dinb(n3274),.dout(n3278),.clk(gclk));
	jand g3224(.dina(n3278),.dinb(n3273),.dout(n3279),.clk(gclk));
	jxor g3225(.dina(n3279),.dinb(w_n1156_7[0]),.dout(n3280),.clk(gclk));
	jand g3226(.dina(w_n3280_0[1]),.dinb(w_n3272_0[1]),.dout(n3281),.clk(gclk));
	jor g3227(.dina(w_n3029_5[2]),.dinb(w_n2836_1[0]),.dout(n3282),.clk(gclk));
	jor g3228(.dina(w_n3210_5[2]),.dinb(w_n2471_4[1]),.dout(n3283),.clk(gclk));
	jor g3229(.dina(w_n3213_5[1]),.dinb(w_n2813_4[0]),.dout(n3284),.clk(gclk));
	jand g3230(.dina(n3284),.dinb(n3283),.dout(n3285),.clk(gclk));
	jor g3231(.dina(w_n3219_5[2]),.dinb(w_n2351_4[2]),.dout(n3286),.clk(gclk));
	jand g3232(.dina(n3286),.dinb(n3285),.dout(n3287),.clk(gclk));
	jand g3233(.dina(n3287),.dinb(n3282),.dout(n3288),.clk(gclk));
	jxor g3234(.dina(n3288),.dinb(w_n1154_5[2]),.dout(n3289),.clk(gclk));
	jnot g3235(.din(w_n3289_0[1]),.dout(n3290),.clk(gclk));
	jor g3236(.dina(w_n2870_0[0]),.dinb(w_n1259_5[1]),.dout(n3291),.clk(gclk));
	jxor g3237(.dina(n3291),.dinb(w_n2878_0[0]),.dout(n3292),.clk(gclk));
	jand g3238(.dina(w_n3292_0[1]),.dinb(n3290),.dout(n3293),.clk(gclk));
	jor g3239(.dina(w_n3029_5[1]),.dinb(w_n2473_0[2]),.dout(n3294),.clk(gclk));
	jor g3240(.dina(w_n3210_5[1]),.dinb(w_n2351_4[1]),.dout(n3295),.clk(gclk));
	jor g3241(.dina(w_n3213_5[0]),.dinb(w_n2471_4[0]),.dout(n3296),.clk(gclk));
	jand g3242(.dina(n3296),.dinb(n3295),.dout(n3297),.clk(gclk));
	jor g3243(.dina(w_n3219_5[1]),.dinb(w_n2256_3[1]),.dout(n3298),.clk(gclk));
	jand g3244(.dina(n3298),.dinb(n3297),.dout(n3299),.clk(gclk));
	jand g3245(.dina(n3299),.dinb(n3294),.dout(n3300),.clk(gclk));
	jxor g3246(.dina(n3300),.dinb(w_n1154_5[1]),.dout(n3301),.clk(gclk));
	jnot g3247(.din(w_n3301_0[1]),.dout(n3302),.clk(gclk));
	jand g3248(.dina(w_n2867_1[0]),.dinb(w_n1257_7[0]),.dout(n3303),.clk(gclk));
	jxor g3249(.dina(n3303),.dinb(w_n2865_0[0]),.dout(n3304),.clk(gclk));
	jand g3250(.dina(w_n3304_0[1]),.dinb(n3302),.dout(n3305),.clk(gclk));
	jand g3251(.dina(w_n3028_1[0]),.dinb(w_n2096_0[1]),.dout(n3306),.clk(gclk));
	jand g3252(.dina(w_n3212_0[1]),.dinb(w_n2094_4[0]),.dout(n3307),.clk(gclk));
	jand g3253(.dina(w_n3209_0[1]),.dinb(w_n1956_3[2]),.dout(n3308),.clk(gclk));
	jor g3254(.dina(n3308),.dinb(n3307),.dout(n3309),.clk(gclk));
	jor g3255(.dina(n3309),.dinb(n3306),.dout(n3310),.clk(gclk));
	jnot g3256(.din(n3310),.dout(n3311),.clk(gclk));
	jand g3257(.dina(w_n3025_0[0]),.dinb(w_n1956_3[1]),.dout(n3312),.clk(gclk));
	jnot g3258(.din(w_n3312_0[2]),.dout(n3313),.clk(gclk));
	jand g3259(.dina(n3313),.dinb(w_n1154_5[0]),.dout(n3314),.clk(gclk));
	jand g3260(.dina(n3314),.dinb(w_n3311_0[1]),.dout(n3315),.clk(gclk));
	jand g3261(.dina(w_n3028_0[2]),.dinb(w_n2238_0[1]),.dout(n3316),.clk(gclk));
	jand g3262(.dina(w_n3212_0[0]),.dinb(w_n2236_3[2]),.dout(n3317),.clk(gclk));
	jand g3263(.dina(w_n3209_0[0]),.dinb(w_n2094_3[2]),.dout(n3318),.clk(gclk));
	jand g3264(.dina(w_n3218_0[1]),.dinb(w_n1956_3[0]),.dout(n3319),.clk(gclk));
	jor g3265(.dina(n3319),.dinb(n3318),.dout(n3320),.clk(gclk));
	jor g3266(.dina(n3320),.dinb(n3317),.dout(n3321),.clk(gclk));
	jor g3267(.dina(n3321),.dinb(n3316),.dout(n3322),.clk(gclk));
	jnot g3268(.din(n3322),.dout(n3323),.clk(gclk));
	jand g3269(.dina(w_n3323_0[1]),.dinb(w_n3315_0[1]),.dout(n3324),.clk(gclk));
	jand g3270(.dina(w_n3324_0[1]),.dinb(w_n2867_0[2]),.dout(n3325),.clk(gclk));
	jxor g3271(.dina(w_n3324_0[0]),.dinb(w_n2867_0[1]),.dout(n3326),.clk(gclk));
	jor g3272(.dina(w_n3029_5[0]),.dinb(w_n2353_1[0]),.dout(n3327),.clk(gclk));
	jor g3273(.dina(w_n3213_4[2]),.dinb(w_n2351_4[0]),.dout(n3328),.clk(gclk));
	jor g3274(.dina(w_n3219_5[0]),.dinb(w_n2116_1[1]),.dout(n3329),.clk(gclk));
	jor g3275(.dina(w_n3210_5[0]),.dinb(w_n2256_3[0]),.dout(n3330),.clk(gclk));
	jand g3276(.dina(n3330),.dinb(n3329),.dout(n3331),.clk(gclk));
	jand g3277(.dina(n3331),.dinb(n3328),.dout(n3332),.clk(gclk));
	jand g3278(.dina(n3332),.dinb(n3327),.dout(n3333),.clk(gclk));
	jxor g3279(.dina(n3333),.dinb(w_n1156_6[2]),.dout(n3334),.clk(gclk));
	jand g3280(.dina(w_n3334_0[1]),.dinb(w_n3326_0[1]),.dout(n3335),.clk(gclk));
	jor g3281(.dina(n3335),.dinb(n3325),.dout(n3336),.clk(gclk));
	jnot g3282(.din(n3336),.dout(n3337),.clk(gclk));
	jxor g3283(.dina(w_n3304_0[0]),.dinb(w_n3301_0[0]),.dout(n3338),.clk(gclk));
	jor g3284(.dina(w_n3338_0[1]),.dinb(w_n3337_0[1]),.dout(n3339),.clk(gclk));
	jnot g3285(.din(n3339),.dout(n3340),.clk(gclk));
	jor g3286(.dina(n3340),.dinb(n3305),.dout(n3341),.clk(gclk));
	jxor g3287(.dina(w_n3292_0[0]),.dinb(w_n3289_0[0]),.dout(n3342),.clk(gclk));
	jnot g3288(.din(n3342),.dout(n3343),.clk(gclk));
	jand g3289(.dina(w_n3343_0[1]),.dinb(w_n3341_0[1]),.dout(n3344),.clk(gclk));
	jor g3290(.dina(n3344),.dinb(n3293),.dout(n3345),.clk(gclk));
	jxor g3291(.dina(w_n3280_0[0]),.dinb(w_n3272_0[0]),.dout(n3346),.clk(gclk));
	jand g3292(.dina(w_n3346_0[1]),.dinb(w_n3345_0[1]),.dout(n3347),.clk(gclk));
	jor g3293(.dina(n3347),.dinb(n3281),.dout(n3348),.clk(gclk));
	jxor g3294(.dina(w_n3270_0[0]),.dinb(w_n3262_0[0]),.dout(n3349),.clk(gclk));
	jand g3295(.dina(w_n3349_0[1]),.dinb(w_n3348_0[1]),.dout(n3350),.clk(gclk));
	jor g3296(.dina(n3350),.dinb(n3271),.dout(n3351),.clk(gclk));
	jxor g3297(.dina(w_n3260_0[0]),.dinb(w_n3252_0[0]),.dout(n3352),.clk(gclk));
	jand g3298(.dina(w_n3352_0[1]),.dinb(w_n3351_0[1]),.dout(n3353),.clk(gclk));
	jor g3299(.dina(n3353),.dinb(n3261),.dout(n3354),.clk(gclk));
	jxor g3300(.dina(w_n3250_0[0]),.dinb(w_n3240_0[0]),.dout(n3355),.clk(gclk));
	jand g3301(.dina(w_n3355_0[1]),.dinb(w_n3354_0[1]),.dout(n3356),.clk(gclk));
	jor g3302(.dina(n3356),.dinb(n3251),.dout(n3357),.clk(gclk));
	jxor g3303(.dina(w_n3237_0[0]),.dinb(w_n3227_0[0]),.dout(n3358),.clk(gclk));
	jand g3304(.dina(w_n3358_0[1]),.dinb(w_n3357_0[1]),.dout(n3359),.clk(gclk));
	jor g3305(.dina(n3359),.dinb(n3239),.dout(n3360),.clk(gclk));
	jxor g3306(.dina(w_n3223_0[0]),.dinb(w_n3020_0[0]),.dout(n3361),.clk(gclk));
	jand g3307(.dina(w_n3361_0[1]),.dinb(w_n3360_0[1]),.dout(n3362),.clk(gclk));
	jor g3308(.dina(n3362),.dinb(n3225),.dout(n3363),.clk(gclk));
	jor g3309(.dina(w_n3018_0[0]),.dinb(w_n2934_0[0]),.dout(n3364),.clk(gclk));
	jnot g3310(.din(n3364),.dout(n3365),.clk(gclk));
	jnot g3311(.din(w_n2906_0[0]),.dout(n3366),.clk(gclk));
	jand g3312(.dina(w_n3019_0[0]),.dinb(n3366),.dout(n3367),.clk(gclk));
	jor g3313(.dina(n3367),.dinb(n3365),.dout(n3368),.clk(gclk));
	jand g3314(.dina(w_n2931_0[0]),.dinb(w_n2918_0[0]),.dout(n3369),.clk(gclk));
	jand g3315(.dina(w_n2932_0[0]),.dinb(w_n2909_0[0]),.dout(n3370),.clk(gclk));
	jor g3316(.dina(n3370),.dinb(n3369),.dout(n3371),.clk(gclk));
	jor g3317(.dina(w_n2825_1[0]),.dinb(w_n2252_6[2]),.dout(n3372),.clk(gclk));
	jor g3318(.dina(w_n2707_4[0]),.dinb(w_n2355_6[1]),.dout(n3373),.clk(gclk));
	jor g3319(.dina(w_n2813_3[2]),.dinb(w_n2359_6[2]),.dout(n3374),.clk(gclk));
	jand g3320(.dina(n3374),.dinb(n3373),.dout(n3375),.clk(gclk));
	jor g3321(.dina(w_n2471_3[2]),.dinb(w_n2357_6[2]),.dout(n3376),.clk(gclk));
	jand g3322(.dina(n3376),.dinb(n3375),.dout(n3377),.clk(gclk));
	jand g3323(.dina(n3377),.dinb(n3372),.dout(n3378),.clk(gclk));
	jxor g3324(.dina(n3378),.dinb(w_n1356_6[1]),.dout(n3379),.clk(gclk));
	jnot g3325(.din(n3379),.dout(n3380),.clk(gclk));
	jnot g3326(.din(w_n2495_0[0]),.dout(n3381),.clk(gclk));
	jor g3327(.dina(w_n2929_0[0]),.dinb(w_n2927_0[0]),.dout(n3382),.clk(gclk));
	jxor g3328(.dina(w_n3382_0[1]),.dinb(w_n3381_0[1]),.dout(n3383),.clk(gclk));
	jnot g3329(.din(w_n2484_1[0]),.dout(n3384),.clk(gclk));
	jor g3330(.dina(w_n3384_7[1]),.dinb(w_n2353_0[2]),.dout(n3385),.clk(gclk));
	jnot g3331(.din(w_n2491_3[0]),.dout(n3386),.clk(gclk));
	jor g3332(.dina(w_n3386_4[1]),.dinb(w_n2351_3[2]),.dout(n3387),.clk(gclk));
	jnot g3333(.din(w_n2923_3[1]),.dout(n3388),.clk(gclk));
	jor g3334(.dina(w_n3388_4[2]),.dinb(w_n2116_1[0]),.dout(n3389),.clk(gclk));
	jnot g3335(.din(w_n2488_3[0]),.dout(n3390),.clk(gclk));
	jor g3336(.dina(w_n3390_4[2]),.dinb(w_n2256_2[2]),.dout(n3391),.clk(gclk));
	jand g3337(.dina(n3391),.dinb(n3389),.dout(n3392),.clk(gclk));
	jand g3338(.dina(n3392),.dinb(n3387),.dout(n3393),.clk(gclk));
	jand g3339(.dina(n3393),.dinb(n3385),.dout(n3394),.clk(gclk));
	jxor g3340(.dina(n3394),.dinb(w_n2051_6[0]),.dout(n3395),.clk(gclk));
	jxor g3341(.dina(w_n3395_0[1]),.dinb(n3383),.dout(n3396),.clk(gclk));
	jxor g3342(.dina(w_n3396_0[1]),.dinb(w_n3380_0[1]),.dout(n3397),.clk(gclk));
	jxor g3343(.dina(w_n3397_0[1]),.dinb(w_n3371_0[1]),.dout(n3398),.clk(gclk));
	jnot g3344(.din(n3398),.dout(n3399),.clk(gclk));
	jor g3345(.dina(w_n3242_1[1]),.dinb(w_n2506_5[2]),.dout(n3400),.clk(gclk));
	jor g3346(.dina(w_n3008_5[1]),.dinb(w_n2807_5[2]),.dout(n3401),.clk(gclk));
	jor g3347(.dina(w_n3216_6[0]),.dinb(w_n2810_5[1]),.dout(n3402),.clk(gclk));
	jand g3348(.dina(n3402),.dinb(n3401),.dout(n3403),.clk(gclk));
	jor g3349(.dina(w_n2816_5[2]),.dinb(w_n2800_4[2]),.dout(n3404),.clk(gclk));
	jand g3350(.dina(n3404),.dinb(n3403),.dout(n3405),.clk(gclk));
	jand g3351(.dina(n3405),.dinb(n3400),.dout(n3406),.clk(gclk));
	jxor g3352(.dina(n3406),.dinb(w_n1257_6[2]),.dout(n3407),.clk(gclk));
	jxor g3353(.dina(w_n3407_0[1]),.dinb(w_n3399_0[1]),.dout(n3408),.clk(gclk));
	jxor g3354(.dina(w_n3408_0[1]),.dinb(w_n3368_0[1]),.dout(n3409),.clk(gclk));
	jnot g3355(.din(w_n3140_0[0]),.dout(n3410),.clk(gclk));
	jxor g3356(.dina(n3410),.dinb(w_n3121_0[0]),.dout(n3411),.clk(gclk));
	jand g3357(.dina(n3411),.dinb(w_n3171_0[0]),.dout(n3412),.clk(gclk));
	jand g3358(.dina(w_n3142_0[0]),.dinb(w_n3093_0[0]),.dout(n3413),.clk(gclk));
	jor g3359(.dina(n3413),.dinb(n3412),.dout(n3414),.clk(gclk));
	jxor g3360(.dina(w_n3202_0[0]),.dinb(w_n3414_0[1]),.dout(n3415),.clk(gclk));
	jand g3361(.dina(w_n3415_1[1]),.dinb(w_n3143_1[0]),.dout(n3416),.clk(gclk));
	jnot g3362(.din(w_n3416_0[1]),.dout(n3417),.clk(gclk));
	jxor g3363(.dina(w_n3203_7[2]),.dinb(w_n3143_0[2]),.dout(n3418),.clk(gclk));
	jor g3364(.dina(w_n3418_0[1]),.dinb(w_n3169_0[0]),.dout(n3419),.clk(gclk));
	jand g3365(.dina(n3419),.dinb(n3417),.dout(n3420),.clk(gclk));
	jand g3366(.dina(w_n1331_0[1]),.dinb(w_n335_0[0]),.dout(n3421),.clk(gclk));
	jand g3367(.dina(w_n436_0[0]),.dinb(w_n218_1[0]),.dout(n3422),.clk(gclk));
	jand g3368(.dina(n3422),.dinb(w_n1385_0[0]),.dout(n3423),.clk(gclk));
	jand g3369(.dina(n3423),.dinb(w_n337_0[2]),.dout(n3424),.clk(gclk));
	jand g3370(.dina(n3424),.dinb(n3421),.dout(n3425),.clk(gclk));
	jand g3371(.dina(w_n1066_0[0]),.dinb(w_n427_1[0]),.dout(n3426),.clk(gclk));
	jand g3372(.dina(w_n283_1[0]),.dinb(w_n215_1[1]),.dout(n3427),.clk(gclk));
	jand g3373(.dina(n3427),.dinb(n3426),.dout(n3428),.clk(gclk));
	jand g3374(.dina(n3428),.dinb(w_n1104_0[0]),.dout(n3429),.clk(gclk));
	jand g3375(.dina(w_n567_0[0]),.dinb(w_n527_1[0]),.dout(n3430),.clk(gclk));
	jand g3376(.dina(n3430),.dinb(w_n378_1[1]),.dout(n3431),.clk(gclk));
	jand g3377(.dina(n3431),.dinb(w_n1987_0[0]),.dout(n3432),.clk(gclk));
	jand g3378(.dina(n3432),.dinb(w_n3429_0[1]),.dout(n3433),.clk(gclk));
	jand g3379(.dina(n3433),.dinb(w_n129_0[1]),.dout(n3434),.clk(gclk));
	jand g3380(.dina(n3434),.dinb(n3425),.dout(n3435),.clk(gclk));
	jnot g3381(.din(w_n3435_0[2]),.dout(n3436),.clk(gclk));
	jor g3382(.dina(w_n3201_0[1]),.dinb(w_n3191_0[1]),.dout(n3437),.clk(gclk));
	jand g3383(.dina(w_n3201_0[0]),.dinb(w_n3191_0[0]),.dout(n3438),.clk(gclk));
	jor g3384(.dina(n3438),.dinb(w_n3414_0[0]),.dout(n3439),.clk(gclk));
	jand g3385(.dina(n3439),.dinb(n3437),.dout(n3440),.clk(gclk));
	jxor g3386(.dina(w_n3440_0[1]),.dinb(n3436),.dout(n3441),.clk(gclk));
	jxor g3387(.dina(w_n3441_7[2]),.dinb(w_n3203_7[1]),.dout(n3442),.clk(gclk));
	jxor g3388(.dina(w_n3442_0[1]),.dinb(w_n3420_0[1]),.dout(n3443),.clk(gclk));
	jor g3389(.dina(w_n3443_1[2]),.dinb(w_n3029_4[2]),.dout(n3444),.clk(gclk));
	jor g3390(.dina(w_n3210_4[2]),.dinb(w_n3203_7[0]),.dout(n3445),.clk(gclk));
	jor g3391(.dina(w_n3441_7[1]),.dinb(w_n3213_4[1]),.dout(n3446),.clk(gclk));
	jor g3392(.dina(w_n3219_4[2]),.dinb(w_n3166_7[0]),.dout(n3447),.clk(gclk));
	jand g3393(.dina(n3447),.dinb(n3446),.dout(n3448),.clk(gclk));
	jand g3394(.dina(n3448),.dinb(n3445),.dout(n3449),.clk(gclk));
	jand g3395(.dina(n3449),.dinb(n3444),.dout(n3450),.clk(gclk));
	jxor g3396(.dina(n3450),.dinb(w_n1156_6[1]),.dout(n3451),.clk(gclk));
	jxor g3397(.dina(w_n3451_0[1]),.dinb(w_n3409_0[1]),.dout(n3452),.clk(gclk));
	jxor g3398(.dina(w_n3452_0[1]),.dinb(w_n3363_0[1]),.dout(n3453),.clk(gclk));
	jnot g3399(.din(n3453),.dout(n3454),.clk(gclk));
	jnot g3400(.din(w_n3023_10[1]),.dout(n3455),.clk(gclk));
	jnot g3401(.din(w_a0_0[1]),.dout(n3456),.clk(gclk));
	jor g3402(.dina(w_a22_0[1]),.dinb(w_n3456_0[2]),.dout(n3457),.clk(gclk));
	jxor g3403(.dina(n3457),.dinb(w_a1_0[1]),.dout(n3458),.clk(gclk));
	jxor g3404(.dina(n3458),.dinb(w_n3023_10[0]),.dout(n3459),.clk(gclk));
	jand g3405(.dina(w_n3459_0[1]),.dinb(w_a0_0[0]),.dout(n3460),.clk(gclk));
	jnot g3406(.din(w_n3460_0[2]),.dout(n3461),.clk(gclk));
	jnot g3407(.din(w_n3200_0[0]),.dout(n3462),.clk(gclk));
	jxor g3408(.dina(n3462),.dinb(w_n3194_0[0]),.dout(n3463),.clk(gclk));
	jand g3409(.dina(w_n3463_0[1]),.dinb(w_n3190_0[1]),.dout(n3464),.clk(gclk));
	jor g3410(.dina(w_n3463_0[0]),.dinb(w_n3190_0[0]),.dout(n3465),.clk(gclk));
	jand g3411(.dina(n3465),.dinb(w_n3174_0[0]),.dout(n3466),.clk(gclk));
	jor g3412(.dina(n3466),.dinb(n3464),.dout(n3467),.clk(gclk));
	jand g3413(.dina(n3467),.dinb(w_n3435_0[1]),.dout(n3468),.clk(gclk));
	jand g3414(.dina(w_n1110_0[0]),.dinb(w_n389_1[2]),.dout(n3469),.clk(gclk));
	jand g3415(.dina(n3469),.dinb(w_n418_0[2]),.dout(n3470),.clk(gclk));
	jand g3416(.dina(w_n3470_0[2]),.dinb(w_n1035_1[0]),.dout(n3471),.clk(gclk));
	jand g3417(.dina(w_n2717_0[0]),.dinb(w_n505_0[0]),.dout(n3472),.clk(gclk));
	jand g3418(.dina(n3472),.dinb(w_n207_1[1]),.dout(n3473),.clk(gclk));
	jand g3419(.dina(n3473),.dinb(n3471),.dout(n3474),.clk(gclk));
	jand g3420(.dina(w_n347_1[0]),.dinb(w_n265_1[0]),.dout(n3475),.clk(gclk));
	jand g3421(.dina(n3475),.dinb(w_n222_1[1]),.dout(n3476),.clk(gclk));
	jand g3422(.dina(w_n462_1[0]),.dinb(w_n434_1[0]),.dout(n3477),.clk(gclk));
	jand g3423(.dina(n3477),.dinb(w_n120_1[0]),.dout(n3478),.clk(gclk));
	jand g3424(.dina(n3478),.dinb(w_n307_0[0]),.dout(n3479),.clk(gclk));
	jand g3425(.dina(n3479),.dinb(n3476),.dout(n3480),.clk(gclk));
	jand g3426(.dina(n3480),.dinb(n3474),.dout(n3481),.clk(gclk));
	jand g3427(.dina(w_n3481_0[2]),.dinb(w_n1032_0[0]),.dout(n3482),.clk(gclk));
	jand g3428(.dina(w_n2394_0[0]),.dinb(w_n190_1[1]),.dout(n3483),.clk(gclk));
	jand g3429(.dina(n3483),.dinb(w_n1009_0[0]),.dout(n3484),.clk(gclk));
	jand g3430(.dina(w_n387_1[2]),.dinb(w_n137_1[1]),.dout(n3485),.clk(gclk));
	jand g3431(.dina(n3485),.dinb(w_n353_1[0]),.dout(n3486),.clk(gclk));
	jand g3432(.dina(n3486),.dinb(n3484),.dout(n3487),.clk(gclk));
	jand g3433(.dina(w_n290_1[1]),.dinb(w_n215_1[0]),.dout(n3488),.clk(gclk));
	jand g3434(.dina(w_n313_0[2]),.dinb(w_n142_1[1]),.dout(n3489),.clk(gclk));
	jand g3435(.dina(w_n3489_0[1]),.dinb(w_n236_0[1]),.dout(n3490),.clk(gclk));
	jand g3436(.dina(n3490),.dinb(w_n3488_0[1]),.dout(n3491),.clk(gclk));
	jand g3437(.dina(n3491),.dinb(w_n435_1[1]),.dout(n3492),.clk(gclk));
	jand g3438(.dina(n3492),.dinb(n3487),.dout(n3493),.clk(gclk));
	jand g3439(.dina(n3493),.dinb(n3482),.dout(n3494),.clk(gclk));
	jxor g3440(.dina(w_n3494_0[2]),.dinb(w_n3468_0[2]),.dout(n3495),.clk(gclk));
	jand g3441(.dina(w_n3494_0[1]),.dinb(w_n3468_0[1]),.dout(n3496),.clk(gclk));
	jnot g3442(.din(w_n1185_0[0]),.dout(n3497),.clk(gclk));
	jand g3443(.dina(w_n2127_1[0]),.dinb(w_n3497_0[2]),.dout(n3498),.clk(gclk));
	jand g3444(.dina(w_n561_0[1]),.dinb(w_n344_1[2]),.dout(n3499),.clk(gclk));
	jand g3445(.dina(n3499),.dinb(w_n1074_1[0]),.dout(n3500),.clk(gclk));
	jand g3446(.dina(n3500),.dinb(n3498),.dout(n3501),.clk(gclk));
	jand g3447(.dina(n3501),.dinb(w_n2968_0[0]),.dout(n3502),.clk(gclk));
	jand g3448(.dina(w_n897_1[0]),.dinb(w_n197_1[1]),.dout(n3503),.clk(gclk));
	jand g3449(.dina(n3503),.dinb(w_n267_1[1]),.dout(n3504),.clk(gclk));
	jand g3450(.dina(n3504),.dinb(w_n248_1[1]),.dout(n3505),.clk(gclk));
	jand g3451(.dina(n3505),.dinb(w_n2134_0[0]),.dout(n3506),.clk(gclk));
	jand g3452(.dina(n3506),.dinb(n3502),.dout(n3507),.clk(gclk));
	jand g3453(.dina(n3507),.dinb(w_n443_1[0]),.dout(n3508),.clk(gclk));
	jand g3454(.dina(n3508),.dinb(w_n1456_0[0]),.dout(n3509),.clk(gclk));
	jxor g3455(.dina(w_n3509_0[2]),.dinb(w_n3496_0[1]),.dout(n3510),.clk(gclk));
	jor g3456(.dina(w_n3510_8[2]),.dinb(w_n3495_8[1]),.dout(n3511),.clk(gclk));
	jor g3457(.dina(w_n3495_8[0]),.dinb(w_n3441_7[0]),.dout(n3512),.clk(gclk));
	jxor g3458(.dina(w_n3440_0[0]),.dinb(w_n3435_0[0]),.dout(n3513),.clk(gclk));
	jand g3459(.dina(w_n3513_1[2]),.dinb(w_n3415_1[0]),.dout(n3514),.clk(gclk));
	jnot g3460(.din(w_n3514_0[1]),.dout(n3515),.clk(gclk));
	jxor g3461(.dina(w_n3441_6[2]),.dinb(w_n3415_0[2]),.dout(n3516),.clk(gclk));
	jor g3462(.dina(n3516),.dinb(w_n3420_0[0]),.dout(n3517),.clk(gclk));
	jand g3463(.dina(n3517),.dinb(n3515),.dout(n3518),.clk(gclk));
	jnot g3464(.din(w_n3494_0[0]),.dout(n3519),.clk(gclk));
	jxor g3465(.dina(w_n3519_0[1]),.dinb(w_n3468_0[0]),.dout(n3520),.clk(gclk));
	jand g3466(.dina(w_n3520_0[2]),.dinb(w_n3513_1[1]),.dout(n3521),.clk(gclk));
	jor g3467(.dina(w_n3519_0[0]),.dinb(w_n3513_1[0]),.dout(n3522),.clk(gclk));
	jnot g3468(.din(w_n3522_0[1]),.dout(n3523),.clk(gclk));
	jor g3469(.dina(n3523),.dinb(w_n3521_0[1]),.dout(n3524),.clk(gclk));
	jor g3470(.dina(n3524),.dinb(w_n3518_0[1]),.dout(n3525),.clk(gclk));
	jand g3471(.dina(n3525),.dinb(w_n3512_0[1]),.dout(n3526),.clk(gclk));
	jand g3472(.dina(w_n3509_0[1]),.dinb(w_n3495_7[2]),.dout(n3527),.clk(gclk));
	jnot g3473(.din(n3527),.dout(n3528),.clk(gclk));
	jand g3474(.dina(n3528),.dinb(w_n3511_0[2]),.dout(n3529),.clk(gclk));
	jnot g3475(.din(w_n3529_0[2]),.dout(n3530),.clk(gclk));
	jor g3476(.dina(n3530),.dinb(w_n3526_0[1]),.dout(n3531),.clk(gclk));
	jand g3477(.dina(n3531),.dinb(w_n3511_0[1]),.dout(n3532),.clk(gclk));
	jand g3478(.dina(w_n1470_0[0]),.dinb(w_n513_0[1]),.dout(n3533),.clk(gclk));
	jand g3479(.dina(n3533),.dinb(w_n459_0[1]),.dout(n3534),.clk(gclk));
	jand g3480(.dina(w_n871_0[0]),.dinb(w_n468_0[0]),.dout(n3535),.clk(gclk));
	jand g3481(.dina(w_n1460_1[0]),.dinb(w_n539_0[2]),.dout(n3536),.clk(gclk));
	jand g3482(.dina(w_n569_1[0]),.dinb(w_n157_1[1]),.dout(n3537),.clk(gclk));
	jand g3483(.dina(w_n3537_1[2]),.dinb(w_n169_1[1]),.dout(n3538),.clk(gclk));
	jand g3484(.dina(n3538),.dinb(n3536),.dout(n3539),.clk(gclk));
	jand g3485(.dina(n3539),.dinb(n3535),.dout(n3540),.clk(gclk));
	jand g3486(.dina(n3540),.dinb(w_n443_0[2]),.dout(n3541),.clk(gclk));
	jand g3487(.dina(n3541),.dinb(w_n1444_0[0]),.dout(n3542),.clk(gclk));
	jand g3488(.dina(n3542),.dinb(n3534),.dout(n3543),.clk(gclk));
	jand g3489(.dina(w_n3543_0[2]),.dinb(w_n3510_8[1]),.dout(n3544),.clk(gclk));
	jnot g3490(.din(n3544),.dout(n3545),.clk(gclk));
	jand g3491(.dina(w_n3509_0[0]),.dinb(w_n3496_0[0]),.dout(n3546),.clk(gclk));
	jxor g3492(.dina(w_n3543_0[1]),.dinb(w_n3546_0[1]),.dout(n3547),.clk(gclk));
	jor g3493(.dina(w_n3547_7[2]),.dinb(w_n3510_8[0]),.dout(n3548),.clk(gclk));
	jand g3494(.dina(w_n3548_0[2]),.dinb(n3545),.dout(n3549),.clk(gclk));
	jxor g3495(.dina(w_n3549_0[2]),.dinb(w_n3532_0[1]),.dout(n3550),.clk(gclk));
	jor g3496(.dina(w_n3550_1[2]),.dinb(w_n3461_8[2]),.dout(n3551),.clk(gclk));
	jor g3497(.dina(w_n50_0[0]),.dinb(w_n3021_0[0]),.dout(n3552),.clk(gclk));
	jor g3498(.dina(w_n3552_7[2]),.dinb(w_n3495_7[1]),.dout(n3553),.clk(gclk));
	jor g3499(.dina(w_n3459_0[0]),.dinb(w_n3456_0[1]),.dout(n3554),.clk(gclk));
	jor g3500(.dina(w_n3554_8[1]),.dinb(w_n3547_7[1]),.dout(n3555),.clk(gclk));
	jand g3501(.dina(n3555),.dinb(n3553),.dout(n3556),.clk(gclk));
	jand g3502(.dina(w_a1_0[0]),.dinb(w_n3456_0[0]),.dout(n3557),.clk(gclk));
	jnot g3503(.din(w_n3557_1[1]),.dout(n3558),.clk(gclk));
	jor g3504(.dina(w_n3558_6[2]),.dinb(w_n3510_7[2]),.dout(n3559),.clk(gclk));
	jand g3505(.dina(n3559),.dinb(n3556),.dout(n3560),.clk(gclk));
	jand g3506(.dina(n3560),.dinb(n3551),.dout(n3561),.clk(gclk));
	jxor g3507(.dina(n3561),.dinb(w_n3455_4[2]),.dout(n3562),.clk(gclk));
	jor g3508(.dina(w_n3562_0[1]),.dinb(w_n3454_0[1]),.dout(n3563),.clk(gclk));
	jnot g3509(.din(w_n3563_0[1]),.dout(n3564),.clk(gclk));
	jxor g3510(.dina(w_n3361_0[0]),.dinb(w_n3360_0[0]),.dout(n3565),.clk(gclk));
	jxor g3511(.dina(w_n3529_0[1]),.dinb(w_n3526_0[0]),.dout(n3566),.clk(gclk));
	jor g3512(.dina(w_n3566_1[2]),.dinb(w_n3461_8[1]),.dout(n3567),.clk(gclk));
	jor g3513(.dina(w_n3554_8[0]),.dinb(w_n3510_7[1]),.dout(n3568),.clk(gclk));
	jor g3514(.dina(w_n3558_6[1]),.dinb(w_n3495_7[0]),.dout(n3569),.clk(gclk));
	jor g3515(.dina(w_n3552_7[1]),.dinb(w_n3441_6[1]),.dout(n3570),.clk(gclk));
	jand g3516(.dina(n3570),.dinb(n3569),.dout(n3571),.clk(gclk));
	jand g3517(.dina(n3571),.dinb(n3568),.dout(n3572),.clk(gclk));
	jand g3518(.dina(n3572),.dinb(n3567),.dout(n3573),.clk(gclk));
	jxor g3519(.dina(n3573),.dinb(w_n3023_9[2]),.dout(n3574),.clk(gclk));
	jand g3520(.dina(w_n3574_0[1]),.dinb(w_n3565_0[1]),.dout(n3575),.clk(gclk));
	jxor g3521(.dina(w_n3574_0[0]),.dinb(w_n3565_0[0]),.dout(n3576),.clk(gclk));
	jxor g3522(.dina(w_n3358_0[0]),.dinb(w_n3357_0[0]),.dout(n3577),.clk(gclk));
	jand g3523(.dina(w_n3522_0[0]),.dinb(w_n3512_0[0]),.dout(n3578),.clk(gclk));
	jxor g3524(.dina(w_n3578_0[1]),.dinb(w_n3518_0[0]),.dout(n3579),.clk(gclk));
	jor g3525(.dina(w_n3579_1[2]),.dinb(w_n3461_8[0]),.dout(n3580),.clk(gclk));
	jor g3526(.dina(w_n3554_7[2]),.dinb(w_n3495_6[2]),.dout(n3581),.clk(gclk));
	jor g3527(.dina(w_n3558_6[0]),.dinb(w_n3441_6[0]),.dout(n3582),.clk(gclk));
	jor g3528(.dina(w_n3552_7[0]),.dinb(w_n3203_6[2]),.dout(n3583),.clk(gclk));
	jand g3529(.dina(n3583),.dinb(n3582),.dout(n3584),.clk(gclk));
	jand g3530(.dina(n3584),.dinb(n3581),.dout(n3585),.clk(gclk));
	jand g3531(.dina(n3585),.dinb(n3580),.dout(n3586),.clk(gclk));
	jxor g3532(.dina(n3586),.dinb(w_n3023_9[1]),.dout(n3587),.clk(gclk));
	jand g3533(.dina(w_n3587_0[1]),.dinb(w_n3577_0[1]),.dout(n3588),.clk(gclk));
	jor g3534(.dina(w_n3587_0[0]),.dinb(w_n3577_0[0]),.dout(n3589),.clk(gclk));
	jxor g3535(.dina(w_n3355_0[0]),.dinb(w_n3354_0[0]),.dout(n3590),.clk(gclk));
	jor g3536(.dina(w_n3461_7[2]),.dinb(w_n3443_1[1]),.dout(n3591),.clk(gclk));
	jor g3537(.dina(w_n3558_5[2]),.dinb(w_n3203_6[1]),.dout(n3592),.clk(gclk));
	jor g3538(.dina(w_n3554_7[1]),.dinb(w_n3441_5[2]),.dout(n3593),.clk(gclk));
	jor g3539(.dina(w_n3552_6[2]),.dinb(w_n3166_6[2]),.dout(n3594),.clk(gclk));
	jand g3540(.dina(n3594),.dinb(n3593),.dout(n3595),.clk(gclk));
	jand g3541(.dina(n3595),.dinb(n3592),.dout(n3596),.clk(gclk));
	jand g3542(.dina(n3596),.dinb(n3591),.dout(n3597),.clk(gclk));
	jxor g3543(.dina(n3597),.dinb(w_n3023_9[0]),.dout(n3598),.clk(gclk));
	jor g3544(.dina(w_n3598_0[1]),.dinb(w_n3590_0[1]),.dout(n3599),.clk(gclk));
	jand g3545(.dina(w_n3598_0[0]),.dinb(w_n3590_0[0]),.dout(n3600),.clk(gclk));
	jxor g3546(.dina(w_n3352_0[0]),.dinb(w_n3351_0[0]),.dout(n3601),.clk(gclk));
	jor g3547(.dina(w_n3461_7[1]),.dinb(w_n3205_1[1]),.dout(n3602),.clk(gclk));
	jor g3548(.dina(w_n3554_7[0]),.dinb(w_n3203_6[0]),.dout(n3603),.clk(gclk));
	jor g3549(.dina(w_n3558_5[1]),.dinb(w_n3166_6[1]),.dout(n3604),.clk(gclk));
	jor g3550(.dina(w_n3552_6[1]),.dinb(w_n3216_5[2]),.dout(n3605),.clk(gclk));
	jand g3551(.dina(n3605),.dinb(n3604),.dout(n3606),.clk(gclk));
	jand g3552(.dina(n3606),.dinb(n3603),.dout(n3607),.clk(gclk));
	jand g3553(.dina(n3607),.dinb(n3602),.dout(n3608),.clk(gclk));
	jxor g3554(.dina(n3608),.dinb(w_n3023_8[2]),.dout(n3609),.clk(gclk));
	jor g3555(.dina(w_n3609_0[1]),.dinb(w_n3601_0[1]),.dout(n3610),.clk(gclk));
	jand g3556(.dina(w_n3609_0[0]),.dinb(w_n3601_0[0]),.dout(n3611),.clk(gclk));
	jxor g3557(.dina(w_n3349_0[0]),.dinb(w_n3348_0[0]),.dout(n3612),.clk(gclk));
	jor g3558(.dina(w_n3461_7[0]),.dinb(w_n3229_1[1]),.dout(n3613),.clk(gclk));
	jor g3559(.dina(w_n3554_6[2]),.dinb(w_n3166_6[0]),.dout(n3614),.clk(gclk));
	jor g3560(.dina(w_n3558_5[0]),.dinb(w_n3216_5[1]),.dout(n3615),.clk(gclk));
	jand g3561(.dina(n3615),.dinb(n3614),.dout(n3616),.clk(gclk));
	jor g3562(.dina(w_n3552_6[0]),.dinb(w_n3008_5[0]),.dout(n3617),.clk(gclk));
	jand g3563(.dina(n3617),.dinb(n3616),.dout(n3618),.clk(gclk));
	jand g3564(.dina(n3618),.dinb(n3613),.dout(n3619),.clk(gclk));
	jxor g3565(.dina(n3619),.dinb(w_n3023_8[1]),.dout(n3620),.clk(gclk));
	jor g3566(.dina(w_n3620_0[1]),.dinb(w_n3612_0[1]),.dout(n3621),.clk(gclk));
	jand g3567(.dina(w_n3620_0[0]),.dinb(w_n3612_0[0]),.dout(n3622),.clk(gclk));
	jxor g3568(.dina(w_n3346_0[0]),.dinb(w_n3345_0[0]),.dout(n3623),.clk(gclk));
	jor g3569(.dina(w_n3461_6[2]),.dinb(w_n3242_1[0]),.dout(n3624),.clk(gclk));
	jor g3570(.dina(w_n3554_6[1]),.dinb(w_n3216_5[0]),.dout(n3625),.clk(gclk));
	jor g3571(.dina(w_n3558_4[2]),.dinb(w_n3008_4[2]),.dout(n3626),.clk(gclk));
	jor g3572(.dina(w_n3552_5[2]),.dinb(w_n2800_4[1]),.dout(n3627),.clk(gclk));
	jand g3573(.dina(n3627),.dinb(n3626),.dout(n3628),.clk(gclk));
	jand g3574(.dina(n3628),.dinb(n3625),.dout(n3629),.clk(gclk));
	jand g3575(.dina(n3629),.dinb(n3624),.dout(n3630),.clk(gclk));
	jxor g3576(.dina(n3630),.dinb(w_n3023_8[0]),.dout(n3631),.clk(gclk));
	jor g3577(.dina(w_n3631_0[1]),.dinb(w_n3623_0[1]),.dout(n3632),.clk(gclk));
	jand g3578(.dina(w_n3631_0[0]),.dinb(w_n3623_0[0]),.dout(n3633),.clk(gclk));
	jxor g3579(.dina(w_n3343_0[0]),.dinb(w_n3341_0[0]),.dout(n3634),.clk(gclk));
	jor g3580(.dina(w_n3461_6[1]),.dinb(w_n3010_1[0]),.dout(n3635),.clk(gclk));
	jor g3581(.dina(w_n3554_6[0]),.dinb(w_n3008_4[1]),.dout(n3636),.clk(gclk));
	jor g3582(.dina(w_n3558_4[1]),.dinb(w_n2800_4[0]),.dout(n3637),.clk(gclk));
	jand g3583(.dina(n3637),.dinb(n3636),.dout(n3638),.clk(gclk));
	jor g3584(.dina(w_n3552_5[1]),.dinb(w_n2707_3[2]),.dout(n3639),.clk(gclk));
	jand g3585(.dina(n3639),.dinb(n3638),.dout(n3640),.clk(gclk));
	jand g3586(.dina(n3640),.dinb(n3635),.dout(n3641),.clk(gclk));
	jxor g3587(.dina(n3641),.dinb(w_n3023_7[2]),.dout(n3642),.clk(gclk));
	jor g3588(.dina(w_n3642_0[1]),.dinb(w_n3634_0[1]),.dout(n3643),.clk(gclk));
	jand g3589(.dina(w_n3642_0[0]),.dinb(w_n3634_0[0]),.dout(n3644),.clk(gclk));
	jxor g3590(.dina(w_n3338_0[0]),.dinb(w_n3337_0[0]),.dout(n3645),.clk(gclk));
	jor g3591(.dina(w_n3461_6[0]),.dinb(w_n2802_1[0]),.dout(n3646),.clk(gclk));
	jor g3592(.dina(w_n3554_5[2]),.dinb(w_n2800_3[2]),.dout(n3647),.clk(gclk));
	jor g3593(.dina(w_n3558_4[0]),.dinb(w_n2707_3[1]),.dout(n3648),.clk(gclk));
	jor g3594(.dina(w_n3552_5[0]),.dinb(w_n2813_3[1]),.dout(n3649),.clk(gclk));
	jand g3595(.dina(n3649),.dinb(n3648),.dout(n3650),.clk(gclk));
	jand g3596(.dina(n3650),.dinb(n3647),.dout(n3651),.clk(gclk));
	jand g3597(.dina(n3651),.dinb(n3646),.dout(n3652),.clk(gclk));
	jxor g3598(.dina(n3652),.dinb(w_n3023_7[1]),.dout(n3653),.clk(gclk));
	jor g3599(.dina(w_n3653_0[1]),.dinb(w_n3645_0[1]),.dout(n3654),.clk(gclk));
	jand g3600(.dina(w_n3653_0[0]),.dinb(w_n3645_0[0]),.dout(n3655),.clk(gclk));
	jxor g3601(.dina(w_n3334_0[0]),.dinb(w_n3326_0[0]),.dout(n3656),.clk(gclk));
	jor g3602(.dina(w_n3461_5[2]),.dinb(w_n2825_0[2]),.dout(n3657),.clk(gclk));
	jor g3603(.dina(w_n3554_5[1]),.dinb(w_n2707_3[0]),.dout(n3658),.clk(gclk));
	jor g3604(.dina(w_n3558_3[2]),.dinb(w_n2813_3[0]),.dout(n3659),.clk(gclk));
	jand g3605(.dina(n3659),.dinb(n3658),.dout(n3660),.clk(gclk));
	jor g3606(.dina(w_n3552_4[2]),.dinb(w_n2471_3[1]),.dout(n3661),.clk(gclk));
	jand g3607(.dina(n3661),.dinb(n3660),.dout(n3662),.clk(gclk));
	jand g3608(.dina(n3662),.dinb(n3657),.dout(n3663),.clk(gclk));
	jxor g3609(.dina(n3663),.dinb(w_n3023_7[0]),.dout(n3664),.clk(gclk));
	jor g3610(.dina(w_n3664_0[1]),.dinb(w_n3656_0[1]),.dout(n3665),.clk(gclk));
	jand g3611(.dina(w_n3557_1[0]),.dinb(w_n2094_3[1]),.dout(n3666),.clk(gclk));
	jor g3612(.dina(n3666),.dinb(w_n3023_6[2]),.dout(n3667),.clk(gclk));
	jor g3613(.dina(n3667),.dinb(w_n1956_2[2]),.dout(n3668),.clk(gclk));
	jnot g3614(.din(n3668),.dout(n3669),.clk(gclk));
	jand g3615(.dina(w_n2256_2[1]),.dinb(w_n2116_0[2]),.dout(n3670),.clk(gclk));
	jor g3616(.dina(n3670),.dinb(w_n3554_5[0]),.dout(n3671),.clk(gclk));
	jand g3617(.dina(w_n2256_2[0]),.dinb(w_n2095_0[0]),.dout(n3672),.clk(gclk));
	jor g3618(.dina(n3672),.dinb(w_n3461_5[1]),.dout(n3673),.clk(gclk));
	jand g3619(.dina(n3673),.dinb(n3671),.dout(n3674),.clk(gclk));
	jand g3620(.dina(n3674),.dinb(n3669),.dout(n3675),.clk(gclk));
	jor g3621(.dina(n3675),.dinb(w_n3312_0[1]),.dout(n3676),.clk(gclk));
	jor g3622(.dina(w_n2236_3[1]),.dinb(w_n1956_2[1]),.dout(n3677),.clk(gclk));
	jand g3623(.dina(n3677),.dinb(w_n2094_3[0]),.dout(n3678),.clk(gclk));
	jxor g3624(.dina(w_n2352_0[1]),.dinb(w_n3678_0[1]),.dout(n3679),.clk(gclk));
	jand g3625(.dina(w_n3460_0[1]),.dinb(n3679),.dout(n3680),.clk(gclk));
	jand g3626(.dina(w_n3557_0[2]),.dinb(w_n2236_3[0]),.dout(n3681),.clk(gclk));
	jnot g3627(.din(w_n3554_4[2]),.dout(n3682),.clk(gclk));
	jand g3628(.dina(w_n3682_0[1]),.dinb(w_n2690_2[1]),.dout(n3683),.clk(gclk));
	jor g3629(.dina(n3683),.dinb(w_n3681_0[1]),.dout(n3684),.clk(gclk));
	jor g3630(.dina(n3684),.dinb(n3680),.dout(n3685),.clk(gclk));
	jnot g3631(.din(w_n3552_4[1]),.dout(n3686),.clk(gclk));
	jand g3632(.dina(w_n3686_0[1]),.dinb(w_n2094_2[2]),.dout(n3687),.clk(gclk));
	jor g3633(.dina(n3687),.dinb(w_n3023_6[1]),.dout(n3688),.clk(gclk));
	jnot g3634(.din(w_n3688_0[1]),.dout(n3689),.clk(gclk));
	jor g3635(.dina(n3689),.dinb(w_n3685_0[1]),.dout(n3690),.clk(gclk));
	jor g3636(.dina(w_n3461_5[0]),.dinb(w_n2353_0[1]),.dout(n3691),.clk(gclk));
	jnot g3637(.din(w_n3681_0[0]),.dout(n3692),.clk(gclk));
	jor g3638(.dina(w_n3554_4[1]),.dinb(w_n2351_3[1]),.dout(n3693),.clk(gclk));
	jand g3639(.dina(n3693),.dinb(n3692),.dout(n3694),.clk(gclk));
	jand g3640(.dina(n3694),.dinb(n3691),.dout(n3695),.clk(gclk));
	jor g3641(.dina(w_n3695_0[1]),.dinb(w_n3023_6[0]),.dout(n3696),.clk(gclk));
	jand g3642(.dina(n3696),.dinb(n3690),.dout(n3697),.clk(gclk));
	jand g3643(.dina(n3697),.dinb(w_n3676_0[1]),.dout(n3698),.clk(gclk));
	jand g3644(.dina(w_n3312_0[0]),.dinb(w_n1154_4[2]),.dout(n3699),.clk(gclk));
	jxor g3645(.dina(n3699),.dinb(w_n3311_0[0]),.dout(n3700),.clk(gclk));
	jnot g3646(.din(w_n3700_0[1]),.dout(n3701),.clk(gclk));
	jand g3647(.dina(w_n3701_0[1]),.dinb(w_n3698_0[1]),.dout(n3702),.clk(gclk));
	jor g3648(.dina(w_n3701_0[0]),.dinb(w_n3698_0[0]),.dout(n3703),.clk(gclk));
	jor g3649(.dina(w_n3461_4[2]),.dinb(w_n2473_0[1]),.dout(n3704),.clk(gclk));
	jand g3650(.dina(w_n3557_0[1]),.dinb(w_n2690_2[0]),.dout(n3705),.clk(gclk));
	jnot g3651(.din(w_n3705_0[1]),.dout(n3706),.clk(gclk));
	jor g3652(.dina(w_n3554_4[0]),.dinb(w_n2471_3[0]),.dout(n3707),.clk(gclk));
	jand g3653(.dina(n3707),.dinb(n3706),.dout(n3708),.clk(gclk));
	jand g3654(.dina(n3708),.dinb(n3704),.dout(n3709),.clk(gclk));
	jor g3655(.dina(w_n3709_0[1]),.dinb(w_n3023_5[2]),.dout(n3710),.clk(gclk));
	jand g3656(.dina(w_n2690_1[2]),.dinb(w_n2236_2[2]),.dout(n3711),.clk(gclk));
	jand g3657(.dina(w_n2352_0[0]),.dinb(w_n3678_0[0]),.dout(n3712),.clk(gclk));
	jor g3658(.dina(n3712),.dinb(n3711),.dout(n3713),.clk(gclk));
	jxor g3659(.dina(w_n2472_0[1]),.dinb(w_n3713_0[1]),.dout(n3714),.clk(gclk));
	jand g3660(.dina(w_n3460_0[0]),.dinb(w_n3714_0[1]),.dout(n3715),.clk(gclk));
	jand g3661(.dina(w_n3682_0[0]),.dinb(w_n2687_2[1]),.dout(n3716),.clk(gclk));
	jor g3662(.dina(n3716),.dinb(w_n3705_0[0]),.dout(n3717),.clk(gclk));
	jor g3663(.dina(n3717),.dinb(n3715),.dout(n3718),.clk(gclk));
	jand g3664(.dina(w_n3686_0[0]),.dinb(w_n2236_2[1]),.dout(n3719),.clk(gclk));
	jor g3665(.dina(n3719),.dinb(w_n3023_5[1]),.dout(n3720),.clk(gclk));
	jnot g3666(.din(w_n3720_0[1]),.dout(n3721),.clk(gclk));
	jor g3667(.dina(n3721),.dinb(w_n3718_0[1]),.dout(n3722),.clk(gclk));
	jand g3668(.dina(n3722),.dinb(n3710),.dout(n3723),.clk(gclk));
	jand g3669(.dina(n3723),.dinb(n3703),.dout(n3724),.clk(gclk));
	jor g3670(.dina(n3724),.dinb(w_n3702_0[1]),.dout(n3725),.clk(gclk));
	jor g3671(.dina(w_n3461_4[1]),.dinb(w_n2836_0[2]),.dout(n3726),.clk(gclk));
	jor g3672(.dina(w_n3554_3[2]),.dinb(w_n2813_2[2]),.dout(n3727),.clk(gclk));
	jor g3673(.dina(w_n3558_3[1]),.dinb(w_n2471_2[2]),.dout(n3728),.clk(gclk));
	jor g3674(.dina(w_n3552_4[0]),.dinb(w_n2351_3[0]),.dout(n3729),.clk(gclk));
	jand g3675(.dina(n3729),.dinb(n3728),.dout(n3730),.clk(gclk));
	jand g3676(.dina(n3730),.dinb(n3727),.dout(n3731),.clk(gclk));
	jand g3677(.dina(n3731),.dinb(n3726),.dout(n3732),.clk(gclk));
	jxor g3678(.dina(n3732),.dinb(w_n3023_5[0]),.dout(n3733),.clk(gclk));
	jor g3679(.dina(w_n3733_0[2]),.dinb(w_n3725_0[1]),.dout(n3734),.clk(gclk));
	jand g3680(.dina(w_n3733_0[1]),.dinb(w_n3725_0[0]),.dout(n3735),.clk(gclk));
	jnot g3681(.din(w_n3315_0[0]),.dout(n3736),.clk(gclk));
	jand g3682(.dina(n3736),.dinb(w_n1154_4[1]),.dout(n3737),.clk(gclk));
	jxor g3683(.dina(n3737),.dinb(w_n3323_0[0]),.dout(n3738),.clk(gclk));
	jnot g3684(.din(w_n3738_0[1]),.dout(n3739),.clk(gclk));
	jor g3685(.dina(n3739),.dinb(n3735),.dout(n3740),.clk(gclk));
	jand g3686(.dina(n3740),.dinb(w_n3734_0[1]),.dout(n3741),.clk(gclk));
	jand g3687(.dina(w_n3664_0[0]),.dinb(w_n3656_0[0]),.dout(n3742),.clk(gclk));
	jor g3688(.dina(w_n3742_0[1]),.dinb(n3741),.dout(n3743),.clk(gclk));
	jand g3689(.dina(n3743),.dinb(w_n3665_0[1]),.dout(n3744),.clk(gclk));
	jor g3690(.dina(n3744),.dinb(w_n3655_0[1]),.dout(n3745),.clk(gclk));
	jand g3691(.dina(n3745),.dinb(w_n3654_0[1]),.dout(n3746),.clk(gclk));
	jor g3692(.dina(n3746),.dinb(w_n3644_0[1]),.dout(n3747),.clk(gclk));
	jand g3693(.dina(n3747),.dinb(w_n3643_0[1]),.dout(n3748),.clk(gclk));
	jor g3694(.dina(n3748),.dinb(w_n3633_0[1]),.dout(n3749),.clk(gclk));
	jand g3695(.dina(n3749),.dinb(w_n3632_0[1]),.dout(n3750),.clk(gclk));
	jor g3696(.dina(n3750),.dinb(w_n3622_0[1]),.dout(n3751),.clk(gclk));
	jand g3697(.dina(n3751),.dinb(w_n3621_0[1]),.dout(n3752),.clk(gclk));
	jor g3698(.dina(n3752),.dinb(w_n3611_0[1]),.dout(n3753),.clk(gclk));
	jand g3699(.dina(n3753),.dinb(w_n3610_0[1]),.dout(n3754),.clk(gclk));
	jor g3700(.dina(n3754),.dinb(w_n3600_0[1]),.dout(n3755),.clk(gclk));
	jand g3701(.dina(n3755),.dinb(w_n3599_0[1]),.dout(n3756),.clk(gclk));
	jand g3702(.dina(n3756),.dinb(w_n3589_0[1]),.dout(n3757),.clk(gclk));
	jor g3703(.dina(n3757),.dinb(w_n3588_0[1]),.dout(n3758),.clk(gclk));
	jand g3704(.dina(n3758),.dinb(w_n3576_0[1]),.dout(n3759),.clk(gclk));
	jor g3705(.dina(n3759),.dinb(w_n3575_0[1]),.dout(n3760),.clk(gclk));
	jxor g3706(.dina(w_n3562_0[0]),.dinb(w_n3454_0[0]),.dout(n3761),.clk(gclk));
	jand g3707(.dina(w_n3761_0[2]),.dinb(w_n3760_0[1]),.dout(n3762),.clk(gclk));
	jor g3708(.dina(n3762),.dinb(n3564),.dout(n3763),.clk(gclk));
	jand g3709(.dina(w_n3451_0[0]),.dinb(w_n3409_0[0]),.dout(n3764),.clk(gclk));
	jand g3710(.dina(w_n3452_0[0]),.dinb(w_n3363_0[0]),.dout(n3765),.clk(gclk));
	jor g3711(.dina(n3765),.dinb(n3764),.dout(n3766),.clk(gclk));
	jor g3712(.dina(w_n3407_0[0]),.dinb(w_n3399_0[0]),.dout(n3767),.clk(gclk));
	jnot g3713(.din(n3767),.dout(n3768),.clk(gclk));
	jand g3714(.dina(w_n3408_0[0]),.dinb(w_n3368_0[0]),.dout(n3769),.clk(gclk));
	jor g3715(.dina(n3769),.dinb(n3768),.dout(n3770),.clk(gclk));
	jand g3716(.dina(w_n3396_0[0]),.dinb(w_n3380_0[0]),.dout(n3771),.clk(gclk));
	jand g3717(.dina(w_n3397_0[0]),.dinb(w_n3371_0[0]),.dout(n3772),.clk(gclk));
	jor g3718(.dina(n3772),.dinb(n3771),.dout(n3773),.clk(gclk));
	jand g3719(.dina(w_n3382_0[0]),.dinb(w_n3381_0[0]),.dout(n3774),.clk(gclk));
	jnot g3720(.din(n3774),.dout(n3775),.clk(gclk));
	jand g3721(.dina(w_n3395_0[0]),.dinb(n3775),.dout(n3779),.clk(gclk));
	jnot g3722(.din(n3779),.dout(n3780),.clk(gclk));
	jand g3723(.dina(w_n2484_0[2]),.dinb(w_n3714_0[0]),.dout(n3781),.clk(gclk));
	jand g3724(.dina(w_n2491_2[2]),.dinb(w_n2687_2[0]),.dout(n3782),.clk(gclk));
	jand g3725(.dina(w_n2488_2[2]),.dinb(w_n2690_1[1]),.dout(n3783),.clk(gclk));
	jand g3726(.dina(w_n2923_3[0]),.dinb(w_n2236_2[0]),.dout(n3784),.clk(gclk));
	jor g3727(.dina(n3784),.dinb(n3783),.dout(n3785),.clk(gclk));
	jor g3728(.dina(n3785),.dinb(n3782),.dout(n3786),.clk(gclk));
	jor g3729(.dina(n3786),.dinb(n3781),.dout(n3787),.clk(gclk));
	jor g3730(.dina(w_n2094_2[1]),.dinb(w_n2051_5[2]),.dout(n3788),.clk(gclk));
	jxor g3731(.dina(n3788),.dinb(w_n3787_0[1]),.dout(n3789),.clk(gclk));
	jxor g3732(.dina(w_n3789_0[1]),.dinb(w_n3780_0[1]),.dout(n3790),.clk(gclk));
	jor g3733(.dina(w_n2802_0[2]),.dinb(w_n2252_6[1]),.dout(n3791),.clk(gclk));
	jor g3734(.dina(w_n2800_3[1]),.dinb(w_n2355_6[0]),.dout(n3792),.clk(gclk));
	jor g3735(.dina(w_n2707_2[2]),.dinb(w_n2359_6[1]),.dout(n3793),.clk(gclk));
	jor g3736(.dina(w_n2813_2[1]),.dinb(w_n2357_6[1]),.dout(n3794),.clk(gclk));
	jand g3737(.dina(n3794),.dinb(n3793),.dout(n3795),.clk(gclk));
	jand g3738(.dina(n3795),.dinb(n3792),.dout(n3796),.clk(gclk));
	jand g3739(.dina(n3796),.dinb(n3791),.dout(n3797),.clk(gclk));
	jxor g3740(.dina(n3797),.dinb(w_n1480_6[0]),.dout(n3798),.clk(gclk));
	jxor g3741(.dina(w_n3798_0[1]),.dinb(w_n3790_0[1]),.dout(n3799),.clk(gclk));
	jxor g3742(.dina(w_n3799_0[1]),.dinb(w_n3773_0[1]),.dout(n3800),.clk(gclk));
	jnot g3743(.din(n3800),.dout(n3801),.clk(gclk));
	jor g3744(.dina(w_n3229_1[0]),.dinb(w_n2506_5[1]),.dout(n3802),.clk(gclk));
	jor g3745(.dina(w_n3166_5[2]),.dinb(w_n2810_5[0]),.dout(n3803),.clk(gclk));
	jor g3746(.dina(w_n3216_4[2]),.dinb(w_n2807_5[1]),.dout(n3804),.clk(gclk));
	jand g3747(.dina(n3804),.dinb(n3803),.dout(n3805),.clk(gclk));
	jor g3748(.dina(w_n3008_4[0]),.dinb(w_n2816_5[1]),.dout(n3806),.clk(gclk));
	jand g3749(.dina(n3806),.dinb(n3805),.dout(n3807),.clk(gclk));
	jand g3750(.dina(n3807),.dinb(n3802),.dout(n3808),.clk(gclk));
	jxor g3751(.dina(n3808),.dinb(w_n1257_6[1]),.dout(n3809),.clk(gclk));
	jxor g3752(.dina(w_n3809_0[1]),.dinb(w_n3801_0[1]),.dout(n3810),.clk(gclk));
	jxor g3753(.dina(w_n3810_0[1]),.dinb(w_n3770_0[1]),.dout(n3811),.clk(gclk));
	jor g3754(.dina(w_n3579_1[1]),.dinb(w_n3029_4[1]),.dout(n3812),.clk(gclk));
	jor g3755(.dina(w_n3495_6[1]),.dinb(w_n3213_4[0]),.dout(n3813),.clk(gclk));
	jor g3756(.dina(w_n3441_5[1]),.dinb(w_n3210_4[1]),.dout(n3814),.clk(gclk));
	jor g3757(.dina(w_n3219_4[1]),.dinb(w_n3203_5[2]),.dout(n3815),.clk(gclk));
	jand g3758(.dina(n3815),.dinb(n3814),.dout(n3816),.clk(gclk));
	jand g3759(.dina(n3816),.dinb(n3813),.dout(n3817),.clk(gclk));
	jand g3760(.dina(n3817),.dinb(n3812),.dout(n3818),.clk(gclk));
	jxor g3761(.dina(n3818),.dinb(w_n1156_6[0]),.dout(n3819),.clk(gclk));
	jxor g3762(.dina(w_n3819_0[1]),.dinb(w_n3811_0[1]),.dout(n3820),.clk(gclk));
	jxor g3763(.dina(w_n3820_0[1]),.dinb(w_n3766_0[1]),.dout(n3821),.clk(gclk));
	jnot g3764(.din(w_n3549_0[1]),.dout(n3822),.clk(gclk));
	jor g3765(.dina(n3822),.dinb(w_n3532_0[0]),.dout(n3823),.clk(gclk));
	jand g3766(.dina(n3823),.dinb(w_n3548_0[1]),.dout(n3824),.clk(gclk));
	jnot g3767(.din(w_n3547_7[0]),.dout(n3825),.clk(gclk));
	jand g3768(.dina(w_n514_0[0]),.dinb(w_n332_1[0]),.dout(n3826),.clk(gclk));
	jand g3769(.dina(w_n1467_0[0]),.dinb(w_n443_0[1]),.dout(n3827),.clk(gclk));
	jand g3770(.dina(n3827),.dinb(w_n3826_0[1]),.dout(n3828),.clk(gclk));
	jand g3771(.dina(w_n232_2[0]),.dinb(w_n213_1[1]),.dout(n3829),.clk(gclk));
	jand g3772(.dina(n3829),.dinb(w_n315_0[2]),.dout(n3830),.clk(gclk));
	jand g3773(.dina(n3830),.dinb(w_n500_0[0]),.dout(n3831),.clk(gclk));
	jand g3774(.dina(n3831),.dinb(w_n1447_0[0]),.dout(n3832),.clk(gclk));
	jand g3775(.dina(n3832),.dinb(n3828),.dout(n3833),.clk(gclk));
	jnot g3776(.din(w_n3833_0[2]),.dout(n3834),.clk(gclk));
	jor g3777(.dina(n3834),.dinb(w_n3825_0[2]),.dout(n3835),.clk(gclk));
	jand g3778(.dina(w_n3543_0[0]),.dinb(w_n3546_0[0]),.dout(n3836),.clk(gclk));
	jxor g3779(.dina(w_n3833_0[1]),.dinb(w_n3836_0[1]),.dout(n3837),.clk(gclk));
	jnot g3780(.din(w_n3837_8[1]),.dout(n3838),.clk(gclk));
	jand g3781(.dina(w_n3838_1[1]),.dinb(w_n3825_0[1]),.dout(n3839),.clk(gclk));
	jnot g3782(.din(w_n3839_0[1]),.dout(n3840),.clk(gclk));
	jand g3783(.dina(w_n3840_0[1]),.dinb(n3835),.dout(n3841),.clk(gclk));
	jxor g3784(.dina(w_n3841_0[2]),.dinb(w_n3824_0[1]),.dout(n3842),.clk(gclk));
	jor g3785(.dina(w_n3842_1[2]),.dinb(w_n3461_4[0]),.dout(n3843),.clk(gclk));
	jor g3786(.dina(w_n3837_8[0]),.dinb(w_n3554_3[1]),.dout(n3844),.clk(gclk));
	jor g3787(.dina(w_n3558_3[0]),.dinb(w_n3547_6[2]),.dout(n3845),.clk(gclk));
	jor g3788(.dina(w_n3552_3[2]),.dinb(w_n3510_7[0]),.dout(n3846),.clk(gclk));
	jand g3789(.dina(n3846),.dinb(n3845),.dout(n3847),.clk(gclk));
	jand g3790(.dina(n3847),.dinb(n3844),.dout(n3848),.clk(gclk));
	jand g3791(.dina(n3848),.dinb(n3843),.dout(n3849),.clk(gclk));
	jxor g3792(.dina(n3849),.dinb(w_n3023_4[2]),.dout(n3850),.clk(gclk));
	jxor g3793(.dina(w_n3850_0[1]),.dinb(w_n3821_0[1]),.dout(n3851),.clk(gclk));
	jxor g3794(.dina(w_n3851_0[2]),.dinb(w_n3763_0[1]),.dout(n3852),.clk(gclk));
	jand g3795(.dina(w_n3852_0[2]),.dinb(w_n325_0[1]),.dout(n3853),.clk(gclk));
	jxor g3796(.dina(w_n3852_0[1]),.dinb(w_n325_0[0]),.dout(n3854),.clk(gclk));
	jand g3797(.dina(w_n344_1[1]),.dinb(w_n152_1[0]),.dout(n3855),.clk(gclk));
	jand g3798(.dina(n3855),.dinb(w_n884_1[0]),.dout(n3856),.clk(gclk));
	jand g3799(.dina(w_n587_1[2]),.dinb(w_n434_0[2]),.dout(n3857),.clk(gclk));
	jand g3800(.dina(n3857),.dinb(w_n446_1[1]),.dout(n3858),.clk(gclk));
	jand g3801(.dina(n3858),.dinb(n3856),.dout(n3859),.clk(gclk));
	jand g3802(.dina(n3859),.dinb(w_n1965_0[0]),.dout(n3860),.clk(gclk));
	jand g3803(.dina(w_n383_1[0]),.dinb(w_n333_1[0]),.dout(n3861),.clk(gclk));
	jand g3804(.dina(n3861),.dinb(w_n241_0[0]),.dout(n3862),.clk(gclk));
	jand g3805(.dina(n3862),.dinb(w_n497_0[2]),.dout(n3863),.clk(gclk));
	jand g3806(.dina(w_n438_0[2]),.dinb(w_n102_1[1]),.dout(n3864),.clk(gclk));
	jand g3807(.dina(n3864),.dinb(w_n600_0[2]),.dout(n3865),.clk(gclk));
	jand g3808(.dina(n3865),.dinb(w_n2377_0[0]),.dout(n3866),.clk(gclk));
	jand g3809(.dina(n3866),.dinb(n3863),.dout(n3867),.clk(gclk));
	jand g3810(.dina(n3867),.dinb(w_n856_0[0]),.dout(n3868),.clk(gclk));
	jand g3811(.dina(w_n1087_0[0]),.dinb(w_n339_2[0]),.dout(n3869),.clk(gclk));
	jand g3812(.dina(n3869),.dinb(w_n361_1[0]),.dout(n3870),.clk(gclk));
	jand g3813(.dina(n3870),.dinb(w_n3868_0[1]),.dout(n3871),.clk(gclk));
	jand g3814(.dina(w_n1072_0[2]),.dinb(w_n166_1[1]),.dout(n3872),.clk(gclk));
	jand g3815(.dina(w_n488_2[0]),.dinb(w_n207_1[0]),.dout(n3873),.clk(gclk));
	jand g3816(.dina(n3873),.dinb(w_n1080_0[0]),.dout(n3874),.clk(gclk));
	jand g3817(.dina(n3874),.dinb(w_n133_0[2]),.dout(n3875),.clk(gclk));
	jand g3818(.dina(w_n3875_0[1]),.dinb(n3872),.dout(n3876),.clk(gclk));
	jand g3819(.dina(w_n510_1[1]),.dinb(w_n384_1[1]),.dout(n3877),.clk(gclk));
	jand g3820(.dina(n3877),.dinb(w_n161_0[0]),.dout(n3878),.clk(gclk));
	jand g3821(.dina(n3878),.dinb(w_n120_0[2]),.dout(n3879),.clk(gclk));
	jand g3822(.dina(n3879),.dinb(w_n3489_0[0]),.dout(n3880),.clk(gclk));
	jand g3823(.dina(n3880),.dinb(n3876),.dout(n3881),.clk(gclk));
	jand g3824(.dina(w_n387_1[1]),.dinb(w_n331_1[0]),.dout(n3882),.clk(gclk));
	jand g3825(.dina(n3882),.dinb(w_n124_1[0]),.dout(n3883),.clk(gclk));
	jand g3826(.dina(n3883),.dinb(w_n94_1[0]),.dout(n3884),.clk(gclk));
	jand g3827(.dina(n3884),.dinb(w_n3881_0[1]),.dout(n3885),.clk(gclk));
	jand g3828(.dina(n3885),.dinb(w_n3871_0[1]),.dout(n3886),.clk(gclk));
	jand g3829(.dina(n3886),.dinb(n3860),.dout(n3887),.clk(gclk));
	jand g3830(.dina(w_n2613_0[0]),.dinb(w_n1332_0[0]),.dout(n3888),.clk(gclk));
	jand g3831(.dina(w_n1460_0[2]),.dinb(w_n173_0[1]),.dout(n3889),.clk(gclk));
	jand g3832(.dina(n3889),.dinb(w_n2142_0[0]),.dout(n3890),.clk(gclk));
	jand g3833(.dina(n3890),.dinb(w_n435_1[0]),.dout(n3891),.clk(gclk));
	jand g3834(.dina(n3891),.dinb(n3888),.dout(n3892),.clk(gclk));
	jand g3835(.dina(w_n152_0[2]),.dinb(w_n136_1[0]),.dout(n3893),.clk(gclk));
	jand g3836(.dina(n3893),.dinb(w_n3185_0[0]),.dout(n3894),.clk(gclk));
	jand g3837(.dina(n3894),.dinb(w_n1078_0[0]),.dout(n3895),.clk(gclk));
	jand g3838(.dina(w_n252_2[1]),.dinb(w_n142_1[0]),.dout(n3896),.clk(gclk));
	jand g3839(.dina(w_n535_1[1]),.dinb(w_n283_0[2]),.dout(n3897),.clk(gclk));
	jand g3840(.dina(w_n347_0[2]),.dinb(w_n232_1[2]),.dout(n3898),.clk(gclk));
	jand g3841(.dina(n3898),.dinb(n3897),.dout(n3899),.clk(gclk));
	jand g3842(.dina(n3899),.dinb(n3896),.dout(n3900),.clk(gclk));
	jand g3843(.dina(w_n463_0[0]),.dinb(w_n382_0[2]),.dout(n3901),.clk(gclk));
	jand g3844(.dina(n3901),.dinb(w_n1366_0[1]),.dout(n3902),.clk(gclk));
	jand g3845(.dina(n3902),.dinb(w_n1961_0[0]),.dout(n3903),.clk(gclk));
	jand g3846(.dina(n3903),.dinb(w_n2155_1[0]),.dout(n3904),.clk(gclk));
	jand g3847(.dina(n3904),.dinb(n3900),.dout(n3905),.clk(gclk));
	jand g3848(.dina(n3905),.dinb(w_n3895_0[1]),.dout(n3906),.clk(gclk));
	jand g3849(.dina(n3906),.dinb(w_n3892_0[2]),.dout(n3907),.clk(gclk));
	jand g3850(.dina(n3907),.dinb(w_n2409_0[0]),.dout(n3908),.clk(gclk));
	jnot g3851(.din(n3908),.dout(n3909),.clk(gclk));
	jnot g3852(.din(w_n3576_0[0]),.dout(n3910),.clk(gclk));
	jnot g3853(.din(w_n3588_0[0]),.dout(n3911),.clk(gclk));
	jnot g3854(.din(w_n3589_0[0]),.dout(n3912),.clk(gclk));
	jnot g3855(.din(w_n3599_0[0]),.dout(n3913),.clk(gclk));
	jnot g3856(.din(w_n3600_0[0]),.dout(n3914),.clk(gclk));
	jnot g3857(.din(w_n3610_0[0]),.dout(n3915),.clk(gclk));
	jnot g3858(.din(w_n3611_0[0]),.dout(n3916),.clk(gclk));
	jnot g3859(.din(w_n3621_0[0]),.dout(n3917),.clk(gclk));
	jnot g3860(.din(w_n3622_0[0]),.dout(n3918),.clk(gclk));
	jnot g3861(.din(w_n3632_0[0]),.dout(n3919),.clk(gclk));
	jnot g3862(.din(w_n3633_0[0]),.dout(n3920),.clk(gclk));
	jnot g3863(.din(w_n3643_0[0]),.dout(n3921),.clk(gclk));
	jnot g3864(.din(w_n3644_0[0]),.dout(n3922),.clk(gclk));
	jnot g3865(.din(w_n3654_0[0]),.dout(n3923),.clk(gclk));
	jnot g3866(.din(w_n3655_0[0]),.dout(n3924),.clk(gclk));
	jnot g3867(.din(w_n3665_0[0]),.dout(n3925),.clk(gclk));
	jnot g3868(.din(w_n3734_0[0]),.dout(n3926),.clk(gclk));
	jnot g3869(.din(w_n3702_0[0]),.dout(n3927),.clk(gclk));
	jnot g3870(.din(w_n3676_0[0]),.dout(n3928),.clk(gclk));
	jand g3871(.dina(w_n3688_0[0]),.dinb(w_n3695_0[0]),.dout(n3929),.clk(gclk));
	jand g3872(.dina(w_n3685_0[0]),.dinb(w_n3455_4[1]),.dout(n3930),.clk(gclk));
	jor g3873(.dina(n3930),.dinb(n3929),.dout(n3931),.clk(gclk));
	jor g3874(.dina(n3931),.dinb(n3928),.dout(n3932),.clk(gclk));
	jand g3875(.dina(w_n3700_0[0]),.dinb(n3932),.dout(n3933),.clk(gclk));
	jand g3876(.dina(w_n3718_0[0]),.dinb(w_n3455_4[0]),.dout(n3934),.clk(gclk));
	jand g3877(.dina(w_n3720_0[0]),.dinb(w_n3709_0[0]),.dout(n3935),.clk(gclk));
	jor g3878(.dina(n3935),.dinb(n3934),.dout(n3936),.clk(gclk));
	jor g3879(.dina(n3936),.dinb(n3933),.dout(n3937),.clk(gclk));
	jand g3880(.dina(n3937),.dinb(n3927),.dout(n3938),.clk(gclk));
	jnot g3881(.din(w_n3733_0[0]),.dout(n3939),.clk(gclk));
	jor g3882(.dina(n3939),.dinb(n3938),.dout(n3940),.clk(gclk));
	jand g3883(.dina(w_n3738_0[0]),.dinb(n3940),.dout(n3941),.clk(gclk));
	jor g3884(.dina(n3941),.dinb(n3926),.dout(n3942),.clk(gclk));
	jnot g3885(.din(w_n3742_0[0]),.dout(n3943),.clk(gclk));
	jand g3886(.dina(n3943),.dinb(n3942),.dout(n3944),.clk(gclk));
	jor g3887(.dina(n3944),.dinb(n3925),.dout(n3945),.clk(gclk));
	jand g3888(.dina(n3945),.dinb(n3924),.dout(n3946),.clk(gclk));
	jor g3889(.dina(n3946),.dinb(n3923),.dout(n3947),.clk(gclk));
	jand g3890(.dina(n3947),.dinb(n3922),.dout(n3948),.clk(gclk));
	jor g3891(.dina(n3948),.dinb(n3921),.dout(n3949),.clk(gclk));
	jand g3892(.dina(n3949),.dinb(n3920),.dout(n3950),.clk(gclk));
	jor g3893(.dina(n3950),.dinb(n3919),.dout(n3951),.clk(gclk));
	jand g3894(.dina(n3951),.dinb(n3918),.dout(n3952),.clk(gclk));
	jor g3895(.dina(n3952),.dinb(n3917),.dout(n3953),.clk(gclk));
	jand g3896(.dina(n3953),.dinb(n3916),.dout(n3954),.clk(gclk));
	jor g3897(.dina(n3954),.dinb(n3915),.dout(n3955),.clk(gclk));
	jand g3898(.dina(n3955),.dinb(n3914),.dout(n3956),.clk(gclk));
	jor g3899(.dina(n3956),.dinb(n3913),.dout(n3957),.clk(gclk));
	jor g3900(.dina(n3957),.dinb(n3912),.dout(n3958),.clk(gclk));
	jand g3901(.dina(n3958),.dinb(n3911),.dout(n3959),.clk(gclk));
	jxor g3902(.dina(w_n3959_0[1]),.dinb(w_n3910_0[1]),.dout(n3960),.clk(gclk));
	jand g3903(.dina(n3960),.dinb(n3909),.dout(n3961),.clk(gclk));
	jnot g3904(.din(w_n3961_0[1]),.dout(n3962),.clk(gclk));
	jand g3905(.dina(n3962),.dinb(w_n3887_0[1]),.dout(n3963),.clk(gclk));
	jnot g3906(.din(w_n3963_0[1]),.dout(n3964),.clk(gclk));
	jnot g3907(.din(w_n3887_0[0]),.dout(n3965),.clk(gclk));
	jand g3908(.dina(w_n3961_0[0]),.dinb(n3965),.dout(n3966),.clk(gclk));
	jxor g3909(.dina(w_n3761_0[1]),.dinb(w_n3760_0[0]),.dout(n3967),.clk(gclk));
	jor g3910(.dina(n3967),.dinb(n3966),.dout(n3968),.clk(gclk));
	jand g3911(.dina(w_n3968_0[1]),.dinb(n3964),.dout(n3969),.clk(gclk));
	jand g3912(.dina(w_n3969_0[1]),.dinb(w_n3854_0[1]),.dout(n3970),.clk(gclk));
	jor g3913(.dina(n3970),.dinb(w_n3853_0[1]),.dout(n3971),.clk(gclk));
	jand g3914(.dina(w_n3850_0[0]),.dinb(w_n3821_0[0]),.dout(n3972),.clk(gclk));
	jnot g3915(.din(w_n3972_0[1]),.dout(n3973),.clk(gclk));
	jnot g3916(.din(w_n3575_0[0]),.dout(n3974),.clk(gclk));
	jor g3917(.dina(w_n3959_0[0]),.dinb(w_n3910_0[0]),.dout(n3975),.clk(gclk));
	jand g3918(.dina(n3975),.dinb(n3974),.dout(n3976),.clk(gclk));
	jnot g3919(.din(w_n3761_0[0]),.dout(n3977),.clk(gclk));
	jor g3920(.dina(n3977),.dinb(n3976),.dout(n3978),.clk(gclk));
	jand g3921(.dina(n3978),.dinb(w_n3563_0[0]),.dout(n3979),.clk(gclk));
	jnot g3922(.din(w_n3851_0[1]),.dout(n3980),.clk(gclk));
	jor g3923(.dina(n3980),.dinb(n3979),.dout(n3981),.clk(gclk));
	jand g3924(.dina(n3981),.dinb(n3973),.dout(n3982),.clk(gclk));
	jand g3925(.dina(w_n3819_0[0]),.dinb(w_n3811_0[0]),.dout(n3983),.clk(gclk));
	jand g3926(.dina(w_n3820_0[0]),.dinb(w_n3766_0[0]),.dout(n3984),.clk(gclk));
	jor g3927(.dina(n3984),.dinb(n3983),.dout(n3985),.clk(gclk));
	jor g3928(.dina(w_n3809_0[0]),.dinb(w_n3801_0[0]),.dout(n3986),.clk(gclk));
	jnot g3929(.din(n3986),.dout(n3987),.clk(gclk));
	jand g3930(.dina(w_n3810_0[0]),.dinb(w_n3770_0[0]),.dout(n3988),.clk(gclk));
	jor g3931(.dina(n3988),.dinb(n3987),.dout(n3989),.clk(gclk));
	jand g3932(.dina(w_n3798_0[0]),.dinb(w_n3790_0[0]),.dout(n3990),.clk(gclk));
	jand g3933(.dina(w_n3799_0[0]),.dinb(w_n3773_0[0]),.dout(n3991),.clk(gclk));
	jor g3934(.dina(n3991),.dinb(n3990),.dout(n3992),.clk(gclk));
	jor g3935(.dina(w_n3789_0[0]),.dinb(w_n3780_0[0]),.dout(n3993),.clk(gclk));
	jnot g3936(.din(w_n3787_0[0]),.dout(n3994),.clk(gclk));
	jand g3937(.dina(n3994),.dinb(w_n1438_15[2]),.dout(n3995),.clk(gclk));
	jand g3938(.dina(n3995),.dinb(w_n2094_2[0]),.dout(n3996),.clk(gclk));
	jnot g3939(.din(n3996),.dout(n3997),.clk(gclk));
	jand g3940(.dina(n3997),.dinb(n3993),.dout(n3998),.clk(gclk));
	jor g3941(.dina(w_n2836_0[1]),.dinb(w_n3384_7[0]),.dout(n3999),.clk(gclk));
	jand g3942(.dina(w_n2684_2[0]),.dinb(w_n2491_2[1]),.dout(n4000),.clk(gclk));
	jand g3943(.dina(w_n2488_2[1]),.dinb(w_n2687_1[2]),.dout(n4001),.clk(gclk));
	jand g3944(.dina(w_n2923_2[2]),.dinb(w_n2690_1[0]),.dout(n4002),.clk(gclk));
	jor g3945(.dina(n4002),.dinb(n4001),.dout(n4003),.clk(gclk));
	jor g3946(.dina(n4003),.dinb(n4000),.dout(n4004),.clk(gclk));
	jnot g3947(.din(n4004),.dout(n4005),.clk(gclk));
	jand g3948(.dina(n4005),.dinb(n3999),.dout(n4006),.clk(gclk));
	jand g3949(.dina(w_n2256_1[2]),.dinb(w_n1438_15[1]),.dout(n4007),.clk(gclk));
	jxor g3950(.dina(n4007),.dinb(w_n4006_0[1]),.dout(n4008),.clk(gclk));
	jxor g3951(.dina(w_n4008_0[1]),.dinb(w_n3998_0[1]),.dout(n4009),.clk(gclk));
	jor g3952(.dina(w_n3010_0[2]),.dinb(w_n2252_6[0]),.dout(n4010),.clk(gclk));
	jor g3953(.dina(w_n2800_3[0]),.dinb(w_n2359_6[0]),.dout(n4011),.clk(gclk));
	jor g3954(.dina(w_n3008_3[2]),.dinb(w_n2355_5[2]),.dout(n4012),.clk(gclk));
	jor g3955(.dina(w_n2707_2[1]),.dinb(w_n2357_6[0]),.dout(n4013),.clk(gclk));
	jand g3956(.dina(n4013),.dinb(n4012),.dout(n4014),.clk(gclk));
	jand g3957(.dina(n4014),.dinb(n4011),.dout(n4015),.clk(gclk));
	jand g3958(.dina(n4015),.dinb(n4010),.dout(n4016),.clk(gclk));
	jxor g3959(.dina(n4016),.dinb(w_n1480_5[2]),.dout(n4017),.clk(gclk));
	jxor g3960(.dina(w_n4017_0[1]),.dinb(w_n4009_0[1]),.dout(n4018),.clk(gclk));
	jxor g3961(.dina(w_n4018_0[1]),.dinb(w_n3992_0[1]),.dout(n4019),.clk(gclk));
	jnot g3962(.din(n4019),.dout(n4020),.clk(gclk));
	jor g3963(.dina(w_n3205_1[0]),.dinb(w_n2506_5[0]),.dout(n4021),.clk(gclk));
	jor g3964(.dina(w_n3166_5[1]),.dinb(w_n2807_5[0]),.dout(n4022),.clk(gclk));
	jor g3965(.dina(w_n3203_5[1]),.dinb(w_n2810_4[2]),.dout(n4023),.clk(gclk));
	jand g3966(.dina(n4023),.dinb(n4022),.dout(n4024),.clk(gclk));
	jor g3967(.dina(w_n3216_4[1]),.dinb(w_n2816_5[0]),.dout(n4025),.clk(gclk));
	jand g3968(.dina(n4025),.dinb(n4024),.dout(n4026),.clk(gclk));
	jand g3969(.dina(n4026),.dinb(n4021),.dout(n4027),.clk(gclk));
	jxor g3970(.dina(n4027),.dinb(w_n1257_6[0]),.dout(n4028),.clk(gclk));
	jxor g3971(.dina(w_n4028_0[1]),.dinb(w_n4020_0[1]),.dout(n4029),.clk(gclk));
	jxor g3972(.dina(w_n4029_0[1]),.dinb(w_n3989_0[1]),.dout(n4030),.clk(gclk));
	jor g3973(.dina(w_n3566_1[1]),.dinb(w_n3029_4[0]),.dout(n4031),.clk(gclk));
	jor g3974(.dina(w_n3510_6[2]),.dinb(w_n3213_3[2]),.dout(n4032),.clk(gclk));
	jor g3975(.dina(w_n3495_6[0]),.dinb(w_n3210_4[0]),.dout(n4033),.clk(gclk));
	jor g3976(.dina(w_n3441_5[0]),.dinb(w_n3219_4[0]),.dout(n4034),.clk(gclk));
	jand g3977(.dina(n4034),.dinb(n4033),.dout(n4035),.clk(gclk));
	jand g3978(.dina(n4035),.dinb(n4032),.dout(n4036),.clk(gclk));
	jand g3979(.dina(n4036),.dinb(n4031),.dout(n4037),.clk(gclk));
	jxor g3980(.dina(n4037),.dinb(w_n1156_5[2]),.dout(n4038),.clk(gclk));
	jxor g3981(.dina(w_n4038_0[1]),.dinb(w_n4030_0[1]),.dout(n4039),.clk(gclk));
	jxor g3982(.dina(w_n4039_0[1]),.dinb(w_n3985_0[1]),.dout(n4040),.clk(gclk));
	jnot g3983(.din(w_n3841_0[1]),.dout(n4041),.clk(gclk));
	jor g3984(.dina(n4041),.dinb(w_n3824_0[0]),.dout(n4042),.clk(gclk));
	jand g3985(.dina(n4042),.dinb(w_n3840_0[0]),.dout(n4043),.clk(gclk));
	jand g3986(.dina(w_n2954_0[0]),.dinb(w_n1133_0[0]),.dout(n4044),.clk(gclk));
	jand g3987(.dina(n4044),.dinb(w_n3177_0[0]),.dout(n4045),.clk(gclk));
	jand g3988(.dina(w_n404_0[1]),.dinb(w_n182_2[1]),.dout(n4046),.clk(gclk));
	jand g3989(.dina(n4046),.dinb(w_n1127_0[0]),.dout(n4047),.clk(gclk));
	jand g3990(.dina(n4047),.dinb(w_n448_0[2]),.dout(n4048),.clk(gclk));
	jand g3991(.dina(w_n385_0[0]),.dinb(w_n251_0[1]),.dout(n4049),.clk(gclk));
	jand g3992(.dina(n4049),.dinb(w_n321_1[0]),.dout(n4050),.clk(gclk));
	jand g3993(.dina(n4050),.dinb(n4048),.dout(n4051),.clk(gclk));
	jand g3994(.dina(w_n4051_0[1]),.dinb(n4045),.dout(n4052),.clk(gclk));
	jand g3995(.dina(w_n2127_0[2]),.dinb(w_n482_0[0]),.dout(n4053),.clk(gclk));
	jand g3996(.dina(n4053),.dinb(w_n252_2[0]),.dout(n4054),.clk(gclk));
	jand g3997(.dina(n4054),.dinb(w_n1023_0[0]),.dout(n4055),.clk(gclk));
	jand g3998(.dina(w_n233_0[2]),.dinb(w_n176_0[2]),.dout(n4056),.clk(gclk));
	jand g3999(.dina(n4056),.dinb(n4055),.dout(n4057),.clk(gclk));
	jand g4000(.dina(n4057),.dinb(n4052),.dout(n4058),.clk(gclk));
	jand g4001(.dina(n4058),.dinb(w_n834_0[0]),.dout(n4059),.clk(gclk));
	jand g4002(.dina(w_n4059_0[2]),.dinb(w_n3837_7[2]),.dout(n4060),.clk(gclk));
	jnot g4003(.din(n4060),.dout(n4061),.clk(gclk));
	jand g4004(.dina(w_n3833_0[0]),.dinb(w_n3836_0[0]),.dout(n4062),.clk(gclk));
	jxor g4005(.dina(w_n4059_0[1]),.dinb(w_n4062_0[1]),.dout(n4063),.clk(gclk));
	jor g4006(.dina(w_n4063_8[1]),.dinb(w_n3837_7[1]),.dout(n4064),.clk(gclk));
	jand g4007(.dina(w_n4064_0[2]),.dinb(n4061),.dout(n4065),.clk(gclk));
	jxor g4008(.dina(w_n4065_0[2]),.dinb(w_n4043_0[1]),.dout(n4066),.clk(gclk));
	jor g4009(.dina(w_n4066_1[2]),.dinb(w_n3461_3[2]),.dout(n4067),.clk(gclk));
	jor g4010(.dina(w_n3552_3[1]),.dinb(w_n3547_6[1]),.dout(n4068),.clk(gclk));
	jor g4011(.dina(w_n3837_7[0]),.dinb(w_n3558_2[2]),.dout(n4069),.clk(gclk));
	jor g4012(.dina(w_n4063_8[0]),.dinb(w_n3554_3[0]),.dout(n4070),.clk(gclk));
	jand g4013(.dina(n4070),.dinb(n4069),.dout(n4071),.clk(gclk));
	jand g4014(.dina(n4071),.dinb(n4068),.dout(n4072),.clk(gclk));
	jand g4015(.dina(n4072),.dinb(n4067),.dout(n4073),.clk(gclk));
	jxor g4016(.dina(n4073),.dinb(w_n3023_4[1]),.dout(n4074),.clk(gclk));
	jxor g4017(.dina(w_n4074_0[1]),.dinb(w_n4040_0[1]),.dout(n4075),.clk(gclk));
	jxor g4018(.dina(w_n4075_1[1]),.dinb(w_n3982_0[1]),.dout(n4076),.clk(gclk));
	jnot g4019(.din(w_n190_1[0]),.dout(n4077),.clk(gclk));
	jor g4020(.dina(w_n1319_0[0]),.dinb(n4077),.dout(n4078),.clk(gclk));
	jor g4021(.dina(n4078),.dinb(w_n628_0[0]),.dout(n4079),.clk(gclk));
	jnot g4022(.din(n4079),.dout(n4080),.clk(gclk));
	jand g4023(.dina(n4080),.dinb(w_n1392_0[0]),.dout(n4081),.clk(gclk));
	jand g4024(.dina(w_n1072_0[1]),.dinb(w_n251_0[0]),.dout(n4082),.clk(gclk));
	jand g4025(.dina(n4082),.dinb(w_n128_1[1]),.dout(n4083),.clk(gclk));
	jand g4026(.dina(w_n825_0[1]),.dinb(w_n102_1[0]),.dout(n4084),.clk(gclk));
	jand g4027(.dina(n4084),.dinb(n4083),.dout(n4085),.clk(gclk));
	jand g4028(.dina(n4085),.dinb(n4081),.dout(n4086),.clk(gclk));
	jand g4029(.dina(w_n2631_0[0]),.dinb(w_n1069_0[0]),.dout(n4087),.clk(gclk));
	jand g4030(.dina(n4087),.dinb(n4086),.dout(n4088),.clk(gclk));
	jxor g4031(.dina(w_n4088_0[2]),.dinb(w_n4076_0[1]),.dout(n4089),.clk(gclk));
	jxor g4032(.dina(w_n4089_0[1]),.dinb(w_n3971_0[1]),.dout(n4090),.clk(gclk));
	jxor g4033(.dina(w_n3969_0[0]),.dinb(w_n3854_0[0]),.dout(n4091),.clk(gclk));
	jxor g4034(.dina(w_n4091_0[1]),.dinb(w_n4090_0[1]),.dout(sin0_fa_),.clk(gclk));
	jxor g4035(.dina(a23),.dinb(w_a22_0[0]),.dout(n4093),.clk(gclk));
	jand g4036(.dina(w_n4093_11[1]),.dinb(w_sin0_0[1]),.dout(n4094),.clk(gclk));
	jnot g4037(.din(w_n4094_0[1]),.dout(n4095),.clk(gclk));
	jand g4038(.dina(w_n4091_0[0]),.dinb(w_n4090_0[0]),.dout(n4096),.clk(gclk));
	jor g4039(.dina(w_n4088_0[1]),.dinb(w_n4076_0[0]),.dout(n4097),.clk(gclk));
	jnot g4040(.din(w_n4097_0[1]),.dout(n4098),.clk(gclk));
	jand g4041(.dina(w_n4089_0[0]),.dinb(w_n3971_0[0]),.dout(n4099),.clk(gclk));
	jor g4042(.dina(n4099),.dinb(n4098),.dout(n4100),.clk(gclk));
	jand g4043(.dina(w_n4074_0[0]),.dinb(w_n4040_0[0]),.dout(n4101),.clk(gclk));
	jnot g4044(.din(w_n4101_0[1]),.dout(n4102),.clk(gclk));
	jnot g4045(.din(w_n4075_1[0]),.dout(n4103),.clk(gclk));
	jor g4046(.dina(n4103),.dinb(w_n3982_0[0]),.dout(n4104),.clk(gclk));
	jand g4047(.dina(n4104),.dinb(n4102),.dout(n4105),.clk(gclk));
	jand g4048(.dina(w_n4038_0[0]),.dinb(w_n4030_0[0]),.dout(n4106),.clk(gclk));
	jand g4049(.dina(w_n4039_0[0]),.dinb(w_n3985_0[0]),.dout(n4107),.clk(gclk));
	jor g4050(.dina(n4107),.dinb(n4106),.dout(n4108),.clk(gclk));
	jor g4051(.dina(w_n4028_0[0]),.dinb(w_n4020_0[0]),.dout(n4109),.clk(gclk));
	jnot g4052(.din(n4109),.dout(n4110),.clk(gclk));
	jand g4053(.dina(w_n4029_0[0]),.dinb(w_n3989_0[0]),.dout(n4111),.clk(gclk));
	jor g4054(.dina(n4111),.dinb(n4110),.dout(n4112),.clk(gclk));
	jand g4055(.dina(w_n4017_0[0]),.dinb(w_n4009_0[0]),.dout(n4113),.clk(gclk));
	jand g4056(.dina(w_n4018_0[0]),.dinb(w_n3992_0[0]),.dout(n4114),.clk(gclk));
	jor g4057(.dina(n4114),.dinb(n4113),.dout(n4115),.clk(gclk));
	jor g4058(.dina(w_n4008_0[0]),.dinb(w_n3998_0[0]),.dout(n4116),.clk(gclk));
	jand g4059(.dina(w_n4006_0[0]),.dinb(w_n1438_15[0]),.dout(n4117),.clk(gclk));
	jand g4060(.dina(n4117),.dinb(w_n2236_1[2]),.dout(n4118),.clk(gclk));
	jnot g4061(.din(n4118),.dout(n4119),.clk(gclk));
	jand g4062(.dina(n4119),.dinb(n4116),.dout(n4120),.clk(gclk));
	jor g4063(.dina(w_n2825_0[1]),.dinb(w_n3384_6[2]),.dout(n4121),.clk(gclk));
	jand g4064(.dina(w_n2684_1[2]),.dinb(w_n2488_2[0]),.dout(n4122),.clk(gclk));
	jand g4065(.dina(w_n2683_1[2]),.dinb(w_n2491_2[0]),.dout(n4123),.clk(gclk));
	jand g4066(.dina(w_n2923_2[1]),.dinb(w_n2687_1[1]),.dout(n4124),.clk(gclk));
	jor g4067(.dina(n4124),.dinb(n4123),.dout(n4125),.clk(gclk));
	jor g4068(.dina(n4125),.dinb(n4122),.dout(n4126),.clk(gclk));
	jnot g4069(.din(n4126),.dout(n4127),.clk(gclk));
	jand g4070(.dina(n4127),.dinb(n4121),.dout(n4128),.clk(gclk));
	jand g4071(.dina(w_n2351_2[2]),.dinb(w_n1438_14[2]),.dout(n4129),.clk(gclk));
	jxor g4072(.dina(n4129),.dinb(w_n4128_0[1]),.dout(n4130),.clk(gclk));
	jxor g4073(.dina(w_n4130_0[1]),.dinb(w_n4120_0[1]),.dout(n4131),.clk(gclk));
	jnot g4074(.din(n4131),.dout(n4132),.clk(gclk));
	jor g4075(.dina(w_n3242_0[2]),.dinb(w_n2252_5[2]),.dout(n4133),.clk(gclk));
	jor g4076(.dina(w_n3008_3[1]),.dinb(w_n2359_5[2]),.dout(n4134),.clk(gclk));
	jor g4077(.dina(w_n3216_4[0]),.dinb(w_n2355_5[1]),.dout(n4135),.clk(gclk));
	jand g4078(.dina(n4135),.dinb(n4134),.dout(n4136),.clk(gclk));
	jor g4079(.dina(w_n2800_2[2]),.dinb(w_n2357_5[2]),.dout(n4137),.clk(gclk));
	jand g4080(.dina(n4137),.dinb(n4136),.dout(n4138),.clk(gclk));
	jand g4081(.dina(n4138),.dinb(n4133),.dout(n4139),.clk(gclk));
	jxor g4082(.dina(n4139),.dinb(w_n1356_6[0]),.dout(n4140),.clk(gclk));
	jxor g4083(.dina(w_n4140_0[1]),.dinb(w_n4132_0[1]),.dout(n4141),.clk(gclk));
	jxor g4084(.dina(w_n4141_0[1]),.dinb(w_n4115_0[1]),.dout(n4142),.clk(gclk));
	jnot g4085(.din(n4142),.dout(n4143),.clk(gclk));
	jor g4086(.dina(w_n3443_1[0]),.dinb(w_n2506_4[2]),.dout(n4144),.clk(gclk));
	jor g4087(.dina(w_n3441_4[2]),.dinb(w_n2810_4[1]),.dout(n4145),.clk(gclk));
	jor g4088(.dina(w_n3203_5[0]),.dinb(w_n2807_4[2]),.dout(n4146),.clk(gclk));
	jand g4089(.dina(n4146),.dinb(n4145),.dout(n4147),.clk(gclk));
	jor g4090(.dina(w_n3166_5[0]),.dinb(w_n2816_4[2]),.dout(n4148),.clk(gclk));
	jand g4091(.dina(n4148),.dinb(n4147),.dout(n4149),.clk(gclk));
	jand g4092(.dina(n4149),.dinb(n4144),.dout(n4150),.clk(gclk));
	jxor g4093(.dina(n4150),.dinb(w_n1257_5[2]),.dout(n4151),.clk(gclk));
	jxor g4094(.dina(w_n4151_0[1]),.dinb(w_n4143_0[1]),.dout(n4152),.clk(gclk));
	jxor g4095(.dina(w_n4152_0[1]),.dinb(w_n4112_0[1]),.dout(n4153),.clk(gclk));
	jor g4096(.dina(w_n3550_1[1]),.dinb(w_n3029_3[2]),.dout(n4154),.clk(gclk));
	jor g4097(.dina(w_n3547_6[0]),.dinb(w_n3213_3[1]),.dout(n4155),.clk(gclk));
	jor g4098(.dina(w_n3510_6[1]),.dinb(w_n3210_3[2]),.dout(n4156),.clk(gclk));
	jor g4099(.dina(w_n3495_5[2]),.dinb(w_n3219_3[2]),.dout(n4157),.clk(gclk));
	jand g4100(.dina(n4157),.dinb(n4156),.dout(n4158),.clk(gclk));
	jand g4101(.dina(n4158),.dinb(n4155),.dout(n4159),.clk(gclk));
	jand g4102(.dina(n4159),.dinb(n4154),.dout(n4160),.clk(gclk));
	jxor g4103(.dina(n4160),.dinb(w_n1156_5[1]),.dout(n4161),.clk(gclk));
	jxor g4104(.dina(w_n4161_0[1]),.dinb(w_n4153_0[1]),.dout(n4162),.clk(gclk));
	jxor g4105(.dina(w_n4162_0[1]),.dinb(w_n4108_0[1]),.dout(n4163),.clk(gclk));
	jnot g4106(.din(w_n4064_0[1]),.dout(n4164),.clk(gclk));
	jnot g4107(.din(w_n3548_0[0]),.dout(n4165),.clk(gclk));
	jnot g4108(.din(w_n3511_0[0]),.dout(n4166),.clk(gclk));
	jand g4109(.dina(w_n2472_0[0]),.dinb(w_n3713_0[0]),.dout(n4167),.clk(gclk));
	jor g4110(.dina(n4167),.dinb(w_n2691_0[0]),.dout(n4168),.clk(gclk));
	jand g4111(.dina(w_n2835_0[0]),.dinb(n4168),.dout(n4169),.clk(gclk));
	jor g4112(.dina(n4169),.dinb(w_n2688_0[0]),.dout(n4170),.clk(gclk));
	jand g4113(.dina(w_n2824_0[0]),.dinb(n4170),.dout(n4171),.clk(gclk));
	jor g4114(.dina(n4171),.dinb(w_n2685_0[0]),.dout(n4172),.clk(gclk));
	jand g4115(.dina(w_n2801_0[0]),.dinb(n4172),.dout(n4173),.clk(gclk));
	jor g4116(.dina(n4173),.dinb(w_n2944_0[0]),.dout(n4174),.clk(gclk));
	jand g4117(.dina(w_n3009_0[0]),.dinb(n4174),.dout(n4175),.clk(gclk));
	jor g4118(.dina(n4175),.dinb(w_n3150_0[0]),.dout(n4176),.clk(gclk));
	jand g4119(.dina(w_n3241_0[0]),.dinb(n4176),.dout(n4177),.clk(gclk));
	jor g4120(.dina(n4177),.dinb(w_n3148_0[0]),.dout(n4178),.clk(gclk));
	jand g4121(.dina(w_n3228_0[0]),.dinb(n4178),.dout(n4179),.clk(gclk));
	jor g4122(.dina(n4179),.dinb(w_n3145_0[0]),.dout(n4180),.clk(gclk));
	jand g4123(.dina(w_n3204_0[0]),.dinb(n4180),.dout(n4181),.clk(gclk));
	jor g4124(.dina(n4181),.dinb(w_n3416_0[0]),.dout(n4182),.clk(gclk));
	jand g4125(.dina(w_n3442_0[0]),.dinb(n4182),.dout(n4183),.clk(gclk));
	jor g4126(.dina(n4183),.dinb(w_n3514_0[0]),.dout(n4184),.clk(gclk));
	jand g4127(.dina(w_n3578_0[0]),.dinb(n4184),.dout(n4185),.clk(gclk));
	jor g4128(.dina(n4185),.dinb(w_n3521_0[0]),.dout(n4186),.clk(gclk));
	jand g4129(.dina(w_n3529_0[0]),.dinb(n4186),.dout(n4187),.clk(gclk));
	jor g4130(.dina(n4187),.dinb(n4166),.dout(n4188),.clk(gclk));
	jand g4131(.dina(w_n3549_0[0]),.dinb(n4188),.dout(n4189),.clk(gclk));
	jor g4132(.dina(n4189),.dinb(n4165),.dout(n4190),.clk(gclk));
	jand g4133(.dina(w_n3841_0[0]),.dinb(n4190),.dout(n4191),.clk(gclk));
	jor g4134(.dina(n4191),.dinb(w_n3839_0[0]),.dout(n4192),.clk(gclk));
	jand g4135(.dina(w_n4065_0[1]),.dinb(n4192),.dout(n4193),.clk(gclk));
	jor g4136(.dina(n4193),.dinb(n4164),.dout(n4194),.clk(gclk));
	jnot g4137(.din(w_n4062_0[0]),.dout(n4195),.clk(gclk));
	jnot g4138(.din(w_n4059_0[0]),.dout(n4196),.clk(gclk));
	jand g4139(.dina(n4196),.dinb(n4195),.dout(n4197),.clk(gclk));
	jand g4140(.dina(w_n2155_0[2]),.dinb(w_n340_0[2]),.dout(n4198),.clk(gclk));
	jand g4141(.dina(w_n310_0[2]),.dinb(w_n114_1[1]),.dout(n4199),.clk(gclk));
	jand g4142(.dina(n4199),.dinb(w_n277_0[0]),.dout(n4200),.clk(gclk));
	jand g4143(.dina(n4200),.dinb(w_n246_0[0]),.dout(n4201),.clk(gclk));
	jand g4144(.dina(n4201),.dinb(w_n477_0[0]),.dout(n4202),.clk(gclk));
	jand g4145(.dina(n4202),.dinb(n4198),.dout(n4203),.clk(gclk));
	jand g4146(.dina(w_n4203_0[1]),.dinb(w_n1079_0[0]),.dout(n4204),.clk(gclk));
	jand g4147(.dina(n4204),.dinb(w_n1339_0[0]),.dout(n4205),.clk(gclk));
	jand g4148(.dina(w_n3497_0[1]),.dinb(w_n439_1[1]),.dout(n4206),.clk(gclk));
	jand g4149(.dina(n4206),.dinb(w_n333_0[2]),.dout(n4207),.clk(gclk));
	jand g4150(.dina(w_n389_1[1]),.dinb(w_n338_0[0]),.dout(n4208),.clk(gclk));
	jand g4151(.dina(w_n540_0[1]),.dinb(w_n446_1[0]),.dout(n4209),.clk(gclk));
	jand g4152(.dina(n4209),.dinb(n4208),.dout(n4210),.clk(gclk));
	jand g4153(.dina(n4210),.dinb(n4207),.dout(n4211),.clk(gclk));
	jand g4154(.dina(n4211),.dinb(w_n2146_0[1]),.dout(n4212),.clk(gclk));
	jand g4155(.dina(n4212),.dinb(n4205),.dout(n4213),.clk(gclk));
	jxor g4156(.dina(w_n4213_6[2]),.dinb(n4197),.dout(n4214),.clk(gclk));
	jxor g4157(.dina(w_n4214_0[2]),.dinb(w_n4194_0[1]),.dout(n4215),.clk(gclk));
	jor g4158(.dina(w_n4215_1[2]),.dinb(w_n3461_3[1]),.dout(n4216),.clk(gclk));
	jor g4159(.dina(w_n4213_6[1]),.dinb(w_n3554_2[2]),.dout(n4219),.clk(gclk));
	jor g4160(.dina(w_n3837_6[2]),.dinb(w_n3552_3[0]),.dout(n4220),.clk(gclk));
	jand g4161(.dina(n4220),.dinb(n4219),.dout(n4221),.clk(gclk));
	jor g4162(.dina(w_n4063_7[2]),.dinb(w_n3558_2[1]),.dout(n4222),.clk(gclk));
	jand g4163(.dina(n4222),.dinb(n4221),.dout(n4223),.clk(gclk));
	jand g4164(.dina(n4223),.dinb(n4216),.dout(n4224),.clk(gclk));
	jxor g4165(.dina(n4224),.dinb(w_n3023_4[0]),.dout(n4225),.clk(gclk));
	jxor g4166(.dina(w_n4225_0[1]),.dinb(w_n4163_0[1]),.dout(n4226),.clk(gclk));
	jxor g4167(.dina(w_n4226_0[2]),.dinb(n4105),.dout(n4227),.clk(gclk));
	jand g4168(.dina(w_n190_0[2]),.dinb(w_n136_0[2]),.dout(n4228),.clk(gclk));
	jand g4169(.dina(n4228),.dinb(w_n3470_0[1]),.dout(n4229),.clk(gclk));
	jand g4170(.dina(w_n2513_1[0]),.dinb(w_n340_0[1]),.dout(n4230),.clk(gclk));
	jand g4171(.dina(w_n383_0[2]),.dinb(w_n286_1[1]),.dout(n4231),.clk(gclk));
	jand g4172(.dina(n4231),.dinb(w_n817_0[1]),.dout(n4232),.clk(gclk));
	jand g4173(.dina(n4232),.dinb(n4230),.dout(n4233),.clk(gclk));
	jand g4174(.dina(n4233),.dinb(w_n305_0[2]),.dout(n4234),.clk(gclk));
	jand g4175(.dina(n4234),.dinb(n4229),.dout(n4235),.clk(gclk));
	jand g4176(.dina(w_n1313_0[0]),.dinb(w_n569_0[2]),.dout(n4236),.clk(gclk));
	jand g4177(.dina(n4236),.dinb(w_n169_1[0]),.dout(n4237),.clk(gclk));
	jand g4178(.dina(w_n4237_0[2]),.dinb(w_n114_1[0]),.dout(n4238),.clk(gclk));
	jand g4179(.dina(n4238),.dinb(w_n587_1[1]),.dout(n4239),.clk(gclk));
	jand g4180(.dina(n4239),.dinb(n4235),.dout(n4240),.clk(gclk));
	jand g4181(.dina(w_n2751_0[0]),.dinb(w_n260_0[0]),.dout(n4241),.clk(gclk));
	jand g4182(.dina(n4241),.dinb(n4240),.dout(n4242),.clk(gclk));
	jxor g4183(.dina(w_n4242_0[2]),.dinb(w_n4227_0[1]),.dout(n4243),.clk(gclk));
	jxor g4184(.dina(w_n4243_0[1]),.dinb(w_n4100_0[1]),.dout(n4244),.clk(gclk));
	jxor g4185(.dina(w_n4244_0[2]),.dinb(w_n4096_0[1]),.dout(n4245),.clk(gclk));
	jand g4186(.dina(w_n4245_0[1]),.dinb(n4095),.dout(n4246),.clk(gclk));
	jnot g4187(.din(w_n4244_0[1]),.dout(n4247),.clk(gclk));
	jand g4188(.dina(n4247),.dinb(w_n4094_0[0]),.dout(n4248),.clk(gclk));
	jor g4189(.dina(n4248),.dinb(n4246),.dout(w_dff_A_aLvUiHOn0_2),.clk(gclk));
	jand g4190(.dina(w_n4244_0[0]),.dinb(w_n4096_0[0]),.dout(n4250),.clk(gclk));
	jor g4191(.dina(w_n4242_0[1]),.dinb(w_n4227_0[0]),.dout(n4251),.clk(gclk));
	jnot g4192(.din(w_n4251_0[1]),.dout(n4252),.clk(gclk));
	jand g4193(.dina(w_n4243_0[0]),.dinb(w_n4100_0[0]),.dout(n4253),.clk(gclk));
	jor g4194(.dina(n4253),.dinb(n4252),.dout(n4254),.clk(gclk));
	jand g4195(.dina(w_n897_0[2]),.dinb(w_n460_1[0]),.dout(n4255),.clk(gclk));
	jand g4196(.dina(n4255),.dinb(w_n389_1[0]),.dout(n4256),.clk(gclk));
	jand g4197(.dina(n4256),.dinb(w_n488_1[2]),.dout(n4257),.clk(gclk));
	jand g4198(.dina(n4257),.dinb(w_n1109_0[0]),.dout(n4258),.clk(gclk));
	jand g4199(.dina(w_n384_1[0]),.dinb(w_n339_1[2]),.dout(n4259),.clk(gclk));
	jand g4200(.dina(n4259),.dinb(w_n1365_0[1]),.dout(n4260),.clk(gclk));
	jand g4201(.dina(n4260),.dinb(w_n124_0[2]),.dout(n4261),.clk(gclk));
	jand g4202(.dina(w_n3179_0[1]),.dinb(w_n176_0[1]),.dout(n4262),.clk(gclk));
	jand g4203(.dina(w_n377_1[1]),.dinb(w_n191_1[1]),.dout(n4263),.clk(gclk));
	jand g4204(.dina(w_n221_1[0]),.dinb(w_n158_0[1]),.dout(n4264),.clk(gclk));
	jand g4205(.dina(n4264),.dinb(n4263),.dout(n4265),.clk(gclk));
	jand g4206(.dina(n4265),.dinb(n4262),.dout(n4266),.clk(gclk));
	jand g4207(.dina(w_n4266_0[1]),.dinb(w_n1448_0[0]),.dout(n4267),.clk(gclk));
	jand g4208(.dina(n4267),.dinb(n4261),.dout(n4268),.clk(gclk));
	jand g4209(.dina(n4268),.dinb(w_n3892_0[1]),.dout(n4269),.clk(gclk));
	jand g4210(.dina(n4269),.dinb(n4258),.dout(n4270),.clk(gclk));
	jnot g4211(.din(w_n4270_0[1]),.dout(n4271),.clk(gclk));
	jand g4212(.dina(w_n4225_0[0]),.dinb(w_n4163_0[0]),.dout(n4272),.clk(gclk));
	jand g4213(.dina(w_n3851_0[0]),.dinb(w_n3763_0[0]),.dout(n4273),.clk(gclk));
	jor g4214(.dina(n4273),.dinb(w_n3972_0[0]),.dout(n4274),.clk(gclk));
	jand g4215(.dina(w_n4075_0[2]),.dinb(w_n4274_0[1]),.dout(n4275),.clk(gclk));
	jor g4216(.dina(n4275),.dinb(w_n4101_0[0]),.dout(n4276),.clk(gclk));
	jand g4217(.dina(w_n4226_0[1]),.dinb(w_n4276_0[1]),.dout(n4277),.clk(gclk));
	jor g4218(.dina(n4277),.dinb(n4272),.dout(n4278),.clk(gclk));
	jand g4219(.dina(w_n4161_0[0]),.dinb(w_n4153_0[0]),.dout(n4279),.clk(gclk));
	jand g4220(.dina(w_n4162_0[0]),.dinb(w_n4108_0[0]),.dout(n4280),.clk(gclk));
	jor g4221(.dina(n4280),.dinb(n4279),.dout(n4281),.clk(gclk));
	jor g4222(.dina(w_n4151_0[0]),.dinb(w_n4143_0[0]),.dout(n4282),.clk(gclk));
	jnot g4223(.din(n4282),.dout(n4283),.clk(gclk));
	jand g4224(.dina(w_n4152_0[0]),.dinb(w_n4112_0[0]),.dout(n4284),.clk(gclk));
	jor g4225(.dina(n4284),.dinb(n4283),.dout(n4285),.clk(gclk));
	jor g4226(.dina(w_n4140_0[0]),.dinb(w_n4132_0[0]),.dout(n4286),.clk(gclk));
	jand g4227(.dina(w_n4141_0[0]),.dinb(w_n4115_0[0]),.dout(n4287),.clk(gclk));
	jnot g4228(.din(n4287),.dout(n4288),.clk(gclk));
	jand g4229(.dina(n4288),.dinb(n4286),.dout(n4289),.clk(gclk));
	jnot g4230(.din(n4289),.dout(n4290),.clk(gclk));
	jor g4231(.dina(w_n4130_0[0]),.dinb(w_n4120_0[0]),.dout(n4291),.clk(gclk));
	jand g4232(.dina(w_n4128_0[0]),.dinb(w_n1438_14[1]),.dout(n4292),.clk(gclk));
	jand g4233(.dina(n4292),.dinb(w_n2690_0[2]),.dout(n4293),.clk(gclk));
	jnot g4234(.din(n4293),.dout(n4294),.clk(gclk));
	jand g4235(.dina(n4294),.dinb(n4291),.dout(n4295),.clk(gclk));
	jor g4236(.dina(w_n2802_0[1]),.dinb(w_n3384_6[1]),.dout(n4296),.clk(gclk));
	jand g4237(.dina(w_n2943_1[1]),.dinb(w_n2491_1[2]),.dout(n4297),.clk(gclk));
	jand g4238(.dina(w_n2683_1[1]),.dinb(w_n2488_1[2]),.dout(n4298),.clk(gclk));
	jand g4239(.dina(w_n2923_2[0]),.dinb(w_n2684_1[1]),.dout(n4299),.clk(gclk));
	jor g4240(.dina(n4299),.dinb(n4298),.dout(n4300),.clk(gclk));
	jor g4241(.dina(n4300),.dinb(n4297),.dout(n4301),.clk(gclk));
	jnot g4242(.din(n4301),.dout(n4302),.clk(gclk));
	jand g4243(.dina(n4302),.dinb(n4296),.dout(n4303),.clk(gclk));
	jand g4244(.dina(w_n2471_2[1]),.dinb(w_n1438_14[0]),.dout(n4304),.clk(gclk));
	jxor g4245(.dina(n4304),.dinb(w_n4303_0[1]),.dout(n4305),.clk(gclk));
	jxor g4246(.dina(w_n4305_0[1]),.dinb(w_n4295_0[1]),.dout(n4306),.clk(gclk));
	jnot g4247(.din(n4306),.dout(n4307),.clk(gclk));
	jor g4248(.dina(w_n3229_0[2]),.dinb(w_n2252_5[1]),.dout(n4308),.clk(gclk));
	jor g4249(.dina(w_n3166_4[2]),.dinb(w_n2355_5[0]),.dout(n4309),.clk(gclk));
	jor g4250(.dina(w_n3216_3[2]),.dinb(w_n2359_5[1]),.dout(n4310),.clk(gclk));
	jand g4251(.dina(n4310),.dinb(n4309),.dout(n4311),.clk(gclk));
	jor g4252(.dina(w_n3008_3[0]),.dinb(w_n2357_5[1]),.dout(n4312),.clk(gclk));
	jand g4253(.dina(n4312),.dinb(n4311),.dout(n4313),.clk(gclk));
	jand g4254(.dina(n4313),.dinb(n4308),.dout(n4314),.clk(gclk));
	jxor g4255(.dina(n4314),.dinb(w_n1356_5[2]),.dout(n4315),.clk(gclk));
	jxor g4256(.dina(w_n4315_0[1]),.dinb(w_n4307_0[1]),.dout(n4316),.clk(gclk));
	jxor g4257(.dina(w_n4316_0[1]),.dinb(w_n4290_0[1]),.dout(n4317),.clk(gclk));
	jor g4258(.dina(w_n3579_1[0]),.dinb(w_n2506_4[1]),.dout(n4318),.clk(gclk));
	jor g4259(.dina(w_n3495_5[1]),.dinb(w_n2810_4[0]),.dout(n4319),.clk(gclk));
	jor g4260(.dina(w_n3203_4[2]),.dinb(w_n2816_4[1]),.dout(n4320),.clk(gclk));
	jor g4261(.dina(w_n3441_4[1]),.dinb(w_n2807_4[1]),.dout(n4321),.clk(gclk));
	jand g4262(.dina(n4321),.dinb(n4320),.dout(n4322),.clk(gclk));
	jand g4263(.dina(n4322),.dinb(n4319),.dout(n4323),.clk(gclk));
	jand g4264(.dina(n4323),.dinb(n4318),.dout(n4324),.clk(gclk));
	jxor g4265(.dina(n4324),.dinb(w_n1259_5[0]),.dout(n4325),.clk(gclk));
	jxor g4266(.dina(w_n4325_0[1]),.dinb(w_n4317_0[1]),.dout(n4326),.clk(gclk));
	jxor g4267(.dina(w_n4326_0[1]),.dinb(w_n4285_0[1]),.dout(n4327),.clk(gclk));
	jor g4268(.dina(w_n3842_1[1]),.dinb(w_n3029_3[1]),.dout(n4328),.clk(gclk));
	jor g4269(.dina(w_n3837_6[1]),.dinb(w_n3213_3[0]),.dout(n4329),.clk(gclk));
	jor g4270(.dina(w_n3547_5[2]),.dinb(w_n3210_3[1]),.dout(n4330),.clk(gclk));
	jor g4271(.dina(w_n3510_6[0]),.dinb(w_n3219_3[1]),.dout(n4331),.clk(gclk));
	jand g4272(.dina(n4331),.dinb(n4330),.dout(n4332),.clk(gclk));
	jand g4273(.dina(n4332),.dinb(n4329),.dout(n4333),.clk(gclk));
	jand g4274(.dina(n4333),.dinb(n4328),.dout(n4334),.clk(gclk));
	jxor g4275(.dina(n4334),.dinb(w_n1156_5[0]),.dout(n4335),.clk(gclk));
	jxor g4276(.dina(w_n4335_0[1]),.dinb(w_n4327_0[1]),.dout(n4336),.clk(gclk));
	jxor g4277(.dina(w_n4336_0[1]),.dinb(w_n4281_0[1]),.dout(n4337),.clk(gclk));
	jnot g4278(.din(w_n4213_6[0]),.dout(n4338),.clk(gclk));
	jnot g4279(.din(w_n4063_7[1]),.dout(n4339),.clk(gclk));
	jnot g4280(.din(w_n4214_0[1]),.dout(n4340),.clk(gclk));
	jand g4281(.dina(n4340),.dinb(w_n4194_0[0]),.dout(n4341),.clk(gclk));
	jor g4282(.dina(n4341),.dinb(n4339),.dout(n4342),.clk(gclk));
	jand g4283(.dina(n4342),.dinb(w_n4338_1[2]),.dout(n4343),.clk(gclk));
	jnot g4284(.din(w_n4065_0[0]),.dout(n4344),.clk(gclk));
	jor g4285(.dina(w_n4344_0[1]),.dinb(w_n4043_0[0]),.dout(n4345),.clk(gclk));
	jand g4286(.dina(n4345),.dinb(w_n4064_0[0]),.dout(n4346),.clk(gclk));
	jor g4287(.dina(w_n4214_0[0]),.dinb(n4346),.dout(n4347),.clk(gclk));
	jand g4288(.dina(w_n4213_5[2]),.dinb(n4347),.dout(n4348),.clk(gclk));
	jor g4289(.dina(n4348),.dinb(w_n4343_2[1]),.dout(n4349),.clk(gclk));
	jor g4290(.dina(w_n4349_1[2]),.dinb(w_n3461_3[0]),.dout(n4350),.clk(gclk));
	jor g4291(.dina(w_n4063_7[0]),.dinb(w_n3552_2[2]),.dout(n4351),.clk(gclk));
	jor g4292(.dina(w_n4213_5[1]),.dinb(w_n3558_2[0]),.dout(n4352),.clk(gclk));
	jand g4293(.dina(n4352),.dinb(n4351),.dout(n4353),.clk(gclk));
	jand g4294(.dina(n4353),.dinb(n4350),.dout(n4354),.clk(gclk));
	jxor g4295(.dina(n4354),.dinb(w_n3023_3[2]),.dout(n4355),.clk(gclk));
	jxor g4296(.dina(w_n4355_0[1]),.dinb(w_n4337_0[1]),.dout(n4356),.clk(gclk));
	jxor g4297(.dina(w_n4356_0[1]),.dinb(w_n4278_0[1]),.dout(n4357),.clk(gclk));
	jxor g4298(.dina(w_n4357_0[2]),.dinb(w_n4271_0[1]),.dout(n4358),.clk(gclk));
	jxor g4299(.dina(w_n4358_0[1]),.dinb(w_n4254_0[1]),.dout(n4359),.clk(gclk));
	jxor g4300(.dina(w_n4359_0[1]),.dinb(w_n4250_0[1]),.dout(n4360),.clk(gclk));
	jor g4301(.dina(w_n4245_0[0]),.dinb(w_sin0_0[0]),.dout(n4361),.clk(gclk));
	jand g4302(.dina(w_n4361_0[1]),.dinb(w_n4093_11[0]),.dout(n4362),.clk(gclk));
	jxor g4303(.dina(n4362),.dinb(w_n4360_0[1]),.dout(w_dff_A_N1eAxMfr7_2),.clk(gclk));
	jor g4304(.dina(w_n4361_0[0]),.dinb(w_n4360_0[0]),.dout(n4364),.clk(gclk));
	jand g4305(.dina(w_n4364_0[1]),.dinb(w_n4093_10[2]),.dout(n4365),.clk(gclk));
	jand g4306(.dina(w_n4359_0[0]),.dinb(w_n4250_0[0]),.dout(n4366),.clk(gclk));
	jand g4307(.dina(w_n4357_0[1]),.dinb(w_n4271_0[0]),.dout(n4367),.clk(gclk));
	jand g4308(.dina(w_n4358_0[0]),.dinb(w_n4254_0[0]),.dout(n4368),.clk(gclk));
	jor g4309(.dina(n4368),.dinb(w_n4367_0[1]),.dout(n4369),.clk(gclk));
	jand g4310(.dina(w_n2964_0[0]),.dinb(w_n535_1[0]),.dout(n4370),.clk(gclk));
	jand g4311(.dina(n4370),.dinb(w_n2513_0[2]),.dout(n4371),.clk(gclk));
	jand g4312(.dina(n4371),.dinb(w_n2738_0[0]),.dout(n4372),.clk(gclk));
	jand g4313(.dina(w_n1460_0[1]),.dinb(w_n462_0[2]),.dout(n4373),.clk(gclk));
	jand g4314(.dina(n4373),.dinb(w_n1135_0[1]),.dout(n4374),.clk(gclk));
	jand g4315(.dina(n4374),.dinb(n4372),.dout(n4375),.clk(gclk));
	jand g4316(.dina(w_n3875_0[0]),.dinb(w_n197_1[0]),.dout(n4376),.clk(gclk));
	jand g4317(.dina(w_n568_0[1]),.dinb(w_n286_1[0]),.dout(n4377),.clk(gclk));
	jand g4318(.dina(n4377),.dinb(w_n1045_0[0]),.dout(n4378),.clk(gclk));
	jand g4319(.dina(n4378),.dinb(n4376),.dout(n4379),.clk(gclk));
	jand g4320(.dina(n4379),.dinb(w_n1331_0[0]),.dout(n4380),.clk(gclk));
	jand g4321(.dina(n4380),.dinb(n4375),.dout(n4381),.clk(gclk));
	jnot g4322(.din(w_n4381_0[1]),.dout(n4382),.clk(gclk));
	jand g4323(.dina(w_n4355_0[0]),.dinb(w_n4337_0[0]),.dout(n4383),.clk(gclk));
	jand g4324(.dina(w_n4356_0[0]),.dinb(w_n4278_0[0]),.dout(n4384),.clk(gclk));
	jor g4325(.dina(n4384),.dinb(n4383),.dout(n4385),.clk(gclk));
	jand g4326(.dina(w_n4335_0[0]),.dinb(w_n4327_0[0]),.dout(n4386),.clk(gclk));
	jand g4327(.dina(w_n4336_0[0]),.dinb(w_n4281_0[0]),.dout(n4387),.clk(gclk));
	jor g4328(.dina(n4387),.dinb(n4386),.dout(n4388),.clk(gclk));
	jand g4329(.dina(w_n4325_0[0]),.dinb(w_n4317_0[0]),.dout(n4389),.clk(gclk));
	jand g4330(.dina(w_n4326_0[0]),.dinb(w_n4285_0[0]),.dout(n4390),.clk(gclk));
	jor g4331(.dina(n4390),.dinb(n4389),.dout(n4391),.clk(gclk));
	jor g4332(.dina(w_n4315_0[0]),.dinb(w_n4307_0[0]),.dout(n4392),.clk(gclk));
	jand g4333(.dina(w_n4316_0[0]),.dinb(w_n4290_0[0]),.dout(n4393),.clk(gclk));
	jnot g4334(.din(n4393),.dout(n4394),.clk(gclk));
	jand g4335(.dina(n4394),.dinb(n4392),.dout(n4395),.clk(gclk));
	jnot g4336(.din(n4395),.dout(n4396),.clk(gclk));
	jor g4337(.dina(w_n4305_0[0]),.dinb(w_n4295_0[0]),.dout(n4397),.clk(gclk));
	jand g4338(.dina(w_n4303_0[0]),.dinb(w_n1438_13[2]),.dout(n4398),.clk(gclk));
	jand g4339(.dina(n4398),.dinb(w_n2687_1[0]),.dout(n4399),.clk(gclk));
	jnot g4340(.din(n4399),.dout(n4400),.clk(gclk));
	jand g4341(.dina(n4400),.dinb(n4397),.dout(n4401),.clk(gclk));
	jor g4342(.dina(w_n3010_0[1]),.dinb(w_n3384_6[0]),.dout(n4402),.clk(gclk));
	jand g4343(.dina(w_n2943_1[0]),.dinb(w_n2488_1[1]),.dout(n4403),.clk(gclk));
	jand g4344(.dina(w_n3147_0[2]),.dinb(w_n2491_1[1]),.dout(n4404),.clk(gclk));
	jand g4345(.dina(w_n2923_1[2]),.dinb(w_n2683_1[0]),.dout(n4405),.clk(gclk));
	jor g4346(.dina(n4405),.dinb(n4404),.dout(n4406),.clk(gclk));
	jor g4347(.dina(n4406),.dinb(n4403),.dout(n4407),.clk(gclk));
	jnot g4348(.din(n4407),.dout(n4408),.clk(gclk));
	jand g4349(.dina(n4408),.dinb(n4402),.dout(n4409),.clk(gclk));
	jand g4350(.dina(w_n2813_2[0]),.dinb(w_n1438_13[1]),.dout(n4410),.clk(gclk));
	jxor g4351(.dina(n4410),.dinb(w_n4409_0[1]),.dout(n4411),.clk(gclk));
	jxor g4352(.dina(w_n4411_0[1]),.dinb(w_n4401_0[1]),.dout(n4412),.clk(gclk));
	jnot g4353(.din(n4412),.dout(n4413),.clk(gclk));
	jor g4354(.dina(w_n3205_0[2]),.dinb(w_n2252_5[0]),.dout(n4414),.clk(gclk));
	jor g4355(.dina(w_n3166_4[1]),.dinb(w_n2359_5[0]),.dout(n4415),.clk(gclk));
	jor g4356(.dina(w_n3203_4[1]),.dinb(w_n2355_4[2]),.dout(n4416),.clk(gclk));
	jand g4357(.dina(n4416),.dinb(n4415),.dout(n4417),.clk(gclk));
	jor g4358(.dina(w_n3216_3[1]),.dinb(w_n2357_5[0]),.dout(n4418),.clk(gclk));
	jand g4359(.dina(n4418),.dinb(n4417),.dout(n4419),.clk(gclk));
	jand g4360(.dina(n4419),.dinb(n4414),.dout(n4420),.clk(gclk));
	jxor g4361(.dina(n4420),.dinb(w_n1356_5[1]),.dout(n4421),.clk(gclk));
	jxor g4362(.dina(w_n4421_0[1]),.dinb(w_n4413_0[1]),.dout(n4422),.clk(gclk));
	jxor g4363(.dina(w_n4422_0[1]),.dinb(w_n4396_0[1]),.dout(n4423),.clk(gclk));
	jnot g4364(.din(n4423),.dout(n4424),.clk(gclk));
	jor g4365(.dina(w_n3566_1[0]),.dinb(w_n2506_4[0]),.dout(n4425),.clk(gclk));
	jor g4366(.dina(w_n3495_5[0]),.dinb(w_n2807_4[0]),.dout(n4426),.clk(gclk));
	jor g4367(.dina(w_n3510_5[2]),.dinb(w_n2810_3[2]),.dout(n4427),.clk(gclk));
	jand g4368(.dina(n4427),.dinb(n4426),.dout(n4428),.clk(gclk));
	jor g4369(.dina(w_n3441_4[0]),.dinb(w_n2816_4[0]),.dout(n4429),.clk(gclk));
	jand g4370(.dina(n4429),.dinb(n4428),.dout(n4430),.clk(gclk));
	jand g4371(.dina(n4430),.dinb(n4425),.dout(n4431),.clk(gclk));
	jxor g4372(.dina(n4431),.dinb(w_n1257_5[1]),.dout(n4432),.clk(gclk));
	jxor g4373(.dina(w_n4432_0[1]),.dinb(w_n4424_0[1]),.dout(n4433),.clk(gclk));
	jxor g4374(.dina(w_n4433_0[1]),.dinb(w_n4391_0[1]),.dout(n4434),.clk(gclk));
	jor g4375(.dina(w_n4066_1[1]),.dinb(w_n3029_3[0]),.dout(n4435),.clk(gclk));
	jor g4376(.dina(w_n3837_6[0]),.dinb(w_n3210_3[0]),.dout(n4436),.clk(gclk));
	jor g4377(.dina(w_n4063_6[2]),.dinb(w_n3213_2[2]),.dout(n4437),.clk(gclk));
	jand g4378(.dina(n4437),.dinb(n4436),.dout(n4438),.clk(gclk));
	jor g4379(.dina(w_n3547_5[1]),.dinb(w_n3219_3[0]),.dout(n4439),.clk(gclk));
	jand g4380(.dina(n4439),.dinb(n4438),.dout(n4440),.clk(gclk));
	jand g4381(.dina(n4440),.dinb(n4435),.dout(n4441),.clk(gclk));
	jxor g4382(.dina(n4441),.dinb(w_n1154_4[0]),.dout(n4442),.clk(gclk));
	jxor g4383(.dina(w_n4442_0[1]),.dinb(w_n4434_0[1]),.dout(n4443),.clk(gclk));
	jor g4384(.dina(w_n4213_5[0]),.dinb(w_n3552_2[1]),.dout(n4444),.clk(gclk));
	jnot g4385(.din(w_n4343_2[0]),.dout(n4445),.clk(gclk));
	jor g4386(.dina(n4445),.dinb(w_n3461_2[2]),.dout(n4446),.clk(gclk));
	jand g4387(.dina(n4446),.dinb(n4444),.dout(n4447),.clk(gclk));
	jxor g4388(.dina(n4447),.dinb(w_n3455_3[2]),.dout(n4448),.clk(gclk));
	jxor g4389(.dina(w_n4448_0[1]),.dinb(w_n4443_0[1]),.dout(n4449),.clk(gclk));
	jxor g4390(.dina(w_n4449_0[1]),.dinb(w_n4388_0[1]),.dout(n4450),.clk(gclk));
	jxor g4391(.dina(w_n4450_0[1]),.dinb(w_n4385_0[1]),.dout(n4451),.clk(gclk));
	jxor g4392(.dina(w_n4451_0[2]),.dinb(w_n4382_0[1]),.dout(n4452),.clk(gclk));
	jxor g4393(.dina(w_n4452_0[1]),.dinb(w_n4369_0[1]),.dout(n4453),.clk(gclk));
	jxor g4394(.dina(w_n4453_0[1]),.dinb(w_n4366_0[1]),.dout(n4454),.clk(gclk));
	jxor g4395(.dina(w_n4454_0[1]),.dinb(n4365),.dout(w_dff_A_GpXyXXB64_2),.clk(gclk));
	jand g4396(.dina(w_n4453_0[0]),.dinb(w_n4366_0[0]),.dout(n4456),.clk(gclk));
	jand g4397(.dina(w_n4451_0[1]),.dinb(w_n4382_0[0]),.dout(n4457),.clk(gclk));
	jand g4398(.dina(w_n4452_0[0]),.dinb(w_n4369_0[0]),.dout(n4458),.clk(gclk));
	jor g4399(.dina(n4458),.dinb(w_n4457_0[1]),.dout(n4459),.clk(gclk));
	jand g4400(.dina(w_n1073_0[1]),.dinb(w_n280_1[0]),.dout(n4460),.clk(gclk));
	jand g4401(.dina(n4460),.dinb(w_n1322_0[1]),.dout(n4461),.clk(gclk));
	jand g4402(.dina(n4461),.dinb(w_n552_0[0]),.dout(n4462),.clk(gclk));
	jand g4403(.dina(n4462),.dinb(w_n300_1[2]),.dout(n4463),.clk(gclk));
	jand g4404(.dina(w_n2127_0[1]),.dinb(w_n904_0[1]),.dout(n4464),.clk(gclk));
	jand g4405(.dina(n4464),.dinb(w_n3179_0[0]),.dout(n4465),.clk(gclk));
	jand g4406(.dina(n4465),.dinb(w_n1235_0[0]),.dout(n4466),.clk(gclk));
	jand g4407(.dina(n4466),.dinb(w_n1974_0[0]),.dout(n4467),.clk(gclk));
	jand g4408(.dina(n4467),.dinb(w_n1016_0[1]),.dout(n4468),.clk(gclk));
	jand g4409(.dina(n4468),.dinb(n4463),.dout(n4469),.clk(gclk));
	jnot g4410(.din(w_n4469_0[1]),.dout(n4470),.clk(gclk));
	jand g4411(.dina(w_n4449_0[0]),.dinb(w_n4388_0[0]),.dout(n4471),.clk(gclk));
	jand g4412(.dina(w_n4450_0[0]),.dinb(w_n4385_0[0]),.dout(n4472),.clk(gclk));
	jor g4413(.dina(n4472),.dinb(n4471),.dout(n4473),.clk(gclk));
	jnot g4414(.din(w_n4434_0[0]),.dout(n4474),.clk(gclk));
	jor g4415(.dina(w_n4442_0[0]),.dinb(n4474),.dout(n4475),.clk(gclk));
	jnot g4416(.din(n4475),.dout(n4476),.clk(gclk));
	jnot g4417(.din(w_n4443_0[0]),.dout(n4477),.clk(gclk));
	jnot g4418(.din(w_n4448_0[0]),.dout(n4478),.clk(gclk));
	jand g4419(.dina(n4478),.dinb(n4477),.dout(n4479),.clk(gclk));
	jor g4420(.dina(n4479),.dinb(n4476),.dout(n4480),.clk(gclk));
	jor g4421(.dina(w_n4432_0[0]),.dinb(w_n4424_0[0]),.dout(n4481),.clk(gclk));
	jand g4422(.dina(w_n4433_0[0]),.dinb(w_n4391_0[0]),.dout(n4482),.clk(gclk));
	jnot g4423(.din(n4482),.dout(n4483),.clk(gclk));
	jand g4424(.dina(n4483),.dinb(n4481),.dout(n4484),.clk(gclk));
	jor g4425(.dina(w_n4421_0[0]),.dinb(w_n4413_0[0]),.dout(n4485),.clk(gclk));
	jand g4426(.dina(w_n4422_0[0]),.dinb(w_n4396_0[0]),.dout(n4486),.clk(gclk));
	jnot g4427(.din(n4486),.dout(n4487),.clk(gclk));
	jand g4428(.dina(n4487),.dinb(n4485),.dout(n4488),.clk(gclk));
	jnot g4429(.din(n4488),.dout(n4489),.clk(gclk));
	jor g4430(.dina(w_n4411_0[0]),.dinb(w_n4401_0[0]),.dout(n4490),.clk(gclk));
	jand g4431(.dina(w_n4409_0[0]),.dinb(w_n1438_13[0]),.dout(n4491),.clk(gclk));
	jand g4432(.dina(n4491),.dinb(w_n2684_1[0]),.dout(n4492),.clk(gclk));
	jnot g4433(.din(n4492),.dout(n4493),.clk(gclk));
	jand g4434(.dina(n4493),.dinb(n4490),.dout(n4494),.clk(gclk));
	jnot g4435(.din(n4494),.dout(n4495),.clk(gclk));
	jand g4436(.dina(w_n2683_0[2]),.dinb(w_n1438_12[2]),.dout(n4496),.clk(gclk));
	jxor g4437(.dina(w_n4496_0[1]),.dinb(w_n3455_3[1]),.dout(n4497),.clk(gclk));
	jor g4438(.dina(w_n3242_0[1]),.dinb(w_n3384_5[2]),.dout(n4498),.clk(gclk));
	jor g4439(.dina(w_n3008_2[2]),.dinb(w_n3390_4[1]),.dout(n4499),.clk(gclk));
	jor g4440(.dina(w_n3216_3[0]),.dinb(w_n3386_4[0]),.dout(n4500),.clk(gclk));
	jand g4441(.dina(n4500),.dinb(n4499),.dout(n4501),.clk(gclk));
	jor g4442(.dina(w_n3388_4[1]),.dinb(w_n2800_2[1]),.dout(n4502),.clk(gclk));
	jand g4443(.dina(n4502),.dinb(n4501),.dout(n4503),.clk(gclk));
	jand g4444(.dina(n4503),.dinb(n4498),.dout(n4504),.clk(gclk));
	jxor g4445(.dina(n4504),.dinb(w_n2051_5[1]),.dout(n4505),.clk(gclk));
	jxor g4446(.dina(w_n4505_0[1]),.dinb(w_n4497_0[1]),.dout(n4506),.clk(gclk));
	jxor g4447(.dina(w_n4506_0[1]),.dinb(w_n4495_0[1]),.dout(n4507),.clk(gclk));
	jnot g4448(.din(n4507),.dout(n4508),.clk(gclk));
	jor g4449(.dina(w_n3443_0[2]),.dinb(w_n2252_4[2]),.dout(n4509),.clk(gclk));
	jor g4450(.dina(w_n3441_3[2]),.dinb(w_n2355_4[1]),.dout(n4510),.clk(gclk));
	jor g4451(.dina(w_n3203_4[0]),.dinb(w_n2359_4[2]),.dout(n4511),.clk(gclk));
	jand g4452(.dina(n4511),.dinb(n4510),.dout(n4512),.clk(gclk));
	jor g4453(.dina(w_n3166_4[0]),.dinb(w_n2357_4[2]),.dout(n4513),.clk(gclk));
	jand g4454(.dina(n4513),.dinb(n4512),.dout(n4514),.clk(gclk));
	jand g4455(.dina(n4514),.dinb(n4509),.dout(n4515),.clk(gclk));
	jxor g4456(.dina(n4515),.dinb(w_n1356_5[0]),.dout(n4516),.clk(gclk));
	jxor g4457(.dina(w_n4516_0[1]),.dinb(w_n4508_0[1]),.dout(n4517),.clk(gclk));
	jxor g4458(.dina(w_n4517_0[1]),.dinb(w_n4489_0[1]),.dout(n4518),.clk(gclk));
	jor g4459(.dina(w_n3550_1[0]),.dinb(w_n2506_3[2]),.dout(n4519),.clk(gclk));
	jor g4460(.dina(w_n3547_5[0]),.dinb(w_n2810_3[1]),.dout(n4520),.clk(gclk));
	jor g4461(.dina(w_n3510_5[1]),.dinb(w_n2807_3[2]),.dout(n4521),.clk(gclk));
	jor g4462(.dina(w_n3495_4[2]),.dinb(w_n2816_3[2]),.dout(n4522),.clk(gclk));
	jand g4463(.dina(n4522),.dinb(n4521),.dout(n4523),.clk(gclk));
	jand g4464(.dina(n4523),.dinb(n4520),.dout(n4524),.clk(gclk));
	jand g4465(.dina(n4524),.dinb(n4519),.dout(n4525),.clk(gclk));
	jxor g4466(.dina(n4525),.dinb(w_n1259_4[2]),.dout(n4526),.clk(gclk));
	jxor g4467(.dina(w_n4526_0[1]),.dinb(w_n4518_0[1]),.dout(n4527),.clk(gclk));
	jxor g4468(.dina(w_n4527_0[1]),.dinb(w_n4484_0[1]),.dout(n4528),.clk(gclk));
	jor g4469(.dina(w_n4215_1[1]),.dinb(w_n3029_2[2]),.dout(n4529),.clk(gclk));
	jor g4470(.dina(w_n4063_6[1]),.dinb(w_n3210_2[2]),.dout(n4530),.clk(gclk));
	jor g4471(.dina(w_n3837_5[2]),.dinb(w_n3219_2[2]),.dout(n4531),.clk(gclk));
	jor g4472(.dina(w_n4213_4[2]),.dinb(w_n3213_2[1]),.dout(n4532),.clk(gclk));
	jand g4473(.dina(n4532),.dinb(n4531),.dout(n4533),.clk(gclk));
	jand g4474(.dina(n4533),.dinb(n4530),.dout(n4534),.clk(gclk));
	jand g4475(.dina(n4534),.dinb(n4529),.dout(n4535),.clk(gclk));
	jxor g4476(.dina(n4535),.dinb(w_n1154_3[2]),.dout(n4536),.clk(gclk));
	jxor g4477(.dina(w_n4536_0[1]),.dinb(w_n4528_0[1]),.dout(n4537),.clk(gclk));
	jxor g4478(.dina(w_n4537_0[1]),.dinb(w_n4480_0[1]),.dout(n4538),.clk(gclk));
	jxor g4479(.dina(w_n4538_0[1]),.dinb(w_n4473_0[1]),.dout(n4539),.clk(gclk));
	jxor g4480(.dina(w_n4539_0[2]),.dinb(w_n4470_0[1]),.dout(n4540),.clk(gclk));
	jxor g4481(.dina(w_n4540_0[1]),.dinb(w_n4459_0[1]),.dout(n4541),.clk(gclk));
	jxor g4482(.dina(w_n4541_0[1]),.dinb(w_n4456_0[1]),.dout(n4542),.clk(gclk));
	jor g4483(.dina(w_n4454_0[0]),.dinb(w_n4364_0[0]),.dout(n4543),.clk(gclk));
	jand g4484(.dina(w_n4543_0[1]),.dinb(w_n4093_10[1]),.dout(n4544),.clk(gclk));
	jxor g4485(.dina(n4544),.dinb(w_n4542_0[1]),.dout(w_dff_A_Kjg55Kq01_2),.clk(gclk));
	jand g4486(.dina(w_n4541_0[0]),.dinb(w_n4456_0[0]),.dout(n4546),.clk(gclk));
	jand g4487(.dina(w_n4539_0[1]),.dinb(w_n4470_0[0]),.dout(n4547),.clk(gclk));
	jand g4488(.dina(w_n4540_0[0]),.dinb(w_n4459_0[0]),.dout(n4548),.clk(gclk));
	jor g4489(.dina(n4548),.dinb(w_n4547_0[1]),.dout(n4549),.clk(gclk));
	jand g4490(.dina(w_n361_0[2]),.dinb(w_n280_0[2]),.dout(n4550),.clk(gclk));
	jand g4491(.dina(w_n2617_0[0]),.dinb(w_n850_0[0]),.dout(n4551),.clk(gclk));
	jand g4492(.dina(n4551),.dinb(n4550),.dout(n4552),.clk(gclk));
	jand g4493(.dina(n4552),.dinb(w_n4203_0[0]),.dout(n4553),.clk(gclk));
	jand g4494(.dina(w_n378_1[0]),.dinb(w_n248_1[0]),.dout(n4554),.clk(gclk));
	jand g4495(.dina(n4554),.dinb(w_n539_0[1]),.dout(n4555),.clk(gclk));
	jand g4496(.dina(w_n2623_0[1]),.dinb(w_n316_0[0]),.dout(n4556),.clk(gclk));
	jand g4497(.dina(w_n510_1[0]),.dinb(w_n411_0[2]),.dout(n4557),.clk(gclk));
	jand g4498(.dina(n4557),.dinb(w_n535_0[2]),.dout(n4558),.clk(gclk));
	jand g4499(.dina(w_n4558_0[2]),.dinb(w_n4556_0[1]),.dout(n4559),.clk(gclk));
	jand g4500(.dina(n4559),.dinb(n4555),.dout(n4560),.clk(gclk));
	jand g4501(.dina(n4560),.dinb(w_n4237_0[1]),.dout(n4561),.clk(gclk));
	jand g4502(.dina(n4561),.dinb(w_n3481_0[1]),.dout(n4562),.clk(gclk));
	jand g4503(.dina(n4562),.dinb(n4553),.dout(n4563),.clk(gclk));
	jnot g4504(.din(w_n4563_0[1]),.dout(n4564),.clk(gclk));
	jand g4505(.dina(w_n4537_0[0]),.dinb(w_n4480_0[0]),.dout(n4565),.clk(gclk));
	jand g4506(.dina(w_n4538_0[0]),.dinb(w_n4473_0[0]),.dout(n4566),.clk(gclk));
	jor g4507(.dina(n4566),.dinb(n4565),.dout(n4567),.clk(gclk));
	jnot g4508(.din(w_n4484_0[0]),.dout(n4568),.clk(gclk));
	jand g4509(.dina(w_n4527_0[0]),.dinb(n4568),.dout(n4569),.clk(gclk));
	jor g4510(.dina(w_n4536_0[0]),.dinb(w_n4528_0[0]),.dout(n4570),.clk(gclk));
	jnot g4511(.din(n4570),.dout(n4571),.clk(gclk));
	jor g4512(.dina(n4571),.dinb(n4569),.dout(n4572),.clk(gclk));
	jand g4513(.dina(w_n4517_0[0]),.dinb(w_n4489_0[0]),.dout(n4573),.clk(gclk));
	jand g4514(.dina(w_n4526_0[0]),.dinb(w_n4518_0[0]),.dout(n4574),.clk(gclk));
	jor g4515(.dina(n4574),.dinb(n4573),.dout(n4575),.clk(gclk));
	jand g4516(.dina(w_n4506_0[0]),.dinb(w_n4495_0[0]),.dout(n4576),.clk(gclk));
	jnot g4517(.din(n4576),.dout(n4577),.clk(gclk));
	jor g4518(.dina(w_n4516_0[0]),.dinb(w_n4508_0[0]),.dout(n4578),.clk(gclk));
	jand g4519(.dina(n4578),.dinb(n4577),.dout(n4579),.clk(gclk));
	jnot g4520(.din(n4579),.dout(n4580),.clk(gclk));
	jand g4521(.dina(w_n4496_0[0]),.dinb(w_n3455_3[0]),.dout(n4581),.clk(gclk));
	jand g4522(.dina(w_n4505_0[0]),.dinb(w_n4497_0[0]),.dout(n4582),.clk(gclk));
	jor g4523(.dina(n4582),.dinb(n4581),.dout(n4583),.clk(gclk));
	jand g4524(.dina(w_n2943_0[2]),.dinb(w_n1438_12[1]),.dout(n4584),.clk(gclk));
	jxor g4525(.dina(w_n4584_0[1]),.dinb(w_n3455_2[2]),.dout(n4585),.clk(gclk));
	jxor g4526(.dina(w_n4585_0[1]),.dinb(w_n4583_0[1]),.dout(n4586),.clk(gclk));
	jor g4527(.dina(w_n3229_0[1]),.dinb(w_n3384_5[1]),.dout(n4587),.clk(gclk));
	jor g4528(.dina(w_n3166_3[2]),.dinb(w_n3386_3[2]),.dout(n4588),.clk(gclk));
	jor g4529(.dina(w_n3216_2[2]),.dinb(w_n3390_4[0]),.dout(n4589),.clk(gclk));
	jand g4530(.dina(n4589),.dinb(n4588),.dout(n4590),.clk(gclk));
	jor g4531(.dina(w_n3008_2[1]),.dinb(w_n3388_4[0]),.dout(n4591),.clk(gclk));
	jand g4532(.dina(n4591),.dinb(n4590),.dout(n4592),.clk(gclk));
	jand g4533(.dina(n4592),.dinb(n4587),.dout(n4593),.clk(gclk));
	jxor g4534(.dina(n4593),.dinb(w_n2051_5[0]),.dout(n4594),.clk(gclk));
	jxor g4535(.dina(w_n4594_0[1]),.dinb(w_n4586_0[1]),.dout(n4595),.clk(gclk));
	jor g4536(.dina(w_n3579_0[2]),.dinb(w_n2252_4[1]),.dout(n4596),.clk(gclk));
	jor g4537(.dina(w_n3495_4[1]),.dinb(w_n2355_4[0]),.dout(n4597),.clk(gclk));
	jor g4538(.dina(w_n3441_3[1]),.dinb(w_n2359_4[1]),.dout(n4598),.clk(gclk));
	jor g4539(.dina(w_n3203_3[2]),.dinb(w_n2357_4[1]),.dout(n4599),.clk(gclk));
	jand g4540(.dina(n4599),.dinb(n4598),.dout(n4600),.clk(gclk));
	jand g4541(.dina(n4600),.dinb(n4597),.dout(n4601),.clk(gclk));
	jand g4542(.dina(n4601),.dinb(n4596),.dout(n4602),.clk(gclk));
	jxor g4543(.dina(n4602),.dinb(w_n1480_5[1]),.dout(n4603),.clk(gclk));
	jxor g4544(.dina(w_n4603_0[1]),.dinb(w_n4595_0[1]),.dout(n4604),.clk(gclk));
	jxor g4545(.dina(w_n4604_0[1]),.dinb(w_n4580_0[1]),.dout(n4605),.clk(gclk));
	jnot g4546(.din(n4605),.dout(n4606),.clk(gclk));
	jor g4547(.dina(w_n3842_1[0]),.dinb(w_n2506_3[1]),.dout(n4607),.clk(gclk));
	jor g4548(.dina(w_n3547_4[2]),.dinb(w_n2807_3[1]),.dout(n4608),.clk(gclk));
	jor g4549(.dina(w_n3837_5[1]),.dinb(w_n2810_3[0]),.dout(n4609),.clk(gclk));
	jand g4550(.dina(n4609),.dinb(n4608),.dout(n4610),.clk(gclk));
	jor g4551(.dina(w_n3510_5[0]),.dinb(w_n2816_3[1]),.dout(n4611),.clk(gclk));
	jand g4552(.dina(n4611),.dinb(n4610),.dout(n4612),.clk(gclk));
	jand g4553(.dina(n4612),.dinb(n4607),.dout(n4613),.clk(gclk));
	jxor g4554(.dina(n4613),.dinb(w_n1257_5[0]),.dout(n4614),.clk(gclk));
	jxor g4555(.dina(w_n4614_0[1]),.dinb(w_n4606_0[1]),.dout(n4615),.clk(gclk));
	jxor g4556(.dina(w_n4615_0[1]),.dinb(w_n4575_0[1]),.dout(n4616),.clk(gclk));
	jor g4557(.dina(w_n4349_1[1]),.dinb(w_n3029_2[1]),.dout(n4617),.clk(gclk));
	jor g4558(.dina(w_n4063_6[0]),.dinb(w_n3219_2[1]),.dout(n4618),.clk(gclk));
	jor g4559(.dina(w_n4213_4[1]),.dinb(w_n3210_2[1]),.dout(n4619),.clk(gclk));
	jand g4560(.dina(n4619),.dinb(n4618),.dout(n4620),.clk(gclk));
	jand g4561(.dina(n4620),.dinb(n4617),.dout(n4621),.clk(gclk));
	jxor g4562(.dina(n4621),.dinb(w_n1156_4[2]),.dout(n4622),.clk(gclk));
	jxor g4563(.dina(w_n4622_0[1]),.dinb(w_n4616_0[1]),.dout(n4623),.clk(gclk));
	jxor g4564(.dina(w_n4623_0[1]),.dinb(w_n4572_0[1]),.dout(n4624),.clk(gclk));
	jxor g4565(.dina(w_n4624_0[1]),.dinb(w_n4567_0[1]),.dout(n4625),.clk(gclk));
	jxor g4566(.dina(w_n4625_0[2]),.dinb(w_n4564_0[1]),.dout(n4626),.clk(gclk));
	jxor g4567(.dina(w_n4626_0[1]),.dinb(w_n4549_0[1]),.dout(n4627),.clk(gclk));
	jxor g4568(.dina(w_n4627_0[1]),.dinb(w_n4546_0[1]),.dout(n4628),.clk(gclk));
	jor g4569(.dina(w_n4543_0[0]),.dinb(w_n4542_0[0]),.dout(n4629),.clk(gclk));
	jand g4570(.dina(w_n4629_0[1]),.dinb(w_n4093_10[0]),.dout(n4630),.clk(gclk));
	jxor g4571(.dina(n4630),.dinb(w_n4628_0[1]),.dout(w_dff_A_jawdh4xz8_2),.clk(gclk));
	jand g4572(.dina(w_n4627_0[0]),.dinb(w_n4546_0[0]),.dout(n4632),.clk(gclk));
	jand g4573(.dina(w_n4625_0[1]),.dinb(w_n4564_0[0]),.dout(n4633),.clk(gclk));
	jand g4574(.dina(w_n4626_0[0]),.dinb(w_n4549_0[0]),.dout(n4634),.clk(gclk));
	jor g4575(.dina(n4634),.dinb(w_n4633_0[1]),.dout(n4635),.clk(gclk));
	jand g4576(.dina(w_n924_0[0]),.dinb(w_n137_1[0]),.dout(n4636),.clk(gclk));
	jand g4577(.dina(n4636),.dinb(w_n2623_0[0]),.dout(n4637),.clk(gclk));
	jand g4578(.dina(w_n2513_0[1]),.dinb(w_n540_0[0]),.dout(n4638),.clk(gclk));
	jand g4579(.dina(n4638),.dinb(n4637),.dout(n4639),.clk(gclk));
	jand g4580(.dina(w_n3497_0[0]),.dinb(w_n489_1[1]),.dout(n4640),.clk(gclk));
	jand g4581(.dina(n4640),.dinb(w_n1122_0[0]),.dout(n4641),.clk(gclk));
	jand g4582(.dina(n4641),.dinb(w_n2130_0[0]),.dout(n4642),.clk(gclk));
	jand g4583(.dina(n4642),.dinb(n4639),.dout(n4643),.clk(gclk));
	jand g4584(.dina(w_n2628_0[0]),.dinb(w_n276_1[1]),.dout(n4644),.clk(gclk));
	jand g4585(.dina(w_n2135_0[1]),.dinb(w_n128_1[0]),.dout(n4645),.clk(gclk));
	jand g4586(.dina(n4645),.dinb(n4644),.dout(n4646),.clk(gclk));
	jand g4587(.dina(n4646),.dinb(w_n1970_0[0]),.dout(n4647),.clk(gclk));
	jand g4588(.dina(w_n3537_1[1]),.dinb(w_n142_0[2]),.dout(n4648),.clk(gclk));
	jand g4589(.dina(n4648),.dinb(w_n288_0[2]),.dout(n4649),.clk(gclk));
	jand g4590(.dina(n4649),.dinb(n4647),.dout(n4650),.clk(gclk));
	jand g4591(.dina(n4650),.dinb(w_n4643_0[1]),.dout(n4651),.clk(gclk));
	jand g4592(.dina(n4651),.dinb(w_n273_0[0]),.dout(n4652),.clk(gclk));
	jnot g4593(.din(w_n4652_0[1]),.dout(n4653),.clk(gclk));
	jand g4594(.dina(w_n4623_0[0]),.dinb(w_n4572_0[0]),.dout(n4654),.clk(gclk));
	jand g4595(.dina(w_n4624_0[0]),.dinb(w_n4567_0[0]),.dout(n4655),.clk(gclk));
	jor g4596(.dina(n4655),.dinb(n4654),.dout(n4656),.clk(gclk));
	jand g4597(.dina(w_n4615_0[0]),.dinb(w_n4575_0[0]),.dout(n4657),.clk(gclk));
	jand g4598(.dina(w_n4622_0[0]),.dinb(w_n4616_0[0]),.dout(n4658),.clk(gclk));
	jor g4599(.dina(n4658),.dinb(n4657),.dout(n4659),.clk(gclk));
	jand g4600(.dina(w_n4604_0[0]),.dinb(w_n4580_0[0]),.dout(n4660),.clk(gclk));
	jnot g4601(.din(n4660),.dout(n4661),.clk(gclk));
	jor g4602(.dina(w_n4614_0[0]),.dinb(w_n4606_0[0]),.dout(n4662),.clk(gclk));
	jand g4603(.dina(n4662),.dinb(n4661),.dout(n4663),.clk(gclk));
	jand g4604(.dina(w_n4338_1[1]),.dinb(w_n3218_0[0]),.dout(n4664),.clk(gclk));
	jand g4605(.dina(w_n4343_1[2]),.dinb(w_n3028_0[1]),.dout(n4665),.clk(gclk));
	jor g4606(.dina(n4665),.dinb(n4664),.dout(n4666),.clk(gclk));
	jxor g4607(.dina(n4666),.dinb(w_n1156_4[1]),.dout(n4667),.clk(gclk));
	jxor g4608(.dina(w_n4667_0[1]),.dinb(w_n4663_0[1]),.dout(n4668),.clk(gclk));
	jand g4609(.dina(w_n4594_0[0]),.dinb(w_n4586_0[0]),.dout(n4669),.clk(gclk));
	jand g4610(.dina(w_n4603_0[0]),.dinb(w_n4595_0[0]),.dout(n4670),.clk(gclk));
	jor g4611(.dina(n4670),.dinb(n4669),.dout(n4671),.clk(gclk));
	jand g4612(.dina(w_n4584_0[0]),.dinb(w_n3455_2[1]),.dout(n4672),.clk(gclk));
	jand g4613(.dina(w_n4585_0[0]),.dinb(w_n4583_0[0]),.dout(n4673),.clk(gclk));
	jor g4614(.dina(n4673),.dinb(n4672),.dout(n4674),.clk(gclk));
	jand g4615(.dina(w_n3147_0[1]),.dinb(w_n1438_12[0]),.dout(n4675),.clk(gclk));
	jxor g4616(.dina(w_n4675_0[1]),.dinb(w_n3455_2[0]),.dout(n4676),.clk(gclk));
	jxor g4617(.dina(w_n4676_0[1]),.dinb(w_n4674_0[1]),.dout(n4677),.clk(gclk));
	jor g4618(.dina(w_n3205_0[1]),.dinb(w_n3384_5[0]),.dout(n4678),.clk(gclk));
	jor g4619(.dina(w_n3166_3[1]),.dinb(w_n3390_3[2]),.dout(n4679),.clk(gclk));
	jor g4620(.dina(w_n3203_3[1]),.dinb(w_n3386_3[1]),.dout(n4680),.clk(gclk));
	jand g4621(.dina(n4680),.dinb(n4679),.dout(n4681),.clk(gclk));
	jor g4622(.dina(w_n3216_2[1]),.dinb(w_n3388_3[2]),.dout(n4682),.clk(gclk));
	jand g4623(.dina(n4682),.dinb(n4681),.dout(n4683),.clk(gclk));
	jand g4624(.dina(n4683),.dinb(n4678),.dout(n4684),.clk(gclk));
	jxor g4625(.dina(n4684),.dinb(w_n2051_4[2]),.dout(n4685),.clk(gclk));
	jxor g4626(.dina(w_n4685_0[1]),.dinb(w_n4677_0[1]),.dout(n4686),.clk(gclk));
	jor g4627(.dina(w_n3566_0[2]),.dinb(w_n2252_4[0]),.dout(n4687),.clk(gclk));
	jor g4628(.dina(w_n3510_4[2]),.dinb(w_n2355_3[2]),.dout(n4688),.clk(gclk));
	jor g4629(.dina(w_n3495_4[0]),.dinb(w_n2359_4[0]),.dout(n4689),.clk(gclk));
	jor g4630(.dina(w_n3441_3[0]),.dinb(w_n2357_4[0]),.dout(n4690),.clk(gclk));
	jand g4631(.dina(n4690),.dinb(n4689),.dout(n4691),.clk(gclk));
	jand g4632(.dina(n4691),.dinb(n4688),.dout(n4692),.clk(gclk));
	jand g4633(.dina(n4692),.dinb(n4687),.dout(n4693),.clk(gclk));
	jxor g4634(.dina(n4693),.dinb(w_n1480_5[0]),.dout(n4694),.clk(gclk));
	jxor g4635(.dina(w_n4694_0[1]),.dinb(w_n4686_0[1]),.dout(n4695),.clk(gclk));
	jxor g4636(.dina(w_n4695_0[1]),.dinb(w_n4671_0[1]),.dout(n4696),.clk(gclk));
	jnot g4637(.din(n4696),.dout(n4697),.clk(gclk));
	jor g4638(.dina(w_n4066_1[0]),.dinb(w_n2506_3[0]),.dout(n4698),.clk(gclk));
	jor g4639(.dina(w_n3837_5[0]),.dinb(w_n2807_3[0]),.dout(n4699),.clk(gclk));
	jor g4640(.dina(w_n4063_5[2]),.dinb(w_n2810_2[2]),.dout(n4700),.clk(gclk));
	jand g4641(.dina(n4700),.dinb(n4699),.dout(n4701),.clk(gclk));
	jor g4642(.dina(w_n3547_4[1]),.dinb(w_n2816_3[0]),.dout(n4702),.clk(gclk));
	jand g4643(.dina(n4702),.dinb(n4701),.dout(n4703),.clk(gclk));
	jand g4644(.dina(n4703),.dinb(n4698),.dout(n4704),.clk(gclk));
	jxor g4645(.dina(n4704),.dinb(w_n1257_4[2]),.dout(n4705),.clk(gclk));
	jxor g4646(.dina(w_n4705_0[1]),.dinb(w_n4697_0[1]),.dout(n4706),.clk(gclk));
	jxor g4647(.dina(w_n4706_0[1]),.dinb(w_n4668_0[1]),.dout(n4707),.clk(gclk));
	jxor g4648(.dina(w_n4707_0[1]),.dinb(w_n4659_0[1]),.dout(n4708),.clk(gclk));
	jxor g4649(.dina(w_n4708_0[1]),.dinb(w_n4656_0[1]),.dout(n4709),.clk(gclk));
	jxor g4650(.dina(w_n4709_0[2]),.dinb(w_n4653_0[1]),.dout(n4710),.clk(gclk));
	jxor g4651(.dina(w_n4710_0[1]),.dinb(w_n4635_0[1]),.dout(n4711),.clk(gclk));
	jxor g4652(.dina(w_n4711_0[1]),.dinb(w_n4632_0[1]),.dout(n4712),.clk(gclk));
	jor g4653(.dina(w_n4629_0[0]),.dinb(w_n4628_0[0]),.dout(n4713),.clk(gclk));
	jand g4654(.dina(w_n4713_0[1]),.dinb(w_n4093_9[2]),.dout(n4714),.clk(gclk));
	jxor g4655(.dina(n4714),.dinb(w_n4712_0[1]),.dout(w_dff_A_Pe38P7pN5_2),.clk(gclk));
	jand g4656(.dina(w_n4711_0[0]),.dinb(w_n4632_0[0]),.dout(n4716),.clk(gclk));
	jand g4657(.dina(w_n4709_0[1]),.dinb(w_n4653_0[0]),.dout(n4717),.clk(gclk));
	jand g4658(.dina(w_n4710_0[0]),.dinb(w_n4635_0[0]),.dout(n4718),.clk(gclk));
	jor g4659(.dina(n4718),.dinb(w_n4717_0[1]),.dout(n4719),.clk(gclk));
	jand g4660(.dina(w_n4707_0[0]),.dinb(w_n4659_0[0]),.dout(n4720),.clk(gclk));
	jand g4661(.dina(w_n4708_0[0]),.dinb(w_n4656_0[0]),.dout(n4721),.clk(gclk));
	jor g4662(.dina(n4721),.dinb(n4720),.dout(n4722),.clk(gclk));
	jor g4663(.dina(w_n4667_0[0]),.dinb(w_n4663_0[0]),.dout(n4723),.clk(gclk));
	jand g4664(.dina(w_n4706_0[0]),.dinb(w_n4668_0[0]),.dout(n4724),.clk(gclk));
	jnot g4665(.din(n4724),.dout(n4725),.clk(gclk));
	jand g4666(.dina(n4725),.dinb(n4723),.dout(n4726),.clk(gclk));
	jnot g4667(.din(n4726),.dout(n4727),.clk(gclk));
	jand g4668(.dina(w_n4695_0[0]),.dinb(w_n4671_0[0]),.dout(n4728),.clk(gclk));
	jnot g4669(.din(n4728),.dout(n4729),.clk(gclk));
	jor g4670(.dina(w_n4705_0[0]),.dinb(w_n4697_0[0]),.dout(n4730),.clk(gclk));
	jand g4671(.dina(n4730),.dinb(n4729),.dout(n4731),.clk(gclk));
	jor g4672(.dina(w_n4215_1[0]),.dinb(w_n2506_2[2]),.dout(n4732),.clk(gclk));
	jor g4673(.dina(w_n4063_5[1]),.dinb(w_n2807_2[2]),.dout(n4733),.clk(gclk));
	jor g4674(.dina(w_n3837_4[2]),.dinb(w_n2816_2[2]),.dout(n4734),.clk(gclk));
	jor g4675(.dina(w_n4213_4[0]),.dinb(w_n2810_2[1]),.dout(n4735),.clk(gclk));
	jand g4676(.dina(n4735),.dinb(n4734),.dout(n4736),.clk(gclk));
	jand g4677(.dina(n4736),.dinb(n4733),.dout(n4737),.clk(gclk));
	jand g4678(.dina(n4737),.dinb(n4732),.dout(n4738),.clk(gclk));
	jxor g4679(.dina(n4738),.dinb(w_n1257_4[1]),.dout(n4739),.clk(gclk));
	jxor g4680(.dina(w_n4739_0[1]),.dinb(w_n4731_0[1]),.dout(n4740),.clk(gclk));
	jand g4681(.dina(w_n4685_0[0]),.dinb(w_n4677_0[0]),.dout(n4741),.clk(gclk));
	jand g4682(.dina(w_n4694_0[0]),.dinb(w_n4686_0[0]),.dout(n4742),.clk(gclk));
	jor g4683(.dina(n4742),.dinb(n4741),.dout(n4743),.clk(gclk));
	jand g4684(.dina(w_n4675_0[0]),.dinb(w_n3455_1[2]),.dout(n4744),.clk(gclk));
	jand g4685(.dina(w_n4676_0[0]),.dinb(w_n4674_0[0]),.dout(n4745),.clk(gclk));
	jor g4686(.dina(n4745),.dinb(n4744),.dout(n4746),.clk(gclk));
	jand g4687(.dina(w_n3144_0[1]),.dinb(w_n1438_11[2]),.dout(n4747),.clk(gclk));
	jxor g4688(.dina(w_n3455_1[1]),.dinb(w_n1154_3[1]),.dout(n4748),.clk(gclk));
	jxor g4689(.dina(w_n4748_0[1]),.dinb(w_n4747_0[1]),.dout(n4749),.clk(gclk));
	jor g4690(.dina(w_n3443_0[1]),.dinb(w_n3384_4[2]),.dout(n4750),.clk(gclk));
	jor g4691(.dina(w_n3203_3[0]),.dinb(w_n3390_3[1]),.dout(n4751),.clk(gclk));
	jor g4692(.dina(w_n3441_2[2]),.dinb(w_n3386_3[0]),.dout(n4752),.clk(gclk));
	jor g4693(.dina(w_n3166_3[0]),.dinb(w_n3388_3[1]),.dout(n4753),.clk(gclk));
	jand g4694(.dina(n4753),.dinb(n4752),.dout(n4754),.clk(gclk));
	jand g4695(.dina(n4754),.dinb(n4751),.dout(n4755),.clk(gclk));
	jand g4696(.dina(n4755),.dinb(n4750),.dout(n4756),.clk(gclk));
	jxor g4697(.dina(n4756),.dinb(w_n2051_4[1]),.dout(n4757),.clk(gclk));
	jxor g4698(.dina(w_n4757_0[1]),.dinb(w_n4749_0[1]),.dout(n4758),.clk(gclk));
	jxor g4699(.dina(w_n4758_0[1]),.dinb(w_n4746_0[1]),.dout(n4759),.clk(gclk));
	jor g4700(.dina(w_n3550_0[2]),.dinb(w_n2252_3[2]),.dout(n4760),.clk(gclk));
	jor g4701(.dina(w_n3547_4[0]),.dinb(w_n2355_3[1]),.dout(n4761),.clk(gclk));
	jor g4702(.dina(w_n3510_4[1]),.dinb(w_n2359_3[2]),.dout(n4762),.clk(gclk));
	jor g4703(.dina(w_n3495_3[2]),.dinb(w_n2357_3[2]),.dout(n4763),.clk(gclk));
	jand g4704(.dina(n4763),.dinb(n4762),.dout(n4764),.clk(gclk));
	jand g4705(.dina(n4764),.dinb(n4761),.dout(n4765),.clk(gclk));
	jand g4706(.dina(n4765),.dinb(n4760),.dout(n4766),.clk(gclk));
	jxor g4707(.dina(n4766),.dinb(w_n1480_4[2]),.dout(n4767),.clk(gclk));
	jxor g4708(.dina(w_n4767_0[1]),.dinb(w_n4759_0[1]),.dout(n4768),.clk(gclk));
	jxor g4709(.dina(w_n4768_0[1]),.dinb(w_n4743_0[1]),.dout(n4769),.clk(gclk));
	jxor g4710(.dina(w_n4769_0[1]),.dinb(w_n4740_0[1]),.dout(n4770),.clk(gclk));
	jxor g4711(.dina(w_n4770_0[1]),.dinb(w_n4727_0[1]),.dout(n4771),.clk(gclk));
	jnot g4712(.din(w_n4771_0[2]),.dout(n4772),.clk(gclk));
	jxor g4713(.dina(n4772),.dinb(w_n4722_0[2]),.dout(n4773),.clk(gclk));
	jand g4714(.dina(w_n2618_0[0]),.dinb(w_n588_0[0]),.dout(n4774),.clk(gclk));
	jand g4715(.dina(n4774),.dinb(w_n4643_0[0]),.dout(n4775),.clk(gclk));
	jand g4716(.dina(w_n1074_0[2]),.dinb(w_n1033_0[0]),.dout(n4776),.clk(gclk));
	jand g4717(.dina(w_n252_1[2]),.dinb(w_n191_1[0]),.dout(n4777),.clk(gclk));
	jand g4718(.dina(n4777),.dinb(n4776),.dout(n4778),.clk(gclk));
	jand g4719(.dina(n4778),.dinb(w_n4558_0[1]),.dout(n4779),.clk(gclk));
	jand g4720(.dina(n4779),.dinb(w_n334_0[0]),.dout(n4780),.clk(gclk));
	jand g4721(.dina(n4780),.dinb(n4775),.dout(n4781),.clk(gclk));
	jand g4722(.dina(n4781),.dinb(w_n2732_0[0]),.dout(n4782),.clk(gclk));
	jxor g4723(.dina(w_n4782_0[2]),.dinb(w_n4773_0[1]),.dout(n4783),.clk(gclk));
	jxor g4724(.dina(w_n4783_0[1]),.dinb(w_n4719_0[1]),.dout(n4784),.clk(gclk));
	jxor g4725(.dina(w_n4784_0[1]),.dinb(w_n4716_0[1]),.dout(n4785),.clk(gclk));
	jor g4726(.dina(w_n4713_0[0]),.dinb(w_n4712_0[0]),.dout(n4786),.clk(gclk));
	jand g4727(.dina(w_n4786_0[1]),.dinb(w_n4093_9[1]),.dout(n4787),.clk(gclk));
	jxor g4728(.dina(n4787),.dinb(w_n4785_0[1]),.dout(w_dff_A_64zGTwWk3_2),.clk(gclk));
	jand g4729(.dina(w_n4784_0[0]),.dinb(w_n4716_0[0]),.dout(n4789),.clk(gclk));
	jor g4730(.dina(w_n4782_0[1]),.dinb(w_n4773_0[0]),.dout(n4790),.clk(gclk));
	jnot g4731(.din(w_n4790_0[1]),.dout(n4791),.clk(gclk));
	jand g4732(.dina(w_n4783_0[0]),.dinb(w_n4719_0[0]),.dout(n4792),.clk(gclk));
	jor g4733(.dina(n4792),.dinb(n4791),.dout(n4793),.clk(gclk));
	jnot g4734(.din(w_n1188_0[0]),.dout(n4794),.clk(gclk));
	jand g4735(.dina(w_n1984_0[0]),.dinb(w_n1192_0[0]),.dout(n4795),.clk(gclk));
	jand g4736(.dina(n4795),.dinb(n4794),.dout(n4796),.clk(gclk));
	jand g4737(.dina(n4796),.dinb(w_n195_0[2]),.dout(n4797),.clk(gclk));
	jand g4738(.dina(w_n353_0[2]),.dinb(w_n213_1[0]),.dout(n4798),.clk(gclk));
	jand g4739(.dina(n4798),.dinb(w_n2510_0[0]),.dout(n4799),.clk(gclk));
	jand g4740(.dina(w_n377_1[0]),.dinb(w_n182_2[0]),.dout(n4800),.clk(gclk));
	jand g4741(.dina(n4800),.dinb(n4799),.dout(n4801),.clk(gclk));
	jand g4742(.dina(n4801),.dinb(n4797),.dout(n4802),.clk(gclk));
	jand g4743(.dina(w_n387_1[0]),.dinb(w_n235_0[2]),.dout(n4803),.clk(gclk));
	jand g4744(.dina(w_n261_1[0]),.dinb(w_n232_1[1]),.dout(n4804),.clk(gclk));
	jand g4745(.dina(n4804),.dinb(w_n309_0[2]),.dout(n4805),.clk(gclk));
	jand g4746(.dina(n4805),.dinb(n4803),.dout(n4806),.clk(gclk));
	jand g4747(.dina(w_n915_0[0]),.dinb(w_n204_0[2]),.dout(n4807),.clk(gclk));
	jand g4748(.dina(n4807),.dinb(w_n226_1[0]),.dout(n4808),.clk(gclk));
	jand g4749(.dina(n4808),.dinb(w_n350_0[0]),.dout(n4809),.clk(gclk));
	jand g4750(.dina(n4809),.dinb(n4806),.dout(n4810),.clk(gclk));
	jand g4751(.dina(n4810),.dinb(w_n180_0[1]),.dout(n4811),.clk(gclk));
	jand g4752(.dina(w_n4811_0[1]),.dinb(w_n3871_0[0]),.dout(n4812),.clk(gclk));
	jand g4753(.dina(n4812),.dinb(n4802),.dout(n4813),.clk(gclk));
	jnot g4754(.din(w_n4813_0[1]),.dout(n4814),.clk(gclk));
	jand g4755(.dina(w_n4770_0[0]),.dinb(w_n4727_0[0]),.dout(n4815),.clk(gclk));
	jand g4756(.dina(w_n4771_0[1]),.dinb(w_n4722_0[1]),.dout(n4816),.clk(gclk));
	jor g4757(.dina(n4816),.dinb(n4815),.dout(n4817),.clk(gclk));
	jor g4758(.dina(w_n4739_0[0]),.dinb(w_n4731_0[0]),.dout(n4818),.clk(gclk));
	jand g4759(.dina(w_n4769_0[0]),.dinb(w_n4740_0[0]),.dout(n4819),.clk(gclk));
	jnot g4760(.din(n4819),.dout(n4820),.clk(gclk));
	jand g4761(.dina(n4820),.dinb(n4818),.dout(n4821),.clk(gclk));
	jnot g4762(.din(n4821),.dout(n4822),.clk(gclk));
	jand g4763(.dina(w_n4767_0[0]),.dinb(w_n4759_0[0]),.dout(n4823),.clk(gclk));
	jand g4764(.dina(w_n4768_0[0]),.dinb(w_n4743_0[0]),.dout(n4824),.clk(gclk));
	jor g4765(.dina(n4824),.dinb(n4823),.dout(n4825),.clk(gclk));
	jand g4766(.dina(w_n4757_0[0]),.dinb(w_n4749_0[0]),.dout(n4826),.clk(gclk));
	jand g4767(.dina(w_n4758_0[0]),.dinb(w_n4746_0[0]),.dout(n4827),.clk(gclk));
	jor g4768(.dina(n4827),.dinb(n4826),.dout(n4828),.clk(gclk));
	jand g4769(.dina(w_n3143_0[1]),.dinb(w_n1438_11[1]),.dout(n4829),.clk(gclk));
	jnot g4770(.din(w_n4829_0[2]),.dout(n4830),.clk(gclk));
	jand g4771(.dina(w_n3023_3[1]),.dinb(w_n1156_4[0]),.dout(n4831),.clk(gclk));
	jand g4772(.dina(w_n4748_0[0]),.dinb(w_n4747_0[0]),.dout(n4832),.clk(gclk));
	jor g4773(.dina(n4832),.dinb(n4831),.dout(n4833),.clk(gclk));
	jxor g4774(.dina(w_n4833_0[1]),.dinb(w_n4830_0[1]),.dout(n4834),.clk(gclk));
	jor g4775(.dina(w_n3579_0[1]),.dinb(w_n3384_4[1]),.dout(n4835),.clk(gclk));
	jor g4776(.dina(w_n3495_3[1]),.dinb(w_n3386_2[2]),.dout(n4836),.clk(gclk));
	jor g4777(.dina(w_n3203_2[2]),.dinb(w_n3388_3[0]),.dout(n4837),.clk(gclk));
	jor g4778(.dina(w_n3441_2[1]),.dinb(w_n3390_3[0]),.dout(n4838),.clk(gclk));
	jand g4779(.dina(n4838),.dinb(n4837),.dout(n4839),.clk(gclk));
	jand g4780(.dina(n4839),.dinb(n4836),.dout(n4840),.clk(gclk));
	jand g4781(.dina(n4840),.dinb(n4835),.dout(n4841),.clk(gclk));
	jxor g4782(.dina(n4841),.dinb(w_n2051_4[0]),.dout(n4842),.clk(gclk));
	jxor g4783(.dina(w_n4842_0[1]),.dinb(w_n4834_0[1]),.dout(n4843),.clk(gclk));
	jxor g4784(.dina(w_n4843_0[1]),.dinb(w_n4828_0[1]),.dout(n4844),.clk(gclk));
	jnot g4785(.din(n4844),.dout(n4845),.clk(gclk));
	jor g4786(.dina(w_n3842_0[2]),.dinb(w_n2252_3[1]),.dout(n4846),.clk(gclk));
	jor g4787(.dina(w_n3547_3[2]),.dinb(w_n2359_3[1]),.dout(n4847),.clk(gclk));
	jor g4788(.dina(w_n3837_4[1]),.dinb(w_n2355_3[0]),.dout(n4848),.clk(gclk));
	jand g4789(.dina(n4848),.dinb(n4847),.dout(n4849),.clk(gclk));
	jor g4790(.dina(w_n3510_4[0]),.dinb(w_n2357_3[1]),.dout(n4850),.clk(gclk));
	jand g4791(.dina(n4850),.dinb(n4849),.dout(n4851),.clk(gclk));
	jand g4792(.dina(n4851),.dinb(n4846),.dout(n4852),.clk(gclk));
	jxor g4793(.dina(n4852),.dinb(w_n1356_4[2]),.dout(n4853),.clk(gclk));
	jxor g4794(.dina(w_n4853_0[1]),.dinb(w_n4845_0[1]),.dout(n4854),.clk(gclk));
	jxor g4795(.dina(w_n4854_0[1]),.dinb(w_n4825_0[1]),.dout(n4855),.clk(gclk));
	jor g4796(.dina(w_n4349_1[0]),.dinb(w_n2506_2[1]),.dout(n4856),.clk(gclk));
	jor g4797(.dina(w_n4063_5[0]),.dinb(w_n2816_2[1]),.dout(n4857),.clk(gclk));
	jor g4798(.dina(w_n4213_3[2]),.dinb(w_n2807_2[1]),.dout(n4858),.clk(gclk));
	jand g4799(.dina(n4858),.dinb(n4857),.dout(n4859),.clk(gclk));
	jand g4800(.dina(n4859),.dinb(n4856),.dout(n4860),.clk(gclk));
	jxor g4801(.dina(n4860),.dinb(w_n1259_4[1]),.dout(n4861),.clk(gclk));
	jxor g4802(.dina(w_n4861_0[1]),.dinb(w_n4855_0[1]),.dout(n4862),.clk(gclk));
	jxor g4803(.dina(w_n4862_0[1]),.dinb(w_n4822_0[1]),.dout(n4863),.clk(gclk));
	jxor g4804(.dina(w_n4863_0[1]),.dinb(w_n4817_0[1]),.dout(n4864),.clk(gclk));
	jxor g4805(.dina(w_n4864_0[2]),.dinb(w_n4814_0[1]),.dout(n4865),.clk(gclk));
	jxor g4806(.dina(w_n4865_0[1]),.dinb(w_n4793_0[1]),.dout(n4866),.clk(gclk));
	jxor g4807(.dina(w_n4866_0[1]),.dinb(w_n4789_0[1]),.dout(n4867),.clk(gclk));
	jor g4808(.dina(w_n4786_0[0]),.dinb(w_n4785_0[0]),.dout(n4868),.clk(gclk));
	jand g4809(.dina(w_n4868_0[1]),.dinb(w_n4093_9[0]),.dout(n4869),.clk(gclk));
	jxor g4810(.dina(n4869),.dinb(w_n4867_0[1]),.dout(w_dff_A_xitZ0m6h4_2),.clk(gclk));
	jand g4811(.dina(w_n4866_0[0]),.dinb(w_n4789_0[0]),.dout(n4871),.clk(gclk));
	jand g4812(.dina(w_n4864_0[1]),.dinb(w_n4814_0[0]),.dout(n4872),.clk(gclk));
	jand g4813(.dina(w_n4865_0[0]),.dinb(w_n4793_0[0]),.dout(n4873),.clk(gclk));
	jor g4814(.dina(n4873),.dinb(w_n4872_0[1]),.dout(n4874),.clk(gclk));
	jand g4815(.dina(w_n3470_0[0]),.dinb(w_n226_0[2]),.dout(n4875),.clk(gclk));
	jand g4816(.dina(w_n1005_1[2]),.dinb(w_n587_1[0]),.dout(n4876),.clk(gclk));
	jand g4817(.dina(w_n346_1[0]),.dinb(w_n160_0[2]),.dout(n4877),.clk(gclk));
	jand g4818(.dina(n4877),.dinb(n4876),.dout(n4878),.clk(gclk));
	jand g4819(.dina(w_n3537_1[0]),.dinb(w_n1074_0[1]),.dout(n4879),.clk(gclk));
	jand g4820(.dina(n4879),.dinb(n4878),.dout(n4880),.clk(gclk));
	jand g4821(.dina(w_n255_0[2]),.dinb(w_n244_1[1]),.dout(n4881),.clk(gclk));
	jand g4822(.dina(n4881),.dinb(w_n1021_0[0]),.dout(n4882),.clk(gclk));
	jand g4823(.dina(n4882),.dinb(n4880),.dout(n4883),.clk(gclk));
	jand g4824(.dina(n4883),.dinb(n4875),.dout(n4884),.clk(gclk));
	jand g4825(.dina(n4884),.dinb(w_n320_0[0]),.dout(n4885),.clk(gclk));
	jand g4826(.dina(n4885),.dinb(w_n2146_0[0]),.dout(n4886),.clk(gclk));
	jnot g4827(.din(w_n4886_0[1]),.dout(n4887),.clk(gclk));
	jand g4828(.dina(w_n4862_0[0]),.dinb(w_n4822_0[0]),.dout(n4888),.clk(gclk));
	jand g4829(.dina(w_n4863_0[0]),.dinb(w_n4817_0[0]),.dout(n4889),.clk(gclk));
	jor g4830(.dina(n4889),.dinb(n4888),.dout(n4890),.clk(gclk));
	jand g4831(.dina(w_n4854_0[0]),.dinb(w_n4825_0[0]),.dout(n4891),.clk(gclk));
	jand g4832(.dina(w_n4861_0[0]),.dinb(w_n4855_0[0]),.dout(n4892),.clk(gclk));
	jor g4833(.dina(n4892),.dinb(n4891),.dout(n4893),.clk(gclk));
	jand g4834(.dina(w_n4843_0[0]),.dinb(w_n4828_0[0]),.dout(n4894),.clk(gclk));
	jnot g4835(.din(n4894),.dout(n4895),.clk(gclk));
	jor g4836(.dina(w_n4853_0[0]),.dinb(w_n4845_0[0]),.dout(n4896),.clk(gclk));
	jand g4837(.dina(n4896),.dinb(n4895),.dout(n4897),.clk(gclk));
	jand g4838(.dina(w_n4338_1[0]),.dinb(w_n2815_0[0]),.dout(n4898),.clk(gclk));
	jand g4839(.dina(w_n4343_1[1]),.dinb(w_n2505_0[1]),.dout(n4899),.clk(gclk));
	jor g4840(.dina(n4899),.dinb(n4898),.dout(n4900),.clk(gclk));
	jxor g4841(.dina(n4900),.dinb(w_n1259_4[0]),.dout(n4901),.clk(gclk));
	jxor g4842(.dina(w_n4901_0[1]),.dinb(w_n4897_0[1]),.dout(n4902),.clk(gclk));
	jand g4843(.dina(w_n4833_0[0]),.dinb(w_n4830_0[0]),.dout(n4903),.clk(gclk));
	jand g4844(.dina(w_n4842_0[0]),.dinb(w_n4834_0[0]),.dout(n4904),.clk(gclk));
	jor g4845(.dina(n4904),.dinb(n4903),.dout(n4905),.clk(gclk));
	jor g4846(.dina(w_n3566_0[1]),.dinb(w_n3384_4[0]),.dout(n4906),.clk(gclk));
	jand g4847(.dina(w_n3520_0[1]),.dinb(w_n2488_1[0]),.dout(n4907),.clk(gclk));
	jnot g4848(.din(w_n3510_3[2]),.dout(n4908),.clk(gclk));
	jand g4849(.dina(w_n4908_0[1]),.dinb(w_n2491_1[0]),.dout(n4909),.clk(gclk));
	jor g4850(.dina(n4909),.dinb(n4907),.dout(n4910),.clk(gclk));
	jand g4851(.dina(w_n3513_0[2]),.dinb(w_n2923_1[1]),.dout(n4911),.clk(gclk));
	jor g4852(.dina(n4911),.dinb(n4910),.dout(n4912),.clk(gclk));
	jnot g4853(.din(n4912),.dout(n4913),.clk(gclk));
	jand g4854(.dina(n4913),.dinb(n4906),.dout(n4914),.clk(gclk));
	jand g4855(.dina(w_n3418_0[0]),.dinb(w_n1438_11[0]),.dout(n4915),.clk(gclk));
	jxor g4856(.dina(w_n4915_0[1]),.dinb(w_n4914_0[2]),.dout(n4916),.clk(gclk));
	jxor g4857(.dina(w_n4916_0[1]),.dinb(w_n4905_0[1]),.dout(n4917),.clk(gclk));
	jnot g4858(.din(n4917),.dout(n4918),.clk(gclk));
	jor g4859(.dina(w_n4066_0[2]),.dinb(w_n2252_3[0]),.dout(n4919),.clk(gclk));
	jor g4860(.dina(w_n3837_4[0]),.dinb(w_n2359_3[0]),.dout(n4920),.clk(gclk));
	jor g4861(.dina(w_n4063_4[2]),.dinb(w_n2355_2[2]),.dout(n4921),.clk(gclk));
	jand g4862(.dina(n4921),.dinb(n4920),.dout(n4922),.clk(gclk));
	jor g4863(.dina(w_n3547_3[1]),.dinb(w_n2357_3[0]),.dout(n4923),.clk(gclk));
	jand g4864(.dina(n4923),.dinb(n4922),.dout(n4924),.clk(gclk));
	jand g4865(.dina(n4924),.dinb(n4919),.dout(n4925),.clk(gclk));
	jxor g4866(.dina(n4925),.dinb(w_n1356_4[1]),.dout(n4926),.clk(gclk));
	jxor g4867(.dina(w_n4926_0[1]),.dinb(w_n4918_0[1]),.dout(n4927),.clk(gclk));
	jxor g4868(.dina(w_n4927_0[1]),.dinb(w_n4902_0[1]),.dout(n4928),.clk(gclk));
	jxor g4869(.dina(w_n4928_0[1]),.dinb(w_n4893_0[1]),.dout(n4929),.clk(gclk));
	jxor g4870(.dina(w_n4929_0[1]),.dinb(w_n4890_0[1]),.dout(n4930),.clk(gclk));
	jxor g4871(.dina(w_n4930_0[2]),.dinb(w_n4887_0[1]),.dout(n4931),.clk(gclk));
	jxor g4872(.dina(w_n4931_0[1]),.dinb(w_n4874_0[1]),.dout(n4932),.clk(gclk));
	jxor g4873(.dina(w_n4932_0[1]),.dinb(w_n4871_0[1]),.dout(n4933),.clk(gclk));
	jor g4874(.dina(w_n4868_0[0]),.dinb(w_n4867_0[0]),.dout(n4934),.clk(gclk));
	jand g4875(.dina(w_n4934_0[1]),.dinb(w_n4093_8[2]),.dout(n4935),.clk(gclk));
	jxor g4876(.dina(n4935),.dinb(w_n4933_0[1]),.dout(w_dff_A_8Yxnvs8b7_2),.clk(gclk));
	jand g4877(.dina(w_n4932_0[0]),.dinb(w_n4871_0[0]),.dout(n4937),.clk(gclk));
	jand g4878(.dina(w_n4930_0[1]),.dinb(w_n4887_0[0]),.dout(n4938),.clk(gclk));
	jand g4879(.dina(w_n4931_0[0]),.dinb(w_n4874_0[0]),.dout(n4939),.clk(gclk));
	jor g4880(.dina(n4939),.dinb(w_n4938_0[1]),.dout(n4940),.clk(gclk));
	jand g4881(.dina(w_n497_0[1]),.dinb(w_n198_0[2]),.dout(n4941),.clk(gclk));
	jand g4882(.dina(w_n3537_0[2]),.dinb(w_n352_0[1]),.dout(n4942),.clk(gclk));
	jand g4883(.dina(n4942),.dinb(n4941),.dout(n4943),.clk(gclk));
	jand g4884(.dina(n4943),.dinb(w_n1387_0[0]),.dout(n4944),.clk(gclk));
	jand g4885(.dina(w_n534_1[0]),.dinb(w_n190_0[1]),.dout(n4945),.clk(gclk));
	jand g4886(.dina(n4945),.dinb(w_n297_0[1]),.dout(n4946),.clk(gclk));
	jnot g4887(.din(w_n1186_0[0]),.dout(n4947),.clk(gclk));
	jand g4888(.dina(n4947),.dinb(w_n506_0[2]),.dout(n4948),.clk(gclk));
	jand g4889(.dina(n4948),.dinb(n4946),.dout(n4949),.clk(gclk));
	jand g4890(.dina(n4949),.dinb(w_n3881_0[0]),.dout(n4950),.clk(gclk));
	jand g4891(.dina(n4950),.dinb(w_n896_0[0]),.dout(n4951),.clk(gclk));
	jand g4892(.dina(n4951),.dinb(n4944),.dout(n4952),.clk(gclk));
	jnot g4893(.din(w_n4952_0[1]),.dout(n4953),.clk(gclk));
	jand g4894(.dina(w_n4928_0[0]),.dinb(w_n4893_0[0]),.dout(n4954),.clk(gclk));
	jand g4895(.dina(w_n4929_0[0]),.dinb(w_n4890_0[0]),.dout(n4955),.clk(gclk));
	jor g4896(.dina(n4955),.dinb(n4954),.dout(n4956),.clk(gclk));
	jor g4897(.dina(w_n4901_0[0]),.dinb(w_n4897_0[0]),.dout(n4957),.clk(gclk));
	jand g4898(.dina(w_n4927_0[0]),.dinb(w_n4902_0[0]),.dout(n4958),.clk(gclk));
	jnot g4899(.din(n4958),.dout(n4959),.clk(gclk));
	jand g4900(.dina(n4959),.dinb(n4957),.dout(n4960),.clk(gclk));
	jnot g4901(.din(n4960),.dout(n4961),.clk(gclk));
	jor g4902(.dina(w_n4914_0[1]),.dinb(w_n1438_10[2]),.dout(n4962),.clk(gclk));
	jand g4903(.dina(w_n4915_0[0]),.dinb(w_n4914_0[0]),.dout(n4963),.clk(gclk));
	jand g4904(.dina(w_n3415_0[1]),.dinb(w_n1438_10[1]),.dout(n4964),.clk(gclk));
	jand g4905(.dina(n4964),.dinb(w_n3166_2[2]),.dout(n4965),.clk(gclk));
	jor g4906(.dina(n4965),.dinb(n4963),.dout(n4966),.clk(gclk));
	jnot g4907(.din(n4966),.dout(n4967),.clk(gclk));
	jand g4908(.dina(n4967),.dinb(n4962),.dout(n4968),.clk(gclk));
	jnot g4909(.din(n4968),.dout(n4969),.clk(gclk));
	jand g4910(.dina(w_n3513_0[1]),.dinb(w_n1438_10[0]),.dout(n4970),.clk(gclk));
	jxor g4911(.dina(w_n4970_0[2]),.dinb(w_n1259_3[2]),.dout(n4971),.clk(gclk));
	jxor g4912(.dina(n4971),.dinb(w_n4829_0[1]),.dout(n4972),.clk(gclk));
	jxor g4913(.dina(w_n4972_0[1]),.dinb(w_n4969_0[1]),.dout(n4973),.clk(gclk));
	jnot g4914(.din(n4973),.dout(n4974),.clk(gclk));
	jor g4915(.dina(w_n3550_0[1]),.dinb(w_n3384_3[2]),.dout(n4975),.clk(gclk));
	jor g4916(.dina(w_n3547_3[0]),.dinb(w_n3386_2[1]),.dout(n4976),.clk(gclk));
	jor g4917(.dina(w_n3510_3[1]),.dinb(w_n3390_2[2]),.dout(n4977),.clk(gclk));
	jor g4918(.dina(w_n3495_3[0]),.dinb(w_n3388_2[2]),.dout(n4978),.clk(gclk));
	jand g4919(.dina(n4978),.dinb(n4977),.dout(n4979),.clk(gclk));
	jand g4920(.dina(n4979),.dinb(n4976),.dout(n4980),.clk(gclk));
	jand g4921(.dina(n4980),.dinb(n4975),.dout(n4981),.clk(gclk));
	jxor g4922(.dina(n4981),.dinb(w_n1438_9[2]),.dout(n4982),.clk(gclk));
	jxor g4923(.dina(w_n4982_0[1]),.dinb(w_n4974_0[1]),.dout(n4983),.clk(gclk));
	jand g4924(.dina(w_n4916_0[0]),.dinb(w_n4905_0[0]),.dout(n4984),.clk(gclk));
	jnot g4925(.din(n4984),.dout(n4985),.clk(gclk));
	jor g4926(.dina(w_n4926_0[0]),.dinb(w_n4918_0[0]),.dout(n4986),.clk(gclk));
	jand g4927(.dina(n4986),.dinb(n4985),.dout(n4987),.clk(gclk));
	jnot g4928(.din(n4987),.dout(n4988),.clk(gclk));
	jor g4929(.dina(w_n4215_0[2]),.dinb(w_n2252_2[2]),.dout(n4989),.clk(gclk));
	jor g4930(.dina(w_n4213_3[1]),.dinb(w_n2355_2[1]),.dout(n4990),.clk(gclk));
	jor g4931(.dina(w_n3837_3[2]),.dinb(w_n2357_2[2]),.dout(n4991),.clk(gclk));
	jand g4932(.dina(n4991),.dinb(n4990),.dout(n4992),.clk(gclk));
	jor g4933(.dina(w_n4063_4[1]),.dinb(w_n2359_2[2]),.dout(n4993),.clk(gclk));
	jand g4934(.dina(n4993),.dinb(n4992),.dout(n4994),.clk(gclk));
	jand g4935(.dina(n4994),.dinb(n4989),.dout(n4995),.clk(gclk));
	jxor g4936(.dina(n4995),.dinb(w_n1480_4[1]),.dout(n4996),.clk(gclk));
	jxor g4937(.dina(w_n4996_0[1]),.dinb(w_n4988_0[1]),.dout(n4997),.clk(gclk));
	jxor g4938(.dina(w_n4997_0[1]),.dinb(w_n4983_0[1]),.dout(n4998),.clk(gclk));
	jxor g4939(.dina(w_n4998_0[1]),.dinb(w_n4961_0[1]),.dout(n4999),.clk(gclk));
	jxor g4940(.dina(w_n4999_0[1]),.dinb(w_n4956_0[1]),.dout(n5000),.clk(gclk));
	jxor g4941(.dina(w_n5000_0[2]),.dinb(w_n4953_0[1]),.dout(n5001),.clk(gclk));
	jxor g4942(.dina(w_n5001_0[1]),.dinb(w_n4940_0[1]),.dout(n5002),.clk(gclk));
	jxor g4943(.dina(w_n5002_0[1]),.dinb(w_n4937_0[1]),.dout(n5003),.clk(gclk));
	jor g4944(.dina(w_n4934_0[0]),.dinb(w_n4933_0[0]),.dout(n5004),.clk(gclk));
	jand g4945(.dina(w_n5004_0[1]),.dinb(w_n4093_8[1]),.dout(n5005),.clk(gclk));
	jxor g4946(.dina(n5005),.dinb(w_n5003_0[1]),.dout(w_dff_A_xTdiVglx2_2),.clk(gclk));
	jand g4947(.dina(w_n5002_0[0]),.dinb(w_n4937_0[0]),.dout(n5007),.clk(gclk));
	jand g4948(.dina(w_n5000_0[1]),.dinb(w_n4953_0[0]),.dout(n5008),.clk(gclk));
	jand g4949(.dina(w_n5001_0[0]),.dinb(w_n4940_0[0]),.dout(n5009),.clk(gclk));
	jor g4950(.dina(n5009),.dinb(w_n5008_0[1]),.dout(n5010),.clk(gclk));
	jand g4951(.dina(w_n816_0[0]),.dinb(w_n717_1[1]),.dout(n5011),.clk(gclk));
	jand g4952(.dina(n5011),.dinb(w_n459_0[0]),.dout(n5012),.clk(gclk));
	jand g4953(.dina(n5012),.dinb(w_n4051_0[0]),.dout(n5013),.clk(gclk));
	jand g4954(.dina(w_n827_0[0]),.dinb(w_n509_0[0]),.dout(n5014),.clk(gclk));
	jand g4955(.dina(n5014),.dinb(n5013),.dout(n5015),.clk(gclk));
	jand g4956(.dina(n5015),.dinb(w_n1381_0[0]),.dout(n5016),.clk(gclk));
	jnot g4957(.din(w_n5016_0[1]),.dout(n5017),.clk(gclk));
	jand g4958(.dina(w_n4998_0[0]),.dinb(w_n4961_0[0]),.dout(n5018),.clk(gclk));
	jand g4959(.dina(w_n4999_0[0]),.dinb(w_n4956_0[0]),.dout(n5019),.clk(gclk));
	jor g4960(.dina(n5019),.dinb(n5018),.dout(n5020),.clk(gclk));
	jand g4961(.dina(w_n4996_0[0]),.dinb(w_n4988_0[0]),.dout(n5021),.clk(gclk));
	jand g4962(.dina(w_n4997_0[0]),.dinb(w_n4983_0[0]),.dout(n5022),.clk(gclk));
	jor g4963(.dina(n5022),.dinb(n5021),.dout(n5023),.clk(gclk));
	jand g4964(.dina(w_n4972_0[0]),.dinb(w_n4969_0[0]),.dout(n5024),.clk(gclk));
	jnot g4965(.din(n5024),.dout(n5025),.clk(gclk));
	jor g4966(.dina(w_n4982_0[0]),.dinb(w_n4974_0[0]),.dout(n5026),.clk(gclk));
	jand g4967(.dina(n5026),.dinb(n5025),.dout(n5027),.clk(gclk));
	jnot g4968(.din(n5027),.dout(n5028),.clk(gclk));
	jand g4969(.dina(w_n3520_0[0]),.dinb(w_n1438_9[1]),.dout(n5029),.clk(gclk));
	jnot g4970(.din(w_n5029_0[1]),.dout(n5030),.clk(gclk));
	jor g4971(.dina(w_n4970_0[1]),.dinb(w_n1259_3[1]),.dout(n5031),.clk(gclk));
	jand g4972(.dina(w_n4970_0[0]),.dinb(w_n1259_3[0]),.dout(n5032),.clk(gclk));
	jor g4973(.dina(n5032),.dinb(w_n4829_0[0]),.dout(n5033),.clk(gclk));
	jand g4974(.dina(n5033),.dinb(n5031),.dout(n5034),.clk(gclk));
	jxor g4975(.dina(w_n5034_0[1]),.dinb(w_n5030_0[1]),.dout(n5035),.clk(gclk));
	jor g4976(.dina(w_n3842_0[1]),.dinb(w_n3384_3[1]),.dout(n5036),.clk(gclk));
	jor g4977(.dina(w_n3837_3[1]),.dinb(w_n3386_2[0]),.dout(n5037),.clk(gclk));
	jor g4978(.dina(w_n3547_2[2]),.dinb(w_n3390_2[1]),.dout(n5038),.clk(gclk));
	jor g4979(.dina(w_n3510_3[0]),.dinb(w_n3388_2[1]),.dout(n5039),.clk(gclk));
	jand g4980(.dina(n5039),.dinb(n5038),.dout(n5040),.clk(gclk));
	jand g4981(.dina(n5040),.dinb(n5037),.dout(n5041),.clk(gclk));
	jand g4982(.dina(n5041),.dinb(n5036),.dout(n5042),.clk(gclk));
	jxor g4983(.dina(n5042),.dinb(w_n2051_3[2]),.dout(n5043),.clk(gclk));
	jxor g4984(.dina(w_n5043_0[1]),.dinb(w_n5035_0[1]),.dout(n5044),.clk(gclk));
	jxor g4985(.dina(w_n5044_0[1]),.dinb(w_n5028_0[1]),.dout(n5045),.clk(gclk));
	jor g4986(.dina(w_n4349_0[2]),.dinb(w_n2252_2[1]),.dout(n5046),.clk(gclk));
	jor g4987(.dina(w_n4063_4[0]),.dinb(w_n2357_2[1]),.dout(n5047),.clk(gclk));
	jor g4988(.dina(w_n4213_3[0]),.dinb(w_n2359_2[1]),.dout(n5048),.clk(gclk));
	jand g4989(.dina(n5048),.dinb(n5047),.dout(n5049),.clk(gclk));
	jand g4990(.dina(n5049),.dinb(n5046),.dout(n5050),.clk(gclk));
	jxor g4991(.dina(n5050),.dinb(w_n1480_4[0]),.dout(n5051),.clk(gclk));
	jxor g4992(.dina(w_n5051_0[1]),.dinb(w_n5045_0[1]),.dout(n5052),.clk(gclk));
	jxor g4993(.dina(w_n5052_0[1]),.dinb(w_n5023_0[1]),.dout(n5053),.clk(gclk));
	jxor g4994(.dina(w_n5053_0[1]),.dinb(w_n5020_0[1]),.dout(n5054),.clk(gclk));
	jxor g4995(.dina(w_n5054_0[2]),.dinb(w_n5017_0[1]),.dout(n5055),.clk(gclk));
	jxor g4996(.dina(w_n5055_0[1]),.dinb(w_n5010_0[1]),.dout(n5056),.clk(gclk));
	jxor g4997(.dina(w_n5056_0[1]),.dinb(w_n5007_0[1]),.dout(n5057),.clk(gclk));
	jor g4998(.dina(w_n5004_0[0]),.dinb(w_n5003_0[0]),.dout(n5058),.clk(gclk));
	jand g4999(.dina(w_n5058_0[1]),.dinb(w_n4093_8[0]),.dout(n5059),.clk(gclk));
	jxor g5000(.dina(n5059),.dinb(w_n5057_0[1]),.dout(w_dff_A_aayeK3ua3_2),.clk(gclk));
	jand g5001(.dina(w_n5056_0[0]),.dinb(w_n5007_0[0]),.dout(n5061),.clk(gclk));
	jand g5002(.dina(w_n5054_0[1]),.dinb(w_n5017_0[0]),.dout(n5062),.clk(gclk));
	jand g5003(.dina(w_n5055_0[0]),.dinb(w_n5010_0[0]),.dout(n5063),.clk(gclk));
	jor g5004(.dina(n5063),.dinb(w_n5062_0[1]),.dout(n5064),.clk(gclk));
	jand g5005(.dina(w_n2395_0[1]),.dinb(w_n261_0[2]),.dout(n5065),.clk(gclk));
	jand g5006(.dina(n5065),.dinb(w_n2971_0[0]),.dout(n5066),.clk(gclk));
	jand g5007(.dina(w_n331_0[2]),.dinb(w_n182_1[2]),.dout(n5067),.clk(gclk));
	jand g5008(.dina(w_n313_0[1]),.dinb(w_n278_0[1]),.dout(n5068),.clk(gclk));
	jand g5009(.dina(n5068),.dinb(w_n244_1[0]),.dout(n5069),.clk(gclk));
	jand g5010(.dina(n5069),.dinb(n5067),.dout(n5070),.clk(gclk));
	jand g5011(.dina(w_n5070_0[1]),.dinb(w_n4266_0[0]),.dout(n5071),.clk(gclk));
	jand g5012(.dina(w_n568_0[0]),.dinb(w_n166_1[0]),.dout(n5072),.clk(gclk));
	jand g5013(.dina(n5072),.dinb(w_n157_1[0]),.dout(n5073),.clk(gclk));
	jand g5014(.dina(n5073),.dinb(n5071),.dout(n5074),.clk(gclk));
	jand g5015(.dina(n5074),.dinb(w_n2384_0[0]),.dout(n5075),.clk(gclk));
	jand g5016(.dina(n5075),.dinb(n5066),.dout(n5076),.clk(gclk));
	jnot g5017(.din(w_n5076_0[1]),.dout(n5077),.clk(gclk));
	jand g5018(.dina(w_n5052_0[0]),.dinb(w_n5023_0[0]),.dout(n5078),.clk(gclk));
	jand g5019(.dina(w_n5053_0[0]),.dinb(w_n5020_0[0]),.dout(n5079),.clk(gclk));
	jor g5020(.dina(n5079),.dinb(n5078),.dout(n5080),.clk(gclk));
	jand g5021(.dina(w_n5044_0[0]),.dinb(w_n5028_0[0]),.dout(n5081),.clk(gclk));
	jand g5022(.dina(w_n5051_0[0]),.dinb(w_n5045_0[0]),.dout(n5082),.clk(gclk));
	jor g5023(.dina(n5082),.dinb(n5081),.dout(n5083),.clk(gclk));
	jand g5024(.dina(w_n4338_0[2]),.dinb(w_n2244_0[0]),.dout(n5084),.clk(gclk));
	jand g5025(.dina(w_n4343_1[0]),.dinb(w_n2101_0[1]),.dout(n5085),.clk(gclk));
	jor g5026(.dina(n5085),.dinb(n5084),.dout(n5086),.clk(gclk));
	jxor g5027(.dina(n5086),.dinb(w_n1356_4[0]),.dout(n5087),.clk(gclk));
	jnot g5028(.din(n5087),.dout(n5088),.clk(gclk));
	jor g5029(.dina(w_n4066_0[1]),.dinb(w_n3384_3[0]),.dout(n5089),.clk(gclk));
	jor g5030(.dina(w_n3547_2[1]),.dinb(w_n3388_2[0]),.dout(n5090),.clk(gclk));
	jor g5031(.dina(w_n3837_3[0]),.dinb(w_n3390_2[0]),.dout(n5091),.clk(gclk));
	jor g5032(.dina(w_n4063_3[2]),.dinb(w_n3386_1[2]),.dout(n5092),.clk(gclk));
	jand g5033(.dina(n5092),.dinb(n5091),.dout(n5093),.clk(gclk));
	jand g5034(.dina(n5093),.dinb(n5090),.dout(n5094),.clk(gclk));
	jand g5035(.dina(n5094),.dinb(n5089),.dout(n5095),.clk(gclk));
	jxor g5036(.dina(n5095),.dinb(w_n1438_9[0]),.dout(n5096),.clk(gclk));
	jxor g5037(.dina(w_n5096_0[1]),.dinb(w_n5088_0[1]),.dout(n5097),.clk(gclk));
	jand g5038(.dina(w_n5034_0[0]),.dinb(w_n5030_0[0]),.dout(n5098),.clk(gclk));
	jand g5039(.dina(w_n5043_0[0]),.dinb(w_n5035_0[0]),.dout(n5099),.clk(gclk));
	jor g5040(.dina(n5099),.dinb(n5098),.dout(n5100),.clk(gclk));
	jand g5041(.dina(w_n5029_0[0]),.dinb(w_n3510_2[2]),.dout(n5101),.clk(gclk));
	jand g5042(.dina(w_n4908_0[0]),.dinb(w_n1438_8[2]),.dout(n5102),.clk(gclk));
	jand g5043(.dina(w_n5102_0[2]),.dinb(w_n3495_2[2]),.dout(n5103),.clk(gclk));
	jor g5044(.dina(n5103),.dinb(w_n5101_0[1]),.dout(n5104),.clk(gclk));
	jnot g5045(.din(n5104),.dout(n5105),.clk(gclk));
	jxor g5046(.dina(w_n5105_0[1]),.dinb(w_n5100_0[1]),.dout(n5106),.clk(gclk));
	jxor g5047(.dina(w_n5106_0[1]),.dinb(w_n5097_0[1]),.dout(n5107),.clk(gclk));
	jxor g5048(.dina(w_n5107_0[1]),.dinb(w_n5083_0[1]),.dout(n5108),.clk(gclk));
	jxor g5049(.dina(w_n5108_0[1]),.dinb(w_n5080_0[1]),.dout(n5109),.clk(gclk));
	jxor g5050(.dina(w_n5109_0[2]),.dinb(w_n5077_0[1]),.dout(n5110),.clk(gclk));
	jxor g5051(.dina(w_n5110_0[1]),.dinb(w_n5064_0[1]),.dout(n5111),.clk(gclk));
	jxor g5052(.dina(w_n5111_0[1]),.dinb(w_n5061_0[1]),.dout(n5112),.clk(gclk));
	jor g5053(.dina(w_n5058_0[0]),.dinb(w_n5057_0[0]),.dout(n5113),.clk(gclk));
	jand g5054(.dina(w_n5113_0[1]),.dinb(w_n4093_7[2]),.dout(n5114),.clk(gclk));
	jxor g5055(.dina(n5114),.dinb(w_n5112_0[1]),.dout(w_dff_A_AXUFYtJ77_2),.clk(gclk));
	jand g5056(.dina(w_n5111_0[0]),.dinb(w_n5061_0[0]),.dout(n5116),.clk(gclk));
	jand g5057(.dina(w_n5109_0[1]),.dinb(w_n5077_0[0]),.dout(n5117),.clk(gclk));
	jand g5058(.dina(w_n5110_0[0]),.dinb(w_n5064_0[0]),.dout(n5118),.clk(gclk));
	jor g5059(.dina(n5118),.dinb(w_n5117_0[1]),.dout(n5119),.clk(gclk));
	jand g5060(.dina(w_n370_1[0]),.dinb(w_n300_1[1]),.dout(n5120),.clk(gclk));
	jand g5061(.dina(w_n2149_0[0]),.dinb(w_n374_1[0]),.dout(n5121),.clk(gclk));
	jand g5062(.dina(n5121),.dinb(n5120),.dout(n5122),.clk(gclk));
	jand g5063(.dina(w_n5122_0[1]),.dinb(w_n4237_0[0]),.dout(n5123),.clk(gclk));
	jand g5064(.dina(n5123),.dinb(w_n415_1[0]),.dout(n5124),.clk(gclk));
	jand g5065(.dina(n5124),.dinb(w_n294_1[0]),.dout(n5125),.clk(gclk));
	jand g5066(.dina(n5125),.dinb(w_n3892_0[0]),.dout(n5126),.clk(gclk));
	jand g5067(.dina(w_n446_0[2]),.dinb(w_n276_1[0]),.dout(n5127),.clk(gclk));
	jand g5068(.dina(n5127),.dinb(w_n1025_0[0]),.dout(n5128),.clk(gclk));
	jand g5069(.dina(n5128),.dinb(w_n884_0[2]),.dout(n5129),.clk(gclk));
	jand g5070(.dina(w_n570_0[2]),.dinb(w_n137_0[2]),.dout(n5130),.clk(gclk));
	jand g5071(.dina(n5130),.dinb(n5129),.dout(n5131),.clk(gclk));
	jand g5072(.dina(w_n3106_0[0]),.dinb(w_n912_0[0]),.dout(n5132),.clk(gclk));
	jand g5073(.dina(n5132),.dinb(n5131),.dout(n5133),.clk(gclk));
	jand g5074(.dina(n5133),.dinb(n5126),.dout(n5134),.clk(gclk));
	jnot g5075(.din(w_n5134_0[1]),.dout(n5135),.clk(gclk));
	jand g5076(.dina(w_n5107_0[0]),.dinb(w_n5083_0[0]),.dout(n5136),.clk(gclk));
	jand g5077(.dina(w_n5108_0[0]),.dinb(w_n5080_0[0]),.dout(n5137),.clk(gclk));
	jor g5078(.dina(n5137),.dinb(n5136),.dout(n5138),.clk(gclk));
	jor g5079(.dina(w_n5096_0[0]),.dinb(w_n5088_0[0]),.dout(n5139),.clk(gclk));
	jand g5080(.dina(w_n5106_0[0]),.dinb(w_n5097_0[0]),.dout(n5140),.clk(gclk));
	jnot g5081(.din(n5140),.dout(n5141),.clk(gclk));
	jand g5082(.dina(n5141),.dinb(n5139),.dout(n5142),.clk(gclk));
	jnot g5083(.din(n5142),.dout(n5143),.clk(gclk));
	jand g5084(.dina(w_n5105_0[0]),.dinb(w_n5100_0[0]),.dout(n5144),.clk(gclk));
	jor g5085(.dina(n5144),.dinb(w_n5101_0[0]),.dout(n5145),.clk(gclk));
	jxor g5086(.dina(w_n5102_0[1]),.dinb(w_n1480_3[2]),.dout(n5146),.clk(gclk));
	jand g5087(.dina(w_n3825_0[0]),.dinb(w_n1438_8[1]),.dout(n5147),.clk(gclk));
	jxor g5088(.dina(w_n5147_0[1]),.dinb(w_n5146_0[1]),.dout(n5148),.clk(gclk));
	jor g5089(.dina(w_n4215_0[1]),.dinb(w_n3384_2[2]),.dout(n5149),.clk(gclk));
	jor g5090(.dina(w_n4213_2[2]),.dinb(w_n3386_1[1]),.dout(n5150),.clk(gclk));
	jor g5091(.dina(w_n3837_2[2]),.dinb(w_n3388_1[2]),.dout(n5151),.clk(gclk));
	jand g5092(.dina(n5151),.dinb(n5150),.dout(n5152),.clk(gclk));
	jor g5093(.dina(w_n4063_3[1]),.dinb(w_n3390_1[2]),.dout(n5153),.clk(gclk));
	jand g5094(.dina(n5153),.dinb(n5152),.dout(n5154),.clk(gclk));
	jand g5095(.dina(n5154),.dinb(n5149),.dout(n5155),.clk(gclk));
	jxor g5096(.dina(n5155),.dinb(w_n2051_3[1]),.dout(n5156),.clk(gclk));
	jxor g5097(.dina(w_n5156_0[1]),.dinb(w_n5148_0[1]),.dout(n5157),.clk(gclk));
	jxor g5098(.dina(w_n5157_0[1]),.dinb(w_n5145_0[1]),.dout(n5158),.clk(gclk));
	jxor g5099(.dina(w_n5158_0[1]),.dinb(w_n5143_0[1]),.dout(n5159),.clk(gclk));
	jxor g5100(.dina(w_n5159_0[1]),.dinb(w_n5138_0[1]),.dout(n5160),.clk(gclk));
	jxor g5101(.dina(w_n5160_0[2]),.dinb(w_n5135_0[1]),.dout(n5161),.clk(gclk));
	jxor g5102(.dina(w_n5161_0[1]),.dinb(w_n5119_0[1]),.dout(n5162),.clk(gclk));
	jxor g5103(.dina(w_n5162_0[1]),.dinb(w_n5116_0[1]),.dout(n5163),.clk(gclk));
	jor g5104(.dina(w_n5113_0[0]),.dinb(w_n5112_0[0]),.dout(n5164),.clk(gclk));
	jand g5105(.dina(w_n5164_0[1]),.dinb(w_n4093_7[1]),.dout(n5165),.clk(gclk));
	jxor g5106(.dina(n5165),.dinb(w_n5163_0[1]),.dout(w_dff_A_i53FbZmW9_2),.clk(gclk));
	jand g5107(.dina(w_n5162_0[0]),.dinb(w_n5116_0[0]),.dout(n5167),.clk(gclk));
	jand g5108(.dina(w_n5160_0[1]),.dinb(w_n5135_0[0]),.dout(n5168),.clk(gclk));
	jand g5109(.dina(w_n5161_0[0]),.dinb(w_n5119_0[0]),.dout(n5169),.clk(gclk));
	jor g5110(.dina(n5169),.dinb(w_n5168_0[1]),.dout(n5170),.clk(gclk));
	jand g5111(.dina(w_n2155_0[1]),.dinb(w_n290_1[0]),.dout(n5171),.clk(gclk));
	jand g5112(.dina(n5171),.dinb(w_n2395_0[0]),.dout(n5172),.clk(gclk));
	jand g5113(.dina(n5172),.dinb(w_n886_0[1]),.dout(n5173),.clk(gclk));
	jand g5114(.dina(n5173),.dinb(w_n1196_0[1]),.dout(n5174),.clk(gclk));
	jand g5115(.dina(w_n1096_0[0]),.dinb(w_n162_0[2]),.dout(n5175),.clk(gclk));
	jand g5116(.dina(n5175),.dinb(n5174),.dout(n5176),.clk(gclk));
	jnot g5117(.din(w_n1312_0[0]),.dout(n5177),.clk(gclk));
	jand g5118(.dina(w_n717_1[0]),.dinb(w_n430_0[1]),.dout(n5178),.clk(gclk));
	jand g5119(.dina(n5178),.dinb(w_n3537_0[1]),.dout(n5179),.clk(gclk));
	jand g5120(.dina(w_n488_1[1]),.dinb(w_n415_0[2]),.dout(n5180),.clk(gclk));
	jand g5121(.dina(n5180),.dinb(n5179),.dout(n5181),.clk(gclk));
	jand g5122(.dina(n5181),.dinb(n5177),.dout(n5182),.clk(gclk));
	jand g5123(.dina(n5182),.dinb(w_n359_0[0]),.dout(n5183),.clk(gclk));
	jand g5124(.dina(n5183),.dinb(n5176),.dout(n5184),.clk(gclk));
	jnot g5125(.din(w_n5184_0[1]),.dout(n5185),.clk(gclk));
	jand g5126(.dina(w_n5158_0[0]),.dinb(w_n5143_0[0]),.dout(n5186),.clk(gclk));
	jand g5127(.dina(w_n5159_0[0]),.dinb(w_n5138_0[0]),.dout(n5187),.clk(gclk));
	jor g5128(.dina(n5187),.dinb(n5186),.dout(n5188),.clk(gclk));
	jand g5129(.dina(w_n5156_0[0]),.dinb(w_n5148_0[0]),.dout(n5189),.clk(gclk));
	jand g5130(.dina(w_n5157_0[0]),.dinb(w_n5145_0[0]),.dout(n5190),.clk(gclk));
	jor g5131(.dina(n5190),.dinb(n5189),.dout(n5191),.clk(gclk));
	jand g5132(.dina(w_n3838_1[0]),.dinb(w_n1438_8[0]),.dout(n5192),.clk(gclk));
	jnot g5133(.din(n5192),.dout(n5193),.clk(gclk));
	jand g5134(.dina(w_n5102_0[0]),.dinb(w_n1480_3[1]),.dout(n5194),.clk(gclk));
	jand g5135(.dina(w_n5147_0[0]),.dinb(w_n5146_0[0]),.dout(n5195),.clk(gclk));
	jor g5136(.dina(n5195),.dinb(n5194),.dout(n5196),.clk(gclk));
	jxor g5137(.dina(w_n5196_0[1]),.dinb(w_n5193_0[1]),.dout(n5197),.clk(gclk));
	jor g5138(.dina(w_n4349_0[1]),.dinb(w_n3384_2[1]),.dout(n5198),.clk(gclk));
	jor g5139(.dina(w_n4063_3[0]),.dinb(w_n3388_1[1]),.dout(n5199),.clk(gclk));
	jor g5140(.dina(w_n4213_2[1]),.dinb(w_n3390_1[1]),.dout(n5200),.clk(gclk));
	jand g5141(.dina(n5200),.dinb(n5199),.dout(n5201),.clk(gclk));
	jand g5142(.dina(n5201),.dinb(n5198),.dout(n5202),.clk(gclk));
	jxor g5143(.dina(n5202),.dinb(w_n2051_3[0]),.dout(n5203),.clk(gclk));
	jxor g5144(.dina(w_n5203_0[1]),.dinb(w_n5197_0[1]),.dout(n5204),.clk(gclk));
	jxor g5145(.dina(w_n5204_0[1]),.dinb(w_n5191_0[1]),.dout(n5205),.clk(gclk));
	jxor g5146(.dina(w_n5205_0[1]),.dinb(w_n5188_0[1]),.dout(n5206),.clk(gclk));
	jxor g5147(.dina(w_n5206_0[2]),.dinb(w_n5185_0[1]),.dout(n5207),.clk(gclk));
	jxor g5148(.dina(w_n5207_0[1]),.dinb(w_n5170_0[1]),.dout(n5208),.clk(gclk));
	jxor g5149(.dina(w_n5208_0[1]),.dinb(w_n5167_0[1]),.dout(n5209),.clk(gclk));
	jor g5150(.dina(w_n5164_0[0]),.dinb(w_n5163_0[0]),.dout(n5210),.clk(gclk));
	jand g5151(.dina(w_n5210_0[1]),.dinb(w_n4093_7[0]),.dout(n5211),.clk(gclk));
	jxor g5152(.dina(n5211),.dinb(w_n5209_0[1]),.dout(w_dff_A_MRzbRLbX5_2),.clk(gclk));
	jand g5153(.dina(w_n5208_0[0]),.dinb(w_n5167_0[0]),.dout(n5213),.clk(gclk));
	jand g5154(.dina(w_n5206_0[1]),.dinb(w_n5185_0[0]),.dout(n5214),.clk(gclk));
	jand g5155(.dina(w_n5207_0[0]),.dinb(w_n5170_0[0]),.dout(n5215),.clk(gclk));
	jor g5156(.dina(n5215),.dinb(w_n5214_0[1]),.dout(n5216),.clk(gclk));
	jand g5157(.dina(w_n1095_0[2]),.dinb(w_n1005_1[1]),.dout(n5217),.clk(gclk));
	jand g5158(.dina(n5217),.dinb(w_n94_0[2]),.dout(n5218),.clk(gclk));
	jand g5159(.dina(n5218),.dinb(w_n858_0[0]),.dout(n5219),.clk(gclk));
	jand g5160(.dina(w_n2402_0[0]),.dinb(w_n206_0[2]),.dout(n5220),.clk(gclk));
	jand g5161(.dina(w_n2135_0[0]),.dinb(w_n395_0[2]),.dout(n5221),.clk(gclk));
	jand g5162(.dina(n5221),.dinb(w_n2508_0[0]),.dout(n5222),.clk(gclk));
	jand g5163(.dina(w_n346_0[2]),.dinb(w_n222_1[0]),.dout(n5223),.clk(gclk));
	jand g5164(.dina(n5223),.dinb(n5222),.dout(n5224),.clk(gclk));
	jand g5165(.dina(n5224),.dinb(w_n903_0[0]),.dout(n5225),.clk(gclk));
	jand g5166(.dina(w_n5070_0[0]),.dinb(w_n488_1[0]),.dout(n5226),.clk(gclk));
	jand g5167(.dina(n5226),.dinb(n5225),.dout(n5227),.clk(gclk));
	jand g5168(.dina(n5227),.dinb(n5220),.dout(n5228),.clk(gclk));
	jand g5169(.dina(n5228),.dinb(w_n5219_0[1]),.dout(n5229),.clk(gclk));
	jnot g5170(.din(w_n5229_0[1]),.dout(n5230),.clk(gclk));
	jand g5171(.dina(w_n5196_0[0]),.dinb(w_n5193_0[0]),.dout(n5231),.clk(gclk));
	jand g5172(.dina(w_n5203_0[0]),.dinb(w_n5197_0[0]),.dout(n5232),.clk(gclk));
	jor g5173(.dina(n5232),.dinb(n5231),.dout(n5233),.clk(gclk));
	jand g5174(.dina(w_n4338_0[1]),.dinb(w_n2923_1[0]),.dout(n5234),.clk(gclk));
	jand g5175(.dina(w_n4343_0[2]),.dinb(w_n2484_0[1]),.dout(n5235),.clk(gclk));
	jor g5176(.dina(n5235),.dinb(n5234),.dout(n5236),.clk(gclk));
	jand g5177(.dina(w_n4344_0[0]),.dinb(w_n1438_7[2]),.dout(n5237),.clk(gclk));
	jnot g5178(.din(n5237),.dout(n5238),.clk(gclk));
	jxor g5179(.dina(w_n5238_0[1]),.dinb(w_n5236_0[2]),.dout(n5239),.clk(gclk));
	jxor g5180(.dina(w_n5239_0[1]),.dinb(w_n5233_0[1]),.dout(n5240),.clk(gclk));
	jand g5181(.dina(w_n5204_0[0]),.dinb(w_n5191_0[0]),.dout(n5241),.clk(gclk));
	jand g5182(.dina(w_n5205_0[0]),.dinb(w_n5188_0[0]),.dout(n5242),.clk(gclk));
	jor g5183(.dina(n5242),.dinb(n5241),.dout(n5243),.clk(gclk));
	jxor g5184(.dina(w_n5243_0[1]),.dinb(w_n5240_0[1]),.dout(n5244),.clk(gclk));
	jxor g5185(.dina(w_n5244_0[2]),.dinb(w_n5230_0[1]),.dout(n5245),.clk(gclk));
	jxor g5186(.dina(w_n5245_0[1]),.dinb(w_n5216_0[1]),.dout(n5246),.clk(gclk));
	jxor g5187(.dina(w_n5246_0[1]),.dinb(w_n5213_0[1]),.dout(n5247),.clk(gclk));
	jor g5188(.dina(w_n5210_0[0]),.dinb(w_n5209_0[0]),.dout(n5248),.clk(gclk));
	jand g5189(.dina(w_n5248_0[1]),.dinb(w_n4093_6[2]),.dout(n5249),.clk(gclk));
	jxor g5190(.dina(n5249),.dinb(w_n5247_0[1]),.dout(w_dff_A_MetX8NB96_2),.clk(gclk));
	jand g5191(.dina(w_n5246_0[0]),.dinb(w_n5213_0[0]),.dout(n5251),.clk(gclk));
	jnot g5192(.din(n5251),.dout(n5252),.clk(gclk));
	jand g5193(.dina(w_n5244_0[1]),.dinb(w_n5230_0[0]),.dout(n5253),.clk(gclk));
	jnot g5194(.din(w_n5253_0[1]),.dout(n5254),.clk(gclk));
	jnot g5195(.din(w_n5214_0[0]),.dout(n5255),.clk(gclk));
	jnot g5196(.din(w_n5168_0[0]),.dout(n5256),.clk(gclk));
	jnot g5197(.din(w_n5117_0[0]),.dout(n5257),.clk(gclk));
	jnot g5198(.din(w_n5062_0[0]),.dout(n5258),.clk(gclk));
	jnot g5199(.din(w_n5008_0[0]),.dout(n5259),.clk(gclk));
	jnot g5200(.din(w_n4938_0[0]),.dout(n5260),.clk(gclk));
	jnot g5201(.din(w_n4872_0[0]),.dout(n5261),.clk(gclk));
	jnot g5202(.din(w_n4717_0[0]),.dout(n5262),.clk(gclk));
	jnot g5203(.din(w_n4633_0[0]),.dout(n5263),.clk(gclk));
	jnot g5204(.din(w_n4547_0[0]),.dout(n5264),.clk(gclk));
	jnot g5205(.din(w_n4457_0[0]),.dout(n5265),.clk(gclk));
	jnot g5206(.din(w_n4367_0[0]),.dout(n5266),.clk(gclk));
	jnot g5207(.din(w_n3853_0[0]),.dout(n5267),.clk(gclk));
	jxor g5208(.dina(w_n3852_0[0]),.dinb(w_n324_0[0]),.dout(n5268),.clk(gclk));
	jnot g5209(.din(w_n3968_0[0]),.dout(n5269),.clk(gclk));
	jor g5210(.dina(n5269),.dinb(w_n3963_0[0]),.dout(n5270),.clk(gclk));
	jor g5211(.dina(n5270),.dinb(n5268),.dout(n5271),.clk(gclk));
	jand g5212(.dina(n5271),.dinb(n5267),.dout(n5272),.clk(gclk));
	jxor g5213(.dina(w_n4075_0[1]),.dinb(w_n4274_0[0]),.dout(n5273),.clk(gclk));
	jxor g5214(.dina(w_n4088_0[0]),.dinb(n5273),.dout(n5274),.clk(gclk));
	jor g5215(.dina(n5274),.dinb(n5272),.dout(n5275),.clk(gclk));
	jand g5216(.dina(n5275),.dinb(w_n4097_0[0]),.dout(n5276),.clk(gclk));
	jxor g5217(.dina(w_n4226_0[0]),.dinb(w_n4276_0[0]),.dout(n5277),.clk(gclk));
	jxor g5218(.dina(w_n4242_0[0]),.dinb(n5277),.dout(n5278),.clk(gclk));
	jor g5219(.dina(n5278),.dinb(n5276),.dout(n5279),.clk(gclk));
	jand g5220(.dina(n5279),.dinb(w_n4251_0[0]),.dout(n5280),.clk(gclk));
	jxor g5221(.dina(w_n4357_0[0]),.dinb(w_n4270_0[0]),.dout(n5281),.clk(gclk));
	jor g5222(.dina(n5281),.dinb(n5280),.dout(n5282),.clk(gclk));
	jand g5223(.dina(n5282),.dinb(n5266),.dout(n5283),.clk(gclk));
	jxor g5224(.dina(w_n4451_0[0]),.dinb(w_n4381_0[0]),.dout(n5284),.clk(gclk));
	jor g5225(.dina(n5284),.dinb(n5283),.dout(n5285),.clk(gclk));
	jand g5226(.dina(n5285),.dinb(n5265),.dout(n5286),.clk(gclk));
	jxor g5227(.dina(w_n4539_0[0]),.dinb(w_n4469_0[0]),.dout(n5287),.clk(gclk));
	jor g5228(.dina(n5287),.dinb(n5286),.dout(n5288),.clk(gclk));
	jand g5229(.dina(n5288),.dinb(n5264),.dout(n5289),.clk(gclk));
	jxor g5230(.dina(w_n4625_0[0]),.dinb(w_n4563_0[0]),.dout(n5290),.clk(gclk));
	jor g5231(.dina(n5290),.dinb(n5289),.dout(n5291),.clk(gclk));
	jand g5232(.dina(n5291),.dinb(n5263),.dout(n5292),.clk(gclk));
	jxor g5233(.dina(w_n4709_0[0]),.dinb(w_n4652_0[0]),.dout(n5293),.clk(gclk));
	jor g5234(.dina(n5293),.dinb(n5292),.dout(n5294),.clk(gclk));
	jand g5235(.dina(n5294),.dinb(n5262),.dout(n5295),.clk(gclk));
	jxor g5236(.dina(w_n4771_0[0]),.dinb(w_n4722_0[0]),.dout(n5296),.clk(gclk));
	jxor g5237(.dina(w_n4782_0[0]),.dinb(n5296),.dout(n5297),.clk(gclk));
	jor g5238(.dina(n5297),.dinb(n5295),.dout(n5298),.clk(gclk));
	jand g5239(.dina(n5298),.dinb(w_n4790_0[0]),.dout(n5299),.clk(gclk));
	jxor g5240(.dina(w_n4864_0[0]),.dinb(w_n4813_0[0]),.dout(n5300),.clk(gclk));
	jor g5241(.dina(n5300),.dinb(n5299),.dout(n5301),.clk(gclk));
	jand g5242(.dina(n5301),.dinb(n5261),.dout(n5302),.clk(gclk));
	jxor g5243(.dina(w_n4930_0[0]),.dinb(w_n4886_0[0]),.dout(n5303),.clk(gclk));
	jor g5244(.dina(n5303),.dinb(n5302),.dout(n5304),.clk(gclk));
	jand g5245(.dina(n5304),.dinb(n5260),.dout(n5305),.clk(gclk));
	jxor g5246(.dina(w_n5000_0[0]),.dinb(w_n4952_0[0]),.dout(n5306),.clk(gclk));
	jor g5247(.dina(n5306),.dinb(n5305),.dout(n5307),.clk(gclk));
	jand g5248(.dina(n5307),.dinb(n5259),.dout(n5308),.clk(gclk));
	jxor g5249(.dina(w_n5054_0[0]),.dinb(w_n5016_0[0]),.dout(n5309),.clk(gclk));
	jor g5250(.dina(n5309),.dinb(n5308),.dout(n5310),.clk(gclk));
	jand g5251(.dina(n5310),.dinb(n5258),.dout(n5311),.clk(gclk));
	jxor g5252(.dina(w_n5109_0[0]),.dinb(w_n5076_0[0]),.dout(n5312),.clk(gclk));
	jor g5253(.dina(n5312),.dinb(n5311),.dout(n5313),.clk(gclk));
	jand g5254(.dina(n5313),.dinb(n5257),.dout(n5314),.clk(gclk));
	jxor g5255(.dina(w_n5160_0[0]),.dinb(w_n5134_0[0]),.dout(n5315),.clk(gclk));
	jor g5256(.dina(n5315),.dinb(n5314),.dout(n5316),.clk(gclk));
	jand g5257(.dina(n5316),.dinb(n5256),.dout(n5317),.clk(gclk));
	jxor g5258(.dina(w_n5206_0[0]),.dinb(w_n5184_0[0]),.dout(n5318),.clk(gclk));
	jor g5259(.dina(n5318),.dinb(n5317),.dout(n5319),.clk(gclk));
	jand g5260(.dina(n5319),.dinb(n5255),.dout(n5320),.clk(gclk));
	jxor g5261(.dina(w_n5244_0[0]),.dinb(w_n5229_0[0]),.dout(n5321),.clk(gclk));
	jor g5262(.dina(n5321),.dinb(n5320),.dout(n5322),.clk(gclk));
	jand g5263(.dina(n5322),.dinb(n5254),.dout(n5323),.clk(gclk));
	jand g5264(.dina(w_n3895_0[0]),.dinb(w_n1035_0[2]),.dout(n5324),.clk(gclk));
	jand g5265(.dina(w_n594_0[0]),.dinb(w_n351_0[1]),.dout(n5325),.clk(gclk));
	jand g5266(.dina(n5325),.dinb(w_n2743_0[0]),.dout(n5326),.clk(gclk));
	jand g5267(.dina(n5326),.dinb(w_n229_0[0]),.dout(n5327),.clk(gclk));
	jand g5268(.dina(n5327),.dinb(w_n435_0[2]),.dout(n5328),.clk(gclk));
	jand g5269(.dina(w_n5122_0[0]),.dinb(w_n188_0[2]),.dout(n5329),.clk(gclk));
	jand g5270(.dina(n5329),.dinb(n5328),.dout(n5330),.clk(gclk));
	jand g5271(.dina(n5330),.dinb(n5324),.dout(n5331),.clk(gclk));
	jand g5272(.dina(n5331),.dinb(w_n2606_0[0]),.dout(n5332),.clk(gclk));
	jxor g5273(.dina(w_n4213_2[0]),.dinb(w_n3838_0[2]),.dout(n5333),.clk(gclk));
	jand g5274(.dina(n5333),.dinb(w_n1438_7[1]),.dout(n5334),.clk(gclk));
	jnot g5275(.din(w_n5334_0[1]),.dout(n5335),.clk(gclk));
	jand g5276(.dina(w_n5239_0[0]),.dinb(w_n5233_0[0]),.dout(n5336),.clk(gclk));
	jand g5277(.dina(w_n5243_0[0]),.dinb(w_n5240_0[0]),.dout(n5337),.clk(gclk));
	jor g5278(.dina(n5337),.dinb(n5336),.dout(n5338),.clk(gclk));
	jor g5279(.dina(w_n5238_0[0]),.dinb(w_n5236_0[1]),.dout(n5339),.clk(gclk));
	jnot g5280(.din(w_n5236_0[0]),.dout(n5340),.clk(gclk));
	jor g5281(.dina(n5340),.dinb(w_n1438_7[0]),.dout(n5341),.clk(gclk));
	jand g5282(.dina(n5341),.dinb(n5339),.dout(n5342),.clk(gclk));
	jor g5283(.dina(w_n4063_2[2]),.dinb(w_n2051_2[2]),.dout(n5343),.clk(gclk));
	jor g5284(.dina(n5343),.dinb(w_n3838_0[1]),.dout(n5344),.clk(gclk));
	jand g5285(.dina(n5344),.dinb(n5342),.dout(n5345),.clk(gclk));
	jxor g5286(.dina(n5345),.dinb(n5338),.dout(n5346),.clk(gclk));
	jxor g5287(.dina(w_n5346_0[1]),.dinb(n5335),.dout(n5347),.clk(gclk));
	jxor g5288(.dina(w_n5347_0[2]),.dinb(w_n5332_1[1]),.dout(n5348),.clk(gclk));
	jxor g5289(.dina(n5348),.dinb(w_n5323_0[1]),.dout(n5349),.clk(gclk));
	jxor g5290(.dina(w_n5349_0[1]),.dinb(w_n5252_0[1]),.dout(n5350),.clk(gclk));
	jor g5291(.dina(w_n5248_0[0]),.dinb(w_n5247_0[0]),.dout(n5351),.clk(gclk));
	jand g5292(.dina(w_n5351_0[1]),.dinb(w_n4093_6[1]),.dout(n5352),.clk(gclk));
	jxor g5293(.dina(w_dff_B_qpX2ZoCZ3_0),.dinb(w_n5350_0[1]),.dout(w_dff_A_HU6Y95fG4_2),.clk(gclk));
	jor g5294(.dina(w_n5351_0[0]),.dinb(w_n5350_0[0]),.dout(n5354),.clk(gclk));
	jand g5295(.dina(w_n5354_0[1]),.dinb(w_n4093_6[0]),.dout(n5355),.clk(gclk));
	jor g5296(.dina(w_n5349_0[0]),.dinb(w_n5252_0[0]),.dout(n5356),.clk(gclk));
	jnot g5297(.din(w_n5356_0[1]),.dout(n5357),.clk(gclk));
	jand g5298(.dina(w_n198_0[1]),.dinb(w_n166_0[2]),.dout(n5358),.clk(gclk));
	jand g5299(.dina(n5358),.dinb(w_n1050_0[0]),.dout(n5359),.clk(gclk));
	jand g5300(.dina(n5359),.dinb(w_n3481_0[0]),.dout(n5360),.clk(gclk));
	jand g5301(.dina(w_n427_0[2]),.dinb(w_n240_0[2]),.dout(n5361),.clk(gclk));
	jand g5302(.dina(n5361),.dinb(w_n388_0[1]),.dout(n5362),.clk(gclk));
	jand g5303(.dina(w_n344_1[0]),.dinb(w_n182_1[1]),.dout(n5363),.clk(gclk));
	jand g5304(.dina(n5363),.dinb(n5362),.dout(n5364),.clk(gclk));
	jand g5305(.dina(n5364),.dinb(w_n150_0[0]),.dout(n5365),.clk(gclk));
	jand g5306(.dina(n5365),.dinb(w_n884_0[1]),.dout(n5366),.clk(gclk));
	jand g5307(.dina(n5366),.dinb(w_n1147_0[0]),.dout(n5367),.clk(gclk));
	jand g5308(.dina(n5367),.dinb(n5360),.dout(n5368),.clk(gclk));
	jnot g5309(.din(w_n5368_0[2]),.dout(n5369),.clk(gclk));
	jnot g5310(.din(w_n5332_1[0]),.dout(n5370),.clk(gclk));
	jxor g5311(.dina(w_n5346_0[0]),.dinb(w_n5334_0[0]),.dout(n5371),.clk(gclk));
	jor g5312(.dina(w_n5371_0[1]),.dinb(w_n5370_0[1]),.dout(n5372),.clk(gclk));
	jand g5313(.dina(w_n5245_0[0]),.dinb(w_n5216_0[0]),.dout(n5373),.clk(gclk));
	jor g5314(.dina(n5373),.dinb(w_n5253_0[0]),.dout(n5374),.clk(gclk));
	jand g5315(.dina(w_n5371_0[0]),.dinb(w_n5370_0[0]),.dout(n5375),.clk(gclk));
	jor g5316(.dina(n5375),.dinb(n5374),.dout(n5376),.clk(gclk));
	jand g5317(.dina(n5376),.dinb(n5372),.dout(n5377),.clk(gclk));
	jxor g5318(.dina(w_n5377_0[2]),.dinb(w_n5369_0[1]),.dout(n5378),.clk(gclk));
	jxor g5319(.dina(w_n5378_0[1]),.dinb(w_n5357_0[1]),.dout(n5379),.clk(gclk));
	jxor g5320(.dina(w_n5379_0[1]),.dinb(n5355),.dout(w_dff_A_GPqiqml02_2),.clk(gclk));
	jand g5321(.dina(w_n489_1[0]),.dinb(w_n250_0[2]),.dout(n5381),.clk(gclk));
	jand g5322(.dina(n5381),.dinb(w_n3488_0[0]),.dout(n5382),.clk(gclk));
	jand g5323(.dina(n5382),.dinb(w_n1365_0[0]),.dout(n5383),.clk(gclk));
	jand g5324(.dina(n5383),.dinb(w_n849_0[0]),.dout(n5384),.clk(gclk));
	jand g5325(.dina(n5384),.dinb(w_n1140_0[0]),.dout(n5385),.clk(gclk));
	jand g5326(.dina(w_n329_0[1]),.dinb(w_n182_1[0]),.dout(n5386),.clk(gclk));
	jand g5327(.dina(n5386),.dinb(w_n3098_0[0]),.dout(n5387),.clk(gclk));
	jand g5328(.dina(w_n3868_0[0]),.dinb(w_n824_0[0]),.dout(n5388),.clk(gclk));
	jand g5329(.dina(n5388),.dinb(n5387),.dout(n5389),.clk(gclk));
	jand g5330(.dina(n5389),.dinb(n5385),.dout(n5390),.clk(gclk));
	jand g5331(.dina(w_n5347_0[1]),.dinb(w_n5332_0[2]),.dout(n5391),.clk(gclk));
	jor g5332(.dina(w_n5347_0[0]),.dinb(w_n5332_0[1]),.dout(n5392),.clk(gclk));
	jand g5333(.dina(n5392),.dinb(w_n5323_0[0]),.dout(n5393),.clk(gclk));
	jor g5334(.dina(n5393),.dinb(n5391),.dout(n5394),.clk(gclk));
	jor g5335(.dina(n5394),.dinb(w_n5368_0[1]),.dout(n5395),.clk(gclk));
	jxor g5336(.dina(w_n5377_0[1]),.dinb(w_n5368_0[0]),.dout(n5396),.clk(gclk));
	jor g5337(.dina(n5396),.dinb(w_n5356_0[0]),.dout(n5397),.clk(gclk));
	jand g5338(.dina(w_n5397_0[1]),.dinb(w_n5395_0[1]),.dout(n5398),.clk(gclk));
	jxor g5339(.dina(w_n5398_0[1]),.dinb(w_n5390_1[1]),.dout(n5399),.clk(gclk));
	jor g5340(.dina(w_n5379_0[0]),.dinb(w_n5354_0[0]),.dout(n5400),.clk(gclk));
	jand g5341(.dina(w_n5400_0[2]),.dinb(w_n4093_5[2]),.dout(n5401),.clk(gclk));
	jxor g5342(.dina(n5401),.dinb(w_n5399_0[1]),.dout(w_dff_A_1nMlhPpu8_2),.clk(gclk));
	jand g5343(.dina(w_n5378_0[0]),.dinb(w_n5357_0[0]),.dout(n5403),.clk(gclk));
	jnot g5344(.din(w_n5390_1[0]),.dout(n5404),.clk(gclk));
	jand g5345(.dina(w_n5404_0[2]),.dinb(n5403),.dout(n5405),.clk(gclk));
	jor g5346(.dina(w_n5390_0[2]),.dinb(w_n5395_0[0]),.dout(n5406),.clk(gclk));
	jand g5347(.dina(w_n5219_0[0]),.dinb(w_n189_0[0]),.dout(n5407),.clk(gclk));
	jand g5348(.dina(w_n4558_0[0]),.dinb(w_n1345_0[1]),.dout(n5408),.clk(gclk));
	jand g5349(.dina(n5408),.dinb(w_n339_1[1]),.dout(n5409),.clk(gclk));
	jand g5350(.dina(n5409),.dinb(w_n3429_0[0]),.dout(n5410),.clk(gclk));
	jand g5351(.dina(n5410),.dinb(w_n598_0[0]),.dout(n5411),.clk(gclk));
	jand g5352(.dina(w_n1178_0[0]),.dinb(w_n169_0[2]),.dout(n5412),.clk(gclk));
	jand g5353(.dina(n5412),.dinb(w_n147_0[2]),.dout(n5413),.clk(gclk));
	jand g5354(.dina(n5413),.dinb(n5411),.dout(n5414),.clk(gclk));
	jand g5355(.dina(n5414),.dinb(n5407),.dout(n5415),.clk(gclk));
	jxor g5356(.dina(w_n5415_1[1]),.dinb(w_n5406_0[1]),.dout(n5416),.clk(gclk));
	jxor g5357(.dina(w_n5416_0[1]),.dinb(w_n5405_0[1]),.dout(n5417),.clk(gclk));
	jor g5358(.dina(w_n5400_0[1]),.dinb(w_n5399_0[0]),.dout(n5418),.clk(gclk));
	jand g5359(.dina(w_n5418_0[1]),.dinb(w_n4093_5[1]),.dout(n5419),.clk(gclk));
	jxor g5360(.dina(n5419),.dinb(w_n5417_0[2]),.dout(w_dff_A_AlCqYWkD8_2),.clk(gclk));
	jor g5361(.dina(w_n5415_1[0]),.dinb(w_n5406_0[0]),.dout(n5421),.clk(gclk));
	jand g5362(.dina(w_n4556_0[0]),.dinb(w_n300_1[0]),.dout(n5422),.clk(gclk));
	jand g5363(.dina(n5422),.dinb(w_n252_1[1]),.dout(n5423),.clk(gclk));
	jand g5364(.dina(w_n1962_0[0]),.dinb(w_n513_0[0]),.dout(n5424),.clk(gclk));
	jand g5365(.dina(w_n534_0[2]),.dinb(w_n267_1[0]),.dout(n5425),.clk(gclk));
	jand g5366(.dina(n5425),.dinb(w_n461_0[0]),.dout(n5426),.clk(gclk));
	jand g5367(.dina(n5426),.dinb(w_n265_0[2]),.dout(n5427),.clk(gclk));
	jand g5368(.dina(n5427),.dinb(n5424),.dout(n5428),.clk(gclk));
	jand g5369(.dina(n5428),.dinb(n5423),.dout(n5429),.clk(gclk));
	jand g5370(.dina(w_n4811_0[0]),.dinb(w_n1250_0[0]),.dout(n5430),.clk(gclk));
	jand g5371(.dina(n5430),.dinb(n5429),.dout(n5431),.clk(gclk));
	jor g5372(.dina(w_n5431_0[2]),.dinb(w_n5421_0[1]),.dout(n5432),.clk(gclk));
	jor g5373(.dina(w_n5390_0[1]),.dinb(w_n5397_0[0]),.dout(n5433),.clk(gclk));
	jand g5374(.dina(w_n5377_0[0]),.dinb(w_n5369_0[0]),.dout(n5434),.clk(gclk));
	jand g5375(.dina(w_n5404_0[1]),.dinb(n5434),.dout(n5435),.clk(gclk));
	jxor g5376(.dina(w_n5415_0[2]),.dinb(w_n5435_0[1]),.dout(n5436),.clk(gclk));
	jor g5377(.dina(n5436),.dinb(n5433),.dout(n5437),.clk(gclk));
	jand g5378(.dina(w_n5431_0[1]),.dinb(w_n5421_0[0]),.dout(n5438),.clk(gclk));
	jxor g5379(.dina(w_n5438_0[2]),.dinb(w_n5437_0[1]),.dout(n5439),.clk(gclk));
	jand g5380(.dina(n5439),.dinb(w_n5432_0[2]),.dout(n5440),.clk(gclk));
	jor g5381(.dina(w_n5418_0[0]),.dinb(w_n5417_0[1]),.dout(n5441),.clk(gclk));
	jand g5382(.dina(w_n5441_0[1]),.dinb(w_n4093_5[0]),.dout(n5442),.clk(gclk));
	jxor g5383(.dina(n5442),.dinb(w_n5440_0[1]),.dout(w_dff_A_QgvCi3b43_2),.clk(gclk));
	jand g5384(.dina(w_n5416_0[0]),.dinb(w_n5405_0[0]),.dout(n5444),.clk(gclk));
	jnot g5385(.din(w_n5415_0[1]),.dout(n5445),.clk(gclk));
	jand g5386(.dina(n5445),.dinb(w_n5435_0[0]),.dout(n5446),.clk(gclk));
	jnot g5387(.din(w_n5431_0[0]),.dout(n5447),.clk(gclk));
	jor g5388(.dina(w_n5447_0[1]),.dinb(w_n5446_0[1]),.dout(n5448),.clk(gclk));
	jand g5389(.dina(n5448),.dinb(w_n5444_0[1]),.dout(n5449),.clk(gclk));
	jand g5390(.dina(w_n452_0[0]),.dinb(w_n373_0[0]),.dout(n5450),.clk(gclk));
	jand g5391(.dina(n5450),.dinb(w_n3826_0[0]),.dout(n5451),.clk(gclk));
	jand g5392(.dina(n5451),.dinb(w_n1474_2[1]),.dout(n5452),.clk(gclk));
	jxor g5393(.dina(w_n5452_1[1]),.dinb(w_n5432_0[1]),.dout(n5453),.clk(gclk));
	jxor g5394(.dina(w_n5453_0[1]),.dinb(w_n5449_0[1]),.dout(n5454),.clk(gclk));
	jor g5395(.dina(w_n5441_0[0]),.dinb(w_n5440_0[0]),.dout(n5455),.clk(gclk));
	jand g5396(.dina(w_n5455_0[1]),.dinb(w_n4093_4[2]),.dout(n5456),.clk(gclk));
	jxor g5397(.dina(n5456),.dinb(w_n5454_0[2]),.dout(w_dff_A_khtMLhmf2_2),.clk(gclk));
	jand g5398(.dina(w_n5453_0[0]),.dinb(w_n5449_0[0]),.dout(n5458),.clk(gclk));
	jand g5399(.dina(w_n5447_0[0]),.dinb(w_n5446_0[0]),.dout(n5459),.clk(gclk));
	jnot g5400(.din(w_n5452_1[0]),.dout(n5460),.clk(gclk));
	jand g5401(.dina(n5460),.dinb(w_n5459_0[2]),.dout(n5461),.clk(gclk));
	jor g5402(.dina(w_n1494_2[0]),.dinb(w_n504_0[0]),.dout(n5462),.clk(gclk));
	jor g5403(.dina(w_n5462_0[2]),.dinb(w_n5461_0[1]),.dout(n5463),.clk(gclk));
	jor g5404(.dina(w_n5463_0[1]),.dinb(w_n5458_0[1]),.dout(n5464),.clk(gclk));
	jor g5405(.dina(w_n5452_0[2]),.dinb(w_n5432_0[0]),.dout(n5465),.clk(gclk));
	jnot g5406(.din(w_n5462_0[1]),.dout(n5466),.clk(gclk));
	jand g5407(.dina(w_n5466_0[1]),.dinb(w_n5465_0[1]),.dout(n5467),.clk(gclk));
	jor g5408(.dina(w_n5438_0[1]),.dinb(w_n5437_0[0]),.dout(n5468),.clk(gclk));
	jxor g5409(.dina(w_n5452_0[1]),.dinb(w_n5459_0[1]),.dout(n5469),.clk(gclk));
	jor g5410(.dina(n5469),.dinb(n5468),.dout(n5470),.clk(gclk));
	jor g5411(.dina(w_n5466_0[0]),.dinb(w_n5465_0[0]),.dout(n5471),.clk(gclk));
	jand g5412(.dina(w_n5471_0[1]),.dinb(w_n5470_0[1]),.dout(n5472),.clk(gclk));
	jor g5413(.dina(n5472),.dinb(n5467),.dout(n5473),.clk(gclk));
	jand g5414(.dina(n5473),.dinb(n5464),.dout(n5474),.clk(gclk));
	jor g5415(.dina(w_n5455_0[0]),.dinb(w_n5454_0[1]),.dout(n5475),.clk(gclk));
	jand g5416(.dina(n5475),.dinb(w_n4093_4[1]),.dout(n5476),.clk(gclk));
	jxor g5417(.dina(w_n5476_0[1]),.dinb(w_n5474_0[1]),.dout(w_dff_A_d1DL4wzM4_2),.clk(gclk));
	jnot g5418(.din(w_n72_0[0]),.dout(n5478),.clk(gclk));
	jand g5419(.dina(n5478),.dinb(w_n49_3[0]),.dout(n5479),.clk(gclk));
	jand g5420(.dina(n5479),.dinb(w_n71_0[0]),.dout(n5480),.clk(gclk));
	jand g5421(.dina(w_n5462_0[0]),.dinb(w_n5461_0[0]),.dout(n5481),.clk(gclk));
	jor g5422(.dina(n5481),.dinb(w_n5458_0[0]),.dout(n5482),.clk(gclk));
	jand g5423(.dina(n5482),.dinb(w_n5463_0[0]),.dout(n5483),.clk(gclk));
	jor g5424(.dina(w_n5471_0[0]),.dinb(w_n5470_0[0]),.dout(n5484),.clk(gclk));
	jand g5425(.dina(w_n5484_0[1]),.dinb(w_n5483_0[1]),.dout(n5485),.clk(gclk));
	jand g5426(.dina(w_n5474_0[0]),.dinb(w_n4093_4[0]),.dout(n5486),.clk(gclk));
	jor g5427(.dina(n5486),.dinb(w_n5476_0[0]),.dout(n5487),.clk(gclk));
	jxor g5428(.dina(w_n5487_0[1]),.dinb(w_dff_B_qjcjo5yK6_1),.dout(n5488),.clk(gclk));
	jor g5429(.dina(n5488),.dinb(w_n5480_0[1]),.dout(sin23),.clk(gclk));
	jand g5430(.dina(w_n5487_0[0]),.dinb(w_n5484_0[0]),.dout(n5490),.clk(gclk));
	jnot g5431(.din(w_n5454_0[0]),.dout(n5491),.clk(gclk));
	jxor g5432(.dina(w_n5438_0[0]),.dinb(w_n5444_0[0]),.dout(n5492),.clk(gclk));
	jor g5433(.dina(n5492),.dinb(w_n5459_0[0]),.dout(n5493),.clk(gclk));
	jnot g5434(.din(w_n5417_0[0]),.dout(n5494),.clk(gclk));
	jxor g5435(.dina(w_n5398_0[0]),.dinb(w_n5404_0[0]),.dout(n5495),.clk(gclk));
	jnot g5436(.din(w_n5400_0[0]),.dout(n5496),.clk(gclk));
	jand g5437(.dina(n5496),.dinb(n5495),.dout(n5497),.clk(gclk));
	jand g5438(.dina(n5497),.dinb(n5494),.dout(n5498),.clk(gclk));
	jand g5439(.dina(n5498),.dinb(n5493),.dout(n5499),.clk(gclk));
	jand g5440(.dina(n5499),.dinb(n5491),.dout(n5500),.clk(gclk));
	jand g5441(.dina(n5500),.dinb(w_n5483_0[0]),.dout(n5501),.clk(gclk));
	jor g5442(.dina(n5501),.dinb(w_n5480_0[0]),.dout(n5502),.clk(gclk));
	jand g5443(.dina(n5502),.dinb(w_n4093_3[2]),.dout(n5503),.clk(gclk));
	jor g5444(.dina(w_dff_B_pNwtQMbW3_0),.dinb(n5490),.dout(sin24),.clk(gclk));
	jspl3 jspl3_w_a0_0(.douta(w_a0_0[0]),.doutb(w_a0_0[1]),.doutc(w_a0_0[2]),.din(a0));
	jspl3 jspl3_w_a1_0(.douta(w_a1_0[0]),.doutb(w_a1_0[1]),.doutc(w_a1_0[2]),.din(a1));
	jspl jspl_w_a2_0(.douta(w_a2_0[0]),.doutb(w_a2_0[1]),.din(a2));
	jspl jspl_w_a3_0(.douta(w_a3_0[0]),.doutb(w_a3_0[1]),.din(a3));
	jspl jspl_w_a4_0(.douta(w_a4_0[0]),.doutb(w_a4_0[1]),.din(a4));
	jspl jspl_w_a5_0(.douta(w_a5_0[0]),.doutb(w_a5_0[1]),.din(a5));
	jspl jspl_w_a6_0(.douta(w_a6_0[0]),.doutb(w_a6_0[1]),.din(a6));
	jspl jspl_w_a7_0(.douta(w_a7_0[0]),.doutb(w_a7_0[1]),.din(a7));
	jspl jspl_w_a8_0(.douta(w_a8_0[0]),.doutb(w_a8_0[1]),.din(a8));
	jspl jspl_w_a9_0(.douta(w_a9_0[0]),.doutb(w_a9_0[1]),.din(a9));
	jspl jspl_w_a10_0(.douta(w_a10_0[0]),.doutb(w_a10_0[1]),.din(a10));
	jspl jspl_w_a11_0(.douta(w_a11_0[0]),.doutb(w_a11_0[1]),.din(a11));
	jspl jspl_w_a12_0(.douta(w_a12_0[0]),.doutb(w_a12_0[1]),.din(a12));
	jspl jspl_w_a13_0(.douta(w_a13_0[0]),.doutb(w_a13_0[1]),.din(a13));
	jspl jspl_w_a14_0(.douta(w_a14_0[0]),.doutb(w_a14_0[1]),.din(a14));
	jspl jspl_w_a15_0(.douta(w_a15_0[0]),.doutb(w_a15_0[1]),.din(a15));
	jspl jspl_w_a16_0(.douta(w_a16_0[0]),.doutb(w_a16_0[1]),.din(a16));
	jspl jspl_w_a17_0(.douta(w_a17_0[0]),.doutb(w_a17_0[1]),.din(a17));
	jspl jspl_w_a18_0(.douta(w_a18_0[0]),.doutb(w_a18_0[1]),.din(a18));
	jspl3 jspl3_w_a19_0(.douta(w_a19_0[0]),.doutb(w_a19_0[1]),.doutc(w_a19_0[2]),.din(a19));
	jspl3 jspl3_w_a20_0(.douta(w_a20_0[0]),.doutb(w_a20_0[1]),.doutc(w_a20_0[2]),.din(a20));
	jspl jspl_w_a21_0(.douta(w_a21_0[0]),.doutb(w_a21_0[1]),.din(a21));
	jspl3 jspl3_w_a22_0(.douta(w_a22_0[0]),.doutb(w_a22_0[1]),.doutc(w_a22_0[2]),.din(a22));
	jspl3 jspl3_w_sin0_0(.douta(w_dff_A_gvfmGipg2_0),.doutb(w_sin0_0[1]),.doutc(w_dff_A_RcIzSiyI2_2),.din(sin0_fa_));
	jspl3 jspl3_w_n49_0(.douta(w_n49_0[0]),.doutb(w_n49_0[1]),.doutc(w_n49_0[2]),.din(n49));
	jspl3 jspl3_w_n49_1(.douta(w_n49_1[0]),.doutb(w_n49_1[1]),.doutc(w_n49_1[2]),.din(w_n49_0[0]));
	jspl3 jspl3_w_n49_2(.douta(w_n49_2[0]),.doutb(w_n49_2[1]),.doutc(w_n49_2[2]),.din(w_n49_0[1]));
	jspl3 jspl3_w_n49_3(.douta(w_n49_3[0]),.doutb(w_n49_3[1]),.doutc(w_n49_3[2]),.din(w_n49_0[2]));
	jspl3 jspl3_w_n49_4(.douta(w_n49_4[0]),.doutb(w_n49_4[1]),.doutc(w_n49_4[2]),.din(w_n49_1[0]));
	jspl3 jspl3_w_n49_5(.douta(w_n49_5[0]),.doutb(w_n49_5[1]),.doutc(w_n49_5[2]),.din(w_n49_1[1]));
	jspl3 jspl3_w_n49_6(.douta(w_n49_6[0]),.doutb(w_n49_6[1]),.doutc(w_n49_6[2]),.din(w_n49_1[2]));
	jspl3 jspl3_w_n49_7(.douta(w_n49_7[0]),.doutb(w_n49_7[1]),.doutc(w_n49_7[2]),.din(w_n49_2[0]));
	jspl3 jspl3_w_n49_8(.douta(w_n49_8[0]),.doutb(w_n49_8[1]),.doutc(w_n49_8[2]),.din(w_n49_2[1]));
	jspl3 jspl3_w_n49_9(.douta(w_n49_9[0]),.doutb(w_n49_9[1]),.doutc(w_n49_9[2]),.din(w_n49_2[2]));
	jspl3 jspl3_w_n50_0(.douta(w_n50_0[0]),.doutb(w_n50_0[1]),.doutc(w_n50_0[2]),.din(n50));
	jspl jspl_w_n51_0(.douta(w_n51_0[0]),.doutb(w_n51_0[1]),.din(n51));
	jspl jspl_w_n52_0(.douta(w_n52_0[0]),.doutb(w_n52_0[1]),.din(n52));
	jspl jspl_w_n53_0(.douta(w_n53_0[0]),.doutb(w_n53_0[1]),.din(n53));
	jspl jspl_w_n54_0(.douta(w_n54_0[0]),.doutb(w_n54_0[1]),.din(n54));
	jspl jspl_w_n55_0(.douta(w_n55_0[0]),.doutb(w_n55_0[1]),.din(n55));
	jspl jspl_w_n56_0(.douta(w_n56_0[0]),.doutb(w_n56_0[1]),.din(n56));
	jspl jspl_w_n57_0(.douta(w_n57_0[0]),.doutb(w_n57_0[1]),.din(n57));
	jspl jspl_w_n58_0(.douta(w_n58_0[0]),.doutb(w_n58_0[1]),.din(n58));
	jspl jspl_w_n59_0(.douta(w_n59_0[0]),.doutb(w_n59_0[1]),.din(n59));
	jspl jspl_w_n60_0(.douta(w_n60_0[0]),.doutb(w_n60_0[1]),.din(n60));
	jspl jspl_w_n61_0(.douta(w_n61_0[0]),.doutb(w_n61_0[1]),.din(n61));
	jspl jspl_w_n62_0(.douta(w_n62_0[0]),.doutb(w_n62_0[1]),.din(n62));
	jspl jspl_w_n63_0(.douta(w_n63_0[0]),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n64_0(.douta(w_n64_0[0]),.doutb(w_n64_0[1]),.din(n64));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n66_0(.douta(w_n66_0[0]),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(n67));
	jspl jspl_w_n68_0(.douta(w_n68_0[0]),.doutb(w_n68_0[1]),.din(n68));
	jspl jspl_w_n69_0(.douta(w_n69_0[0]),.doutb(w_n69_0[1]),.din(n69));
	jspl3 jspl3_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.doutc(w_n70_0[2]),.din(n70));
	jspl jspl_w_n70_1(.douta(w_n70_1[0]),.doutb(w_n70_1[1]),.din(w_n70_0[0]));
	jspl jspl_w_n71_0(.douta(w_n71_0[0]),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n72_0(.douta(w_n72_0[0]),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.din(n73));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.doutc(w_n75_0[2]),.din(n75));
	jspl3 jspl3_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.doutc(w_n75_1[2]),.din(w_n75_0[0]));
	jspl jspl_w_n75_2(.douta(w_n75_2[0]),.doutb(w_n75_2[1]),.din(w_n75_0[1]));
	jspl3 jspl3_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.doutc(w_n77_0[2]),.din(n77));
	jspl3 jspl3_w_n77_1(.douta(w_n77_1[0]),.doutb(w_n77_1[1]),.doutc(w_n77_1[2]),.din(w_n77_0[0]));
	jspl3 jspl3_w_n77_2(.douta(w_n77_2[0]),.doutb(w_n77_2[1]),.doutc(w_n77_2[2]),.din(w_n77_0[1]));
	jspl3 jspl3_w_n77_3(.douta(w_n77_3[0]),.doutb(w_n77_3[1]),.doutc(w_n77_3[2]),.din(w_n77_0[2]));
	jspl3 jspl3_w_n77_4(.douta(w_n77_4[0]),.doutb(w_n77_4[1]),.doutc(w_n77_4[2]),.din(w_n77_1[0]));
	jspl3 jspl3_w_n77_5(.douta(w_n77_5[0]),.doutb(w_n77_5[1]),.doutc(w_n77_5[2]),.din(w_n77_1[1]));
	jspl3 jspl3_w_n77_6(.douta(w_n77_6[0]),.doutb(w_n77_6[1]),.doutc(w_n77_6[2]),.din(w_n77_1[2]));
	jspl3 jspl3_w_n77_7(.douta(w_n77_7[0]),.doutb(w_n77_7[1]),.doutc(w_n77_7[2]),.din(w_n77_2[0]));
	jspl3 jspl3_w_n77_8(.douta(w_n77_8[0]),.doutb(w_n77_8[1]),.doutc(w_n77_8[2]),.din(w_n77_2[1]));
	jspl3 jspl3_w_n77_9(.douta(w_n77_9[0]),.doutb(w_n77_9[1]),.doutc(w_n77_9[2]),.din(w_n77_2[2]));
	jspl3 jspl3_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.doutc(w_n78_0[2]),.din(n78));
	jspl3 jspl3_w_n78_1(.douta(w_n78_1[0]),.doutb(w_n78_1[1]),.doutc(w_n78_1[2]),.din(w_n78_0[0]));
	jspl3 jspl3_w_n78_2(.douta(w_n78_2[0]),.doutb(w_n78_2[1]),.doutc(w_n78_2[2]),.din(w_n78_0[1]));
	jspl3 jspl3_w_n78_3(.douta(w_n78_3[0]),.doutb(w_n78_3[1]),.doutc(w_n78_3[2]),.din(w_n78_0[2]));
	jspl jspl_w_n80_0(.douta(w_n80_0[0]),.doutb(w_n80_0[1]),.din(n80));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl3 jspl3_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.doutc(w_n83_0[2]),.din(n83));
	jspl3 jspl3_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.doutc(w_n84_0[2]),.din(n84));
	jspl3 jspl3_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.doutc(w_n85_0[2]),.din(n85));
	jspl jspl_w_n85_1(.douta(w_n85_1[0]),.doutb(w_n85_1[1]),.din(w_n85_0[0]));
	jspl3 jspl3_w_n87_0(.douta(w_n87_0[0]),.doutb(w_n87_0[1]),.doutc(w_n87_0[2]),.din(n87));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.doutc(w_n90_0[2]),.din(n90));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.doutc(w_n91_0[2]),.din(n91));
	jspl jspl_w_n91_1(.douta(w_n91_1[0]),.doutb(w_n91_1[1]),.din(w_n91_0[0]));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl3 jspl3_w_n92_1(.douta(w_n92_1[0]),.doutb(w_n92_1[1]),.doutc(w_n92_1[2]),.din(w_n92_0[0]));
	jspl3 jspl3_w_n92_2(.douta(w_n92_2[0]),.doutb(w_n92_2[1]),.doutc(w_n92_2[2]),.din(w_n92_0[1]));
	jspl3 jspl3_w_n92_3(.douta(w_n92_3[0]),.doutb(w_n92_3[1]),.doutc(w_n92_3[2]),.din(w_n92_0[2]));
	jspl3 jspl3_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.doutc(w_n93_0[2]),.din(n93));
	jspl3 jspl3_w_n93_1(.douta(w_n93_1[0]),.doutb(w_n93_1[1]),.doutc(w_n93_1[2]),.din(w_n93_0[0]));
	jspl3 jspl3_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl3 jspl3_w_n94_1(.douta(w_n94_1[0]),.doutb(w_n94_1[1]),.doutc(w_n94_1[2]),.din(w_n94_0[0]));
	jspl3 jspl3_w_n94_2(.douta(w_n94_2[0]),.doutb(w_n94_2[1]),.doutc(w_n94_2[2]),.din(w_n94_0[1]));
	jspl jspl_w_n95_0(.douta(w_n95_0[0]),.doutb(w_n95_0[1]),.din(n95));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.doutc(w_n96_0[2]),.din(n96));
	jspl jspl_w_n96_1(.douta(w_n96_1[0]),.doutb(w_n96_1[1]),.din(w_n96_0[0]));
	jspl3 jspl3_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.doutc(w_n97_0[2]),.din(n97));
	jspl jspl_w_n97_1(.douta(w_n97_1[0]),.doutb(w_n97_1[1]),.din(w_n97_0[0]));
	jspl3 jspl3_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.doutc(w_n98_0[2]),.din(n98));
	jspl3 jspl3_w_n98_1(.douta(w_n98_1[0]),.doutb(w_n98_1[1]),.doutc(w_n98_1[2]),.din(w_n98_0[0]));
	jspl3 jspl3_w_n98_2(.douta(w_n98_2[0]),.doutb(w_n98_2[1]),.doutc(w_n98_2[2]),.din(w_n98_0[1]));
	jspl3 jspl3_w_n98_3(.douta(w_n98_3[0]),.doutb(w_n98_3[1]),.doutc(w_n98_3[2]),.din(w_n98_0[2]));
	jspl3 jspl3_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.doutc(w_n99_0[2]),.din(n99));
	jspl3 jspl3_w_n99_1(.douta(w_n99_1[0]),.doutb(w_n99_1[1]),.doutc(w_n99_1[2]),.din(w_n99_0[0]));
	jspl3 jspl3_w_n99_2(.douta(w_n99_2[0]),.doutb(w_n99_2[1]),.doutc(w_n99_2[2]),.din(w_n99_0[1]));
	jspl jspl_w_n99_3(.douta(w_n99_3[0]),.doutb(w_n99_3[1]),.din(w_n99_0[2]));
	jspl3 jspl3_w_n100_0(.douta(w_n100_0[0]),.doutb(w_n100_0[1]),.doutc(w_n100_0[2]),.din(n100));
	jspl3 jspl3_w_n100_1(.douta(w_n100_1[0]),.doutb(w_n100_1[1]),.doutc(w_n100_1[2]),.din(w_n100_0[0]));
	jspl3 jspl3_w_n100_2(.douta(w_n100_2[0]),.doutb(w_n100_2[1]),.doutc(w_n100_2[2]),.din(w_n100_0[1]));
	jspl3 jspl3_w_n100_3(.douta(w_n100_3[0]),.doutb(w_n100_3[1]),.doutc(w_n100_3[2]),.din(w_n100_0[2]));
	jspl3 jspl3_w_n100_4(.douta(w_n100_4[0]),.doutb(w_n100_4[1]),.doutc(w_n100_4[2]),.din(w_n100_1[0]));
	jspl3 jspl3_w_n100_5(.douta(w_n100_5[0]),.doutb(w_n100_5[1]),.doutc(w_n100_5[2]),.din(w_n100_1[1]));
	jspl3 jspl3_w_n100_6(.douta(w_n100_6[0]),.doutb(w_n100_6[1]),.doutc(w_n100_6[2]),.din(w_n100_1[2]));
	jspl3 jspl3_w_n100_7(.douta(w_n100_7[0]),.doutb(w_n100_7[1]),.doutc(w_n100_7[2]),.din(w_n100_2[0]));
	jspl3 jspl3_w_n100_8(.douta(w_n100_8[0]),.doutb(w_n100_8[1]),.doutc(w_n100_8[2]),.din(w_n100_2[1]));
	jspl3 jspl3_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl3 jspl3_w_n101_1(.douta(w_n101_1[0]),.doutb(w_n101_1[1]),.doutc(w_n101_1[2]),.din(w_n101_0[0]));
	jspl3 jspl3_w_n101_2(.douta(w_n101_2[0]),.doutb(w_n101_2[1]),.doutc(w_n101_2[2]),.din(w_n101_0[1]));
	jspl3 jspl3_w_n101_3(.douta(w_n101_3[0]),.doutb(w_n101_3[1]),.doutc(w_n101_3[2]),.din(w_n101_0[2]));
	jspl3 jspl3_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.doutc(w_n102_0[2]),.din(n102));
	jspl3 jspl3_w_n102_1(.douta(w_n102_1[0]),.doutb(w_n102_1[1]),.doutc(w_n102_1[2]),.din(w_n102_0[0]));
	jspl3 jspl3_w_n102_2(.douta(w_n102_2[0]),.doutb(w_n102_2[1]),.doutc(w_n102_2[2]),.din(w_n102_0[1]));
	jspl jspl_w_n102_3(.douta(w_n102_3[0]),.doutb(w_n102_3[1]),.din(w_n102_0[2]));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.doutc(w_n103_0[2]),.din(n103));
	jspl jspl_w_n103_1(.douta(w_n103_1[0]),.doutb(w_n103_1[1]),.din(w_n103_0[0]));
	jspl3 jspl3_w_n105_0(.douta(w_n105_0[0]),.doutb(w_n105_0[1]),.doutc(w_n105_0[2]),.din(n105));
	jspl jspl_w_n105_1(.douta(w_n105_1[0]),.doutb(w_n105_1[1]),.din(w_n105_0[0]));
	jspl3 jspl3_w_n106_0(.douta(w_n106_0[0]),.doutb(w_n106_0[1]),.doutc(w_n106_0[2]),.din(n106));
	jspl jspl_w_n106_1(.douta(w_n106_1[0]),.doutb(w_n106_1[1]),.din(w_n106_0[0]));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl3 jspl3_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.doutc(w_n108_0[2]),.din(n108));
	jspl3 jspl3_w_n108_1(.douta(w_n108_1[0]),.doutb(w_n108_1[1]),.doutc(w_n108_1[2]),.din(w_n108_0[0]));
	jspl3 jspl3_w_n108_2(.douta(w_n108_2[0]),.doutb(w_n108_2[1]),.doutc(w_n108_2[2]),.din(w_n108_0[1]));
	jspl3 jspl3_w_n108_3(.douta(w_n108_3[0]),.doutb(w_n108_3[1]),.doutc(w_n108_3[2]),.din(w_n108_0[2]));
	jspl3 jspl3_w_n108_4(.douta(w_n108_4[0]),.doutb(w_n108_4[1]),.doutc(w_n108_4[2]),.din(w_n108_1[0]));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n110_0(.douta(w_n110_0[0]),.doutb(w_n110_0[1]),.doutc(w_n110_0[2]),.din(n110));
	jspl3 jspl3_w_n110_1(.douta(w_n110_1[0]),.doutb(w_n110_1[1]),.doutc(w_n110_1[2]),.din(w_n110_0[0]));
	jspl3 jspl3_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.doutc(w_n111_0[2]),.din(n111));
	jspl jspl_w_n111_1(.douta(w_n111_1[0]),.doutb(w_n111_1[1]),.din(w_n111_0[0]));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl3 jspl3_w_n112_3(.douta(w_n112_3[0]),.doutb(w_n112_3[1]),.doutc(w_n112_3[2]),.din(w_n112_0[2]));
	jspl jspl_w_n112_4(.douta(w_n112_4[0]),.doutb(w_n112_4[1]),.din(w_n112_1[0]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.doutc(w_n113_0[2]),.din(n113));
	jspl3 jspl3_w_n113_1(.douta(w_n113_1[0]),.doutb(w_n113_1[1]),.doutc(w_n113_1[2]),.din(w_n113_0[0]));
	jspl3 jspl3_w_n113_2(.douta(w_n113_2[0]),.doutb(w_n113_2[1]),.doutc(w_n113_2[2]),.din(w_n113_0[1]));
	jspl3 jspl3_w_n114_0(.douta(w_n114_0[0]),.doutb(w_n114_0[1]),.doutc(w_n114_0[2]),.din(n114));
	jspl3 jspl3_w_n114_1(.douta(w_n114_1[0]),.doutb(w_n114_1[1]),.doutc(w_n114_1[2]),.din(w_n114_0[0]));
	jspl3 jspl3_w_n114_2(.douta(w_n114_2[0]),.doutb(w_n114_2[1]),.doutc(w_n114_2[2]),.din(w_n114_0[1]));
	jspl3 jspl3_w_n114_3(.douta(w_n114_3[0]),.doutb(w_n114_3[1]),.doutc(w_n114_3[2]),.din(w_n114_0[2]));
	jspl3 jspl3_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.doutc(w_n115_0[2]),.din(n115));
	jspl jspl_w_n115_1(.douta(w_n115_1[0]),.doutb(w_n115_1[1]),.din(w_n115_0[0]));
	jspl3 jspl3_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.doutc(w_n116_0[2]),.din(n116));
	jspl3 jspl3_w_n116_1(.douta(w_n116_1[0]),.doutb(w_n116_1[1]),.doutc(w_n116_1[2]),.din(w_n116_0[0]));
	jspl3 jspl3_w_n116_2(.douta(w_n116_2[0]),.doutb(w_n116_2[1]),.doutc(w_n116_2[2]),.din(w_n116_0[1]));
	jspl jspl_w_n116_3(.douta(w_n116_3[0]),.doutb(w_n116_3[1]),.din(w_n116_0[2]));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n117_1(.douta(w_n117_1[0]),.doutb(w_n117_1[1]),.din(w_n117_0[0]));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl3 jspl3_w_n118_1(.douta(w_n118_1[0]),.doutb(w_n118_1[1]),.doutc(w_n118_1[2]),.din(w_n118_0[0]));
	jspl3 jspl3_w_n118_2(.douta(w_n118_2[0]),.doutb(w_n118_2[1]),.doutc(w_n118_2[2]),.din(w_n118_0[1]));
	jspl3 jspl3_w_n118_3(.douta(w_n118_3[0]),.doutb(w_n118_3[1]),.doutc(w_n118_3[2]),.din(w_n118_0[2]));
	jspl3 jspl3_w_n118_4(.douta(w_n118_4[0]),.doutb(w_n118_4[1]),.doutc(w_n118_4[2]),.din(w_n118_1[0]));
	jspl3 jspl3_w_n118_5(.douta(w_n118_5[0]),.doutb(w_n118_5[1]),.doutc(w_n118_5[2]),.din(w_n118_1[1]));
	jspl3 jspl3_w_n118_6(.douta(w_n118_6[0]),.doutb(w_n118_6[1]),.doutc(w_n118_6[2]),.din(w_n118_1[2]));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl3 jspl3_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.doutc(w_n120_0[2]),.din(n120));
	jspl3 jspl3_w_n120_1(.douta(w_n120_1[0]),.doutb(w_n120_1[1]),.doutc(w_n120_1[2]),.din(w_n120_0[0]));
	jspl3 jspl3_w_n120_2(.douta(w_n120_2[0]),.doutb(w_n120_2[1]),.doutc(w_n120_2[2]),.din(w_n120_0[1]));
	jspl3 jspl3_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.doutc(w_n123_0[2]),.din(n123));
	jspl3 jspl3_w_n123_1(.douta(w_n123_1[0]),.doutb(w_n123_1[1]),.doutc(w_n123_1[2]),.din(w_n123_0[0]));
	jspl jspl_w_n123_2(.douta(w_n123_2[0]),.doutb(w_n123_2[1]),.din(w_n123_0[1]));
	jspl3 jspl3_w_n124_0(.douta(w_n124_0[0]),.doutb(w_n124_0[1]),.doutc(w_n124_0[2]),.din(n124));
	jspl3 jspl3_w_n124_1(.douta(w_n124_1[0]),.doutb(w_n124_1[1]),.doutc(w_n124_1[2]),.din(w_n124_0[0]));
	jspl3 jspl3_w_n124_2(.douta(w_n124_2[0]),.doutb(w_n124_2[1]),.doutc(w_n124_2[2]),.din(w_n124_0[1]));
	jspl3 jspl3_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.doutc(w_n125_0[2]),.din(n125));
	jspl3 jspl3_w_n125_1(.douta(w_n125_1[0]),.doutb(w_n125_1[1]),.doutc(w_n125_1[2]),.din(w_n125_0[0]));
	jspl3 jspl3_w_n125_2(.douta(w_n125_2[0]),.doutb(w_n125_2[1]),.doutc(w_n125_2[2]),.din(w_n125_0[1]));
	jspl3 jspl3_w_n125_3(.douta(w_n125_3[0]),.doutb(w_n125_3[1]),.doutc(w_n125_3[2]),.din(w_n125_0[2]));
	jspl3 jspl3_w_n125_4(.douta(w_n125_4[0]),.doutb(w_n125_4[1]),.doutc(w_n125_4[2]),.din(w_n125_1[0]));
	jspl jspl_w_n125_5(.douta(w_n125_5[0]),.doutb(w_n125_5[1]),.din(w_n125_1[1]));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl3 jspl3_w_n126_1(.douta(w_n126_1[0]),.doutb(w_n126_1[1]),.doutc(w_n126_1[2]),.din(w_n126_0[0]));
	jspl3 jspl3_w_n126_2(.douta(w_n126_2[0]),.doutb(w_n126_2[1]),.doutc(w_n126_2[2]),.din(w_n126_0[1]));
	jspl3 jspl3_w_n126_3(.douta(w_n126_3[0]),.doutb(w_n126_3[1]),.doutc(w_n126_3[2]),.din(w_n126_0[2]));
	jspl jspl_w_n126_4(.douta(w_n126_4[0]),.doutb(w_n126_4[1]),.din(w_n126_1[0]));
	jspl3 jspl3_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.doutc(w_n127_0[2]),.din(n127));
	jspl3 jspl3_w_n127_1(.douta(w_n127_1[0]),.doutb(w_n127_1[1]),.doutc(w_n127_1[2]),.din(w_n127_0[0]));
	jspl3 jspl3_w_n127_2(.douta(w_n127_2[0]),.doutb(w_n127_2[1]),.doutc(w_n127_2[2]),.din(w_n127_0[1]));
	jspl jspl_w_n127_3(.douta(w_n127_3[0]),.doutb(w_n127_3[1]),.din(w_n127_0[2]));
	jspl3 jspl3_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.doutc(w_n128_0[2]),.din(n128));
	jspl3 jspl3_w_n128_1(.douta(w_n128_1[0]),.doutb(w_n128_1[1]),.doutc(w_n128_1[2]),.din(w_n128_0[0]));
	jspl3 jspl3_w_n128_2(.douta(w_n128_2[0]),.doutb(w_n128_2[1]),.doutc(w_n128_2[2]),.din(w_n128_0[1]));
	jspl jspl_w_n128_3(.douta(w_n128_3[0]),.doutb(w_n128_3[1]),.din(w_n128_0[2]));
	jspl3 jspl3_w_n129_0(.douta(w_n129_0[0]),.doutb(w_n129_0[1]),.doutc(w_n129_0[2]),.din(n129));
	jspl3 jspl3_w_n129_1(.douta(w_n129_1[0]),.doutb(w_n129_1[1]),.doutc(w_n129_1[2]),.din(w_n129_0[0]));
	jspl3 jspl3_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.doutc(w_n130_0[2]),.din(n130));
	jspl3 jspl3_w_n130_1(.douta(w_n130_1[0]),.doutb(w_n130_1[1]),.doutc(w_n130_1[2]),.din(w_n130_0[0]));
	jspl3 jspl3_w_n130_2(.douta(w_n130_2[0]),.doutb(w_n130_2[1]),.doutc(w_n130_2[2]),.din(w_n130_0[1]));
	jspl jspl_w_n130_3(.douta(w_n130_3[0]),.doutb(w_n130_3[1]),.din(w_n130_0[2]));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_n132_0[1]),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.doutc(w_n133_0[2]),.din(n133));
	jspl3 jspl3_w_n133_1(.douta(w_n133_1[0]),.doutb(w_n133_1[1]),.doutc(w_n133_1[2]),.din(w_n133_0[0]));
	jspl jspl_w_n133_2(.douta(w_n133_2[0]),.doutb(w_n133_2[1]),.din(w_n133_0[1]));
	jspl3 jspl3_w_n134_0(.douta(w_n134_0[0]),.doutb(w_n134_0[1]),.doutc(w_n134_0[2]),.din(n134));
	jspl jspl_w_n134_1(.douta(w_n134_1[0]),.doutb(w_n134_1[1]),.din(w_n134_0[0]));
	jspl3 jspl3_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.doutc(w_n135_0[2]),.din(n135));
	jspl3 jspl3_w_n135_1(.douta(w_n135_1[0]),.doutb(w_n135_1[1]),.doutc(w_n135_1[2]),.din(w_n135_0[0]));
	jspl3 jspl3_w_n135_2(.douta(w_n135_2[0]),.doutb(w_n135_2[1]),.doutc(w_n135_2[2]),.din(w_n135_0[1]));
	jspl3 jspl3_w_n135_3(.douta(w_n135_3[0]),.doutb(w_n135_3[1]),.doutc(w_n135_3[2]),.din(w_n135_0[2]));
	jspl3 jspl3_w_n135_4(.douta(w_n135_4[0]),.doutb(w_n135_4[1]),.doutc(w_n135_4[2]),.din(w_n135_1[0]));
	jspl3 jspl3_w_n136_0(.douta(w_n136_0[0]),.doutb(w_n136_0[1]),.doutc(w_n136_0[2]),.din(n136));
	jspl3 jspl3_w_n136_1(.douta(w_n136_1[0]),.doutb(w_n136_1[1]),.doutc(w_n136_1[2]),.din(w_n136_0[0]));
	jspl jspl_w_n136_2(.douta(w_n136_2[0]),.doutb(w_n136_2[1]),.din(w_n136_0[1]));
	jspl3 jspl3_w_n137_0(.douta(w_n137_0[0]),.doutb(w_n137_0[1]),.doutc(w_n137_0[2]),.din(n137));
	jspl3 jspl3_w_n137_1(.douta(w_n137_1[0]),.doutb(w_n137_1[1]),.doutc(w_n137_1[2]),.din(w_n137_0[0]));
	jspl jspl_w_n137_2(.douta(w_n137_2[0]),.doutb(w_n137_2[1]),.din(w_n137_0[1]));
	jspl3 jspl3_w_n138_0(.douta(w_n138_0[0]),.doutb(w_n138_0[1]),.doutc(w_n138_0[2]),.din(n138));
	jspl3 jspl3_w_n138_1(.douta(w_n138_1[0]),.doutb(w_n138_1[1]),.doutc(w_n138_1[2]),.din(w_n138_0[0]));
	jspl3 jspl3_w_n138_2(.douta(w_n138_2[0]),.doutb(w_n138_2[1]),.doutc(w_n138_2[2]),.din(w_n138_0[1]));
	jspl3 jspl3_w_n138_3(.douta(w_n138_3[0]),.doutb(w_n138_3[1]),.doutc(w_n138_3[2]),.din(w_n138_0[2]));
	jspl jspl_w_n138_4(.douta(w_n138_4[0]),.doutb(w_n138_4[1]),.din(w_n138_1[0]));
	jspl3 jspl3_w_n139_0(.douta(w_n139_0[0]),.doutb(w_n139_0[1]),.doutc(w_n139_0[2]),.din(n139));
	jspl jspl_w_n139_1(.douta(w_n139_1[0]),.doutb(w_n139_1[1]),.din(w_n139_0[0]));
	jspl3 jspl3_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.doutc(w_n140_0[2]),.din(n140));
	jspl3 jspl3_w_n140_1(.douta(w_n140_1[0]),.doutb(w_n140_1[1]),.doutc(w_n140_1[2]),.din(w_n140_0[0]));
	jspl3 jspl3_w_n140_2(.douta(w_n140_2[0]),.doutb(w_n140_2[1]),.doutc(w_n140_2[2]),.din(w_n140_0[1]));
	jspl jspl_w_n140_3(.douta(w_n140_3[0]),.doutb(w_n140_3[1]),.din(w_n140_0[2]));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl3 jspl3_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.doutc(w_n142_0[2]),.din(n142));
	jspl3 jspl3_w_n142_1(.douta(w_n142_1[0]),.doutb(w_n142_1[1]),.doutc(w_n142_1[2]),.din(w_n142_0[0]));
	jspl jspl_w_n142_2(.douta(w_n142_2[0]),.doutb(w_n142_2[1]),.din(w_n142_0[1]));
	jspl3 jspl3_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.doutc(w_n143_0[2]),.din(n143));
	jspl jspl_w_n143_1(.douta(w_n143_1[0]),.doutb(w_n143_1[1]),.din(w_n143_0[0]));
	jspl3 jspl3_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.doutc(w_n144_0[2]),.din(n144));
	jspl3 jspl3_w_n144_1(.douta(w_n144_1[0]),.doutb(w_n144_1[1]),.doutc(w_n144_1[2]),.din(w_n144_0[0]));
	jspl3 jspl3_w_n144_2(.douta(w_n144_2[0]),.doutb(w_n144_2[1]),.doutc(w_n144_2[2]),.din(w_n144_0[1]));
	jspl3 jspl3_w_n144_3(.douta(w_n144_3[0]),.doutb(w_n144_3[1]),.doutc(w_n144_3[2]),.din(w_n144_0[2]));
	jspl3 jspl3_w_n144_4(.douta(w_n144_4[0]),.doutb(w_n144_4[1]),.doutc(w_n144_4[2]),.din(w_n144_1[0]));
	jspl3 jspl3_w_n144_5(.douta(w_n144_5[0]),.doutb(w_n144_5[1]),.doutc(w_n144_5[2]),.din(w_n144_1[1]));
	jspl3 jspl3_w_n144_6(.douta(w_n144_6[0]),.doutb(w_n144_6[1]),.doutc(w_n144_6[2]),.din(w_n144_1[2]));
	jspl3 jspl3_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.doutc(w_n145_0[2]),.din(n145));
	jspl3 jspl3_w_n145_1(.douta(w_n145_1[0]),.doutb(w_n145_1[1]),.doutc(w_n145_1[2]),.din(w_n145_0[0]));
	jspl3 jspl3_w_n145_2(.douta(w_n145_2[0]),.doutb(w_n145_2[1]),.doutc(w_n145_2[2]),.din(w_n145_0[1]));
	jspl jspl_w_n145_3(.douta(w_n145_3[0]),.doutb(w_n145_3[1]),.din(w_n145_0[2]));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.doutc(w_n147_0[2]),.din(n147));
	jspl3 jspl3_w_n147_1(.douta(w_n147_1[0]),.doutb(w_n147_1[1]),.doutc(w_n147_1[2]),.din(w_n147_0[0]));
	jspl jspl_w_n147_2(.douta(w_n147_2[0]),.doutb(w_n147_2[1]),.din(w_n147_0[1]));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl jspl_w_n148_1(.douta(w_n148_1[0]),.doutb(w_n148_1[1]),.din(w_n148_0[0]));
	jspl jspl_w_n150_0(.douta(w_n150_0[0]),.doutb(w_n150_0[1]),.din(n150));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_n151_0[1]),.doutc(w_n151_0[2]),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_n151_1[1]),.doutc(w_n151_1[2]),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_n151_2[0]),.doutb(w_n151_2[1]),.doutc(w_n151_2[2]),.din(w_n151_0[1]));
	jspl3 jspl3_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.doutc(w_n152_0[2]),.din(n152));
	jspl3 jspl3_w_n152_1(.douta(w_n152_1[0]),.doutb(w_n152_1[1]),.doutc(w_n152_1[2]),.din(w_n152_0[0]));
	jspl3 jspl3_w_n152_2(.douta(w_n152_2[0]),.doutb(w_n152_2[1]),.doutc(w_n152_2[2]),.din(w_n152_0[1]));
	jspl3 jspl3_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.doutc(w_n154_0[2]),.din(n154));
	jspl3 jspl3_w_n154_1(.douta(w_n154_1[0]),.doutb(w_n154_1[1]),.doutc(w_n154_1[2]),.din(w_n154_0[0]));
	jspl3 jspl3_w_n154_2(.douta(w_n154_2[0]),.doutb(w_n154_2[1]),.doutc(w_n154_2[2]),.din(w_n154_0[1]));
	jspl3 jspl3_w_n154_3(.douta(w_n154_3[0]),.doutb(w_n154_3[1]),.doutc(w_n154_3[2]),.din(w_n154_0[2]));
	jspl3 jspl3_w_n154_4(.douta(w_n154_4[0]),.doutb(w_n154_4[1]),.doutc(w_n154_4[2]),.din(w_n154_1[0]));
	jspl3 jspl3_w_n154_5(.douta(w_n154_5[0]),.doutb(w_n154_5[1]),.doutc(w_n154_5[2]),.din(w_n154_1[1]));
	jspl3 jspl3_w_n154_6(.douta(w_n154_6[0]),.doutb(w_n154_6[1]),.doutc(w_n154_6[2]),.din(w_n154_1[2]));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl3 jspl3_w_n155_1(.douta(w_n155_1[0]),.doutb(w_n155_1[1]),.doutc(w_n155_1[2]),.din(w_n155_0[0]));
	jspl3 jspl3_w_n155_2(.douta(w_n155_2[0]),.doutb(w_n155_2[1]),.doutc(w_n155_2[2]),.din(w_n155_0[1]));
	jspl3 jspl3_w_n155_3(.douta(w_n155_3[0]),.doutb(w_n155_3[1]),.doutc(w_n155_3[2]),.din(w_n155_0[2]));
	jspl3 jspl3_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.doutc(w_n157_0[2]),.din(n157));
	jspl3 jspl3_w_n157_1(.douta(w_n157_1[0]),.doutb(w_n157_1[1]),.doutc(w_n157_1[2]),.din(w_n157_0[0]));
	jspl3 jspl3_w_n157_2(.douta(w_n157_2[0]),.doutb(w_n157_2[1]),.doutc(w_n157_2[2]),.din(w_n157_0[1]));
	jspl jspl_w_n157_3(.douta(w_n157_3[0]),.doutb(w_n157_3[1]),.din(w_n157_0[2]));
	jspl3 jspl3_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.doutc(w_n158_0[2]),.din(n158));
	jspl3 jspl3_w_n158_1(.douta(w_n158_1[0]),.doutb(w_n158_1[1]),.doutc(w_n158_1[2]),.din(w_n158_0[0]));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl3 jspl3_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.doutc(w_n160_0[2]),.din(n160));
	jspl3 jspl3_w_n160_1(.douta(w_n160_1[0]),.doutb(w_n160_1[1]),.doutc(w_n160_1[2]),.din(w_n160_0[0]));
	jspl3 jspl3_w_n160_2(.douta(w_n160_2[0]),.doutb(w_n160_2[1]),.doutc(w_n160_2[2]),.din(w_n160_0[1]));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_n161_0[2]),.din(n161));
	jspl3 jspl3_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.doutc(w_n162_0[2]),.din(n162));
	jspl3 jspl3_w_n162_1(.douta(w_n162_1[0]),.doutb(w_n162_1[1]),.doutc(w_n162_1[2]),.din(w_n162_0[0]));
	jspl jspl_w_n162_2(.douta(w_n162_2[0]),.doutb(w_n162_2[1]),.din(w_n162_0[1]));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.doutc(w_n165_0[2]),.din(n165));
	jspl3 jspl3_w_n165_1(.douta(w_n165_1[0]),.doutb(w_n165_1[1]),.doutc(w_n165_1[2]),.din(w_n165_0[0]));
	jspl3 jspl3_w_n165_2(.douta(w_n165_2[0]),.doutb(w_n165_2[1]),.doutc(w_n165_2[2]),.din(w_n165_0[1]));
	jspl3 jspl3_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_n166_1[1]),.doutc(w_n166_1[2]),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_n166_2[2]),.din(w_n166_0[1]));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.doutc(w_n167_0[2]),.din(n167));
	jspl3 jspl3_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.doutc(w_n167_1[2]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n167_2(.douta(w_n167_2[0]),.doutb(w_n167_2[1]),.doutc(w_n167_2[2]),.din(w_n167_0[1]));
	jspl3 jspl3_w_n167_3(.douta(w_n167_3[0]),.doutb(w_n167_3[1]),.doutc(w_n167_3[2]),.din(w_n167_0[2]));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl3 jspl3_w_n168_1(.douta(w_n168_1[0]),.doutb(w_n168_1[1]),.doutc(w_n168_1[2]),.din(w_n168_0[0]));
	jspl jspl_w_n168_2(.douta(w_n168_2[0]),.doutb(w_n168_2[1]),.din(w_n168_0[1]));
	jspl3 jspl3_w_n169_0(.douta(w_n169_0[0]),.doutb(w_n169_0[1]),.doutc(w_n169_0[2]),.din(n169));
	jspl3 jspl3_w_n169_1(.douta(w_n169_1[0]),.doutb(w_n169_1[1]),.doutc(w_n169_1[2]),.din(w_n169_0[0]));
	jspl jspl_w_n169_2(.douta(w_n169_2[0]),.doutb(w_n169_2[1]),.din(w_n169_0[1]));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl3 jspl3_w_n170_1(.douta(w_n170_1[0]),.doutb(w_n170_1[1]),.doutc(w_n170_1[2]),.din(w_n170_0[0]));
	jspl3 jspl3_w_n170_2(.douta(w_n170_2[0]),.doutb(w_n170_2[1]),.doutc(w_n170_2[2]),.din(w_n170_0[1]));
	jspl jspl_w_n170_3(.douta(w_n170_3[0]),.doutb(w_n170_3[1]),.din(w_n170_0[2]));
	jspl3 jspl3_w_n171_0(.douta(w_n171_0[0]),.doutb(w_n171_0[1]),.doutc(w_n171_0[2]),.din(n171));
	jspl3 jspl3_w_n171_1(.douta(w_n171_1[0]),.doutb(w_n171_1[1]),.doutc(w_n171_1[2]),.din(w_n171_0[0]));
	jspl3 jspl3_w_n171_2(.douta(w_n171_2[0]),.doutb(w_n171_2[1]),.doutc(w_n171_2[2]),.din(w_n171_0[1]));
	jspl3 jspl3_w_n171_3(.douta(w_n171_3[0]),.doutb(w_n171_3[1]),.doutc(w_n171_3[2]),.din(w_n171_0[2]));
	jspl jspl_w_n171_4(.douta(w_n171_4[0]),.doutb(w_n171_4[1]),.din(w_n171_1[0]));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl3 jspl3_w_n173_1(.douta(w_n173_1[0]),.doutb(w_n173_1[1]),.doutc(w_n173_1[2]),.din(w_n173_0[0]));
	jspl3 jspl3_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.doutc(w_n174_0[2]),.din(n174));
	jspl3 jspl3_w_n174_1(.douta(w_n174_1[0]),.doutb(w_n174_1[1]),.doutc(w_n174_1[2]),.din(w_n174_0[0]));
	jspl3 jspl3_w_n174_2(.douta(w_n174_2[0]),.doutb(w_n174_2[1]),.doutc(w_n174_2[2]),.din(w_n174_0[1]));
	jspl3 jspl3_w_n174_3(.douta(w_n174_3[0]),.doutb(w_n174_3[1]),.doutc(w_n174_3[2]),.din(w_n174_0[2]));
	jspl3 jspl3_w_n174_4(.douta(w_n174_4[0]),.doutb(w_n174_4[1]),.doutc(w_n174_4[2]),.din(w_n174_1[0]));
	jspl3 jspl3_w_n174_5(.douta(w_n174_5[0]),.doutb(w_n174_5[1]),.doutc(w_n174_5[2]),.din(w_n174_1[1]));
	jspl3 jspl3_w_n174_6(.douta(w_n174_6[0]),.doutb(w_n174_6[1]),.doutc(w_n174_6[2]),.din(w_n174_1[2]));
	jspl3 jspl3_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.doutc(w_n176_0[2]),.din(n176));
	jspl3 jspl3_w_n176_1(.douta(w_n176_1[0]),.doutb(w_n176_1[1]),.doutc(w_n176_1[2]),.din(w_n176_0[0]));
	jspl jspl_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.doutc(w_n180_0[2]),.din(n180));
	jspl jspl_w_n180_1(.douta(w_n180_1[0]),.doutb(w_n180_1[1]),.din(w_n180_0[0]));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n182_2(.douta(w_n182_2[0]),.doutb(w_n182_2[1]),.doutc(w_n182_2[2]),.din(w_n182_0[1]));
	jspl jspl_w_n182_3(.douta(w_n182_3[0]),.doutb(w_n182_3[1]),.din(w_n182_0[2]));
	jspl3 jspl3_w_n183_0(.douta(w_n183_0[0]),.doutb(w_n183_0[1]),.doutc(w_n183_0[2]),.din(n183));
	jspl3 jspl3_w_n184_0(.douta(w_n184_0[0]),.doutb(w_n184_0[1]),.doutc(w_n184_0[2]),.din(n184));
	jspl3 jspl3_w_n184_1(.douta(w_n184_1[0]),.doutb(w_n184_1[1]),.doutc(w_n184_1[2]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n184_2(.douta(w_n184_2[0]),.doutb(w_n184_2[1]),.doutc(w_n184_2[2]),.din(w_n184_0[1]));
	jspl3 jspl3_w_n184_3(.douta(w_n184_3[0]),.doutb(w_n184_3[1]),.doutc(w_n184_3[2]),.din(w_n184_0[2]));
	jspl3 jspl3_w_n184_4(.douta(w_n184_4[0]),.doutb(w_n184_4[1]),.doutc(w_n184_4[2]),.din(w_n184_1[0]));
	jspl3 jspl3_w_n184_5(.douta(w_n184_5[0]),.doutb(w_n184_5[1]),.doutc(w_n184_5[2]),.din(w_n184_1[1]));
	jspl3 jspl3_w_n184_6(.douta(w_n184_6[0]),.doutb(w_n184_6[1]),.doutc(w_n184_6[2]),.din(w_n184_1[2]));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.doutc(w_n185_0[2]),.din(n185));
	jspl3 jspl3_w_n185_1(.douta(w_n185_1[0]),.doutb(w_n185_1[1]),.doutc(w_n185_1[2]),.din(w_n185_0[0]));
	jspl3 jspl3_w_n185_2(.douta(w_n185_2[0]),.doutb(w_n185_2[1]),.doutc(w_n185_2[2]),.din(w_n185_0[1]));
	jspl3 jspl3_w_n185_3(.douta(w_n185_3[0]),.doutb(w_n185_3[1]),.doutc(w_n185_3[2]),.din(w_n185_0[2]));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl3 jspl3_w_n187_0(.douta(w_n187_0[0]),.doutb(w_n187_0[1]),.doutc(w_n187_0[2]),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_n187_1[0]),.doutb(w_n187_1[1]),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n187_2(.douta(w_n187_2[0]),.doutb(w_n187_2[1]),.din(w_n187_0[1]));
	jspl3 jspl3_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.doutc(w_n188_0[2]),.din(n188));
	jspl3 jspl3_w_n188_1(.douta(w_n188_1[0]),.doutb(w_n188_1[1]),.doutc(w_n188_1[2]),.din(w_n188_0[0]));
	jspl jspl_w_n188_2(.douta(w_n188_2[0]),.doutb(w_n188_2[1]),.din(w_n188_0[1]));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.doutc(w_n190_0[2]),.din(n190));
	jspl3 jspl3_w_n190_1(.douta(w_n190_1[0]),.doutb(w_n190_1[1]),.doutc(w_n190_1[2]),.din(w_n190_0[0]));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl3 jspl3_w_n191_1(.douta(w_n191_1[0]),.doutb(w_n191_1[1]),.doutc(w_n191_1[2]),.din(w_n191_0[0]));
	jspl3 jspl3_w_n191_2(.douta(w_n191_2[0]),.doutb(w_n191_2[1]),.doutc(w_n191_2[2]),.din(w_n191_0[1]));
	jspl3 jspl3_w_n191_3(.douta(w_n191_3[0]),.doutb(w_n191_3[1]),.doutc(w_n191_3[2]),.din(w_n191_0[2]));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.doutc(w_n192_0[2]),.din(n192));
	jspl3 jspl3_w_n192_1(.douta(w_n192_1[0]),.doutb(w_n192_1[1]),.doutc(w_n192_1[2]),.din(w_n192_0[0]));
	jspl3 jspl3_w_n192_2(.douta(w_n192_2[0]),.doutb(w_n192_2[1]),.doutc(w_n192_2[2]),.din(w_n192_0[1]));
	jspl jspl_w_n192_3(.douta(w_n192_3[0]),.doutb(w_n192_3[1]),.din(w_n192_0[2]));
	jspl3 jspl3_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.doutc(w_n193_0[2]),.din(n193));
	jspl3 jspl3_w_n193_1(.douta(w_n193_1[0]),.doutb(w_n193_1[1]),.doutc(w_n193_1[2]),.din(w_n193_0[0]));
	jspl jspl_w_n193_2(.douta(w_n193_2[0]),.doutb(w_n193_2[1]),.din(w_n193_0[1]));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.doutc(w_n194_0[2]),.din(n194));
	jspl3 jspl3_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.doutc(w_n195_0[2]),.din(n195));
	jspl3 jspl3_w_n195_1(.douta(w_n195_1[0]),.doutb(w_n195_1[1]),.doutc(w_n195_1[2]),.din(w_n195_0[0]));
	jspl jspl_w_n195_2(.douta(w_n195_2[0]),.doutb(w_n195_2[1]),.din(w_n195_0[1]));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl3 jspl3_w_n197_1(.douta(w_n197_1[0]),.doutb(w_n197_1[1]),.doutc(w_n197_1[2]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n197_2(.douta(w_n197_2[0]),.doutb(w_n197_2[1]),.doutc(w_n197_2[2]),.din(w_n197_0[1]));
	jspl jspl_w_n197_3(.douta(w_n197_3[0]),.doutb(w_n197_3[1]),.din(w_n197_0[2]));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_n198_0[2]),.din(n198));
	jspl jspl_w_n198_1(.douta(w_n198_1[0]),.doutb(w_n198_1[1]),.din(w_n198_0[0]));
	jspl3 jspl3_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.doutc(w_n203_0[2]),.din(n203));
	jspl jspl_w_n203_1(.douta(w_n203_1[0]),.doutb(w_n203_1[1]),.din(w_n203_0[0]));
	jspl3 jspl3_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.doutc(w_n204_0[2]),.din(n204));
	jspl3 jspl3_w_n204_1(.douta(w_n204_1[0]),.doutb(w_n204_1[1]),.doutc(w_n204_1[2]),.din(w_n204_0[0]));
	jspl3 jspl3_w_n204_2(.douta(w_n204_2[0]),.doutb(w_n204_2[1]),.doutc(w_n204_2[2]),.din(w_n204_0[1]));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl3 jspl3_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.doutc(w_n206_0[2]),.din(n206));
	jspl3 jspl3_w_n206_1(.douta(w_n206_1[0]),.doutb(w_n206_1[1]),.doutc(w_n206_1[2]),.din(w_n206_0[0]));
	jspl jspl_w_n206_2(.douta(w_n206_2[0]),.doutb(w_n206_2[1]),.din(w_n206_0[1]));
	jspl3 jspl3_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.doutc(w_n207_0[2]),.din(n207));
	jspl3 jspl3_w_n207_1(.douta(w_n207_1[0]),.doutb(w_n207_1[1]),.doutc(w_n207_1[2]),.din(w_n207_0[0]));
	jspl3 jspl3_w_n207_2(.douta(w_n207_2[0]),.doutb(w_n207_2[1]),.doutc(w_n207_2[2]),.din(w_n207_0[1]));
	jspl jspl_w_n207_3(.douta(w_n207_3[0]),.doutb(w_n207_3[1]),.din(w_n207_0[2]));
	jspl jspl_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.din(n212));
	jspl3 jspl3_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.doutc(w_n213_0[2]),.din(n213));
	jspl3 jspl3_w_n213_1(.douta(w_n213_1[0]),.doutb(w_n213_1[1]),.doutc(w_n213_1[2]),.din(w_n213_0[0]));
	jspl3 jspl3_w_n213_2(.douta(w_n213_2[0]),.doutb(w_n213_2[1]),.doutc(w_n213_2[2]),.din(w_n213_0[1]));
	jspl jspl_w_n213_3(.douta(w_n213_3[0]),.doutb(w_n213_3[1]),.din(w_n213_0[2]));
	jspl jspl_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.din(n214));
	jspl3 jspl3_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.doutc(w_n215_0[2]),.din(n215));
	jspl3 jspl3_w_n215_1(.douta(w_n215_1[0]),.doutb(w_n215_1[1]),.doutc(w_n215_1[2]),.din(w_n215_0[0]));
	jspl3 jspl3_w_n215_2(.douta(w_n215_2[0]),.doutb(w_n215_2[1]),.doutc(w_n215_2[2]),.din(w_n215_0[1]));
	jspl3 jspl3_w_n215_3(.douta(w_n215_3[0]),.doutb(w_n215_3[1]),.doutc(w_n215_3[2]),.din(w_n215_0[2]));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.doutc(w_n216_0[2]),.din(n216));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl3 jspl3_w_n217_1(.douta(w_n217_1[0]),.doutb(w_n217_1[1]),.doutc(w_n217_1[2]),.din(w_n217_0[0]));
	jspl3 jspl3_w_n217_2(.douta(w_n217_2[0]),.doutb(w_n217_2[1]),.doutc(w_n217_2[2]),.din(w_n217_0[1]));
	jspl3 jspl3_w_n217_3(.douta(w_n217_3[0]),.doutb(w_n217_3[1]),.doutc(w_n217_3[2]),.din(w_n217_0[2]));
	jspl jspl_w_n217_4(.douta(w_n217_4[0]),.doutb(w_n217_4[1]),.din(w_n217_1[0]));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_n218_0[2]),.din(n218));
	jspl3 jspl3_w_n218_1(.douta(w_n218_1[0]),.doutb(w_n218_1[1]),.doutc(w_n218_1[2]),.din(w_n218_0[0]));
	jspl3 jspl3_w_n218_2(.douta(w_n218_2[0]),.doutb(w_n218_2[1]),.doutc(w_n218_2[2]),.din(w_n218_0[1]));
	jspl3 jspl3_w_n218_3(.douta(w_n218_3[0]),.doutb(w_n218_3[1]),.doutc(w_n218_3[2]),.din(w_n218_0[2]));
	jspl3 jspl3_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.doutc(w_n221_0[2]),.din(n221));
	jspl3 jspl3_w_n221_1(.douta(w_n221_1[0]),.doutb(w_n221_1[1]),.doutc(w_n221_1[2]),.din(w_n221_0[0]));
	jspl3 jspl3_w_n221_2(.douta(w_n221_2[0]),.doutb(w_n221_2[1]),.doutc(w_n221_2[2]),.din(w_n221_0[1]));
	jspl3 jspl3_w_n221_3(.douta(w_n221_3[0]),.doutb(w_n221_3[1]),.doutc(w_n221_3[2]),.din(w_n221_0[2]));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.doutc(w_n222_0[2]),.din(n222));
	jspl3 jspl3_w_n222_1(.douta(w_n222_1[0]),.doutb(w_n222_1[1]),.doutc(w_n222_1[2]),.din(w_n222_0[0]));
	jspl3 jspl3_w_n222_2(.douta(w_n222_2[0]),.doutb(w_n222_2[1]),.doutc(w_n222_2[2]),.din(w_n222_0[1]));
	jspl jspl_w_n222_3(.douta(w_n222_3[0]),.doutb(w_n222_3[1]),.din(w_n222_0[2]));
	jspl3 jspl3_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.doutc(w_n223_0[2]),.din(n223));
	jspl3 jspl3_w_n223_1(.douta(w_n223_1[0]),.doutb(w_n223_1[1]),.doutc(w_n223_1[2]),.din(w_n223_0[0]));
	jspl3 jspl3_w_n223_2(.douta(w_n223_2[0]),.doutb(w_n223_2[1]),.doutc(w_n223_2[2]),.din(w_n223_0[1]));
	jspl jspl_w_n223_3(.douta(w_n223_3[0]),.doutb(w_n223_3[1]),.din(w_n223_0[2]));
	jspl3 jspl3_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.doutc(w_n224_0[2]),.din(n224));
	jspl3 jspl3_w_n224_1(.douta(w_n224_1[0]),.doutb(w_n224_1[1]),.doutc(w_n224_1[2]),.din(w_n224_0[0]));
	jspl3 jspl3_w_n224_2(.douta(w_n224_2[0]),.doutb(w_n224_2[1]),.doutc(w_n224_2[2]),.din(w_n224_0[1]));
	jspl3 jspl3_w_n224_3(.douta(w_n224_3[0]),.doutb(w_n224_3[1]),.doutc(w_n224_3[2]),.din(w_n224_0[2]));
	jspl3 jspl3_w_n224_4(.douta(w_n224_4[0]),.doutb(w_n224_4[1]),.doutc(w_n224_4[2]),.din(w_n224_1[0]));
	jspl jspl_w_n224_5(.douta(w_n224_5[0]),.doutb(w_n224_5[1]),.din(w_n224_1[1]));
	jspl3 jspl3_w_n226_0(.douta(w_n226_0[0]),.doutb(w_n226_0[1]),.doutc(w_n226_0[2]),.din(n226));
	jspl3 jspl3_w_n226_1(.douta(w_n226_1[0]),.doutb(w_n226_1[1]),.doutc(w_n226_1[2]),.din(w_n226_0[0]));
	jspl3 jspl3_w_n226_2(.douta(w_n226_2[0]),.doutb(w_n226_2[1]),.doutc(w_n226_2[2]),.din(w_n226_0[1]));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.din(n229));
	jspl3 jspl3_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.doutc(w_n230_0[2]),.din(n230));
	jspl3 jspl3_w_n230_1(.douta(w_n230_1[0]),.doutb(w_n230_1[1]),.doutc(w_n230_1[2]),.din(w_n230_0[0]));
	jspl3 jspl3_w_n230_2(.douta(w_n230_2[0]),.doutb(w_n230_2[1]),.doutc(w_n230_2[2]),.din(w_n230_0[1]));
	jspl jspl_w_n230_3(.douta(w_n230_3[0]),.doutb(w_n230_3[1]),.din(w_n230_0[2]));
	jspl3 jspl3_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.doutc(w_n231_0[2]),.din(n231));
	jspl jspl_w_n231_1(.douta(w_n231_1[0]),.doutb(w_n231_1[1]),.din(w_n231_0[0]));
	jspl3 jspl3_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.doutc(w_n232_0[2]),.din(n232));
	jspl3 jspl3_w_n232_1(.douta(w_n232_1[0]),.doutb(w_n232_1[1]),.doutc(w_n232_1[2]),.din(w_n232_0[0]));
	jspl3 jspl3_w_n232_2(.douta(w_n232_2[0]),.doutb(w_n232_2[1]),.doutc(w_n232_2[2]),.din(w_n232_0[1]));
	jspl3 jspl3_w_n232_3(.douta(w_n232_3[0]),.doutb(w_n232_3[1]),.doutc(w_n232_3[2]),.din(w_n232_0[2]));
	jspl3 jspl3_w_n232_4(.douta(w_n232_4[0]),.doutb(w_n232_4[1]),.doutc(w_n232_4[2]),.din(w_n232_1[0]));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl3 jspl3_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.doutc(w_n233_1[2]),.din(w_n233_0[0]));
	jspl jspl_w_n233_2(.douta(w_n233_2[0]),.doutb(w_n233_2[1]),.din(w_n233_0[1]));
	jspl3 jspl3_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.doutc(w_n234_0[2]),.din(n234));
	jspl3 jspl3_w_n235_0(.douta(w_n235_0[0]),.doutb(w_n235_0[1]),.doutc(w_n235_0[2]),.din(n235));
	jspl3 jspl3_w_n235_1(.douta(w_n235_1[0]),.doutb(w_n235_1[1]),.doutc(w_n235_1[2]),.din(w_n235_0[0]));
	jspl jspl_w_n235_2(.douta(w_n235_2[0]),.doutb(w_n235_2[1]),.din(w_n235_0[1]));
	jspl3 jspl3_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.doutc(w_n236_0[2]),.din(n236));
	jspl3 jspl3_w_n236_1(.douta(w_n236_1[0]),.doutb(w_n236_1[1]),.doutc(w_n236_1[2]),.din(w_n236_0[0]));
	jspl3 jspl3_w_n238_0(.douta(w_n238_0[0]),.doutb(w_n238_0[1]),.doutc(w_n238_0[2]),.din(n238));
	jspl3 jspl3_w_n238_1(.douta(w_n238_1[0]),.doutb(w_n238_1[1]),.doutc(w_n238_1[2]),.din(w_n238_0[0]));
	jspl jspl_w_n238_2(.douta(w_n238_2[0]),.doutb(w_n238_2[1]),.din(w_n238_0[1]));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(n239));
	jspl3 jspl3_w_n240_0(.douta(w_n240_0[0]),.doutb(w_n240_0[1]),.doutc(w_n240_0[2]),.din(n240));
	jspl3 jspl3_w_n240_1(.douta(w_n240_1[0]),.doutb(w_n240_1[1]),.doutc(w_n240_1[2]),.din(w_n240_0[0]));
	jspl jspl_w_n240_2(.douta(w_n240_2[0]),.doutb(w_n240_2[1]),.din(w_n240_0[1]));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(n241));
	jspl3 jspl3_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.doutc(w_n244_0[2]),.din(n244));
	jspl3 jspl3_w_n244_1(.douta(w_n244_1[0]),.doutb(w_n244_1[1]),.doutc(w_n244_1[2]),.din(w_n244_0[0]));
	jspl3 jspl3_w_n244_2(.douta(w_n244_2[0]),.doutb(w_n244_2[1]),.doutc(w_n244_2[2]),.din(w_n244_0[1]));
	jspl jspl_w_n244_3(.douta(w_n244_3[0]),.doutb(w_n244_3[1]),.din(w_n244_0[2]));
	jspl3 jspl3_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.doutc(w_n245_0[2]),.din(n245));
	jspl3 jspl3_w_n245_1(.douta(w_n245_1[0]),.doutb(w_n245_1[1]),.doutc(w_n245_1[2]),.din(w_n245_0[0]));
	jspl jspl_w_n245_2(.douta(w_n245_2[0]),.doutb(w_n245_2[1]),.din(w_n245_0[1]));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl3 jspl3_w_n248_0(.douta(w_n248_0[0]),.doutb(w_n248_0[1]),.doutc(w_n248_0[2]),.din(n248));
	jspl3 jspl3_w_n248_1(.douta(w_n248_1[0]),.doutb(w_n248_1[1]),.doutc(w_n248_1[2]),.din(w_n248_0[0]));
	jspl3 jspl3_w_n248_2(.douta(w_n248_2[0]),.doutb(w_n248_2[1]),.doutc(w_n248_2[2]),.din(w_n248_0[1]));
	jspl3 jspl3_w_n248_3(.douta(w_n248_3[0]),.doutb(w_n248_3[1]),.doutc(w_n248_3[2]),.din(w_n248_0[2]));
	jspl3 jspl3_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.doutc(w_n249_0[2]),.din(n249));
	jspl3 jspl3_w_n249_1(.douta(w_n249_1[0]),.doutb(w_n249_1[1]),.doutc(w_n249_1[2]),.din(w_n249_0[0]));
	jspl jspl_w_n249_2(.douta(w_n249_2[0]),.doutb(w_n249_2[1]),.din(w_n249_0[1]));
	jspl3 jspl3_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.doutc(w_n250_0[2]),.din(n250));
	jspl3 jspl3_w_n250_1(.douta(w_n250_1[0]),.doutb(w_n250_1[1]),.doutc(w_n250_1[2]),.din(w_n250_0[0]));
	jspl3 jspl3_w_n250_2(.douta(w_n250_2[0]),.doutb(w_n250_2[1]),.doutc(w_n250_2[2]),.din(w_n250_0[1]));
	jspl3 jspl3_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.doutc(w_n251_0[2]),.din(n251));
	jspl3 jspl3_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.doutc(w_n252_0[2]),.din(n252));
	jspl3 jspl3_w_n252_1(.douta(w_n252_1[0]),.doutb(w_n252_1[1]),.doutc(w_n252_1[2]),.din(w_n252_0[0]));
	jspl3 jspl3_w_n252_2(.douta(w_n252_2[0]),.doutb(w_n252_2[1]),.doutc(w_n252_2[2]),.din(w_n252_0[1]));
	jspl3 jspl3_w_n252_3(.douta(w_n252_3[0]),.doutb(w_n252_3[1]),.doutc(w_n252_3[2]),.din(w_n252_0[2]));
	jspl jspl_w_n252_4(.douta(w_n252_4[0]),.doutb(w_n252_4[1]),.din(w_n252_1[0]));
	jspl3 jspl3_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.doutc(w_n253_0[2]),.din(n253));
	jspl3 jspl3_w_n253_1(.douta(w_n253_1[0]),.doutb(w_n253_1[1]),.doutc(w_n253_1[2]),.din(w_n253_0[0]));
	jspl3 jspl3_w_n253_2(.douta(w_n253_2[0]),.doutb(w_n253_2[1]),.doutc(w_n253_2[2]),.din(w_n253_0[1]));
	jspl3 jspl3_w_n253_3(.douta(w_n253_3[0]),.doutb(w_n253_3[1]),.doutc(w_n253_3[2]),.din(w_n253_0[2]));
	jspl3 jspl3_w_n253_4(.douta(w_n253_4[0]),.doutb(w_n253_4[1]),.doutc(w_n253_4[2]),.din(w_n253_1[0]));
	jspl3 jspl3_w_n253_5(.douta(w_n253_5[0]),.doutb(w_n253_5[1]),.doutc(w_n253_5[2]),.din(w_n253_1[1]));
	jspl3 jspl3_w_n253_6(.douta(w_n253_6[0]),.doutb(w_n253_6[1]),.doutc(w_n253_6[2]),.din(w_n253_1[2]));
	jspl3 jspl3_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.doutc(w_n254_0[2]),.din(n254));
	jspl3 jspl3_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.doutc(w_n255_0[2]),.din(n255));
	jspl3 jspl3_w_n255_1(.douta(w_n255_1[0]),.doutb(w_n255_1[1]),.doutc(w_n255_1[2]),.din(w_n255_0[0]));
	jspl jspl_w_n255_2(.douta(w_n255_2[0]),.doutb(w_n255_2[1]),.din(w_n255_0[1]));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl3 jspl3_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.doutc(w_n261_0[2]),.din(n261));
	jspl3 jspl3_w_n261_1(.douta(w_n261_1[0]),.doutb(w_n261_1[1]),.doutc(w_n261_1[2]),.din(w_n261_0[0]));
	jspl3 jspl3_w_n261_2(.douta(w_n261_2[0]),.doutb(w_n261_2[1]),.doutc(w_n261_2[2]),.din(w_n261_0[1]));
	jspl3 jspl3_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.doutc(w_n262_0[2]),.din(n262));
	jspl3 jspl3_w_n262_1(.douta(w_n262_1[0]),.doutb(w_n262_1[1]),.doutc(w_n262_1[2]),.din(w_n262_0[0]));
	jspl3 jspl3_w_n262_2(.douta(w_n262_2[0]),.doutb(w_n262_2[1]),.doutc(w_n262_2[2]),.din(w_n262_0[1]));
	jspl3 jspl3_w_n262_3(.douta(w_n262_3[0]),.doutb(w_n262_3[1]),.doutc(w_n262_3[2]),.din(w_n262_0[2]));
	jspl3 jspl3_w_n262_4(.douta(w_n262_4[0]),.doutb(w_n262_4[1]),.doutc(w_n262_4[2]),.din(w_n262_1[0]));
	jspl jspl_w_n262_5(.douta(w_n262_5[0]),.doutb(w_n262_5[1]),.din(w_n262_1[1]));
	jspl3 jspl3_w_n263_0(.douta(w_n263_0[0]),.doutb(w_n263_0[1]),.doutc(w_n263_0[2]),.din(n263));
	jspl3 jspl3_w_n263_1(.douta(w_n263_1[0]),.doutb(w_n263_1[1]),.doutc(w_n263_1[2]),.din(w_n263_0[0]));
	jspl3 jspl3_w_n263_2(.douta(w_n263_2[0]),.doutb(w_n263_2[1]),.doutc(w_n263_2[2]),.din(w_n263_0[1]));
	jspl3 jspl3_w_n263_3(.douta(w_n263_3[0]),.doutb(w_n263_3[1]),.doutc(w_n263_3[2]),.din(w_n263_0[2]));
	jspl jspl_w_n263_4(.douta(w_n263_4[0]),.doutb(w_n263_4[1]),.din(w_n263_1[0]));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl3 jspl3_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.doutc(w_n265_0[2]),.din(n265));
	jspl3 jspl3_w_n265_1(.douta(w_n265_1[0]),.doutb(w_n265_1[1]),.doutc(w_n265_1[2]),.din(w_n265_0[0]));
	jspl jspl_w_n265_2(.douta(w_n265_2[0]),.doutb(w_n265_2[1]),.din(w_n265_0[1]));
	jspl3 jspl3_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.doutc(w_n266_0[2]),.din(n266));
	jspl3 jspl3_w_n266_1(.douta(w_n266_1[0]),.doutb(w_n266_1[1]),.doutc(w_n266_1[2]),.din(w_n266_0[0]));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.doutc(w_n267_0[2]),.din(n267));
	jspl3 jspl3_w_n267_1(.douta(w_n267_1[0]),.doutb(w_n267_1[1]),.doutc(w_n267_1[2]),.din(w_n267_0[0]));
	jspl3 jspl3_w_n267_2(.douta(w_n267_2[0]),.doutb(w_n267_2[1]),.doutc(w_n267_2[2]),.din(w_n267_0[1]));
	jspl jspl_w_n267_3(.douta(w_n267_3[0]),.doutb(w_n267_3[1]),.din(w_n267_0[2]));
	jspl3 jspl3_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.doutc(w_n268_0[2]),.din(n268));
	jspl3 jspl3_w_n268_1(.douta(w_n268_1[0]),.doutb(w_n268_1[1]),.doutc(w_n268_1[2]),.din(w_n268_0[0]));
	jspl jspl_w_n268_2(.douta(w_n268_2[0]),.doutb(w_n268_2[1]),.din(w_n268_0[1]));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.doutc(w_n269_1[2]),.din(w_n269_0[0]));
	jspl3 jspl3_w_n269_2(.douta(w_n269_2[0]),.doutb(w_n269_2[1]),.doutc(w_n269_2[2]),.din(w_n269_0[1]));
	jspl jspl_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.din(n273));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl3 jspl3_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.doutc(w_n275_0[2]),.din(n275));
	jspl3 jspl3_w_n275_1(.douta(w_n275_1[0]),.doutb(w_n275_1[1]),.doutc(w_n275_1[2]),.din(w_n275_0[0]));
	jspl jspl_w_n275_2(.douta(w_n275_2[0]),.doutb(w_n275_2[1]),.din(w_n275_0[1]));
	jspl3 jspl3_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.doutc(w_n276_0[2]),.din(n276));
	jspl3 jspl3_w_n276_1(.douta(w_n276_1[0]),.doutb(w_n276_1[1]),.doutc(w_n276_1[2]),.din(w_n276_0[0]));
	jspl3 jspl3_w_n276_2(.douta(w_n276_2[0]),.doutb(w_n276_2[1]),.doutc(w_n276_2[2]),.din(w_n276_0[1]));
	jspl3 jspl3_w_n276_3(.douta(w_n276_3[0]),.doutb(w_n276_3[1]),.doutc(w_n276_3[2]),.din(w_n276_0[2]));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl3 jspl3_w_n278_0(.douta(w_n278_0[0]),.doutb(w_n278_0[1]),.doutc(w_n278_0[2]),.din(n278));
	jspl3 jspl3_w_n278_1(.douta(w_n278_1[0]),.doutb(w_n278_1[1]),.doutc(w_n278_1[2]),.din(w_n278_0[0]));
	jspl3 jspl3_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.doutc(w_n279_0[2]),.din(n279));
	jspl3 jspl3_w_n280_0(.douta(w_n280_0[0]),.doutb(w_n280_0[1]),.doutc(w_n280_0[2]),.din(n280));
	jspl3 jspl3_w_n280_1(.douta(w_n280_1[0]),.doutb(w_n280_1[1]),.doutc(w_n280_1[2]),.din(w_n280_0[0]));
	jspl3 jspl3_w_n280_2(.douta(w_n280_2[0]),.doutb(w_n280_2[1]),.doutc(w_n280_2[2]),.din(w_n280_0[1]));
	jspl3 jspl3_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.doutc(w_n281_0[2]),.din(n281));
	jspl3 jspl3_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.doutc(w_n282_0[2]),.din(n282));
	jspl3 jspl3_w_n282_1(.douta(w_n282_1[0]),.doutb(w_n282_1[1]),.doutc(w_n282_1[2]),.din(w_n282_0[0]));
	jspl3 jspl3_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.doutc(w_n283_0[2]),.din(n283));
	jspl3 jspl3_w_n283_1(.douta(w_n283_1[0]),.doutb(w_n283_1[1]),.doutc(w_n283_1[2]),.din(w_n283_0[0]));
	jspl jspl_w_n283_2(.douta(w_n283_2[0]),.doutb(w_n283_2[1]),.din(w_n283_0[1]));
	jspl3 jspl3_w_n286_0(.douta(w_n286_0[0]),.doutb(w_n286_0[1]),.doutc(w_n286_0[2]),.din(n286));
	jspl3 jspl3_w_n286_1(.douta(w_n286_1[0]),.doutb(w_n286_1[1]),.doutc(w_n286_1[2]),.din(w_n286_0[0]));
	jspl3 jspl3_w_n286_2(.douta(w_n286_2[0]),.doutb(w_n286_2[1]),.doutc(w_n286_2[2]),.din(w_n286_0[1]));
	jspl jspl_w_n286_3(.douta(w_n286_3[0]),.doutb(w_n286_3[1]),.din(w_n286_0[2]));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl3 jspl3_w_n288_1(.douta(w_n288_1[0]),.doutb(w_n288_1[1]),.doutc(w_n288_1[2]),.din(w_n288_0[0]));
	jspl jspl_w_n288_2(.douta(w_n288_2[0]),.doutb(w_n288_2[1]),.din(w_n288_0[1]));
	jspl3 jspl3_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.doutc(w_n289_0[2]),.din(n289));
	jspl jspl_w_n289_1(.douta(w_n289_1[0]),.doutb(w_n289_1[1]),.din(w_n289_0[0]));
	jspl3 jspl3_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.doutc(w_n290_0[2]),.din(n290));
	jspl3 jspl3_w_n290_1(.douta(w_n290_1[0]),.doutb(w_n290_1[1]),.doutc(w_n290_1[2]),.din(w_n290_0[0]));
	jspl3 jspl3_w_n290_2(.douta(w_n290_2[0]),.doutb(w_n290_2[1]),.doutc(w_n290_2[2]),.din(w_n290_0[1]));
	jspl3 jspl3_w_n290_3(.douta(w_n290_3[0]),.doutb(w_n290_3[1]),.doutc(w_n290_3[2]),.din(w_n290_0[2]));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl3 jspl3_w_n294_0(.douta(w_n294_0[0]),.doutb(w_n294_0[1]),.doutc(w_n294_0[2]),.din(n294));
	jspl3 jspl3_w_n294_1(.douta(w_n294_1[0]),.doutb(w_n294_1[1]),.doutc(w_n294_1[2]),.din(w_n294_0[0]));
	jspl3 jspl3_w_n294_2(.douta(w_n294_2[0]),.doutb(w_n294_2[1]),.doutc(w_n294_2[2]),.din(w_n294_0[1]));
	jspl3 jspl3_w_n294_3(.douta(w_n294_3[0]),.doutb(w_n294_3[1]),.doutc(w_n294_3[2]),.din(w_n294_0[2]));
	jspl3 jspl3_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.doutc(w_n295_0[2]),.din(n295));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl3 jspl3_w_n297_0(.douta(w_n297_0[0]),.doutb(w_n297_0[1]),.doutc(w_n297_0[2]),.din(n297));
	jspl3 jspl3_w_n297_1(.douta(w_n297_1[0]),.doutb(w_n297_1[1]),.doutc(w_n297_1[2]),.din(w_n297_0[0]));
	jspl jspl_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.din(n299));
	jspl3 jspl3_w_n300_0(.douta(w_n300_0[0]),.doutb(w_n300_0[1]),.doutc(w_n300_0[2]),.din(n300));
	jspl3 jspl3_w_n300_1(.douta(w_n300_1[0]),.doutb(w_n300_1[1]),.doutc(w_n300_1[2]),.din(w_n300_0[0]));
	jspl3 jspl3_w_n300_2(.douta(w_n300_2[0]),.doutb(w_n300_2[1]),.doutc(w_n300_2[2]),.din(w_n300_0[1]));
	jspl jspl_w_n300_3(.douta(w_n300_3[0]),.doutb(w_n300_3[1]),.din(w_n300_0[2]));
	jspl3 jspl3_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.doutc(w_n301_0[2]),.din(n301));
	jspl jspl_w_n301_1(.douta(w_n301_1[0]),.doutb(w_n301_1[1]),.din(w_n301_0[0]));
	jspl3 jspl3_w_n302_0(.douta(w_n302_0[0]),.doutb(w_n302_0[1]),.doutc(w_n302_0[2]),.din(n302));
	jspl3 jspl3_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.doutc(w_n303_0[2]),.din(n303));
	jspl3 jspl3_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.doutc(w_n305_0[2]),.din(n305));
	jspl3 jspl3_w_n305_1(.douta(w_n305_1[0]),.doutb(w_n305_1[1]),.doutc(w_n305_1[2]),.din(w_n305_0[0]));
	jspl3 jspl3_w_n305_2(.douta(w_n305_2[0]),.doutb(w_n305_2[1]),.doutc(w_n305_2[2]),.din(w_n305_0[1]));
	jspl jspl_w_n307_0(.douta(w_n307_0[0]),.doutb(w_n307_0[1]),.din(n307));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl3 jspl3_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.doutc(w_n309_0[2]),.din(n309));
	jspl3 jspl3_w_n309_1(.douta(w_n309_1[0]),.doutb(w_n309_1[1]),.doutc(w_n309_1[2]),.din(w_n309_0[0]));
	jspl3 jspl3_w_n309_2(.douta(w_n309_2[0]),.doutb(w_n309_2[1]),.doutc(w_n309_2[2]),.din(w_n309_0[1]));
	jspl3 jspl3_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.doutc(w_n310_0[2]),.din(n310));
	jspl3 jspl3_w_n310_1(.douta(w_n310_1[0]),.doutb(w_n310_1[1]),.doutc(w_n310_1[2]),.din(w_n310_0[0]));
	jspl3 jspl3_w_n310_2(.douta(w_n310_2[0]),.doutb(w_n310_2[1]),.doutc(w_n310_2[2]),.din(w_n310_0[1]));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.doutc(w_n311_0[2]),.din(n311));
	jspl3 jspl3_w_n311_1(.douta(w_n311_1[0]),.doutb(w_n311_1[1]),.doutc(w_n311_1[2]),.din(w_n311_0[0]));
	jspl3 jspl3_w_n311_2(.douta(w_n311_2[0]),.doutb(w_n311_2[1]),.doutc(w_n311_2[2]),.din(w_n311_0[1]));
	jspl jspl_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.din(n312));
	jspl3 jspl3_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.doutc(w_n313_0[2]),.din(n313));
	jspl3 jspl3_w_n313_1(.douta(w_n313_1[0]),.doutb(w_n313_1[1]),.doutc(w_n313_1[2]),.din(w_n313_0[0]));
	jspl3 jspl3_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.doutc(w_n314_0[2]),.din(n314));
	jspl3 jspl3_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.doutc(w_n315_0[2]),.din(n315));
	jspl3 jspl3_w_n315_1(.douta(w_n315_1[0]),.doutb(w_n315_1[1]),.doutc(w_n315_1[2]),.din(w_n315_0[0]));
	jspl jspl_w_n315_2(.douta(w_n315_2[0]),.doutb(w_n315_2[1]),.din(w_n315_0[1]));
	jspl3 jspl3_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.doutc(w_n316_0[2]),.din(n316));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl3 jspl3_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.doutc(w_n321_0[2]),.din(n321));
	jspl3 jspl3_w_n321_1(.douta(w_n321_1[0]),.doutb(w_n321_1[1]),.doutc(w_n321_1[2]),.din(w_n321_0[0]));
	jspl3 jspl3_w_n321_2(.douta(w_n321_2[0]),.doutb(w_n321_2[1]),.doutc(w_n321_2[2]),.din(w_n321_0[1]));
	jspl jspl_w_n321_3(.douta(w_n321_3[0]),.doutb(w_n321_3[1]),.din(w_n321_0[2]));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl3 jspl3_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.doutc(w_n327_0[2]),.din(n327));
	jspl3 jspl3_w_n327_1(.douta(w_n327_1[0]),.doutb(w_n327_1[1]),.doutc(w_n327_1[2]),.din(w_n327_0[0]));
	jspl3 jspl3_w_n329_0(.douta(w_n329_0[0]),.doutb(w_n329_0[1]),.doutc(w_n329_0[2]),.din(n329));
	jspl jspl_w_n329_1(.douta(w_n329_1[0]),.doutb(w_n329_1[1]),.din(w_n329_0[0]));
	jspl3 jspl3_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.doutc(w_n330_0[2]),.din(n330));
	jspl3 jspl3_w_n331_0(.douta(w_n331_0[0]),.doutb(w_n331_0[1]),.doutc(w_n331_0[2]),.din(n331));
	jspl3 jspl3_w_n331_1(.douta(w_n331_1[0]),.doutb(w_n331_1[1]),.doutc(w_n331_1[2]),.din(w_n331_0[0]));
	jspl3 jspl3_w_n331_2(.douta(w_n331_2[0]),.doutb(w_n331_2[1]),.doutc(w_n331_2[2]),.din(w_n331_0[1]));
	jspl3 jspl3_w_n332_0(.douta(w_n332_0[0]),.doutb(w_n332_0[1]),.doutc(w_n332_0[2]),.din(n332));
	jspl3 jspl3_w_n332_1(.douta(w_n332_1[0]),.doutb(w_n332_1[1]),.doutc(w_n332_1[2]),.din(w_n332_0[0]));
	jspl3 jspl3_w_n332_2(.douta(w_n332_2[0]),.doutb(w_n332_2[1]),.doutc(w_n332_2[2]),.din(w_n332_0[1]));
	jspl jspl_w_n332_3(.douta(w_n332_3[0]),.doutb(w_n332_3[1]),.din(w_n332_0[2]));
	jspl3 jspl3_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.doutc(w_n333_0[2]),.din(n333));
	jspl3 jspl3_w_n333_1(.douta(w_n333_1[0]),.doutb(w_n333_1[1]),.doutc(w_n333_1[2]),.din(w_n333_0[0]));
	jspl jspl_w_n333_2(.douta(w_n333_2[0]),.doutb(w_n333_2[1]),.din(w_n333_0[1]));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.doutc(w_n336_0[2]),.din(n336));
	jspl3 jspl3_w_n336_1(.douta(w_n336_1[0]),.doutb(w_n336_1[1]),.doutc(w_n336_1[2]),.din(w_n336_0[0]));
	jspl3 jspl3_w_n336_2(.douta(w_n336_2[0]),.doutb(w_n336_2[1]),.doutc(w_n336_2[2]),.din(w_n336_0[1]));
	jspl3 jspl3_w_n337_0(.douta(w_n337_0[0]),.doutb(w_n337_0[1]),.doutc(w_n337_0[2]),.din(n337));
	jspl3 jspl3_w_n337_1(.douta(w_n337_1[0]),.doutb(w_n337_1[1]),.doutc(w_n337_1[2]),.din(w_n337_0[0]));
	jspl3 jspl3_w_n337_2(.douta(w_n337_2[0]),.doutb(w_n337_2[1]),.doutc(w_n337_2[2]),.din(w_n337_0[1]));
	jspl3 jspl3_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.doutc(w_n338_0[2]),.din(n338));
	jspl3 jspl3_w_n339_0(.douta(w_n339_0[0]),.doutb(w_n339_0[1]),.doutc(w_n339_0[2]),.din(n339));
	jspl3 jspl3_w_n339_1(.douta(w_n339_1[0]),.doutb(w_n339_1[1]),.doutc(w_n339_1[2]),.din(w_n339_0[0]));
	jspl3 jspl3_w_n339_2(.douta(w_n339_2[0]),.doutb(w_n339_2[1]),.doutc(w_n339_2[2]),.din(w_n339_0[1]));
	jspl3 jspl3_w_n339_3(.douta(w_n339_3[0]),.doutb(w_n339_3[1]),.doutc(w_n339_3[2]),.din(w_n339_0[2]));
	jspl jspl_w_n339_4(.douta(w_n339_4[0]),.doutb(w_n339_4[1]),.din(w_n339_1[0]));
	jspl3 jspl3_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.doutc(w_n340_0[2]),.din(n340));
	jspl3 jspl3_w_n340_1(.douta(w_n340_1[0]),.doutb(w_n340_1[1]),.doutc(w_n340_1[2]),.din(w_n340_0[0]));
	jspl3 jspl3_w_n344_0(.douta(w_n344_0[0]),.doutb(w_n344_0[1]),.doutc(w_n344_0[2]),.din(n344));
	jspl3 jspl3_w_n344_1(.douta(w_n344_1[0]),.doutb(w_n344_1[1]),.doutc(w_n344_1[2]),.din(w_n344_0[0]));
	jspl3 jspl3_w_n344_2(.douta(w_n344_2[0]),.doutb(w_n344_2[1]),.doutc(w_n344_2[2]),.din(w_n344_0[1]));
	jspl jspl_w_n344_3(.douta(w_n344_3[0]),.doutb(w_n344_3[1]),.din(w_n344_0[2]));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(n345));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl3 jspl3_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.doutc(w_n346_1[2]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n346_2(.douta(w_n346_2[0]),.doutb(w_n346_2[1]),.doutc(w_n346_2[2]),.din(w_n346_0[1]));
	jspl3 jspl3_w_n347_0(.douta(w_n347_0[0]),.doutb(w_n347_0[1]),.doutc(w_n347_0[2]),.din(n347));
	jspl3 jspl3_w_n347_1(.douta(w_n347_1[0]),.doutb(w_n347_1[1]),.doutc(w_n347_1[2]),.din(w_n347_0[0]));
	jspl3 jspl3_w_n347_2(.douta(w_n347_2[0]),.doutb(w_n347_2[1]),.doutc(w_n347_2[2]),.din(w_n347_0[1]));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl3 jspl3_w_n351_0(.douta(w_n351_0[0]),.doutb(w_n351_0[1]),.doutc(w_n351_0[2]),.din(n351));
	jspl jspl_w_n351_1(.douta(w_n351_1[0]),.doutb(w_n351_1[1]),.din(w_n351_0[0]));
	jspl3 jspl3_w_n352_0(.douta(w_n352_0[0]),.doutb(w_n352_0[1]),.doutc(w_n352_0[2]),.din(n352));
	jspl jspl_w_n352_1(.douta(w_n352_1[0]),.doutb(w_n352_1[1]),.din(w_n352_0[0]));
	jspl3 jspl3_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.doutc(w_n353_0[2]),.din(n353));
	jspl3 jspl3_w_n353_1(.douta(w_n353_1[0]),.doutb(w_n353_1[1]),.doutc(w_n353_1[2]),.din(w_n353_0[0]));
	jspl3 jspl3_w_n353_2(.douta(w_n353_2[0]),.doutb(w_n353_2[1]),.doutc(w_n353_2[2]),.din(w_n353_0[1]));
	jspl jspl_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.din(n355));
	jspl3 jspl3_w_n359_0(.douta(w_n359_0[0]),.doutb(w_n359_0[1]),.doutc(w_n359_0[2]),.din(n359));
	jspl3 jspl3_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.doutc(w_n360_0[2]),.din(n360));
	jspl3 jspl3_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.doutc(w_n361_0[2]),.din(n361));
	jspl3 jspl3_w_n361_1(.douta(w_n361_1[0]),.doutb(w_n361_1[1]),.doutc(w_n361_1[2]),.din(w_n361_0[0]));
	jspl3 jspl3_w_n361_2(.douta(w_n361_2[0]),.doutb(w_n361_2[1]),.doutc(w_n361_2[2]),.din(w_n361_0[1]));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n366_2(.douta(w_n366_2[0]),.doutb(w_n366_2[1]),.doutc(w_n366_2[2]),.din(w_n366_0[1]));
	jspl jspl_w_n366_3(.douta(w_n366_3[0]),.doutb(w_n366_3[1]),.din(w_n366_0[2]));
	jspl3 jspl3_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.doutc(w_n370_0[2]),.din(n370));
	jspl3 jspl3_w_n370_1(.douta(w_n370_1[0]),.doutb(w_n370_1[1]),.doutc(w_n370_1[2]),.din(w_n370_0[0]));
	jspl3 jspl3_w_n370_2(.douta(w_n370_2[0]),.doutb(w_n370_2[1]),.doutc(w_n370_2[2]),.din(w_n370_0[1]));
	jspl jspl_w_n370_3(.douta(w_n370_3[0]),.doutb(w_n370_3[1]),.din(w_n370_0[2]));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl3 jspl3_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.doutc(w_n373_0[2]),.din(n373));
	jspl3 jspl3_w_n374_0(.douta(w_n374_0[0]),.doutb(w_n374_0[1]),.doutc(w_n374_0[2]),.din(n374));
	jspl3 jspl3_w_n374_1(.douta(w_n374_1[0]),.doutb(w_n374_1[1]),.doutc(w_n374_1[2]),.din(w_n374_0[0]));
	jspl3 jspl3_w_n374_2(.douta(w_n374_2[0]),.doutb(w_n374_2[1]),.doutc(w_n374_2[2]),.din(w_n374_0[1]));
	jspl jspl_w_n374_3(.douta(w_n374_3[0]),.doutb(w_n374_3[1]),.din(w_n374_0[2]));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_n377_0[2]),.din(n377));
	jspl3 jspl3_w_n377_1(.douta(w_n377_1[0]),.doutb(w_n377_1[1]),.doutc(w_n377_1[2]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n377_2(.douta(w_n377_2[0]),.doutb(w_n377_2[1]),.doutc(w_n377_2[2]),.din(w_n377_0[1]));
	jspl3 jspl3_w_n377_3(.douta(w_n377_3[0]),.doutb(w_n377_3[1]),.doutc(w_n377_3[2]),.din(w_n377_0[2]));
	jspl3 jspl3_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.doutc(w_n378_0[2]),.din(n378));
	jspl3 jspl3_w_n378_1(.douta(w_n378_1[0]),.doutb(w_n378_1[1]),.doutc(w_n378_1[2]),.din(w_n378_0[0]));
	jspl3 jspl3_w_n378_2(.douta(w_n378_2[0]),.doutb(w_n378_2[1]),.doutc(w_n378_2[2]),.din(w_n378_0[1]));
	jspl jspl_w_n378_3(.douta(w_n378_3[0]),.doutb(w_n378_3[1]),.din(w_n378_0[2]));
	jspl jspl_w_n381_0(.douta(w_n381_0[0]),.doutb(w_n381_0[1]),.din(n381));
	jspl3 jspl3_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.doutc(w_n382_0[2]),.din(n382));
	jspl3 jspl3_w_n382_1(.douta(w_n382_1[0]),.doutb(w_n382_1[1]),.doutc(w_n382_1[2]),.din(w_n382_0[0]));
	jspl jspl_w_n382_2(.douta(w_n382_2[0]),.doutb(w_n382_2[1]),.din(w_n382_0[1]));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n383_1(.douta(w_n383_1[0]),.doutb(w_n383_1[1]),.doutc(w_n383_1[2]),.din(w_n383_0[0]));
	jspl3 jspl3_w_n383_2(.douta(w_n383_2[0]),.doutb(w_n383_2[1]),.doutc(w_n383_2[2]),.din(w_n383_0[1]));
	jspl3 jspl3_w_n384_0(.douta(w_n384_0[0]),.doutb(w_n384_0[1]),.doutc(w_n384_0[2]),.din(n384));
	jspl3 jspl3_w_n384_1(.douta(w_n384_1[0]),.doutb(w_n384_1[1]),.doutc(w_n384_1[2]),.din(w_n384_0[0]));
	jspl3 jspl3_w_n384_2(.douta(w_n384_2[0]),.doutb(w_n384_2[1]),.doutc(w_n384_2[2]),.din(w_n384_0[1]));
	jspl jspl_w_n384_3(.douta(w_n384_3[0]),.doutb(w_n384_3[1]),.din(w_n384_0[2]));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl3 jspl3_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.doutc(w_n387_1[2]),.din(w_n387_0[0]));
	jspl3 jspl3_w_n387_2(.douta(w_n387_2[0]),.doutb(w_n387_2[1]),.doutc(w_n387_2[2]),.din(w_n387_0[1]));
	jspl jspl_w_n387_3(.douta(w_n387_3[0]),.doutb(w_n387_3[1]),.din(w_n387_0[2]));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_n388_0[2]),.din(n388));
	jspl jspl_w_n388_1(.douta(w_n388_1[0]),.doutb(w_n388_1[1]),.din(w_n388_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_n389_0[2]),.din(n389));
	jspl3 jspl3_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.doutc(w_n389_1[2]),.din(w_n389_0[0]));
	jspl3 jspl3_w_n389_2(.douta(w_n389_2[0]),.doutb(w_n389_2[1]),.doutc(w_n389_2[2]),.din(w_n389_0[1]));
	jspl3 jspl3_w_n389_3(.douta(w_n389_3[0]),.doutb(w_n389_3[1]),.doutc(w_n389_3[2]),.din(w_n389_0[2]));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl3 jspl3_w_n395_0(.douta(w_n395_0[0]),.doutb(w_n395_0[1]),.doutc(w_n395_0[2]),.din(n395));
	jspl3 jspl3_w_n395_1(.douta(w_n395_1[0]),.doutb(w_n395_1[1]),.doutc(w_n395_1[2]),.din(w_n395_0[0]));
	jspl3 jspl3_w_n395_2(.douta(w_n395_2[0]),.doutb(w_n395_2[1]),.doutc(w_n395_2[2]),.din(w_n395_0[1]));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.din(n396));
	jspl3 jspl3_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.doutc(w_n398_0[2]),.din(n398));
	jspl3 jspl3_w_n399_0(.douta(w_n399_0[0]),.doutb(w_n399_0[1]),.doutc(w_n399_0[2]),.din(n399));
	jspl3 jspl3_w_n400_0(.douta(w_n400_0[0]),.doutb(w_n400_0[1]),.doutc(w_n400_0[2]),.din(n400));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.doutc(w_n401_0[2]),.din(n401));
	jspl jspl_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.din(n402));
	jspl3 jspl3_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.doutc(w_n403_0[2]),.din(n403));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl3 jspl3_w_n404_1(.douta(w_n404_1[0]),.doutb(w_n404_1[1]),.doutc(w_n404_1[2]),.din(w_n404_0[0]));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl3 jspl3_w_n409_0(.douta(w_n409_0[0]),.doutb(w_n409_0[1]),.doutc(w_n409_0[2]),.din(n409));
	jspl3 jspl3_w_n409_1(.douta(w_n409_1[0]),.doutb(w_n409_1[1]),.doutc(w_n409_1[2]),.din(w_n409_0[0]));
	jspl3 jspl3_w_n409_2(.douta(w_n409_2[0]),.doutb(w_n409_2[1]),.doutc(w_n409_2[2]),.din(w_n409_0[1]));
	jspl jspl_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.din(n410));
	jspl3 jspl3_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.doutc(w_n411_0[2]),.din(n411));
	jspl3 jspl3_w_n411_1(.douta(w_n411_1[0]),.doutb(w_n411_1[1]),.doutc(w_n411_1[2]),.din(w_n411_0[0]));
	jspl jspl_w_n411_2(.douta(w_n411_2[0]),.doutb(w_n411_2[1]),.din(w_n411_0[1]));
	jspl jspl_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.din(n413));
	jspl3 jspl3_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.doutc(w_n415_0[2]),.din(n415));
	jspl3 jspl3_w_n415_1(.douta(w_n415_1[0]),.doutb(w_n415_1[1]),.doutc(w_n415_1[2]),.din(w_n415_0[0]));
	jspl3 jspl3_w_n415_2(.douta(w_n415_2[0]),.doutb(w_n415_2[1]),.doutc(w_n415_2[2]),.din(w_n415_0[1]));
	jspl3 jspl3_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.doutc(w_n417_0[2]),.din(n417));
	jspl3 jspl3_w_n418_0(.douta(w_n418_0[0]),.doutb(w_n418_0[1]),.doutc(w_n418_0[2]),.din(n418));
	jspl3 jspl3_w_n418_1(.douta(w_n418_1[0]),.doutb(w_n418_1[1]),.doutc(w_n418_1[2]),.din(w_n418_0[0]));
	jspl jspl_w_n418_2(.douta(w_n418_2[0]),.doutb(w_n418_2[1]),.din(w_n418_0[1]));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.din(n420));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl3 jspl3_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.doutc(w_n426_0[2]),.din(n426));
	jspl3 jspl3_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.doutc(w_n427_0[2]),.din(n427));
	jspl3 jspl3_w_n427_1(.douta(w_n427_1[0]),.doutb(w_n427_1[1]),.doutc(w_n427_1[2]),.din(w_n427_0[0]));
	jspl3 jspl3_w_n427_2(.douta(w_n427_2[0]),.doutb(w_n427_2[1]),.doutc(w_n427_2[2]),.din(w_n427_0[1]));
	jspl3 jspl3_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.doutc(w_n429_0[2]),.din(n429));
	jspl3 jspl3_w_n429_1(.douta(w_n429_1[0]),.doutb(w_n429_1[1]),.doutc(w_n429_1[2]),.din(w_n429_0[0]));
	jspl3 jspl3_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.doutc(w_n430_0[2]),.din(n430));
	jspl jspl_w_n430_1(.douta(w_n430_1[0]),.doutb(w_n430_1[1]),.din(w_n430_0[0]));
	jspl jspl_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.din(n433));
	jspl3 jspl3_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.doutc(w_n434_0[2]),.din(n434));
	jspl3 jspl3_w_n434_1(.douta(w_n434_1[0]),.doutb(w_n434_1[1]),.doutc(w_n434_1[2]),.din(w_n434_0[0]));
	jspl3 jspl3_w_n434_2(.douta(w_n434_2[0]),.doutb(w_n434_2[1]),.doutc(w_n434_2[2]),.din(w_n434_0[1]));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl3 jspl3_w_n435_2(.douta(w_n435_2[0]),.doutb(w_n435_2[1]),.doutc(w_n435_2[2]),.din(w_n435_0[1]));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.doutc(w_n437_0[2]),.din(n437));
	jspl3 jspl3_w_n437_1(.douta(w_n437_1[0]),.doutb(w_n437_1[1]),.doutc(w_n437_1[2]),.din(w_n437_0[0]));
	jspl3 jspl3_w_n438_0(.douta(w_n438_0[0]),.doutb(w_n438_0[1]),.doutc(w_n438_0[2]),.din(n438));
	jspl3 jspl3_w_n438_1(.douta(w_n438_1[0]),.doutb(w_n438_1[1]),.doutc(w_n438_1[2]),.din(w_n438_0[0]));
	jspl jspl_w_n438_2(.douta(w_n438_2[0]),.doutb(w_n438_2[1]),.din(w_n438_0[1]));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.doutc(w_n439_0[2]),.din(n439));
	jspl3 jspl3_w_n439_1(.douta(w_n439_1[0]),.doutb(w_n439_1[1]),.doutc(w_n439_1[2]),.din(w_n439_0[0]));
	jspl3 jspl3_w_n439_2(.douta(w_n439_2[0]),.doutb(w_n439_2[1]),.doutc(w_n439_2[2]),.din(w_n439_0[1]));
	jspl3 jspl3_w_n439_3(.douta(w_n439_3[0]),.doutb(w_n439_3[1]),.doutc(w_n439_3[2]),.din(w_n439_0[2]));
	jspl jspl_w_n439_4(.douta(w_n439_4[0]),.doutb(w_n439_4[1]),.din(w_n439_1[0]));
	jspl3 jspl3_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.doutc(w_n443_0[2]),.din(n443));
	jspl jspl_w_n443_1(.douta(w_n443_1[0]),.doutb(w_n443_1[1]),.din(w_n443_0[0]));
	jspl3 jspl3_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.doutc(w_n445_0[2]),.din(n445));
	jspl3 jspl3_w_n445_1(.douta(w_n445_1[0]),.doutb(w_n445_1[1]),.doutc(w_n445_1[2]),.din(w_n445_0[0]));
	jspl3 jspl3_w_n445_2(.douta(w_n445_2[0]),.doutb(w_n445_2[1]),.doutc(w_n445_2[2]),.din(w_n445_0[1]));
	jspl3 jspl3_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.doutc(w_n446_0[2]),.din(n446));
	jspl3 jspl3_w_n446_1(.douta(w_n446_1[0]),.doutb(w_n446_1[1]),.doutc(w_n446_1[2]),.din(w_n446_0[0]));
	jspl jspl_w_n446_2(.douta(w_n446_2[0]),.doutb(w_n446_2[1]),.din(w_n446_0[1]));
	jspl3 jspl3_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.doutc(w_n447_0[2]),.din(n447));
	jspl3 jspl3_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.doutc(w_n448_0[2]),.din(n448));
	jspl3 jspl3_w_n448_1(.douta(w_n448_1[0]),.doutb(w_n448_1[1]),.doutc(w_n448_1[2]),.din(w_n448_0[0]));
	jspl jspl_w_n448_2(.douta(w_n448_2[0]),.doutb(w_n448_2[1]),.din(w_n448_0[1]));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.din(n455));
	jspl3 jspl3_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.doutc(w_n456_0[2]),.din(n456));
	jspl3 jspl3_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.doutc(w_n457_0[2]),.din(n457));
	jspl3 jspl3_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.doutc(w_n459_0[2]),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n460_2(.douta(w_n460_2[0]),.doutb(w_n460_2[1]),.doutc(w_n460_2[2]),.din(w_n460_0[1]));
	jspl jspl_w_n460_3(.douta(w_n460_3[0]),.doutb(w_n460_3[1]),.din(w_n460_0[2]));
	jspl3 jspl3_w_n461_0(.douta(w_n461_0[0]),.doutb(w_n461_0[1]),.doutc(w_n461_0[2]),.din(n461));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl3 jspl3_w_n462_1(.douta(w_n462_1[0]),.doutb(w_n462_1[1]),.doutc(w_n462_1[2]),.din(w_n462_0[0]));
	jspl jspl_w_n462_2(.douta(w_n462_2[0]),.doutb(w_n462_2[1]),.din(w_n462_0[1]));
	jspl3 jspl3_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.doutc(w_n463_0[2]),.din(n463));
	jspl3 jspl3_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.doutc(w_n467_0[2]),.din(n467));
	jspl3 jspl3_w_n467_1(.douta(w_n467_1[0]),.doutb(w_n467_1[1]),.doutc(w_n467_1[2]),.din(w_n467_0[0]));
	jspl3 jspl3_w_n467_2(.douta(w_n467_2[0]),.doutb(w_n467_2[1]),.doutc(w_n467_2[2]),.din(w_n467_0[1]));
	jspl3 jspl3_w_n468_0(.douta(w_n468_0[0]),.doutb(w_n468_0[1]),.doutc(w_n468_0[2]),.din(n468));
	jspl3 jspl3_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.doutc(w_n470_0[2]),.din(n470));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n480_0(.douta(w_n480_0[0]),.doutb(w_n480_0[1]),.din(n480));
	jspl3 jspl3_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.doutc(w_n481_0[2]),.din(n481));
	jspl jspl_w_n481_1(.douta(w_n481_1[0]),.doutb(w_n481_1[1]),.din(w_n481_0[0]));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(n482));
	jspl3 jspl3_w_n486_0(.douta(w_n486_0[0]),.doutb(w_n486_0[1]),.doutc(w_n486_0[2]),.din(n486));
	jspl3 jspl3_w_n486_1(.douta(w_n486_1[0]),.doutb(w_n486_1[1]),.doutc(w_n486_1[2]),.din(w_n486_0[0]));
	jspl3 jspl3_w_n488_0(.douta(w_n488_0[0]),.doutb(w_n488_0[1]),.doutc(w_n488_0[2]),.din(n488));
	jspl3 jspl3_w_n488_1(.douta(w_n488_1[0]),.doutb(w_n488_1[1]),.doutc(w_n488_1[2]),.din(w_n488_0[0]));
	jspl3 jspl3_w_n488_2(.douta(w_n488_2[0]),.doutb(w_n488_2[1]),.doutc(w_n488_2[2]),.din(w_n488_0[1]));
	jspl jspl_w_n488_3(.douta(w_n488_3[0]),.doutb(w_n488_3[1]),.din(w_n488_0[2]));
	jspl3 jspl3_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.doutc(w_n489_0[2]),.din(n489));
	jspl3 jspl3_w_n489_1(.douta(w_n489_1[0]),.doutb(w_n489_1[1]),.doutc(w_n489_1[2]),.din(w_n489_0[0]));
	jspl3 jspl3_w_n489_2(.douta(w_n489_2[0]),.doutb(w_n489_2[1]),.doutc(w_n489_2[2]),.din(w_n489_0[1]));
	jspl jspl_w_n489_3(.douta(w_n489_3[0]),.doutb(w_n489_3[1]),.din(w_n489_0[2]));
	jspl jspl_w_n491_0(.douta(w_n491_0[0]),.doutb(w_n491_0[1]),.din(n491));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl3 jspl3_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.doutc(w_n495_0[2]),.din(n495));
	jspl jspl_w_n496_0(.douta(w_n496_0[0]),.doutb(w_n496_0[1]),.din(n496));
	jspl3 jspl3_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.doutc(w_n497_0[2]),.din(n497));
	jspl jspl_w_n497_1(.douta(w_n497_1[0]),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl jspl_w_n500_0(.douta(w_n500_0[0]),.doutb(w_n500_0[1]),.din(n500));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl3 jspl3_w_n506_0(.douta(w_n506_0[0]),.doutb(w_n506_0[1]),.doutc(w_n506_0[2]),.din(n506));
	jspl3 jspl3_w_n506_1(.douta(w_n506_1[0]),.doutb(w_n506_1[1]),.doutc(w_n506_1[2]),.din(w_n506_0[0]));
	jspl3 jspl3_w_n506_2(.douta(w_n506_2[0]),.doutb(w_n506_2[1]),.doutc(w_n506_2[2]),.din(w_n506_0[1]));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(n509));
	jspl3 jspl3_w_n510_0(.douta(w_n510_0[0]),.doutb(w_n510_0[1]),.doutc(w_n510_0[2]),.din(n510));
	jspl3 jspl3_w_n510_1(.douta(w_n510_1[0]),.doutb(w_n510_1[1]),.doutc(w_n510_1[2]),.din(w_n510_0[0]));
	jspl3 jspl3_w_n510_2(.douta(w_n510_2[0]),.doutb(w_n510_2[1]),.doutc(w_n510_2[2]),.din(w_n510_0[1]));
	jspl jspl_w_n510_3(.douta(w_n510_3[0]),.doutb(w_n510_3[1]),.din(w_n510_0[2]));
	jspl3 jspl3_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.doutc(w_n513_0[2]),.din(n513));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl3 jspl3_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.doutc(w_n516_0[2]),.din(n516));
	jspl3 jspl3_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.doutc(w_n517_0[2]),.din(n517));
	jspl3 jspl3_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.doutc(w_n519_0[2]),.din(n519));
	jspl3 jspl3_w_n519_1(.douta(w_n519_1[0]),.doutb(w_n519_1[1]),.doutc(w_n519_1[2]),.din(w_n519_0[0]));
	jspl3 jspl3_w_n519_2(.douta(w_n519_2[0]),.doutb(w_n519_2[1]),.doutc(w_n519_2[2]),.din(w_n519_0[1]));
	jspl3 jspl3_w_n519_3(.douta(w_n519_3[0]),.doutb(w_n519_3[1]),.doutc(w_n519_3[2]),.din(w_n519_0[2]));
	jspl3 jspl3_w_n519_4(.douta(w_n519_4[0]),.doutb(w_n519_4[1]),.doutc(w_n519_4[2]),.din(w_n519_1[0]));
	jspl3 jspl3_w_n519_5(.douta(w_n519_5[0]),.doutb(w_n519_5[1]),.doutc(w_n519_5[2]),.din(w_n519_1[1]));
	jspl jspl_w_n521_0(.douta(w_n521_0[0]),.doutb(w_n521_0[1]),.din(n521));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl jspl_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n525_0(.douta(w_n525_0[0]),.doutb(w_n525_0[1]),.din(n525));
	jspl jspl_w_n526_0(.douta(w_n526_0[0]),.doutb(w_n526_0[1]),.din(n526));
	jspl3 jspl3_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.doutc(w_n527_0[2]),.din(n527));
	jspl3 jspl3_w_n527_1(.douta(w_n527_1[0]),.doutb(w_n527_1[1]),.doutc(w_n527_1[2]),.din(w_n527_0[0]));
	jspl3 jspl3_w_n527_2(.douta(w_n527_2[0]),.doutb(w_n527_2[1]),.doutc(w_n527_2[2]),.din(w_n527_0[1]));
	jspl3 jspl3_w_n527_3(.douta(w_n527_3[0]),.doutb(w_n527_3[1]),.doutc(w_n527_3[2]),.din(w_n527_0[2]));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(n530));
	jspl jspl_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.din(n531));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(n532));
	jspl3 jspl3_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.doutc(w_n534_0[2]),.din(n534));
	jspl3 jspl3_w_n534_1(.douta(w_n534_1[0]),.doutb(w_n534_1[1]),.doutc(w_n534_1[2]),.din(w_n534_0[0]));
	jspl3 jspl3_w_n534_2(.douta(w_n534_2[0]),.doutb(w_n534_2[1]),.doutc(w_n534_2[2]),.din(w_n534_0[1]));
	jspl3 jspl3_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.doutc(w_n535_0[2]),.din(n535));
	jspl3 jspl3_w_n535_1(.douta(w_n535_1[0]),.doutb(w_n535_1[1]),.doutc(w_n535_1[2]),.din(w_n535_0[0]));
	jspl jspl_w_n535_2(.douta(w_n535_2[0]),.doutb(w_n535_2[1]),.din(w_n535_0[1]));
	jspl jspl_w_n537_0(.douta(w_n537_0[0]),.doutb(w_n537_0[1]),.din(n537));
	jspl3 jspl3_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.doutc(w_n539_0[2]),.din(n539));
	jspl3 jspl3_w_n539_1(.douta(w_n539_1[0]),.doutb(w_n539_1[1]),.doutc(w_n539_1[2]),.din(w_n539_0[0]));
	jspl3 jspl3_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.doutc(w_n540_0[2]),.din(n540));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(n544));
	jspl3 jspl3_w_n546_0(.douta(w_n546_0[0]),.doutb(w_n546_0[1]),.doutc(w_n546_0[2]),.din(n546));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl3 jspl3_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.doutc(w_n552_0[2]),.din(n552));
	jspl jspl_w_n553_0(.douta(w_n553_0[0]),.doutb(w_n553_0[1]),.din(n553));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_n559_0[1]),.din(n559));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n561_1(.douta(w_n561_1[0]),.doutb(w_n561_1[1]),.din(w_n561_0[0]));
	jspl3 jspl3_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.doutc(w_n562_0[2]),.din(n562));
	jspl jspl_w_n562_1(.douta(w_n562_1[0]),.doutb(w_n562_1[1]),.din(w_n562_0[0]));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(n563));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(n567));
	jspl3 jspl3_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.doutc(w_n568_0[2]),.din(n568));
	jspl3 jspl3_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.doutc(w_n569_0[2]),.din(n569));
	jspl3 jspl3_w_n569_1(.douta(w_n569_1[0]),.doutb(w_n569_1[1]),.doutc(w_n569_1[2]),.din(w_n569_0[0]));
	jspl jspl_w_n569_2(.douta(w_n569_2[0]),.doutb(w_n569_2[1]),.din(w_n569_0[1]));
	jspl3 jspl3_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.doutc(w_n570_0[2]),.din(n570));
	jspl3 jspl3_w_n570_1(.douta(w_n570_1[0]),.doutb(w_n570_1[1]),.doutc(w_n570_1[2]),.din(w_n570_0[0]));
	jspl jspl_w_n570_2(.douta(w_n570_2[0]),.doutb(w_n570_2[1]),.din(w_n570_0[1]));
	jspl jspl_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.din(n572));
	jspl jspl_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.din(n574));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(n577));
	jspl jspl_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.din(n579));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.din(n583));
	jspl3 jspl3_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.doutc(w_n586_0[2]),.din(n586));
	jspl3 jspl3_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.doutc(w_n587_0[2]),.din(n587));
	jspl3 jspl3_w_n587_1(.douta(w_n587_1[0]),.doutb(w_n587_1[1]),.doutc(w_n587_1[2]),.din(w_n587_0[0]));
	jspl3 jspl3_w_n587_2(.douta(w_n587_2[0]),.doutb(w_n587_2[1]),.doutc(w_n587_2[2]),.din(w_n587_0[1]));
	jspl jspl_w_n587_3(.douta(w_n587_3[0]),.doutb(w_n587_3[1]),.din(w_n587_0[2]));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl3 jspl3_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.doutc(w_n594_0[2]),.din(n594));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl jspl_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.din(n599));
	jspl3 jspl3_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.doutc(w_n600_0[2]),.din(n600));
	jspl3 jspl3_w_n600_1(.douta(w_n600_1[0]),.doutb(w_n600_1[1]),.doutc(w_n600_1[2]),.din(w_n600_0[0]));
	jspl3 jspl3_w_n600_2(.douta(w_n600_2[0]),.doutb(w_n600_2[1]),.doutc(w_n600_2[2]),.din(w_n600_0[1]));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.doutc(w_n607_0[2]),.din(n607));
	jspl3 jspl3_w_n607_1(.douta(w_n607_1[0]),.doutb(w_n607_1[1]),.doutc(w_n607_1[2]),.din(w_n607_0[0]));
	jspl jspl_w_n607_2(.douta(w_n607_2[0]),.doutb(w_n607_2[1]),.din(w_n607_0[1]));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.din(n609));
	jspl jspl_w_n610_0(.douta(w_n610_0[0]),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl jspl_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.din(n613));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl3 jspl3_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.doutc(w_n624_0[2]),.din(n624));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.din(n625));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(n628));
	jspl3 jspl3_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.doutc(w_n630_0[2]),.din(n630));
	jspl3 jspl3_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.doutc(w_n634_0[2]),.din(n634));
	jspl jspl_w_n644_0(.douta(w_n644_0[0]),.doutb(w_n644_0[1]),.din(n644));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n646_0(.douta(w_n646_0[0]),.doutb(w_n646_0[1]),.din(n646));
	jspl jspl_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.din(n648));
	jspl3 jspl3_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.doutc(w_n652_0[2]),.din(n652));
	jspl3 jspl3_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.doutc(w_n654_0[2]),.din(n654));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl jspl_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.din(n660));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl jspl_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.din(n663));
	jspl jspl_w_n666_0(.douta(w_n666_0[0]),.doutb(w_n666_0[1]),.din(n666));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(n667));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(n669));
	jspl jspl_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.din(n673));
	jspl3 jspl3_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.doutc(w_n676_0[2]),.din(n676));
	jspl3 jspl3_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.doutc(w_n677_0[2]),.din(n677));
	jspl jspl_w_n677_1(.douta(w_n677_1[0]),.doutb(w_n677_1[1]),.din(w_n677_0[0]));
	jspl3 jspl3_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.doutc(w_n684_0[2]),.din(n684));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(n686));
	jspl3 jspl3_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.doutc(w_n689_0[2]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_n700_0[1]),.din(n700));
	jspl jspl_w_n702_0(.douta(w_n702_0[0]),.doutb(w_n702_0[1]),.din(n702));
	jspl3 jspl3_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.doutc(w_n705_0[2]),.din(n705));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.din(n708));
	jspl3 jspl3_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.doutc(w_n716_0[2]),.din(n716));
	jspl3 jspl3_w_n716_1(.douta(w_n716_1[0]),.doutb(w_n716_1[1]),.doutc(w_n716_1[2]),.din(w_n716_0[0]));
	jspl3 jspl3_w_n716_2(.douta(w_n716_2[0]),.doutb(w_n716_2[1]),.doutc(w_n716_2[2]),.din(w_n716_0[1]));
	jspl3 jspl3_w_n716_3(.douta(w_n716_3[0]),.doutb(w_n716_3[1]),.doutc(w_n716_3[2]),.din(w_n716_0[2]));
	jspl3 jspl3_w_n716_4(.douta(w_n716_4[0]),.doutb(w_n716_4[1]),.doutc(w_n716_4[2]),.din(w_n716_1[0]));
	jspl3 jspl3_w_n716_5(.douta(w_n716_5[0]),.doutb(w_n716_5[1]),.doutc(w_n716_5[2]),.din(w_n716_1[1]));
	jspl3 jspl3_w_n716_6(.douta(w_n716_6[0]),.doutb(w_n716_6[1]),.doutc(w_n716_6[2]),.din(w_n716_1[2]));
	jspl3 jspl3_w_n716_7(.douta(w_n716_7[0]),.doutb(w_n716_7[1]),.doutc(w_n716_7[2]),.din(w_n716_2[0]));
	jspl3 jspl3_w_n716_8(.douta(w_n716_8[0]),.doutb(w_n716_8[1]),.doutc(w_n716_8[2]),.din(w_n716_2[1]));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.doutc(w_n717_0[2]),.din(n717));
	jspl3 jspl3_w_n717_1(.douta(w_n717_1[0]),.doutb(w_n717_1[1]),.doutc(w_n717_1[2]),.din(w_n717_0[0]));
	jspl3 jspl3_w_n717_2(.douta(w_n717_2[0]),.doutb(w_n717_2[1]),.doutc(w_n717_2[2]),.din(w_n717_0[1]));
	jspl jspl_w_n717_3(.douta(w_n717_3[0]),.doutb(w_n717_3[1]),.din(w_n717_0[2]));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl jspl_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.din(n725));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.din(n744));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(n749));
	jspl jspl_w_n751_0(.douta(w_n751_0[0]),.doutb(w_n751_0[1]),.din(n751));
	jspl3 jspl3_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.doutc(w_n752_0[2]),.din(n752));
	jspl jspl_w_n766_0(.douta(w_n766_0[0]),.doutb(w_n766_0[1]),.din(n766));
	jspl3 jspl3_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.doutc(w_n777_0[2]),.din(n777));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(n787));
	jspl jspl_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.din(n788));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(n803));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl jspl_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.din(n814));
	jspl3 jspl3_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.doutc(w_n815_0[2]),.din(n815));
	jspl jspl_w_n815_1(.douta(w_n815_1[0]),.doutb(w_n815_1[1]),.din(w_n815_0[0]));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl3 jspl3_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.doutc(w_n817_0[2]),.din(n817));
	jspl3 jspl3_w_n817_1(.douta(w_n817_1[0]),.doutb(w_n817_1[1]),.doutc(w_n817_1[2]),.din(w_n817_0[0]));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl3 jspl3_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.doutc(w_n825_0[2]),.din(n825));
	jspl3 jspl3_w_n825_1(.douta(w_n825_1[0]),.doutb(w_n825_1[1]),.doutc(w_n825_1[2]),.din(w_n825_0[0]));
	jspl jspl_w_n826_0(.douta(w_n826_0[0]),.doutb(w_n826_0[1]),.din(n826));
	jspl3 jspl3_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.doutc(w_n827_0[2]),.din(n827));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl jspl_w_n841_0(.douta(w_n841_0[0]),.doutb(w_n841_0[1]),.din(n841));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(n842));
	jspl jspl_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.din(n847));
	jspl3 jspl3_w_n849_0(.douta(w_n849_0[0]),.doutb(w_n849_0[1]),.doutc(w_n849_0[2]),.din(n849));
	jspl3 jspl3_w_n850_0(.douta(w_n850_0[0]),.doutb(w_n850_0[1]),.doutc(w_n850_0[2]),.din(n850));
	jspl3 jspl3_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.doutc(w_n852_0[2]),.din(n852));
	jspl jspl_w_n852_1(.douta(w_n852_1[0]),.doutb(w_n852_1[1]),.din(w_n852_0[0]));
	jspl3 jspl3_w_n853_0(.douta(w_n853_0[0]),.doutb(w_n853_0[1]),.doutc(w_n853_0[2]),.din(n853));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl jspl_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.din(n858));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(n862));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.din(n863));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(n866));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl3 jspl3_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.doutc(w_n876_0[2]),.din(n876));
	jspl jspl_w_n876_1(.douta(w_n876_1[0]),.doutb(w_n876_1[1]),.din(w_n876_0[0]));
	jspl3 jspl3_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.doutc(w_n877_0[2]),.din(n877));
	jspl3 jspl3_w_n878_0(.douta(w_n878_0[0]),.doutb(w_n878_0[1]),.doutc(w_n878_0[2]),.din(n878));
	jspl3 jspl3_w_n878_1(.douta(w_n878_1[0]),.doutb(w_n878_1[1]),.doutc(w_n878_1[2]),.din(w_n878_0[0]));
	jspl3 jspl3_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.doutc(w_n880_0[2]),.din(n880));
	jspl3 jspl3_w_n880_1(.douta(w_n880_1[0]),.doutb(w_n880_1[1]),.doutc(w_n880_1[2]),.din(w_n880_0[0]));
	jspl3 jspl3_w_n880_2(.douta(w_n880_2[0]),.doutb(w_n880_2[1]),.doutc(w_n880_2[2]),.din(w_n880_0[1]));
	jspl3 jspl3_w_n880_3(.douta(w_n880_3[0]),.doutb(w_n880_3[1]),.doutc(w_n880_3[2]),.din(w_n880_0[2]));
	jspl3 jspl3_w_n880_4(.douta(w_n880_4[0]),.doutb(w_n880_4[1]),.doutc(w_n880_4[2]),.din(w_n880_1[0]));
	jspl3 jspl3_w_n880_5(.douta(w_n880_5[0]),.doutb(w_n880_5[1]),.doutc(w_n880_5[2]),.din(w_n880_1[1]));
	jspl jspl_w_n880_6(.douta(w_n880_6[0]),.doutb(w_n880_6[1]),.din(w_n880_1[2]));
	jspl3 jspl3_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.doutc(w_n881_0[2]),.din(n881));
	jspl3 jspl3_w_n881_1(.douta(w_n881_1[0]),.doutb(w_n881_1[1]),.doutc(w_n881_1[2]),.din(w_n881_0[0]));
	jspl3 jspl3_w_n881_2(.douta(w_n881_2[0]),.doutb(w_n881_2[1]),.doutc(w_n881_2[2]),.din(w_n881_0[1]));
	jspl3 jspl3_w_n881_3(.douta(w_n881_3[0]),.doutb(w_n881_3[1]),.doutc(w_n881_3[2]),.din(w_n881_0[2]));
	jspl3 jspl3_w_n881_4(.douta(w_n881_4[0]),.doutb(w_n881_4[1]),.doutc(w_n881_4[2]),.din(w_n881_1[0]));
	jspl3 jspl3_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.doutc(w_n884_0[2]),.din(n884));
	jspl jspl_w_n884_1(.douta(w_n884_1[0]),.doutb(w_n884_1[1]),.din(w_n884_0[0]));
	jspl3 jspl3_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.doutc(w_n886_0[2]),.din(n886));
	jspl jspl_w_n886_1(.douta(w_n886_1[0]),.doutb(w_n886_1[1]),.din(w_n886_0[0]));
	jspl3 jspl3_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.doutc(w_n896_0[2]),.din(n896));
	jspl3 jspl3_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.doutc(w_n897_0[2]),.din(n897));
	jspl3 jspl3_w_n897_1(.douta(w_n897_1[0]),.doutb(w_n897_1[1]),.doutc(w_n897_1[2]),.din(w_n897_0[0]));
	jspl jspl_w_n897_2(.douta(w_n897_2[0]),.doutb(w_n897_2[1]),.din(w_n897_0[1]));
	jspl jspl_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.din(n903));
	jspl3 jspl3_w_n904_0(.douta(w_n904_0[0]),.doutb(w_n904_0[1]),.doutc(w_n904_0[2]),.din(n904));
	jspl jspl_w_n904_1(.douta(w_n904_1[0]),.doutb(w_n904_1[1]),.din(w_n904_0[0]));
	jspl3 jspl3_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.doutc(w_n912_0[2]),.din(n912));
	jspl3 jspl3_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.doutc(w_n915_0[2]),.din(n915));
	jspl jspl_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.din(n919));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl3 jspl3_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.doutc(w_n924_0[2]),.din(n924));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_n930_0[2]),.din(n930));
	jspl3 jspl3_w_n930_1(.douta(w_n930_1[0]),.doutb(w_n930_1[1]),.doutc(w_n930_1[2]),.din(w_n930_0[0]));
	jspl jspl_w_n930_2(.douta(w_n930_2[0]),.doutb(w_n930_2[1]),.din(w_n930_0[1]));
	jspl jspl_w_n931_0(.douta(w_n931_0[0]),.doutb(w_n931_0[1]),.din(n931));
	jspl jspl_w_n965_0(.douta(w_n965_0[0]),.doutb(w_n965_0[1]),.din(n965));
	jspl jspl_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.din(n966));
	jspl jspl_w_n968_0(.douta(w_n968_0[0]),.doutb(w_n968_0[1]),.din(n968));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n975_0(.douta(w_n975_0[0]),.doutb(w_n975_0[1]),.din(n975));
	jspl3 jspl3_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.doutc(w_n987_0[2]),.din(n987));
	jspl jspl_w_n987_1(.douta(w_n987_1[0]),.doutb(w_n987_1[1]),.din(w_n987_0[0]));
	jspl3 jspl3_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.doutc(w_n989_0[2]),.din(n989));
	jspl3 jspl3_w_n989_1(.douta(w_n989_1[0]),.doutb(w_n989_1[1]),.doutc(w_n989_1[2]),.din(w_n989_0[0]));
	jspl jspl_w_n989_2(.douta(w_n989_2[0]),.doutb(w_n989_2[1]),.din(w_n989_0[1]));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl3 jspl3_w_n992_1(.douta(w_n992_1[0]),.doutb(w_n992_1[1]),.doutc(w_n992_1[2]),.din(w_n992_0[0]));
	jspl3 jspl3_w_n992_2(.douta(w_n992_2[0]),.doutb(w_n992_2[1]),.doutc(w_n992_2[2]),.din(w_n992_0[1]));
	jspl3 jspl3_w_n992_3(.douta(w_n992_3[0]),.doutb(w_n992_3[1]),.doutc(w_n992_3[2]),.din(w_n992_0[2]));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n994_1(.douta(w_n994_1[0]),.doutb(w_n994_1[1]),.doutc(w_n994_1[2]),.din(w_n994_0[0]));
	jspl3 jspl3_w_n994_2(.douta(w_n994_2[0]),.doutb(w_n994_2[1]),.doutc(w_n994_2[2]),.din(w_n994_0[1]));
	jspl3 jspl3_w_n994_3(.douta(w_n994_3[0]),.doutb(w_n994_3[1]),.doutc(w_n994_3[2]),.din(w_n994_0[2]));
	jspl3 jspl3_w_n994_4(.douta(w_n994_4[0]),.doutb(w_n994_4[1]),.doutc(w_n994_4[2]),.din(w_n994_1[0]));
	jspl3 jspl3_w_n994_5(.douta(w_n994_5[0]),.doutb(w_n994_5[1]),.doutc(w_n994_5[2]),.din(w_n994_1[1]));
	jspl jspl_w_n994_6(.douta(w_n994_6[0]),.doutb(w_n994_6[1]),.din(w_n994_1[2]));
	jspl3 jspl3_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.doutc(w_n996_0[2]),.din(n996));
	jspl3 jspl3_w_n996_1(.douta(w_n996_1[0]),.doutb(w_n996_1[1]),.doutc(w_n996_1[2]),.din(w_n996_0[0]));
	jspl3 jspl3_w_n996_2(.douta(w_n996_2[0]),.doutb(w_n996_2[1]),.doutc(w_n996_2[2]),.din(w_n996_0[1]));
	jspl3 jspl3_w_n996_3(.douta(w_n996_3[0]),.doutb(w_n996_3[1]),.doutc(w_n996_3[2]),.din(w_n996_0[2]));
	jspl3 jspl3_w_n996_4(.douta(w_n996_4[0]),.doutb(w_n996_4[1]),.doutc(w_n996_4[2]),.din(w_n996_1[0]));
	jspl3 jspl3_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.doutc(w_n997_0[2]),.din(n997));
	jspl3 jspl3_w_n997_1(.douta(w_n997_1[0]),.doutb(w_n997_1[1]),.doutc(w_n997_1[2]),.din(w_n997_0[0]));
	jspl3 jspl3_w_n997_2(.douta(w_n997_2[0]),.doutb(w_n997_2[1]),.doutc(w_n997_2[2]),.din(w_n997_0[1]));
	jspl3 jspl3_w_n997_3(.douta(w_n997_3[0]),.doutb(w_n997_3[1]),.doutc(w_n997_3[2]),.din(w_n997_0[2]));
	jspl jspl_w_n997_4(.douta(w_n997_4[0]),.doutb(w_n997_4[1]),.din(w_n997_1[0]));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl jspl_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.din(n1002));
	jspl3 jspl3_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.doutc(w_n1005_0[2]),.din(n1005));
	jspl3 jspl3_w_n1005_1(.douta(w_n1005_1[0]),.doutb(w_n1005_1[1]),.doutc(w_n1005_1[2]),.din(w_n1005_0[0]));
	jspl3 jspl3_w_n1005_2(.douta(w_n1005_2[0]),.doutb(w_n1005_2[1]),.doutc(w_n1005_2[2]),.din(w_n1005_0[1]));
	jspl3 jspl3_w_n1005_3(.douta(w_n1005_3[0]),.doutb(w_n1005_3[1]),.doutc(w_n1005_3[2]),.din(w_n1005_0[2]));
	jspl jspl_w_n1005_4(.douta(w_n1005_4[0]),.doutb(w_n1005_4[1]),.din(w_n1005_1[0]));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.din(n1006));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.din(n1012));
	jspl3 jspl3_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.doutc(w_n1016_0[2]),.din(n1016));
	jspl jspl_w_n1016_1(.douta(w_n1016_1[0]),.doutb(w_n1016_1[1]),.din(w_n1016_0[0]));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.din(n1019));
	jspl jspl_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.din(n1021));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(n1023));
	jspl3 jspl3_w_n1024_0(.douta(w_n1024_0[0]),.doutb(w_n1024_0[1]),.doutc(w_n1024_0[2]),.din(n1024));
	jspl3 jspl3_w_n1025_0(.douta(w_n1025_0[0]),.doutb(w_n1025_0[1]),.doutc(w_n1025_0[2]),.din(n1025));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.din(n1030));
	jspl jspl_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.din(n1032));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl3 jspl3_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.doutc(w_n1035_0[2]),.din(n1035));
	jspl3 jspl3_w_n1035_1(.douta(w_n1035_1[0]),.doutb(w_n1035_1[1]),.doutc(w_n1035_1[2]),.din(w_n1035_0[0]));
	jspl3 jspl3_w_n1035_2(.douta(w_n1035_2[0]),.doutb(w_n1035_2[1]),.doutc(w_n1035_2[2]),.din(w_n1035_0[1]));
	jspl3 jspl3_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.doutc(w_n1039_0[2]),.din(n1039));
	jspl jspl_w_n1040_0(.douta(w_n1040_0[0]),.doutb(w_n1040_0[1]),.din(n1040));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(n1043));
	jspl jspl_w_n1045_0(.douta(w_n1045_0[0]),.doutb(w_n1045_0[1]),.din(n1045));
	jspl jspl_w_n1050_0(.douta(w_n1050_0[0]),.doutb(w_n1050_0[1]),.din(n1050));
	jspl jspl_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.din(n1053));
	jspl3 jspl3_w_n1055_0(.douta(w_n1055_0[0]),.doutb(w_n1055_0[1]),.doutc(w_n1055_0[2]),.din(n1055));
	jspl3 jspl3_w_n1055_1(.douta(w_n1055_1[0]),.doutb(w_n1055_1[1]),.doutc(w_n1055_1[2]),.din(w_n1055_0[0]));
	jspl jspl_w_n1055_2(.douta(w_n1055_2[0]),.doutb(w_n1055_2[1]),.din(w_n1055_0[1]));
	jspl jspl_w_n1056_0(.douta(w_n1056_0[0]),.doutb(w_n1056_0[1]),.din(n1056));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.din(n1057));
	jspl jspl_w_n1060_0(.douta(w_n1060_0[0]),.doutb(w_n1060_0[1]),.din(n1060));
	jspl3 jspl3_w_n1064_0(.douta(w_n1064_0[0]),.doutb(w_n1064_0[1]),.doutc(w_n1064_0[2]),.din(n1064));
	jspl jspl_w_n1064_1(.douta(w_n1064_1[0]),.doutb(w_n1064_1[1]),.din(w_n1064_0[0]));
	jspl jspl_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.din(n1066));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(n1069));
	jspl jspl_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.din(n1071));
	jspl3 jspl3_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.doutc(w_n1072_0[2]),.din(n1072));
	jspl jspl_w_n1072_1(.douta(w_n1072_1[0]),.doutb(w_n1072_1[1]),.din(w_n1072_0[0]));
	jspl3 jspl3_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.doutc(w_n1073_0[2]),.din(n1073));
	jspl jspl_w_n1073_1(.douta(w_n1073_1[0]),.doutb(w_n1073_1[1]),.din(w_n1073_0[0]));
	jspl3 jspl3_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.doutc(w_n1074_0[2]),.din(n1074));
	jspl3 jspl3_w_n1074_1(.douta(w_n1074_1[0]),.doutb(w_n1074_1[1]),.doutc(w_n1074_1[2]),.din(w_n1074_0[0]));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(n1078));
	jspl jspl_w_n1079_0(.douta(w_n1079_0[0]),.doutb(w_n1079_0[1]),.din(n1079));
	jspl jspl_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.din(n1080));
	jspl jspl_w_n1085_0(.douta(w_n1085_0[0]),.doutb(w_n1085_0[1]),.din(n1085));
	jspl3 jspl3_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.doutc(w_n1087_0[2]),.din(n1087));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl jspl_w_n1093_0(.douta(w_n1093_0[0]),.doutb(w_n1093_0[1]),.din(n1093));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(n1094));
	jspl3 jspl3_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.doutc(w_n1095_0[2]),.din(n1095));
	jspl3 jspl3_w_n1095_1(.douta(w_n1095_1[0]),.doutb(w_n1095_1[1]),.doutc(w_n1095_1[2]),.din(w_n1095_0[0]));
	jspl3 jspl3_w_n1095_2(.douta(w_n1095_2[0]),.doutb(w_n1095_2[1]),.doutc(w_n1095_2[2]),.din(w_n1095_0[1]));
	jspl3 jspl3_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.doutc(w_n1096_0[2]),.din(n1096));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1104_0(.douta(w_n1104_0[0]),.doutb(w_n1104_0[1]),.din(n1104));
	jspl3 jspl3_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.doutc(w_n1105_0[2]),.din(n1105));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl3 jspl3_w_n1110_0(.douta(w_n1110_0[0]),.doutb(w_n1110_0[1]),.doutc(w_n1110_0[2]),.din(n1110));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl3 jspl3_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.doutc(w_n1115_0[2]),.din(n1115));
	jspl jspl_w_n1115_1(.douta(w_n1115_1[0]),.doutb(w_n1115_1[1]),.din(w_n1115_0[0]));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl jspl_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.din(n1122));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl3 jspl3_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.doutc(w_n1127_0[2]),.din(n1127));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.din(n1133));
	jspl3 jspl3_w_n1135_0(.douta(w_n1135_0[0]),.doutb(w_n1135_0[1]),.doutc(w_n1135_0[2]),.din(n1135));
	jspl jspl_w_n1135_1(.douta(w_n1135_1[0]),.doutb(w_n1135_1[1]),.din(w_n1135_0[0]));
	jspl jspl_w_n1140_0(.douta(w_n1140_0[0]),.doutb(w_n1140_0[1]),.din(n1140));
	jspl jspl_w_n1147_0(.douta(w_n1147_0[0]),.doutb(w_n1147_0[1]),.din(n1147));
	jspl3 jspl3_w_n1149_0(.douta(w_n1149_0[0]),.doutb(w_n1149_0[1]),.doutc(w_n1149_0[2]),.din(n1149));
	jspl3 jspl3_w_n1149_1(.douta(w_n1149_1[0]),.doutb(w_n1149_1[1]),.doutc(w_n1149_1[2]),.din(w_n1149_0[0]));
	jspl jspl_w_n1150_0(.douta(w_n1150_0[0]),.doutb(w_n1150_0[1]),.din(n1150));
	jspl3 jspl3_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.doutc(w_n1151_0[2]),.din(n1151));
	jspl3 jspl3_w_n1151_1(.douta(w_n1151_1[0]),.doutb(w_n1151_1[1]),.doutc(w_n1151_1[2]),.din(w_n1151_0[0]));
	jspl3 jspl3_w_n1152_0(.douta(w_n1152_0[0]),.doutb(w_n1152_0[1]),.doutc(w_n1152_0[2]),.din(n1152));
	jspl3 jspl3_w_n1152_1(.douta(w_n1152_1[0]),.doutb(w_n1152_1[1]),.doutc(w_n1152_1[2]),.din(w_n1152_0[0]));
	jspl jspl_w_n1152_2(.douta(w_n1152_2[0]),.doutb(w_n1152_2[1]),.din(w_n1152_0[1]));
	jspl3 jspl3_w_n1154_0(.douta(w_n1154_0[0]),.doutb(w_n1154_0[1]),.doutc(w_n1154_0[2]),.din(n1154));
	jspl3 jspl3_w_n1154_1(.douta(w_n1154_1[0]),.doutb(w_n1154_1[1]),.doutc(w_n1154_1[2]),.din(w_n1154_0[0]));
	jspl3 jspl3_w_n1154_2(.douta(w_n1154_2[0]),.doutb(w_n1154_2[1]),.doutc(w_n1154_2[2]),.din(w_n1154_0[1]));
	jspl3 jspl3_w_n1154_3(.douta(w_n1154_3[0]),.doutb(w_n1154_3[1]),.doutc(w_n1154_3[2]),.din(w_n1154_0[2]));
	jspl3 jspl3_w_n1154_4(.douta(w_n1154_4[0]),.doutb(w_n1154_4[1]),.doutc(w_n1154_4[2]),.din(w_n1154_1[0]));
	jspl3 jspl3_w_n1154_5(.douta(w_n1154_5[0]),.doutb(w_n1154_5[1]),.doutc(w_n1154_5[2]),.din(w_n1154_1[1]));
	jspl3 jspl3_w_n1154_6(.douta(w_n1154_6[0]),.doutb(w_n1154_6[1]),.doutc(w_n1154_6[2]),.din(w_n1154_1[2]));
	jspl3 jspl3_w_n1154_7(.douta(w_n1154_7[0]),.doutb(w_n1154_7[1]),.doutc(w_n1154_7[2]),.din(w_n1154_2[0]));
	jspl3 jspl3_w_n1154_8(.douta(w_n1154_8[0]),.doutb(w_n1154_8[1]),.doutc(w_n1154_8[2]),.din(w_n1154_2[1]));
	jspl3 jspl3_w_n1154_9(.douta(w_n1154_9[0]),.doutb(w_n1154_9[1]),.doutc(w_n1154_9[2]),.din(w_n1154_2[2]));
	jspl3 jspl3_w_n1154_10(.douta(w_n1154_10[0]),.doutb(w_n1154_10[1]),.doutc(w_n1154_10[2]),.din(w_n1154_3[0]));
	jspl3 jspl3_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.doutc(w_n1156_0[2]),.din(n1156));
	jspl3 jspl3_w_n1156_1(.douta(w_n1156_1[0]),.doutb(w_n1156_1[1]),.doutc(w_n1156_1[2]),.din(w_n1156_0[0]));
	jspl3 jspl3_w_n1156_2(.douta(w_n1156_2[0]),.doutb(w_n1156_2[1]),.doutc(w_n1156_2[2]),.din(w_n1156_0[1]));
	jspl3 jspl3_w_n1156_3(.douta(w_n1156_3[0]),.doutb(w_n1156_3[1]),.doutc(w_n1156_3[2]),.din(w_n1156_0[2]));
	jspl3 jspl3_w_n1156_4(.douta(w_n1156_4[0]),.doutb(w_n1156_4[1]),.doutc(w_n1156_4[2]),.din(w_n1156_1[0]));
	jspl3 jspl3_w_n1156_5(.douta(w_n1156_5[0]),.doutb(w_n1156_5[1]),.doutc(w_n1156_5[2]),.din(w_n1156_1[1]));
	jspl3 jspl3_w_n1156_6(.douta(w_n1156_6[0]),.doutb(w_n1156_6[1]),.doutc(w_n1156_6[2]),.din(w_n1156_1[2]));
	jspl3 jspl3_w_n1156_7(.douta(w_n1156_7[0]),.doutb(w_n1156_7[1]),.doutc(w_n1156_7[2]),.din(w_n1156_2[0]));
	jspl3 jspl3_w_n1156_8(.douta(w_n1156_8[0]),.doutb(w_n1156_8[1]),.doutc(w_n1156_8[2]),.din(w_n1156_2[1]));
	jspl3 jspl3_w_n1156_9(.douta(w_n1156_9[0]),.doutb(w_n1156_9[1]),.doutc(w_n1156_9[2]),.din(w_n1156_2[2]));
	jspl3 jspl3_w_n1156_10(.douta(w_n1156_10[0]),.doutb(w_n1156_10[1]),.doutc(w_n1156_10[2]),.din(w_n1156_3[0]));
	jspl3 jspl3_w_n1156_11(.douta(w_n1156_11[0]),.doutb(w_n1156_11[1]),.doutc(w_n1156_11[2]),.din(w_n1156_3[1]));
	jspl jspl_w_n1156_12(.douta(w_n1156_12[0]),.doutb(w_n1156_12[1]),.din(w_n1156_3[2]));
	jspl jspl_w_n1158_0(.douta(w_n1158_0[0]),.doutb(w_n1158_0[1]),.din(n1158));
	jspl3 jspl3_w_n1160_0(.douta(w_n1160_0[0]),.doutb(w_n1160_0[1]),.doutc(w_n1160_0[2]),.din(n1160));
	jspl3 jspl3_w_n1160_1(.douta(w_n1160_1[0]),.doutb(w_n1160_1[1]),.doutc(w_n1160_1[2]),.din(w_n1160_0[0]));
	jspl jspl_w_n1160_2(.douta(w_n1160_2[0]),.doutb(w_n1160_2[1]),.din(w_n1160_0[1]));
	jspl3 jspl3_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.doutc(w_n1163_0[2]),.din(n1163));
	jspl3 jspl3_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.doutc(w_n1164_0[2]),.din(n1164));
	jspl3 jspl3_w_n1164_1(.douta(w_n1164_1[0]),.doutb(w_n1164_1[1]),.doutc(w_n1164_1[2]),.din(w_n1164_0[0]));
	jspl3 jspl3_w_n1164_2(.douta(w_n1164_2[0]),.doutb(w_n1164_2[1]),.doutc(w_n1164_2[2]),.din(w_n1164_0[1]));
	jspl3 jspl3_w_n1164_3(.douta(w_n1164_3[0]),.doutb(w_n1164_3[1]),.doutc(w_n1164_3[2]),.din(w_n1164_0[2]));
	jspl3 jspl3_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.doutc(w_n1166_0[2]),.din(n1166));
	jspl3 jspl3_w_n1166_1(.douta(w_n1166_1[0]),.doutb(w_n1166_1[1]),.doutc(w_n1166_1[2]),.din(w_n1166_0[0]));
	jspl3 jspl3_w_n1166_2(.douta(w_n1166_2[0]),.doutb(w_n1166_2[1]),.doutc(w_n1166_2[2]),.din(w_n1166_0[1]));
	jspl3 jspl3_w_n1166_3(.douta(w_n1166_3[0]),.doutb(w_n1166_3[1]),.doutc(w_n1166_3[2]),.din(w_n1166_0[2]));
	jspl3 jspl3_w_n1166_4(.douta(w_n1166_4[0]),.doutb(w_n1166_4[1]),.doutc(w_n1166_4[2]),.din(w_n1166_1[0]));
	jspl3 jspl3_w_n1166_5(.douta(w_n1166_5[0]),.doutb(w_n1166_5[1]),.doutc(w_n1166_5[2]),.din(w_n1166_1[1]));
	jspl jspl_w_n1166_6(.douta(w_n1166_6[0]),.doutb(w_n1166_6[1]),.din(w_n1166_1[2]));
	jspl3 jspl3_w_n1168_0(.douta(w_n1168_0[0]),.doutb(w_n1168_0[1]),.doutc(w_n1168_0[2]),.din(n1168));
	jspl3 jspl3_w_n1168_1(.douta(w_n1168_1[0]),.doutb(w_n1168_1[1]),.doutc(w_n1168_1[2]),.din(w_n1168_0[0]));
	jspl3 jspl3_w_n1168_2(.douta(w_n1168_2[0]),.doutb(w_n1168_2[1]),.doutc(w_n1168_2[2]),.din(w_n1168_0[1]));
	jspl3 jspl3_w_n1168_3(.douta(w_n1168_3[0]),.doutb(w_n1168_3[1]),.doutc(w_n1168_3[2]),.din(w_n1168_0[2]));
	jspl3 jspl3_w_n1168_4(.douta(w_n1168_4[0]),.doutb(w_n1168_4[1]),.doutc(w_n1168_4[2]),.din(w_n1168_1[0]));
	jspl3 jspl3_w_n1170_0(.douta(w_n1170_0[0]),.doutb(w_n1170_0[1]),.doutc(w_n1170_0[2]),.din(n1170));
	jspl3 jspl3_w_n1170_1(.douta(w_n1170_1[0]),.doutb(w_n1170_1[1]),.doutc(w_n1170_1[2]),.din(w_n1170_0[0]));
	jspl3 jspl3_w_n1170_2(.douta(w_n1170_2[0]),.doutb(w_n1170_2[1]),.doutc(w_n1170_2[2]),.din(w_n1170_0[1]));
	jspl3 jspl3_w_n1170_3(.douta(w_n1170_3[0]),.doutb(w_n1170_3[1]),.doutc(w_n1170_3[2]),.din(w_n1170_0[2]));
	jspl jspl_w_n1170_4(.douta(w_n1170_4[0]),.doutb(w_n1170_4[1]),.din(w_n1170_1[0]));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(n1173));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(n1176));
	jspl3 jspl3_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.doutc(w_n1178_0[2]),.din(n1178));
	jspl jspl_w_n1180_0(.douta(w_n1180_0[0]),.doutb(w_n1180_0[1]),.din(n1180));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(n1186));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(n1188));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1192_0(.douta(w_n1192_0[0]),.doutb(w_n1192_0[1]),.din(n1192));
	jspl3 jspl3_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.doutc(w_n1196_0[2]),.din(n1196));
	jspl jspl_w_n1196_1(.douta(w_n1196_1[0]),.doutb(w_n1196_1[1]),.din(w_n1196_0[0]));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.din(n1215));
	jspl jspl_w_n1226_0(.douta(w_n1226_0[0]),.doutb(w_n1226_0[1]),.din(n1226));
	jspl3 jspl3_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.doutc(w_n1232_0[2]),.din(n1232));
	jspl jspl_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.din(n1235));
	jspl jspl_w_n1243_0(.douta(w_n1243_0[0]),.doutb(w_n1243_0[1]),.din(n1243));
	jspl jspl_w_n1249_0(.douta(w_n1249_0[0]),.doutb(w_n1249_0[1]),.din(n1249));
	jspl jspl_w_n1250_0(.douta(w_n1250_0[0]),.doutb(w_n1250_0[1]),.din(n1250));
	jspl3 jspl3_w_n1252_0(.douta(w_n1252_0[0]),.doutb(w_n1252_0[1]),.doutc(w_n1252_0[2]),.din(n1252));
	jspl jspl_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.din(n1253));
	jspl3 jspl3_w_n1254_0(.douta(w_n1254_0[0]),.doutb(w_n1254_0[1]),.doutc(w_n1254_0[2]),.din(n1254));
	jspl3 jspl3_w_n1254_1(.douta(w_n1254_1[0]),.doutb(w_n1254_1[1]),.doutc(w_n1254_1[2]),.din(w_n1254_0[0]));
	jspl jspl_w_n1254_2(.douta(w_n1254_2[0]),.doutb(w_n1254_2[1]),.din(w_n1254_0[1]));
	jspl3 jspl3_w_n1255_0(.douta(w_n1255_0[0]),.doutb(w_n1255_0[1]),.doutc(w_n1255_0[2]),.din(n1255));
	jspl3 jspl3_w_n1255_1(.douta(w_n1255_1[0]),.doutb(w_n1255_1[1]),.doutc(w_n1255_1[2]),.din(w_n1255_0[0]));
	jspl jspl_w_n1255_2(.douta(w_n1255_2[0]),.doutb(w_n1255_2[1]),.din(w_n1255_0[1]));
	jspl3 jspl3_w_n1257_0(.douta(w_n1257_0[0]),.doutb(w_n1257_0[1]),.doutc(w_n1257_0[2]),.din(n1257));
	jspl3 jspl3_w_n1257_1(.douta(w_n1257_1[0]),.doutb(w_n1257_1[1]),.doutc(w_n1257_1[2]),.din(w_n1257_0[0]));
	jspl3 jspl3_w_n1257_2(.douta(w_n1257_2[0]),.doutb(w_n1257_2[1]),.doutc(w_n1257_2[2]),.din(w_n1257_0[1]));
	jspl3 jspl3_w_n1257_3(.douta(w_n1257_3[0]),.doutb(w_n1257_3[1]),.doutc(w_n1257_3[2]),.din(w_n1257_0[2]));
	jspl3 jspl3_w_n1257_4(.douta(w_n1257_4[0]),.doutb(w_n1257_4[1]),.doutc(w_n1257_4[2]),.din(w_n1257_1[0]));
	jspl3 jspl3_w_n1257_5(.douta(w_n1257_5[0]),.doutb(w_n1257_5[1]),.doutc(w_n1257_5[2]),.din(w_n1257_1[1]));
	jspl3 jspl3_w_n1257_6(.douta(w_n1257_6[0]),.doutb(w_n1257_6[1]),.doutc(w_n1257_6[2]),.din(w_n1257_1[2]));
	jspl3 jspl3_w_n1257_7(.douta(w_n1257_7[0]),.doutb(w_n1257_7[1]),.doutc(w_n1257_7[2]),.din(w_n1257_2[0]));
	jspl3 jspl3_w_n1257_8(.douta(w_n1257_8[0]),.doutb(w_n1257_8[1]),.doutc(w_n1257_8[2]),.din(w_n1257_2[1]));
	jspl3 jspl3_w_n1257_9(.douta(w_n1257_9[0]),.doutb(w_n1257_9[1]),.doutc(w_n1257_9[2]),.din(w_n1257_2[2]));
	jspl3 jspl3_w_n1257_10(.douta(w_n1257_10[0]),.doutb(w_n1257_10[1]),.doutc(w_n1257_10[2]),.din(w_n1257_3[0]));
	jspl3 jspl3_w_n1257_11(.douta(w_n1257_11[0]),.doutb(w_n1257_11[1]),.doutc(w_n1257_11[2]),.din(w_n1257_3[1]));
	jspl3 jspl3_w_n1257_12(.douta(w_n1257_12[0]),.doutb(w_n1257_12[1]),.doutc(w_n1257_12[2]),.din(w_n1257_3[2]));
	jspl3 jspl3_w_n1257_13(.douta(w_n1257_13[0]),.doutb(w_n1257_13[1]),.doutc(w_n1257_13[2]),.din(w_n1257_4[0]));
	jspl3 jspl3_w_n1259_0(.douta(w_n1259_0[0]),.doutb(w_n1259_0[1]),.doutc(w_n1259_0[2]),.din(n1259));
	jspl3 jspl3_w_n1259_1(.douta(w_n1259_1[0]),.doutb(w_n1259_1[1]),.doutc(w_n1259_1[2]),.din(w_n1259_0[0]));
	jspl3 jspl3_w_n1259_2(.douta(w_n1259_2[0]),.doutb(w_n1259_2[1]),.doutc(w_n1259_2[2]),.din(w_n1259_0[1]));
	jspl3 jspl3_w_n1259_3(.douta(w_n1259_3[0]),.doutb(w_n1259_3[1]),.doutc(w_n1259_3[2]),.din(w_n1259_0[2]));
	jspl3 jspl3_w_n1259_4(.douta(w_n1259_4[0]),.doutb(w_n1259_4[1]),.doutc(w_n1259_4[2]),.din(w_n1259_1[0]));
	jspl3 jspl3_w_n1259_5(.douta(w_n1259_5[0]),.doutb(w_n1259_5[1]),.doutc(w_n1259_5[2]),.din(w_n1259_1[1]));
	jspl3 jspl3_w_n1259_6(.douta(w_n1259_6[0]),.doutb(w_n1259_6[1]),.doutc(w_n1259_6[2]),.din(w_n1259_1[2]));
	jspl3 jspl3_w_n1259_7(.douta(w_n1259_7[0]),.doutb(w_n1259_7[1]),.doutc(w_n1259_7[2]),.din(w_n1259_2[0]));
	jspl3 jspl3_w_n1259_8(.douta(w_n1259_8[0]),.doutb(w_n1259_8[1]),.doutc(w_n1259_8[2]),.din(w_n1259_2[1]));
	jspl jspl_w_n1259_9(.douta(w_n1259_9[0]),.doutb(w_n1259_9[1]),.din(w_n1259_2[2]));
	jspl3 jspl3_w_n1260_0(.douta(w_n1260_0[0]),.doutb(w_n1260_0[1]),.doutc(w_n1260_0[2]),.din(n1260));
	jspl3 jspl3_w_n1261_0(.douta(w_n1261_0[0]),.doutb(w_n1261_0[1]),.doutc(w_n1261_0[2]),.din(n1261));
	jspl3 jspl3_w_n1261_1(.douta(w_n1261_1[0]),.doutb(w_n1261_1[1]),.doutc(w_n1261_1[2]),.din(w_n1261_0[0]));
	jspl3 jspl3_w_n1261_2(.douta(w_n1261_2[0]),.doutb(w_n1261_2[1]),.doutc(w_n1261_2[2]),.din(w_n1261_0[1]));
	jspl3 jspl3_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.doutc(w_n1266_0[2]),.din(n1266));
	jspl3 jspl3_w_n1266_1(.douta(w_n1266_1[0]),.doutb(w_n1266_1[1]),.doutc(w_n1266_1[2]),.din(w_n1266_0[0]));
	jspl3 jspl3_w_n1266_2(.douta(w_n1266_2[0]),.doutb(w_n1266_2[1]),.doutc(w_n1266_2[2]),.din(w_n1266_0[1]));
	jspl3 jspl3_w_n1266_3(.douta(w_n1266_3[0]),.doutb(w_n1266_3[1]),.doutc(w_n1266_3[2]),.din(w_n1266_0[2]));
	jspl3 jspl3_w_n1266_4(.douta(w_n1266_4[0]),.doutb(w_n1266_4[1]),.doutc(w_n1266_4[2]),.din(w_n1266_1[0]));
	jspl3 jspl3_w_n1266_5(.douta(w_n1266_5[0]),.doutb(w_n1266_5[1]),.doutc(w_n1266_5[2]),.din(w_n1266_1[1]));
	jspl jspl_w_n1266_6(.douta(w_n1266_6[0]),.doutb(w_n1266_6[1]),.din(w_n1266_1[2]));
	jspl jspl_w_n1268_0(.douta(w_n1268_0[0]),.doutb(w_n1268_0[1]),.din(n1268));
	jspl3 jspl3_w_n1270_0(.douta(w_n1270_0[0]),.doutb(w_n1270_0[1]),.doutc(w_n1270_0[2]),.din(n1270));
	jspl3 jspl3_w_n1270_1(.douta(w_n1270_1[0]),.doutb(w_n1270_1[1]),.doutc(w_n1270_1[2]),.din(w_n1270_0[0]));
	jspl3 jspl3_w_n1270_2(.douta(w_n1270_2[0]),.doutb(w_n1270_2[1]),.doutc(w_n1270_2[2]),.din(w_n1270_0[1]));
	jspl3 jspl3_w_n1270_3(.douta(w_n1270_3[0]),.doutb(w_n1270_3[1]),.doutc(w_n1270_3[2]),.din(w_n1270_0[2]));
	jspl3 jspl3_w_n1272_0(.douta(w_n1272_0[0]),.doutb(w_n1272_0[1]),.doutc(w_n1272_0[2]),.din(n1272));
	jspl3 jspl3_w_n1272_1(.douta(w_n1272_1[0]),.doutb(w_n1272_1[1]),.doutc(w_n1272_1[2]),.din(w_n1272_0[0]));
	jspl3 jspl3_w_n1272_2(.douta(w_n1272_2[0]),.doutb(w_n1272_2[1]),.doutc(w_n1272_2[2]),.din(w_n1272_0[1]));
	jspl3 jspl3_w_n1272_3(.douta(w_n1272_3[0]),.doutb(w_n1272_3[1]),.doutc(w_n1272_3[2]),.din(w_n1272_0[2]));
	jspl3 jspl3_w_n1272_4(.douta(w_n1272_4[0]),.doutb(w_n1272_4[1]),.doutc(w_n1272_4[2]),.din(w_n1272_1[0]));
	jspl3 jspl3_w_n1294_0(.douta(w_n1294_0[0]),.doutb(w_n1294_0[1]),.doutc(w_n1294_0[2]),.din(n1294));
	jspl3 jspl3_w_n1295_0(.douta(w_n1295_0[0]),.doutb(w_n1295_0[1]),.doutc(w_n1295_0[2]),.din(n1295));
	jspl3 jspl3_w_n1295_1(.douta(w_n1295_1[0]),.doutb(w_n1295_1[1]),.doutc(w_n1295_1[2]),.din(w_n1295_0[0]));
	jspl3 jspl3_w_n1295_2(.douta(w_n1295_2[0]),.doutb(w_n1295_2[1]),.doutc(w_n1295_2[2]),.din(w_n1295_0[1]));
	jspl3 jspl3_w_n1295_3(.douta(w_n1295_3[0]),.doutb(w_n1295_3[1]),.doutc(w_n1295_3[2]),.din(w_n1295_0[2]));
	jspl jspl_w_n1299_0(.douta(w_n1299_0[0]),.doutb(w_n1299_0[1]),.din(n1299));
	jspl jspl_w_n1300_0(.douta(w_n1300_0[0]),.doutb(w_n1300_0[1]),.din(n1300));
	jspl jspl_w_n1302_0(.douta(w_n1302_0[0]),.doutb(w_n1302_0[1]),.din(n1302));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(n1312));
	jspl jspl_w_n1313_0(.douta(w_n1313_0[0]),.doutb(w_n1313_0[1]),.din(n1313));
	jspl jspl_w_n1319_0(.douta(w_n1319_0[0]),.doutb(w_n1319_0[1]),.din(n1319));
	jspl3 jspl3_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.doutc(w_n1322_0[2]),.din(n1322));
	jspl3 jspl3_w_n1322_1(.douta(w_n1322_1[0]),.doutb(w_n1322_1[1]),.doutc(w_n1322_1[2]),.din(w_n1322_0[0]));
	jspl3 jspl3_w_n1331_0(.douta(w_n1331_0[0]),.doutb(w_n1331_0[1]),.doutc(w_n1331_0[2]),.din(n1331));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(n1332));
	jspl jspl_w_n1339_0(.douta(w_n1339_0[0]),.doutb(w_n1339_0[1]),.din(n1339));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(n1343));
	jspl3 jspl3_w_n1345_0(.douta(w_n1345_0[0]),.doutb(w_n1345_0[1]),.doutc(w_n1345_0[2]),.din(n1345));
	jspl3 jspl3_w_n1345_1(.douta(w_n1345_1[0]),.doutb(w_n1345_1[1]),.doutc(w_n1345_1[2]),.din(w_n1345_0[0]));
	jspl jspl_w_n1346_0(.douta(w_n1346_0[0]),.doutb(w_n1346_0[1]),.din(n1346));
	jspl3 jspl3_w_n1353_0(.douta(w_n1353_0[0]),.doutb(w_n1353_0[1]),.doutc(w_n1353_0[2]),.din(n1353));
	jspl3 jspl3_w_n1353_1(.douta(w_n1353_1[0]),.doutb(w_n1353_1[1]),.doutc(w_n1353_1[2]),.din(w_n1353_0[0]));
	jspl3 jspl3_w_n1353_2(.douta(w_n1353_2[0]),.doutb(w_n1353_2[1]),.doutc(w_n1353_2[2]),.din(w_n1353_0[1]));
	jspl3 jspl3_w_n1353_3(.douta(w_n1353_3[0]),.doutb(w_n1353_3[1]),.doutc(w_n1353_3[2]),.din(w_n1353_0[2]));
	jspl3 jspl3_w_n1353_4(.douta(w_n1353_4[0]),.doutb(w_n1353_4[1]),.doutc(w_n1353_4[2]),.din(w_n1353_1[0]));
	jspl3 jspl3_w_n1353_5(.douta(w_n1353_5[0]),.doutb(w_n1353_5[1]),.doutc(w_n1353_5[2]),.din(w_n1353_1[1]));
	jspl3 jspl3_w_n1354_0(.douta(w_n1354_0[0]),.doutb(w_n1354_0[1]),.doutc(w_n1354_0[2]),.din(n1354));
	jspl3 jspl3_w_n1354_1(.douta(w_n1354_1[0]),.doutb(w_n1354_1[1]),.doutc(w_n1354_1[2]),.din(w_n1354_0[0]));
	jspl3 jspl3_w_n1354_2(.douta(w_n1354_2[0]),.doutb(w_n1354_2[1]),.doutc(w_n1354_2[2]),.din(w_n1354_0[1]));
	jspl3 jspl3_w_n1354_3(.douta(w_n1354_3[0]),.doutb(w_n1354_3[1]),.doutc(w_n1354_3[2]),.din(w_n1354_0[2]));
	jspl3 jspl3_w_n1356_0(.douta(w_n1356_0[0]),.doutb(w_n1356_0[1]),.doutc(w_n1356_0[2]),.din(n1356));
	jspl3 jspl3_w_n1356_1(.douta(w_n1356_1[0]),.doutb(w_n1356_1[1]),.doutc(w_n1356_1[2]),.din(w_n1356_0[0]));
	jspl3 jspl3_w_n1356_2(.douta(w_n1356_2[0]),.doutb(w_n1356_2[1]),.doutc(w_n1356_2[2]),.din(w_n1356_0[1]));
	jspl3 jspl3_w_n1356_3(.douta(w_n1356_3[0]),.doutb(w_n1356_3[1]),.doutc(w_n1356_3[2]),.din(w_n1356_0[2]));
	jspl3 jspl3_w_n1356_4(.douta(w_n1356_4[0]),.doutb(w_n1356_4[1]),.doutc(w_n1356_4[2]),.din(w_n1356_1[0]));
	jspl3 jspl3_w_n1356_5(.douta(w_n1356_5[0]),.doutb(w_n1356_5[1]),.doutc(w_n1356_5[2]),.din(w_n1356_1[1]));
	jspl3 jspl3_w_n1356_6(.douta(w_n1356_6[0]),.doutb(w_n1356_6[1]),.doutc(w_n1356_6[2]),.din(w_n1356_1[2]));
	jspl3 jspl3_w_n1356_7(.douta(w_n1356_7[0]),.doutb(w_n1356_7[1]),.doutc(w_n1356_7[2]),.din(w_n1356_2[0]));
	jspl3 jspl3_w_n1356_8(.douta(w_n1356_8[0]),.doutb(w_n1356_8[1]),.doutc(w_n1356_8[2]),.din(w_n1356_2[1]));
	jspl3 jspl3_w_n1356_9(.douta(w_n1356_9[0]),.doutb(w_n1356_9[1]),.doutc(w_n1356_9[2]),.din(w_n1356_2[2]));
	jspl3 jspl3_w_n1356_10(.douta(w_n1356_10[0]),.doutb(w_n1356_10[1]),.doutc(w_n1356_10[2]),.din(w_n1356_3[0]));
	jspl3 jspl3_w_n1356_11(.douta(w_n1356_11[0]),.doutb(w_n1356_11[1]),.doutc(w_n1356_11[2]),.din(w_n1356_3[1]));
	jspl jspl_w_n1356_12(.douta(w_n1356_12[0]),.doutb(w_n1356_12[1]),.din(w_n1356_3[2]));
	jspl3 jspl3_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.doutc(w_n1360_0[2]),.din(n1360));
	jspl3 jspl3_w_n1360_1(.douta(w_n1360_1[0]),.doutb(w_n1360_1[1]),.doutc(w_n1360_1[2]),.din(w_n1360_0[0]));
	jspl3 jspl3_w_n1360_2(.douta(w_n1360_2[0]),.doutb(w_n1360_2[1]),.doutc(w_n1360_2[2]),.din(w_n1360_0[1]));
	jspl3 jspl3_w_n1360_3(.douta(w_n1360_3[0]),.doutb(w_n1360_3[1]),.doutc(w_n1360_3[2]),.din(w_n1360_0[2]));
	jspl3 jspl3_w_n1360_4(.douta(w_n1360_4[0]),.doutb(w_n1360_4[1]),.doutc(w_n1360_4[2]),.din(w_n1360_1[0]));
	jspl3 jspl3_w_n1360_5(.douta(w_n1360_5[0]),.doutb(w_n1360_5[1]),.doutc(w_n1360_5[2]),.din(w_n1360_1[1]));
	jspl jspl_w_n1360_6(.douta(w_n1360_6[0]),.doutb(w_n1360_6[1]),.din(w_n1360_1[2]));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(n1363));
	jspl3 jspl3_w_n1365_0(.douta(w_n1365_0[0]),.doutb(w_n1365_0[1]),.doutc(w_n1365_0[2]),.din(n1365));
	jspl3 jspl3_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.doutc(w_n1366_0[2]),.din(n1366));
	jspl jspl_w_n1366_1(.douta(w_n1366_1[0]),.doutb(w_n1366_1[1]),.din(w_n1366_0[0]));
	jspl jspl_w_n1375_0(.douta(w_n1375_0[0]),.doutb(w_n1375_0[1]),.din(n1375));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(n1378));
	jspl jspl_w_n1381_0(.douta(w_n1381_0[0]),.doutb(w_n1381_0[1]),.din(n1381));
	jspl jspl_w_n1385_0(.douta(w_n1385_0[0]),.doutb(w_n1385_0[1]),.din(n1385));
	jspl jspl_w_n1387_0(.douta(w_n1387_0[0]),.doutb(w_n1387_0[1]),.din(n1387));
	jspl jspl_w_n1392_0(.douta(w_n1392_0[0]),.doutb(w_n1392_0[1]),.din(n1392));
	jspl3 jspl3_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.doutc(w_n1400_0[2]),.din(n1400));
	jspl3 jspl3_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_n1402_0[1]),.doutc(w_n1402_0[2]),.din(n1402));
	jspl3 jspl3_w_n1402_1(.douta(w_n1402_1[0]),.doutb(w_n1402_1[1]),.doutc(w_n1402_1[2]),.din(w_n1402_0[0]));
	jspl3 jspl3_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.doutc(w_n1403_0[2]),.din(n1403));
	jspl jspl_w_n1403_1(.douta(w_n1403_1[0]),.doutb(w_n1403_1[1]),.din(w_n1403_0[0]));
	jspl3 jspl3_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_n1404_0[1]),.doutc(w_n1404_0[2]),.din(n1404));
	jspl jspl_w_n1406_0(.douta(w_n1406_0[0]),.doutb(w_n1406_0[1]),.din(n1406));
	jspl jspl_w_n1407_0(.douta(w_n1407_0[0]),.doutb(w_n1407_0[1]),.din(n1407));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(n1415));
	jspl3 jspl3_w_n1416_0(.douta(w_n1416_0[0]),.doutb(w_n1416_0[1]),.doutc(w_n1416_0[2]),.din(n1416));
	jspl3 jspl3_w_n1416_1(.douta(w_n1416_1[0]),.doutb(w_n1416_1[1]),.doutc(w_n1416_1[2]),.din(w_n1416_0[0]));
	jspl jspl_w_n1416_2(.douta(w_n1416_2[0]),.doutb(w_n1416_2[1]),.din(w_n1416_0[1]));
	jspl3 jspl3_w_n1418_0(.douta(w_n1418_0[0]),.doutb(w_n1418_0[1]),.doutc(w_n1418_0[2]),.din(n1418));
	jspl3 jspl3_w_n1418_1(.douta(w_n1418_1[0]),.doutb(w_n1418_1[1]),.doutc(w_n1418_1[2]),.din(w_n1418_0[0]));
	jspl3 jspl3_w_n1418_2(.douta(w_n1418_2[0]),.doutb(w_n1418_2[1]),.doutc(w_n1418_2[2]),.din(w_n1418_0[1]));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(n1426));
	jspl jspl_w_n1427_0(.douta(w_n1427_0[0]),.doutb(w_n1427_0[1]),.din(n1427));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1432_0(.douta(w_n1432_0[0]),.doutb(w_n1432_0[1]),.din(n1432));
	jspl3 jspl3_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.doutc(w_n1434_0[2]),.din(n1434));
	jspl3 jspl3_w_n1434_1(.douta(w_n1434_1[0]),.doutb(w_n1434_1[1]),.doutc(w_n1434_1[2]),.din(w_n1434_0[0]));
	jspl3 jspl3_w_n1434_2(.douta(w_n1434_2[0]),.doutb(w_n1434_2[1]),.doutc(w_n1434_2[2]),.din(w_n1434_0[1]));
	jspl3 jspl3_w_n1434_3(.douta(w_n1434_3[0]),.doutb(w_n1434_3[1]),.doutc(w_n1434_3[2]),.din(w_n1434_0[2]));
	jspl3 jspl3_w_n1434_4(.douta(w_n1434_4[0]),.doutb(w_n1434_4[1]),.doutc(w_n1434_4[2]),.din(w_n1434_1[0]));
	jspl3 jspl3_w_n1434_5(.douta(w_n1434_5[0]),.doutb(w_n1434_5[1]),.doutc(w_n1434_5[2]),.din(w_n1434_1[1]));
	jspl3 jspl3_w_n1434_6(.douta(w_n1434_6[0]),.doutb(w_n1434_6[1]),.doutc(w_n1434_6[2]),.din(w_n1434_1[2]));
	jspl3 jspl3_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_n1438_0[1]),.doutc(w_n1438_0[2]),.din(n1438));
	jspl3 jspl3_w_n1438_1(.douta(w_n1438_1[0]),.doutb(w_n1438_1[1]),.doutc(w_n1438_1[2]),.din(w_n1438_0[0]));
	jspl3 jspl3_w_n1438_2(.douta(w_n1438_2[0]),.doutb(w_n1438_2[1]),.doutc(w_n1438_2[2]),.din(w_n1438_0[1]));
	jspl3 jspl3_w_n1438_3(.douta(w_n1438_3[0]),.doutb(w_n1438_3[1]),.doutc(w_n1438_3[2]),.din(w_n1438_0[2]));
	jspl3 jspl3_w_n1438_4(.douta(w_n1438_4[0]),.doutb(w_n1438_4[1]),.doutc(w_n1438_4[2]),.din(w_n1438_1[0]));
	jspl3 jspl3_w_n1438_5(.douta(w_n1438_5[0]),.doutb(w_n1438_5[1]),.doutc(w_n1438_5[2]),.din(w_n1438_1[1]));
	jspl3 jspl3_w_n1438_6(.douta(w_n1438_6[0]),.doutb(w_n1438_6[1]),.doutc(w_n1438_6[2]),.din(w_n1438_1[2]));
	jspl3 jspl3_w_n1438_7(.douta(w_n1438_7[0]),.doutb(w_n1438_7[1]),.doutc(w_n1438_7[2]),.din(w_n1438_2[0]));
	jspl3 jspl3_w_n1438_8(.douta(w_n1438_8[0]),.doutb(w_n1438_8[1]),.doutc(w_n1438_8[2]),.din(w_n1438_2[1]));
	jspl3 jspl3_w_n1438_9(.douta(w_n1438_9[0]),.doutb(w_n1438_9[1]),.doutc(w_n1438_9[2]),.din(w_n1438_2[2]));
	jspl3 jspl3_w_n1438_10(.douta(w_n1438_10[0]),.doutb(w_n1438_10[1]),.doutc(w_n1438_10[2]),.din(w_n1438_3[0]));
	jspl3 jspl3_w_n1438_11(.douta(w_n1438_11[0]),.doutb(w_n1438_11[1]),.doutc(w_n1438_11[2]),.din(w_n1438_3[1]));
	jspl3 jspl3_w_n1438_12(.douta(w_n1438_12[0]),.doutb(w_n1438_12[1]),.doutc(w_n1438_12[2]),.din(w_n1438_3[2]));
	jspl3 jspl3_w_n1438_13(.douta(w_n1438_13[0]),.doutb(w_n1438_13[1]),.doutc(w_n1438_13[2]),.din(w_n1438_4[0]));
	jspl3 jspl3_w_n1438_14(.douta(w_n1438_14[0]),.doutb(w_n1438_14[1]),.doutc(w_n1438_14[2]),.din(w_n1438_4[1]));
	jspl3 jspl3_w_n1438_15(.douta(w_n1438_15[0]),.doutb(w_n1438_15[1]),.doutc(w_n1438_15[2]),.din(w_n1438_4[2]));
	jspl3 jspl3_w_n1438_16(.douta(w_n1438_16[0]),.doutb(w_n1438_16[1]),.doutc(w_n1438_16[2]),.din(w_n1438_5[0]));
	jspl3 jspl3_w_n1438_17(.douta(w_n1438_17[0]),.doutb(w_n1438_17[1]),.doutc(w_n1438_17[2]),.din(w_n1438_5[1]));
	jspl3 jspl3_w_n1438_18(.douta(w_n1438_18[0]),.doutb(w_n1438_18[1]),.doutc(w_n1438_18[2]),.din(w_n1438_5[2]));
	jspl3 jspl3_w_n1438_19(.douta(w_n1438_19[0]),.doutb(w_n1438_19[1]),.doutc(w_n1438_19[2]),.din(w_n1438_6[0]));
	jspl3 jspl3_w_n1438_20(.douta(w_n1438_20[0]),.doutb(w_n1438_20[1]),.doutc(w_n1438_20[2]),.din(w_n1438_6[1]));
	jspl jspl_w_n1438_21(.douta(w_n1438_21[0]),.doutb(w_n1438_21[1]),.din(w_n1438_6[2]));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(n1444));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1448_0(.douta(w_n1448_0[0]),.doutb(w_n1448_0[1]),.din(n1448));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1456_0(.douta(w_n1456_0[0]),.doutb(w_n1456_0[1]),.din(n1456));
	jspl3 jspl3_w_n1459_0(.douta(w_n1459_0[0]),.doutb(w_n1459_0[1]),.doutc(w_n1459_0[2]),.din(n1459));
	jspl3 jspl3_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.doutc(w_n1460_0[2]),.din(n1460));
	jspl3 jspl3_w_n1460_1(.douta(w_n1460_1[0]),.doutb(w_n1460_1[1]),.doutc(w_n1460_1[2]),.din(w_n1460_0[0]));
	jspl jspl_w_n1467_0(.douta(w_n1467_0[0]),.doutb(w_n1467_0[1]),.din(n1467));
	jspl jspl_w_n1470_0(.douta(w_n1470_0[0]),.doutb(w_n1470_0[1]),.din(n1470));
	jspl3 jspl3_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.doutc(w_n1474_0[2]),.din(n1474));
	jspl3 jspl3_w_n1474_1(.douta(w_n1474_1[0]),.doutb(w_n1474_1[1]),.doutc(w_n1474_1[2]),.din(w_n1474_0[0]));
	jspl3 jspl3_w_n1474_2(.douta(w_n1474_2[0]),.doutb(w_n1474_2[1]),.doutc(w_n1474_2[2]),.din(w_n1474_0[1]));
	jspl3 jspl3_w_n1474_3(.douta(w_n1474_3[0]),.doutb(w_n1474_3[1]),.doutc(w_n1474_3[2]),.din(w_n1474_0[2]));
	jspl3 jspl3_w_n1474_4(.douta(w_n1474_4[0]),.doutb(w_n1474_4[1]),.doutc(w_n1474_4[2]),.din(w_n1474_1[0]));
	jspl3 jspl3_w_n1474_5(.douta(w_n1474_5[0]),.doutb(w_n1474_5[1]),.doutc(w_n1474_5[2]),.din(w_n1474_1[1]));
	jspl3 jspl3_w_n1474_6(.douta(w_n1474_6[0]),.doutb(w_n1474_6[1]),.doutc(w_n1474_6[2]),.din(w_n1474_1[2]));
	jspl jspl_w_n1474_7(.douta(w_n1474_7[0]),.doutb(w_n1474_7[1]),.din(w_n1474_2[0]));
	jspl jspl_w_n1478_0(.douta(w_n1478_0[0]),.doutb(w_n1478_0[1]),.din(n1478));
	jspl3 jspl3_w_n1480_0(.douta(w_n1480_0[0]),.doutb(w_n1480_0[1]),.doutc(w_n1480_0[2]),.din(n1480));
	jspl3 jspl3_w_n1480_1(.douta(w_n1480_1[0]),.doutb(w_n1480_1[1]),.doutc(w_n1480_1[2]),.din(w_n1480_0[0]));
	jspl3 jspl3_w_n1480_2(.douta(w_n1480_2[0]),.doutb(w_n1480_2[1]),.doutc(w_n1480_2[2]),.din(w_n1480_0[1]));
	jspl3 jspl3_w_n1480_3(.douta(w_n1480_3[0]),.doutb(w_n1480_3[1]),.doutc(w_n1480_3[2]),.din(w_n1480_0[2]));
	jspl3 jspl3_w_n1480_4(.douta(w_n1480_4[0]),.doutb(w_n1480_4[1]),.doutc(w_n1480_4[2]),.din(w_n1480_1[0]));
	jspl3 jspl3_w_n1480_5(.douta(w_n1480_5[0]),.doutb(w_n1480_5[1]),.doutc(w_n1480_5[2]),.din(w_n1480_1[1]));
	jspl3 jspl3_w_n1480_6(.douta(w_n1480_6[0]),.doutb(w_n1480_6[1]),.doutc(w_n1480_6[2]),.din(w_n1480_1[2]));
	jspl3 jspl3_w_n1480_7(.douta(w_n1480_7[0]),.doutb(w_n1480_7[1]),.doutc(w_n1480_7[2]),.din(w_n1480_2[0]));
	jspl3 jspl3_w_n1480_8(.douta(w_n1480_8[0]),.doutb(w_n1480_8[1]),.doutc(w_n1480_8[2]),.din(w_n1480_2[1]));
	jspl3 jspl3_w_n1480_9(.douta(w_n1480_9[0]),.doutb(w_n1480_9[1]),.doutc(w_n1480_9[2]),.din(w_n1480_2[2]));
	jspl jspl_w_n1480_10(.douta(w_n1480_10[0]),.doutb(w_n1480_10[1]),.din(w_n1480_3[0]));
	jspl3 jspl3_w_n1485_0(.douta(w_n1485_0[0]),.doutb(w_n1485_0[1]),.doutc(w_n1485_0[2]),.din(n1485));
	jspl3 jspl3_w_n1485_1(.douta(w_n1485_1[0]),.doutb(w_n1485_1[1]),.doutc(w_n1485_1[2]),.din(w_n1485_0[0]));
	jspl3 jspl3_w_n1485_2(.douta(w_n1485_2[0]),.doutb(w_n1485_2[1]),.doutc(w_n1485_2[2]),.din(w_n1485_0[1]));
	jspl3 jspl3_w_n1485_3(.douta(w_n1485_3[0]),.doutb(w_n1485_3[1]),.doutc(w_n1485_3[2]),.din(w_n1485_0[2]));
	jspl3 jspl3_w_n1485_4(.douta(w_n1485_4[0]),.doutb(w_n1485_4[1]),.doutc(w_n1485_4[2]),.din(w_n1485_1[0]));
	jspl jspl_w_n1489_0(.douta(w_n1489_0[0]),.doutb(w_n1489_0[1]),.din(n1489));
	jspl3 jspl3_w_n1490_0(.douta(w_n1490_0[0]),.doutb(w_n1490_0[1]),.doutc(w_n1490_0[2]),.din(n1490));
	jspl3 jspl3_w_n1490_1(.douta(w_n1490_1[0]),.doutb(w_n1490_1[1]),.doutc(w_n1490_1[2]),.din(w_n1490_0[0]));
	jspl3 jspl3_w_n1490_2(.douta(w_n1490_2[0]),.doutb(w_n1490_2[1]),.doutc(w_n1490_2[2]),.din(w_n1490_0[1]));
	jspl3 jspl3_w_n1490_3(.douta(w_n1490_3[0]),.doutb(w_n1490_3[1]),.doutc(w_n1490_3[2]),.din(w_n1490_0[2]));
	jspl3 jspl3_w_n1490_4(.douta(w_n1490_4[0]),.doutb(w_n1490_4[1]),.doutc(w_n1490_4[2]),.din(w_n1490_1[0]));
	jspl jspl_w_n1490_5(.douta(w_n1490_5[0]),.doutb(w_n1490_5[1]),.din(w_n1490_1[1]));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(n1491));
	jspl3 jspl3_w_n1493_0(.douta(w_n1493_0[0]),.doutb(w_n1493_0[1]),.doutc(w_n1493_0[2]),.din(n1493));
	jspl3 jspl3_w_n1493_1(.douta(w_n1493_1[0]),.doutb(w_n1493_1[1]),.doutc(w_n1493_1[2]),.din(w_n1493_0[0]));
	jspl3 jspl3_w_n1493_2(.douta(w_n1493_2[0]),.doutb(w_n1493_2[1]),.doutc(w_n1493_2[2]),.din(w_n1493_0[1]));
	jspl3 jspl3_w_n1493_3(.douta(w_n1493_3[0]),.doutb(w_n1493_3[1]),.doutc(w_n1493_3[2]),.din(w_n1493_0[2]));
	jspl3 jspl3_w_n1493_4(.douta(w_n1493_4[0]),.doutb(w_n1493_4[1]),.doutc(w_n1493_4[2]),.din(w_n1493_1[0]));
	jspl jspl_w_n1493_5(.douta(w_n1493_5[0]),.doutb(w_n1493_5[1]),.din(w_n1493_1[1]));
	jspl3 jspl3_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.doutc(w_n1494_0[2]),.din(n1494));
	jspl3 jspl3_w_n1494_1(.douta(w_n1494_1[0]),.doutb(w_n1494_1[1]),.doutc(w_n1494_1[2]),.din(w_n1494_0[0]));
	jspl3 jspl3_w_n1494_2(.douta(w_n1494_2[0]),.doutb(w_n1494_2[1]),.doutc(w_n1494_2[2]),.din(w_n1494_0[1]));
	jspl3 jspl3_w_n1494_3(.douta(w_n1494_3[0]),.doutb(w_n1494_3[1]),.doutc(w_n1494_3[2]),.din(w_n1494_0[2]));
	jspl3 jspl3_w_n1494_4(.douta(w_n1494_4[0]),.doutb(w_n1494_4[1]),.doutc(w_n1494_4[2]),.din(w_n1494_1[0]));
	jspl3 jspl3_w_n1494_5(.douta(w_n1494_5[0]),.doutb(w_n1494_5[1]),.doutc(w_n1494_5[2]),.din(w_n1494_1[1]));
	jspl jspl_w_n1494_6(.douta(w_n1494_6[0]),.doutb(w_n1494_6[1]),.din(w_n1494_1[2]));
	jspl3 jspl3_w_n1499_0(.douta(w_n1499_0[0]),.doutb(w_n1499_0[1]),.doutc(w_n1499_0[2]),.din(n1499));
	jspl3 jspl3_w_n1499_1(.douta(w_n1499_1[0]),.doutb(w_n1499_1[1]),.doutc(w_n1499_1[2]),.din(w_n1499_0[0]));
	jspl3 jspl3_w_n1499_2(.douta(w_n1499_2[0]),.doutb(w_n1499_2[1]),.doutc(w_n1499_2[2]),.din(w_n1499_0[1]));
	jspl3 jspl3_w_n1499_3(.douta(w_n1499_3[0]),.doutb(w_n1499_3[1]),.doutc(w_n1499_3[2]),.din(w_n1499_0[2]));
	jspl3 jspl3_w_n1499_4(.douta(w_n1499_4[0]),.doutb(w_n1499_4[1]),.doutc(w_n1499_4[2]),.din(w_n1499_1[0]));
	jspl3 jspl3_w_n1499_5(.douta(w_n1499_5[0]),.doutb(w_n1499_5[1]),.doutc(w_n1499_5[2]),.din(w_n1499_1[1]));
	jspl3 jspl3_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.doutc(w_n1500_0[2]),.din(n1500));
	jspl3 jspl3_w_n1500_1(.douta(w_n1500_1[0]),.doutb(w_n1500_1[1]),.doutc(w_n1500_1[2]),.din(w_n1500_0[0]));
	jspl3 jspl3_w_n1500_2(.douta(w_n1500_2[0]),.doutb(w_n1500_2[1]),.doutc(w_n1500_2[2]),.din(w_n1500_0[1]));
	jspl3 jspl3_w_n1500_3(.douta(w_n1500_3[0]),.doutb(w_n1500_3[1]),.doutc(w_n1500_3[2]),.din(w_n1500_0[2]));
	jspl3 jspl3_w_n1500_4(.douta(w_n1500_4[0]),.doutb(w_n1500_4[1]),.doutc(w_n1500_4[2]),.din(w_n1500_1[0]));
	jspl jspl_w_n1500_5(.douta(w_n1500_5[0]),.doutb(w_n1500_5[1]),.din(w_n1500_1[1]));
	jspl3 jspl3_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.doutc(w_n1504_0[2]),.din(n1504));
	jspl3 jspl3_w_n1504_1(.douta(w_n1504_1[0]),.doutb(w_n1504_1[1]),.doutc(w_n1504_1[2]),.din(w_n1504_0[0]));
	jspl3 jspl3_w_n1504_2(.douta(w_n1504_2[0]),.doutb(w_n1504_2[1]),.doutc(w_n1504_2[2]),.din(w_n1504_0[1]));
	jspl3 jspl3_w_n1504_3(.douta(w_n1504_3[0]),.doutb(w_n1504_3[1]),.doutc(w_n1504_3[2]),.din(w_n1504_0[2]));
	jspl3 jspl3_w_n1505_0(.douta(w_n1505_0[0]),.doutb(w_n1505_0[1]),.doutc(w_n1505_0[2]),.din(n1505));
	jspl3 jspl3_w_n1505_1(.douta(w_n1505_1[0]),.doutb(w_n1505_1[1]),.doutc(w_n1505_1[2]),.din(w_n1505_0[0]));
	jspl3 jspl3_w_n1505_2(.douta(w_n1505_2[0]),.doutb(w_n1505_2[1]),.doutc(w_n1505_2[2]),.din(w_n1505_0[1]));
	jspl3 jspl3_w_n1505_3(.douta(w_n1505_3[0]),.doutb(w_n1505_3[1]),.doutc(w_n1505_3[2]),.din(w_n1505_0[2]));
	jspl3 jspl3_w_n1505_4(.douta(w_n1505_4[0]),.doutb(w_n1505_4[1]),.doutc(w_n1505_4[2]),.din(w_n1505_1[0]));
	jspl jspl_w_n1508_0(.douta(w_n1508_0[0]),.doutb(w_n1508_0[1]),.din(n1508));
	jspl jspl_w_n1509_0(.douta(w_n1509_0[0]),.doutb(w_n1509_0[1]),.din(n1509));
	jspl jspl_w_n1511_0(.douta(w_n1511_0[0]),.doutb(w_n1511_0[1]),.din(n1511));
	jspl jspl_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.din(n1513));
	jspl3 jspl3_w_n1516_0(.douta(w_n1516_0[0]),.doutb(w_n1516_0[1]),.doutc(w_n1516_0[2]),.din(n1516));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.din(n1520));
	jspl jspl_w_n1523_0(.douta(w_n1523_0[0]),.doutb(w_n1523_0[1]),.din(n1523));
	jspl jspl_w_n1528_0(.douta(w_n1528_0[0]),.doutb(w_n1528_0[1]),.din(n1528));
	jspl3 jspl3_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.doutc(w_n1529_0[2]),.din(n1529));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(n1531));
	jspl3 jspl3_w_n1532_0(.douta(w_n1532_0[0]),.doutb(w_n1532_0[1]),.doutc(w_n1532_0[2]),.din(n1532));
	jspl jspl_w_n1533_0(.douta(w_n1533_0[0]),.doutb(w_n1533_0[1]),.din(n1533));
	jspl3 jspl3_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.doutc(w_n1534_0[2]),.din(n1534));
	jspl3 jspl3_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.doutc(w_n1539_0[2]),.din(n1539));
	jspl3 jspl3_w_n1539_1(.douta(w_n1539_1[0]),.doutb(w_n1539_1[1]),.doutc(w_n1539_1[2]),.din(w_n1539_0[0]));
	jspl3 jspl3_w_n1539_2(.douta(w_n1539_2[0]),.doutb(w_n1539_2[1]),.doutc(w_n1539_2[2]),.din(w_n1539_0[1]));
	jspl jspl_w_n1541_0(.douta(w_n1541_0[0]),.doutb(w_n1541_0[1]),.din(n1541));
	jspl3 jspl3_w_n1542_0(.douta(w_n1542_0[0]),.doutb(w_n1542_0[1]),.doutc(w_n1542_0[2]),.din(n1542));
	jspl3 jspl3_w_n1542_1(.douta(w_n1542_1[0]),.doutb(w_n1542_1[1]),.doutc(w_n1542_1[2]),.din(w_n1542_0[0]));
	jspl3 jspl3_w_n1542_2(.douta(w_n1542_2[0]),.doutb(w_n1542_2[1]),.doutc(w_n1542_2[2]),.din(w_n1542_0[1]));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1547_0(.douta(w_n1547_0[0]),.doutb(w_n1547_0[1]),.din(n1547));
	jspl3 jspl3_w_n1549_0(.douta(w_n1549_0[0]),.doutb(w_n1549_0[1]),.doutc(w_n1549_0[2]),.din(n1549));
	jspl3 jspl3_w_n1549_1(.douta(w_n1549_1[0]),.doutb(w_n1549_1[1]),.doutc(w_n1549_1[2]),.din(w_n1549_0[0]));
	jspl3 jspl3_w_n1549_2(.douta(w_n1549_2[0]),.doutb(w_n1549_2[1]),.doutc(w_n1549_2[2]),.din(w_n1549_0[1]));
	jspl3 jspl3_w_n1549_3(.douta(w_n1549_3[0]),.doutb(w_n1549_3[1]),.doutc(w_n1549_3[2]),.din(w_n1549_0[2]));
	jspl3 jspl3_w_n1549_4(.douta(w_n1549_4[0]),.doutb(w_n1549_4[1]),.doutc(w_n1549_4[2]),.din(w_n1549_1[0]));
	jspl3 jspl3_w_n1551_0(.douta(w_n1551_0[0]),.doutb(w_n1551_0[1]),.doutc(w_n1551_0[2]),.din(n1551));
	jspl3 jspl3_w_n1551_1(.douta(w_n1551_1[0]),.doutb(w_n1551_1[1]),.doutc(w_n1551_1[2]),.din(w_n1551_0[0]));
	jspl3 jspl3_w_n1551_2(.douta(w_n1551_2[0]),.doutb(w_n1551_2[1]),.doutc(w_n1551_2[2]),.din(w_n1551_0[1]));
	jspl3 jspl3_w_n1551_3(.douta(w_n1551_3[0]),.doutb(w_n1551_3[1]),.doutc(w_n1551_3[2]),.din(w_n1551_0[2]));
	jspl3 jspl3_w_n1551_4(.douta(w_n1551_4[0]),.doutb(w_n1551_4[1]),.doutc(w_n1551_4[2]),.din(w_n1551_1[0]));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(n1555));
	jspl jspl_w_n1556_0(.douta(w_n1556_0[0]),.doutb(w_n1556_0[1]),.din(n1556));
	jspl jspl_w_n1557_0(.douta(w_n1557_0[0]),.doutb(w_n1557_0[1]),.din(n1557));
	jspl3 jspl3_w_n1558_0(.douta(w_n1558_0[0]),.doutb(w_n1558_0[1]),.doutc(w_n1558_0[2]),.din(n1558));
	jspl3 jspl3_w_n1558_1(.douta(w_n1558_1[0]),.doutb(w_n1558_1[1]),.doutc(w_n1558_1[2]),.din(w_n1558_0[0]));
	jspl3 jspl3_w_n1558_2(.douta(w_n1558_2[0]),.doutb(w_n1558_2[1]),.doutc(w_n1558_2[2]),.din(w_n1558_0[1]));
	jspl3 jspl3_w_n1558_3(.douta(w_n1558_3[0]),.doutb(w_n1558_3[1]),.doutc(w_n1558_3[2]),.din(w_n1558_0[2]));
	jspl jspl_w_n1558_4(.douta(w_n1558_4[0]),.doutb(w_n1558_4[1]),.din(w_n1558_1[0]));
	jspl3 jspl3_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.doutc(w_n1560_0[2]),.din(n1560));
	jspl3 jspl3_w_n1560_1(.douta(w_n1560_1[0]),.doutb(w_n1560_1[1]),.doutc(w_n1560_1[2]),.din(w_n1560_0[0]));
	jspl3 jspl3_w_n1560_2(.douta(w_n1560_2[0]),.doutb(w_n1560_2[1]),.doutc(w_n1560_2[2]),.din(w_n1560_0[1]));
	jspl3 jspl3_w_n1560_3(.douta(w_n1560_3[0]),.doutb(w_n1560_3[1]),.doutc(w_n1560_3[2]),.din(w_n1560_0[2]));
	jspl3 jspl3_w_n1560_4(.douta(w_n1560_4[0]),.doutb(w_n1560_4[1]),.doutc(w_n1560_4[2]),.din(w_n1560_1[0]));
	jspl jspl_w_n1563_0(.douta(w_n1563_0[0]),.doutb(w_n1563_0[1]),.din(n1563));
	jspl jspl_w_n1564_0(.douta(w_n1564_0[0]),.doutb(w_n1564_0[1]),.din(n1564));
	jspl jspl_w_n1566_0(.douta(w_n1566_0[0]),.doutb(w_n1566_0[1]),.din(n1566));
	jspl jspl_w_n1567_0(.douta(w_n1567_0[0]),.doutb(w_n1567_0[1]),.din(n1567));
	jspl jspl_w_n1575_0(.douta(w_n1575_0[0]),.doutb(w_n1575_0[1]),.din(n1575));
	jspl3 jspl3_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.doutc(w_n1576_0[2]),.din(n1576));
	jspl jspl_w_n1584_0(.douta(w_n1584_0[0]),.doutb(w_n1584_0[1]),.din(n1584));
	jspl jspl_w_n1592_0(.douta(w_n1592_0[0]),.doutb(w_n1592_0[1]),.din(n1592));
	jspl jspl_w_n1593_0(.douta(w_n1593_0[0]),.doutb(w_n1593_0[1]),.din(n1593));
	jspl jspl_w_n1594_0(.douta(w_n1594_0[0]),.doutb(w_n1594_0[1]),.din(n1594));
	jspl jspl_w_n1595_0(.douta(w_n1595_0[0]),.doutb(w_n1595_0[1]),.din(n1595));
	jspl jspl_w_n1598_0(.douta(w_n1598_0[0]),.doutb(w_n1598_0[1]),.din(n1598));
	jspl jspl_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.din(n1601));
	jspl jspl_w_n1604_0(.douta(w_n1604_0[0]),.doutb(w_n1604_0[1]),.din(n1604));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1613_0(.douta(w_n1613_0[0]),.doutb(w_n1613_0[1]),.din(n1613));
	jspl jspl_w_n1614_0(.douta(w_n1614_0[0]),.doutb(w_n1614_0[1]),.din(n1614));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(n1615));
	jspl jspl_w_n1616_0(.douta(w_n1616_0[0]),.doutb(w_n1616_0[1]),.din(n1616));
	jspl3 jspl3_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.doutc(w_n1622_0[2]),.din(n1622));
	jspl3 jspl3_w_n1622_1(.douta(w_n1622_1[0]),.doutb(w_n1622_1[1]),.doutc(w_n1622_1[2]),.din(w_n1622_0[0]));
	jspl3 jspl3_w_n1622_2(.douta(w_n1622_2[0]),.doutb(w_n1622_2[1]),.doutc(w_n1622_2[2]),.din(w_n1622_0[1]));
	jspl3 jspl3_w_n1622_3(.douta(w_n1622_3[0]),.doutb(w_n1622_3[1]),.doutc(w_n1622_3[2]),.din(w_n1622_0[2]));
	jspl jspl_w_n1622_4(.douta(w_n1622_4[0]),.doutb(w_n1622_4[1]),.din(w_n1622_1[0]));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl jspl_w_n1626_0(.douta(w_n1626_0[0]),.doutb(w_n1626_0[1]),.din(n1626));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1630_0(.douta(w_n1630_0[0]),.doutb(w_n1630_0[1]),.din(n1630));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(n1631));
	jspl jspl_w_n1632_0(.douta(w_n1632_0[0]),.doutb(w_n1632_0[1]),.din(n1632));
	jspl jspl_w_n1640_0(.douta(w_n1640_0[0]),.doutb(w_n1640_0[1]),.din(n1640));
	jspl jspl_w_n1648_0(.douta(w_n1648_0[0]),.doutb(w_n1648_0[1]),.din(n1648));
	jspl3 jspl3_w_n1649_0(.douta(w_n1649_0[0]),.doutb(w_n1649_0[1]),.doutc(w_n1649_0[2]),.din(n1649));
	jspl3 jspl3_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.doutc(w_n1651_0[2]),.din(n1651));
	jspl jspl_w_n1651_1(.douta(w_n1651_1[0]),.doutb(w_n1651_1[1]),.din(w_n1651_0[0]));
	jspl3 jspl3_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.doutc(w_n1656_0[2]),.din(n1656));
	jspl3 jspl3_w_n1656_1(.douta(w_n1656_1[0]),.doutb(w_n1656_1[1]),.doutc(w_n1656_1[2]),.din(w_n1656_0[0]));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1660_0(.douta(w_n1660_0[0]),.doutb(w_n1660_0[1]),.din(n1660));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(n1661));
	jspl jspl_w_n1662_0(.douta(w_n1662_0[0]),.doutb(w_n1662_0[1]),.din(n1662));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(n1663));
	jspl3 jspl3_w_n1664_0(.douta(w_n1664_0[0]),.doutb(w_n1664_0[1]),.doutc(w_n1664_0[2]),.din(n1664));
	jspl jspl_w_n1673_0(.douta(w_n1673_0[0]),.doutb(w_n1673_0[1]),.din(n1673));
	jspl jspl_w_n1674_0(.douta(w_n1674_0[0]),.doutb(w_n1674_0[1]),.din(n1674));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_n1687_0[1]),.din(n1687));
	jspl jspl_w_n1696_0(.douta(w_n1696_0[0]),.doutb(w_n1696_0[1]),.din(n1696));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_n1697_0[1]),.din(n1697));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(n1699));
	jspl jspl_w_n1700_0(.douta(w_n1700_0[0]),.doutb(w_n1700_0[1]),.din(n1700));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(n1702));
	jspl jspl_w_n1703_0(.douta(w_n1703_0[0]),.doutb(w_n1703_0[1]),.din(n1703));
	jspl jspl_w_n1705_0(.douta(w_n1705_0[0]),.doutb(w_n1705_0[1]),.din(n1705));
	jspl jspl_w_n1706_0(.douta(w_n1706_0[0]),.doutb(w_n1706_0[1]),.din(n1706));
	jspl jspl_w_n1708_0(.douta(w_n1708_0[0]),.doutb(w_n1708_0[1]),.din(n1708));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(n1709));
	jspl jspl_w_n1710_0(.douta(w_n1710_0[0]),.doutb(w_n1710_0[1]),.din(n1710));
	jspl jspl_w_n1718_0(.douta(w_n1718_0[0]),.doutb(w_n1718_0[1]),.din(n1718));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1733_0(.douta(w_n1733_0[0]),.doutb(w_n1733_0[1]),.din(n1733));
	jspl jspl_w_n1734_0(.douta(w_n1734_0[0]),.doutb(w_n1734_0[1]),.din(n1734));
	jspl jspl_w_n1736_0(.douta(w_n1736_0[0]),.doutb(w_n1736_0[1]),.din(n1736));
	jspl jspl_w_n1737_0(.douta(w_n1737_0[0]),.doutb(w_n1737_0[1]),.din(n1737));
	jspl jspl_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.din(n1743));
	jspl3 jspl3_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.doutc(w_n1744_0[2]),.din(n1744));
	jspl jspl_w_n1746_0(.douta(w_n1746_0[0]),.doutb(w_n1746_0[1]),.din(n1746));
	jspl jspl_w_n1747_0(.douta(w_n1747_0[0]),.doutb(w_n1747_0[1]),.din(n1747));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1759_0(.douta(w_n1759_0[0]),.doutb(w_n1759_0[1]),.din(n1759));
	jspl jspl_w_n1763_0(.douta(w_n1763_0[0]),.doutb(w_n1763_0[1]),.din(n1763));
	jspl jspl_w_n1764_0(.douta(w_n1764_0[0]),.doutb(w_n1764_0[1]),.din(n1764));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl jspl_w_n1766_0(.douta(w_n1766_0[0]),.doutb(w_n1766_0[1]),.din(n1766));
	jspl3 jspl3_w_n1767_0(.douta(w_n1767_0[0]),.doutb(w_n1767_0[1]),.doutc(w_n1767_0[2]),.din(n1767));
	jspl jspl_w_n1768_0(.douta(w_n1768_0[0]),.doutb(w_n1768_0[1]),.din(n1768));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(n1770));
	jspl jspl_w_n1778_0(.douta(w_n1778_0[0]),.doutb(w_n1778_0[1]),.din(n1778));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1793_0(.douta(w_n1793_0[0]),.doutb(w_n1793_0[1]),.din(n1793));
	jspl jspl_w_n1794_0(.douta(w_n1794_0[0]),.doutb(w_n1794_0[1]),.din(n1794));
	jspl jspl_w_n1796_0(.douta(w_n1796_0[0]),.doutb(w_n1796_0[1]),.din(n1796));
	jspl jspl_w_n1799_0(.douta(w_n1799_0[0]),.doutb(w_n1799_0[1]),.din(n1799));
	jspl jspl_w_n1800_0(.douta(w_n1800_0[0]),.doutb(w_n1800_0[1]),.din(n1800));
	jspl jspl_w_n1802_0(.douta(w_n1802_0[0]),.doutb(w_n1802_0[1]),.din(n1802));
	jspl jspl_w_n1804_0(.douta(w_n1804_0[0]),.doutb(w_n1804_0[1]),.din(n1804));
	jspl jspl_w_n1806_0(.douta(w_n1806_0[0]),.doutb(w_n1806_0[1]),.din(n1806));
	jspl jspl_w_n1811_0(.douta(w_n1811_0[0]),.doutb(w_n1811_0[1]),.din(n1811));
	jspl jspl_w_n1812_0(.douta(w_n1812_0[0]),.doutb(w_n1812_0[1]),.din(n1812));
	jspl3 jspl3_w_n1813_0(.douta(w_n1813_0[0]),.doutb(w_n1813_0[1]),.doutc(w_n1813_0[2]),.din(n1813));
	jspl jspl_w_n1813_1(.douta(w_n1813_1[0]),.doutb(w_n1813_1[1]),.din(w_n1813_0[0]));
	jspl jspl_w_n1814_0(.douta(w_n1814_0[0]),.doutb(w_n1814_0[1]),.din(n1814));
	jspl jspl_w_n1815_0(.douta(w_n1815_0[0]),.doutb(w_n1815_0[1]),.din(n1815));
	jspl jspl_w_n1823_0(.douta(w_n1823_0[0]),.doutb(w_n1823_0[1]),.din(n1823));
	jspl jspl_w_n1830_0(.douta(w_n1830_0[0]),.doutb(w_n1830_0[1]),.din(n1830));
	jspl jspl_w_n1832_0(.douta(w_n1832_0[0]),.doutb(w_n1832_0[1]),.din(n1832));
	jspl jspl_w_n1833_0(.douta(w_n1833_0[0]),.doutb(w_n1833_0[1]),.din(n1833));
	jspl jspl_w_n1835_0(.douta(w_n1835_0[0]),.doutb(w_n1835_0[1]),.din(n1835));
	jspl jspl_w_n1836_0(.douta(w_n1836_0[0]),.doutb(w_n1836_0[1]),.din(n1836));
	jspl jspl_w_n1838_0(.douta(w_n1838_0[0]),.doutb(w_n1838_0[1]),.din(n1838));
	jspl jspl_w_n1839_0(.douta(w_n1839_0[0]),.doutb(w_n1839_0[1]),.din(n1839));
	jspl jspl_w_n1840_0(.douta(w_n1840_0[0]),.doutb(w_n1840_0[1]),.din(n1840));
	jspl jspl_w_n1842_0(.douta(w_n1842_0[0]),.doutb(w_n1842_0[1]),.din(n1842));
	jspl jspl_w_n1843_0(.douta(w_n1843_0[0]),.doutb(w_n1843_0[1]),.din(n1843));
	jspl jspl_w_n1844_0(.douta(w_n1844_0[0]),.doutb(w_n1844_0[1]),.din(n1844));
	jspl jspl_w_n1846_0(.douta(w_n1846_0[0]),.doutb(w_n1846_0[1]),.din(n1846));
	jspl jspl_w_n1850_0(.douta(w_n1850_0[0]),.doutb(w_n1850_0[1]),.din(n1850));
	jspl jspl_w_n1860_0(.douta(w_n1860_0[0]),.doutb(w_n1860_0[1]),.din(n1860));
	jspl jspl_w_n1865_0(.douta(w_n1865_0[0]),.doutb(w_n1865_0[1]),.din(n1865));
	jspl jspl_w_n1867_0(.douta(w_n1867_0[0]),.doutb(w_n1867_0[1]),.din(n1867));
	jspl3 jspl3_w_n1868_0(.douta(w_n1868_0[0]),.doutb(w_n1868_0[1]),.doutc(w_n1868_0[2]),.din(n1868));
	jspl jspl_w_n1873_0(.douta(w_n1873_0[0]),.doutb(w_n1873_0[1]),.din(n1873));
	jspl jspl_w_n1885_0(.douta(w_n1885_0[0]),.doutb(w_n1885_0[1]),.din(n1885));
	jspl jspl_w_n1886_0(.douta(w_n1886_0[0]),.doutb(w_n1886_0[1]),.din(n1886));
	jspl jspl_w_n1888_0(.douta(w_n1888_0[0]),.doutb(w_n1888_0[1]),.din(n1888));
	jspl3 jspl3_w_n1890_0(.douta(w_n1890_0[0]),.doutb(w_n1890_0[1]),.doutc(w_n1890_0[2]),.din(n1890));
	jspl3 jspl3_w_n1895_0(.douta(w_n1895_0[0]),.doutb(w_n1895_0[1]),.doutc(w_n1895_0[2]),.din(n1895));
	jspl3 jspl3_w_n1902_0(.douta(w_n1902_0[0]),.doutb(w_n1902_0[1]),.doutc(w_n1902_0[2]),.din(n1902));
	jspl jspl_w_n1903_0(.douta(w_n1903_0[0]),.doutb(w_n1903_0[1]),.din(n1903));
	jspl jspl_w_n1904_0(.douta(w_n1904_0[0]),.doutb(w_n1904_0[1]),.din(n1904));
	jspl3 jspl3_w_n1908_0(.douta(w_n1908_0[0]),.doutb(w_n1908_0[1]),.doutc(w_n1908_0[2]),.din(n1908));
	jspl jspl_w_n1910_0(.douta(w_n1910_0[0]),.doutb(w_n1910_0[1]),.din(n1910));
	jspl jspl_w_n1921_0(.douta(w_n1921_0[0]),.doutb(w_n1921_0[1]),.din(n1921));
	jspl jspl_w_n1922_0(.douta(w_n1922_0[0]),.doutb(w_n1922_0[1]),.din(n1922));
	jspl jspl_w_n1930_0(.douta(w_n1930_0[0]),.doutb(w_n1930_0[1]),.din(n1930));
	jspl jspl_w_n1933_0(.douta(w_n1933_0[0]),.doutb(w_n1933_0[1]),.din(n1933));
	jspl jspl_w_n1938_0(.douta(w_n1938_0[0]),.doutb(w_n1938_0[1]),.din(n1938));
	jspl jspl_w_n1939_0(.douta(w_n1939_0[0]),.doutb(w_n1939_0[1]),.din(n1939));
	jspl jspl_w_n1940_0(.douta(w_n1940_0[0]),.doutb(w_n1940_0[1]),.din(n1940));
	jspl jspl_w_n1950_0(.douta(w_n1950_0[0]),.doutb(w_n1950_0[1]),.din(n1950));
	jspl jspl_w_n1953_0(.douta(w_n1953_0[0]),.doutb(w_n1953_0[1]),.din(n1953));
	jspl jspl_w_n1954_0(.douta(w_n1954_0[0]),.doutb(w_n1954_0[1]),.din(n1954));
	jspl3 jspl3_w_n1955_0(.douta(w_n1955_0[0]),.doutb(w_n1955_0[1]),.doutc(w_n1955_0[2]),.din(n1955));
	jspl3 jspl3_w_n1956_0(.douta(w_n1956_0[0]),.doutb(w_n1956_0[1]),.doutc(w_n1956_0[2]),.din(n1956));
	jspl3 jspl3_w_n1956_1(.douta(w_n1956_1[0]),.doutb(w_n1956_1[1]),.doutc(w_n1956_1[2]),.din(w_n1956_0[0]));
	jspl3 jspl3_w_n1956_2(.douta(w_n1956_2[0]),.doutb(w_n1956_2[1]),.doutc(w_n1956_2[2]),.din(w_n1956_0[1]));
	jspl3 jspl3_w_n1956_3(.douta(w_n1956_3[0]),.doutb(w_n1956_3[1]),.doutc(w_n1956_3[2]),.din(w_n1956_0[2]));
	jspl3 jspl3_w_n1956_4(.douta(w_n1956_4[0]),.doutb(w_n1956_4[1]),.doutc(w_n1956_4[2]),.din(w_n1956_1[0]));
	jspl3 jspl3_w_n1956_5(.douta(w_n1956_5[0]),.doutb(w_n1956_5[1]),.doutc(w_n1956_5[2]),.din(w_n1956_1[1]));
	jspl3 jspl3_w_n1956_6(.douta(w_n1956_6[0]),.doutb(w_n1956_6[1]),.doutc(w_n1956_6[2]),.din(w_n1956_1[2]));
	jspl jspl_w_n1956_7(.douta(w_n1956_7[0]),.doutb(w_n1956_7[1]),.din(w_n1956_2[0]));
	jspl3 jspl3_w_n1957_0(.douta(w_n1957_0[0]),.doutb(w_n1957_0[1]),.doutc(w_n1957_0[2]),.din(n1957));
	jspl3 jspl3_w_n1958_0(.douta(w_n1958_0[0]),.doutb(w_n1958_0[1]),.doutc(w_n1958_0[2]),.din(n1958));
	jspl jspl_w_n1958_1(.douta(w_n1958_1[0]),.doutb(w_n1958_1[1]),.din(w_n1958_0[0]));
	jspl3 jspl3_w_n1959_0(.douta(w_n1959_0[0]),.doutb(w_n1959_0[1]),.doutc(w_n1959_0[2]),.din(n1959));
	jspl3 jspl3_w_n1960_0(.douta(w_n1960_0[0]),.doutb(w_n1960_0[1]),.doutc(w_n1960_0[2]),.din(n1960));
	jspl3 jspl3_w_n1961_0(.douta(w_n1961_0[0]),.doutb(w_n1961_0[1]),.doutc(w_n1961_0[2]),.din(n1961));
	jspl jspl_w_n1962_0(.douta(w_n1962_0[0]),.doutb(w_n1962_0[1]),.din(n1962));
	jspl jspl_w_n1965_0(.douta(w_n1965_0[0]),.doutb(w_n1965_0[1]),.din(n1965));
	jspl jspl_w_n1970_0(.douta(w_n1970_0[0]),.doutb(w_n1970_0[1]),.din(n1970));
	jspl jspl_w_n1974_0(.douta(w_n1974_0[0]),.doutb(w_n1974_0[1]),.din(n1974));
	jspl jspl_w_n1979_0(.douta(w_n1979_0[0]),.doutb(w_n1979_0[1]),.din(n1979));
	jspl jspl_w_n1984_0(.douta(w_n1984_0[0]),.doutb(w_n1984_0[1]),.din(n1984));
	jspl3 jspl3_w_n1987_0(.douta(w_n1987_0[0]),.doutb(w_n1987_0[1]),.doutc(w_n1987_0[2]),.din(n1987));
	jspl3 jspl3_w_n1993_0(.douta(w_n1993_0[0]),.doutb(w_n1993_0[1]),.doutc(w_n1993_0[2]),.din(n1993));
	jspl jspl_w_n1994_0(.douta(w_n1994_0[0]),.doutb(w_n1994_0[1]),.din(n1994));
	jspl jspl_w_n1996_0(.douta(w_n1996_0[0]),.doutb(w_n1996_0[1]),.din(n1996));
	jspl jspl_w_n1999_0(.douta(w_n1999_0[0]),.doutb(w_n1999_0[1]),.din(n1999));
	jspl jspl_w_n2002_0(.douta(w_n2002_0[0]),.doutb(w_n2002_0[1]),.din(n2002));
	jspl jspl_w_n2014_0(.douta(w_n2014_0[0]),.doutb(w_n2014_0[1]),.din(n2014));
	jspl jspl_w_n2023_0(.douta(w_n2023_0[0]),.doutb(w_n2023_0[1]),.din(n2023));
	jspl jspl_w_n2026_0(.douta(w_n2026_0[0]),.doutb(w_n2026_0[1]),.din(n2026));
	jspl jspl_w_n2029_0(.douta(w_n2029_0[0]),.doutb(w_n2029_0[1]),.din(n2029));
	jspl jspl_w_n2037_0(.douta(w_n2037_0[0]),.doutb(w_n2037_0[1]),.din(n2037));
	jspl jspl_w_n2040_0(.douta(w_n2040_0[0]),.doutb(w_n2040_0[1]),.din(n2040));
	jspl jspl_w_n2041_0(.douta(w_n2041_0[0]),.doutb(w_n2041_0[1]),.din(n2041));
	jspl jspl_w_n2044_0(.douta(w_n2044_0[0]),.doutb(w_n2044_0[1]),.din(n2044));
	jspl jspl_w_n2045_0(.douta(w_n2045_0[0]),.doutb(w_n2045_0[1]),.din(n2045));
	jspl jspl_w_n2046_0(.douta(w_n2046_0[0]),.doutb(w_n2046_0[1]),.din(n2046));
	jspl jspl_w_n2049_0(.douta(w_n2049_0[0]),.doutb(w_n2049_0[1]),.din(n2049));
	jspl3 jspl3_w_n2051_0(.douta(w_n2051_0[0]),.doutb(w_n2051_0[1]),.doutc(w_n2051_0[2]),.din(n2051));
	jspl3 jspl3_w_n2051_1(.douta(w_n2051_1[0]),.doutb(w_n2051_1[1]),.doutc(w_n2051_1[2]),.din(w_n2051_0[0]));
	jspl3 jspl3_w_n2051_2(.douta(w_n2051_2[0]),.doutb(w_n2051_2[1]),.doutc(w_n2051_2[2]),.din(w_n2051_0[1]));
	jspl3 jspl3_w_n2051_3(.douta(w_n2051_3[0]),.doutb(w_n2051_3[1]),.doutc(w_n2051_3[2]),.din(w_n2051_0[2]));
	jspl3 jspl3_w_n2051_4(.douta(w_n2051_4[0]),.doutb(w_n2051_4[1]),.doutc(w_n2051_4[2]),.din(w_n2051_1[0]));
	jspl3 jspl3_w_n2051_5(.douta(w_n2051_5[0]),.doutb(w_n2051_5[1]),.doutc(w_n2051_5[2]),.din(w_n2051_1[1]));
	jspl3 jspl3_w_n2051_6(.douta(w_n2051_6[0]),.doutb(w_n2051_6[1]),.doutc(w_n2051_6[2]),.din(w_n2051_1[2]));
	jspl3 jspl3_w_n2051_7(.douta(w_n2051_7[0]),.doutb(w_n2051_7[1]),.doutc(w_n2051_7[2]),.din(w_n2051_2[0]));
	jspl jspl_w_n2051_8(.douta(w_n2051_8[0]),.doutb(w_n2051_8[1]),.din(w_n2051_2[1]));
	jspl jspl_w_n2058_0(.douta(w_n2058_0[0]),.doutb(w_n2058_0[1]),.din(n2058));
	jspl jspl_w_n2059_0(.douta(w_n2059_0[0]),.doutb(w_n2059_0[1]),.din(n2059));
	jspl jspl_w_n2060_0(.douta(w_n2060_0[0]),.doutb(w_n2060_0[1]),.din(n2060));
	jspl jspl_w_n2061_0(.douta(w_n2061_0[0]),.doutb(w_n2061_0[1]),.din(n2061));
	jspl jspl_w_n2062_0(.douta(w_n2062_0[0]),.doutb(w_n2062_0[1]),.din(n2062));
	jspl jspl_w_n2070_0(.douta(w_n2070_0[0]),.doutb(w_n2070_0[1]),.din(n2070));
	jspl jspl_w_n2078_0(.douta(w_n2078_0[0]),.doutb(w_n2078_0[1]),.din(n2078));
	jspl jspl_w_n2086_0(.douta(w_n2086_0[0]),.doutb(w_n2086_0[1]),.din(n2086));
	jspl jspl_w_n2087_0(.douta(w_n2087_0[0]),.doutb(w_n2087_0[1]),.din(n2087));
	jspl jspl_w_n2088_0(.douta(w_n2088_0[0]),.doutb(w_n2088_0[1]),.din(n2088));
	jspl jspl_w_n2089_0(.douta(w_n2089_0[0]),.doutb(w_n2089_0[1]),.din(n2089));
	jspl jspl_w_n2090_0(.douta(w_n2090_0[0]),.doutb(w_n2090_0[1]),.din(n2090));
	jspl3 jspl3_w_n2091_0(.douta(w_n2091_0[0]),.doutb(w_n2091_0[1]),.doutc(w_n2091_0[2]),.din(n2091));
	jspl jspl_w_n2091_1(.douta(w_n2091_1[0]),.doutb(w_n2091_1[1]),.din(w_n2091_0[0]));
	jspl3 jspl3_w_n2092_0(.douta(w_n2092_0[0]),.doutb(w_n2092_0[1]),.doutc(w_n2092_0[2]),.din(n2092));
	jspl jspl_w_n2093_0(.douta(w_n2093_0[0]),.doutb(w_n2093_0[1]),.din(n2093));
	jspl3 jspl3_w_n2094_0(.douta(w_n2094_0[0]),.doutb(w_n2094_0[1]),.doutc(w_n2094_0[2]),.din(n2094));
	jspl3 jspl3_w_n2094_1(.douta(w_n2094_1[0]),.doutb(w_n2094_1[1]),.doutc(w_n2094_1[2]),.din(w_n2094_0[0]));
	jspl3 jspl3_w_n2094_2(.douta(w_n2094_2[0]),.doutb(w_n2094_2[1]),.doutc(w_n2094_2[2]),.din(w_n2094_0[1]));
	jspl3 jspl3_w_n2094_3(.douta(w_n2094_3[0]),.doutb(w_n2094_3[1]),.doutc(w_n2094_3[2]),.din(w_n2094_0[2]));
	jspl3 jspl3_w_n2094_4(.douta(w_n2094_4[0]),.doutb(w_n2094_4[1]),.doutc(w_n2094_4[2]),.din(w_n2094_1[0]));
	jspl3 jspl3_w_n2094_5(.douta(w_n2094_5[0]),.doutb(w_n2094_5[1]),.doutc(w_n2094_5[2]),.din(w_n2094_1[1]));
	jspl3 jspl3_w_n2094_6(.douta(w_n2094_6[0]),.doutb(w_n2094_6[1]),.doutc(w_n2094_6[2]),.din(w_n2094_1[2]));
	jspl jspl_w_n2095_0(.douta(w_n2095_0[0]),.doutb(w_n2095_0[1]),.din(n2095));
	jspl3 jspl3_w_n2096_0(.douta(w_n2096_0[0]),.doutb(w_n2096_0[1]),.doutc(w_n2096_0[2]),.din(n2096));
	jspl jspl_w_n2096_1(.douta(w_n2096_1[0]),.doutb(w_n2096_1[1]),.din(w_n2096_0[0]));
	jspl3 jspl3_w_n2097_0(.douta(w_n2097_0[0]),.doutb(w_n2097_0[1]),.doutc(w_n2097_0[2]),.din(n2097));
	jspl3 jspl3_w_n2098_0(.douta(w_n2098_0[0]),.doutb(w_n2098_0[1]),.doutc(w_n2098_0[2]),.din(n2098));
	jspl jspl_w_n2099_0(.douta(w_n2099_0[0]),.doutb(w_n2099_0[1]),.din(n2099));
	jspl jspl_w_n2100_0(.douta(w_n2100_0[0]),.doutb(w_n2100_0[1]),.din(n2100));
	jspl3 jspl3_w_n2101_0(.douta(w_n2101_0[0]),.doutb(w_n2101_0[1]),.doutc(w_n2101_0[2]),.din(n2101));
	jspl jspl_w_n2101_1(.douta(w_n2101_1[0]),.doutb(w_n2101_1[1]),.din(w_n2101_0[0]));
	jspl3 jspl3_w_n2103_0(.douta(w_n2103_0[0]),.doutb(w_n2103_0[1]),.doutc(w_n2103_0[2]),.din(n2103));
	jspl jspl_w_n2105_0(.douta(w_n2105_0[0]),.doutb(w_n2105_0[1]),.din(n2105));
	jspl3 jspl3_w_n2107_0(.douta(w_n2107_0[0]),.doutb(w_n2107_0[1]),.doutc(w_n2107_0[2]),.din(n2107));
	jspl jspl_w_n2110_0(.douta(w_n2110_0[0]),.doutb(w_n2110_0[1]),.din(n2110));
	jspl3 jspl3_w_n2112_0(.douta(w_n2112_0[0]),.doutb(w_n2112_0[1]),.doutc(w_n2112_0[2]),.din(n2112));
	jspl jspl_w_n2112_1(.douta(w_n2112_1[0]),.doutb(w_n2112_1[1]),.din(w_n2112_0[0]));
	jspl jspl_w_n2115_0(.douta(w_n2115_0[0]),.doutb(w_n2115_0[1]),.din(n2115));
	jspl3 jspl3_w_n2116_0(.douta(w_n2116_0[0]),.doutb(w_n2116_0[1]),.doutc(w_n2116_0[2]),.din(n2116));
	jspl3 jspl3_w_n2116_1(.douta(w_n2116_1[0]),.doutb(w_n2116_1[1]),.doutc(w_n2116_1[2]),.din(w_n2116_0[0]));
	jspl3 jspl3_w_n2116_2(.douta(w_n2116_2[0]),.doutb(w_n2116_2[1]),.doutc(w_n2116_2[2]),.din(w_n2116_0[1]));
	jspl jspl_w_n2120_0(.douta(w_n2120_0[0]),.doutb(w_n2120_0[1]),.din(n2120));
	jspl jspl_w_n2126_0(.douta(w_n2126_0[0]),.doutb(w_n2126_0[1]),.din(n2126));
	jspl3 jspl3_w_n2127_0(.douta(w_n2127_0[0]),.doutb(w_n2127_0[1]),.doutc(w_n2127_0[2]),.din(n2127));
	jspl jspl_w_n2127_1(.douta(w_n2127_1[0]),.doutb(w_n2127_1[1]),.din(w_n2127_0[0]));
	jspl jspl_w_n2130_0(.douta(w_n2130_0[0]),.doutb(w_n2130_0[1]),.din(n2130));
	jspl3 jspl3_w_n2134_0(.douta(w_n2134_0[0]),.doutb(w_n2134_0[1]),.doutc(w_n2134_0[2]),.din(n2134));
	jspl3 jspl3_w_n2135_0(.douta(w_n2135_0[0]),.doutb(w_n2135_0[1]),.doutc(w_n2135_0[2]),.din(n2135));
	jspl3 jspl3_w_n2142_0(.douta(w_n2142_0[0]),.doutb(w_n2142_0[1]),.doutc(w_n2142_0[2]),.din(n2142));
	jspl3 jspl3_w_n2146_0(.douta(w_n2146_0[0]),.doutb(w_n2146_0[1]),.doutc(w_n2146_0[2]),.din(n2146));
	jspl jspl_w_n2147_0(.douta(w_n2147_0[0]),.doutb(w_n2147_0[1]),.din(n2147));
	jspl jspl_w_n2149_0(.douta(w_n2149_0[0]),.doutb(w_n2149_0[1]),.din(n2149));
	jspl jspl_w_n2154_0(.douta(w_n2154_0[0]),.doutb(w_n2154_0[1]),.din(n2154));
	jspl3 jspl3_w_n2155_0(.douta(w_n2155_0[0]),.doutb(w_n2155_0[1]),.doutc(w_n2155_0[2]),.din(n2155));
	jspl jspl_w_n2155_1(.douta(w_n2155_1[0]),.doutb(w_n2155_1[1]),.din(w_n2155_0[0]));
	jspl3 jspl3_w_n2166_0(.douta(w_n2166_0[0]),.doutb(w_n2166_0[1]),.doutc(w_n2166_0[2]),.din(n2166));
	jspl jspl_w_n2167_0(.douta(w_n2167_0[0]),.doutb(w_n2167_0[1]),.din(n2167));
	jspl jspl_w_n2169_0(.douta(w_n2169_0[0]),.doutb(w_n2169_0[1]),.din(n2169));
	jspl jspl_w_n2172_0(.douta(w_n2172_0[0]),.doutb(w_n2172_0[1]),.din(n2172));
	jspl jspl_w_n2175_0(.douta(w_n2175_0[0]),.doutb(w_n2175_0[1]),.din(n2175));
	jspl jspl_w_n2183_0(.douta(w_n2183_0[0]),.doutb(w_n2183_0[1]),.din(n2183));
	jspl jspl_w_n2186_0(.douta(w_n2186_0[0]),.doutb(w_n2186_0[1]),.din(n2186));
	jspl jspl_w_n2187_0(.douta(w_n2187_0[0]),.doutb(w_n2187_0[1]),.din(n2187));
	jspl jspl_w_n2190_0(.douta(w_n2190_0[0]),.doutb(w_n2190_0[1]),.din(n2190));
	jspl jspl_w_n2191_0(.douta(w_n2191_0[0]),.doutb(w_n2191_0[1]),.din(n2191));
	jspl jspl_w_n2192_0(.douta(w_n2192_0[0]),.doutb(w_n2192_0[1]),.din(n2192));
	jspl jspl_w_n2195_0(.douta(w_n2195_0[0]),.doutb(w_n2195_0[1]),.din(n2195));
	jspl jspl_w_n2203_0(.douta(w_n2203_0[0]),.doutb(w_n2203_0[1]),.din(n2203));
	jspl jspl_w_n2211_0(.douta(w_n2211_0[0]),.doutb(w_n2211_0[1]),.din(n2211));
	jspl jspl_w_n2219_0(.douta(w_n2219_0[0]),.doutb(w_n2219_0[1]),.din(n2219));
	jspl jspl_w_n2220_0(.douta(w_n2220_0[0]),.doutb(w_n2220_0[1]),.din(n2220));
	jspl jspl_w_n2221_0(.douta(w_n2221_0[0]),.doutb(w_n2221_0[1]),.din(n2221));
	jspl jspl_w_n2226_0(.douta(w_n2226_0[0]),.doutb(w_n2226_0[1]),.din(n2226));
	jspl jspl_w_n2227_0(.douta(w_n2227_0[0]),.doutb(w_n2227_0[1]),.din(n2227));
	jspl jspl_w_n2228_0(.douta(w_n2228_0[0]),.doutb(w_n2228_0[1]),.din(n2228));
	jspl jspl_w_n2229_0(.douta(w_n2229_0[0]),.doutb(w_n2229_0[1]),.din(n2229));
	jspl jspl_w_n2230_0(.douta(w_n2230_0[0]),.doutb(w_n2230_0[1]),.din(n2230));
	jspl jspl_w_n2231_0(.douta(w_n2231_0[0]),.doutb(w_n2231_0[1]),.din(n2231));
	jspl jspl_w_n2232_0(.douta(w_n2232_0[0]),.doutb(w_n2232_0[1]),.din(n2232));
	jspl3 jspl3_w_n2233_0(.douta(w_n2233_0[0]),.doutb(w_n2233_0[1]),.doutc(w_n2233_0[2]),.din(n2233));
	jspl jspl_w_n2233_1(.douta(w_n2233_1[0]),.doutb(w_n2233_1[1]),.din(w_n2233_0[0]));
	jspl3 jspl3_w_n2234_0(.douta(w_n2234_0[0]),.doutb(w_n2234_0[1]),.doutc(w_n2234_0[2]),.din(n2234));
	jspl3 jspl3_w_n2235_0(.douta(w_n2235_0[0]),.doutb(w_n2235_0[1]),.doutc(w_n2235_0[2]),.din(n2235));
	jspl3 jspl3_w_n2236_0(.douta(w_n2236_0[0]),.doutb(w_n2236_0[1]),.doutc(w_n2236_0[2]),.din(n2236));
	jspl3 jspl3_w_n2236_1(.douta(w_n2236_1[0]),.doutb(w_n2236_1[1]),.doutc(w_n2236_1[2]),.din(w_n2236_0[0]));
	jspl3 jspl3_w_n2236_2(.douta(w_n2236_2[0]),.doutb(w_n2236_2[1]),.doutc(w_n2236_2[2]),.din(w_n2236_0[1]));
	jspl3 jspl3_w_n2236_3(.douta(w_n2236_3[0]),.doutb(w_n2236_3[1]),.doutc(w_n2236_3[2]),.din(w_n2236_0[2]));
	jspl3 jspl3_w_n2236_4(.douta(w_n2236_4[0]),.doutb(w_n2236_4[1]),.doutc(w_n2236_4[2]),.din(w_n2236_1[0]));
	jspl jspl_w_n2236_5(.douta(w_n2236_5[0]),.doutb(w_n2236_5[1]),.din(w_n2236_1[1]));
	jspl3 jspl3_w_n2238_0(.douta(w_n2238_0[0]),.doutb(w_n2238_0[1]),.doutc(w_n2238_0[2]),.din(n2238));
	jspl jspl_w_n2238_1(.douta(w_n2238_1[0]),.doutb(w_n2238_1[1]),.din(w_n2238_0[0]));
	jspl3 jspl3_w_n2244_0(.douta(w_n2244_0[0]),.doutb(w_n2244_0[1]),.doutc(w_n2244_0[2]),.din(n2244));
	jspl jspl_w_n2248_0(.douta(w_n2248_0[0]),.doutb(w_n2248_0[1]),.din(n2248));
	jspl jspl_w_n2249_0(.douta(w_n2249_0[0]),.doutb(w_n2249_0[1]),.din(n2249));
	jspl jspl_w_n2251_0(.douta(w_n2251_0[0]),.doutb(w_n2251_0[1]),.din(n2251));
	jspl3 jspl3_w_n2252_0(.douta(w_n2252_0[0]),.doutb(w_n2252_0[1]),.doutc(w_n2252_0[2]),.din(n2252));
	jspl3 jspl3_w_n2252_1(.douta(w_n2252_1[0]),.doutb(w_n2252_1[1]),.doutc(w_n2252_1[2]),.din(w_n2252_0[0]));
	jspl3 jspl3_w_n2252_2(.douta(w_n2252_2[0]),.doutb(w_n2252_2[1]),.doutc(w_n2252_2[2]),.din(w_n2252_0[1]));
	jspl3 jspl3_w_n2252_3(.douta(w_n2252_3[0]),.doutb(w_n2252_3[1]),.doutc(w_n2252_3[2]),.din(w_n2252_0[2]));
	jspl3 jspl3_w_n2252_4(.douta(w_n2252_4[0]),.doutb(w_n2252_4[1]),.doutc(w_n2252_4[2]),.din(w_n2252_1[0]));
	jspl3 jspl3_w_n2252_5(.douta(w_n2252_5[0]),.doutb(w_n2252_5[1]),.doutc(w_n2252_5[2]),.din(w_n2252_1[1]));
	jspl3 jspl3_w_n2252_6(.douta(w_n2252_6[0]),.doutb(w_n2252_6[1]),.doutc(w_n2252_6[2]),.din(w_n2252_1[2]));
	jspl3 jspl3_w_n2252_7(.douta(w_n2252_7[0]),.doutb(w_n2252_7[1]),.doutc(w_n2252_7[2]),.din(w_n2252_2[0]));
	jspl jspl_w_n2255_0(.douta(w_n2255_0[0]),.doutb(w_n2255_0[1]),.din(n2255));
	jspl3 jspl3_w_n2256_0(.douta(w_n2256_0[0]),.doutb(w_n2256_0[1]),.doutc(w_n2256_0[2]),.din(n2256));
	jspl3 jspl3_w_n2256_1(.douta(w_n2256_1[0]),.doutb(w_n2256_1[1]),.doutc(w_n2256_1[2]),.din(w_n2256_0[0]));
	jspl3 jspl3_w_n2256_2(.douta(w_n2256_2[0]),.doutb(w_n2256_2[1]),.doutc(w_n2256_2[2]),.din(w_n2256_0[1]));
	jspl3 jspl3_w_n2256_3(.douta(w_n2256_3[0]),.doutb(w_n2256_3[1]),.doutc(w_n2256_3[2]),.din(w_n2256_0[2]));
	jspl3 jspl3_w_n2256_4(.douta(w_n2256_4[0]),.doutb(w_n2256_4[1]),.doutc(w_n2256_4[2]),.din(w_n2256_1[0]));
	jspl3 jspl3_w_n2256_5(.douta(w_n2256_5[0]),.doutb(w_n2256_5[1]),.doutc(w_n2256_5[2]),.din(w_n2256_1[1]));
	jspl jspl_w_n2258_0(.douta(w_n2258_0[0]),.doutb(w_n2258_0[1]),.din(n2258));
	jspl jspl_w_n2260_0(.douta(w_n2260_0[0]),.doutb(w_n2260_0[1]),.din(n2260));
	jspl jspl_w_n2263_0(.douta(w_n2263_0[0]),.doutb(w_n2263_0[1]),.din(n2263));
	jspl3 jspl3_w_n2277_0(.douta(w_n2277_0[0]),.doutb(w_n2277_0[1]),.doutc(w_n2277_0[2]),.din(n2277));
	jspl jspl_w_n2278_0(.douta(w_n2278_0[0]),.doutb(w_n2278_0[1]),.din(n2278));
	jspl jspl_w_n2280_0(.douta(w_n2280_0[0]),.doutb(w_n2280_0[1]),.din(n2280));
	jspl jspl_w_n2283_0(.douta(w_n2283_0[0]),.doutb(w_n2283_0[1]),.din(n2283));
	jspl jspl_w_n2286_0(.douta(w_n2286_0[0]),.doutb(w_n2286_0[1]),.din(n2286));
	jspl jspl_w_n2289_0(.douta(w_n2289_0[0]),.doutb(w_n2289_0[1]),.din(n2289));
	jspl jspl_w_n2297_0(.douta(w_n2297_0[0]),.doutb(w_n2297_0[1]),.din(n2297));
	jspl jspl_w_n2299_0(.douta(w_n2299_0[0]),.doutb(w_n2299_0[1]),.din(n2299));
	jspl jspl_w_n2301_0(.douta(w_n2301_0[0]),.doutb(w_n2301_0[1]),.din(n2301));
	jspl jspl_w_n2302_0(.douta(w_n2302_0[0]),.doutb(w_n2302_0[1]),.din(n2302));
	jspl jspl_w_n2305_0(.douta(w_n2305_0[0]),.doutb(w_n2305_0[1]),.din(n2305));
	jspl jspl_w_n2306_0(.douta(w_n2306_0[0]),.doutb(w_n2306_0[1]),.din(n2306));
	jspl jspl_w_n2309_0(.douta(w_n2309_0[0]),.doutb(w_n2309_0[1]),.din(n2309));
	jspl jspl_w_n2310_0(.douta(w_n2310_0[0]),.doutb(w_n2310_0[1]),.din(n2310));
	jspl jspl_w_n2311_0(.douta(w_n2311_0[0]),.doutb(w_n2311_0[1]),.din(n2311));
	jspl jspl_w_n2312_0(.douta(w_n2312_0[0]),.doutb(w_n2312_0[1]),.din(n2312));
	jspl jspl_w_n2315_0(.douta(w_n2315_0[0]),.doutb(w_n2315_0[1]),.din(n2315));
	jspl jspl_w_n2318_0(.douta(w_n2318_0[0]),.doutb(w_n2318_0[1]),.din(n2318));
	jspl jspl_w_n2326_0(.douta(w_n2326_0[0]),.doutb(w_n2326_0[1]),.din(n2326));
	jspl jspl_w_n2334_0(.douta(w_n2334_0[0]),.doutb(w_n2334_0[1]),.din(n2334));
	jspl jspl_w_n2342_0(.douta(w_n2342_0[0]),.doutb(w_n2342_0[1]),.din(n2342));
	jspl jspl_w_n2343_0(.douta(w_n2343_0[0]),.doutb(w_n2343_0[1]),.din(n2343));
	jspl jspl_w_n2344_0(.douta(w_n2344_0[0]),.doutb(w_n2344_0[1]),.din(n2344));
	jspl jspl_w_n2345_0(.douta(w_n2345_0[0]),.doutb(w_n2345_0[1]),.din(n2345));
	jspl jspl_w_n2346_0(.douta(w_n2346_0[0]),.doutb(w_n2346_0[1]),.din(n2346));
	jspl jspl_w_n2347_0(.douta(w_n2347_0[0]),.doutb(w_n2347_0[1]),.din(n2347));
	jspl3 jspl3_w_n2348_0(.douta(w_n2348_0[0]),.doutb(w_n2348_0[1]),.doutc(w_n2348_0[2]),.din(n2348));
	jspl jspl_w_n2348_1(.douta(w_n2348_1[0]),.doutb(w_n2348_1[1]),.din(w_n2348_0[0]));
	jspl3 jspl3_w_n2349_0(.douta(w_n2349_0[0]),.doutb(w_n2349_0[1]),.doutc(w_n2349_0[2]),.din(n2349));
	jspl3 jspl3_w_n2350_0(.douta(w_n2350_0[0]),.doutb(w_n2350_0[1]),.doutc(w_n2350_0[2]),.din(n2350));
	jspl3 jspl3_w_n2351_0(.douta(w_n2351_0[0]),.doutb(w_n2351_0[1]),.doutc(w_n2351_0[2]),.din(n2351));
	jspl3 jspl3_w_n2351_1(.douta(w_n2351_1[0]),.doutb(w_n2351_1[1]),.doutc(w_n2351_1[2]),.din(w_n2351_0[0]));
	jspl3 jspl3_w_n2351_2(.douta(w_n2351_2[0]),.doutb(w_n2351_2[1]),.doutc(w_n2351_2[2]),.din(w_n2351_0[1]));
	jspl3 jspl3_w_n2351_3(.douta(w_n2351_3[0]),.doutb(w_n2351_3[1]),.doutc(w_n2351_3[2]),.din(w_n2351_0[2]));
	jspl3 jspl3_w_n2351_4(.douta(w_n2351_4[0]),.doutb(w_n2351_4[1]),.doutc(w_n2351_4[2]),.din(w_n2351_1[0]));
	jspl3 jspl3_w_n2351_5(.douta(w_n2351_5[0]),.doutb(w_n2351_5[1]),.doutc(w_n2351_5[2]),.din(w_n2351_1[1]));
	jspl3 jspl3_w_n2351_6(.douta(w_n2351_6[0]),.doutb(w_n2351_6[1]),.doutc(w_n2351_6[2]),.din(w_n2351_1[2]));
	jspl3 jspl3_w_n2351_7(.douta(w_n2351_7[0]),.doutb(w_n2351_7[1]),.doutc(w_n2351_7[2]),.din(w_n2351_2[0]));
	jspl jspl_w_n2351_8(.douta(w_n2351_8[0]),.doutb(w_n2351_8[1]),.din(w_n2351_2[1]));
	jspl3 jspl3_w_n2352_0(.douta(w_n2352_0[0]),.doutb(w_n2352_0[1]),.doutc(w_n2352_0[2]),.din(n2352));
	jspl3 jspl3_w_n2353_0(.douta(w_n2353_0[0]),.doutb(w_n2353_0[1]),.doutc(w_n2353_0[2]),.din(n2353));
	jspl3 jspl3_w_n2353_1(.douta(w_n2353_1[0]),.doutb(w_n2353_1[1]),.doutc(w_n2353_1[2]),.din(w_n2353_0[0]));
	jspl3 jspl3_w_n2355_0(.douta(w_n2355_0[0]),.doutb(w_n2355_0[1]),.doutc(w_n2355_0[2]),.din(n2355));
	jspl3 jspl3_w_n2355_1(.douta(w_n2355_1[0]),.doutb(w_n2355_1[1]),.doutc(w_n2355_1[2]),.din(w_n2355_0[0]));
	jspl3 jspl3_w_n2355_2(.douta(w_n2355_2[0]),.doutb(w_n2355_2[1]),.doutc(w_n2355_2[2]),.din(w_n2355_0[1]));
	jspl3 jspl3_w_n2355_3(.douta(w_n2355_3[0]),.doutb(w_n2355_3[1]),.doutc(w_n2355_3[2]),.din(w_n2355_0[2]));
	jspl3 jspl3_w_n2355_4(.douta(w_n2355_4[0]),.doutb(w_n2355_4[1]),.doutc(w_n2355_4[2]),.din(w_n2355_1[0]));
	jspl3 jspl3_w_n2355_5(.douta(w_n2355_5[0]),.doutb(w_n2355_5[1]),.doutc(w_n2355_5[2]),.din(w_n2355_1[1]));
	jspl3 jspl3_w_n2355_6(.douta(w_n2355_6[0]),.doutb(w_n2355_6[1]),.doutc(w_n2355_6[2]),.din(w_n2355_1[2]));
	jspl jspl_w_n2355_7(.douta(w_n2355_7[0]),.doutb(w_n2355_7[1]),.din(w_n2355_2[0]));
	jspl3 jspl3_w_n2357_0(.douta(w_n2357_0[0]),.doutb(w_n2357_0[1]),.doutc(w_n2357_0[2]),.din(n2357));
	jspl3 jspl3_w_n2357_1(.douta(w_n2357_1[0]),.doutb(w_n2357_1[1]),.doutc(w_n2357_1[2]),.din(w_n2357_0[0]));
	jspl3 jspl3_w_n2357_2(.douta(w_n2357_2[0]),.doutb(w_n2357_2[1]),.doutc(w_n2357_2[2]),.din(w_n2357_0[1]));
	jspl3 jspl3_w_n2357_3(.douta(w_n2357_3[0]),.doutb(w_n2357_3[1]),.doutc(w_n2357_3[2]),.din(w_n2357_0[2]));
	jspl3 jspl3_w_n2357_4(.douta(w_n2357_4[0]),.doutb(w_n2357_4[1]),.doutc(w_n2357_4[2]),.din(w_n2357_1[0]));
	jspl3 jspl3_w_n2357_5(.douta(w_n2357_5[0]),.doutb(w_n2357_5[1]),.doutc(w_n2357_5[2]),.din(w_n2357_1[1]));
	jspl3 jspl3_w_n2357_6(.douta(w_n2357_6[0]),.doutb(w_n2357_6[1]),.doutc(w_n2357_6[2]),.din(w_n2357_1[2]));
	jspl3 jspl3_w_n2357_7(.douta(w_n2357_7[0]),.doutb(w_n2357_7[1]),.doutc(w_n2357_7[2]),.din(w_n2357_2[0]));
	jspl3 jspl3_w_n2359_0(.douta(w_n2359_0[0]),.doutb(w_n2359_0[1]),.doutc(w_n2359_0[2]),.din(n2359));
	jspl3 jspl3_w_n2359_1(.douta(w_n2359_1[0]),.doutb(w_n2359_1[1]),.doutc(w_n2359_1[2]),.din(w_n2359_0[0]));
	jspl3 jspl3_w_n2359_2(.douta(w_n2359_2[0]),.doutb(w_n2359_2[1]),.doutc(w_n2359_2[2]),.din(w_n2359_0[1]));
	jspl3 jspl3_w_n2359_3(.douta(w_n2359_3[0]),.doutb(w_n2359_3[1]),.doutc(w_n2359_3[2]),.din(w_n2359_0[2]));
	jspl3 jspl3_w_n2359_4(.douta(w_n2359_4[0]),.doutb(w_n2359_4[1]),.doutc(w_n2359_4[2]),.din(w_n2359_1[0]));
	jspl3 jspl3_w_n2359_5(.douta(w_n2359_5[0]),.doutb(w_n2359_5[1]),.doutc(w_n2359_5[2]),.din(w_n2359_1[1]));
	jspl3 jspl3_w_n2359_6(.douta(w_n2359_6[0]),.doutb(w_n2359_6[1]),.doutc(w_n2359_6[2]),.din(w_n2359_1[2]));
	jspl3 jspl3_w_n2359_7(.douta(w_n2359_7[0]),.doutb(w_n2359_7[1]),.doutc(w_n2359_7[2]),.din(w_n2359_2[0]));
	jspl jspl_w_n2364_0(.douta(w_n2364_0[0]),.doutb(w_n2364_0[1]),.din(n2364));
	jspl jspl_w_n2366_0(.douta(w_n2366_0[0]),.doutb(w_n2366_0[1]),.din(n2366));
	jspl jspl_w_n2370_0(.douta(w_n2370_0[0]),.doutb(w_n2370_0[1]),.din(n2370));
	jspl jspl_w_n2372_0(.douta(w_n2372_0[0]),.doutb(w_n2372_0[1]),.din(n2372));
	jspl jspl_w_n2375_0(.douta(w_n2375_0[0]),.doutb(w_n2375_0[1]),.din(n2375));
	jspl jspl_w_n2377_0(.douta(w_n2377_0[0]),.doutb(w_n2377_0[1]),.din(n2377));
	jspl jspl_w_n2384_0(.douta(w_n2384_0[0]),.doutb(w_n2384_0[1]),.din(n2384));
	jspl jspl_w_n2386_0(.douta(w_n2386_0[0]),.doutb(w_n2386_0[1]),.din(n2386));
	jspl jspl_w_n2394_0(.douta(w_n2394_0[0]),.doutb(w_n2394_0[1]),.din(n2394));
	jspl3 jspl3_w_n2395_0(.douta(w_n2395_0[0]),.doutb(w_n2395_0[1]),.doutc(w_n2395_0[2]),.din(n2395));
	jspl jspl_w_n2402_0(.douta(w_n2402_0[0]),.doutb(w_n2402_0[1]),.din(n2402));
	jspl jspl_w_n2409_0(.douta(w_n2409_0[0]),.doutb(w_n2409_0[1]),.din(n2409));
	jspl3 jspl3_w_n2412_0(.douta(w_n2412_0[0]),.doutb(w_n2412_0[1]),.doutc(w_n2412_0[2]),.din(n2412));
	jspl jspl_w_n2413_0(.douta(w_n2413_0[0]),.doutb(w_n2413_0[1]),.din(n2413));
	jspl jspl_w_n2415_0(.douta(w_n2415_0[0]),.doutb(w_n2415_0[1]),.din(n2415));
	jspl jspl_w_n2418_0(.douta(w_n2418_0[0]),.doutb(w_n2418_0[1]),.din(n2418));
	jspl jspl_w_n2421_0(.douta(w_n2421_0[0]),.doutb(w_n2421_0[1]),.din(n2421));
	jspl jspl_w_n2424_0(.douta(w_n2424_0[0]),.doutb(w_n2424_0[1]),.din(n2424));
	jspl jspl_w_n2425_0(.douta(w_n2425_0[0]),.doutb(w_n2425_0[1]),.din(n2425));
	jspl jspl_w_n2426_0(.douta(w_n2426_0[0]),.doutb(w_n2426_0[1]),.din(n2426));
	jspl jspl_w_n2434_0(.douta(w_n2434_0[0]),.doutb(w_n2434_0[1]),.din(n2434));
	jspl jspl_w_n2442_0(.douta(w_n2442_0[0]),.doutb(w_n2442_0[1]),.din(n2442));
	jspl jspl_w_n2443_0(.douta(w_n2443_0[0]),.doutb(w_n2443_0[1]),.din(n2443));
	jspl jspl_w_n2444_0(.douta(w_n2444_0[0]),.doutb(w_n2444_0[1]),.din(n2444));
	jspl jspl_w_n2447_0(.douta(w_n2447_0[0]),.doutb(w_n2447_0[1]),.din(n2447));
	jspl jspl_w_n2455_0(.douta(w_n2455_0[0]),.doutb(w_n2455_0[1]),.din(n2455));
	jspl3 jspl3_w_n2456_0(.douta(w_n2456_0[0]),.doutb(w_n2456_0[1]),.doutc(w_n2456_0[2]),.din(n2456));
	jspl jspl_w_n2457_0(.douta(w_n2457_0[0]),.doutb(w_n2457_0[1]),.din(n2457));
	jspl jspl_w_n2462_0(.douta(w_n2462_0[0]),.doutb(w_n2462_0[1]),.din(n2462));
	jspl jspl_w_n2463_0(.douta(w_n2463_0[0]),.doutb(w_n2463_0[1]),.din(n2463));
	jspl jspl_w_n2464_0(.douta(w_n2464_0[0]),.doutb(w_n2464_0[1]),.din(n2464));
	jspl jspl_w_n2465_0(.douta(w_n2465_0[0]),.doutb(w_n2465_0[1]),.din(n2465));
	jspl jspl_w_n2466_0(.douta(w_n2466_0[0]),.doutb(w_n2466_0[1]),.din(n2466));
	jspl jspl_w_n2467_0(.douta(w_n2467_0[0]),.doutb(w_n2467_0[1]),.din(n2467));
	jspl3 jspl3_w_n2468_0(.douta(w_n2468_0[0]),.doutb(w_n2468_0[1]),.doutc(w_n2468_0[2]),.din(n2468));
	jspl jspl_w_n2468_1(.douta(w_n2468_1[0]),.doutb(w_n2468_1[1]),.din(w_n2468_0[0]));
	jspl3 jspl3_w_n2469_0(.douta(w_n2469_0[0]),.doutb(w_n2469_0[1]),.doutc(w_n2469_0[2]),.din(n2469));
	jspl3 jspl3_w_n2470_0(.douta(w_n2470_0[0]),.doutb(w_n2470_0[1]),.doutc(w_n2470_0[2]),.din(n2470));
	jspl3 jspl3_w_n2471_0(.douta(w_n2471_0[0]),.doutb(w_n2471_0[1]),.doutc(w_n2471_0[2]),.din(n2471));
	jspl3 jspl3_w_n2471_1(.douta(w_n2471_1[0]),.doutb(w_n2471_1[1]),.doutc(w_n2471_1[2]),.din(w_n2471_0[0]));
	jspl3 jspl3_w_n2471_2(.douta(w_n2471_2[0]),.doutb(w_n2471_2[1]),.doutc(w_n2471_2[2]),.din(w_n2471_0[1]));
	jspl3 jspl3_w_n2471_3(.douta(w_n2471_3[0]),.doutb(w_n2471_3[1]),.doutc(w_n2471_3[2]),.din(w_n2471_0[2]));
	jspl3 jspl3_w_n2471_4(.douta(w_n2471_4[0]),.doutb(w_n2471_4[1]),.doutc(w_n2471_4[2]),.din(w_n2471_1[0]));
	jspl3 jspl3_w_n2471_5(.douta(w_n2471_5[0]),.doutb(w_n2471_5[1]),.doutc(w_n2471_5[2]),.din(w_n2471_1[1]));
	jspl3 jspl3_w_n2471_6(.douta(w_n2471_6[0]),.doutb(w_n2471_6[1]),.doutc(w_n2471_6[2]),.din(w_n2471_1[2]));
	jspl jspl_w_n2471_7(.douta(w_n2471_7[0]),.doutb(w_n2471_7[1]),.din(w_n2471_2[0]));
	jspl3 jspl3_w_n2472_0(.douta(w_n2472_0[0]),.doutb(w_n2472_0[1]),.doutc(w_n2472_0[2]),.din(n2472));
	jspl3 jspl3_w_n2473_0(.douta(w_n2473_0[0]),.doutb(w_n2473_0[1]),.doutc(w_n2473_0[2]),.din(n2473));
	jspl jspl_w_n2473_1(.douta(w_n2473_1[0]),.doutb(w_n2473_1[1]),.din(w_n2473_0[0]));
	jspl jspl_w_n2482_0(.douta(w_n2482_0[0]),.doutb(w_n2482_0[1]),.din(n2482));
	jspl3 jspl3_w_n2483_0(.douta(w_n2483_0[0]),.doutb(w_n2483_0[1]),.doutc(w_n2483_0[2]),.din(n2483));
	jspl jspl_w_n2483_1(.douta(w_n2483_1[0]),.doutb(w_n2483_1[1]),.din(w_n2483_0[0]));
	jspl3 jspl3_w_n2484_0(.douta(w_n2484_0[0]),.doutb(w_n2484_0[1]),.doutc(w_n2484_0[2]),.din(n2484));
	jspl3 jspl3_w_n2484_1(.douta(w_n2484_1[0]),.doutb(w_n2484_1[1]),.doutc(w_n2484_1[2]),.din(w_n2484_0[0]));
	jspl jspl_w_n2486_0(.douta(w_n2486_0[0]),.doutb(w_n2486_0[1]),.din(n2486));
	jspl3 jspl3_w_n2488_0(.douta(w_n2488_0[0]),.doutb(w_n2488_0[1]),.doutc(w_n2488_0[2]),.din(n2488));
	jspl3 jspl3_w_n2488_1(.douta(w_n2488_1[0]),.doutb(w_n2488_1[1]),.doutc(w_n2488_1[2]),.din(w_n2488_0[0]));
	jspl3 jspl3_w_n2488_2(.douta(w_n2488_2[0]),.doutb(w_n2488_2[1]),.doutc(w_n2488_2[2]),.din(w_n2488_0[1]));
	jspl3 jspl3_w_n2488_3(.douta(w_n2488_3[0]),.doutb(w_n2488_3[1]),.doutc(w_n2488_3[2]),.din(w_n2488_0[2]));
	jspl3 jspl3_w_n2491_0(.douta(w_n2491_0[0]),.doutb(w_n2491_0[1]),.doutc(w_n2491_0[2]),.din(n2491));
	jspl3 jspl3_w_n2491_1(.douta(w_n2491_1[0]),.doutb(w_n2491_1[1]),.doutc(w_n2491_1[2]),.din(w_n2491_0[0]));
	jspl3 jspl3_w_n2491_2(.douta(w_n2491_2[0]),.doutb(w_n2491_2[1]),.doutc(w_n2491_2[2]),.din(w_n2491_0[1]));
	jspl3 jspl3_w_n2491_3(.douta(w_n2491_3[0]),.doutb(w_n2491_3[1]),.doutc(w_n2491_3[2]),.din(w_n2491_0[2]));
	jspl jspl_w_n2494_0(.douta(w_n2494_0[0]),.doutb(w_n2494_0[1]),.din(n2494));
	jspl jspl_w_n2495_0(.douta(w_n2495_0[0]),.doutb(w_n2495_0[1]),.din(n2495));
	jspl jspl_w_n2497_0(.douta(w_n2497_0[0]),.doutb(w_n2497_0[1]),.din(n2497));
	jspl jspl_w_n2498_0(.douta(w_n2498_0[0]),.doutb(w_n2498_0[1]),.din(n2498));
	jspl jspl_w_n2500_0(.douta(w_n2500_0[0]),.doutb(w_n2500_0[1]),.din(n2500));
	jspl3 jspl3_w_n2501_0(.douta(w_n2501_0[0]),.doutb(w_n2501_0[1]),.doutc(w_n2501_0[2]),.din(n2501));
	jspl3 jspl3_w_n2502_0(.douta(w_n2502_0[0]),.doutb(w_n2502_0[1]),.doutc(w_n2502_0[2]),.din(n2502));
	jspl jspl_w_n2503_0(.douta(w_n2503_0[0]),.doutb(w_n2503_0[1]),.din(n2503));
	jspl jspl_w_n2504_0(.douta(w_n2504_0[0]),.doutb(w_n2504_0[1]),.din(n2504));
	jspl3 jspl3_w_n2505_0(.douta(w_n2505_0[0]),.doutb(w_n2505_0[1]),.doutc(w_n2505_0[2]),.din(n2505));
	jspl jspl_w_n2505_1(.douta(w_n2505_1[0]),.doutb(w_n2505_1[1]),.din(w_n2505_0[0]));
	jspl3 jspl3_w_n2506_0(.douta(w_n2506_0[0]),.doutb(w_n2506_0[1]),.doutc(w_n2506_0[2]),.din(n2506));
	jspl3 jspl3_w_n2506_1(.douta(w_n2506_1[0]),.doutb(w_n2506_1[1]),.doutc(w_n2506_1[2]),.din(w_n2506_0[0]));
	jspl3 jspl3_w_n2506_2(.douta(w_n2506_2[0]),.doutb(w_n2506_2[1]),.doutc(w_n2506_2[2]),.din(w_n2506_0[1]));
	jspl3 jspl3_w_n2506_3(.douta(w_n2506_3[0]),.doutb(w_n2506_3[1]),.doutc(w_n2506_3[2]),.din(w_n2506_0[2]));
	jspl3 jspl3_w_n2506_4(.douta(w_n2506_4[0]),.doutb(w_n2506_4[1]),.doutc(w_n2506_4[2]),.din(w_n2506_1[0]));
	jspl3 jspl3_w_n2506_5(.douta(w_n2506_5[0]),.doutb(w_n2506_5[1]),.doutc(w_n2506_5[2]),.din(w_n2506_1[1]));
	jspl3 jspl3_w_n2506_6(.douta(w_n2506_6[0]),.doutb(w_n2506_6[1]),.doutc(w_n2506_6[2]),.din(w_n2506_1[2]));
	jspl3 jspl3_w_n2506_7(.douta(w_n2506_7[0]),.doutb(w_n2506_7[1]),.doutc(w_n2506_7[2]),.din(w_n2506_2[0]));
	jspl jspl_w_n2508_0(.douta(w_n2508_0[0]),.doutb(w_n2508_0[1]),.din(n2508));
	jspl jspl_w_n2510_0(.douta(w_n2510_0[0]),.doutb(w_n2510_0[1]),.din(n2510));
	jspl3 jspl3_w_n2513_0(.douta(w_n2513_0[0]),.doutb(w_n2513_0[1]),.doutc(w_n2513_0[2]),.din(n2513));
	jspl jspl_w_n2513_1(.douta(w_n2513_1[0]),.doutb(w_n2513_1[1]),.din(w_n2513_0[0]));
	jspl3 jspl3_w_n2519_0(.douta(w_n2519_0[0]),.doutb(w_n2519_0[1]),.doutc(w_n2519_0[2]),.din(n2519));
	jspl jspl_w_n2520_0(.douta(w_n2520_0[0]),.doutb(w_n2520_0[1]),.din(n2520));
	jspl jspl_w_n2521_0(.douta(w_n2521_0[0]),.doutb(w_n2521_0[1]),.din(n2521));
	jspl jspl_w_n2528_0(.douta(w_n2528_0[0]),.doutb(w_n2528_0[1]),.din(n2528));
	jspl jspl_w_n2531_0(.douta(w_n2531_0[0]),.doutb(w_n2531_0[1]),.din(n2531));
	jspl jspl_w_n2534_0(.douta(w_n2534_0[0]),.doutb(w_n2534_0[1]),.din(n2534));
	jspl jspl_w_n2537_0(.douta(w_n2537_0[0]),.doutb(w_n2537_0[1]),.din(n2537));
	jspl jspl_w_n2540_0(.douta(w_n2540_0[0]),.doutb(w_n2540_0[1]),.din(n2540));
	jspl jspl_w_n2543_0(.douta(w_n2543_0[0]),.doutb(w_n2543_0[1]),.din(n2543));
	jspl jspl_w_n2551_0(.douta(w_n2551_0[0]),.doutb(w_n2551_0[1]),.din(n2551));
	jspl jspl_w_n2559_0(.douta(w_n2559_0[0]),.doutb(w_n2559_0[1]),.din(n2559));
	jspl jspl_w_n2567_0(.douta(w_n2567_0[0]),.doutb(w_n2567_0[1]),.din(n2567));
	jspl jspl_w_n2568_0(.douta(w_n2568_0[0]),.doutb(w_n2568_0[1]),.din(n2568));
	jspl jspl_w_n2569_0(.douta(w_n2569_0[0]),.doutb(w_n2569_0[1]),.din(n2569));
	jspl jspl_w_n2570_0(.douta(w_n2570_0[0]),.doutb(w_n2570_0[1]),.din(n2570));
	jspl jspl_w_n2573_0(.douta(w_n2573_0[0]),.doutb(w_n2573_0[1]),.din(n2573));
	jspl jspl_w_n2576_0(.douta(w_n2576_0[0]),.doutb(w_n2576_0[1]),.din(n2576));
	jspl jspl_w_n2577_0(.douta(w_n2577_0[0]),.doutb(w_n2577_0[1]),.din(n2577));
	jspl jspl_w_n2578_0(.douta(w_n2578_0[0]),.doutb(w_n2578_0[1]),.din(n2578));
	jspl jspl_w_n2579_0(.douta(w_n2579_0[0]),.doutb(w_n2579_0[1]),.din(n2579));
	jspl jspl_w_n2580_0(.douta(w_n2580_0[0]),.doutb(w_n2580_0[1]),.din(n2580));
	jspl jspl_w_n2581_0(.douta(w_n2581_0[0]),.doutb(w_n2581_0[1]),.din(n2581));
	jspl jspl_w_n2582_0(.douta(w_n2582_0[0]),.doutb(w_n2582_0[1]),.din(n2582));
	jspl3 jspl3_w_n2583_0(.douta(w_n2583_0[0]),.doutb(w_n2583_0[1]),.doutc(w_n2583_0[2]),.din(n2583));
	jspl jspl_w_n2583_1(.douta(w_n2583_1[0]),.doutb(w_n2583_1[1]),.din(w_n2583_0[0]));
	jspl jspl_w_n2586_0(.douta(w_n2586_0[0]),.doutb(w_n2586_0[1]),.din(n2586));
	jspl jspl_w_n2594_0(.douta(w_n2594_0[0]),.doutb(w_n2594_0[1]),.din(n2594));
	jspl jspl_w_n2596_0(.douta(w_n2596_0[0]),.doutb(w_n2596_0[1]),.din(n2596));
	jspl jspl_w_n2598_0(.douta(w_n2598_0[0]),.doutb(w_n2598_0[1]),.din(n2598));
	jspl jspl_w_n2600_0(.douta(w_n2600_0[0]),.doutb(w_n2600_0[1]),.din(n2600));
	jspl3 jspl3_w_n2601_0(.douta(w_n2601_0[0]),.doutb(w_n2601_0[1]),.doutc(w_n2601_0[2]),.din(n2601));
	jspl3 jspl3_w_n2602_0(.douta(w_n2602_0[0]),.doutb(w_n2602_0[1]),.doutc(w_n2602_0[2]),.din(n2602));
	jspl jspl_w_n2604_0(.douta(w_n2604_0[0]),.doutb(w_n2604_0[1]),.din(n2604));
	jspl jspl_w_n2606_0(.douta(w_n2606_0[0]),.doutb(w_n2606_0[1]),.din(n2606));
	jspl jspl_w_n2613_0(.douta(w_n2613_0[0]),.doutb(w_n2613_0[1]),.din(n2613));
	jspl jspl_w_n2617_0(.douta(w_n2617_0[0]),.doutb(w_n2617_0[1]),.din(n2617));
	jspl jspl_w_n2618_0(.douta(w_n2618_0[0]),.doutb(w_n2618_0[1]),.din(n2618));
	jspl3 jspl3_w_n2623_0(.douta(w_n2623_0[0]),.doutb(w_n2623_0[1]),.doutc(w_n2623_0[2]),.din(n2623));
	jspl jspl_w_n2628_0(.douta(w_n2628_0[0]),.doutb(w_n2628_0[1]),.din(n2628));
	jspl jspl_w_n2631_0(.douta(w_n2631_0[0]),.doutb(w_n2631_0[1]),.din(n2631));
	jspl3 jspl3_w_n2636_0(.douta(w_n2636_0[0]),.doutb(w_n2636_0[1]),.doutc(w_n2636_0[2]),.din(n2636));
	jspl jspl_w_n2637_0(.douta(w_n2637_0[0]),.doutb(w_n2637_0[1]),.din(n2637));
	jspl jspl_w_n2639_0(.douta(w_n2639_0[0]),.doutb(w_n2639_0[1]),.din(n2639));
	jspl jspl_w_n2642_0(.douta(w_n2642_0[0]),.doutb(w_n2642_0[1]),.din(n2642));
	jspl jspl_w_n2645_0(.douta(w_n2645_0[0]),.doutb(w_n2645_0[1]),.din(n2645));
	jspl jspl_w_n2653_0(.douta(w_n2653_0[0]),.doutb(w_n2653_0[1]),.din(n2653));
	jspl3 jspl3_w_n2654_0(.douta(w_n2654_0[0]),.doutb(w_n2654_0[1]),.doutc(w_n2654_0[2]),.din(n2654));
	jspl jspl_w_n2655_0(.douta(w_n2655_0[0]),.doutb(w_n2655_0[1]),.din(n2655));
	jspl jspl_w_n2659_0(.douta(w_n2659_0[0]),.doutb(w_n2659_0[1]),.din(n2659));
	jspl jspl_w_n2660_0(.douta(w_n2660_0[0]),.doutb(w_n2660_0[1]),.din(n2660));
	jspl jspl_w_n2661_0(.douta(w_n2661_0[0]),.doutb(w_n2661_0[1]),.din(n2661));
	jspl jspl_w_n2662_0(.douta(w_n2662_0[0]),.doutb(w_n2662_0[1]),.din(n2662));
	jspl jspl_w_n2665_0(.douta(w_n2665_0[0]),.doutb(w_n2665_0[1]),.din(n2665));
	jspl jspl_w_n2673_0(.douta(w_n2673_0[0]),.doutb(w_n2673_0[1]),.din(n2673));
	jspl jspl_w_n2676_0(.douta(w_n2676_0[0]),.doutb(w_n2676_0[1]),.din(n2676));
	jspl jspl_w_n2677_0(.douta(w_n2677_0[0]),.doutb(w_n2677_0[1]),.din(n2677));
	jspl jspl_w_n2678_0(.douta(w_n2678_0[0]),.doutb(w_n2678_0[1]),.din(n2678));
	jspl jspl_w_n2679_0(.douta(w_n2679_0[0]),.doutb(w_n2679_0[1]),.din(n2679));
	jspl3 jspl3_w_n2680_0(.douta(w_n2680_0[0]),.doutb(w_n2680_0[1]),.doutc(w_n2680_0[2]),.din(n2680));
	jspl jspl_w_n2680_1(.douta(w_n2680_1[0]),.doutb(w_n2680_1[1]),.din(w_n2680_0[0]));
	jspl3 jspl3_w_n2681_0(.douta(w_n2681_0[0]),.doutb(w_n2681_0[1]),.doutc(w_n2681_0[2]),.din(n2681));
	jspl3 jspl3_w_n2682_0(.douta(w_n2682_0[0]),.doutb(w_n2682_0[1]),.doutc(w_n2682_0[2]),.din(n2682));
	jspl3 jspl3_w_n2683_0(.douta(w_n2683_0[0]),.doutb(w_n2683_0[1]),.doutc(w_n2683_0[2]),.din(n2683));
	jspl3 jspl3_w_n2683_1(.douta(w_n2683_1[0]),.doutb(w_n2683_1[1]),.doutc(w_n2683_1[2]),.din(w_n2683_0[0]));
	jspl jspl_w_n2683_2(.douta(w_n2683_2[0]),.doutb(w_n2683_2[1]),.din(w_n2683_0[1]));
	jspl3 jspl3_w_n2684_0(.douta(w_n2684_0[0]),.doutb(w_n2684_0[1]),.doutc(w_n2684_0[2]),.din(n2684));
	jspl3 jspl3_w_n2684_1(.douta(w_n2684_1[0]),.doutb(w_n2684_1[1]),.doutc(w_n2684_1[2]),.din(w_n2684_0[0]));
	jspl3 jspl3_w_n2684_2(.douta(w_n2684_2[0]),.doutb(w_n2684_2[1]),.doutc(w_n2684_2[2]),.din(w_n2684_0[1]));
	jspl jspl_w_n2684_3(.douta(w_n2684_3[0]),.doutb(w_n2684_3[1]),.din(w_n2684_0[2]));
	jspl jspl_w_n2685_0(.douta(w_n2685_0[0]),.doutb(w_n2685_0[1]),.din(n2685));
	jspl3 jspl3_w_n2687_0(.douta(w_n2687_0[0]),.doutb(w_n2687_0[1]),.doutc(w_n2687_0[2]),.din(n2687));
	jspl3 jspl3_w_n2687_1(.douta(w_n2687_1[0]),.doutb(w_n2687_1[1]),.doutc(w_n2687_1[2]),.din(w_n2687_0[0]));
	jspl3 jspl3_w_n2687_2(.douta(w_n2687_2[0]),.doutb(w_n2687_2[1]),.doutc(w_n2687_2[2]),.din(w_n2687_0[1]));
	jspl jspl_w_n2687_3(.douta(w_n2687_3[0]),.doutb(w_n2687_3[1]),.din(w_n2687_0[2]));
	jspl jspl_w_n2688_0(.douta(w_n2688_0[0]),.doutb(w_n2688_0[1]),.din(n2688));
	jspl3 jspl3_w_n2690_0(.douta(w_n2690_0[0]),.doutb(w_n2690_0[1]),.doutc(w_n2690_0[2]),.din(n2690));
	jspl3 jspl3_w_n2690_1(.douta(w_n2690_1[0]),.doutb(w_n2690_1[1]),.doutc(w_n2690_1[2]),.din(w_n2690_0[0]));
	jspl3 jspl3_w_n2690_2(.douta(w_n2690_2[0]),.doutb(w_n2690_2[1]),.doutc(w_n2690_2[2]),.din(w_n2690_0[1]));
	jspl jspl_w_n2691_0(.douta(w_n2691_0[0]),.doutb(w_n2691_0[1]),.din(n2691));
	jspl jspl_w_n2695_0(.douta(w_n2695_0[0]),.doutb(w_n2695_0[1]),.din(n2695));
	jspl jspl_w_n2698_0(.douta(w_n2698_0[0]),.doutb(w_n2698_0[1]),.din(n2698));
	jspl jspl_w_n2703_0(.douta(w_n2703_0[0]),.doutb(w_n2703_0[1]),.din(n2703));
	jspl jspl_w_n2706_0(.douta(w_n2706_0[0]),.doutb(w_n2706_0[1]),.din(n2706));
	jspl3 jspl3_w_n2707_0(.douta(w_n2707_0[0]),.doutb(w_n2707_0[1]),.doutc(w_n2707_0[2]),.din(n2707));
	jspl3 jspl3_w_n2707_1(.douta(w_n2707_1[0]),.doutb(w_n2707_1[1]),.doutc(w_n2707_1[2]),.din(w_n2707_0[0]));
	jspl3 jspl3_w_n2707_2(.douta(w_n2707_2[0]),.doutb(w_n2707_2[1]),.doutc(w_n2707_2[2]),.din(w_n2707_0[1]));
	jspl3 jspl3_w_n2707_3(.douta(w_n2707_3[0]),.doutb(w_n2707_3[1]),.doutc(w_n2707_3[2]),.din(w_n2707_0[2]));
	jspl3 jspl3_w_n2707_4(.douta(w_n2707_4[0]),.doutb(w_n2707_4[1]),.doutc(w_n2707_4[2]),.din(w_n2707_1[0]));
	jspl3 jspl3_w_n2707_5(.douta(w_n2707_5[0]),.doutb(w_n2707_5[1]),.doutc(w_n2707_5[2]),.din(w_n2707_1[1]));
	jspl3 jspl3_w_n2707_6(.douta(w_n2707_6[0]),.doutb(w_n2707_6[1]),.doutc(w_n2707_6[2]),.din(w_n2707_1[2]));
	jspl jspl_w_n2707_7(.douta(w_n2707_7[0]),.doutb(w_n2707_7[1]),.din(w_n2707_2[0]));
	jspl jspl_w_n2710_0(.douta(w_n2710_0[0]),.doutb(w_n2710_0[1]),.din(n2710));
	jspl jspl_w_n2712_0(.douta(w_n2712_0[0]),.doutb(w_n2712_0[1]),.din(n2712));
	jspl jspl_w_n2715_0(.douta(w_n2715_0[0]),.doutb(w_n2715_0[1]),.din(n2715));
	jspl3 jspl3_w_n2717_0(.douta(w_n2717_0[0]),.doutb(w_n2717_0[1]),.doutc(w_n2717_0[2]),.din(n2717));
	jspl jspl_w_n2725_0(.douta(w_n2725_0[0]),.doutb(w_n2725_0[1]),.din(n2725));
	jspl jspl_w_n2729_0(.douta(w_n2729_0[0]),.doutb(w_n2729_0[1]),.din(n2729));
	jspl jspl_w_n2732_0(.douta(w_n2732_0[0]),.doutb(w_n2732_0[1]),.din(n2732));
	jspl3 jspl3_w_n2738_0(.douta(w_n2738_0[0]),.doutb(w_n2738_0[1]),.doutc(w_n2738_0[2]),.din(n2738));
	jspl3 jspl3_w_n2743_0(.douta(w_n2743_0[0]),.doutb(w_n2743_0[1]),.doutc(w_n2743_0[2]),.din(n2743));
	jspl jspl_w_n2744_0(.douta(w_n2744_0[0]),.doutb(w_n2744_0[1]),.din(n2744));
	jspl jspl_w_n2751_0(.douta(w_n2751_0[0]),.doutb(w_n2751_0[1]),.din(n2751));
	jspl3 jspl3_w_n2759_0(.douta(w_n2759_0[0]),.doutb(w_n2759_0[1]),.doutc(w_n2759_0[2]),.din(n2759));
	jspl jspl_w_n2760_0(.douta(w_n2760_0[0]),.doutb(w_n2760_0[1]),.din(n2760));
	jspl jspl_w_n2762_0(.douta(w_n2762_0[0]),.doutb(w_n2762_0[1]),.din(n2762));
	jspl jspl_w_n2765_0(.douta(w_n2765_0[0]),.doutb(w_n2765_0[1]),.din(n2765));
	jspl jspl_w_n2768_0(.douta(w_n2768_0[0]),.doutb(w_n2768_0[1]),.din(n2768));
	jspl jspl_w_n2769_0(.douta(w_n2769_0[0]),.doutb(w_n2769_0[1]),.din(n2769));
	jspl jspl_w_n2770_0(.douta(w_n2770_0[0]),.doutb(w_n2770_0[1]),.din(n2770));
	jspl jspl_w_n2771_0(.douta(w_n2771_0[0]),.doutb(w_n2771_0[1]),.din(n2771));
	jspl jspl_w_n2772_0(.douta(w_n2772_0[0]),.doutb(w_n2772_0[1]),.din(n2772));
	jspl jspl_w_n2773_0(.douta(w_n2773_0[0]),.doutb(w_n2773_0[1]),.din(n2773));
	jspl jspl_w_n2777_0(.douta(w_n2777_0[0]),.doutb(w_n2777_0[1]),.din(n2777));
	jspl jspl_w_n2785_0(.douta(w_n2785_0[0]),.doutb(w_n2785_0[1]),.din(n2785));
	jspl jspl_w_n2793_0(.douta(w_n2793_0[0]),.doutb(w_n2793_0[1]),.din(n2793));
	jspl jspl_w_n2794_0(.douta(w_n2794_0[0]),.doutb(w_n2794_0[1]),.din(n2794));
	jspl jspl_w_n2795_0(.douta(w_n2795_0[0]),.doutb(w_n2795_0[1]),.din(n2795));
	jspl jspl_w_n2796_0(.douta(w_n2796_0[0]),.doutb(w_n2796_0[1]),.din(n2796));
	jspl3 jspl3_w_n2797_0(.douta(w_n2797_0[0]),.doutb(w_n2797_0[1]),.doutc(w_n2797_0[2]),.din(n2797));
	jspl jspl_w_n2797_1(.douta(w_n2797_1[0]),.doutb(w_n2797_1[1]),.din(w_n2797_0[0]));
	jspl3 jspl3_w_n2798_0(.douta(w_n2798_0[0]),.doutb(w_n2798_0[1]),.doutc(w_n2798_0[2]),.din(n2798));
	jspl3 jspl3_w_n2799_0(.douta(w_n2799_0[0]),.doutb(w_n2799_0[1]),.doutc(w_n2799_0[2]),.din(n2799));
	jspl3 jspl3_w_n2800_0(.douta(w_n2800_0[0]),.doutb(w_n2800_0[1]),.doutc(w_n2800_0[2]),.din(n2800));
	jspl3 jspl3_w_n2800_1(.douta(w_n2800_1[0]),.doutb(w_n2800_1[1]),.doutc(w_n2800_1[2]),.din(w_n2800_0[0]));
	jspl3 jspl3_w_n2800_2(.douta(w_n2800_2[0]),.doutb(w_n2800_2[1]),.doutc(w_n2800_2[2]),.din(w_n2800_0[1]));
	jspl3 jspl3_w_n2800_3(.douta(w_n2800_3[0]),.doutb(w_n2800_3[1]),.doutc(w_n2800_3[2]),.din(w_n2800_0[2]));
	jspl3 jspl3_w_n2800_4(.douta(w_n2800_4[0]),.doutb(w_n2800_4[1]),.doutc(w_n2800_4[2]),.din(w_n2800_1[0]));
	jspl3 jspl3_w_n2800_5(.douta(w_n2800_5[0]),.doutb(w_n2800_5[1]),.doutc(w_n2800_5[2]),.din(w_n2800_1[1]));
	jspl3 jspl3_w_n2800_6(.douta(w_n2800_6[0]),.doutb(w_n2800_6[1]),.doutc(w_n2800_6[2]),.din(w_n2800_1[2]));
	jspl jspl_w_n2800_7(.douta(w_n2800_7[0]),.doutb(w_n2800_7[1]),.din(w_n2800_2[0]));
	jspl jspl_w_n2801_0(.douta(w_n2801_0[0]),.doutb(w_n2801_0[1]),.din(n2801));
	jspl3 jspl3_w_n2802_0(.douta(w_n2802_0[0]),.doutb(w_n2802_0[1]),.doutc(w_n2802_0[2]),.din(n2802));
	jspl3 jspl3_w_n2802_1(.douta(w_n2802_1[0]),.doutb(w_n2802_1[1]),.doutc(w_n2802_1[2]),.din(w_n2802_0[0]));
	jspl jspl_w_n2804_0(.douta(w_n2804_0[0]),.doutb(w_n2804_0[1]),.din(n2804));
	jspl3 jspl3_w_n2806_0(.douta(w_n2806_0[0]),.doutb(w_n2806_0[1]),.doutc(w_n2806_0[2]),.din(n2806));
	jspl3 jspl3_w_n2807_0(.douta(w_n2807_0[0]),.doutb(w_n2807_0[1]),.doutc(w_n2807_0[2]),.din(n2807));
	jspl3 jspl3_w_n2807_1(.douta(w_n2807_1[0]),.doutb(w_n2807_1[1]),.doutc(w_n2807_1[2]),.din(w_n2807_0[0]));
	jspl3 jspl3_w_n2807_2(.douta(w_n2807_2[0]),.doutb(w_n2807_2[1]),.doutc(w_n2807_2[2]),.din(w_n2807_0[1]));
	jspl3 jspl3_w_n2807_3(.douta(w_n2807_3[0]),.doutb(w_n2807_3[1]),.doutc(w_n2807_3[2]),.din(w_n2807_0[2]));
	jspl3 jspl3_w_n2807_4(.douta(w_n2807_4[0]),.doutb(w_n2807_4[1]),.doutc(w_n2807_4[2]),.din(w_n2807_1[0]));
	jspl3 jspl3_w_n2807_5(.douta(w_n2807_5[0]),.doutb(w_n2807_5[1]),.doutc(w_n2807_5[2]),.din(w_n2807_1[1]));
	jspl3 jspl3_w_n2807_6(.douta(w_n2807_6[0]),.doutb(w_n2807_6[1]),.doutc(w_n2807_6[2]),.din(w_n2807_1[2]));
	jspl3 jspl3_w_n2807_7(.douta(w_n2807_7[0]),.doutb(w_n2807_7[1]),.doutc(w_n2807_7[2]),.din(w_n2807_2[0]));
	jspl3 jspl3_w_n2809_0(.douta(w_n2809_0[0]),.doutb(w_n2809_0[1]),.doutc(w_n2809_0[2]),.din(n2809));
	jspl3 jspl3_w_n2810_0(.douta(w_n2810_0[0]),.doutb(w_n2810_0[1]),.doutc(w_n2810_0[2]),.din(n2810));
	jspl3 jspl3_w_n2810_1(.douta(w_n2810_1[0]),.doutb(w_n2810_1[1]),.doutc(w_n2810_1[2]),.din(w_n2810_0[0]));
	jspl3 jspl3_w_n2810_2(.douta(w_n2810_2[0]),.doutb(w_n2810_2[1]),.doutc(w_n2810_2[2]),.din(w_n2810_0[1]));
	jspl3 jspl3_w_n2810_3(.douta(w_n2810_3[0]),.doutb(w_n2810_3[1]),.doutc(w_n2810_3[2]),.din(w_n2810_0[2]));
	jspl3 jspl3_w_n2810_4(.douta(w_n2810_4[0]),.doutb(w_n2810_4[1]),.doutc(w_n2810_4[2]),.din(w_n2810_1[0]));
	jspl3 jspl3_w_n2810_5(.douta(w_n2810_5[0]),.doutb(w_n2810_5[1]),.doutc(w_n2810_5[2]),.din(w_n2810_1[1]));
	jspl3 jspl3_w_n2810_6(.douta(w_n2810_6[0]),.doutb(w_n2810_6[1]),.doutc(w_n2810_6[2]),.din(w_n2810_1[2]));
	jspl jspl_w_n2810_7(.douta(w_n2810_7[0]),.doutb(w_n2810_7[1]),.din(w_n2810_2[0]));
	jspl3 jspl3_w_n2813_0(.douta(w_n2813_0[0]),.doutb(w_n2813_0[1]),.doutc(w_n2813_0[2]),.din(n2813));
	jspl3 jspl3_w_n2813_1(.douta(w_n2813_1[0]),.doutb(w_n2813_1[1]),.doutc(w_n2813_1[2]),.din(w_n2813_0[0]));
	jspl3 jspl3_w_n2813_2(.douta(w_n2813_2[0]),.doutb(w_n2813_2[1]),.doutc(w_n2813_2[2]),.din(w_n2813_0[1]));
	jspl3 jspl3_w_n2813_3(.douta(w_n2813_3[0]),.doutb(w_n2813_3[1]),.doutc(w_n2813_3[2]),.din(w_n2813_0[2]));
	jspl3 jspl3_w_n2813_4(.douta(w_n2813_4[0]),.doutb(w_n2813_4[1]),.doutc(w_n2813_4[2]),.din(w_n2813_1[0]));
	jspl3 jspl3_w_n2813_5(.douta(w_n2813_5[0]),.doutb(w_n2813_5[1]),.doutc(w_n2813_5[2]),.din(w_n2813_1[1]));
	jspl3 jspl3_w_n2813_6(.douta(w_n2813_6[0]),.doutb(w_n2813_6[1]),.doutc(w_n2813_6[2]),.din(w_n2813_1[2]));
	jspl3 jspl3_w_n2815_0(.douta(w_n2815_0[0]),.doutb(w_n2815_0[1]),.doutc(w_n2815_0[2]),.din(n2815));
	jspl3 jspl3_w_n2816_0(.douta(w_n2816_0[0]),.doutb(w_n2816_0[1]),.doutc(w_n2816_0[2]),.din(n2816));
	jspl3 jspl3_w_n2816_1(.douta(w_n2816_1[0]),.doutb(w_n2816_1[1]),.doutc(w_n2816_1[2]),.din(w_n2816_0[0]));
	jspl3 jspl3_w_n2816_2(.douta(w_n2816_2[0]),.doutb(w_n2816_2[1]),.doutc(w_n2816_2[2]),.din(w_n2816_0[1]));
	jspl3 jspl3_w_n2816_3(.douta(w_n2816_3[0]),.doutb(w_n2816_3[1]),.doutc(w_n2816_3[2]),.din(w_n2816_0[2]));
	jspl3 jspl3_w_n2816_4(.douta(w_n2816_4[0]),.doutb(w_n2816_4[1]),.doutc(w_n2816_4[2]),.din(w_n2816_1[0]));
	jspl3 jspl3_w_n2816_5(.douta(w_n2816_5[0]),.doutb(w_n2816_5[1]),.doutc(w_n2816_5[2]),.din(w_n2816_1[1]));
	jspl3 jspl3_w_n2816_6(.douta(w_n2816_6[0]),.doutb(w_n2816_6[1]),.doutc(w_n2816_6[2]),.din(w_n2816_1[2]));
	jspl3 jspl3_w_n2816_7(.douta(w_n2816_7[0]),.doutb(w_n2816_7[1]),.doutc(w_n2816_7[2]),.din(w_n2816_2[0]));
	jspl jspl_w_n2820_0(.douta(w_n2820_0[0]),.doutb(w_n2820_0[1]),.din(n2820));
	jspl jspl_w_n2823_0(.douta(w_n2823_0[0]),.doutb(w_n2823_0[1]),.din(n2823));
	jspl jspl_w_n2824_0(.douta(w_n2824_0[0]),.doutb(w_n2824_0[1]),.din(n2824));
	jspl3 jspl3_w_n2825_0(.douta(w_n2825_0[0]),.doutb(w_n2825_0[1]),.doutc(w_n2825_0[2]),.din(n2825));
	jspl3 jspl3_w_n2825_1(.douta(w_n2825_1[0]),.doutb(w_n2825_1[1]),.doutc(w_n2825_1[2]),.din(w_n2825_0[0]));
	jspl jspl_w_n2833_0(.douta(w_n2833_0[0]),.doutb(w_n2833_0[1]),.din(n2833));
	jspl jspl_w_n2835_0(.douta(w_n2835_0[0]),.doutb(w_n2835_0[1]),.din(n2835));
	jspl3 jspl3_w_n2836_0(.douta(w_n2836_0[0]),.doutb(w_n2836_0[1]),.doutc(w_n2836_0[2]),.din(n2836));
	jspl3 jspl3_w_n2836_1(.douta(w_n2836_1[0]),.doutb(w_n2836_1[1]),.doutc(w_n2836_1[2]),.din(w_n2836_0[0]));
	jspl jspl_w_n2845_0(.douta(w_n2845_0[0]),.doutb(w_n2845_0[1]),.din(n2845));
	jspl jspl_w_n2847_0(.douta(w_n2847_0[0]),.doutb(w_n2847_0[1]),.din(n2847));
	jspl jspl_w_n2857_0(.douta(w_n2857_0[0]),.doutb(w_n2857_0[1]),.din(n2857));
	jspl jspl_w_n2859_0(.douta(w_n2859_0[0]),.doutb(w_n2859_0[1]),.din(n2859));
	jspl jspl_w_n2865_0(.douta(w_n2865_0[0]),.doutb(w_n2865_0[1]),.din(n2865));
	jspl3 jspl3_w_n2867_0(.douta(w_n2867_0[0]),.doutb(w_n2867_0[1]),.doutc(w_n2867_0[2]),.din(n2867));
	jspl jspl_w_n2867_1(.douta(w_n2867_1[0]),.doutb(w_n2867_1[1]),.din(w_n2867_0[0]));
	jspl jspl_w_n2870_0(.douta(w_n2870_0[0]),.doutb(w_n2870_0[1]),.din(n2870));
	jspl jspl_w_n2878_0(.douta(w_n2878_0[0]),.doutb(w_n2878_0[1]),.din(n2878));
	jspl jspl_w_n2879_0(.douta(w_n2879_0[0]),.doutb(w_n2879_0[1]),.din(n2879));
	jspl jspl_w_n2881_0(.douta(w_n2881_0[0]),.doutb(w_n2881_0[1]),.din(n2881));
	jspl jspl_w_n2889_0(.douta(w_n2889_0[0]),.doutb(w_n2889_0[1]),.din(n2889));
	jspl jspl_w_n2891_0(.douta(w_n2891_0[0]),.doutb(w_n2891_0[1]),.din(n2891));
	jspl jspl_w_n2892_0(.douta(w_n2892_0[0]),.doutb(w_n2892_0[1]),.din(n2892));
	jspl jspl_w_n2894_0(.douta(w_n2894_0[0]),.doutb(w_n2894_0[1]),.din(n2894));
	jspl jspl_w_n2895_0(.douta(w_n2895_0[0]),.doutb(w_n2895_0[1]),.din(n2895));
	jspl jspl_w_n2897_0(.douta(w_n2897_0[0]),.doutb(w_n2897_0[1]),.din(n2897));
	jspl jspl_w_n2898_0(.douta(w_n2898_0[0]),.doutb(w_n2898_0[1]),.din(n2898));
	jspl jspl_w_n2902_0(.douta(w_n2902_0[0]),.doutb(w_n2902_0[1]),.din(n2902));
	jspl jspl_w_n2903_0(.douta(w_n2903_0[0]),.doutb(w_n2903_0[1]),.din(n2903));
	jspl jspl_w_n2906_0(.douta(w_n2906_0[0]),.doutb(w_n2906_0[1]),.din(n2906));
	jspl jspl_w_n2909_0(.douta(w_n2909_0[0]),.doutb(w_n2909_0[1]),.din(n2909));
	jspl jspl_w_n2918_0(.douta(w_n2918_0[0]),.doutb(w_n2918_0[1]),.din(n2918));
	jspl3 jspl3_w_n2923_0(.douta(w_n2923_0[0]),.doutb(w_n2923_0[1]),.doutc(w_n2923_0[2]),.din(n2923));
	jspl3 jspl3_w_n2923_1(.douta(w_n2923_1[0]),.doutb(w_n2923_1[1]),.doutc(w_n2923_1[2]),.din(w_n2923_0[0]));
	jspl3 jspl3_w_n2923_2(.douta(w_n2923_2[0]),.doutb(w_n2923_2[1]),.doutc(w_n2923_2[2]),.din(w_n2923_0[1]));
	jspl3 jspl3_w_n2923_3(.douta(w_n2923_3[0]),.doutb(w_n2923_3[1]),.doutc(w_n2923_3[2]),.din(w_n2923_0[2]));
	jspl jspl_w_n2927_0(.douta(w_n2927_0[0]),.doutb(w_n2927_0[1]),.din(n2927));
	jspl jspl_w_n2929_0(.douta(w_n2929_0[0]),.doutb(w_n2929_0[1]),.din(n2929));
	jspl jspl_w_n2931_0(.douta(w_n2931_0[0]),.doutb(w_n2931_0[1]),.din(n2931));
	jspl jspl_w_n2932_0(.douta(w_n2932_0[0]),.doutb(w_n2932_0[1]),.din(n2932));
	jspl jspl_w_n2934_0(.douta(w_n2934_0[0]),.doutb(w_n2934_0[1]),.din(n2934));
	jspl jspl_w_n2938_0(.douta(w_n2938_0[0]),.doutb(w_n2938_0[1]),.din(n2938));
	jspl jspl_w_n2942_0(.douta(w_n2942_0[0]),.doutb(w_n2942_0[1]),.din(n2942));
	jspl3 jspl3_w_n2943_0(.douta(w_n2943_0[0]),.doutb(w_n2943_0[1]),.doutc(w_n2943_0[2]),.din(n2943));
	jspl3 jspl3_w_n2943_1(.douta(w_n2943_1[0]),.doutb(w_n2943_1[1]),.doutc(w_n2943_1[2]),.din(w_n2943_0[0]));
	jspl jspl_w_n2943_2(.douta(w_n2943_2[0]),.doutb(w_n2943_2[1]),.din(w_n2943_0[1]));
	jspl jspl_w_n2944_0(.douta(w_n2944_0[0]),.doutb(w_n2944_0[1]),.din(n2944));
	jspl jspl_w_n2948_0(.douta(w_n2948_0[0]),.doutb(w_n2948_0[1]),.din(n2948));
	jspl jspl_w_n2950_0(.douta(w_n2950_0[0]),.doutb(w_n2950_0[1]),.din(n2950));
	jspl jspl_w_n2953_0(.douta(w_n2953_0[0]),.doutb(w_n2953_0[1]),.din(n2953));
	jspl jspl_w_n2954_0(.douta(w_n2954_0[0]),.doutb(w_n2954_0[1]),.din(n2954));
	jspl jspl_w_n2964_0(.douta(w_n2964_0[0]),.doutb(w_n2964_0[1]),.din(n2964));
	jspl jspl_w_n2968_0(.douta(w_n2968_0[0]),.doutb(w_n2968_0[1]),.din(n2968));
	jspl jspl_w_n2971_0(.douta(w_n2971_0[0]),.doutb(w_n2971_0[1]),.din(n2971));
	jspl3 jspl3_w_n2973_0(.douta(w_n2973_0[0]),.doutb(w_n2973_0[1]),.doutc(w_n2973_0[2]),.din(n2973));
	jspl jspl_w_n2974_0(.douta(w_n2974_0[0]),.doutb(w_n2974_0[1]),.din(n2974));
	jspl jspl_w_n2976_0(.douta(w_n2976_0[0]),.doutb(w_n2976_0[1]),.din(n2976));
	jspl jspl_w_n2979_0(.douta(w_n2979_0[0]),.doutb(w_n2979_0[1]),.din(n2979));
	jspl jspl_w_n2987_0(.douta(w_n2987_0[0]),.doutb(w_n2987_0[1]),.din(n2987));
	jspl3 jspl3_w_n2988_0(.douta(w_n2988_0[0]),.doutb(w_n2988_0[1]),.doutc(w_n2988_0[2]),.din(n2988));
	jspl jspl_w_n2990_0(.douta(w_n2990_0[0]),.doutb(w_n2990_0[1]),.din(n2990));
	jspl jspl_w_n2994_0(.douta(w_n2994_0[0]),.doutb(w_n2994_0[1]),.din(n2994));
	jspl jspl_w_n2995_0(.douta(w_n2995_0[0]),.doutb(w_n2995_0[1]),.din(n2995));
	jspl jspl_w_n2996_0(.douta(w_n2996_0[0]),.doutb(w_n2996_0[1]),.din(n2996));
	jspl jspl_w_n2999_0(.douta(w_n2999_0[0]),.doutb(w_n2999_0[1]),.din(n2999));
	jspl jspl_w_n3002_0(.douta(w_n3002_0[0]),.doutb(w_n3002_0[1]),.din(n3002));
	jspl jspl_w_n3003_0(.douta(w_n3003_0[0]),.doutb(w_n3003_0[1]),.din(n3003));
	jspl jspl_w_n3004_0(.douta(w_n3004_0[0]),.doutb(w_n3004_0[1]),.din(n3004));
	jspl3 jspl3_w_n3005_0(.douta(w_n3005_0[0]),.doutb(w_n3005_0[1]),.doutc(w_n3005_0[2]),.din(n3005));
	jspl jspl_w_n3005_1(.douta(w_n3005_1[0]),.doutb(w_n3005_1[1]),.din(w_n3005_0[0]));
	jspl3 jspl3_w_n3006_0(.douta(w_n3006_0[0]),.doutb(w_n3006_0[1]),.doutc(w_n3006_0[2]),.din(n3006));
	jspl3 jspl3_w_n3007_0(.douta(w_n3007_0[0]),.doutb(w_n3007_0[1]),.doutc(w_n3007_0[2]),.din(n3007));
	jspl3 jspl3_w_n3008_0(.douta(w_n3008_0[0]),.doutb(w_n3008_0[1]),.doutc(w_n3008_0[2]),.din(n3008));
	jspl3 jspl3_w_n3008_1(.douta(w_n3008_1[0]),.doutb(w_n3008_1[1]),.doutc(w_n3008_1[2]),.din(w_n3008_0[0]));
	jspl3 jspl3_w_n3008_2(.douta(w_n3008_2[0]),.doutb(w_n3008_2[1]),.doutc(w_n3008_2[2]),.din(w_n3008_0[1]));
	jspl3 jspl3_w_n3008_3(.douta(w_n3008_3[0]),.doutb(w_n3008_3[1]),.doutc(w_n3008_3[2]),.din(w_n3008_0[2]));
	jspl3 jspl3_w_n3008_4(.douta(w_n3008_4[0]),.doutb(w_n3008_4[1]),.doutc(w_n3008_4[2]),.din(w_n3008_1[0]));
	jspl3 jspl3_w_n3008_5(.douta(w_n3008_5[0]),.doutb(w_n3008_5[1]),.doutc(w_n3008_5[2]),.din(w_n3008_1[1]));
	jspl3 jspl3_w_n3008_6(.douta(w_n3008_6[0]),.doutb(w_n3008_6[1]),.doutc(w_n3008_6[2]),.din(w_n3008_1[2]));
	jspl3 jspl3_w_n3008_7(.douta(w_n3008_7[0]),.doutb(w_n3008_7[1]),.doutc(w_n3008_7[2]),.din(w_n3008_2[0]));
	jspl jspl_w_n3009_0(.douta(w_n3009_0[0]),.doutb(w_n3009_0[1]),.din(n3009));
	jspl3 jspl3_w_n3010_0(.douta(w_n3010_0[0]),.doutb(w_n3010_0[1]),.doutc(w_n3010_0[2]),.din(n3010));
	jspl3 jspl3_w_n3010_1(.douta(w_n3010_1[0]),.doutb(w_n3010_1[1]),.doutc(w_n3010_1[2]),.din(w_n3010_0[0]));
	jspl jspl_w_n3018_0(.douta(w_n3018_0[0]),.doutb(w_n3018_0[1]),.din(n3018));
	jspl jspl_w_n3019_0(.douta(w_n3019_0[0]),.doutb(w_n3019_0[1]),.din(n3019));
	jspl jspl_w_n3020_0(.douta(w_n3020_0[0]),.doutb(w_n3020_0[1]),.din(n3020));
	jspl jspl_w_n3021_0(.douta(w_n3021_0[0]),.doutb(w_n3021_0[1]),.din(n3021));
	jspl3 jspl3_w_n3023_0(.douta(w_n3023_0[0]),.doutb(w_n3023_0[1]),.doutc(w_n3023_0[2]),.din(n3023));
	jspl3 jspl3_w_n3023_1(.douta(w_n3023_1[0]),.doutb(w_n3023_1[1]),.doutc(w_n3023_1[2]),.din(w_n3023_0[0]));
	jspl3 jspl3_w_n3023_2(.douta(w_n3023_2[0]),.doutb(w_n3023_2[1]),.doutc(w_n3023_2[2]),.din(w_n3023_0[1]));
	jspl3 jspl3_w_n3023_3(.douta(w_n3023_3[0]),.doutb(w_n3023_3[1]),.doutc(w_n3023_3[2]),.din(w_n3023_0[2]));
	jspl3 jspl3_w_n3023_4(.douta(w_n3023_4[0]),.doutb(w_n3023_4[1]),.doutc(w_n3023_4[2]),.din(w_n3023_1[0]));
	jspl3 jspl3_w_n3023_5(.douta(w_n3023_5[0]),.doutb(w_n3023_5[1]),.doutc(w_n3023_5[2]),.din(w_n3023_1[1]));
	jspl3 jspl3_w_n3023_6(.douta(w_n3023_6[0]),.doutb(w_n3023_6[1]),.doutc(w_n3023_6[2]),.din(w_n3023_1[2]));
	jspl3 jspl3_w_n3023_7(.douta(w_n3023_7[0]),.doutb(w_n3023_7[1]),.doutc(w_n3023_7[2]),.din(w_n3023_2[0]));
	jspl3 jspl3_w_n3023_8(.douta(w_n3023_8[0]),.doutb(w_n3023_8[1]),.doutc(w_n3023_8[2]),.din(w_n3023_2[1]));
	jspl3 jspl3_w_n3023_9(.douta(w_n3023_9[0]),.doutb(w_n3023_9[1]),.doutc(w_n3023_9[2]),.din(w_n3023_2[2]));
	jspl3 jspl3_w_n3023_10(.douta(w_n3023_10[0]),.doutb(w_n3023_10[1]),.doutc(w_n3023_10[2]),.din(w_n3023_3[0]));
	jspl3 jspl3_w_n3024_0(.douta(w_n3024_0[0]),.doutb(w_n3024_0[1]),.doutc(w_n3024_0[2]),.din(n3024));
	jspl3 jspl3_w_n3025_0(.douta(w_n3025_0[0]),.doutb(w_n3025_0[1]),.doutc(w_n3025_0[2]),.din(n3025));
	jspl jspl_w_n3026_0(.douta(w_n3026_0[0]),.doutb(w_n3026_0[1]),.din(n3026));
	jspl jspl_w_n3027_0(.douta(w_n3027_0[0]),.doutb(w_n3027_0[1]),.din(n3027));
	jspl3 jspl3_w_n3028_0(.douta(w_n3028_0[0]),.doutb(w_n3028_0[1]),.doutc(w_n3028_0[2]),.din(n3028));
	jspl jspl_w_n3028_1(.douta(w_n3028_1[0]),.doutb(w_n3028_1[1]),.din(w_n3028_0[0]));
	jspl3 jspl3_w_n3029_0(.douta(w_n3029_0[0]),.doutb(w_n3029_0[1]),.doutc(w_n3029_0[2]),.din(n3029));
	jspl3 jspl3_w_n3029_1(.douta(w_n3029_1[0]),.doutb(w_n3029_1[1]),.doutc(w_n3029_1[2]),.din(w_n3029_0[0]));
	jspl3 jspl3_w_n3029_2(.douta(w_n3029_2[0]),.doutb(w_n3029_2[1]),.doutc(w_n3029_2[2]),.din(w_n3029_0[1]));
	jspl3 jspl3_w_n3029_3(.douta(w_n3029_3[0]),.doutb(w_n3029_3[1]),.doutc(w_n3029_3[2]),.din(w_n3029_0[2]));
	jspl3 jspl3_w_n3029_4(.douta(w_n3029_4[0]),.doutb(w_n3029_4[1]),.doutc(w_n3029_4[2]),.din(w_n3029_1[0]));
	jspl3 jspl3_w_n3029_5(.douta(w_n3029_5[0]),.doutb(w_n3029_5[1]),.doutc(w_n3029_5[2]),.din(w_n3029_1[1]));
	jspl3 jspl3_w_n3029_6(.douta(w_n3029_6[0]),.doutb(w_n3029_6[1]),.doutc(w_n3029_6[2]),.din(w_n3029_1[2]));
	jspl3 jspl3_w_n3029_7(.douta(w_n3029_7[0]),.doutb(w_n3029_7[1]),.doutc(w_n3029_7[2]),.din(w_n3029_2[0]));
	jspl3 jspl3_w_n3042_0(.douta(w_n3042_0[0]),.doutb(w_n3042_0[1]),.doutc(w_n3042_0[2]),.din(n3042));
	jspl jspl_w_n3043_0(.douta(w_n3043_0[0]),.doutb(w_n3043_0[1]),.din(n3043));
	jspl jspl_w_n3044_0(.douta(w_n3044_0[0]),.doutb(w_n3044_0[1]),.din(n3044));
	jspl jspl_w_n3050_0(.douta(w_n3050_0[0]),.doutb(w_n3050_0[1]),.din(n3050));
	jspl jspl_w_n3053_0(.douta(w_n3053_0[0]),.doutb(w_n3053_0[1]),.din(n3053));
	jspl jspl_w_n3059_0(.douta(w_n3059_0[0]),.doutb(w_n3059_0[1]),.din(n3059));
	jspl jspl_w_n3065_0(.douta(w_n3065_0[0]),.doutb(w_n3065_0[1]),.din(n3065));
	jspl jspl_w_n3069_0(.douta(w_n3069_0[0]),.doutb(w_n3069_0[1]),.din(n3069));
	jspl jspl_w_n3070_0(.douta(w_n3070_0[0]),.doutb(w_n3070_0[1]),.din(n3070));
	jspl jspl_w_n3071_0(.douta(w_n3071_0[0]),.doutb(w_n3071_0[1]),.din(n3071));
	jspl jspl_w_n3072_0(.douta(w_n3072_0[0]),.doutb(w_n3072_0[1]),.din(n3072));
	jspl jspl_w_n3073_0(.douta(w_n3073_0[0]),.doutb(w_n3073_0[1]),.din(n3073));
	jspl jspl_w_n3074_0(.douta(w_n3074_0[0]),.doutb(w_n3074_0[1]),.din(n3074));
	jspl jspl_w_n3075_0(.douta(w_n3075_0[0]),.doutb(w_n3075_0[1]),.din(n3075));
	jspl3 jspl3_w_n3076_0(.douta(w_n3076_0[0]),.doutb(w_n3076_0[1]),.doutc(w_n3076_0[2]),.din(n3076));
	jspl jspl_w_n3079_0(.douta(w_n3079_0[0]),.doutb(w_n3079_0[1]),.din(n3079));
	jspl jspl_w_n3085_0(.douta(w_n3085_0[0]),.doutb(w_n3085_0[1]),.din(n3085));
	jspl jspl_w_n3087_0(.douta(w_n3087_0[0]),.doutb(w_n3087_0[1]),.din(n3087));
	jspl jspl_w_n3089_0(.douta(w_n3089_0[0]),.doutb(w_n3089_0[1]),.din(n3089));
	jspl3 jspl3_w_n3090_0(.douta(w_n3090_0[0]),.doutb(w_n3090_0[1]),.doutc(w_n3090_0[2]),.din(n3090));
	jspl3 jspl3_w_n3091_0(.douta(w_n3091_0[0]),.doutb(w_n3091_0[1]),.doutc(w_n3091_0[2]),.din(n3091));
	jspl jspl_w_n3093_0(.douta(w_n3093_0[0]),.doutb(w_n3093_0[1]),.din(n3093));
	jspl jspl_w_n3098_0(.douta(w_n3098_0[0]),.doutb(w_n3098_0[1]),.din(n3098));
	jspl jspl_w_n3106_0(.douta(w_n3106_0[0]),.doutb(w_n3106_0[1]),.din(n3106));
	jspl3 jspl3_w_n3118_0(.douta(w_n3118_0[0]),.doutb(w_n3118_0[1]),.doutc(w_n3118_0[2]),.din(n3118));
	jspl3 jspl3_w_n3121_0(.douta(w_n3121_0[0]),.doutb(w_n3121_0[1]),.doutc(w_n3121_0[2]),.din(n3121));
	jspl jspl_w_n3126_0(.douta(w_n3126_0[0]),.doutb(w_n3126_0[1]),.din(n3126));
	jspl jspl_w_n3130_0(.douta(w_n3130_0[0]),.doutb(w_n3130_0[1]),.din(n3130));
	jspl jspl_w_n3131_0(.douta(w_n3131_0[0]),.doutb(w_n3131_0[1]),.din(n3131));
	jspl jspl_w_n3132_0(.douta(w_n3132_0[0]),.doutb(w_n3132_0[1]),.din(n3132));
	jspl jspl_w_n3136_0(.douta(w_n3136_0[0]),.doutb(w_n3136_0[1]),.din(n3136));
	jspl jspl_w_n3138_0(.douta(w_n3138_0[0]),.doutb(w_n3138_0[1]),.din(n3138));
	jspl jspl_w_n3139_0(.douta(w_n3139_0[0]),.doutb(w_n3139_0[1]),.din(n3139));
	jspl3 jspl3_w_n3140_0(.douta(w_n3140_0[0]),.doutb(w_n3140_0[1]),.doutc(w_n3140_0[2]),.din(n3140));
	jspl3 jspl3_w_n3141_0(.douta(w_n3141_0[0]),.doutb(w_n3141_0[1]),.doutc(w_n3141_0[2]),.din(n3141));
	jspl3 jspl3_w_n3142_0(.douta(w_n3142_0[0]),.doutb(w_n3142_0[1]),.doutc(w_n3142_0[2]),.din(n3142));
	jspl3 jspl3_w_n3143_0(.douta(w_n3143_0[0]),.doutb(w_n3143_0[1]),.doutc(w_n3143_0[2]),.din(n3143));
	jspl jspl_w_n3143_1(.douta(w_n3143_1[0]),.doutb(w_n3143_1[1]),.din(w_n3143_0[0]));
	jspl3 jspl3_w_n3144_0(.douta(w_n3144_0[0]),.doutb(w_n3144_0[1]),.doutc(w_n3144_0[2]),.din(n3144));
	jspl3 jspl3_w_n3144_1(.douta(w_n3144_1[0]),.doutb(w_n3144_1[1]),.doutc(w_n3144_1[2]),.din(w_n3144_0[0]));
	jspl jspl_w_n3145_0(.douta(w_n3145_0[0]),.doutb(w_n3145_0[1]),.din(n3145));
	jspl3 jspl3_w_n3147_0(.douta(w_n3147_0[0]),.doutb(w_n3147_0[1]),.doutc(w_n3147_0[2]),.din(n3147));
	jspl3 jspl3_w_n3147_1(.douta(w_n3147_1[0]),.doutb(w_n3147_1[1]),.doutc(w_n3147_1[2]),.din(w_n3147_0[0]));
	jspl jspl_w_n3148_0(.douta(w_n3148_0[0]),.doutb(w_n3148_0[1]),.din(n3148));
	jspl jspl_w_n3150_0(.douta(w_n3150_0[0]),.doutb(w_n3150_0[1]),.din(n3150));
	jspl jspl_w_n3154_0(.douta(w_n3154_0[0]),.doutb(w_n3154_0[1]),.din(n3154));
	jspl jspl_w_n3157_0(.douta(w_n3157_0[0]),.doutb(w_n3157_0[1]),.din(n3157));
	jspl jspl_w_n3162_0(.douta(w_n3162_0[0]),.doutb(w_n3162_0[1]),.din(n3162));
	jspl jspl_w_n3165_0(.douta(w_n3165_0[0]),.doutb(w_n3165_0[1]),.din(n3165));
	jspl3 jspl3_w_n3166_0(.douta(w_n3166_0[0]),.doutb(w_n3166_0[1]),.doutc(w_n3166_0[2]),.din(n3166));
	jspl3 jspl3_w_n3166_1(.douta(w_n3166_1[0]),.doutb(w_n3166_1[1]),.doutc(w_n3166_1[2]),.din(w_n3166_0[0]));
	jspl3 jspl3_w_n3166_2(.douta(w_n3166_2[0]),.doutb(w_n3166_2[1]),.doutc(w_n3166_2[2]),.din(w_n3166_0[1]));
	jspl3 jspl3_w_n3166_3(.douta(w_n3166_3[0]),.doutb(w_n3166_3[1]),.doutc(w_n3166_3[2]),.din(w_n3166_0[2]));
	jspl3 jspl3_w_n3166_4(.douta(w_n3166_4[0]),.doutb(w_n3166_4[1]),.doutc(w_n3166_4[2]),.din(w_n3166_1[0]));
	jspl3 jspl3_w_n3166_5(.douta(w_n3166_5[0]),.doutb(w_n3166_5[1]),.doutc(w_n3166_5[2]),.din(w_n3166_1[1]));
	jspl3 jspl3_w_n3166_6(.douta(w_n3166_6[0]),.doutb(w_n3166_6[1]),.doutc(w_n3166_6[2]),.din(w_n3166_1[2]));
	jspl3 jspl3_w_n3166_7(.douta(w_n3166_7[0]),.doutb(w_n3166_7[1]),.doutc(w_n3166_7[2]),.din(w_n3166_2[0]));
	jspl3 jspl3_w_n3166_8(.douta(w_n3166_8[0]),.doutb(w_n3166_8[1]),.doutc(w_n3166_8[2]),.din(w_n3166_2[1]));
	jspl jspl_w_n3169_0(.douta(w_n3169_0[0]),.doutb(w_n3169_0[1]),.din(n3169));
	jspl jspl_w_n3171_0(.douta(w_n3171_0[0]),.doutb(w_n3171_0[1]),.din(n3171));
	jspl jspl_w_n3174_0(.douta(w_n3174_0[0]),.doutb(w_n3174_0[1]),.din(n3174));
	jspl jspl_w_n3177_0(.douta(w_n3177_0[0]),.doutb(w_n3177_0[1]),.din(n3177));
	jspl3 jspl3_w_n3179_0(.douta(w_n3179_0[0]),.doutb(w_n3179_0[1]),.doutc(w_n3179_0[2]),.din(n3179));
	jspl jspl_w_n3185_0(.douta(w_n3185_0[0]),.doutb(w_n3185_0[1]),.din(n3185));
	jspl3 jspl3_w_n3190_0(.douta(w_n3190_0[0]),.doutb(w_n3190_0[1]),.doutc(w_n3190_0[2]),.din(n3190));
	jspl3 jspl3_w_n3191_0(.douta(w_n3191_0[0]),.doutb(w_n3191_0[1]),.doutc(w_n3191_0[2]),.din(n3191));
	jspl jspl_w_n3194_0(.douta(w_n3194_0[0]),.doutb(w_n3194_0[1]),.din(n3194));
	jspl jspl_w_n3200_0(.douta(w_n3200_0[0]),.doutb(w_n3200_0[1]),.din(n3200));
	jspl3 jspl3_w_n3201_0(.douta(w_n3201_0[0]),.doutb(w_n3201_0[1]),.doutc(w_n3201_0[2]),.din(n3201));
	jspl jspl_w_n3202_0(.douta(w_n3202_0[0]),.doutb(w_n3202_0[1]),.din(n3202));
	jspl3 jspl3_w_n3203_0(.douta(w_n3203_0[0]),.doutb(w_n3203_0[1]),.doutc(w_n3203_0[2]),.din(n3203));
	jspl3 jspl3_w_n3203_1(.douta(w_n3203_1[0]),.doutb(w_n3203_1[1]),.doutc(w_n3203_1[2]),.din(w_n3203_0[0]));
	jspl3 jspl3_w_n3203_2(.douta(w_n3203_2[0]),.doutb(w_n3203_2[1]),.doutc(w_n3203_2[2]),.din(w_n3203_0[1]));
	jspl3 jspl3_w_n3203_3(.douta(w_n3203_3[0]),.doutb(w_n3203_3[1]),.doutc(w_n3203_3[2]),.din(w_n3203_0[2]));
	jspl3 jspl3_w_n3203_4(.douta(w_n3203_4[0]),.doutb(w_n3203_4[1]),.doutc(w_n3203_4[2]),.din(w_n3203_1[0]));
	jspl3 jspl3_w_n3203_5(.douta(w_n3203_5[0]),.doutb(w_n3203_5[1]),.doutc(w_n3203_5[2]),.din(w_n3203_1[1]));
	jspl3 jspl3_w_n3203_6(.douta(w_n3203_6[0]),.doutb(w_n3203_6[1]),.doutc(w_n3203_6[2]),.din(w_n3203_1[2]));
	jspl3 jspl3_w_n3203_7(.douta(w_n3203_7[0]),.doutb(w_n3203_7[1]),.doutc(w_n3203_7[2]),.din(w_n3203_2[0]));
	jspl jspl_w_n3203_8(.douta(w_n3203_8[0]),.doutb(w_n3203_8[1]),.din(w_n3203_2[1]));
	jspl jspl_w_n3204_0(.douta(w_n3204_0[0]),.doutb(w_n3204_0[1]),.din(n3204));
	jspl3 jspl3_w_n3205_0(.douta(w_n3205_0[0]),.doutb(w_n3205_0[1]),.doutc(w_n3205_0[2]),.din(n3205));
	jspl3 jspl3_w_n3205_1(.douta(w_n3205_1[0]),.doutb(w_n3205_1[1]),.doutc(w_n3205_1[2]),.din(w_n3205_0[0]));
	jspl jspl_w_n3207_0(.douta(w_n3207_0[0]),.doutb(w_n3207_0[1]),.din(n3207));
	jspl3 jspl3_w_n3209_0(.douta(w_n3209_0[0]),.doutb(w_n3209_0[1]),.doutc(w_n3209_0[2]),.din(n3209));
	jspl3 jspl3_w_n3210_0(.douta(w_n3210_0[0]),.doutb(w_n3210_0[1]),.doutc(w_n3210_0[2]),.din(n3210));
	jspl3 jspl3_w_n3210_1(.douta(w_n3210_1[0]),.doutb(w_n3210_1[1]),.doutc(w_n3210_1[2]),.din(w_n3210_0[0]));
	jspl3 jspl3_w_n3210_2(.douta(w_n3210_2[0]),.doutb(w_n3210_2[1]),.doutc(w_n3210_2[2]),.din(w_n3210_0[1]));
	jspl3 jspl3_w_n3210_3(.douta(w_n3210_3[0]),.doutb(w_n3210_3[1]),.doutc(w_n3210_3[2]),.din(w_n3210_0[2]));
	jspl3 jspl3_w_n3210_4(.douta(w_n3210_4[0]),.doutb(w_n3210_4[1]),.doutc(w_n3210_4[2]),.din(w_n3210_1[0]));
	jspl3 jspl3_w_n3210_5(.douta(w_n3210_5[0]),.doutb(w_n3210_5[1]),.doutc(w_n3210_5[2]),.din(w_n3210_1[1]));
	jspl3 jspl3_w_n3210_6(.douta(w_n3210_6[0]),.doutb(w_n3210_6[1]),.doutc(w_n3210_6[2]),.din(w_n3210_1[2]));
	jspl3 jspl3_w_n3210_7(.douta(w_n3210_7[0]),.doutb(w_n3210_7[1]),.doutc(w_n3210_7[2]),.din(w_n3210_2[0]));
	jspl3 jspl3_w_n3212_0(.douta(w_n3212_0[0]),.doutb(w_n3212_0[1]),.doutc(w_n3212_0[2]),.din(n3212));
	jspl3 jspl3_w_n3213_0(.douta(w_n3213_0[0]),.doutb(w_n3213_0[1]),.doutc(w_n3213_0[2]),.din(n3213));
	jspl3 jspl3_w_n3213_1(.douta(w_n3213_1[0]),.doutb(w_n3213_1[1]),.doutc(w_n3213_1[2]),.din(w_n3213_0[0]));
	jspl3 jspl3_w_n3213_2(.douta(w_n3213_2[0]),.doutb(w_n3213_2[1]),.doutc(w_n3213_2[2]),.din(w_n3213_0[1]));
	jspl3 jspl3_w_n3213_3(.douta(w_n3213_3[0]),.doutb(w_n3213_3[1]),.doutc(w_n3213_3[2]),.din(w_n3213_0[2]));
	jspl3 jspl3_w_n3213_4(.douta(w_n3213_4[0]),.doutb(w_n3213_4[1]),.doutc(w_n3213_4[2]),.din(w_n3213_1[0]));
	jspl3 jspl3_w_n3213_5(.douta(w_n3213_5[0]),.doutb(w_n3213_5[1]),.doutc(w_n3213_5[2]),.din(w_n3213_1[1]));
	jspl3 jspl3_w_n3213_6(.douta(w_n3213_6[0]),.doutb(w_n3213_6[1]),.doutc(w_n3213_6[2]),.din(w_n3213_1[2]));
	jspl jspl_w_n3213_7(.douta(w_n3213_7[0]),.doutb(w_n3213_7[1]),.din(w_n3213_2[0]));
	jspl3 jspl3_w_n3216_0(.douta(w_n3216_0[0]),.doutb(w_n3216_0[1]),.doutc(w_n3216_0[2]),.din(n3216));
	jspl3 jspl3_w_n3216_1(.douta(w_n3216_1[0]),.doutb(w_n3216_1[1]),.doutc(w_n3216_1[2]),.din(w_n3216_0[0]));
	jspl3 jspl3_w_n3216_2(.douta(w_n3216_2[0]),.doutb(w_n3216_2[1]),.doutc(w_n3216_2[2]),.din(w_n3216_0[1]));
	jspl3 jspl3_w_n3216_3(.douta(w_n3216_3[0]),.doutb(w_n3216_3[1]),.doutc(w_n3216_3[2]),.din(w_n3216_0[2]));
	jspl3 jspl3_w_n3216_4(.douta(w_n3216_4[0]),.doutb(w_n3216_4[1]),.doutc(w_n3216_4[2]),.din(w_n3216_1[0]));
	jspl3 jspl3_w_n3216_5(.douta(w_n3216_5[0]),.doutb(w_n3216_5[1]),.doutc(w_n3216_5[2]),.din(w_n3216_1[1]));
	jspl3 jspl3_w_n3216_6(.douta(w_n3216_6[0]),.doutb(w_n3216_6[1]),.doutc(w_n3216_6[2]),.din(w_n3216_1[2]));
	jspl3 jspl3_w_n3216_7(.douta(w_n3216_7[0]),.doutb(w_n3216_7[1]),.doutc(w_n3216_7[2]),.din(w_n3216_2[0]));
	jspl3 jspl3_w_n3218_0(.douta(w_n3218_0[0]),.doutb(w_n3218_0[1]),.doutc(w_n3218_0[2]),.din(n3218));
	jspl3 jspl3_w_n3219_0(.douta(w_n3219_0[0]),.doutb(w_n3219_0[1]),.doutc(w_n3219_0[2]),.din(n3219));
	jspl3 jspl3_w_n3219_1(.douta(w_n3219_1[0]),.doutb(w_n3219_1[1]),.doutc(w_n3219_1[2]),.din(w_n3219_0[0]));
	jspl3 jspl3_w_n3219_2(.douta(w_n3219_2[0]),.doutb(w_n3219_2[1]),.doutc(w_n3219_2[2]),.din(w_n3219_0[1]));
	jspl3 jspl3_w_n3219_3(.douta(w_n3219_3[0]),.doutb(w_n3219_3[1]),.doutc(w_n3219_3[2]),.din(w_n3219_0[2]));
	jspl3 jspl3_w_n3219_4(.douta(w_n3219_4[0]),.doutb(w_n3219_4[1]),.doutc(w_n3219_4[2]),.din(w_n3219_1[0]));
	jspl3 jspl3_w_n3219_5(.douta(w_n3219_5[0]),.doutb(w_n3219_5[1]),.doutc(w_n3219_5[2]),.din(w_n3219_1[1]));
	jspl3 jspl3_w_n3219_6(.douta(w_n3219_6[0]),.doutb(w_n3219_6[1]),.doutc(w_n3219_6[2]),.din(w_n3219_1[2]));
	jspl3 jspl3_w_n3219_7(.douta(w_n3219_7[0]),.doutb(w_n3219_7[1]),.doutc(w_n3219_7[2]),.din(w_n3219_2[0]));
	jspl jspl_w_n3223_0(.douta(w_n3223_0[0]),.doutb(w_n3223_0[1]),.din(n3223));
	jspl jspl_w_n3227_0(.douta(w_n3227_0[0]),.doutb(w_n3227_0[1]),.din(n3227));
	jspl jspl_w_n3228_0(.douta(w_n3228_0[0]),.doutb(w_n3228_0[1]),.din(n3228));
	jspl3 jspl3_w_n3229_0(.douta(w_n3229_0[0]),.doutb(w_n3229_0[1]),.doutc(w_n3229_0[2]),.din(n3229));
	jspl3 jspl3_w_n3229_1(.douta(w_n3229_1[0]),.doutb(w_n3229_1[1]),.doutc(w_n3229_1[2]),.din(w_n3229_0[0]));
	jspl jspl_w_n3237_0(.douta(w_n3237_0[0]),.doutb(w_n3237_0[1]),.din(n3237));
	jspl jspl_w_n3240_0(.douta(w_n3240_0[0]),.doutb(w_n3240_0[1]),.din(n3240));
	jspl jspl_w_n3241_0(.douta(w_n3241_0[0]),.doutb(w_n3241_0[1]),.din(n3241));
	jspl3 jspl3_w_n3242_0(.douta(w_n3242_0[0]),.doutb(w_n3242_0[1]),.doutc(w_n3242_0[2]),.din(n3242));
	jspl3 jspl3_w_n3242_1(.douta(w_n3242_1[0]),.doutb(w_n3242_1[1]),.doutc(w_n3242_1[2]),.din(w_n3242_0[0]));
	jspl jspl_w_n3250_0(.douta(w_n3250_0[0]),.doutb(w_n3250_0[1]),.din(n3250));
	jspl jspl_w_n3252_0(.douta(w_n3252_0[0]),.doutb(w_n3252_0[1]),.din(n3252));
	jspl jspl_w_n3260_0(.douta(w_n3260_0[0]),.doutb(w_n3260_0[1]),.din(n3260));
	jspl jspl_w_n3262_0(.douta(w_n3262_0[0]),.doutb(w_n3262_0[1]),.din(n3262));
	jspl jspl_w_n3270_0(.douta(w_n3270_0[0]),.doutb(w_n3270_0[1]),.din(n3270));
	jspl jspl_w_n3272_0(.douta(w_n3272_0[0]),.doutb(w_n3272_0[1]),.din(n3272));
	jspl jspl_w_n3280_0(.douta(w_n3280_0[0]),.doutb(w_n3280_0[1]),.din(n3280));
	jspl jspl_w_n3289_0(.douta(w_n3289_0[0]),.doutb(w_n3289_0[1]),.din(n3289));
	jspl jspl_w_n3292_0(.douta(w_n3292_0[0]),.doutb(w_n3292_0[1]),.din(n3292));
	jspl jspl_w_n3301_0(.douta(w_n3301_0[0]),.doutb(w_n3301_0[1]),.din(n3301));
	jspl jspl_w_n3304_0(.douta(w_n3304_0[0]),.doutb(w_n3304_0[1]),.din(n3304));
	jspl jspl_w_n3311_0(.douta(w_n3311_0[0]),.doutb(w_n3311_0[1]),.din(n3311));
	jspl3 jspl3_w_n3312_0(.douta(w_n3312_0[0]),.doutb(w_n3312_0[1]),.doutc(w_n3312_0[2]),.din(n3312));
	jspl jspl_w_n3315_0(.douta(w_n3315_0[0]),.doutb(w_n3315_0[1]),.din(n3315));
	jspl jspl_w_n3323_0(.douta(w_n3323_0[0]),.doutb(w_n3323_0[1]),.din(n3323));
	jspl jspl_w_n3324_0(.douta(w_n3324_0[0]),.doutb(w_n3324_0[1]),.din(n3324));
	jspl jspl_w_n3326_0(.douta(w_n3326_0[0]),.doutb(w_n3326_0[1]),.din(n3326));
	jspl jspl_w_n3334_0(.douta(w_n3334_0[0]),.doutb(w_n3334_0[1]),.din(n3334));
	jspl jspl_w_n3337_0(.douta(w_n3337_0[0]),.doutb(w_n3337_0[1]),.din(n3337));
	jspl jspl_w_n3338_0(.douta(w_n3338_0[0]),.doutb(w_n3338_0[1]),.din(n3338));
	jspl jspl_w_n3341_0(.douta(w_n3341_0[0]),.doutb(w_n3341_0[1]),.din(n3341));
	jspl jspl_w_n3343_0(.douta(w_n3343_0[0]),.doutb(w_n3343_0[1]),.din(n3343));
	jspl jspl_w_n3345_0(.douta(w_n3345_0[0]),.doutb(w_n3345_0[1]),.din(n3345));
	jspl jspl_w_n3346_0(.douta(w_n3346_0[0]),.doutb(w_n3346_0[1]),.din(n3346));
	jspl jspl_w_n3348_0(.douta(w_n3348_0[0]),.doutb(w_n3348_0[1]),.din(n3348));
	jspl jspl_w_n3349_0(.douta(w_n3349_0[0]),.doutb(w_n3349_0[1]),.din(n3349));
	jspl jspl_w_n3351_0(.douta(w_n3351_0[0]),.doutb(w_n3351_0[1]),.din(n3351));
	jspl jspl_w_n3352_0(.douta(w_n3352_0[0]),.doutb(w_n3352_0[1]),.din(n3352));
	jspl jspl_w_n3354_0(.douta(w_n3354_0[0]),.doutb(w_n3354_0[1]),.din(n3354));
	jspl jspl_w_n3355_0(.douta(w_n3355_0[0]),.doutb(w_n3355_0[1]),.din(n3355));
	jspl jspl_w_n3357_0(.douta(w_n3357_0[0]),.doutb(w_n3357_0[1]),.din(n3357));
	jspl jspl_w_n3358_0(.douta(w_n3358_0[0]),.doutb(w_n3358_0[1]),.din(n3358));
	jspl jspl_w_n3360_0(.douta(w_n3360_0[0]),.doutb(w_n3360_0[1]),.din(n3360));
	jspl jspl_w_n3361_0(.douta(w_n3361_0[0]),.doutb(w_n3361_0[1]),.din(n3361));
	jspl jspl_w_n3363_0(.douta(w_n3363_0[0]),.doutb(w_n3363_0[1]),.din(n3363));
	jspl jspl_w_n3368_0(.douta(w_n3368_0[0]),.doutb(w_n3368_0[1]),.din(n3368));
	jspl jspl_w_n3371_0(.douta(w_n3371_0[0]),.doutb(w_n3371_0[1]),.din(n3371));
	jspl jspl_w_n3380_0(.douta(w_n3380_0[0]),.doutb(w_n3380_0[1]),.din(n3380));
	jspl jspl_w_n3381_0(.douta(w_n3381_0[0]),.doutb(w_n3381_0[1]),.din(n3381));
	jspl jspl_w_n3382_0(.douta(w_n3382_0[0]),.doutb(w_n3382_0[1]),.din(n3382));
	jspl3 jspl3_w_n3384_0(.douta(w_n3384_0[0]),.doutb(w_n3384_0[1]),.doutc(w_n3384_0[2]),.din(n3384));
	jspl3 jspl3_w_n3384_1(.douta(w_n3384_1[0]),.doutb(w_n3384_1[1]),.doutc(w_n3384_1[2]),.din(w_n3384_0[0]));
	jspl3 jspl3_w_n3384_2(.douta(w_n3384_2[0]),.doutb(w_n3384_2[1]),.doutc(w_n3384_2[2]),.din(w_n3384_0[1]));
	jspl3 jspl3_w_n3384_3(.douta(w_n3384_3[0]),.doutb(w_n3384_3[1]),.doutc(w_n3384_3[2]),.din(w_n3384_0[2]));
	jspl3 jspl3_w_n3384_4(.douta(w_n3384_4[0]),.doutb(w_n3384_4[1]),.doutc(w_n3384_4[2]),.din(w_n3384_1[0]));
	jspl3 jspl3_w_n3384_5(.douta(w_n3384_5[0]),.doutb(w_n3384_5[1]),.doutc(w_n3384_5[2]),.din(w_n3384_1[1]));
	jspl3 jspl3_w_n3384_6(.douta(w_n3384_6[0]),.doutb(w_n3384_6[1]),.doutc(w_n3384_6[2]),.din(w_n3384_1[2]));
	jspl jspl_w_n3384_7(.douta(w_n3384_7[0]),.doutb(w_n3384_7[1]),.din(w_n3384_2[0]));
	jspl3 jspl3_w_n3386_0(.douta(w_n3386_0[0]),.doutb(w_n3386_0[1]),.doutc(w_n3386_0[2]),.din(n3386));
	jspl3 jspl3_w_n3386_1(.douta(w_n3386_1[0]),.doutb(w_n3386_1[1]),.doutc(w_n3386_1[2]),.din(w_n3386_0[0]));
	jspl3 jspl3_w_n3386_2(.douta(w_n3386_2[0]),.doutb(w_n3386_2[1]),.doutc(w_n3386_2[2]),.din(w_n3386_0[1]));
	jspl3 jspl3_w_n3386_3(.douta(w_n3386_3[0]),.doutb(w_n3386_3[1]),.doutc(w_n3386_3[2]),.din(w_n3386_0[2]));
	jspl jspl_w_n3386_4(.douta(w_n3386_4[0]),.doutb(w_n3386_4[1]),.din(w_n3386_1[0]));
	jspl3 jspl3_w_n3388_0(.douta(w_n3388_0[0]),.doutb(w_n3388_0[1]),.doutc(w_n3388_0[2]),.din(n3388));
	jspl3 jspl3_w_n3388_1(.douta(w_n3388_1[0]),.doutb(w_n3388_1[1]),.doutc(w_n3388_1[2]),.din(w_n3388_0[0]));
	jspl3 jspl3_w_n3388_2(.douta(w_n3388_2[0]),.doutb(w_n3388_2[1]),.doutc(w_n3388_2[2]),.din(w_n3388_0[1]));
	jspl3 jspl3_w_n3388_3(.douta(w_n3388_3[0]),.doutb(w_n3388_3[1]),.doutc(w_n3388_3[2]),.din(w_n3388_0[2]));
	jspl3 jspl3_w_n3388_4(.douta(w_n3388_4[0]),.doutb(w_n3388_4[1]),.doutc(w_n3388_4[2]),.din(w_n3388_1[0]));
	jspl3 jspl3_w_n3390_0(.douta(w_n3390_0[0]),.doutb(w_n3390_0[1]),.doutc(w_n3390_0[2]),.din(n3390));
	jspl3 jspl3_w_n3390_1(.douta(w_n3390_1[0]),.doutb(w_n3390_1[1]),.doutc(w_n3390_1[2]),.din(w_n3390_0[0]));
	jspl3 jspl3_w_n3390_2(.douta(w_n3390_2[0]),.doutb(w_n3390_2[1]),.doutc(w_n3390_2[2]),.din(w_n3390_0[1]));
	jspl3 jspl3_w_n3390_3(.douta(w_n3390_3[0]),.doutb(w_n3390_3[1]),.doutc(w_n3390_3[2]),.din(w_n3390_0[2]));
	jspl3 jspl3_w_n3390_4(.douta(w_n3390_4[0]),.doutb(w_n3390_4[1]),.doutc(w_n3390_4[2]),.din(w_n3390_1[0]));
	jspl jspl_w_n3395_0(.douta(w_n3395_0[0]),.doutb(w_n3395_0[1]),.din(n3395));
	jspl jspl_w_n3396_0(.douta(w_n3396_0[0]),.doutb(w_n3396_0[1]),.din(n3396));
	jspl jspl_w_n3397_0(.douta(w_n3397_0[0]),.doutb(w_n3397_0[1]),.din(n3397));
	jspl jspl_w_n3399_0(.douta(w_n3399_0[0]),.doutb(w_n3399_0[1]),.din(n3399));
	jspl jspl_w_n3407_0(.douta(w_n3407_0[0]),.doutb(w_n3407_0[1]),.din(n3407));
	jspl jspl_w_n3408_0(.douta(w_n3408_0[0]),.doutb(w_n3408_0[1]),.din(n3408));
	jspl jspl_w_n3409_0(.douta(w_n3409_0[0]),.doutb(w_n3409_0[1]),.din(n3409));
	jspl jspl_w_n3414_0(.douta(w_n3414_0[0]),.doutb(w_n3414_0[1]),.din(n3414));
	jspl3 jspl3_w_n3415_0(.douta(w_n3415_0[0]),.doutb(w_n3415_0[1]),.doutc(w_n3415_0[2]),.din(n3415));
	jspl jspl_w_n3415_1(.douta(w_n3415_1[0]),.doutb(w_n3415_1[1]),.din(w_n3415_0[0]));
	jspl jspl_w_n3416_0(.douta(w_n3416_0[0]),.doutb(w_n3416_0[1]),.din(n3416));
	jspl jspl_w_n3418_0(.douta(w_n3418_0[0]),.doutb(w_n3418_0[1]),.din(n3418));
	jspl jspl_w_n3420_0(.douta(w_n3420_0[0]),.doutb(w_n3420_0[1]),.din(n3420));
	jspl jspl_w_n3429_0(.douta(w_n3429_0[0]),.doutb(w_n3429_0[1]),.din(n3429));
	jspl3 jspl3_w_n3435_0(.douta(w_n3435_0[0]),.doutb(w_n3435_0[1]),.doutc(w_n3435_0[2]),.din(n3435));
	jspl jspl_w_n3440_0(.douta(w_n3440_0[0]),.doutb(w_n3440_0[1]),.din(n3440));
	jspl3 jspl3_w_n3441_0(.douta(w_n3441_0[0]),.doutb(w_n3441_0[1]),.doutc(w_n3441_0[2]),.din(n3441));
	jspl3 jspl3_w_n3441_1(.douta(w_n3441_1[0]),.doutb(w_n3441_1[1]),.doutc(w_n3441_1[2]),.din(w_n3441_0[0]));
	jspl3 jspl3_w_n3441_2(.douta(w_n3441_2[0]),.doutb(w_n3441_2[1]),.doutc(w_n3441_2[2]),.din(w_n3441_0[1]));
	jspl3 jspl3_w_n3441_3(.douta(w_n3441_3[0]),.doutb(w_n3441_3[1]),.doutc(w_n3441_3[2]),.din(w_n3441_0[2]));
	jspl3 jspl3_w_n3441_4(.douta(w_n3441_4[0]),.doutb(w_n3441_4[1]),.doutc(w_n3441_4[2]),.din(w_n3441_1[0]));
	jspl3 jspl3_w_n3441_5(.douta(w_n3441_5[0]),.doutb(w_n3441_5[1]),.doutc(w_n3441_5[2]),.din(w_n3441_1[1]));
	jspl3 jspl3_w_n3441_6(.douta(w_n3441_6[0]),.doutb(w_n3441_6[1]),.doutc(w_n3441_6[2]),.din(w_n3441_1[2]));
	jspl3 jspl3_w_n3441_7(.douta(w_n3441_7[0]),.doutb(w_n3441_7[1]),.doutc(w_n3441_7[2]),.din(w_n3441_2[0]));
	jspl jspl_w_n3442_0(.douta(w_n3442_0[0]),.doutb(w_n3442_0[1]),.din(n3442));
	jspl3 jspl3_w_n3443_0(.douta(w_n3443_0[0]),.doutb(w_n3443_0[1]),.doutc(w_n3443_0[2]),.din(n3443));
	jspl3 jspl3_w_n3443_1(.douta(w_n3443_1[0]),.doutb(w_n3443_1[1]),.doutc(w_n3443_1[2]),.din(w_n3443_0[0]));
	jspl jspl_w_n3451_0(.douta(w_n3451_0[0]),.doutb(w_n3451_0[1]),.din(n3451));
	jspl jspl_w_n3452_0(.douta(w_n3452_0[0]),.doutb(w_n3452_0[1]),.din(n3452));
	jspl jspl_w_n3454_0(.douta(w_n3454_0[0]),.doutb(w_n3454_0[1]),.din(n3454));
	jspl3 jspl3_w_n3455_0(.douta(w_n3455_0[0]),.doutb(w_n3455_0[1]),.doutc(w_n3455_0[2]),.din(n3455));
	jspl3 jspl3_w_n3455_1(.douta(w_n3455_1[0]),.doutb(w_n3455_1[1]),.doutc(w_n3455_1[2]),.din(w_n3455_0[0]));
	jspl3 jspl3_w_n3455_2(.douta(w_n3455_2[0]),.doutb(w_n3455_2[1]),.doutc(w_n3455_2[2]),.din(w_n3455_0[1]));
	jspl3 jspl3_w_n3455_3(.douta(w_n3455_3[0]),.doutb(w_n3455_3[1]),.doutc(w_n3455_3[2]),.din(w_n3455_0[2]));
	jspl3 jspl3_w_n3455_4(.douta(w_n3455_4[0]),.doutb(w_n3455_4[1]),.doutc(w_n3455_4[2]),.din(w_n3455_1[0]));
	jspl3 jspl3_w_n3456_0(.douta(w_n3456_0[0]),.doutb(w_n3456_0[1]),.doutc(w_n3456_0[2]),.din(n3456));
	jspl jspl_w_n3459_0(.douta(w_n3459_0[0]),.doutb(w_n3459_0[1]),.din(n3459));
	jspl3 jspl3_w_n3460_0(.douta(w_n3460_0[0]),.doutb(w_n3460_0[1]),.doutc(w_n3460_0[2]),.din(n3460));
	jspl3 jspl3_w_n3461_0(.douta(w_n3461_0[0]),.doutb(w_n3461_0[1]),.doutc(w_n3461_0[2]),.din(n3461));
	jspl3 jspl3_w_n3461_1(.douta(w_n3461_1[0]),.doutb(w_n3461_1[1]),.doutc(w_n3461_1[2]),.din(w_n3461_0[0]));
	jspl3 jspl3_w_n3461_2(.douta(w_n3461_2[0]),.doutb(w_n3461_2[1]),.doutc(w_n3461_2[2]),.din(w_n3461_0[1]));
	jspl3 jspl3_w_n3461_3(.douta(w_n3461_3[0]),.doutb(w_n3461_3[1]),.doutc(w_n3461_3[2]),.din(w_n3461_0[2]));
	jspl3 jspl3_w_n3461_4(.douta(w_n3461_4[0]),.doutb(w_n3461_4[1]),.doutc(w_n3461_4[2]),.din(w_n3461_1[0]));
	jspl3 jspl3_w_n3461_5(.douta(w_n3461_5[0]),.doutb(w_n3461_5[1]),.doutc(w_n3461_5[2]),.din(w_n3461_1[1]));
	jspl3 jspl3_w_n3461_6(.douta(w_n3461_6[0]),.doutb(w_n3461_6[1]),.doutc(w_n3461_6[2]),.din(w_n3461_1[2]));
	jspl3 jspl3_w_n3461_7(.douta(w_n3461_7[0]),.doutb(w_n3461_7[1]),.doutc(w_n3461_7[2]),.din(w_n3461_2[0]));
	jspl3 jspl3_w_n3461_8(.douta(w_n3461_8[0]),.doutb(w_n3461_8[1]),.doutc(w_n3461_8[2]),.din(w_n3461_2[1]));
	jspl jspl_w_n3463_0(.douta(w_n3463_0[0]),.doutb(w_n3463_0[1]),.din(n3463));
	jspl3 jspl3_w_n3468_0(.douta(w_n3468_0[0]),.doutb(w_n3468_0[1]),.doutc(w_n3468_0[2]),.din(n3468));
	jspl3 jspl3_w_n3470_0(.douta(w_n3470_0[0]),.doutb(w_n3470_0[1]),.doutc(w_n3470_0[2]),.din(n3470));
	jspl3 jspl3_w_n3481_0(.douta(w_n3481_0[0]),.doutb(w_n3481_0[1]),.doutc(w_n3481_0[2]),.din(n3481));
	jspl jspl_w_n3488_0(.douta(w_n3488_0[0]),.doutb(w_n3488_0[1]),.din(n3488));
	jspl jspl_w_n3489_0(.douta(w_n3489_0[0]),.doutb(w_n3489_0[1]),.din(n3489));
	jspl3 jspl3_w_n3494_0(.douta(w_n3494_0[0]),.doutb(w_n3494_0[1]),.doutc(w_n3494_0[2]),.din(n3494));
	jspl3 jspl3_w_n3495_0(.douta(w_n3495_0[0]),.doutb(w_n3495_0[1]),.doutc(w_n3495_0[2]),.din(n3495));
	jspl3 jspl3_w_n3495_1(.douta(w_n3495_1[0]),.doutb(w_n3495_1[1]),.doutc(w_n3495_1[2]),.din(w_n3495_0[0]));
	jspl3 jspl3_w_n3495_2(.douta(w_n3495_2[0]),.doutb(w_n3495_2[1]),.doutc(w_n3495_2[2]),.din(w_n3495_0[1]));
	jspl3 jspl3_w_n3495_3(.douta(w_n3495_3[0]),.doutb(w_n3495_3[1]),.doutc(w_n3495_3[2]),.din(w_n3495_0[2]));
	jspl3 jspl3_w_n3495_4(.douta(w_n3495_4[0]),.doutb(w_n3495_4[1]),.doutc(w_n3495_4[2]),.din(w_n3495_1[0]));
	jspl3 jspl3_w_n3495_5(.douta(w_n3495_5[0]),.doutb(w_n3495_5[1]),.doutc(w_n3495_5[2]),.din(w_n3495_1[1]));
	jspl3 jspl3_w_n3495_6(.douta(w_n3495_6[0]),.doutb(w_n3495_6[1]),.doutc(w_n3495_6[2]),.din(w_n3495_1[2]));
	jspl3 jspl3_w_n3495_7(.douta(w_n3495_7[0]),.doutb(w_n3495_7[1]),.doutc(w_n3495_7[2]),.din(w_n3495_2[0]));
	jspl jspl_w_n3495_8(.douta(w_n3495_8[0]),.doutb(w_n3495_8[1]),.din(w_n3495_2[1]));
	jspl jspl_w_n3496_0(.douta(w_n3496_0[0]),.doutb(w_n3496_0[1]),.din(n3496));
	jspl3 jspl3_w_n3497_0(.douta(w_n3497_0[0]),.doutb(w_n3497_0[1]),.doutc(w_n3497_0[2]),.din(n3497));
	jspl3 jspl3_w_n3509_0(.douta(w_n3509_0[0]),.doutb(w_n3509_0[1]),.doutc(w_n3509_0[2]),.din(n3509));
	jspl3 jspl3_w_n3510_0(.douta(w_n3510_0[0]),.doutb(w_n3510_0[1]),.doutc(w_n3510_0[2]),.din(n3510));
	jspl3 jspl3_w_n3510_1(.douta(w_n3510_1[0]),.doutb(w_n3510_1[1]),.doutc(w_n3510_1[2]),.din(w_n3510_0[0]));
	jspl3 jspl3_w_n3510_2(.douta(w_n3510_2[0]),.doutb(w_n3510_2[1]),.doutc(w_n3510_2[2]),.din(w_n3510_0[1]));
	jspl3 jspl3_w_n3510_3(.douta(w_n3510_3[0]),.doutb(w_n3510_3[1]),.doutc(w_n3510_3[2]),.din(w_n3510_0[2]));
	jspl3 jspl3_w_n3510_4(.douta(w_n3510_4[0]),.doutb(w_n3510_4[1]),.doutc(w_n3510_4[2]),.din(w_n3510_1[0]));
	jspl3 jspl3_w_n3510_5(.douta(w_n3510_5[0]),.doutb(w_n3510_5[1]),.doutc(w_n3510_5[2]),.din(w_n3510_1[1]));
	jspl3 jspl3_w_n3510_6(.douta(w_n3510_6[0]),.doutb(w_n3510_6[1]),.doutc(w_n3510_6[2]),.din(w_n3510_1[2]));
	jspl3 jspl3_w_n3510_7(.douta(w_n3510_7[0]),.doutb(w_n3510_7[1]),.doutc(w_n3510_7[2]),.din(w_n3510_2[0]));
	jspl3 jspl3_w_n3510_8(.douta(w_n3510_8[0]),.doutb(w_n3510_8[1]),.doutc(w_n3510_8[2]),.din(w_n3510_2[1]));
	jspl3 jspl3_w_n3511_0(.douta(w_n3511_0[0]),.doutb(w_n3511_0[1]),.doutc(w_n3511_0[2]),.din(n3511));
	jspl jspl_w_n3512_0(.douta(w_n3512_0[0]),.doutb(w_n3512_0[1]),.din(n3512));
	jspl3 jspl3_w_n3513_0(.douta(w_n3513_0[0]),.doutb(w_n3513_0[1]),.doutc(w_n3513_0[2]),.din(n3513));
	jspl3 jspl3_w_n3513_1(.douta(w_n3513_1[0]),.doutb(w_n3513_1[1]),.doutc(w_n3513_1[2]),.din(w_n3513_0[0]));
	jspl jspl_w_n3514_0(.douta(w_n3514_0[0]),.doutb(w_n3514_0[1]),.din(n3514));
	jspl jspl_w_n3518_0(.douta(w_n3518_0[0]),.doutb(w_n3518_0[1]),.din(n3518));
	jspl jspl_w_n3519_0(.douta(w_n3519_0[0]),.doutb(w_n3519_0[1]),.din(n3519));
	jspl3 jspl3_w_n3520_0(.douta(w_n3520_0[0]),.doutb(w_n3520_0[1]),.doutc(w_n3520_0[2]),.din(n3520));
	jspl jspl_w_n3521_0(.douta(w_n3521_0[0]),.doutb(w_n3521_0[1]),.din(n3521));
	jspl jspl_w_n3522_0(.douta(w_n3522_0[0]),.doutb(w_n3522_0[1]),.din(n3522));
	jspl jspl_w_n3526_0(.douta(w_n3526_0[0]),.doutb(w_n3526_0[1]),.din(n3526));
	jspl3 jspl3_w_n3529_0(.douta(w_n3529_0[0]),.doutb(w_n3529_0[1]),.doutc(w_n3529_0[2]),.din(n3529));
	jspl jspl_w_n3532_0(.douta(w_n3532_0[0]),.doutb(w_n3532_0[1]),.din(n3532));
	jspl3 jspl3_w_n3537_0(.douta(w_n3537_0[0]),.doutb(w_n3537_0[1]),.doutc(w_n3537_0[2]),.din(n3537));
	jspl3 jspl3_w_n3537_1(.douta(w_n3537_1[0]),.doutb(w_n3537_1[1]),.doutc(w_n3537_1[2]),.din(w_n3537_0[0]));
	jspl3 jspl3_w_n3543_0(.douta(w_n3543_0[0]),.doutb(w_n3543_0[1]),.doutc(w_n3543_0[2]),.din(n3543));
	jspl jspl_w_n3546_0(.douta(w_n3546_0[0]),.doutb(w_n3546_0[1]),.din(n3546));
	jspl3 jspl3_w_n3547_0(.douta(w_n3547_0[0]),.doutb(w_n3547_0[1]),.doutc(w_n3547_0[2]),.din(n3547));
	jspl3 jspl3_w_n3547_1(.douta(w_n3547_1[0]),.doutb(w_n3547_1[1]),.doutc(w_n3547_1[2]),.din(w_n3547_0[0]));
	jspl3 jspl3_w_n3547_2(.douta(w_n3547_2[0]),.doutb(w_n3547_2[1]),.doutc(w_n3547_2[2]),.din(w_n3547_0[1]));
	jspl3 jspl3_w_n3547_3(.douta(w_n3547_3[0]),.doutb(w_n3547_3[1]),.doutc(w_n3547_3[2]),.din(w_n3547_0[2]));
	jspl3 jspl3_w_n3547_4(.douta(w_n3547_4[0]),.doutb(w_n3547_4[1]),.doutc(w_n3547_4[2]),.din(w_n3547_1[0]));
	jspl3 jspl3_w_n3547_5(.douta(w_n3547_5[0]),.doutb(w_n3547_5[1]),.doutc(w_n3547_5[2]),.din(w_n3547_1[1]));
	jspl3 jspl3_w_n3547_6(.douta(w_n3547_6[0]),.doutb(w_n3547_6[1]),.doutc(w_n3547_6[2]),.din(w_n3547_1[2]));
	jspl3 jspl3_w_n3547_7(.douta(w_n3547_7[0]),.doutb(w_n3547_7[1]),.doutc(w_n3547_7[2]),.din(w_n3547_2[0]));
	jspl3 jspl3_w_n3548_0(.douta(w_n3548_0[0]),.doutb(w_n3548_0[1]),.doutc(w_n3548_0[2]),.din(n3548));
	jspl3 jspl3_w_n3549_0(.douta(w_n3549_0[0]),.doutb(w_n3549_0[1]),.doutc(w_n3549_0[2]),.din(n3549));
	jspl3 jspl3_w_n3550_0(.douta(w_n3550_0[0]),.doutb(w_n3550_0[1]),.doutc(w_n3550_0[2]),.din(n3550));
	jspl3 jspl3_w_n3550_1(.douta(w_n3550_1[0]),.doutb(w_n3550_1[1]),.doutc(w_n3550_1[2]),.din(w_n3550_0[0]));
	jspl3 jspl3_w_n3552_0(.douta(w_n3552_0[0]),.doutb(w_n3552_0[1]),.doutc(w_n3552_0[2]),.din(n3552));
	jspl3 jspl3_w_n3552_1(.douta(w_n3552_1[0]),.doutb(w_n3552_1[1]),.doutc(w_n3552_1[2]),.din(w_n3552_0[0]));
	jspl3 jspl3_w_n3552_2(.douta(w_n3552_2[0]),.doutb(w_n3552_2[1]),.doutc(w_n3552_2[2]),.din(w_n3552_0[1]));
	jspl3 jspl3_w_n3552_3(.douta(w_n3552_3[0]),.doutb(w_n3552_3[1]),.doutc(w_n3552_3[2]),.din(w_n3552_0[2]));
	jspl3 jspl3_w_n3552_4(.douta(w_n3552_4[0]),.doutb(w_n3552_4[1]),.doutc(w_n3552_4[2]),.din(w_n3552_1[0]));
	jspl3 jspl3_w_n3552_5(.douta(w_n3552_5[0]),.doutb(w_n3552_5[1]),.doutc(w_n3552_5[2]),.din(w_n3552_1[1]));
	jspl3 jspl3_w_n3552_6(.douta(w_n3552_6[0]),.doutb(w_n3552_6[1]),.doutc(w_n3552_6[2]),.din(w_n3552_1[2]));
	jspl3 jspl3_w_n3552_7(.douta(w_n3552_7[0]),.doutb(w_n3552_7[1]),.doutc(w_n3552_7[2]),.din(w_n3552_2[0]));
	jspl3 jspl3_w_n3554_0(.douta(w_n3554_0[0]),.doutb(w_n3554_0[1]),.doutc(w_n3554_0[2]),.din(n3554));
	jspl3 jspl3_w_n3554_1(.douta(w_n3554_1[0]),.doutb(w_n3554_1[1]),.doutc(w_n3554_1[2]),.din(w_n3554_0[0]));
	jspl3 jspl3_w_n3554_2(.douta(w_n3554_2[0]),.doutb(w_n3554_2[1]),.doutc(w_n3554_2[2]),.din(w_n3554_0[1]));
	jspl3 jspl3_w_n3554_3(.douta(w_n3554_3[0]),.doutb(w_n3554_3[1]),.doutc(w_n3554_3[2]),.din(w_n3554_0[2]));
	jspl3 jspl3_w_n3554_4(.douta(w_n3554_4[0]),.doutb(w_n3554_4[1]),.doutc(w_n3554_4[2]),.din(w_n3554_1[0]));
	jspl3 jspl3_w_n3554_5(.douta(w_n3554_5[0]),.doutb(w_n3554_5[1]),.doutc(w_n3554_5[2]),.din(w_n3554_1[1]));
	jspl3 jspl3_w_n3554_6(.douta(w_n3554_6[0]),.doutb(w_n3554_6[1]),.doutc(w_n3554_6[2]),.din(w_n3554_1[2]));
	jspl3 jspl3_w_n3554_7(.douta(w_n3554_7[0]),.doutb(w_n3554_7[1]),.doutc(w_n3554_7[2]),.din(w_n3554_2[0]));
	jspl jspl_w_n3554_8(.douta(w_n3554_8[0]),.doutb(w_n3554_8[1]),.din(w_n3554_2[1]));
	jspl3 jspl3_w_n3557_0(.douta(w_n3557_0[0]),.doutb(w_n3557_0[1]),.doutc(w_n3557_0[2]),.din(n3557));
	jspl jspl_w_n3557_1(.douta(w_n3557_1[0]),.doutb(w_n3557_1[1]),.din(w_n3557_0[0]));
	jspl3 jspl3_w_n3558_0(.douta(w_n3558_0[0]),.doutb(w_n3558_0[1]),.doutc(w_n3558_0[2]),.din(n3558));
	jspl3 jspl3_w_n3558_1(.douta(w_n3558_1[0]),.doutb(w_n3558_1[1]),.doutc(w_n3558_1[2]),.din(w_n3558_0[0]));
	jspl3 jspl3_w_n3558_2(.douta(w_n3558_2[0]),.doutb(w_n3558_2[1]),.doutc(w_n3558_2[2]),.din(w_n3558_0[1]));
	jspl3 jspl3_w_n3558_3(.douta(w_n3558_3[0]),.doutb(w_n3558_3[1]),.doutc(w_n3558_3[2]),.din(w_n3558_0[2]));
	jspl3 jspl3_w_n3558_4(.douta(w_n3558_4[0]),.doutb(w_n3558_4[1]),.doutc(w_n3558_4[2]),.din(w_n3558_1[0]));
	jspl3 jspl3_w_n3558_5(.douta(w_n3558_5[0]),.doutb(w_n3558_5[1]),.doutc(w_n3558_5[2]),.din(w_n3558_1[1]));
	jspl3 jspl3_w_n3558_6(.douta(w_n3558_6[0]),.doutb(w_n3558_6[1]),.doutc(w_n3558_6[2]),.din(w_n3558_1[2]));
	jspl jspl_w_n3562_0(.douta(w_n3562_0[0]),.doutb(w_n3562_0[1]),.din(n3562));
	jspl jspl_w_n3563_0(.douta(w_n3563_0[0]),.doutb(w_n3563_0[1]),.din(n3563));
	jspl jspl_w_n3565_0(.douta(w_n3565_0[0]),.doutb(w_n3565_0[1]),.din(n3565));
	jspl3 jspl3_w_n3566_0(.douta(w_n3566_0[0]),.doutb(w_n3566_0[1]),.doutc(w_n3566_0[2]),.din(n3566));
	jspl3 jspl3_w_n3566_1(.douta(w_n3566_1[0]),.doutb(w_n3566_1[1]),.doutc(w_n3566_1[2]),.din(w_n3566_0[0]));
	jspl jspl_w_n3574_0(.douta(w_n3574_0[0]),.doutb(w_n3574_0[1]),.din(n3574));
	jspl jspl_w_n3575_0(.douta(w_n3575_0[0]),.doutb(w_n3575_0[1]),.din(n3575));
	jspl jspl_w_n3576_0(.douta(w_n3576_0[0]),.doutb(w_n3576_0[1]),.din(n3576));
	jspl jspl_w_n3577_0(.douta(w_n3577_0[0]),.doutb(w_n3577_0[1]),.din(n3577));
	jspl jspl_w_n3578_0(.douta(w_n3578_0[0]),.doutb(w_n3578_0[1]),.din(n3578));
	jspl3 jspl3_w_n3579_0(.douta(w_n3579_0[0]),.doutb(w_n3579_0[1]),.doutc(w_n3579_0[2]),.din(n3579));
	jspl3 jspl3_w_n3579_1(.douta(w_n3579_1[0]),.doutb(w_n3579_1[1]),.doutc(w_n3579_1[2]),.din(w_n3579_0[0]));
	jspl jspl_w_n3587_0(.douta(w_n3587_0[0]),.doutb(w_n3587_0[1]),.din(n3587));
	jspl jspl_w_n3588_0(.douta(w_n3588_0[0]),.doutb(w_n3588_0[1]),.din(n3588));
	jspl jspl_w_n3589_0(.douta(w_n3589_0[0]),.doutb(w_n3589_0[1]),.din(n3589));
	jspl jspl_w_n3590_0(.douta(w_n3590_0[0]),.doutb(w_n3590_0[1]),.din(n3590));
	jspl jspl_w_n3598_0(.douta(w_n3598_0[0]),.doutb(w_n3598_0[1]),.din(n3598));
	jspl jspl_w_n3599_0(.douta(w_n3599_0[0]),.doutb(w_n3599_0[1]),.din(n3599));
	jspl jspl_w_n3600_0(.douta(w_n3600_0[0]),.doutb(w_n3600_0[1]),.din(n3600));
	jspl jspl_w_n3601_0(.douta(w_n3601_0[0]),.doutb(w_n3601_0[1]),.din(n3601));
	jspl jspl_w_n3609_0(.douta(w_n3609_0[0]),.doutb(w_n3609_0[1]),.din(n3609));
	jspl jspl_w_n3610_0(.douta(w_n3610_0[0]),.doutb(w_n3610_0[1]),.din(n3610));
	jspl jspl_w_n3611_0(.douta(w_n3611_0[0]),.doutb(w_n3611_0[1]),.din(n3611));
	jspl jspl_w_n3612_0(.douta(w_n3612_0[0]),.doutb(w_n3612_0[1]),.din(n3612));
	jspl jspl_w_n3620_0(.douta(w_n3620_0[0]),.doutb(w_n3620_0[1]),.din(n3620));
	jspl jspl_w_n3621_0(.douta(w_n3621_0[0]),.doutb(w_n3621_0[1]),.din(n3621));
	jspl jspl_w_n3622_0(.douta(w_n3622_0[0]),.doutb(w_n3622_0[1]),.din(n3622));
	jspl jspl_w_n3623_0(.douta(w_n3623_0[0]),.doutb(w_n3623_0[1]),.din(n3623));
	jspl jspl_w_n3631_0(.douta(w_n3631_0[0]),.doutb(w_n3631_0[1]),.din(n3631));
	jspl jspl_w_n3632_0(.douta(w_n3632_0[0]),.doutb(w_n3632_0[1]),.din(n3632));
	jspl jspl_w_n3633_0(.douta(w_n3633_0[0]),.doutb(w_n3633_0[1]),.din(n3633));
	jspl jspl_w_n3634_0(.douta(w_n3634_0[0]),.doutb(w_n3634_0[1]),.din(n3634));
	jspl jspl_w_n3642_0(.douta(w_n3642_0[0]),.doutb(w_n3642_0[1]),.din(n3642));
	jspl jspl_w_n3643_0(.douta(w_n3643_0[0]),.doutb(w_n3643_0[1]),.din(n3643));
	jspl jspl_w_n3644_0(.douta(w_n3644_0[0]),.doutb(w_n3644_0[1]),.din(n3644));
	jspl jspl_w_n3645_0(.douta(w_n3645_0[0]),.doutb(w_n3645_0[1]),.din(n3645));
	jspl jspl_w_n3653_0(.douta(w_n3653_0[0]),.doutb(w_n3653_0[1]),.din(n3653));
	jspl jspl_w_n3654_0(.douta(w_n3654_0[0]),.doutb(w_n3654_0[1]),.din(n3654));
	jspl jspl_w_n3655_0(.douta(w_n3655_0[0]),.doutb(w_n3655_0[1]),.din(n3655));
	jspl jspl_w_n3656_0(.douta(w_n3656_0[0]),.doutb(w_n3656_0[1]),.din(n3656));
	jspl jspl_w_n3664_0(.douta(w_n3664_0[0]),.doutb(w_n3664_0[1]),.din(n3664));
	jspl jspl_w_n3665_0(.douta(w_n3665_0[0]),.doutb(w_n3665_0[1]),.din(n3665));
	jspl jspl_w_n3676_0(.douta(w_n3676_0[0]),.doutb(w_n3676_0[1]),.din(n3676));
	jspl jspl_w_n3678_0(.douta(w_n3678_0[0]),.doutb(w_n3678_0[1]),.din(n3678));
	jspl jspl_w_n3681_0(.douta(w_n3681_0[0]),.doutb(w_n3681_0[1]),.din(n3681));
	jspl jspl_w_n3682_0(.douta(w_n3682_0[0]),.doutb(w_n3682_0[1]),.din(n3682));
	jspl jspl_w_n3685_0(.douta(w_n3685_0[0]),.doutb(w_n3685_0[1]),.din(n3685));
	jspl jspl_w_n3686_0(.douta(w_n3686_0[0]),.doutb(w_n3686_0[1]),.din(n3686));
	jspl jspl_w_n3688_0(.douta(w_n3688_0[0]),.doutb(w_n3688_0[1]),.din(n3688));
	jspl jspl_w_n3695_0(.douta(w_n3695_0[0]),.doutb(w_n3695_0[1]),.din(n3695));
	jspl jspl_w_n3698_0(.douta(w_n3698_0[0]),.doutb(w_n3698_0[1]),.din(n3698));
	jspl jspl_w_n3700_0(.douta(w_n3700_0[0]),.doutb(w_n3700_0[1]),.din(n3700));
	jspl jspl_w_n3701_0(.douta(w_n3701_0[0]),.doutb(w_n3701_0[1]),.din(n3701));
	jspl jspl_w_n3702_0(.douta(w_n3702_0[0]),.doutb(w_n3702_0[1]),.din(n3702));
	jspl jspl_w_n3705_0(.douta(w_n3705_0[0]),.doutb(w_n3705_0[1]),.din(n3705));
	jspl jspl_w_n3709_0(.douta(w_n3709_0[0]),.doutb(w_n3709_0[1]),.din(n3709));
	jspl jspl_w_n3713_0(.douta(w_n3713_0[0]),.doutb(w_n3713_0[1]),.din(n3713));
	jspl jspl_w_n3714_0(.douta(w_n3714_0[0]),.doutb(w_n3714_0[1]),.din(n3714));
	jspl jspl_w_n3718_0(.douta(w_n3718_0[0]),.doutb(w_n3718_0[1]),.din(n3718));
	jspl jspl_w_n3720_0(.douta(w_n3720_0[0]),.doutb(w_n3720_0[1]),.din(n3720));
	jspl jspl_w_n3725_0(.douta(w_n3725_0[0]),.doutb(w_n3725_0[1]),.din(n3725));
	jspl3 jspl3_w_n3733_0(.douta(w_n3733_0[0]),.doutb(w_n3733_0[1]),.doutc(w_n3733_0[2]),.din(n3733));
	jspl jspl_w_n3734_0(.douta(w_n3734_0[0]),.doutb(w_n3734_0[1]),.din(n3734));
	jspl jspl_w_n3738_0(.douta(w_n3738_0[0]),.doutb(w_n3738_0[1]),.din(n3738));
	jspl jspl_w_n3742_0(.douta(w_n3742_0[0]),.doutb(w_n3742_0[1]),.din(n3742));
	jspl jspl_w_n3760_0(.douta(w_n3760_0[0]),.doutb(w_n3760_0[1]),.din(n3760));
	jspl3 jspl3_w_n3761_0(.douta(w_n3761_0[0]),.doutb(w_n3761_0[1]),.doutc(w_n3761_0[2]),.din(n3761));
	jspl jspl_w_n3763_0(.douta(w_n3763_0[0]),.doutb(w_n3763_0[1]),.din(n3763));
	jspl jspl_w_n3766_0(.douta(w_n3766_0[0]),.doutb(w_n3766_0[1]),.din(n3766));
	jspl jspl_w_n3770_0(.douta(w_n3770_0[0]),.doutb(w_n3770_0[1]),.din(n3770));
	jspl jspl_w_n3773_0(.douta(w_n3773_0[0]),.doutb(w_n3773_0[1]),.din(n3773));
	jspl jspl_w_n3780_0(.douta(w_n3780_0[0]),.doutb(w_n3780_0[1]),.din(n3780));
	jspl jspl_w_n3787_0(.douta(w_n3787_0[0]),.doutb(w_n3787_0[1]),.din(n3787));
	jspl jspl_w_n3789_0(.douta(w_n3789_0[0]),.doutb(w_n3789_0[1]),.din(n3789));
	jspl jspl_w_n3790_0(.douta(w_n3790_0[0]),.doutb(w_n3790_0[1]),.din(n3790));
	jspl jspl_w_n3798_0(.douta(w_n3798_0[0]),.doutb(w_n3798_0[1]),.din(n3798));
	jspl jspl_w_n3799_0(.douta(w_n3799_0[0]),.doutb(w_n3799_0[1]),.din(n3799));
	jspl jspl_w_n3801_0(.douta(w_n3801_0[0]),.doutb(w_n3801_0[1]),.din(n3801));
	jspl jspl_w_n3809_0(.douta(w_n3809_0[0]),.doutb(w_n3809_0[1]),.din(n3809));
	jspl jspl_w_n3810_0(.douta(w_n3810_0[0]),.doutb(w_n3810_0[1]),.din(n3810));
	jspl jspl_w_n3811_0(.douta(w_n3811_0[0]),.doutb(w_n3811_0[1]),.din(n3811));
	jspl jspl_w_n3819_0(.douta(w_n3819_0[0]),.doutb(w_n3819_0[1]),.din(n3819));
	jspl jspl_w_n3820_0(.douta(w_n3820_0[0]),.doutb(w_n3820_0[1]),.din(n3820));
	jspl jspl_w_n3821_0(.douta(w_n3821_0[0]),.doutb(w_n3821_0[1]),.din(n3821));
	jspl jspl_w_n3824_0(.douta(w_n3824_0[0]),.doutb(w_n3824_0[1]),.din(n3824));
	jspl3 jspl3_w_n3825_0(.douta(w_n3825_0[0]),.doutb(w_n3825_0[1]),.doutc(w_n3825_0[2]),.din(n3825));
	jspl jspl_w_n3826_0(.douta(w_n3826_0[0]),.doutb(w_n3826_0[1]),.din(n3826));
	jspl3 jspl3_w_n3833_0(.douta(w_n3833_0[0]),.doutb(w_n3833_0[1]),.doutc(w_n3833_0[2]),.din(n3833));
	jspl jspl_w_n3836_0(.douta(w_n3836_0[0]),.doutb(w_n3836_0[1]),.din(n3836));
	jspl3 jspl3_w_n3837_0(.douta(w_n3837_0[0]),.doutb(w_n3837_0[1]),.doutc(w_n3837_0[2]),.din(n3837));
	jspl3 jspl3_w_n3837_1(.douta(w_n3837_1[0]),.doutb(w_n3837_1[1]),.doutc(w_n3837_1[2]),.din(w_n3837_0[0]));
	jspl3 jspl3_w_n3837_2(.douta(w_n3837_2[0]),.doutb(w_n3837_2[1]),.doutc(w_n3837_2[2]),.din(w_n3837_0[1]));
	jspl3 jspl3_w_n3837_3(.douta(w_n3837_3[0]),.doutb(w_n3837_3[1]),.doutc(w_n3837_3[2]),.din(w_n3837_0[2]));
	jspl3 jspl3_w_n3837_4(.douta(w_n3837_4[0]),.doutb(w_n3837_4[1]),.doutc(w_n3837_4[2]),.din(w_n3837_1[0]));
	jspl3 jspl3_w_n3837_5(.douta(w_n3837_5[0]),.doutb(w_n3837_5[1]),.doutc(w_n3837_5[2]),.din(w_n3837_1[1]));
	jspl3 jspl3_w_n3837_6(.douta(w_n3837_6[0]),.doutb(w_n3837_6[1]),.doutc(w_n3837_6[2]),.din(w_n3837_1[2]));
	jspl3 jspl3_w_n3837_7(.douta(w_n3837_7[0]),.doutb(w_n3837_7[1]),.doutc(w_n3837_7[2]),.din(w_n3837_2[0]));
	jspl jspl_w_n3837_8(.douta(w_n3837_8[0]),.doutb(w_n3837_8[1]),.din(w_n3837_2[1]));
	jspl3 jspl3_w_n3838_0(.douta(w_n3838_0[0]),.doutb(w_n3838_0[1]),.doutc(w_n3838_0[2]),.din(n3838));
	jspl jspl_w_n3838_1(.douta(w_n3838_1[0]),.doutb(w_n3838_1[1]),.din(w_n3838_0[0]));
	jspl jspl_w_n3839_0(.douta(w_n3839_0[0]),.doutb(w_n3839_0[1]),.din(n3839));
	jspl jspl_w_n3840_0(.douta(w_n3840_0[0]),.doutb(w_n3840_0[1]),.din(n3840));
	jspl3 jspl3_w_n3841_0(.douta(w_n3841_0[0]),.doutb(w_n3841_0[1]),.doutc(w_n3841_0[2]),.din(n3841));
	jspl3 jspl3_w_n3842_0(.douta(w_n3842_0[0]),.doutb(w_n3842_0[1]),.doutc(w_n3842_0[2]),.din(n3842));
	jspl3 jspl3_w_n3842_1(.douta(w_n3842_1[0]),.doutb(w_n3842_1[1]),.doutc(w_n3842_1[2]),.din(w_n3842_0[0]));
	jspl jspl_w_n3850_0(.douta(w_n3850_0[0]),.doutb(w_n3850_0[1]),.din(n3850));
	jspl3 jspl3_w_n3851_0(.douta(w_n3851_0[0]),.doutb(w_n3851_0[1]),.doutc(w_n3851_0[2]),.din(n3851));
	jspl3 jspl3_w_n3852_0(.douta(w_n3852_0[0]),.doutb(w_n3852_0[1]),.doutc(w_n3852_0[2]),.din(n3852));
	jspl jspl_w_n3853_0(.douta(w_n3853_0[0]),.doutb(w_n3853_0[1]),.din(n3853));
	jspl jspl_w_n3854_0(.douta(w_n3854_0[0]),.doutb(w_n3854_0[1]),.din(n3854));
	jspl jspl_w_n3868_0(.douta(w_n3868_0[0]),.doutb(w_n3868_0[1]),.din(n3868));
	jspl jspl_w_n3871_0(.douta(w_n3871_0[0]),.doutb(w_n3871_0[1]),.din(n3871));
	jspl jspl_w_n3875_0(.douta(w_n3875_0[0]),.doutb(w_n3875_0[1]),.din(n3875));
	jspl jspl_w_n3881_0(.douta(w_n3881_0[0]),.doutb(w_n3881_0[1]),.din(n3881));
	jspl jspl_w_n3887_0(.douta(w_n3887_0[0]),.doutb(w_n3887_0[1]),.din(n3887));
	jspl3 jspl3_w_n3892_0(.douta(w_n3892_0[0]),.doutb(w_n3892_0[1]),.doutc(w_n3892_0[2]),.din(n3892));
	jspl jspl_w_n3895_0(.douta(w_n3895_0[0]),.doutb(w_n3895_0[1]),.din(n3895));
	jspl jspl_w_n3910_0(.douta(w_n3910_0[0]),.doutb(w_n3910_0[1]),.din(n3910));
	jspl jspl_w_n3959_0(.douta(w_n3959_0[0]),.doutb(w_n3959_0[1]),.din(n3959));
	jspl jspl_w_n3961_0(.douta(w_n3961_0[0]),.doutb(w_n3961_0[1]),.din(n3961));
	jspl jspl_w_n3963_0(.douta(w_n3963_0[0]),.doutb(w_n3963_0[1]),.din(n3963));
	jspl jspl_w_n3968_0(.douta(w_n3968_0[0]),.doutb(w_n3968_0[1]),.din(n3968));
	jspl jspl_w_n3969_0(.douta(w_n3969_0[0]),.doutb(w_n3969_0[1]),.din(n3969));
	jspl jspl_w_n3971_0(.douta(w_n3971_0[0]),.doutb(w_n3971_0[1]),.din(n3971));
	jspl jspl_w_n3972_0(.douta(w_n3972_0[0]),.doutb(w_n3972_0[1]),.din(n3972));
	jspl jspl_w_n3982_0(.douta(w_n3982_0[0]),.doutb(w_n3982_0[1]),.din(n3982));
	jspl jspl_w_n3985_0(.douta(w_n3985_0[0]),.doutb(w_n3985_0[1]),.din(n3985));
	jspl jspl_w_n3989_0(.douta(w_n3989_0[0]),.doutb(w_n3989_0[1]),.din(n3989));
	jspl jspl_w_n3992_0(.douta(w_n3992_0[0]),.doutb(w_n3992_0[1]),.din(n3992));
	jspl jspl_w_n3998_0(.douta(w_n3998_0[0]),.doutb(w_n3998_0[1]),.din(n3998));
	jspl jspl_w_n4006_0(.douta(w_n4006_0[0]),.doutb(w_n4006_0[1]),.din(n4006));
	jspl jspl_w_n4008_0(.douta(w_n4008_0[0]),.doutb(w_n4008_0[1]),.din(n4008));
	jspl jspl_w_n4009_0(.douta(w_n4009_0[0]),.doutb(w_n4009_0[1]),.din(n4009));
	jspl jspl_w_n4017_0(.douta(w_n4017_0[0]),.doutb(w_n4017_0[1]),.din(n4017));
	jspl jspl_w_n4018_0(.douta(w_n4018_0[0]),.doutb(w_n4018_0[1]),.din(n4018));
	jspl jspl_w_n4020_0(.douta(w_n4020_0[0]),.doutb(w_n4020_0[1]),.din(n4020));
	jspl jspl_w_n4028_0(.douta(w_n4028_0[0]),.doutb(w_n4028_0[1]),.din(n4028));
	jspl jspl_w_n4029_0(.douta(w_n4029_0[0]),.doutb(w_n4029_0[1]),.din(n4029));
	jspl jspl_w_n4030_0(.douta(w_n4030_0[0]),.doutb(w_n4030_0[1]),.din(n4030));
	jspl jspl_w_n4038_0(.douta(w_n4038_0[0]),.doutb(w_n4038_0[1]),.din(n4038));
	jspl jspl_w_n4039_0(.douta(w_n4039_0[0]),.doutb(w_n4039_0[1]),.din(n4039));
	jspl jspl_w_n4040_0(.douta(w_n4040_0[0]),.doutb(w_n4040_0[1]),.din(n4040));
	jspl jspl_w_n4043_0(.douta(w_n4043_0[0]),.doutb(w_n4043_0[1]),.din(n4043));
	jspl jspl_w_n4051_0(.douta(w_n4051_0[0]),.doutb(w_n4051_0[1]),.din(n4051));
	jspl3 jspl3_w_n4059_0(.douta(w_n4059_0[0]),.doutb(w_n4059_0[1]),.doutc(w_n4059_0[2]),.din(n4059));
	jspl jspl_w_n4062_0(.douta(w_n4062_0[0]),.doutb(w_n4062_0[1]),.din(n4062));
	jspl3 jspl3_w_n4063_0(.douta(w_n4063_0[0]),.doutb(w_n4063_0[1]),.doutc(w_n4063_0[2]),.din(n4063));
	jspl3 jspl3_w_n4063_1(.douta(w_n4063_1[0]),.doutb(w_n4063_1[1]),.doutc(w_n4063_1[2]),.din(w_n4063_0[0]));
	jspl3 jspl3_w_n4063_2(.douta(w_n4063_2[0]),.doutb(w_n4063_2[1]),.doutc(w_n4063_2[2]),.din(w_n4063_0[1]));
	jspl3 jspl3_w_n4063_3(.douta(w_n4063_3[0]),.doutb(w_n4063_3[1]),.doutc(w_n4063_3[2]),.din(w_n4063_0[2]));
	jspl3 jspl3_w_n4063_4(.douta(w_n4063_4[0]),.doutb(w_n4063_4[1]),.doutc(w_n4063_4[2]),.din(w_n4063_1[0]));
	jspl3 jspl3_w_n4063_5(.douta(w_n4063_5[0]),.doutb(w_n4063_5[1]),.doutc(w_n4063_5[2]),.din(w_n4063_1[1]));
	jspl3 jspl3_w_n4063_6(.douta(w_n4063_6[0]),.doutb(w_n4063_6[1]),.doutc(w_n4063_6[2]),.din(w_n4063_1[2]));
	jspl3 jspl3_w_n4063_7(.douta(w_n4063_7[0]),.doutb(w_n4063_7[1]),.doutc(w_n4063_7[2]),.din(w_n4063_2[0]));
	jspl jspl_w_n4063_8(.douta(w_n4063_8[0]),.doutb(w_n4063_8[1]),.din(w_n4063_2[1]));
	jspl3 jspl3_w_n4064_0(.douta(w_n4064_0[0]),.doutb(w_n4064_0[1]),.doutc(w_n4064_0[2]),.din(n4064));
	jspl3 jspl3_w_n4065_0(.douta(w_n4065_0[0]),.doutb(w_n4065_0[1]),.doutc(w_n4065_0[2]),.din(n4065));
	jspl3 jspl3_w_n4066_0(.douta(w_n4066_0[0]),.doutb(w_n4066_0[1]),.doutc(w_n4066_0[2]),.din(n4066));
	jspl3 jspl3_w_n4066_1(.douta(w_n4066_1[0]),.doutb(w_n4066_1[1]),.doutc(w_n4066_1[2]),.din(w_n4066_0[0]));
	jspl jspl_w_n4074_0(.douta(w_n4074_0[0]),.doutb(w_n4074_0[1]),.din(n4074));
	jspl3 jspl3_w_n4075_0(.douta(w_n4075_0[0]),.doutb(w_n4075_0[1]),.doutc(w_n4075_0[2]),.din(n4075));
	jspl jspl_w_n4075_1(.douta(w_n4075_1[0]),.doutb(w_n4075_1[1]),.din(w_n4075_0[0]));
	jspl jspl_w_n4076_0(.douta(w_n4076_0[0]),.doutb(w_n4076_0[1]),.din(n4076));
	jspl3 jspl3_w_n4088_0(.douta(w_n4088_0[0]),.doutb(w_n4088_0[1]),.doutc(w_n4088_0[2]),.din(n4088));
	jspl jspl_w_n4089_0(.douta(w_n4089_0[0]),.doutb(w_n4089_0[1]),.din(n4089));
	jspl jspl_w_n4090_0(.douta(w_n4090_0[0]),.doutb(w_n4090_0[1]),.din(n4090));
	jspl jspl_w_n4091_0(.douta(w_n4091_0[0]),.doutb(w_n4091_0[1]),.din(n4091));
	jspl3 jspl3_w_n4093_0(.douta(w_n4093_0[0]),.doutb(w_n4093_0[1]),.doutc(w_n4093_0[2]),.din(n4093));
	jspl3 jspl3_w_n4093_1(.douta(w_n4093_1[0]),.doutb(w_n4093_1[1]),.doutc(w_n4093_1[2]),.din(w_n4093_0[0]));
	jspl3 jspl3_w_n4093_2(.douta(w_dff_A_fbO785X92_0),.doutb(w_dff_A_9NWZDZCv5_1),.doutc(w_n4093_2[2]),.din(w_n4093_0[1]));
	jspl3 jspl3_w_n4093_3(.douta(w_dff_A_SAnq582t7_0),.doutb(w_n4093_3[1]),.doutc(w_dff_A_IxICBTvT9_2),.din(w_n4093_0[2]));
	jspl3 jspl3_w_n4093_4(.douta(w_n4093_4[0]),.doutb(w_n4093_4[1]),.doutc(w_n4093_4[2]),.din(w_n4093_1[0]));
	jspl3 jspl3_w_n4093_5(.douta(w_dff_A_Iu0AqP8D9_0),.doutb(w_dff_A_suv5RVkp5_1),.doutc(w_n4093_5[2]),.din(w_n4093_1[1]));
	jspl3 jspl3_w_n4093_6(.douta(w_dff_A_8BQJrza76_0),.doutb(w_dff_A_imlgG5NP4_1),.doutc(w_n4093_6[2]),.din(w_n4093_1[2]));
	jspl3 jspl3_w_n4093_7(.douta(w_dff_A_xH2PJntQ0_0),.doutb(w_dff_A_55rtkZ763_1),.doutc(w_n4093_7[2]),.din(w_n4093_2[0]));
	jspl3 jspl3_w_n4093_8(.douta(w_dff_A_cUDtSJyJ3_0),.doutb(w_dff_A_BPbGrQYz5_1),.doutc(w_n4093_8[2]),.din(w_n4093_2[1]));
	jspl3 jspl3_w_n4093_9(.douta(w_dff_A_AZO8FXmC7_0),.doutb(w_dff_A_wpA3GKq05_1),.doutc(w_n4093_9[2]),.din(w_n4093_2[2]));
	jspl3 jspl3_w_n4093_10(.douta(w_dff_A_k4Whxaqa7_0),.doutb(w_dff_A_8u2TGooJ9_1),.doutc(w_n4093_10[2]),.din(w_n4093_3[0]));
	jspl jspl_w_n4093_11(.douta(w_dff_A_9OrtdDC35_0),.doutb(w_n4093_11[1]),.din(w_n4093_3[1]));
	jspl jspl_w_n4094_0(.douta(w_dff_A_nhphmE1W6_0),.doutb(w_n4094_0[1]),.din(n4094));
	jspl jspl_w_n4096_0(.douta(w_n4096_0[0]),.doutb(w_n4096_0[1]),.din(n4096));
	jspl jspl_w_n4097_0(.douta(w_n4097_0[0]),.doutb(w_n4097_0[1]),.din(n4097));
	jspl jspl_w_n4100_0(.douta(w_n4100_0[0]),.doutb(w_n4100_0[1]),.din(n4100));
	jspl jspl_w_n4101_0(.douta(w_n4101_0[0]),.doutb(w_n4101_0[1]),.din(n4101));
	jspl jspl_w_n4108_0(.douta(w_n4108_0[0]),.doutb(w_n4108_0[1]),.din(n4108));
	jspl jspl_w_n4112_0(.douta(w_n4112_0[0]),.doutb(w_n4112_0[1]),.din(n4112));
	jspl jspl_w_n4115_0(.douta(w_n4115_0[0]),.doutb(w_n4115_0[1]),.din(n4115));
	jspl jspl_w_n4120_0(.douta(w_n4120_0[0]),.doutb(w_n4120_0[1]),.din(n4120));
	jspl jspl_w_n4128_0(.douta(w_n4128_0[0]),.doutb(w_n4128_0[1]),.din(n4128));
	jspl jspl_w_n4130_0(.douta(w_n4130_0[0]),.doutb(w_n4130_0[1]),.din(n4130));
	jspl jspl_w_n4132_0(.douta(w_n4132_0[0]),.doutb(w_n4132_0[1]),.din(n4132));
	jspl jspl_w_n4140_0(.douta(w_n4140_0[0]),.doutb(w_n4140_0[1]),.din(n4140));
	jspl jspl_w_n4141_0(.douta(w_n4141_0[0]),.doutb(w_n4141_0[1]),.din(n4141));
	jspl jspl_w_n4143_0(.douta(w_n4143_0[0]),.doutb(w_n4143_0[1]),.din(n4143));
	jspl jspl_w_n4151_0(.douta(w_n4151_0[0]),.doutb(w_n4151_0[1]),.din(n4151));
	jspl jspl_w_n4152_0(.douta(w_n4152_0[0]),.doutb(w_n4152_0[1]),.din(n4152));
	jspl jspl_w_n4153_0(.douta(w_n4153_0[0]),.doutb(w_n4153_0[1]),.din(n4153));
	jspl jspl_w_n4161_0(.douta(w_n4161_0[0]),.doutb(w_n4161_0[1]),.din(n4161));
	jspl jspl_w_n4162_0(.douta(w_n4162_0[0]),.doutb(w_n4162_0[1]),.din(n4162));
	jspl jspl_w_n4163_0(.douta(w_n4163_0[0]),.doutb(w_n4163_0[1]),.din(n4163));
	jspl jspl_w_n4194_0(.douta(w_n4194_0[0]),.doutb(w_n4194_0[1]),.din(n4194));
	jspl jspl_w_n4203_0(.douta(w_n4203_0[0]),.doutb(w_n4203_0[1]),.din(n4203));
	jspl3 jspl3_w_n4213_0(.douta(w_n4213_0[0]),.doutb(w_n4213_0[1]),.doutc(w_n4213_0[2]),.din(n4213));
	jspl3 jspl3_w_n4213_1(.douta(w_n4213_1[0]),.doutb(w_n4213_1[1]),.doutc(w_n4213_1[2]),.din(w_n4213_0[0]));
	jspl3 jspl3_w_n4213_2(.douta(w_n4213_2[0]),.doutb(w_n4213_2[1]),.doutc(w_n4213_2[2]),.din(w_n4213_0[1]));
	jspl3 jspl3_w_n4213_3(.douta(w_n4213_3[0]),.doutb(w_n4213_3[1]),.doutc(w_n4213_3[2]),.din(w_n4213_0[2]));
	jspl3 jspl3_w_n4213_4(.douta(w_n4213_4[0]),.doutb(w_n4213_4[1]),.doutc(w_n4213_4[2]),.din(w_n4213_1[0]));
	jspl3 jspl3_w_n4213_5(.douta(w_n4213_5[0]),.doutb(w_n4213_5[1]),.doutc(w_n4213_5[2]),.din(w_n4213_1[1]));
	jspl3 jspl3_w_n4213_6(.douta(w_n4213_6[0]),.doutb(w_n4213_6[1]),.doutc(w_n4213_6[2]),.din(w_n4213_1[2]));
	jspl3 jspl3_w_n4214_0(.douta(w_n4214_0[0]),.doutb(w_n4214_0[1]),.doutc(w_n4214_0[2]),.din(n4214));
	jspl3 jspl3_w_n4215_0(.douta(w_n4215_0[0]),.doutb(w_n4215_0[1]),.doutc(w_n4215_0[2]),.din(n4215));
	jspl3 jspl3_w_n4215_1(.douta(w_n4215_1[0]),.doutb(w_n4215_1[1]),.doutc(w_n4215_1[2]),.din(w_n4215_0[0]));
	jspl jspl_w_n4225_0(.douta(w_n4225_0[0]),.doutb(w_n4225_0[1]),.din(n4225));
	jspl3 jspl3_w_n4226_0(.douta(w_n4226_0[0]),.doutb(w_n4226_0[1]),.doutc(w_n4226_0[2]),.din(n4226));
	jspl jspl_w_n4227_0(.douta(w_n4227_0[0]),.doutb(w_n4227_0[1]),.din(n4227));
	jspl3 jspl3_w_n4237_0(.douta(w_n4237_0[0]),.doutb(w_n4237_0[1]),.doutc(w_n4237_0[2]),.din(n4237));
	jspl3 jspl3_w_n4242_0(.douta(w_n4242_0[0]),.doutb(w_n4242_0[1]),.doutc(w_n4242_0[2]),.din(n4242));
	jspl jspl_w_n4243_0(.douta(w_n4243_0[0]),.doutb(w_n4243_0[1]),.din(n4243));
	jspl3 jspl3_w_n4244_0(.douta(w_n4244_0[0]),.doutb(w_n4244_0[1]),.doutc(w_n4244_0[2]),.din(n4244));
	jspl jspl_w_n4245_0(.douta(w_n4245_0[0]),.doutb(w_n4245_0[1]),.din(n4245));
	jspl jspl_w_n4250_0(.douta(w_n4250_0[0]),.doutb(w_n4250_0[1]),.din(n4250));
	jspl jspl_w_n4251_0(.douta(w_n4251_0[0]),.doutb(w_n4251_0[1]),.din(n4251));
	jspl jspl_w_n4254_0(.douta(w_n4254_0[0]),.doutb(w_n4254_0[1]),.din(n4254));
	jspl jspl_w_n4266_0(.douta(w_n4266_0[0]),.doutb(w_n4266_0[1]),.din(n4266));
	jspl jspl_w_n4270_0(.douta(w_n4270_0[0]),.doutb(w_n4270_0[1]),.din(n4270));
	jspl jspl_w_n4271_0(.douta(w_n4271_0[0]),.doutb(w_n4271_0[1]),.din(n4271));
	jspl jspl_w_n4274_0(.douta(w_n4274_0[0]),.doutb(w_n4274_0[1]),.din(n4274));
	jspl jspl_w_n4276_0(.douta(w_n4276_0[0]),.doutb(w_n4276_0[1]),.din(n4276));
	jspl jspl_w_n4278_0(.douta(w_n4278_0[0]),.doutb(w_n4278_0[1]),.din(n4278));
	jspl jspl_w_n4281_0(.douta(w_n4281_0[0]),.doutb(w_n4281_0[1]),.din(n4281));
	jspl jspl_w_n4285_0(.douta(w_n4285_0[0]),.doutb(w_n4285_0[1]),.din(n4285));
	jspl jspl_w_n4290_0(.douta(w_n4290_0[0]),.doutb(w_n4290_0[1]),.din(n4290));
	jspl jspl_w_n4295_0(.douta(w_n4295_0[0]),.doutb(w_n4295_0[1]),.din(n4295));
	jspl jspl_w_n4303_0(.douta(w_n4303_0[0]),.doutb(w_n4303_0[1]),.din(n4303));
	jspl jspl_w_n4305_0(.douta(w_n4305_0[0]),.doutb(w_n4305_0[1]),.din(n4305));
	jspl jspl_w_n4307_0(.douta(w_n4307_0[0]),.doutb(w_n4307_0[1]),.din(n4307));
	jspl jspl_w_n4315_0(.douta(w_n4315_0[0]),.doutb(w_n4315_0[1]),.din(n4315));
	jspl jspl_w_n4316_0(.douta(w_n4316_0[0]),.doutb(w_n4316_0[1]),.din(n4316));
	jspl jspl_w_n4317_0(.douta(w_n4317_0[0]),.doutb(w_n4317_0[1]),.din(n4317));
	jspl jspl_w_n4325_0(.douta(w_n4325_0[0]),.doutb(w_n4325_0[1]),.din(n4325));
	jspl jspl_w_n4326_0(.douta(w_n4326_0[0]),.doutb(w_n4326_0[1]),.din(n4326));
	jspl jspl_w_n4327_0(.douta(w_n4327_0[0]),.doutb(w_n4327_0[1]),.din(n4327));
	jspl jspl_w_n4335_0(.douta(w_n4335_0[0]),.doutb(w_n4335_0[1]),.din(n4335));
	jspl jspl_w_n4336_0(.douta(w_n4336_0[0]),.doutb(w_n4336_0[1]),.din(n4336));
	jspl jspl_w_n4337_0(.douta(w_n4337_0[0]),.doutb(w_n4337_0[1]),.din(n4337));
	jspl3 jspl3_w_n4338_0(.douta(w_n4338_0[0]),.doutb(w_n4338_0[1]),.doutc(w_n4338_0[2]),.din(n4338));
	jspl3 jspl3_w_n4338_1(.douta(w_n4338_1[0]),.doutb(w_n4338_1[1]),.doutc(w_n4338_1[2]),.din(w_n4338_0[0]));
	jspl3 jspl3_w_n4343_0(.douta(w_n4343_0[0]),.doutb(w_n4343_0[1]),.doutc(w_n4343_0[2]),.din(n4343));
	jspl3 jspl3_w_n4343_1(.douta(w_n4343_1[0]),.doutb(w_n4343_1[1]),.doutc(w_n4343_1[2]),.din(w_n4343_0[0]));
	jspl jspl_w_n4343_2(.douta(w_n4343_2[0]),.doutb(w_n4343_2[1]),.din(w_n4343_0[1]));
	jspl jspl_w_n4344_0(.douta(w_n4344_0[0]),.doutb(w_n4344_0[1]),.din(n4344));
	jspl3 jspl3_w_n4349_0(.douta(w_n4349_0[0]),.doutb(w_n4349_0[1]),.doutc(w_n4349_0[2]),.din(n4349));
	jspl3 jspl3_w_n4349_1(.douta(w_n4349_1[0]),.doutb(w_n4349_1[1]),.doutc(w_n4349_1[2]),.din(w_n4349_0[0]));
	jspl jspl_w_n4355_0(.douta(w_n4355_0[0]),.doutb(w_n4355_0[1]),.din(n4355));
	jspl jspl_w_n4356_0(.douta(w_n4356_0[0]),.doutb(w_n4356_0[1]),.din(n4356));
	jspl3 jspl3_w_n4357_0(.douta(w_n4357_0[0]),.doutb(w_n4357_0[1]),.doutc(w_n4357_0[2]),.din(n4357));
	jspl jspl_w_n4358_0(.douta(w_n4358_0[0]),.doutb(w_n4358_0[1]),.din(n4358));
	jspl jspl_w_n4359_0(.douta(w_n4359_0[0]),.doutb(w_n4359_0[1]),.din(n4359));
	jspl jspl_w_n4360_0(.douta(w_n4360_0[0]),.doutb(w_n4360_0[1]),.din(n4360));
	jspl jspl_w_n4361_0(.douta(w_dff_A_nhCEAzVC8_0),.doutb(w_n4361_0[1]),.din(n4361));
	jspl jspl_w_n4364_0(.douta(w_dff_A_y8pPL52h4_0),.doutb(w_n4364_0[1]),.din(n4364));
	jspl jspl_w_n4366_0(.douta(w_n4366_0[0]),.doutb(w_n4366_0[1]),.din(n4366));
	jspl jspl_w_n4367_0(.douta(w_n4367_0[0]),.doutb(w_n4367_0[1]),.din(n4367));
	jspl jspl_w_n4369_0(.douta(w_n4369_0[0]),.doutb(w_n4369_0[1]),.din(n4369));
	jspl jspl_w_n4381_0(.douta(w_n4381_0[0]),.doutb(w_n4381_0[1]),.din(n4381));
	jspl jspl_w_n4382_0(.douta(w_n4382_0[0]),.doutb(w_n4382_0[1]),.din(n4382));
	jspl jspl_w_n4385_0(.douta(w_n4385_0[0]),.doutb(w_n4385_0[1]),.din(n4385));
	jspl jspl_w_n4388_0(.douta(w_n4388_0[0]),.doutb(w_n4388_0[1]),.din(n4388));
	jspl jspl_w_n4391_0(.douta(w_n4391_0[0]),.doutb(w_n4391_0[1]),.din(n4391));
	jspl jspl_w_n4396_0(.douta(w_n4396_0[0]),.doutb(w_n4396_0[1]),.din(n4396));
	jspl jspl_w_n4401_0(.douta(w_n4401_0[0]),.doutb(w_n4401_0[1]),.din(n4401));
	jspl jspl_w_n4409_0(.douta(w_n4409_0[0]),.doutb(w_n4409_0[1]),.din(n4409));
	jspl jspl_w_n4411_0(.douta(w_n4411_0[0]),.doutb(w_n4411_0[1]),.din(n4411));
	jspl jspl_w_n4413_0(.douta(w_n4413_0[0]),.doutb(w_n4413_0[1]),.din(n4413));
	jspl jspl_w_n4421_0(.douta(w_n4421_0[0]),.doutb(w_n4421_0[1]),.din(n4421));
	jspl jspl_w_n4422_0(.douta(w_n4422_0[0]),.doutb(w_n4422_0[1]),.din(n4422));
	jspl jspl_w_n4424_0(.douta(w_n4424_0[0]),.doutb(w_n4424_0[1]),.din(n4424));
	jspl jspl_w_n4432_0(.douta(w_n4432_0[0]),.doutb(w_n4432_0[1]),.din(n4432));
	jspl jspl_w_n4433_0(.douta(w_n4433_0[0]),.doutb(w_n4433_0[1]),.din(n4433));
	jspl jspl_w_n4434_0(.douta(w_n4434_0[0]),.doutb(w_n4434_0[1]),.din(n4434));
	jspl jspl_w_n4442_0(.douta(w_n4442_0[0]),.doutb(w_n4442_0[1]),.din(n4442));
	jspl jspl_w_n4443_0(.douta(w_n4443_0[0]),.doutb(w_n4443_0[1]),.din(n4443));
	jspl jspl_w_n4448_0(.douta(w_n4448_0[0]),.doutb(w_n4448_0[1]),.din(n4448));
	jspl jspl_w_n4449_0(.douta(w_n4449_0[0]),.doutb(w_n4449_0[1]),.din(n4449));
	jspl jspl_w_n4450_0(.douta(w_n4450_0[0]),.doutb(w_n4450_0[1]),.din(n4450));
	jspl3 jspl3_w_n4451_0(.douta(w_n4451_0[0]),.doutb(w_n4451_0[1]),.doutc(w_n4451_0[2]),.din(n4451));
	jspl jspl_w_n4452_0(.douta(w_n4452_0[0]),.doutb(w_n4452_0[1]),.din(n4452));
	jspl jspl_w_n4453_0(.douta(w_n4453_0[0]),.doutb(w_n4453_0[1]),.din(n4453));
	jspl jspl_w_n4454_0(.douta(w_n4454_0[0]),.doutb(w_n4454_0[1]),.din(n4454));
	jspl jspl_w_n4456_0(.douta(w_n4456_0[0]),.doutb(w_n4456_0[1]),.din(n4456));
	jspl jspl_w_n4457_0(.douta(w_n4457_0[0]),.doutb(w_n4457_0[1]),.din(n4457));
	jspl jspl_w_n4459_0(.douta(w_n4459_0[0]),.doutb(w_n4459_0[1]),.din(n4459));
	jspl jspl_w_n4469_0(.douta(w_n4469_0[0]),.doutb(w_n4469_0[1]),.din(n4469));
	jspl jspl_w_n4470_0(.douta(w_n4470_0[0]),.doutb(w_n4470_0[1]),.din(n4470));
	jspl jspl_w_n4473_0(.douta(w_n4473_0[0]),.doutb(w_n4473_0[1]),.din(n4473));
	jspl jspl_w_n4480_0(.douta(w_n4480_0[0]),.doutb(w_n4480_0[1]),.din(n4480));
	jspl jspl_w_n4484_0(.douta(w_n4484_0[0]),.doutb(w_n4484_0[1]),.din(n4484));
	jspl jspl_w_n4489_0(.douta(w_n4489_0[0]),.doutb(w_n4489_0[1]),.din(n4489));
	jspl jspl_w_n4495_0(.douta(w_n4495_0[0]),.doutb(w_n4495_0[1]),.din(n4495));
	jspl jspl_w_n4496_0(.douta(w_n4496_0[0]),.doutb(w_n4496_0[1]),.din(n4496));
	jspl jspl_w_n4497_0(.douta(w_n4497_0[0]),.doutb(w_n4497_0[1]),.din(n4497));
	jspl jspl_w_n4505_0(.douta(w_n4505_0[0]),.doutb(w_n4505_0[1]),.din(n4505));
	jspl jspl_w_n4506_0(.douta(w_n4506_0[0]),.doutb(w_n4506_0[1]),.din(n4506));
	jspl jspl_w_n4508_0(.douta(w_n4508_0[0]),.doutb(w_n4508_0[1]),.din(n4508));
	jspl jspl_w_n4516_0(.douta(w_n4516_0[0]),.doutb(w_n4516_0[1]),.din(n4516));
	jspl jspl_w_n4517_0(.douta(w_n4517_0[0]),.doutb(w_n4517_0[1]),.din(n4517));
	jspl jspl_w_n4518_0(.douta(w_n4518_0[0]),.doutb(w_n4518_0[1]),.din(n4518));
	jspl jspl_w_n4526_0(.douta(w_n4526_0[0]),.doutb(w_n4526_0[1]),.din(n4526));
	jspl jspl_w_n4527_0(.douta(w_n4527_0[0]),.doutb(w_n4527_0[1]),.din(n4527));
	jspl jspl_w_n4528_0(.douta(w_n4528_0[0]),.doutb(w_n4528_0[1]),.din(n4528));
	jspl jspl_w_n4536_0(.douta(w_n4536_0[0]),.doutb(w_n4536_0[1]),.din(n4536));
	jspl jspl_w_n4537_0(.douta(w_n4537_0[0]),.doutb(w_n4537_0[1]),.din(n4537));
	jspl jspl_w_n4538_0(.douta(w_n4538_0[0]),.doutb(w_n4538_0[1]),.din(n4538));
	jspl3 jspl3_w_n4539_0(.douta(w_n4539_0[0]),.doutb(w_n4539_0[1]),.doutc(w_n4539_0[2]),.din(n4539));
	jspl jspl_w_n4540_0(.douta(w_n4540_0[0]),.doutb(w_n4540_0[1]),.din(n4540));
	jspl jspl_w_n4541_0(.douta(w_n4541_0[0]),.doutb(w_n4541_0[1]),.din(n4541));
	jspl jspl_w_n4542_0(.douta(w_n4542_0[0]),.doutb(w_n4542_0[1]),.din(n4542));
	jspl jspl_w_n4543_0(.douta(w_dff_A_rxmmLz2D9_0),.doutb(w_n4543_0[1]),.din(n4543));
	jspl jspl_w_n4546_0(.douta(w_n4546_0[0]),.doutb(w_n4546_0[1]),.din(n4546));
	jspl jspl_w_n4547_0(.douta(w_n4547_0[0]),.doutb(w_n4547_0[1]),.din(n4547));
	jspl jspl_w_n4549_0(.douta(w_n4549_0[0]),.doutb(w_n4549_0[1]),.din(n4549));
	jspl jspl_w_n4556_0(.douta(w_n4556_0[0]),.doutb(w_n4556_0[1]),.din(n4556));
	jspl3 jspl3_w_n4558_0(.douta(w_n4558_0[0]),.doutb(w_n4558_0[1]),.doutc(w_n4558_0[2]),.din(n4558));
	jspl jspl_w_n4563_0(.douta(w_n4563_0[0]),.doutb(w_n4563_0[1]),.din(n4563));
	jspl jspl_w_n4564_0(.douta(w_n4564_0[0]),.doutb(w_n4564_0[1]),.din(n4564));
	jspl jspl_w_n4567_0(.douta(w_n4567_0[0]),.doutb(w_n4567_0[1]),.din(n4567));
	jspl jspl_w_n4572_0(.douta(w_n4572_0[0]),.doutb(w_n4572_0[1]),.din(n4572));
	jspl jspl_w_n4575_0(.douta(w_n4575_0[0]),.doutb(w_n4575_0[1]),.din(n4575));
	jspl jspl_w_n4580_0(.douta(w_n4580_0[0]),.doutb(w_n4580_0[1]),.din(n4580));
	jspl jspl_w_n4583_0(.douta(w_n4583_0[0]),.doutb(w_n4583_0[1]),.din(n4583));
	jspl jspl_w_n4584_0(.douta(w_n4584_0[0]),.doutb(w_n4584_0[1]),.din(n4584));
	jspl jspl_w_n4585_0(.douta(w_n4585_0[0]),.doutb(w_n4585_0[1]),.din(n4585));
	jspl jspl_w_n4586_0(.douta(w_n4586_0[0]),.doutb(w_n4586_0[1]),.din(n4586));
	jspl jspl_w_n4594_0(.douta(w_n4594_0[0]),.doutb(w_n4594_0[1]),.din(n4594));
	jspl jspl_w_n4595_0(.douta(w_n4595_0[0]),.doutb(w_n4595_0[1]),.din(n4595));
	jspl jspl_w_n4603_0(.douta(w_n4603_0[0]),.doutb(w_n4603_0[1]),.din(n4603));
	jspl jspl_w_n4604_0(.douta(w_n4604_0[0]),.doutb(w_n4604_0[1]),.din(n4604));
	jspl jspl_w_n4606_0(.douta(w_n4606_0[0]),.doutb(w_n4606_0[1]),.din(n4606));
	jspl jspl_w_n4614_0(.douta(w_n4614_0[0]),.doutb(w_n4614_0[1]),.din(n4614));
	jspl jspl_w_n4615_0(.douta(w_n4615_0[0]),.doutb(w_n4615_0[1]),.din(n4615));
	jspl jspl_w_n4616_0(.douta(w_n4616_0[0]),.doutb(w_n4616_0[1]),.din(n4616));
	jspl jspl_w_n4622_0(.douta(w_n4622_0[0]),.doutb(w_n4622_0[1]),.din(n4622));
	jspl jspl_w_n4623_0(.douta(w_n4623_0[0]),.doutb(w_n4623_0[1]),.din(n4623));
	jspl jspl_w_n4624_0(.douta(w_n4624_0[0]),.doutb(w_n4624_0[1]),.din(n4624));
	jspl3 jspl3_w_n4625_0(.douta(w_n4625_0[0]),.doutb(w_n4625_0[1]),.doutc(w_n4625_0[2]),.din(n4625));
	jspl jspl_w_n4626_0(.douta(w_n4626_0[0]),.doutb(w_n4626_0[1]),.din(n4626));
	jspl jspl_w_n4627_0(.douta(w_n4627_0[0]),.doutb(w_n4627_0[1]),.din(n4627));
	jspl jspl_w_n4628_0(.douta(w_n4628_0[0]),.doutb(w_n4628_0[1]),.din(n4628));
	jspl jspl_w_n4629_0(.douta(w_dff_A_kXRcecfy2_0),.doutb(w_n4629_0[1]),.din(n4629));
	jspl jspl_w_n4632_0(.douta(w_n4632_0[0]),.doutb(w_n4632_0[1]),.din(n4632));
	jspl jspl_w_n4633_0(.douta(w_n4633_0[0]),.doutb(w_n4633_0[1]),.din(n4633));
	jspl jspl_w_n4635_0(.douta(w_n4635_0[0]),.doutb(w_n4635_0[1]),.din(n4635));
	jspl jspl_w_n4643_0(.douta(w_n4643_0[0]),.doutb(w_n4643_0[1]),.din(n4643));
	jspl jspl_w_n4652_0(.douta(w_n4652_0[0]),.doutb(w_n4652_0[1]),.din(n4652));
	jspl jspl_w_n4653_0(.douta(w_n4653_0[0]),.doutb(w_n4653_0[1]),.din(n4653));
	jspl jspl_w_n4656_0(.douta(w_n4656_0[0]),.doutb(w_n4656_0[1]),.din(n4656));
	jspl jspl_w_n4659_0(.douta(w_n4659_0[0]),.doutb(w_n4659_0[1]),.din(n4659));
	jspl jspl_w_n4663_0(.douta(w_n4663_0[0]),.doutb(w_n4663_0[1]),.din(n4663));
	jspl jspl_w_n4667_0(.douta(w_n4667_0[0]),.doutb(w_n4667_0[1]),.din(n4667));
	jspl jspl_w_n4668_0(.douta(w_n4668_0[0]),.doutb(w_n4668_0[1]),.din(n4668));
	jspl jspl_w_n4671_0(.douta(w_n4671_0[0]),.doutb(w_n4671_0[1]),.din(n4671));
	jspl jspl_w_n4674_0(.douta(w_n4674_0[0]),.doutb(w_n4674_0[1]),.din(n4674));
	jspl jspl_w_n4675_0(.douta(w_n4675_0[0]),.doutb(w_n4675_0[1]),.din(n4675));
	jspl jspl_w_n4676_0(.douta(w_n4676_0[0]),.doutb(w_n4676_0[1]),.din(n4676));
	jspl jspl_w_n4677_0(.douta(w_n4677_0[0]),.doutb(w_n4677_0[1]),.din(n4677));
	jspl jspl_w_n4685_0(.douta(w_n4685_0[0]),.doutb(w_n4685_0[1]),.din(n4685));
	jspl jspl_w_n4686_0(.douta(w_n4686_0[0]),.doutb(w_n4686_0[1]),.din(n4686));
	jspl jspl_w_n4694_0(.douta(w_n4694_0[0]),.doutb(w_n4694_0[1]),.din(n4694));
	jspl jspl_w_n4695_0(.douta(w_n4695_0[0]),.doutb(w_n4695_0[1]),.din(n4695));
	jspl jspl_w_n4697_0(.douta(w_n4697_0[0]),.doutb(w_n4697_0[1]),.din(n4697));
	jspl jspl_w_n4705_0(.douta(w_n4705_0[0]),.doutb(w_n4705_0[1]),.din(n4705));
	jspl jspl_w_n4706_0(.douta(w_n4706_0[0]),.doutb(w_n4706_0[1]),.din(n4706));
	jspl jspl_w_n4707_0(.douta(w_n4707_0[0]),.doutb(w_n4707_0[1]),.din(n4707));
	jspl jspl_w_n4708_0(.douta(w_n4708_0[0]),.doutb(w_n4708_0[1]),.din(n4708));
	jspl3 jspl3_w_n4709_0(.douta(w_n4709_0[0]),.doutb(w_n4709_0[1]),.doutc(w_n4709_0[2]),.din(n4709));
	jspl jspl_w_n4710_0(.douta(w_n4710_0[0]),.doutb(w_n4710_0[1]),.din(n4710));
	jspl jspl_w_n4711_0(.douta(w_n4711_0[0]),.doutb(w_n4711_0[1]),.din(n4711));
	jspl jspl_w_n4712_0(.douta(w_n4712_0[0]),.doutb(w_n4712_0[1]),.din(n4712));
	jspl jspl_w_n4713_0(.douta(w_dff_A_CepdS1678_0),.doutb(w_n4713_0[1]),.din(n4713));
	jspl jspl_w_n4716_0(.douta(w_n4716_0[0]),.doutb(w_n4716_0[1]),.din(n4716));
	jspl jspl_w_n4717_0(.douta(w_n4717_0[0]),.doutb(w_n4717_0[1]),.din(n4717));
	jspl jspl_w_n4719_0(.douta(w_n4719_0[0]),.doutb(w_n4719_0[1]),.din(n4719));
	jspl3 jspl3_w_n4722_0(.douta(w_n4722_0[0]),.doutb(w_n4722_0[1]),.doutc(w_n4722_0[2]),.din(n4722));
	jspl jspl_w_n4727_0(.douta(w_n4727_0[0]),.doutb(w_n4727_0[1]),.din(n4727));
	jspl jspl_w_n4731_0(.douta(w_n4731_0[0]),.doutb(w_n4731_0[1]),.din(n4731));
	jspl jspl_w_n4739_0(.douta(w_n4739_0[0]),.doutb(w_n4739_0[1]),.din(n4739));
	jspl jspl_w_n4740_0(.douta(w_n4740_0[0]),.doutb(w_n4740_0[1]),.din(n4740));
	jspl jspl_w_n4743_0(.douta(w_n4743_0[0]),.doutb(w_n4743_0[1]),.din(n4743));
	jspl jspl_w_n4746_0(.douta(w_n4746_0[0]),.doutb(w_n4746_0[1]),.din(n4746));
	jspl jspl_w_n4747_0(.douta(w_n4747_0[0]),.doutb(w_n4747_0[1]),.din(n4747));
	jspl jspl_w_n4748_0(.douta(w_n4748_0[0]),.doutb(w_n4748_0[1]),.din(n4748));
	jspl jspl_w_n4749_0(.douta(w_n4749_0[0]),.doutb(w_n4749_0[1]),.din(n4749));
	jspl jspl_w_n4757_0(.douta(w_n4757_0[0]),.doutb(w_n4757_0[1]),.din(n4757));
	jspl jspl_w_n4758_0(.douta(w_n4758_0[0]),.doutb(w_n4758_0[1]),.din(n4758));
	jspl jspl_w_n4759_0(.douta(w_n4759_0[0]),.doutb(w_n4759_0[1]),.din(n4759));
	jspl jspl_w_n4767_0(.douta(w_n4767_0[0]),.doutb(w_n4767_0[1]),.din(n4767));
	jspl jspl_w_n4768_0(.douta(w_n4768_0[0]),.doutb(w_n4768_0[1]),.din(n4768));
	jspl jspl_w_n4769_0(.douta(w_n4769_0[0]),.doutb(w_n4769_0[1]),.din(n4769));
	jspl jspl_w_n4770_0(.douta(w_n4770_0[0]),.doutb(w_n4770_0[1]),.din(n4770));
	jspl3 jspl3_w_n4771_0(.douta(w_n4771_0[0]),.doutb(w_n4771_0[1]),.doutc(w_n4771_0[2]),.din(n4771));
	jspl jspl_w_n4773_0(.douta(w_n4773_0[0]),.doutb(w_n4773_0[1]),.din(n4773));
	jspl3 jspl3_w_n4782_0(.douta(w_n4782_0[0]),.doutb(w_n4782_0[1]),.doutc(w_n4782_0[2]),.din(n4782));
	jspl jspl_w_n4783_0(.douta(w_n4783_0[0]),.doutb(w_n4783_0[1]),.din(n4783));
	jspl jspl_w_n4784_0(.douta(w_n4784_0[0]),.doutb(w_n4784_0[1]),.din(n4784));
	jspl jspl_w_n4785_0(.douta(w_n4785_0[0]),.doutb(w_n4785_0[1]),.din(n4785));
	jspl jspl_w_n4786_0(.douta(w_dff_A_ws4tWc4i8_0),.doutb(w_n4786_0[1]),.din(n4786));
	jspl jspl_w_n4789_0(.douta(w_n4789_0[0]),.doutb(w_n4789_0[1]),.din(n4789));
	jspl jspl_w_n4790_0(.douta(w_n4790_0[0]),.doutb(w_n4790_0[1]),.din(n4790));
	jspl jspl_w_n4793_0(.douta(w_n4793_0[0]),.doutb(w_n4793_0[1]),.din(n4793));
	jspl jspl_w_n4811_0(.douta(w_n4811_0[0]),.doutb(w_n4811_0[1]),.din(n4811));
	jspl jspl_w_n4813_0(.douta(w_n4813_0[0]),.doutb(w_n4813_0[1]),.din(n4813));
	jspl jspl_w_n4814_0(.douta(w_n4814_0[0]),.doutb(w_n4814_0[1]),.din(n4814));
	jspl jspl_w_n4817_0(.douta(w_n4817_0[0]),.doutb(w_n4817_0[1]),.din(n4817));
	jspl jspl_w_n4822_0(.douta(w_n4822_0[0]),.doutb(w_n4822_0[1]),.din(n4822));
	jspl jspl_w_n4825_0(.douta(w_n4825_0[0]),.doutb(w_n4825_0[1]),.din(n4825));
	jspl jspl_w_n4828_0(.douta(w_n4828_0[0]),.doutb(w_n4828_0[1]),.din(n4828));
	jspl3 jspl3_w_n4829_0(.douta(w_n4829_0[0]),.doutb(w_n4829_0[1]),.doutc(w_n4829_0[2]),.din(n4829));
	jspl jspl_w_n4830_0(.douta(w_n4830_0[0]),.doutb(w_n4830_0[1]),.din(n4830));
	jspl jspl_w_n4833_0(.douta(w_n4833_0[0]),.doutb(w_n4833_0[1]),.din(n4833));
	jspl jspl_w_n4834_0(.douta(w_n4834_0[0]),.doutb(w_n4834_0[1]),.din(n4834));
	jspl jspl_w_n4842_0(.douta(w_n4842_0[0]),.doutb(w_n4842_0[1]),.din(n4842));
	jspl jspl_w_n4843_0(.douta(w_n4843_0[0]),.doutb(w_n4843_0[1]),.din(n4843));
	jspl jspl_w_n4845_0(.douta(w_n4845_0[0]),.doutb(w_n4845_0[1]),.din(n4845));
	jspl jspl_w_n4853_0(.douta(w_n4853_0[0]),.doutb(w_n4853_0[1]),.din(n4853));
	jspl jspl_w_n4854_0(.douta(w_n4854_0[0]),.doutb(w_n4854_0[1]),.din(n4854));
	jspl jspl_w_n4855_0(.douta(w_n4855_0[0]),.doutb(w_n4855_0[1]),.din(n4855));
	jspl jspl_w_n4861_0(.douta(w_n4861_0[0]),.doutb(w_n4861_0[1]),.din(n4861));
	jspl jspl_w_n4862_0(.douta(w_n4862_0[0]),.doutb(w_n4862_0[1]),.din(n4862));
	jspl jspl_w_n4863_0(.douta(w_n4863_0[0]),.doutb(w_n4863_0[1]),.din(n4863));
	jspl3 jspl3_w_n4864_0(.douta(w_n4864_0[0]),.doutb(w_n4864_0[1]),.doutc(w_n4864_0[2]),.din(n4864));
	jspl jspl_w_n4865_0(.douta(w_n4865_0[0]),.doutb(w_n4865_0[1]),.din(n4865));
	jspl jspl_w_n4866_0(.douta(w_n4866_0[0]),.doutb(w_n4866_0[1]),.din(n4866));
	jspl jspl_w_n4867_0(.douta(w_n4867_0[0]),.doutb(w_n4867_0[1]),.din(n4867));
	jspl jspl_w_n4868_0(.douta(w_dff_A_qqLHRbws4_0),.doutb(w_n4868_0[1]),.din(n4868));
	jspl jspl_w_n4871_0(.douta(w_n4871_0[0]),.doutb(w_n4871_0[1]),.din(n4871));
	jspl jspl_w_n4872_0(.douta(w_n4872_0[0]),.doutb(w_n4872_0[1]),.din(n4872));
	jspl jspl_w_n4874_0(.douta(w_n4874_0[0]),.doutb(w_n4874_0[1]),.din(n4874));
	jspl jspl_w_n4886_0(.douta(w_n4886_0[0]),.doutb(w_n4886_0[1]),.din(n4886));
	jspl jspl_w_n4887_0(.douta(w_n4887_0[0]),.doutb(w_n4887_0[1]),.din(n4887));
	jspl jspl_w_n4890_0(.douta(w_n4890_0[0]),.doutb(w_n4890_0[1]),.din(n4890));
	jspl jspl_w_n4893_0(.douta(w_n4893_0[0]),.doutb(w_n4893_0[1]),.din(n4893));
	jspl jspl_w_n4897_0(.douta(w_n4897_0[0]),.doutb(w_n4897_0[1]),.din(n4897));
	jspl jspl_w_n4901_0(.douta(w_n4901_0[0]),.doutb(w_n4901_0[1]),.din(n4901));
	jspl jspl_w_n4902_0(.douta(w_n4902_0[0]),.doutb(w_n4902_0[1]),.din(n4902));
	jspl jspl_w_n4905_0(.douta(w_n4905_0[0]),.doutb(w_n4905_0[1]),.din(n4905));
	jspl jspl_w_n4908_0(.douta(w_n4908_0[0]),.doutb(w_n4908_0[1]),.din(n4908));
	jspl3 jspl3_w_n4914_0(.douta(w_n4914_0[0]),.doutb(w_n4914_0[1]),.doutc(w_n4914_0[2]),.din(n4914));
	jspl jspl_w_n4915_0(.douta(w_n4915_0[0]),.doutb(w_n4915_0[1]),.din(n4915));
	jspl jspl_w_n4916_0(.douta(w_n4916_0[0]),.doutb(w_n4916_0[1]),.din(n4916));
	jspl jspl_w_n4918_0(.douta(w_n4918_0[0]),.doutb(w_n4918_0[1]),.din(n4918));
	jspl jspl_w_n4926_0(.douta(w_n4926_0[0]),.doutb(w_n4926_0[1]),.din(n4926));
	jspl jspl_w_n4927_0(.douta(w_n4927_0[0]),.doutb(w_n4927_0[1]),.din(n4927));
	jspl jspl_w_n4928_0(.douta(w_n4928_0[0]),.doutb(w_n4928_0[1]),.din(n4928));
	jspl jspl_w_n4929_0(.douta(w_n4929_0[0]),.doutb(w_n4929_0[1]),.din(n4929));
	jspl3 jspl3_w_n4930_0(.douta(w_n4930_0[0]),.doutb(w_n4930_0[1]),.doutc(w_n4930_0[2]),.din(n4930));
	jspl jspl_w_n4931_0(.douta(w_n4931_0[0]),.doutb(w_n4931_0[1]),.din(n4931));
	jspl jspl_w_n4932_0(.douta(w_n4932_0[0]),.doutb(w_n4932_0[1]),.din(n4932));
	jspl jspl_w_n4933_0(.douta(w_n4933_0[0]),.doutb(w_n4933_0[1]),.din(n4933));
	jspl jspl_w_n4934_0(.douta(w_dff_A_c4lpFFo59_0),.doutb(w_n4934_0[1]),.din(n4934));
	jspl jspl_w_n4937_0(.douta(w_n4937_0[0]),.doutb(w_n4937_0[1]),.din(n4937));
	jspl jspl_w_n4938_0(.douta(w_n4938_0[0]),.doutb(w_n4938_0[1]),.din(n4938));
	jspl jspl_w_n4940_0(.douta(w_n4940_0[0]),.doutb(w_n4940_0[1]),.din(n4940));
	jspl jspl_w_n4952_0(.douta(w_n4952_0[0]),.doutb(w_n4952_0[1]),.din(n4952));
	jspl jspl_w_n4953_0(.douta(w_n4953_0[0]),.doutb(w_n4953_0[1]),.din(n4953));
	jspl jspl_w_n4956_0(.douta(w_n4956_0[0]),.doutb(w_n4956_0[1]),.din(n4956));
	jspl jspl_w_n4961_0(.douta(w_n4961_0[0]),.doutb(w_n4961_0[1]),.din(n4961));
	jspl jspl_w_n4969_0(.douta(w_n4969_0[0]),.doutb(w_n4969_0[1]),.din(n4969));
	jspl3 jspl3_w_n4970_0(.douta(w_n4970_0[0]),.doutb(w_n4970_0[1]),.doutc(w_n4970_0[2]),.din(n4970));
	jspl jspl_w_n4972_0(.douta(w_n4972_0[0]),.doutb(w_n4972_0[1]),.din(n4972));
	jspl jspl_w_n4974_0(.douta(w_n4974_0[0]),.doutb(w_n4974_0[1]),.din(n4974));
	jspl jspl_w_n4982_0(.douta(w_n4982_0[0]),.doutb(w_n4982_0[1]),.din(n4982));
	jspl jspl_w_n4983_0(.douta(w_n4983_0[0]),.doutb(w_n4983_0[1]),.din(n4983));
	jspl jspl_w_n4988_0(.douta(w_n4988_0[0]),.doutb(w_n4988_0[1]),.din(n4988));
	jspl jspl_w_n4996_0(.douta(w_n4996_0[0]),.doutb(w_n4996_0[1]),.din(n4996));
	jspl jspl_w_n4997_0(.douta(w_n4997_0[0]),.doutb(w_n4997_0[1]),.din(n4997));
	jspl jspl_w_n4998_0(.douta(w_n4998_0[0]),.doutb(w_n4998_0[1]),.din(n4998));
	jspl jspl_w_n4999_0(.douta(w_n4999_0[0]),.doutb(w_n4999_0[1]),.din(n4999));
	jspl3 jspl3_w_n5000_0(.douta(w_n5000_0[0]),.doutb(w_n5000_0[1]),.doutc(w_n5000_0[2]),.din(n5000));
	jspl jspl_w_n5001_0(.douta(w_n5001_0[0]),.doutb(w_n5001_0[1]),.din(n5001));
	jspl jspl_w_n5002_0(.douta(w_n5002_0[0]),.doutb(w_n5002_0[1]),.din(n5002));
	jspl jspl_w_n5003_0(.douta(w_n5003_0[0]),.doutb(w_n5003_0[1]),.din(n5003));
	jspl jspl_w_n5004_0(.douta(w_dff_A_AlQfCFvp1_0),.doutb(w_n5004_0[1]),.din(n5004));
	jspl jspl_w_n5007_0(.douta(w_n5007_0[0]),.doutb(w_n5007_0[1]),.din(n5007));
	jspl jspl_w_n5008_0(.douta(w_n5008_0[0]),.doutb(w_n5008_0[1]),.din(n5008));
	jspl jspl_w_n5010_0(.douta(w_n5010_0[0]),.doutb(w_n5010_0[1]),.din(n5010));
	jspl jspl_w_n5016_0(.douta(w_n5016_0[0]),.doutb(w_n5016_0[1]),.din(n5016));
	jspl jspl_w_n5017_0(.douta(w_n5017_0[0]),.doutb(w_n5017_0[1]),.din(n5017));
	jspl jspl_w_n5020_0(.douta(w_n5020_0[0]),.doutb(w_n5020_0[1]),.din(n5020));
	jspl jspl_w_n5023_0(.douta(w_n5023_0[0]),.doutb(w_n5023_0[1]),.din(n5023));
	jspl jspl_w_n5028_0(.douta(w_n5028_0[0]),.doutb(w_n5028_0[1]),.din(n5028));
	jspl jspl_w_n5029_0(.douta(w_n5029_0[0]),.doutb(w_n5029_0[1]),.din(n5029));
	jspl jspl_w_n5030_0(.douta(w_n5030_0[0]),.doutb(w_n5030_0[1]),.din(n5030));
	jspl jspl_w_n5034_0(.douta(w_n5034_0[0]),.doutb(w_n5034_0[1]),.din(n5034));
	jspl jspl_w_n5035_0(.douta(w_n5035_0[0]),.doutb(w_n5035_0[1]),.din(n5035));
	jspl jspl_w_n5043_0(.douta(w_n5043_0[0]),.doutb(w_n5043_0[1]),.din(n5043));
	jspl jspl_w_n5044_0(.douta(w_n5044_0[0]),.doutb(w_n5044_0[1]),.din(n5044));
	jspl jspl_w_n5045_0(.douta(w_n5045_0[0]),.doutb(w_n5045_0[1]),.din(n5045));
	jspl jspl_w_n5051_0(.douta(w_n5051_0[0]),.doutb(w_n5051_0[1]),.din(n5051));
	jspl jspl_w_n5052_0(.douta(w_n5052_0[0]),.doutb(w_n5052_0[1]),.din(n5052));
	jspl jspl_w_n5053_0(.douta(w_n5053_0[0]),.doutb(w_n5053_0[1]),.din(n5053));
	jspl3 jspl3_w_n5054_0(.douta(w_n5054_0[0]),.doutb(w_n5054_0[1]),.doutc(w_n5054_0[2]),.din(n5054));
	jspl jspl_w_n5055_0(.douta(w_n5055_0[0]),.doutb(w_n5055_0[1]),.din(n5055));
	jspl jspl_w_n5056_0(.douta(w_n5056_0[0]),.doutb(w_n5056_0[1]),.din(n5056));
	jspl jspl_w_n5057_0(.douta(w_n5057_0[0]),.doutb(w_n5057_0[1]),.din(n5057));
	jspl jspl_w_n5058_0(.douta(w_dff_A_vrPoZQgf4_0),.doutb(w_n5058_0[1]),.din(n5058));
	jspl jspl_w_n5061_0(.douta(w_n5061_0[0]),.doutb(w_n5061_0[1]),.din(n5061));
	jspl jspl_w_n5062_0(.douta(w_n5062_0[0]),.doutb(w_n5062_0[1]),.din(n5062));
	jspl jspl_w_n5064_0(.douta(w_n5064_0[0]),.doutb(w_n5064_0[1]),.din(n5064));
	jspl jspl_w_n5070_0(.douta(w_n5070_0[0]),.doutb(w_n5070_0[1]),.din(n5070));
	jspl jspl_w_n5076_0(.douta(w_n5076_0[0]),.doutb(w_n5076_0[1]),.din(n5076));
	jspl jspl_w_n5077_0(.douta(w_n5077_0[0]),.doutb(w_n5077_0[1]),.din(n5077));
	jspl jspl_w_n5080_0(.douta(w_n5080_0[0]),.doutb(w_n5080_0[1]),.din(n5080));
	jspl jspl_w_n5083_0(.douta(w_n5083_0[0]),.doutb(w_n5083_0[1]),.din(n5083));
	jspl jspl_w_n5088_0(.douta(w_n5088_0[0]),.doutb(w_n5088_0[1]),.din(n5088));
	jspl jspl_w_n5096_0(.douta(w_n5096_0[0]),.doutb(w_n5096_0[1]),.din(n5096));
	jspl jspl_w_n5097_0(.douta(w_n5097_0[0]),.doutb(w_n5097_0[1]),.din(n5097));
	jspl jspl_w_n5100_0(.douta(w_n5100_0[0]),.doutb(w_n5100_0[1]),.din(n5100));
	jspl jspl_w_n5101_0(.douta(w_n5101_0[0]),.doutb(w_n5101_0[1]),.din(n5101));
	jspl3 jspl3_w_n5102_0(.douta(w_n5102_0[0]),.doutb(w_n5102_0[1]),.doutc(w_n5102_0[2]),.din(n5102));
	jspl jspl_w_n5105_0(.douta(w_n5105_0[0]),.doutb(w_n5105_0[1]),.din(n5105));
	jspl jspl_w_n5106_0(.douta(w_n5106_0[0]),.doutb(w_n5106_0[1]),.din(n5106));
	jspl jspl_w_n5107_0(.douta(w_n5107_0[0]),.doutb(w_n5107_0[1]),.din(n5107));
	jspl jspl_w_n5108_0(.douta(w_n5108_0[0]),.doutb(w_n5108_0[1]),.din(n5108));
	jspl3 jspl3_w_n5109_0(.douta(w_n5109_0[0]),.doutb(w_n5109_0[1]),.doutc(w_n5109_0[2]),.din(n5109));
	jspl jspl_w_n5110_0(.douta(w_n5110_0[0]),.doutb(w_n5110_0[1]),.din(n5110));
	jspl jspl_w_n5111_0(.douta(w_n5111_0[0]),.doutb(w_n5111_0[1]),.din(n5111));
	jspl jspl_w_n5112_0(.douta(w_n5112_0[0]),.doutb(w_n5112_0[1]),.din(n5112));
	jspl jspl_w_n5113_0(.douta(w_dff_A_A2xONnuD7_0),.doutb(w_n5113_0[1]),.din(n5113));
	jspl jspl_w_n5116_0(.douta(w_n5116_0[0]),.doutb(w_n5116_0[1]),.din(n5116));
	jspl jspl_w_n5117_0(.douta(w_n5117_0[0]),.doutb(w_n5117_0[1]),.din(n5117));
	jspl jspl_w_n5119_0(.douta(w_n5119_0[0]),.doutb(w_n5119_0[1]),.din(n5119));
	jspl jspl_w_n5122_0(.douta(w_n5122_0[0]),.doutb(w_n5122_0[1]),.din(n5122));
	jspl jspl_w_n5134_0(.douta(w_n5134_0[0]),.doutb(w_n5134_0[1]),.din(n5134));
	jspl jspl_w_n5135_0(.douta(w_n5135_0[0]),.doutb(w_n5135_0[1]),.din(n5135));
	jspl jspl_w_n5138_0(.douta(w_n5138_0[0]),.doutb(w_n5138_0[1]),.din(n5138));
	jspl jspl_w_n5143_0(.douta(w_n5143_0[0]),.doutb(w_n5143_0[1]),.din(n5143));
	jspl jspl_w_n5145_0(.douta(w_n5145_0[0]),.doutb(w_n5145_0[1]),.din(n5145));
	jspl jspl_w_n5146_0(.douta(w_n5146_0[0]),.doutb(w_n5146_0[1]),.din(n5146));
	jspl jspl_w_n5147_0(.douta(w_n5147_0[0]),.doutb(w_n5147_0[1]),.din(n5147));
	jspl jspl_w_n5148_0(.douta(w_n5148_0[0]),.doutb(w_n5148_0[1]),.din(n5148));
	jspl jspl_w_n5156_0(.douta(w_n5156_0[0]),.doutb(w_n5156_0[1]),.din(n5156));
	jspl jspl_w_n5157_0(.douta(w_n5157_0[0]),.doutb(w_n5157_0[1]),.din(n5157));
	jspl jspl_w_n5158_0(.douta(w_n5158_0[0]),.doutb(w_n5158_0[1]),.din(n5158));
	jspl jspl_w_n5159_0(.douta(w_n5159_0[0]),.doutb(w_n5159_0[1]),.din(n5159));
	jspl3 jspl3_w_n5160_0(.douta(w_n5160_0[0]),.doutb(w_n5160_0[1]),.doutc(w_n5160_0[2]),.din(n5160));
	jspl jspl_w_n5161_0(.douta(w_n5161_0[0]),.doutb(w_n5161_0[1]),.din(n5161));
	jspl jspl_w_n5162_0(.douta(w_n5162_0[0]),.doutb(w_n5162_0[1]),.din(n5162));
	jspl jspl_w_n5163_0(.douta(w_n5163_0[0]),.doutb(w_n5163_0[1]),.din(n5163));
	jspl jspl_w_n5164_0(.douta(w_dff_A_zf31BzpE2_0),.doutb(w_n5164_0[1]),.din(n5164));
	jspl jspl_w_n5167_0(.douta(w_n5167_0[0]),.doutb(w_n5167_0[1]),.din(n5167));
	jspl jspl_w_n5168_0(.douta(w_n5168_0[0]),.doutb(w_n5168_0[1]),.din(n5168));
	jspl jspl_w_n5170_0(.douta(w_n5170_0[0]),.doutb(w_n5170_0[1]),.din(n5170));
	jspl jspl_w_n5184_0(.douta(w_n5184_0[0]),.doutb(w_n5184_0[1]),.din(n5184));
	jspl jspl_w_n5185_0(.douta(w_n5185_0[0]),.doutb(w_n5185_0[1]),.din(n5185));
	jspl jspl_w_n5188_0(.douta(w_n5188_0[0]),.doutb(w_n5188_0[1]),.din(n5188));
	jspl jspl_w_n5191_0(.douta(w_n5191_0[0]),.doutb(w_n5191_0[1]),.din(n5191));
	jspl jspl_w_n5193_0(.douta(w_n5193_0[0]),.doutb(w_n5193_0[1]),.din(n5193));
	jspl jspl_w_n5196_0(.douta(w_n5196_0[0]),.doutb(w_n5196_0[1]),.din(n5196));
	jspl jspl_w_n5197_0(.douta(w_n5197_0[0]),.doutb(w_n5197_0[1]),.din(n5197));
	jspl jspl_w_n5203_0(.douta(w_n5203_0[0]),.doutb(w_n5203_0[1]),.din(n5203));
	jspl jspl_w_n5204_0(.douta(w_n5204_0[0]),.doutb(w_n5204_0[1]),.din(n5204));
	jspl jspl_w_n5205_0(.douta(w_n5205_0[0]),.doutb(w_n5205_0[1]),.din(n5205));
	jspl3 jspl3_w_n5206_0(.douta(w_n5206_0[0]),.doutb(w_n5206_0[1]),.doutc(w_n5206_0[2]),.din(n5206));
	jspl jspl_w_n5207_0(.douta(w_n5207_0[0]),.doutb(w_n5207_0[1]),.din(n5207));
	jspl jspl_w_n5208_0(.douta(w_n5208_0[0]),.doutb(w_n5208_0[1]),.din(n5208));
	jspl jspl_w_n5209_0(.douta(w_n5209_0[0]),.doutb(w_n5209_0[1]),.din(n5209));
	jspl jspl_w_n5210_0(.douta(w_dff_A_bxvqYTYx4_0),.doutb(w_n5210_0[1]),.din(n5210));
	jspl jspl_w_n5213_0(.douta(w_n5213_0[0]),.doutb(w_n5213_0[1]),.din(n5213));
	jspl jspl_w_n5214_0(.douta(w_n5214_0[0]),.doutb(w_n5214_0[1]),.din(n5214));
	jspl jspl_w_n5216_0(.douta(w_n5216_0[0]),.doutb(w_n5216_0[1]),.din(n5216));
	jspl jspl_w_n5219_0(.douta(w_n5219_0[0]),.doutb(w_n5219_0[1]),.din(n5219));
	jspl jspl_w_n5229_0(.douta(w_n5229_0[0]),.doutb(w_n5229_0[1]),.din(n5229));
	jspl jspl_w_n5230_0(.douta(w_n5230_0[0]),.doutb(w_n5230_0[1]),.din(n5230));
	jspl jspl_w_n5233_0(.douta(w_n5233_0[0]),.doutb(w_n5233_0[1]),.din(n5233));
	jspl3 jspl3_w_n5236_0(.douta(w_n5236_0[0]),.doutb(w_n5236_0[1]),.doutc(w_n5236_0[2]),.din(n5236));
	jspl jspl_w_n5238_0(.douta(w_n5238_0[0]),.doutb(w_n5238_0[1]),.din(n5238));
	jspl jspl_w_n5239_0(.douta(w_n5239_0[0]),.doutb(w_n5239_0[1]),.din(n5239));
	jspl jspl_w_n5240_0(.douta(w_n5240_0[0]),.doutb(w_n5240_0[1]),.din(n5240));
	jspl jspl_w_n5243_0(.douta(w_n5243_0[0]),.doutb(w_n5243_0[1]),.din(n5243));
	jspl3 jspl3_w_n5244_0(.douta(w_n5244_0[0]),.doutb(w_n5244_0[1]),.doutc(w_n5244_0[2]),.din(n5244));
	jspl jspl_w_n5245_0(.douta(w_n5245_0[0]),.doutb(w_n5245_0[1]),.din(n5245));
	jspl jspl_w_n5246_0(.douta(w_n5246_0[0]),.doutb(w_n5246_0[1]),.din(n5246));
	jspl jspl_w_n5247_0(.douta(w_n5247_0[0]),.doutb(w_n5247_0[1]),.din(n5247));
	jspl jspl_w_n5248_0(.douta(w_dff_A_ruo15GOT6_0),.doutb(w_n5248_0[1]),.din(n5248));
	jspl jspl_w_n5252_0(.douta(w_n5252_0[0]),.doutb(w_n5252_0[1]),.din(n5252));
	jspl jspl_w_n5253_0(.douta(w_n5253_0[0]),.doutb(w_n5253_0[1]),.din(n5253));
	jspl jspl_w_n5323_0(.douta(w_n5323_0[0]),.doutb(w_n5323_0[1]),.din(n5323));
	jspl3 jspl3_w_n5332_0(.douta(w_n5332_0[0]),.doutb(w_n5332_0[1]),.doutc(w_n5332_0[2]),.din(n5332));
	jspl jspl_w_n5332_1(.douta(w_n5332_1[0]),.doutb(w_n5332_1[1]),.din(w_n5332_0[0]));
	jspl jspl_w_n5334_0(.douta(w_n5334_0[0]),.doutb(w_n5334_0[1]),.din(n5334));
	jspl jspl_w_n5346_0(.douta(w_n5346_0[0]),.doutb(w_n5346_0[1]),.din(n5346));
	jspl3 jspl3_w_n5347_0(.douta(w_n5347_0[0]),.doutb(w_n5347_0[1]),.doutc(w_n5347_0[2]),.din(n5347));
	jspl jspl_w_n5349_0(.douta(w_n5349_0[0]),.doutb(w_n5349_0[1]),.din(n5349));
	jspl jspl_w_n5350_0(.douta(w_n5350_0[0]),.doutb(w_n5350_0[1]),.din(n5350));
	jspl jspl_w_n5351_0(.douta(w_dff_A_ghwMUcgR8_0),.doutb(w_n5351_0[1]),.din(n5351));
	jspl jspl_w_n5354_0(.douta(w_dff_A_0wlIeazr9_0),.doutb(w_n5354_0[1]),.din(n5354));
	jspl jspl_w_n5356_0(.douta(w_n5356_0[0]),.doutb(w_n5356_0[1]),.din(n5356));
	jspl jspl_w_n5357_0(.douta(w_n5357_0[0]),.doutb(w_n5357_0[1]),.din(n5357));
	jspl3 jspl3_w_n5368_0(.douta(w_n5368_0[0]),.doutb(w_n5368_0[1]),.doutc(w_n5368_0[2]),.din(n5368));
	jspl jspl_w_n5369_0(.douta(w_n5369_0[0]),.doutb(w_n5369_0[1]),.din(n5369));
	jspl jspl_w_n5370_0(.douta(w_n5370_0[0]),.doutb(w_n5370_0[1]),.din(n5370));
	jspl jspl_w_n5371_0(.douta(w_n5371_0[0]),.doutb(w_n5371_0[1]),.din(n5371));
	jspl3 jspl3_w_n5377_0(.douta(w_n5377_0[0]),.doutb(w_n5377_0[1]),.doutc(w_n5377_0[2]),.din(n5377));
	jspl jspl_w_n5378_0(.douta(w_n5378_0[0]),.doutb(w_n5378_0[1]),.din(n5378));
	jspl jspl_w_n5379_0(.douta(w_n5379_0[0]),.doutb(w_n5379_0[1]),.din(n5379));
	jspl3 jspl3_w_n5390_0(.douta(w_n5390_0[0]),.doutb(w_n5390_0[1]),.doutc(w_n5390_0[2]),.din(n5390));
	jspl jspl_w_n5390_1(.douta(w_n5390_1[0]),.doutb(w_n5390_1[1]),.din(w_n5390_0[0]));
	jspl jspl_w_n5395_0(.douta(w_n5395_0[0]),.doutb(w_n5395_0[1]),.din(n5395));
	jspl jspl_w_n5397_0(.douta(w_n5397_0[0]),.doutb(w_n5397_0[1]),.din(n5397));
	jspl jspl_w_n5398_0(.douta(w_n5398_0[0]),.doutb(w_n5398_0[1]),.din(n5398));
	jspl jspl_w_n5399_0(.douta(w_n5399_0[0]),.doutb(w_n5399_0[1]),.din(n5399));
	jspl3 jspl3_w_n5400_0(.douta(w_n5400_0[0]),.doutb(w_dff_A_jveqLtSa7_1),.doutc(w_n5400_0[2]),.din(n5400));
	jspl3 jspl3_w_n5404_0(.douta(w_n5404_0[0]),.doutb(w_n5404_0[1]),.doutc(w_n5404_0[2]),.din(n5404));
	jspl jspl_w_n5405_0(.douta(w_n5405_0[0]),.doutb(w_n5405_0[1]),.din(n5405));
	jspl jspl_w_n5406_0(.douta(w_n5406_0[0]),.doutb(w_n5406_0[1]),.din(n5406));
	jspl3 jspl3_w_n5415_0(.douta(w_n5415_0[0]),.doutb(w_n5415_0[1]),.doutc(w_n5415_0[2]),.din(n5415));
	jspl jspl_w_n5415_1(.douta(w_n5415_1[0]),.doutb(w_n5415_1[1]),.din(w_n5415_0[0]));
	jspl jspl_w_n5416_0(.douta(w_n5416_0[0]),.doutb(w_n5416_0[1]),.din(n5416));
	jspl3 jspl3_w_n5417_0(.douta(w_n5417_0[0]),.doutb(w_n5417_0[1]),.doutc(w_n5417_0[2]),.din(n5417));
	jspl jspl_w_n5418_0(.douta(w_n5418_0[0]),.doutb(w_n5418_0[1]),.din(n5418));
	jspl jspl_w_n5421_0(.douta(w_n5421_0[0]),.doutb(w_n5421_0[1]),.din(n5421));
	jspl3 jspl3_w_n5431_0(.douta(w_n5431_0[0]),.doutb(w_n5431_0[1]),.doutc(w_n5431_0[2]),.din(n5431));
	jspl3 jspl3_w_n5432_0(.douta(w_n5432_0[0]),.doutb(w_n5432_0[1]),.doutc(w_n5432_0[2]),.din(n5432));
	jspl jspl_w_n5435_0(.douta(w_n5435_0[0]),.doutb(w_n5435_0[1]),.din(n5435));
	jspl jspl_w_n5437_0(.douta(w_n5437_0[0]),.doutb(w_n5437_0[1]),.din(n5437));
	jspl3 jspl3_w_n5438_0(.douta(w_n5438_0[0]),.doutb(w_n5438_0[1]),.doutc(w_n5438_0[2]),.din(n5438));
	jspl jspl_w_n5440_0(.douta(w_n5440_0[0]),.doutb(w_dff_A_JzuBWyFX9_1),.din(n5440));
	jspl jspl_w_n5441_0(.douta(w_n5441_0[0]),.doutb(w_n5441_0[1]),.din(n5441));
	jspl jspl_w_n5444_0(.douta(w_n5444_0[0]),.doutb(w_n5444_0[1]),.din(n5444));
	jspl jspl_w_n5446_0(.douta(w_n5446_0[0]),.doutb(w_n5446_0[1]),.din(n5446));
	jspl jspl_w_n5447_0(.douta(w_n5447_0[0]),.doutb(w_n5447_0[1]),.din(n5447));
	jspl jspl_w_n5449_0(.douta(w_n5449_0[0]),.doutb(w_n5449_0[1]),.din(n5449));
	jspl3 jspl3_w_n5452_0(.douta(w_n5452_0[0]),.doutb(w_n5452_0[1]),.doutc(w_n5452_0[2]),.din(n5452));
	jspl jspl_w_n5452_1(.douta(w_n5452_1[0]),.doutb(w_n5452_1[1]),.din(w_n5452_0[0]));
	jspl jspl_w_n5453_0(.douta(w_n5453_0[0]),.doutb(w_n5453_0[1]),.din(n5453));
	jspl3 jspl3_w_n5454_0(.douta(w_n5454_0[0]),.doutb(w_n5454_0[1]),.doutc(w_n5454_0[2]),.din(n5454));
	jspl jspl_w_n5455_0(.douta(w_n5455_0[0]),.doutb(w_n5455_0[1]),.din(n5455));
	jspl jspl_w_n5458_0(.douta(w_n5458_0[0]),.doutb(w_n5458_0[1]),.din(n5458));
	jspl3 jspl3_w_n5459_0(.douta(w_n5459_0[0]),.doutb(w_n5459_0[1]),.doutc(w_n5459_0[2]),.din(n5459));
	jspl jspl_w_n5461_0(.douta(w_n5461_0[0]),.doutb(w_n5461_0[1]),.din(n5461));
	jspl3 jspl3_w_n5462_0(.douta(w_n5462_0[0]),.doutb(w_n5462_0[1]),.doutc(w_n5462_0[2]),.din(n5462));
	jspl jspl_w_n5463_0(.douta(w_n5463_0[0]),.doutb(w_n5463_0[1]),.din(n5463));
	jspl jspl_w_n5465_0(.douta(w_n5465_0[0]),.doutb(w_n5465_0[1]),.din(n5465));
	jspl jspl_w_n5466_0(.douta(w_n5466_0[0]),.doutb(w_n5466_0[1]),.din(n5466));
	jspl jspl_w_n5470_0(.douta(w_n5470_0[0]),.doutb(w_n5470_0[1]),.din(n5470));
	jspl jspl_w_n5471_0(.douta(w_n5471_0[0]),.doutb(w_n5471_0[1]),.din(n5471));
	jspl jspl_w_n5474_0(.douta(w_n5474_0[0]),.doutb(w_n5474_0[1]),.din(n5474));
	jspl jspl_w_n5476_0(.douta(w_dff_A_9fZQPXhh0_0),.doutb(w_n5476_0[1]),.din(n5476));
	jspl jspl_w_n5480_0(.douta(w_n5480_0[0]),.doutb(w_dff_A_Ms0ywCUm8_1),.din(w_dff_B_rKPkvx055_2));
	jspl jspl_w_n5483_0(.douta(w_n5483_0[0]),.doutb(w_n5483_0[1]),.din(n5483));
	jspl jspl_w_n5484_0(.douta(w_n5484_0[0]),.doutb(w_n5484_0[1]),.din(n5484));
	jspl jspl_w_n5487_0(.douta(w_n5487_0[0]),.doutb(w_n5487_0[1]),.din(n5487));
	jdff dff_A_nhphmE1W6_0(.dout(w_n4094_0[0]),.din(w_dff_A_nhphmE1W6_0),.clk(gclk));
	jdff dff_A_aq1r8Nrv9_0(.dout(w_n4093_11[0]),.din(w_dff_A_aq1r8Nrv9_0),.clk(gclk));
	jdff dff_A_BnrGsSKY8_0(.dout(w_dff_A_aq1r8Nrv9_0),.din(w_dff_A_BnrGsSKY8_0),.clk(gclk));
	jdff dff_A_9OrtdDC35_0(.dout(w_dff_A_BnrGsSKY8_0),.din(w_dff_A_9OrtdDC35_0),.clk(gclk));
	jdff dff_A_GI8REpUn5_0(.dout(w_n4093_10[0]),.din(w_dff_A_GI8REpUn5_0),.clk(gclk));
	jdff dff_A_i9IctGI95_0(.dout(w_dff_A_GI8REpUn5_0),.din(w_dff_A_i9IctGI95_0),.clk(gclk));
	jdff dff_A_IuwzUmsQ4_0(.dout(w_dff_A_i9IctGI95_0),.din(w_dff_A_IuwzUmsQ4_0),.clk(gclk));
	jdff dff_A_k4Whxaqa7_0(.dout(w_dff_A_IuwzUmsQ4_0),.din(w_dff_A_k4Whxaqa7_0),.clk(gclk));
	jdff dff_A_H7NfKn0e1_1(.dout(w_n4093_10[1]),.din(w_dff_A_H7NfKn0e1_1),.clk(gclk));
	jdff dff_A_8u2TGooJ9_1(.dout(w_dff_A_H7NfKn0e1_1),.din(w_dff_A_8u2TGooJ9_1),.clk(gclk));
	jdff dff_A_zthfvi4X4_0(.dout(w_n4093_9[0]),.din(w_dff_A_zthfvi4X4_0),.clk(gclk));
	jdff dff_A_STnUsJAO6_0(.dout(w_dff_A_zthfvi4X4_0),.din(w_dff_A_STnUsJAO6_0),.clk(gclk));
	jdff dff_A_MPoSOk006_0(.dout(w_dff_A_STnUsJAO6_0),.din(w_dff_A_MPoSOk006_0),.clk(gclk));
	jdff dff_A_AZO8FXmC7_0(.dout(w_dff_A_MPoSOk006_0),.din(w_dff_A_AZO8FXmC7_0),.clk(gclk));
	jdff dff_A_mfNsh70O0_1(.dout(w_n4093_9[1]),.din(w_dff_A_mfNsh70O0_1),.clk(gclk));
	jdff dff_A_wpA3GKq05_1(.dout(w_dff_A_mfNsh70O0_1),.din(w_dff_A_wpA3GKq05_1),.clk(gclk));
	jdff dff_A_MITM5qKS5_0(.dout(w_n4093_8[0]),.din(w_dff_A_MITM5qKS5_0),.clk(gclk));
	jdff dff_A_CfbEZi267_0(.dout(w_dff_A_MITM5qKS5_0),.din(w_dff_A_CfbEZi267_0),.clk(gclk));
	jdff dff_A_Ee8k0hks1_0(.dout(w_dff_A_CfbEZi267_0),.din(w_dff_A_Ee8k0hks1_0),.clk(gclk));
	jdff dff_A_cUDtSJyJ3_0(.dout(w_dff_A_Ee8k0hks1_0),.din(w_dff_A_cUDtSJyJ3_0),.clk(gclk));
	jdff dff_A_DRpHc2cG9_1(.dout(w_n4093_8[1]),.din(w_dff_A_DRpHc2cG9_1),.clk(gclk));
	jdff dff_A_BPbGrQYz5_1(.dout(w_dff_A_DRpHc2cG9_1),.din(w_dff_A_BPbGrQYz5_1),.clk(gclk));
	jdff dff_A_Dd9u7gyD3_0(.dout(w_n4093_7[0]),.din(w_dff_A_Dd9u7gyD3_0),.clk(gclk));
	jdff dff_A_lq02Zg2a4_0(.dout(w_dff_A_Dd9u7gyD3_0),.din(w_dff_A_lq02Zg2a4_0),.clk(gclk));
	jdff dff_A_KCQwo8UC3_0(.dout(w_dff_A_lq02Zg2a4_0),.din(w_dff_A_KCQwo8UC3_0),.clk(gclk));
	jdff dff_A_xH2PJntQ0_0(.dout(w_dff_A_KCQwo8UC3_0),.din(w_dff_A_xH2PJntQ0_0),.clk(gclk));
	jdff dff_A_TJ7EiHcb4_1(.dout(w_n4093_7[1]),.din(w_dff_A_TJ7EiHcb4_1),.clk(gclk));
	jdff dff_A_55rtkZ763_1(.dout(w_dff_A_TJ7EiHcb4_1),.din(w_dff_A_55rtkZ763_1),.clk(gclk));
	jdff dff_A_Bg5Nu4RH8_0(.dout(w_n4093_2[0]),.din(w_dff_A_Bg5Nu4RH8_0),.clk(gclk));
	jdff dff_A_pThksnDn4_0(.dout(w_dff_A_Bg5Nu4RH8_0),.din(w_dff_A_pThksnDn4_0),.clk(gclk));
	jdff dff_A_yQupp8fW5_0(.dout(w_dff_A_pThksnDn4_0),.din(w_dff_A_yQupp8fW5_0),.clk(gclk));
	jdff dff_A_B2o3GbHy5_0(.dout(w_dff_A_yQupp8fW5_0),.din(w_dff_A_B2o3GbHy5_0),.clk(gclk));
	jdff dff_A_ppYAdYzc9_0(.dout(w_dff_A_B2o3GbHy5_0),.din(w_dff_A_ppYAdYzc9_0),.clk(gclk));
	jdff dff_A_ygimsAm25_0(.dout(w_dff_A_ppYAdYzc9_0),.din(w_dff_A_ygimsAm25_0),.clk(gclk));
	jdff dff_A_GkIFZOZv8_0(.dout(w_dff_A_ygimsAm25_0),.din(w_dff_A_GkIFZOZv8_0),.clk(gclk));
	jdff dff_A_MzbPBSaa5_0(.dout(w_dff_A_GkIFZOZv8_0),.din(w_dff_A_MzbPBSaa5_0),.clk(gclk));
	jdff dff_A_xKT4koJY9_0(.dout(w_dff_A_MzbPBSaa5_0),.din(w_dff_A_xKT4koJY9_0),.clk(gclk));
	jdff dff_A_lykm64H75_0(.dout(w_dff_A_xKT4koJY9_0),.din(w_dff_A_lykm64H75_0),.clk(gclk));
	jdff dff_A_rj3wy9UT4_0(.dout(w_dff_A_lykm64H75_0),.din(w_dff_A_rj3wy9UT4_0),.clk(gclk));
	jdff dff_A_fbO785X92_0(.dout(w_dff_A_rj3wy9UT4_0),.din(w_dff_A_fbO785X92_0),.clk(gclk));
	jdff dff_A_Bppkcx0L3_1(.dout(w_n4093_2[1]),.din(w_dff_A_Bppkcx0L3_1),.clk(gclk));
	jdff dff_A_bDwv7Pyo2_1(.dout(w_dff_A_Bppkcx0L3_1),.din(w_dff_A_bDwv7Pyo2_1),.clk(gclk));
	jdff dff_A_EdZtp1rz5_1(.dout(w_dff_A_bDwv7Pyo2_1),.din(w_dff_A_EdZtp1rz5_1),.clk(gclk));
	jdff dff_A_Yd2y2bpJ5_1(.dout(w_dff_A_EdZtp1rz5_1),.din(w_dff_A_Yd2y2bpJ5_1),.clk(gclk));
	jdff dff_A_TQJu4EWX8_1(.dout(w_dff_A_Yd2y2bpJ5_1),.din(w_dff_A_TQJu4EWX8_1),.clk(gclk));
	jdff dff_A_9NWZDZCv5_1(.dout(w_dff_A_TQJu4EWX8_1),.din(w_dff_A_9NWZDZCv5_1),.clk(gclk));
	jdff dff_B_qpX2ZoCZ3_0(.din(n5352),.dout(w_dff_B_qpX2ZoCZ3_0),.clk(gclk));
	jdff dff_A_g1w0aTHP1_0(.dout(w_n4093_6[0]),.din(w_dff_A_g1w0aTHP1_0),.clk(gclk));
	jdff dff_A_urx9Osvr5_0(.dout(w_dff_A_g1w0aTHP1_0),.din(w_dff_A_urx9Osvr5_0),.clk(gclk));
	jdff dff_A_XhYdEVGP9_0(.dout(w_dff_A_urx9Osvr5_0),.din(w_dff_A_XhYdEVGP9_0),.clk(gclk));
	jdff dff_A_cAl4L0fX0_0(.dout(w_dff_A_XhYdEVGP9_0),.din(w_dff_A_cAl4L0fX0_0),.clk(gclk));
	jdff dff_A_8BQJrza76_0(.dout(w_dff_A_cAl4L0fX0_0),.din(w_dff_A_8BQJrza76_0),.clk(gclk));
	jdff dff_A_uFawYx0e7_1(.dout(w_n4093_6[1]),.din(w_dff_A_uFawYx0e7_1),.clk(gclk));
	jdff dff_A_imlgG5NP4_1(.dout(w_dff_A_uFawYx0e7_1),.din(w_dff_A_imlgG5NP4_1),.clk(gclk));
	jdff dff_A_KitWvW7m5_0(.dout(w_n4093_5[0]),.din(w_dff_A_KitWvW7m5_0),.clk(gclk));
	jdff dff_A_EUkGuJ364_0(.dout(w_dff_A_KitWvW7m5_0),.din(w_dff_A_EUkGuJ364_0),.clk(gclk));
	jdff dff_A_Iu0AqP8D9_0(.dout(w_dff_A_EUkGuJ364_0),.din(w_dff_A_Iu0AqP8D9_0),.clk(gclk));
	jdff dff_A_wOYd2JLH5_1(.dout(w_n4093_5[1]),.din(w_dff_A_wOYd2JLH5_1),.clk(gclk));
	jdff dff_A_suv5RVkp5_1(.dout(w_dff_A_wOYd2JLH5_1),.din(w_dff_A_suv5RVkp5_1),.clk(gclk));
	jdff dff_B_79XZBc8E3_1(.din(n5485),.dout(w_dff_B_79XZBc8E3_1),.clk(gclk));
	jdff dff_B_qjcjo5yK6_1(.din(w_dff_B_79XZBc8E3_1),.dout(w_dff_B_qjcjo5yK6_1),.clk(gclk));
	jdff dff_B_pNwtQMbW3_0(.din(n5503),.dout(w_dff_B_pNwtQMbW3_0),.clk(gclk));
	jdff dff_A_wA1LpPh75_1(.dout(w_n5480_0[1]),.din(w_dff_A_wA1LpPh75_1),.clk(gclk));
	jdff dff_A_rXux2KXN2_1(.dout(w_dff_A_wA1LpPh75_1),.din(w_dff_A_rXux2KXN2_1),.clk(gclk));
	jdff dff_A_Ms0ywCUm8_1(.dout(w_dff_A_rXux2KXN2_1),.din(w_dff_A_Ms0ywCUm8_1),.clk(gclk));
	jdff dff_B_1F1gfXBh4_2(.din(n5480),.dout(w_dff_B_1F1gfXBh4_2),.clk(gclk));
	jdff dff_B_VKoVih2S8_2(.din(w_dff_B_1F1gfXBh4_2),.dout(w_dff_B_VKoVih2S8_2),.clk(gclk));
	jdff dff_B_zipXXgMG7_2(.din(w_dff_B_VKoVih2S8_2),.dout(w_dff_B_zipXXgMG7_2),.clk(gclk));
	jdff dff_B_3Y7HE1ps2_2(.din(w_dff_B_zipXXgMG7_2),.dout(w_dff_B_3Y7HE1ps2_2),.clk(gclk));
	jdff dff_B_r7mfL8Xx3_2(.din(w_dff_B_3Y7HE1ps2_2),.dout(w_dff_B_r7mfL8Xx3_2),.clk(gclk));
	jdff dff_B_2ZCumULd4_2(.din(w_dff_B_r7mfL8Xx3_2),.dout(w_dff_B_2ZCumULd4_2),.clk(gclk));
	jdff dff_B_lgQ2CJpm0_2(.din(w_dff_B_2ZCumULd4_2),.dout(w_dff_B_lgQ2CJpm0_2),.clk(gclk));
	jdff dff_B_tCtVDcet3_2(.din(w_dff_B_lgQ2CJpm0_2),.dout(w_dff_B_tCtVDcet3_2),.clk(gclk));
	jdff dff_B_f8hVMZUo0_2(.din(w_dff_B_tCtVDcet3_2),.dout(w_dff_B_f8hVMZUo0_2),.clk(gclk));
	jdff dff_B_KcdrDF0c4_2(.din(w_dff_B_f8hVMZUo0_2),.dout(w_dff_B_KcdrDF0c4_2),.clk(gclk));
	jdff dff_B_TAg8WBza2_2(.din(w_dff_B_KcdrDF0c4_2),.dout(w_dff_B_TAg8WBza2_2),.clk(gclk));
	jdff dff_B_KrYqum444_2(.din(w_dff_B_TAg8WBza2_2),.dout(w_dff_B_KrYqum444_2),.clk(gclk));
	jdff dff_B_QG15WaUo1_2(.din(w_dff_B_KrYqum444_2),.dout(w_dff_B_QG15WaUo1_2),.clk(gclk));
	jdff dff_B_nx4o88U60_2(.din(w_dff_B_QG15WaUo1_2),.dout(w_dff_B_nx4o88U60_2),.clk(gclk));
	jdff dff_B_UhS4FA638_2(.din(w_dff_B_nx4o88U60_2),.dout(w_dff_B_UhS4FA638_2),.clk(gclk));
	jdff dff_B_JDNh7iiZ2_2(.din(w_dff_B_UhS4FA638_2),.dout(w_dff_B_JDNh7iiZ2_2),.clk(gclk));
	jdff dff_B_OxKRY7227_2(.din(w_dff_B_JDNh7iiZ2_2),.dout(w_dff_B_OxKRY7227_2),.clk(gclk));
	jdff dff_B_AU3fIqR25_2(.din(w_dff_B_OxKRY7227_2),.dout(w_dff_B_AU3fIqR25_2),.clk(gclk));
	jdff dff_B_Kth0DFSO8_2(.din(w_dff_B_AU3fIqR25_2),.dout(w_dff_B_Kth0DFSO8_2),.clk(gclk));
	jdff dff_B_g0gyRwvL0_2(.din(w_dff_B_Kth0DFSO8_2),.dout(w_dff_B_g0gyRwvL0_2),.clk(gclk));
	jdff dff_B_sHUH4X1Q0_2(.din(w_dff_B_g0gyRwvL0_2),.dout(w_dff_B_sHUH4X1Q0_2),.clk(gclk));
	jdff dff_B_DNAmQGUn9_2(.din(w_dff_B_sHUH4X1Q0_2),.dout(w_dff_B_DNAmQGUn9_2),.clk(gclk));
	jdff dff_B_aV2a0Cps4_2(.din(w_dff_B_DNAmQGUn9_2),.dout(w_dff_B_aV2a0Cps4_2),.clk(gclk));
	jdff dff_B_tZeRuOxq7_2(.din(w_dff_B_aV2a0Cps4_2),.dout(w_dff_B_tZeRuOxq7_2),.clk(gclk));
	jdff dff_B_3sZmPu2P2_2(.din(w_dff_B_tZeRuOxq7_2),.dout(w_dff_B_3sZmPu2P2_2),.clk(gclk));
	jdff dff_B_ZePAYJ262_2(.din(w_dff_B_3sZmPu2P2_2),.dout(w_dff_B_ZePAYJ262_2),.clk(gclk));
	jdff dff_B_T8xTOSvj0_2(.din(w_dff_B_ZePAYJ262_2),.dout(w_dff_B_T8xTOSvj0_2),.clk(gclk));
	jdff dff_B_n7qHaveF2_2(.din(w_dff_B_T8xTOSvj0_2),.dout(w_dff_B_n7qHaveF2_2),.clk(gclk));
	jdff dff_B_zzK0lWC83_2(.din(w_dff_B_n7qHaveF2_2),.dout(w_dff_B_zzK0lWC83_2),.clk(gclk));
	jdff dff_B_WAsBDibx6_2(.din(w_dff_B_zzK0lWC83_2),.dout(w_dff_B_WAsBDibx6_2),.clk(gclk));
	jdff dff_B_YtehPBPw5_2(.din(w_dff_B_WAsBDibx6_2),.dout(w_dff_B_YtehPBPw5_2),.clk(gclk));
	jdff dff_B_ZCj9Sgpe9_2(.din(w_dff_B_YtehPBPw5_2),.dout(w_dff_B_ZCj9Sgpe9_2),.clk(gclk));
	jdff dff_B_R9p6zXHr1_2(.din(w_dff_B_ZCj9Sgpe9_2),.dout(w_dff_B_R9p6zXHr1_2),.clk(gclk));
	jdff dff_B_rfl1FEMf9_2(.din(w_dff_B_R9p6zXHr1_2),.dout(w_dff_B_rfl1FEMf9_2),.clk(gclk));
	jdff dff_B_F7eW0GgV7_2(.din(w_dff_B_rfl1FEMf9_2),.dout(w_dff_B_F7eW0GgV7_2),.clk(gclk));
	jdff dff_B_aeFwX27L8_2(.din(w_dff_B_F7eW0GgV7_2),.dout(w_dff_B_aeFwX27L8_2),.clk(gclk));
	jdff dff_B_VRSTJzhP5_2(.din(w_dff_B_aeFwX27L8_2),.dout(w_dff_B_VRSTJzhP5_2),.clk(gclk));
	jdff dff_B_o3Y9g7EF3_2(.din(w_dff_B_VRSTJzhP5_2),.dout(w_dff_B_o3Y9g7EF3_2),.clk(gclk));
	jdff dff_B_jLQg0u2Q6_2(.din(w_dff_B_o3Y9g7EF3_2),.dout(w_dff_B_jLQg0u2Q6_2),.clk(gclk));
	jdff dff_B_GcjS3Fik0_2(.din(w_dff_B_jLQg0u2Q6_2),.dout(w_dff_B_GcjS3Fik0_2),.clk(gclk));
	jdff dff_B_gCZ78ql51_2(.din(w_dff_B_GcjS3Fik0_2),.dout(w_dff_B_gCZ78ql51_2),.clk(gclk));
	jdff dff_B_O8Z66YzX5_2(.din(w_dff_B_gCZ78ql51_2),.dout(w_dff_B_O8Z66YzX5_2),.clk(gclk));
	jdff dff_B_SZI9QF5N6_2(.din(w_dff_B_O8Z66YzX5_2),.dout(w_dff_B_SZI9QF5N6_2),.clk(gclk));
	jdff dff_B_FX9Tqe2G0_2(.din(w_dff_B_SZI9QF5N6_2),.dout(w_dff_B_FX9Tqe2G0_2),.clk(gclk));
	jdff dff_B_Vf48OteZ5_2(.din(w_dff_B_FX9Tqe2G0_2),.dout(w_dff_B_Vf48OteZ5_2),.clk(gclk));
	jdff dff_B_BjWISscr8_2(.din(w_dff_B_Vf48OteZ5_2),.dout(w_dff_B_BjWISscr8_2),.clk(gclk));
	jdff dff_B_vj2wDx672_2(.din(w_dff_B_BjWISscr8_2),.dout(w_dff_B_vj2wDx672_2),.clk(gclk));
	jdff dff_B_wDPUzVfv3_2(.din(w_dff_B_vj2wDx672_2),.dout(w_dff_B_wDPUzVfv3_2),.clk(gclk));
	jdff dff_B_qjQmfUAx7_2(.din(w_dff_B_wDPUzVfv3_2),.dout(w_dff_B_qjQmfUAx7_2),.clk(gclk));
	jdff dff_B_Azfpz1S68_2(.din(w_dff_B_qjQmfUAx7_2),.dout(w_dff_B_Azfpz1S68_2),.clk(gclk));
	jdff dff_B_hcgaCqcM6_2(.din(w_dff_B_Azfpz1S68_2),.dout(w_dff_B_hcgaCqcM6_2),.clk(gclk));
	jdff dff_B_3UeVQoDM4_2(.din(w_dff_B_hcgaCqcM6_2),.dout(w_dff_B_3UeVQoDM4_2),.clk(gclk));
	jdff dff_B_Q4AQdZVD8_2(.din(w_dff_B_3UeVQoDM4_2),.dout(w_dff_B_Q4AQdZVD8_2),.clk(gclk));
	jdff dff_B_mHlD39nI3_2(.din(w_dff_B_Q4AQdZVD8_2),.dout(w_dff_B_mHlD39nI3_2),.clk(gclk));
	jdff dff_B_iEZyaL1c4_2(.din(w_dff_B_mHlD39nI3_2),.dout(w_dff_B_iEZyaL1c4_2),.clk(gclk));
	jdff dff_B_XbZFELvh9_2(.din(w_dff_B_iEZyaL1c4_2),.dout(w_dff_B_XbZFELvh9_2),.clk(gclk));
	jdff dff_B_mPS8lHRW8_2(.din(w_dff_B_XbZFELvh9_2),.dout(w_dff_B_mPS8lHRW8_2),.clk(gclk));
	jdff dff_B_HcZRw80p2_2(.din(w_dff_B_mPS8lHRW8_2),.dout(w_dff_B_HcZRw80p2_2),.clk(gclk));
	jdff dff_B_OmqXnA2Q9_2(.din(w_dff_B_HcZRw80p2_2),.dout(w_dff_B_OmqXnA2Q9_2),.clk(gclk));
	jdff dff_B_DYxtLUtm1_2(.din(w_dff_B_OmqXnA2Q9_2),.dout(w_dff_B_DYxtLUtm1_2),.clk(gclk));
	jdff dff_B_D1Vf5IR67_2(.din(w_dff_B_DYxtLUtm1_2),.dout(w_dff_B_D1Vf5IR67_2),.clk(gclk));
	jdff dff_B_YaBbk4dy6_2(.din(w_dff_B_D1Vf5IR67_2),.dout(w_dff_B_YaBbk4dy6_2),.clk(gclk));
	jdff dff_B_skCxo6cn5_2(.din(w_dff_B_YaBbk4dy6_2),.dout(w_dff_B_skCxo6cn5_2),.clk(gclk));
	jdff dff_B_oLai4ogo7_2(.din(w_dff_B_skCxo6cn5_2),.dout(w_dff_B_oLai4ogo7_2),.clk(gclk));
	jdff dff_B_oCqZeK9A2_2(.din(w_dff_B_oLai4ogo7_2),.dout(w_dff_B_oCqZeK9A2_2),.clk(gclk));
	jdff dff_B_t8rZiQpd3_2(.din(w_dff_B_oCqZeK9A2_2),.dout(w_dff_B_t8rZiQpd3_2),.clk(gclk));
	jdff dff_B_g8A50B8m5_2(.din(w_dff_B_t8rZiQpd3_2),.dout(w_dff_B_g8A50B8m5_2),.clk(gclk));
	jdff dff_B_dWR5q1Fo9_2(.din(w_dff_B_g8A50B8m5_2),.dout(w_dff_B_dWR5q1Fo9_2),.clk(gclk));
	jdff dff_B_pHDyiLtD2_2(.din(w_dff_B_dWR5q1Fo9_2),.dout(w_dff_B_pHDyiLtD2_2),.clk(gclk));
	jdff dff_B_NMNpQCzb9_2(.din(w_dff_B_pHDyiLtD2_2),.dout(w_dff_B_NMNpQCzb9_2),.clk(gclk));
	jdff dff_B_l40YQyJq7_2(.din(w_dff_B_NMNpQCzb9_2),.dout(w_dff_B_l40YQyJq7_2),.clk(gclk));
	jdff dff_B_BT3ftis21_2(.din(w_dff_B_l40YQyJq7_2),.dout(w_dff_B_BT3ftis21_2),.clk(gclk));
	jdff dff_B_piv4UxAW4_2(.din(w_dff_B_BT3ftis21_2),.dout(w_dff_B_piv4UxAW4_2),.clk(gclk));
	jdff dff_B_YaZOEOUM2_2(.din(w_dff_B_piv4UxAW4_2),.dout(w_dff_B_YaZOEOUM2_2),.clk(gclk));
	jdff dff_B_7yHGmmnQ4_2(.din(w_dff_B_YaZOEOUM2_2),.dout(w_dff_B_7yHGmmnQ4_2),.clk(gclk));
	jdff dff_B_Eqw1Eoid2_2(.din(w_dff_B_7yHGmmnQ4_2),.dout(w_dff_B_Eqw1Eoid2_2),.clk(gclk));
	jdff dff_B_gxMfK08z8_2(.din(w_dff_B_Eqw1Eoid2_2),.dout(w_dff_B_gxMfK08z8_2),.clk(gclk));
	jdff dff_B_wrNl0mPO3_2(.din(w_dff_B_gxMfK08z8_2),.dout(w_dff_B_wrNl0mPO3_2),.clk(gclk));
	jdff dff_B_5wg4ZqNC2_2(.din(w_dff_B_wrNl0mPO3_2),.dout(w_dff_B_5wg4ZqNC2_2),.clk(gclk));
	jdff dff_B_QZ2jD26B7_2(.din(w_dff_B_5wg4ZqNC2_2),.dout(w_dff_B_QZ2jD26B7_2),.clk(gclk));
	jdff dff_B_mgLcBMrq0_2(.din(w_dff_B_QZ2jD26B7_2),.dout(w_dff_B_mgLcBMrq0_2),.clk(gclk));
	jdff dff_B_oqKx0yJG3_2(.din(w_dff_B_mgLcBMrq0_2),.dout(w_dff_B_oqKx0yJG3_2),.clk(gclk));
	jdff dff_B_a5YMA9Xd5_2(.din(w_dff_B_oqKx0yJG3_2),.dout(w_dff_B_a5YMA9Xd5_2),.clk(gclk));
	jdff dff_B_nj95YJpD7_2(.din(w_dff_B_a5YMA9Xd5_2),.dout(w_dff_B_nj95YJpD7_2),.clk(gclk));
	jdff dff_B_ic5w4RTK2_2(.din(w_dff_B_nj95YJpD7_2),.dout(w_dff_B_ic5w4RTK2_2),.clk(gclk));
	jdff dff_B_dXIi2qk55_2(.din(w_dff_B_ic5w4RTK2_2),.dout(w_dff_B_dXIi2qk55_2),.clk(gclk));
	jdff dff_B_esowjK944_2(.din(w_dff_B_dXIi2qk55_2),.dout(w_dff_B_esowjK944_2),.clk(gclk));
	jdff dff_B_lV2zAyrv2_2(.din(w_dff_B_esowjK944_2),.dout(w_dff_B_lV2zAyrv2_2),.clk(gclk));
	jdff dff_B_wdHBHGlt9_2(.din(w_dff_B_lV2zAyrv2_2),.dout(w_dff_B_wdHBHGlt9_2),.clk(gclk));
	jdff dff_B_12H6lgze3_2(.din(w_dff_B_wdHBHGlt9_2),.dout(w_dff_B_12H6lgze3_2),.clk(gclk));
	jdff dff_B_cfAJE7kt4_2(.din(w_dff_B_12H6lgze3_2),.dout(w_dff_B_cfAJE7kt4_2),.clk(gclk));
	jdff dff_B_6uoYTNQ31_2(.din(w_dff_B_cfAJE7kt4_2),.dout(w_dff_B_6uoYTNQ31_2),.clk(gclk));
	jdff dff_B_T5nNgsKl4_2(.din(w_dff_B_6uoYTNQ31_2),.dout(w_dff_B_T5nNgsKl4_2),.clk(gclk));
	jdff dff_B_2an2B9t30_2(.din(w_dff_B_T5nNgsKl4_2),.dout(w_dff_B_2an2B9t30_2),.clk(gclk));
	jdff dff_B_hHzmKy4M6_2(.din(w_dff_B_2an2B9t30_2),.dout(w_dff_B_hHzmKy4M6_2),.clk(gclk));
	jdff dff_B_cRoA1fFK0_2(.din(w_dff_B_hHzmKy4M6_2),.dout(w_dff_B_cRoA1fFK0_2),.clk(gclk));
	jdff dff_B_hTwIDE0m7_2(.din(w_dff_B_cRoA1fFK0_2),.dout(w_dff_B_hTwIDE0m7_2),.clk(gclk));
	jdff dff_B_Guqptcbx6_2(.din(w_dff_B_hTwIDE0m7_2),.dout(w_dff_B_Guqptcbx6_2),.clk(gclk));
	jdff dff_B_VCH2f1942_2(.din(w_dff_B_Guqptcbx6_2),.dout(w_dff_B_VCH2f1942_2),.clk(gclk));
	jdff dff_B_IANTEjUk4_2(.din(w_dff_B_VCH2f1942_2),.dout(w_dff_B_IANTEjUk4_2),.clk(gclk));
	jdff dff_B_jUUEGEbz3_2(.din(w_dff_B_IANTEjUk4_2),.dout(w_dff_B_jUUEGEbz3_2),.clk(gclk));
	jdff dff_B_5ILDH56V2_2(.din(w_dff_B_jUUEGEbz3_2),.dout(w_dff_B_5ILDH56V2_2),.clk(gclk));
	jdff dff_B_fSqyH1h07_2(.din(w_dff_B_5ILDH56V2_2),.dout(w_dff_B_fSqyH1h07_2),.clk(gclk));
	jdff dff_B_66DMoCJC3_2(.din(w_dff_B_fSqyH1h07_2),.dout(w_dff_B_66DMoCJC3_2),.clk(gclk));
	jdff dff_B_0HtgoPMs5_2(.din(w_dff_B_66DMoCJC3_2),.dout(w_dff_B_0HtgoPMs5_2),.clk(gclk));
	jdff dff_B_Vtxq4e4r5_2(.din(w_dff_B_0HtgoPMs5_2),.dout(w_dff_B_Vtxq4e4r5_2),.clk(gclk));
	jdff dff_B_xGEbT75K7_2(.din(w_dff_B_Vtxq4e4r5_2),.dout(w_dff_B_xGEbT75K7_2),.clk(gclk));
	jdff dff_B_vH0bzWc02_2(.din(w_dff_B_xGEbT75K7_2),.dout(w_dff_B_vH0bzWc02_2),.clk(gclk));
	jdff dff_B_w7n94gEX8_2(.din(w_dff_B_vH0bzWc02_2),.dout(w_dff_B_w7n94gEX8_2),.clk(gclk));
	jdff dff_B_YFN78Xne8_2(.din(w_dff_B_w7n94gEX8_2),.dout(w_dff_B_YFN78Xne8_2),.clk(gclk));
	jdff dff_B_G3xf6Y8X5_2(.din(w_dff_B_YFN78Xne8_2),.dout(w_dff_B_G3xf6Y8X5_2),.clk(gclk));
	jdff dff_B_WeiAwsGA5_2(.din(w_dff_B_G3xf6Y8X5_2),.dout(w_dff_B_WeiAwsGA5_2),.clk(gclk));
	jdff dff_B_AJtHLJFq3_2(.din(w_dff_B_WeiAwsGA5_2),.dout(w_dff_B_AJtHLJFq3_2),.clk(gclk));
	jdff dff_B_sgIIXb0q8_2(.din(w_dff_B_AJtHLJFq3_2),.dout(w_dff_B_sgIIXb0q8_2),.clk(gclk));
	jdff dff_B_rsT1Gty44_2(.din(w_dff_B_sgIIXb0q8_2),.dout(w_dff_B_rsT1Gty44_2),.clk(gclk));
	jdff dff_B_trnnJA641_2(.din(w_dff_B_rsT1Gty44_2),.dout(w_dff_B_trnnJA641_2),.clk(gclk));
	jdff dff_B_uHnlTEZm1_2(.din(w_dff_B_trnnJA641_2),.dout(w_dff_B_uHnlTEZm1_2),.clk(gclk));
	jdff dff_B_uipMsoLk5_2(.din(w_dff_B_uHnlTEZm1_2),.dout(w_dff_B_uipMsoLk5_2),.clk(gclk));
	jdff dff_B_cdI1whfO0_2(.din(w_dff_B_uipMsoLk5_2),.dout(w_dff_B_cdI1whfO0_2),.clk(gclk));
	jdff dff_B_68oxuLKL0_2(.din(w_dff_B_cdI1whfO0_2),.dout(w_dff_B_68oxuLKL0_2),.clk(gclk));
	jdff dff_B_hdmnGyEV0_2(.din(w_dff_B_68oxuLKL0_2),.dout(w_dff_B_hdmnGyEV0_2),.clk(gclk));
	jdff dff_B_6F56Vpri7_2(.din(w_dff_B_hdmnGyEV0_2),.dout(w_dff_B_6F56Vpri7_2),.clk(gclk));
	jdff dff_B_rKPkvx055_2(.din(w_dff_B_6F56Vpri7_2),.dout(w_dff_B_rKPkvx055_2),.clk(gclk));
	jdff dff_A_L0OSZQeM0_0(.dout(w_n4093_3[0]),.din(w_dff_A_L0OSZQeM0_0),.clk(gclk));
	jdff dff_A_EzVOOBro3_0(.dout(w_dff_A_L0OSZQeM0_0),.din(w_dff_A_EzVOOBro3_0),.clk(gclk));
	jdff dff_A_S76g9eo65_0(.dout(w_dff_A_EzVOOBro3_0),.din(w_dff_A_S76g9eo65_0),.clk(gclk));
	jdff dff_A_ym8OQgjx3_0(.dout(w_dff_A_S76g9eo65_0),.din(w_dff_A_ym8OQgjx3_0),.clk(gclk));
	jdff dff_A_SAnq582t7_0(.dout(w_dff_A_ym8OQgjx3_0),.din(w_dff_A_SAnq582t7_0),.clk(gclk));
	jdff dff_A_3DhaB3OS0_2(.dout(w_n4093_3[2]),.din(w_dff_A_3DhaB3OS0_2),.clk(gclk));
	jdff dff_A_kWqmFeRs7_2(.dout(w_dff_A_3DhaB3OS0_2),.din(w_dff_A_kWqmFeRs7_2),.clk(gclk));
	jdff dff_A_srR7HyzS7_2(.dout(w_dff_A_kWqmFeRs7_2),.din(w_dff_A_srR7HyzS7_2),.clk(gclk));
	jdff dff_A_OBpDxHwd5_2(.dout(w_dff_A_srR7HyzS7_2),.din(w_dff_A_OBpDxHwd5_2),.clk(gclk));
	jdff dff_A_Dhx2dUCK6_2(.dout(w_dff_A_OBpDxHwd5_2),.din(w_dff_A_Dhx2dUCK6_2),.clk(gclk));
	jdff dff_A_SBZ1jIyq3_2(.dout(w_dff_A_Dhx2dUCK6_2),.din(w_dff_A_SBZ1jIyq3_2),.clk(gclk));
	jdff dff_A_reKGcl5w9_2(.dout(w_dff_A_SBZ1jIyq3_2),.din(w_dff_A_reKGcl5w9_2),.clk(gclk));
	jdff dff_A_3CAYALH19_2(.dout(w_dff_A_reKGcl5w9_2),.din(w_dff_A_3CAYALH19_2),.clk(gclk));
	jdff dff_A_3WCqoWx00_2(.dout(w_dff_A_3CAYALH19_2),.din(w_dff_A_3WCqoWx00_2),.clk(gclk));
	jdff dff_A_WClAtgeI0_2(.dout(w_dff_A_3WCqoWx00_2),.din(w_dff_A_WClAtgeI0_2),.clk(gclk));
	jdff dff_A_41HVUZn98_2(.dout(w_dff_A_WClAtgeI0_2),.din(w_dff_A_41HVUZn98_2),.clk(gclk));
	jdff dff_A_mLXrjMgu6_2(.dout(w_dff_A_41HVUZn98_2),.din(w_dff_A_mLXrjMgu6_2),.clk(gclk));
	jdff dff_A_RYsBOHbI4_2(.dout(w_dff_A_mLXrjMgu6_2),.din(w_dff_A_RYsBOHbI4_2),.clk(gclk));
	jdff dff_A_dLlsKCHL4_2(.dout(w_dff_A_RYsBOHbI4_2),.din(w_dff_A_dLlsKCHL4_2),.clk(gclk));
	jdff dff_A_NX8QHL285_2(.dout(w_dff_A_dLlsKCHL4_2),.din(w_dff_A_NX8QHL285_2),.clk(gclk));
	jdff dff_A_xRtQnvNO0_2(.dout(w_dff_A_NX8QHL285_2),.din(w_dff_A_xRtQnvNO0_2),.clk(gclk));
	jdff dff_A_0QscNQfu9_2(.dout(w_dff_A_xRtQnvNO0_2),.din(w_dff_A_0QscNQfu9_2),.clk(gclk));
	jdff dff_A_5TgjVQ6D2_2(.dout(w_dff_A_0QscNQfu9_2),.din(w_dff_A_5TgjVQ6D2_2),.clk(gclk));
	jdff dff_A_wdCcFoKc2_2(.dout(w_dff_A_5TgjVQ6D2_2),.din(w_dff_A_wdCcFoKc2_2),.clk(gclk));
	jdff dff_A_7nV63SFc6_2(.dout(w_dff_A_wdCcFoKc2_2),.din(w_dff_A_7nV63SFc6_2),.clk(gclk));
	jdff dff_A_F9b0VBf80_2(.dout(w_dff_A_7nV63SFc6_2),.din(w_dff_A_F9b0VBf80_2),.clk(gclk));
	jdff dff_A_D1Do9hXi2_2(.dout(w_dff_A_F9b0VBf80_2),.din(w_dff_A_D1Do9hXi2_2),.clk(gclk));
	jdff dff_A_Wr6rtGAY9_2(.dout(w_dff_A_D1Do9hXi2_2),.din(w_dff_A_Wr6rtGAY9_2),.clk(gclk));
	jdff dff_A_51A04pXA4_2(.dout(w_dff_A_Wr6rtGAY9_2),.din(w_dff_A_51A04pXA4_2),.clk(gclk));
	jdff dff_A_Hfc4Msnq2_2(.dout(w_dff_A_51A04pXA4_2),.din(w_dff_A_Hfc4Msnq2_2),.clk(gclk));
	jdff dff_A_WbIvKlhB1_2(.dout(w_dff_A_Hfc4Msnq2_2),.din(w_dff_A_WbIvKlhB1_2),.clk(gclk));
	jdff dff_A_KiShnFwz1_2(.dout(w_dff_A_WbIvKlhB1_2),.din(w_dff_A_KiShnFwz1_2),.clk(gclk));
	jdff dff_A_ON4G458g6_2(.dout(w_dff_A_KiShnFwz1_2),.din(w_dff_A_ON4G458g6_2),.clk(gclk));
	jdff dff_A_yEunRhnk7_2(.dout(w_dff_A_ON4G458g6_2),.din(w_dff_A_yEunRhnk7_2),.clk(gclk));
	jdff dff_A_S1qxlL0P9_2(.dout(w_dff_A_yEunRhnk7_2),.din(w_dff_A_S1qxlL0P9_2),.clk(gclk));
	jdff dff_A_SdjizuFJ5_2(.dout(w_dff_A_S1qxlL0P9_2),.din(w_dff_A_SdjizuFJ5_2),.clk(gclk));
	jdff dff_A_DqhU2h8p0_2(.dout(w_dff_A_SdjizuFJ5_2),.din(w_dff_A_DqhU2h8p0_2),.clk(gclk));
	jdff dff_A_6KqLycjQ3_2(.dout(w_dff_A_DqhU2h8p0_2),.din(w_dff_A_6KqLycjQ3_2),.clk(gclk));
	jdff dff_A_s366T35O6_2(.dout(w_dff_A_6KqLycjQ3_2),.din(w_dff_A_s366T35O6_2),.clk(gclk));
	jdff dff_A_NpGDyYQY8_2(.dout(w_dff_A_s366T35O6_2),.din(w_dff_A_NpGDyYQY8_2),.clk(gclk));
	jdff dff_A_bbaWNdBH9_2(.dout(w_dff_A_NpGDyYQY8_2),.din(w_dff_A_bbaWNdBH9_2),.clk(gclk));
	jdff dff_A_1rxV4xZO2_2(.dout(w_dff_A_bbaWNdBH9_2),.din(w_dff_A_1rxV4xZO2_2),.clk(gclk));
	jdff dff_A_IOp0rUXs9_2(.dout(w_dff_A_1rxV4xZO2_2),.din(w_dff_A_IOp0rUXs9_2),.clk(gclk));
	jdff dff_A_YwlGR1es5_2(.dout(w_dff_A_IOp0rUXs9_2),.din(w_dff_A_YwlGR1es5_2),.clk(gclk));
	jdff dff_A_6OZN7T3U7_2(.dout(w_dff_A_YwlGR1es5_2),.din(w_dff_A_6OZN7T3U7_2),.clk(gclk));
	jdff dff_A_qPkaeIQa7_2(.dout(w_dff_A_6OZN7T3U7_2),.din(w_dff_A_qPkaeIQa7_2),.clk(gclk));
	jdff dff_A_TbPrP1sW3_2(.dout(w_dff_A_qPkaeIQa7_2),.din(w_dff_A_TbPrP1sW3_2),.clk(gclk));
	jdff dff_A_IxICBTvT9_2(.dout(w_dff_A_TbPrP1sW3_2),.din(w_dff_A_IxICBTvT9_2),.clk(gclk));
	jdff dff_A_9fZQPXhh0_0(.dout(w_n5476_0[0]),.din(w_dff_A_9fZQPXhh0_0),.clk(gclk));
	jdff dff_A_jveqLtSa7_1(.dout(w_n5400_0[1]),.din(w_dff_A_jveqLtSa7_1),.clk(gclk));
	jdff dff_A_0wlIeazr9_0(.dout(w_n5354_0[0]),.din(w_dff_A_0wlIeazr9_0),.clk(gclk));
	jdff dff_A_xMHNluYy5_0(.dout(w_n5351_0[0]),.din(w_dff_A_xMHNluYy5_0),.clk(gclk));
	jdff dff_A_ghwMUcgR8_0(.dout(w_dff_A_xMHNluYy5_0),.din(w_dff_A_ghwMUcgR8_0),.clk(gclk));
	jdff dff_A_ruo15GOT6_0(.dout(w_n5248_0[0]),.din(w_dff_A_ruo15GOT6_0),.clk(gclk));
	jdff dff_A_bxvqYTYx4_0(.dout(w_n5210_0[0]),.din(w_dff_A_bxvqYTYx4_0),.clk(gclk));
	jdff dff_A_zf31BzpE2_0(.dout(w_n5164_0[0]),.din(w_dff_A_zf31BzpE2_0),.clk(gclk));
	jdff dff_A_A2xONnuD7_0(.dout(w_n5113_0[0]),.din(w_dff_A_A2xONnuD7_0),.clk(gclk));
	jdff dff_A_vrPoZQgf4_0(.dout(w_n5058_0[0]),.din(w_dff_A_vrPoZQgf4_0),.clk(gclk));
	jdff dff_A_AlQfCFvp1_0(.dout(w_n5004_0[0]),.din(w_dff_A_AlQfCFvp1_0),.clk(gclk));
	jdff dff_A_c4lpFFo59_0(.dout(w_n4934_0[0]),.din(w_dff_A_c4lpFFo59_0),.clk(gclk));
	jdff dff_A_qqLHRbws4_0(.dout(w_n4868_0[0]),.din(w_dff_A_qqLHRbws4_0),.clk(gclk));
	jdff dff_A_ws4tWc4i8_0(.dout(w_n4786_0[0]),.din(w_dff_A_ws4tWc4i8_0),.clk(gclk));
	jdff dff_A_CepdS1678_0(.dout(w_n4713_0[0]),.din(w_dff_A_CepdS1678_0),.clk(gclk));
	jdff dff_A_kXRcecfy2_0(.dout(w_n4629_0[0]),.din(w_dff_A_kXRcecfy2_0),.clk(gclk));
	jdff dff_A_rxmmLz2D9_0(.dout(w_n4543_0[0]),.din(w_dff_A_rxmmLz2D9_0),.clk(gclk));
	jdff dff_A_y8pPL52h4_0(.dout(w_n4364_0[0]),.din(w_dff_A_y8pPL52h4_0),.clk(gclk));
	jdff dff_A_nhCEAzVC8_0(.dout(w_n4361_0[0]),.din(w_dff_A_nhCEAzVC8_0),.clk(gclk));
	jdff dff_A_4X71YBkO2_0(.dout(w_sin0_0[0]),.din(w_dff_A_4X71YBkO2_0),.clk(gclk));
	jdff dff_A_gvfmGipg2_0(.dout(w_dff_A_4X71YBkO2_0),.din(w_dff_A_gvfmGipg2_0),.clk(gclk));
	jdff dff_A_JzuBWyFX9_1(.dout(w_n5440_0[1]),.din(w_dff_A_JzuBWyFX9_1),.clk(gclk));
	jdff dff_A_RcIzSiyI2_2(.dout(w_dff_A_e7OvVlbE3_0),.din(w_dff_A_RcIzSiyI2_2),.clk(gclk));
	jdff dff_A_e7OvVlbE3_0(.dout(w_dff_A_x8u3rqMD0_0),.din(w_dff_A_e7OvVlbE3_0),.clk(gclk));
	jdff dff_A_x8u3rqMD0_0(.dout(w_dff_A_P2fU1v5w1_0),.din(w_dff_A_x8u3rqMD0_0),.clk(gclk));
	jdff dff_A_P2fU1v5w1_0(.dout(w_dff_A_3xwklP8D3_0),.din(w_dff_A_P2fU1v5w1_0),.clk(gclk));
	jdff dff_A_3xwklP8D3_0(.dout(w_dff_A_1GEFQsI24_0),.din(w_dff_A_3xwklP8D3_0),.clk(gclk));
	jdff dff_A_1GEFQsI24_0(.dout(w_dff_A_e2sVsjtH3_0),.din(w_dff_A_1GEFQsI24_0),.clk(gclk));
	jdff dff_A_e2sVsjtH3_0(.dout(w_dff_A_O2BO2SuL6_0),.din(w_dff_A_e2sVsjtH3_0),.clk(gclk));
	jdff dff_A_O2BO2SuL6_0(.dout(w_dff_A_ZJQET9YO9_0),.din(w_dff_A_O2BO2SuL6_0),.clk(gclk));
	jdff dff_A_ZJQET9YO9_0(.dout(w_dff_A_mc8ahk2U2_0),.din(w_dff_A_ZJQET9YO9_0),.clk(gclk));
	jdff dff_A_mc8ahk2U2_0(.dout(w_dff_A_49KuOZhG8_0),.din(w_dff_A_mc8ahk2U2_0),.clk(gclk));
	jdff dff_A_49KuOZhG8_0(.dout(w_dff_A_GCpml2Rb2_0),.din(w_dff_A_49KuOZhG8_0),.clk(gclk));
	jdff dff_A_GCpml2Rb2_0(.dout(w_dff_A_9FdPHtPY2_0),.din(w_dff_A_GCpml2Rb2_0),.clk(gclk));
	jdff dff_A_9FdPHtPY2_0(.dout(w_dff_A_mSsyGlbX9_0),.din(w_dff_A_9FdPHtPY2_0),.clk(gclk));
	jdff dff_A_mSsyGlbX9_0(.dout(w_dff_A_HLhGPyqR3_0),.din(w_dff_A_mSsyGlbX9_0),.clk(gclk));
	jdff dff_A_HLhGPyqR3_0(.dout(w_dff_A_1O6kJoWc7_0),.din(w_dff_A_HLhGPyqR3_0),.clk(gclk));
	jdff dff_A_1O6kJoWc7_0(.dout(w_dff_A_w2WYrEui2_0),.din(w_dff_A_1O6kJoWc7_0),.clk(gclk));
	jdff dff_A_w2WYrEui2_0(.dout(w_dff_A_lAXy6uRz5_0),.din(w_dff_A_w2WYrEui2_0),.clk(gclk));
	jdff dff_A_lAXy6uRz5_0(.dout(w_dff_A_AftDaAqX0_0),.din(w_dff_A_lAXy6uRz5_0),.clk(gclk));
	jdff dff_A_AftDaAqX0_0(.dout(w_dff_A_7Fzu6oUl4_0),.din(w_dff_A_AftDaAqX0_0),.clk(gclk));
	jdff dff_A_7Fzu6oUl4_0(.dout(w_dff_A_zlRC7fJ27_0),.din(w_dff_A_7Fzu6oUl4_0),.clk(gclk));
	jdff dff_A_zlRC7fJ27_0(.dout(w_dff_A_eAGqGZV06_0),.din(w_dff_A_zlRC7fJ27_0),.clk(gclk));
	jdff dff_A_eAGqGZV06_0(.dout(w_dff_A_VdNX6NyX9_0),.din(w_dff_A_eAGqGZV06_0),.clk(gclk));
	jdff dff_A_VdNX6NyX9_0(.dout(w_dff_A_MT890JFd0_0),.din(w_dff_A_VdNX6NyX9_0),.clk(gclk));
	jdff dff_A_MT890JFd0_0(.dout(w_dff_A_11Rao2mE8_0),.din(w_dff_A_MT890JFd0_0),.clk(gclk));
	jdff dff_A_11Rao2mE8_0(.dout(w_dff_A_Sb9gVHhB4_0),.din(w_dff_A_11Rao2mE8_0),.clk(gclk));
	jdff dff_A_Sb9gVHhB4_0(.dout(w_dff_A_hvUl05Pf1_0),.din(w_dff_A_Sb9gVHhB4_0),.clk(gclk));
	jdff dff_A_hvUl05Pf1_0(.dout(w_dff_A_9OZLVE5l3_0),.din(w_dff_A_hvUl05Pf1_0),.clk(gclk));
	jdff dff_A_9OZLVE5l3_0(.dout(w_dff_A_jtnIGmFe4_0),.din(w_dff_A_9OZLVE5l3_0),.clk(gclk));
	jdff dff_A_jtnIGmFe4_0(.dout(w_dff_A_zUG6Bm9Q7_0),.din(w_dff_A_jtnIGmFe4_0),.clk(gclk));
	jdff dff_A_zUG6Bm9Q7_0(.dout(w_dff_A_XxcD9WVy3_0),.din(w_dff_A_zUG6Bm9Q7_0),.clk(gclk));
	jdff dff_A_XxcD9WVy3_0(.dout(w_dff_A_RyqwCY9u2_0),.din(w_dff_A_XxcD9WVy3_0),.clk(gclk));
	jdff dff_A_RyqwCY9u2_0(.dout(w_dff_A_FxOhrNQK7_0),.din(w_dff_A_RyqwCY9u2_0),.clk(gclk));
	jdff dff_A_FxOhrNQK7_0(.dout(w_dff_A_Qn7JLtK60_0),.din(w_dff_A_FxOhrNQK7_0),.clk(gclk));
	jdff dff_A_Qn7JLtK60_0(.dout(w_dff_A_oSQJc16z0_0),.din(w_dff_A_Qn7JLtK60_0),.clk(gclk));
	jdff dff_A_oSQJc16z0_0(.dout(w_dff_A_FKebBWTn9_0),.din(w_dff_A_oSQJc16z0_0),.clk(gclk));
	jdff dff_A_FKebBWTn9_0(.dout(w_dff_A_Yzu5N13E9_0),.din(w_dff_A_FKebBWTn9_0),.clk(gclk));
	jdff dff_A_Yzu5N13E9_0(.dout(w_dff_A_ckZ4nhGs3_0),.din(w_dff_A_Yzu5N13E9_0),.clk(gclk));
	jdff dff_A_ckZ4nhGs3_0(.dout(w_dff_A_rRcHmzzS2_0),.din(w_dff_A_ckZ4nhGs3_0),.clk(gclk));
	jdff dff_A_rRcHmzzS2_0(.dout(w_dff_A_SFMSlVxD8_0),.din(w_dff_A_rRcHmzzS2_0),.clk(gclk));
	jdff dff_A_SFMSlVxD8_0(.dout(w_dff_A_cUSIBKFX0_0),.din(w_dff_A_SFMSlVxD8_0),.clk(gclk));
	jdff dff_A_cUSIBKFX0_0(.dout(w_dff_A_zCNYNeL25_0),.din(w_dff_A_cUSIBKFX0_0),.clk(gclk));
	jdff dff_A_zCNYNeL25_0(.dout(w_dff_A_d8buYoeM8_0),.din(w_dff_A_zCNYNeL25_0),.clk(gclk));
	jdff dff_A_d8buYoeM8_0(.dout(w_dff_A_LSNUlBTH4_0),.din(w_dff_A_d8buYoeM8_0),.clk(gclk));
	jdff dff_A_LSNUlBTH4_0(.dout(w_dff_A_UEaQSzRB1_0),.din(w_dff_A_LSNUlBTH4_0),.clk(gclk));
	jdff dff_A_UEaQSzRB1_0(.dout(w_dff_A_lqrq3xOV2_0),.din(w_dff_A_UEaQSzRB1_0),.clk(gclk));
	jdff dff_A_lqrq3xOV2_0(.dout(sin0),.din(w_dff_A_lqrq3xOV2_0),.clk(gclk));
	jdff dff_A_aLvUiHOn0_2(.dout(w_dff_A_36xkr33S4_0),.din(w_dff_A_aLvUiHOn0_2),.clk(gclk));
	jdff dff_A_36xkr33S4_0(.dout(w_dff_A_o55eBeBQ4_0),.din(w_dff_A_36xkr33S4_0),.clk(gclk));
	jdff dff_A_o55eBeBQ4_0(.dout(w_dff_A_I44ZRdTT2_0),.din(w_dff_A_o55eBeBQ4_0),.clk(gclk));
	jdff dff_A_I44ZRdTT2_0(.dout(w_dff_A_BBmXfpbl4_0),.din(w_dff_A_I44ZRdTT2_0),.clk(gclk));
	jdff dff_A_BBmXfpbl4_0(.dout(w_dff_A_0ub60h0U0_0),.din(w_dff_A_BBmXfpbl4_0),.clk(gclk));
	jdff dff_A_0ub60h0U0_0(.dout(w_dff_A_MZFFVovT9_0),.din(w_dff_A_0ub60h0U0_0),.clk(gclk));
	jdff dff_A_MZFFVovT9_0(.dout(w_dff_A_IHLM9I733_0),.din(w_dff_A_MZFFVovT9_0),.clk(gclk));
	jdff dff_A_IHLM9I733_0(.dout(w_dff_A_KLHWcDfI4_0),.din(w_dff_A_IHLM9I733_0),.clk(gclk));
	jdff dff_A_KLHWcDfI4_0(.dout(w_dff_A_Hd0B8Jnf1_0),.din(w_dff_A_KLHWcDfI4_0),.clk(gclk));
	jdff dff_A_Hd0B8Jnf1_0(.dout(w_dff_A_2vEbmlFC5_0),.din(w_dff_A_Hd0B8Jnf1_0),.clk(gclk));
	jdff dff_A_2vEbmlFC5_0(.dout(w_dff_A_hSQHa8jX8_0),.din(w_dff_A_2vEbmlFC5_0),.clk(gclk));
	jdff dff_A_hSQHa8jX8_0(.dout(w_dff_A_3RiqyP598_0),.din(w_dff_A_hSQHa8jX8_0),.clk(gclk));
	jdff dff_A_3RiqyP598_0(.dout(w_dff_A_m7toEkNz9_0),.din(w_dff_A_3RiqyP598_0),.clk(gclk));
	jdff dff_A_m7toEkNz9_0(.dout(w_dff_A_g8OhgRoj8_0),.din(w_dff_A_m7toEkNz9_0),.clk(gclk));
	jdff dff_A_g8OhgRoj8_0(.dout(w_dff_A_nigqpQkF5_0),.din(w_dff_A_g8OhgRoj8_0),.clk(gclk));
	jdff dff_A_nigqpQkF5_0(.dout(w_dff_A_A1jV4zv96_0),.din(w_dff_A_nigqpQkF5_0),.clk(gclk));
	jdff dff_A_A1jV4zv96_0(.dout(w_dff_A_2I9T2eCA4_0),.din(w_dff_A_A1jV4zv96_0),.clk(gclk));
	jdff dff_A_2I9T2eCA4_0(.dout(w_dff_A_KicReXWK1_0),.din(w_dff_A_2I9T2eCA4_0),.clk(gclk));
	jdff dff_A_KicReXWK1_0(.dout(w_dff_A_3XaUSEr87_0),.din(w_dff_A_KicReXWK1_0),.clk(gclk));
	jdff dff_A_3XaUSEr87_0(.dout(w_dff_A_NkYjzl1y2_0),.din(w_dff_A_3XaUSEr87_0),.clk(gclk));
	jdff dff_A_NkYjzl1y2_0(.dout(w_dff_A_KnkghA6m8_0),.din(w_dff_A_NkYjzl1y2_0),.clk(gclk));
	jdff dff_A_KnkghA6m8_0(.dout(w_dff_A_fIQ9wPgT5_0),.din(w_dff_A_KnkghA6m8_0),.clk(gclk));
	jdff dff_A_fIQ9wPgT5_0(.dout(w_dff_A_sYPqM0Ne0_0),.din(w_dff_A_fIQ9wPgT5_0),.clk(gclk));
	jdff dff_A_sYPqM0Ne0_0(.dout(w_dff_A_1dBbuaDt8_0),.din(w_dff_A_sYPqM0Ne0_0),.clk(gclk));
	jdff dff_A_1dBbuaDt8_0(.dout(w_dff_A_ddmVdl7d3_0),.din(w_dff_A_1dBbuaDt8_0),.clk(gclk));
	jdff dff_A_ddmVdl7d3_0(.dout(w_dff_A_MltskOaQ4_0),.din(w_dff_A_ddmVdl7d3_0),.clk(gclk));
	jdff dff_A_MltskOaQ4_0(.dout(w_dff_A_dLbVsA956_0),.din(w_dff_A_MltskOaQ4_0),.clk(gclk));
	jdff dff_A_dLbVsA956_0(.dout(w_dff_A_byJOwl0s0_0),.din(w_dff_A_dLbVsA956_0),.clk(gclk));
	jdff dff_A_byJOwl0s0_0(.dout(w_dff_A_KwEVwRUv5_0),.din(w_dff_A_byJOwl0s0_0),.clk(gclk));
	jdff dff_A_KwEVwRUv5_0(.dout(w_dff_A_QujEOu9A6_0),.din(w_dff_A_KwEVwRUv5_0),.clk(gclk));
	jdff dff_A_QujEOu9A6_0(.dout(w_dff_A_c53COlZH7_0),.din(w_dff_A_QujEOu9A6_0),.clk(gclk));
	jdff dff_A_c53COlZH7_0(.dout(w_dff_A_EkkJoVIu3_0),.din(w_dff_A_c53COlZH7_0),.clk(gclk));
	jdff dff_A_EkkJoVIu3_0(.dout(w_dff_A_FtCXtbQg9_0),.din(w_dff_A_EkkJoVIu3_0),.clk(gclk));
	jdff dff_A_FtCXtbQg9_0(.dout(w_dff_A_vAmYOYGm1_0),.din(w_dff_A_FtCXtbQg9_0),.clk(gclk));
	jdff dff_A_vAmYOYGm1_0(.dout(w_dff_A_ZESBphvC5_0),.din(w_dff_A_vAmYOYGm1_0),.clk(gclk));
	jdff dff_A_ZESBphvC5_0(.dout(w_dff_A_uRDFrFV11_0),.din(w_dff_A_ZESBphvC5_0),.clk(gclk));
	jdff dff_A_uRDFrFV11_0(.dout(w_dff_A_JJxzZPom5_0),.din(w_dff_A_uRDFrFV11_0),.clk(gclk));
	jdff dff_A_JJxzZPom5_0(.dout(w_dff_A_zLTGmJ074_0),.din(w_dff_A_JJxzZPom5_0),.clk(gclk));
	jdff dff_A_zLTGmJ074_0(.dout(w_dff_A_6Q65BMSk9_0),.din(w_dff_A_zLTGmJ074_0),.clk(gclk));
	jdff dff_A_6Q65BMSk9_0(.dout(w_dff_A_g2OhW2KO0_0),.din(w_dff_A_6Q65BMSk9_0),.clk(gclk));
	jdff dff_A_g2OhW2KO0_0(.dout(w_dff_A_MkI2c3Bi5_0),.din(w_dff_A_g2OhW2KO0_0),.clk(gclk));
	jdff dff_A_MkI2c3Bi5_0(.dout(sin1),.din(w_dff_A_MkI2c3Bi5_0),.clk(gclk));
	jdff dff_A_N1eAxMfr7_2(.dout(w_dff_A_Rq5spMDm0_0),.din(w_dff_A_N1eAxMfr7_2),.clk(gclk));
	jdff dff_A_Rq5spMDm0_0(.dout(w_dff_A_i9nintPf9_0),.din(w_dff_A_Rq5spMDm0_0),.clk(gclk));
	jdff dff_A_i9nintPf9_0(.dout(w_dff_A_AblW14053_0),.din(w_dff_A_i9nintPf9_0),.clk(gclk));
	jdff dff_A_AblW14053_0(.dout(w_dff_A_6dVfI5uI0_0),.din(w_dff_A_AblW14053_0),.clk(gclk));
	jdff dff_A_6dVfI5uI0_0(.dout(w_dff_A_n8tTywNa8_0),.din(w_dff_A_6dVfI5uI0_0),.clk(gclk));
	jdff dff_A_n8tTywNa8_0(.dout(w_dff_A_UMCcn4bR2_0),.din(w_dff_A_n8tTywNa8_0),.clk(gclk));
	jdff dff_A_UMCcn4bR2_0(.dout(w_dff_A_NUur3pNc7_0),.din(w_dff_A_UMCcn4bR2_0),.clk(gclk));
	jdff dff_A_NUur3pNc7_0(.dout(w_dff_A_p3ALE3In6_0),.din(w_dff_A_NUur3pNc7_0),.clk(gclk));
	jdff dff_A_p3ALE3In6_0(.dout(w_dff_A_NNjP8ur99_0),.din(w_dff_A_p3ALE3In6_0),.clk(gclk));
	jdff dff_A_NNjP8ur99_0(.dout(w_dff_A_I6THQCKm2_0),.din(w_dff_A_NNjP8ur99_0),.clk(gclk));
	jdff dff_A_I6THQCKm2_0(.dout(w_dff_A_oDiZMTry0_0),.din(w_dff_A_I6THQCKm2_0),.clk(gclk));
	jdff dff_A_oDiZMTry0_0(.dout(w_dff_A_T9qHtUv04_0),.din(w_dff_A_oDiZMTry0_0),.clk(gclk));
	jdff dff_A_T9qHtUv04_0(.dout(w_dff_A_J261o2Ss1_0),.din(w_dff_A_T9qHtUv04_0),.clk(gclk));
	jdff dff_A_J261o2Ss1_0(.dout(w_dff_A_gb1thYBX5_0),.din(w_dff_A_J261o2Ss1_0),.clk(gclk));
	jdff dff_A_gb1thYBX5_0(.dout(w_dff_A_OOVB7UZJ9_0),.din(w_dff_A_gb1thYBX5_0),.clk(gclk));
	jdff dff_A_OOVB7UZJ9_0(.dout(w_dff_A_PduTcBVN6_0),.din(w_dff_A_OOVB7UZJ9_0),.clk(gclk));
	jdff dff_A_PduTcBVN6_0(.dout(w_dff_A_2Rx7qi8X1_0),.din(w_dff_A_PduTcBVN6_0),.clk(gclk));
	jdff dff_A_2Rx7qi8X1_0(.dout(w_dff_A_ibZGM0ph6_0),.din(w_dff_A_2Rx7qi8X1_0),.clk(gclk));
	jdff dff_A_ibZGM0ph6_0(.dout(w_dff_A_LlfKHEXB0_0),.din(w_dff_A_ibZGM0ph6_0),.clk(gclk));
	jdff dff_A_LlfKHEXB0_0(.dout(w_dff_A_dZYeahfo5_0),.din(w_dff_A_LlfKHEXB0_0),.clk(gclk));
	jdff dff_A_dZYeahfo5_0(.dout(w_dff_A_MVwpyAgL3_0),.din(w_dff_A_dZYeahfo5_0),.clk(gclk));
	jdff dff_A_MVwpyAgL3_0(.dout(w_dff_A_Dxjd7JBQ6_0),.din(w_dff_A_MVwpyAgL3_0),.clk(gclk));
	jdff dff_A_Dxjd7JBQ6_0(.dout(w_dff_A_Z7ToR5508_0),.din(w_dff_A_Dxjd7JBQ6_0),.clk(gclk));
	jdff dff_A_Z7ToR5508_0(.dout(w_dff_A_xr2NpMAe7_0),.din(w_dff_A_Z7ToR5508_0),.clk(gclk));
	jdff dff_A_xr2NpMAe7_0(.dout(w_dff_A_B2LKw6Hh0_0),.din(w_dff_A_xr2NpMAe7_0),.clk(gclk));
	jdff dff_A_B2LKw6Hh0_0(.dout(w_dff_A_ny4AM0fk2_0),.din(w_dff_A_B2LKw6Hh0_0),.clk(gclk));
	jdff dff_A_ny4AM0fk2_0(.dout(w_dff_A_jNH3n5Mv4_0),.din(w_dff_A_ny4AM0fk2_0),.clk(gclk));
	jdff dff_A_jNH3n5Mv4_0(.dout(w_dff_A_B1EZ8cCP3_0),.din(w_dff_A_jNH3n5Mv4_0),.clk(gclk));
	jdff dff_A_B1EZ8cCP3_0(.dout(w_dff_A_gZpOUTGo5_0),.din(w_dff_A_B1EZ8cCP3_0),.clk(gclk));
	jdff dff_A_gZpOUTGo5_0(.dout(w_dff_A_ns0uvPKF4_0),.din(w_dff_A_gZpOUTGo5_0),.clk(gclk));
	jdff dff_A_ns0uvPKF4_0(.dout(w_dff_A_D5etW4Tb0_0),.din(w_dff_A_ns0uvPKF4_0),.clk(gclk));
	jdff dff_A_D5etW4Tb0_0(.dout(w_dff_A_TMcxvjUk7_0),.din(w_dff_A_D5etW4Tb0_0),.clk(gclk));
	jdff dff_A_TMcxvjUk7_0(.dout(w_dff_A_wuUwQJDP6_0),.din(w_dff_A_TMcxvjUk7_0),.clk(gclk));
	jdff dff_A_wuUwQJDP6_0(.dout(w_dff_A_ZnA4sBYo1_0),.din(w_dff_A_wuUwQJDP6_0),.clk(gclk));
	jdff dff_A_ZnA4sBYo1_0(.dout(w_dff_A_qmQpENUI5_0),.din(w_dff_A_ZnA4sBYo1_0),.clk(gclk));
	jdff dff_A_qmQpENUI5_0(.dout(w_dff_A_UmRC19KI8_0),.din(w_dff_A_qmQpENUI5_0),.clk(gclk));
	jdff dff_A_UmRC19KI8_0(.dout(w_dff_A_UhCzM3vJ9_0),.din(w_dff_A_UmRC19KI8_0),.clk(gclk));
	jdff dff_A_UhCzM3vJ9_0(.dout(w_dff_A_9rl593Pk8_0),.din(w_dff_A_UhCzM3vJ9_0),.clk(gclk));
	jdff dff_A_9rl593Pk8_0(.dout(w_dff_A_Qcnenz3c3_0),.din(w_dff_A_9rl593Pk8_0),.clk(gclk));
	jdff dff_A_Qcnenz3c3_0(.dout(w_dff_A_GzWX4srB6_0),.din(w_dff_A_Qcnenz3c3_0),.clk(gclk));
	jdff dff_A_GzWX4srB6_0(.dout(sin2),.din(w_dff_A_GzWX4srB6_0),.clk(gclk));
	jdff dff_A_GpXyXXB64_2(.dout(w_dff_A_ALipnorC1_0),.din(w_dff_A_GpXyXXB64_2),.clk(gclk));
	jdff dff_A_ALipnorC1_0(.dout(w_dff_A_XhjQDMNB6_0),.din(w_dff_A_ALipnorC1_0),.clk(gclk));
	jdff dff_A_XhjQDMNB6_0(.dout(w_dff_A_7H1A6hjr8_0),.din(w_dff_A_XhjQDMNB6_0),.clk(gclk));
	jdff dff_A_7H1A6hjr8_0(.dout(w_dff_A_84qVARgy6_0),.din(w_dff_A_7H1A6hjr8_0),.clk(gclk));
	jdff dff_A_84qVARgy6_0(.dout(w_dff_A_cwKIrz4B6_0),.din(w_dff_A_84qVARgy6_0),.clk(gclk));
	jdff dff_A_cwKIrz4B6_0(.dout(w_dff_A_9YKuMTny4_0),.din(w_dff_A_cwKIrz4B6_0),.clk(gclk));
	jdff dff_A_9YKuMTny4_0(.dout(w_dff_A_kAOXuQAV5_0),.din(w_dff_A_9YKuMTny4_0),.clk(gclk));
	jdff dff_A_kAOXuQAV5_0(.dout(w_dff_A_PeA6fPhU6_0),.din(w_dff_A_kAOXuQAV5_0),.clk(gclk));
	jdff dff_A_PeA6fPhU6_0(.dout(w_dff_A_D7FMRUwh7_0),.din(w_dff_A_PeA6fPhU6_0),.clk(gclk));
	jdff dff_A_D7FMRUwh7_0(.dout(w_dff_A_miLhcljX0_0),.din(w_dff_A_D7FMRUwh7_0),.clk(gclk));
	jdff dff_A_miLhcljX0_0(.dout(w_dff_A_fa7iecpj0_0),.din(w_dff_A_miLhcljX0_0),.clk(gclk));
	jdff dff_A_fa7iecpj0_0(.dout(w_dff_A_r0qUSK9q1_0),.din(w_dff_A_fa7iecpj0_0),.clk(gclk));
	jdff dff_A_r0qUSK9q1_0(.dout(w_dff_A_7AXVUXh24_0),.din(w_dff_A_r0qUSK9q1_0),.clk(gclk));
	jdff dff_A_7AXVUXh24_0(.dout(w_dff_A_v9AKyfJg1_0),.din(w_dff_A_7AXVUXh24_0),.clk(gclk));
	jdff dff_A_v9AKyfJg1_0(.dout(w_dff_A_h3u6UiJg2_0),.din(w_dff_A_v9AKyfJg1_0),.clk(gclk));
	jdff dff_A_h3u6UiJg2_0(.dout(w_dff_A_88rRlTUG7_0),.din(w_dff_A_h3u6UiJg2_0),.clk(gclk));
	jdff dff_A_88rRlTUG7_0(.dout(w_dff_A_UlO6ny3g1_0),.din(w_dff_A_88rRlTUG7_0),.clk(gclk));
	jdff dff_A_UlO6ny3g1_0(.dout(w_dff_A_EW0FfGZY6_0),.din(w_dff_A_UlO6ny3g1_0),.clk(gclk));
	jdff dff_A_EW0FfGZY6_0(.dout(w_dff_A_JhvnjQke7_0),.din(w_dff_A_EW0FfGZY6_0),.clk(gclk));
	jdff dff_A_JhvnjQke7_0(.dout(w_dff_A_lGeebp1P5_0),.din(w_dff_A_JhvnjQke7_0),.clk(gclk));
	jdff dff_A_lGeebp1P5_0(.dout(w_dff_A_DAsj5WNq9_0),.din(w_dff_A_lGeebp1P5_0),.clk(gclk));
	jdff dff_A_DAsj5WNq9_0(.dout(w_dff_A_joayAzx24_0),.din(w_dff_A_DAsj5WNq9_0),.clk(gclk));
	jdff dff_A_joayAzx24_0(.dout(w_dff_A_8D4lveQN6_0),.din(w_dff_A_joayAzx24_0),.clk(gclk));
	jdff dff_A_8D4lveQN6_0(.dout(w_dff_A_uVeIlb1G3_0),.din(w_dff_A_8D4lveQN6_0),.clk(gclk));
	jdff dff_A_uVeIlb1G3_0(.dout(w_dff_A_7uCWuWUr2_0),.din(w_dff_A_uVeIlb1G3_0),.clk(gclk));
	jdff dff_A_7uCWuWUr2_0(.dout(w_dff_A_Mq2S7sZk4_0),.din(w_dff_A_7uCWuWUr2_0),.clk(gclk));
	jdff dff_A_Mq2S7sZk4_0(.dout(w_dff_A_nER4U6K48_0),.din(w_dff_A_Mq2S7sZk4_0),.clk(gclk));
	jdff dff_A_nER4U6K48_0(.dout(w_dff_A_IZv0YM7F1_0),.din(w_dff_A_nER4U6K48_0),.clk(gclk));
	jdff dff_A_IZv0YM7F1_0(.dout(w_dff_A_crm6Esgu7_0),.din(w_dff_A_IZv0YM7F1_0),.clk(gclk));
	jdff dff_A_crm6Esgu7_0(.dout(w_dff_A_OFoQEhMQ7_0),.din(w_dff_A_crm6Esgu7_0),.clk(gclk));
	jdff dff_A_OFoQEhMQ7_0(.dout(w_dff_A_T3cjDN794_0),.din(w_dff_A_OFoQEhMQ7_0),.clk(gclk));
	jdff dff_A_T3cjDN794_0(.dout(w_dff_A_70WuzKR46_0),.din(w_dff_A_T3cjDN794_0),.clk(gclk));
	jdff dff_A_70WuzKR46_0(.dout(w_dff_A_17BjVtui6_0),.din(w_dff_A_70WuzKR46_0),.clk(gclk));
	jdff dff_A_17BjVtui6_0(.dout(w_dff_A_A6PQVR7i4_0),.din(w_dff_A_17BjVtui6_0),.clk(gclk));
	jdff dff_A_A6PQVR7i4_0(.dout(w_dff_A_azR70T864_0),.din(w_dff_A_A6PQVR7i4_0),.clk(gclk));
	jdff dff_A_azR70T864_0(.dout(w_dff_A_6eS7l4G83_0),.din(w_dff_A_azR70T864_0),.clk(gclk));
	jdff dff_A_6eS7l4G83_0(.dout(w_dff_A_rreE02PC5_0),.din(w_dff_A_6eS7l4G83_0),.clk(gclk));
	jdff dff_A_rreE02PC5_0(.dout(w_dff_A_e5QaUZSQ6_0),.din(w_dff_A_rreE02PC5_0),.clk(gclk));
	jdff dff_A_e5QaUZSQ6_0(.dout(sin3),.din(w_dff_A_e5QaUZSQ6_0),.clk(gclk));
	jdff dff_A_Kjg55Kq01_2(.dout(w_dff_A_exl6Wb7n2_0),.din(w_dff_A_Kjg55Kq01_2),.clk(gclk));
	jdff dff_A_exl6Wb7n2_0(.dout(w_dff_A_ClGP5wdM3_0),.din(w_dff_A_exl6Wb7n2_0),.clk(gclk));
	jdff dff_A_ClGP5wdM3_0(.dout(w_dff_A_u3xdwEuT4_0),.din(w_dff_A_ClGP5wdM3_0),.clk(gclk));
	jdff dff_A_u3xdwEuT4_0(.dout(w_dff_A_iEubiO8B1_0),.din(w_dff_A_u3xdwEuT4_0),.clk(gclk));
	jdff dff_A_iEubiO8B1_0(.dout(w_dff_A_ruNAGpa23_0),.din(w_dff_A_iEubiO8B1_0),.clk(gclk));
	jdff dff_A_ruNAGpa23_0(.dout(w_dff_A_mCcryNGs9_0),.din(w_dff_A_ruNAGpa23_0),.clk(gclk));
	jdff dff_A_mCcryNGs9_0(.dout(w_dff_A_NCFpvP1o3_0),.din(w_dff_A_mCcryNGs9_0),.clk(gclk));
	jdff dff_A_NCFpvP1o3_0(.dout(w_dff_A_KIkikeco2_0),.din(w_dff_A_NCFpvP1o3_0),.clk(gclk));
	jdff dff_A_KIkikeco2_0(.dout(w_dff_A_e1vnGn374_0),.din(w_dff_A_KIkikeco2_0),.clk(gclk));
	jdff dff_A_e1vnGn374_0(.dout(w_dff_A_sMop9cDf7_0),.din(w_dff_A_e1vnGn374_0),.clk(gclk));
	jdff dff_A_sMop9cDf7_0(.dout(w_dff_A_r2Fd3AFe4_0),.din(w_dff_A_sMop9cDf7_0),.clk(gclk));
	jdff dff_A_r2Fd3AFe4_0(.dout(w_dff_A_z2psqKaj4_0),.din(w_dff_A_r2Fd3AFe4_0),.clk(gclk));
	jdff dff_A_z2psqKaj4_0(.dout(w_dff_A_dza0UVxx8_0),.din(w_dff_A_z2psqKaj4_0),.clk(gclk));
	jdff dff_A_dza0UVxx8_0(.dout(w_dff_A_Xq7W6AMn2_0),.din(w_dff_A_dza0UVxx8_0),.clk(gclk));
	jdff dff_A_Xq7W6AMn2_0(.dout(w_dff_A_FY2QkzWg3_0),.din(w_dff_A_Xq7W6AMn2_0),.clk(gclk));
	jdff dff_A_FY2QkzWg3_0(.dout(w_dff_A_HqbCpj6h4_0),.din(w_dff_A_FY2QkzWg3_0),.clk(gclk));
	jdff dff_A_HqbCpj6h4_0(.dout(w_dff_A_FVmRCHvx7_0),.din(w_dff_A_HqbCpj6h4_0),.clk(gclk));
	jdff dff_A_FVmRCHvx7_0(.dout(w_dff_A_YeI9e0lF3_0),.din(w_dff_A_FVmRCHvx7_0),.clk(gclk));
	jdff dff_A_YeI9e0lF3_0(.dout(w_dff_A_izyZBich0_0),.din(w_dff_A_YeI9e0lF3_0),.clk(gclk));
	jdff dff_A_izyZBich0_0(.dout(w_dff_A_8tKQAvOq7_0),.din(w_dff_A_izyZBich0_0),.clk(gclk));
	jdff dff_A_8tKQAvOq7_0(.dout(w_dff_A_YXYPFMNK8_0),.din(w_dff_A_8tKQAvOq7_0),.clk(gclk));
	jdff dff_A_YXYPFMNK8_0(.dout(w_dff_A_BPX4faWu2_0),.din(w_dff_A_YXYPFMNK8_0),.clk(gclk));
	jdff dff_A_BPX4faWu2_0(.dout(w_dff_A_gAdfh5234_0),.din(w_dff_A_BPX4faWu2_0),.clk(gclk));
	jdff dff_A_gAdfh5234_0(.dout(w_dff_A_Af6nxECs9_0),.din(w_dff_A_gAdfh5234_0),.clk(gclk));
	jdff dff_A_Af6nxECs9_0(.dout(w_dff_A_3xZjHrmI4_0),.din(w_dff_A_Af6nxECs9_0),.clk(gclk));
	jdff dff_A_3xZjHrmI4_0(.dout(w_dff_A_Oy88hPKX9_0),.din(w_dff_A_3xZjHrmI4_0),.clk(gclk));
	jdff dff_A_Oy88hPKX9_0(.dout(w_dff_A_nE3iIpth5_0),.din(w_dff_A_Oy88hPKX9_0),.clk(gclk));
	jdff dff_A_nE3iIpth5_0(.dout(w_dff_A_tMJTaLlv9_0),.din(w_dff_A_nE3iIpth5_0),.clk(gclk));
	jdff dff_A_tMJTaLlv9_0(.dout(w_dff_A_n8Gz5rOt8_0),.din(w_dff_A_tMJTaLlv9_0),.clk(gclk));
	jdff dff_A_n8Gz5rOt8_0(.dout(w_dff_A_bgY8fUOw5_0),.din(w_dff_A_n8Gz5rOt8_0),.clk(gclk));
	jdff dff_A_bgY8fUOw5_0(.dout(w_dff_A_S6B5c8LW1_0),.din(w_dff_A_bgY8fUOw5_0),.clk(gclk));
	jdff dff_A_S6B5c8LW1_0(.dout(w_dff_A_rGTXUjBc0_0),.din(w_dff_A_S6B5c8LW1_0),.clk(gclk));
	jdff dff_A_rGTXUjBc0_0(.dout(w_dff_A_svb5edEV5_0),.din(w_dff_A_rGTXUjBc0_0),.clk(gclk));
	jdff dff_A_svb5edEV5_0(.dout(w_dff_A_QJRbqGjc5_0),.din(w_dff_A_svb5edEV5_0),.clk(gclk));
	jdff dff_A_QJRbqGjc5_0(.dout(w_dff_A_TXtnJcIN5_0),.din(w_dff_A_QJRbqGjc5_0),.clk(gclk));
	jdff dff_A_TXtnJcIN5_0(.dout(w_dff_A_hqtUx4ZL7_0),.din(w_dff_A_TXtnJcIN5_0),.clk(gclk));
	jdff dff_A_hqtUx4ZL7_0(.dout(sin4),.din(w_dff_A_hqtUx4ZL7_0),.clk(gclk));
	jdff dff_A_jawdh4xz8_2(.dout(w_dff_A_9iV3vboV8_0),.din(w_dff_A_jawdh4xz8_2),.clk(gclk));
	jdff dff_A_9iV3vboV8_0(.dout(w_dff_A_mUGqYtG34_0),.din(w_dff_A_9iV3vboV8_0),.clk(gclk));
	jdff dff_A_mUGqYtG34_0(.dout(w_dff_A_PHsUUrIT5_0),.din(w_dff_A_mUGqYtG34_0),.clk(gclk));
	jdff dff_A_PHsUUrIT5_0(.dout(w_dff_A_5dj5NOr98_0),.din(w_dff_A_PHsUUrIT5_0),.clk(gclk));
	jdff dff_A_5dj5NOr98_0(.dout(w_dff_A_9epO0p3g9_0),.din(w_dff_A_5dj5NOr98_0),.clk(gclk));
	jdff dff_A_9epO0p3g9_0(.dout(w_dff_A_JduSHjIT0_0),.din(w_dff_A_9epO0p3g9_0),.clk(gclk));
	jdff dff_A_JduSHjIT0_0(.dout(w_dff_A_9iJivsOC3_0),.din(w_dff_A_JduSHjIT0_0),.clk(gclk));
	jdff dff_A_9iJivsOC3_0(.dout(w_dff_A_Ym1Im8Jw5_0),.din(w_dff_A_9iJivsOC3_0),.clk(gclk));
	jdff dff_A_Ym1Im8Jw5_0(.dout(w_dff_A_S5O0Fwqf6_0),.din(w_dff_A_Ym1Im8Jw5_0),.clk(gclk));
	jdff dff_A_S5O0Fwqf6_0(.dout(w_dff_A_R9HyIRHj3_0),.din(w_dff_A_S5O0Fwqf6_0),.clk(gclk));
	jdff dff_A_R9HyIRHj3_0(.dout(w_dff_A_BiKzDwcT5_0),.din(w_dff_A_R9HyIRHj3_0),.clk(gclk));
	jdff dff_A_BiKzDwcT5_0(.dout(w_dff_A_OsQhl5lF6_0),.din(w_dff_A_BiKzDwcT5_0),.clk(gclk));
	jdff dff_A_OsQhl5lF6_0(.dout(w_dff_A_pzaFM3mo6_0),.din(w_dff_A_OsQhl5lF6_0),.clk(gclk));
	jdff dff_A_pzaFM3mo6_0(.dout(w_dff_A_n0WZ2Xct9_0),.din(w_dff_A_pzaFM3mo6_0),.clk(gclk));
	jdff dff_A_n0WZ2Xct9_0(.dout(w_dff_A_VqCDgc329_0),.din(w_dff_A_n0WZ2Xct9_0),.clk(gclk));
	jdff dff_A_VqCDgc329_0(.dout(w_dff_A_3Uak3UhB5_0),.din(w_dff_A_VqCDgc329_0),.clk(gclk));
	jdff dff_A_3Uak3UhB5_0(.dout(w_dff_A_LxsMLQuO6_0),.din(w_dff_A_3Uak3UhB5_0),.clk(gclk));
	jdff dff_A_LxsMLQuO6_0(.dout(w_dff_A_5ZFq95xx6_0),.din(w_dff_A_LxsMLQuO6_0),.clk(gclk));
	jdff dff_A_5ZFq95xx6_0(.dout(w_dff_A_2cwPZCds0_0),.din(w_dff_A_5ZFq95xx6_0),.clk(gclk));
	jdff dff_A_2cwPZCds0_0(.dout(w_dff_A_zSbL8nS36_0),.din(w_dff_A_2cwPZCds0_0),.clk(gclk));
	jdff dff_A_zSbL8nS36_0(.dout(w_dff_A_fhU1izvd1_0),.din(w_dff_A_zSbL8nS36_0),.clk(gclk));
	jdff dff_A_fhU1izvd1_0(.dout(w_dff_A_JmUqeRJK8_0),.din(w_dff_A_fhU1izvd1_0),.clk(gclk));
	jdff dff_A_JmUqeRJK8_0(.dout(w_dff_A_D73D64gy7_0),.din(w_dff_A_JmUqeRJK8_0),.clk(gclk));
	jdff dff_A_D73D64gy7_0(.dout(w_dff_A_1zth1a1g5_0),.din(w_dff_A_D73D64gy7_0),.clk(gclk));
	jdff dff_A_1zth1a1g5_0(.dout(w_dff_A_Qx9kCEGX2_0),.din(w_dff_A_1zth1a1g5_0),.clk(gclk));
	jdff dff_A_Qx9kCEGX2_0(.dout(w_dff_A_EpvSigF52_0),.din(w_dff_A_Qx9kCEGX2_0),.clk(gclk));
	jdff dff_A_EpvSigF52_0(.dout(w_dff_A_DtBBIc706_0),.din(w_dff_A_EpvSigF52_0),.clk(gclk));
	jdff dff_A_DtBBIc706_0(.dout(w_dff_A_uGsoqZmV7_0),.din(w_dff_A_DtBBIc706_0),.clk(gclk));
	jdff dff_A_uGsoqZmV7_0(.dout(w_dff_A_x4HO3zVQ9_0),.din(w_dff_A_uGsoqZmV7_0),.clk(gclk));
	jdff dff_A_x4HO3zVQ9_0(.dout(w_dff_A_fMOgHJeK9_0),.din(w_dff_A_x4HO3zVQ9_0),.clk(gclk));
	jdff dff_A_fMOgHJeK9_0(.dout(w_dff_A_B6YdI7do9_0),.din(w_dff_A_fMOgHJeK9_0),.clk(gclk));
	jdff dff_A_B6YdI7do9_0(.dout(w_dff_A_gHKRirfE3_0),.din(w_dff_A_B6YdI7do9_0),.clk(gclk));
	jdff dff_A_gHKRirfE3_0(.dout(w_dff_A_Cn401hVH9_0),.din(w_dff_A_gHKRirfE3_0),.clk(gclk));
	jdff dff_A_Cn401hVH9_0(.dout(w_dff_A_D333eUok3_0),.din(w_dff_A_Cn401hVH9_0),.clk(gclk));
	jdff dff_A_D333eUok3_0(.dout(sin5),.din(w_dff_A_D333eUok3_0),.clk(gclk));
	jdff dff_A_Pe38P7pN5_2(.dout(w_dff_A_nCtEnPSJ2_0),.din(w_dff_A_Pe38P7pN5_2),.clk(gclk));
	jdff dff_A_nCtEnPSJ2_0(.dout(w_dff_A_Ma3O3KvU1_0),.din(w_dff_A_nCtEnPSJ2_0),.clk(gclk));
	jdff dff_A_Ma3O3KvU1_0(.dout(w_dff_A_Ep7KrQup3_0),.din(w_dff_A_Ma3O3KvU1_0),.clk(gclk));
	jdff dff_A_Ep7KrQup3_0(.dout(w_dff_A_e6ZbUdPx9_0),.din(w_dff_A_Ep7KrQup3_0),.clk(gclk));
	jdff dff_A_e6ZbUdPx9_0(.dout(w_dff_A_msOno7Ka6_0),.din(w_dff_A_e6ZbUdPx9_0),.clk(gclk));
	jdff dff_A_msOno7Ka6_0(.dout(w_dff_A_tqzbhEqh8_0),.din(w_dff_A_msOno7Ka6_0),.clk(gclk));
	jdff dff_A_tqzbhEqh8_0(.dout(w_dff_A_fsO3fsos1_0),.din(w_dff_A_tqzbhEqh8_0),.clk(gclk));
	jdff dff_A_fsO3fsos1_0(.dout(w_dff_A_ghzjACQP6_0),.din(w_dff_A_fsO3fsos1_0),.clk(gclk));
	jdff dff_A_ghzjACQP6_0(.dout(w_dff_A_TDvTJT7n3_0),.din(w_dff_A_ghzjACQP6_0),.clk(gclk));
	jdff dff_A_TDvTJT7n3_0(.dout(w_dff_A_CXJZvFPU5_0),.din(w_dff_A_TDvTJT7n3_0),.clk(gclk));
	jdff dff_A_CXJZvFPU5_0(.dout(w_dff_A_uyTcqu9B1_0),.din(w_dff_A_CXJZvFPU5_0),.clk(gclk));
	jdff dff_A_uyTcqu9B1_0(.dout(w_dff_A_Q2bnUvrU5_0),.din(w_dff_A_uyTcqu9B1_0),.clk(gclk));
	jdff dff_A_Q2bnUvrU5_0(.dout(w_dff_A_wbCW6RWZ7_0),.din(w_dff_A_Q2bnUvrU5_0),.clk(gclk));
	jdff dff_A_wbCW6RWZ7_0(.dout(w_dff_A_zU6d6cKq6_0),.din(w_dff_A_wbCW6RWZ7_0),.clk(gclk));
	jdff dff_A_zU6d6cKq6_0(.dout(w_dff_A_5b9FxAtZ5_0),.din(w_dff_A_zU6d6cKq6_0),.clk(gclk));
	jdff dff_A_5b9FxAtZ5_0(.dout(w_dff_A_IDaLhTdA5_0),.din(w_dff_A_5b9FxAtZ5_0),.clk(gclk));
	jdff dff_A_IDaLhTdA5_0(.dout(w_dff_A_VT3BquvT5_0),.din(w_dff_A_IDaLhTdA5_0),.clk(gclk));
	jdff dff_A_VT3BquvT5_0(.dout(w_dff_A_f21aEBkc3_0),.din(w_dff_A_VT3BquvT5_0),.clk(gclk));
	jdff dff_A_f21aEBkc3_0(.dout(w_dff_A_mMSm4fmZ2_0),.din(w_dff_A_f21aEBkc3_0),.clk(gclk));
	jdff dff_A_mMSm4fmZ2_0(.dout(w_dff_A_g14aAOT03_0),.din(w_dff_A_mMSm4fmZ2_0),.clk(gclk));
	jdff dff_A_g14aAOT03_0(.dout(w_dff_A_tAQiefrK0_0),.din(w_dff_A_g14aAOT03_0),.clk(gclk));
	jdff dff_A_tAQiefrK0_0(.dout(w_dff_A_XNb9bnLK7_0),.din(w_dff_A_tAQiefrK0_0),.clk(gclk));
	jdff dff_A_XNb9bnLK7_0(.dout(w_dff_A_Z4LR6hMY9_0),.din(w_dff_A_XNb9bnLK7_0),.clk(gclk));
	jdff dff_A_Z4LR6hMY9_0(.dout(w_dff_A_8XUyS7db8_0),.din(w_dff_A_Z4LR6hMY9_0),.clk(gclk));
	jdff dff_A_8XUyS7db8_0(.dout(w_dff_A_jjEQFNqj1_0),.din(w_dff_A_8XUyS7db8_0),.clk(gclk));
	jdff dff_A_jjEQFNqj1_0(.dout(w_dff_A_1troq28w6_0),.din(w_dff_A_jjEQFNqj1_0),.clk(gclk));
	jdff dff_A_1troq28w6_0(.dout(w_dff_A_VYoYmtW93_0),.din(w_dff_A_1troq28w6_0),.clk(gclk));
	jdff dff_A_VYoYmtW93_0(.dout(w_dff_A_GPXb8OUm1_0),.din(w_dff_A_VYoYmtW93_0),.clk(gclk));
	jdff dff_A_GPXb8OUm1_0(.dout(w_dff_A_uZYSGDVi8_0),.din(w_dff_A_GPXb8OUm1_0),.clk(gclk));
	jdff dff_A_uZYSGDVi8_0(.dout(w_dff_A_2VRka1ES2_0),.din(w_dff_A_uZYSGDVi8_0),.clk(gclk));
	jdff dff_A_2VRka1ES2_0(.dout(w_dff_A_YkMkjnyG3_0),.din(w_dff_A_2VRka1ES2_0),.clk(gclk));
	jdff dff_A_YkMkjnyG3_0(.dout(w_dff_A_gSW324tT4_0),.din(w_dff_A_YkMkjnyG3_0),.clk(gclk));
	jdff dff_A_gSW324tT4_0(.dout(sin6),.din(w_dff_A_gSW324tT4_0),.clk(gclk));
	jdff dff_A_64zGTwWk3_2(.dout(w_dff_A_uoBovu303_0),.din(w_dff_A_64zGTwWk3_2),.clk(gclk));
	jdff dff_A_uoBovu303_0(.dout(w_dff_A_lWdZZcdk5_0),.din(w_dff_A_uoBovu303_0),.clk(gclk));
	jdff dff_A_lWdZZcdk5_0(.dout(w_dff_A_XBM05sUU2_0),.din(w_dff_A_lWdZZcdk5_0),.clk(gclk));
	jdff dff_A_XBM05sUU2_0(.dout(w_dff_A_DO1RDvC50_0),.din(w_dff_A_XBM05sUU2_0),.clk(gclk));
	jdff dff_A_DO1RDvC50_0(.dout(w_dff_A_AjYtVRkR7_0),.din(w_dff_A_DO1RDvC50_0),.clk(gclk));
	jdff dff_A_AjYtVRkR7_0(.dout(w_dff_A_bK1kIERF9_0),.din(w_dff_A_AjYtVRkR7_0),.clk(gclk));
	jdff dff_A_bK1kIERF9_0(.dout(w_dff_A_AKHF9kOM8_0),.din(w_dff_A_bK1kIERF9_0),.clk(gclk));
	jdff dff_A_AKHF9kOM8_0(.dout(w_dff_A_KhCy3EHF8_0),.din(w_dff_A_AKHF9kOM8_0),.clk(gclk));
	jdff dff_A_KhCy3EHF8_0(.dout(w_dff_A_glSHPEDr3_0),.din(w_dff_A_KhCy3EHF8_0),.clk(gclk));
	jdff dff_A_glSHPEDr3_0(.dout(w_dff_A_hxHpYU7r5_0),.din(w_dff_A_glSHPEDr3_0),.clk(gclk));
	jdff dff_A_hxHpYU7r5_0(.dout(w_dff_A_8GHlr7Q89_0),.din(w_dff_A_hxHpYU7r5_0),.clk(gclk));
	jdff dff_A_8GHlr7Q89_0(.dout(w_dff_A_VOejKKPC9_0),.din(w_dff_A_8GHlr7Q89_0),.clk(gclk));
	jdff dff_A_VOejKKPC9_0(.dout(w_dff_A_7pUuxhwX7_0),.din(w_dff_A_VOejKKPC9_0),.clk(gclk));
	jdff dff_A_7pUuxhwX7_0(.dout(w_dff_A_P99XQ2265_0),.din(w_dff_A_7pUuxhwX7_0),.clk(gclk));
	jdff dff_A_P99XQ2265_0(.dout(w_dff_A_VF9FwnGg7_0),.din(w_dff_A_P99XQ2265_0),.clk(gclk));
	jdff dff_A_VF9FwnGg7_0(.dout(w_dff_A_DdghD26L5_0),.din(w_dff_A_VF9FwnGg7_0),.clk(gclk));
	jdff dff_A_DdghD26L5_0(.dout(w_dff_A_BDvvNO2J5_0),.din(w_dff_A_DdghD26L5_0),.clk(gclk));
	jdff dff_A_BDvvNO2J5_0(.dout(w_dff_A_hCOdVZp18_0),.din(w_dff_A_BDvvNO2J5_0),.clk(gclk));
	jdff dff_A_hCOdVZp18_0(.dout(w_dff_A_4hSfu2Ow5_0),.din(w_dff_A_hCOdVZp18_0),.clk(gclk));
	jdff dff_A_4hSfu2Ow5_0(.dout(w_dff_A_DYm5XO3d1_0),.din(w_dff_A_4hSfu2Ow5_0),.clk(gclk));
	jdff dff_A_DYm5XO3d1_0(.dout(w_dff_A_gpyHIEUg6_0),.din(w_dff_A_DYm5XO3d1_0),.clk(gclk));
	jdff dff_A_gpyHIEUg6_0(.dout(w_dff_A_ag1chzb80_0),.din(w_dff_A_gpyHIEUg6_0),.clk(gclk));
	jdff dff_A_ag1chzb80_0(.dout(w_dff_A_b8ff46Sh1_0),.din(w_dff_A_ag1chzb80_0),.clk(gclk));
	jdff dff_A_b8ff46Sh1_0(.dout(w_dff_A_5RXLLOWz5_0),.din(w_dff_A_b8ff46Sh1_0),.clk(gclk));
	jdff dff_A_5RXLLOWz5_0(.dout(w_dff_A_Q9sgvRmZ2_0),.din(w_dff_A_5RXLLOWz5_0),.clk(gclk));
	jdff dff_A_Q9sgvRmZ2_0(.dout(w_dff_A_GaacqGqW2_0),.din(w_dff_A_Q9sgvRmZ2_0),.clk(gclk));
	jdff dff_A_GaacqGqW2_0(.dout(w_dff_A_LWnl3p6B3_0),.din(w_dff_A_GaacqGqW2_0),.clk(gclk));
	jdff dff_A_LWnl3p6B3_0(.dout(w_dff_A_wFRmwx9C7_0),.din(w_dff_A_LWnl3p6B3_0),.clk(gclk));
	jdff dff_A_wFRmwx9C7_0(.dout(w_dff_A_YDV1FGeX0_0),.din(w_dff_A_wFRmwx9C7_0),.clk(gclk));
	jdff dff_A_YDV1FGeX0_0(.dout(w_dff_A_kHcegJFv5_0),.din(w_dff_A_YDV1FGeX0_0),.clk(gclk));
	jdff dff_A_kHcegJFv5_0(.dout(sin7),.din(w_dff_A_kHcegJFv5_0),.clk(gclk));
	jdff dff_A_xitZ0m6h4_2(.dout(w_dff_A_GFtWDc9i0_0),.din(w_dff_A_xitZ0m6h4_2),.clk(gclk));
	jdff dff_A_GFtWDc9i0_0(.dout(w_dff_A_yD4fRJtr7_0),.din(w_dff_A_GFtWDc9i0_0),.clk(gclk));
	jdff dff_A_yD4fRJtr7_0(.dout(w_dff_A_6U0Wy77e6_0),.din(w_dff_A_yD4fRJtr7_0),.clk(gclk));
	jdff dff_A_6U0Wy77e6_0(.dout(w_dff_A_eIl7S7ze6_0),.din(w_dff_A_6U0Wy77e6_0),.clk(gclk));
	jdff dff_A_eIl7S7ze6_0(.dout(w_dff_A_33AONRCr6_0),.din(w_dff_A_eIl7S7ze6_0),.clk(gclk));
	jdff dff_A_33AONRCr6_0(.dout(w_dff_A_rk23tv952_0),.din(w_dff_A_33AONRCr6_0),.clk(gclk));
	jdff dff_A_rk23tv952_0(.dout(w_dff_A_PDy9BJo49_0),.din(w_dff_A_rk23tv952_0),.clk(gclk));
	jdff dff_A_PDy9BJo49_0(.dout(w_dff_A_IrWmIFaR5_0),.din(w_dff_A_PDy9BJo49_0),.clk(gclk));
	jdff dff_A_IrWmIFaR5_0(.dout(w_dff_A_dkMNYgt21_0),.din(w_dff_A_IrWmIFaR5_0),.clk(gclk));
	jdff dff_A_dkMNYgt21_0(.dout(w_dff_A_oj0DwjpZ0_0),.din(w_dff_A_dkMNYgt21_0),.clk(gclk));
	jdff dff_A_oj0DwjpZ0_0(.dout(w_dff_A_PYfLi9Z31_0),.din(w_dff_A_oj0DwjpZ0_0),.clk(gclk));
	jdff dff_A_PYfLi9Z31_0(.dout(w_dff_A_MPxYtxEM6_0),.din(w_dff_A_PYfLi9Z31_0),.clk(gclk));
	jdff dff_A_MPxYtxEM6_0(.dout(w_dff_A_71LUllYi9_0),.din(w_dff_A_MPxYtxEM6_0),.clk(gclk));
	jdff dff_A_71LUllYi9_0(.dout(w_dff_A_4JHIOQn55_0),.din(w_dff_A_71LUllYi9_0),.clk(gclk));
	jdff dff_A_4JHIOQn55_0(.dout(w_dff_A_PBGcaEpT1_0),.din(w_dff_A_4JHIOQn55_0),.clk(gclk));
	jdff dff_A_PBGcaEpT1_0(.dout(w_dff_A_S3P1buBC1_0),.din(w_dff_A_PBGcaEpT1_0),.clk(gclk));
	jdff dff_A_S3P1buBC1_0(.dout(w_dff_A_jaYVMiG42_0),.din(w_dff_A_S3P1buBC1_0),.clk(gclk));
	jdff dff_A_jaYVMiG42_0(.dout(w_dff_A_aXInF5FS1_0),.din(w_dff_A_jaYVMiG42_0),.clk(gclk));
	jdff dff_A_aXInF5FS1_0(.dout(w_dff_A_iY0Av4zl2_0),.din(w_dff_A_aXInF5FS1_0),.clk(gclk));
	jdff dff_A_iY0Av4zl2_0(.dout(w_dff_A_baKc940N6_0),.din(w_dff_A_iY0Av4zl2_0),.clk(gclk));
	jdff dff_A_baKc940N6_0(.dout(w_dff_A_1w93GRRl7_0),.din(w_dff_A_baKc940N6_0),.clk(gclk));
	jdff dff_A_1w93GRRl7_0(.dout(w_dff_A_bilfhlDs8_0),.din(w_dff_A_1w93GRRl7_0),.clk(gclk));
	jdff dff_A_bilfhlDs8_0(.dout(w_dff_A_kgM4MgPf9_0),.din(w_dff_A_bilfhlDs8_0),.clk(gclk));
	jdff dff_A_kgM4MgPf9_0(.dout(w_dff_A_W4XVNCal3_0),.din(w_dff_A_kgM4MgPf9_0),.clk(gclk));
	jdff dff_A_W4XVNCal3_0(.dout(w_dff_A_HOYph2ei1_0),.din(w_dff_A_W4XVNCal3_0),.clk(gclk));
	jdff dff_A_HOYph2ei1_0(.dout(w_dff_A_kkT9ksFJ8_0),.din(w_dff_A_HOYph2ei1_0),.clk(gclk));
	jdff dff_A_kkT9ksFJ8_0(.dout(w_dff_A_7wsIWUxq1_0),.din(w_dff_A_kkT9ksFJ8_0),.clk(gclk));
	jdff dff_A_7wsIWUxq1_0(.dout(w_dff_A_ds9s3jEa9_0),.din(w_dff_A_7wsIWUxq1_0),.clk(gclk));
	jdff dff_A_ds9s3jEa9_0(.dout(sin8),.din(w_dff_A_ds9s3jEa9_0),.clk(gclk));
	jdff dff_A_8Yxnvs8b7_2(.dout(w_dff_A_SYPWSNcc7_0),.din(w_dff_A_8Yxnvs8b7_2),.clk(gclk));
	jdff dff_A_SYPWSNcc7_0(.dout(w_dff_A_mFPo1r7P1_0),.din(w_dff_A_SYPWSNcc7_0),.clk(gclk));
	jdff dff_A_mFPo1r7P1_0(.dout(w_dff_A_2qRNLAHc7_0),.din(w_dff_A_mFPo1r7P1_0),.clk(gclk));
	jdff dff_A_2qRNLAHc7_0(.dout(w_dff_A_0TrraRCu0_0),.din(w_dff_A_2qRNLAHc7_0),.clk(gclk));
	jdff dff_A_0TrraRCu0_0(.dout(w_dff_A_DNxIYxTd3_0),.din(w_dff_A_0TrraRCu0_0),.clk(gclk));
	jdff dff_A_DNxIYxTd3_0(.dout(w_dff_A_o9SgQY2c2_0),.din(w_dff_A_DNxIYxTd3_0),.clk(gclk));
	jdff dff_A_o9SgQY2c2_0(.dout(w_dff_A_SdQ2osBz4_0),.din(w_dff_A_o9SgQY2c2_0),.clk(gclk));
	jdff dff_A_SdQ2osBz4_0(.dout(w_dff_A_ormlNuEr7_0),.din(w_dff_A_SdQ2osBz4_0),.clk(gclk));
	jdff dff_A_ormlNuEr7_0(.dout(w_dff_A_y88nNxrE7_0),.din(w_dff_A_ormlNuEr7_0),.clk(gclk));
	jdff dff_A_y88nNxrE7_0(.dout(w_dff_A_bJsBhGGJ6_0),.din(w_dff_A_y88nNxrE7_0),.clk(gclk));
	jdff dff_A_bJsBhGGJ6_0(.dout(w_dff_A_gsNmYIGd5_0),.din(w_dff_A_bJsBhGGJ6_0),.clk(gclk));
	jdff dff_A_gsNmYIGd5_0(.dout(w_dff_A_307EDnhC9_0),.din(w_dff_A_gsNmYIGd5_0),.clk(gclk));
	jdff dff_A_307EDnhC9_0(.dout(w_dff_A_ruBncPID5_0),.din(w_dff_A_307EDnhC9_0),.clk(gclk));
	jdff dff_A_ruBncPID5_0(.dout(w_dff_A_SuvKsSB52_0),.din(w_dff_A_ruBncPID5_0),.clk(gclk));
	jdff dff_A_SuvKsSB52_0(.dout(w_dff_A_dy3ZYaHg3_0),.din(w_dff_A_SuvKsSB52_0),.clk(gclk));
	jdff dff_A_dy3ZYaHg3_0(.dout(w_dff_A_h3PoJ9bF4_0),.din(w_dff_A_dy3ZYaHg3_0),.clk(gclk));
	jdff dff_A_h3PoJ9bF4_0(.dout(w_dff_A_moWmkxYx5_0),.din(w_dff_A_h3PoJ9bF4_0),.clk(gclk));
	jdff dff_A_moWmkxYx5_0(.dout(w_dff_A_3AYTVXA91_0),.din(w_dff_A_moWmkxYx5_0),.clk(gclk));
	jdff dff_A_3AYTVXA91_0(.dout(w_dff_A_KQIyPtLu6_0),.din(w_dff_A_3AYTVXA91_0),.clk(gclk));
	jdff dff_A_KQIyPtLu6_0(.dout(w_dff_A_WOFOicfO2_0),.din(w_dff_A_KQIyPtLu6_0),.clk(gclk));
	jdff dff_A_WOFOicfO2_0(.dout(w_dff_A_3FiKsycw7_0),.din(w_dff_A_WOFOicfO2_0),.clk(gclk));
	jdff dff_A_3FiKsycw7_0(.dout(w_dff_A_2K98D7ug1_0),.din(w_dff_A_3FiKsycw7_0),.clk(gclk));
	jdff dff_A_2K98D7ug1_0(.dout(w_dff_A_bX9MNSnE5_0),.din(w_dff_A_2K98D7ug1_0),.clk(gclk));
	jdff dff_A_bX9MNSnE5_0(.dout(w_dff_A_Dz8B5NhD2_0),.din(w_dff_A_bX9MNSnE5_0),.clk(gclk));
	jdff dff_A_Dz8B5NhD2_0(.dout(w_dff_A_yfk4EEVA6_0),.din(w_dff_A_Dz8B5NhD2_0),.clk(gclk));
	jdff dff_A_yfk4EEVA6_0(.dout(w_dff_A_dWWTNci52_0),.din(w_dff_A_yfk4EEVA6_0),.clk(gclk));
	jdff dff_A_dWWTNci52_0(.dout(sin9),.din(w_dff_A_dWWTNci52_0),.clk(gclk));
	jdff dff_A_xTdiVglx2_2(.dout(w_dff_A_iKz2u3Ft2_0),.din(w_dff_A_xTdiVglx2_2),.clk(gclk));
	jdff dff_A_iKz2u3Ft2_0(.dout(w_dff_A_Kv10FGAn7_0),.din(w_dff_A_iKz2u3Ft2_0),.clk(gclk));
	jdff dff_A_Kv10FGAn7_0(.dout(w_dff_A_MdLREMMe9_0),.din(w_dff_A_Kv10FGAn7_0),.clk(gclk));
	jdff dff_A_MdLREMMe9_0(.dout(w_dff_A_ynVVe63h9_0),.din(w_dff_A_MdLREMMe9_0),.clk(gclk));
	jdff dff_A_ynVVe63h9_0(.dout(w_dff_A_c0lGk08l2_0),.din(w_dff_A_ynVVe63h9_0),.clk(gclk));
	jdff dff_A_c0lGk08l2_0(.dout(w_dff_A_4VhsE6I25_0),.din(w_dff_A_c0lGk08l2_0),.clk(gclk));
	jdff dff_A_4VhsE6I25_0(.dout(w_dff_A_bz8fAUZd0_0),.din(w_dff_A_4VhsE6I25_0),.clk(gclk));
	jdff dff_A_bz8fAUZd0_0(.dout(w_dff_A_PXFejuCE3_0),.din(w_dff_A_bz8fAUZd0_0),.clk(gclk));
	jdff dff_A_PXFejuCE3_0(.dout(w_dff_A_LpZgHsik2_0),.din(w_dff_A_PXFejuCE3_0),.clk(gclk));
	jdff dff_A_LpZgHsik2_0(.dout(w_dff_A_h4NgCVKe9_0),.din(w_dff_A_LpZgHsik2_0),.clk(gclk));
	jdff dff_A_h4NgCVKe9_0(.dout(w_dff_A_oSsmJyKB3_0),.din(w_dff_A_h4NgCVKe9_0),.clk(gclk));
	jdff dff_A_oSsmJyKB3_0(.dout(w_dff_A_AOWMjE2N9_0),.din(w_dff_A_oSsmJyKB3_0),.clk(gclk));
	jdff dff_A_AOWMjE2N9_0(.dout(w_dff_A_eypCkUHH9_0),.din(w_dff_A_AOWMjE2N9_0),.clk(gclk));
	jdff dff_A_eypCkUHH9_0(.dout(w_dff_A_4tRQtxpw5_0),.din(w_dff_A_eypCkUHH9_0),.clk(gclk));
	jdff dff_A_4tRQtxpw5_0(.dout(w_dff_A_eRIEMAlA4_0),.din(w_dff_A_4tRQtxpw5_0),.clk(gclk));
	jdff dff_A_eRIEMAlA4_0(.dout(w_dff_A_k8ncxhei8_0),.din(w_dff_A_eRIEMAlA4_0),.clk(gclk));
	jdff dff_A_k8ncxhei8_0(.dout(w_dff_A_1WFopbwc6_0),.din(w_dff_A_k8ncxhei8_0),.clk(gclk));
	jdff dff_A_1WFopbwc6_0(.dout(w_dff_A_Urc2OIlf8_0),.din(w_dff_A_1WFopbwc6_0),.clk(gclk));
	jdff dff_A_Urc2OIlf8_0(.dout(w_dff_A_rrE04nif2_0),.din(w_dff_A_Urc2OIlf8_0),.clk(gclk));
	jdff dff_A_rrE04nif2_0(.dout(w_dff_A_8WsMtF2e0_0),.din(w_dff_A_rrE04nif2_0),.clk(gclk));
	jdff dff_A_8WsMtF2e0_0(.dout(w_dff_A_dqTM58VY9_0),.din(w_dff_A_8WsMtF2e0_0),.clk(gclk));
	jdff dff_A_dqTM58VY9_0(.dout(w_dff_A_jBCqwqHM5_0),.din(w_dff_A_dqTM58VY9_0),.clk(gclk));
	jdff dff_A_jBCqwqHM5_0(.dout(w_dff_A_p10qzOdw2_0),.din(w_dff_A_jBCqwqHM5_0),.clk(gclk));
	jdff dff_A_p10qzOdw2_0(.dout(w_dff_A_kZdX2cu59_0),.din(w_dff_A_p10qzOdw2_0),.clk(gclk));
	jdff dff_A_kZdX2cu59_0(.dout(sin10),.din(w_dff_A_kZdX2cu59_0),.clk(gclk));
	jdff dff_A_aayeK3ua3_2(.dout(w_dff_A_VGdSfmU19_0),.din(w_dff_A_aayeK3ua3_2),.clk(gclk));
	jdff dff_A_VGdSfmU19_0(.dout(w_dff_A_V5ASmAJW4_0),.din(w_dff_A_VGdSfmU19_0),.clk(gclk));
	jdff dff_A_V5ASmAJW4_0(.dout(w_dff_A_G7f3wmJt0_0),.din(w_dff_A_V5ASmAJW4_0),.clk(gclk));
	jdff dff_A_G7f3wmJt0_0(.dout(w_dff_A_jtyFGDub8_0),.din(w_dff_A_G7f3wmJt0_0),.clk(gclk));
	jdff dff_A_jtyFGDub8_0(.dout(w_dff_A_f84gTufo3_0),.din(w_dff_A_jtyFGDub8_0),.clk(gclk));
	jdff dff_A_f84gTufo3_0(.dout(w_dff_A_75J3istD6_0),.din(w_dff_A_f84gTufo3_0),.clk(gclk));
	jdff dff_A_75J3istD6_0(.dout(w_dff_A_zZaK0t8K5_0),.din(w_dff_A_75J3istD6_0),.clk(gclk));
	jdff dff_A_zZaK0t8K5_0(.dout(w_dff_A_cc09lsfE2_0),.din(w_dff_A_zZaK0t8K5_0),.clk(gclk));
	jdff dff_A_cc09lsfE2_0(.dout(w_dff_A_Cm7P6Bt25_0),.din(w_dff_A_cc09lsfE2_0),.clk(gclk));
	jdff dff_A_Cm7P6Bt25_0(.dout(w_dff_A_O2tfOzqU8_0),.din(w_dff_A_Cm7P6Bt25_0),.clk(gclk));
	jdff dff_A_O2tfOzqU8_0(.dout(w_dff_A_qFyzp0X27_0),.din(w_dff_A_O2tfOzqU8_0),.clk(gclk));
	jdff dff_A_qFyzp0X27_0(.dout(w_dff_A_zoeSuDYo6_0),.din(w_dff_A_qFyzp0X27_0),.clk(gclk));
	jdff dff_A_zoeSuDYo6_0(.dout(w_dff_A_vYCuIY6O1_0),.din(w_dff_A_zoeSuDYo6_0),.clk(gclk));
	jdff dff_A_vYCuIY6O1_0(.dout(w_dff_A_qvYGC0N36_0),.din(w_dff_A_vYCuIY6O1_0),.clk(gclk));
	jdff dff_A_qvYGC0N36_0(.dout(w_dff_A_IHTE9jDe2_0),.din(w_dff_A_qvYGC0N36_0),.clk(gclk));
	jdff dff_A_IHTE9jDe2_0(.dout(w_dff_A_HTxnzyPQ0_0),.din(w_dff_A_IHTE9jDe2_0),.clk(gclk));
	jdff dff_A_HTxnzyPQ0_0(.dout(w_dff_A_eJSGrcMc5_0),.din(w_dff_A_HTxnzyPQ0_0),.clk(gclk));
	jdff dff_A_eJSGrcMc5_0(.dout(w_dff_A_IlR0jRwe6_0),.din(w_dff_A_eJSGrcMc5_0),.clk(gclk));
	jdff dff_A_IlR0jRwe6_0(.dout(w_dff_A_rEIHsrsR0_0),.din(w_dff_A_IlR0jRwe6_0),.clk(gclk));
	jdff dff_A_rEIHsrsR0_0(.dout(w_dff_A_SLBpBbuv5_0),.din(w_dff_A_rEIHsrsR0_0),.clk(gclk));
	jdff dff_A_SLBpBbuv5_0(.dout(w_dff_A_2Pm6Yf1P8_0),.din(w_dff_A_SLBpBbuv5_0),.clk(gclk));
	jdff dff_A_2Pm6Yf1P8_0(.dout(w_dff_A_iRJl67vO2_0),.din(w_dff_A_2Pm6Yf1P8_0),.clk(gclk));
	jdff dff_A_iRJl67vO2_0(.dout(sin11),.din(w_dff_A_iRJl67vO2_0),.clk(gclk));
	jdff dff_A_AXUFYtJ77_2(.dout(w_dff_A_5TAVS12D0_0),.din(w_dff_A_AXUFYtJ77_2),.clk(gclk));
	jdff dff_A_5TAVS12D0_0(.dout(w_dff_A_vLnUZfVP7_0),.din(w_dff_A_5TAVS12D0_0),.clk(gclk));
	jdff dff_A_vLnUZfVP7_0(.dout(w_dff_A_Kqhxnf8I0_0),.din(w_dff_A_vLnUZfVP7_0),.clk(gclk));
	jdff dff_A_Kqhxnf8I0_0(.dout(w_dff_A_uF89uJ3j4_0),.din(w_dff_A_Kqhxnf8I0_0),.clk(gclk));
	jdff dff_A_uF89uJ3j4_0(.dout(w_dff_A_3bidzuuM6_0),.din(w_dff_A_uF89uJ3j4_0),.clk(gclk));
	jdff dff_A_3bidzuuM6_0(.dout(w_dff_A_Pp8SQXoO2_0),.din(w_dff_A_3bidzuuM6_0),.clk(gclk));
	jdff dff_A_Pp8SQXoO2_0(.dout(w_dff_A_MFRpCeGw4_0),.din(w_dff_A_Pp8SQXoO2_0),.clk(gclk));
	jdff dff_A_MFRpCeGw4_0(.dout(w_dff_A_3IOEKufs7_0),.din(w_dff_A_MFRpCeGw4_0),.clk(gclk));
	jdff dff_A_3IOEKufs7_0(.dout(w_dff_A_R0rBZZB28_0),.din(w_dff_A_3IOEKufs7_0),.clk(gclk));
	jdff dff_A_R0rBZZB28_0(.dout(w_dff_A_16JrRSM28_0),.din(w_dff_A_R0rBZZB28_0),.clk(gclk));
	jdff dff_A_16JrRSM28_0(.dout(w_dff_A_GngooLNm4_0),.din(w_dff_A_16JrRSM28_0),.clk(gclk));
	jdff dff_A_GngooLNm4_0(.dout(w_dff_A_n1YSv8a61_0),.din(w_dff_A_GngooLNm4_0),.clk(gclk));
	jdff dff_A_n1YSv8a61_0(.dout(w_dff_A_jdCWc5VP2_0),.din(w_dff_A_n1YSv8a61_0),.clk(gclk));
	jdff dff_A_jdCWc5VP2_0(.dout(w_dff_A_1T4GIvtJ0_0),.din(w_dff_A_jdCWc5VP2_0),.clk(gclk));
	jdff dff_A_1T4GIvtJ0_0(.dout(w_dff_A_Ti15zLwd1_0),.din(w_dff_A_1T4GIvtJ0_0),.clk(gclk));
	jdff dff_A_Ti15zLwd1_0(.dout(w_dff_A_RgMAxGqo5_0),.din(w_dff_A_Ti15zLwd1_0),.clk(gclk));
	jdff dff_A_RgMAxGqo5_0(.dout(w_dff_A_BEXiJ5Yu3_0),.din(w_dff_A_RgMAxGqo5_0),.clk(gclk));
	jdff dff_A_BEXiJ5Yu3_0(.dout(w_dff_A_7DylCnW46_0),.din(w_dff_A_BEXiJ5Yu3_0),.clk(gclk));
	jdff dff_A_7DylCnW46_0(.dout(w_dff_A_ziewSLq43_0),.din(w_dff_A_7DylCnW46_0),.clk(gclk));
	jdff dff_A_ziewSLq43_0(.dout(w_dff_A_eolJeCl28_0),.din(w_dff_A_ziewSLq43_0),.clk(gclk));
	jdff dff_A_eolJeCl28_0(.dout(sin12),.din(w_dff_A_eolJeCl28_0),.clk(gclk));
	jdff dff_A_i53FbZmW9_2(.dout(w_dff_A_hVj1eVRn2_0),.din(w_dff_A_i53FbZmW9_2),.clk(gclk));
	jdff dff_A_hVj1eVRn2_0(.dout(w_dff_A_czrKWigV5_0),.din(w_dff_A_hVj1eVRn2_0),.clk(gclk));
	jdff dff_A_czrKWigV5_0(.dout(w_dff_A_OguOl2FX5_0),.din(w_dff_A_czrKWigV5_0),.clk(gclk));
	jdff dff_A_OguOl2FX5_0(.dout(w_dff_A_NBsStWDP9_0),.din(w_dff_A_OguOl2FX5_0),.clk(gclk));
	jdff dff_A_NBsStWDP9_0(.dout(w_dff_A_0NaOZ1y67_0),.din(w_dff_A_NBsStWDP9_0),.clk(gclk));
	jdff dff_A_0NaOZ1y67_0(.dout(w_dff_A_AfnOP99w3_0),.din(w_dff_A_0NaOZ1y67_0),.clk(gclk));
	jdff dff_A_AfnOP99w3_0(.dout(w_dff_A_AwtUWFMI1_0),.din(w_dff_A_AfnOP99w3_0),.clk(gclk));
	jdff dff_A_AwtUWFMI1_0(.dout(w_dff_A_M5tqbj6J2_0),.din(w_dff_A_AwtUWFMI1_0),.clk(gclk));
	jdff dff_A_M5tqbj6J2_0(.dout(w_dff_A_GiTQ42wU7_0),.din(w_dff_A_M5tqbj6J2_0),.clk(gclk));
	jdff dff_A_GiTQ42wU7_0(.dout(w_dff_A_aW7cCnZQ8_0),.din(w_dff_A_GiTQ42wU7_0),.clk(gclk));
	jdff dff_A_aW7cCnZQ8_0(.dout(w_dff_A_fVmUA1oC1_0),.din(w_dff_A_aW7cCnZQ8_0),.clk(gclk));
	jdff dff_A_fVmUA1oC1_0(.dout(w_dff_A_oeUyyrxc7_0),.din(w_dff_A_fVmUA1oC1_0),.clk(gclk));
	jdff dff_A_oeUyyrxc7_0(.dout(w_dff_A_ThJfWili0_0),.din(w_dff_A_oeUyyrxc7_0),.clk(gclk));
	jdff dff_A_ThJfWili0_0(.dout(w_dff_A_S99gi9db1_0),.din(w_dff_A_ThJfWili0_0),.clk(gclk));
	jdff dff_A_S99gi9db1_0(.dout(w_dff_A_HbdVtext7_0),.din(w_dff_A_S99gi9db1_0),.clk(gclk));
	jdff dff_A_HbdVtext7_0(.dout(w_dff_A_XnyY5NX66_0),.din(w_dff_A_HbdVtext7_0),.clk(gclk));
	jdff dff_A_XnyY5NX66_0(.dout(w_dff_A_f9nbxHLb0_0),.din(w_dff_A_XnyY5NX66_0),.clk(gclk));
	jdff dff_A_f9nbxHLb0_0(.dout(w_dff_A_9hSL2wJF7_0),.din(w_dff_A_f9nbxHLb0_0),.clk(gclk));
	jdff dff_A_9hSL2wJF7_0(.dout(sin13),.din(w_dff_A_9hSL2wJF7_0),.clk(gclk));
	jdff dff_A_MRzbRLbX5_2(.dout(w_dff_A_bmcMeNgS4_0),.din(w_dff_A_MRzbRLbX5_2),.clk(gclk));
	jdff dff_A_bmcMeNgS4_0(.dout(w_dff_A_wDSIqWH43_0),.din(w_dff_A_bmcMeNgS4_0),.clk(gclk));
	jdff dff_A_wDSIqWH43_0(.dout(w_dff_A_mgBB9fcK0_0),.din(w_dff_A_wDSIqWH43_0),.clk(gclk));
	jdff dff_A_mgBB9fcK0_0(.dout(w_dff_A_CVdXtpmj5_0),.din(w_dff_A_mgBB9fcK0_0),.clk(gclk));
	jdff dff_A_CVdXtpmj5_0(.dout(w_dff_A_wkRbPaiG1_0),.din(w_dff_A_CVdXtpmj5_0),.clk(gclk));
	jdff dff_A_wkRbPaiG1_0(.dout(w_dff_A_79qiRzi08_0),.din(w_dff_A_wkRbPaiG1_0),.clk(gclk));
	jdff dff_A_79qiRzi08_0(.dout(w_dff_A_yCs0SDH25_0),.din(w_dff_A_79qiRzi08_0),.clk(gclk));
	jdff dff_A_yCs0SDH25_0(.dout(w_dff_A_Tbr0acDy0_0),.din(w_dff_A_yCs0SDH25_0),.clk(gclk));
	jdff dff_A_Tbr0acDy0_0(.dout(w_dff_A_JLox2jbS0_0),.din(w_dff_A_Tbr0acDy0_0),.clk(gclk));
	jdff dff_A_JLox2jbS0_0(.dout(w_dff_A_K8h2N7414_0),.din(w_dff_A_JLox2jbS0_0),.clk(gclk));
	jdff dff_A_K8h2N7414_0(.dout(w_dff_A_aOa6z9ue3_0),.din(w_dff_A_K8h2N7414_0),.clk(gclk));
	jdff dff_A_aOa6z9ue3_0(.dout(w_dff_A_P17RISnR3_0),.din(w_dff_A_aOa6z9ue3_0),.clk(gclk));
	jdff dff_A_P17RISnR3_0(.dout(w_dff_A_pW5IAoT87_0),.din(w_dff_A_P17RISnR3_0),.clk(gclk));
	jdff dff_A_pW5IAoT87_0(.dout(w_dff_A_bBrHfNIo9_0),.din(w_dff_A_pW5IAoT87_0),.clk(gclk));
	jdff dff_A_bBrHfNIo9_0(.dout(w_dff_A_JrSD9GXH9_0),.din(w_dff_A_bBrHfNIo9_0),.clk(gclk));
	jdff dff_A_JrSD9GXH9_0(.dout(w_dff_A_lnGqSLfY2_0),.din(w_dff_A_JrSD9GXH9_0),.clk(gclk));
	jdff dff_A_lnGqSLfY2_0(.dout(sin14),.din(w_dff_A_lnGqSLfY2_0),.clk(gclk));
	jdff dff_A_MetX8NB96_2(.dout(w_dff_A_kFCIRYxd1_0),.din(w_dff_A_MetX8NB96_2),.clk(gclk));
	jdff dff_A_kFCIRYxd1_0(.dout(w_dff_A_6Y8hv5bq5_0),.din(w_dff_A_kFCIRYxd1_0),.clk(gclk));
	jdff dff_A_6Y8hv5bq5_0(.dout(w_dff_A_ZQME5H1p6_0),.din(w_dff_A_6Y8hv5bq5_0),.clk(gclk));
	jdff dff_A_ZQME5H1p6_0(.dout(w_dff_A_qgc6oGFr0_0),.din(w_dff_A_ZQME5H1p6_0),.clk(gclk));
	jdff dff_A_qgc6oGFr0_0(.dout(w_dff_A_bPL7G4gV4_0),.din(w_dff_A_qgc6oGFr0_0),.clk(gclk));
	jdff dff_A_bPL7G4gV4_0(.dout(w_dff_A_7xpwiQHR9_0),.din(w_dff_A_bPL7G4gV4_0),.clk(gclk));
	jdff dff_A_7xpwiQHR9_0(.dout(w_dff_A_5GHgZTa38_0),.din(w_dff_A_7xpwiQHR9_0),.clk(gclk));
	jdff dff_A_5GHgZTa38_0(.dout(w_dff_A_rJ46syzs8_0),.din(w_dff_A_5GHgZTa38_0),.clk(gclk));
	jdff dff_A_rJ46syzs8_0(.dout(w_dff_A_OTlabvXC5_0),.din(w_dff_A_rJ46syzs8_0),.clk(gclk));
	jdff dff_A_OTlabvXC5_0(.dout(w_dff_A_1I877Ghn7_0),.din(w_dff_A_OTlabvXC5_0),.clk(gclk));
	jdff dff_A_1I877Ghn7_0(.dout(w_dff_A_vzSImIZ66_0),.din(w_dff_A_1I877Ghn7_0),.clk(gclk));
	jdff dff_A_vzSImIZ66_0(.dout(w_dff_A_T2c3bCeS4_0),.din(w_dff_A_vzSImIZ66_0),.clk(gclk));
	jdff dff_A_T2c3bCeS4_0(.dout(w_dff_A_HbkmqjKA8_0),.din(w_dff_A_T2c3bCeS4_0),.clk(gclk));
	jdff dff_A_HbkmqjKA8_0(.dout(w_dff_A_XEFqRjOB6_0),.din(w_dff_A_HbkmqjKA8_0),.clk(gclk));
	jdff dff_A_XEFqRjOB6_0(.dout(sin15),.din(w_dff_A_XEFqRjOB6_0),.clk(gclk));
	jdff dff_A_HU6Y95fG4_2(.dout(w_dff_A_fkSelirA5_0),.din(w_dff_A_HU6Y95fG4_2),.clk(gclk));
	jdff dff_A_fkSelirA5_0(.dout(w_dff_A_s9XgZCGz4_0),.din(w_dff_A_fkSelirA5_0),.clk(gclk));
	jdff dff_A_s9XgZCGz4_0(.dout(w_dff_A_ldn8tt7l8_0),.din(w_dff_A_s9XgZCGz4_0),.clk(gclk));
	jdff dff_A_ldn8tt7l8_0(.dout(w_dff_A_tooFhoxr9_0),.din(w_dff_A_ldn8tt7l8_0),.clk(gclk));
	jdff dff_A_tooFhoxr9_0(.dout(w_dff_A_dC4MAl1s5_0),.din(w_dff_A_tooFhoxr9_0),.clk(gclk));
	jdff dff_A_dC4MAl1s5_0(.dout(w_dff_A_FmpBvojb2_0),.din(w_dff_A_dC4MAl1s5_0),.clk(gclk));
	jdff dff_A_FmpBvojb2_0(.dout(w_dff_A_UAdGPHSE4_0),.din(w_dff_A_FmpBvojb2_0),.clk(gclk));
	jdff dff_A_UAdGPHSE4_0(.dout(w_dff_A_TKRQg00C4_0),.din(w_dff_A_UAdGPHSE4_0),.clk(gclk));
	jdff dff_A_TKRQg00C4_0(.dout(w_dff_A_tPk8mCWW7_0),.din(w_dff_A_TKRQg00C4_0),.clk(gclk));
	jdff dff_A_tPk8mCWW7_0(.dout(w_dff_A_FeGbU0Yv3_0),.din(w_dff_A_tPk8mCWW7_0),.clk(gclk));
	jdff dff_A_FeGbU0Yv3_0(.dout(w_dff_A_fhuCuywo1_0),.din(w_dff_A_FeGbU0Yv3_0),.clk(gclk));
	jdff dff_A_fhuCuywo1_0(.dout(sin16),.din(w_dff_A_fhuCuywo1_0),.clk(gclk));
	jdff dff_A_GPqiqml02_2(.dout(w_dff_A_yfQkah866_0),.din(w_dff_A_GPqiqml02_2),.clk(gclk));
	jdff dff_A_yfQkah866_0(.dout(w_dff_A_bUPQneH97_0),.din(w_dff_A_yfQkah866_0),.clk(gclk));
	jdff dff_A_bUPQneH97_0(.dout(w_dff_A_KFuKxUiF3_0),.din(w_dff_A_bUPQneH97_0),.clk(gclk));
	jdff dff_A_KFuKxUiF3_0(.dout(w_dff_A_XiktjTX59_0),.din(w_dff_A_KFuKxUiF3_0),.clk(gclk));
	jdff dff_A_XiktjTX59_0(.dout(w_dff_A_8MC6z9Bx5_0),.din(w_dff_A_XiktjTX59_0),.clk(gclk));
	jdff dff_A_8MC6z9Bx5_0(.dout(w_dff_A_BR5L0SJE6_0),.din(w_dff_A_8MC6z9Bx5_0),.clk(gclk));
	jdff dff_A_BR5L0SJE6_0(.dout(w_dff_A_RyEZ8Cq11_0),.din(w_dff_A_BR5L0SJE6_0),.clk(gclk));
	jdff dff_A_RyEZ8Cq11_0(.dout(w_dff_A_VKAVuqlZ6_0),.din(w_dff_A_RyEZ8Cq11_0),.clk(gclk));
	jdff dff_A_VKAVuqlZ6_0(.dout(w_dff_A_MLj3FGzh5_0),.din(w_dff_A_VKAVuqlZ6_0),.clk(gclk));
	jdff dff_A_MLj3FGzh5_0(.dout(sin17),.din(w_dff_A_MLj3FGzh5_0),.clk(gclk));
	jdff dff_A_1nMlhPpu8_2(.dout(w_dff_A_w7E0o7ab6_0),.din(w_dff_A_1nMlhPpu8_2),.clk(gclk));
	jdff dff_A_w7E0o7ab6_0(.dout(w_dff_A_V4HYM5qa8_0),.din(w_dff_A_w7E0o7ab6_0),.clk(gclk));
	jdff dff_A_V4HYM5qa8_0(.dout(w_dff_A_Zk6ZIW6G3_0),.din(w_dff_A_V4HYM5qa8_0),.clk(gclk));
	jdff dff_A_Zk6ZIW6G3_0(.dout(w_dff_A_Nng9uJFY2_0),.din(w_dff_A_Zk6ZIW6G3_0),.clk(gclk));
	jdff dff_A_Nng9uJFY2_0(.dout(w_dff_A_svTt3Rct3_0),.din(w_dff_A_Nng9uJFY2_0),.clk(gclk));
	jdff dff_A_svTt3Rct3_0(.dout(w_dff_A_6A34fKVP7_0),.din(w_dff_A_svTt3Rct3_0),.clk(gclk));
	jdff dff_A_6A34fKVP7_0(.dout(w_dff_A_5DqkBfTU6_0),.din(w_dff_A_6A34fKVP7_0),.clk(gclk));
	jdff dff_A_5DqkBfTU6_0(.dout(sin18),.din(w_dff_A_5DqkBfTU6_0),.clk(gclk));
	jdff dff_A_AlCqYWkD8_2(.dout(w_dff_A_gNv4B3hs4_0),.din(w_dff_A_AlCqYWkD8_2),.clk(gclk));
	jdff dff_A_gNv4B3hs4_0(.dout(w_dff_A_zJu0IT1w5_0),.din(w_dff_A_gNv4B3hs4_0),.clk(gclk));
	jdff dff_A_zJu0IT1w5_0(.dout(w_dff_A_M6b6oqqB4_0),.din(w_dff_A_zJu0IT1w5_0),.clk(gclk));
	jdff dff_A_M6b6oqqB4_0(.dout(w_dff_A_OJtixmIZ4_0),.din(w_dff_A_M6b6oqqB4_0),.clk(gclk));
	jdff dff_A_OJtixmIZ4_0(.dout(w_dff_A_wcSxKrSD1_0),.din(w_dff_A_OJtixmIZ4_0),.clk(gclk));
	jdff dff_A_wcSxKrSD1_0(.dout(sin19),.din(w_dff_A_wcSxKrSD1_0),.clk(gclk));
	jdff dff_A_QgvCi3b43_2(.dout(w_dff_A_nRfPDqbs5_0),.din(w_dff_A_QgvCi3b43_2),.clk(gclk));
	jdff dff_A_nRfPDqbs5_0(.dout(w_dff_A_vzTX9Gql9_0),.din(w_dff_A_nRfPDqbs5_0),.clk(gclk));
	jdff dff_A_vzTX9Gql9_0(.dout(w_dff_A_eEF03FKE6_0),.din(w_dff_A_vzTX9Gql9_0),.clk(gclk));
	jdff dff_A_eEF03FKE6_0(.dout(w_dff_A_S1RJz5WQ3_0),.din(w_dff_A_eEF03FKE6_0),.clk(gclk));
	jdff dff_A_S1RJz5WQ3_0(.dout(sin20),.din(w_dff_A_S1RJz5WQ3_0),.clk(gclk));
	jdff dff_A_khtMLhmf2_2(.dout(w_dff_A_ufMNppQ99_0),.din(w_dff_A_khtMLhmf2_2),.clk(gclk));
	jdff dff_A_ufMNppQ99_0(.dout(w_dff_A_JKLHkgMy0_0),.din(w_dff_A_ufMNppQ99_0),.clk(gclk));
	jdff dff_A_JKLHkgMy0_0(.dout(w_dff_A_WEvisCtm5_0),.din(w_dff_A_JKLHkgMy0_0),.clk(gclk));
	jdff dff_A_WEvisCtm5_0(.dout(sin21),.din(w_dff_A_WEvisCtm5_0),.clk(gclk));
	jdff dff_A_d1DL4wzM4_2(.dout(w_dff_A_6D1oDIwG4_0),.din(w_dff_A_d1DL4wzM4_2),.clk(gclk));
	jdff dff_A_6D1oDIwG4_0(.dout(w_dff_A_xOJ1iUnI3_0),.din(w_dff_A_6D1oDIwG4_0),.clk(gclk));
	jdff dff_A_xOJ1iUnI3_0(.dout(sin22),.din(w_dff_A_xOJ1iUnI3_0),.clk(gclk));
endmodule

