/*
rf_c7552:
	jxor: 228
	jspl: 345
	jspl3: 346
	jnot: 270
	jdff: 4170
	jor: 395
	jand: 513

Summary:
	jxor: 228
	jspl: 345
	jspl3: 346
	jnot: 270
	jdff: 4170
	jor: 395
	jand: 513

The maximum logic level gap of any gate:
	rf_c7552: 21
*/

module rf_c7552(gclk, G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526, G4528, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399);
	input gclk;
	input G1;
	input G5;
	input G9;
	input G12;
	input G15;
	input G18;
	input G23;
	input G26;
	input G29;
	input G32;
	input G35;
	input G38;
	input G41;
	input G44;
	input G47;
	input G50;
	input G53;
	input G54;
	input G55;
	input G56;
	input G57;
	input G58;
	input G59;
	input G60;
	input G61;
	input G62;
	input G63;
	input G64;
	input G65;
	input G66;
	input G69;
	input G70;
	input G73;
	input G74;
	input G75;
	input G76;
	input G77;
	input G78;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G84;
	input G85;
	input G86;
	input G87;
	input G88;
	input G89;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G110;
	input G111;
	input G112;
	input G113;
	input G114;
	input G115;
	input G118;
	input G121;
	input G124;
	input G127;
	input G130;
	input G133;
	input G134;
	input G135;
	input G138;
	input G141;
	input G144;
	input G147;
	input G150;
	input G151;
	input G152;
	input G153;
	input G154;
	input G155;
	input G156;
	input G157;
	input G158;
	input G159;
	input G160;
	input G161;
	input G162;
	input G163;
	input G164;
	input G165;
	input G166;
	input G167;
	input G168;
	input G169;
	input G170;
	input G171;
	input G172;
	input G173;
	input G174;
	input G175;
	input G176;
	input G177;
	input G178;
	input G179;
	input G180;
	input G181;
	input G182;
	input G183;
	input G184;
	input G185;
	input G186;
	input G187;
	input G188;
	input G189;
	input G190;
	input G191;
	input G192;
	input G193;
	input G194;
	input G195;
	input G196;
	input G197;
	input G198;
	input G199;
	input G200;
	input G201;
	input G202;
	input G203;
	input G204;
	input G205;
	input G206;
	input G207;
	input G208;
	input G209;
	input G210;
	input G211;
	input G212;
	input G213;
	input G214;
	input G215;
	input G216;
	input G217;
	input G218;
	input G219;
	input G220;
	input G221;
	input G222;
	input G223;
	input G224;
	input G225;
	input G226;
	input G227;
	input G228;
	input G229;
	input G230;
	input G231;
	input G232;
	input G233;
	input G234;
	input G235;
	input G236;
	input G237;
	input G238;
	input G239;
	input G240;
	input G339;
	input G1197;
	input G1455;
	input G1459;
	input G1462;
	input G1469;
	input G1480;
	input G1486;
	input G1492;
	input G1496;
	input G2204;
	input G2208;
	input G2211;
	input G2218;
	input G2224;
	input G2230;
	input G2236;
	input G2239;
	input G2247;
	input G2253;
	input G2256;
	input G3698;
	input G3701;
	input G3705;
	input G3711;
	input G3717;
	input G3723;
	input G3729;
	input G3737;
	input G3743;
	input G3749;
	input G4393;
	input G4394;
	input G4400;
	input G4405;
	input G4410;
	input G4415;
	input G4420;
	input G4427;
	input G4432;
	input G4437;
	input G4526;
	input G4528;
	output G2;
	output G3;
	output G450;
	output G448;
	output G444;
	output G442;
	output G440;
	output G438;
	output G496;
	output G494;
	output G492;
	output G490;
	output G488;
	output G486;
	output G484;
	output G482;
	output G480;
	output G560;
	output G542;
	output G558;
	output G556;
	output G554;
	output G552;
	output G550;
	output G548;
	output G546;
	output G544;
	output G540;
	output G538;
	output G536;
	output G534;
	output G532;
	output G530;
	output G528;
	output G526;
	output G524;
	output G279;
	output G436;
	output G478;
	output G522;
	output G402;
	output G404;
	output G406;
	output G408;
	output G410;
	output G432;
	output G446;
	output G284;
	output G286;
	output G289;
	output G292;
	output G341;
	output G281;
	output G453;
	output G278;
	output G373;
	output G246;
	output G258;
	output G264;
	output G270;
	output G388;
	output G391;
	output G394;
	output G397;
	output G376;
	output G379;
	output G382;
	output G385;
	output G412;
	output G414;
	output G416;
	output G249;
	output G295;
	output G324;
	output G252;
	output G276;
	output G310;
	output G313;
	output G316;
	output G319;
	output G327;
	output G330;
	output G333;
	output G336;
	output G418;
	output G273;
	output G298;
	output G301;
	output G304;
	output G307;
	output G344;
	output G422;
	output G469;
	output G419;
	output G471;
	output G359;
	output G362;
	output G365;
	output G368;
	output G347;
	output G350;
	output G353;
	output G356;
	output G321;
	output G338;
	output G370;
	output G399;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n347;
	wire n348;
	wire n349;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1134;
	wire n1136;
	wire n1137;
	wire n1139;
	wire n1140;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1146;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1410;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1417;
	wire n1418;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1429;
	wire n1430;
	wire n1432;
	wire n1433;
	wire n1435;
	wire n1436;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1451;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1477;
	wire n1479;
	wire n1480;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1490;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [2:0] w_G5_0;
	wire [2:0] w_G5_1;
	wire [2:0] w_G15_0;
	wire [2:0] w_G18_0;
	wire [2:0] w_G18_1;
	wire [2:0] w_G18_2;
	wire [2:0] w_G18_3;
	wire [2:0] w_G18_4;
	wire [2:0] w_G18_5;
	wire [2:0] w_G18_6;
	wire [2:0] w_G18_7;
	wire [2:0] w_G18_8;
	wire [2:0] w_G18_9;
	wire [2:0] w_G18_10;
	wire [2:0] w_G18_11;
	wire [2:0] w_G18_12;
	wire [2:0] w_G18_13;
	wire [2:0] w_G18_14;
	wire [2:0] w_G18_15;
	wire [2:0] w_G18_16;
	wire [2:0] w_G18_17;
	wire [2:0] w_G18_18;
	wire [2:0] w_G18_19;
	wire [2:0] w_G18_20;
	wire [2:0] w_G18_21;
	wire [2:0] w_G18_22;
	wire [2:0] w_G18_23;
	wire [2:0] w_G18_24;
	wire [2:0] w_G18_25;
	wire [2:0] w_G18_26;
	wire [2:0] w_G18_27;
	wire [2:0] w_G18_28;
	wire [2:0] w_G18_29;
	wire [2:0] w_G18_30;
	wire [2:0] w_G18_31;
	wire [2:0] w_G18_32;
	wire [2:0] w_G18_33;
	wire [2:0] w_G18_34;
	wire [2:0] w_G18_35;
	wire [2:0] w_G18_36;
	wire [2:0] w_G18_37;
	wire [2:0] w_G18_38;
	wire [2:0] w_G18_39;
	wire [2:0] w_G18_40;
	wire [2:0] w_G18_41;
	wire [2:0] w_G18_42;
	wire [2:0] w_G18_43;
	wire [2:0] w_G18_44;
	wire [2:0] w_G18_45;
	wire [2:0] w_G18_46;
	wire [2:0] w_G18_47;
	wire [2:0] w_G18_48;
	wire [2:0] w_G18_49;
	wire [2:0] w_G18_50;
	wire [2:0] w_G18_51;
	wire [2:0] w_G18_52;
	wire [2:0] w_G18_53;
	wire [2:0] w_G18_54;
	wire [2:0] w_G18_55;
	wire [2:0] w_G18_56;
	wire [2:0] w_G18_57;
	wire [2:0] w_G18_58;
	wire [2:0] w_G38_0;
	wire [2:0] w_G38_1;
	wire [2:0] w_G41_0;
	wire [1:0] w_G69_0;
	wire [1:0] w_G70_0;
	wire [2:0] w_G106_0;
	wire [1:0] w_G106_1;
	wire [1:0] w_G229_0;
	wire [2:0] w_G1455_0;
	wire [1:0] w_G1459_0;
	wire [2:0] w_G1462_0;
	wire [2:0] w_G1469_0;
	wire [1:0] w_G1469_1;
	wire [2:0] w_G1480_0;
	wire [2:0] w_G1486_0;
	wire [2:0] w_G1492_0;
	wire [1:0] w_G1492_1;
	wire [2:0] w_G1496_0;
	wire [2:0] w_G2204_0;
	wire [1:0] w_G2208_0;
	wire [2:0] w_G2211_0;
	wire [2:0] w_G2218_0;
	wire [2:0] w_G2224_0;
	wire [1:0] w_G2224_1;
	wire [2:0] w_G2230_0;
	wire [1:0] w_G2230_1;
	wire [2:0] w_G2236_0;
	wire [1:0] w_G2236_1;
	wire [2:0] w_G2239_0;
	wire [2:0] w_G2247_0;
	wire [2:0] w_G2253_0;
	wire [1:0] w_G2253_1;
	wire [2:0] w_G2256_0;
	wire [1:0] w_G2256_1;
	wire [1:0] w_G3698_0;
	wire [2:0] w_G3701_0;
	wire [1:0] w_G3701_1;
	wire [2:0] w_G3705_0;
	wire [2:0] w_G3705_1;
	wire [1:0] w_G3705_2;
	wire [2:0] w_G3711_0;
	wire [1:0] w_G3711_1;
	wire [2:0] w_G3717_0;
	wire [2:0] w_G3717_1;
	wire [1:0] w_G3717_2;
	wire [2:0] w_G3723_0;
	wire [1:0] w_G3723_1;
	wire [2:0] w_G3729_0;
	wire [1:0] w_G3729_1;
	wire [2:0] w_G3737_0;
	wire [1:0] w_G3737_1;
	wire [2:0] w_G3743_0;
	wire [2:0] w_G3743_1;
	wire [2:0] w_G3749_0;
	wire [1:0] w_G3749_1;
	wire [1:0] w_G4393_0;
	wire [2:0] w_G4394_0;
	wire [1:0] w_G4394_1;
	wire [2:0] w_G4400_0;
	wire [2:0] w_G4405_0;
	wire [2:0] w_G4405_1;
	wire [2:0] w_G4410_0;
	wire [1:0] w_G4410_1;
	wire [2:0] w_G4415_0;
	wire [1:0] w_G4415_1;
	wire [2:0] w_G4420_0;
	wire [1:0] w_G4427_0;
	wire [2:0] w_G4432_0;
	wire [1:0] w_G4432_1;
	wire [2:0] w_G4437_0;
	wire [2:0] w_G4526_0;
	wire [1:0] w_G4526_1;
	wire [2:0] w_G4528_0;
	wire w_G404_0;
	wire G404_fa_;
	wire w_G406_0;
	wire G406_fa_;
	wire w_G408_0;
	wire G408_fa_;
	wire w_G410_0;
	wire G410_fa_;
	wire w_G412_0;
	wire G412_fa_;
	wire w_G414_0;
	wire G414_fa_;
	wire w_G416_0;
	wire G416_fa_;
	wire [1:0] w_n345_0;
	wire [1:0] w_n349_0;
	wire [2:0] w_n353_0;
	wire [2:0] w_n354_0;
	wire [2:0] w_n354_1;
	wire [2:0] w_n355_0;
	wire [2:0] w_n355_1;
	wire [2:0] w_n355_2;
	wire [2:0] w_n355_3;
	wire [2:0] w_n355_4;
	wire [2:0] w_n355_5;
	wire [2:0] w_n355_6;
	wire [2:0] w_n355_7;
	wire [2:0] w_n355_8;
	wire [2:0] w_n355_9;
	wire [2:0] w_n355_10;
	wire [2:0] w_n355_11;
	wire [2:0] w_n355_12;
	wire [2:0] w_n355_13;
	wire [2:0] w_n355_14;
	wire [2:0] w_n355_15;
	wire [2:0] w_n355_16;
	wire [2:0] w_n355_17;
	wire [2:0] w_n355_18;
	wire [2:0] w_n355_19;
	wire [2:0] w_n355_20;
	wire [2:0] w_n355_21;
	wire [2:0] w_n355_22;
	wire [2:0] w_n355_23;
	wire [2:0] w_n355_24;
	wire [2:0] w_n355_25;
	wire [1:0] w_n355_26;
	wire [2:0] w_n356_0;
	wire [1:0] w_n358_0;
	wire [1:0] w_n359_0;
	wire [2:0] w_n362_0;
	wire [1:0] w_n364_0;
	wire [1:0] w_n365_0;
	wire [1:0] w_n366_0;
	wire [1:0] w_n370_0;
	wire [2:0] w_n371_0;
	wire [1:0] w_n371_1;
	wire [2:0] w_n372_0;
	wire [2:0] w_n372_1;
	wire [1:0] w_n376_0;
	wire [2:0] w_n377_0;
	wire [2:0] w_n377_1;
	wire [2:0] w_n379_0;
	wire [1:0] w_n379_1;
	wire [2:0] w_n380_0;
	wire [1:0] w_n385_0;
	wire [2:0] w_n386_0;
	wire [2:0] w_n387_0;
	wire [2:0] w_n387_1;
	wire [2:0] w_n388_0;
	wire [1:0] w_n389_0;
	wire [2:0] w_n390_0;
	wire [1:0] w_n390_1;
	wire [2:0] w_n395_0;
	wire [1:0] w_n400_0;
	wire [2:0] w_n401_0;
	wire [2:0] w_n401_1;
	wire [2:0] w_n402_0;
	wire [1:0] w_n402_1;
	wire [1:0] w_n403_0;
	wire [1:0] w_n404_0;
	wire [2:0] w_n405_0;
	wire [2:0] w_n407_0;
	wire [1:0] w_n408_0;
	wire [1:0] w_n410_0;
	wire [2:0] w_n412_0;
	wire [2:0] w_n413_0;
	wire [1:0] w_n413_1;
	wire [2:0] w_n417_0;
	wire [1:0] w_n419_0;
	wire [2:0] w_n422_0;
	wire [2:0] w_n422_1;
	wire [1:0] w_n427_0;
	wire [2:0] w_n428_0;
	wire [2:0] w_n429_0;
	wire [2:0] w_n429_1;
	wire [1:0] w_n429_2;
	wire [1:0] w_n430_0;
	wire [1:0] w_n434_0;
	wire [2:0] w_n435_0;
	wire [1:0] w_n435_1;
	wire [1:0] w_n436_0;
	wire [1:0] w_n437_0;
	wire [1:0] w_n441_0;
	wire [2:0] w_n442_0;
	wire [1:0] w_n443_0;
	wire [1:0] w_n445_0;
	wire [2:0] w_n446_0;
	wire [1:0] w_n446_1;
	wire [1:0] w_n448_0;
	wire [2:0] w_n449_0;
	wire [2:0] w_n450_0;
	wire [1:0] w_n452_0;
	wire [1:0] w_n454_0;
	wire [1:0] w_n455_0;
	wire [2:0] w_n456_0;
	wire [1:0] w_n457_0;
	wire [2:0] w_n458_0;
	wire [2:0] w_n460_0;
	wire [1:0] w_n461_0;
	wire [2:0] w_n462_0;
	wire [1:0] w_n464_0;
	wire [2:0] w_n465_0;
	wire [1:0] w_n466_0;
	wire [1:0] w_n468_0;
	wire [2:0] w_n469_0;
	wire [1:0] w_n469_1;
	wire [2:0] w_n470_0;
	wire [2:0] w_n471_0;
	wire [1:0] w_n473_0;
	wire [2:0] w_n474_0;
	wire [1:0] w_n474_1;
	wire [2:0] w_n475_0;
	wire [1:0] w_n475_1;
	wire [1:0] w_n477_0;
	wire [1:0] w_n478_0;
	wire [1:0] w_n479_0;
	wire [2:0] w_n480_0;
	wire [1:0] w_n480_1;
	wire [2:0] w_n481_0;
	wire [1:0] w_n482_0;
	wire [1:0] w_n484_0;
	wire [2:0] w_n485_0;
	wire [2:0] w_n486_0;
	wire [1:0] w_n488_0;
	wire [1:0] w_n489_0;
	wire [2:0] w_n490_0;
	wire [2:0] w_n491_0;
	wire [1:0] w_n491_1;
	wire [1:0] w_n493_0;
	wire [1:0] w_n494_0;
	wire [1:0] w_n502_0;
	wire [1:0] w_n503_0;
	wire [1:0] w_n505_0;
	wire [2:0] w_n507_0;
	wire [2:0] w_n507_1;
	wire [1:0] w_n508_0;
	wire [1:0] w_n509_0;
	wire [1:0] w_n510_0;
	wire [1:0] w_n512_0;
	wire [2:0] w_n514_0;
	wire [2:0] w_n516_0;
	wire [1:0] w_n518_0;
	wire [1:0] w_n519_0;
	wire [2:0] w_n520_0;
	wire [1:0] w_n522_0;
	wire [2:0] w_n523_0;
	wire [2:0] w_n524_0;
	wire [2:0] w_n524_1;
	wire [1:0] w_n524_2;
	wire [2:0] w_n525_0;
	wire [1:0] w_n527_0;
	wire [2:0] w_n528_0;
	wire [1:0] w_n528_1;
	wire [1:0] w_n529_0;
	wire [1:0] w_n530_0;
	wire [2:0] w_n531_0;
	wire [1:0] w_n533_0;
	wire [2:0] w_n534_0;
	wire [1:0] w_n534_1;
	wire [2:0] w_n535_0;
	wire [1:0] w_n535_1;
	wire [1:0] w_n536_0;
	wire [1:0] w_n538_0;
	wire [2:0] w_n539_0;
	wire [1:0] w_n539_1;
	wire [2:0] w_n540_0;
	wire [1:0] w_n542_0;
	wire [1:0] w_n549_0;
	wire [1:0] w_n551_0;
	wire [1:0] w_n552_0;
	wire [1:0] w_n553_0;
	wire [2:0] w_n554_0;
	wire [2:0] w_n556_0;
	wire [1:0] w_n557_0;
	wire [2:0] w_n558_0;
	wire [1:0] w_n560_0;
	wire [2:0] w_n562_0;
	wire [1:0] w_n563_0;
	wire [2:0] w_n564_0;
	wire [2:0] w_n565_0;
	wire [2:0] w_n565_1;
	wire [2:0] w_n565_2;
	wire [2:0] w_n565_3;
	wire [2:0] w_n565_4;
	wire [2:0] w_n565_5;
	wire [2:0] w_n565_6;
	wire [2:0] w_n565_7;
	wire [2:0] w_n565_8;
	wire [2:0] w_n565_9;
	wire [1:0] w_n565_10;
	wire [2:0] w_n567_0;
	wire [1:0] w_n567_1;
	wire [2:0] w_n568_0;
	wire [2:0] w_n569_0;
	wire [1:0] w_n570_0;
	wire [2:0] w_n572_0;
	wire [1:0] w_n572_1;
	wire [2:0] w_n573_0;
	wire [1:0] w_n573_1;
	wire [1:0] w_n574_0;
	wire [1:0] w_n575_0;
	wire [2:0] w_n577_0;
	wire [2:0] w_n578_0;
	wire [1:0] w_n578_1;
	wire [2:0] w_n579_0;
	wire [1:0] w_n580_0;
	wire [1:0] w_n581_0;
	wire [2:0] w_n583_0;
	wire [1:0] w_n583_1;
	wire [2:0] w_n584_0;
	wire [1:0] w_n585_0;
	wire [1:0] w_n586_0;
	wire [2:0] w_n588_0;
	wire [1:0] w_n588_1;
	wire [2:0] w_n589_0;
	wire [1:0] w_n589_1;
	wire [1:0] w_n591_0;
	wire [1:0] w_n592_0;
	wire [1:0] w_n599_0;
	wire [1:0] w_n605_0;
	wire [2:0] w_n606_0;
	wire [2:0] w_n606_1;
	wire [1:0] w_n607_0;
	wire [2:0] w_n608_0;
	wire [1:0] w_n610_0;
	wire [1:0] w_n612_0;
	wire [2:0] w_n613_0;
	wire [2:0] w_n615_0;
	wire [1:0] w_n615_1;
	wire [1:0] w_n617_0;
	wire [2:0] w_n618_0;
	wire [1:0] w_n619_0;
	wire [1:0] w_n620_0;
	wire [2:0] w_n621_0;
	wire [2:0] w_n622_0;
	wire [1:0] w_n622_1;
	wire [2:0] w_n623_0;
	wire [1:0] w_n624_0;
	wire [2:0] w_n625_0;
	wire [1:0] w_n626_0;
	wire [1:0] w_n627_0;
	wire [1:0] w_n628_0;
	wire [1:0] w_n629_0;
	wire [2:0] w_n630_0;
	wire [1:0] w_n631_0;
	wire [1:0] w_n632_0;
	wire [1:0] w_n633_0;
	wire [2:0] w_n634_0;
	wire [2:0] w_n635_0;
	wire [1:0] w_n637_0;
	wire [1:0] w_n642_0;
	wire [1:0] w_n643_0;
	wire [2:0] w_n645_0;
	wire [1:0] w_n647_0;
	wire [2:0] w_n648_0;
	wire [1:0] w_n649_0;
	wire [1:0] w_n650_0;
	wire [1:0] w_n652_0;
	wire [2:0] w_n653_0;
	wire [1:0] w_n653_1;
	wire [1:0] w_n656_0;
	wire [2:0] w_n657_0;
	wire [1:0] w_n657_1;
	wire [2:0] w_n658_0;
	wire [1:0] w_n659_0;
	wire [2:0] w_n660_0;
	wire [1:0] w_n660_1;
	wire [1:0] w_n661_0;
	wire [2:0] w_n662_0;
	wire [1:0] w_n663_0;
	wire [2:0] w_n664_0;
	wire [1:0] w_n664_1;
	wire [2:0] w_n665_0;
	wire [1:0] w_n666_0;
	wire [1:0] w_n667_0;
	wire [2:0] w_n668_0;
	wire [2:0] w_n669_0;
	wire [1:0] w_n671_0;
	wire [1:0] w_n672_0;
	wire [2:0] w_n673_0;
	wire [2:0] w_n674_0;
	wire [1:0] w_n674_1;
	wire [2:0] w_n675_0;
	wire [1:0] w_n676_0;
	wire [2:0] w_n677_0;
	wire [2:0] w_n678_0;
	wire [2:0] w_n679_0;
	wire [1:0] w_n679_1;
	wire [1:0] w_n680_0;
	wire [1:0] w_n683_0;
	wire [1:0] w_n686_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n690_0;
	wire [1:0] w_n692_0;
	wire [1:0] w_n693_0;
	wire [2:0] w_n697_0;
	wire [2:0] w_n699_0;
	wire [1:0] w_n699_1;
	wire [2:0] w_n701_0;
	wire [1:0] w_n701_1;
	wire [1:0] w_n703_0;
	wire [1:0] w_n704_0;
	wire [1:0] w_n705_0;
	wire [2:0] w_n707_0;
	wire [1:0] w_n708_0;
	wire [2:0] w_n709_0;
	wire [1:0] w_n709_1;
	wire [1:0] w_n710_0;
	wire [1:0] w_n711_0;
	wire [1:0] w_n712_0;
	wire [2:0] w_n713_0;
	wire [1:0] w_n713_1;
	wire [1:0] w_n714_0;
	wire [2:0] w_n715_0;
	wire [2:0] w_n716_0;
	wire [1:0] w_n716_1;
	wire [2:0] w_n720_0;
	wire [1:0] w_n720_1;
	wire [2:0] w_n723_0;
	wire [2:0] w_n727_0;
	wire [1:0] w_n728_0;
	wire [2:0] w_n730_0;
	wire [2:0] w_n734_0;
	wire [1:0] w_n735_0;
	wire [2:0] w_n737_0;
	wire [2:0] w_n741_0;
	wire [1:0] w_n742_0;
	wire [2:0] w_n744_0;
	wire [2:0] w_n748_0;
	wire [1:0] w_n751_0;
	wire [1:0] w_n752_0;
	wire [2:0] w_n754_0;
	wire [2:0] w_n758_0;
	wire [1:0] w_n759_0;
	wire [1:0] w_n764_0;
	wire [1:0] w_n765_0;
	wire [1:0] w_n782_0;
	wire [2:0] w_n784_0;
	wire [2:0] w_n787_0;
	wire [2:0] w_n790_0;
	wire [1:0] w_n790_1;
	wire [2:0] w_n793_0;
	wire [1:0] w_n793_1;
	wire [1:0] w_n795_0;
	wire [2:0] w_n797_0;
	wire [1:0] w_n797_1;
	wire [2:0] w_n801_0;
	wire [1:0] w_n801_1;
	wire [1:0] w_n802_0;
	wire [2:0] w_n804_0;
	wire [2:0] w_n807_0;
	wire [2:0] w_n810_0;
	wire [2:0] w_n812_0;
	wire [2:0] w_n816_0;
	wire [1:0] w_n817_0;
	wire [2:0] w_n819_0;
	wire [2:0] w_n823_0;
	wire [1:0] w_n824_0;
	wire [2:0] w_n827_0;
	wire [2:0] w_n831_0;
	wire [1:0] w_n832_0;
	wire [1:0] w_n834_0;
	wire [1:0] w_n838_0;
	wire [2:0] w_n843_0;
	wire [2:0] w_n847_0;
	wire [1:0] w_n848_0;
	wire [2:0] w_n851_0;
	wire [2:0] w_n855_0;
	wire [1:0] w_n856_0;
	wire [2:0] w_n858_0;
	wire [1:0] w_n859_0;
	wire [1:0] w_n864_0;
	wire [1:0] w_n865_0;
	wire [2:0] w_n869_0;
	wire [2:0] w_n873_0;
	wire [1:0] w_n874_0;
	wire [2:0] w_n878_0;
	wire [2:0] w_n882_0;
	wire [1:0] w_n885_0;
	wire [1:0] w_n887_0;
	wire [1:0] w_n889_0;
	wire [2:0] w_n891_0;
	wire [1:0] w_n891_1;
	wire [2:0] w_n895_0;
	wire [1:0] w_n895_1;
	wire [1:0] w_n896_0;
	wire [2:0] w_n899_0;
	wire [2:0] w_n902_0;
	wire [2:0] w_n905_0;
	wire [2:0] w_n908_0;
	wire [2:0] w_n912_0;
	wire [1:0] w_n913_0;
	wire [2:0] w_n916_0;
	wire [2:0] w_n920_0;
	wire [1:0] w_n921_0;
	wire [1:0] w_n923_0;
	wire [2:0] w_n927_0;
	wire [2:0] w_n931_0;
	wire [1:0] w_n932_0;
	wire [1:0] w_n935_0;
	wire [1:0] w_n937_0;
	wire [1:0] w_n939_0;
	wire [2:0] w_n945_0;
	wire [1:0] w_n945_1;
	wire [2:0] w_n948_0;
	wire [1:0] w_n948_1;
	wire [1:0] w_n950_0;
	wire [1:0] w_n952_0;
	wire [1:0] w_n957_0;
	wire [1:0] w_n972_0;
	wire [1:0] w_n981_0;
	wire [1:0] w_n987_0;
	wire [2:0] w_n988_0;
	wire [2:0] w_n992_0;
	wire [1:0] w_n993_0;
	wire [1:0] w_n994_0;
	wire [2:0] w_n995_0;
	wire [2:0] w_n999_0;
	wire [1:0] w_n1000_0;
	wire [1:0] w_n1003_0;
	wire [1:0] w_n1007_0;
	wire [1:0] w_n1008_0;
	wire [2:0] w_n1009_0;
	wire [1:0] w_n1009_1;
	wire [2:0] w_n1013_0;
	wire [1:0] w_n1013_1;
	wire [1:0] w_n1014_0;
	wire [1:0] w_n1015_0;
	wire [2:0] w_n1016_0;
	wire [2:0] w_n1019_0;
	wire [1:0] w_n1022_0;
	wire [1:0] w_n1033_0;
	wire [1:0] w_n1044_0;
	wire [2:0] w_n1061_0;
	wire [1:0] w_n1062_0;
	wire [2:0] w_n1066_0;
	wire [1:0] w_n1068_0;
	wire [1:0] w_n1069_0;
	wire [2:0] w_n1073_0;
	wire [1:0] w_n1075_0;
	wire [1:0] w_n1076_0;
	wire [2:0] w_n1077_0;
	wire [2:0] w_n1081_0;
	wire [1:0] w_n1082_0;
	wire [2:0] w_n1086_0;
	wire [1:0] w_n1092_0;
	wire [1:0] w_n1095_0;
	wire [2:0] w_n1096_0;
	wire [2:0] w_n1100_0;
	wire [1:0] w_n1102_0;
	wire [1:0] w_n1104_0;
	wire [1:0] w_n1105_0;
	wire [1:0] w_n1116_0;
	wire [2:0] w_n1122_0;
	wire [2:0] w_n1125_0;
	wire [1:0] w_n1127_0;
	wire [2:0] w_n1128_0;
	wire [1:0] w_n1128_1;
	wire [1:0] w_n1130_0;
	wire [1:0] w_n1136_0;
	wire [1:0] w_n1142_0;
	wire [2:0] w_n1148_0;
	wire [1:0] w_n1156_0;
	wire [1:0] w_n1166_0;
	wire [1:0] w_n1173_0;
	wire [1:0] w_n1189_0;
	wire [1:0] w_n1205_0;
	wire [1:0] w_n1236_0;
	wire [1:0] w_n1244_0;
	wire [1:0] w_n1283_0;
	wire [1:0] w_n1301_0;
	wire [1:0] w_n1309_0;
	wire [1:0] w_n1317_0;
	wire [1:0] w_n1325_0;
	wire [2:0] w_n1359_0;
	wire [2:0] w_n1360_0;
	wire [1:0] w_n1360_1;
	wire [1:0] w_n1361_0;
	wire [1:0] w_n1362_0;
	wire [1:0] w_n1376_0;
	wire [2:0] w_n1380_0;
	wire [1:0] w_n1380_1;
	wire [2:0] w_n1383_0;
	wire [2:0] w_n1383_1;
	wire [2:0] w_n1385_0;
	wire [1:0] w_n1385_1;
	wire [2:0] w_n1389_0;
	wire [1:0] w_n1389_1;
	wire [2:0] w_n1392_0;
	wire [1:0] w_n1392_1;
	wire [1:0] w_n1401_0;
	wire [1:0] w_n1402_0;
	wire [1:0] w_n1403_0;
	wire [1:0] w_n1404_0;
	wire [1:0] w_n1405_0;
	wire [1:0] w_n1406_0;
	wire [1:0] w_n1414_0;
	wire [2:0] w_n1420_0;
	wire [1:0] w_n1421_0;
	wire [1:0] w_n1422_0;
	wire [1:0] w_n1424_0;
	wire [1:0] w_n1425_0;
	wire [2:0] w_n1444_0;
	wire [1:0] w_n1445_0;
	wire [1:0] w_n1447_0;
	wire [1:0] w_n1454_0;
	wire [2:0] w_n1463_0;
	wire [1:0] w_n1464_0;
	wire [1:0] w_n1465_0;
	wire [1:0] w_n1468_0;
	wire [1:0] w_n1469_0;
	wire [1:0] w_n1470_0;
	wire [1:0] w_n1471_0;
	wire [1:0] w_n1472_0;
	wire [1:0] w_n1473_0;
	wire [1:0] w_n1479_0;
	wire [1:0] w_n1482_0;
	wire [1:0] w_n1486_0;
	wire [2:0] w_n1494_0;
	wire [1:0] w_n1501_0;
	wire [1:0] w_n1510_0;
	wire [1:0] w_n1520_0;
	wire [1:0] w_n1536_0;
	wire [1:0] w_n1571_0;
	wire [1:0] w_n1599_0;
	wire [1:0] w_n1610_0;
	wire [1:0] w_n1611_0;
	wire [1:0] w_n1625_0;
	wire [1:0] w_n1642_0;
	wire [1:0] w_n1644_0;
	wire [1:0] w_n1651_0;
	wire [1:0] w_n1654_0;
	wire [1:0] w_n1659_0;
	wire [1:0] w_n1667_0;
	wire [1:0] w_n1670_0;
	wire [1:0] w_n1672_0;
	wire [1:0] w_n1675_0;
	wire [1:0] w_n1680_0;
	wire [1:0] w_n1687_0;
	wire [1:0] w_n1689_0;
	wire [1:0] w_n1699_0;
	wire w_dff_A_H1x1fNcX7_0;
	wire w_dff_A_LJ5eExnU7_0;
	wire w_dff_A_2Rxoc2Fc8_1;
	wire w_dff_A_DJsdh6RM2_1;
	wire w_dff_A_Csyy1rkH6_1;
	wire w_dff_A_FaHfh2fO1_2;
	wire w_dff_B_aOYLngUM6_0;
	wire w_dff_B_8GT5GJoe7_3;
	wire w_dff_B_Fh6oaYhI2_3;
	wire w_dff_B_PdMoONtd1_3;
	wire w_dff_B_p4BRydNP0_3;
	wire w_dff_B_ZthGTssf3_3;
	wire w_dff_B_o9rZ0ppE2_3;
	wire w_dff_B_uBKdNDcH8_3;
	wire w_dff_B_Obt8tKE48_3;
	wire w_dff_B_1hfgjHjp7_3;
	wire w_dff_B_pSXeCuZx2_3;
	wire w_dff_B_SkkVDdcH5_3;
	wire w_dff_B_oos6ncU33_3;
	wire w_dff_B_aX6FGgSH8_3;
	wire w_dff_B_2zK51HxV0_3;
	wire w_dff_B_dPUIaYT13_3;
	wire w_dff_B_4GVNBzqu1_3;
	wire w_dff_B_nmwzeh3H7_1;
	wire w_dff_B_zluYwsbb9_0;
	wire w_dff_B_kmsBd3pO9_0;
	wire w_dff_B_LJchpJ413_0;
	wire w_dff_B_ZknSM7Q69_0;
	wire w_dff_B_tPUdWo8h1_0;
	wire w_dff_B_Jg7oXZfN3_0;
	wire w_dff_B_O9PQ5rko9_0;
	wire w_dff_B_IKeI7tOk1_0;
	wire w_dff_B_eaos86KW9_0;
	wire w_dff_B_CmYdmzaQ9_0;
	wire w_dff_B_RqVXRd1E5_0;
	wire w_dff_B_PlJ4JVtI2_0;
	wire w_dff_B_xZjP3xbI8_0;
	wire w_dff_B_rgTnpi6f8_0;
	wire w_dff_B_5b8wHGdI0_0;
	wire w_dff_B_cx1mKahK3_0;
	wire w_dff_B_sOzLRDlF8_0;
	wire w_dff_B_RPVfbBDI2_0;
	wire w_dff_B_lbPZEWeQ2_0;
	wire w_dff_B_YzKhEAQz8_0;
	wire w_dff_B_sybW8anM3_0;
	wire w_dff_B_LoxfYKrX8_1;
	wire w_dff_B_Taz8ROiW9_1;
	wire w_dff_B_ucUW0KpF7_1;
	wire w_dff_A_dNJIceBS3_1;
	wire w_dff_A_W8W1Fbec0_0;
	wire w_dff_A_JEJp4n9Z2_0;
	wire w_dff_A_wZ1bMUCk5_0;
	wire w_dff_B_clBketc26_0;
	wire w_dff_B_owubJqtn6_0;
	wire w_dff_B_uGdKD9RF0_0;
	wire w_dff_B_3YcnjEPM0_0;
	wire w_dff_B_Ke6pguCj6_0;
	wire w_dff_B_Qusatsm47_0;
	wire w_dff_B_xLARylk14_0;
	wire w_dff_B_Y78YgRbs9_0;
	wire w_dff_B_Szp1HVeJ0_0;
	wire w_dff_B_yrJTjGSX8_0;
	wire w_dff_A_wKweXwCq6_1;
	wire w_dff_A_JYNCkgNE3_1;
	wire w_dff_A_29vt0Iai6_1;
	wire w_dff_A_upaUkcFz2_1;
	wire w_dff_A_xwS9Vmph3_1;
	wire w_dff_A_QwCMM5pe6_1;
	wire w_dff_B_RBqfXNkC9_2;
	wire w_dff_B_M2eV6rMb1_0;
	wire w_dff_B_fECzl2j29_0;
	wire w_dff_B_A2vgLadr0_0;
	wire w_dff_A_1Do7kB6g2_0;
	wire w_dff_A_hFQ53zNg9_0;
	wire w_dff_A_TnOnyZIt6_1;
	wire w_dff_B_vsnB5BLX1_1;
	wire w_dff_B_Hlblfcs99_1;
	wire w_dff_B_CF1uAkos3_1;
	wire w_dff_B_omwt6g2n2_1;
	wire w_dff_B_zEB8zR890_0;
	wire w_dff_B_X0fm0r7M0_0;
	wire w_dff_A_b3Ut7UhH7_1;
	wire w_dff_A_op38Mzqe5_1;
	wire w_dff_A_uxOA9Led6_1;
	wire w_dff_A_TXy3bDe50_1;
	wire w_dff_A_u8gNdpKz3_1;
	wire w_dff_B_NjHQMahz2_1;
	wire w_dff_B_UQ2eWhvW8_0;
	wire w_dff_B_rz3yo8bX1_0;
	wire w_dff_B_pgl8Hcza8_0;
	wire w_dff_B_iEn66Zu24_0;
	wire w_dff_A_9oY2BN3F2_0;
	wire w_dff_A_nSYGefZu7_0;
	wire w_dff_A_YZHuPk2K1_1;
	wire w_dff_A_WfDfgt2O1_1;
	wire w_dff_A_F4VMf2ru8_1;
	wire w_dff_A_HiQIEYI01_1;
	wire w_dff_B_zZtQAI2w2_2;
	wire w_dff_A_9nUYdiC35_1;
	wire w_dff_A_jmBMnJRL4_1;
	wire w_dff_A_c7cyeEG07_1;
	wire w_dff_A_oja2GgdL4_1;
	wire w_dff_B_qex5kdE77_2;
	wire w_dff_B_E2BqAmmD6_1;
	wire w_dff_B_hlUP6DoB9_1;
	wire w_dff_B_gUT1FJ6E2_1;
	wire w_dff_B_VebpQi8Y0_1;
	wire w_dff_B_Iv8egv9x3_0;
	wire w_dff_B_QS8e2wgJ2_0;
	wire w_dff_B_0r9OQegj7_0;
	wire w_dff_B_cf8N8jNw3_1;
	wire w_dff_B_hzR408JK2_1;
	wire w_dff_B_dHwOYEWc2_1;
	wire w_dff_B_jbgvIvE76_1;
	wire w_dff_B_gUelUwAH4_1;
	wire w_dff_B_DjlADNOI5_1;
	wire w_dff_B_Jfuhpsui9_1;
	wire w_dff_B_vti9Bbka6_1;
	wire w_dff_B_K6n9Gu5M3_1;
	wire w_dff_B_oKPFqOOM6_1;
	wire w_dff_B_zGP8pgHY2_1;
	wire w_dff_A_Dbnl3XpI9_0;
	wire w_dff_B_La6IPfwy8_1;
	wire w_dff_A_hfnE4kP47_1;
	wire w_dff_A_DYqfH4B18_0;
	wire w_dff_B_mUrVDMiY4_3;
	wire w_dff_B_NunZNfAB4_0;
	wire w_dff_B_UPaggQHO7_0;
	wire w_dff_A_yVSrZYYS8_0;
	wire w_dff_B_JyTawwKo8_2;
	wire w_dff_B_73b3XT5p2_0;
	wire w_dff_B_yYE49MnY2_0;
	wire w_dff_B_bSp9X1LY2_0;
	wire w_dff_B_Crt9Bh7Q1_0;
	wire w_dff_B_ipreZXo37_0;
	wire w_dff_B_E1vqs5So6_2;
	wire w_dff_A_FaUhQEIr8_1;
	wire w_dff_B_oyvPw3HP8_0;
	wire w_dff_A_uSouiXpl1_0;
	wire w_dff_A_kpWQCibZ0_0;
	wire w_dff_A_KeBEqL1b9_0;
	wire w_dff_A_eXNx4TLQ8_0;
	wire w_dff_A_7geiDjfL8_0;
	wire w_dff_A_x8erXmeB9_0;
	wire w_dff_B_olKMC4kn6_1;
	wire w_dff_B_BB9j9eEC6_1;
	wire w_dff_B_eyGmmzk53_0;
	wire w_dff_B_hc7iIvA21_1;
	wire w_dff_A_4emVkdrr4_0;
	wire w_dff_A_34VAu1QY2_0;
	wire w_dff_A_ZsIGRV5g6_0;
	wire w_dff_A_DxoGZ2jD9_0;
	wire w_dff_A_KOtvCfEw3_0;
	wire w_dff_A_FS4dxPOV8_0;
	wire w_dff_B_BaWeFQ4N1_0;
	wire w_dff_A_KD4wimPd0_0;
	wire w_dff_A_IUzccUPO8_2;
	wire w_dff_A_YBvaUdOP4_1;
	wire w_dff_A_wB9sN0yI0_0;
	wire w_dff_A_cZ3tvlSy3_0;
	wire w_dff_A_30epYld30_0;
	wire w_dff_A_tK5Ktzi97_0;
	wire w_dff_A_tNzfigGw5_0;
	wire w_dff_A_M6GKYzr27_0;
	wire w_dff_A_yE9Belt04_0;
	wire w_dff_A_NdAjGV575_0;
	wire w_dff_A_n3OppnbW5_2;
	wire w_dff_B_0A8unDCZ9_3;
	wire w_dff_B_EsG6Kwdn3_3;
	wire w_dff_A_BxmbYe4G3_0;
	wire w_dff_A_vxfEyPsa7_0;
	wire w_dff_A_DoJtKWku7_0;
	wire w_dff_A_wblS193s2_0;
	wire w_dff_A_ioM7agik6_0;
	wire w_dff_A_a30oBt2Z5_0;
	wire w_dff_A_olH5ydUu8_0;
	wire w_dff_B_BGQRYwhH0_2;
	wire w_dff_B_ocApAAlI3_1;
	wire w_dff_B_hntVSUkP1_1;
	wire w_dff_B_HRf6BwCS8_1;
	wire w_dff_A_rQDQa0fV1_0;
	wire w_dff_B_Qcden2jP5_2;
	wire w_dff_B_VOOtMusF2_2;
	wire w_dff_B_IblNFaSL7_2;
	wire w_dff_B_KxNlxfcE2_2;
	wire w_dff_B_x5jDJCzn2_2;
	wire w_dff_B_RwQl9RZp8_2;
	wire w_dff_B_wQV5JdOo7_2;
	wire w_dff_B_WKJbX2TY6_2;
	wire w_dff_B_YJqjLwA85_2;
	wire w_dff_B_UJMbps260_2;
	wire w_dff_B_H8qyBEwP5_2;
	wire w_dff_B_eQgywDC07_2;
	wire w_dff_B_zDz5HAab4_2;
	wire w_dff_A_U5A0OWvQ2_0;
	wire w_dff_B_8OKTv9XE9_2;
	wire w_dff_B_GD9uVb5h8_2;
	wire w_dff_B_U2Q129iN0_2;
	wire w_dff_B_NgjrwS3f3_2;
	wire w_dff_B_EM70p3Km8_2;
	wire w_dff_B_xayyrLPC6_2;
	wire w_dff_B_0gN2yr7p2_2;
	wire w_dff_B_Eo2L0ZQs7_2;
	wire w_dff_B_ps9EMUV09_2;
	wire w_dff_B_w6PwYQ2n3_2;
	wire w_dff_B_SITQzVFv6_2;
	wire w_dff_B_0l4IU0o40_2;
	wire w_dff_B_mKUwH91I0_1;
	wire w_dff_B_kdpLK6Ir2_1;
	wire w_dff_B_pKPkoAf66_1;
	wire w_dff_B_7X10Oy2z1_1;
	wire w_dff_B_YHswpmBN6_1;
	wire w_dff_B_hTLr99948_1;
	wire w_dff_B_kh0mG0oH5_1;
	wire w_dff_B_UXERPa0q1_1;
	wire w_dff_B_wiYCOpmh7_1;
	wire w_dff_B_YnIuCaKP6_1;
	wire w_dff_B_NWEmCtOZ2_1;
	wire w_dff_B_wCjmDPvJ6_1;
	wire w_dff_A_D6vLbTgQ8_0;
	wire w_dff_B_53fwDjvP2_2;
	wire w_dff_B_QOYar6qD9_2;
	wire w_dff_B_vleLRqDg6_2;
	wire w_dff_B_3bb3j1dn9_2;
	wire w_dff_B_IPMENRrq7_2;
	wire w_dff_B_o3Jo6RyQ2_2;
	wire w_dff_B_jhaJRz5v8_2;
	wire w_dff_B_LDnfabSV4_2;
	wire w_dff_B_LU6tQWlE5_2;
	wire w_dff_B_koyHqIvp9_2;
	wire w_dff_B_uYehnKMl7_2;
	wire w_dff_B_XagOhMGU8_2;
	wire w_dff_B_WRvEsVRJ4_2;
	wire w_dff_B_0DdkLjYW4_2;
	wire w_dff_B_KFLkPMMh7_2;
	wire w_dff_B_NaOW4y5v8_2;
	wire w_dff_B_6nDF9O8S7_2;
	wire w_dff_B_x5PVJcHZ1_1;
	wire w_dff_B_EhEJoKax5_1;
	wire w_dff_B_gh8Zhfvx7_1;
	wire w_dff_B_cZNQdkW77_1;
	wire w_dff_B_I7eyIFiw4_1;
	wire w_dff_B_zZiQPSHB6_1;
	wire w_dff_B_MkJ4RXvv1_1;
	wire w_dff_B_N3I8Jjz22_1;
	wire w_dff_B_f0Uny1RB5_1;
	wire w_dff_B_asBaZ9r35_1;
	wire w_dff_B_BeNWbI3f0_1;
	wire w_dff_B_latO3i3i6_1;
	wire w_dff_B_nxH7yyo68_1;
	wire w_dff_B_KQXKqvIk2_0;
	wire w_dff_B_IZwVng5o1_0;
	wire w_dff_B_vzpbRXCp6_0;
	wire w_dff_B_2Bc6UJop7_0;
	wire w_dff_B_sqMfXfB26_0;
	wire w_dff_B_okDF1nOz8_0;
	wire w_dff_B_3Hwed9uF8_0;
	wire w_dff_B_gce3rBAo9_0;
	wire w_dff_B_PrrVwQBD1_0;
	wire w_dff_B_mhxu8Eq72_0;
	wire w_dff_B_2ErCsl821_0;
	wire w_dff_B_09oTuabG4_0;
	wire w_dff_B_HjQBwVVw1_0;
	wire w_dff_B_KHPRBnxK0_0;
	wire w_dff_A_0Tg0GVpc8_0;
	wire w_dff_B_NpolJDHj7_2;
	wire w_dff_B_aTtyaxgO4_2;
	wire w_dff_B_cvk4diKq2_2;
	wire w_dff_B_XN4lpS7F4_2;
	wire w_dff_B_VzR6Q3Nw9_2;
	wire w_dff_B_WaMjxWFi9_2;
	wire w_dff_B_wzO7q3NX5_2;
	wire w_dff_B_EljRkBnR8_2;
	wire w_dff_B_FjHYRCtP3_2;
	wire w_dff_B_Wyodgqcx1_2;
	wire w_dff_B_5WyXIVz35_2;
	wire w_dff_B_CvXfG5r89_2;
	wire w_dff_B_mbFam3nO9_2;
	wire w_dff_B_XHdLJZGC4_2;
	wire w_dff_B_UQDYOXCH3_2;
	wire w_dff_B_Hq71TNA62_2;
	wire w_dff_B_mr5mYk7H5_0;
	wire w_dff_B_QD0a7OGU7_0;
	wire w_dff_B_P52bzwOL2_0;
	wire w_dff_B_6E67m9nk2_0;
	wire w_dff_B_o6C0FC1J8_0;
	wire w_dff_B_gmsbbxjL8_0;
	wire w_dff_B_pP0s51ua1_0;
	wire w_dff_B_173T7hMJ2_0;
	wire w_dff_B_Q74RQj760_0;
	wire w_dff_B_HWQXCFiG4_1;
	wire w_dff_B_NHTV8UlK1_1;
	wire w_dff_B_fWbOweMG4_0;
	wire w_dff_B_fjEFjj683_1;
	wire w_dff_B_EhhukHxl3_1;
	wire w_dff_B_uzyJlzBQ0_1;
	wire w_dff_B_9IECpHVC3_1;
	wire w_dff_B_Wv8yPjb91_1;
	wire w_dff_B_pSO67Ttc4_1;
	wire w_dff_B_Y3DHXPlw4_1;
	wire w_dff_B_DJ4w6L5y8_1;
	wire w_dff_B_OGURsFGT2_1;
	wire w_dff_B_W377iLEv9_1;
	wire w_dff_B_SyQToNJc4_1;
	wire w_dff_B_BdmlA7k07_1;
	wire w_dff_B_9gASExGS4_0;
	wire w_dff_B_tDGVdp7M2_0;
	wire w_dff_B_sVv5WnBc8_1;
	wire w_dff_B_rqPeaL4Q4_1;
	wire w_dff_B_UYU4h3RQ3_1;
	wire w_dff_B_oe85dSHx4_1;
	wire w_dff_B_Z1bZWMPx7_1;
	wire w_dff_B_TvFokxhq6_1;
	wire w_dff_B_xHL8bKfi8_1;
	wire w_dff_B_ORUhP1w48_1;
	wire w_dff_B_boMQhpJ27_0;
	wire w_dff_B_Mq6MvMiN9_0;
	wire w_dff_B_opeCNCVQ1_0;
	wire w_dff_B_bpWNMMEc7_0;
	wire w_dff_B_cRJVO95d6_0;
	wire w_dff_B_B2EznjiX3_0;
	wire w_dff_B_gjvsLsyS4_0;
	wire w_dff_B_WHtaxa8G1_1;
	wire w_dff_B_nlwoff1o3_1;
	wire w_dff_B_0ZQfZymY9_1;
	wire w_dff_B_BRbGO4Yg4_1;
	wire w_dff_B_cIktG6lr3_1;
	wire w_dff_B_LfJWX3D13_1;
	wire w_dff_B_MCaZvy6c3_0;
	wire w_dff_B_2hXY8mZJ4_0;
	wire w_dff_B_uQvFpwT72_0;
	wire w_dff_B_ZhNlUfdm8_0;
	wire w_dff_B_OEvkFNga5_0;
	wire w_dff_B_bRo8Z4hO6_0;
	wire w_dff_B_kwT9n1fz3_0;
	wire w_dff_B_jMZecd1B1_0;
	wire w_dff_B_xFKgSs601_0;
	wire w_dff_B_mds2AIK08_0;
	wire w_dff_B_2pGwruPz1_0;
	wire w_dff_A_FCPrPmIm8_0;
	wire w_dff_B_uYOex2N95_0;
	wire w_dff_B_1NXFRMjk4_1;
	wire w_dff_B_rreQ0XYf0_1;
	wire w_dff_B_gICgOpXL2_1;
	wire w_dff_B_yLk5tBE51_1;
	wire w_dff_B_p3lLlLER1_1;
	wire w_dff_B_Ua5UgG9c8_0;
	wire w_dff_B_N64ZuN0W7_0;
	wire w_dff_B_rtQVUCQU1_0;
	wire w_dff_B_fPYqTgMv3_0;
	wire w_dff_B_83WXd5ql7_0;
	wire w_dff_B_ppmXzpJe8_0;
	wire w_dff_B_1MoapjDq3_0;
	wire w_dff_B_PhDfeFx85_0;
	wire w_dff_B_rf7vgArF7_0;
	wire w_dff_B_rVvKV7Bp3_0;
	wire w_dff_B_n43mFXus8_1;
	wire w_dff_B_lQ8Q3Dii3_1;
	wire w_dff_B_v0ffNHLM7_1;
	wire w_dff_B_CN1hRy5D4_0;
	wire w_dff_B_7XSr0N1X0_0;
	wire w_dff_A_xTpTo3FQ6_1;
	wire w_dff_B_8XEg0JBA1_0;
	wire w_dff_B_0p1asTaz8_0;
	wire w_dff_B_GHMBKMEz3_0;
	wire w_dff_B_3u7H70DV1_0;
	wire w_dff_B_ACQkRp2d8_0;
	wire w_dff_B_ZkCoSXX81_0;
	wire w_dff_B_lXAUZjrw9_0;
	wire w_dff_B_FVEpOpmI2_0;
	wire w_dff_B_Cq4SEy4M3_0;
	wire w_dff_B_VWQRY0eh8_0;
	wire w_dff_B_pEGy5yFX6_0;
	wire w_dff_B_QcCZd2tT0_0;
	wire w_dff_B_lMdIjjqA3_0;
	wire w_dff_A_jov50joB5_1;
	wire w_dff_B_y2mL8afH4_0;
	wire w_dff_B_yCOS2wms3_0;
	wire w_dff_B_BdF6J7Nd9_0;
	wire w_dff_B_UYt0YtB46_0;
	wire w_dff_A_VL9wH6h17_0;
	wire w_dff_A_XC64y0ZQ7_0;
	wire w_dff_B_h00Pwn007_0;
	wire w_dff_B_fIb3v3qv5_1;
	wire w_dff_B_xEb6tKc84_0;
	wire w_dff_B_P2YIAgvt6_0;
	wire w_dff_B_4Ng3MVty1_0;
	wire w_dff_B_mxs537I87_0;
	wire w_dff_A_2DeFixeh3_2;
	wire w_dff_A_p6fYGlLf3_2;
	wire w_dff_A_n6hM84nC4_0;
	wire w_dff_A_VqC2Fu7o5_0;
	wire w_dff_B_7fLkiLQM3_0;
	wire w_dff_A_c2BPqbnV3_0;
	wire w_dff_A_v1DXBwy66_0;
	wire w_dff_B_t28gJu808_0;
	wire w_dff_A_tvyGr8hS2_0;
	wire w_dff_A_mwjuaXS58_1;
	wire w_dff_B_cmy3iLci6_1;
	wire w_dff_B_b19WWDy46_0;
	wire w_dff_A_RBRzs81B1_0;
	wire w_dff_B_FnEjt97S5_0;
	wire w_dff_A_L9yEVs9h8_0;
	wire w_dff_A_GksR6ZpJ8_0;
	wire w_dff_A_CfZ6Oqln4_0;
	wire w_dff_B_64dqJnW15_1;
	wire w_dff_B_W3BPbTjj3_1;
	wire w_dff_B_OP2RUF7k2_0;
	wire w_dff_B_Lcgy86XL0_0;
	wire w_dff_B_U1958RBQ3_0;
	wire w_dff_B_hfEIVdUV0_1;
	wire w_dff_B_ZvV1HQX72_0;
	wire w_dff_B_m2voZ3vE6_0;
	wire w_dff_A_xccNKG1p6_1;
	wire w_dff_B_UY3GNvtW9_0;
	wire w_dff_B_eCcZfGh83_0;
	wire w_dff_B_gbjOsGnH4_0;
	wire w_dff_B_l5t1Lzlf2_0;
	wire w_dff_A_81yKPvvS6_0;
	wire w_dff_A_MOHz5gvg5_0;
	wire w_dff_B_Ys5oJSE10_0;
	wire w_dff_B_NBUZtjFn9_1;
	wire w_dff_B_Q9WaGEmw0_0;
	wire w_dff_B_9hGaIqOb4_0;
	wire w_dff_B_R6DqXCQT1_0;
	wire w_dff_A_1y77Buen6_0;
	wire w_dff_B_FkoeeYcx3_0;
	wire w_dff_A_Um3i6k0s2_0;
	wire w_dff_B_zwpHeb496_0;
	wire w_dff_B_hCoIS9vy3_1;
	wire w_dff_B_4F3mVGZg2_0;
	wire w_dff_B_6eM1AfF22_0;
	wire w_dff_A_Aax5Nc2t1_1;
	wire w_dff_B_AqWoWdRJ9_1;
	wire w_dff_B_1rCp1k1u8_1;
	wire w_dff_B_UT9nz9814_1;
	wire w_dff_B_fsMbef7P3_1;
	wire w_dff_B_aLTbXciP5_1;
	wire w_dff_A_Rjv8E4uC9_1;
	wire w_dff_A_DWrTK79g5_2;
	wire w_dff_B_IUEL5QAU1_1;
	wire w_dff_B_hNhDWOew7_1;
	wire w_dff_A_8QpsK7Yt1_1;
	wire w_dff_A_5CD2Eegm4_2;
	wire w_dff_B_PUf4qp3b3_1;
	wire w_dff_A_1PkpiUyh1_1;
	wire w_dff_A_QYNBPp378_2;
	wire w_dff_B_JfloGEvr0_1;
	wire w_dff_A_SJRSbQzT0_1;
	wire w_dff_A_M23IpCZd7_2;
	wire w_dff_B_uXICOqHD1_1;
	wire w_dff_A_Omj3E1au7_0;
	wire w_dff_A_OMALyz483_2;
	wire w_dff_B_tcaMqhgn1_1;
	wire w_dff_A_d6l7CZCQ0_1;
	wire w_dff_A_r5guVyE14_2;
	wire w_dff_B_zE8vol1i0_1;
	wire w_dff_A_IJjwYJTk3_0;
	wire w_dff_A_MeVxKv7k8_0;
	wire w_dff_A_ZmKoTLCU6_1;
	wire w_dff_B_CzetVjBx0_3;
	wire w_dff_B_Bh5QiV947_1;
	wire w_dff_B_pos8EslO2_1;
	wire w_dff_B_bgi1gc382_1;
	wire w_dff_B_DbGk8HA50_1;
	wire w_dff_B_SJTdq7ix4_1;
	wire w_dff_B_GSjpiOkW6_0;
	wire w_dff_B_8LCFIIXv6_0;
	wire w_dff_A_8eJPHOff4_1;
	wire w_dff_A_3iXJCCI03_1;
	wire w_dff_B_aDgzSQ3W6_1;
	wire w_dff_B_sNtu3yve4_1;
	wire w_dff_B_XUlCmyH13_1;
	wire w_dff_B_B0owYQxb4_1;
	wire w_dff_B_F9BIbIMB5_1;
	wire w_dff_B_WDAEk5L34_1;
	wire w_dff_A_bQRHzGDs9_0;
	wire w_dff_B_02keszY75_1;
	wire w_dff_B_DAJuA5HC0_1;
	wire w_dff_B_P2O9N3ze6_1;
	wire w_dff_B_WBgQZcFf6_3;
	wire w_dff_B_Bcaf6cA64_3;
	wire w_dff_B_3eVDKZ8r3_3;
	wire w_dff_B_lqrthS1O3_3;
	wire w_dff_B_Jj3NHDP84_3;
	wire w_dff_B_KXnUiTzW5_3;
	wire w_dff_B_JD2Rz16V0_3;
	wire w_dff_B_aR637i0J9_3;
	wire w_dff_B_TJ6EZ4fW9_3;
	wire w_dff_B_uJQ2eOXl4_3;
	wire w_dff_B_0CMEndwP5_3;
	wire w_dff_B_V69zn5WE9_3;
	wire w_dff_B_SbyWKT4c1_3;
	wire w_dff_B_b5gDHqmV4_3;
	wire w_dff_B_kkRlhK8R5_3;
	wire w_dff_B_CXby5lLn8_3;
	wire w_dff_B_jh6Pz9Zb5_3;
	wire w_dff_B_5R7QQSBq3_3;
	wire w_dff_B_cB0oiWbK4_3;
	wire w_dff_B_ohEwP5um6_3;
	wire w_dff_B_fJVRGy5q8_3;
	wire w_dff_B_2oZZjT7X1_1;
	wire w_dff_B_KgojfExN2_1;
	wire w_dff_B_8UnFFy893_1;
	wire w_dff_B_tuSUn7M79_1;
	wire w_dff_B_bOcn9bFA5_1;
	wire w_dff_B_rCxV8oK94_1;
	wire w_dff_B_pXv33GAe6_1;
	wire w_dff_B_YSYV19dJ5_1;
	wire w_dff_B_ATGUKbGM5_1;
	wire w_dff_B_SzUDHR6b7_1;
	wire w_dff_B_LpWTZVwP6_1;
	wire w_dff_B_p6Dvi9i21_1;
	wire w_dff_B_oUEGXJvf0_1;
	wire w_dff_B_5FxkY6i03_1;
	wire w_dff_B_z5Hs1uc00_1;
	wire w_dff_B_yo79W8XW9_1;
	wire w_dff_A_X8KAt6jb7_0;
	wire w_dff_A_mNktjaKO5_1;
	wire w_dff_A_lX3g4Itf2_0;
	wire w_dff_B_dM42cA8C7_2;
	wire w_dff_B_MJTYYIxQ6_2;
	wire w_dff_B_GXOXjQLM0_2;
	wire w_dff_B_zEDiIaCw9_2;
	wire w_dff_B_G2n4ifS46_2;
	wire w_dff_B_yjrW8SYW8_2;
	wire w_dff_B_ldsqRPJP1_2;
	wire w_dff_B_AU69szzi5_2;
	wire w_dff_B_R8RVR4Em2_2;
	wire w_dff_A_ltbWdfQG3_0;
	wire w_dff_B_44HkEJvN5_2;
	wire w_dff_B_Qogw2FEU5_2;
	wire w_dff_B_c373aXyp3_2;
	wire w_dff_B_G54LPRDw9_2;
	wire w_dff_B_XD9VrQfq4_2;
	wire w_dff_B_BBr7EVxo5_2;
	wire w_dff_B_EsLk7yv80_2;
	wire w_dff_B_t0V9Cd6B6_1;
	wire w_dff_B_KUAIJL757_1;
	wire w_dff_B_oFG2qDPi6_1;
	wire w_dff_B_qu9AU5DH7_1;
	wire w_dff_B_e1LrZ9FG8_1;
	wire w_dff_B_Kqxsl6xq7_1;
	wire w_dff_B_0BdZoDHv6_1;
	wire w_dff_B_HtZdZ1D74_1;
	wire w_dff_B_iCMngwBU5_1;
	wire w_dff_B_d5fv3hk86_1;
	wire w_dff_B_SoWd5YXX4_1;
	wire w_dff_B_ryspUru82_1;
	wire w_dff_B_aYOpmNQu3_1;
	wire w_dff_B_9zrF3Isv5_1;
	wire w_dff_B_U8EmEL2h4_1;
	wire w_dff_B_LNzOzkYx4_0;
	wire w_dff_B_gnBCZDhH4_0;
	wire w_dff_B_J5xJEgnn2_0;
	wire w_dff_B_QTp7Gtxt6_0;
	wire w_dff_B_xR1d7E2a2_1;
	wire w_dff_B_u3cQHpfZ3_1;
	wire w_dff_B_AM7IyKHC6_1;
	wire w_dff_B_aI1HuN814_1;
	wire w_dff_B_HkRHqI9f6_1;
	wire w_dff_B_V4RiUXRg5_1;
	wire w_dff_B_AF1N2f3f8_1;
	wire w_dff_B_RAz5LPa67_1;
	wire w_dff_B_PSFf9n4w9_1;
	wire w_dff_B_HFTzXLQg0_1;
	wire w_dff_B_PYhRQtCE6_1;
	wire w_dff_B_X1okK80g2_1;
	wire w_dff_B_aeoxuii34_0;
	wire w_dff_B_Nh6WyFZo2_1;
	wire w_dff_B_xVxqDQz99_0;
	wire w_dff_A_189A6ZlH4_1;
	wire w_dff_A_eTuTsUzN9_1;
	wire w_dff_A_YeVLCuEd5_1;
	wire w_dff_A_7Sb9knEw0_1;
	wire w_dff_A_sBamll1V9_1;
	wire w_dff_A_pWlNBqqc1_1;
	wire w_dff_A_HTXHixWY6_1;
	wire w_dff_A_qm6gHRym3_1;
	wire w_dff_A_buTZcA207_1;
	wire w_dff_A_gQJETuFf1_1;
	wire w_dff_B_Qst8B18I0_1;
	wire w_dff_A_WVjGtuSH1_1;
	wire w_dff_A_mLbPJ5GU7_1;
	wire w_dff_A_OEGK5aPO0_1;
	wire w_dff_A_cA44UuRA4_1;
	wire w_dff_A_dtyJ8XnP2_1;
	wire w_dff_A_JTWpSgbv7_1;
	wire w_dff_A_TMhhQwq76_1;
	wire w_dff_A_sy9AdmYK5_1;
	wire w_dff_A_SuUZyTFP8_1;
	wire w_dff_B_KlXKBtaX3_2;
	wire w_dff_B_cUKLYI2q2_0;
	wire w_dff_B_LMw4H1BS8_0;
	wire w_dff_B_nHV2rcZB0_0;
	wire w_dff_B_3Z2683L62_1;
	wire w_dff_B_INRxn0Zf8_1;
	wire w_dff_B_qYyCQUq50_0;
	wire w_dff_B_puz4657M8_0;
	wire w_dff_B_h1hNkmOI9_0;
	wire w_dff_B_WS9Io77u8_1;
	wire w_dff_A_t08G5Bbe2_1;
	wire w_dff_A_LJD4TZIk5_1;
	wire w_dff_A_N9e8tcqr4_1;
	wire w_dff_A_F0FfSBz80_1;
	wire w_dff_A_B62EhZho3_1;
	wire w_dff_A_gKREzjCS2_1;
	wire w_dff_A_iasVbBSK8_1;
	wire w_dff_A_zCPEnLGe2_1;
	wire w_dff_A_HnnnsTka4_1;
	wire w_dff_B_kXOVzd9I2_2;
	wire w_dff_B_HTieYIFO7_2;
	wire w_dff_B_nevWWI0v8_2;
	wire w_dff_B_iSRBWQMZ6_2;
	wire w_dff_B_NIXbY9Ao0_2;
	wire w_dff_B_WUarIzIc6_2;
	wire w_dff_A_kUmEGgAQ2_1;
	wire w_dff_B_bKnFP9Jd3_0;
	wire w_dff_B_majlC20b5_0;
	wire w_dff_B_gLo6NdRF1_0;
	wire w_dff_B_Mm9GiAn24_0;
	wire w_dff_B_qRoOA2Qd9_0;
	wire w_dff_B_UMNJLbhl3_1;
	wire w_dff_B_4Vp9XJcD5_1;
	wire w_dff_B_9THo75lP0_1;
	wire w_dff_B_7Hmehq3E6_1;
	wire w_dff_B_r8AFxmE49_1;
	wire w_dff_B_jMIpVqyN4_1;
	wire w_dff_B_WfMAqJW37_0;
	wire w_dff_A_wXk9aqtR3_1;
	wire w_dff_A_C957GCgo6_1;
	wire w_dff_A_4vVxTJGK5_1;
	wire w_dff_A_fBWZPxuy6_1;
	wire w_dff_A_fTYnZjd86_1;
	wire w_dff_A_twiNsobd1_1;
	wire w_dff_A_Ad1WD2fp6_1;
	wire w_dff_A_se79etU97_1;
	wire w_dff_A_pOl1XUOm4_1;
	wire w_dff_A_JL2dJkcJ1_1;
	wire w_dff_A_vE50oDBr4_1;
	wire w_dff_B_UthSIp5O4_2;
	wire w_dff_B_8ozVRkdB5_0;
	wire w_dff_B_eAaxFN4c8_0;
	wire w_dff_B_GRpiWZ8t0_0;
	wire w_dff_B_sJXleZJV5_0;
	wire w_dff_B_82qNFKIF8_0;
	wire w_dff_B_B5qAVPdK2_0;
	wire w_dff_B_KoHBeDLk7_0;
	wire w_dff_A_xqicetMq9_0;
	wire w_dff_A_tj41q6wh8_0;
	wire w_dff_A_E6LFlpmq0_2;
	wire w_dff_A_k9KSXCIp0_2;
	wire w_dff_A_VYR4DypP3_2;
	wire w_dff_A_73fzXHMZ8_2;
	wire w_dff_A_PxD9yZqd5_2;
	wire w_dff_A_w0Iz6dlr5_2;
	wire w_dff_A_XqWRHUXo0_2;
	wire w_dff_A_DW5A0erl8_2;
	wire w_dff_A_BwmJgd5x7_2;
	wire w_dff_A_SLMe2BuB5_2;
	wire w_dff_A_uAmDQLEZ8_2;
	wire w_dff_A_NSIIuSUk2_2;
	wire w_dff_A_dlooAmvU0_2;
	wire w_dff_B_bRi3SU7w6_3;
	wire w_dff_B_Mb7QQDlE8_3;
	wire w_dff_B_atMmZB8Y1_3;
	wire w_dff_B_SI0CUn5e3_3;
	wire w_dff_A_BIyh4ZNm7_1;
	wire w_dff_A_bU0yKjex8_1;
	wire w_dff_A_garw6vSx8_1;
	wire w_dff_A_0bdyKZb81_1;
	wire w_dff_A_iatti9uZ2_1;
	wire w_dff_A_2EEXSPAA6_1;
	wire w_dff_A_54ofLsbF8_1;
	wire w_dff_A_7jKDsxoq3_1;
	wire w_dff_A_O2xzF8Dh2_1;
	wire w_dff_A_8QDMDMFw1_1;
	wire w_dff_A_mvDqumTc6_1;
	wire w_dff_A_uX2DG70z2_1;
	wire w_dff_B_jNmrxi3S8_2;
	wire w_dff_B_cZdZCxDD9_2;
	wire w_dff_B_Nc8LrthW4_2;
	wire w_dff_B_sThnjLOW4_2;
	wire w_dff_B_2jMqZwdh5_2;
	wire w_dff_B_kyfv9RBk3_0;
	wire w_dff_B_qMcc0HEP6_0;
	wire w_dff_B_YLdHd6tD0_0;
	wire w_dff_B_9YfKdWK08_1;
	wire w_dff_B_UQKYH9Ol9_1;
	wire w_dff_B_zccf1NQR1_1;
	wire w_dff_B_DsDLv6TT5_1;
	wire w_dff_B_Kf49E3wu8_1;
	wire w_dff_B_XjMt2yO34_1;
	wire w_dff_B_SySFhhGT3_1;
	wire w_dff_B_cNLpmMdh9_1;
	wire w_dff_B_MGzbcxmn3_1;
	wire w_dff_B_JUnEuirv2_1;
	wire w_dff_B_BhTQqvKk4_1;
	wire w_dff_B_OKiIDr9X6_1;
	wire w_dff_B_2O444AIl1_1;
	wire w_dff_B_EsPNKSXH3_1;
	wire w_dff_B_p4HONLhX2_1;
	wire w_dff_B_x2kVBAV96_1;
	wire w_dff_B_8qb9JnrM6_1;
	wire w_dff_B_bVCbw5jP6_0;
	wire w_dff_B_7FIOKbKe8_0;
	wire w_dff_B_9zCOOAxD2_0;
	wire w_dff_B_92bLwit86_0;
	wire w_dff_B_1nNq9ubr4_0;
	wire w_dff_B_WYKqQNdS8_0;
	wire w_dff_B_jgRtkKpr3_0;
	wire w_dff_B_E5nqfP4x2_0;
	wire w_dff_B_F2TP6eVx6_1;
	wire w_dff_B_cPEWPHhX5_1;
	wire w_dff_B_AQXSGaOY9_1;
	wire w_dff_B_Jdd7TguC6_0;
	wire w_dff_B_AsBXhVOA6_0;
	wire w_dff_B_gtqeDLaA1_0;
	wire w_dff_B_qUMsoeRw8_0;
	wire w_dff_B_54ePHx2p1_0;
	wire w_dff_B_VuDupfmp4_0;
	wire w_dff_B_UXMno1W47_0;
	wire w_dff_B_eqgWUqGr2_0;
	wire w_dff_B_d7qp4tb85_0;
	wire w_dff_B_11Q2SXGH8_0;
	wire w_dff_B_g6FwZoqP4_0;
	wire w_dff_B_oJAojJul3_0;
	wire w_dff_B_7T2CMOVL2_0;
	wire w_dff_B_qqXNUt202_0;
	wire w_dff_B_ESh5Qf9G8_0;
	wire w_dff_B_zxuyijCv3_0;
	wire w_dff_B_XZZm6ftf0_0;
	wire w_dff_A_PXGPS2LS4_1;
	wire w_dff_A_1W9ogM5S2_1;
	wire w_dff_A_YAhy02zL6_1;
	wire w_dff_A_hJn7yT7j7_1;
	wire w_dff_A_KuhxwjDN7_2;
	wire w_dff_A_9B3hDVd52_2;
	wire w_dff_A_VRs2VgW55_2;
	wire w_dff_A_uEyEvH4i8_2;
	wire w_dff_A_mTIZ4Kb78_2;
	wire w_dff_A_TwBweXs65_2;
	wire w_dff_A_yFR6T61W9_2;
	wire w_dff_A_LOyNwaeG2_2;
	wire w_dff_A_0VUNrvOx1_2;
	wire w_dff_A_K9bwiR2B9_2;
	wire w_dff_A_o0RjupcQ4_2;
	wire w_dff_A_5Ppzryr87_2;
	wire w_dff_A_D2lhm79R9_2;
	wire w_dff_A_whQeeJ9W9_2;
	wire w_dff_A_LDUmc2re1_2;
	wire w_dff_A_t7v2Foso9_2;
	wire w_dff_B_riTkMIhQ1_3;
	wire w_dff_B_BA6ypliL0_3;
	wire w_dff_B_prn8QpJd1_3;
	wire w_dff_B_uP0Es38F6_0;
	wire w_dff_B_ySHsmOrS1_0;
	wire w_dff_B_p8TN8DnC6_0;
	wire w_dff_B_PI4UAjCe7_0;
	wire w_dff_B_ULeS2Hdb5_0;
	wire w_dff_B_8MufqKta2_0;
	wire w_dff_B_BFXyUr5n4_0;
	wire w_dff_B_xS7EoXhY9_0;
	wire w_dff_B_M7sTA4wo4_0;
	wire w_dff_B_WMdstgmH6_0;
	wire w_dff_B_dQ2XVzZb1_0;
	wire w_dff_B_pBDQt7Fm1_0;
	wire w_dff_A_hYRC2GmT0_1;
	wire w_dff_A_ETdLGiEY0_1;
	wire w_dff_A_csLbnYY68_1;
	wire w_dff_A_KbhxKYfc1_1;
	wire w_dff_A_KIdcbo8U6_1;
	wire w_dff_A_cIAROaMX8_1;
	wire w_dff_A_ykPomkwX5_1;
	wire w_dff_B_wrLotaPu8_2;
	wire w_dff_B_qlpbRo6X8_2;
	wire w_dff_B_OslxSPui1_2;
	wire w_dff_B_LMZAH95D2_2;
	wire w_dff_B_W7sI2l7y4_2;
	wire w_dff_B_jY4d4e6v0_2;
	wire w_dff_B_xfjsJTi02_2;
	wire w_dff_B_MZyPwBM32_2;
	wire w_dff_B_XHc56SKP0_2;
	wire w_dff_B_ixzvRv4d5_2;
	wire w_dff_B_Ue1tB1dW8_2;
	wire w_dff_B_2rNbrDSn7_2;
	wire w_dff_B_HuXvoX1q7_0;
	wire w_dff_B_wIXhcqSn5_0;
	wire w_dff_B_AnSrUlyW8_0;
	wire w_dff_B_oUAMA5Bw9_0;
	wire w_dff_B_blBRfFA76_0;
	wire w_dff_B_RVNBsr5A7_0;
	wire w_dff_B_Feo5D2xO0_0;
	wire w_dff_B_vdXXe8U12_0;
	wire w_dff_B_mecUcKPL7_0;
	wire w_dff_B_6JClkLPU5_0;
	wire w_dff_B_iot4Zr9i4_0;
	wire w_dff_B_o9eZOgmS1_0;
	wire w_dff_B_GIOaFgy69_3;
	wire w_dff_B_AthcAGN26_3;
	wire w_dff_B_02lejIxl3_3;
	wire w_dff_B_Xp3YSTii9_3;
	wire w_dff_B_WHQ1Ggsp6_3;
	wire w_dff_B_CsnQHbpm0_3;
	wire w_dff_B_lLWNjJ9j3_3;
	wire w_dff_B_y3fjucnV8_3;
	wire w_dff_B_qJra4Pqc5_3;
	wire w_dff_B_l1SLN5z83_3;
	wire w_dff_B_vBcehRgJ4_3;
	wire w_dff_B_syuzaC8i3_3;
	wire w_dff_B_xWHdXOLP2_3;
	wire w_dff_B_fQZma7k94_3;
	wire w_dff_B_nKlIzAtF4_3;
	wire w_dff_B_fiaUomy91_3;
	wire w_dff_B_1rzDFzsj1_3;
	wire w_dff_B_wcNfDzhL9_3;
	wire w_dff_B_FivChyJd2_3;
	wire w_dff_A_2pLA6sGi2_0;
	wire w_dff_A_IScrSnDp4_0;
	wire w_dff_A_RIj09X6r4_0;
	wire w_dff_A_5miIlYs52_0;
	wire w_dff_A_8S2mVXtp5_0;
	wire w_dff_A_bVnIap0S4_0;
	wire w_dff_A_RUIAskX05_0;
	wire w_dff_A_bqr44H7R8_0;
	wire w_dff_A_s2bnclLQ6_0;
	wire w_dff_A_NKs9K9fI5_0;
	wire w_dff_A_rVwvjIRN8_0;
	wire w_dff_A_TEOTdLan2_0;
	wire w_dff_A_4pEt9iRe8_0;
	wire w_dff_A_2fsMJv6Z9_0;
	wire w_dff_A_rYs4GucR6_1;
	wire w_dff_A_DSUFAiTB4_1;
	wire w_dff_A_AAIVqFnq0_1;
	wire w_dff_A_aKdzrLD49_1;
	wire w_dff_A_93P75Fw56_1;
	wire w_dff_A_63JeO8yX5_1;
	wire w_dff_A_RToS7jYS6_1;
	wire w_dff_A_0N8FCyks1_1;
	wire w_dff_A_6EiRPQPw6_1;
	wire w_dff_A_DUwVtVMp5_1;
	wire w_dff_B_5GJbIelO2_1;
	wire w_dff_B_6QqI81sW6_1;
	wire w_dff_B_31axOZ779_1;
	wire w_dff_B_WcgBQG6L5_1;
	wire w_dff_B_AW24cn5E4_1;
	wire w_dff_B_98DFixQV3_1;
	wire w_dff_B_6CyJdoem4_1;
	wire w_dff_B_j5sFEgj30_1;
	wire w_dff_B_nBGwLroT7_1;
	wire w_dff_B_dBcfTNrF6_1;
	wire w_dff_B_QSBeyMPl2_1;
	wire w_dff_B_31TRHZrU5_1;
	wire w_dff_B_j117HOou5_1;
	wire w_dff_B_nAACLr1z2_1;
	wire w_dff_B_DQ1EHF7V3_1;
	wire w_dff_B_xJnr10EK2_1;
	wire w_dff_B_qnY7mpwh9_1;
	wire w_dff_B_CrkyE9VK5_1;
	wire w_dff_B_R8R1GegZ9_1;
	wire w_dff_A_b3NQQGGA8_0;
	wire w_dff_A_QP6gin3t0_0;
	wire w_dff_A_Cy4gb3jU5_0;
	wire w_dff_A_XtNZ2cwT4_0;
	wire w_dff_A_uztjHBXS0_0;
	wire w_dff_A_AFbJ8nJ87_0;
	wire w_dff_A_F2FgUrfK6_0;
	wire w_dff_A_0ehuDGa37_0;
	wire w_dff_A_geo1gBGY6_0;
	wire w_dff_A_QVllah6X5_0;
	wire w_dff_A_W7cqJDbd8_0;
	wire w_dff_B_mMspoOhi8_1;
	wire w_dff_B_SbXtGPCx1_1;
	wire w_dff_B_3RZrnDtC6_1;
	wire w_dff_B_k26eojcT9_1;
	wire w_dff_B_eirtcAzx3_1;
	wire w_dff_B_USI1XqZs9_1;
	wire w_dff_B_lbDXiSBl2_1;
	wire w_dff_B_c7vP74jz2_1;
	wire w_dff_B_fuS5g3We1_1;
	wire w_dff_B_ZrU08K1A0_0;
	wire w_dff_A_pDvDnkNp0_0;
	wire w_dff_A_VHmyh0658_0;
	wire w_dff_A_llREnJMm9_0;
	wire w_dff_A_5plgl53j5_0;
	wire w_dff_A_FUNQwxCo7_0;
	wire w_dff_A_rFRXfMHw8_0;
	wire w_dff_A_Heppkal78_0;
	wire w_dff_A_S98k5jCQ7_0;
	wire w_dff_A_yGyzPe4B2_0;
	wire w_dff_A_7FMjB3Vu6_0;
	wire w_dff_A_63wWsD236_0;
	wire w_dff_A_VnPbcDzP7_0;
	wire w_dff_A_u7F2Q8m55_1;
	wire w_dff_A_OXz8K64H4_1;
	wire w_dff_A_h6WxvGi87_1;
	wire w_dff_A_N1hFQIAX4_1;
	wire w_dff_A_kqHA7SEI9_1;
	wire w_dff_A_OHcH1tg02_1;
	wire w_dff_A_pIWS2X621_1;
	wire w_dff_A_Cy9aYAbq4_1;
	wire w_dff_A_fSmbRiGw6_1;
	wire w_dff_A_ntRiys6G6_1;
	wire w_dff_A_GtSFQ6Iu6_1;
	wire w_dff_A_NxWtbGzu4_1;
	wire w_dff_A_h48hVY0p1_1;
	wire w_dff_A_39wYxN6T5_1;
	wire w_dff_A_ywic1fHk4_1;
	wire w_dff_A_ohcuHZ8E6_1;
	wire w_dff_A_T8J0NI7b7_1;
	wire w_dff_A_N0r6384D1_1;
	wire w_dff_A_1IQtyevN2_1;
	wire w_dff_B_3CWIUYUh5_2;
	wire w_dff_B_ZSb2eyue1_2;
	wire w_dff_B_UEr6zIbv1_2;
	wire w_dff_B_JqLPROAF1_2;
	wire w_dff_B_FRjIx0s29_2;
	wire w_dff_A_0uQLXxFj7_0;
	wire w_dff_A_se3lgJdO6_0;
	wire w_dff_A_tw1W2qY31_0;
	wire w_dff_A_HijjC0fh7_0;
	wire w_dff_A_OzFdgeut2_0;
	wire w_dff_B_a6vI01Xa7_0;
	wire w_dff_B_PbVZSAaj7_0;
	wire w_dff_B_zoGqrCsr9_0;
	wire w_dff_B_8TrRRcVy0_0;
	wire w_dff_B_UD8zV4Fo8_0;
	wire w_dff_B_3vhR5FRd5_0;
	wire w_dff_B_egxG1bLp0_0;
	wire w_dff_B_wzsIbGOs3_0;
	wire w_dff_B_M597tXan2_0;
	wire w_dff_B_oSwk6T4H0_0;
	wire w_dff_B_lbYoKhjc4_0;
	wire w_dff_B_v6k1PaaS2_0;
	wire w_dff_A_nRk0F1yu3_0;
	wire w_dff_A_9F0lqJYL3_0;
	wire w_dff_A_ahdHbyKk0_0;
	wire w_dff_A_BsN9hC1e8_0;
	wire w_dff_A_bmHVwHPA3_0;
	wire w_dff_A_8v14q7Rr6_1;
	wire w_dff_A_bxt3cWg04_1;
	wire w_dff_A_ROvKrg5y1_2;
	wire w_dff_A_IUaQs51h2_0;
	wire w_dff_A_RQV5umD88_0;
	wire w_dff_A_DZvNQCFr8_0;
	wire w_dff_A_Efe0r4uT8_0;
	wire w_dff_A_BOeQg6d50_0;
	wire w_dff_A_mcxyT3IL0_0;
	wire w_dff_A_83idBDcV2_0;
	wire w_dff_A_1SOOwDKX2_0;
	wire w_dff_A_GfgfAQdm0_0;
	wire w_dff_A_qN9E9QMu1_0;
	wire w_dff_A_SZwoJk737_0;
	wire w_dff_A_FoAN2lGm2_0;
	wire w_dff_A_U9khHxe71_0;
	wire w_dff_A_LOgY3SDJ6_0;
	wire w_dff_A_24HZQlwX4_0;
	wire w_dff_A_Hk3heCbt6_0;
	wire w_dff_A_dy8idU0p2_1;
	wire w_dff_A_0k3ywTYN8_1;
	wire w_dff_A_FfUNx92S1_1;
	wire w_dff_A_xeqNNqnp7_1;
	wire w_dff_A_uhzyLWyT7_1;
	wire w_dff_A_yI1dmKmU2_1;
	wire w_dff_A_7ed9KzhY5_1;
	wire w_dff_A_g9dXKNb59_1;
	wire w_dff_A_fivInbil4_1;
	wire w_dff_A_TuC4Q1IY3_1;
	wire w_dff_A_zHTplkiB0_1;
	wire w_dff_A_HCOkP9kF2_1;
	wire w_dff_A_pFcKP18F0_1;
	wire w_dff_A_aQekNMNG6_1;
	wire w_dff_A_BrggSZaM2_1;
	wire w_dff_A_ksJ7tGhk9_1;
	wire w_dff_B_ntO3dZxz6_0;
	wire w_dff_B_Eb137lpD7_3;
	wire w_dff_B_1b42s4Cf3_3;
	wire w_dff_A_FXzQTZBz9_0;
	wire w_dff_A_W3wYQSli9_0;
	wire w_dff_A_JXQWSPKi0_0;
	wire w_dff_A_Vtxl6EgM4_0;
	wire w_dff_A_IS4t9m6n0_0;
	wire w_dff_A_qnmJzlNA5_0;
	wire w_dff_A_traQn1J99_0;
	wire w_dff_A_0KY4L7qb6_0;
	wire w_dff_A_cLN2eEGx0_0;
	wire w_dff_A_J3qQsUsv8_0;
	wire w_dff_A_hpwijWbA4_0;
	wire w_dff_A_w8FTFYUL0_0;
	wire w_dff_A_6Hl9xR1E1_0;
	wire w_dff_A_jPop937a0_0;
	wire w_dff_A_csVXd10E6_0;
	wire w_dff_A_m1C0VH770_0;
	wire w_dff_A_CIVjT5VM8_0;
	wire w_dff_A_v7RfquDs0_0;
	wire w_dff_A_QUy4eyxe1_1;
	wire w_dff_A_phBDlMg71_1;
	wire w_dff_A_fIC2p0Xx1_1;
	wire w_dff_A_uCNOdBRd7_1;
	wire w_dff_A_A0vxmUpU9_1;
	wire w_dff_A_TxJfzI5u1_1;
	wire w_dff_A_9Q4iBcA39_1;
	wire w_dff_A_OKZphSOh1_1;
	wire w_dff_A_pVVPqvYX2_1;
	wire w_dff_A_QZfrvL4I7_1;
	wire w_dff_A_8O7LrDql9_1;
	wire w_dff_A_FhDUAYYh0_1;
	wire w_dff_A_mzieiADk9_1;
	wire w_dff_A_ohXg0I1s7_0;
	wire w_dff_A_1aqJqf1o2_0;
	wire w_dff_B_k0FUDk4O7_0;
	wire w_dff_B_UFEOpjR45_2;
	wire w_dff_B_xfvM5hH19_2;
	wire w_dff_A_D4pDAyua3_0;
	wire w_dff_A_dA0aAkgi9_0;
	wire w_dff_A_66mRX9688_0;
	wire w_dff_A_6HCsU9672_0;
	wire w_dff_A_iVqUbNYz1_0;
	wire w_dff_A_Rt6Qggwj7_0;
	wire w_dff_B_XHcYUwEC3_0;
	wire w_dff_B_ZdNvDYb41_2;
	wire w_dff_B_xceFMOFW7_2;
	wire w_dff_A_IuovkDfs4_0;
	wire w_dff_A_A3N2WasT5_0;
	wire w_dff_A_v0z01ZgM1_0;
	wire w_dff_A_pPlrvx5T9_0;
	wire w_dff_B_n7oZ3W448_0;
	wire w_dff_B_rNlhbg6w2_3;
	wire w_dff_B_pmxFTMoD6_3;
	wire w_dff_A_N0kDuRwy6_1;
	wire w_dff_A_Ivn3BrT31_1;
	wire w_dff_B_tR2LbQ4n4_0;
	wire w_dff_B_z6Iml3TC6_3;
	wire w_dff_B_VXaHy9Hx2_3;
	wire w_dff_A_LhYOVxyI5_1;
	wire w_dff_A_Ug3mK5NG0_1;
	wire w_dff_A_7wd10qIo0_1;
	wire w_dff_A_EAb3kC1d5_1;
	wire w_dff_A_MAQeO5oo4_1;
	wire w_dff_A_B6LaQCym1_1;
	wire w_dff_A_mRWBJonj2_1;
	wire w_dff_A_15KflhwZ3_1;
	wire w_dff_A_HSuaGMv20_1;
	wire w_dff_B_fVfsT3JD2_1;
	wire w_dff_B_Mkxo0zjz7_1;
	wire w_dff_B_Z7mHQ0hz1_1;
	wire w_dff_B_M9KreNBI5_1;
	wire w_dff_B_hAhFDvod4_0;
	wire w_dff_B_QRx72X1R3_0;
	wire w_dff_A_nx74sppU0_0;
	wire w_dff_A_pLdcDt4v1_0;
	wire w_dff_A_UmgNyxXY9_0;
	wire w_dff_A_whLRc9xJ3_0;
	wire w_dff_A_mdlHZwOP4_0;
	wire w_dff_A_1lprh0ls4_0;
	wire w_dff_A_afMyLor28_0;
	wire w_dff_A_vQHn923G0_0;
	wire w_dff_A_H5ozfvEf8_0;
	wire w_dff_A_Bn4mYZrY0_0;
	wire w_dff_A_1fPSTm731_0;
	wire w_dff_A_hPBh4mk55_0;
	wire w_dff_A_LAnBHev18_0;
	wire w_dff_A_N85r8T5u6_0;
	wire w_dff_A_bYH1Yk4w1_0;
	wire w_dff_A_piWLtxRU3_1;
	wire w_dff_A_wne7cskn8_1;
	wire w_dff_A_sUtFUMxE0_1;
	wire w_dff_A_mni2gDwA4_1;
	wire w_dff_A_9qscZx968_1;
	wire w_dff_A_DOr04mro5_1;
	wire w_dff_A_VTSm0hsC0_1;
	wire w_dff_A_ZCxDpFtE6_1;
	wire w_dff_A_ucRnVag98_1;
	wire w_dff_A_0EK1odHV0_1;
	wire w_dff_A_PMyYqndW8_1;
	wire w_dff_A_DB7tKIUf7_1;
	wire w_dff_A_YR6YSlRF7_1;
	wire w_dff_A_IpbrTOhL4_1;
	wire w_dff_A_LnBaAuQd1_1;
	wire w_dff_B_C4tzDZ6m2_1;
	wire w_dff_A_NlXmhPtA6_0;
	wire w_dff_A_qb3jlVHQ1_1;
	wire w_dff_A_imvC1xlh9_1;
	wire w_dff_A_SlLxopcg6_1;
	wire w_dff_A_SntQfvgC6_1;
	wire w_dff_A_rORgkK0L6_1;
	wire w_dff_A_i8Ge2UoJ1_1;
	wire w_dff_A_xTDhwCkA7_1;
	wire w_dff_A_u1XntUmo6_1;
	wire w_dff_A_A3w1LbOh4_1;
	wire w_dff_A_hAcYqbdW5_1;
	wire w_dff_A_URvGaDG78_1;
	wire w_dff_A_o77milgf7_1;
	wire w_dff_A_UkMHL19G4_1;
	wire w_dff_A_TYce3fmA5_1;
	wire w_dff_A_xKhpYeJo3_1;
	wire w_dff_A_TF2dRplP6_0;
	wire w_dff_A_NSQ0FXRP2_0;
	wire w_dff_A_xjREGCon4_0;
	wire w_dff_A_gTFgY2Nd6_0;
	wire w_dff_A_YdIucaZ67_0;
	wire w_dff_A_WVB6Expa2_0;
	wire w_dff_A_b9qFrL5p4_0;
	wire w_dff_A_kZNUPEa16_0;
	wire w_dff_A_UzbzHfDK9_0;
	wire w_dff_A_bO5DoJI41_0;
	wire w_dff_A_BhdhF3A34_0;
	wire w_dff_A_H378nXVf0_0;
	wire w_dff_A_xApNFDDi8_0;
	wire w_dff_A_htWSNZ0U3_0;
	wire w_dff_B_8bzvD6Xj6_2;
	wire w_dff_B_64BnYiHV3_2;
	wire w_dff_A_kTkwB2Kb6_0;
	wire w_dff_A_g5E6Xoil8_0;
	wire w_dff_A_PxZd0RBT7_0;
	wire w_dff_A_e1l956lS8_0;
	wire w_dff_A_8nXhsAqp5_0;
	wire w_dff_B_ePSTFwxn2_0;
	wire w_dff_B_dZZlInJA2_0;
	wire w_dff_B_5FdAPyX25_0;
	wire w_dff_B_yE7AFs3X2_0;
	wire w_dff_B_P4AxfDd10_0;
	wire w_dff_B_2dTI95Ag6_0;
	wire w_dff_B_GJhZjZyj5_0;
	wire w_dff_B_GF1bxYkC6_0;
	wire w_dff_B_cDhyUstl7_0;
	wire w_dff_B_hyaXkRZh4_0;
	wire w_dff_B_5bVHzCoB6_0;
	wire w_dff_A_dI8kEoUQ0_0;
	wire w_dff_A_v283yLyc2_0;
	wire w_dff_A_9CzZbaMW0_0;
	wire w_dff_A_PTXyHzPb2_0;
	wire w_dff_A_7yrQxVyh3_0;
	wire w_dff_A_hXgRrwjt0_0;
	wire w_dff_A_mQ7JHL7A0_0;
	wire w_dff_A_jJWjSZLk1_0;
	wire w_dff_A_tGKiAFJ45_0;
	wire w_dff_A_OAwK0ZCv7_0;
	wire w_dff_A_GJ4scgZd6_0;
	wire w_dff_A_YBLe62Qq7_0;
	wire w_dff_A_U3iOSSB60_0;
	wire w_dff_A_BhhxFeUR3_0;
	wire w_dff_A_z6Z7PJLr0_0;
	wire w_dff_B_gmR2tVV00_0;
	wire w_dff_B_Wun7VePb7_2;
	wire w_dff_B_TLKxVHrz8_2;
	wire w_dff_A_5KOVEoVw7_0;
	wire w_dff_A_ZMWNQO8U4_0;
	wire w_dff_A_MwA18U3m5_0;
	wire w_dff_A_9uuk3uJU2_0;
	wire w_dff_A_PlpkORAv3_0;
	wire w_dff_A_EX3ZzQQk9_0;
	wire w_dff_B_9U7qMuqH0_0;
	wire w_dff_B_wkLN8WmT3_2;
	wire w_dff_B_KqGlf3EU9_2;
	wire w_dff_A_H4W4do6z0_0;
	wire w_dff_A_oif6KGoZ0_0;
	wire w_dff_A_8cHYjrwL0_0;
	wire w_dff_A_Of6m4djP1_0;
	wire w_dff_A_s8YrdGsc3_0;
	wire w_dff_A_RnCEZq7s6_0;
	wire w_dff_A_tjQ9oybE9_0;
	wire w_dff_A_CWdmyTBg6_0;
	wire w_dff_A_xgzkMFPV2_0;
	wire w_dff_A_n6EGCexi3_0;
	wire w_dff_A_Lyuesbap7_0;
	wire w_dff_A_UaKZasdC2_0;
	wire w_dff_A_xVfsRKwD1_0;
	wire w_dff_A_I12FHI8l0_0;
	wire w_dff_A_NRpGR77t6_0;
	wire w_dff_A_kOdyl9j68_0;
	wire w_dff_A_YcCrtlXV4_0;
	wire w_dff_A_DqfIZIe95_0;
	wire w_dff_A_OnR7F0Ov0_0;
	wire w_dff_A_xUWqSw9H1_0;
	wire w_dff_B_q90zLv3b6_0;
	wire w_dff_A_8IlHPIpi6_1;
	wire w_dff_A_hhuo9bPa3_1;
	wire w_dff_A_jOYC5UJN4_2;
	wire w_dff_A_82enB9Zl4_2;
	wire w_dff_A_K6kRUXt23_1;
	wire w_dff_A_lzE1Hsi35_1;
	wire w_dff_A_L8NjtLMm4_1;
	wire w_dff_A_mBJGbxOA3_1;
	wire w_dff_A_Jx6Nmo0H4_2;
	wire w_dff_A_Inpx9wdH7_2;
	wire w_dff_A_1sTzqk7F1_2;
	wire w_dff_A_n9sFzddv8_2;
	wire w_dff_A_5hBpT9Dg3_2;
	wire w_dff_A_H9zOAFHx9_2;
	wire w_dff_A_DepeEy322_2;
	wire w_dff_A_xiHKryJN7_2;
	wire w_dff_A_zCrUtDH90_2;
	wire w_dff_A_eN39hUaF2_2;
	wire w_dff_A_pLg4OBT42_2;
	wire w_dff_A_66N60CTd1_2;
	wire w_dff_A_famUi9Ow7_2;
	wire w_dff_A_FlQ3axMt0_2;
	wire w_dff_A_w0z19Z6F8_2;
	wire w_dff_A_QOjGnQml7_2;
	wire w_dff_A_j7dIH2GR1_0;
	wire w_dff_A_Kir7Rrku2_0;
	wire w_dff_B_ushaR9vI3_0;
	wire w_dff_B_g6uKnzF50_2;
	wire w_dff_B_an6MDwmU2_2;
	wire w_dff_A_7hEVAEFb8_1;
	wire w_dff_A_HWHE1biM3_1;
	wire w_dff_A_prTVDyTp7_1;
	wire w_dff_A_8ufHP8OR6_1;
	wire w_dff_A_6arFQ3iJ3_1;
	wire w_dff_B_7BmYyDMm7_1;
	wire w_dff_B_SlYEXmrL8_1;
	wire w_dff_B_xlCfDRVl8_1;
	wire w_dff_B_LHWRhSg61_1;
	wire w_dff_B_bOwuuzCy2_1;
	wire w_dff_B_9fDOTzUJ0_1;
	wire w_dff_B_D5Q2xOZA1_1;
	wire w_dff_B_yME1aZo34_1;
	wire w_dff_B_rpVKhQ6F6_1;
	wire w_dff_B_l3n405Ep5_1;
	wire w_dff_B_IFTfh1mX6_1;
	wire w_dff_A_81XBlqvm4_0;
	wire w_dff_A_D1phObl95_0;
	wire w_dff_A_uHmO9OH33_0;
	wire w_dff_A_h3AVsrzd6_0;
	wire w_dff_A_REXG7Zhp7_0;
	wire w_dff_A_vklsPczg5_0;
	wire w_dff_A_4QMJZCK65_0;
	wire w_dff_A_VsAIbkmZ9_0;
	wire w_dff_A_KrygBMp55_0;
	wire w_dff_B_6pPOnS6H0_1;
	wire w_dff_B_TlsEcBTW6_1;
	wire w_dff_B_iTUWS4sz1_1;
	wire w_dff_B_bO2tCcQc4_1;
	wire w_dff_B_x1Yl5yVa8_1;
	wire w_dff_B_wFDA0cag7_1;
	wire w_dff_B_PSNRXKgT4_1;
	wire w_dff_A_wjUihQaD1_1;
	wire w_dff_A_x70VSDT46_1;
	wire w_dff_A_KmiCco6I6_1;
	wire w_dff_A_JyowotkQ5_1;
	wire w_dff_A_5jgCpFzy0_1;
	wire w_dff_A_AmXvraAA1_1;
	wire w_dff_A_8UQcol652_1;
	wire w_dff_A_WbBHUvTq9_1;
	wire w_dff_A_9cezoIdV4_1;
	wire w_dff_A_AeGQcbZC4_1;
	wire w_dff_A_JOD0nreV1_0;
	wire w_dff_A_Nei84SfY4_0;
	wire w_dff_A_OyMjnSER3_0;
	wire w_dff_A_nv66cA3z1_0;
	wire w_dff_A_PGBKZuMi7_0;
	wire w_dff_A_D2YnCEkM4_0;
	wire w_dff_A_FuQ2lwZi3_0;
	wire w_dff_A_8CDfmc8z6_0;
	wire w_dff_A_gFW2FglF0_1;
	wire w_dff_A_MfH5EZsL5_1;
	wire w_dff_A_OgMELuPM1_1;
	wire w_dff_A_lI0VZls23_1;
	wire w_dff_A_y36RNCp36_1;
	wire w_dff_A_auSOT7Ez1_1;
	wire w_dff_A_07zLDTuy0_1;
	wire w_dff_A_3Gaffbtx8_1;
	wire w_dff_A_Legihi8a8_1;
	wire w_dff_A_pRiVCr5C8_1;
	wire w_dff_A_nQrK5SOy7_1;
	wire w_dff_A_90PfBetN6_1;
	wire w_dff_A_sIc5B8IA5_1;
	wire w_dff_A_bpIZOWyw1_0;
	wire w_dff_A_gsuy1xhg7_0;
	wire w_dff_A_NVkVw5Rr0_0;
	wire w_dff_A_9kPS5u6Z9_0;
	wire w_dff_A_cOrKHC8r7_0;
	wire w_dff_B_ALmpcn5E2_0;
	wire w_dff_B_8DMOOf4i3_0;
	wire w_dff_B_m293t9WZ8_0;
	wire w_dff_B_gmoTMHaR0_0;
	wire w_dff_B_d5sNZA4I3_0;
	wire w_dff_B_IDfMCid82_0;
	wire w_dff_B_3MDwyOK57_0;
	wire w_dff_B_fuApnOfa2_0;
	wire w_dff_A_zcwsYSNy8_0;
	wire w_dff_A_lLbhIJXG0_0;
	wire w_dff_A_pM3KtXqT8_0;
	wire w_dff_A_ps7QqfkW5_0;
	wire w_dff_A_z7tTAFy69_0;
	wire w_dff_A_No7cUPur3_0;
	wire w_dff_A_PTQffy812_0;
	wire w_dff_A_6lDzlWRP6_0;
	wire w_dff_A_LwVKvSsc3_0;
	wire w_dff_A_VcZ0ObV67_1;
	wire w_dff_B_DeBhIout9_0;
	wire w_dff_B_lV3ChrZN8_0;
	wire w_dff_B_xZ08vA4y3_2;
	wire w_dff_B_WDEbrLem7_2;
	wire w_dff_A_fzbjfxrA9_0;
	wire w_dff_A_479Mr7cO0_0;
	wire w_dff_A_W3X3aebx9_0;
	wire w_dff_A_mm6HwVJP0_0;
	wire w_dff_B_D5js8nOw4_0;
	wire w_dff_B_1N5R0yCL3_0;
	wire w_dff_B_0K0C5rfL1_2;
	wire w_dff_B_0BNgGgMg3_2;
	wire w_dff_A_cm1WQzw24_0;
	wire w_dff_A_AxAcsGCx7_0;
	wire w_dff_A_UmwWKvEW7_0;
	wire w_dff_A_1rQxkaMZ6_0;
	wire w_dff_A_zXQNcWHq8_0;
	wire w_dff_A_LZhMNDa49_0;
	wire w_dff_A_IYbuSqnC5_0;
	wire w_dff_A_hTIxALdH9_0;
	wire w_dff_A_MKUfhvux9_0;
	wire w_dff_A_2mCGjD1i9_0;
	wire w_dff_A_QL5ApbaD7_0;
	wire w_dff_A_Gz8E25yi4_0;
	wire w_dff_A_iuTt8jDK2_0;
	wire w_dff_A_4Px20A4r9_0;
	wire w_dff_A_iK6pO9725_0;
	wire w_dff_A_BLNwJD364_0;
	wire w_dff_A_GcFNFohd4_1;
	wire w_dff_A_GipSjDUt4_1;
	wire w_dff_A_OP4lTLMV3_1;
	wire w_dff_A_qtJnsGNi4_1;
	wire w_dff_A_q2fnkuVw8_2;
	wire w_dff_A_batIeYWG1_2;
	wire w_dff_A_OINP2Htl1_2;
	wire w_dff_A_f7oh9e0H0_2;
	wire w_dff_A_7qcirIbk1_2;
	wire w_dff_A_NZAOmBEF5_2;
	wire w_dff_A_Z41uG3Qb5_2;
	wire w_dff_A_dct5lZS76_2;
	wire w_dff_A_6B2059224_2;
	wire w_dff_A_kTiYQC3z8_2;
	wire w_dff_A_1G46lzN70_2;
	wire w_dff_A_AR6PB7eS3_2;
	wire w_dff_B_3C2QXZfv3_0;
	wire w_dff_B_rnocEosP8_0;
	wire w_dff_B_77YsmIWU1_2;
	wire w_dff_B_sKxW7ouH5_2;
	wire w_dff_A_wILlbT7T3_2;
	wire w_dff_A_4YWfzSay5_2;
	wire w_dff_A_Kne2JWyF3_2;
	wire w_dff_A_6MKETmv02_2;
	wire w_dff_A_BFa9jBAm4_2;
	wire w_dff_A_UZhSkQ3u9_2;
	wire w_dff_A_QcSwRD9w2_2;
	wire w_dff_A_zFfFWEtR2_2;
	wire w_dff_A_yICARhwM9_2;
	wire w_dff_A_SW4xabWb7_2;
	wire w_dff_A_rpso9bRS2_2;
	wire w_dff_A_gRtxQXhT5_2;
	wire w_dff_A_txnbFa000_2;
	wire w_dff_A_xnCWaTuR7_2;
	wire w_dff_A_Ao79kSAN0_2;
	wire w_dff_B_KhfQAqlt3_0;
	wire w_dff_B_3uEs4dVE0_0;
	wire w_dff_B_oNNov6Cs0_3;
	wire w_dff_B_syGTL4xv9_3;
	wire w_dff_A_iL4NUDBV5_0;
	wire w_dff_A_kb6YfBSF5_0;
	wire w_dff_A_bUkzMEKL9_0;
	wire w_dff_A_7k2u0Uhk4_0;
	wire w_dff_A_mBGChZA09_2;
	wire w_dff_A_KB6PSNHp2_2;
	wire w_dff_B_gkRoOqZ43_0;
	wire w_dff_A_FdM5IzSU3_0;
	wire w_dff_A_yGaO7Vih8_0;
	wire w_dff_A_VMS3oj4g6_0;
	wire w_dff_A_d8qwEVrX0_1;
	wire w_dff_B_yVkI5nMr4_2;
	wire w_dff_B_YAXYqcGI0_2;
	wire w_dff_A_u6ht5Zzm1_0;
	wire w_dff_A_fPsIodG79_0;
	wire w_dff_A_soUu5tBA0_0;
	wire w_dff_A_j7vDye4R5_0;
	wire w_dff_B_6qNqKJ7I7_0;
	wire w_dff_B_zhQ5zoaN3_0;
	wire w_dff_B_oZxpILHP5_0;
	wire w_dff_B_eqNB2x3B1_0;
	wire w_dff_A_pf5blDt83_0;
	wire w_dff_A_GJmzwBgT8_0;
	wire w_dff_A_j8v0MkH30_0;
	wire w_dff_A_ugtOsKZg0_0;
	wire w_dff_A_GOtlVnN46_0;
	wire w_dff_B_j2k8mZZE5_1;
	wire w_dff_B_v4dk76pM1_1;
	wire w_dff_B_INxAodTD2_1;
	wire w_dff_B_3EeUhV7m3_1;
	wire w_dff_B_4KCJDPpx6_1;
	wire w_dff_B_YYMfaYUU9_1;
	wire w_dff_B_bU2JFqUT9_1;
	wire w_dff_B_DTSOZ4kH2_0;
	wire w_dff_B_HVTNJEOF6_0;
	wire w_dff_B_SnIFAloN7_0;
	wire w_dff_B_6UuhMnFy3_0;
	wire w_dff_B_6h0p151i4_0;
	wire w_dff_B_g93XN7Hd9_0;
	wire w_dff_B_Cd0jMb9i0_0;
	wire w_dff_A_0tNitACA4_0;
	wire w_dff_A_NqvdE97N4_0;
	wire w_dff_A_V0ljnoLg8_0;
	wire w_dff_A_ccNtsWX08_0;
	wire w_dff_A_FIyJsI0G3_0;
	wire w_dff_A_xnYzgbV02_0;
	wire w_dff_A_5Z8h4EPz9_0;
	wire w_dff_A_DjpXitUl9_0;
	wire w_dff_A_JovB0lwN3_0;
	wire w_dff_A_E5K7alzc4_0;
	wire w_dff_A_KJ3vDEya8_0;
	wire w_dff_A_eheffV112_0;
	wire w_dff_A_joYyMP7n7_0;
	wire w_dff_A_KU3rHIqv9_0;
	wire w_dff_A_hB3e9Lal8_0;
	wire w_dff_A_czRxNlFA7_0;
	wire w_dff_A_xfECxXcF3_0;
	wire w_dff_A_PJSjd5ZO0_0;
	wire w_dff_A_EXpZaSpZ3_0;
	wire w_dff_A_R5aBBOiV2_0;
	wire w_dff_A_1GIilQCR3_0;
	wire w_dff_A_px7SGiXE3_0;
	wire w_dff_A_m3rSiGQ31_0;
	wire w_dff_A_suR2No9l5_0;
	wire w_dff_A_0NvkXn7P2_0;
	wire w_dff_A_Mk4ll8HJ2_0;
	wire w_dff_A_G0ExnXCE7_0;
	wire w_dff_A_niLYAnRN9_0;
	wire w_dff_A_BFIbBuJj1_0;
	wire w_dff_A_CmHLRX2u3_0;
	wire w_dff_A_CJ2XfhFk2_0;
	wire w_dff_A_VCRb9KBz1_0;
	wire w_dff_A_wh4rldlH9_0;
	wire w_dff_A_kusIEkBs1_0;
	wire w_dff_A_DpbZDXwP0_0;
	wire w_dff_A_lPdV6RPk9_0;
	wire w_dff_A_dDUxUmdE1_0;
	wire w_dff_A_mmuEb3QL8_0;
	wire w_dff_A_AhamDzMV9_0;
	wire w_dff_A_CscisU493_0;
	wire w_dff_A_vO6IatWr4_0;
	wire w_dff_A_rJFI9lK38_0;
	wire w_dff_A_qKcgb3jQ7_0;
	wire w_dff_A_gDjcuU4m7_0;
	wire w_dff_A_KfEs8R6r0_0;
	wire w_dff_A_kRLrKGtV7_0;
	wire w_dff_A_HiBM4pVC7_0;
	wire w_dff_A_EGetv3MI1_0;
	wire w_dff_A_cKy94sAX5_0;
	wire w_dff_A_tXHQJMnv0_0;
	wire w_dff_A_ZxbK0vmW0_0;
	wire w_dff_A_gMf7R9sU2_1;
	wire w_dff_A_D5fs9vIB1_1;
	wire w_dff_A_3K7rC5Qk6_1;
	wire w_dff_A_WiNWTh6M3_1;
	wire w_dff_A_AZaIBfQd3_1;
	wire w_dff_A_0gFLWxzC7_1;
	wire w_dff_A_ranaJklK5_1;
	wire w_dff_A_4FRVz7XB5_1;
	wire w_dff_A_jEvkwzsX6_1;
	wire w_dff_A_t6sEAL5Z8_1;
	wire w_dff_A_iwIUXNDC4_1;
	wire w_dff_A_MbKVSPC10_1;
	wire w_dff_A_hfE9EebZ0_1;
	wire w_dff_A_2LREpPro2_1;
	wire w_dff_A_GAxHeVLN5_1;
	wire w_dff_A_bvKcreuB4_1;
	wire w_dff_A_hIUtR8a03_1;
	wire w_dff_A_PBd0LuDz8_1;
	wire w_dff_A_RGme1VQO3_1;
	wire w_dff_B_uHLU5VDr0_0;
	wire w_dff_A_eAUesVzk7_1;
	wire w_dff_A_xFztVBjF1_1;
	wire w_dff_A_xmevM6pX6_1;
	wire w_dff_A_IjN4mPtd6_1;
	wire w_dff_A_5KN7Waln8_1;
	wire w_dff_A_oeUb5HEf1_1;
	wire w_dff_A_WgF7CZ8P1_1;
	wire w_dff_A_2VlzlvdJ3_1;
	wire w_dff_A_aeGU1Iix2_1;
	wire w_dff_A_t5iGKbeR6_1;
	wire w_dff_A_gx9i3qNR3_1;
	wire w_dff_A_6aVfz3u40_1;
	wire w_dff_A_DrolHScC2_1;
	wire w_dff_A_S4OE00AN7_1;
	wire w_dff_A_R9H01SW31_1;
	wire w_dff_A_n78vXkR71_1;
	wire w_dff_A_eagtifbf5_1;
	wire w_dff_A_DInUTTPn0_1;
	wire w_dff_A_dzkYWVGd4_1;
	wire w_dff_A_EvcAKS2p6_1;
	wire w_dff_A_9zWEW9xr4_1;
	wire w_dff_A_FDYHxj9q1_0;
	wire w_dff_A_YVjUeDoE8_0;
	wire w_dff_A_5gGa3kNr3_0;
	wire w_dff_A_VmzUsI6k4_2;
	wire w_dff_A_WJWqTm6j3_1;
	wire w_dff_A_GrQxdQNd2_2;
	wire w_dff_A_DvvVmoVy6_2;
	wire w_dff_B_H54XB8QL4_1;
	wire w_dff_B_kEK1mXdw5_1;
	wire w_dff_B_5dHBPNPx4_1;
	wire w_dff_B_mIULG2T30_1;
	wire w_dff_B_2zhiKpty8_1;
	wire w_dff_B_4A3Dnlax8_1;
	wire w_dff_B_pA6yzUWF7_1;
	wire w_dff_B_60QWl5sd9_1;
	wire w_dff_B_xqiXDl2v5_1;
	wire w_dff_B_ceOtUC3a3_1;
	wire w_dff_B_WPeyNfHw0_1;
	wire w_dff_B_ASHbUCWz7_1;
	wire w_dff_B_OKEBBw1v9_1;
	wire w_dff_B_xMBW8gtM9_1;
	wire w_dff_B_ez4oe8O89_1;
	wire w_dff_B_tP5QGGy90_1;
	wire w_dff_B_4Gm3sYUt8_1;
	wire w_dff_B_FUVbq3kE0_1;
	wire w_dff_B_82E0SqC84_1;
	wire w_dff_B_H0YLKs2Y6_1;
	wire w_dff_B_AMKVK5VG7_1;
	wire w_dff_B_79HMWNLb4_1;
	wire w_dff_B_nw132nbh3_1;
	wire w_dff_B_wwJVCGX44_1;
	wire w_dff_B_MkWhOmse4_1;
	wire w_dff_B_MjDQdwRa4_1;
	wire w_dff_B_1UGtU2pP1_1;
	wire w_dff_B_eYsFY6Dz2_1;
	wire w_dff_B_ldlJ2nWL0_1;
	wire w_dff_B_lxx2CanO3_1;
	wire w_dff_B_tmvJ6XVG7_1;
	wire w_dff_B_nGaZYB9h6_1;
	wire w_dff_B_9XJZ6PK16_0;
	wire w_dff_B_4stDTBS90_0;
	wire w_dff_A_g0sE4gYu5_1;
	wire w_dff_A_WG64xLY17_1;
	wire w_dff_A_sjwH9waE9_1;
	wire w_dff_A_Qzifh2BF2_1;
	wire w_dff_A_XyOJ4ZVF4_1;
	wire w_dff_A_KtsyxYg13_1;
	wire w_dff_A_Ed8GysSM6_1;
	wire w_dff_A_VkjFpfeo2_1;
	wire w_dff_A_L9MFRLub6_1;
	wire w_dff_A_t1OorFeT8_1;
	wire w_dff_A_pJKJ5JGS9_1;
	wire w_dff_B_AFVHb2Dm8_1;
	wire w_dff_B_VTOZJaWd5_1;
	wire w_dff_B_zMT5VBaP1_1;
	wire w_dff_B_Jmwo1Vpq5_1;
	wire w_dff_B_hIlveP8D7_1;
	wire w_dff_B_2yNwb2Rz4_1;
	wire w_dff_B_XKqHvp1z8_0;
	wire w_dff_A_KjU7AqUT0_1;
	wire w_dff_A_tLo5OXNk5_1;
	wire w_dff_A_5lvn2ewi5_1;
	wire w_dff_A_W1Q2ulZp0_1;
	wire w_dff_A_iO7mZrfs7_1;
	wire w_dff_A_Y5jRghTd6_1;
	wire w_dff_A_0WAxktpG4_1;
	wire w_dff_A_syDZq2026_1;
	wire w_dff_A_F77pSxzR3_1;
	wire w_dff_A_jLvMlcrl4_1;
	wire w_dff_A_JR4JKGp92_1;
	wire w_dff_A_vaUUkInl2_1;
	wire w_dff_B_donYkLVC3_2;
	wire w_dff_B_mbjCN1LT8_2;
	wire w_dff_B_IoS9XBZo6_2;
	wire w_dff_B_WdTyTBTI2_2;
	wire w_dff_B_p5naMZBK5_2;
	wire w_dff_B_jllnJNpC9_2;
	wire w_dff_B_2ZlPMjFp5_2;
	wire w_dff_B_4ORWPjYZ0_1;
	wire w_dff_B_IERriCYy9_0;
	wire w_dff_B_EjHF14WT6_0;
	wire w_dff_B_ornnWYyA2_1;
	wire w_dff_B_IDeAhHgO2_1;
	wire w_dff_B_86ioJiNl5_1;
	wire w_dff_B_DpYNnzbp2_1;
	wire w_dff_B_1DOt81Ad4_1;
	wire w_dff_B_sel0X8RR9_0;
	wire w_dff_A_FnpgA7eZ4_0;
	wire w_dff_A_Ng5qy9pI2_1;
	wire w_dff_A_kUyaWBU63_1;
	wire w_dff_A_lRVvlXKr1_1;
	wire w_dff_A_4BSE3NL41_1;
	wire w_dff_A_bHanTw4u7_1;
	wire w_dff_A_P3pamEE47_1;
	wire w_dff_A_5E4wL1zE3_1;
	wire w_dff_A_XixEvbBh8_1;
	wire w_dff_A_IynqEskC4_1;
	wire w_dff_A_0gA4mnx75_1;
	wire w_dff_B_vi9gKCrh7_0;
	wire w_dff_B_Pr4cRVXm5_0;
	wire w_dff_B_Eh2Rk16E7_0;
	wire w_dff_B_VkEavW1t2_0;
	wire w_dff_B_9ZpuAkHu2_0;
	wire w_dff_B_RjQZLPU06_0;
	wire w_dff_B_XX9PT8uf5_0;
	wire w_dff_A_CMDxxD1q7_2;
	wire w_dff_A_CCfkFeBt8_2;
	wire w_dff_A_4GL5I2FX7_2;
	wire w_dff_A_9C6nb4KK7_2;
	wire w_dff_A_CHLv29ha1_2;
	wire w_dff_A_27sUQoDV3_2;
	wire w_dff_A_I8542ZhQ6_2;
	wire w_dff_A_IGyUEtNS0_2;
	wire w_dff_A_opi42OKV6_1;
	wire w_dff_A_50Pk9rpa7_1;
	wire w_dff_A_h97gtSDy3_2;
	wire w_dff_A_KDwJqF2U7_2;
	wire w_dff_A_nyalX7Vu4_2;
	wire w_dff_A_EJWBJjO24_2;
	wire w_dff_A_kyC7fiAW9_2;
	wire w_dff_A_gSCgWGLe3_2;
	wire w_dff_A_UasxrxzM1_2;
	wire w_dff_A_3loQDpa12_2;
	wire w_dff_A_tJTwwsdY4_2;
	wire w_dff_A_RAC4MjRG2_2;
	wire w_dff_A_ihl4IpdQ5_2;
	wire w_dff_A_GMvBdxUO4_2;
	wire w_dff_B_OIKxCJxU6_1;
	wire w_dff_B_GJv8SWDd3_1;
	wire w_dff_B_xgc1Od2f3_1;
	wire w_dff_B_mm7fPUEe4_1;
	wire w_dff_B_2DsdV5O88_0;
	wire w_dff_A_x19YsS0i6_1;
	wire w_dff_B_SAlCeFYl0_2;
	wire w_dff_B_rFAGAFOx4_2;
	wire w_dff_A_fzKjvWig5_1;
	wire w_dff_A_HtvCpDy58_1;
	wire w_dff_A_Ns2WddQp2_1;
	wire w_dff_A_s7orHyME7_1;
	wire w_dff_A_9BI1CyFY4_1;
	wire w_dff_A_sKP7S97R2_1;
	wire w_dff_A_7MI3tEFm7_1;
	wire w_dff_A_lwZauxQ99_1;
	wire w_dff_A_W9Oe9Irk5_1;
	wire w_dff_A_nCU9MRR05_1;
	wire w_dff_A_hHJMPfl68_1;
	wire w_dff_A_UqO1TnTV9_1;
	wire w_dff_A_iGjyd2mM3_1;
	wire w_dff_A_fNXRIG3F4_1;
	wire w_dff_A_6qYis3IZ4_1;
	wire w_dff_A_GIqro3PQ5_1;
	wire w_dff_A_pvqZuXdk9_1;
	wire w_dff_A_TcSk9PEH7_1;
	wire w_dff_A_fIfmGo6g3_1;
	wire w_dff_A_ck0iszft9_1;
	wire w_dff_B_PcBIj1gP7_1;
	wire w_dff_B_4FoRgvuD6_0;
	wire w_dff_A_AqZSHEOy8_1;
	wire w_dff_A_4E7K3r0y5_1;
	wire w_dff_A_EiVtXFOz7_2;
	wire w_dff_A_JIK2jnnq1_2;
	wire w_dff_A_lAvt5qLZ3_1;
	wire w_dff_A_KCyLF0xG5_1;
	wire w_dff_A_3jSymNVW0_1;
	wire w_dff_A_8eBzixrq7_1;
	wire w_dff_A_DgDAJlvf3_2;
	wire w_dff_A_Iuxr2gKJ8_2;
	wire w_dff_A_pE32UJ6Y0_0;
	wire w_dff_A_5dgnjyY68_0;
	wire w_dff_B_JGSCKHOj3_2;
	wire w_dff_B_fzUH6Gwg3_1;
	wire w_dff_B_AJSqunPQ4_0;
	wire w_dff_A_EhA8q3zh6_1;
	wire w_dff_A_rPxpNk2v5_1;
	wire w_dff_A_6cgcbzJM4_2;
	wire w_dff_A_t8sJnWpR2_2;
	wire w_dff_A_fDzA0mv00_0;
	wire w_dff_A_o5zNdw3o6_0;
	wire w_dff_A_Q9lzvkjn7_0;
	wire w_dff_A_gCT6V1oP9_0;
	wire w_dff_A_o1KJXdOF0_0;
	wire w_dff_A_DSPztC9M3_0;
	wire w_dff_A_4Jyj9n3U1_0;
	wire w_dff_A_v7Y8xzsW1_0;
	wire w_dff_A_EZo0lXF13_0;
	wire w_dff_A_wUx0yTa09_0;
	wire w_dff_A_UzABrpJR6_0;
	wire w_dff_A_EYlpZPJq4_0;
	wire w_dff_A_egm8n0ej7_1;
	wire w_dff_B_yAKEZt6k3_1;
	wire w_dff_B_84iRtvq86_0;
	wire w_dff_A_0iBeJp9B8_1;
	wire w_dff_A_T9rOa2NS6_1;
	wire w_dff_A_6gtT0VQr7_2;
	wire w_dff_A_bcAtzUew4_2;
	wire w_dff_A_XB3GkqvB2_1;
	wire w_dff_A_r1Eae4on4_1;
	wire w_dff_A_BKMaKKir6_1;
	wire w_dff_A_VgHUHFeN3_1;
	wire w_dff_A_5nLHnB6C4_1;
	wire w_dff_B_nM3yZrsY8_1;
	wire w_dff_B_lUP2YVfW1_1;
	wire w_dff_B_B0NN0BAE9_1;
	wire w_dff_B_FX4kO5pn5_1;
	wire w_dff_B_G3a7yDBn7_1;
	wire w_dff_B_ReywKQIc6_1;
	wire w_dff_B_4c1rMKSY1_1;
	wire w_dff_B_kVQlZe7Y6_1;
	wire w_dff_B_VV4ipEa63_1;
	wire w_dff_B_NU9PT9Tc7_1;
	wire w_dff_B_7bPW3G278_1;
	wire w_dff_A_u77RTt2G0_1;
	wire w_dff_A_qgFMoNKm5_1;
	wire w_dff_A_XTAzeNi84_1;
	wire w_dff_A_0LzmGCC08_1;
	wire w_dff_A_5qzCAV2S8_1;
	wire w_dff_B_uW98lKMF6_1;
	wire w_dff_B_wJZHFkYc5_1;
	wire w_dff_B_RSpnqIE92_1;
	wire w_dff_A_GsSCDuzU2_1;
	wire w_dff_A_Lh6XoaEJ7_1;
	wire w_dff_A_vznTILIU3_1;
	wire w_dff_A_DMkJGa9p8_1;
	wire w_dff_A_xvBOGYZI5_1;
	wire w_dff_A_pH4My2IA7_1;
	wire w_dff_A_NdcOEkCb6_0;
	wire w_dff_A_6U1UqLW16_0;
	wire w_dff_A_xxOlJ3CW8_0;
	wire w_dff_A_U0hXA5h91_0;
	wire w_dff_A_JE9mLRAe8_2;
	wire w_dff_A_YOXyXLCP3_2;
	wire w_dff_A_QXQ9j92N2_2;
	wire w_dff_A_zIdw6yhx1_2;
	wire w_dff_A_L8v9zKPK0_1;
	wire w_dff_B_BpLrxlZp9_2;
	wire w_dff_A_zzibIUZP2_0;
	wire w_dff_A_WeQLK4OR9_0;
	wire w_dff_B_KV71pfwJ2_2;
	wire w_dff_B_pMrX8p496_2;
	wire w_dff_B_EYruc3vf3_2;
	wire w_dff_B_Kmrt3sfJ7_2;
	wire w_dff_B_VVfKKsny1_0;
	wire w_dff_B_vqSnrWII8_0;
	wire w_dff_B_2GNWMdUI1_0;
	wire w_dff_A_u1xDV8Vf1_0;
	wire w_dff_A_iRiUx5rP2_0;
	wire w_dff_A_0siaQzSh6_0;
	wire w_dff_A_tOfU8hJU1_0;
	wire w_dff_A_6t7b2Fct8_0;
	wire w_dff_A_5pYyDCjl1_0;
	wire w_dff_A_F5L11Xlj2_0;
	wire w_dff_A_ajUlbdyL5_0;
	wire w_dff_A_ldFYse3U6_0;
	wire w_dff_A_8uUtDvTF5_0;
	wire w_dff_A_tTHkCHta4_0;
	wire w_dff_A_kwfy8KXb7_0;
	wire w_dff_A_kqH5AU9u5_0;
	wire w_dff_A_qEgsXavU1_0;
	wire w_dff_A_PXkeGuLe9_0;
	wire w_dff_A_fdpewNTe8_1;
	wire w_dff_A_WvhCOYmd0_1;
	wire w_dff_A_tVXKqJGB9_1;
	wire w_dff_A_EP0sGnie1_2;
	wire w_dff_A_hKmYyrgv9_2;
	wire w_dff_A_p77vMcCr0_2;
	wire w_dff_A_ojFg92OK0_2;
	wire w_dff_A_VvOpbdxn0_2;
	wire w_dff_A_ENMNb7XV9_2;
	wire w_dff_A_NwdEVlzB8_2;
	wire w_dff_B_I7HteV6h8_1;
	wire w_dff_B_EYX6X5V06_0;
	wire w_dff_A_TDelmwbm7_0;
	wire w_dff_A_okpQ7hcA6_0;
	wire w_dff_A_o0jEiWOW7_0;
	wire w_dff_A_F6zSoCrM3_0;
	wire w_dff_A_UMlRGQE61_1;
	wire w_dff_A_Ar2t3l8F8_1;
	wire w_dff_A_ZtNUuRnv6_2;
	wire w_dff_A_3o7m0Os36_2;
	wire w_dff_A_k7JJI3cr8_2;
	wire w_dff_A_atQfae210_2;
	wire w_dff_A_1iOGvwmI5_2;
	wire w_dff_A_sdAdEEBW6_2;
	wire w_dff_A_gk9VVL3Z7_2;
	wire w_dff_A_CUvmDf5J0_2;
	wire w_dff_A_abvw01o64_2;
	wire w_dff_A_KGEqSJ7R2_2;
	wire w_dff_B_QMTRnMAr5_1;
	wire w_dff_B_Y2u8jKVw1_0;
	wire w_dff_B_T69QBFzD0_3;
	wire w_dff_B_QCLCXMcC4_3;
	wire w_dff_A_TnqZL3N03_0;
	wire w_dff_A_3WBdhEWs9_0;
	wire w_dff_A_vmr5aENK6_0;
	wire w_dff_A_R0cohlg94_0;
	wire w_dff_A_azehETn11_2;
	wire w_dff_A_sclD5zdd4_2;
	wire w_dff_A_Iu8Av3AH3_2;
	wire w_dff_B_wSeJvHvY2_1;
	wire w_dff_B_Bzm4aaA47_0;
	wire w_dff_B_G4bOJIy79_2;
	wire w_dff_B_jr5IL4iN8_2;
	wire w_dff_A_yoOFCVWY1_0;
	wire w_dff_A_1ETaXjQF7_0;
	wire w_dff_A_70SR8ZAK3_0;
	wire w_dff_A_YppMUfdg6_0;
	wire w_dff_A_4OlQz9K68_0;
	wire w_dff_A_o4THdZ0n0_0;
	wire w_dff_A_plzDQIpw4_0;
	wire w_dff_A_b5VbxXny3_0;
	wire w_dff_A_GO7S0n6C9_1;
	wire w_dff_A_sqp9Njm17_1;
	wire w_dff_A_ayvScaaT2_1;
	wire w_dff_A_dfPLcqln1_0;
	wire w_dff_A_kXBd5JXl6_0;
	wire w_dff_A_mjnJcMV75_0;
	wire w_dff_A_ttlRrIgr0_0;
	wire w_dff_A_0szJyxE99_0;
	wire w_dff_A_WJQMmuie9_0;
	wire w_dff_A_NBaBoVcZ7_0;
	wire w_dff_A_IiN5JI5s8_0;
	wire w_dff_A_W5tLDX4L7_0;
	wire w_dff_A_7zf17ZJ46_0;
	wire w_dff_B_XJUEGaX61_2;
	wire w_dff_B_cteXpGLd6_2;
	wire w_dff_A_rYZP6bhc0_0;
	wire w_dff_A_lXbV1seQ8_0;
	wire w_dff_A_OloIHzAR1_0;
	wire w_dff_A_T2HkbbHv0_0;
	wire w_dff_A_GTbnRU559_0;
	wire w_dff_A_mtPxmBZR7_0;
	wire w_dff_A_p7UtFTKd6_1;
	wire w_dff_A_zUKcF8oA4_1;
	wire w_dff_A_IxiQpLBq7_1;
	wire w_dff_B_5hU4vHiZ8_1;
	wire w_dff_B_0QEtDJod2_0;
	wire w_dff_A_bIhfmbo90_0;
	wire w_dff_A_mdiprYfS9_0;
	wire w_dff_A_mb7C1QHa8_0;
	wire w_dff_A_J2qPaUXQ6_0;
	wire w_dff_A_xdlzvDjW9_0;
	wire w_dff_A_x71sLdCq3_2;
	wire w_dff_B_JjtPmCHB3_1;
	wire w_dff_B_r7ZZahyA5_0;
	wire w_dff_B_vh3Uguei7_2;
	wire w_dff_B_2P58I5eT7_2;
	wire w_dff_A_vIvxKYgN7_0;
	wire w_dff_A_U9HEbJgo5_0;
	wire w_dff_A_K48xyCr10_0;
	wire w_dff_A_6pxG1Fq52_0;
	wire w_dff_A_5EbDisAo9_0;
	wire w_dff_A_IlnJLqiF5_0;
	wire w_dff_A_TzbzIG4M8_1;
	wire w_dff_A_9LNjiWNT4_1;
	wire w_dff_A_TO5rHO6z6_1;
	wire w_dff_A_xb40rgLK8_1;
	wire w_dff_A_3bsSzGkA5_1;
	wire w_dff_A_OL3a0SAZ9_1;
	wire w_dff_A_LqKGtasU1_1;
	wire w_dff_A_NdTm2IRH8_1;
	wire w_dff_A_UIODt7P69_1;
	wire w_dff_A_KJ01KZjo3_1;
	wire w_dff_A_HpI7Zu6e0_1;
	wire w_dff_A_nW4mItQv2_1;
	wire w_dff_B_Uq25joIQ0_1;
	wire w_dff_B_RbOHchf68_0;
	wire w_dff_B_Th2dA3IE6_2;
	wire w_dff_B_clWffWiI2_2;
	wire w_dff_A_232Wcgk02_0;
	wire w_dff_A_h4ekmAyz2_0;
	wire w_dff_A_MAUrdrhs9_0;
	wire w_dff_A_vK1SaVCu5_0;
	wire w_dff_B_zr9TvNSk1_1;
	wire w_dff_B_Wfe7UT0x5_1;
	wire w_dff_B_KqnuhGgy5_1;
	wire w_dff_B_kmOdv2Jc1_1;
	wire w_dff_B_2iXF6qVS1_1;
	wire w_dff_B_VR6pvUXp8_1;
	wire w_dff_B_Z8lwB16C9_1;
	wire w_dff_B_aMHTsw7C1_1;
	wire w_dff_B_NpLUcPD67_1;
	wire w_dff_B_KBuj21bs4_1;
	wire w_dff_B_VzJehx210_1;
	wire w_dff_B_U7wBcD9C1_1;
	wire w_dff_B_iXzO8Qrp3_1;
	wire w_dff_B_KiFOFoT63_1;
	wire w_dff_B_3LGbg9YE5_1;
	wire w_dff_B_YN8G514S2_1;
	wire w_dff_B_Ot2uxS2b8_1;
	wire w_dff_B_LqYwp0DK4_1;
	wire w_dff_B_cC0B5eQI6_0;
	wire w_dff_B_mHSsPA474_1;
	wire w_dff_B_FqaGOYoO0_1;
	wire w_dff_B_29kOIiyV1_0;
	wire w_dff_B_AOo5QAEB4_0;
	wire w_dff_B_4WpU1ehT3_0;
	wire w_dff_B_fvd44txS3_0;
	wire w_dff_B_H5omkcwW9_0;
	wire w_dff_B_ryHRoTbl5_0;
	wire w_dff_B_tUAfxP7n4_0;
	wire w_dff_B_H0K3lUBb0_1;
	wire w_dff_B_xleab02x0_1;
	wire w_dff_B_tuMJqVnd7_1;
	wire w_dff_B_2bGQ9w4O4_1;
	wire w_dff_B_FuQFIgH88_1;
	wire w_dff_B_CIsA5jLb0_1;
	wire w_dff_B_hWdk9Lp90_1;
	wire w_dff_B_v2w6Y5368_1;
	wire w_dff_B_BaY2riKL9_1;
	wire w_dff_A_I1cbKSU18_1;
	wire w_dff_A_qiZJRdEy0_1;
	wire w_dff_A_riHYd6Xt7_1;
	wire w_dff_A_ybqhCZ7i9_1;
	wire w_dff_B_yaGAndz76_1;
	wire w_dff_A_qRjD17OP6_0;
	wire w_dff_A_dTfLmEGw5_0;
	wire w_dff_A_azqyXgUa4_0;
	wire w_dff_B_78qQyTrY1_2;
	wire w_dff_B_zFxoyLqs4_2;
	wire w_dff_B_yKeTjvzk6_2;
	wire w_dff_B_pfOlVf9R1_2;
	wire w_dff_A_T06DSO181_1;
	wire w_dff_A_bUccLvCp0_1;
	wire w_dff_A_4DWiGXIG0_1;
	wire w_dff_B_OGgUC0wS8_1;
	wire w_dff_B_REeW9gvT5_1;
	wire w_dff_B_psoXIpxT9_0;
	wire w_dff_B_jxRLmfFY1_0;
	wire w_dff_A_ZJHbP3dP6_0;
	wire w_dff_A_CBVuSnub1_0;
	wire w_dff_A_ZPEdoOs90_0;
	wire w_dff_A_vpVwBZGG7_1;
	wire w_dff_B_rjvqatEd1_1;
	wire w_dff_B_wHCiczz55_1;
	wire w_dff_B_JRcaNep85_1;
	wire w_dff_B_QUIsBXBh1_1;
	wire w_dff_B_j4SVgvbl0_1;
	wire w_dff_B_4Wj5yp2j5_1;
	wire w_dff_B_qAlmacbT0_1;
	wire w_dff_B_Lzk0vi2H7_1;
	wire w_dff_B_zd0yajDr0_1;
	wire w_dff_B_lbznyI1u1_1;
	wire w_dff_A_9qZgzsNs9_0;
	wire w_dff_A_TdBdHRL18_0;
	wire w_dff_A_9yFEB4Tk7_0;
	wire w_dff_A_6Yzdt3Ak2_0;
	wire w_dff_B_o9uY41Ac7_1;
	wire w_dff_A_cV1ghasb7_1;
	wire w_dff_A_MK79zHne4_0;
	wire w_dff_A_mqnS2Z4X2_0;
	wire w_dff_A_Pbera6bC7_0;
	wire w_dff_A_MV8HZdIY7_1;
	wire w_dff_A_wEcAMxBO0_1;
	wire w_dff_A_r4uRtzhq8_1;
	wire w_dff_A_kNbcT2hR0_0;
	wire w_dff_A_BXHabmH63_0;
	wire w_dff_A_CszolQZC5_0;
	wire w_dff_A_7BAqe4RH3_0;
	wire w_dff_A_sOHOWnrF9_0;
	wire w_dff_B_qH8YMZAq3_0;
	wire w_dff_A_zgO2fUiT9_1;
	wire w_dff_A_5wPFBUs39_1;
	wire w_dff_A_YU2PxwHh9_1;
	wire w_dff_A_u9w86PM44_2;
	wire w_dff_A_1fPZMeRr7_2;
	wire w_dff_B_P9QBsc5k9_0;
	wire w_dff_A_8VN8W2Jp5_0;
	wire w_dff_A_FFoxzIYb8_0;
	wire w_dff_A_fUSrVCF72_0;
	wire w_dff_A_UZkBPwWu9_1;
	wire w_dff_A_BRbsPw8B7_1;
	wire w_dff_A_SXnMlaJE4_1;
	wire w_dff_B_vA4D5r9z7_0;
	wire w_dff_B_wtTzXQZ68_0;
	wire w_dff_B_5MKJui9C7_0;
	wire w_dff_B_iWkXe2AJ4_0;
	wire w_dff_A_BxX42A2O3_1;
	wire w_dff_A_5gRjoGy61_1;
	wire w_dff_A_0WhToFMW5_1;
	wire w_dff_A_fDmLV9JP5_1;
	wire w_dff_A_wWhXJe5g4_1;
	wire w_dff_A_oqZruxcR8_1;
	wire w_dff_A_PKKRSAtR4_1;
	wire w_dff_A_DOXs29d90_1;
	wire w_dff_A_X1w6X3UH9_1;
	wire w_dff_A_oJGc6wik0_1;
	wire w_dff_A_tvCdJFBR8_1;
	wire w_dff_A_bMRYvsgy9_1;
	wire w_dff_B_KeNprzu58_0;
	wire w_dff_A_sTYy0b9H1_1;
	wire w_dff_A_sBgJxJKt1_1;
	wire w_dff_B_5GHdNSKJ6_1;
	wire w_dff_A_Oh3JpdHS7_0;
	wire w_dff_A_6M5Ju3np0_0;
	wire w_dff_A_5vS2KP6j3_0;
	wire w_dff_A_uuWTafWp4_0;
	wire w_dff_A_iqDMWr1G8_0;
	wire w_dff_A_2ORK7MJ96_0;
	wire w_dff_A_ruTERdd65_0;
	wire w_dff_A_PFrRtPz72_0;
	wire w_dff_A_v76VSXqZ6_1;
	wire w_dff_A_JAoynUOq8_1;
	wire w_dff_A_rShiufyc4_1;
	wire w_dff_A_u95AvtUA5_1;
	wire w_dff_A_Mu6B6EbU7_1;
	wire w_dff_A_8TRro6Rh2_0;
	wire w_dff_A_74cnW4016_0;
	wire w_dff_A_qPeJQYRD1_0;
	wire w_dff_A_9H4knwf08_1;
	wire w_dff_A_AIM5S5t53_0;
	wire w_dff_A_5gSkhRnC7_0;
	wire w_dff_A_TbXBDE7v1_2;
	wire w_dff_A_68KSUdat4_2;
	wire w_dff_A_B6Cf6Acw1_2;
	wire w_dff_A_WFaEeLe79_2;
	wire w_dff_A_8oLxctnW1_2;
	wire w_dff_A_G9vcx2wh9_2;
	wire w_dff_A_36dz6SZj6_2;
	wire w_dff_A_PWZDMPJl4_2;
	wire w_dff_A_WWKtgBrA9_2;
	wire w_dff_A_b2eYmO4R5_2;
	wire w_dff_B_KidPtzUp6_3;
	wire w_dff_A_wN9Pvajd7_2;
	wire w_dff_A_VW7Yj6298_2;
	wire w_dff_A_DknvD8Cx1_1;
	wire w_dff_A_hy19a9jk7_1;
	wire w_dff_A_UK6liytN6_1;
	wire w_dff_A_Y35dsLT03_1;
	wire w_dff_A_NW0XW22D6_1;
	wire w_dff_A_5hMSZaFC4_1;
	wire w_dff_A_JmylGvGX8_1;
	wire w_dff_A_GRIDOSq39_1;
	wire w_dff_A_0cOZA6cA9_1;
	wire w_dff_A_7gf8DVbR1_1;
	wire w_dff_A_fn373POl2_2;
	wire w_dff_A_Agm25rVm7_2;
	wire w_dff_A_QTlFZtkZ7_2;
	wire w_dff_B_ijgckosu9_1;
	wire w_dff_B_sTsRkrCo0_1;
	wire w_dff_A_0fReXTFg6_0;
	wire w_dff_A_kVT3uzCz5_0;
	wire w_dff_A_MeHNMQtc8_0;
	wire w_dff_A_uSWqszjk6_0;
	wire w_dff_A_sK9IWy2v7_0;
	wire w_dff_A_MSVHLPQs9_1;
	wire w_dff_A_ZxAd4Hdj4_2;
	wire w_dff_A_xb6S6qui0_2;
	wire w_dff_A_nMiP9VN05_2;
	wire w_dff_A_fNiV9ITl2_2;
	wire w_dff_A_oaivMi756_2;
	wire w_dff_B_26IBZNyP1_3;
	wire w_dff_A_5Sf6yYef6_0;
	wire w_dff_A_DItjsZtr7_0;
	wire w_dff_A_aE5bhzcy6_0;
	wire w_dff_A_VMwgvIR75_0;
	wire w_dff_A_1JWV0Pyl7_1;
	wire w_dff_A_NVapzCBn3_1;
	wire w_dff_A_iUgl4et14_0;
	wire w_dff_A_7xgMrx8f8_0;
	wire w_dff_A_L8oEP3pi9_0;
	wire w_dff_A_CM5uF7Q79_0;
	wire w_dff_A_jQm4POQd1_0;
	wire w_dff_A_ueMveMMH3_0;
	wire w_dff_A_7njmmzcU3_0;
	wire w_dff_A_JivydptM7_0;
	wire w_dff_A_FHod2HfN7_0;
	wire w_dff_A_n9lY1H8r0_0;
	wire w_dff_A_DsbOikcy1_0;
	wire w_dff_A_QLd0u7Pk2_0;
	wire w_dff_A_t2vvxLIv2_2;
	wire w_dff_B_P9oTzFiG0_3;
	wire w_dff_B_pLDP2Vqt9_3;
	wire w_dff_B_TBNi1hV02_3;
	wire w_dff_B_mLOxX17m9_3;
	wire w_dff_A_X2hJZbNH9_1;
	wire w_dff_A_rTCYYuTb9_1;
	wire w_dff_A_MJsQ6nGm6_1;
	wire w_dff_A_BpQsFthV1_1;
	wire w_dff_A_ms5Q6tOQ7_1;
	wire w_dff_A_9PM9D7hK7_1;
	wire w_dff_A_WKlATLgI7_1;
	wire w_dff_A_fy6nSdI54_1;
	wire w_dff_A_PgvoQJuA2_1;
	wire w_dff_A_UdbUjPSL4_1;
	wire w_dff_A_VpOZSvnH0_1;
	wire w_dff_A_PRsLHwbW7_1;
	wire w_dff_A_VDwri5zt0_1;
	wire w_dff_A_6LaLYoZz7_1;
	wire w_dff_A_XDKhkYet6_1;
	wire w_dff_A_DLlCpuQU8_1;
	wire w_dff_A_Vvn0hPCn1_1;
	wire w_dff_A_YOC4rDdX5_1;
	wire w_dff_A_2bAkTEUW4_1;
	wire w_dff_A_d505jNZO2_1;
	wire w_dff_A_9M9WJaAl2_2;
	wire w_dff_A_vPudiIHb7_2;
	wire w_dff_A_nuR6vZS55_2;
	wire w_dff_A_u6pCXeVY1_2;
	wire w_dff_A_FlXCStQ04_2;
	wire w_dff_A_CGzIPUJQ0_2;
	wire w_dff_A_fptldo2Z1_1;
	wire w_dff_A_UfqrjIig3_2;
	wire w_dff_A_XjEUdPLg8_2;
	wire w_dff_A_8zOw0JFN9_2;
	wire w_dff_A_ujmd7dth2_1;
	wire w_dff_A_fxhrM4H85_2;
	wire w_dff_A_QCnVwtnx0_2;
	wire w_dff_A_NsVQY6dY5_0;
	wire w_dff_A_tlg9K5ml4_0;
	wire w_dff_A_uFNboZ7w4_0;
	wire w_dff_A_KIbxWG680_1;
	wire w_dff_A_nsY4tZgM7_1;
	wire w_dff_A_T4oDNzeA1_1;
	wire w_dff_A_lAUA7D2V6_1;
	wire w_dff_A_E1HN2sYi3_1;
	wire w_dff_A_gi09h5j40_1;
	wire w_dff_A_AiXPINR31_1;
	wire w_dff_A_c0J9rYi81_1;
	wire w_dff_A_wDZaEiJY1_1;
	wire w_dff_A_YFnBr3dz8_1;
	wire w_dff_A_rLEOKtgO7_1;
	wire w_dff_A_Y7XVqhIw2_1;
	wire w_dff_A_2xgicKFQ5_1;
	wire w_dff_A_k9uy9nRV1_1;
	wire w_dff_A_lxXH7riZ8_2;
	wire w_dff_A_isE6yyPm5_2;
	wire w_dff_A_yXdKgWiP7_2;
	wire w_dff_A_JeDlUWyh1_2;
	wire w_dff_A_pzV3NkDf7_2;
	wire w_dff_A_Y5zX2Jn48_1;
	wire w_dff_A_Awt1ZS5b6_1;
	wire w_dff_A_f4GZOwov5_1;
	wire w_dff_A_MjfUwtZn7_1;
	wire w_dff_A_QzaHcTNw8_1;
	wire w_dff_A_xNRUv05R1_1;
	wire w_dff_A_zfdkBFJC6_1;
	wire w_dff_A_qxygZq8W6_1;
	wire w_dff_A_viZejYLv6_1;
	wire w_dff_A_xBUmBKqi3_1;
	wire w_dff_A_aPEOWLYQ7_1;
	wire w_dff_A_sCnlMVHi9_2;
	wire w_dff_A_O1OWSXsT9_1;
	wire w_dff_A_O09Sv88N4_1;
	wire w_dff_A_myC7Op7m9_1;
	wire w_dff_A_lVTS1oef4_1;
	wire w_dff_A_1F408bzs9_1;
	wire w_dff_A_OvmsPZXt0_1;
	wire w_dff_A_kGUs8Ygl7_2;
	wire w_dff_A_2PKsHjju1_2;
	wire w_dff_A_O3pZ11if4_2;
	wire w_dff_A_G4vODcwN8_2;
	wire w_dff_A_BfEahovQ1_2;
	wire w_dff_A_IPFhCnFv0_2;
	wire w_dff_A_bUV5ZSHt7_2;
	wire w_dff_A_nvfLFF5L2_2;
	wire w_dff_A_siTTxv4V7_1;
	wire w_dff_A_7OWMYmKc6_1;
	wire w_dff_A_rkwUqV5s2_1;
	wire w_dff_A_A0c8EOMR5_0;
	wire w_dff_A_oT3PokxN3_0;
	wire w_dff_A_WhROGiIe9_0;
	wire w_dff_A_9SzzS9C42_2;
	wire w_dff_A_9IeOG2S09_2;
	wire w_dff_A_heDmG2sM6_2;
	wire w_dff_B_IDWVY7Qp0_0;
	wire w_dff_B_HKpF9qpd8_0;
	wire w_dff_B_glvbTKBU9_0;
	wire w_dff_B_M0X3wcWY0_0;
	wire w_dff_B_XYYkBOti0_0;
	wire w_dff_A_bxT6hRH78_0;
	wire w_dff_A_n78Njfyl6_0;
	wire w_dff_A_c3nTc5gs1_0;
	wire w_dff_A_J4TEJD776_0;
	wire w_dff_A_N99NFegW8_0;
	wire w_dff_A_srNQeTzb1_2;
	wire w_dff_A_O97I3AvY0_2;
	wire w_dff_A_epmZ90cf7_2;
	wire w_dff_A_ORIrRChN2_2;
	wire w_dff_A_nkNKKBf63_2;
	wire w_dff_A_ua17eETB6_2;
	wire w_dff_A_Z8dSX2lB7_2;
	wire w_dff_A_N77G8Ucv9_2;
	wire w_dff_A_7gOmAGjr3_2;
	wire w_dff_A_ZIz1Wk376_2;
	wire w_dff_A_a9jK7E3F3_2;
	wire w_dff_A_jj0BgXic4_2;
	wire w_dff_A_M2sNt5aJ0_2;
	wire w_dff_A_SuogiHgF1_2;
	wire w_dff_B_8HgM9npp3_1;
	wire w_dff_A_WQ7rGcbR6_1;
	wire w_dff_A_7KKGRqGr4_1;
	wire w_dff_A_Eo8pjj496_0;
	wire w_dff_A_iiFUvMV99_1;
	wire w_dff_A_e9pqetUX0_1;
	wire w_dff_A_BI8gDIYZ4_1;
	wire w_dff_A_c1RFncXA6_1;
	wire w_dff_A_UFFdpIeU1_1;
	wire w_dff_A_Ei9lQM4A3_1;
	wire w_dff_A_VNLWXNkb2_1;
	wire w_dff_A_EnvjuNp65_1;
	wire w_dff_A_UKT2WkAc4_1;
	wire w_dff_A_x11vc7E51_1;
	wire w_dff_A_3lQu6qF98_1;
	wire w_dff_A_v5z2xYqi5_1;
	wire w_dff_A_Pa5T8Khv1_0;
	wire w_dff_A_8LcK8OjW1_0;
	wire w_dff_A_FABQIxU61_0;
	wire w_dff_A_oU161Ncu3_2;
	wire w_dff_A_PsQowceb7_2;
	wire w_dff_A_aF5AZzhG1_2;
	wire w_dff_B_h21CaGwJ6_1;
	wire w_dff_B_l6O1nGen5_1;
	wire w_dff_B_aoQ4cO6G4_2;
	wire w_dff_A_Ez3fDP7O2_0;
	wire w_dff_A_LnfPSjCj1_2;
	wire w_dff_A_5wOY19y38_0;
	wire w_dff_A_TwEkicrX2_0;
	wire w_dff_A_HfR9wvXH0_0;
	wire w_dff_A_xFFZkzla9_1;
	wire w_dff_A_l1nYXMXi6_1;
	wire w_dff_A_S887kdNf8_1;
	wire w_dff_A_ldZ1KY7c8_1;
	wire w_dff_A_YkCQntDW9_1;
	wire w_dff_A_41bqDbRo2_1;
	wire w_dff_A_fSaZrFse3_2;
	wire w_dff_A_zlrFOdIx5_2;
	wire w_dff_A_Oh7A8BMG5_2;
	wire w_dff_A_Mbxmu5IA8_2;
	wire w_dff_A_7nHzeAQE8_0;
	wire w_dff_A_i8MxtEqX8_0;
	wire w_dff_A_gJo61eAj1_0;
	wire w_dff_A_jCSaDnGt3_0;
	wire w_dff_B_PlwNksKA7_2;
	wire w_dff_A_UiYgcqjj0_0;
	wire w_dff_A_4K5YfUEq1_0;
	wire w_dff_A_qYFnchSb5_0;
	wire w_dff_A_qg2u1FFT9_0;
	wire w_dff_A_NME46QeS8_1;
	wire w_dff_A_hrTl2yRI2_0;
	wire w_dff_A_ZBdNzVag3_0;
	wire w_dff_A_6QumpSRY2_0;
	wire w_dff_A_zAZyEvqU4_1;
	wire w_dff_A_S2y8jGwy7_1;
	wire w_dff_A_eBkTexpT7_1;
	wire w_dff_A_1GyyuEdD3_1;
	wire w_dff_A_7Jc62E2n3_1;
	wire w_dff_A_Pgbhg1V60_1;
	wire w_dff_A_yGPNZGOU3_1;
	wire w_dff_A_DQ9xXhsI5_2;
	wire w_dff_B_JFMYzIFG6_3;
	wire w_dff_B_44dd0rRk9_1;
	wire w_dff_B_hcyQBnBz9_0;
	wire w_dff_A_JffuGsQJ7_2;
	wire w_dff_A_cXHyq6OK4_1;
	wire w_dff_A_984qphLh4_2;
	wire w_dff_A_n0yhwvps7_2;
	wire w_dff_A_yxDm7fX93_0;
	wire w_dff_A_j8emn42k0_1;
	wire w_dff_A_Mop6iPGY8_0;
	wire w_dff_A_WIVPdZkN8_0;
	wire w_dff_A_vVahhG232_0;
	wire w_dff_A_hSoXGY9p8_1;
	wire w_dff_A_rsI4cXCp7_2;
	wire w_dff_A_s7ItAJyX3_2;
	wire w_dff_A_EagitJIb6_2;
	wire w_dff_A_GOOt5XX88_2;
	wire w_dff_B_8A4vRwvi3_1;
	wire w_dff_B_Lmpe7ff84_1;
	wire w_dff_A_g8Yd2so27_0;
	wire w_dff_A_e7OVtupO2_2;
	wire w_dff_A_DIwKuMg99_0;
	wire w_dff_A_7OXfBqVa7_0;
	wire w_dff_A_nDhm2kq96_0;
	wire w_dff_A_Lj9zbcUa6_1;
	wire w_dff_A_ywehXCUa1_0;
	wire w_dff_A_hpZHBmGS3_0;
	wire w_dff_A_sfSARdCR5_0;
	wire w_dff_A_nBd1YF5H6_0;
	wire w_dff_A_M3jxpyfz4_0;
	wire w_dff_A_PFYmG4hZ5_0;
	wire w_dff_A_eiOEw5107_0;
	wire w_dff_A_YXbuUOnv8_0;
	wire w_dff_A_XCVPSGM95_0;
	wire w_dff_A_ZX6fe0lf9_0;
	wire w_dff_A_uWzz0TLL9_0;
	wire w_dff_A_EfuQuOuc9_0;
	wire w_dff_A_hgvHOupC1_0;
	wire w_dff_A_wtqYKzGc1_0;
	wire w_dff_A_7XduDj1U7_0;
	wire w_dff_A_A7GNF2XS4_0;
	wire w_dff_A_CEmI8Lxr6_0;
	wire w_dff_A_5PrQnNSk7_0;
	wire w_dff_A_2sPFJEsh9_0;
	wire w_dff_A_9b6dwdyC6_0;
	wire w_dff_A_aZWE634o2_0;
	wire w_dff_A_BEWgpPnm6_0;
	wire w_dff_A_MNU1QNoV9_0;
	wire w_dff_A_LX11k00f7_0;
	wire w_dff_A_iNnnpCsJ0_0;
	wire w_dff_A_bKUyBodi8_1;
	wire w_dff_A_v285L7xL5_0;
	wire w_dff_A_rUDYX13a7_0;
	wire w_dff_A_4tDnO5nJ5_0;
	wire w_dff_A_h0o3o1xr8_0;
	wire w_dff_A_OYeP2yOu7_0;
	wire w_dff_A_uKTFaQJ35_0;
	wire w_dff_A_eUrAMSmT5_0;
	wire w_dff_A_yHDXYlgH7_0;
	wire w_dff_A_TMxFEqwz9_0;
	wire w_dff_A_tVliGP8n1_0;
	wire w_dff_A_nt2KtYtx8_0;
	wire w_dff_A_8p4nqR3a8_0;
	wire w_dff_A_BKsLBISq9_0;
	wire w_dff_A_YZsBBmMq7_0;
	wire w_dff_A_lSdz3bWj1_0;
	wire w_dff_A_C3PejpNi8_0;
	wire w_dff_A_1tqrNl0d8_0;
	wire w_dff_A_7dJI4oOY1_0;
	wire w_dff_A_JG1vOCvW3_0;
	wire w_dff_A_MdcULH4j6_0;
	wire w_dff_A_rnzCGt0E3_0;
	wire w_dff_A_LpNmMvXA5_0;
	wire w_dff_A_8pPVXDib0_0;
	wire w_dff_A_wOKaWCPZ0_0;
	wire w_dff_A_4RoSXpPO6_0;
	wire w_dff_A_ykkR7BTX5_1;
	wire w_dff_A_EpDTHM1d0_0;
	wire w_dff_A_brZ3xIhE2_0;
	wire w_dff_A_mqLJ9KNt3_0;
	wire w_dff_A_ToyAXf8w3_0;
	wire w_dff_A_LuN51aD65_0;
	wire w_dff_A_XH5w1yxR1_0;
	wire w_dff_A_3nAWI0la7_0;
	wire w_dff_A_ZRPZAtOX5_0;
	wire w_dff_A_c7HJVQT50_0;
	wire w_dff_A_7wrTDaOS1_0;
	wire w_dff_A_VAz7b4Gi5_0;
	wire w_dff_A_6SFwqig01_0;
	wire w_dff_A_IOVpHB1G7_0;
	wire w_dff_A_RyEOauqP4_0;
	wire w_dff_A_6ZTgUnNV6_0;
	wire w_dff_A_VThvqpi84_0;
	wire w_dff_A_K5pe7vPB7_0;
	wire w_dff_A_K3AtxB7M4_0;
	wire w_dff_A_A9TpM5qa7_0;
	wire w_dff_A_jhEdUKFC0_0;
	wire w_dff_A_Coq6BMl46_0;
	wire w_dff_A_hv1lnQ6D7_0;
	wire w_dff_A_AVvk53uu6_0;
	wire w_dff_A_zRW9CPGS3_0;
	wire w_dff_A_teD8M2gk8_0;
	wire w_dff_A_5BZl4JPk1_1;
	wire w_dff_A_PIJL7jhG7_0;
	wire w_dff_A_FnQYp6ul2_0;
	wire w_dff_A_i4X35nkB3_0;
	wire w_dff_A_X1aQbOx61_0;
	wire w_dff_A_Tz9Ll54v1_0;
	wire w_dff_A_N9m2u4dY9_0;
	wire w_dff_A_xSNJ1BTN8_0;
	wire w_dff_A_4kKgQLrM4_0;
	wire w_dff_A_h1PCNJ8L1_0;
	wire w_dff_A_LWfeLkUz3_0;
	wire w_dff_A_XFMDUF8M2_0;
	wire w_dff_A_USC1GW618_0;
	wire w_dff_A_f0pTPOsW2_0;
	wire w_dff_A_6dARqQ2a3_0;
	wire w_dff_A_svgvGrkX3_0;
	wire w_dff_A_qZKJUXgl6_0;
	wire w_dff_A_aw2zk8MI0_0;
	wire w_dff_A_FnH9o1Tb4_0;
	wire w_dff_A_eOlFEr7z1_0;
	wire w_dff_A_bVOZMBm67_0;
	wire w_dff_A_14yrAvKb5_0;
	wire w_dff_A_lkSNs8He8_0;
	wire w_dff_A_vvfK3lCp9_0;
	wire w_dff_A_v2yELCdE9_0;
	wire w_dff_A_3PEnCtBv8_0;
	wire w_dff_A_lpzyHoCB3_1;
	wire w_dff_A_oDbiegJ57_0;
	wire w_dff_A_Hhzsciea1_0;
	wire w_dff_A_YwcUCT5Z8_0;
	wire w_dff_A_n817RTmT7_0;
	wire w_dff_A_nxrsyCh59_0;
	wire w_dff_A_7voHvPDZ3_0;
	wire w_dff_A_UqJ05x1V3_0;
	wire w_dff_A_5n1Pyn2d8_0;
	wire w_dff_A_u8dNkfQO1_0;
	wire w_dff_A_1yUxlyNT3_0;
	wire w_dff_A_0N75zwGr0_0;
	wire w_dff_A_1rln8GPN5_0;
	wire w_dff_A_9yOpdUW36_0;
	wire w_dff_A_FdeNCbK17_0;
	wire w_dff_A_SWqyt6at7_0;
	wire w_dff_A_JZ3Vvpni9_0;
	wire w_dff_A_i8ZCNfUd9_0;
	wire w_dff_A_0lmWSpFa0_0;
	wire w_dff_A_3j3Lnv4x0_0;
	wire w_dff_A_fqLPO4jp5_0;
	wire w_dff_A_y7pZHwE02_0;
	wire w_dff_A_sUDznM3e7_0;
	wire w_dff_A_4KUrw3ax4_0;
	wire w_dff_A_9XzUPOPa3_0;
	wire w_dff_A_LrxXiihK5_0;
	wire w_dff_A_rEh14yc44_1;
	wire w_dff_A_WHwPWy2u7_0;
	wire w_dff_A_u3PY3FCf3_0;
	wire w_dff_A_IAxjzWOd2_0;
	wire w_dff_A_tkmeiAQe7_0;
	wire w_dff_A_E7tDs0jO9_0;
	wire w_dff_A_PvvokCLV7_0;
	wire w_dff_A_UjGj5Ycc8_0;
	wire w_dff_A_1F61HQYx6_0;
	wire w_dff_A_ixNBkNpN0_0;
	wire w_dff_A_VrxocDes2_0;
	wire w_dff_A_wT6ECk2p1_0;
	wire w_dff_A_Oq07xbS00_0;
	wire w_dff_A_2CA241fZ3_0;
	wire w_dff_A_nDr6tM732_0;
	wire w_dff_A_zvMdIWmt8_0;
	wire w_dff_A_0BcZrKz53_0;
	wire w_dff_A_XcAMIdEi2_0;
	wire w_dff_A_EK9vnq0r5_0;
	wire w_dff_A_M64VN9N93_0;
	wire w_dff_A_PXIRguxK4_0;
	wire w_dff_A_1dGvCvkD2_0;
	wire w_dff_A_aGWXHUdU9_0;
	wire w_dff_A_oKOQuPsj7_0;
	wire w_dff_A_PMovNCDZ8_0;
	wire w_dff_A_RUro9E0k3_0;
	wire w_dff_A_Qb2jOS5o0_1;
	wire w_dff_A_tIWBtJn27_0;
	wire w_dff_A_OA0wYm853_0;
	wire w_dff_A_G3QHnqgV6_0;
	wire w_dff_A_gFSGMReh4_0;
	wire w_dff_A_XM9QDtR27_0;
	wire w_dff_A_F7xGfi0s8_0;
	wire w_dff_A_OWvvromt7_0;
	wire w_dff_A_PX9v89ft9_0;
	wire w_dff_A_piwCPmhX3_0;
	wire w_dff_A_NO5XX01t3_0;
	wire w_dff_A_5f7o3nb18_0;
	wire w_dff_A_2oEv4P7U4_0;
	wire w_dff_A_SlzhVd5S8_0;
	wire w_dff_A_cSzB5Gr83_0;
	wire w_dff_A_t2p3AynC4_0;
	wire w_dff_A_fE6VYTnp9_0;
	wire w_dff_A_KIr9fKK00_0;
	wire w_dff_A_rDeUE6176_0;
	wire w_dff_A_HaGEhSji1_0;
	wire w_dff_A_Inbqn0dD7_0;
	wire w_dff_A_3q9vZQW89_0;
	wire w_dff_A_IGygduFJ1_0;
	wire w_dff_A_Bv5RYsxJ9_0;
	wire w_dff_A_zDxST4zS3_0;
	wire w_dff_A_bZbRI6vH5_0;
	wire w_dff_A_lmpG2qDt1_1;
	wire w_dff_A_uNDxEd1U6_0;
	wire w_dff_A_goDTdAAp2_0;
	wire w_dff_A_XRqvAbIk7_0;
	wire w_dff_A_gsrNM9RN2_0;
	wire w_dff_A_guYgLIJS6_0;
	wire w_dff_A_9AMwW71b3_0;
	wire w_dff_A_ykmvIyn41_0;
	wire w_dff_A_xoOlKdZ24_0;
	wire w_dff_A_GburK90B9_0;
	wire w_dff_A_OeN8qLYi2_0;
	wire w_dff_A_EvhxFCeK1_0;
	wire w_dff_A_O203UWHR0_0;
	wire w_dff_A_FeU06reW0_0;
	wire w_dff_A_ZBYZw6Ck2_0;
	wire w_dff_A_KQ5R8WS64_0;
	wire w_dff_A_paOEspV96_0;
	wire w_dff_A_sjJDN5VP2_0;
	wire w_dff_A_QS5hikjm0_0;
	wire w_dff_A_pS4Sz9By5_0;
	wire w_dff_A_U3z2FtCz3_0;
	wire w_dff_A_FrdDRHar5_0;
	wire w_dff_A_r8DucLA32_0;
	wire w_dff_A_pX4mqxh24_0;
	wire w_dff_A_0BrYTy6u5_0;
	wire w_dff_A_6BcXm8jQ7_0;
	wire w_dff_A_6XQh2fku4_1;
	wire w_dff_A_refaBZnK1_0;
	wire w_dff_A_v7pSivbv4_0;
	wire w_dff_A_5WO8c8WX3_0;
	wire w_dff_A_9ctrAMm45_0;
	wire w_dff_A_XG5Z3lUp0_0;
	wire w_dff_A_mIdx8PiL0_0;
	wire w_dff_A_s97xlK6J4_0;
	wire w_dff_A_MgW2xVXs6_0;
	wire w_dff_A_hYAfsJQT8_0;
	wire w_dff_A_4HD76SjN7_0;
	wire w_dff_A_lmRroHVc8_0;
	wire w_dff_A_Y5QSLk240_0;
	wire w_dff_A_850XsCfT5_0;
	wire w_dff_A_JBpYG9X07_0;
	wire w_dff_A_WjllqeKO9_0;
	wire w_dff_A_i7k7jgCg0_0;
	wire w_dff_A_yloCJqOE0_0;
	wire w_dff_A_0OnIPhgy8_0;
	wire w_dff_A_z8RBLO0Y4_0;
	wire w_dff_A_4ecQ7nfB0_0;
	wire w_dff_A_3C99x4QS6_0;
	wire w_dff_A_FP1CR0gh5_0;
	wire w_dff_A_xSRs55z35_0;
	wire w_dff_A_skyWf8pi4_0;
	wire w_dff_A_9kzeriYN3_0;
	wire w_dff_A_hlgqtfXa0_1;
	wire w_dff_A_tbOYvf3p0_0;
	wire w_dff_A_hLJMW56M1_0;
	wire w_dff_A_dejgQg8S3_0;
	wire w_dff_A_ps2e0bHv0_0;
	wire w_dff_A_eStmDrLs9_0;
	wire w_dff_A_m7KfGna07_0;
	wire w_dff_A_3SlH0Ty24_0;
	wire w_dff_A_oG9KUfTy3_0;
	wire w_dff_A_wjNvo2rN9_0;
	wire w_dff_A_2TqheRFW2_0;
	wire w_dff_A_NoRlpiHW3_0;
	wire w_dff_A_YGEGc6Wu1_0;
	wire w_dff_A_4iv8EiES8_0;
	wire w_dff_A_74ndzxJd2_0;
	wire w_dff_A_6UgmVWUd7_0;
	wire w_dff_A_BrI94TK16_0;
	wire w_dff_A_UKYlCVZ00_0;
	wire w_dff_A_0CxWStX33_0;
	wire w_dff_A_1cE0Kbcx5_0;
	wire w_dff_A_Bc9wqrlK4_0;
	wire w_dff_A_pgItJNNg9_0;
	wire w_dff_A_CTE9SC373_0;
	wire w_dff_A_0b5GBUFN6_0;
	wire w_dff_A_iTnffcDf9_0;
	wire w_dff_A_plhMp4FJ4_0;
	wire w_dff_A_k7VluDx66_1;
	wire w_dff_A_4JCyLnPT8_0;
	wire w_dff_A_CqQVVofU5_0;
	wire w_dff_A_0tGO98om5_0;
	wire w_dff_A_cus2wNyR3_0;
	wire w_dff_A_ykwg2N3S4_0;
	wire w_dff_A_rHEvjDg05_0;
	wire w_dff_A_Nr2H2tn92_0;
	wire w_dff_A_OWbhJzUE5_0;
	wire w_dff_A_SyABLrul8_0;
	wire w_dff_A_oAEcGWz79_0;
	wire w_dff_A_1JtRs0mg6_0;
	wire w_dff_A_QvhOosfP7_0;
	wire w_dff_A_cldCjiAI9_0;
	wire w_dff_A_2dCumnk10_0;
	wire w_dff_A_drQEzZcd0_0;
	wire w_dff_A_6m0xKfwG8_0;
	wire w_dff_A_EMeWYtEd7_0;
	wire w_dff_A_mq1eryS33_0;
	wire w_dff_A_vw7Fow2q3_0;
	wire w_dff_A_7X219nVw4_0;
	wire w_dff_A_zTqGXTec1_0;
	wire w_dff_A_SVAf83Wu1_0;
	wire w_dff_A_GYtMXHAg0_0;
	wire w_dff_A_Lg75cSrF3_0;
	wire w_dff_A_7Aqi7KFB9_0;
	wire w_dff_A_f0loBwmj7_1;
	wire w_dff_A_UA06XAEd3_0;
	wire w_dff_A_KQkcnd6s5_0;
	wire w_dff_A_Xebfgn7k8_0;
	wire w_dff_A_Kb6DbJdl0_0;
	wire w_dff_A_oiQwF4St6_0;
	wire w_dff_A_7LVfNoyI8_0;
	wire w_dff_A_fbw2mTka4_0;
	wire w_dff_A_sguDky4c4_0;
	wire w_dff_A_6G8WXdwX6_0;
	wire w_dff_A_uVPYL2Fk3_0;
	wire w_dff_A_4VR2xzza4_0;
	wire w_dff_A_3c7hkXfT7_0;
	wire w_dff_A_PLL3p1Ae0_0;
	wire w_dff_A_UDPIlZY19_0;
	wire w_dff_A_gPGJ0XNR6_0;
	wire w_dff_A_VApq8idV0_0;
	wire w_dff_A_PCnDiEUn8_0;
	wire w_dff_A_QcPzhlbh9_0;
	wire w_dff_A_PErFiEsZ7_0;
	wire w_dff_A_LPQLaZXx8_0;
	wire w_dff_A_nU3rmj2L1_0;
	wire w_dff_A_K9Z7zOhI0_0;
	wire w_dff_A_5J3jbhlA4_0;
	wire w_dff_A_qfbcGDFo5_0;
	wire w_dff_A_W040WQg59_0;
	wire w_dff_A_KZTb2yWC7_1;
	wire w_dff_A_9m7fLkwH1_0;
	wire w_dff_A_9o66xI0j9_0;
	wire w_dff_A_74RbtHo87_0;
	wire w_dff_A_SJrsLISZ6_0;
	wire w_dff_A_YDCImGTg2_0;
	wire w_dff_A_pKIbaLtX3_0;
	wire w_dff_A_8u03lCP34_0;
	wire w_dff_A_XAn5zpBf1_0;
	wire w_dff_A_ji7vzwIU7_0;
	wire w_dff_A_0CFrNTyK3_0;
	wire w_dff_A_SpUmqvJX4_0;
	wire w_dff_A_JFCxMApy4_0;
	wire w_dff_A_2o52tIzB6_0;
	wire w_dff_A_X0IpWm9L2_0;
	wire w_dff_A_67dkHOgN2_0;
	wire w_dff_A_gC4IHWYU7_0;
	wire w_dff_A_NuZIAZZe1_0;
	wire w_dff_A_YurapNLy8_0;
	wire w_dff_A_BLCgKjbE5_0;
	wire w_dff_A_nHtR25q09_0;
	wire w_dff_A_5m64xqTj3_0;
	wire w_dff_A_C39eLG786_0;
	wire w_dff_A_Z5fCVx9H0_0;
	wire w_dff_A_Ypbcdhpv7_0;
	wire w_dff_A_Qm1nj8Uz2_0;
	wire w_dff_A_QLfkh51b8_1;
	wire w_dff_A_DUa9HZnC3_0;
	wire w_dff_A_UlCDh2JK1_0;
	wire w_dff_A_N2V6AKne6_0;
	wire w_dff_A_cG8znGBF0_0;
	wire w_dff_A_jU9dvUXv4_0;
	wire w_dff_A_6cpxOmBw2_0;
	wire w_dff_A_mc0wcpd06_0;
	wire w_dff_A_LHj9tWjm9_0;
	wire w_dff_A_1hts7Ibg8_0;
	wire w_dff_A_oB5odyPv2_0;
	wire w_dff_A_MKcANnJ04_0;
	wire w_dff_A_9CFgohJx4_0;
	wire w_dff_A_QwEVE3bG8_0;
	wire w_dff_A_vd3cvdKb9_0;
	wire w_dff_A_f0Zkd5IP9_0;
	wire w_dff_A_W3zNEd0U5_0;
	wire w_dff_A_z1aJ5j6L9_0;
	wire w_dff_A_FjTypjNG6_0;
	wire w_dff_A_G7vqqoYa4_0;
	wire w_dff_A_xw6jvl1U5_0;
	wire w_dff_A_SDEeN8se9_0;
	wire w_dff_A_bIifVykH6_0;
	wire w_dff_A_CtIWqBnI8_0;
	wire w_dff_A_5PdX3Cv19_0;
	wire w_dff_A_RIUIkOOA8_0;
	wire w_dff_A_OfURwhBQ4_1;
	wire w_dff_A_ytSQMmZV7_0;
	wire w_dff_A_yINPCqiF1_0;
	wire w_dff_A_aX0zZrfI5_0;
	wire w_dff_A_Z4owilih7_0;
	wire w_dff_A_tA2mEIM04_0;
	wire w_dff_A_RNvZio891_0;
	wire w_dff_A_7PgBZI536_0;
	wire w_dff_A_ZMV5J3RQ6_0;
	wire w_dff_A_zDAudBa62_0;
	wire w_dff_A_drX3DFpO8_0;
	wire w_dff_A_iwCJhtCM6_0;
	wire w_dff_A_VnZKnpWY9_0;
	wire w_dff_A_uRyf39Wa0_0;
	wire w_dff_A_XCCaCKBf8_0;
	wire w_dff_A_0RZ9zW1X4_0;
	wire w_dff_A_WfZcjshR7_0;
	wire w_dff_A_B88VNbXs3_0;
	wire w_dff_A_YkKK2TBb4_0;
	wire w_dff_A_3JpGJlkj6_0;
	wire w_dff_A_aRnGBIFF9_0;
	wire w_dff_A_9LIutuJ13_0;
	wire w_dff_A_AagqdROk1_0;
	wire w_dff_A_QmDodXM35_0;
	wire w_dff_A_9HjBWwfe6_0;
	wire w_dff_A_980EDFiP5_0;
	wire w_dff_A_fIekaECE3_1;
	wire w_dff_A_bk775PTy5_0;
	wire w_dff_A_IIfDcN731_0;
	wire w_dff_A_5PMu0ONu2_0;
	wire w_dff_A_eLol9rpd9_0;
	wire w_dff_A_PLHaiAic9_0;
	wire w_dff_A_mZTV7jyz6_0;
	wire w_dff_A_lcJl65Ah2_0;
	wire w_dff_A_6QXCIqm39_0;
	wire w_dff_A_dSNySXUc9_0;
	wire w_dff_A_7l5v8nxi4_0;
	wire w_dff_A_rNrrtCYT4_0;
	wire w_dff_A_CHI7qLaG5_0;
	wire w_dff_A_sELod8Nb5_0;
	wire w_dff_A_xf27V03z0_0;
	wire w_dff_A_7tmE429A8_0;
	wire w_dff_A_MESAuxb88_0;
	wire w_dff_A_vwHscXbt7_0;
	wire w_dff_A_PLGKFfh65_0;
	wire w_dff_A_d75bt1mm2_0;
	wire w_dff_A_etmB4GOC4_0;
	wire w_dff_A_sBArkJi94_0;
	wire w_dff_A_Z8MyH8wl9_0;
	wire w_dff_A_Z2kC9TQE6_0;
	wire w_dff_A_nLGhbYri1_0;
	wire w_dff_A_CCE3pTEC0_0;
	wire w_dff_A_gOv57F6o7_1;
	wire w_dff_A_4ycNk5ue3_0;
	wire w_dff_A_kQb6alwb4_0;
	wire w_dff_A_750YHGfC0_0;
	wire w_dff_A_1jsP5YW74_0;
	wire w_dff_A_rQRGYg105_0;
	wire w_dff_A_pGGC2MO08_0;
	wire w_dff_A_hz0j8EbO0_0;
	wire w_dff_A_wvPlMp6f5_0;
	wire w_dff_A_te0lC6vD2_0;
	wire w_dff_A_lTnOwFar8_0;
	wire w_dff_A_axSqLTYo9_0;
	wire w_dff_A_vVKtUhnG0_0;
	wire w_dff_A_gKwZEhym9_0;
	wire w_dff_A_SQYHVqPZ2_0;
	wire w_dff_A_GszOT3Ft5_0;
	wire w_dff_A_1KIl7Y784_0;
	wire w_dff_A_HGmNnvMP1_0;
	wire w_dff_A_fjvhIx1R6_0;
	wire w_dff_A_VKCNYq9P8_0;
	wire w_dff_A_lM8MGmMt3_0;
	wire w_dff_A_N8yYnooQ6_0;
	wire w_dff_A_NSmpGyrU1_0;
	wire w_dff_A_PWWzkdMT3_0;
	wire w_dff_A_AcKnVu8F1_0;
	wire w_dff_A_1IMPCMjz6_0;
	wire w_dff_A_11QQyRH85_1;
	wire w_dff_A_UjXJohJy7_0;
	wire w_dff_A_ShEUuRJO0_0;
	wire w_dff_A_tg3mlVew4_0;
	wire w_dff_A_4J1i6TzQ3_0;
	wire w_dff_A_7ZwDlCyW6_0;
	wire w_dff_A_VXPcrupP7_0;
	wire w_dff_A_Itga5flg1_0;
	wire w_dff_A_VwnCLoSN9_0;
	wire w_dff_A_91dpDgg91_0;
	wire w_dff_A_UpWY8KVq9_0;
	wire w_dff_A_bAoMvQUp4_0;
	wire w_dff_A_UgK6i5xj8_0;
	wire w_dff_A_3H0IbKDz8_0;
	wire w_dff_A_wbSVtmAL5_0;
	wire w_dff_A_83nN3jnE0_0;
	wire w_dff_A_52jTadLY9_0;
	wire w_dff_A_Bt01Oqwz6_0;
	wire w_dff_A_BAh45ch20_0;
	wire w_dff_A_lVSsa0Tp3_0;
	wire w_dff_A_WlWbRkXP1_0;
	wire w_dff_A_P2OROSa06_0;
	wire w_dff_A_SxaMNOeq4_0;
	wire w_dff_A_yA0kOM8s5_0;
	wire w_dff_A_2QpzgJ2M6_0;
	wire w_dff_A_Cnhvxw4A4_0;
	wire w_dff_A_9okMP1UV2_1;
	wire w_dff_A_W0z5pZCe5_0;
	wire w_dff_A_tqrobSO45_0;
	wire w_dff_A_olNmtkdm8_0;
	wire w_dff_A_vckhYKQb4_0;
	wire w_dff_A_kBPXqeMc7_0;
	wire w_dff_A_g3WJ2c3N6_0;
	wire w_dff_A_wM3Xz4T23_0;
	wire w_dff_A_CCiZ0XNY6_0;
	wire w_dff_A_xLCoukH15_0;
	wire w_dff_A_XGY4ms5n3_0;
	wire w_dff_A_G41BNQGi2_0;
	wire w_dff_A_FL7zkHKh0_0;
	wire w_dff_A_3HXQdHjF9_0;
	wire w_dff_A_5gDjCqpK0_0;
	wire w_dff_A_nOXzo6UW1_0;
	wire w_dff_A_9zHsPENT5_0;
	wire w_dff_A_SSqTzJ4a8_0;
	wire w_dff_A_WC0oSFax0_0;
	wire w_dff_A_Nw7VJFwA3_0;
	wire w_dff_A_a2kMC4mj5_0;
	wire w_dff_A_FMGgHupn6_0;
	wire w_dff_A_F6impo4g7_0;
	wire w_dff_A_T8b8AyAx1_0;
	wire w_dff_A_B7P0jwiJ3_0;
	wire w_dff_A_QByHr7ms8_0;
	wire w_dff_A_XMLPmksm8_1;
	wire w_dff_A_nXCBi7Zg4_0;
	wire w_dff_A_vata1kJy9_0;
	wire w_dff_A_X5xU5kKc2_0;
	wire w_dff_A_OcHyEATI4_0;
	wire w_dff_A_xtrwPTaF7_0;
	wire w_dff_A_TuikUtQJ5_0;
	wire w_dff_A_ScJYNUfR6_0;
	wire w_dff_A_EFkx2fPr0_0;
	wire w_dff_A_05fRovvS0_0;
	wire w_dff_A_gOoMGAOP1_0;
	wire w_dff_A_6CdV0Dx76_0;
	wire w_dff_A_vhsbPAM43_0;
	wire w_dff_A_U2PW0Nf06_0;
	wire w_dff_A_x6PQxXnG6_0;
	wire w_dff_A_g1Ki7iYn5_0;
	wire w_dff_A_LSN81seR6_0;
	wire w_dff_A_umLDc4e32_0;
	wire w_dff_A_D3Z8w65C0_0;
	wire w_dff_A_kZ0VP6MF3_0;
	wire w_dff_A_9MQfuMzn7_0;
	wire w_dff_A_Q4hBb8IV3_0;
	wire w_dff_A_zSXUF6JB8_0;
	wire w_dff_A_FxPuHxzq9_0;
	wire w_dff_A_fIEu4iUG2_0;
	wire w_dff_A_aSYzNRAE5_0;
	wire w_dff_A_RwGKFHG76_1;
	wire w_dff_A_pSsJqAGi2_0;
	wire w_dff_A_QTQ3LRou3_0;
	wire w_dff_A_zHpTy2Ma4_0;
	wire w_dff_A_6U9Q47tX8_0;
	wire w_dff_A_vQSlVRYl5_0;
	wire w_dff_A_lqbPE6rA9_0;
	wire w_dff_A_DhQ8CBJN5_0;
	wire w_dff_A_0mmd6iAP6_0;
	wire w_dff_A_B4B3iqNi7_0;
	wire w_dff_A_6V3SgN718_0;
	wire w_dff_A_xPzwMw5Y4_0;
	wire w_dff_A_pFhm7M850_0;
	wire w_dff_A_DHgizohK1_0;
	wire w_dff_A_QoKQdfTy8_0;
	wire w_dff_A_xdsvHBIa9_0;
	wire w_dff_A_FqKVM69n1_0;
	wire w_dff_A_z73PWgP01_0;
	wire w_dff_A_KZNvMPRo8_0;
	wire w_dff_A_DDY7NAzT2_0;
	wire w_dff_A_WmMGUKcV8_0;
	wire w_dff_A_Eu8t7ZoD2_0;
	wire w_dff_A_Ui7AEILB9_0;
	wire w_dff_A_MXzLsN6d8_0;
	wire w_dff_A_uaTHpDKo8_0;
	wire w_dff_A_yI6apG2r3_0;
	wire w_dff_A_o7j95bj09_1;
	wire w_dff_A_RCk2tpz64_0;
	wire w_dff_A_9iGhDWcK7_0;
	wire w_dff_A_dsHEauon1_0;
	wire w_dff_A_8AZu8qJD2_0;
	wire w_dff_A_7uOv7Jir4_0;
	wire w_dff_A_0Cliso2d7_0;
	wire w_dff_A_1qFCwSei7_0;
	wire w_dff_A_G4vSpu0G5_0;
	wire w_dff_A_wE2z1JIn6_0;
	wire w_dff_A_bcaSGDxa1_0;
	wire w_dff_A_JKQi14PJ0_0;
	wire w_dff_A_C0DiUZfg5_0;
	wire w_dff_A_XkoFf4qk1_0;
	wire w_dff_A_Sb6cXqc88_0;
	wire w_dff_A_HXKwbOBe7_0;
	wire w_dff_A_SsSbmzrP0_0;
	wire w_dff_A_fT3hszoY9_0;
	wire w_dff_A_4jYnIGsu8_0;
	wire w_dff_A_mSQhwvnh6_0;
	wire w_dff_A_R2BG7Hr51_0;
	wire w_dff_A_qiy3e5fv6_0;
	wire w_dff_A_v4Qi1qBk1_0;
	wire w_dff_A_DZwuPhxq7_0;
	wire w_dff_A_gcSvZpbq3_0;
	wire w_dff_A_h2PKgTfh5_0;
	wire w_dff_A_SwcSZ5mu2_1;
	wire w_dff_A_I5TtFsPO3_0;
	wire w_dff_A_I7sBW1ym7_0;
	wire w_dff_A_8nuYlqo78_0;
	wire w_dff_A_H1pT0KGG1_0;
	wire w_dff_A_mTgeVoxi5_0;
	wire w_dff_A_r4j6ACKh3_0;
	wire w_dff_A_OpoqpKPM1_0;
	wire w_dff_A_JlLzhrCR7_0;
	wire w_dff_A_1NKXrdeO7_0;
	wire w_dff_A_FY8pf0bB7_0;
	wire w_dff_A_qNhI5oZQ8_0;
	wire w_dff_A_ex65tSP45_0;
	wire w_dff_A_LzjMLhai6_0;
	wire w_dff_A_0s70ksDY3_0;
	wire w_dff_A_eahvI2Tw5_0;
	wire w_dff_A_O5ChEaQ90_0;
	wire w_dff_A_xUzzNqTC1_0;
	wire w_dff_A_JTDcJUGE2_0;
	wire w_dff_A_OrQMIMW96_0;
	wire w_dff_A_Z0MWjToV7_0;
	wire w_dff_A_asxkmu0C6_0;
	wire w_dff_A_CnTbIlim7_0;
	wire w_dff_A_5eOxR1ck5_0;
	wire w_dff_A_YRco1Ivp7_0;
	wire w_dff_A_WqGolFye2_0;
	wire w_dff_A_UOFpF7hR0_1;
	wire w_dff_A_DFmfw6vG3_0;
	wire w_dff_A_ne2TrUOm7_0;
	wire w_dff_A_HixFBzjI3_0;
	wire w_dff_A_NtJ9bVEG1_0;
	wire w_dff_A_QP80W6xl8_0;
	wire w_dff_A_sufIrqeR3_0;
	wire w_dff_A_QHxrtEBw3_0;
	wire w_dff_A_RmGhJCkc5_0;
	wire w_dff_A_gjMK7HsI2_0;
	wire w_dff_A_63XSR0MP2_0;
	wire w_dff_A_ldZWNcFg1_0;
	wire w_dff_A_sgeEwrXI0_0;
	wire w_dff_A_T1s58ywb7_0;
	wire w_dff_A_cS2UAUHB4_0;
	wire w_dff_A_hHRRzcPO5_0;
	wire w_dff_A_GMB2abC96_0;
	wire w_dff_A_SUMRqDyo5_0;
	wire w_dff_A_bdWj76Op9_0;
	wire w_dff_A_DqUTDiHQ6_0;
	wire w_dff_A_2reMXbBq1_0;
	wire w_dff_A_h7KHJgaO4_0;
	wire w_dff_A_dwLIIFPH4_0;
	wire w_dff_A_1Wbd86ql5_0;
	wire w_dff_A_E6XSqH0Y5_0;
	wire w_dff_A_XzveyaxA5_0;
	wire w_dff_A_3rAom8zd6_1;
	wire w_dff_A_fYXRzNNc1_0;
	wire w_dff_A_Mtc00sxC0_0;
	wire w_dff_A_t5bc0efI2_0;
	wire w_dff_A_C3oAI2Fi4_0;
	wire w_dff_A_FH2lil4W1_0;
	wire w_dff_A_QqZeptEe5_0;
	wire w_dff_A_BvkR98yw1_0;
	wire w_dff_A_wBytA4eS0_0;
	wire w_dff_A_W1Nj9btQ3_0;
	wire w_dff_A_WIoNprCO3_0;
	wire w_dff_A_oTH6z8ii4_0;
	wire w_dff_A_iNIdyMhq9_0;
	wire w_dff_A_wr3GPQIf2_0;
	wire w_dff_A_RN5oxCKr4_0;
	wire w_dff_A_GBLQJdzc8_0;
	wire w_dff_A_6GrH231a8_0;
	wire w_dff_A_LzCj4MQa3_0;
	wire w_dff_A_YNuIQ53q7_0;
	wire w_dff_A_Qv19K5je0_0;
	wire w_dff_A_uVgXRt9m1_0;
	wire w_dff_A_0fqMLhtF9_0;
	wire w_dff_A_IxknPB2B0_0;
	wire w_dff_A_lDRYKVjv0_0;
	wire w_dff_A_rfayoZ0G4_0;
	wire w_dff_A_HGvALjB69_0;
	wire w_dff_A_jC7At71Q2_1;
	wire w_dff_A_LxBBIU8o3_0;
	wire w_dff_A_r9UDQrDN1_0;
	wire w_dff_A_FkUvftfL8_0;
	wire w_dff_A_tDVD6uAd0_0;
	wire w_dff_A_ujznNtWB1_0;
	wire w_dff_A_9u2bSJuP0_0;
	wire w_dff_A_6A8laloR9_0;
	wire w_dff_A_4bnnsnk34_0;
	wire w_dff_A_hCILH0XJ5_0;
	wire w_dff_A_8E1PgMP80_0;
	wire w_dff_A_cOc4c2bI7_0;
	wire w_dff_A_it3y7hed1_0;
	wire w_dff_A_GhWC7yu38_0;
	wire w_dff_A_H5skBDB29_0;
	wire w_dff_A_6obFelOy3_0;
	wire w_dff_A_cJ7KDIQ20_0;
	wire w_dff_A_9qrHKiPs2_0;
	wire w_dff_A_yclbE7nM1_0;
	wire w_dff_A_WHkxj6nR7_0;
	wire w_dff_A_ADqu8nAL5_0;
	wire w_dff_A_wvVlABbh6_0;
	wire w_dff_A_V6m99F9k9_0;
	wire w_dff_A_iGzYGW3S4_0;
	wire w_dff_A_L4fSNyRt2_0;
	wire w_dff_A_Cu3qY5nH9_0;
	wire w_dff_A_O7RMNuf06_1;
	wire w_dff_A_doiTLMWg7_0;
	wire w_dff_A_pg5VpNzU3_0;
	wire w_dff_A_uWjlNu2E3_0;
	wire w_dff_A_ljXNqORV6_0;
	wire w_dff_A_WqFnMp7F1_0;
	wire w_dff_A_yIgB1hws4_0;
	wire w_dff_A_3Mn7T0Mc1_0;
	wire w_dff_A_vKDjREg19_0;
	wire w_dff_A_y6BvsBzb5_0;
	wire w_dff_A_JefxyndS9_0;
	wire w_dff_A_OWHgQ3gL0_0;
	wire w_dff_A_w8U8XJOq5_0;
	wire w_dff_A_QbVkguio0_0;
	wire w_dff_A_NT8Dk4SR2_0;
	wire w_dff_A_aRnnqE9j7_0;
	wire w_dff_A_jkl0cphT9_0;
	wire w_dff_A_MIVY0kBj5_0;
	wire w_dff_A_I2AoVKde4_0;
	wire w_dff_A_4pytqjya8_0;
	wire w_dff_A_EP2uysYu8_0;
	wire w_dff_A_OylISZWJ4_0;
	wire w_dff_A_U3RlEzgC0_0;
	wire w_dff_A_SkPYBmGP8_0;
	wire w_dff_A_fDWQvJ6h5_0;
	wire w_dff_A_6MiqYO5M0_0;
	wire w_dff_A_cykvuITa8_1;
	wire w_dff_A_770ukYv22_0;
	wire w_dff_A_aJRWQdhK0_0;
	wire w_dff_A_lKFzJtcr0_0;
	wire w_dff_A_q9bJKAqu5_0;
	wire w_dff_A_zVZkXWJq6_0;
	wire w_dff_A_xo0s4Jdx9_0;
	wire w_dff_A_qYZ9UaqO6_0;
	wire w_dff_A_zeNUlbEx4_0;
	wire w_dff_A_WqjG7eI77_0;
	wire w_dff_A_1Zn3Ue1k8_0;
	wire w_dff_A_u1bfDX7C2_0;
	wire w_dff_A_E1CkVYeH5_0;
	wire w_dff_A_TymXuwcy5_0;
	wire w_dff_A_wG4UJRUV2_0;
	wire w_dff_A_DMadvdJh4_0;
	wire w_dff_A_bM89scTp8_0;
	wire w_dff_A_jUY7NL5b5_0;
	wire w_dff_A_aMmGBlsD6_0;
	wire w_dff_A_s7grm0hQ4_0;
	wire w_dff_A_56FFMSOa8_0;
	wire w_dff_A_VhFAjZOL5_0;
	wire w_dff_A_rSbD6nUO1_0;
	wire w_dff_A_4S3Q3aPN4_0;
	wire w_dff_A_f2bmOJli8_0;
	wire w_dff_A_Ub6SdZnE2_0;
	wire w_dff_A_ZmdyHmdd8_1;
	wire w_dff_A_mcWpOpJu8_0;
	wire w_dff_A_JAMipuF20_0;
	wire w_dff_A_lcdRUCoI8_0;
	wire w_dff_A_l0sFi7ci9_0;
	wire w_dff_A_14pZ2zFV1_0;
	wire w_dff_A_kM4IefWL3_0;
	wire w_dff_A_3SC9EuCc1_0;
	wire w_dff_A_p9rERASQ0_0;
	wire w_dff_A_w18NPP820_0;
	wire w_dff_A_xQNOfzUB7_0;
	wire w_dff_A_z1NqDnVO2_0;
	wire w_dff_A_Pznzn9Fh9_0;
	wire w_dff_A_RnIBIxir5_0;
	wire w_dff_A_bilz34lm8_0;
	wire w_dff_A_AefvOYKG9_0;
	wire w_dff_A_DhX6PBLq1_0;
	wire w_dff_A_7kpp6Y2X0_0;
	wire w_dff_A_il0yoA8c2_0;
	wire w_dff_A_VNUV6xRn4_0;
	wire w_dff_A_UsKiHWMT2_0;
	wire w_dff_A_RhI2wq0z5_0;
	wire w_dff_A_NTf5VPGD7_0;
	wire w_dff_A_bTcdFqlR5_0;
	wire w_dff_A_1E3cOk3U5_0;
	wire w_dff_A_6latRHez4_0;
	wire w_dff_A_bVT2Wp258_1;
	wire w_dff_A_TWjxMiy76_0;
	wire w_dff_A_ZEcQB5Jl7_0;
	wire w_dff_A_DNfbcwZX4_0;
	wire w_dff_A_rt1KetpS8_0;
	wire w_dff_A_d83EbDdg2_0;
	wire w_dff_A_3bZAt0Hm5_0;
	wire w_dff_A_gBrCuvdu4_0;
	wire w_dff_A_W5yMHXz95_0;
	wire w_dff_A_ZZ9zmRnp3_0;
	wire w_dff_A_31WN9WR89_0;
	wire w_dff_A_dGioZHas1_0;
	wire w_dff_A_NP4F7CHk5_0;
	wire w_dff_A_txfAdmnr5_0;
	wire w_dff_A_dE6GOoFS8_0;
	wire w_dff_A_bL9jkJr21_0;
	wire w_dff_A_PCsnKyw47_0;
	wire w_dff_A_WKZ7MFIb3_0;
	wire w_dff_A_dehq0JxD4_0;
	wire w_dff_A_PRdaNg3o0_0;
	wire w_dff_A_73lR5fPK3_0;
	wire w_dff_A_BwZ9htRo1_0;
	wire w_dff_A_VUwT3GaX3_0;
	wire w_dff_A_apxQIS8p5_0;
	wire w_dff_A_CK0UtfAN4_0;
	wire w_dff_A_9vdyOd9n5_0;
	wire w_dff_A_1ISwIh973_1;
	wire w_dff_A_xxcJnGPc1_0;
	wire w_dff_A_1f89aRfw3_0;
	wire w_dff_A_zaiDhMWa6_0;
	wire w_dff_A_xlZk6Hun3_0;
	wire w_dff_A_IiRPdPLX1_0;
	wire w_dff_A_AmsLyTTL7_0;
	wire w_dff_A_UYH5WbYg5_0;
	wire w_dff_A_xzCKYHee1_0;
	wire w_dff_A_F0ydn2vw7_0;
	wire w_dff_A_lf1zOueQ8_0;
	wire w_dff_A_mrDtIXis0_0;
	wire w_dff_A_CiyHWuyA4_0;
	wire w_dff_A_5yH4yel01_0;
	wire w_dff_A_zLGMLEYs7_0;
	wire w_dff_A_V1JJ2rO97_0;
	wire w_dff_A_4oZSJe060_0;
	wire w_dff_A_t118G6i42_0;
	wire w_dff_A_Ot5bP7Dg0_0;
	wire w_dff_A_Ty92eDGb9_0;
	wire w_dff_A_qKlU8vAu5_0;
	wire w_dff_A_qzBzlYFR7_0;
	wire w_dff_A_qOnaJgEF2_0;
	wire w_dff_A_rP1B7lWF8_0;
	wire w_dff_A_qbRmjG5t1_0;
	wire w_dff_A_CAN7PF2s2_0;
	wire w_dff_A_uyVV29G02_1;
	wire w_dff_A_YpAS42Pd0_0;
	wire w_dff_A_aABiHqDV8_0;
	wire w_dff_A_wUqlU6bb6_0;
	wire w_dff_A_HpeNI6hu8_0;
	wire w_dff_A_31ifhgLe3_0;
	wire w_dff_A_20LL0kXl3_0;
	wire w_dff_A_5frTfrNj9_0;
	wire w_dff_A_MnRCGrLU2_0;
	wire w_dff_A_iyKzf2e81_0;
	wire w_dff_A_bHVODOSr4_0;
	wire w_dff_A_BgMe5zfd0_0;
	wire w_dff_A_IYQi4gKK1_0;
	wire w_dff_A_vyipA3Is1_0;
	wire w_dff_A_QQxLPPac5_0;
	wire w_dff_A_bYELoScb0_0;
	wire w_dff_A_zy7vFfa32_0;
	wire w_dff_A_JDIrwvVA2_0;
	wire w_dff_A_627Yje469_0;
	wire w_dff_A_TMA9OBaf5_0;
	wire w_dff_A_O8OwSJCu5_0;
	wire w_dff_A_wsyX4SW31_0;
	wire w_dff_A_Y70sezAz6_0;
	wire w_dff_A_dc3tr08t9_0;
	wire w_dff_A_C1dJ18Gh8_0;
	wire w_dff_A_XzuygA3z9_0;
	wire w_dff_A_paBQc1dR5_1;
	wire w_dff_A_KrKWbOFh4_0;
	wire w_dff_A_owVCqCIt3_0;
	wire w_dff_A_8tjNKYJW7_0;
	wire w_dff_A_IKRWkruj3_0;
	wire w_dff_A_7ILXqpvi9_0;
	wire w_dff_A_9ssq8esx2_0;
	wire w_dff_A_mz5ZwWi41_0;
	wire w_dff_A_S3H3brTp1_0;
	wire w_dff_A_R3hJPeZ30_0;
	wire w_dff_A_M19Bz4np1_0;
	wire w_dff_A_1xd8j4TM9_0;
	wire w_dff_A_bjysYcGH5_0;
	wire w_dff_A_yFlYAY4Q1_0;
	wire w_dff_A_Itab8r2P7_0;
	wire w_dff_A_nxHJwfuq2_0;
	wire w_dff_A_qjpSuRHT0_0;
	wire w_dff_A_M21h6pYF5_0;
	wire w_dff_A_meqkVuQd2_0;
	wire w_dff_A_1SqBkC2z1_0;
	wire w_dff_A_mfmqXWB09_0;
	wire w_dff_A_wkbJbniV5_0;
	wire w_dff_A_bDCKCygv0_0;
	wire w_dff_A_tRoI4P0z5_0;
	wire w_dff_A_Ulamf9mu4_0;
	wire w_dff_A_DLzrrKos7_0;
	wire w_dff_A_BhtDhst74_1;
	wire w_dff_A_PAVZXrKf0_0;
	wire w_dff_A_01cYpg8b6_0;
	wire w_dff_A_fajuVp6Z6_0;
	wire w_dff_A_DJXiWyPe2_0;
	wire w_dff_A_dlsyUagO4_0;
	wire w_dff_A_vmKx730D5_0;
	wire w_dff_A_0RmeoFv85_0;
	wire w_dff_A_IZaZ4JT98_0;
	wire w_dff_A_o7wAR7Kf5_0;
	wire w_dff_A_ZWrN8TAT6_0;
	wire w_dff_A_GC1pX1l39_0;
	wire w_dff_A_DAT3tjR14_0;
	wire w_dff_A_Lp3fWjAx2_0;
	wire w_dff_A_HhyK5uS78_0;
	wire w_dff_A_I6VdQDZF7_0;
	wire w_dff_A_sBPhlIxo5_0;
	wire w_dff_A_gZb17gAj1_0;
	wire w_dff_A_3eYdNwvV9_0;
	wire w_dff_A_hKabU6aP9_0;
	wire w_dff_A_GRmOsZCc2_0;
	wire w_dff_A_jOt2u3W90_0;
	wire w_dff_A_2nW35xZC6_0;
	wire w_dff_A_pEyMk4PZ2_0;
	wire w_dff_A_Ef2unXg22_0;
	wire w_dff_A_f6nhjreC0_0;
	wire w_dff_A_xoVdo85w5_1;
	wire w_dff_A_5gDDdwws1_0;
	wire w_dff_A_tDSURJ8L5_0;
	wire w_dff_A_7T47Z8Ee6_0;
	wire w_dff_A_0qzoXbNm6_0;
	wire w_dff_A_emAtNjXO1_0;
	wire w_dff_A_Gm5iDwRD3_0;
	wire w_dff_A_ijIOBYxc4_0;
	wire w_dff_A_jFEJhcw94_0;
	wire w_dff_A_JVvijcYU1_0;
	wire w_dff_A_yGx7oG0K3_0;
	wire w_dff_A_FHiqnv7H8_0;
	wire w_dff_A_f0gM1s5W2_0;
	wire w_dff_A_4iHu8ezz9_0;
	wire w_dff_A_mJY6w7js8_0;
	wire w_dff_A_LD26rznv4_0;
	wire w_dff_A_HNHrvkNo8_0;
	wire w_dff_A_Qj9BCZR75_0;
	wire w_dff_A_5czEvGOu2_0;
	wire w_dff_A_nsgSRCgU3_0;
	wire w_dff_A_okbHxb314_0;
	wire w_dff_A_5ZmMUI1l1_0;
	wire w_dff_A_6hMGT60p9_0;
	wire w_dff_A_HuYc30OT2_0;
	wire w_dff_A_NbavnChT7_0;
	wire w_dff_A_xNJ98UHb0_0;
	wire w_dff_A_7CNN2QGj1_1;
	wire w_dff_A_wPADSHmc3_0;
	wire w_dff_A_UfqHfyUg4_0;
	wire w_dff_A_XLoXWYXv6_0;
	wire w_dff_A_9CZaF95Y6_0;
	wire w_dff_A_fXX5esH14_0;
	wire w_dff_A_H6sED84P5_0;
	wire w_dff_A_ixSHJUKU4_0;
	wire w_dff_A_Ax5ViNf71_0;
	wire w_dff_A_xIk4ZfjZ1_0;
	wire w_dff_A_ww5h3tzY7_0;
	wire w_dff_A_T2WSgOqE8_0;
	wire w_dff_A_H7KwQJ684_0;
	wire w_dff_A_AB3GZso39_0;
	wire w_dff_A_tEJ9L1XR0_0;
	wire w_dff_A_XObD0KSJ3_0;
	wire w_dff_A_ftVRf9Jn2_0;
	wire w_dff_A_VfMZnpqv9_0;
	wire w_dff_A_CzQ4pz1a5_0;
	wire w_dff_A_OOAtbI1m4_0;
	wire w_dff_A_Gsx3K5yd6_0;
	wire w_dff_A_FESGzfjc1_0;
	wire w_dff_A_4E4cdKaC4_0;
	wire w_dff_A_gYgrfdEk4_0;
	wire w_dff_A_EVpZsa9A0_0;
	wire w_dff_A_kLXAngYK6_0;
	wire w_dff_A_rfiYBFTn8_1;
	wire w_dff_A_KBv17TNX9_0;
	wire w_dff_A_eYF8b48w9_0;
	wire w_dff_A_Bws8PJEh4_0;
	wire w_dff_A_3DAFSLe24_0;
	wire w_dff_A_EqiYcGl26_0;
	wire w_dff_A_kvlIc9Fz3_0;
	wire w_dff_A_6Z60N6TK4_0;
	wire w_dff_A_6FalZRrc5_0;
	wire w_dff_A_v7Zzebew6_0;
	wire w_dff_A_lDTvXDzZ3_0;
	wire w_dff_A_8yNCk5pb1_0;
	wire w_dff_A_HXlHmMDz8_0;
	wire w_dff_A_YAQm3VGj2_0;
	wire w_dff_A_TyTEpEEQ6_0;
	wire w_dff_A_GnILxcXe2_0;
	wire w_dff_A_BjlgeGGf3_0;
	wire w_dff_A_LWN4IjBz3_0;
	wire w_dff_A_7CQEVQDv5_0;
	wire w_dff_A_Svu2ui5v0_0;
	wire w_dff_A_5SUASKkG3_0;
	wire w_dff_A_vEzzzN135_0;
	wire w_dff_A_GvabwsAo3_0;
	wire w_dff_A_srrWgsu77_0;
	wire w_dff_A_o1tEZ4r95_0;
	wire w_dff_A_NhoOKTcF7_0;
	wire w_dff_A_vzwKrL7w6_1;
	wire w_dff_A_6JOIMAZh5_0;
	wire w_dff_A_HXCK9GeG6_0;
	wire w_dff_A_jnAEY3hC4_0;
	wire w_dff_A_5T71wfnt9_0;
	wire w_dff_A_RSOKYoRU9_0;
	wire w_dff_A_kMdOAi0x2_0;
	wire w_dff_A_J3I9FHX88_0;
	wire w_dff_A_zerZj92j0_0;
	wire w_dff_A_pox6fFuC4_0;
	wire w_dff_A_Duz2K8qb1_0;
	wire w_dff_A_sCyRjIMc0_0;
	wire w_dff_A_cq5ftkKE6_0;
	wire w_dff_A_YLNZXz9w3_0;
	wire w_dff_A_iEgz1ea65_0;
	wire w_dff_A_cw8y85bi0_0;
	wire w_dff_A_Uslt2Quc2_0;
	wire w_dff_A_nczOkbvE2_0;
	wire w_dff_A_LMIHyfFj4_0;
	wire w_dff_A_6chGvKM88_0;
	wire w_dff_A_bRBAi5Lb3_0;
	wire w_dff_A_OW8nLXc88_0;
	wire w_dff_A_3TrrA0Ne9_0;
	wire w_dff_A_ISuiKvfN8_0;
	wire w_dff_A_ctXFwlbt2_0;
	wire w_dff_A_7eIriKKN8_0;
	wire w_dff_A_FaNycJh43_1;
	wire w_dff_A_qGY3H2J69_0;
	wire w_dff_A_lsSkBHxA3_0;
	wire w_dff_A_GcliZzoZ7_0;
	wire w_dff_A_vV6ldDxr2_0;
	wire w_dff_A_YWZF2o7m3_0;
	wire w_dff_A_ySXUJJNC7_0;
	wire w_dff_A_HgFrOgpO1_0;
	wire w_dff_A_MCzTh2bB6_0;
	wire w_dff_A_KecxzNaP9_0;
	wire w_dff_A_BORnleMq9_0;
	wire w_dff_A_cssMt9s20_0;
	wire w_dff_A_ZnpVQHlJ1_0;
	wire w_dff_A_deleM0tD5_0;
	wire w_dff_A_ErLBn5y45_0;
	wire w_dff_A_55Q1owVA1_0;
	wire w_dff_A_LbLt0Dhv2_0;
	wire w_dff_A_LstWs4qX6_0;
	wire w_dff_A_NACdGWnd0_0;
	wire w_dff_A_O7Pr7R1k4_0;
	wire w_dff_A_GjOo3sNm4_0;
	wire w_dff_A_K2M5jAHP2_0;
	wire w_dff_A_MJuuir9n5_0;
	wire w_dff_A_robZoaqS9_0;
	wire w_dff_A_gAIBCOyk9_0;
	wire w_dff_A_AMKGO00a5_0;
	wire w_dff_A_brqg9SVn2_1;
	wire w_dff_A_i2nClWBd8_0;
	wire w_dff_A_rjGy2gj30_0;
	wire w_dff_A_8a2xj6IU7_0;
	wire w_dff_A_SIGElxjj8_0;
	wire w_dff_A_wJTkngWn6_0;
	wire w_dff_A_mLbAkSGR0_0;
	wire w_dff_A_klxBYdW41_0;
	wire w_dff_A_Xbv4C9a58_0;
	wire w_dff_A_aoc4nmTr8_0;
	wire w_dff_A_ZSaE2QXU7_0;
	wire w_dff_A_266lQG9v2_0;
	wire w_dff_A_ACClf9oO2_0;
	wire w_dff_A_xt4hKMK18_0;
	wire w_dff_A_8EV2gJwp6_0;
	wire w_dff_A_0qYkfXI60_0;
	wire w_dff_A_3JpaDPRG0_0;
	wire w_dff_A_29vsu59F3_0;
	wire w_dff_A_9K2fRsf20_0;
	wire w_dff_A_wexf8Kp48_0;
	wire w_dff_A_MOslUsCL4_0;
	wire w_dff_A_wtQqCkoa2_0;
	wire w_dff_A_JpM7Yh8f2_0;
	wire w_dff_A_WozjK2822_0;
	wire w_dff_A_oR7RuUwk7_0;
	wire w_dff_A_UJXTa3yz1_0;
	wire w_dff_A_ZwI2TXIA4_2;
	wire w_dff_A_sYOBUnNc1_0;
	wire w_dff_A_SWDkKvin7_0;
	wire w_dff_A_JjIlIpCG1_0;
	wire w_dff_A_ABN2chsT9_0;
	wire w_dff_A_Btkxkv7A9_0;
	wire w_dff_A_cwgUJgkC7_0;
	wire w_dff_A_vipA9yt70_0;
	wire w_dff_A_OdKV93LJ2_0;
	wire w_dff_A_kSn5jDc07_0;
	wire w_dff_A_KNQPhlBV5_0;
	wire w_dff_A_ZrlN9XDj7_0;
	wire w_dff_A_qHJFyHS24_0;
	wire w_dff_A_8CNmKfhf2_0;
	wire w_dff_A_zWxyZbO43_0;
	wire w_dff_A_2c8CazQk6_0;
	wire w_dff_A_3Ah7ubNf7_0;
	wire w_dff_A_m0PycPBr2_0;
	wire w_dff_A_3errfxBV5_0;
	wire w_dff_A_4lcwrkSK1_0;
	wire w_dff_A_O2j4AT3g2_0;
	wire w_dff_A_Apx7J8mW7_0;
	wire w_dff_A_e7RAeC0K0_0;
	wire w_dff_A_QjToOTvY1_0;
	wire w_dff_A_tVxoQLMN0_0;
	wire w_dff_A_7lcWiGlO9_0;
	wire w_dff_A_amYEkAj00_1;
	wire w_dff_A_LaqWwdLI9_0;
	wire w_dff_A_AKECcuck3_0;
	wire w_dff_A_RpsUUWyQ1_0;
	wire w_dff_A_eROdEdx10_0;
	wire w_dff_A_4DHT6LpY4_0;
	wire w_dff_A_5mDj9NIa8_0;
	wire w_dff_A_bw0vr69i8_0;
	wire w_dff_A_dLmmBDjx3_0;
	wire w_dff_A_vPFBJJbJ9_0;
	wire w_dff_A_Twal4M3a4_0;
	wire w_dff_A_oqWc8lh36_0;
	wire w_dff_A_U6HvmVBJ8_0;
	wire w_dff_A_aoOGWk9v8_0;
	wire w_dff_A_1Jo9rpXr5_0;
	wire w_dff_A_xQ9nMkpX1_0;
	wire w_dff_A_5SbnuXRR1_0;
	wire w_dff_A_w3mJGjV52_0;
	wire w_dff_A_7gPHDzAO7_0;
	wire w_dff_A_fUfY2IBG8_0;
	wire w_dff_A_WkWstzRA6_0;
	wire w_dff_A_8QG85tXQ5_0;
	wire w_dff_A_rPwfwKyQ7_0;
	wire w_dff_A_GnEmrQDq6_0;
	wire w_dff_A_t6zLtL210_1;
	wire w_dff_A_0GahgdHp1_0;
	wire w_dff_A_jMA16JGn6_0;
	wire w_dff_A_TDTUcUn22_0;
	wire w_dff_A_jWjxuwBj5_0;
	wire w_dff_A_lkwW53Hb9_0;
	wire w_dff_A_WpFj8LLB2_0;
	wire w_dff_A_aolWF1GW7_0;
	wire w_dff_A_GWLXQRzp2_0;
	wire w_dff_A_qO5YtnWr3_0;
	wire w_dff_A_BSs8seSw3_0;
	wire w_dff_A_OWT6ucqT4_0;
	wire w_dff_A_z4W6vr4U3_0;
	wire w_dff_A_E9n4eXgP9_0;
	wire w_dff_A_w3jBFa2V8_0;
	wire w_dff_A_OYdpdVrd2_0;
	wire w_dff_A_7wJGjD7S5_0;
	wire w_dff_A_8KaPnuhh1_0;
	wire w_dff_A_eIuhuls23_0;
	wire w_dff_A_4UfwIdWz5_0;
	wire w_dff_A_6pgKHLx60_0;
	wire w_dff_A_uyafAuev0_0;
	wire w_dff_A_ZvUt2NIY0_0;
	wire w_dff_A_Chpxamw89_0;
	wire w_dff_A_08FIgT3x3_1;
	wire w_dff_A_DEWlQHHu2_0;
	wire w_dff_A_NMtfxNaz9_0;
	wire w_dff_A_QEoySopq9_0;
	wire w_dff_A_8Q0uVE093_0;
	wire w_dff_A_ZFv72X4T8_0;
	wire w_dff_A_CXac6MEm2_0;
	wire w_dff_A_DMK9C7R25_0;
	wire w_dff_A_LQkf1OU52_0;
	wire w_dff_A_1GojHfPY9_0;
	wire w_dff_A_qRdmqRbv7_0;
	wire w_dff_A_K6kgOyaC8_0;
	wire w_dff_A_z9ssNojK7_0;
	wire w_dff_A_D9iUZg1s9_0;
	wire w_dff_A_d5h4aF7y9_0;
	wire w_dff_A_p4SBo7ed9_0;
	wire w_dff_A_OUFQjWLF5_0;
	wire w_dff_A_GKB4SBDy1_0;
	wire w_dff_A_pBwVRTGm3_0;
	wire w_dff_A_Y2ftOXnw3_0;
	wire w_dff_A_rycyxBW90_0;
	wire w_dff_A_6Hi7eGz54_0;
	wire w_dff_A_cm03bSxK5_0;
	wire w_dff_A_HanoiqVF5_0;
	wire w_dff_A_OYPAWhe44_1;
	wire w_dff_A_Dp7qLDe60_0;
	wire w_dff_A_RQOGItHR2_0;
	wire w_dff_A_qsVKNdr56_0;
	wire w_dff_A_1VrXme1e0_0;
	wire w_dff_A_Z7DtqWKy9_0;
	wire w_dff_A_AyOK5qy39_0;
	wire w_dff_A_XHSITl1N6_0;
	wire w_dff_A_25gz9LWm6_0;
	wire w_dff_A_tMyhFtJO9_0;
	wire w_dff_A_CxaKyIIo8_0;
	wire w_dff_A_CnP9KI3A0_0;
	wire w_dff_A_zsbHjANn7_0;
	wire w_dff_A_8CoC8X014_0;
	wire w_dff_A_XhWbLnqH2_0;
	wire w_dff_A_T0i8zvlZ5_0;
	wire w_dff_A_Gqjgf0B03_0;
	wire w_dff_A_vMeWpli98_0;
	wire w_dff_A_Uz9TNndU9_0;
	wire w_dff_A_XvS0LSSn0_0;
	wire w_dff_A_PPBrGKr10_0;
	wire w_dff_A_rM2fcNiD2_0;
	wire w_dff_A_OP2oINcU6_0;
	wire w_dff_A_0x6LqtEa7_0;
	wire w_dff_A_72jiinuu9_1;
	wire w_dff_A_9EfaEjWq2_0;
	wire w_dff_A_JJ9ymX5w3_0;
	wire w_dff_A_oIQSNchm2_0;
	wire w_dff_A_6GloHEU80_0;
	wire w_dff_A_dKoQ4bme0_0;
	wire w_dff_A_foZ7Xmps6_0;
	wire w_dff_A_hs7SzKHx5_0;
	wire w_dff_A_aABwAC8k3_0;
	wire w_dff_A_987uaKlJ6_0;
	wire w_dff_A_RIApDNOh1_0;
	wire w_dff_A_fFDtMKm58_0;
	wire w_dff_A_zvFqjdZP1_0;
	wire w_dff_A_F14rt1un7_0;
	wire w_dff_A_1fxqwxrk0_0;
	wire w_dff_A_rqv531aD1_0;
	wire w_dff_A_M9RJhOXS1_0;
	wire w_dff_A_s7dAlhV41_0;
	wire w_dff_A_bZDnzNKi7_0;
	wire w_dff_A_pPf9xNxG2_0;
	wire w_dff_A_YO1pMBP66_0;
	wire w_dff_A_7F4X4YAc1_0;
	wire w_dff_A_PoAmZBwf0_0;
	wire w_dff_A_bFsmNfY29_0;
	wire w_dff_A_bLpXWvvb6_0;
	wire w_dff_A_OvPuv0aa0_0;
	wire w_dff_A_VcYMcl4d4_1;
	wire w_dff_A_Yf6Mekoh8_0;
	wire w_dff_A_Yzq3GCri5_0;
	wire w_dff_A_FzC9c08i2_0;
	wire w_dff_A_BLjghiPx3_0;
	wire w_dff_A_D2MU0aDz7_0;
	wire w_dff_A_mPT6bhaT9_0;
	wire w_dff_A_yB4gbMmo9_0;
	wire w_dff_A_tF0P8ENf7_0;
	wire w_dff_A_jVbVynpX2_0;
	wire w_dff_A_sR8KRVtc9_0;
	wire w_dff_A_zYfAKsO99_0;
	wire w_dff_A_InB5Ribs0_0;
	wire w_dff_A_0lDEJ6Vf9_0;
	wire w_dff_A_uqtJAVxu4_0;
	wire w_dff_A_lackjnTj4_0;
	wire w_dff_A_C3Wea6Qn8_0;
	wire w_dff_A_INP3Vl365_0;
	wire w_dff_A_2h5znEYC7_0;
	wire w_dff_A_pDkLOFAW9_0;
	wire w_dff_A_Xovkznt48_0;
	wire w_dff_A_rR1PNAVS2_0;
	wire w_dff_A_KqK4n9an8_0;
	wire w_dff_A_zWXHBiP27_0;
	wire w_dff_A_BiNXUr146_0;
	wire w_dff_A_nbWEwK1h1_0;
	wire w_dff_A_g7IbVewx2_2;
	wire w_dff_A_5wY67q0c8_0;
	wire w_dff_A_pwJQ3Uk11_0;
	wire w_dff_A_2KxLRPgB1_0;
	wire w_dff_A_c9WI7ptW7_0;
	wire w_dff_A_l6Mr2j9G6_0;
	wire w_dff_A_gg64z5bj4_0;
	wire w_dff_A_08gqP7Sd4_0;
	wire w_dff_A_BkYoCBqS3_0;
	wire w_dff_A_4GXBB69u9_0;
	wire w_dff_A_gMYI0Bi43_0;
	wire w_dff_A_nZpA95Uc8_0;
	wire w_dff_A_xcBzd2uN8_0;
	wire w_dff_A_ZDQDla7X1_0;
	wire w_dff_A_JaYtXLZq9_0;
	wire w_dff_A_ehqFbnaG5_0;
	wire w_dff_A_B6PFfiDO5_0;
	wire w_dff_A_bt8591e34_0;
	wire w_dff_A_wtQeivoA9_0;
	wire w_dff_A_jQaCBwwH6_0;
	wire w_dff_A_JZoykD9o0_0;
	wire w_dff_A_HEctrAiX7_0;
	wire w_dff_A_8ky1ZFCm5_0;
	wire w_dff_A_N445o3Rm9_0;
	wire w_dff_A_X9VjWtUB8_0;
	wire w_dff_A_X70tw3Lb1_1;
	wire w_dff_A_ivQxTsSS9_0;
	wire w_dff_A_bbtb0N6U5_0;
	wire w_dff_A_hPzLgahQ0_0;
	wire w_dff_A_2Nla7SxG5_0;
	wire w_dff_A_mVvi4glR3_0;
	wire w_dff_A_Dzv8NsPq9_0;
	wire w_dff_A_22z3wZQn7_0;
	wire w_dff_A_s9tWOigg2_0;
	wire w_dff_A_H3DCpLJK0_0;
	wire w_dff_A_s43xw4uT1_0;
	wire w_dff_A_pywCpTOG2_0;
	wire w_dff_A_fXXipKZO0_0;
	wire w_dff_A_1Vhkare43_0;
	wire w_dff_A_3tbOnTc90_0;
	wire w_dff_A_IVfxt1M71_0;
	wire w_dff_A_SAgrBDqA8_0;
	wire w_dff_A_gruBKQpP1_0;
	wire w_dff_A_QIAjReQU7_0;
	wire w_dff_A_jUh98gZM4_0;
	wire w_dff_A_YX9ndtTA1_0;
	wire w_dff_A_AMOmrFv77_0;
	wire w_dff_A_vmednM2Z1_0;
	wire w_dff_A_9t4FJwtc1_0;
	wire w_dff_A_JqeIkt3S9_0;
	wire w_dff_A_bJdDKUnI4_0;
	wire w_dff_A_B1dnqkxZ4_2;
	wire w_dff_A_FjlWCj2b4_0;
	wire w_dff_A_Ob68xE3g0_0;
	wire w_dff_A_SRZrteZt4_0;
	wire w_dff_A_BjoHQKXg5_0;
	wire w_dff_A_Ys4vWhET0_0;
	wire w_dff_A_9U4sHRSA4_0;
	wire w_dff_A_RiaeiVOj0_0;
	wire w_dff_A_tqr91HKx9_0;
	wire w_dff_A_td3SoSxZ4_0;
	wire w_dff_A_B5xA7uuC2_0;
	wire w_dff_A_7i0u7VnG0_0;
	wire w_dff_A_uvS5cts93_0;
	wire w_dff_A_jtelvk5G4_0;
	wire w_dff_A_ffF48l0z7_0;
	wire w_dff_A_PFBddvsS8_0;
	wire w_dff_A_EoD8049A5_0;
	wire w_dff_A_qO8Kzqhg2_0;
	wire w_dff_A_K8MY7GbE9_0;
	wire w_dff_A_RVwgB2Tj4_0;
	wire w_dff_A_MQJAntPL9_0;
	wire w_dff_A_nPVIIYij4_0;
	wire w_dff_A_mpA9ibvw3_0;
	wire w_dff_A_r6dNMP9X2_0;
	wire w_dff_A_jzj3M23R2_0;
	wire w_dff_A_Ti7Z5XKL2_2;
	wire w_dff_A_XZJSgp7Q0_0;
	wire w_dff_A_6uYZIZJe3_0;
	wire w_dff_A_kWDoJ2f79_0;
	wire w_dff_A_HwwT2VBs3_0;
	wire w_dff_A_0IYeoJO08_0;
	wire w_dff_A_jYew3Hxd8_0;
	wire w_dff_A_3Q53PGQx6_0;
	wire w_dff_A_DzcVN8oE2_0;
	wire w_dff_A_atxPUGMS8_0;
	wire w_dff_A_jbFWPGkK0_0;
	wire w_dff_A_uYEAjJdY3_0;
	wire w_dff_A_WltOxQ4d6_0;
	wire w_dff_A_yq4ktUSW8_0;
	wire w_dff_A_Xr7dG80L3_0;
	wire w_dff_A_3NTHNzxg5_0;
	wire w_dff_A_eCEWwOLG8_0;
	wire w_dff_A_BQ2wGKp42_0;
	wire w_dff_A_uKEtiqzL7_0;
	wire w_dff_A_WB6mi2477_0;
	wire w_dff_A_mTDUt9HN2_0;
	wire w_dff_A_4UzhitIC0_0;
	wire w_dff_A_tVeKdouP0_0;
	wire w_dff_A_sSTDtCZF9_0;
	wire w_dff_A_w5MdrG526_1;
	wire w_dff_A_ZmDIu1cI5_0;
	wire w_dff_A_RGEZTkao7_0;
	wire w_dff_A_RowHP7Ov6_0;
	wire w_dff_A_KQ3zL1Bu0_0;
	wire w_dff_A_Z58CL2R31_0;
	wire w_dff_A_vL7Wn4443_0;
	wire w_dff_A_x2gAadT62_0;
	wire w_dff_A_frIeChTW7_0;
	wire w_dff_A_Z2Wsc5eu7_0;
	wire w_dff_A_re6X1cVW3_0;
	wire w_dff_A_mwV8252j8_0;
	wire w_dff_A_oNmloiZZ7_0;
	wire w_dff_A_7bf8dao58_0;
	wire w_dff_A_I6Pd9k5c6_0;
	wire w_dff_A_VFB3a0un3_0;
	wire w_dff_A_bnM2uTsC1_0;
	wire w_dff_A_qKiuXRsu4_0;
	wire w_dff_A_Px8UShAx9_0;
	wire w_dff_A_PDcYMmLt2_0;
	wire w_dff_A_IJyfc8eZ7_0;
	wire w_dff_A_Rau2rxJ47_0;
	wire w_dff_A_CHKqgrw39_0;
	wire w_dff_A_jJFIApff5_0;
	wire w_dff_A_TUnYOaP23_0;
	wire w_dff_A_ypRPQATu8_0;
	wire w_dff_A_KrEOdKkt7_2;
	wire w_dff_A_mVZ1O6Hg3_0;
	wire w_dff_A_OgrGov5P8_0;
	wire w_dff_A_CCfZjVuf9_0;
	wire w_dff_A_JBkwmDO49_0;
	wire w_dff_A_dd5Lt2ZD9_0;
	wire w_dff_A_JnR1XVpz2_0;
	wire w_dff_A_mfh1uOZu7_0;
	wire w_dff_A_qdpVz5IX4_0;
	wire w_dff_A_CDgFEVpt9_0;
	wire w_dff_A_aZe4e1ew5_0;
	wire w_dff_A_TGP3O5wA8_0;
	wire w_dff_A_1CjAG2pP2_0;
	wire w_dff_A_euzOGjlo0_0;
	wire w_dff_A_Vf3PdFCW9_0;
	wire w_dff_A_WuzeQQ1s7_0;
	wire w_dff_A_t8W8UlgB0_0;
	wire w_dff_A_LtRtOvmL0_0;
	wire w_dff_A_ItvX0lT74_0;
	wire w_dff_A_vLeYnClR3_0;
	wire w_dff_A_cuKXS15k1_0;
	wire w_dff_A_ERkJuYSS5_0;
	wire w_dff_A_JU682vyY6_0;
	wire w_dff_A_iq9tyi289_0;
	wire w_dff_A_WfeN12RN7_1;
	wire w_dff_A_tZyf03n89_0;
	wire w_dff_A_Gjvg1V2t4_0;
	wire w_dff_A_azWxccFr5_0;
	wire w_dff_A_CtB9QTOK3_0;
	wire w_dff_A_8ZxcYVqP1_0;
	wire w_dff_A_NtXSZeMD2_0;
	wire w_dff_A_IFbVjk4p0_0;
	wire w_dff_A_tmjihczE0_0;
	wire w_dff_A_mJaz4RL47_0;
	wire w_dff_A_jGsiy5Vs4_0;
	wire w_dff_A_cWKhQbOq7_0;
	wire w_dff_A_l2yFXSXP9_0;
	wire w_dff_A_4AJOowQ61_0;
	wire w_dff_A_Ggj6PLQA7_0;
	wire w_dff_A_sCvFeNMs8_0;
	wire w_dff_A_Pr7Qdmus9_0;
	wire w_dff_A_828TThmF2_0;
	wire w_dff_A_kMdQl0sT9_0;
	wire w_dff_A_rw9JupFW6_0;
	wire w_dff_A_6YDxurMj0_0;
	wire w_dff_A_nJBLzrFr4_0;
	wire w_dff_A_jI5PA4cr5_0;
	wire w_dff_A_8JYjHguq9_0;
	wire w_dff_A_LnjKUAvC2_0;
	wire w_dff_A_ZsdjeHLx7_0;
	wire w_dff_A_NHAxy8Qq4_2;
	wire w_dff_A_Ed2rPu1D0_0;
	wire w_dff_A_5GKxlkRZ6_0;
	wire w_dff_A_12W7fw4g4_0;
	wire w_dff_A_qnwoH1QE8_0;
	wire w_dff_A_l4jzBRgz9_0;
	wire w_dff_A_g855YBmC2_0;
	wire w_dff_A_9HW4GkQG2_0;
	wire w_dff_A_lpZiuo7Q5_0;
	wire w_dff_A_Vywao6KF8_0;
	wire w_dff_A_uB2ThT4B7_0;
	wire w_dff_A_EKIfQgUg4_0;
	wire w_dff_A_rFhaQCry4_0;
	wire w_dff_A_4lu8Ud9g5_0;
	wire w_dff_A_NsMAW75Q4_0;
	wire w_dff_A_u37X9amP7_0;
	wire w_dff_A_hIO7XOSO3_0;
	wire w_dff_A_juM6jieX6_0;
	wire w_dff_A_Kk3CIjBV7_0;
	wire w_dff_A_FvC1yZEg1_0;
	wire w_dff_A_6uv0cKzz0_0;
	wire w_dff_A_1KH2B4jk1_0;
	wire w_dff_A_aRdiGPis4_0;
	wire w_dff_A_g3TADX9Q0_0;
	wire w_dff_A_FTt1kzgv0_0;
	wire w_dff_A_616RzkKH1_0;
	wire w_dff_A_CGluyyLx8_2;
	wire w_dff_A_7g34HPfj9_0;
	wire w_dff_A_VHezfZ6H0_0;
	wire w_dff_A_AW4dAvYN2_0;
	wire w_dff_A_k30oTUpH7_0;
	wire w_dff_A_RViSHWIa6_0;
	wire w_dff_A_UkK3hfsn5_0;
	wire w_dff_A_cRyE3iZd2_0;
	wire w_dff_A_0FfUMgF40_0;
	wire w_dff_A_ffppzAl97_0;
	wire w_dff_A_7lvWxaUV1_0;
	wire w_dff_A_rDQulIv00_0;
	wire w_dff_A_2K8I8pYJ2_0;
	wire w_dff_A_duZ6ox7B9_0;
	wire w_dff_A_J9CsCj704_0;
	wire w_dff_A_IZKCF9bv4_0;
	wire w_dff_A_tUg9irBn6_0;
	wire w_dff_A_aOg81CMv9_0;
	wire w_dff_A_AOegXKqA3_0;
	wire w_dff_A_wt6Hobxm6_0;
	wire w_dff_A_Vdzrohec1_0;
	wire w_dff_A_R2YdaLCt7_2;
	wire w_dff_A_Q0JJXQ6q2_2;
	wire w_dff_A_EolVQK7x9_0;
	wire w_dff_A_sC8XpTxb0_0;
	wire w_dff_A_mlraThnj5_0;
	wire w_dff_A_hqOvNHIe1_0;
	wire w_dff_A_xBLn3BnK2_0;
	wire w_dff_A_VxpAgs9w9_0;
	wire w_dff_A_A5XS2GlF0_2;
	wire w_dff_A_NfaO50cd0_0;
	wire w_dff_A_WaQ6FwW05_0;
	wire w_dff_A_XCW9JrQp7_0;
	wire w_dff_A_B7VaiMwO9_0;
	wire w_dff_A_0qrM3nOe3_0;
	wire w_dff_A_k292zF0g9_0;
	wire w_dff_A_nl5Rctji5_2;
	wire w_dff_A_l9LCgxGv9_2;
	wire w_dff_A_kyTaRLFF9_0;
	wire w_dff_A_cYIudUaM3_0;
	wire w_dff_A_LfJ9L3gi7_0;
	wire w_dff_A_DstrArim9_0;
	wire w_dff_A_CRC1ax6O2_0;
	wire w_dff_A_RgXVgALg9_0;
	wire w_dff_A_RL0IalGz4_0;
	wire w_dff_A_lfTIEuZs4_0;
	wire w_dff_A_AXXGvaV37_0;
	wire w_dff_A_REsitmqL9_0;
	wire w_dff_A_PBnnuB6u7_0;
	wire w_dff_A_XE6rjJ8Q7_0;
	wire w_dff_A_Uw3YYzYS7_0;
	wire w_dff_A_iTOYy22w6_0;
	wire w_dff_A_f4MjxiJZ3_2;
	wire w_dff_A_YjJZ0vk19_0;
	wire w_dff_A_evzt3vR01_0;
	wire w_dff_A_jJkwxnye2_0;
	wire w_dff_A_nwtmSoKe8_0;
	wire w_dff_A_h9k8PZIV0_0;
	wire w_dff_A_L7xEiLZH9_0;
	wire w_dff_A_fOBBr3vE7_0;
	wire w_dff_A_5Dx3uy0W1_0;
	wire w_dff_A_RUKf3Paw2_0;
	wire w_dff_A_5OJnOWhJ3_0;
	wire w_dff_A_B1GN1IsM6_0;
	wire w_dff_A_mRydFenQ2_0;
	wire w_dff_A_bUZ8UM2f2_0;
	wire w_dff_A_hMRbFHPt0_0;
	wire w_dff_A_ahq94RXh2_0;
	wire w_dff_A_xb28ihKw9_0;
	wire w_dff_A_wd3queQl0_2;
	wire w_dff_A_bGy4FE5o1_0;
	wire w_dff_A_JvoLXZv29_0;
	wire w_dff_A_nc2zuewP2_0;
	wire w_dff_A_fEJYJaC64_0;
	wire w_dff_A_Bqrd55ic6_0;
	wire w_dff_A_6pg4YxwW2_0;
	wire w_dff_A_JFg8rEiJ6_0;
	wire w_dff_A_OcCMQ68y4_0;
	wire w_dff_A_pUlb9P5P1_0;
	wire w_dff_A_wSkeehsm1_0;
	wire w_dff_A_Ly7xUSq95_0;
	wire w_dff_A_r8yX35OL0_0;
	wire w_dff_A_OvuI36Xm3_0;
	wire w_dff_A_b4esieFH2_0;
	wire w_dff_A_rGQ9rEbx1_0;
	wire w_dff_A_bA3xXtm41_0;
	wire w_dff_A_fqNnckpX0_0;
	wire w_dff_A_vEddeJa75_2;
	wire w_dff_A_vmdaJfph6_0;
	wire w_dff_A_FMvSAZ0R2_0;
	wire w_dff_A_iLpUerIY1_0;
	wire w_dff_A_ZUoOI0BO5_0;
	wire w_dff_A_VYie8oKZ4_0;
	wire w_dff_A_D8skds636_0;
	wire w_dff_A_GNuP6mjp8_0;
	wire w_dff_A_z1gzQNb06_0;
	wire w_dff_A_OSTDsA4W7_0;
	wire w_dff_A_3WbuAF9l4_0;
	wire w_dff_A_xfZCYeKO1_0;
	wire w_dff_A_yg8BF1l82_0;
	wire w_dff_A_wXGwjV8M1_0;
	wire w_dff_A_4J9jGk8k2_0;
	wire w_dff_A_nYIGNC6q8_0;
	wire w_dff_A_paqg3lvO4_0;
	wire w_dff_A_STpoYxwp4_0;
	wire w_dff_A_2FJp0xsN4_0;
	wire w_dff_A_KMCbaGeF1_2;
	wire w_dff_A_q36PlStj3_0;
	wire w_dff_A_dBqpDcpe0_0;
	wire w_dff_A_hvDXOGaJ2_0;
	wire w_dff_A_Qfzya5Ze6_0;
	wire w_dff_A_bv59T8UL8_0;
	wire w_dff_A_Gd6waxCM1_0;
	wire w_dff_A_hMo2T9ni6_0;
	wire w_dff_A_IOOoSHDD5_0;
	wire w_dff_A_MJlkpX5O9_0;
	wire w_dff_A_MqYYqK3a1_0;
	wire w_dff_A_RuO7mcqB9_0;
	wire w_dff_A_dUxt6AWx7_0;
	wire w_dff_A_8VidLIuF6_2;
	wire w_dff_A_dnP6G8TY7_0;
	wire w_dff_A_FmiXhclr4_0;
	wire w_dff_A_OMstosv94_0;
	wire w_dff_A_vsPVKiou5_0;
	wire w_dff_A_1wUGljjO2_0;
	wire w_dff_A_rdtp5aFN2_0;
	wire w_dff_A_p8pYFDhF7_0;
	wire w_dff_A_aXzsrJp07_0;
	wire w_dff_A_0Bx1f9IE1_0;
	wire w_dff_A_I4jCtoFc9_0;
	wire w_dff_A_57TMX5lc6_0;
	wire w_dff_A_SJ3isSEu3_0;
	wire w_dff_A_M1p3FErj9_0;
	wire w_dff_A_f3sHIXSK4_2;
	wire w_dff_A_9WmLhrWF7_0;
	wire w_dff_A_8nnZTuLO6_0;
	wire w_dff_A_ao8l4W4i3_0;
	wire w_dff_A_NdYWOdoP6_0;
	wire w_dff_A_SeZHf1mh4_0;
	wire w_dff_A_mVqDdQf03_0;
	wire w_dff_A_Rz8PGoUa2_0;
	wire w_dff_A_MRYJka3J2_0;
	wire w_dff_A_Mzv24KvU8_0;
	wire w_dff_A_BbYuBmPy4_0;
	wire w_dff_A_E0shbqX76_0;
	wire w_dff_A_MZeBBfbI7_0;
	wire w_dff_A_zOjJnjDn1_0;
	wire w_dff_A_H03IRAWS8_2;
	wire w_dff_A_NxRbqHJi1_0;
	wire w_dff_A_kn56FF7D5_0;
	wire w_dff_A_Do8OgmES8_0;
	wire w_dff_A_507IISw87_0;
	wire w_dff_A_19jiPMKQ0_0;
	wire w_dff_A_udbXHxti9_0;
	wire w_dff_A_wfrMokYK3_0;
	wire w_dff_A_3oRT5DHU4_0;
	wire w_dff_A_MmLIGxEI6_0;
	wire w_dff_A_kT2xvXs51_0;
	wire w_dff_A_bwfAXsGr4_0;
	wire w_dff_A_La0VcisY5_0;
	wire w_dff_A_DzVLEwtQ3_0;
	wire w_dff_A_G4xBhRH19_0;
	wire w_dff_A_Z4ta4T7k2_0;
	wire w_dff_A_wykqDbm08_1;
	wire w_dff_A_9zPqFGQz7_0;
	wire w_dff_A_wc9ihYAb6_0;
	wire w_dff_A_KSSYnzCg4_0;
	wire w_dff_A_JEMkHivD3_0;
	wire w_dff_A_wwXYz9bQ8_0;
	wire w_dff_A_fJtPq6tq7_0;
	wire w_dff_A_1EZv6f307_0;
	wire w_dff_A_W2Pe5qtY8_0;
	wire w_dff_A_lpC5Yjxz4_0;
	wire w_dff_A_AXYOX6if8_0;
	wire w_dff_A_zoXH8DyH0_0;
	wire w_dff_A_AYx6ANXW1_0;
	wire w_dff_A_bCsRiVss5_0;
	wire w_dff_A_12cptL5E3_0;
	wire w_dff_A_tgV96mPK7_0;
	wire w_dff_A_nyyEt9jd2_1;
	wire w_dff_A_pkJ0GkZQ3_0;
	wire w_dff_A_trM5DOrX7_0;
	wire w_dff_A_ZHXGwIji4_0;
	wire w_dff_A_ydPQZw6P4_0;
	wire w_dff_A_KZ876fa08_0;
	wire w_dff_A_KCQfCrxM3_0;
	wire w_dff_A_8I9NFbmK2_0;
	wire w_dff_A_2VFTo9823_0;
	wire w_dff_A_f8kk55bC7_0;
	wire w_dff_A_E0G0wta24_0;
	wire w_dff_A_AJCzSzAi8_0;
	wire w_dff_A_uu30PPq45_0;
	wire w_dff_A_l36IXXuE2_0;
	wire w_dff_A_7yOlvR0b9_0;
	wire w_dff_A_cJ8tRCMf1_0;
	wire w_dff_A_5Phao2qY9_1;
	wire w_dff_A_SlpxzlWo9_0;
	wire w_dff_A_IPLLeTBj4_0;
	wire w_dff_A_9HxK52q10_0;
	wire w_dff_A_ZIlnqiwe7_0;
	wire w_dff_A_Y6Rgkjl59_0;
	wire w_dff_A_BLZDHSPz7_0;
	wire w_dff_A_dtQrnXPr1_0;
	wire w_dff_A_xtdju5j15_0;
	wire w_dff_A_RUF0Bp9h5_0;
	wire w_dff_A_gGKKYrL76_0;
	wire w_dff_A_eZsSL7no0_0;
	wire w_dff_A_JgCU2Fav8_0;
	wire w_dff_A_IFN6ScqP4_0;
	wire w_dff_A_hMJWlTAb8_2;
	wire w_dff_A_7iyGzNrG8_0;
	wire w_dff_A_HRHixrIo2_0;
	wire w_dff_A_IShvtZLt9_0;
	wire w_dff_A_AACjyD1C0_0;
	wire w_dff_A_dz6pocrP5_0;
	wire w_dff_A_oXOkdpwq9_0;
	wire w_dff_A_k8fwsG6X8_2;
	wire w_dff_A_GI0MnWIo1_0;
	wire w_dff_A_Otjvdvdr9_0;
	wire w_dff_A_EZQyUxsP2_0;
	wire w_dff_A_e9EVMRV11_0;
	wire w_dff_A_nvdRjiDF3_0;
	wire w_dff_A_kdjx6fiP2_0;
	wire w_dff_A_r89USscb9_0;
	wire w_dff_A_6if8DXLV5_0;
	wire w_dff_A_ncsEIN7l2_0;
	wire w_dff_A_ouDDPZkR1_2;
	wire w_dff_A_I97Xg4N51_0;
	wire w_dff_A_zYoIwaxo4_0;
	wire w_dff_A_Cle7SSIO7_0;
	wire w_dff_A_rf51OD4G6_0;
	wire w_dff_A_6x2DiZCh2_0;
	wire w_dff_A_y1lICjJJ6_2;
	wire w_dff_A_xV6enaR67_0;
	wire w_dff_A_aYv5HA7j9_0;
	wire w_dff_A_V1Y6LPsY3_0;
	wire w_dff_A_Uy4DScXa9_0;
	wire w_dff_A_r0NcR0A47_0;
	wire w_dff_A_lgpTcbSX8_0;
	wire w_dff_A_jsap1kaJ3_0;
	wire w_dff_A_Tsmut07i4_0;
	wire w_dff_A_NfzkrZUl7_0;
	wire w_dff_A_kfLFkw6M5_2;
	wire w_dff_A_ACqslBCv7_2;
	wire w_dff_A_Y4t8sdBm8_0;
	wire w_dff_A_kifR7LAe6_0;
	wire w_dff_A_uw9UyzKk2_0;
	wire w_dff_A_Bo9l5qom6_0;
	wire w_dff_A_pHtuYwCX5_0;
	wire w_dff_A_u94kLzpL1_2;
	wire w_dff_A_7l6AgJFW3_0;
	wire w_dff_A_ruIjEfsc5_0;
	wire w_dff_A_eGCBi7UI3_0;
	wire w_dff_A_IMsKFPMu0_0;
	wire w_dff_A_BkSUfK953_0;
	wire w_dff_A_S7sW2fzJ2_0;
	wire w_dff_A_iJCHvIYW2_2;
	wire w_dff_A_DwVU4p0z8_0;
	wire w_dff_A_RxdP6a0E7_0;
	wire w_dff_A_t5Uihtn31_0;
	wire w_dff_A_THjpltkp3_0;
	wire w_dff_A_a5BYp71V9_0;
	wire w_dff_A_eKNM7vN50_0;
	wire w_dff_A_7WMxIowz2_0;
	wire w_dff_A_IhK2kk8i6_2;
	wire w_dff_A_KDAv0QYT0_0;
	wire w_dff_A_j0C65L6g2_0;
	wire w_dff_A_aVSyyIGQ5_0;
	wire w_dff_A_4AYGEmap7_0;
	wire w_dff_A_xI4IW2bo6_0;
	wire w_dff_A_h8Q04HCz0_0;
	wire w_dff_A_yZTlQUTQ7_0;
	wire w_dff_A_IyoCa8wx8_2;
	wire w_dff_A_NvrgdMKU2_0;
	wire w_dff_A_HUfgb5F17_2;
	wire w_dff_A_WZFDRTZ02_0;
	wire w_dff_A_UgHHmDTh0_0;
	wire w_dff_A_56MDtBHq7_2;
	wire w_dff_A_YMbsQHww3_0;
	wire w_dff_A_eoKninLD1_0;
	wire w_dff_A_jVNl1AUr1_0;
	wire w_dff_A_bmy2DIyV3_2;
	wire w_dff_A_DmiOXxqU7_0;
	wire w_dff_A_MrFmcRjM9_0;
	wire w_dff_A_Faa1tfed9_0;
	wire w_dff_A_jhWvCLTd0_2;
	wire w_dff_A_DOhhlZFY7_0;
	wire w_dff_A_IydLM9Go8_0;
	wire w_dff_A_r7pMVeiv4_0;
	wire w_dff_A_W32TXfhs9_0;
	wire w_dff_A_89CIiKXN0_0;
	wire w_dff_A_yTIIXXdG2_0;
	wire w_dff_A_n4QvVDPh2_0;
	wire w_dff_A_DmSxY9v33_0;
	wire w_dff_A_JZZMLKg54_0;
	wire w_dff_A_mmQlEfuy6_0;
	wire w_dff_A_8zlm28G46_0;
	wire w_dff_A_FoWZznBm6_2;
	wire w_dff_A_bXHu9UF51_2;
	wire w_dff_A_Yexk4taD4_0;
	wire w_dff_A_9IN6LYZ30_0;
	wire w_dff_A_3ubhS1Ve3_0;
	wire w_dff_A_kO1eFYA95_2;
	wire w_dff_A_KvSYlQtB0_0;
	wire w_dff_A_2e7Pzvlt4_0;
	wire w_dff_A_wI0jkKM02_0;
	wire w_dff_A_pq520oT52_0;
	wire w_dff_A_FQeftoZR1_0;
	wire w_dff_A_QNPL4Nn99_2;
	wire w_dff_A_eF8HMsmM0_0;
	wire w_dff_A_nVo2cKWp6_0;
	wire w_dff_A_wMRy0g015_0;
	wire w_dff_A_JqoY9hF47_0;
	wire w_dff_A_15EPoaaV9_0;
	wire w_dff_A_GtDw502C2_2;
	wire w_dff_A_idBcVgJA1_0;
	wire w_dff_A_QW7ti7wh7_0;
	wire w_dff_A_F74uv20G6_0;
	wire w_dff_A_4at4GPYc7_0;
	wire w_dff_A_gmPvQ6Lp0_0;
	wire w_dff_A_7tF7lrrX4_0;
	wire w_dff_A_CLY8YUQh0_0;
	wire w_dff_A_u2VS0eu85_2;
	wire w_dff_A_0WEmXAVP9_0;
	wire w_dff_A_AmHEvaNU2_0;
	wire w_dff_A_DVNHGDkx9_0;
	wire w_dff_A_PZYJlCxG8_0;
	wire w_dff_A_hgG319v29_0;
	wire w_dff_A_XGIEQCg10_0;
	wire w_dff_A_SpyAcNEH9_0;
	wire w_dff_A_nRWXLRke4_0;
	wire w_dff_A_r2jAo6Mu9_0;
	wire w_dff_A_vN0bMFAx7_0;
	wire w_dff_A_dGxuGP4h3_0;
	wire w_dff_A_dflpMAFK7_0;
	wire w_dff_A_d63CencI3_0;
	wire w_dff_A_u8189vHk1_2;
	wire w_dff_A_KJykaV3M0_2;
	wire w_dff_A_pN6IxNGh5_2;
	wire w_dff_A_TeChXTMa7_0;
	wire w_dff_A_ikIdkQUw3_0;
	wire w_dff_A_EoeqTSWy8_0;
	wire w_dff_A_E8jalRTs2_2;
	wire w_dff_A_wfUaDLW66_0;
	wire w_dff_A_arKIhtye4_0;
	wire w_dff_A_QzOwvaFh3_0;
	wire w_dff_A_Qutbbi7W3_2;
	wire w_dff_A_j9wtRz0k2_0;
	wire w_dff_A_zB9ZqTqK2_0;
	wire w_dff_A_bwLEuQlq6_0;
	wire w_dff_A_U7c5MoiX0_0;
	wire w_dff_A_gi4w7YCi8_0;
	wire w_dff_A_J5yOHCRL9_0;
	wire w_dff_A_i45KJBzy6_0;
	wire w_dff_A_AQx62qQL1_0;
	wire w_dff_A_Xe1ad79S1_0;
	wire w_dff_A_QxgVD2QB2_2;
	wire w_dff_A_zgWesmuJ1_0;
	wire w_dff_A_aaoXjhMP0_0;
	wire w_dff_A_FiiC9BSW1_0;
	wire w_dff_A_m5y08wEu6_0;
	wire w_dff_A_5dlFzehl4_0;
	wire w_dff_A_HRaAPMWW8_0;
	wire w_dff_A_z4W1hAW05_0;
	wire w_dff_A_SphUPevv8_0;
	wire w_dff_A_dqPJ984U6_0;
	wire w_dff_A_6FJsb1lw2_0;
	wire w_dff_A_OEN3E7xB2_2;
	wire w_dff_A_FBPSAZrq3_0;
	wire w_dff_A_73WPHF0a8_0;
	wire w_dff_A_ugyj3iQ65_0;
	wire w_dff_A_ZZ2Y7ZiW0_0;
	wire w_dff_A_EklCC1Fx2_0;
	wire w_dff_A_hdHDfOPH7_0;
	wire w_dff_A_Gb0kjhg59_0;
	wire w_dff_A_oQuZ9C3o7_0;
	wire w_dff_A_HdHLYKd25_0;
	wire w_dff_A_4YZ7HJAB9_0;
	wire w_dff_A_LLUDcLli2_0;
	wire w_dff_A_BRr7V1Dd0_2;
	wire w_dff_A_bTLj5nNy8_0;
	wire w_dff_A_5waj8wW36_0;
	wire w_dff_A_RMkVxy4D8_0;
	wire w_dff_A_jVXSzJcQ9_0;
	wire w_dff_A_AOsmoC2R4_0;
	wire w_dff_A_3e1Lm0s86_0;
	wire w_dff_A_1HCHJbDg8_0;
	wire w_dff_A_0T8uOQtH3_0;
	wire w_dff_A_kJM8BYLq2_0;
	wire w_dff_A_cHjh7vKg0_0;
	wire w_dff_A_mPaS6Mha1_0;
	wire w_dff_A_VimgZs4n3_2;
	wire w_dff_A_3PbZ1Jbq8_0;
	wire w_dff_A_zXS4Xfyi0_0;
	wire w_dff_A_GRpvyfWq5_0;
	wire w_dff_A_psKGp7Cq9_0;
	wire w_dff_A_lxkcQEtM0_0;
	wire w_dff_A_Q58gQSBR2_0;
	wire w_dff_A_ekUOwAko3_0;
	wire w_dff_A_dx0HSNzG9_0;
	wire w_dff_A_djG7tKrZ7_2;
	wire w_dff_A_ghteABgK6_0;
	wire w_dff_A_Ab0KCW1j2_0;
	wire w_dff_A_pZELC5nk3_0;
	wire w_dff_A_9iZodpNr8_0;
	wire w_dff_A_IVFAHnMD3_0;
	wire w_dff_A_VIktzUjc1_0;
	wire w_dff_A_GjlOPqmp8_0;
	wire w_dff_A_6Y8UhFqg3_0;
	wire w_dff_A_CzzP5pjZ0_0;
	wire w_dff_A_P8hPtzqU4_2;
	wire w_dff_A_9ybG1xG72_0;
	wire w_dff_A_21VOdRlb4_0;
	wire w_dff_A_ALy7YhUb2_0;
	wire w_dff_A_WrKJH55W6_0;
	wire w_dff_A_ieoW1bNp6_0;
	wire w_dff_A_ea7jBFts1_0;
	wire w_dff_A_0iF253ta6_0;
	wire w_dff_A_Z3sOWuaz0_0;
	wire w_dff_A_rw5qINAa0_0;
	wire w_dff_A_ypcAw9sg9_2;
	wire w_dff_A_mOswMUxg3_0;
	wire w_dff_A_tIzFAeLt4_0;
	wire w_dff_A_7BPlkgWi9_0;
	wire w_dff_A_dAgHZCA45_0;
	wire w_dff_A_QWZOHusX0_0;
	wire w_dff_A_E1az6nZ82_0;
	wire w_dff_A_XiIHYqRH8_0;
	wire w_dff_A_OsqvV3eo7_0;
	wire w_dff_A_38FS1zn56_0;
	wire w_dff_A_y6MjP8Qb8_0;
	wire w_dff_A_nv0Y42PX8_0;
	wire w_dff_A_O0ichDPW1_2;
	wire w_dff_A_PtgjT43b1_0;
	wire w_dff_A_IOZH2WS93_0;
	wire w_dff_A_jfawbR8f2_0;
	wire w_dff_A_LEzamXti6_0;
	wire w_dff_A_p7vnaGTp4_2;
	wire w_dff_A_yDtmijmt8_0;
	wire w_dff_A_5B511Ywc8_0;
	wire w_dff_A_Y0TP6KzS4_0;
	wire w_dff_A_8x9IJLGt1_0;
	wire w_dff_A_reD76IVv3_0;
	wire w_dff_A_T0RPmTc91_0;
	wire w_dff_A_neBD5Ml89_2;
	wire w_dff_A_LeXqoUCC1_0;
	wire w_dff_A_tlVoCh1Z5_0;
	wire w_dff_A_uh82oImW5_0;
	wire w_dff_A_BG2uy8SX9_0;
	jnot g0000(.din(w_G15_0[2]),.dout(w_dff_A_rfiYBFTn8_1),.clk(gclk));
	jor g0001(.dina(G57),.dinb(w_G5_1[2]),.dout(w_dff_A_ZwI2TXIA4_2),.clk(gclk));
	jnot g0002(.din(G184),.dout(n317),.clk(gclk));
	jnot g0003(.din(G228),.dout(n318),.clk(gclk));
	jor g0004(.dina(n318),.dinb(n317),.dout(n319),.clk(gclk));
	jnot g0005(.din(G150),.dout(n320),.clk(gclk));
	jnot g0006(.din(G240),.dout(n321),.clk(gclk));
	jor g0007(.dina(n321),.dinb(n320),.dout(n322),.clk(gclk));
	jor g0008(.dina(n322),.dinb(n319),.dout(G404_fa_),.clk(gclk));
	jnot g0009(.din(G210),.dout(n324),.clk(gclk));
	jnot g0010(.din(G218),.dout(n325),.clk(gclk));
	jor g0011(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jnot g0012(.din(G152),.dout(n327),.clk(gclk));
	jnot g0013(.din(G230),.dout(n328),.clk(gclk));
	jor g0014(.dina(n328),.dinb(n327),.dout(n329),.clk(gclk));
	jor g0015(.dina(n329),.dinb(n326),.dout(G406_fa_),.clk(gclk));
	jnot g0016(.din(G183),.dout(n331),.clk(gclk));
	jnot g0017(.din(G185),.dout(n332),.clk(gclk));
	jor g0018(.dina(n332),.dinb(n331),.dout(n333),.clk(gclk));
	jnot g0019(.din(G182),.dout(n334),.clk(gclk));
	jnot g0020(.din(G186),.dout(n335),.clk(gclk));
	jor g0021(.dina(n335),.dinb(n334),.dout(n336),.clk(gclk));
	jor g0022(.dina(n336),.dinb(n333),.dout(G408_fa_),.clk(gclk));
	jnot g0023(.din(G172),.dout(n338),.clk(gclk));
	jnot g0024(.din(G188),.dout(n339),.clk(gclk));
	jor g0025(.dina(n339),.dinb(n338),.dout(n340),.clk(gclk));
	jnot g0026(.din(G162),.dout(n341),.clk(gclk));
	jnot g0027(.din(G199),.dout(n342),.clk(gclk));
	jor g0028(.dina(n342),.dinb(n341),.dout(n343),.clk(gclk));
	jor g0029(.dina(n343),.dinb(n340),.dout(G410_fa_),.clk(gclk));
	jnot g0030(.din(G1197),.dout(n345),.clk(gclk));
	jor g0031(.dina(w_n345_0[1]),.dinb(w_G5_1[1]),.dout(w_dff_A_g7IbVewx2_2),.clk(gclk));
	jnot g0032(.din(G133),.dout(n347),.clk(gclk));
	jdff g0033(.din(G134),.dout(n348),.clk(gclk));
	jor g0034(.dina(n348),.dinb(n347),.dout(n349),.clk(gclk));
	jor g0035(.dina(w_n349_0[1]),.dinb(w_G5_1[0]),.dout(w_dff_A_Ti7Z5XKL2_2),.clk(gclk));
	jand g0036(.dina(G163),.dinb(w_G1_1[2]),.dout(w_dff_A_NHAxy8Qq4_2),.clk(gclk));
	jnot g0037(.din(w_G41_0[2]),.dout(n352),.clk(gclk));
	jor g0038(.dina(n352),.dinb(w_G18_58[2]),.dout(n353),.clk(gclk));
	jor g0039(.dina(w_n353_0[2]),.dinb(w_G3701_1[1]),.dout(n354),.clk(gclk));
	jnot g0040(.din(w_G18_58[1]),.dout(n355),.clk(gclk));
	jand g0041(.dina(w_G41_0[1]),.dinb(w_n355_26[1]),.dout(n356),.clk(gclk));
	jor g0042(.dina(w_G229_0[1]),.dinb(w_G18_58[0]),.dout(n357),.clk(gclk));
	jor g0043(.dina(w_dff_B_qH8YMZAq3_0),.dinb(w_n356_0[2]),.dout(n358),.clk(gclk));
	jand g0044(.dina(w_G3701_1[0]),.dinb(w_n355_26[0]),.dout(n359),.clk(gclk));
	jnot g0045(.din(w_n359_0[1]),.dout(n360),.clk(gclk));
	jor g0046(.dina(n360),.dinb(w_n358_0[1]),.dout(n361),.clk(gclk));
	jand g0047(.dina(n361),.dinb(w_n354_1[2]),.dout(n362),.clk(gclk));
	jxor g0048(.dina(w_n362_0[2]),.dinb(w_G4526_1[1]),.dout(w_dff_A_CGluyyLx8_2),.clk(gclk));
	jand g0049(.dina(w_G4528_0[2]),.dinb(w_G1496_0[2]),.dout(n364),.clk(gclk));
	jxor g0050(.dina(w_n364_0[1]),.dinb(w_G38_1[2]),.dout(n365),.clk(gclk));
	jnot g0051(.din(w_G3723_1[1]),.dout(n366),.clk(gclk));
	jand g0052(.dina(G235),.dinb(w_G18_57[2]),.dout(n367),.clk(gclk));
	jnot g0053(.din(n367),.dout(n368),.clk(gclk));
	jnot g0054(.din(G103),.dout(n369),.clk(gclk));
	jor g0055(.dina(n369),.dinb(w_G18_57[1]),.dout(n370),.clk(gclk));
	jand g0056(.dina(w_n370_0[1]),.dinb(n368),.dout(n371),.clk(gclk));
	jxor g0057(.dina(w_n371_1[1]),.dinb(w_n366_0[1]),.dout(n372),.clk(gclk));
	jand g0058(.dina(G236),.dinb(w_G18_57[0]),.dout(n373),.clk(gclk));
	jnot g0059(.din(n373),.dout(n374),.clk(gclk));
	jnot g0060(.din(G23),.dout(n375),.clk(gclk));
	jor g0061(.dina(n375),.dinb(w_G18_56[2]),.dout(n376),.clk(gclk));
	jand g0062(.dina(w_n376_0[1]),.dinb(n374),.dout(n377),.clk(gclk));
	jnot g0063(.din(w_n377_1[2]),.dout(n378),.clk(gclk));
	jxor g0064(.dina(n378),.dinb(w_G3717_2[1]),.dout(n379),.clk(gclk));
	jor g0065(.dina(w_n379_1[1]),.dinb(w_n372_1[2]),.dout(n380),.clk(gclk));
	jnot g0066(.din(w_G3711_1[1]),.dout(n381),.clk(gclk));
	jand g0067(.dina(G237),.dinb(w_G18_56[1]),.dout(n382),.clk(gclk));
	jnot g0068(.din(n382),.dout(n383),.clk(gclk));
	jnot g0069(.din(G26),.dout(n384),.clk(gclk));
	jor g0070(.dina(n384),.dinb(w_G18_56[0]),.dout(n385),.clk(gclk));
	jand g0071(.dina(w_n385_0[1]),.dinb(n383),.dout(n386),.clk(gclk));
	jxor g0072(.dina(w_n386_0[2]),.dinb(w_dff_B_Lmpe7ff84_1),.dout(n387),.clk(gclk));
	jnot g0073(.din(w_G4526_1[0]),.dout(n388),.clk(gclk));
	jnot g0074(.din(w_G3701_0[2]),.dout(n389),.clk(gclk));
	jand g0075(.dina(w_n356_0[1]),.dinb(w_n389_0[1]),.dout(n390),.clk(gclk));
	jnot g0076(.din(w_G229_0[0]),.dout(n391),.clk(gclk));
	jor g0077(.dina(n391),.dinb(w_n355_25[2]),.dout(n392),.clk(gclk));
	jand g0078(.dina(n392),.dinb(w_n353_0[1]),.dout(n393),.clk(gclk));
	jand g0079(.dina(w_n359_0[0]),.dinb(n393),.dout(n394),.clk(gclk));
	jor g0080(.dina(n394),.dinb(w_n390_1[1]),.dout(n395),.clk(gclk));
	jnot g0081(.din(w_G3705_2[1]),.dout(n396),.clk(gclk));
	jnot g0082(.din(G238),.dout(n397),.clk(gclk));
	jor g0083(.dina(n397),.dinb(w_n355_25[1]),.dout(n398),.clk(gclk));
	jnot g0084(.din(G29),.dout(n399),.clk(gclk));
	jor g0085(.dina(n399),.dinb(w_G18_55[2]),.dout(n400),.clk(gclk));
	jand g0086(.dina(w_n400_0[1]),.dinb(n398),.dout(n401),.clk(gclk));
	jxor g0087(.dina(w_n401_1[2]),.dinb(w_dff_B_sTsRkrCo0_1),.dout(n402),.clk(gclk));
	jor g0088(.dina(w_n402_1[1]),.dinb(w_n395_0[2]),.dout(n403),.clk(gclk));
	jor g0089(.dina(w_n403_0[1]),.dinb(w_n388_0[2]),.dout(n404),.clk(gclk));
	jor g0090(.dina(w_n404_0[1]),.dinb(w_n387_1[2]),.dout(n405),.clk(gclk));
	jor g0091(.dina(w_n405_0[2]),.dinb(w_n380_0[2]),.dout(n406),.clk(gclk));
	jor g0092(.dina(w_n386_0[1]),.dinb(w_G3711_1[0]),.dout(n407),.clk(gclk));
	jor g0093(.dina(w_n402_1[0]),.dinb(w_n354_1[1]),.dout(n408),.clk(gclk));
	jor g0094(.dina(w_n408_0[1]),.dinb(w_n387_1[1]),.dout(n409),.clk(gclk));
	jand g0095(.dina(n409),.dinb(w_n407_0[2]),.dout(n410),.clk(gclk));
	jor g0096(.dina(w_n410_0[1]),.dinb(w_n380_0[1]),.dout(n411),.clk(gclk));
	jor g0097(.dina(w_n401_1[1]),.dinb(w_G3705_2[0]),.dout(n412),.clk(gclk));
	jor g0098(.dina(w_n412_0[2]),.dinb(w_n387_1[0]),.dout(n413),.clk(gclk));
	jor g0099(.dina(w_n413_1[1]),.dinb(w_n380_0[0]),.dout(n414),.clk(gclk));
	jor g0100(.dina(w_n371_1[0]),.dinb(w_G3723_1[0]),.dout(n415),.clk(gclk));
	jand g0101(.dina(w_n371_0[2]),.dinb(w_G3723_0[2]),.dout(n416),.clk(gclk));
	jor g0102(.dina(w_n377_1[1]),.dinb(w_G3717_2[0]),.dout(n417),.clk(gclk));
	jor g0103(.dina(w_n417_0[2]),.dinb(n416),.dout(n418),.clk(gclk));
	jand g0104(.dina(n418),.dinb(w_dff_B_5GHdNSKJ6_1),.dout(n419),.clk(gclk));
	jand g0105(.dina(w_n419_0[1]),.dinb(n414),.dout(n420),.clk(gclk));
	jand g0106(.dina(n420),.dinb(n411),.dout(n421),.clk(gclk));
	jand g0107(.dina(n421),.dinb(n406),.dout(n422),.clk(gclk));
	jnot g0108(.din(w_G3737_1[1]),.dout(n423),.clk(gclk));
	jand g0109(.dina(G233),.dinb(w_G18_55[1]),.dout(n424),.clk(gclk));
	jnot g0110(.din(n424),.dout(n425),.clk(gclk));
	jnot g0111(.din(G127),.dout(n426),.clk(gclk));
	jor g0112(.dina(n426),.dinb(w_G18_55[0]),.dout(n427),.clk(gclk));
	jand g0113(.dina(w_n427_0[1]),.dinb(n425),.dout(n428),.clk(gclk));
	jxor g0114(.dina(w_n428_0[2]),.dinb(w_dff_B_l6O1nGen5_1),.dout(n429),.clk(gclk));
	jnot g0115(.din(w_G3729_1[1]),.dout(n430),.clk(gclk));
	jand g0116(.dina(G234),.dinb(w_G18_54[2]),.dout(n431),.clk(gclk));
	jnot g0117(.din(n431),.dout(n432),.clk(gclk));
	jnot g0118(.din(G130),.dout(n433),.clk(gclk));
	jor g0119(.dina(n433),.dinb(w_G18_54[1]),.dout(n434),.clk(gclk));
	jand g0120(.dina(w_n434_0[1]),.dinb(n432),.dout(n435),.clk(gclk));
	jxor g0121(.dina(w_n435_1[1]),.dinb(w_n430_0[1]),.dout(n436),.clk(gclk));
	jor g0122(.dina(w_n436_0[1]),.dinb(w_n429_2[1]),.dout(n437),.clk(gclk));
	jand g0123(.dina(G231),.dinb(w_G18_54[0]),.dout(n438),.clk(gclk));
	jnot g0124(.din(n438),.dout(n439),.clk(gclk));
	jnot g0125(.din(G100),.dout(n440),.clk(gclk));
	jor g0126(.dina(n440),.dinb(w_G18_53[2]),.dout(n441),.clk(gclk));
	jand g0127(.dina(w_n441_0[1]),.dinb(n439),.dout(n442),.clk(gclk));
	jor g0128(.dina(w_n442_0[2]),.dinb(w_G3749_1[1]),.dout(n443),.clk(gclk));
	jnot g0129(.din(w_n443_0[1]),.dout(n444),.clk(gclk));
	jand g0130(.dina(w_n442_0[1]),.dinb(w_G3749_1[0]),.dout(n445),.clk(gclk));
	jor g0131(.dina(w_n445_0[1]),.dinb(n444),.dout(n446),.clk(gclk));
	jand g0132(.dina(G232),.dinb(w_G18_53[1]),.dout(n447),.clk(gclk));
	jand g0133(.dina(w_dff_B_hcyQBnBz9_0),.dinb(w_n355_25[0]),.dout(n448),.clk(gclk));
	jor g0134(.dina(w_n448_0[1]),.dinb(w_dff_B_44dd0rRk9_1),.dout(n449),.clk(gclk));
	jxor g0135(.dina(w_n449_0[2]),.dinb(w_G3743_1[2]),.dout(n450),.clk(gclk));
	jor g0136(.dina(w_n450_0[2]),.dinb(w_n446_1[1]),.dout(n451),.clk(gclk));
	jor g0137(.dina(n451),.dinb(w_n437_0[1]),.dout(n452),.clk(gclk));
	jor g0138(.dina(w_n452_0[1]),.dinb(w_n422_1[2]),.dout(n453),.clk(gclk));
	jnot g0139(.din(w_n449_0[1]),.dout(n454),.clk(gclk));
	jor g0140(.dina(w_n454_0[1]),.dinb(w_G3743_1[1]),.dout(n455),.clk(gclk));
	jand g0141(.dina(w_n454_0[0]),.dinb(w_G3743_1[0]),.dout(n456),.clk(gclk));
	jor g0142(.dina(w_n428_0[1]),.dinb(w_G3737_1[0]),.dout(n457),.clk(gclk));
	jor g0143(.dina(w_n435_1[0]),.dinb(w_G3729_1[0]),.dout(n458),.clk(gclk));
	jor g0144(.dina(w_n458_0[2]),.dinb(w_n429_2[0]),.dout(n459),.clk(gclk));
	jand g0145(.dina(n459),.dinb(w_n457_0[1]),.dout(n460),.clk(gclk));
	jor g0146(.dina(w_n460_0[2]),.dinb(w_n456_0[2]),.dout(n461),.clk(gclk));
	jand g0147(.dina(w_n461_0[1]),.dinb(w_n455_0[1]),.dout(n462),.clk(gclk));
	jand g0148(.dina(w_n462_0[2]),.dinb(w_n443_0[0]),.dout(n463),.clk(gclk));
	jor g0149(.dina(n463),.dinb(w_n445_0[0]),.dout(n464),.clk(gclk));
	jand g0150(.dina(w_n464_0[1]),.dinb(n453),.dout(n465),.clk(gclk));
	jnot g0151(.din(w_G4415_1[1]),.dout(n466),.clk(gclk));
	jand g0152(.dina(G223),.dinb(w_G18_53[0]),.dout(n467),.clk(gclk));
	jand g0153(.dina(w_dff_B_Bzm4aaA47_0),.dinb(w_n355_24[2]),.dout(n468),.clk(gclk));
	jor g0154(.dina(w_n468_0[1]),.dinb(w_dff_B_wSeJvHvY2_1),.dout(n469),.clk(gclk));
	jxor g0155(.dina(w_n469_1[1]),.dinb(w_n466_0[1]),.dout(n470),.clk(gclk));
	jnot g0156(.din(w_G4400_0[2]),.dout(n471),.clk(gclk));
	jand g0157(.dina(G226),.dinb(w_G18_52[2]),.dout(n472),.clk(gclk));
	jand g0158(.dina(w_dff_B_Y2u8jKVw1_0),.dinb(w_n355_24[1]),.dout(n473),.clk(gclk));
	jor g0159(.dina(w_n473_0[1]),.dinb(w_dff_B_QMTRnMAr5_1),.dout(n474),.clk(gclk));
	jxor g0160(.dina(w_n474_1[1]),.dinb(w_n471_0[2]),.dout(n475),.clk(gclk));
	jand g0161(.dina(G217),.dinb(w_G18_52[1]),.dout(n476),.clk(gclk));
	jand g0162(.dina(w_dff_B_EYX6X5V06_0),.dinb(w_n355_24[0]),.dout(n477),.clk(gclk));
	jor g0163(.dina(w_n477_0[1]),.dinb(w_dff_B_I7HteV6h8_1),.dout(n478),.clk(gclk));
	jnot g0164(.din(w_n478_0[1]),.dout(n479),.clk(gclk));
	jxor g0165(.dina(w_n479_0[1]),.dinb(w_G4394_1[1]),.dout(n480),.clk(gclk));
	jand g0166(.dina(w_n480_1[1]),.dinb(w_n475_1[1]),.dout(n481),.clk(gclk));
	jnot g0167(.din(w_G4410_1[1]),.dout(n482),.clk(gclk));
	jand g0168(.dina(G224),.dinb(w_G18_52[0]),.dout(n483),.clk(gclk));
	jand g0169(.dina(w_dff_B_r7ZZahyA5_0),.dinb(w_n355_23[2]),.dout(n484),.clk(gclk));
	jor g0170(.dina(w_n484_0[1]),.dinb(w_dff_B_JjtPmCHB3_1),.dout(n485),.clk(gclk));
	jxor g0171(.dina(w_n485_0[2]),.dinb(w_n482_0[1]),.dout(n486),.clk(gclk));
	jand g0172(.dina(G225),.dinb(w_G18_51[2]),.dout(n487),.clk(gclk));
	jand g0173(.dina(w_dff_B_0QEtDJod2_0),.dinb(w_n355_23[1]),.dout(n488),.clk(gclk));
	jor g0174(.dina(w_n488_0[1]),.dinb(w_dff_B_5hU4vHiZ8_1),.dout(n489),.clk(gclk));
	jnot g0175(.din(w_n489_0[1]),.dout(n490),.clk(gclk));
	jxor g0176(.dina(w_n490_0[2]),.dinb(w_G4405_1[2]),.dout(n491),.clk(gclk));
	jand g0177(.dina(w_n491_1[1]),.dinb(w_n486_0[2]),.dout(n492),.clk(gclk));
	jand g0178(.dina(n492),.dinb(w_n481_0[2]),.dout(n493),.clk(gclk));
	jand g0179(.dina(w_n493_0[1]),.dinb(w_n470_0[2]),.dout(n494),.clk(gclk));
	jnot g0180(.din(w_n494_0[1]),.dout(n495),.clk(gclk));
	jor g0181(.dina(w_dff_B_2GNWMdUI1_0),.dinb(w_n465_0[2]),.dout(n496),.clk(gclk));
	jnot g0182(.din(w_n469_1[0]),.dout(n497),.clk(gclk));
	jand g0183(.dina(n497),.dinb(w_G4415_1[0]),.dout(n498),.clk(gclk));
	jand g0184(.dina(w_n469_0[2]),.dinb(w_n466_0[0]),.dout(n499),.clk(gclk));
	jnot g0185(.din(n499),.dout(n500),.clk(gclk));
	jand g0186(.dina(w_n485_0[1]),.dinb(w_n482_0[0]),.dout(n501),.clk(gclk));
	jnot g0187(.din(n501),.dout(n502),.clk(gclk));
	jnot g0188(.din(w_n485_0[0]),.dout(n503),.clk(gclk));
	jand g0189(.dina(w_n503_0[1]),.dinb(w_G4410_1[0]),.dout(n504),.clk(gclk));
	jand g0190(.dina(w_n490_0[1]),.dinb(w_G4405_1[1]),.dout(n505),.clk(gclk));
	jnot g0191(.din(w_n475_1[0]),.dout(n506),.clk(gclk));
	jor g0192(.dina(w_n479_0[0]),.dinb(w_G4394_1[0]),.dout(n507),.clk(gclk));
	jor g0193(.dina(w_n507_1[2]),.dinb(n506),.dout(n508),.clk(gclk));
	jand g0194(.dina(w_n474_1[0]),.dinb(w_n471_0[1]),.dout(n509),.clk(gclk));
	jnot g0195(.din(w_n509_0[1]),.dout(n510),.clk(gclk));
	jor g0196(.dina(w_n490_0[0]),.dinb(w_G4405_1[0]),.dout(n511),.clk(gclk));
	jand g0197(.dina(n511),.dinb(w_n510_0[1]),.dout(n512),.clk(gclk));
	jand g0198(.dina(w_n512_0[1]),.dinb(w_n508_0[1]),.dout(n513),.clk(gclk));
	jor g0199(.dina(n513),.dinb(w_n505_0[1]),.dout(n514),.clk(gclk));
	jor g0200(.dina(w_n514_0[2]),.dinb(w_dff_B_RSpnqIE92_1),.dout(n515),.clk(gclk));
	jand g0201(.dina(n515),.dinb(w_n502_0[1]),.dout(n516),.clk(gclk));
	jand g0202(.dina(w_n516_0[2]),.dinb(w_dff_B_7bPW3G278_1),.dout(n517),.clk(gclk));
	jor g0203(.dina(n517),.dinb(w_dff_B_ReywKQIc6_1),.dout(n518),.clk(gclk));
	jand g0204(.dina(w_n518_0[1]),.dinb(n496),.dout(n519),.clk(gclk));
	jnot g0205(.din(w_G4427_0[1]),.dout(n520),.clk(gclk));
	jand g0206(.dina(G221),.dinb(w_G18_51[1]),.dout(n521),.clk(gclk));
	jand g0207(.dina(w_dff_B_AJSqunPQ4_0),.dinb(w_n355_23[0]),.dout(n522),.clk(gclk));
	jor g0208(.dina(w_n522_0[1]),.dinb(w_dff_B_fzUH6Gwg3_1),.dout(n523),.clk(gclk));
	jxor g0209(.dina(w_n523_0[2]),.dinb(w_n520_0[2]),.dout(n524),.clk(gclk));
	jnot g0210(.din(w_G4420_0[2]),.dout(n525),.clk(gclk));
	jand g0211(.dina(G222),.dinb(w_G18_51[0]),.dout(n526),.clk(gclk));
	jand g0212(.dina(w_dff_B_4FoRgvuD6_0),.dinb(w_n355_22[2]),.dout(n527),.clk(gclk));
	jor g0213(.dina(w_n527_0[1]),.dinb(w_dff_B_PcBIj1gP7_1),.dout(n528),.clk(gclk));
	jxor g0214(.dina(w_n528_1[1]),.dinb(w_n525_0[2]),.dout(n529),.clk(gclk));
	jand g0215(.dina(w_n529_0[1]),.dinb(w_n524_2[1]),.dout(n530),.clk(gclk));
	jnot g0216(.din(w_G4437_0[2]),.dout(n531),.clk(gclk));
	jand g0217(.dina(G219),.dinb(w_G18_50[2]),.dout(n532),.clk(gclk));
	jand g0218(.dina(w_dff_B_84iRtvq86_0),.dinb(w_n355_22[1]),.dout(n533),.clk(gclk));
	jor g0219(.dina(w_n533_0[1]),.dinb(w_dff_B_yAKEZt6k3_1),.dout(n534),.clk(gclk));
	jxor g0220(.dina(w_n534_1[1]),.dinb(w_n531_0[2]),.dout(n535),.clk(gclk));
	jnot g0221(.din(w_G4432_1[1]),.dout(n536),.clk(gclk));
	jand g0222(.dina(G220),.dinb(w_G18_50[1]),.dout(n537),.clk(gclk));
	jand g0223(.dina(w_dff_B_RbOHchf68_0),.dinb(w_n355_22[0]),.dout(n538),.clk(gclk));
	jor g0224(.dina(w_n538_0[1]),.dinb(w_dff_B_Uq25joIQ0_1),.dout(n539),.clk(gclk));
	jxor g0225(.dina(w_n539_1[1]),.dinb(w_n536_0[1]),.dout(n540),.clk(gclk));
	jand g0226(.dina(w_n540_0[2]),.dinb(w_n535_1[1]),.dout(n541),.clk(gclk));
	jand g0227(.dina(n541),.dinb(w_n530_0[1]),.dout(n542),.clk(gclk));
	jnot g0228(.din(w_n542_0[1]),.dout(n543),.clk(gclk));
	jor g0229(.dina(w_dff_B_Cd0jMb9i0_0),.dinb(w_n519_0[1]),.dout(n544),.clk(gclk));
	jnot g0230(.din(w_n534_1[0]),.dout(n545),.clk(gclk));
	jand g0231(.dina(n545),.dinb(w_G4437_0[1]),.dout(n546),.clk(gclk));
	jnot g0232(.din(n546),.dout(n547),.clk(gclk));
	jand g0233(.dina(w_n534_0[2]),.dinb(w_n531_0[1]),.dout(n548),.clk(gclk));
	jand g0234(.dina(w_n539_1[0]),.dinb(w_n536_0[0]),.dout(n549),.clk(gclk));
	jnot g0235(.din(w_n539_0[2]),.dout(n550),.clk(gclk));
	jand g0236(.dina(n550),.dinb(w_G4432_1[0]),.dout(n551),.clk(gclk));
	jnot g0237(.din(w_n551_0[1]),.dout(n552),.clk(gclk));
	jand g0238(.dina(w_n523_0[1]),.dinb(w_n520_0[1]),.dout(n553),.clk(gclk));
	jand g0239(.dina(w_n528_1[0]),.dinb(w_n525_0[1]),.dout(n554),.clk(gclk));
	jand g0240(.dina(w_n554_0[2]),.dinb(w_n524_2[0]),.dout(n555),.clk(gclk));
	jor g0241(.dina(n555),.dinb(w_n553_0[1]),.dout(n556),.clk(gclk));
	jand g0242(.dina(w_n556_0[2]),.dinb(w_n552_0[1]),.dout(n557),.clk(gclk));
	jor g0243(.dina(w_n557_0[1]),.dinb(w_n549_0[1]),.dout(n558),.clk(gclk));
	jor g0244(.dina(w_n558_0[2]),.dinb(w_dff_B_bU2JFqUT9_1),.dout(n559),.clk(gclk));
	jand g0245(.dina(n559),.dinb(w_dff_B_INxAodTD2_1),.dout(n560),.clk(gclk));
	jnot g0246(.din(w_n560_0[1]),.dout(n561),.clk(gclk));
	jand g0247(.dina(w_dff_B_eqNB2x3B1_0),.dinb(n544),.dout(n562),.clk(gclk));
	jnot g0248(.din(w_G2236_1[1]),.dout(n563),.clk(gclk));
	jand g0249(.dina(G12),.dinb(G9),.dout(n564),.clk(gclk));
	jnot g0250(.din(w_n564_0[2]),.dout(n565),.clk(gclk));
	jor g0251(.dina(w_dff_B_gkRoOqZ43_0),.dinb(w_n355_21[2]),.dout(n566),.clk(gclk));
	jand g0252(.dina(n566),.dinb(w_n565_10[1]),.dout(n567),.clk(gclk));
	jxor g0253(.dina(w_n567_1[1]),.dinb(w_n563_0[1]),.dout(n568),.clk(gclk));
	jnot g0254(.din(w_G2218_0[2]),.dout(n569),.clk(gclk));
	jand g0255(.dina(w_dff_B_3uEs4dVE0_0),.dinb(w_n355_21[1]),.dout(n570),.clk(gclk));
	jand g0256(.dina(G160),.dinb(w_G18_50[0]),.dout(n571),.clk(gclk));
	jor g0257(.dina(w_dff_B_KhfQAqlt3_0),.dinb(w_n570_0[1]),.dout(n572),.clk(gclk));
	jxor g0258(.dina(w_n572_1[1]),.dinb(w_n569_0[2]),.dout(n573),.clk(gclk));
	jnot g0259(.din(w_G2211_0[2]),.dout(n574),.clk(gclk));
	jand g0260(.dina(w_dff_B_rnocEosP8_0),.dinb(w_n355_21[0]),.dout(n575),.clk(gclk));
	jand g0261(.dina(G151),.dinb(w_G18_49[2]),.dout(n576),.clk(gclk));
	jor g0262(.dina(w_dff_B_3C2QXZfv3_0),.dinb(w_n575_0[1]),.dout(n577),.clk(gclk));
	jxor g0263(.dina(w_n577_0[2]),.dinb(w_n574_0[1]),.dout(n578),.clk(gclk));
	jand g0264(.dina(w_n578_1[1]),.dinb(w_n573_1[1]),.dout(n579),.clk(gclk));
	jnot g0265(.din(w_G2230_1[1]),.dout(n580),.clk(gclk));
	jand g0266(.dina(w_dff_B_1N5R0yCL3_0),.dinb(w_n355_20[2]),.dout(n581),.clk(gclk));
	jand g0267(.dina(G158),.dinb(w_G18_49[1]),.dout(n582),.clk(gclk));
	jor g0268(.dina(w_dff_B_D5js8nOw4_0),.dinb(w_n581_0[1]),.dout(n583),.clk(gclk));
	jxor g0269(.dina(w_n583_1[1]),.dinb(w_n580_0[1]),.dout(n584),.clk(gclk));
	jnot g0270(.din(w_G2224_1[1]),.dout(n585),.clk(gclk));
	jand g0271(.dina(w_dff_B_lV3ChrZN8_0),.dinb(w_n355_20[1]),.dout(n586),.clk(gclk));
	jand g0272(.dina(G159),.dinb(w_G18_49[0]),.dout(n587),.clk(gclk));
	jor g0273(.dina(w_dff_B_DeBhIout9_0),.dinb(w_n586_0[1]),.dout(n588),.clk(gclk));
	jxor g0274(.dina(w_n588_1[1]),.dinb(w_n585_0[1]),.dout(n589),.clk(gclk));
	jand g0275(.dina(w_n589_1[1]),.dinb(w_n584_0[2]),.dout(n590),.clk(gclk));
	jand g0276(.dina(n590),.dinb(w_n579_0[2]),.dout(n591),.clk(gclk));
	jand g0277(.dina(w_n591_0[1]),.dinb(w_n568_0[2]),.dout(n592),.clk(gclk));
	jnot g0278(.din(w_n592_0[1]),.dout(n593),.clk(gclk));
	jor g0279(.dina(w_dff_B_fuApnOfa2_0),.dinb(w_n562_0[2]),.dout(n594),.clk(gclk));
	jand g0280(.dina(w_n567_1[0]),.dinb(w_n563_0[0]),.dout(n595),.clk(gclk));
	jnot g0281(.din(n595),.dout(n596),.clk(gclk));
	jnot g0282(.din(w_n567_0[2]),.dout(n597),.clk(gclk));
	jand g0283(.dina(n597),.dinb(w_G2236_1[0]),.dout(n598),.clk(gclk));
	jand g0284(.dina(w_n583_1[0]),.dinb(w_n580_0[0]),.dout(n599),.clk(gclk));
	jnot g0285(.din(w_n599_0[1]),.dout(n600),.clk(gclk));
	jnot g0286(.din(w_n583_0[2]),.dout(n601),.clk(gclk));
	jand g0287(.dina(n601),.dinb(w_G2230_1[0]),.dout(n602),.clk(gclk));
	jnot g0288(.din(w_n588_1[0]),.dout(n603),.clk(gclk));
	jand g0289(.dina(n603),.dinb(w_G2224_1[0]),.dout(n604),.clk(gclk));
	jnot g0290(.din(n604),.dout(n605),.clk(gclk));
	jand g0291(.dina(w_n577_0[1]),.dinb(w_n574_0[0]),.dout(n606),.clk(gclk));
	jand g0292(.dina(w_n606_1[2]),.dinb(w_n573_1[0]),.dout(n607),.clk(gclk));
	jand g0293(.dina(w_n572_1[0]),.dinb(w_n569_0[1]),.dout(n608),.clk(gclk));
	jand g0294(.dina(w_n588_0[2]),.dinb(w_n585_0[0]),.dout(n609),.clk(gclk));
	jor g0295(.dina(n609),.dinb(w_n608_0[2]),.dout(n610),.clk(gclk));
	jor g0296(.dina(w_n610_0[1]),.dinb(w_n607_0[1]),.dout(n611),.clk(gclk));
	jand g0297(.dina(n611),.dinb(w_n605_0[1]),.dout(n612),.clk(gclk));
	jnot g0298(.din(w_n612_0[1]),.dout(n613),.clk(gclk));
	jor g0299(.dina(w_n613_0[2]),.dinb(w_dff_B_PSNRXKgT4_1),.dout(n614),.clk(gclk));
	jand g0300(.dina(n614),.dinb(w_dff_B_bO2tCcQc4_1),.dout(n615),.clk(gclk));
	jor g0301(.dina(w_n615_1[1]),.dinb(w_dff_B_IFTfh1mX6_1),.dout(n616),.clk(gclk));
	jand g0302(.dina(n616),.dinb(w_dff_B_9fDOTzUJ0_1),.dout(n617),.clk(gclk));
	jand g0303(.dina(w_n617_0[1]),.dinb(n594),.dout(n618),.clk(gclk));
	jnot g0304(.din(w_G2247_0[2]),.dout(n619),.clk(gclk));
	jor g0305(.dina(w_dff_B_ushaR9vI3_0),.dinb(w_n355_20[0]),.dout(n620),.clk(gclk));
	jand g0306(.dina(w_n620_0[1]),.dinb(w_n565_10[0]),.dout(n621),.clk(gclk));
	jxor g0307(.dina(w_n621_0[2]),.dinb(w_n619_0[1]),.dout(n622),.clk(gclk));
	jnot g0308(.din(w_G2239_0[2]),.dout(n623),.clk(gclk));
	jor g0309(.dina(w_dff_B_q90zLv3b6_0),.dinb(w_n355_19[2]),.dout(n624),.clk(gclk));
	jand g0310(.dina(w_n624_0[1]),.dinb(w_n565_9[2]),.dout(n625),.clk(gclk));
	jxor g0311(.dina(w_n625_0[2]),.dinb(w_n623_0[2]),.dout(n626),.clk(gclk));
	jand g0312(.dina(w_n626_0[1]),.dinb(w_n622_1[1]),.dout(n627),.clk(gclk));
	jnot g0313(.din(w_G2256_1[1]),.dout(n628),.clk(gclk));
	jor g0314(.dina(w_dff_B_9U7qMuqH0_0),.dinb(w_n355_19[1]),.dout(n629),.clk(gclk));
	jand g0315(.dina(w_n629_0[1]),.dinb(w_n565_9[1]),.dout(n630),.clk(gclk));
	jxor g0316(.dina(w_n630_0[2]),.dinb(w_n628_0[1]),.dout(n631),.clk(gclk));
	jnot g0317(.din(w_G2253_1[1]),.dout(n632),.clk(gclk));
	jor g0318(.dina(w_dff_B_gmR2tVV00_0),.dinb(w_n355_19[0]),.dout(n633),.clk(gclk));
	jand g0319(.dina(w_n633_0[1]),.dinb(w_n565_9[0]),.dout(n634),.clk(gclk));
	jxor g0320(.dina(w_n634_0[2]),.dinb(w_n632_0[1]),.dout(n635),.clk(gclk));
	jand g0321(.dina(w_n635_0[2]),.dinb(w_n631_0[1]),.dout(n636),.clk(gclk));
	jand g0322(.dina(n636),.dinb(w_n627_0[1]),.dout(n637),.clk(gclk));
	jnot g0323(.din(w_n637_0[1]),.dout(n638),.clk(gclk));
	jor g0324(.dina(w_dff_B_5bVHzCoB6_0),.dinb(w_n618_0[2]),.dout(n639),.clk(gclk));
	jand g0325(.dina(w_n630_0[1]),.dinb(w_n628_0[0]),.dout(n640),.clk(gclk));
	jnot g0326(.din(n640),.dout(n641),.clk(gclk));
	jand g0327(.dina(w_n634_0[1]),.dinb(w_n632_0[0]),.dout(n642),.clk(gclk));
	jnot g0328(.din(w_n642_0[1]),.dout(n643),.clk(gclk));
	jand g0329(.dina(w_n621_0[1]),.dinb(w_n619_0[0]),.dout(n644),.clk(gclk));
	jand g0330(.dina(w_n625_0[1]),.dinb(w_n623_0[1]),.dout(n645),.clk(gclk));
	jand g0331(.dina(w_n645_0[2]),.dinb(w_n622_1[0]),.dout(n646),.clk(gclk));
	jor g0332(.dina(n646),.dinb(w_dff_B_C4tzDZ6m2_1),.dout(n647),.clk(gclk));
	jnot g0333(.din(w_n647_0[1]),.dout(n648),.clk(gclk));
	jand g0334(.dina(w_n648_0[2]),.dinb(w_n643_0[1]),.dout(n649),.clk(gclk));
	jnot g0335(.din(w_n630_0[0]),.dout(n650),.clk(gclk));
	jand g0336(.dina(w_n650_0[1]),.dinb(w_G2256_1[0]),.dout(n651),.clk(gclk));
	jnot g0337(.din(w_n634_0[0]),.dout(n652),.clk(gclk));
	jand g0338(.dina(w_n652_0[1]),.dinb(w_G2253_1[0]),.dout(n653),.clk(gclk));
	jor g0339(.dina(w_n653_1[1]),.dinb(n651),.dout(n654),.clk(gclk));
	jor g0340(.dina(w_dff_B_QRx72X1R3_0),.dinb(w_n649_0[1]),.dout(n655),.clk(gclk));
	jand g0341(.dina(n655),.dinb(w_dff_B_M9KreNBI5_1),.dout(n656),.clk(gclk));
	jand g0342(.dina(w_n656_0[1]),.dinb(n639),.dout(n657),.clk(gclk));
	jnot g0343(.din(w_G1486_0[2]),.dout(n658),.clk(gclk));
	jor g0344(.dina(w_dff_B_tR2LbQ4n4_0),.dinb(w_n355_18[2]),.dout(n659),.clk(gclk));
	jand g0345(.dina(w_n659_0[1]),.dinb(w_n565_8[2]),.dout(n660),.clk(gclk));
	jxor g0346(.dina(w_n660_1[1]),.dinb(w_n658_0[2]),.dout(n661),.clk(gclk));
	jnot g0347(.din(w_G1480_0[2]),.dout(n662),.clk(gclk));
	jor g0348(.dina(w_dff_B_n7oZ3W448_0),.dinb(w_n355_18[1]),.dout(n663),.clk(gclk));
	jand g0349(.dina(w_n663_0[1]),.dinb(w_n565_8[1]),.dout(n664),.clk(gclk));
	jxor g0350(.dina(w_n664_1[1]),.dinb(w_n662_0[2]),.dout(n665),.clk(gclk));
	jnot g0351(.din(w_G106_1[1]),.dout(n666),.clk(gclk));
	jor g0352(.dina(w_dff_B_XHcYUwEC3_0),.dinb(w_n355_18[0]),.dout(n667),.clk(gclk));
	jand g0353(.dina(w_n667_0[1]),.dinb(w_n565_8[0]),.dout(n668),.clk(gclk));
	jxor g0354(.dina(w_n668_0[2]),.dinb(w_n666_0[1]),.dout(n669),.clk(gclk));
	jand g0355(.dina(w_n669_0[2]),.dinb(w_n665_0[2]),.dout(n670),.clk(gclk));
	jnot g0356(.din(w_G1469_1[1]),.dout(n671),.clk(gclk));
	jor g0357(.dina(w_dff_B_k0FUDk4O7_0),.dinb(w_n355_17[2]),.dout(n672),.clk(gclk));
	jand g0358(.dina(w_n672_0[1]),.dinb(w_n565_7[2]),.dout(n673),.clk(gclk));
	jxor g0359(.dina(w_n673_0[2]),.dinb(w_n671_0[1]),.dout(n674),.clk(gclk));
	jnot g0360(.din(w_G1462_0[2]),.dout(n675),.clk(gclk));
	jor g0361(.dina(w_dff_B_ntO3dZxz6_0),.dinb(w_n355_17[1]),.dout(n676),.clk(gclk));
	jand g0362(.dina(w_n676_0[1]),.dinb(w_n565_7[1]),.dout(n677),.clk(gclk));
	jxor g0363(.dina(w_n677_0[2]),.dinb(w_n675_0[2]),.dout(n678),.clk(gclk));
	jand g0364(.dina(w_n678_0[2]),.dinb(w_n674_1[1]),.dout(n679),.clk(gclk));
	jand g0365(.dina(w_n679_1[1]),.dinb(n670),.dout(n680),.clk(gclk));
	jand g0366(.dina(w_n680_0[1]),.dinb(w_n661_0[1]),.dout(n681),.clk(gclk));
	jnot g0367(.din(n681),.dout(n682),.clk(gclk));
	jor g0368(.dina(w_dff_B_v6k1PaaS2_0),.dinb(w_n657_1[1]),.dout(n683),.clk(gclk));
	jand g0369(.dina(w_n660_1[0]),.dinb(w_n658_0[1]),.dout(n684),.clk(gclk));
	jor g0370(.dina(w_n660_0[2]),.dinb(w_n658_0[0]),.dout(n685),.clk(gclk));
	jand g0371(.dina(w_n664_1[0]),.dinb(w_n662_0[1]),.dout(n686),.clk(gclk));
	jnot g0372(.din(w_n686_0[1]),.dout(n687),.clk(gclk));
	jor g0373(.dina(w_n664_0[2]),.dinb(w_n662_0[0]),.dout(n688),.clk(gclk));
	jand g0374(.dina(w_n668_0[1]),.dinb(w_n666_0[0]),.dout(n689),.clk(gclk));
	jnot g0375(.din(w_n668_0[0]),.dout(n690),.clk(gclk));
	jand g0376(.dina(w_n690_0[1]),.dinb(w_G106_1[0]),.dout(n691),.clk(gclk));
	jnot g0377(.din(n691),.dout(n692),.clk(gclk));
	jnot g0378(.din(w_n673_0[1]),.dout(n693),.clk(gclk));
	jand g0379(.dina(w_n693_0[1]),.dinb(w_G1469_1[0]),.dout(n694),.clk(gclk));
	jnot g0380(.din(n694),.dout(n695),.clk(gclk));
	jand g0381(.dina(w_n673_0[0]),.dinb(w_n671_0[0]),.dout(n696),.clk(gclk));
	jand g0382(.dina(w_n677_0[1]),.dinb(w_n675_0[1]),.dout(n697),.clk(gclk));
	jor g0383(.dina(w_n697_0[2]),.dinb(n696),.dout(n698),.clk(gclk));
	jand g0384(.dina(w_dff_B_ZrU08K1A0_0),.dinb(n695),.dout(n699),.clk(gclk));
	jand g0385(.dina(w_n699_1[1]),.dinb(w_n692_0[1]),.dout(n700),.clk(gclk));
	jor g0386(.dina(n700),.dinb(w_dff_B_fuS5g3We1_1),.dout(n701),.clk(gclk));
	jand g0387(.dina(w_n701_1[1]),.dinb(w_dff_B_eirtcAzx3_1),.dout(n702),.clk(gclk));
	jnot g0388(.din(n702),.dout(n703),.clk(gclk));
	jand g0389(.dina(w_n703_0[1]),.dinb(w_n687_0[1]),.dout(n704),.clk(gclk));
	jnot g0390(.din(w_n704_0[1]),.dout(n705),.clk(gclk));
	jand g0391(.dina(w_n705_0[1]),.dinb(w_dff_B_R8R1GegZ9_1),.dout(n706),.clk(gclk));
	jor g0392(.dina(n706),.dinb(w_dff_B_dBcfTNrF6_1),.dout(n707),.clk(gclk));
	jnot g0393(.din(w_n707_0[2]),.dout(n708),.clk(gclk));
	jand g0394(.dina(w_n708_0[1]),.dinb(w_n683_0[1]),.dout(n709),.clk(gclk));
	jnot g0395(.din(w_G38_1[1]),.dout(n710),.clk(gclk));
	jand g0396(.dina(w_G4528_0[1]),.dinb(w_G1492_1[1]),.dout(n711),.clk(gclk));
	jxor g0397(.dina(w_n711_0[1]),.dinb(w_n710_0[1]),.dout(n712),.clk(gclk));
	jnot g0398(.din(w_n712_0[1]),.dout(n713),.clk(gclk));
	jor g0399(.dina(w_n713_1[1]),.dinb(w_n709_1[1]),.dout(n714),.clk(gclk));
	jor g0400(.dina(w_n714_0[1]),.dinb(w_n365_0[1]),.dout(n715),.clk(gclk));
	jnot g0401(.din(w_n715_0[2]),.dout(n716),.clk(gclk));
	jnot g0402(.din(w_G1492_1[0]),.dout(n717),.clk(gclk));
	jnot g0403(.din(w_n364_0[0]),.dout(n718),.clk(gclk));
	jor g0404(.dina(n718),.dinb(w_dff_B_2oZZjT7X1_1),.dout(n719),.clk(gclk));
	jand g0405(.dina(n719),.dinb(w_G38_1[0]),.dout(n720),.clk(gclk));
	jor g0406(.dina(w_n720_1[1]),.dinb(w_n716_1[1]),.dout(w_dff_A_R2YdaLCt7_2),.clk(gclk));
	jor g0407(.dina(w_dff_B_xFKgSs601_0),.dinb(w_n355_17[0]),.dout(n722),.clk(gclk));
	jand g0408(.dina(n722),.dinb(w_n565_7[0]),.dout(n723),.clk(gclk));
	jand g0409(.dina(w_G2236_0[2]),.dinb(w_G18_48[2]),.dout(n724),.clk(gclk));
	jnot g0410(.din(n724),.dout(n725),.clk(gclk));
	jor g0411(.dina(G64),.dinb(w_G18_48[1]),.dout(n726),.clk(gclk));
	jand g0412(.dina(w_dff_B_Ys5oJSE10_0),.dinb(n725),.dout(n727),.clk(gclk));
	jor g0413(.dina(w_n727_0[2]),.dinb(w_n723_0[2]),.dout(n728),.clk(gclk));
	jand g0414(.dina(G178),.dinb(w_G18_48[0]),.dout(n729),.clk(gclk));
	jor g0415(.dina(w_dff_B_2pGwruPz1_0),.dinb(w_n581_0[0]),.dout(n730),.clk(gclk));
	jand g0416(.dina(w_G2230_0[2]),.dinb(w_G18_47[2]),.dout(n731),.clk(gclk));
	jnot g0417(.din(n731),.dout(n732),.clk(gclk));
	jor g0418(.dina(G85),.dinb(w_G18_47[1]),.dout(n733),.clk(gclk));
	jand g0419(.dina(w_dff_B_U1958RBQ3_0),.dinb(n732),.dout(n734),.clk(gclk));
	jor g0420(.dina(w_n734_0[2]),.dinb(w_n730_0[2]),.dout(n735),.clk(gclk));
	jand g0421(.dina(G179),.dinb(w_G18_47[0]),.dout(n736),.clk(gclk));
	jor g0422(.dina(w_dff_B_uYOex2N95_0),.dinb(w_n586_0[0]),.dout(n737),.clk(gclk));
	jand g0423(.dina(w_G2224_0[2]),.dinb(w_G18_46[2]),.dout(n738),.clk(gclk));
	jnot g0424(.din(n738),.dout(n739),.clk(gclk));
	jor g0425(.dina(G84),.dinb(w_G18_46[1]),.dout(n740),.clk(gclk));
	jand g0426(.dina(w_dff_B_Lcgy86XL0_0),.dinb(n739),.dout(n741),.clk(gclk));
	jand g0427(.dina(w_n741_0[2]),.dinb(w_n737_0[2]),.dout(n742),.clk(gclk));
	jand g0428(.dina(G180),.dinb(w_G18_46[0]),.dout(n743),.clk(gclk));
	jor g0429(.dina(w_dff_B_mds2AIK08_0),.dinb(w_n570_0[0]),.dout(n744),.clk(gclk));
	jand g0430(.dina(w_G2218_0[1]),.dinb(w_G18_45[2]),.dout(n745),.clk(gclk));
	jnot g0431(.din(n745),.dout(n746),.clk(gclk));
	jor g0432(.dina(G83),.dinb(w_G18_45[1]),.dout(n747),.clk(gclk));
	jand g0433(.dina(w_dff_B_m2voZ3vE6_0),.dinb(n746),.dout(n748),.clk(gclk));
	jor g0434(.dina(w_n748_0[2]),.dinb(w_n744_0[2]),.dout(n749),.clk(gclk));
	jor g0435(.dina(w_n741_0[1]),.dinb(w_n737_0[1]),.dout(n750),.clk(gclk));
	jand g0436(.dina(n750),.dinb(n749),.dout(n751),.clk(gclk));
	jand g0437(.dina(w_n748_0[1]),.dinb(w_n744_0[1]),.dout(n752),.clk(gclk));
	jand g0438(.dina(G171),.dinb(w_G18_45[0]),.dout(n753),.clk(gclk));
	jor g0439(.dina(w_dff_B_jMZecd1B1_0),.dinb(w_n575_0[0]),.dout(n754),.clk(gclk));
	jand g0440(.dina(w_G2211_0[1]),.dinb(w_G18_44[2]),.dout(n755),.clk(gclk));
	jnot g0441(.din(n755),.dout(n756),.clk(gclk));
	jor g0442(.dina(G65),.dinb(w_G18_44[1]),.dout(n757),.clk(gclk));
	jand g0443(.dina(w_dff_B_ZvV1HQX72_0),.dinb(n756),.dout(n758),.clk(gclk));
	jand g0444(.dina(w_n758_0[2]),.dinb(w_n754_0[2]),.dout(n759),.clk(gclk));
	jor g0445(.dina(w_n759_0[1]),.dinb(w_n752_0[1]),.dout(n760),.clk(gclk));
	jand g0446(.dina(n760),.dinb(w_n751_0[1]),.dout(n761),.clk(gclk));
	jor g0447(.dina(n761),.dinb(w_n742_0[1]),.dout(n762),.clk(gclk));
	jand g0448(.dina(n762),.dinb(w_n735_0[1]),.dout(n763),.clk(gclk));
	jand g0449(.dina(w_n734_0[1]),.dinb(w_n730_0[1]),.dout(n764),.clk(gclk));
	jand g0450(.dina(w_n727_0[1]),.dinb(w_n723_0[1]),.dout(n765),.clk(gclk));
	jor g0451(.dina(w_n765_0[1]),.dinb(w_n764_0[1]),.dout(n766),.clk(gclk));
	jor g0452(.dina(w_dff_B_iEn66Zu24_0),.dinb(n763),.dout(n767),.clk(gclk));
	jand g0453(.dina(n767),.dinb(w_n728_0[1]),.dout(n768),.clk(gclk));
	jnot g0454(.din(w_n752_0[0]),.dout(n769),.clk(gclk));
	jand g0455(.dina(n769),.dinb(w_n735_0[0]),.dout(n770),.clk(gclk));
	jnot g0456(.din(w_n742_0[0]),.dout(n771),.clk(gclk));
	jnot g0457(.din(w_n759_0[0]),.dout(n772),.clk(gclk));
	jand g0458(.dina(n772),.dinb(n771),.dout(n773),.clk(gclk));
	jand g0459(.dina(n773),.dinb(n770),.dout(n774),.clk(gclk));
	jnot g0460(.din(w_n765_0[0]),.dout(n775),.clk(gclk));
	jor g0461(.dina(w_n758_0[1]),.dinb(w_n754_0[1]),.dout(n776),.clk(gclk));
	jand g0462(.dina(w_dff_B_UQ2eWhvW8_0),.dinb(n775),.dout(n777),.clk(gclk));
	jnot g0463(.din(w_n764_0[0]),.dout(n778),.clk(gclk));
	jand g0464(.dina(n778),.dinb(w_n728_0[0]),.dout(n779),.clk(gclk));
	jand g0465(.dina(n779),.dinb(n777),.dout(n780),.clk(gclk));
	jand g0466(.dina(n780),.dinb(w_n751_0[0]),.dout(n781),.clk(gclk));
	jand g0467(.dina(n781),.dinb(w_dff_B_NjHQMahz2_1),.dout(n782),.clk(gclk));
	jand g0468(.dina(G191),.dinb(w_G18_44[0]),.dout(n783),.clk(gclk));
	jor g0469(.dina(w_dff_B_UYt0YtB46_0),.dinb(w_n522_0[0]),.dout(n784),.clk(gclk));
	jor g0470(.dina(G60),.dinb(w_G18_43[2]),.dout(n785),.clk(gclk));
	jor g0471(.dina(w_n520_0[0]),.dinb(w_n355_16[2]),.dout(n786),.clk(gclk));
	jand g0472(.dina(n786),.dinb(w_dff_B_B0owYQxb4_1),.dout(n787),.clk(gclk));
	jxor g0473(.dina(w_n787_0[2]),.dinb(w_n784_0[2]),.dout(n788),.clk(gclk));
	jand g0474(.dina(G189),.dinb(w_G18_43[1]),.dout(n789),.clk(gclk));
	jor g0475(.dina(w_dff_B_BdF6J7Nd9_0),.dinb(w_n533_0[0]),.dout(n790),.clk(gclk));
	jor g0476(.dina(G62),.dinb(w_G18_43[0]),.dout(n791),.clk(gclk));
	jor g0477(.dina(w_n531_0[0]),.dinb(w_n355_16[1]),.dout(n792),.clk(gclk));
	jand g0478(.dina(n792),.dinb(w_dff_B_XUlCmyH13_1),.dout(n793),.clk(gclk));
	jxor g0479(.dina(w_n793_1[1]),.dinb(w_n790_1[1]),.dout(n794),.clk(gclk));
	jand g0480(.dina(n794),.dinb(n788),.dout(n795),.clk(gclk));
	jand g0481(.dina(G190),.dinb(w_G18_42[2]),.dout(n796),.clk(gclk));
	jor g0482(.dina(w_dff_B_yCOS2wms3_0),.dinb(w_n538_0[0]),.dout(n797),.clk(gclk));
	jor g0483(.dina(G61),.dinb(w_G18_42[1]),.dout(n798),.clk(gclk));
	jand g0484(.dina(w_G4432_0[2]),.dinb(w_G18_42[0]),.dout(n799),.clk(gclk));
	jnot g0485(.din(n799),.dout(n800),.clk(gclk));
	jand g0486(.dina(n800),.dinb(w_dff_B_sNtu3yve4_1),.dout(n801),.clk(gclk));
	jxor g0487(.dina(w_n801_1[1]),.dinb(w_n797_1[1]),.dout(n802),.clk(gclk));
	jand g0488(.dina(G192),.dinb(w_G18_41[2]),.dout(n803),.clk(gclk));
	jor g0489(.dina(w_dff_B_y2mL8afH4_0),.dinb(w_n527_0[0]),.dout(n804),.clk(gclk));
	jor g0490(.dina(G79),.dinb(w_G18_41[1]),.dout(n805),.clk(gclk));
	jor g0491(.dina(w_n525_0[0]),.dinb(w_n355_16[0]),.dout(n806),.clk(gclk));
	jand g0492(.dina(n806),.dinb(w_dff_B_aDgzSQ3W6_1),.dout(n807),.clk(gclk));
	jxor g0493(.dina(w_n807_0[2]),.dinb(w_n804_0[2]),.dout(n808),.clk(gclk));
	jand g0494(.dina(n808),.dinb(w_n802_0[1]),.dout(n809),.clk(gclk));
	jand g0495(.dina(n809),.dinb(w_n795_0[1]),.dout(n810),.clk(gclk));
	jand g0496(.dina(G196),.dinb(w_G18_41[0]),.dout(n811),.clk(gclk));
	jor g0497(.dina(w_dff_B_Cq4SEy4M3_0),.dinb(w_n473_0[0]),.dout(n812),.clk(gclk));
	jor g0498(.dina(G78),.dinb(w_G18_40[2]),.dout(n813),.clk(gclk));
	jand g0499(.dina(w_G4400_0[1]),.dinb(w_G18_40[1]),.dout(n814),.clk(gclk));
	jnot g0500(.din(n814),.dout(n815),.clk(gclk));
	jand g0501(.dina(n815),.dinb(w_dff_B_WDAEk5L34_1),.dout(n816),.clk(gclk));
	jor g0502(.dina(w_n816_0[2]),.dinb(w_n812_0[2]),.dout(n817),.clk(gclk));
	jand g0503(.dina(G195),.dinb(w_G18_40[0]),.dout(n818),.clk(gclk));
	jor g0504(.dina(w_dff_B_pEGy5yFX6_0),.dinb(w_n488_0[0]),.dout(n819),.clk(gclk));
	jor g0505(.dina(G59),.dinb(w_G18_39[2]),.dout(n820),.clk(gclk));
	jand g0506(.dina(w_G4405_0[2]),.dinb(w_G18_39[1]),.dout(n821),.clk(gclk));
	jnot g0507(.din(n821),.dout(n822),.clk(gclk));
	jand g0508(.dina(n822),.dinb(w_dff_B_P2O9N3ze6_1),.dout(n823),.clk(gclk));
	jor g0509(.dina(w_n823_0[2]),.dinb(w_n819_0[2]),.dout(n824),.clk(gclk));
	jand g0510(.dina(w_n824_0[1]),.dinb(w_n817_0[1]),.dout(n825),.clk(gclk));
	jand g0511(.dina(G187),.dinb(w_G18_39[0]),.dout(n826),.clk(gclk));
	jor g0512(.dina(w_dff_B_VWQRY0eh8_0),.dinb(w_n477_0[0]),.dout(n827),.clk(gclk));
	jor g0513(.dina(G77),.dinb(w_G18_38[2]),.dout(n828),.clk(gclk));
	jand g0514(.dina(w_G4394_0[2]),.dinb(w_G18_38[1]),.dout(n829),.clk(gclk));
	jnot g0515(.din(n829),.dout(n830),.clk(gclk));
	jand g0516(.dina(n830),.dinb(w_dff_B_DAJuA5HC0_1),.dout(n831),.clk(gclk));
	jand g0517(.dina(w_n831_0[2]),.dinb(w_n827_0[2]),.dout(n832),.clk(gclk));
	jnot g0518(.din(w_n832_0[1]),.dout(n833),.clk(gclk));
	jand g0519(.dina(w_n823_0[1]),.dinb(w_n819_0[1]),.dout(n834),.clk(gclk));
	jnot g0520(.din(w_n834_0[1]),.dout(n835),.clk(gclk));
	jand g0521(.dina(n835),.dinb(n833),.dout(n836),.clk(gclk));
	jand g0522(.dina(n836),.dinb(w_dff_B_hc7iIvA21_1),.dout(n837),.clk(gclk));
	jand g0523(.dina(w_n816_0[1]),.dinb(w_n812_0[1]),.dout(n838),.clk(gclk));
	jnot g0524(.din(w_n838_0[1]),.dout(n839),.clk(gclk));
	jor g0525(.dina(w_n831_0[1]),.dinb(w_n827_0[1]),.dout(n840),.clk(gclk));
	jand g0526(.dina(w_dff_B_eyGmmzk53_0),.dinb(n839),.dout(n841),.clk(gclk));
	jand g0527(.dina(G193),.dinb(w_G18_38[0]),.dout(n842),.clk(gclk));
	jor g0528(.dina(w_dff_B_FVEpOpmI2_0),.dinb(w_n468_0[0]),.dout(n843),.clk(gclk));
	jor g0529(.dina(G80),.dinb(w_G18_37[2]),.dout(n844),.clk(gclk));
	jand g0530(.dina(w_G4415_0[2]),.dinb(w_G18_37[1]),.dout(n845),.clk(gclk));
	jnot g0531(.din(n845),.dout(n846),.clk(gclk));
	jand g0532(.dina(n846),.dinb(w_dff_B_F9BIbIMB5_1),.dout(n847),.clk(gclk));
	jand g0533(.dina(w_n847_0[2]),.dinb(w_n843_0[2]),.dout(n848),.clk(gclk));
	jnot g0534(.din(w_n848_0[1]),.dout(n849),.clk(gclk));
	jand g0535(.dina(G194),.dinb(w_G18_37[0]),.dout(n850),.clk(gclk));
	jor g0536(.dina(w_dff_B_h00Pwn007_0),.dinb(w_n484_0[0]),.dout(n851),.clk(gclk));
	jor g0537(.dina(G81),.dinb(w_G18_36[2]),.dout(n852),.clk(gclk));
	jand g0538(.dina(w_G4410_0[2]),.dinb(w_G18_36[1]),.dout(n853),.clk(gclk));
	jnot g0539(.din(n853),.dout(n854),.clk(gclk));
	jand g0540(.dina(n854),.dinb(w_dff_B_02keszY75_1),.dout(n855),.clk(gclk));
	jor g0541(.dina(w_n855_0[2]),.dinb(w_n851_0[2]),.dout(n856),.clk(gclk));
	jand g0542(.dina(w_n856_0[1]),.dinb(n849),.dout(n857),.clk(gclk));
	jor g0543(.dina(w_n847_0[1]),.dinb(w_n843_0[1]),.dout(n858),.clk(gclk));
	jand g0544(.dina(w_n855_0[1]),.dinb(w_n851_0[1]),.dout(n859),.clk(gclk));
	jnot g0545(.din(w_n859_0[1]),.dout(n860),.clk(gclk));
	jand g0546(.dina(n860),.dinb(w_n858_0[2]),.dout(n861),.clk(gclk));
	jand g0547(.dina(n861),.dinb(n857),.dout(n862),.clk(gclk));
	jand g0548(.dina(n862),.dinb(w_dff_B_BB9j9eEC6_1),.dout(n863),.clk(gclk));
	jand g0549(.dina(n863),.dinb(w_dff_B_olKMC4kn6_1),.dout(n864),.clk(gclk));
	jand g0550(.dina(w_n864_0[1]),.dinb(w_n810_0[2]),.dout(n865),.clk(gclk));
	jand g0551(.dina(G200),.dinb(w_G18_36[0]),.dout(n866),.clk(gclk));
	jnot g0552(.din(n866),.dout(n867),.clk(gclk));
	jand g0553(.dina(n867),.dinb(w_n441_0[0]),.dout(n868),.clk(gclk));
	jnot g0554(.din(n868),.dout(n869),.clk(gclk));
	jor g0555(.dina(G56),.dinb(w_G18_35[2]),.dout(n870),.clk(gclk));
	jand g0556(.dina(w_G3749_0[2]),.dinb(w_G18_35[1]),.dout(n871),.clk(gclk));
	jnot g0557(.din(n871),.dout(n872),.clk(gclk));
	jand g0558(.dina(n872),.dinb(w_dff_B_JfloGEvr0_1),.dout(n873),.clk(gclk));
	jand g0559(.dina(w_n873_0[2]),.dinb(w_n869_0[2]),.dout(n874),.clk(gclk));
	jnot g0560(.din(w_n874_0[1]),.dout(n875),.clk(gclk));
	jnot g0561(.din(w_n427_0[0]),.dout(n876),.clk(gclk));
	jand g0562(.dina(G202),.dinb(w_G18_35[0]),.dout(n877),.clk(gclk));
	jor g0563(.dina(w_dff_B_GHMBKMEz3_0),.dinb(n876),.dout(n878),.clk(gclk));
	jor g0564(.dina(G54),.dinb(w_G18_34[2]),.dout(n879),.clk(gclk));
	jand g0565(.dina(w_G3737_0[2]),.dinb(w_G18_34[1]),.dout(n880),.clk(gclk));
	jnot g0566(.din(n880),.dout(n881),.clk(gclk));
	jand g0567(.dina(n881),.dinb(w_dff_B_PUf4qp3b3_1),.dout(n882),.clk(gclk));
	jor g0568(.dina(w_n882_0[2]),.dinb(w_n878_0[2]),.dout(n883),.clk(gclk));
	jand g0569(.dina(w_dff_B_oyvPw3HP8_0),.dinb(n875),.dout(n884),.clk(gclk));
	jand g0570(.dina(w_n882_0[1]),.dinb(w_n878_0[1]),.dout(n885),.clk(gclk));
	jnot g0571(.din(w_n885_0[1]),.dout(n886),.clk(gclk));
	jor g0572(.dina(w_n873_0[1]),.dinb(w_n869_0[1]),.dout(n887),.clk(gclk));
	jand g0573(.dina(w_n887_0[1]),.dinb(n886),.dout(n888),.clk(gclk));
	jand g0574(.dina(n888),.dinb(n884),.dout(n889),.clk(gclk));
	jand g0575(.dina(G201),.dinb(w_G18_34[0]),.dout(n890),.clk(gclk));
	jor g0576(.dina(w_dff_B_8XEg0JBA1_0),.dinb(w_n448_0[0]),.dout(n891),.clk(gclk));
	jor g0577(.dina(G55),.dinb(w_G18_33[2]),.dout(n892),.clk(gclk));
	jand g0578(.dina(w_G3743_0[2]),.dinb(w_G18_33[1]),.dout(n893),.clk(gclk));
	jnot g0579(.din(n893),.dout(n894),.clk(gclk));
	jand g0580(.dina(n894),.dinb(w_dff_B_hNhDWOew7_1),.dout(n895),.clk(gclk));
	jxor g0581(.dina(w_n895_1[1]),.dinb(w_n891_1[1]),.dout(n896),.clk(gclk));
	jnot g0582(.din(w_n434_0[0]),.dout(n897),.clk(gclk));
	jand g0583(.dina(G203),.dinb(w_G18_33[0]),.dout(n898),.clk(gclk));
	jor g0584(.dina(w_dff_B_7XSr0N1X0_0),.dinb(n897),.dout(n899),.clk(gclk));
	jor g0585(.dina(G53),.dinb(w_G18_32[2]),.dout(n900),.clk(gclk));
	jor g0586(.dina(w_n430_0[0]),.dinb(w_n355_15[2]),.dout(n901),.clk(gclk));
	jand g0587(.dina(n901),.dinb(w_dff_B_IUEL5QAU1_1),.dout(n902),.clk(gclk));
	jxor g0588(.dina(w_n902_0[2]),.dinb(w_n899_0[2]),.dout(n903),.clk(gclk));
	jand g0589(.dina(n903),.dinb(w_n896_0[1]),.dout(n904),.clk(gclk));
	jand g0590(.dina(w_dff_B_UPaggQHO7_0),.dinb(w_n889_0[1]),.dout(n905),.clk(gclk));
	jnot g0591(.din(w_n400_0[0]),.dout(n906),.clk(gclk));
	jand g0592(.dina(G207),.dinb(w_G18_32[1]),.dout(n907),.clk(gclk));
	jor g0593(.dina(w_dff_B_fPYqTgMv3_0),.dinb(n906),.dout(n908),.clk(gclk));
	jor g0594(.dina(G74),.dinb(w_G18_32[0]),.dout(n909),.clk(gclk));
	jand g0595(.dina(w_G3705_1[2]),.dinb(w_G18_31[2]),.dout(n910),.clk(gclk));
	jnot g0596(.din(n910),.dout(n911),.clk(gclk));
	jand g0597(.dina(n911),.dinb(w_dff_B_Bh5QiV947_1),.dout(n912),.clk(gclk));
	jor g0598(.dina(w_n912_0[2]),.dinb(w_n908_0[2]),.dout(n913),.clk(gclk));
	jnot g0599(.din(w_n376_0[0]),.dout(n914),.clk(gclk));
	jand g0600(.dina(G205),.dinb(w_G18_31[1]),.dout(n915),.clk(gclk));
	jor g0601(.dina(w_dff_B_rVvKV7Bp3_0),.dinb(n914),.dout(n916),.clk(gclk));
	jor g0602(.dina(G75),.dinb(w_G18_31[0]),.dout(n917),.clk(gclk));
	jand g0603(.dina(w_G3717_1[2]),.dinb(w_G18_30[2]),.dout(n918),.clk(gclk));
	jnot g0604(.din(n918),.dout(n919),.clk(gclk));
	jand g0605(.dina(n919),.dinb(w_dff_B_uXICOqHD1_1),.dout(n920),.clk(gclk));
	jor g0606(.dina(w_n920_0[2]),.dinb(w_n916_0[2]),.dout(n921),.clk(gclk));
	jand g0607(.dina(w_n921_0[1]),.dinb(w_n913_0[1]),.dout(n922),.clk(gclk));
	jand g0608(.dina(w_n920_0[1]),.dinb(w_n916_0[1]),.dout(n923),.clk(gclk));
	jnot g0609(.din(w_n923_0[1]),.dout(n924),.clk(gclk));
	jnot g0610(.din(w_n385_0[0]),.dout(n925),.clk(gclk));
	jand g0611(.dina(G206),.dinb(w_G18_30[1]),.dout(n926),.clk(gclk));
	jor g0612(.dina(w_dff_B_PhDfeFx85_0),.dinb(n925),.dout(n927),.clk(gclk));
	jor g0613(.dina(G76),.dinb(w_G18_30[0]),.dout(n928),.clk(gclk));
	jand g0614(.dina(w_G3711_0[2]),.dinb(w_G18_29[2]),.dout(n929),.clk(gclk));
	jnot g0615(.din(n929),.dout(n930),.clk(gclk));
	jand g0616(.dina(n930),.dinb(w_dff_B_zE8vol1i0_1),.dout(n931),.clk(gclk));
	jor g0617(.dina(w_n931_0[2]),.dinb(w_n927_0[2]),.dout(n932),.clk(gclk));
	jand g0618(.dina(w_n932_0[1]),.dinb(n924),.dout(n933),.clk(gclk));
	jand g0619(.dina(n933),.dinb(w_dff_B_La6IPfwy8_1),.dout(n934),.clk(gclk));
	jnot g0620(.din(w_G70_0[1]),.dout(n935),.clk(gclk));
	jand g0621(.dina(w_n935_0[1]),.dinb(w_n355_15[1]),.dout(n936),.clk(gclk));
	jnot g0622(.din(n936),.dout(n937),.clk(gclk));
	jor g0623(.dina(w_n937_0[1]),.dinb(w_G41_0[0]),.dout(n938),.clk(gclk));
	jand g0624(.dina(w_n937_0[0]),.dinb(w_n356_0[0]),.dout(n939),.clk(gclk));
	jnot g0625(.din(w_n939_0[1]),.dout(n940),.clk(gclk));
	jand g0626(.dina(n940),.dinb(w_dff_B_zGP8pgHY2_1),.dout(n941),.clk(gclk));
	jand g0627(.dina(n941),.dinb(w_dff_B_DjlADNOI5_1),.dout(n942),.clk(gclk));
	jnot g0628(.din(w_n370_0[0]),.dout(n943),.clk(gclk));
	jand g0629(.dina(G204),.dinb(w_G18_29[1]),.dout(n944),.clk(gclk));
	jor g0630(.dina(w_dff_B_ppmXzpJe8_0),.dinb(n943),.dout(n945),.clk(gclk));
	jor g0631(.dina(G73),.dinb(w_G18_29[0]),.dout(n946),.clk(gclk));
	jor g0632(.dina(w_n366_0[0]),.dinb(w_n355_15[0]),.dout(n947),.clk(gclk));
	jand g0633(.dina(n947),.dinb(w_dff_B_tcaMqhgn1_1),.dout(n948),.clk(gclk));
	jxor g0634(.dina(w_n948_1[1]),.dinb(w_n945_1[1]),.dout(n949),.clk(gclk));
	jand g0635(.dina(w_n912_0[1]),.dinb(w_n908_0[1]),.dout(n950),.clk(gclk));
	jnot g0636(.din(w_n950_0[1]),.dout(n951),.clk(gclk));
	jand g0637(.dina(w_n931_0[1]),.dinb(w_n927_0[1]),.dout(n952),.clk(gclk));
	jnot g0638(.din(w_n952_0[1]),.dout(n953),.clk(gclk));
	jand g0639(.dina(n953),.dinb(n951),.dout(n954),.clk(gclk));
	jand g0640(.dina(n954),.dinb(w_dff_B_jbgvIvE76_1),.dout(n955),.clk(gclk));
	jand g0641(.dina(n955),.dinb(w_dff_B_hzR408JK2_1),.dout(n956),.clk(gclk));
	jand g0642(.dina(n956),.dinb(w_dff_B_cf8N8jNw3_1),.dout(n957),.clk(gclk));
	jand g0643(.dina(w_n957_0[1]),.dinb(w_n905_0[2]),.dout(n958),.clk(gclk));
	jand g0644(.dina(n958),.dinb(w_n865_0[1]),.dout(n959),.clk(gclk));
	jand g0645(.dina(w_n807_0[1]),.dinb(w_n804_0[1]),.dout(n960),.clk(gclk));
	jand g0646(.dina(n960),.dinb(w_n802_0[0]),.dout(n961),.clk(gclk));
	jand g0647(.dina(n961),.dinb(w_n795_0[0]),.dout(n962),.clk(gclk));
	jand g0648(.dina(w_n793_1[0]),.dinb(w_n790_1[0]),.dout(n963),.clk(gclk));
	jand g0649(.dina(w_n787_0[1]),.dinb(w_n784_0[1]),.dout(n964),.clk(gclk));
	jand g0650(.dina(w_n801_1[0]),.dinb(w_n797_1[0]),.dout(n965),.clk(gclk));
	jor g0651(.dina(n965),.dinb(n964),.dout(n966),.clk(gclk));
	jor g0652(.dina(w_n793_0[2]),.dinb(w_n790_0[2]),.dout(n967),.clk(gclk));
	jor g0653(.dina(w_n801_0[2]),.dinb(w_n797_0[2]),.dout(n968),.clk(gclk));
	jand g0654(.dina(n968),.dinb(n967),.dout(n969),.clk(gclk));
	jand g0655(.dina(n969),.dinb(n966),.dout(n970),.clk(gclk));
	jor g0656(.dina(n970),.dinb(w_dff_B_HRf6BwCS8_1),.dout(n971),.clk(gclk));
	jor g0657(.dina(n971),.dinb(w_dff_B_ocApAAlI3_1),.dout(n972),.clk(gclk));
	jand g0658(.dina(w_n832_0[0]),.dinb(w_n817_0[0]),.dout(n973),.clk(gclk));
	jor g0659(.dina(w_n838_0[0]),.dinb(w_n834_0[0]),.dout(n974),.clk(gclk));
	jor g0660(.dina(n974),.dinb(n973),.dout(n975),.clk(gclk));
	jand g0661(.dina(w_n858_0[1]),.dinb(w_n856_0[0]),.dout(n976),.clk(gclk));
	jand g0662(.dina(n976),.dinb(w_n824_0[0]),.dout(n977),.clk(gclk));
	jand g0663(.dina(n977),.dinb(n975),.dout(n978),.clk(gclk));
	jand g0664(.dina(w_n859_0[0]),.dinb(w_n858_0[0]),.dout(n979),.clk(gclk));
	jor g0665(.dina(n979),.dinb(w_n848_0[0]),.dout(n980),.clk(gclk));
	jor g0666(.dina(w_dff_B_BaWeFQ4N1_0),.dinb(n978),.dout(n981),.clk(gclk));
	jand g0667(.dina(w_n981_0[1]),.dinb(w_n810_0[1]),.dout(n982),.clk(gclk));
	jor g0668(.dina(n982),.dinb(w_n972_0[1]),.dout(n983),.clk(gclk));
	jor g0669(.dina(w_dff_B_X0fm0r7M0_0),.dinb(n959),.dout(n984),.clk(gclk));
	jand g0670(.dina(n984),.dinb(w_n782_0[1]),.dout(n985),.clk(gclk));
	jor g0671(.dina(n985),.dinb(w_dff_B_omwt6g2n2_1),.dout(n986),.clk(gclk));
	jor g0672(.dina(w_dff_B_OEvkFNga5_0),.dinb(w_n355_14[2]),.dout(n987),.clk(gclk));
	jand g0673(.dina(w_n987_0[1]),.dinb(w_n565_6[2]),.dout(n988),.clk(gclk));
	jand g0674(.dina(w_G2256_0[2]),.dinb(w_G18_28[2]),.dout(n989),.clk(gclk));
	jnot g0675(.din(n989),.dout(n990),.clk(gclk));
	jor g0676(.dina(G110),.dinb(w_G18_28[1]),.dout(n991),.clk(gclk));
	jand g0677(.dina(w_dff_B_l5t1Lzlf2_0),.dinb(n990),.dout(n992),.clk(gclk));
	jor g0678(.dina(w_n992_0[2]),.dinb(w_n988_0[2]),.dout(n993),.clk(gclk));
	jor g0679(.dina(w_dff_B_kwT9n1fz3_0),.dinb(w_n355_14[1]),.dout(n994),.clk(gclk));
	jand g0680(.dina(w_n994_0[1]),.dinb(w_n565_6[1]),.dout(n995),.clk(gclk));
	jand g0681(.dina(w_G2247_0[1]),.dinb(w_G18_28[0]),.dout(n996),.clk(gclk));
	jnot g0682(.din(n996),.dout(n997),.clk(gclk));
	jor g0683(.dina(G86),.dinb(w_G18_27[2]),.dout(n998),.clk(gclk));
	jand g0684(.dina(w_dff_B_gbjOsGnH4_0),.dinb(n997),.dout(n999),.clk(gclk));
	jand g0685(.dina(w_n999_0[2]),.dinb(w_n995_0[2]),.dout(n1000),.clk(gclk));
	jnot g0686(.din(w_n1000_0[1]),.dout(n1001),.clk(gclk));
	jand g0687(.dina(n1001),.dinb(w_n993_0[1]),.dout(n1002),.clk(gclk));
	jand g0688(.dina(w_n992_0[1]),.dinb(w_n988_0[1]),.dout(n1003),.clk(gclk));
	jnot g0689(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jor g0690(.dina(w_n999_0[1]),.dinb(w_n995_0[1]),.dout(n1005),.clk(gclk));
	jand g0691(.dina(w_dff_B_A2vgLadr0_0),.dinb(n1004),.dout(n1006),.clk(gclk));
	jand g0692(.dina(n1006),.dinb(n1002),.dout(n1007),.clk(gclk));
	jor g0693(.dina(w_dff_B_ZhNlUfdm8_0),.dinb(w_n355_14[0]),.dout(n1008),.clk(gclk));
	jand g0694(.dina(w_n1008_0[1]),.dinb(w_n565_6[0]),.dout(n1009),.clk(gclk));
	jand g0695(.dina(w_G2253_0[2]),.dinb(w_G18_27[1]),.dout(n1010),.clk(gclk));
	jnot g0696(.din(n1010),.dout(n1011),.clk(gclk));
	jor g0697(.dina(G109),.dinb(w_G18_27[0]),.dout(n1012),.clk(gclk));
	jand g0698(.dina(w_dff_B_eCcZfGh83_0),.dinb(n1011),.dout(n1013),.clk(gclk));
	jxor g0699(.dina(w_n1013_1[1]),.dinb(w_n1009_1[1]),.dout(n1014),.clk(gclk));
	jor g0700(.dina(w_dff_B_bRo8Z4hO6_0),.dinb(w_n355_13[2]),.dout(n1015),.clk(gclk));
	jand g0701(.dina(w_n1015_0[1]),.dinb(w_n565_5[2]),.dout(n1016),.clk(gclk));
	jor g0702(.dina(w_n623_0[0]),.dinb(w_n355_13[1]),.dout(n1017),.clk(gclk));
	jor g0703(.dina(G63),.dinb(w_G18_26[2]),.dout(n1018),.clk(gclk));
	jand g0704(.dina(w_dff_B_UY3GNvtW9_0),.dinb(n1017),.dout(n1019),.clk(gclk));
	jxor g0705(.dina(w_n1019_0[2]),.dinb(w_n1016_0[2]),.dout(n1020),.clk(gclk));
	jand g0706(.dina(n1020),.dinb(w_n1014_0[1]),.dout(n1021),.clk(gclk));
	jand g0707(.dina(w_dff_B_fECzl2j29_0),.dinb(w_n1007_0[1]),.dout(n1022),.clk(gclk));
	jand g0708(.dina(w_n1022_0[1]),.dinb(n986),.dout(n1023),.clk(gclk));
	jand g0709(.dina(w_n948_1[0]),.dinb(w_n945_1[0]),.dout(n1024),.clk(gclk));
	jor g0710(.dina(w_n950_0[0]),.dinb(w_n939_0[0]),.dout(n1025),.clk(gclk));
	jand g0711(.dina(w_n932_0[0]),.dinb(w_n913_0[0]),.dout(n1026),.clk(gclk));
	jand g0712(.dina(n1026),.dinb(n1025),.dout(n1027),.clk(gclk));
	jor g0713(.dina(w_n952_0[0]),.dinb(w_n923_0[0]),.dout(n1028),.clk(gclk));
	jor g0714(.dina(w_dff_B_0r9OQegj7_0),.dinb(n1027),.dout(n1029),.clk(gclk));
	jor g0715(.dina(w_n948_0[2]),.dinb(w_n945_0[2]),.dout(n1030),.clk(gclk));
	jand g0716(.dina(n1030),.dinb(w_n921_0[0]),.dout(n1031),.clk(gclk));
	jand g0717(.dina(w_dff_B_QS8e2wgJ2_0),.dinb(n1029),.dout(n1032),.clk(gclk));
	jor g0718(.dina(n1032),.dinb(w_dff_B_VebpQi8Y0_1),.dout(n1033),.clk(gclk));
	jand g0719(.dina(w_n1033_0[1]),.dinb(w_n905_0[1]),.dout(n1034),.clk(gclk));
	jand g0720(.dina(w_n902_0[1]),.dinb(w_n899_0[1]),.dout(n1035),.clk(gclk));
	jand g0721(.dina(n1035),.dinb(w_n896_0[0]),.dout(n1036),.clk(gclk));
	jand g0722(.dina(w_dff_B_ipreZXo37_0),.dinb(w_n889_0[0]),.dout(n1037),.clk(gclk));
	jand g0723(.dina(w_n895_1[0]),.dinb(w_n891_1[0]),.dout(n1038),.clk(gclk));
	jor g0724(.dina(w_dff_B_bSp9X1LY2_0),.dinb(w_n885_0[0]),.dout(n1039),.clk(gclk));
	jor g0725(.dina(w_n895_0[2]),.dinb(w_n891_0[2]),.dout(n1040),.clk(gclk));
	jand g0726(.dina(w_dff_B_yYE49MnY2_0),.dinb(w_n887_0[0]),.dout(n1041),.clk(gclk));
	jand g0727(.dina(n1041),.dinb(n1039),.dout(n1042),.clk(gclk));
	jor g0728(.dina(n1042),.dinb(w_n874_0[0]),.dout(n1043),.clk(gclk));
	jor g0729(.dina(w_dff_B_73b3XT5p2_0),.dinb(n1037),.dout(n1044),.clk(gclk));
	jor g0730(.dina(w_n1044_0[1]),.dinb(n1034),.dout(n1045),.clk(gclk));
	jand g0731(.dina(w_n1022_0[0]),.dinb(w_n782_0[0]),.dout(n1046),.clk(gclk));
	jand g0732(.dina(n1046),.dinb(w_n865_0[0]),.dout(n1047),.clk(gclk));
	jand g0733(.dina(w_dff_B_yrJTjGSX8_0),.dinb(n1045),.dout(n1048),.clk(gclk));
	jand g0734(.dina(w_n1019_0[1]),.dinb(w_n1016_0[1]),.dout(n1049),.clk(gclk));
	jand g0735(.dina(n1049),.dinb(w_n1014_0[0]),.dout(n1050),.clk(gclk));
	jand g0736(.dina(w_dff_B_Szp1HVeJ0_0),.dinb(w_n1007_0[0]),.dout(n1051),.clk(gclk));
	jand g0737(.dina(w_n1013_1[0]),.dinb(w_n1009_1[0]),.dout(n1052),.clk(gclk));
	jor g0738(.dina(n1052),.dinb(w_n1000_0[0]),.dout(n1053),.clk(gclk));
	jor g0739(.dina(w_n1013_0[2]),.dinb(w_n1009_0[2]),.dout(n1054),.clk(gclk));
	jand g0740(.dina(n1054),.dinb(w_n993_0[0]),.dout(n1055),.clk(gclk));
	jand g0741(.dina(n1055),.dinb(n1053),.dout(n1056),.clk(gclk));
	jor g0742(.dina(n1056),.dinb(w_n1003_0[0]),.dout(n1057),.clk(gclk));
	jor g0743(.dina(w_dff_B_xLARylk14_0),.dinb(n1051),.dout(n1058),.clk(gclk));
	jor g0744(.dina(w_dff_B_Qusatsm47_0),.dinb(n1048),.dout(n1059),.clk(gclk));
	jor g0745(.dina(w_dff_B_owubJqtn6_0),.dinb(n1023),.dout(n1060),.clk(gclk));
	jor g0746(.dina(w_dff_B_FnEjt97S5_0),.dinb(w_n355_13[0]),.dout(n1061),.clk(gclk));
	jand g0747(.dina(w_n1061_0[2]),.dinb(w_n565_5[1]),.dout(n1062),.clk(gclk));
	jand g0748(.dina(w_G1480_0[1]),.dinb(w_G18_26[1]),.dout(n1063),.clk(gclk));
	jnot g0749(.din(n1063),.dout(n1064),.clk(gclk));
	jor g0750(.dina(G112),.dinb(w_G18_26[0]),.dout(n1065),.clk(gclk));
	jand g0751(.dina(w_dff_B_zwpHeb496_0),.dinb(n1064),.dout(n1066),.clk(gclk));
	jor g0752(.dina(w_n1066_0[2]),.dinb(w_n1062_0[1]),.dout(n1067),.clk(gclk));
	jor g0753(.dina(w_dff_B_b19WWDy46_0),.dinb(w_n355_12[2]),.dout(n1068),.clk(gclk));
	jand g0754(.dina(w_n1068_0[1]),.dinb(w_n565_5[0]),.dout(n1069),.clk(gclk));
	jand g0755(.dina(w_G1486_0[1]),.dinb(w_G18_25[2]),.dout(n1070),.clk(gclk));
	jnot g0756(.din(n1070),.dout(n1071),.clk(gclk));
	jor g0757(.dina(G88),.dinb(w_G18_25[1]),.dout(n1072),.clk(gclk));
	jand g0758(.dina(w_dff_B_FkoeeYcx3_0),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0759(.dina(w_n1073_0[2]),.dinb(w_n1069_0[1]),.dout(n1074),.clk(gclk));
	jand g0760(.dina(n1074),.dinb(n1067),.dout(n1075),.clk(gclk));
	jor g0761(.dina(w_dff_B_t28gJu808_0),.dinb(w_n355_12[1]),.dout(n1076),.clk(gclk));
	jand g0762(.dina(w_n1076_0[1]),.dinb(w_n565_4[2]),.dout(n1077),.clk(gclk));
	jand g0763(.dina(w_G1469_0[2]),.dinb(w_G18_25[0]),.dout(n1078),.clk(gclk));
	jnot g0764(.din(n1078),.dout(n1079),.clk(gclk));
	jor g0765(.dina(G111),.dinb(w_G18_24[2]),.dout(n1080),.clk(gclk));
	jand g0766(.dina(w_dff_B_6eM1AfF22_0),.dinb(n1079),.dout(n1081),.clk(gclk));
	jor g0767(.dina(w_n1081_0[2]),.dinb(w_n1077_0[2]),.dout(n1082),.clk(gclk));
	jand g0768(.dina(w_G1462_0[1]),.dinb(w_G18_24[1]),.dout(n1083),.clk(gclk));
	jnot g0769(.din(n1083),.dout(n1084),.clk(gclk));
	jor g0770(.dina(G113),.dinb(w_G18_24[0]),.dout(n1085),.clk(gclk));
	jand g0771(.dina(w_dff_B_4F3mVGZg2_0),.dinb(n1084),.dout(n1086),.clk(gclk));
	jor g0772(.dina(w_n1086_0[2]),.dinb(w_n565_4[1]),.dout(n1087),.clk(gclk));
	jand g0773(.dina(n1087),.dinb(w_n1082_0[1]),.dout(n1088),.clk(gclk));
	jand g0774(.dina(n1088),.dinb(w_n1075_0[1]),.dout(n1089),.clk(gclk));
	jand g0775(.dina(w_n1081_0[1]),.dinb(w_n1077_0[1]),.dout(n1090),.clk(gclk));
	jand g0776(.dina(w_n1086_0[1]),.dinb(w_n565_4[0]),.dout(n1091),.clk(gclk));
	jor g0777(.dina(n1091),.dinb(n1090),.dout(n1092),.clk(gclk));
	jnot g0778(.din(w_n1092_0[1]),.dout(n1093),.clk(gclk));
	jand g0779(.dina(w_n1066_0[1]),.dinb(w_n1062_0[0]),.dout(n1094),.clk(gclk));
	jor g0780(.dina(w_dff_B_7fLkiLQM3_0),.dinb(w_n355_12[0]),.dout(n1095),.clk(gclk));
	jand g0781(.dina(w_n1095_0[1]),.dinb(w_n565_3[2]),.dout(n1096),.clk(gclk));
	jand g0782(.dina(w_G106_0[2]),.dinb(w_G18_23[2]),.dout(n1097),.clk(gclk));
	jnot g0783(.din(n1097),.dout(n1098),.clk(gclk));
	jor g0784(.dina(G87),.dinb(w_G18_23[1]),.dout(n1099),.clk(gclk));
	jand g0785(.dina(w_dff_B_R6DqXCQT1_0),.dinb(n1098),.dout(n1100),.clk(gclk));
	jand g0786(.dina(w_n1100_0[2]),.dinb(w_n1096_0[2]),.dout(n1101),.clk(gclk));
	jor g0787(.dina(n1101),.dinb(n1094),.dout(n1102),.clk(gclk));
	jnot g0788(.din(w_n1102_0[1]),.dout(n1103),.clk(gclk));
	jor g0789(.dina(w_n1100_0[1]),.dinb(w_n1096_0[1]),.dout(n1104),.clk(gclk));
	jand g0790(.dina(w_n1073_0[1]),.dinb(w_n1069_0[0]),.dout(n1105),.clk(gclk));
	jnot g0791(.din(w_n1105_0[1]),.dout(n1106),.clk(gclk));
	jand g0792(.dina(n1106),.dinb(w_n1104_0[1]),.dout(n1107),.clk(gclk));
	jand g0793(.dina(n1107),.dinb(n1103),.dout(n1108),.clk(gclk));
	jand g0794(.dina(n1108),.dinb(w_dff_B_ucUW0KpF7_1),.dout(n1109),.clk(gclk));
	jand g0795(.dina(n1109),.dinb(w_dff_B_Taz8ROiW9_1),.dout(n1110),.clk(gclk));
	jand g0796(.dina(w_dff_B_sybW8anM3_0),.dinb(n1060),.dout(n1111),.clk(gclk));
	jand g0797(.dina(w_n1104_0[0]),.dinb(w_n1082_0[0]),.dout(n1112),.clk(gclk));
	jand g0798(.dina(n1112),.dinb(w_n1092_0[0]),.dout(n1113),.clk(gclk));
	jor g0799(.dina(n1113),.dinb(w_n1102_0[0]),.dout(n1114),.clk(gclk));
	jand g0800(.dina(n1114),.dinb(w_n1075_0[0]),.dout(n1115),.clk(gclk));
	jnot g0801(.din(w_G4528_0[0]),.dout(n1116),.clk(gclk));
	jor g0802(.dina(w_G2204_0[2]),.dinb(w_G1455_0[2]),.dout(n1117),.clk(gclk));
	jor g0803(.dina(n1117),.dinb(w_n1116_0[1]),.dout(n1118),.clk(gclk));
	jand g0804(.dina(n1118),.dinb(w_G38_0[2]),.dout(n1119),.clk(gclk));
	jor g0805(.dina(w_dff_B_xZjP3xbI8_0),.dinb(w_n1105_0[0]),.dout(n1120),.clk(gclk));
	jor g0806(.dina(w_dff_B_PlJ4JVtI2_0),.dinb(n1115),.dout(n1121),.clk(gclk));
	jor g0807(.dina(w_dff_B_eaos86KW9_0),.dinb(n1111),.dout(n1122),.clk(gclk));
	jand g0808(.dina(w_G2204_0[1]),.dinb(w_G1455_0[1]),.dout(n1123),.clk(gclk));
	jor g0809(.dina(w_n1116_0[0]),.dinb(w_G38_0[1]),.dout(n1124),.clk(gclk));
	jor g0810(.dina(n1124),.dinb(w_dff_B_nmwzeh3H7_1),.dout(n1125),.clk(gclk));
	jand g0811(.dina(w_n1125_0[2]),.dinb(w_n1122_0[2]),.dout(w_dff_A_Q0JJXQ6q2_2),.clk(gclk));
	jand g0812(.dina(w_n377_1[0]),.dinb(w_G3717_1[1]),.dout(n1127),.clk(gclk));
	jand g0813(.dina(w_n413_1[0]),.dinb(w_n410_0[0]),.dout(n1128),.clk(gclk));
	jor g0814(.dina(w_n1128_1[1]),.dinb(w_n1127_0[1]),.dout(n1129),.clk(gclk));
	jand g0815(.dina(n1129),.dinb(w_n417_0[1]),.dout(n1130),.clk(gclk));
	jor g0816(.dina(w_n405_0[1]),.dinb(w_n379_1[0]),.dout(n1131),.clk(gclk));
	jand g0817(.dina(w_dff_B_aOYLngUM6_0),.dinb(w_n1130_0[1]),.dout(n1132),.clk(gclk));
	jxor g0818(.dina(n1132),.dinb(w_n372_1[1]),.dout(w_dff_A_l9LCgxGv9_2),.clk(gclk));
	jand g0819(.dina(w_n1128_1[0]),.dinb(w_n405_0[0]),.dout(n1134),.clk(gclk));
	jxor g0820(.dina(n1134),.dinb(w_n379_0[2]),.dout(w_dff_A_f4MjxiJZ3_2),.clk(gclk));
	jand g0821(.dina(w_n408_0[0]),.dinb(w_n412_0[1]),.dout(n1136),.clk(gclk));
	jand g0822(.dina(w_n1136_0[1]),.dinb(w_n404_0[0]),.dout(n1137),.clk(gclk));
	jxor g0823(.dina(n1137),.dinb(w_n387_0[2]),.dout(w_dff_A_wd3queQl0_2),.clk(gclk));
	jor g0824(.dina(w_n395_0[1]),.dinb(w_n388_0[1]),.dout(n1139),.clk(gclk));
	jand g0825(.dina(n1139),.dinb(w_n354_1[0]),.dout(n1140),.clk(gclk));
	jxor g0826(.dina(n1140),.dinb(w_n402_0[2]),.dout(w_dff_A_vEddeJa75_2),.clk(gclk));
	jor g0827(.dina(w_n437_0[0]),.dinb(w_n422_1[1]),.dout(n1142),.clk(gclk));
	jor g0828(.dina(w_n1142_0[1]),.dinb(w_n456_0[1]),.dout(n1143),.clk(gclk));
	jand g0829(.dina(n1143),.dinb(w_n462_0[1]),.dout(n1144),.clk(gclk));
	jxor g0830(.dina(n1144),.dinb(w_n446_1[0]),.dout(w_dff_A_KMCbaGeF1_2),.clk(gclk));
	jand g0831(.dina(w_n1142_0[0]),.dinb(w_n460_0[1]),.dout(n1146),.clk(gclk));
	jxor g0832(.dina(n1146),.dinb(w_n450_0[1]),.dout(w_dff_A_8VidLIuF6_2),.clk(gclk));
	jand g0833(.dina(w_n435_0[2]),.dinb(w_G3729_0[2]),.dout(n1148),.clk(gclk));
	jor g0834(.dina(w_n1148_0[2]),.dinb(w_n422_1[0]),.dout(n1149),.clk(gclk));
	jand g0835(.dina(n1149),.dinb(w_n458_0[1]),.dout(n1150),.clk(gclk));
	jxor g0836(.dina(n1150),.dinb(w_n429_1[2]),.dout(w_dff_A_f3sHIXSK4_2),.clk(gclk));
	jxor g0837(.dina(w_n436_0[0]),.dinb(w_n422_0[2]),.dout(w_dff_A_H03IRAWS8_2),.clk(gclk));
	jxor g0838(.dina(w_n583_0[1]),.dinb(w_n577_0[0]),.dout(n1153),.clk(gclk));
	jxor g0839(.dina(w_n588_0[1]),.dinb(w_n567_0[1]),.dout(n1154),.clk(gclk));
	jxor g0840(.dina(n1154),.dinb(w_n572_0[2]),.dout(n1155),.clk(gclk));
	jnot g0841(.din(w_n625_0[0]),.dout(n1156),.clk(gclk));
	jor g0842(.dina(w_n1156_0[1]),.dinb(w_n620_0[0]),.dout(n1157),.clk(gclk));
	jnot g0843(.din(w_n621_0[0]),.dout(n1158),.clk(gclk));
	jor g0844(.dina(w_n624_0[0]),.dinb(n1158),.dout(n1159),.clk(gclk));
	jand g0845(.dina(n1159),.dinb(n1157),.dout(n1160),.clk(gclk));
	jor g0846(.dina(w_n652_0[0]),.dinb(w_n629_0[0]),.dout(n1161),.clk(gclk));
	jor g0847(.dina(w_n633_0[0]),.dinb(w_n650_0[0]),.dout(n1162),.clk(gclk));
	jand g0848(.dina(n1162),.dinb(n1161),.dout(n1163),.clk(gclk));
	jxor g0849(.dina(n1163),.dinb(n1160),.dout(n1164),.clk(gclk));
	jnot g0850(.din(G141),.dout(n1165),.clk(gclk));
	jor g0851(.dina(n1165),.dinb(w_G18_23[0]),.dout(n1166),.clk(gclk));
	jnot g0852(.din(G161),.dout(n1167),.clk(gclk));
	jor g0853(.dina(n1167),.dinb(w_n355_11[2]),.dout(n1168),.clk(gclk));
	jand g0854(.dina(n1168),.dinb(w_n1166_0[1]),.dout(n1169),.clk(gclk));
	jxor g0855(.dina(w_dff_B_bpWNMMEc7_0),.dinb(n1164),.dout(n1170),.clk(gclk));
	jxor g0856(.dina(n1170),.dinb(w_dff_B_ORUhP1w48_1),.dout(n1171),.clk(gclk));
	jxor g0857(.dina(n1171),.dinb(w_dff_B_Z1bZWMPx7_1),.dout(n1172),.clk(gclk));
	jand g0858(.dina(w_n565_3[1]),.dinb(w_G18_22[2]),.dout(n1173),.clk(gclk));
	jxor g0859(.dina(G212),.dinb(G211),.dout(n1174),.clk(gclk));
	jand g0860(.dina(w_dff_B_tDGVdp7M2_0),.dinb(w_n1173_0[1]),.dout(n1175),.clk(gclk));
	jor g0861(.dina(w_n676_0[0]),.dinb(w_n564_0[1]),.dout(n1176),.clk(gclk));
	jnot g0862(.din(w_n659_0[0]),.dout(n1177),.clk(gclk));
	jand g0863(.dina(w_n664_0[1]),.dinb(n1177),.dout(n1178),.clk(gclk));
	jnot g0864(.din(w_n663_0[0]),.dout(n1179),.clk(gclk));
	jand g0865(.dina(n1179),.dinb(w_n660_0[1]),.dout(n1180),.clk(gclk));
	jor g0866(.dina(n1180),.dinb(n1178),.dout(n1181),.clk(gclk));
	jor g0867(.dina(w_n693_0[0]),.dinb(w_n667_0[0]),.dout(n1182),.clk(gclk));
	jor g0868(.dina(w_n672_0[0]),.dinb(w_n690_0[0]),.dout(n1183),.clk(gclk));
	jand g0869(.dina(n1183),.dinb(n1182),.dout(n1184),.clk(gclk));
	jxor g0870(.dina(n1184),.dinb(w_dff_B_BdmlA7k07_1),.dout(n1185),.clk(gclk));
	jxor g0871(.dina(n1185),.dinb(w_dff_B_SyQToNJc4_1),.dout(n1186),.clk(gclk));
	jxor g0872(.dina(n1186),.dinb(w_dff_B_Y3DHXPlw4_1),.dout(n1187),.clk(gclk));
	jand g0873(.dina(G239),.dinb(w_G18_22[1]),.dout(n1188),.clk(gclk));
	jand g0874(.dina(w_dff_B_ACQkRp2d8_0),.dinb(w_n355_11[1]),.dout(n1189),.clk(gclk));
	jor g0875(.dina(w_n1189_0[1]),.dinb(w_dff_B_uzyJlzBQ0_1),.dout(n1190),.clk(gclk));
	jxor g0876(.dina(w_n442_0[0]),.dinb(w_n428_0[0]),.dout(n1191),.clk(gclk));
	jxor g0877(.dina(w_n449_0[0]),.dinb(w_n435_0[1]),.dout(n1192),.clk(gclk));
	jxor g0878(.dina(n1192),.dinb(n1191),.dout(n1193),.clk(gclk));
	jxor g0879(.dina(n1193),.dinb(w_dff_B_EhhukHxl3_1),.dout(n1194),.clk(gclk));
	jxor g0880(.dina(w_n401_1[0]),.dinb(w_n371_0[1]),.dout(n1195),.clk(gclk));
	jxor g0881(.dina(n1195),.dinb(w_n377_0[2]),.dout(n1196),.clk(gclk));
	jxor g0882(.dina(w_n386_0[0]),.dinb(w_n358_0[0]),.dout(n1197),.clk(gclk));
	jxor g0883(.dina(w_dff_B_fWbOweMG4_0),.dinb(n1196),.dout(n1198),.clk(gclk));
	jxor g0884(.dina(n1198),.dinb(n1194),.dout(n1199),.clk(gclk));
	jxor g0885(.dina(w_n534_0[1]),.dinb(w_n523_0[0]),.dout(n1200),.clk(gclk));
	jxor g0886(.dina(w_n539_0[1]),.dinb(w_n528_0[2]),.dout(n1201),.clk(gclk));
	jxor g0887(.dina(n1201),.dinb(n1200),.dout(n1202),.clk(gclk));
	jxor g0888(.dina(n1202),.dinb(w_n503_0[0]),.dout(n1203),.clk(gclk));
	jand g0889(.dina(G227),.dinb(w_G18_22[0]),.dout(n1204),.clk(gclk));
	jand g0890(.dina(w_dff_B_lMdIjjqA3_0),.dinb(w_n355_11[0]),.dout(n1205),.clk(gclk));
	jor g0891(.dina(w_n1205_0[1]),.dinb(w_dff_B_NHTV8UlK1_1),.dout(n1206),.clk(gclk));
	jxor g0892(.dina(w_n489_0[0]),.dinb(w_n478_0[0]),.dout(n1207),.clk(gclk));
	jxor g0893(.dina(n1207),.dinb(w_dff_B_HWQXCFiG4_1),.dout(n1208),.clk(gclk));
	jxor g0894(.dina(w_n474_0[2]),.dinb(w_n469_0[1]),.dout(n1209),.clk(gclk));
	jxor g0895(.dina(w_dff_B_Q74RQj760_0),.dinb(n1208),.dout(n1210),.clk(gclk));
	jxor g0896(.dina(n1210),.dinb(n1203),.dout(n1211),.clk(gclk));
	jor g0897(.dina(n1211),.dinb(n1199),.dout(n1212),.clk(gclk));
	jor g0898(.dina(w_dff_B_173T7hMJ2_0),.dinb(n1187),.dout(n1213),.clk(gclk));
	jor g0899(.dina(n1213),.dinb(n1172),.dout(G412_fa_),.clk(gclk));
	jxor g0900(.dina(w_n831_0[0]),.dinb(w_n823_0[0]),.dout(n1215),.clk(gclk));
	jxor g0901(.dina(w_n847_0[0]),.dinb(w_n816_0[0]),.dout(n1216),.clk(gclk));
	jxor g0902(.dina(n1216),.dinb(w_n855_0[0]),.dout(n1217),.clk(gclk));
	jxor g0903(.dina(w_n793_0[1]),.dinb(w_n787_0[0]),.dout(n1218),.clk(gclk));
	jxor g0904(.dina(w_n807_0[0]),.dinb(w_n801_0[1]),.dout(n1219),.clk(gclk));
	jxor g0905(.dina(n1219),.dinb(n1218),.dout(n1220),.clk(gclk));
	jor g0906(.dina(w_G4393_0[1]),.dinb(w_n355_10[2]),.dout(n1221),.clk(gclk));
	jnot g0907(.din(G58),.dout(n1222),.clk(gclk));
	jor g0908(.dina(n1222),.dinb(w_G18_21[2]),.dout(n1223),.clk(gclk));
	jand g0909(.dina(n1223),.dinb(n1221),.dout(n1224),.clk(gclk));
	jxor g0910(.dina(w_dff_B_8LCFIIXv6_0),.dinb(n1220),.dout(n1225),.clk(gclk));
	jxor g0911(.dina(n1225),.dinb(w_dff_B_SJTdq7ix4_1),.dout(n1226),.clk(gclk));
	jxor g0912(.dina(n1226),.dinb(w_dff_B_DbGk8HA50_1),.dout(n1227),.clk(gclk));
	jxor g0913(.dina(w_n389_0[0]),.dinb(w_G3698_0[1]),.dout(n1228),.clk(gclk));
	jor g0914(.dina(n1228),.dinb(w_n355_10[1]),.dout(n1229),.clk(gclk));
	jnot g0915(.din(w_G69_0[1]),.dout(n1230),.clk(gclk));
	jand g0916(.dina(w_n935_0[0]),.dinb(n1230),.dout(n1231),.clk(gclk));
	jand g0917(.dina(w_G70_0[0]),.dinb(w_G69_0[0]),.dout(n1232),.clk(gclk));
	jor g0918(.dina(n1232),.dinb(w_G18_21[1]),.dout(n1233),.clk(gclk));
	jor g0919(.dina(n1233),.dinb(n1231),.dout(n1234),.clk(gclk));
	jand g0920(.dina(n1234),.dinb(n1229),.dout(n1235),.clk(gclk));
	jxor g0921(.dina(n1235),.dinb(w_n912_0[0]),.dout(n1236),.clk(gclk));
	jnot g0922(.din(w_n1236_0[1]),.dout(n1237),.clk(gclk));
	jxor g0923(.dina(w_n948_0[1]),.dinb(w_n931_0[0]),.dout(n1238),.clk(gclk));
	jnot g0924(.din(w_n920_0[0]),.dout(n1239),.clk(gclk));
	jxor g0925(.dina(w_n882_0[0]),.dinb(w_n873_0[0]),.dout(n1240),.clk(gclk));
	jxor g0926(.dina(w_n902_0[0]),.dinb(w_n895_0[1]),.dout(n1241),.clk(gclk));
	jxor g0927(.dina(n1241),.dinb(n1240),.dout(n1242),.clk(gclk));
	jxor g0928(.dina(n1242),.dinb(w_dff_B_aLTbXciP5_1),.dout(n1243),.clk(gclk));
	jxor g0929(.dina(n1243),.dinb(w_dff_B_fsMbef7P3_1),.dout(n1244),.clk(gclk));
	jnot g0930(.din(w_n1244_0[1]),.dout(n1245),.clk(gclk));
	jand g0931(.dina(n1245),.dinb(w_dff_B_1rCp1k1u8_1),.dout(n1246),.clk(gclk));
	jand g0932(.dina(w_n1244_0[0]),.dinb(w_n1236_0[0]),.dout(n1247),.clk(gclk));
	jor g0933(.dina(w_G1459_0[1]),.dinb(w_n355_10[0]),.dout(n1248),.clk(gclk));
	jnot g0934(.din(G114),.dout(n1249),.clk(gclk));
	jor g0935(.dina(n1249),.dinb(w_G18_21[0]),.dout(n1250),.clk(gclk));
	jand g0936(.dina(n1250),.dinb(n1248),.dout(n1251),.clk(gclk));
	jxor g0937(.dina(w_n1086_0[0]),.dinb(w_n1081_0[0]),.dout(n1252),.clk(gclk));
	jxor g0938(.dina(n1252),.dinb(w_dff_B_hCoIS9vy3_1),.dout(n1253),.clk(gclk));
	jxor g0939(.dina(w_n1100_0[0]),.dinb(w_n1073_0[0]),.dout(n1254),.clk(gclk));
	jxor g0940(.dina(n1254),.dinb(w_n1066_0[0]),.dout(n1255),.clk(gclk));
	jxor g0941(.dina(w_G1496_0[1]),.dinb(w_G1492_0[2]),.dout(n1256),.clk(gclk));
	jor g0942(.dina(n1256),.dinb(w_n355_9[2]),.dout(n1257),.clk(gclk));
	jxor g0943(.dina(w_G2204_0[0]),.dinb(w_G1455_0[0]),.dout(n1258),.clk(gclk));
	jor g0944(.dina(n1258),.dinb(w_G18_20[2]),.dout(n1259),.clk(gclk));
	jand g0945(.dina(n1259),.dinb(n1257),.dout(n1260),.clk(gclk));
	jxor g0946(.dina(w_dff_B_9hGaIqOb4_0),.dinb(n1255),.dout(n1261),.clk(gclk));
	jxor g0947(.dina(n1261),.dinb(w_dff_B_NBUZtjFn9_1),.dout(n1262),.clk(gclk));
	jxor g0948(.dina(w_n999_0[0]),.dinb(w_n992_0[0]),.dout(n1263),.clk(gclk));
	jxor g0949(.dina(w_n1019_0[0]),.dinb(w_n1013_0[1]),.dout(n1264),.clk(gclk));
	jxor g0950(.dina(n1264),.dinb(n1263),.dout(n1265),.clk(gclk));
	jxor g0951(.dina(n1265),.dinb(w_n727_0[0]),.dout(n1266),.clk(gclk));
	jor g0952(.dina(w_G2208_0[1]),.dinb(w_n355_9[1]),.dout(n1267),.clk(gclk));
	jnot g0953(.din(G82),.dout(n1268),.clk(gclk));
	jor g0954(.dina(n1268),.dinb(w_G18_20[1]),.dout(n1269),.clk(gclk));
	jand g0955(.dina(n1269),.dinb(n1267),.dout(n1270),.clk(gclk));
	jxor g0956(.dina(w_n758_0[0]),.dinb(w_n748_0[0]),.dout(n1271),.clk(gclk));
	jxor g0957(.dina(n1271),.dinb(w_dff_B_hfEIVdUV0_1),.dout(n1272),.clk(gclk));
	jxor g0958(.dina(w_n741_0[0]),.dinb(w_n734_0[0]),.dout(n1273),.clk(gclk));
	jxor g0959(.dina(w_dff_B_OP2RUF7k2_0),.dinb(n1272),.dout(n1274),.clk(gclk));
	jxor g0960(.dina(n1274),.dinb(n1266),.dout(n1275),.clk(gclk));
	jor g0961(.dina(n1275),.dinb(n1262),.dout(n1276),.clk(gclk));
	jor g0962(.dina(n1276),.dinb(n1247),.dout(n1277),.clk(gclk));
	jor g0963(.dina(n1277),.dinb(n1246),.dout(n1278),.clk(gclk));
	jor g0964(.dina(n1278),.dinb(w_dff_B_W3BPbTjj3_1),.dout(G414_fa_),.clk(gclk));
	jnot g0965(.din(w_n1061_0[1]),.dout(n1280),.clk(gclk));
	jnot g0966(.din(G170),.dout(n1281),.clk(gclk));
	jand g0967(.dina(n1281),.dinb(w_G18_20[0]),.dout(n1282),.clk(gclk));
	jxor g0968(.dina(n1282),.dinb(w_n1068_0[0]),.dout(n1283),.clk(gclk));
	jnot g0969(.din(w_n1283_0[1]),.dout(n1284),.clk(gclk));
	jand g0970(.dina(n1284),.dinb(w_dff_B_cmy3iLci6_1),.dout(n1285),.clk(gclk));
	jand g0971(.dina(w_n1283_0[0]),.dinb(w_n1061_0[0]),.dout(n1286),.clk(gclk));
	jor g0972(.dina(n1286),.dinb(w_n564_0[0]),.dout(n1287),.clk(gclk));
	jor g0973(.dina(n1287),.dinb(n1285),.dout(n1288),.clk(gclk));
	jnot g0974(.din(w_n1077_0[0]),.dout(n1289),.clk(gclk));
	jor g0975(.dina(w_n1095_0[0]),.dinb(n1289),.dout(n1290),.clk(gclk));
	jnot g0976(.din(w_n1096_0[0]),.dout(n1291),.clk(gclk));
	jor g0977(.dina(n1291),.dinb(w_n1076_0[0]),.dout(n1292),.clk(gclk));
	jand g0978(.dina(n1292),.dinb(n1290),.dout(n1293),.clk(gclk));
	jxor g0979(.dina(G165),.dinb(G164),.dout(n1294),.clk(gclk));
	jand g0980(.dina(w_dff_B_mxs537I87_0),.dinb(w_n1173_0[0]),.dout(n1295),.clk(gclk));
	jxor g0981(.dina(w_dff_B_P2YIAgvt6_0),.dinb(n1293),.dout(n1296),.clk(gclk));
	jxor g0982(.dina(n1296),.dinb(w_dff_B_fIb3v3qv5_1),.dout(n1297),.clk(gclk));
	jxor g0983(.dina(w_n790_0[1]),.dinb(w_n784_0[0]),.dout(n1298),.clk(gclk));
	jxor g0984(.dina(w_n804_0[0]),.dinb(w_n797_0[1]),.dout(n1299),.clk(gclk));
	jxor g0985(.dina(n1299),.dinb(n1298),.dout(n1300),.clk(gclk));
	jxor g0986(.dina(n1300),.dinb(w_n851_0[0]),.dout(n1301),.clk(gclk));
	jand g0987(.dina(G197),.dinb(w_G18_19[2]),.dout(n1302),.clk(gclk));
	jor g0988(.dina(w_dff_B_QcCZd2tT0_0),.dinb(w_n1205_0[0]),.dout(n1303),.clk(gclk));
	jnot g0989(.din(n1303),.dout(n1304),.clk(gclk));
	jxor g0990(.dina(w_n827_0[0]),.dinb(w_n819_0[0]),.dout(n1305),.clk(gclk));
	jxor g0991(.dina(n1305),.dinb(n1304),.dout(n1306),.clk(gclk));
	jnot g0992(.din(n1306),.dout(n1307),.clk(gclk));
	jxor g0993(.dina(w_n843_0[0]),.dinb(w_n812_0[0]),.dout(n1308),.clk(gclk));
	jxor g0994(.dina(w_dff_B_lXAUZjrw9_0),.dinb(n1307),.dout(n1309),.clk(gclk));
	jand g0995(.dina(w_n1309_0[1]),.dinb(w_n1301_0[1]),.dout(n1310),.clk(gclk));
	jor g0996(.dina(n1310),.dinb(n1297),.dout(n1311),.clk(gclk));
	jand g0997(.dina(G208),.dinb(w_G18_19[1]),.dout(n1312),.clk(gclk));
	jor g0998(.dina(w_dff_B_3u7H70DV1_0),.dinb(w_n1189_0[0]),.dout(n1313),.clk(gclk));
	jxor g0999(.dina(w_n878_0[0]),.dinb(w_n869_0[0]),.dout(n1314),.clk(gclk));
	jxor g1000(.dina(w_n899_0[0]),.dinb(w_n891_0[1]),.dout(n1315),.clk(gclk));
	jxor g1001(.dina(n1315),.dinb(n1314),.dout(n1316),.clk(gclk));
	jxor g1002(.dina(n1316),.dinb(w_dff_B_v0ffNHLM7_1),.dout(n1317),.clk(gclk));
	jnot g1003(.din(w_n916_0[0]),.dout(n1318),.clk(gclk));
	jxor g1004(.dina(w_n945_0[1]),.dinb(w_n927_0[0]),.dout(n1319),.clk(gclk));
	jxor g1005(.dina(n1319),.dinb(n1318),.dout(n1320),.clk(gclk));
	jnot g1006(.din(G198),.dout(n1321),.clk(gclk));
	jor g1007(.dina(n1321),.dinb(w_n355_9[0]),.dout(n1322),.clk(gclk));
	jand g1008(.dina(n1322),.dinb(w_n353_0[0]),.dout(n1323),.clk(gclk));
	jxor g1009(.dina(w_dff_B_N64ZuN0W7_0),.dinb(w_n908_0[0]),.dout(n1324),.clk(gclk));
	jxor g1010(.dina(w_dff_B_Ua5UgG9c8_0),.dinb(n1320),.dout(n1325),.clk(gclk));
	jand g1011(.dina(w_n1325_0[1]),.dinb(w_n1317_0[1]),.dout(n1326),.clk(gclk));
	jnot g1012(.din(w_n1301_0[0]),.dout(n1327),.clk(gclk));
	jnot g1013(.din(w_n1309_0[0]),.dout(n1328),.clk(gclk));
	jand g1014(.dina(n1328),.dinb(w_dff_B_p3lLlLER1_1),.dout(n1329),.clk(gclk));
	jnot g1015(.din(w_n1317_0[0]),.dout(n1330),.clk(gclk));
	jnot g1016(.din(w_n1325_0[0]),.dout(n1331),.clk(gclk));
	jand g1017(.dina(n1331),.dinb(n1330),.dout(n1332),.clk(gclk));
	jor g1018(.dina(n1332),.dinb(n1329),.dout(n1333),.clk(gclk));
	jor g1019(.dina(n1333),.dinb(w_dff_B_yLk5tBE51_1),.dout(n1334),.clk(gclk));
	jor g1020(.dina(n1334),.dinb(w_dff_B_rreQ0XYf0_1),.dout(n1335),.clk(gclk));
	jxor g1021(.dina(w_n744_0[0]),.dinb(w_n730_0[0]),.dout(n1336),.clk(gclk));
	jxor g1022(.dina(n1336),.dinb(w_n737_0[0]),.dout(n1337),.clk(gclk));
	jxor g1023(.dina(w_n754_0[0]),.dinb(w_n723_0[0]),.dout(n1338),.clk(gclk));
	jnot g1024(.din(w_n994_0[0]),.dout(n1339),.clk(gclk));
	jand g1025(.dina(w_n1016_0[0]),.dinb(n1339),.dout(n1340),.clk(gclk));
	jnot g1026(.din(w_n1015_0[0]),.dout(n1341),.clk(gclk));
	jand g1027(.dina(n1341),.dinb(w_n995_0[0]),.dout(n1342),.clk(gclk));
	jor g1028(.dina(n1342),.dinb(n1340),.dout(n1343),.clk(gclk));
	jnot g1029(.din(w_n987_0[0]),.dout(n1344),.clk(gclk));
	jand g1030(.dina(w_n1009_0[1]),.dinb(n1344),.dout(n1345),.clk(gclk));
	jnot g1031(.din(w_n1008_0[0]),.dout(n1346),.clk(gclk));
	jand g1032(.dina(n1346),.dinb(w_n988_0[0]),.dout(n1347),.clk(gclk));
	jor g1033(.dina(n1347),.dinb(n1345),.dout(n1348),.clk(gclk));
	jxor g1034(.dina(n1348),.dinb(n1343),.dout(n1349),.clk(gclk));
	jnot g1035(.din(G181),.dout(n1350),.clk(gclk));
	jor g1036(.dina(n1350),.dinb(w_n355_8[2]),.dout(n1351),.clk(gclk));
	jand g1037(.dina(n1351),.dinb(w_n1166_0[0]),.dout(n1352),.clk(gclk));
	jxor g1038(.dina(w_dff_B_uQvFpwT72_0),.dinb(n1349),.dout(n1353),.clk(gclk));
	jxor g1039(.dina(n1353),.dinb(w_dff_B_LfJWX3D13_1),.dout(n1354),.clk(gclk));
	jxor g1040(.dina(n1354),.dinb(w_dff_B_0ZQfZymY9_1),.dout(n1355),.clk(gclk));
	jor g1041(.dina(w_dff_B_gjvsLsyS4_0),.dinb(n1335),.dout(G416_fa_),.clk(gclk));
	jnot g1042(.din(w_n372_1[0]),.dout(n1357),.clk(gclk));
	jxor g1043(.dina(w_n377_0[1]),.dinb(w_G3717_1[0]),.dout(n1358),.clk(gclk));
	jand g1044(.dina(w_dff_B_P9QBsc5k9_0),.dinb(n1357),.dout(n1359),.clk(gclk));
	jnot g1045(.din(w_n387_0[1]),.dout(n1360),.clk(gclk));
	jxor g1046(.dina(w_n401_0[2]),.dinb(w_G3705_1[1]),.dout(n1361),.clk(gclk));
	jand g1047(.dina(w_n1361_0[1]),.dinb(w_n362_0[1]),.dout(n1362),.clk(gclk));
	jand g1048(.dina(w_n1362_0[1]),.dinb(w_G4526_0[2]),.dout(n1363),.clk(gclk));
	jand g1049(.dina(n1363),.dinb(w_n1360_1[1]),.dout(n1364),.clk(gclk));
	jand g1050(.dina(n1364),.dinb(w_n1359_0[2]),.dout(n1365),.clk(gclk));
	jnot g1051(.din(w_n407_0[1]),.dout(n1366),.clk(gclk));
	jand g1052(.dina(w_n1361_0[0]),.dinb(w_n390_1[0]),.dout(n1367),.clk(gclk));
	jand g1053(.dina(n1367),.dinb(w_n1360_1[0]),.dout(n1368),.clk(gclk));
	jor g1054(.dina(n1368),.dinb(w_dff_B_o9uY41Ac7_1),.dout(n1369),.clk(gclk));
	jand g1055(.dina(n1369),.dinb(w_n1359_0[1]),.dout(n1370),.clk(gclk));
	jnot g1056(.din(w_n413_0[2]),.dout(n1371),.clk(gclk));
	jand g1057(.dina(n1371),.dinb(w_n1359_0[0]),.dout(n1372),.clk(gclk));
	jnot g1058(.din(w_n419_0[0]),.dout(n1373),.clk(gclk));
	jor g1059(.dina(n1373),.dinb(n1372),.dout(n1374),.clk(gclk));
	jor g1060(.dina(n1374),.dinb(n1370),.dout(n1375),.clk(gclk));
	jor g1061(.dina(n1375),.dinb(n1365),.dout(n1376),.clk(gclk));
	jnot g1062(.din(w_n452_0[0]),.dout(n1377),.clk(gclk));
	jand g1063(.dina(w_dff_B_vi9gKCrh7_0),.dinb(w_n1376_0[1]),.dout(n1378),.clk(gclk));
	jnot g1064(.din(w_n464_0[0]),.dout(n1379),.clk(gclk));
	jor g1065(.dina(n1379),.dinb(n1378),.dout(n1380),.clk(gclk));
	jand g1066(.dina(w_n494_0[0]),.dinb(w_n1380_1[1]),.dout(n1381),.clk(gclk));
	jnot g1067(.din(w_n518_0[0]),.dout(n1382),.clk(gclk));
	jor g1068(.dina(n1382),.dinb(n1381),.dout(n1383),.clk(gclk));
	jand g1069(.dina(w_n542_0[0]),.dinb(w_n1383_1[2]),.dout(n1384),.clk(gclk));
	jor g1070(.dina(w_n560_0[0]),.dinb(n1384),.dout(n1385),.clk(gclk));
	jxor g1071(.dina(w_n578_1[0]),.dinb(w_n1385_1[1]),.dout(w_dff_A_k8fwsG6X8_2),.clk(gclk));
	jand g1072(.dina(w_n592_0[0]),.dinb(w_n1385_1[0]),.dout(n1387),.clk(gclk));
	jnot g1073(.din(w_n617_0[0]),.dout(n1388),.clk(gclk));
	jor g1074(.dina(w_dff_B_o9eZOgmS1_0),.dinb(n1387),.dout(n1389),.clk(gclk));
	jand g1075(.dina(w_n637_0[0]),.dinb(w_n1389_1[1]),.dout(n1390),.clk(gclk));
	jnot g1076(.din(w_n656_0[0]),.dout(n1391),.clk(gclk));
	jor g1077(.dina(w_dff_B_vdXXe8U12_0),.dinb(n1390),.dout(n1392),.clk(gclk));
	jxor g1078(.dina(w_n678_0[1]),.dinb(w_n1392_1[1]),.dout(w_dff_A_ouDDPZkR1_2),.clk(gclk));
	jor g1079(.dina(w_n1033_0[0]),.dinb(w_n957_0[0]),.dout(n1394),.clk(gclk));
	jand g1080(.dina(n1394),.dinb(w_n905_0[0]),.dout(n1395),.clk(gclk));
	jor g1081(.dina(n1395),.dinb(w_n1044_0[0]),.dout(n1396),.clk(gclk));
	jand g1082(.dina(n1396),.dinb(w_n864_0[0]),.dout(n1397),.clk(gclk));
	jor g1083(.dina(n1397),.dinb(w_n981_0[0]),.dout(n1398),.clk(gclk));
	jand g1084(.dina(n1398),.dinb(w_n810_0[0]),.dout(n1399),.clk(gclk));
	jor g1085(.dina(n1399),.dinb(w_n972_0[0]),.dout(w_dff_A_y1lICjJJ6_2),.clk(gclk));
	jnot g1086(.din(w_n568_0[1]),.dout(n1401),.clk(gclk));
	jnot g1087(.din(w_n584_0[1]),.dout(n1402),.clk(gclk));
	jnot g1088(.din(w_n589_1[0]),.dout(n1403),.clk(gclk));
	jnot g1089(.din(w_n579_0[1]),.dout(n1404),.clk(gclk));
	jor g1090(.dina(w_n1404_0[1]),.dinb(w_n562_0[1]),.dout(n1405),.clk(gclk));
	jor g1091(.dina(w_n1405_0[1]),.dinb(w_n1403_0[1]),.dout(n1406),.clk(gclk));
	jor g1092(.dina(w_n1406_0[1]),.dinb(w_n1402_0[1]),.dout(n1407),.clk(gclk));
	jand g1093(.dina(n1407),.dinb(w_n615_1[0]),.dout(n1408),.clk(gclk));
	jxor g1094(.dina(n1408),.dinb(w_n1401_0[1]),.dout(w_dff_A_ACqslBCv7_2),.clk(gclk));
	jand g1095(.dina(w_n1406_0[0]),.dinb(w_n613_0[1]),.dout(n1410),.clk(gclk));
	jxor g1096(.dina(n1410),.dinb(w_n1402_0[0]),.dout(w_dff_A_u94kLzpL1_2),.clk(gclk));
	jnot g1097(.din(w_n608_0[1]),.dout(n1412),.clk(gclk));
	jnot g1098(.din(w_n607_0[0]),.dout(n1413),.clk(gclk));
	jand g1099(.dina(n1413),.dinb(w_dff_B_Qst8B18I0_1),.dout(n1414),.clk(gclk));
	jand g1100(.dina(w_n1414_0[1]),.dinb(w_n1405_0[0]),.dout(n1415),.clk(gclk));
	jxor g1101(.dina(n1415),.dinb(w_n1403_0[0]),.dout(w_dff_A_iJCHvIYW2_2),.clk(gclk));
	jand g1102(.dina(w_n578_0[2]),.dinb(w_n1385_0[2]),.dout(n1417),.clk(gclk));
	jor g1103(.dina(n1417),.dinb(w_n606_1[1]),.dout(n1418),.clk(gclk));
	jxor g1104(.dina(n1418),.dinb(w_n573_0[2]),.dout(w_dff_A_IhK2kk8i6_2),.clk(gclk));
	jnot g1105(.din(w_n661_0[0]),.dout(n1420),.clk(gclk));
	jnot g1106(.din(w_n665_0[1]),.dout(n1421),.clk(gclk));
	jnot g1107(.din(w_n669_0[1]),.dout(n1422),.clk(gclk));
	jnot g1108(.din(w_n679_1[0]),.dout(n1423),.clk(gclk));
	jor g1109(.dina(w_dff_B_KHPRBnxK0_0),.dinb(w_n657_1[0]),.dout(n1424),.clk(gclk));
	jor g1110(.dina(w_n1424_0[1]),.dinb(w_n1422_0[1]),.dout(n1425),.clk(gclk));
	jor g1111(.dina(w_n1425_0[1]),.dinb(w_n1421_0[1]),.dout(n1426),.clk(gclk));
	jand g1112(.dina(n1426),.dinb(w_n704_0[0]),.dout(n1427),.clk(gclk));
	jxor g1113(.dina(n1427),.dinb(w_n1420_0[2]),.dout(w_dff_A_IyoCa8wx8_2),.clk(gclk));
	jnot g1114(.din(w_n701_1[0]),.dout(n1429),.clk(gclk));
	jand g1115(.dina(w_n1425_0[0]),.dinb(w_dff_B_wCjmDPvJ6_1),.dout(n1430),.clk(gclk));
	jxor g1116(.dina(n1430),.dinb(w_n1421_0[0]),.dout(w_dff_A_HUfgb5F17_2),.clk(gclk));
	jnot g1117(.din(w_n699_1[0]),.dout(n1432),.clk(gclk));
	jand g1118(.dina(w_n1424_0[0]),.dinb(w_dff_B_nxH7yyo68_1),.dout(n1433),.clk(gclk));
	jxor g1119(.dina(n1433),.dinb(w_n1422_0[0]),.dout(w_dff_A_56MDtBHq7_2),.clk(gclk));
	jand g1120(.dina(w_n678_0[0]),.dinb(w_n1392_1[0]),.dout(n1435),.clk(gclk));
	jor g1121(.dina(n1435),.dinb(w_n697_0[1]),.dout(n1436),.clk(gclk));
	jxor g1122(.dina(n1436),.dinb(w_n674_1[0]),.dout(w_dff_A_bmy2DIyV3_2),.clk(gclk));
	jor g1123(.dina(w_G408_0),.dinb(w_G404_0),.dout(n1438),.clk(gclk));
	jor g1124(.dina(w_G410_0),.dinb(w_G406_0),.dout(n1439),.clk(gclk));
	jor g1125(.dina(n1439),.dinb(n1438),.dout(n1440),.clk(gclk));
	jor g1126(.dina(w_dff_B_pP0s51ua1_0),.dinb(w_G412_0),.dout(n1441),.clk(gclk));
	jor g1127(.dina(w_dff_B_mr5mYk7H5_0),.dinb(w_G416_0),.dout(n1442),.clk(gclk));
	jor g1128(.dina(n1442),.dinb(w_G414_0),.dout(w_dff_A_jhWvCLTd0_2),.clk(gclk));
	jnot g1129(.din(w_n631_0[0]),.dout(n1444),.clk(gclk));
	jnot g1130(.din(w_n627_0[0]),.dout(n1445),.clk(gclk));
	jor g1131(.dina(w_n1445_0[1]),.dinb(w_n618_0[1]),.dout(n1446),.clk(gclk));
	jand g1132(.dina(n1446),.dinb(w_n648_0[1]),.dout(n1447),.clk(gclk));
	jor g1133(.dina(w_n1447_0[1]),.dinb(w_n653_1[0]),.dout(n1448),.clk(gclk));
	jand g1134(.dina(n1448),.dinb(w_n643_0[0]),.dout(n1449),.clk(gclk));
	jxor g1135(.dina(n1449),.dinb(w_n1444_0[2]),.dout(w_dff_A_bXHu9UF51_2),.clk(gclk));
	jnot g1136(.din(w_n635_0[1]),.dout(n1451),.clk(gclk));
	jxor g1137(.dina(w_n1447_0[0]),.dinb(w_dff_B_yo79W8XW9_1),.dout(w_dff_A_kO1eFYA95_2),.clk(gclk));
	jand g1138(.dina(w_n1156_0[0]),.dinb(w_G2239_0[1]),.dout(n1453),.clk(gclk));
	jnot g1139(.din(n1453),.dout(n1454),.clk(gclk));
	jand g1140(.dina(w_n1454_0[1]),.dinb(w_n1389_1[0]),.dout(n1455),.clk(gclk));
	jor g1141(.dina(n1455),.dinb(w_n645_0[1]),.dout(n1456),.clk(gclk));
	jxor g1142(.dina(n1456),.dinb(w_n622_0[2]),.dout(w_dff_A_QNPL4Nn99_2),.clk(gclk));
	jxor g1143(.dina(w_n626_0[0]),.dinb(w_n1389_0[2]),.dout(w_dff_A_GtDw502C2_2),.clk(gclk));
	jxor g1144(.dina(w_n480_1[0]),.dinb(w_n1380_1[0]),.dout(w_dff_A_u2VS0eu85_2),.clk(gclk));
	jnot g1145(.din(w_n714_0[0]),.dout(n1460),.clk(gclk));
	jnot g1146(.din(w_n365_0[0]),.dout(n1461),.clk(gclk));
	jor g1147(.dina(w_n711_0[0]),.dinb(w_n710_0[0]),.dout(n1462),.clk(gclk));
	jxor g1148(.dina(w_dff_B_uHLU5VDr0_0),.dinb(n1461),.dout(n1463),.clk(gclk));
	jnot g1149(.din(w_n1463_0[2]),.dout(n1464),.clk(gclk));
	jor g1150(.dina(w_n1464_0[1]),.dinb(n1460),.dout(n1465),.clk(gclk));
	jand g1151(.dina(w_n1465_0[1]),.dinb(w_n715_0[1]),.dout(w_dff_A_u8189vHk1_2),.clk(gclk));
	jxor g1152(.dina(w_n713_1[0]),.dinb(w_n709_1[0]),.dout(w_dff_A_pN6IxNGh5_2),.clk(gclk));
	jnot g1153(.din(w_n470_0[1]),.dout(n1468),.clk(gclk));
	jnot g1154(.din(w_n486_0[1]),.dout(n1469),.clk(gclk));
	jnot g1155(.din(w_n491_1[0]),.dout(n1470),.clk(gclk));
	jnot g1156(.din(w_n481_0[1]),.dout(n1471),.clk(gclk));
	jor g1157(.dina(w_n1471_0[1]),.dinb(w_n465_0[1]),.dout(n1472),.clk(gclk));
	jor g1158(.dina(w_n1472_0[1]),.dinb(w_n1470_0[1]),.dout(n1473),.clk(gclk));
	jor g1159(.dina(w_n1473_0[1]),.dinb(w_n1469_0[1]),.dout(n1474),.clk(gclk));
	jand g1160(.dina(n1474),.dinb(w_n516_0[1]),.dout(n1475),.clk(gclk));
	jxor g1161(.dina(n1475),.dinb(w_n1468_0[1]),.dout(w_dff_A_Qutbbi7W3_2),.clk(gclk));
	jand g1162(.dina(w_n1473_0[0]),.dinb(w_n514_0[1]),.dout(n1477),.clk(gclk));
	jxor g1163(.dina(n1477),.dinb(w_n1469_0[0]),.dout(w_dff_A_QxgVD2QB2_2),.clk(gclk));
	jand g1164(.dina(w_n508_0[0]),.dinb(w_n510_0[0]),.dout(n1479),.clk(gclk));
	jand g1165(.dina(w_n1479_0[1]),.dinb(w_n1472_0[0]),.dout(n1480),.clk(gclk));
	jxor g1166(.dina(n1480),.dinb(w_n1470_0[0]),.dout(w_dff_A_OEN3E7xB2_2),.clk(gclk));
	jnot g1167(.din(w_n507_1[1]),.dout(n1482),.clk(gclk));
	jand g1168(.dina(w_n480_0[2]),.dinb(w_n1380_0[2]),.dout(n1483),.clk(gclk));
	jor g1169(.dina(n1483),.dinb(w_n1482_0[1]),.dout(n1484),.clk(gclk));
	jxor g1170(.dina(n1484),.dinb(w_n475_0[2]),.dout(w_dff_A_BRr7V1Dd0_2),.clk(gclk));
	jand g1171(.dina(w_n530_0[0]),.dinb(w_n1383_1[1]),.dout(n1486),.clk(gclk));
	jand g1172(.dina(w_n1486_0[1]),.dinb(w_n552_0[0]),.dout(n1487),.clk(gclk));
	jor g1173(.dina(n1487),.dinb(w_n558_0[1]),.dout(n1488),.clk(gclk));
	jxor g1174(.dina(n1488),.dinb(w_n535_1[0]),.dout(w_dff_A_VimgZs4n3_2),.clk(gclk));
	jor g1175(.dina(w_n1486_0[0]),.dinb(w_n556_0[1]),.dout(n1490),.clk(gclk));
	jxor g1176(.dina(n1490),.dinb(w_n540_0[1]),.dout(w_dff_A_djG7tKrZ7_2),.clk(gclk));
	jnot g1177(.din(w_n528_0[1]),.dout(n1492),.clk(gclk));
	jand g1178(.dina(n1492),.dinb(w_G4420_0[1]),.dout(n1493),.clk(gclk));
	jnot g1179(.din(n1493),.dout(n1494),.clk(gclk));
	jand g1180(.dina(w_n1494_0[2]),.dinb(w_n1383_1[0]),.dout(n1495),.clk(gclk));
	jor g1181(.dina(n1495),.dinb(w_n554_0[1]),.dout(n1496),.clk(gclk));
	jxor g1182(.dina(n1496),.dinb(w_n524_1[2]),.dout(w_dff_A_P8hPtzqU4_2),.clk(gclk));
	jxor g1183(.dina(w_n529_0[0]),.dinb(w_n1383_0[2]),.dout(w_dff_A_ypcAw9sg9_2),.clk(gclk));
	jxor g1184(.dina(w_n589_0[2]),.dinb(w_n584_0[0]),.dout(n1499),.clk(gclk));
	jxor g1185(.dina(n1499),.dinb(w_n635_0[0]),.dout(n1500),.clk(gclk));
	jnot g1186(.din(w_n622_0[1]),.dout(n1501),.clk(gclk));
	jnot g1187(.din(w_n653_0[2]),.dout(n1502),.clk(gclk));
	jand g1188(.dina(w_n647_0[0]),.dinb(n1502),.dout(n1503),.clk(gclk));
	jor g1189(.dina(w_dff_B_KoHBeDLk7_0),.dinb(w_n649_0[0]),.dout(n1504),.clk(gclk));
	jxor g1190(.dina(n1504),.dinb(w_n1444_0[1]),.dout(n1505),.clk(gclk));
	jxor g1191(.dina(n1505),.dinb(w_n1501_0[1]),.dout(n1506),.clk(gclk));
	jxor g1192(.dina(n1506),.dinb(w_n1454_0[0]),.dout(n1507),.clk(gclk));
	jand g1193(.dina(w_dff_B_B5qAVPdK2_0),.dinb(w_n618_0[0]),.dout(n1508),.clk(gclk));
	jxor g1194(.dina(w_n645_0[0]),.dinb(w_n1501_0[0]),.dout(n1509),.clk(gclk));
	jand g1195(.dina(w_n648_0[0]),.dinb(w_n1445_0[0]),.dout(n1510),.clk(gclk));
	jnot g1196(.din(w_n1510_0[1]),.dout(n1511),.clk(gclk));
	jor g1197(.dina(n1511),.dinb(w_n642_0[0]),.dout(n1512),.clk(gclk));
	jor g1198(.dina(w_n1510_0[0]),.dinb(w_n653_0[1]),.dout(n1513),.clk(gclk));
	jand g1199(.dina(w_dff_B_WfMAqJW37_0),.dinb(n1512),.dout(n1514),.clk(gclk));
	jxor g1200(.dina(n1514),.dinb(w_n1444_0[0]),.dout(n1515),.clk(gclk));
	jxor g1201(.dina(n1515),.dinb(w_dff_B_jMIpVqyN4_1),.dout(n1516),.clk(gclk));
	jand g1202(.dina(w_dff_B_qRoOA2Qd9_0),.dinb(w_n1389_0[1]),.dout(n1517),.clk(gclk));
	jor g1203(.dina(n1517),.dinb(n1508),.dout(n1518),.clk(gclk));
	jand g1204(.dina(w_n613_0[0]),.dinb(w_n606_1[0]),.dout(n1519),.clk(gclk));
	jnot g1205(.din(w_n606_0[2]),.dout(n1520),.clk(gclk));
	jand g1206(.dina(w_n605_0[0]),.dinb(w_n1520_0[1]),.dout(n1521),.clk(gclk));
	jand g1207(.dina(n1521),.dinb(w_n610_0[0]),.dout(n1522),.clk(gclk));
	jxor g1208(.dina(n1522),.dinb(w_n578_0[1]),.dout(n1523),.clk(gclk));
	jor g1209(.dina(n1523),.dinb(n1519),.dout(n1524),.clk(gclk));
	jor g1210(.dina(w_n572_0[1]),.dinb(w_n569_0[0]),.dout(n1525),.clk(gclk));
	jand g1211(.dina(w_n1520_0[0]),.dinb(w_dff_B_WS9Io77u8_1),.dout(n1526),.clk(gclk));
	jor g1212(.dina(n1526),.dinb(w_n608_0[0]),.dout(n1527),.clk(gclk));
	jxor g1213(.dina(w_dff_B_h1hNkmOI9_0),.dinb(w_n615_0[2]),.dout(n1528),.clk(gclk));
	jxor g1214(.dina(n1528),.dinb(w_n1401_0[0]),.dout(n1529),.clk(gclk));
	jxor g1215(.dina(n1529),.dinb(w_dff_B_INRxn0Zf8_1),.dout(n1530),.clk(gclk));
	jor g1216(.dina(w_dff_B_nHV2rcZB0_0),.dinb(w_n1385_0[1]),.dout(n1531),.clk(gclk));
	jand g1217(.dina(w_n1414_0[0]),.dinb(w_n1404_0[0]),.dout(n1532),.clk(gclk));
	jxor g1218(.dina(n1532),.dinb(w_n568_0[0]),.dout(n1533),.clk(gclk));
	jxor g1219(.dina(w_n606_0[1]),.dinb(w_n573_0[1]),.dout(n1534),.clk(gclk));
	jand g1220(.dina(w_n589_0[1]),.dinb(w_n579_0[0]),.dout(n1535),.clk(gclk));
	jor g1221(.dina(w_dff_B_xVxqDQz99_0),.dinb(w_n612_0[0]),.dout(n1536),.clk(gclk));
	jnot g1222(.din(w_n1536_0[1]),.dout(n1537),.clk(gclk));
	jand g1223(.dina(n1537),.dinb(w_n599_0[0]),.dout(n1538),.clk(gclk));
	jnot g1224(.din(w_n591_0[0]),.dout(n1539),.clk(gclk));
	jand g1225(.dina(w_n1536_0[0]),.dinb(w_dff_B_Nh6WyFZo2_1),.dout(n1540),.clk(gclk));
	jand g1226(.dina(w_dff_B_aeoxuii34_0),.dinb(w_n615_0[1]),.dout(n1541),.clk(gclk));
	jor g1227(.dina(n1541),.dinb(w_dff_B_X1okK80g2_1),.dout(n1542),.clk(gclk));
	jxor g1228(.dina(n1542),.dinb(w_dff_B_PYhRQtCE6_1),.dout(n1543),.clk(gclk));
	jxor g1229(.dina(n1543),.dinb(w_dff_B_aI1HuN814_1),.dout(n1544),.clk(gclk));
	jor g1230(.dina(w_dff_B_QTp7Gtxt6_0),.dinb(w_n562_0[0]),.dout(n1545),.clk(gclk));
	jand g1231(.dina(n1545),.dinb(n1531),.dout(n1546),.clk(gclk));
	jxor g1232(.dina(w_dff_B_gnBCZDhH4_0),.dinb(n1518),.dout(n1547),.clk(gclk));
	jxor g1233(.dina(n1547),.dinb(w_dff_B_U8EmEL2h4_1),.dout(w_dff_A_O0ichDPW1_2),.clk(gclk));
	jand g1234(.dina(w_n713_0[2]),.dinb(w_n709_0[2]),.dout(n1549),.clk(gclk));
	jor g1235(.dina(n1549),.dinb(w_n1463_0[1]),.dout(n1550),.clk(gclk));
	jnot g1236(.din(w_n683_0[0]),.dout(n1551),.clk(gclk));
	jand g1237(.dina(w_n707_0[1]),.dinb(w_n1392_0[2]),.dout(n1552),.clk(gclk));
	jand g1238(.dina(w_n712_0[0]),.dinb(w_n708_0[0]),.dout(n1553),.clk(gclk));
	jor g1239(.dina(n1553),.dinb(w_n1464_0[0]),.dout(n1554),.clk(gclk));
	jor g1240(.dina(w_dff_B_pBDQt7Fm1_0),.dinb(n1552),.dout(n1555),.clk(gclk));
	jor g1241(.dina(n1555),.dinb(n1551),.dout(n1556),.clk(gclk));
	jand g1242(.dina(w_dff_B_M7sTA4wo4_0),.dinb(n1550),.dout(n1557),.clk(gclk));
	jand g1243(.dina(w_n1463_0[0]),.dinb(w_n707_0[0]),.dout(n1558),.clk(gclk));
	jand g1244(.dina(w_dff_B_xS7EoXhY9_0),.dinb(w_n657_0[2]),.dout(n1559),.clk(gclk));
	jor g1245(.dina(w_dff_B_PI4UAjCe7_0),.dinb(n1557),.dout(n1560),.clk(gclk));
	jxor g1246(.dina(w_n669_0[0]),.dinb(w_n665_0[0]),.dout(n1561),.clk(gclk));
	jor g1247(.dina(w_n701_0[2]),.dinb(w_n686_0[0]),.dout(n1562),.clk(gclk));
	jand g1248(.dina(w_dff_B_XZZm6ftf0_0),.dinb(w_n703_0[0]),.dout(n1563),.clk(gclk));
	jxor g1249(.dina(n1563),.dinb(w_n1420_0[1]),.dout(n1564),.clk(gclk));
	jor g1250(.dina(w_n677_0[0]),.dinb(w_n675_0[0]),.dout(n1565),.clk(gclk));
	jxor g1251(.dina(n1565),.dinb(w_n674_0[2]),.dout(n1566),.clk(gclk));
	jxor g1252(.dina(w_dff_B_zxuyijCv3_0),.dinb(w_n699_0[2]),.dout(n1567),.clk(gclk));
	jxor g1253(.dina(w_dff_B_qqXNUt202_0),.dinb(n1564),.dout(n1568),.clk(gclk));
	jand g1254(.dina(w_dff_B_d7qp4tb85_0),.dinb(w_n657_0[1]),.dout(n1569),.clk(gclk));
	jand g1255(.dina(w_n679_0[2]),.dinb(w_n692_0[0]),.dout(n1570),.clk(gclk));
	jor g1256(.dina(w_dff_B_gtqeDLaA1_0),.dinb(w_n701_0[1]),.dout(n1571),.clk(gclk));
	jor g1257(.dina(w_n1571_0[1]),.dinb(w_n687_0[0]),.dout(n1572),.clk(gclk));
	jnot g1258(.din(w_n1571_0[0]),.dout(n1573),.clk(gclk));
	jor g1259(.dina(n1573),.dinb(w_n680_0[0]),.dout(n1574),.clk(gclk));
	jor g1260(.dina(w_dff_B_Jdd7TguC6_0),.dinb(w_n705_0[0]),.dout(n1575),.clk(gclk));
	jand g1261(.dina(n1575),.dinb(w_dff_B_AQXSGaOY9_1),.dout(n1576),.clk(gclk));
	jor g1262(.dina(w_n699_0[1]),.dinb(w_n679_0[1]),.dout(n1577),.clk(gclk));
	jxor g1263(.dina(n1577),.dinb(w_n1420_0[0]),.dout(n1578),.clk(gclk));
	jxor g1264(.dina(w_dff_B_E5nqfP4x2_0),.dinb(n1576),.dout(n1579),.clk(gclk));
	jxor g1265(.dina(n1579),.dinb(w_n697_0[0]),.dout(n1580),.clk(gclk));
	jxor g1266(.dina(n1580),.dinb(w_n674_0[1]),.dout(n1581),.clk(gclk));
	jand g1267(.dina(w_dff_B_7FIOKbKe8_0),.dinb(w_n1392_0[1]),.dout(n1582),.clk(gclk));
	jor g1268(.dina(n1582),.dinb(n1569),.dout(n1583),.clk(gclk));
	jxor g1269(.dina(n1583),.dinb(w_dff_B_8qb9JnrM6_1),.dout(n1584),.clk(gclk));
	jxor g1270(.dina(w_dff_B_YLdHd6tD0_0),.dinb(n1560),.dout(G338),.clk(gclk));
	jxor g1271(.dina(w_n491_0[2]),.dinb(w_n486_0[0]),.dout(n1586),.clk(gclk));
	jxor g1272(.dina(n1586),.dinb(w_n540_0[0]),.dout(n1587),.clk(gclk));
	jnot g1273(.din(w_n535_0[2]),.dout(n1588),.clk(gclk));
	jnot g1274(.din(w_n557_0[0]),.dout(n1589),.clk(gclk));
	jor g1275(.dina(w_n556_0[0]),.dinb(w_n549_0[0]),.dout(n1590),.clk(gclk));
	jand g1276(.dina(w_dff_B_2DsdV5O88_0),.dinb(n1589),.dout(n1591),.clk(gclk));
	jxor g1277(.dina(n1591),.dinb(w_dff_B_mm7fPUEe4_1),.dout(n1592),.clk(gclk));
	jxor g1278(.dina(w_n1494_0[1]),.dinb(w_n524_1[1]),.dout(n1593),.clk(gclk));
	jxor g1279(.dina(w_dff_B_XX9PT8uf5_0),.dinb(n1592),.dout(n1594),.clk(gclk));
	jand g1280(.dina(w_dff_B_VkEavW1t2_0),.dinb(w_n519_0[0]),.dout(n1595),.clk(gclk));
	jxor g1281(.dina(w_n554_0[0]),.dinb(w_n524_1[0]),.dout(n1596),.clk(gclk));
	jxor g1282(.dina(n1596),.dinb(w_n535_0[1]),.dout(n1597),.clk(gclk));
	jand g1283(.dina(w_n1494_0[0]),.dinb(w_n524_0[2]),.dout(n1598),.clk(gclk));
	jor g1284(.dina(n1598),.dinb(w_n553_0[0]),.dout(n1599),.clk(gclk));
	jnot g1285(.din(w_n1599_0[1]),.dout(n1600),.clk(gclk));
	jand g1286(.dina(n1600),.dinb(w_n558_0[0]),.dout(n1601),.clk(gclk));
	jand g1287(.dina(w_n1599_0[0]),.dinb(w_n551_0[0]),.dout(n1602),.clk(gclk));
	jor g1288(.dina(w_dff_B_sel0X8RR9_0),.dinb(n1601),.dout(n1603),.clk(gclk));
	jxor g1289(.dina(n1603),.dinb(w_dff_B_1DOt81Ad4_1),.dout(n1604),.clk(gclk));
	jand g1290(.dina(w_dff_B_EjHF14WT6_0),.dinb(w_n1383_0[1]),.dout(n1605),.clk(gclk));
	jor g1291(.dina(n1605),.dinb(n1595),.dout(n1606),.clk(gclk));
	jor g1292(.dina(w_n474_0[1]),.dinb(w_n471_0[0]),.dout(n1607),.clk(gclk));
	jand g1293(.dina(w_n507_1[0]),.dinb(w_dff_B_4ORWPjYZ0_1),.dout(n1608),.clk(gclk));
	jor g1294(.dina(n1608),.dinb(w_n509_0[0]),.dout(n1609),.clk(gclk));
	jnot g1295(.din(w_n516_0[0]),.dout(n1610),.clk(gclk));
	jnot g1296(.din(w_n514_0[0]),.dout(n1611),.clk(gclk));
	jor g1297(.dina(w_n1611_0[1]),.dinb(w_n507_0[2]),.dout(n1612),.clk(gclk));
	jor g1298(.dina(w_n505_0[0]),.dinb(w_n1482_0[0]),.dout(n1613),.clk(gclk));
	jor g1299(.dina(n1613),.dinb(w_n512_0[0]),.dout(n1614),.clk(gclk));
	jxor g1300(.dina(n1614),.dinb(w_n480_0[1]),.dout(n1615),.clk(gclk));
	jand g1301(.dina(w_dff_B_XKqHvp1z8_0),.dinb(n1612),.dout(n1616),.clk(gclk));
	jxor g1302(.dina(n1616),.dinb(w_n1468_0[0]),.dout(n1617),.clk(gclk));
	jxor g1303(.dina(n1617),.dinb(w_n1610_0[1]),.dout(n1618),.clk(gclk));
	jxor g1304(.dina(n1618),.dinb(w_dff_B_2yNwb2Rz4_1),.dout(n1619),.clk(gclk));
	jor g1305(.dina(n1619),.dinb(w_n1380_0[1]),.dout(n1620),.clk(gclk));
	jand g1306(.dina(w_n1479_0[0]),.dinb(w_n1471_0[0]),.dout(n1621),.clk(gclk));
	jxor g1307(.dina(n1621),.dinb(w_n470_0[0]),.dout(n1622),.clk(gclk));
	jxor g1308(.dina(w_n507_0[1]),.dinb(w_n475_0[1]),.dout(n1623),.clk(gclk));
	jand g1309(.dina(w_n491_0[1]),.dinb(w_n481_0[0]),.dout(n1624),.clk(gclk));
	jor g1310(.dina(w_dff_B_4stDTBS90_0),.dinb(w_n1611_0[0]),.dout(n1625),.clk(gclk));
	jor g1311(.dina(w_n1625_0[1]),.dinb(w_n502_0[0]),.dout(n1626),.clk(gclk));
	jnot g1312(.din(w_n1625_0[0]),.dout(n1627),.clk(gclk));
	jor g1313(.dina(n1627),.dinb(w_n493_0[0]),.dout(n1628),.clk(gclk));
	jor g1314(.dina(n1628),.dinb(w_n1610_0[0]),.dout(n1629),.clk(gclk));
	jand g1315(.dina(n1629),.dinb(w_dff_B_nGaZYB9h6_1),.dout(n1630),.clk(gclk));
	jxor g1316(.dina(n1630),.dinb(w_dff_B_lxx2CanO3_1),.dout(n1631),.clk(gclk));
	jxor g1317(.dina(n1631),.dinb(w_dff_B_79HMWNLb4_1),.dout(n1632),.clk(gclk));
	jor g1318(.dina(n1632),.dinb(w_n465_0[0]),.dout(n1633),.clk(gclk));
	jand g1319(.dina(n1633),.dinb(w_dff_B_tP5QGGy90_1),.dout(n1634),.clk(gclk));
	jxor g1320(.dina(n1634),.dinb(w_dff_B_xMBW8gtM9_1),.dout(n1635),.clk(gclk));
	jxor g1321(.dina(n1635),.dinb(w_dff_B_ASHbUCWz7_1),.dout(w_dff_A_p7vnaGTp4_2),.clk(gclk));
	jxor g1322(.dina(w_n450_0[0]),.dinb(w_n1360_0[2]),.dout(n1637),.clk(gclk));
	jnot g1323(.din(w_n455_0[0]),.dout(n1638),.clk(gclk));
	jnot g1324(.din(w_n460_0[0]),.dout(n1639),.clk(gclk));
	jor g1325(.dina(n1639),.dinb(w_dff_B_8HgM9npp3_1),.dout(n1640),.clk(gclk));
	jand g1326(.dina(n1640),.dinb(w_n461_0[0]),.dout(n1641),.clk(gclk));
	jxor g1327(.dina(n1641),.dinb(w_n446_0[2]),.dout(n1642),.clk(gclk));
	jnot g1328(.din(w_n1642_0[1]),.dout(n1643),.clk(gclk));
	jxor g1329(.dina(w_n1148_0[1]),.dinb(w_n429_1[1]),.dout(n1644),.clk(gclk));
	jnot g1330(.din(w_n1644_0[1]),.dout(n1645),.clk(gclk));
	jor g1331(.dina(w_dff_B_XYYkBOti0_0),.dinb(n1643),.dout(n1646),.clk(gclk));
	jor g1332(.dina(w_n1644_0[0]),.dinb(w_n1642_0[0]),.dout(n1647),.clk(gclk));
	jand g1333(.dina(n1647),.dinb(w_n422_0[1]),.dout(n1648),.clk(gclk));
	jand g1334(.dina(n1648),.dinb(n1646),.dout(n1649),.clk(gclk));
	jxor g1335(.dina(w_n458_0[0]),.dinb(w_n429_1[0]),.dout(n1650),.clk(gclk));
	jxor g1336(.dina(w_dff_B_KeNprzu58_0),.dinb(w_n446_0[1]),.dout(n1651),.clk(gclk));
	jnot g1337(.din(w_n462_0[0]),.dout(n1652),.clk(gclk));
	jor g1338(.dina(w_n1148_0[0]),.dinb(w_n429_0[2]),.dout(n1653),.clk(gclk));
	jand g1339(.dina(n1653),.dinb(w_n457_0[0]),.dout(n1654),.clk(gclk));
	jand g1340(.dina(w_n1654_0[1]),.dinb(n1652),.dout(n1655),.clk(gclk));
	jnot g1341(.din(n1655),.dout(n1656),.clk(gclk));
	jnot g1342(.din(w_n456_0[0]),.dout(n1657),.clk(gclk));
	jor g1343(.dina(w_n1654_0[0]),.dinb(n1657),.dout(n1658),.clk(gclk));
	jand g1344(.dina(w_dff_B_iWkXe2AJ4_0),.dinb(n1656),.dout(n1659),.clk(gclk));
	jor g1345(.dina(w_n1659_0[1]),.dinb(w_n1651_0[1]),.dout(n1660),.clk(gclk));
	jnot g1346(.din(w_n1651_0[0]),.dout(n1661),.clk(gclk));
	jnot g1347(.din(w_n1659_0[0]),.dout(n1662),.clk(gclk));
	jor g1348(.dina(n1662),.dinb(w_dff_B_lbznyI1u1_1),.dout(n1663),.clk(gclk));
	jand g1349(.dina(n1663),.dinb(w_n1376_0[0]),.dout(n1664),.clk(gclk));
	jand g1350(.dina(n1664),.dinb(w_dff_B_j4SVgvbl0_1),.dout(n1665),.clk(gclk));
	jor g1351(.dina(n1665),.dinb(w_dff_B_JRcaNep85_1),.dout(n1666),.clk(gclk));
	jand g1352(.dina(w_n1136_0[0]),.dinb(w_n403_0[0]),.dout(n1667),.clk(gclk));
	jnot g1353(.din(w_n1667_0[1]),.dout(n1668),.clk(gclk));
	jor g1354(.dina(n1668),.dinb(w_n1128_0[2]),.dout(n1669),.clk(gclk));
	jnot g1355(.din(w_n1128_0[1]),.dout(n1670),.clk(gclk));
	jand g1356(.dina(w_n1362_0[0]),.dinb(w_n1360_0[1]),.dout(n1671),.clk(gclk));
	jor g1357(.dina(w_dff_B_jxRLmfFY1_0),.dinb(w_n1670_0[1]),.dout(n1672),.clk(gclk));
	jor g1358(.dina(w_n1672_0[1]),.dinb(w_n1667_0[0]),.dout(n1673),.clk(gclk));
	jand g1359(.dina(n1673),.dinb(w_dff_B_REeW9gvT5_1),.dout(n1674),.clk(gclk));
	jxor g1360(.dina(n1674),.dinb(w_n372_0[2]),.dout(n1675),.clk(gclk));
	jnot g1361(.din(w_n1672_0[0]),.dout(n1676),.clk(gclk));
	jor g1362(.dina(n1676),.dinb(w_n1127_0[0]),.dout(n1677),.clk(gclk));
	jand g1363(.dina(n1677),.dinb(w_n417_0[0]),.dout(n1678),.clk(gclk));
	jxor g1364(.dina(n1678),.dinb(w_n402_0[1]),.dout(n1679),.clk(gclk));
	jxor g1365(.dina(n1679),.dinb(w_n354_0[2]),.dout(n1680),.clk(gclk));
	jnot g1366(.din(w_n1680_0[1]),.dout(n1681),.clk(gclk));
	jand g1367(.dina(n1681),.dinb(w_n1675_0[1]),.dout(n1682),.clk(gclk));
	jnot g1368(.din(w_n1675_0[0]),.dout(n1683),.clk(gclk));
	jand g1369(.dina(w_n1680_0[0]),.dinb(w_dff_B_yaGAndz76_1),.dout(n1684),.clk(gclk));
	jor g1370(.dina(n1684),.dinb(w_n388_0[0]),.dout(n1685),.clk(gclk));
	jor g1371(.dina(n1685),.dinb(n1682),.dout(n1686),.clk(gclk));
	jxor g1372(.dina(w_n1130_0[0]),.dinb(w_n372_0[1]),.dout(n1687),.clk(gclk));
	jand g1373(.dina(w_n407_0[0]),.dinb(w_n354_0[1]),.dout(n1688),.clk(gclk));
	jand g1374(.dina(n1688),.dinb(w_n413_0[1]),.dout(n1689),.clk(gclk));
	jand g1375(.dina(w_n1689_0[1]),.dinb(w_n395_0[0]),.dout(n1690),.clk(gclk));
	jnot g1376(.din(w_n1689_0[0]),.dout(n1691),.clk(gclk));
	jand g1377(.dina(w_n1670_0[0]),.dinb(w_n390_0[2]),.dout(n1692),.clk(gclk));
	jor g1378(.dina(n1692),.dinb(w_n362_0[0]),.dout(n1693),.clk(gclk));
	jand g1379(.dina(n1693),.dinb(w_dff_B_BaY2riKL9_1),.dout(n1694),.clk(gclk));
	jor g1380(.dina(n1694),.dinb(w_dff_B_FuQFIgH88_1),.dout(n1695),.clk(gclk));
	jand g1381(.dina(w_n401_0[1]),.dinb(w_G3705_1[0]),.dout(n1696),.clk(gclk));
	jor g1382(.dina(n1696),.dinb(w_n390_0[1]),.dout(n1697),.clk(gclk));
	jand g1383(.dina(n1697),.dinb(w_n412_0[0]),.dout(n1698),.clk(gclk));
	jxor g1384(.dina(w_dff_B_tUAfxP7n4_0),.dinb(n1695),.dout(n1699),.clk(gclk));
	jnot g1385(.din(w_n1699_0[1]),.dout(n1700),.clk(gclk));
	jand g1386(.dina(n1700),.dinb(w_n1687_0[1]),.dout(n1701),.clk(gclk));
	jnot g1387(.din(w_n1687_0[0]),.dout(n1702),.clk(gclk));
	jand g1388(.dina(w_n1699_0[0]),.dinb(w_dff_B_FqaGOYoO0_1),.dout(n1703),.clk(gclk));
	jor g1389(.dina(n1703),.dinb(w_G4526_0[1]),.dout(n1704),.clk(gclk));
	jor g1390(.dina(n1704),.dinb(n1701),.dout(n1705),.clk(gclk));
	jand g1391(.dina(w_dff_B_cC0B5eQI6_0),.dinb(n1686),.dout(n1706),.clk(gclk));
	jxor g1392(.dina(n1706),.dinb(w_n379_0[1]),.dout(n1707),.clk(gclk));
	jxor g1393(.dina(n1707),.dinb(w_dff_B_LqYwp0DK4_1),.dout(n1708),.clk(gclk));
	jxor g1394(.dina(n1708),.dinb(w_dff_B_3LGbg9YE5_1),.dout(w_dff_A_neBD5Ml89_2),.clk(gclk));
	jdff g1395(.din(w_G1_1[1]),.dout(w_dff_A_Lj9zbcUa6_1),.clk(gclk));
	jdff g1396(.din(w_G1_1[0]),.dout(w_dff_A_bKUyBodi8_1),.clk(gclk));
	jdff g1397(.din(w_G1459_0[0]),.dout(w_dff_A_ykkR7BTX5_1),.clk(gclk));
	jdff g1398(.din(w_G1469_0[1]),.dout(w_dff_A_5BZl4JPk1_1),.clk(gclk));
	jdff g1399(.din(w_G1480_0[0]),.dout(w_dff_A_lpzyHoCB3_1),.clk(gclk));
	jdff g1400(.din(w_G1486_0[0]),.dout(w_dff_A_rEh14yc44_1),.clk(gclk));
	jdff g1401(.din(w_G1492_0[1]),.dout(w_dff_A_Qb2jOS5o0_1),.clk(gclk));
	jdff g1402(.din(w_G1496_0[0]),.dout(w_dff_A_lmpG2qDt1_1),.clk(gclk));
	jdff g1403(.din(w_G2208_0[0]),.dout(w_dff_A_6XQh2fku4_1),.clk(gclk));
	jdff g1404(.din(w_G2218_0[0]),.dout(w_dff_A_hlgqtfXa0_1),.clk(gclk));
	jdff g1405(.din(w_G2224_0[1]),.dout(w_dff_A_k7VluDx66_1),.clk(gclk));
	jdff g1406(.din(w_G2230_0[1]),.dout(w_dff_A_f0loBwmj7_1),.clk(gclk));
	jdff g1407(.din(w_G2236_0[1]),.dout(w_dff_A_KZTb2yWC7_1),.clk(gclk));
	jdff g1408(.din(w_G2239_0[0]),.dout(w_dff_A_QLfkh51b8_1),.clk(gclk));
	jdff g1409(.din(w_G2247_0[0]),.dout(w_dff_A_OfURwhBQ4_1),.clk(gclk));
	jdff g1410(.din(w_G2253_0[1]),.dout(w_dff_A_fIekaECE3_1),.clk(gclk));
	jdff g1411(.din(w_G2256_0[1]),.dout(w_dff_A_gOv57F6o7_1),.clk(gclk));
	jdff g1412(.din(w_G3698_0[0]),.dout(w_dff_A_11QQyRH85_1),.clk(gclk));
	jdff g1413(.din(w_G3701_0[1]),.dout(w_dff_A_9okMP1UV2_1),.clk(gclk));
	jdff g1414(.din(w_G3705_0[2]),.dout(w_dff_A_XMLPmksm8_1),.clk(gclk));
	jdff g1415(.din(w_G3711_0[1]),.dout(w_dff_A_RwGKFHG76_1),.clk(gclk));
	jdff g1416(.din(w_G3717_0[2]),.dout(w_dff_A_o7j95bj09_1),.clk(gclk));
	jdff g1417(.din(w_G3723_0[1]),.dout(w_dff_A_SwcSZ5mu2_1),.clk(gclk));
	jdff g1418(.din(w_G3729_0[1]),.dout(w_dff_A_UOFpF7hR0_1),.clk(gclk));
	jdff g1419(.din(w_G3737_0[1]),.dout(w_dff_A_3rAom8zd6_1),.clk(gclk));
	jdff g1420(.din(w_G3743_0[1]),.dout(w_dff_A_jC7At71Q2_1),.clk(gclk));
	jdff g1421(.din(w_G3749_0[1]),.dout(w_dff_A_O7RMNuf06_1),.clk(gclk));
	jdff g1422(.din(w_G4393_0[0]),.dout(w_dff_A_cykvuITa8_1),.clk(gclk));
	jdff g1423(.din(w_G4400_0[0]),.dout(w_dff_A_ZmdyHmdd8_1),.clk(gclk));
	jdff g1424(.din(w_G4405_0[1]),.dout(w_dff_A_bVT2Wp258_1),.clk(gclk));
	jdff g1425(.din(w_G4410_0[1]),.dout(w_dff_A_1ISwIh973_1),.clk(gclk));
	jdff g1426(.din(w_G4415_0[1]),.dout(w_dff_A_uyVV29G02_1),.clk(gclk));
	jdff g1427(.din(w_G4420_0[0]),.dout(w_dff_A_paBQc1dR5_1),.clk(gclk));
	jdff g1428(.din(w_G4427_0[0]),.dout(w_dff_A_BhtDhst74_1),.clk(gclk));
	jdff g1429(.din(w_G4432_0[1]),.dout(w_dff_A_xoVdo85w5_1),.clk(gclk));
	jdff g1430(.din(w_G4437_0[0]),.dout(w_dff_A_7CNN2QGj1_1),.clk(gclk));
	jdff g1431(.din(w_G1462_0[0]),.dout(w_dff_A_vzwKrL7w6_1),.clk(gclk));
	jdff g1432(.din(w_G2211_0[0]),.dout(w_dff_A_FaNycJh43_1),.clk(gclk));
	jdff g1433(.din(w_G4394_0[1]),.dout(w_dff_A_brqg9SVn2_1),.clk(gclk));
	jdff g1434(.din(w_G1_0[2]),.dout(w_dff_A_72jiinuu9_1),.clk(gclk));
	jdff g1435(.din(w_G106_0[1]),.dout(w_dff_A_VcYMcl4d4_1),.clk(gclk));
	jnot g1436(.din(w_G15_0[1]),.dout(w_dff_A_X70tw3Lb1_1),.clk(gclk));
	jor g1437(.dina(w_n345_0[0]),.dinb(w_G5_0[2]),.dout(w_dff_A_B1dnqkxZ4_2),.clk(gclk));
	jnot g1438(.din(w_G15_0[0]),.dout(w_dff_A_w5MdrG526_1),.clk(gclk));
	jor g1439(.dina(w_n349_0[0]),.dinb(w_G5_0[1]),.dout(w_dff_A_KrEOdKkt7_2),.clk(gclk));
	jdff g1440(.din(w_G1_0[1]),.dout(w_dff_A_WfeN12RN7_1),.clk(gclk));
	jand g1441(.dina(w_n1125_0[1]),.dinb(w_n1122_0[1]),.dout(w_dff_A_A5XS2GlF0_2),.clk(gclk));
	jor g1442(.dina(w_n720_1[0]),.dinb(w_n716_1[0]),.dout(w_dff_A_nl5Rctji5_2),.clk(gclk));
	jand g1443(.dina(w_n1125_0[0]),.dinb(w_n1122_0[0]),.dout(w_dff_A_hMJWlTAb8_2),.clk(gclk));
	jor g1444(.dina(w_n720_0[2]),.dinb(w_n716_0[2]),.dout(w_dff_A_kfLFkw6M5_2),.clk(gclk));
	jor g1445(.dina(w_n720_0[1]),.dinb(w_n716_0[1]),.dout(w_dff_A_FoWZznBm6_2),.clk(gclk));
	jand g1446(.dina(w_n1465_0[0]),.dinb(w_n715_0[0]),.dout(w_dff_A_KJykaV3M0_2),.clk(gclk));
	jxor g1447(.dina(w_n713_0[1]),.dinb(w_n709_0[1]),.dout(w_dff_A_E8jalRTs2_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G5_0(.douta(w_G5_0[0]),.doutb(w_dff_A_Csyy1rkH6_1),.doutc(w_dff_A_FaHfh2fO1_2),.din(G5));
	jspl3 jspl3_w_G5_1(.douta(w_dff_A_LJ5eExnU7_0),.doutb(w_dff_A_2Rxoc2Fc8_1),.doutc(w_G5_1[2]),.din(w_G5_0[0]));
	jspl3 jspl3_w_G15_0(.douta(w_G15_0[0]),.doutb(w_G15_0[1]),.doutc(w_G15_0[2]),.din(G15));
	jspl3 jspl3_w_G18_0(.douta(w_G18_0[0]),.doutb(w_G18_0[1]),.doutc(w_G18_0[2]),.din(G18));
	jspl3 jspl3_w_G18_1(.douta(w_G18_1[0]),.doutb(w_G18_1[1]),.doutc(w_G18_1[2]),.din(w_G18_0[0]));
	jspl3 jspl3_w_G18_2(.douta(w_G18_2[0]),.doutb(w_G18_2[1]),.doutc(w_G18_2[2]),.din(w_G18_0[1]));
	jspl3 jspl3_w_G18_3(.douta(w_G18_3[0]),.doutb(w_G18_3[1]),.doutc(w_G18_3[2]),.din(w_G18_0[2]));
	jspl3 jspl3_w_G18_4(.douta(w_G18_4[0]),.doutb(w_G18_4[1]),.doutc(w_G18_4[2]),.din(w_G18_1[0]));
	jspl3 jspl3_w_G18_5(.douta(w_G18_5[0]),.doutb(w_G18_5[1]),.doutc(w_G18_5[2]),.din(w_G18_1[1]));
	jspl3 jspl3_w_G18_6(.douta(w_G18_6[0]),.doutb(w_dff_A_cXHyq6OK4_1),.doutc(w_dff_A_984qphLh4_2),.din(w_G18_1[2]));
	jspl3 jspl3_w_G18_7(.douta(w_G18_7[0]),.doutb(w_G18_7[1]),.doutc(w_G18_7[2]),.din(w_G18_2[0]));
	jspl3 jspl3_w_G18_8(.douta(w_G18_8[0]),.doutb(w_G18_8[1]),.doutc(w_G18_8[2]),.din(w_G18_2[1]));
	jspl3 jspl3_w_G18_9(.douta(w_G18_9[0]),.doutb(w_G18_9[1]),.doutc(w_G18_9[2]),.din(w_G18_2[2]));
	jspl3 jspl3_w_G18_10(.douta(w_G18_10[0]),.doutb(w_G18_10[1]),.doutc(w_G18_10[2]),.din(w_G18_3[0]));
	jspl3 jspl3_w_G18_11(.douta(w_G18_11[0]),.doutb(w_G18_11[1]),.doutc(w_G18_11[2]),.din(w_G18_3[1]));
	jspl3 jspl3_w_G18_12(.douta(w_G18_12[0]),.doutb(w_G18_12[1]),.doutc(w_G18_12[2]),.din(w_G18_3[2]));
	jspl3 jspl3_w_G18_13(.douta(w_G18_13[0]),.doutb(w_G18_13[1]),.doutc(w_G18_13[2]),.din(w_G18_4[0]));
	jspl3 jspl3_w_G18_14(.douta(w_G18_14[0]),.doutb(w_G18_14[1]),.doutc(w_G18_14[2]),.din(w_G18_4[1]));
	jspl3 jspl3_w_G18_15(.douta(w_G18_15[0]),.doutb(w_G18_15[1]),.doutc(w_G18_15[2]),.din(w_G18_4[2]));
	jspl3 jspl3_w_G18_16(.douta(w_G18_16[0]),.doutb(w_G18_16[1]),.doutc(w_G18_16[2]),.din(w_G18_5[0]));
	jspl3 jspl3_w_G18_17(.douta(w_G18_17[0]),.doutb(w_G18_17[1]),.doutc(w_G18_17[2]),.din(w_G18_5[1]));
	jspl3 jspl3_w_G18_18(.douta(w_G18_18[0]),.doutb(w_G18_18[1]),.doutc(w_G18_18[2]),.din(w_G18_5[2]));
	jspl3 jspl3_w_G18_19(.douta(w_G18_19[0]),.doutb(w_G18_19[1]),.doutc(w_G18_19[2]),.din(w_G18_6[0]));
	jspl3 jspl3_w_G18_20(.douta(w_G18_20[0]),.doutb(w_G18_20[1]),.doutc(w_G18_20[2]),.din(w_G18_6[1]));
	jspl3 jspl3_w_G18_21(.douta(w_G18_21[0]),.doutb(w_G18_21[1]),.doutc(w_G18_21[2]),.din(w_G18_6[2]));
	jspl3 jspl3_w_G18_22(.douta(w_G18_22[0]),.doutb(w_G18_22[1]),.doutc(w_dff_A_p6fYGlLf3_2),.din(w_G18_7[0]));
	jspl3 jspl3_w_G18_23(.douta(w_dff_A_1y77Buen6_0),.doutb(w_G18_23[1]),.doutc(w_G18_23[2]),.din(w_G18_7[1]));
	jspl3 jspl3_w_G18_24(.douta(w_G18_24[0]),.doutb(w_G18_24[1]),.doutc(w_G18_24[2]),.din(w_G18_7[2]));
	jspl3 jspl3_w_G18_25(.douta(w_G18_25[0]),.doutb(w_G18_25[1]),.doutc(w_G18_25[2]),.din(w_G18_8[0]));
	jspl3 jspl3_w_G18_26(.douta(w_G18_26[0]),.doutb(w_G18_26[1]),.doutc(w_G18_26[2]),.din(w_G18_8[1]));
	jspl3 jspl3_w_G18_27(.douta(w_G18_27[0]),.doutb(w_G18_27[1]),.doutc(w_G18_27[2]),.din(w_G18_8[2]));
	jspl3 jspl3_w_G18_28(.douta(w_G18_28[0]),.doutb(w_G18_28[1]),.doutc(w_G18_28[2]),.din(w_G18_9[0]));
	jspl3 jspl3_w_G18_29(.douta(w_G18_29[0]),.doutb(w_G18_29[1]),.doutc(w_G18_29[2]),.din(w_G18_9[1]));
	jspl3 jspl3_w_G18_30(.douta(w_G18_30[0]),.doutb(w_G18_30[1]),.doutc(w_G18_30[2]),.din(w_G18_9[2]));
	jspl3 jspl3_w_G18_31(.douta(w_G18_31[0]),.doutb(w_G18_31[1]),.doutc(w_G18_31[2]),.din(w_G18_10[0]));
	jspl3 jspl3_w_G18_32(.douta(w_G18_32[0]),.doutb(w_G18_32[1]),.doutc(w_G18_32[2]),.din(w_G18_10[1]));
	jspl3 jspl3_w_G18_33(.douta(w_G18_33[0]),.doutb(w_G18_33[1]),.doutc(w_G18_33[2]),.din(w_G18_10[2]));
	jspl3 jspl3_w_G18_34(.douta(w_G18_34[0]),.doutb(w_G18_34[1]),.doutc(w_G18_34[2]),.din(w_G18_11[0]));
	jspl3 jspl3_w_G18_35(.douta(w_G18_35[0]),.doutb(w_G18_35[1]),.doutc(w_G18_35[2]),.din(w_G18_11[1]));
	jspl3 jspl3_w_G18_36(.douta(w_G18_36[0]),.doutb(w_G18_36[1]),.doutc(w_G18_36[2]),.din(w_G18_11[2]));
	jspl3 jspl3_w_G18_37(.douta(w_G18_37[0]),.doutb(w_G18_37[1]),.doutc(w_G18_37[2]),.din(w_G18_12[0]));
	jspl3 jspl3_w_G18_38(.douta(w_G18_38[0]),.doutb(w_G18_38[1]),.doutc(w_G18_38[2]),.din(w_G18_12[1]));
	jspl3 jspl3_w_G18_39(.douta(w_G18_39[0]),.doutb(w_G18_39[1]),.doutc(w_G18_39[2]),.din(w_G18_12[2]));
	jspl3 jspl3_w_G18_40(.douta(w_G18_40[0]),.doutb(w_G18_40[1]),.doutc(w_G18_40[2]),.din(w_G18_13[0]));
	jspl3 jspl3_w_G18_41(.douta(w_G18_41[0]),.doutb(w_G18_41[1]),.doutc(w_G18_41[2]),.din(w_G18_13[1]));
	jspl3 jspl3_w_G18_42(.douta(w_G18_42[0]),.doutb(w_G18_42[1]),.doutc(w_G18_42[2]),.din(w_G18_13[2]));
	jspl3 jspl3_w_G18_43(.douta(w_G18_43[0]),.doutb(w_G18_43[1]),.doutc(w_G18_43[2]),.din(w_G18_14[0]));
	jspl3 jspl3_w_G18_44(.douta(w_G18_44[0]),.doutb(w_G18_44[1]),.doutc(w_G18_44[2]),.din(w_G18_14[1]));
	jspl3 jspl3_w_G18_45(.douta(w_G18_45[0]),.doutb(w_G18_45[1]),.doutc(w_G18_45[2]),.din(w_G18_14[2]));
	jspl3 jspl3_w_G18_46(.douta(w_G18_46[0]),.doutb(w_G18_46[1]),.doutc(w_G18_46[2]),.din(w_G18_15[0]));
	jspl3 jspl3_w_G18_47(.douta(w_G18_47[0]),.doutb(w_G18_47[1]),.doutc(w_G18_47[2]),.din(w_G18_15[1]));
	jspl3 jspl3_w_G18_48(.douta(w_G18_48[0]),.doutb(w_G18_48[1]),.doutc(w_G18_48[2]),.din(w_G18_15[2]));
	jspl3 jspl3_w_G18_49(.douta(w_G18_49[0]),.doutb(w_G18_49[1]),.doutc(w_G18_49[2]),.din(w_G18_16[0]));
	jspl3 jspl3_w_G18_50(.douta(w_G18_50[0]),.doutb(w_G18_50[1]),.doutc(w_G18_50[2]),.din(w_G18_16[1]));
	jspl3 jspl3_w_G18_51(.douta(w_G18_51[0]),.doutb(w_G18_51[1]),.doutc(w_G18_51[2]),.din(w_G18_16[2]));
	jspl3 jspl3_w_G18_52(.douta(w_G18_52[0]),.doutb(w_G18_52[1]),.doutc(w_G18_52[2]),.din(w_G18_17[0]));
	jspl3 jspl3_w_G18_53(.douta(w_G18_53[0]),.doutb(w_G18_53[1]),.doutc(w_dff_A_n0yhwvps7_2),.din(w_G18_17[1]));
	jspl3 jspl3_w_G18_54(.douta(w_G18_54[0]),.doutb(w_dff_A_NME46QeS8_1),.doutc(w_G18_54[2]),.din(w_G18_17[2]));
	jspl3 jspl3_w_G18_55(.douta(w_dff_A_Ez3fDP7O2_0),.doutb(w_G18_55[1]),.doutc(w_dff_A_LnfPSjCj1_2),.din(w_G18_18[0]));
	jspl3 jspl3_w_G18_56(.douta(w_dff_A_g8Yd2so27_0),.doutb(w_G18_56[1]),.doutc(w_dff_A_e7OVtupO2_2),.din(w_G18_18[1]));
	jspl3 jspl3_w_G18_57(.douta(w_G18_57[0]),.doutb(w_dff_A_siTTxv4V7_1),.doutc(w_G18_57[2]),.din(w_G18_18[2]));
	jspl3 jspl3_w_G18_58(.douta(w_G18_58[0]),.doutb(w_G18_58[1]),.doutc(w_dff_A_JffuGsQJ7_2),.din(w_G18_19[0]));
	jspl3 jspl3_w_G38_0(.douta(w_G38_0[0]),.doutb(w_dff_A_WJWqTm6j3_1),.doutc(w_dff_A_DvvVmoVy6_2),.din(G38));
	jspl3 jspl3_w_G38_1(.douta(w_dff_A_5gGa3kNr3_0),.doutb(w_G38_1[1]),.doutc(w_dff_A_VmzUsI6k4_2),.din(w_G38_0[0]));
	jspl3 jspl3_w_G41_0(.douta(w_dff_A_VMwgvIR75_0),.doutb(w_dff_A_1JWV0Pyl7_1),.doutc(w_G41_0[2]),.din(G41));
	jspl jspl_w_G69_0(.douta(w_G69_0[0]),.doutb(w_G69_0[1]),.din(G69));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(G70));
	jspl3 jspl3_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.doutc(w_G106_0[2]),.din(G106));
	jspl jspl_w_G106_1(.douta(w_dff_A_pPlrvx5T9_0),.doutb(w_G106_1[1]),.din(w_G106_0[0]));
	jspl jspl_w_G229_0(.douta(w_G229_0[0]),.doutb(w_G229_0[1]),.din(G229));
	jspl3 jspl3_w_G1455_0(.douta(w_G1455_0[0]),.doutb(w_G1455_0[1]),.doutc(w_G1455_0[2]),.din(G1455));
	jspl jspl_w_G1459_0(.douta(w_G1459_0[0]),.doutb(w_dff_A_Aax5Nc2t1_1),.din(G1459));
	jspl3 jspl3_w_G1462_0(.douta(w_G1462_0[0]),.doutb(w_G1462_0[1]),.doutc(w_G1462_0[2]),.din(G1462));
	jspl3 jspl3_w_G1469_0(.douta(w_G1469_0[0]),.doutb(w_G1469_0[1]),.doutc(w_G1469_0[2]),.din(G1469));
	jspl jspl_w_G1469_1(.douta(w_dff_A_6HCsU9672_0),.doutb(w_G1469_1[1]),.din(w_G1469_0[0]));
	jspl3 jspl3_w_G1480_0(.douta(w_G1480_0[0]),.doutb(w_G1480_0[1]),.doutc(w_G1480_0[2]),.din(G1480));
	jspl3 jspl3_w_G1486_0(.douta(w_G1486_0[0]),.doutb(w_G1486_0[1]),.doutc(w_G1486_0[2]),.din(G1486));
	jspl3 jspl3_w_G1492_0(.douta(w_G1492_0[0]),.doutb(w_G1492_0[1]),.doutc(w_G1492_0[2]),.din(G1492));
	jspl jspl_w_G1492_1(.douta(w_G1492_1[0]),.doutb(w_G1492_1[1]),.din(w_G1492_0[0]));
	jspl3 jspl3_w_G1496_0(.douta(w_G1496_0[0]),.doutb(w_G1496_0[1]),.doutc(w_G1496_0[2]),.din(G1496));
	jspl3 jspl3_w_G2204_0(.douta(w_G2204_0[0]),.doutb(w_G2204_0[1]),.doutc(w_G2204_0[2]),.din(G2204));
	jspl jspl_w_G2208_0(.douta(w_G2208_0[0]),.doutb(w_dff_A_xccNKG1p6_1),.din(G2208));
	jspl3 jspl3_w_G2211_0(.douta(w_G2211_0[0]),.doutb(w_G2211_0[1]),.doutc(w_G2211_0[2]),.din(G2211));
	jspl3 jspl3_w_G2218_0(.douta(w_G2218_0[0]),.doutb(w_G2218_0[1]),.doutc(w_G2218_0[2]),.din(G2218));
	jspl3 jspl3_w_G2224_0(.douta(w_G2224_0[0]),.doutb(w_G2224_0[1]),.doutc(w_G2224_0[2]),.din(G2224));
	jspl jspl_w_G2224_1(.douta(w_dff_A_mm6HwVJP0_0),.doutb(w_G2224_1[1]),.din(w_G2224_0[0]));
	jspl3 jspl3_w_G2230_0(.douta(w_G2230_0[0]),.doutb(w_G2230_0[1]),.doutc(w_G2230_0[2]),.din(G2230));
	jspl jspl_w_G2230_1(.douta(w_dff_A_1rQxkaMZ6_0),.doutb(w_G2230_1[1]),.din(w_G2230_0[0]));
	jspl3 jspl3_w_G2236_0(.douta(w_G2236_0[0]),.doutb(w_G2236_0[1]),.doutc(w_G2236_0[2]),.din(G2236));
	jspl jspl_w_G2236_1(.douta(w_dff_A_j7vDye4R5_0),.doutb(w_G2236_1[1]),.din(w_G2236_0[0]));
	jspl3 jspl3_w_G2239_0(.douta(w_G2239_0[0]),.doutb(w_dff_A_mBJGbxOA3_1),.doutc(w_G2239_0[2]),.din(G2239));
	jspl3 jspl3_w_G2247_0(.douta(w_G2247_0[0]),.doutb(w_G2247_0[1]),.doutc(w_G2247_0[2]),.din(G2247));
	jspl3 jspl3_w_G2253_0(.douta(w_G2253_0[0]),.doutb(w_G2253_0[1]),.doutc(w_G2253_0[2]),.din(G2253));
	jspl jspl_w_G2253_1(.douta(w_dff_A_9uuk3uJU2_0),.doutb(w_G2253_1[1]),.din(w_G2253_0[0]));
	jspl3 jspl3_w_G2256_0(.douta(w_G2256_0[0]),.doutb(w_G2256_0[1]),.doutc(w_G2256_0[2]),.din(G2256));
	jspl jspl_w_G2256_1(.douta(w_dff_A_Of6m4djP1_0),.doutb(w_G2256_1[1]),.din(w_G2256_0[0]));
	jspl jspl_w_G3698_0(.douta(w_G3698_0[0]),.doutb(w_dff_A_ZmKoTLCU6_1),.din(G3698));
	jspl3 jspl3_w_G3701_0(.douta(w_dff_A_iUgl4et14_0),.doutb(w_G3701_0[1]),.doutc(w_G3701_0[2]),.din(G3701));
	jspl jspl_w_G3701_1(.douta(w_G3701_1[0]),.doutb(w_dff_A_MSVHLPQs9_1),.din(w_G3701_0[0]));
	jspl3 jspl3_w_G3705_0(.douta(w_G3705_0[0]),.doutb(w_G3705_0[1]),.doutc(w_G3705_0[2]),.din(G3705));
	jspl3 jspl3_w_G3705_1(.douta(w_dff_A_Pbera6bC7_0),.doutb(w_dff_A_r4uRtzhq8_1),.doutc(w_G3705_1[2]),.din(w_G3705_0[0]));
	jspl jspl_w_G3705_2(.douta(w_dff_A_MeHNMQtc8_0),.doutb(w_G3705_2[1]),.din(w_G3705_0[1]));
	jspl3 jspl3_w_G3711_0(.douta(w_G3711_0[0]),.doutb(w_G3711_0[1]),.doutc(w_G3711_0[2]),.din(G3711));
	jspl jspl_w_G3711_1(.douta(w_dff_A_nDhm2kq96_0),.doutb(w_G3711_1[1]),.din(w_G3711_0[0]));
	jspl3 jspl3_w_G3717_0(.douta(w_G3717_0[0]),.doutb(w_dff_A_MjfUwtZn7_1),.doutc(w_G3717_0[2]),.din(G3717));
	jspl3 jspl3_w_G3717_1(.douta(w_dff_A_fUSrVCF72_0),.doutb(w_dff_A_SXnMlaJE4_1),.doutc(w_G3717_1[2]),.din(w_G3717_0[0]));
	jspl jspl_w_G3717_2(.douta(w_G3717_2[0]),.doutb(w_dff_A_Y5zX2Jn48_1),.din(w_G3717_0[1]));
	jspl3 jspl3_w_G3723_0(.douta(w_G3723_0[0]),.doutb(w_G3723_0[1]),.doutc(w_dff_A_heDmG2sM6_2),.din(G3723));
	jspl jspl_w_G3723_1(.douta(w_dff_A_WhROGiIe9_0),.doutb(w_G3723_1[1]),.din(w_G3723_0[0]));
	jspl3 jspl3_w_G3729_0(.douta(w_G3729_0[0]),.doutb(w_G3729_0[1]),.doutc(w_dff_A_aF5AZzhG1_2),.din(G3729));
	jspl jspl_w_G3729_1(.douta(w_dff_A_FABQIxU61_0),.doutb(w_G3729_1[1]),.din(w_G3729_0[0]));
	jspl3 jspl3_w_G3737_0(.douta(w_G3737_0[0]),.doutb(w_G3737_0[1]),.doutc(w_G3737_0[2]),.din(G3737));
	jspl jspl_w_G3737_1(.douta(w_dff_A_HfR9wvXH0_0),.doutb(w_G3737_1[1]),.din(w_G3737_0[0]));
	jspl3 jspl3_w_G3743_0(.douta(w_dff_A_vVahhG232_0),.doutb(w_G3743_0[1]),.doutc(w_G3743_0[2]),.din(G3743));
	jspl3 jspl3_w_G3743_1(.douta(w_dff_A_yxDm7fX93_0),.doutb(w_dff_A_j8emn42k0_1),.doutc(w_G3743_1[2]),.din(w_G3743_0[0]));
	jspl3 jspl3_w_G3749_0(.douta(w_dff_A_6QumpSRY2_0),.doutb(w_G3749_0[1]),.doutc(w_G3749_0[2]),.din(G3749));
	jspl jspl_w_G3749_1(.douta(w_G3749_1[0]),.doutb(w_G3749_1[1]),.din(w_G3749_0[0]));
	jspl jspl_w_G4393_0(.douta(w_G4393_0[0]),.doutb(w_dff_A_8eJPHOff4_1),.din(G4393));
	jspl3 jspl3_w_G4394_0(.douta(w_dff_A_F6zSoCrM3_0),.doutb(w_G4394_0[1]),.doutc(w_G4394_0[2]),.din(G4394));
	jspl jspl_w_G4394_1(.douta(w_G4394_1[0]),.doutb(w_G4394_1[1]),.din(w_G4394_0[0]));
	jspl3 jspl3_w_G4400_0(.douta(w_G4400_0[0]),.doutb(w_G4400_0[1]),.doutc(w_G4400_0[2]),.din(G4400));
	jspl3 jspl3_w_G4405_0(.douta(w_dff_A_J2qPaUXQ6_0),.doutb(w_G4405_0[1]),.doutc(w_G4405_0[2]),.din(G4405));
	jspl3 jspl3_w_G4405_1(.douta(w_G4405_1[0]),.doutb(w_G4405_1[1]),.doutc(w_G4405_1[2]),.din(w_G4405_0[0]));
	jspl3 jspl3_w_G4410_0(.douta(w_G4410_0[0]),.doutb(w_G4410_0[1]),.doutc(w_G4410_0[2]),.din(G4410));
	jspl jspl_w_G4410_1(.douta(w_dff_A_6pxG1Fq52_0),.doutb(w_G4410_1[1]),.din(w_G4410_0[0]));
	jspl3 jspl3_w_G4415_0(.douta(w_G4415_0[0]),.doutb(w_G4415_0[1]),.doutc(w_G4415_0[2]),.din(G4415));
	jspl jspl_w_G4415_1(.douta(w_dff_A_YppMUfdg6_0),.doutb(w_G4415_1[1]),.din(w_G4415_0[0]));
	jspl3 jspl3_w_G4420_0(.douta(w_G4420_0[0]),.doutb(w_dff_A_8eBzixrq7_1),.doutc(w_G4420_0[2]),.din(G4420));
	jspl jspl_w_G4427_0(.douta(w_G4427_0[0]),.doutb(w_G4427_0[1]),.din(G4427));
	jspl3 jspl3_w_G4432_0(.douta(w_G4432_0[0]),.doutb(w_G4432_0[1]),.doutc(w_G4432_0[2]),.din(G4432));
	jspl jspl_w_G4432_1(.douta(w_dff_A_vK1SaVCu5_0),.doutb(w_G4432_1[1]),.din(w_G4432_0[0]));
	jspl3 jspl3_w_G4437_0(.douta(w_G4437_0[0]),.doutb(w_dff_A_VgHUHFeN3_1),.doutc(w_G4437_0[2]),.din(G4437));
	jspl3 jspl3_w_G4526_0(.douta(w_G4526_0[0]),.doutb(w_dff_A_d505jNZO2_1),.doutc(w_dff_A_CGzIPUJQ0_2),.din(G4526));
	jspl jspl_w_G4526_1(.douta(w_G4526_1[0]),.doutb(w_dff_A_ms5Q6tOQ7_1),.din(w_G4526_0[0]));
	jspl3 jspl3_w_G4528_0(.douta(w_G4528_0[0]),.doutb(w_G4528_0[1]),.doutc(w_G4528_0[2]),.din(G4528));
	jspl jspl_w_G404_0(.douta(w_G404_0),.doutb(w_dff_A_amYEkAj00_1),.din(G404_fa_));
	jspl jspl_w_G406_0(.douta(w_G406_0),.doutb(w_dff_A_t6zLtL210_1),.din(G406_fa_));
	jspl jspl_w_G408_0(.douta(w_G408_0),.doutb(w_dff_A_08FIgT3x3_1),.din(G408_fa_));
	jspl jspl_w_G410_0(.douta(w_G410_0),.doutb(w_dff_A_OYPAWhe44_1),.din(G410_fa_));
	jspl jspl_w_G412_0(.douta(w_G412_0),.doutb(w_dff_A_wykqDbm08_1),.din(G412_fa_));
	jspl jspl_w_G414_0(.douta(w_dff_A_CfZ6Oqln4_0),.doutb(w_dff_A_nyyEt9jd2_1),.din(G414_fa_));
	jspl jspl_w_G416_0(.douta(w_G416_0),.doutb(w_dff_A_5Phao2qY9_1),.din(G416_fa_));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(n345));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl3 jspl3_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.doutc(w_n353_0[2]),.din(n353));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_dff_A_b2eYmO4R5_2),.din(w_dff_B_KidPtzUp6_3));
	jspl3 jspl3_w_n354_1(.douta(w_dff_A_5gSkhRnC7_0),.doutb(w_n354_1[1]),.doutc(w_n354_1[2]),.din(w_n354_0[0]));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl3 jspl3_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.doutc(w_n355_1[2]),.din(w_n355_0[0]));
	jspl3 jspl3_w_n355_2(.douta(w_n355_2[0]),.doutb(w_n355_2[1]),.doutc(w_n355_2[2]),.din(w_n355_0[1]));
	jspl3 jspl3_w_n355_3(.douta(w_n355_3[0]),.doutb(w_n355_3[1]),.doutc(w_n355_3[2]),.din(w_n355_0[2]));
	jspl3 jspl3_w_n355_4(.douta(w_n355_4[0]),.doutb(w_n355_4[1]),.doutc(w_n355_4[2]),.din(w_n355_1[0]));
	jspl3 jspl3_w_n355_5(.douta(w_n355_5[0]),.doutb(w_n355_5[1]),.doutc(w_n355_5[2]),.din(w_n355_1[1]));
	jspl3 jspl3_w_n355_6(.douta(w_n355_6[0]),.doutb(w_n355_6[1]),.doutc(w_n355_6[2]),.din(w_n355_1[2]));
	jspl3 jspl3_w_n355_7(.douta(w_n355_7[0]),.doutb(w_n355_7[1]),.doutc(w_n355_7[2]),.din(w_n355_2[0]));
	jspl3 jspl3_w_n355_8(.douta(w_n355_8[0]),.doutb(w_n355_8[1]),.doutc(w_n355_8[2]),.din(w_n355_2[1]));
	jspl3 jspl3_w_n355_9(.douta(w_n355_9[0]),.doutb(w_n355_9[1]),.doutc(w_n355_9[2]),.din(w_n355_2[2]));
	jspl3 jspl3_w_n355_10(.douta(w_n355_10[0]),.doutb(w_dff_A_3iXJCCI03_1),.doutc(w_n355_10[2]),.din(w_n355_3[0]));
	jspl3 jspl3_w_n355_11(.douta(w_n355_11[0]),.doutb(w_n355_11[1]),.doutc(w_n355_11[2]),.din(w_n355_3[1]));
	jspl3 jspl3_w_n355_12(.douta(w_n355_12[0]),.doutb(w_n355_12[1]),.doutc(w_n355_12[2]),.din(w_n355_3[2]));
	jspl3 jspl3_w_n355_13(.douta(w_n355_13[0]),.doutb(w_n355_13[1]),.doutc(w_n355_13[2]),.din(w_n355_4[0]));
	jspl3 jspl3_w_n355_14(.douta(w_n355_14[0]),.doutb(w_n355_14[1]),.doutc(w_n355_14[2]),.din(w_n355_4[1]));
	jspl3 jspl3_w_n355_15(.douta(w_n355_15[0]),.doutb(w_n355_15[1]),.doutc(w_n355_15[2]),.din(w_n355_4[2]));
	jspl3 jspl3_w_n355_16(.douta(w_n355_16[0]),.doutb(w_n355_16[1]),.doutc(w_n355_16[2]),.din(w_n355_5[0]));
	jspl3 jspl3_w_n355_17(.douta(w_n355_17[0]),.doutb(w_n355_17[1]),.doutc(w_n355_17[2]),.din(w_n355_5[1]));
	jspl3 jspl3_w_n355_18(.douta(w_n355_18[0]),.doutb(w_n355_18[1]),.doutc(w_n355_18[2]),.din(w_n355_5[2]));
	jspl3 jspl3_w_n355_19(.douta(w_n355_19[0]),.doutb(w_n355_19[1]),.doutc(w_n355_19[2]),.din(w_n355_6[0]));
	jspl3 jspl3_w_n355_20(.douta(w_n355_20[0]),.doutb(w_n355_20[1]),.doutc(w_n355_20[2]),.din(w_n355_6[1]));
	jspl3 jspl3_w_n355_21(.douta(w_n355_21[0]),.doutb(w_n355_21[1]),.doutc(w_n355_21[2]),.din(w_n355_6[2]));
	jspl3 jspl3_w_n355_22(.douta(w_n355_22[0]),.doutb(w_n355_22[1]),.doutc(w_n355_22[2]),.din(w_n355_7[0]));
	jspl3 jspl3_w_n355_23(.douta(w_n355_23[0]),.doutb(w_n355_23[1]),.doutc(w_n355_23[2]),.din(w_n355_7[1]));
	jspl3 jspl3_w_n355_24(.douta(w_n355_24[0]),.doutb(w_n355_24[1]),.doutc(w_n355_24[2]),.din(w_n355_7[2]));
	jspl3 jspl3_w_n355_25(.douta(w_n355_25[0]),.doutb(w_n355_25[1]),.doutc(w_n355_25[2]),.din(w_n355_8[0]));
	jspl jspl_w_n355_26(.douta(w_n355_26[0]),.doutb(w_n355_26[1]),.din(w_n355_8[1]));
	jspl3 jspl3_w_n356_0(.douta(w_dff_A_5Sf6yYef6_0),.doutb(w_n356_0[1]),.doutc(w_n356_0[2]),.din(n356));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(n358));
	jspl jspl_w_n359_0(.douta(w_dff_A_sK9IWy2v7_0),.doutb(w_n359_0[1]),.din(n359));
	jspl3 jspl3_w_n362_0(.douta(w_dff_A_sOHOWnrF9_0),.doutb(w_n362_0[1]),.doutc(w_n362_0[2]),.din(n362));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_dff_A_9zWEW9xr4_1),.din(n365));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_dff_A_rkwUqV5s2_1),.din(n366));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(n370));
	jspl3 jspl3_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.doutc(w_n371_0[2]),.din(n371));
	jspl jspl_w_n371_1(.douta(w_n371_1[0]),.doutb(w_n371_1[1]),.din(w_n371_0[0]));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_OvmsPZXt0_1),.doutc(w_dff_A_nvfLFF5L2_2),.din(n372));
	jspl3 jspl3_w_n372_1(.douta(w_n372_1[0]),.doutb(w_dff_A_aPEOWLYQ7_1),.doutc(w_dff_A_sCnlMVHi9_2),.din(w_n372_0[0]));
	jspl jspl_w_n376_0(.douta(w_n376_0[0]),.doutb(w_n376_0[1]),.din(n376));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_dff_A_pzV3NkDf7_2),.din(n377));
	jspl3 jspl3_w_n377_1(.douta(w_n377_1[0]),.doutb(w_n377_1[1]),.doutc(w_n377_1[2]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n379_0(.douta(w_n379_0[0]),.doutb(w_dff_A_k9uy9nRV1_1),.doutc(w_dff_A_JeDlUWyh1_2),.din(n379));
	jspl jspl_w_n379_1(.douta(w_dff_A_uFNboZ7w4_0),.doutb(w_n379_1[1]),.din(w_n379_0[0]));
	jspl3 jspl3_w_n380_0(.douta(w_n380_0[0]),.doutb(w_dff_A_ujmd7dth2_1),.doutc(w_dff_A_QCnVwtnx0_2),.din(n380));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_dff_A_GOOt5XX88_2),.din(n387));
	jspl3 jspl3_w_n387_1(.douta(w_n387_1[0]),.doutb(w_dff_A_fptldo2Z1_1),.doutc(w_dff_A_8zOw0JFN9_2),.din(w_n387_0[0]));
	jspl3 jspl3_w_n388_0(.douta(w_dff_A_QLd0u7Pk2_0),.doutb(w_n388_0[1]),.doutc(w_dff_A_t2vvxLIv2_2),.din(w_dff_B_mLOxX17m9_3));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_dff_A_NVapzCBn3_1),.din(n389));
	jspl3 jspl3_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.doutc(w_dff_A_oaivMi756_2),.din(w_dff_B_26IBZNyP1_3));
	jspl jspl_w_n390_1(.douta(w_n390_1[0]),.doutb(w_n390_1[1]),.din(w_n390_0[0]));
	jspl3 jspl3_w_n395_0(.douta(w_dff_A_uSWqszjk6_0),.doutb(w_n395_0[1]),.doutc(w_n395_0[2]),.din(n395));
	jspl jspl_w_n400_0(.douta(w_n400_0[0]),.doutb(w_n400_0[1]),.din(n400));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n401_1(.douta(w_n401_1[0]),.doutb(w_n401_1[1]),.doutc(w_n401_1[2]),.din(w_n401_0[0]));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_dff_A_7gf8DVbR1_1),.doutc(w_dff_A_QTlFZtkZ7_2),.din(n402));
	jspl jspl_w_n402_1(.douta(w_n402_1[0]),.doutb(w_dff_A_DknvD8Cx1_1),.din(w_n402_0[0]));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl jspl_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.din(n404));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl3 jspl3_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.doutc(w_dff_A_VW7Yj6298_2),.din(n407));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl jspl_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.din(n410));
	jspl3 jspl3_w_n412_0(.douta(w_dff_A_qPeJQYRD1_0),.doutb(w_dff_A_9H4knwf08_1),.doutc(w_n412_0[2]),.din(n412));
	jspl3 jspl3_w_n413_0(.douta(w_dff_A_74cnW4016_0),.doutb(w_n413_0[1]),.doutc(w_n413_0[2]),.din(n413));
	jspl jspl_w_n413_1(.douta(w_dff_A_8TRro6Rh2_0),.doutb(w_n413_1[1]),.din(w_n413_0[0]));
	jspl3 jspl3_w_n417_0(.douta(w_dff_A_PFrRtPz72_0),.doutb(w_dff_A_Mu6B6EbU7_1),.doutc(w_n417_0[2]),.din(n417));
	jspl jspl_w_n419_0(.douta(w_n419_0[0]),.doutb(w_dff_A_sBgJxJKt1_1),.din(n419));
	jspl3 jspl3_w_n422_0(.douta(w_n422_0[0]),.doutb(w_dff_A_sTYy0b9H1_1),.doutc(w_n422_0[2]),.din(n422));
	jspl3 jspl3_w_n422_1(.douta(w_n422_1[0]),.doutb(w_n422_1[1]),.doutc(w_n422_1[2]),.din(w_n422_0[0]));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(n427));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.doutc(w_n428_0[2]),.din(n428));
	jspl3 jspl3_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.doutc(w_n429_0[2]),.din(n429));
	jspl3 jspl3_w_n429_1(.douta(w_n429_1[0]),.doutb(w_n429_1[1]),.doutc(w_dff_A_SuogiHgF1_2),.din(w_n429_0[0]));
	jspl jspl_w_n429_2(.douta(w_n429_2[0]),.doutb(w_n429_2[1]),.din(w_n429_0[1]));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_dff_A_zUKcF8oA4_1),.din(n430));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl jspl_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.din(w_n435_0[0]));
	jspl jspl_w_n436_0(.douta(w_dff_A_mtPxmBZR7_0),.doutb(w_n436_0[1]),.din(n436));
	jspl jspl_w_n437_0(.douta(w_dff_A_7zf17ZJ46_0),.doutb(w_n437_0[1]),.din(w_dff_B_cteXpGLd6_2));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl3 jspl3_w_n442_0(.douta(w_n442_0[0]),.doutb(w_n442_0[1]),.doutc(w_n442_0[2]),.din(n442));
	jspl jspl_w_n443_0(.douta(w_dff_A_qg2u1FFT9_0),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n445_0(.douta(w_dff_A_jCSaDnGt3_0),.doutb(w_n445_0[1]),.din(w_dff_B_PlwNksKA7_2));
	jspl3 jspl3_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.doutc(w_dff_A_Mbxmu5IA8_2),.din(n446));
	jspl jspl_w_n446_1(.douta(w_dff_A_NBaBoVcZ7_0),.doutb(w_n446_1[1]),.din(w_n446_0[0]));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.din(n448));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n450_0(.douta(w_n450_0[0]),.doutb(w_dff_A_yGPNZGOU3_1),.doutc(w_dff_A_DQ9xXhsI5_2),.din(w_dff_B_JFMYzIFG6_3));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_dff_A_ayvScaaT2_1),.din(n452));
	jspl jspl_w_n454_0(.douta(w_n454_0[0]),.doutb(w_n454_0[1]),.din(n454));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_dff_A_7KKGRqGr4_1),.din(n455));
	jspl3 jspl3_w_n456_0(.douta(w_n456_0[0]),.doutb(w_dff_A_41bqDbRo2_1),.doutc(w_dff_A_fSaZrFse3_2),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(w_dff_B_aoQ4cO6G4_2));
	jspl3 jspl3_w_n458_0(.douta(w_n458_0[0]),.doutb(w_dff_A_v5z2xYqi5_1),.doutc(w_n458_0[2]),.din(n458));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_dff_A_UFFdpIeU1_1),.doutc(w_n460_0[2]),.din(n460));
	jspl jspl_w_n461_0(.douta(w_dff_A_Eo8pjj496_0),.doutb(w_n461_0[1]),.din(n461));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_PKKRSAtR4_1),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_dff_A_GO7S0n6C9_1),.din(n464));
	jspl3 jspl3_w_n465_0(.douta(w_dff_A_b5VbxXny3_0),.doutb(w_n465_0[1]),.doutc(w_n465_0[2]),.din(n465));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(w_dff_B_jr5IL4iN8_2));
	jspl jspl_w_n468_0(.douta(w_n468_0[0]),.doutb(w_n468_0[1]),.din(n468));
	jspl3 jspl3_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.doutc(w_n469_0[2]),.din(n469));
	jspl jspl_w_n469_1(.douta(w_n469_1[0]),.doutb(w_n469_1[1]),.din(w_n469_0[0]));
	jspl3 jspl3_w_n470_0(.douta(w_dff_A_R0cohlg94_0),.doutb(w_n470_0[1]),.doutc(w_dff_A_Iu8Av3AH3_2),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(w_dff_B_QCLCXMcC4_3));
	jspl jspl_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.din(n473));
	jspl3 jspl3_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.doutc(w_n474_0[2]),.din(n474));
	jspl jspl_w_n474_1(.douta(w_n474_1[0]),.doutb(w_n474_1[1]),.din(w_n474_0[0]));
	jspl3 jspl3_w_n475_0(.douta(w_n475_0[0]),.doutb(w_dff_A_Ar2t3l8F8_1),.doutc(w_dff_A_KGEqSJ7R2_2),.din(n475));
	jspl jspl_w_n475_1(.douta(w_n475_1[0]),.doutb(w_dff_A_UMlRGQE61_1),.din(w_n475_0[0]));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(n479));
	jspl3 jspl3_w_n480_0(.douta(w_n480_0[0]),.doutb(w_dff_A_tVXKqJGB9_1),.doutc(w_dff_A_NwdEVlzB8_2),.din(n480));
	jspl jspl_w_n480_1(.douta(w_dff_A_PXkeGuLe9_0),.doutb(w_n480_1[1]),.din(w_n480_0[0]));
	jspl3 jspl3_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.doutc(w_n481_0[2]),.din(n481));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(w_dff_B_2P58I5eT7_2));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl3 jspl3_w_n485_0(.douta(w_n485_0[0]),.doutb(w_n485_0[1]),.doutc(w_n485_0[2]),.din(n485));
	jspl3 jspl3_w_n486_0(.douta(w_dff_A_xdlzvDjW9_0),.doutb(w_n486_0[1]),.doutc(w_dff_A_x71sLdCq3_2),.din(n486));
	jspl jspl_w_n488_0(.douta(w_n488_0[0]),.doutb(w_n488_0[1]),.din(n488));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(n489));
	jspl3 jspl3_w_n490_0(.douta(w_n490_0[0]),.doutb(w_n490_0[1]),.doutc(w_n490_0[2]),.din(n490));
	jspl3 jspl3_w_n491_0(.douta(w_n491_0[0]),.doutb(w_dff_A_IxiQpLBq7_1),.doutc(w_n491_0[2]),.din(n491));
	jspl jspl_w_n491_1(.douta(w_n491_1[0]),.doutb(w_n491_1[1]),.din(w_n491_0[0]));
	jspl jspl_w_n493_0(.douta(w_dff_A_ajUlbdyL5_0),.doutb(w_n493_0[1]),.din(n493));
	jspl jspl_w_n494_0(.douta(w_dff_A_tOfU8hJU1_0),.doutb(w_n494_0[1]),.din(n494));
	jspl jspl_w_n502_0(.douta(w_dff_A_WeQLK4OR9_0),.doutb(w_n502_0[1]),.din(w_dff_B_Kmrt3sfJ7_2));
	jspl jspl_w_n503_0(.douta(w_dff_A_zzibIUZP2_0),.doutb(w_n503_0[1]),.din(n503));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_dff_A_L8v9zKPK0_1),.din(w_dff_B_BpLrxlZp9_2));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_dff_A_zIdw6yhx1_2),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n509_0(.douta(w_dff_A_U0hXA5h91_0),.doutb(w_n509_0[1]),.din(n509));
	jspl jspl_w_n510_0(.douta(w_dff_A_6U1UqLW16_0),.doutb(w_n510_0[1]),.din(n510));
	jspl jspl_w_n512_0(.douta(w_dff_A_NdcOEkCb6_0),.doutb(w_n512_0[1]),.din(n512));
	jspl3 jspl3_w_n514_0(.douta(w_n514_0[0]),.doutb(w_dff_A_pH4My2IA7_1),.doutc(w_n514_0[2]),.din(n514));
	jspl3 jspl3_w_n516_0(.douta(w_n516_0[0]),.doutb(w_dff_A_5qzCAV2S8_1),.doutc(w_n516_0[2]),.din(n516));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_dff_A_5nLHnB6C4_1),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(n519));
	jspl3 jspl3_w_n520_0(.douta(w_n520_0[0]),.doutb(w_dff_A_rPxpNk2v5_1),.doutc(w_dff_A_t8sJnWpR2_2),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.doutc(w_n523_0[2]),.din(n523));
	jspl3 jspl3_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.doutc(w_dff_A_Iuxr2gKJ8_2),.din(n524));
	jspl3 jspl3_w_n524_1(.douta(w_n524_1[0]),.doutb(w_dff_A_50Pk9rpa7_1),.doutc(w_dff_A_GMvBdxUO4_2),.din(w_n524_0[0]));
	jspl jspl_w_n524_2(.douta(w_n524_2[0]),.doutb(w_n524_2[1]),.din(w_n524_0[1]));
	jspl3 jspl3_w_n525_0(.douta(w_n525_0[0]),.doutb(w_dff_A_4E7K3r0y5_1),.doutc(w_dff_A_JIK2jnnq1_2),.din(n525));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl3 jspl3_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.doutc(w_n528_0[2]),.din(n528));
	jspl jspl_w_n528_1(.douta(w_n528_1[0]),.doutb(w_n528_1[1]),.din(w_n528_0[0]));
	jspl jspl_w_n529_0(.douta(w_dff_A_CscisU493_0),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n530_0(.douta(w_dff_A_CmHLRX2u3_0),.doutb(w_n530_0[1]),.din(n530));
	jspl3 jspl3_w_n531_0(.douta(w_n531_0[0]),.doutb(w_dff_A_T9rOa2NS6_1),.doutc(w_dff_A_bcAtzUew4_2),.din(n531));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl3 jspl3_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.doutc(w_n534_0[2]),.din(n534));
	jspl jspl_w_n534_1(.douta(w_n534_1[0]),.doutb(w_n534_1[1]),.din(w_n534_0[0]));
	jspl3 jspl3_w_n535_0(.douta(w_n535_0[0]),.doutb(w_dff_A_egm8n0ej7_1),.doutc(w_n535_0[2]),.din(n535));
	jspl jspl_w_n535_1(.douta(w_dff_A_1GIilQCR3_0),.doutb(w_n535_1[1]),.din(w_n535_0[0]));
	jspl jspl_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.din(w_dff_B_clWffWiI2_2));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl3 jspl3_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.doutc(w_n539_0[2]),.din(n539));
	jspl jspl_w_n539_1(.douta(w_n539_1[0]),.doutb(w_n539_1[1]),.din(w_n539_0[0]));
	jspl3 jspl3_w_n540_0(.douta(w_dff_A_IlnJLqiF5_0),.doutb(w_dff_A_nW4mItQv2_1),.doutc(w_n540_0[2]),.din(n540));
	jspl jspl_w_n542_0(.douta(w_dff_A_DjpXitUl9_0),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n549_0(.douta(w_n549_0[0]),.doutb(w_dff_A_x19YsS0i6_1),.din(w_dff_B_rFAGAFOx4_2));
	jspl jspl_w_n551_0(.douta(w_dff_A_EYlpZPJq4_0),.doutb(w_n551_0[1]),.din(n551));
	jspl jspl_w_n552_0(.douta(w_dff_A_EZo0lXF13_0),.doutb(w_n552_0[1]),.din(n552));
	jspl jspl_w_n553_0(.douta(w_dff_A_5dgnjyY68_0),.doutb(w_n553_0[1]),.din(w_dff_B_JGSCKHOj3_2));
	jspl3 jspl3_w_n554_0(.douta(w_n554_0[0]),.doutb(w_dff_A_ck0iszft9_1),.doutc(w_n554_0[2]),.din(n554));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_dff_A_W9Oe9Irk5_1),.doutc(w_n556_0[2]),.din(n556));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl3 jspl3_w_n558_0(.douta(w_dff_A_FnpgA7eZ4_0),.doutb(w_dff_A_XixEvbBh8_1),.doutc(w_n558_0[2]),.din(n558));
	jspl jspl_w_n560_0(.douta(w_dff_A_GOtlVnN46_0),.doutb(w_n560_0[1]),.din(n560));
	jspl3 jspl3_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.doutc(w_n562_0[2]),.din(n562));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(w_dff_B_YAXYqcGI0_2));
	jspl3 jspl3_w_n564_0(.douta(w_dff_A_VMS3oj4g6_0),.doutb(w_dff_A_d8qwEVrX0_1),.doutc(w_n564_0[2]),.din(n564));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl3 jspl3_w_n565_1(.douta(w_n565_1[0]),.doutb(w_n565_1[1]),.doutc(w_n565_1[2]),.din(w_n565_0[0]));
	jspl3 jspl3_w_n565_2(.douta(w_n565_2[0]),.doutb(w_n565_2[1]),.doutc(w_n565_2[2]),.din(w_n565_0[1]));
	jspl3 jspl3_w_n565_3(.douta(w_n565_3[0]),.doutb(w_n565_3[1]),.doutc(w_n565_3[2]),.din(w_n565_0[2]));
	jspl3 jspl3_w_n565_4(.douta(w_dff_A_tvyGr8hS2_0),.doutb(w_dff_A_mwjuaXS58_1),.doutc(w_n565_4[2]),.din(w_n565_1[0]));
	jspl3 jspl3_w_n565_5(.douta(w_n565_5[0]),.doutb(w_n565_5[1]),.doutc(w_n565_5[2]),.din(w_n565_1[1]));
	jspl3 jspl3_w_n565_6(.douta(w_n565_6[0]),.doutb(w_n565_6[1]),.doutc(w_n565_6[2]),.din(w_n565_1[2]));
	jspl3 jspl3_w_n565_7(.douta(w_n565_7[0]),.doutb(w_n565_7[1]),.doutc(w_n565_7[2]),.din(w_n565_2[0]));
	jspl3 jspl3_w_n565_8(.douta(w_n565_8[0]),.doutb(w_n565_8[1]),.doutc(w_n565_8[2]),.din(w_n565_2[1]));
	jspl3 jspl3_w_n565_9(.douta(w_n565_9[0]),.doutb(w_n565_9[1]),.doutc(w_n565_9[2]),.din(w_n565_2[2]));
	jspl jspl_w_n565_10(.douta(w_n565_10[0]),.doutb(w_n565_10[1]),.din(w_n565_3[0]));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n567_1(.douta(w_n567_1[0]),.doutb(w_n567_1[1]),.din(w_n567_0[0]));
	jspl3 jspl3_w_n568_0(.douta(w_dff_A_7k2u0Uhk4_0),.doutb(w_n568_0[1]),.doutc(w_dff_A_KB6PSNHp2_2),.din(n568));
	jspl3 jspl3_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.doutc(w_n569_0[2]),.din(w_dff_B_syGTL4xv9_3));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_dff_A_Ao79kSAN0_2),.din(n572));
	jspl jspl_w_n572_1(.douta(w_n572_1[0]),.doutb(w_n572_1[1]),.din(w_n572_0[0]));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_dff_A_xnCWaTuR7_2),.din(n573));
	jspl jspl_w_n573_1(.douta(w_n573_1[0]),.doutb(w_n573_1[1]),.din(w_n573_0[0]));
	jspl jspl_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.din(w_dff_B_sKxW7ouH5_2));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl3 jspl3_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.doutc(w_n577_0[2]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_dff_A_qtJnsGNi4_1),.doutc(w_dff_A_AR6PB7eS3_2),.din(n578));
	jspl jspl_w_n578_1(.douta(w_dff_A_BLNwJD364_0),.doutb(w_n578_1[1]),.din(w_n578_0[0]));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.doutc(w_n579_0[2]),.din(n579));
	jspl jspl_w_n580_0(.douta(w_n580_0[0]),.doutb(w_n580_0[1]),.din(w_dff_B_0BNgGgMg3_2));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl3 jspl3_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.doutc(w_n583_0[2]),.din(n583));
	jspl jspl_w_n583_1(.douta(w_n583_1[0]),.doutb(w_n583_1[1]),.din(w_n583_0[0]));
	jspl3 jspl3_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.doutc(w_n584_0[2]),.din(n584));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(w_dff_B_WDEbrLem7_2));
	jspl jspl_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.din(n586));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n589_0(.douta(w_n589_0[0]),.doutb(w_dff_A_VcZ0ObV67_1),.doutc(w_n589_0[2]),.din(n589));
	jspl jspl_w_n589_1(.douta(w_n589_1[0]),.doutb(w_n589_1[1]),.din(w_n589_0[0]));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n592_0(.douta(w_dff_A_LwVKvSsc3_0),.doutb(w_n592_0[1]),.din(n592));
	jspl jspl_w_n599_0(.douta(w_dff_A_cOrKHC8r7_0),.doutb(w_n599_0[1]),.din(n599));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl3 jspl3_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.doutc(w_n606_0[2]),.din(n606));
	jspl3 jspl3_w_n606_1(.douta(w_dff_A_8CDfmc8z6_0),.doutb(w_dff_A_sIc5B8IA5_1),.doutc(w_n606_1[2]),.din(w_n606_0[0]));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl3 jspl3_w_n608_0(.douta(w_dff_A_nv66cA3z1_0),.doutb(w_n608_0[1]),.doutc(w_n608_0[2]),.din(n608));
	jspl jspl_w_n610_0(.douta(w_dff_A_Nei84SfY4_0),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_dff_A_AeGQcbZC4_1),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.doutc(w_n615_0[2]),.din(n615));
	jspl jspl_w_n615_1(.douta(w_dff_A_KrygBMp55_0),.doutb(w_n615_1[1]),.din(w_n615_0[0]));
	jspl jspl_w_n617_0(.douta(w_n617_0[0]),.doutb(w_dff_A_6arFQ3iJ3_1),.din(n617));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(w_dff_B_an6MDwmU2_2));
	jspl jspl_w_n620_0(.douta(w_dff_A_Kir7Rrku2_0),.doutb(w_n620_0[1]),.din(n620));
	jspl3 jspl3_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.doutc(w_n621_0[2]),.din(n621));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_dff_A_QOjGnQml7_2),.din(n622));
	jspl jspl_w_n622_1(.douta(w_n622_1[0]),.doutb(w_n622_1[1]),.din(w_n622_0[0]));
	jspl3 jspl3_w_n623_0(.douta(w_n623_0[0]),.doutb(w_dff_A_hhuo9bPa3_1),.doutc(w_dff_A_82enB9Zl4_2),.din(n623));
	jspl jspl_w_n624_0(.douta(w_dff_A_xUWqSw9H1_0),.doutb(w_n624_0[1]),.din(n624));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n626_0(.douta(w_dff_A_DqfIZIe95_0),.doutb(w_n626_0[1]),.din(n626));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(w_dff_B_KqGlf3EU9_2));
	jspl jspl_w_n629_0(.douta(w_dff_A_EX3ZzQQk9_0),.doutb(w_n629_0[1]),.din(n629));
	jspl3 jspl3_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.doutc(w_n630_0[2]),.din(n630));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(w_dff_B_TLKxVHrz8_2));
	jspl jspl_w_n633_0(.douta(w_dff_A_z6Z7PJLr0_0),.doutb(w_n633_0[1]),.din(n633));
	jspl3 jspl3_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.doutc(w_n634_0[2]),.din(n634));
	jspl3 jspl3_w_n635_0(.douta(w_dff_A_U3iOSSB60_0),.doutb(w_n635_0[1]),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n637_0(.douta(w_dff_A_YBLe62Qq7_0),.doutb(w_n637_0[1]),.din(n637));
	jspl jspl_w_n642_0(.douta(w_dff_A_8nXhsAqp5_0),.doutb(w_n642_0[1]),.din(n642));
	jspl jspl_w_n643_0(.douta(w_dff_A_htWSNZ0U3_0),.doutb(w_n643_0[1]),.din(w_dff_B_64BnYiHV3_2));
	jspl3 jspl3_w_n645_0(.douta(w_dff_A_NlXmhPtA6_0),.doutb(w_dff_A_xKhpYeJo3_1),.doutc(w_n645_0[2]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(n647));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_dff_A_LnBaAuQd1_1),.doutc(w_n648_0[2]),.din(n648));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl3 jspl3_w_n653_0(.douta(w_n653_0[0]),.doutb(w_dff_A_sUtFUMxE0_1),.doutc(w_n653_0[2]),.din(n653));
	jspl jspl_w_n653_1(.douta(w_dff_A_bYH1Yk4w1_0),.doutb(w_n653_1[1]),.din(w_n653_0[0]));
	jspl jspl_w_n656_0(.douta(w_n656_0[0]),.doutb(w_dff_A_HSuaGMv20_1),.din(n656));
	jspl3 jspl3_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.doutc(w_n657_0[2]),.din(n657));
	jspl jspl_w_n657_1(.douta(w_n657_1[0]),.doutb(w_n657_1[1]),.din(w_n657_0[0]));
	jspl3 jspl3_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.doutc(w_n658_0[2]),.din(w_dff_B_VXaHy9Hx2_3));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_n660_0[2]),.din(n660));
	jspl jspl_w_n660_1(.douta(w_n660_1[0]),.doutb(w_n660_1[1]),.din(w_n660_0[0]));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_dff_A_Ivn3BrT31_1),.din(n661));
	jspl3 jspl3_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.doutc(w_n662_0[2]),.din(w_dff_B_pmxFTMoD6_3));
	jspl jspl_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.din(n663));
	jspl3 jspl3_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.doutc(w_n664_0[2]),.din(n664));
	jspl jspl_w_n664_1(.douta(w_n664_1[0]),.doutb(w_n664_1[1]),.din(w_n664_0[0]));
	jspl3 jspl3_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.doutc(w_n665_0[2]),.din(n665));
	jspl jspl_w_n666_0(.douta(w_n666_0[0]),.doutb(w_n666_0[1]),.din(w_dff_B_xceFMOFW7_2));
	jspl jspl_w_n667_0(.douta(w_dff_A_Rt6Qggwj7_0),.doutb(w_n667_0[1]),.din(n667));
	jspl3 jspl3_w_n668_0(.douta(w_n668_0[0]),.doutb(w_n668_0[1]),.doutc(w_n668_0[2]),.din(n668));
	jspl3 jspl3_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.doutc(w_n669_0[2]),.din(n669));
	jspl jspl_w_n671_0(.douta(w_n671_0[0]),.doutb(w_n671_0[1]),.din(w_dff_B_xfvM5hH19_2));
	jspl jspl_w_n672_0(.douta(w_dff_A_1aqJqf1o2_0),.doutb(w_n672_0[1]),.din(n672));
	jspl3 jspl3_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.doutc(w_n673_0[2]),.din(n673));
	jspl3 jspl3_w_n674_0(.douta(w_n674_0[0]),.doutb(w_dff_A_mzieiADk9_1),.doutc(w_n674_0[2]),.din(n674));
	jspl jspl_w_n674_1(.douta(w_dff_A_v7RfquDs0_0),.doutb(w_n674_1[1]),.din(w_n674_0[0]));
	jspl3 jspl3_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.doutc(w_n675_0[2]),.din(w_dff_B_1b42s4Cf3_3));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl3 jspl3_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.doutc(w_n677_0[2]),.din(n677));
	jspl3 jspl3_w_n678_0(.douta(w_dff_A_Hk3heCbt6_0),.doutb(w_dff_A_ksJ7tGhk9_1),.doutc(w_n678_0[2]),.din(n678));
	jspl3 jspl3_w_n679_0(.douta(w_n679_0[0]),.doutb(w_dff_A_bxt3cWg04_1),.doutc(w_dff_A_ROvKrg5y1_2),.din(n679));
	jspl jspl_w_n679_1(.douta(w_n679_1[0]),.doutb(w_n679_1[1]),.din(w_n679_0[0]));
	jspl jspl_w_n680_0(.douta(w_dff_A_bmHVwHPA3_0),.doutb(w_n680_0[1]),.din(n680));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n686_0(.douta(w_dff_A_OzFdgeut2_0),.doutb(w_n686_0[1]),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_dff_A_1IQtyevN2_1),.din(w_dff_B_FRjIx0s29_2));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_dff_A_N0r6384D1_1),.din(n692));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl3 jspl3_w_n697_0(.douta(w_dff_A_VnPbcDzP7_0),.doutb(w_dff_A_T8J0NI7b7_1),.doutc(w_n697_0[2]),.din(n697));
	jspl3 jspl3_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.doutc(w_n699_0[2]),.din(n699));
	jspl jspl_w_n699_1(.douta(w_n699_1[0]),.doutb(w_n699_1[1]),.din(w_n699_0[0]));
	jspl3 jspl3_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.doutc(w_n701_0[2]),.din(n701));
	jspl jspl_w_n701_1(.douta(w_n701_1[0]),.doutb(w_n701_1[1]),.din(w_n701_0[0]));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_dff_A_W7cqJDbd8_0),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_dff_A_DUwVtVMp5_1),.doutc(w_n707_0[2]),.din(n707));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_dff_A_93P75Fw56_1),.din(n708));
	jspl3 jspl3_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.doutc(w_n709_0[2]),.din(n709));
	jspl jspl_w_n709_1(.douta(w_n709_1[0]),.doutb(w_n709_1[1]),.din(w_n709_0[0]));
	jspl jspl_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_dff_A_2fsMJv6Z9_0),.doutb(w_n712_0[1]),.din(n712));
	jspl3 jspl3_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.doutc(w_n713_0[2]),.din(w_dff_B_FivChyJd2_3));
	jspl jspl_w_n713_1(.douta(w_n713_1[0]),.doutb(w_n713_1[1]),.din(w_n713_0[0]));
	jspl jspl_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.din(n714));
	jspl3 jspl3_w_n715_0(.douta(w_dff_A_X8KAt6jb7_0),.doutb(w_dff_A_mNktjaKO5_1),.doutc(w_n715_0[2]),.din(n715));
	jspl3 jspl3_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.doutc(w_n716_0[2]),.din(n716));
	jspl jspl_w_n716_1(.douta(w_n716_1[0]),.doutb(w_n716_1[1]),.din(w_n716_0[0]));
	jspl3 jspl3_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.doutc(w_n720_0[2]),.din(w_dff_B_fJVRGy5q8_3));
	jspl jspl_w_n720_1(.douta(w_n720_1[0]),.doutb(w_n720_1[1]),.din(w_n720_0[0]));
	jspl3 jspl3_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.doutc(w_n723_0[2]),.din(n723));
	jspl3 jspl3_w_n727_0(.douta(w_dff_A_MOHz5gvg5_0),.doutb(w_n727_0[1]),.doutc(w_n727_0[2]),.din(n727));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_dff_A_oja2GgdL4_1),.din(w_dff_B_qex5kdE77_2));
	jspl3 jspl3_w_n730_0(.douta(w_n730_0[0]),.doutb(w_n730_0[1]),.doutc(w_n730_0[2]),.din(n730));
	jspl3 jspl3_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.doutc(w_n734_0[2]),.din(n734));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_dff_A_HiQIEYI01_1),.din(w_dff_B_zZtQAI2w2_2));
	jspl3 jspl3_w_n737_0(.douta(w_dff_A_FCPrPmIm8_0),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_dff_A_WfDfgt2O1_1),.din(n742));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_n744_0[2]),.din(n744));
	jspl3 jspl3_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.doutc(w_n748_0[2]),.din(n748));
	jspl jspl_w_n751_0(.douta(w_dff_A_nSYGefZu7_0),.doutb(w_n751_0[1]),.din(n751));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl3 jspl3_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.doutc(w_n754_0[2]),.din(n754));
	jspl3 jspl3_w_n758_0(.douta(w_n758_0[0]),.doutb(w_n758_0[1]),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(n764));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_dff_A_u8gNdpKz3_1),.din(n782));
	jspl3 jspl3_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.doutc(w_n784_0[2]),.din(n784));
	jspl3 jspl3_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.doutc(w_n787_0[2]),.din(n787));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.doutc(w_n790_0[2]),.din(n790));
	jspl jspl_w_n790_1(.douta(w_n790_1[0]),.doutb(w_n790_1[1]),.din(w_n790_0[0]));
	jspl3 jspl3_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.doutc(w_n793_0[2]),.din(n793));
	jspl jspl_w_n793_1(.douta(w_n793_1[0]),.doutb(w_n793_1[1]),.din(w_n793_0[0]));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl jspl_w_n797_1(.douta(w_n797_1[0]),.doutb(w_n797_1[1]),.din(w_n797_0[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl jspl_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.din(w_n801_0[0]));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl3 jspl3_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.doutc(w_n804_0[2]),.din(n804));
	jspl3 jspl3_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.doutc(w_n807_0[2]),.din(n807));
	jspl3 jspl3_w_n810_0(.douta(w_dff_A_NdAjGV575_0),.doutb(w_n810_0[1]),.doutc(w_dff_A_n3OppnbW5_2),.din(w_dff_B_EsG6Kwdn3_3));
	jspl3 jspl3_w_n812_0(.douta(w_n812_0[0]),.doutb(w_n812_0[1]),.doutc(w_n812_0[2]),.din(n812));
	jspl3 jspl3_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.doutc(w_n816_0[2]),.din(n816));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(n817));
	jspl3 jspl3_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.doutc(w_n819_0[2]),.din(n819));
	jspl3 jspl3_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.doutc(w_n823_0[2]),.din(n823));
	jspl jspl_w_n824_0(.douta(w_dff_A_wB9sN0yI0_0),.doutb(w_n824_0[1]),.din(n824));
	jspl3 jspl3_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.doutc(w_n827_0[2]),.din(n827));
	jspl3 jspl3_w_n831_0(.douta(w_n831_0[0]),.doutb(w_n831_0[1]),.doutc(w_n831_0[2]),.din(n831));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n838_0(.douta(w_n838_0[0]),.doutb(w_n838_0[1]),.din(n838));
	jspl3 jspl3_w_n843_0(.douta(w_n843_0[0]),.doutb(w_n843_0[1]),.doutc(w_n843_0[2]),.din(n843));
	jspl3 jspl3_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.doutc(w_n847_0[2]),.din(n847));
	jspl jspl_w_n848_0(.douta(w_dff_A_KD4wimPd0_0),.doutb(w_n848_0[1]),.din(n848));
	jspl3 jspl3_w_n851_0(.douta(w_dff_A_XC64y0ZQ7_0),.doutb(w_n851_0[1]),.doutc(w_n851_0[2]),.din(n851));
	jspl3 jspl3_w_n855_0(.douta(w_dff_A_bQRHzGDs9_0),.doutb(w_n855_0[1]),.doutc(w_n855_0[2]),.din(n855));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_dff_A_YBvaUdOP4_1),.din(n856));
	jspl3 jspl3_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.doutc(w_dff_A_IUzccUPO8_2),.din(n858));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n864_0(.douta(w_dff_A_x8erXmeB9_0),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_dff_A_b3Ut7UhH7_1),.din(n865));
	jspl3 jspl3_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.doutc(w_n869_0[2]),.din(n869));
	jspl3 jspl3_w_n873_0(.douta(w_n873_0[0]),.doutb(w_dff_A_1PkpiUyh1_1),.doutc(w_dff_A_QYNBPp378_2),.din(n873));
	jspl jspl_w_n874_0(.douta(w_dff_A_kpWQCibZ0_0),.doutb(w_n874_0[1]),.din(n874));
	jspl3 jspl3_w_n878_0(.douta(w_n878_0[0]),.doutb(w_n878_0[1]),.doutc(w_n878_0[2]),.din(n878));
	jspl3 jspl3_w_n882_0(.douta(w_n882_0[0]),.doutb(w_dff_A_8QpsK7Yt1_1),.doutc(w_dff_A_5CD2Eegm4_2),.din(n882));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_dff_A_FaUhQEIr8_1),.din(n887));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl3 jspl3_w_n891_0(.douta(w_n891_0[0]),.doutb(w_dff_A_xTpTo3FQ6_1),.doutc(w_n891_0[2]),.din(n891));
	jspl jspl_w_n891_1(.douta(w_n891_1[0]),.doutb(w_n891_1[1]),.din(w_n891_0[0]));
	jspl3 jspl3_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.doutc(w_n895_0[2]),.din(n895));
	jspl jspl_w_n895_1(.douta(w_n895_1[0]),.doutb(w_n895_1[1]),.din(w_n895_0[0]));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(w_dff_B_E1vqs5So6_2));
	jspl3 jspl3_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.doutc(w_n899_0[2]),.din(n899));
	jspl3 jspl3_w_n902_0(.douta(w_n902_0[0]),.doutb(w_dff_A_Rjv8E4uC9_1),.doutc(w_dff_A_DWrTK79g5_2),.din(n902));
	jspl3 jspl3_w_n905_0(.douta(w_dff_A_DYqfH4B18_0),.doutb(w_n905_0[1]),.doutc(w_n905_0[2]),.din(w_dff_B_mUrVDMiY4_3));
	jspl3 jspl3_w_n908_0(.douta(w_n908_0[0]),.doutb(w_n908_0[1]),.doutc(w_n908_0[2]),.din(n908));
	jspl3 jspl3_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.doutc(w_n912_0[2]),.din(w_dff_B_CzetVjBx0_3));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(n913));
	jspl3 jspl3_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.doutc(w_n916_0[2]),.din(n916));
	jspl3 jspl3_w_n920_0(.douta(w_n920_0[0]),.doutb(w_dff_A_SJRSbQzT0_1),.doutc(w_dff_A_M23IpCZd7_2),.din(n920));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(n923));
	jspl3 jspl3_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.doutc(w_n927_0[2]),.din(n927));
	jspl3 jspl3_w_n931_0(.douta(w_n931_0[0]),.doutb(w_dff_A_d6l7CZCQ0_1),.doutc(w_dff_A_r5guVyE14_2),.din(n931));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_dff_A_hfnE4kP47_1),.din(n932));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n939_0(.douta(w_dff_A_Dbnl3XpI9_0),.doutb(w_n939_0[1]),.din(n939));
	jspl3 jspl3_w_n945_0(.douta(w_n945_0[0]),.doutb(w_n945_0[1]),.doutc(w_n945_0[2]),.din(n945));
	jspl jspl_w_n945_1(.douta(w_n945_1[0]),.doutb(w_n945_1[1]),.din(w_n945_0[0]));
	jspl3 jspl3_w_n948_0(.douta(w_dff_A_Omj3E1au7_0),.doutb(w_n948_0[1]),.doutc(w_dff_A_OMALyz483_2),.din(n948));
	jspl jspl_w_n948_1(.douta(w_n948_1[0]),.doutb(w_n948_1[1]),.din(w_n948_0[0]));
	jspl jspl_w_n950_0(.douta(w_n950_0[0]),.doutb(w_n950_0[1]),.din(n950));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n972_0(.douta(w_dff_A_olH5ydUu8_0),.doutb(w_n972_0[1]),.din(w_dff_B_BGQRYwhH0_2));
	jspl jspl_w_n981_0(.douta(w_dff_A_FS4dxPOV8_0),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.doutc(w_n988_0[2]),.din(n988));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_dff_A_TnOnyZIt6_1),.din(n993));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl3 jspl3_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.doutc(w_n995_0[2]),.din(n995));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.doutc(w_n999_0[2]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1003_0(.douta(w_dff_A_hFQ53zNg9_0),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.din(n1008));
	jspl3 jspl3_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.doutc(w_n1009_0[2]),.din(n1009));
	jspl jspl_w_n1009_1(.douta(w_n1009_1[0]),.doutb(w_n1009_1[1]),.din(w_n1009_0[0]));
	jspl3 jspl3_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.doutc(w_n1013_0[2]),.din(n1013));
	jspl jspl_w_n1013_1(.douta(w_n1013_1[0]),.doutb(w_n1013_1[1]),.din(w_n1013_0[0]));
	jspl jspl_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.din(n1014));
	jspl jspl_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.din(n1015));
	jspl3 jspl3_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.doutc(w_n1016_0[2]),.din(n1016));
	jspl3 jspl3_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.doutc(w_n1019_0[2]),.din(n1019));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_dff_A_QwCMM5pe6_1),.din(w_dff_B_RBqfXNkC9_2));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1044_0(.douta(w_dff_A_yVSrZYYS8_0),.doutb(w_n1044_0[1]),.din(w_dff_B_JyTawwKo8_2));
	jspl3 jspl3_w_n1061_0(.douta(w_dff_A_RBRzs81B1_0),.doutb(w_n1061_0[1]),.doutc(w_n1061_0[2]),.din(n1061));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.din(n1062));
	jspl3 jspl3_w_n1066_0(.douta(w_dff_A_Um3i6k0s2_0),.doutb(w_n1066_0[1]),.doutc(w_n1066_0[2]),.din(n1066));
	jspl jspl_w_n1068_0(.douta(w_n1068_0[0]),.doutb(w_n1068_0[1]),.din(n1068));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(n1069));
	jspl3 jspl3_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.doutc(w_n1073_0[2]),.din(n1073));
	jspl jspl_w_n1075_0(.douta(w_dff_A_wZ1bMUCk5_0),.doutb(w_n1075_0[1]),.din(n1075));
	jspl jspl_w_n1076_0(.douta(w_dff_A_v1DXBwy66_0),.doutb(w_n1076_0[1]),.din(n1076));
	jspl3 jspl3_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.doutc(w_n1077_0[2]),.din(n1077));
	jspl3 jspl3_w_n1081_0(.douta(w_n1081_0[0]),.doutb(w_n1081_0[1]),.doutc(w_n1081_0[2]),.din(n1081));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl3 jspl3_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.doutc(w_n1086_0[2]),.din(n1086));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1095_0(.douta(w_dff_A_VqC2Fu7o5_0),.doutb(w_n1095_0[1]),.din(n1095));
	jspl3 jspl3_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.doutc(w_n1096_0[2]),.din(n1096));
	jspl3 jspl3_w_n1100_0(.douta(w_n1100_0[0]),.doutb(w_n1100_0[1]),.doutc(w_n1100_0[2]),.din(n1100));
	jspl jspl_w_n1102_0(.douta(w_dff_A_W8W1Fbec0_0),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1104_0(.douta(w_n1104_0[0]),.doutb(w_dff_A_dNJIceBS3_1),.din(n1104));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.din(n1105));
	jspl jspl_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.din(n1116));
	jspl3 jspl3_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.doutc(w_n1122_0[2]),.din(n1122));
	jspl3 jspl3_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.doutc(w_n1125_0[2]),.din(w_dff_B_4GVNBzqu1_3));
	jspl jspl_w_n1127_0(.douta(w_dff_A_azqyXgUa4_0),.doutb(w_n1127_0[1]),.din(w_dff_B_pfOlVf9R1_2));
	jspl3 jspl3_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.doutc(w_n1128_0[2]),.din(n1128));
	jspl jspl_w_n1128_1(.douta(w_n1128_1[0]),.doutb(w_n1128_1[1]),.din(w_n1128_0[0]));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1136_0(.douta(w_n1136_0[0]),.doutb(w_dff_A_vpVwBZGG7_1),.din(n1136));
	jspl jspl_w_n1142_0(.douta(w_n1142_0[0]),.doutb(w_n1142_0[1]),.din(n1142));
	jspl3 jspl3_w_n1148_0(.douta(w_n1148_0[0]),.doutb(w_n1148_0[1]),.doutc(w_dff_A_ua17eETB6_2),.din(n1148));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(n1156));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(n1173));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1236_0(.douta(w_dff_A_MeVxKv7k8_0),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(n1283));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_dff_A_jov50joB5_1),.din(n1301));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl3 jspl3_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_dff_A_YU2PxwHh9_1),.doutc(w_dff_A_1fPZMeRr7_2),.din(n1359));
	jspl3 jspl3_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_dff_A_hSoXGY9p8_1),.doutc(w_n1360_0[2]),.din(n1360));
	jspl jspl_w_n1360_1(.douta(w_n1360_1[0]),.doutb(w_dff_A_5wPFBUs39_1),.din(w_n1360_0[0]));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_dff_A_cV1ghasb7_1),.din(n1361));
	jspl jspl_w_n1362_0(.douta(w_n1362_0[0]),.doutb(w_n1362_0[1]),.din(n1362));
	jspl jspl_w_n1376_0(.douta(w_dff_A_6Yzdt3Ak2_0),.doutb(w_n1376_0[1]),.din(n1376));
	jspl3 jspl3_w_n1380_0(.douta(w_n1380_0[0]),.doutb(w_dff_A_0gA4mnx75_1),.doutc(w_n1380_0[2]),.din(n1380));
	jspl jspl_w_n1380_1(.douta(w_n1380_1[0]),.doutb(w_n1380_1[1]),.din(w_n1380_0[0]));
	jspl3 jspl3_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.doutc(w_n1383_0[2]),.din(n1383));
	jspl3 jspl3_w_n1383_1(.douta(w_n1383_1[0]),.doutb(w_n1383_1[1]),.doutc(w_n1383_1[2]),.din(w_n1383_0[0]));
	jspl3 jspl3_w_n1385_0(.douta(w_n1385_0[0]),.doutb(w_n1385_0[1]),.doutc(w_n1385_0[2]),.din(n1385));
	jspl jspl_w_n1385_1(.douta(w_n1385_1[0]),.doutb(w_n1385_1[1]),.din(w_n1385_0[0]));
	jspl3 jspl3_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.doutc(w_n1389_0[2]),.din(n1389));
	jspl jspl_w_n1389_1(.douta(w_n1389_1[0]),.doutb(w_n1389_1[1]),.din(w_n1389_0[0]));
	jspl3 jspl3_w_n1392_0(.douta(w_n1392_0[0]),.doutb(w_n1392_0[1]),.doutc(w_n1392_0[2]),.din(n1392));
	jspl jspl_w_n1392_1(.douta(w_n1392_1[0]),.doutb(w_n1392_1[1]),.din(w_n1392_0[0]));
	jspl jspl_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_dff_A_HnnnsTka4_1),.din(w_dff_B_WUarIzIc6_2));
	jspl jspl_w_n1402_0(.douta(w_dff_A_rQDQa0fV1_0),.doutb(w_n1402_0[1]),.din(w_dff_B_zDz5HAab4_2));
	jspl jspl_w_n1403_0(.douta(w_dff_A_U5A0OWvQ2_0),.doutb(w_n1403_0[1]),.din(w_dff_B_0l4IU0o40_2));
	jspl jspl_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_dff_A_SuUZyTFP8_1),.din(w_dff_B_KlXKBtaX3_2));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl jspl_w_n1406_0(.douta(w_n1406_0[0]),.doutb(w_n1406_0[1]),.din(n1406));
	jspl jspl_w_n1414_0(.douta(w_n1414_0[0]),.doutb(w_dff_A_gQJETuFf1_1),.din(n1414));
	jspl3 jspl3_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_dff_A_hJn7yT7j7_1),.doutc(w_dff_A_t7v2Foso9_2),.din(w_dff_B_prn8QpJd1_3));
	jspl jspl_w_n1421_0(.douta(w_dff_A_D6vLbTgQ8_0),.doutb(w_n1421_0[1]),.din(w_dff_B_6nDF9O8S7_2));
	jspl jspl_w_n1422_0(.douta(w_dff_A_0Tg0GVpc8_0),.doutb(w_n1422_0[1]),.din(w_dff_B_Hq71TNA62_2));
	jspl jspl_w_n1424_0(.douta(w_n1424_0[0]),.doutb(w_n1424_0[1]),.din(n1424));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl3 jspl3_w_n1444_0(.douta(w_dff_A_tj41q6wh8_0),.doutb(w_n1444_0[1]),.doutc(w_dff_A_dlooAmvU0_2),.din(w_dff_B_SI0CUn5e3_3));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_dff_A_vE50oDBr4_1),.din(w_dff_B_UthSIp5O4_2));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_dff_A_uX2DG70z2_1),.din(w_dff_B_2jMqZwdh5_2));
	jspl3 jspl3_w_n1463_0(.douta(w_dff_A_ZxbK0vmW0_0),.doutb(w_dff_A_RGme1VQO3_1),.doutc(w_n1463_0[2]),.din(n1463));
	jspl jspl_w_n1464_0(.douta(w_n1464_0[0]),.doutb(w_dff_A_ykPomkwX5_1),.din(w_dff_B_2rNbrDSn7_2));
	jspl jspl_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.din(n1465));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_dff_A_vaUUkInl2_1),.din(w_dff_B_jllnJNpC9_2));
	jspl jspl_w_n1469_0(.douta(w_dff_A_lX3g4Itf2_0),.doutb(w_n1469_0[1]),.din(w_dff_B_R8RVR4Em2_2));
	jspl jspl_w_n1470_0(.douta(w_dff_A_ltbWdfQG3_0),.doutb(w_n1470_0[1]),.din(w_dff_B_EsLk7yv80_2));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_dff_A_pJKJ5JGS9_1),.din(n1471));
	jspl jspl_w_n1472_0(.douta(w_n1472_0[0]),.doutb(w_n1472_0[1]),.din(n1472));
	jspl jspl_w_n1473_0(.douta(w_n1473_0[0]),.doutb(w_n1473_0[1]),.din(n1473));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_dff_A_KtsyxYg13_1),.din(n1479));
	jspl jspl_w_n1482_0(.douta(w_n1482_0[0]),.doutb(w_dff_A_0WAxktpG4_1),.din(n1482));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(n1486));
	jspl3 jspl3_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.doutc(w_dff_A_IGyUEtNS0_2),.din(n1494));
	jspl jspl_w_n1501_0(.douta(w_n1501_0[0]),.doutb(w_dff_A_iatti9uZ2_1),.din(n1501));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_dff_A_kUmEGgAQ2_1),.din(n1520));
	jspl jspl_w_n1536_0(.douta(w_n1536_0[0]),.doutb(w_n1536_0[1]),.din(n1536));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(n1571));
	jspl jspl_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(w_dff_B_2ZlPMjFp5_2));
	jspl jspl_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.din(n1611));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl jspl_w_n1642_0(.douta(w_n1642_0[0]),.doutb(w_n1642_0[1]),.din(n1642));
	jspl jspl_w_n1644_0(.douta(w_dff_A_N99NFegW8_0),.doutb(w_n1644_0[1]),.din(n1644));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_dff_A_bMRYvsgy9_1),.din(n1651));
	jspl jspl_w_n1654_0(.douta(w_n1654_0[0]),.doutb(w_dff_A_0WhToFMW5_1),.din(n1654));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1667_0(.douta(w_dff_A_ZPEdoOs90_0),.doutb(w_n1667_0[1]),.din(n1667));
	jspl jspl_w_n1670_0(.douta(w_n1670_0[0]),.doutb(w_n1670_0[1]),.din(n1670));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(n1672));
	jspl jspl_w_n1675_0(.douta(w_n1675_0[0]),.doutb(w_dff_A_4DWiGXIG0_1),.din(n1675));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_dff_A_ybqhCZ7i9_1),.din(n1687));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(n1689));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(n1699));
	jdff dff_A_H1x1fNcX7_0(.dout(w_G5_1[0]),.din(w_dff_A_H1x1fNcX7_0),.clk(gclk));
	jdff dff_A_LJ5eExnU7_0(.dout(w_dff_A_H1x1fNcX7_0),.din(w_dff_A_LJ5eExnU7_0),.clk(gclk));
	jdff dff_A_2Rxoc2Fc8_1(.dout(w_G5_1[1]),.din(w_dff_A_2Rxoc2Fc8_1),.clk(gclk));
	jdff dff_A_DJsdh6RM2_1(.dout(w_G5_0[1]),.din(w_dff_A_DJsdh6RM2_1),.clk(gclk));
	jdff dff_A_Csyy1rkH6_1(.dout(w_dff_A_DJsdh6RM2_1),.din(w_dff_A_Csyy1rkH6_1),.clk(gclk));
	jdff dff_A_FaHfh2fO1_2(.dout(w_G5_0[2]),.din(w_dff_A_FaHfh2fO1_2),.clk(gclk));
	jdff dff_B_aOYLngUM6_0(.din(n1131),.dout(w_dff_B_aOYLngUM6_0),.clk(gclk));
	jdff dff_B_8GT5GJoe7_3(.din(n1125),.dout(w_dff_B_8GT5GJoe7_3),.clk(gclk));
	jdff dff_B_Fh6oaYhI2_3(.din(w_dff_B_8GT5GJoe7_3),.dout(w_dff_B_Fh6oaYhI2_3),.clk(gclk));
	jdff dff_B_PdMoONtd1_3(.din(w_dff_B_Fh6oaYhI2_3),.dout(w_dff_B_PdMoONtd1_3),.clk(gclk));
	jdff dff_B_p4BRydNP0_3(.din(w_dff_B_PdMoONtd1_3),.dout(w_dff_B_p4BRydNP0_3),.clk(gclk));
	jdff dff_B_ZthGTssf3_3(.din(w_dff_B_p4BRydNP0_3),.dout(w_dff_B_ZthGTssf3_3),.clk(gclk));
	jdff dff_B_o9rZ0ppE2_3(.din(w_dff_B_ZthGTssf3_3),.dout(w_dff_B_o9rZ0ppE2_3),.clk(gclk));
	jdff dff_B_uBKdNDcH8_3(.din(w_dff_B_o9rZ0ppE2_3),.dout(w_dff_B_uBKdNDcH8_3),.clk(gclk));
	jdff dff_B_Obt8tKE48_3(.din(w_dff_B_uBKdNDcH8_3),.dout(w_dff_B_Obt8tKE48_3),.clk(gclk));
	jdff dff_B_1hfgjHjp7_3(.din(w_dff_B_Obt8tKE48_3),.dout(w_dff_B_1hfgjHjp7_3),.clk(gclk));
	jdff dff_B_pSXeCuZx2_3(.din(w_dff_B_1hfgjHjp7_3),.dout(w_dff_B_pSXeCuZx2_3),.clk(gclk));
	jdff dff_B_SkkVDdcH5_3(.din(w_dff_B_pSXeCuZx2_3),.dout(w_dff_B_SkkVDdcH5_3),.clk(gclk));
	jdff dff_B_oos6ncU33_3(.din(w_dff_B_SkkVDdcH5_3),.dout(w_dff_B_oos6ncU33_3),.clk(gclk));
	jdff dff_B_aX6FGgSH8_3(.din(w_dff_B_oos6ncU33_3),.dout(w_dff_B_aX6FGgSH8_3),.clk(gclk));
	jdff dff_B_2zK51HxV0_3(.din(w_dff_B_aX6FGgSH8_3),.dout(w_dff_B_2zK51HxV0_3),.clk(gclk));
	jdff dff_B_dPUIaYT13_3(.din(w_dff_B_2zK51HxV0_3),.dout(w_dff_B_dPUIaYT13_3),.clk(gclk));
	jdff dff_B_4GVNBzqu1_3(.din(w_dff_B_dPUIaYT13_3),.dout(w_dff_B_4GVNBzqu1_3),.clk(gclk));
	jdff dff_B_nmwzeh3H7_1(.din(n1123),.dout(w_dff_B_nmwzeh3H7_1),.clk(gclk));
	jdff dff_B_zluYwsbb9_0(.din(n1121),.dout(w_dff_B_zluYwsbb9_0),.clk(gclk));
	jdff dff_B_kmsBd3pO9_0(.din(w_dff_B_zluYwsbb9_0),.dout(w_dff_B_kmsBd3pO9_0),.clk(gclk));
	jdff dff_B_LJchpJ413_0(.din(w_dff_B_kmsBd3pO9_0),.dout(w_dff_B_LJchpJ413_0),.clk(gclk));
	jdff dff_B_ZknSM7Q69_0(.din(w_dff_B_LJchpJ413_0),.dout(w_dff_B_ZknSM7Q69_0),.clk(gclk));
	jdff dff_B_tPUdWo8h1_0(.din(w_dff_B_ZknSM7Q69_0),.dout(w_dff_B_tPUdWo8h1_0),.clk(gclk));
	jdff dff_B_Jg7oXZfN3_0(.din(w_dff_B_tPUdWo8h1_0),.dout(w_dff_B_Jg7oXZfN3_0),.clk(gclk));
	jdff dff_B_O9PQ5rko9_0(.din(w_dff_B_Jg7oXZfN3_0),.dout(w_dff_B_O9PQ5rko9_0),.clk(gclk));
	jdff dff_B_IKeI7tOk1_0(.din(w_dff_B_O9PQ5rko9_0),.dout(w_dff_B_IKeI7tOk1_0),.clk(gclk));
	jdff dff_B_eaos86KW9_0(.din(w_dff_B_IKeI7tOk1_0),.dout(w_dff_B_eaos86KW9_0),.clk(gclk));
	jdff dff_B_CmYdmzaQ9_0(.din(n1120),.dout(w_dff_B_CmYdmzaQ9_0),.clk(gclk));
	jdff dff_B_RqVXRd1E5_0(.din(w_dff_B_CmYdmzaQ9_0),.dout(w_dff_B_RqVXRd1E5_0),.clk(gclk));
	jdff dff_B_PlJ4JVtI2_0(.din(w_dff_B_RqVXRd1E5_0),.dout(w_dff_B_PlJ4JVtI2_0),.clk(gclk));
	jdff dff_B_xZjP3xbI8_0(.din(n1119),.dout(w_dff_B_xZjP3xbI8_0),.clk(gclk));
	jdff dff_B_rgTnpi6f8_0(.din(n1110),.dout(w_dff_B_rgTnpi6f8_0),.clk(gclk));
	jdff dff_B_5b8wHGdI0_0(.din(w_dff_B_rgTnpi6f8_0),.dout(w_dff_B_5b8wHGdI0_0),.clk(gclk));
	jdff dff_B_cx1mKahK3_0(.din(w_dff_B_5b8wHGdI0_0),.dout(w_dff_B_cx1mKahK3_0),.clk(gclk));
	jdff dff_B_sOzLRDlF8_0(.din(w_dff_B_cx1mKahK3_0),.dout(w_dff_B_sOzLRDlF8_0),.clk(gclk));
	jdff dff_B_RPVfbBDI2_0(.din(w_dff_B_sOzLRDlF8_0),.dout(w_dff_B_RPVfbBDI2_0),.clk(gclk));
	jdff dff_B_lbPZEWeQ2_0(.din(w_dff_B_RPVfbBDI2_0),.dout(w_dff_B_lbPZEWeQ2_0),.clk(gclk));
	jdff dff_B_YzKhEAQz8_0(.din(w_dff_B_lbPZEWeQ2_0),.dout(w_dff_B_YzKhEAQz8_0),.clk(gclk));
	jdff dff_B_sybW8anM3_0(.din(w_dff_B_YzKhEAQz8_0),.dout(w_dff_B_sybW8anM3_0),.clk(gclk));
	jdff dff_B_LoxfYKrX8_1(.din(n1089),.dout(w_dff_B_LoxfYKrX8_1),.clk(gclk));
	jdff dff_B_Taz8ROiW9_1(.din(w_dff_B_LoxfYKrX8_1),.dout(w_dff_B_Taz8ROiW9_1),.clk(gclk));
	jdff dff_B_ucUW0KpF7_1(.din(n1093),.dout(w_dff_B_ucUW0KpF7_1),.clk(gclk));
	jdff dff_A_dNJIceBS3_1(.dout(w_n1104_0[1]),.din(w_dff_A_dNJIceBS3_1),.clk(gclk));
	jdff dff_A_W8W1Fbec0_0(.dout(w_n1102_0[0]),.din(w_dff_A_W8W1Fbec0_0),.clk(gclk));
	jdff dff_A_JEJp4n9Z2_0(.dout(w_n1075_0[0]),.din(w_dff_A_JEJp4n9Z2_0),.clk(gclk));
	jdff dff_A_wZ1bMUCk5_0(.dout(w_dff_A_JEJp4n9Z2_0),.din(w_dff_A_wZ1bMUCk5_0),.clk(gclk));
	jdff dff_B_clBketc26_0(.din(n1059),.dout(w_dff_B_clBketc26_0),.clk(gclk));
	jdff dff_B_owubJqtn6_0(.din(w_dff_B_clBketc26_0),.dout(w_dff_B_owubJqtn6_0),.clk(gclk));
	jdff dff_B_uGdKD9RF0_0(.din(n1058),.dout(w_dff_B_uGdKD9RF0_0),.clk(gclk));
	jdff dff_B_3YcnjEPM0_0(.din(w_dff_B_uGdKD9RF0_0),.dout(w_dff_B_3YcnjEPM0_0),.clk(gclk));
	jdff dff_B_Ke6pguCj6_0(.din(w_dff_B_3YcnjEPM0_0),.dout(w_dff_B_Ke6pguCj6_0),.clk(gclk));
	jdff dff_B_Qusatsm47_0(.din(w_dff_B_Ke6pguCj6_0),.dout(w_dff_B_Qusatsm47_0),.clk(gclk));
	jdff dff_B_xLARylk14_0(.din(n1057),.dout(w_dff_B_xLARylk14_0),.clk(gclk));
	jdff dff_B_Y78YgRbs9_0(.din(n1050),.dout(w_dff_B_Y78YgRbs9_0),.clk(gclk));
	jdff dff_B_Szp1HVeJ0_0(.din(w_dff_B_Y78YgRbs9_0),.dout(w_dff_B_Szp1HVeJ0_0),.clk(gclk));
	jdff dff_B_yrJTjGSX8_0(.din(n1047),.dout(w_dff_B_yrJTjGSX8_0),.clk(gclk));
	jdff dff_A_wKweXwCq6_1(.dout(w_n1022_0[1]),.din(w_dff_A_wKweXwCq6_1),.clk(gclk));
	jdff dff_A_JYNCkgNE3_1(.dout(w_dff_A_wKweXwCq6_1),.din(w_dff_A_JYNCkgNE3_1),.clk(gclk));
	jdff dff_A_29vt0Iai6_1(.dout(w_dff_A_JYNCkgNE3_1),.din(w_dff_A_29vt0Iai6_1),.clk(gclk));
	jdff dff_A_upaUkcFz2_1(.dout(w_dff_A_29vt0Iai6_1),.din(w_dff_A_upaUkcFz2_1),.clk(gclk));
	jdff dff_A_xwS9Vmph3_1(.dout(w_dff_A_upaUkcFz2_1),.din(w_dff_A_xwS9Vmph3_1),.clk(gclk));
	jdff dff_A_QwCMM5pe6_1(.dout(w_dff_A_xwS9Vmph3_1),.din(w_dff_A_QwCMM5pe6_1),.clk(gclk));
	jdff dff_B_RBqfXNkC9_2(.din(n1022),.dout(w_dff_B_RBqfXNkC9_2),.clk(gclk));
	jdff dff_B_M2eV6rMb1_0(.din(n1021),.dout(w_dff_B_M2eV6rMb1_0),.clk(gclk));
	jdff dff_B_fECzl2j29_0(.din(w_dff_B_M2eV6rMb1_0),.dout(w_dff_B_fECzl2j29_0),.clk(gclk));
	jdff dff_B_A2vgLadr0_0(.din(n1005),.dout(w_dff_B_A2vgLadr0_0),.clk(gclk));
	jdff dff_A_1Do7kB6g2_0(.dout(w_n1003_0[0]),.din(w_dff_A_1Do7kB6g2_0),.clk(gclk));
	jdff dff_A_hFQ53zNg9_0(.dout(w_dff_A_1Do7kB6g2_0),.din(w_dff_A_hFQ53zNg9_0),.clk(gclk));
	jdff dff_A_TnOnyZIt6_1(.dout(w_n993_0[1]),.din(w_dff_A_TnOnyZIt6_1),.clk(gclk));
	jdff dff_B_vsnB5BLX1_1(.din(n768),.dout(w_dff_B_vsnB5BLX1_1),.clk(gclk));
	jdff dff_B_Hlblfcs99_1(.din(w_dff_B_vsnB5BLX1_1),.dout(w_dff_B_Hlblfcs99_1),.clk(gclk));
	jdff dff_B_CF1uAkos3_1(.din(w_dff_B_Hlblfcs99_1),.dout(w_dff_B_CF1uAkos3_1),.clk(gclk));
	jdff dff_B_omwt6g2n2_1(.din(w_dff_B_CF1uAkos3_1),.dout(w_dff_B_omwt6g2n2_1),.clk(gclk));
	jdff dff_B_zEB8zR890_0(.din(n983),.dout(w_dff_B_zEB8zR890_0),.clk(gclk));
	jdff dff_B_X0fm0r7M0_0(.din(w_dff_B_zEB8zR890_0),.dout(w_dff_B_X0fm0r7M0_0),.clk(gclk));
	jdff dff_A_b3Ut7UhH7_1(.dout(w_n865_0[1]),.din(w_dff_A_b3Ut7UhH7_1),.clk(gclk));
	jdff dff_A_op38Mzqe5_1(.dout(w_n782_0[1]),.din(w_dff_A_op38Mzqe5_1),.clk(gclk));
	jdff dff_A_uxOA9Led6_1(.dout(w_dff_A_op38Mzqe5_1),.din(w_dff_A_uxOA9Led6_1),.clk(gclk));
	jdff dff_A_TXy3bDe50_1(.dout(w_dff_A_uxOA9Led6_1),.din(w_dff_A_TXy3bDe50_1),.clk(gclk));
	jdff dff_A_u8gNdpKz3_1(.dout(w_dff_A_TXy3bDe50_1),.din(w_dff_A_u8gNdpKz3_1),.clk(gclk));
	jdff dff_B_NjHQMahz2_1(.din(n774),.dout(w_dff_B_NjHQMahz2_1),.clk(gclk));
	jdff dff_B_UQ2eWhvW8_0(.din(n776),.dout(w_dff_B_UQ2eWhvW8_0),.clk(gclk));
	jdff dff_B_rz3yo8bX1_0(.din(n766),.dout(w_dff_B_rz3yo8bX1_0),.clk(gclk));
	jdff dff_B_pgl8Hcza8_0(.din(w_dff_B_rz3yo8bX1_0),.dout(w_dff_B_pgl8Hcza8_0),.clk(gclk));
	jdff dff_B_iEn66Zu24_0(.din(w_dff_B_pgl8Hcza8_0),.dout(w_dff_B_iEn66Zu24_0),.clk(gclk));
	jdff dff_A_9oY2BN3F2_0(.dout(w_n751_0[0]),.din(w_dff_A_9oY2BN3F2_0),.clk(gclk));
	jdff dff_A_nSYGefZu7_0(.dout(w_dff_A_9oY2BN3F2_0),.din(w_dff_A_nSYGefZu7_0),.clk(gclk));
	jdff dff_A_YZHuPk2K1_1(.dout(w_n742_0[1]),.din(w_dff_A_YZHuPk2K1_1),.clk(gclk));
	jdff dff_A_WfDfgt2O1_1(.dout(w_dff_A_YZHuPk2K1_1),.din(w_dff_A_WfDfgt2O1_1),.clk(gclk));
	jdff dff_A_F4VMf2ru8_1(.dout(w_n735_0[1]),.din(w_dff_A_F4VMf2ru8_1),.clk(gclk));
	jdff dff_A_HiQIEYI01_1(.dout(w_dff_A_F4VMf2ru8_1),.din(w_dff_A_HiQIEYI01_1),.clk(gclk));
	jdff dff_B_zZtQAI2w2_2(.din(n735),.dout(w_dff_B_zZtQAI2w2_2),.clk(gclk));
	jdff dff_A_9nUYdiC35_1(.dout(w_n728_0[1]),.din(w_dff_A_9nUYdiC35_1),.clk(gclk));
	jdff dff_A_jmBMnJRL4_1(.dout(w_dff_A_9nUYdiC35_1),.din(w_dff_A_jmBMnJRL4_1),.clk(gclk));
	jdff dff_A_c7cyeEG07_1(.dout(w_dff_A_jmBMnJRL4_1),.din(w_dff_A_c7cyeEG07_1),.clk(gclk));
	jdff dff_A_oja2GgdL4_1(.dout(w_dff_A_c7cyeEG07_1),.din(w_dff_A_oja2GgdL4_1),.clk(gclk));
	jdff dff_B_qex5kdE77_2(.din(n728),.dout(w_dff_B_qex5kdE77_2),.clk(gclk));
	jdff dff_B_E2BqAmmD6_1(.din(n1024),.dout(w_dff_B_E2BqAmmD6_1),.clk(gclk));
	jdff dff_B_hlUP6DoB9_1(.din(w_dff_B_E2BqAmmD6_1),.dout(w_dff_B_hlUP6DoB9_1),.clk(gclk));
	jdff dff_B_gUT1FJ6E2_1(.din(w_dff_B_hlUP6DoB9_1),.dout(w_dff_B_gUT1FJ6E2_1),.clk(gclk));
	jdff dff_B_VebpQi8Y0_1(.din(w_dff_B_gUT1FJ6E2_1),.dout(w_dff_B_VebpQi8Y0_1),.clk(gclk));
	jdff dff_B_Iv8egv9x3_0(.din(n1031),.dout(w_dff_B_Iv8egv9x3_0),.clk(gclk));
	jdff dff_B_QS8e2wgJ2_0(.din(w_dff_B_Iv8egv9x3_0),.dout(w_dff_B_QS8e2wgJ2_0),.clk(gclk));
	jdff dff_B_0r9OQegj7_0(.din(n1028),.dout(w_dff_B_0r9OQegj7_0),.clk(gclk));
	jdff dff_B_cf8N8jNw3_1(.din(n934),.dout(w_dff_B_cf8N8jNw3_1),.clk(gclk));
	jdff dff_B_hzR408JK2_1(.din(n942),.dout(w_dff_B_hzR408JK2_1),.clk(gclk));
	jdff dff_B_dHwOYEWc2_1(.din(n949),.dout(w_dff_B_dHwOYEWc2_1),.clk(gclk));
	jdff dff_B_jbgvIvE76_1(.din(w_dff_B_dHwOYEWc2_1),.dout(w_dff_B_jbgvIvE76_1),.clk(gclk));
	jdff dff_B_gUelUwAH4_1(.din(n938),.dout(w_dff_B_gUelUwAH4_1),.clk(gclk));
	jdff dff_B_DjlADNOI5_1(.din(w_dff_B_gUelUwAH4_1),.dout(w_dff_B_DjlADNOI5_1),.clk(gclk));
	jdff dff_B_Jfuhpsui9_1(.din(G89),.dout(w_dff_B_Jfuhpsui9_1),.clk(gclk));
	jdff dff_B_vti9Bbka6_1(.din(w_dff_B_Jfuhpsui9_1),.dout(w_dff_B_vti9Bbka6_1),.clk(gclk));
	jdff dff_B_K6n9Gu5M3_1(.din(w_dff_B_vti9Bbka6_1),.dout(w_dff_B_K6n9Gu5M3_1),.clk(gclk));
	jdff dff_B_oKPFqOOM6_1(.din(w_dff_B_K6n9Gu5M3_1),.dout(w_dff_B_oKPFqOOM6_1),.clk(gclk));
	jdff dff_B_zGP8pgHY2_1(.din(w_dff_B_oKPFqOOM6_1),.dout(w_dff_B_zGP8pgHY2_1),.clk(gclk));
	jdff dff_A_Dbnl3XpI9_0(.dout(w_n939_0[0]),.din(w_dff_A_Dbnl3XpI9_0),.clk(gclk));
	jdff dff_B_La6IPfwy8_1(.din(n922),.dout(w_dff_B_La6IPfwy8_1),.clk(gclk));
	jdff dff_A_hfnE4kP47_1(.dout(w_n932_0[1]),.din(w_dff_A_hfnE4kP47_1),.clk(gclk));
	jdff dff_A_DYqfH4B18_0(.dout(w_n905_0[0]),.din(w_dff_A_DYqfH4B18_0),.clk(gclk));
	jdff dff_B_mUrVDMiY4_3(.din(n905),.dout(w_dff_B_mUrVDMiY4_3),.clk(gclk));
	jdff dff_B_NunZNfAB4_0(.din(n904),.dout(w_dff_B_NunZNfAB4_0),.clk(gclk));
	jdff dff_B_UPaggQHO7_0(.din(w_dff_B_NunZNfAB4_0),.dout(w_dff_B_UPaggQHO7_0),.clk(gclk));
	jdff dff_A_yVSrZYYS8_0(.dout(w_n1044_0[0]),.din(w_dff_A_yVSrZYYS8_0),.clk(gclk));
	jdff dff_B_JyTawwKo8_2(.din(n1044),.dout(w_dff_B_JyTawwKo8_2),.clk(gclk));
	jdff dff_B_73b3XT5p2_0(.din(n1043),.dout(w_dff_B_73b3XT5p2_0),.clk(gclk));
	jdff dff_B_yYE49MnY2_0(.din(n1040),.dout(w_dff_B_yYE49MnY2_0),.clk(gclk));
	jdff dff_B_bSp9X1LY2_0(.din(n1038),.dout(w_dff_B_bSp9X1LY2_0),.clk(gclk));
	jdff dff_B_Crt9Bh7Q1_0(.din(n1036),.dout(w_dff_B_Crt9Bh7Q1_0),.clk(gclk));
	jdff dff_B_ipreZXo37_0(.din(w_dff_B_Crt9Bh7Q1_0),.dout(w_dff_B_ipreZXo37_0),.clk(gclk));
	jdff dff_B_E1vqs5So6_2(.din(n896),.dout(w_dff_B_E1vqs5So6_2),.clk(gclk));
	jdff dff_A_FaUhQEIr8_1(.dout(w_n887_0[1]),.din(w_dff_A_FaUhQEIr8_1),.clk(gclk));
	jdff dff_B_oyvPw3HP8_0(.din(n883),.dout(w_dff_B_oyvPw3HP8_0),.clk(gclk));
	jdff dff_A_uSouiXpl1_0(.dout(w_n874_0[0]),.din(w_dff_A_uSouiXpl1_0),.clk(gclk));
	jdff dff_A_kpWQCibZ0_0(.dout(w_dff_A_uSouiXpl1_0),.din(w_dff_A_kpWQCibZ0_0),.clk(gclk));
	jdff dff_A_KeBEqL1b9_0(.dout(w_n864_0[0]),.din(w_dff_A_KeBEqL1b9_0),.clk(gclk));
	jdff dff_A_eXNx4TLQ8_0(.dout(w_dff_A_KeBEqL1b9_0),.din(w_dff_A_eXNx4TLQ8_0),.clk(gclk));
	jdff dff_A_7geiDjfL8_0(.dout(w_dff_A_eXNx4TLQ8_0),.din(w_dff_A_7geiDjfL8_0),.clk(gclk));
	jdff dff_A_x8erXmeB9_0(.dout(w_dff_A_7geiDjfL8_0),.din(w_dff_A_x8erXmeB9_0),.clk(gclk));
	jdff dff_B_olKMC4kn6_1(.din(n837),.dout(w_dff_B_olKMC4kn6_1),.clk(gclk));
	jdff dff_B_BB9j9eEC6_1(.din(n841),.dout(w_dff_B_BB9j9eEC6_1),.clk(gclk));
	jdff dff_B_eyGmmzk53_0(.din(n840),.dout(w_dff_B_eyGmmzk53_0),.clk(gclk));
	jdff dff_B_hc7iIvA21_1(.din(n825),.dout(w_dff_B_hc7iIvA21_1),.clk(gclk));
	jdff dff_A_4emVkdrr4_0(.dout(w_n981_0[0]),.din(w_dff_A_4emVkdrr4_0),.clk(gclk));
	jdff dff_A_34VAu1QY2_0(.dout(w_dff_A_4emVkdrr4_0),.din(w_dff_A_34VAu1QY2_0),.clk(gclk));
	jdff dff_A_ZsIGRV5g6_0(.dout(w_dff_A_34VAu1QY2_0),.din(w_dff_A_ZsIGRV5g6_0),.clk(gclk));
	jdff dff_A_DxoGZ2jD9_0(.dout(w_dff_A_ZsIGRV5g6_0),.din(w_dff_A_DxoGZ2jD9_0),.clk(gclk));
	jdff dff_A_KOtvCfEw3_0(.dout(w_dff_A_DxoGZ2jD9_0),.din(w_dff_A_KOtvCfEw3_0),.clk(gclk));
	jdff dff_A_FS4dxPOV8_0(.dout(w_dff_A_KOtvCfEw3_0),.din(w_dff_A_FS4dxPOV8_0),.clk(gclk));
	jdff dff_B_BaWeFQ4N1_0(.din(n980),.dout(w_dff_B_BaWeFQ4N1_0),.clk(gclk));
	jdff dff_A_KD4wimPd0_0(.dout(w_n848_0[0]),.din(w_dff_A_KD4wimPd0_0),.clk(gclk));
	jdff dff_A_IUzccUPO8_2(.dout(w_n858_0[2]),.din(w_dff_A_IUzccUPO8_2),.clk(gclk));
	jdff dff_A_YBvaUdOP4_1(.dout(w_n856_0[1]),.din(w_dff_A_YBvaUdOP4_1),.clk(gclk));
	jdff dff_A_wB9sN0yI0_0(.dout(w_n824_0[0]),.din(w_dff_A_wB9sN0yI0_0),.clk(gclk));
	jdff dff_A_cZ3tvlSy3_0(.dout(w_n810_0[0]),.din(w_dff_A_cZ3tvlSy3_0),.clk(gclk));
	jdff dff_A_30epYld30_0(.dout(w_dff_A_cZ3tvlSy3_0),.din(w_dff_A_30epYld30_0),.clk(gclk));
	jdff dff_A_tK5Ktzi97_0(.dout(w_dff_A_30epYld30_0),.din(w_dff_A_tK5Ktzi97_0),.clk(gclk));
	jdff dff_A_tNzfigGw5_0(.dout(w_dff_A_tK5Ktzi97_0),.din(w_dff_A_tNzfigGw5_0),.clk(gclk));
	jdff dff_A_M6GKYzr27_0(.dout(w_dff_A_tNzfigGw5_0),.din(w_dff_A_M6GKYzr27_0),.clk(gclk));
	jdff dff_A_yE9Belt04_0(.dout(w_dff_A_M6GKYzr27_0),.din(w_dff_A_yE9Belt04_0),.clk(gclk));
	jdff dff_A_NdAjGV575_0(.dout(w_dff_A_yE9Belt04_0),.din(w_dff_A_NdAjGV575_0),.clk(gclk));
	jdff dff_A_n3OppnbW5_2(.dout(w_n810_0[2]),.din(w_dff_A_n3OppnbW5_2),.clk(gclk));
	jdff dff_B_0A8unDCZ9_3(.din(n810),.dout(w_dff_B_0A8unDCZ9_3),.clk(gclk));
	jdff dff_B_EsG6Kwdn3_3(.din(w_dff_B_0A8unDCZ9_3),.dout(w_dff_B_EsG6Kwdn3_3),.clk(gclk));
	jdff dff_A_BxmbYe4G3_0(.dout(w_n972_0[0]),.din(w_dff_A_BxmbYe4G3_0),.clk(gclk));
	jdff dff_A_vxfEyPsa7_0(.dout(w_dff_A_BxmbYe4G3_0),.din(w_dff_A_vxfEyPsa7_0),.clk(gclk));
	jdff dff_A_DoJtKWku7_0(.dout(w_dff_A_vxfEyPsa7_0),.din(w_dff_A_DoJtKWku7_0),.clk(gclk));
	jdff dff_A_wblS193s2_0(.dout(w_dff_A_DoJtKWku7_0),.din(w_dff_A_wblS193s2_0),.clk(gclk));
	jdff dff_A_ioM7agik6_0(.dout(w_dff_A_wblS193s2_0),.din(w_dff_A_ioM7agik6_0),.clk(gclk));
	jdff dff_A_a30oBt2Z5_0(.dout(w_dff_A_ioM7agik6_0),.din(w_dff_A_a30oBt2Z5_0),.clk(gclk));
	jdff dff_A_olH5ydUu8_0(.dout(w_dff_A_a30oBt2Z5_0),.din(w_dff_A_olH5ydUu8_0),.clk(gclk));
	jdff dff_B_BGQRYwhH0_2(.din(n972),.dout(w_dff_B_BGQRYwhH0_2),.clk(gclk));
	jdff dff_B_ocApAAlI3_1(.din(n962),.dout(w_dff_B_ocApAAlI3_1),.clk(gclk));
	jdff dff_B_hntVSUkP1_1(.din(n963),.dout(w_dff_B_hntVSUkP1_1),.clk(gclk));
	jdff dff_B_HRf6BwCS8_1(.din(w_dff_B_hntVSUkP1_1),.dout(w_dff_B_HRf6BwCS8_1),.clk(gclk));
	jdff dff_A_rQDQa0fV1_0(.dout(w_n1402_0[0]),.din(w_dff_A_rQDQa0fV1_0),.clk(gclk));
	jdff dff_B_Qcden2jP5_2(.din(n1402),.dout(w_dff_B_Qcden2jP5_2),.clk(gclk));
	jdff dff_B_VOOtMusF2_2(.din(w_dff_B_Qcden2jP5_2),.dout(w_dff_B_VOOtMusF2_2),.clk(gclk));
	jdff dff_B_IblNFaSL7_2(.din(w_dff_B_VOOtMusF2_2),.dout(w_dff_B_IblNFaSL7_2),.clk(gclk));
	jdff dff_B_KxNlxfcE2_2(.din(w_dff_B_IblNFaSL7_2),.dout(w_dff_B_KxNlxfcE2_2),.clk(gclk));
	jdff dff_B_x5jDJCzn2_2(.din(w_dff_B_KxNlxfcE2_2),.dout(w_dff_B_x5jDJCzn2_2),.clk(gclk));
	jdff dff_B_RwQl9RZp8_2(.din(w_dff_B_x5jDJCzn2_2),.dout(w_dff_B_RwQl9RZp8_2),.clk(gclk));
	jdff dff_B_wQV5JdOo7_2(.din(w_dff_B_RwQl9RZp8_2),.dout(w_dff_B_wQV5JdOo7_2),.clk(gclk));
	jdff dff_B_WKJbX2TY6_2(.din(w_dff_B_wQV5JdOo7_2),.dout(w_dff_B_WKJbX2TY6_2),.clk(gclk));
	jdff dff_B_YJqjLwA85_2(.din(w_dff_B_WKJbX2TY6_2),.dout(w_dff_B_YJqjLwA85_2),.clk(gclk));
	jdff dff_B_UJMbps260_2(.din(w_dff_B_YJqjLwA85_2),.dout(w_dff_B_UJMbps260_2),.clk(gclk));
	jdff dff_B_H8qyBEwP5_2(.din(w_dff_B_UJMbps260_2),.dout(w_dff_B_H8qyBEwP5_2),.clk(gclk));
	jdff dff_B_eQgywDC07_2(.din(w_dff_B_H8qyBEwP5_2),.dout(w_dff_B_eQgywDC07_2),.clk(gclk));
	jdff dff_B_zDz5HAab4_2(.din(w_dff_B_eQgywDC07_2),.dout(w_dff_B_zDz5HAab4_2),.clk(gclk));
	jdff dff_A_U5A0OWvQ2_0(.dout(w_n1403_0[0]),.din(w_dff_A_U5A0OWvQ2_0),.clk(gclk));
	jdff dff_B_8OKTv9XE9_2(.din(n1403),.dout(w_dff_B_8OKTv9XE9_2),.clk(gclk));
	jdff dff_B_GD9uVb5h8_2(.din(w_dff_B_8OKTv9XE9_2),.dout(w_dff_B_GD9uVb5h8_2),.clk(gclk));
	jdff dff_B_U2Q129iN0_2(.din(w_dff_B_GD9uVb5h8_2),.dout(w_dff_B_U2Q129iN0_2),.clk(gclk));
	jdff dff_B_NgjrwS3f3_2(.din(w_dff_B_U2Q129iN0_2),.dout(w_dff_B_NgjrwS3f3_2),.clk(gclk));
	jdff dff_B_EM70p3Km8_2(.din(w_dff_B_NgjrwS3f3_2),.dout(w_dff_B_EM70p3Km8_2),.clk(gclk));
	jdff dff_B_xayyrLPC6_2(.din(w_dff_B_EM70p3Km8_2),.dout(w_dff_B_xayyrLPC6_2),.clk(gclk));
	jdff dff_B_0gN2yr7p2_2(.din(w_dff_B_xayyrLPC6_2),.dout(w_dff_B_0gN2yr7p2_2),.clk(gclk));
	jdff dff_B_Eo2L0ZQs7_2(.din(w_dff_B_0gN2yr7p2_2),.dout(w_dff_B_Eo2L0ZQs7_2),.clk(gclk));
	jdff dff_B_ps9EMUV09_2(.din(w_dff_B_Eo2L0ZQs7_2),.dout(w_dff_B_ps9EMUV09_2),.clk(gclk));
	jdff dff_B_w6PwYQ2n3_2(.din(w_dff_B_ps9EMUV09_2),.dout(w_dff_B_w6PwYQ2n3_2),.clk(gclk));
	jdff dff_B_SITQzVFv6_2(.din(w_dff_B_w6PwYQ2n3_2),.dout(w_dff_B_SITQzVFv6_2),.clk(gclk));
	jdff dff_B_0l4IU0o40_2(.din(w_dff_B_SITQzVFv6_2),.dout(w_dff_B_0l4IU0o40_2),.clk(gclk));
	jdff dff_B_mKUwH91I0_1(.din(n1429),.dout(w_dff_B_mKUwH91I0_1),.clk(gclk));
	jdff dff_B_kdpLK6Ir2_1(.din(w_dff_B_mKUwH91I0_1),.dout(w_dff_B_kdpLK6Ir2_1),.clk(gclk));
	jdff dff_B_pKPkoAf66_1(.din(w_dff_B_kdpLK6Ir2_1),.dout(w_dff_B_pKPkoAf66_1),.clk(gclk));
	jdff dff_B_7X10Oy2z1_1(.din(w_dff_B_pKPkoAf66_1),.dout(w_dff_B_7X10Oy2z1_1),.clk(gclk));
	jdff dff_B_YHswpmBN6_1(.din(w_dff_B_7X10Oy2z1_1),.dout(w_dff_B_YHswpmBN6_1),.clk(gclk));
	jdff dff_B_hTLr99948_1(.din(w_dff_B_YHswpmBN6_1),.dout(w_dff_B_hTLr99948_1),.clk(gclk));
	jdff dff_B_kh0mG0oH5_1(.din(w_dff_B_hTLr99948_1),.dout(w_dff_B_kh0mG0oH5_1),.clk(gclk));
	jdff dff_B_UXERPa0q1_1(.din(w_dff_B_kh0mG0oH5_1),.dout(w_dff_B_UXERPa0q1_1),.clk(gclk));
	jdff dff_B_wiYCOpmh7_1(.din(w_dff_B_UXERPa0q1_1),.dout(w_dff_B_wiYCOpmh7_1),.clk(gclk));
	jdff dff_B_YnIuCaKP6_1(.din(w_dff_B_wiYCOpmh7_1),.dout(w_dff_B_YnIuCaKP6_1),.clk(gclk));
	jdff dff_B_NWEmCtOZ2_1(.din(w_dff_B_YnIuCaKP6_1),.dout(w_dff_B_NWEmCtOZ2_1),.clk(gclk));
	jdff dff_B_wCjmDPvJ6_1(.din(w_dff_B_NWEmCtOZ2_1),.dout(w_dff_B_wCjmDPvJ6_1),.clk(gclk));
	jdff dff_A_D6vLbTgQ8_0(.dout(w_n1421_0[0]),.din(w_dff_A_D6vLbTgQ8_0),.clk(gclk));
	jdff dff_B_53fwDjvP2_2(.din(n1421),.dout(w_dff_B_53fwDjvP2_2),.clk(gclk));
	jdff dff_B_QOYar6qD9_2(.din(w_dff_B_53fwDjvP2_2),.dout(w_dff_B_QOYar6qD9_2),.clk(gclk));
	jdff dff_B_vleLRqDg6_2(.din(w_dff_B_QOYar6qD9_2),.dout(w_dff_B_vleLRqDg6_2),.clk(gclk));
	jdff dff_B_3bb3j1dn9_2(.din(w_dff_B_vleLRqDg6_2),.dout(w_dff_B_3bb3j1dn9_2),.clk(gclk));
	jdff dff_B_IPMENRrq7_2(.din(w_dff_B_3bb3j1dn9_2),.dout(w_dff_B_IPMENRrq7_2),.clk(gclk));
	jdff dff_B_o3Jo6RyQ2_2(.din(w_dff_B_IPMENRrq7_2),.dout(w_dff_B_o3Jo6RyQ2_2),.clk(gclk));
	jdff dff_B_jhaJRz5v8_2(.din(w_dff_B_o3Jo6RyQ2_2),.dout(w_dff_B_jhaJRz5v8_2),.clk(gclk));
	jdff dff_B_LDnfabSV4_2(.din(w_dff_B_jhaJRz5v8_2),.dout(w_dff_B_LDnfabSV4_2),.clk(gclk));
	jdff dff_B_LU6tQWlE5_2(.din(w_dff_B_LDnfabSV4_2),.dout(w_dff_B_LU6tQWlE5_2),.clk(gclk));
	jdff dff_B_koyHqIvp9_2(.din(w_dff_B_LU6tQWlE5_2),.dout(w_dff_B_koyHqIvp9_2),.clk(gclk));
	jdff dff_B_uYehnKMl7_2(.din(w_dff_B_koyHqIvp9_2),.dout(w_dff_B_uYehnKMl7_2),.clk(gclk));
	jdff dff_B_XagOhMGU8_2(.din(w_dff_B_uYehnKMl7_2),.dout(w_dff_B_XagOhMGU8_2),.clk(gclk));
	jdff dff_B_WRvEsVRJ4_2(.din(w_dff_B_XagOhMGU8_2),.dout(w_dff_B_WRvEsVRJ4_2),.clk(gclk));
	jdff dff_B_0DdkLjYW4_2(.din(w_dff_B_WRvEsVRJ4_2),.dout(w_dff_B_0DdkLjYW4_2),.clk(gclk));
	jdff dff_B_KFLkPMMh7_2(.din(w_dff_B_0DdkLjYW4_2),.dout(w_dff_B_KFLkPMMh7_2),.clk(gclk));
	jdff dff_B_NaOW4y5v8_2(.din(w_dff_B_KFLkPMMh7_2),.dout(w_dff_B_NaOW4y5v8_2),.clk(gclk));
	jdff dff_B_6nDF9O8S7_2(.din(w_dff_B_NaOW4y5v8_2),.dout(w_dff_B_6nDF9O8S7_2),.clk(gclk));
	jdff dff_B_x5PVJcHZ1_1(.din(n1432),.dout(w_dff_B_x5PVJcHZ1_1),.clk(gclk));
	jdff dff_B_EhEJoKax5_1(.din(w_dff_B_x5PVJcHZ1_1),.dout(w_dff_B_EhEJoKax5_1),.clk(gclk));
	jdff dff_B_gh8Zhfvx7_1(.din(w_dff_B_EhEJoKax5_1),.dout(w_dff_B_gh8Zhfvx7_1),.clk(gclk));
	jdff dff_B_cZNQdkW77_1(.din(w_dff_B_gh8Zhfvx7_1),.dout(w_dff_B_cZNQdkW77_1),.clk(gclk));
	jdff dff_B_I7eyIFiw4_1(.din(w_dff_B_cZNQdkW77_1),.dout(w_dff_B_I7eyIFiw4_1),.clk(gclk));
	jdff dff_B_zZiQPSHB6_1(.din(w_dff_B_I7eyIFiw4_1),.dout(w_dff_B_zZiQPSHB6_1),.clk(gclk));
	jdff dff_B_MkJ4RXvv1_1(.din(w_dff_B_zZiQPSHB6_1),.dout(w_dff_B_MkJ4RXvv1_1),.clk(gclk));
	jdff dff_B_N3I8Jjz22_1(.din(w_dff_B_MkJ4RXvv1_1),.dout(w_dff_B_N3I8Jjz22_1),.clk(gclk));
	jdff dff_B_f0Uny1RB5_1(.din(w_dff_B_N3I8Jjz22_1),.dout(w_dff_B_f0Uny1RB5_1),.clk(gclk));
	jdff dff_B_asBaZ9r35_1(.din(w_dff_B_f0Uny1RB5_1),.dout(w_dff_B_asBaZ9r35_1),.clk(gclk));
	jdff dff_B_BeNWbI3f0_1(.din(w_dff_B_asBaZ9r35_1),.dout(w_dff_B_BeNWbI3f0_1),.clk(gclk));
	jdff dff_B_latO3i3i6_1(.din(w_dff_B_BeNWbI3f0_1),.dout(w_dff_B_latO3i3i6_1),.clk(gclk));
	jdff dff_B_nxH7yyo68_1(.din(w_dff_B_latO3i3i6_1),.dout(w_dff_B_nxH7yyo68_1),.clk(gclk));
	jdff dff_B_KQXKqvIk2_0(.din(n1423),.dout(w_dff_B_KQXKqvIk2_0),.clk(gclk));
	jdff dff_B_IZwVng5o1_0(.din(w_dff_B_KQXKqvIk2_0),.dout(w_dff_B_IZwVng5o1_0),.clk(gclk));
	jdff dff_B_vzpbRXCp6_0(.din(w_dff_B_IZwVng5o1_0),.dout(w_dff_B_vzpbRXCp6_0),.clk(gclk));
	jdff dff_B_2Bc6UJop7_0(.din(w_dff_B_vzpbRXCp6_0),.dout(w_dff_B_2Bc6UJop7_0),.clk(gclk));
	jdff dff_B_sqMfXfB26_0(.din(w_dff_B_2Bc6UJop7_0),.dout(w_dff_B_sqMfXfB26_0),.clk(gclk));
	jdff dff_B_okDF1nOz8_0(.din(w_dff_B_sqMfXfB26_0),.dout(w_dff_B_okDF1nOz8_0),.clk(gclk));
	jdff dff_B_3Hwed9uF8_0(.din(w_dff_B_okDF1nOz8_0),.dout(w_dff_B_3Hwed9uF8_0),.clk(gclk));
	jdff dff_B_gce3rBAo9_0(.din(w_dff_B_3Hwed9uF8_0),.dout(w_dff_B_gce3rBAo9_0),.clk(gclk));
	jdff dff_B_PrrVwQBD1_0(.din(w_dff_B_gce3rBAo9_0),.dout(w_dff_B_PrrVwQBD1_0),.clk(gclk));
	jdff dff_B_mhxu8Eq72_0(.din(w_dff_B_PrrVwQBD1_0),.dout(w_dff_B_mhxu8Eq72_0),.clk(gclk));
	jdff dff_B_2ErCsl821_0(.din(w_dff_B_mhxu8Eq72_0),.dout(w_dff_B_2ErCsl821_0),.clk(gclk));
	jdff dff_B_09oTuabG4_0(.din(w_dff_B_2ErCsl821_0),.dout(w_dff_B_09oTuabG4_0),.clk(gclk));
	jdff dff_B_HjQBwVVw1_0(.din(w_dff_B_09oTuabG4_0),.dout(w_dff_B_HjQBwVVw1_0),.clk(gclk));
	jdff dff_B_KHPRBnxK0_0(.din(w_dff_B_HjQBwVVw1_0),.dout(w_dff_B_KHPRBnxK0_0),.clk(gclk));
	jdff dff_A_0Tg0GVpc8_0(.dout(w_n1422_0[0]),.din(w_dff_A_0Tg0GVpc8_0),.clk(gclk));
	jdff dff_B_NpolJDHj7_2(.din(n1422),.dout(w_dff_B_NpolJDHj7_2),.clk(gclk));
	jdff dff_B_aTtyaxgO4_2(.din(w_dff_B_NpolJDHj7_2),.dout(w_dff_B_aTtyaxgO4_2),.clk(gclk));
	jdff dff_B_cvk4diKq2_2(.din(w_dff_B_aTtyaxgO4_2),.dout(w_dff_B_cvk4diKq2_2),.clk(gclk));
	jdff dff_B_XN4lpS7F4_2(.din(w_dff_B_cvk4diKq2_2),.dout(w_dff_B_XN4lpS7F4_2),.clk(gclk));
	jdff dff_B_VzR6Q3Nw9_2(.din(w_dff_B_XN4lpS7F4_2),.dout(w_dff_B_VzR6Q3Nw9_2),.clk(gclk));
	jdff dff_B_WaMjxWFi9_2(.din(w_dff_B_VzR6Q3Nw9_2),.dout(w_dff_B_WaMjxWFi9_2),.clk(gclk));
	jdff dff_B_wzO7q3NX5_2(.din(w_dff_B_WaMjxWFi9_2),.dout(w_dff_B_wzO7q3NX5_2),.clk(gclk));
	jdff dff_B_EljRkBnR8_2(.din(w_dff_B_wzO7q3NX5_2),.dout(w_dff_B_EljRkBnR8_2),.clk(gclk));
	jdff dff_B_FjHYRCtP3_2(.din(w_dff_B_EljRkBnR8_2),.dout(w_dff_B_FjHYRCtP3_2),.clk(gclk));
	jdff dff_B_Wyodgqcx1_2(.din(w_dff_B_FjHYRCtP3_2),.dout(w_dff_B_Wyodgqcx1_2),.clk(gclk));
	jdff dff_B_5WyXIVz35_2(.din(w_dff_B_Wyodgqcx1_2),.dout(w_dff_B_5WyXIVz35_2),.clk(gclk));
	jdff dff_B_CvXfG5r89_2(.din(w_dff_B_5WyXIVz35_2),.dout(w_dff_B_CvXfG5r89_2),.clk(gclk));
	jdff dff_B_mbFam3nO9_2(.din(w_dff_B_CvXfG5r89_2),.dout(w_dff_B_mbFam3nO9_2),.clk(gclk));
	jdff dff_B_XHdLJZGC4_2(.din(w_dff_B_mbFam3nO9_2),.dout(w_dff_B_XHdLJZGC4_2),.clk(gclk));
	jdff dff_B_UQDYOXCH3_2(.din(w_dff_B_XHdLJZGC4_2),.dout(w_dff_B_UQDYOXCH3_2),.clk(gclk));
	jdff dff_B_Hq71TNA62_2(.din(w_dff_B_UQDYOXCH3_2),.dout(w_dff_B_Hq71TNA62_2),.clk(gclk));
	jdff dff_B_mr5mYk7H5_0(.din(n1441),.dout(w_dff_B_mr5mYk7H5_0),.clk(gclk));
	jdff dff_B_QD0a7OGU7_0(.din(n1440),.dout(w_dff_B_QD0a7OGU7_0),.clk(gclk));
	jdff dff_B_P52bzwOL2_0(.din(w_dff_B_QD0a7OGU7_0),.dout(w_dff_B_P52bzwOL2_0),.clk(gclk));
	jdff dff_B_6E67m9nk2_0(.din(w_dff_B_P52bzwOL2_0),.dout(w_dff_B_6E67m9nk2_0),.clk(gclk));
	jdff dff_B_o6C0FC1J8_0(.din(w_dff_B_6E67m9nk2_0),.dout(w_dff_B_o6C0FC1J8_0),.clk(gclk));
	jdff dff_B_gmsbbxjL8_0(.din(w_dff_B_o6C0FC1J8_0),.dout(w_dff_B_gmsbbxjL8_0),.clk(gclk));
	jdff dff_B_pP0s51ua1_0(.din(w_dff_B_gmsbbxjL8_0),.dout(w_dff_B_pP0s51ua1_0),.clk(gclk));
	jdff dff_B_173T7hMJ2_0(.din(n1212),.dout(w_dff_B_173T7hMJ2_0),.clk(gclk));
	jdff dff_B_Q74RQj760_0(.din(n1209),.dout(w_dff_B_Q74RQj760_0),.clk(gclk));
	jdff dff_B_HWQXCFiG4_1(.din(n1206),.dout(w_dff_B_HWQXCFiG4_1),.clk(gclk));
	jdff dff_B_NHTV8UlK1_1(.din(n1204),.dout(w_dff_B_NHTV8UlK1_1),.clk(gclk));
	jdff dff_B_fWbOweMG4_0(.din(n1197),.dout(w_dff_B_fWbOweMG4_0),.clk(gclk));
	jdff dff_B_fjEFjj683_1(.din(n1190),.dout(w_dff_B_fjEFjj683_1),.clk(gclk));
	jdff dff_B_EhhukHxl3_1(.din(w_dff_B_fjEFjj683_1),.dout(w_dff_B_EhhukHxl3_1),.clk(gclk));
	jdff dff_B_uzyJlzBQ0_1(.din(n1188),.dout(w_dff_B_uzyJlzBQ0_1),.clk(gclk));
	jdff dff_B_9IECpHVC3_1(.din(n1175),.dout(w_dff_B_9IECpHVC3_1),.clk(gclk));
	jdff dff_B_Wv8yPjb91_1(.din(w_dff_B_9IECpHVC3_1),.dout(w_dff_B_Wv8yPjb91_1),.clk(gclk));
	jdff dff_B_pSO67Ttc4_1(.din(w_dff_B_Wv8yPjb91_1),.dout(w_dff_B_pSO67Ttc4_1),.clk(gclk));
	jdff dff_B_Y3DHXPlw4_1(.din(w_dff_B_pSO67Ttc4_1),.dout(w_dff_B_Y3DHXPlw4_1),.clk(gclk));
	jdff dff_B_DJ4w6L5y8_1(.din(n1176),.dout(w_dff_B_DJ4w6L5y8_1),.clk(gclk));
	jdff dff_B_OGURsFGT2_1(.din(w_dff_B_DJ4w6L5y8_1),.dout(w_dff_B_OGURsFGT2_1),.clk(gclk));
	jdff dff_B_W377iLEv9_1(.din(w_dff_B_OGURsFGT2_1),.dout(w_dff_B_W377iLEv9_1),.clk(gclk));
	jdff dff_B_SyQToNJc4_1(.din(w_dff_B_W377iLEv9_1),.dout(w_dff_B_SyQToNJc4_1),.clk(gclk));
	jdff dff_B_BdmlA7k07_1(.din(n1181),.dout(w_dff_B_BdmlA7k07_1),.clk(gclk));
	jdff dff_B_9gASExGS4_0(.din(n1174),.dout(w_dff_B_9gASExGS4_0),.clk(gclk));
	jdff dff_B_tDGVdp7M2_0(.din(w_dff_B_9gASExGS4_0),.dout(w_dff_B_tDGVdp7M2_0),.clk(gclk));
	jdff dff_B_sVv5WnBc8_1(.din(n1153),.dout(w_dff_B_sVv5WnBc8_1),.clk(gclk));
	jdff dff_B_rqPeaL4Q4_1(.din(w_dff_B_sVv5WnBc8_1),.dout(w_dff_B_rqPeaL4Q4_1),.clk(gclk));
	jdff dff_B_UYU4h3RQ3_1(.din(w_dff_B_rqPeaL4Q4_1),.dout(w_dff_B_UYU4h3RQ3_1),.clk(gclk));
	jdff dff_B_oe85dSHx4_1(.din(w_dff_B_UYU4h3RQ3_1),.dout(w_dff_B_oe85dSHx4_1),.clk(gclk));
	jdff dff_B_Z1bZWMPx7_1(.din(w_dff_B_oe85dSHx4_1),.dout(w_dff_B_Z1bZWMPx7_1),.clk(gclk));
	jdff dff_B_TvFokxhq6_1(.din(n1155),.dout(w_dff_B_TvFokxhq6_1),.clk(gclk));
	jdff dff_B_xHL8bKfi8_1(.din(w_dff_B_TvFokxhq6_1),.dout(w_dff_B_xHL8bKfi8_1),.clk(gclk));
	jdff dff_B_ORUhP1w48_1(.din(w_dff_B_xHL8bKfi8_1),.dout(w_dff_B_ORUhP1w48_1),.clk(gclk));
	jdff dff_B_boMQhpJ27_0(.din(n1169),.dout(w_dff_B_boMQhpJ27_0),.clk(gclk));
	jdff dff_B_Mq6MvMiN9_0(.din(w_dff_B_boMQhpJ27_0),.dout(w_dff_B_Mq6MvMiN9_0),.clk(gclk));
	jdff dff_B_opeCNCVQ1_0(.din(w_dff_B_Mq6MvMiN9_0),.dout(w_dff_B_opeCNCVQ1_0),.clk(gclk));
	jdff dff_B_bpWNMMEc7_0(.din(w_dff_B_opeCNCVQ1_0),.dout(w_dff_B_bpWNMMEc7_0),.clk(gclk));
	jdff dff_B_cRJVO95d6_0(.din(n1355),.dout(w_dff_B_cRJVO95d6_0),.clk(gclk));
	jdff dff_B_B2EznjiX3_0(.din(w_dff_B_cRJVO95d6_0),.dout(w_dff_B_B2EznjiX3_0),.clk(gclk));
	jdff dff_B_gjvsLsyS4_0(.din(w_dff_B_B2EznjiX3_0),.dout(w_dff_B_gjvsLsyS4_0),.clk(gclk));
	jdff dff_B_WHtaxa8G1_1(.din(n1337),.dout(w_dff_B_WHtaxa8G1_1),.clk(gclk));
	jdff dff_B_nlwoff1o3_1(.din(w_dff_B_WHtaxa8G1_1),.dout(w_dff_B_nlwoff1o3_1),.clk(gclk));
	jdff dff_B_0ZQfZymY9_1(.din(w_dff_B_nlwoff1o3_1),.dout(w_dff_B_0ZQfZymY9_1),.clk(gclk));
	jdff dff_B_BRbGO4Yg4_1(.din(n1338),.dout(w_dff_B_BRbGO4Yg4_1),.clk(gclk));
	jdff dff_B_cIktG6lr3_1(.din(w_dff_B_BRbGO4Yg4_1),.dout(w_dff_B_cIktG6lr3_1),.clk(gclk));
	jdff dff_B_LfJWX3D13_1(.din(w_dff_B_cIktG6lr3_1),.dout(w_dff_B_LfJWX3D13_1),.clk(gclk));
	jdff dff_B_MCaZvy6c3_0(.din(n1352),.dout(w_dff_B_MCaZvy6c3_0),.clk(gclk));
	jdff dff_B_2hXY8mZJ4_0(.din(w_dff_B_MCaZvy6c3_0),.dout(w_dff_B_2hXY8mZJ4_0),.clk(gclk));
	jdff dff_B_uQvFpwT72_0(.din(w_dff_B_2hXY8mZJ4_0),.dout(w_dff_B_uQvFpwT72_0),.clk(gclk));
	jdff dff_B_ZhNlUfdm8_0(.din(G174),.dout(w_dff_B_ZhNlUfdm8_0),.clk(gclk));
	jdff dff_B_OEvkFNga5_0(.din(G173),.dout(w_dff_B_OEvkFNga5_0),.clk(gclk));
	jdff dff_B_bRo8Z4hO6_0(.din(G176),.dout(w_dff_B_bRo8Z4hO6_0),.clk(gclk));
	jdff dff_B_kwT9n1fz3_0(.din(G175),.dout(w_dff_B_kwT9n1fz3_0),.clk(gclk));
	jdff dff_B_jMZecd1B1_0(.din(n753),.dout(w_dff_B_jMZecd1B1_0),.clk(gclk));
	jdff dff_B_xFKgSs601_0(.din(G177),.dout(w_dff_B_xFKgSs601_0),.clk(gclk));
	jdff dff_B_mds2AIK08_0(.din(n743),.dout(w_dff_B_mds2AIK08_0),.clk(gclk));
	jdff dff_B_2pGwruPz1_0(.din(n729),.dout(w_dff_B_2pGwruPz1_0),.clk(gclk));
	jdff dff_A_FCPrPmIm8_0(.dout(w_n737_0[0]),.din(w_dff_A_FCPrPmIm8_0),.clk(gclk));
	jdff dff_B_uYOex2N95_0(.din(n736),.dout(w_dff_B_uYOex2N95_0),.clk(gclk));
	jdff dff_B_1NXFRMjk4_1(.din(n1311),.dout(w_dff_B_1NXFRMjk4_1),.clk(gclk));
	jdff dff_B_rreQ0XYf0_1(.din(w_dff_B_1NXFRMjk4_1),.dout(w_dff_B_rreQ0XYf0_1),.clk(gclk));
	jdff dff_B_gICgOpXL2_1(.din(n1326),.dout(w_dff_B_gICgOpXL2_1),.clk(gclk));
	jdff dff_B_yLk5tBE51_1(.din(w_dff_B_gICgOpXL2_1),.dout(w_dff_B_yLk5tBE51_1),.clk(gclk));
	jdff dff_B_p3lLlLER1_1(.din(n1327),.dout(w_dff_B_p3lLlLER1_1),.clk(gclk));
	jdff dff_B_Ua5UgG9c8_0(.din(n1324),.dout(w_dff_B_Ua5UgG9c8_0),.clk(gclk));
	jdff dff_B_N64ZuN0W7_0(.din(n1323),.dout(w_dff_B_N64ZuN0W7_0),.clk(gclk));
	jdff dff_B_rtQVUCQU1_0(.din(n907),.dout(w_dff_B_rtQVUCQU1_0),.clk(gclk));
	jdff dff_B_fPYqTgMv3_0(.din(w_dff_B_rtQVUCQU1_0),.dout(w_dff_B_fPYqTgMv3_0),.clk(gclk));
	jdff dff_B_83WXd5ql7_0(.din(n944),.dout(w_dff_B_83WXd5ql7_0),.clk(gclk));
	jdff dff_B_ppmXzpJe8_0(.din(w_dff_B_83WXd5ql7_0),.dout(w_dff_B_ppmXzpJe8_0),.clk(gclk));
	jdff dff_B_1MoapjDq3_0(.din(n926),.dout(w_dff_B_1MoapjDq3_0),.clk(gclk));
	jdff dff_B_PhDfeFx85_0(.din(w_dff_B_1MoapjDq3_0),.dout(w_dff_B_PhDfeFx85_0),.clk(gclk));
	jdff dff_B_rf7vgArF7_0(.din(n915),.dout(w_dff_B_rf7vgArF7_0),.clk(gclk));
	jdff dff_B_rVvKV7Bp3_0(.din(w_dff_B_rf7vgArF7_0),.dout(w_dff_B_rVvKV7Bp3_0),.clk(gclk));
	jdff dff_B_n43mFXus8_1(.din(n1313),.dout(w_dff_B_n43mFXus8_1),.clk(gclk));
	jdff dff_B_lQ8Q3Dii3_1(.din(w_dff_B_n43mFXus8_1),.dout(w_dff_B_lQ8Q3Dii3_1),.clk(gclk));
	jdff dff_B_v0ffNHLM7_1(.din(w_dff_B_lQ8Q3Dii3_1),.dout(w_dff_B_v0ffNHLM7_1),.clk(gclk));
	jdff dff_B_CN1hRy5D4_0(.din(n898),.dout(w_dff_B_CN1hRy5D4_0),.clk(gclk));
	jdff dff_B_7XSr0N1X0_0(.din(w_dff_B_CN1hRy5D4_0),.dout(w_dff_B_7XSr0N1X0_0),.clk(gclk));
	jdff dff_A_xTpTo3FQ6_1(.dout(w_n891_0[1]),.din(w_dff_A_xTpTo3FQ6_1),.clk(gclk));
	jdff dff_B_8XEg0JBA1_0(.din(n890),.dout(w_dff_B_8XEg0JBA1_0),.clk(gclk));
	jdff dff_B_0p1asTaz8_0(.din(n877),.dout(w_dff_B_0p1asTaz8_0),.clk(gclk));
	jdff dff_B_GHMBKMEz3_0(.din(w_dff_B_0p1asTaz8_0),.dout(w_dff_B_GHMBKMEz3_0),.clk(gclk));
	jdff dff_B_3u7H70DV1_0(.din(n1312),.dout(w_dff_B_3u7H70DV1_0),.clk(gclk));
	jdff dff_B_ACQkRp2d8_0(.din(G44),.dout(w_dff_B_ACQkRp2d8_0),.clk(gclk));
	jdff dff_B_ZkCoSXX81_0(.din(n1308),.dout(w_dff_B_ZkCoSXX81_0),.clk(gclk));
	jdff dff_B_lXAUZjrw9_0(.din(w_dff_B_ZkCoSXX81_0),.dout(w_dff_B_lXAUZjrw9_0),.clk(gclk));
	jdff dff_B_FVEpOpmI2_0(.din(n842),.dout(w_dff_B_FVEpOpmI2_0),.clk(gclk));
	jdff dff_B_Cq4SEy4M3_0(.din(n811),.dout(w_dff_B_Cq4SEy4M3_0),.clk(gclk));
	jdff dff_B_VWQRY0eh8_0(.din(n826),.dout(w_dff_B_VWQRY0eh8_0),.clk(gclk));
	jdff dff_B_pEGy5yFX6_0(.din(n818),.dout(w_dff_B_pEGy5yFX6_0),.clk(gclk));
	jdff dff_B_QcCZd2tT0_0(.din(n1302),.dout(w_dff_B_QcCZd2tT0_0),.clk(gclk));
	jdff dff_B_lMdIjjqA3_0(.din(G115),.dout(w_dff_B_lMdIjjqA3_0),.clk(gclk));
	jdff dff_A_jov50joB5_1(.dout(w_n1301_0[1]),.din(w_dff_A_jov50joB5_1),.clk(gclk));
	jdff dff_B_y2mL8afH4_0(.din(n803),.dout(w_dff_B_y2mL8afH4_0),.clk(gclk));
	jdff dff_B_yCOS2wms3_0(.din(n796),.dout(w_dff_B_yCOS2wms3_0),.clk(gclk));
	jdff dff_B_BdF6J7Nd9_0(.din(n789),.dout(w_dff_B_BdF6J7Nd9_0),.clk(gclk));
	jdff dff_B_UYt0YtB46_0(.din(n783),.dout(w_dff_B_UYt0YtB46_0),.clk(gclk));
	jdff dff_A_VL9wH6h17_0(.dout(w_n851_0[0]),.din(w_dff_A_VL9wH6h17_0),.clk(gclk));
	jdff dff_A_XC64y0ZQ7_0(.dout(w_dff_A_VL9wH6h17_0),.din(w_dff_A_XC64y0ZQ7_0),.clk(gclk));
	jdff dff_B_h00Pwn007_0(.din(n850),.dout(w_dff_B_h00Pwn007_0),.clk(gclk));
	jdff dff_B_fIb3v3qv5_1(.din(n1288),.dout(w_dff_B_fIb3v3qv5_1),.clk(gclk));
	jdff dff_B_xEb6tKc84_0(.din(n1295),.dout(w_dff_B_xEb6tKc84_0),.clk(gclk));
	jdff dff_B_P2YIAgvt6_0(.din(w_dff_B_xEb6tKc84_0),.dout(w_dff_B_P2YIAgvt6_0),.clk(gclk));
	jdff dff_B_4Ng3MVty1_0(.din(n1294),.dout(w_dff_B_4Ng3MVty1_0),.clk(gclk));
	jdff dff_B_mxs537I87_0(.din(w_dff_B_4Ng3MVty1_0),.dout(w_dff_B_mxs537I87_0),.clk(gclk));
	jdff dff_A_2DeFixeh3_2(.dout(w_G18_22[2]),.din(w_dff_A_2DeFixeh3_2),.clk(gclk));
	jdff dff_A_p6fYGlLf3_2(.dout(w_dff_A_2DeFixeh3_2),.din(w_dff_A_p6fYGlLf3_2),.clk(gclk));
	jdff dff_A_n6hM84nC4_0(.dout(w_n1095_0[0]),.din(w_dff_A_n6hM84nC4_0),.clk(gclk));
	jdff dff_A_VqC2Fu7o5_0(.dout(w_dff_A_n6hM84nC4_0),.din(w_dff_A_VqC2Fu7o5_0),.clk(gclk));
	jdff dff_B_7fLkiLQM3_0(.din(G168),.dout(w_dff_B_7fLkiLQM3_0),.clk(gclk));
	jdff dff_A_c2BPqbnV3_0(.dout(w_n1076_0[0]),.din(w_dff_A_c2BPqbnV3_0),.clk(gclk));
	jdff dff_A_v1DXBwy66_0(.dout(w_dff_A_c2BPqbnV3_0),.din(w_dff_A_v1DXBwy66_0),.clk(gclk));
	jdff dff_B_t28gJu808_0(.din(G169),.dout(w_dff_B_t28gJu808_0),.clk(gclk));
	jdff dff_A_tvyGr8hS2_0(.dout(w_n565_4[0]),.din(w_dff_A_tvyGr8hS2_0),.clk(gclk));
	jdff dff_A_mwjuaXS58_1(.dout(w_n565_4[1]),.din(w_dff_A_mwjuaXS58_1),.clk(gclk));
	jdff dff_B_cmy3iLci6_1(.din(n1280),.dout(w_dff_B_cmy3iLci6_1),.clk(gclk));
	jdff dff_B_b19WWDy46_0(.din(G166),.dout(w_dff_B_b19WWDy46_0),.clk(gclk));
	jdff dff_A_RBRzs81B1_0(.dout(w_n1061_0[0]),.din(w_dff_A_RBRzs81B1_0),.clk(gclk));
	jdff dff_B_FnEjt97S5_0(.din(G167),.dout(w_dff_B_FnEjt97S5_0),.clk(gclk));
	jdff dff_A_L9yEVs9h8_0(.dout(w_G414_0),.din(w_dff_A_L9yEVs9h8_0),.clk(gclk));
	jdff dff_A_GksR6ZpJ8_0(.dout(w_dff_A_L9yEVs9h8_0),.din(w_dff_A_GksR6ZpJ8_0),.clk(gclk));
	jdff dff_A_CfZ6Oqln4_0(.dout(w_dff_A_GksR6ZpJ8_0),.din(w_dff_A_CfZ6Oqln4_0),.clk(gclk));
	jdff dff_B_64dqJnW15_1(.din(n1227),.dout(w_dff_B_64dqJnW15_1),.clk(gclk));
	jdff dff_B_W3BPbTjj3_1(.din(w_dff_B_64dqJnW15_1),.dout(w_dff_B_W3BPbTjj3_1),.clk(gclk));
	jdff dff_B_OP2RUF7k2_0(.din(n1273),.dout(w_dff_B_OP2RUF7k2_0),.clk(gclk));
	jdff dff_B_Lcgy86XL0_0(.din(n740),.dout(w_dff_B_Lcgy86XL0_0),.clk(gclk));
	jdff dff_B_U1958RBQ3_0(.din(n733),.dout(w_dff_B_U1958RBQ3_0),.clk(gclk));
	jdff dff_B_hfEIVdUV0_1(.din(n1270),.dout(w_dff_B_hfEIVdUV0_1),.clk(gclk));
	jdff dff_B_ZvV1HQX72_0(.din(n757),.dout(w_dff_B_ZvV1HQX72_0),.clk(gclk));
	jdff dff_B_m2voZ3vE6_0(.din(n747),.dout(w_dff_B_m2voZ3vE6_0),.clk(gclk));
	jdff dff_A_xccNKG1p6_1(.dout(w_G2208_0[1]),.din(w_dff_A_xccNKG1p6_1),.clk(gclk));
	jdff dff_B_UY3GNvtW9_0(.din(n1018),.dout(w_dff_B_UY3GNvtW9_0),.clk(gclk));
	jdff dff_B_eCcZfGh83_0(.din(n1012),.dout(w_dff_B_eCcZfGh83_0),.clk(gclk));
	jdff dff_B_gbjOsGnH4_0(.din(n998),.dout(w_dff_B_gbjOsGnH4_0),.clk(gclk));
	jdff dff_B_l5t1Lzlf2_0(.din(n991),.dout(w_dff_B_l5t1Lzlf2_0),.clk(gclk));
	jdff dff_A_81yKPvvS6_0(.dout(w_n727_0[0]),.din(w_dff_A_81yKPvvS6_0),.clk(gclk));
	jdff dff_A_MOHz5gvg5_0(.dout(w_dff_A_81yKPvvS6_0),.din(w_dff_A_MOHz5gvg5_0),.clk(gclk));
	jdff dff_B_Ys5oJSE10_0(.din(n726),.dout(w_dff_B_Ys5oJSE10_0),.clk(gclk));
	jdff dff_B_NBUZtjFn9_1(.din(n1253),.dout(w_dff_B_NBUZtjFn9_1),.clk(gclk));
	jdff dff_B_Q9WaGEmw0_0(.din(n1260),.dout(w_dff_B_Q9WaGEmw0_0),.clk(gclk));
	jdff dff_B_9hGaIqOb4_0(.din(w_dff_B_Q9WaGEmw0_0),.dout(w_dff_B_9hGaIqOb4_0),.clk(gclk));
	jdff dff_B_R6DqXCQT1_0(.din(n1099),.dout(w_dff_B_R6DqXCQT1_0),.clk(gclk));
	jdff dff_A_1y77Buen6_0(.dout(w_G18_23[0]),.din(w_dff_A_1y77Buen6_0),.clk(gclk));
	jdff dff_B_FkoeeYcx3_0(.din(n1072),.dout(w_dff_B_FkoeeYcx3_0),.clk(gclk));
	jdff dff_A_Um3i6k0s2_0(.dout(w_n1066_0[0]),.din(w_dff_A_Um3i6k0s2_0),.clk(gclk));
	jdff dff_B_zwpHeb496_0(.din(n1065),.dout(w_dff_B_zwpHeb496_0),.clk(gclk));
	jdff dff_B_hCoIS9vy3_1(.din(n1251),.dout(w_dff_B_hCoIS9vy3_1),.clk(gclk));
	jdff dff_B_4F3mVGZg2_0(.din(n1085),.dout(w_dff_B_4F3mVGZg2_0),.clk(gclk));
	jdff dff_B_6eM1AfF22_0(.din(n1080),.dout(w_dff_B_6eM1AfF22_0),.clk(gclk));
	jdff dff_A_Aax5Nc2t1_1(.dout(w_G1459_0[1]),.din(w_dff_A_Aax5Nc2t1_1),.clk(gclk));
	jdff dff_B_AqWoWdRJ9_1(.din(n1237),.dout(w_dff_B_AqWoWdRJ9_1),.clk(gclk));
	jdff dff_B_1rCp1k1u8_1(.din(w_dff_B_AqWoWdRJ9_1),.dout(w_dff_B_1rCp1k1u8_1),.clk(gclk));
	jdff dff_B_UT9nz9814_1(.din(n1238),.dout(w_dff_B_UT9nz9814_1),.clk(gclk));
	jdff dff_B_fsMbef7P3_1(.din(w_dff_B_UT9nz9814_1),.dout(w_dff_B_fsMbef7P3_1),.clk(gclk));
	jdff dff_B_aLTbXciP5_1(.din(n1239),.dout(w_dff_B_aLTbXciP5_1),.clk(gclk));
	jdff dff_A_Rjv8E4uC9_1(.dout(w_n902_0[1]),.din(w_dff_A_Rjv8E4uC9_1),.clk(gclk));
	jdff dff_A_DWrTK79g5_2(.dout(w_n902_0[2]),.din(w_dff_A_DWrTK79g5_2),.clk(gclk));
	jdff dff_B_IUEL5QAU1_1(.din(n900),.dout(w_dff_B_IUEL5QAU1_1),.clk(gclk));
	jdff dff_B_hNhDWOew7_1(.din(n892),.dout(w_dff_B_hNhDWOew7_1),.clk(gclk));
	jdff dff_A_8QpsK7Yt1_1(.dout(w_n882_0[1]),.din(w_dff_A_8QpsK7Yt1_1),.clk(gclk));
	jdff dff_A_5CD2Eegm4_2(.dout(w_n882_0[2]),.din(w_dff_A_5CD2Eegm4_2),.clk(gclk));
	jdff dff_B_PUf4qp3b3_1(.din(n879),.dout(w_dff_B_PUf4qp3b3_1),.clk(gclk));
	jdff dff_A_1PkpiUyh1_1(.dout(w_n873_0[1]),.din(w_dff_A_1PkpiUyh1_1),.clk(gclk));
	jdff dff_A_QYNBPp378_2(.dout(w_n873_0[2]),.din(w_dff_A_QYNBPp378_2),.clk(gclk));
	jdff dff_B_JfloGEvr0_1(.din(n870),.dout(w_dff_B_JfloGEvr0_1),.clk(gclk));
	jdff dff_A_SJRSbQzT0_1(.dout(w_n920_0[1]),.din(w_dff_A_SJRSbQzT0_1),.clk(gclk));
	jdff dff_A_M23IpCZd7_2(.dout(w_n920_0[2]),.din(w_dff_A_M23IpCZd7_2),.clk(gclk));
	jdff dff_B_uXICOqHD1_1(.din(n917),.dout(w_dff_B_uXICOqHD1_1),.clk(gclk));
	jdff dff_A_Omj3E1au7_0(.dout(w_n948_0[0]),.din(w_dff_A_Omj3E1au7_0),.clk(gclk));
	jdff dff_A_OMALyz483_2(.dout(w_n948_0[2]),.din(w_dff_A_OMALyz483_2),.clk(gclk));
	jdff dff_B_tcaMqhgn1_1(.din(n946),.dout(w_dff_B_tcaMqhgn1_1),.clk(gclk));
	jdff dff_A_d6l7CZCQ0_1(.dout(w_n931_0[1]),.din(w_dff_A_d6l7CZCQ0_1),.clk(gclk));
	jdff dff_A_r5guVyE14_2(.dout(w_n931_0[2]),.din(w_dff_A_r5guVyE14_2),.clk(gclk));
	jdff dff_B_zE8vol1i0_1(.din(n928),.dout(w_dff_B_zE8vol1i0_1),.clk(gclk));
	jdff dff_A_IJjwYJTk3_0(.dout(w_n1236_0[0]),.din(w_dff_A_IJjwYJTk3_0),.clk(gclk));
	jdff dff_A_MeVxKv7k8_0(.dout(w_dff_A_IJjwYJTk3_0),.din(w_dff_A_MeVxKv7k8_0),.clk(gclk));
	jdff dff_A_ZmKoTLCU6_1(.dout(w_G3698_0[1]),.din(w_dff_A_ZmKoTLCU6_1),.clk(gclk));
	jdff dff_B_CzetVjBx0_3(.din(n912),.dout(w_dff_B_CzetVjBx0_3),.clk(gclk));
	jdff dff_B_Bh5QiV947_1(.din(n909),.dout(w_dff_B_Bh5QiV947_1),.clk(gclk));
	jdff dff_B_pos8EslO2_1(.din(n1215),.dout(w_dff_B_pos8EslO2_1),.clk(gclk));
	jdff dff_B_bgi1gc382_1(.din(w_dff_B_pos8EslO2_1),.dout(w_dff_B_bgi1gc382_1),.clk(gclk));
	jdff dff_B_DbGk8HA50_1(.din(w_dff_B_bgi1gc382_1),.dout(w_dff_B_DbGk8HA50_1),.clk(gclk));
	jdff dff_B_SJTdq7ix4_1(.din(n1217),.dout(w_dff_B_SJTdq7ix4_1),.clk(gclk));
	jdff dff_B_GSjpiOkW6_0(.din(n1224),.dout(w_dff_B_GSjpiOkW6_0),.clk(gclk));
	jdff dff_B_8LCFIIXv6_0(.din(w_dff_B_GSjpiOkW6_0),.dout(w_dff_B_8LCFIIXv6_0),.clk(gclk));
	jdff dff_A_8eJPHOff4_1(.dout(w_G4393_0[1]),.din(w_dff_A_8eJPHOff4_1),.clk(gclk));
	jdff dff_A_3iXJCCI03_1(.dout(w_n355_10[1]),.din(w_dff_A_3iXJCCI03_1),.clk(gclk));
	jdff dff_B_aDgzSQ3W6_1(.din(n805),.dout(w_dff_B_aDgzSQ3W6_1),.clk(gclk));
	jdff dff_B_sNtu3yve4_1(.din(n798),.dout(w_dff_B_sNtu3yve4_1),.clk(gclk));
	jdff dff_B_XUlCmyH13_1(.din(n791),.dout(w_dff_B_XUlCmyH13_1),.clk(gclk));
	jdff dff_B_B0owYQxb4_1(.din(n785),.dout(w_dff_B_B0owYQxb4_1),.clk(gclk));
	jdff dff_B_F9BIbIMB5_1(.din(n844),.dout(w_dff_B_F9BIbIMB5_1),.clk(gclk));
	jdff dff_B_WDAEk5L34_1(.din(n813),.dout(w_dff_B_WDAEk5L34_1),.clk(gclk));
	jdff dff_A_bQRHzGDs9_0(.dout(w_n855_0[0]),.din(w_dff_A_bQRHzGDs9_0),.clk(gclk));
	jdff dff_B_02keszY75_1(.din(n852),.dout(w_dff_B_02keszY75_1),.clk(gclk));
	jdff dff_B_DAJuA5HC0_1(.din(n828),.dout(w_dff_B_DAJuA5HC0_1),.clk(gclk));
	jdff dff_B_P2O9N3ze6_1(.din(n820),.dout(w_dff_B_P2O9N3ze6_1),.clk(gclk));
	jdff dff_B_WBgQZcFf6_3(.din(n720),.dout(w_dff_B_WBgQZcFf6_3),.clk(gclk));
	jdff dff_B_Bcaf6cA64_3(.din(w_dff_B_WBgQZcFf6_3),.dout(w_dff_B_Bcaf6cA64_3),.clk(gclk));
	jdff dff_B_3eVDKZ8r3_3(.din(w_dff_B_Bcaf6cA64_3),.dout(w_dff_B_3eVDKZ8r3_3),.clk(gclk));
	jdff dff_B_lqrthS1O3_3(.din(w_dff_B_3eVDKZ8r3_3),.dout(w_dff_B_lqrthS1O3_3),.clk(gclk));
	jdff dff_B_Jj3NHDP84_3(.din(w_dff_B_lqrthS1O3_3),.dout(w_dff_B_Jj3NHDP84_3),.clk(gclk));
	jdff dff_B_KXnUiTzW5_3(.din(w_dff_B_Jj3NHDP84_3),.dout(w_dff_B_KXnUiTzW5_3),.clk(gclk));
	jdff dff_B_JD2Rz16V0_3(.din(w_dff_B_KXnUiTzW5_3),.dout(w_dff_B_JD2Rz16V0_3),.clk(gclk));
	jdff dff_B_aR637i0J9_3(.din(w_dff_B_JD2Rz16V0_3),.dout(w_dff_B_aR637i0J9_3),.clk(gclk));
	jdff dff_B_TJ6EZ4fW9_3(.din(w_dff_B_aR637i0J9_3),.dout(w_dff_B_TJ6EZ4fW9_3),.clk(gclk));
	jdff dff_B_uJQ2eOXl4_3(.din(w_dff_B_TJ6EZ4fW9_3),.dout(w_dff_B_uJQ2eOXl4_3),.clk(gclk));
	jdff dff_B_0CMEndwP5_3(.din(w_dff_B_uJQ2eOXl4_3),.dout(w_dff_B_0CMEndwP5_3),.clk(gclk));
	jdff dff_B_V69zn5WE9_3(.din(w_dff_B_0CMEndwP5_3),.dout(w_dff_B_V69zn5WE9_3),.clk(gclk));
	jdff dff_B_SbyWKT4c1_3(.din(w_dff_B_V69zn5WE9_3),.dout(w_dff_B_SbyWKT4c1_3),.clk(gclk));
	jdff dff_B_b5gDHqmV4_3(.din(w_dff_B_SbyWKT4c1_3),.dout(w_dff_B_b5gDHqmV4_3),.clk(gclk));
	jdff dff_B_kkRlhK8R5_3(.din(w_dff_B_b5gDHqmV4_3),.dout(w_dff_B_kkRlhK8R5_3),.clk(gclk));
	jdff dff_B_CXby5lLn8_3(.din(w_dff_B_kkRlhK8R5_3),.dout(w_dff_B_CXby5lLn8_3),.clk(gclk));
	jdff dff_B_jh6Pz9Zb5_3(.din(w_dff_B_CXby5lLn8_3),.dout(w_dff_B_jh6Pz9Zb5_3),.clk(gclk));
	jdff dff_B_5R7QQSBq3_3(.din(w_dff_B_jh6Pz9Zb5_3),.dout(w_dff_B_5R7QQSBq3_3),.clk(gclk));
	jdff dff_B_cB0oiWbK4_3(.din(w_dff_B_5R7QQSBq3_3),.dout(w_dff_B_cB0oiWbK4_3),.clk(gclk));
	jdff dff_B_ohEwP5um6_3(.din(w_dff_B_cB0oiWbK4_3),.dout(w_dff_B_ohEwP5um6_3),.clk(gclk));
	jdff dff_B_fJVRGy5q8_3(.din(w_dff_B_ohEwP5um6_3),.dout(w_dff_B_fJVRGy5q8_3),.clk(gclk));
	jdff dff_B_2oZZjT7X1_1(.din(n717),.dout(w_dff_B_2oZZjT7X1_1),.clk(gclk));
	jdff dff_B_KgojfExN2_1(.din(n1451),.dout(w_dff_B_KgojfExN2_1),.clk(gclk));
	jdff dff_B_8UnFFy893_1(.din(w_dff_B_KgojfExN2_1),.dout(w_dff_B_8UnFFy893_1),.clk(gclk));
	jdff dff_B_tuSUn7M79_1(.din(w_dff_B_8UnFFy893_1),.dout(w_dff_B_tuSUn7M79_1),.clk(gclk));
	jdff dff_B_bOcn9bFA5_1(.din(w_dff_B_tuSUn7M79_1),.dout(w_dff_B_bOcn9bFA5_1),.clk(gclk));
	jdff dff_B_rCxV8oK94_1(.din(w_dff_B_bOcn9bFA5_1),.dout(w_dff_B_rCxV8oK94_1),.clk(gclk));
	jdff dff_B_pXv33GAe6_1(.din(w_dff_B_rCxV8oK94_1),.dout(w_dff_B_pXv33GAe6_1),.clk(gclk));
	jdff dff_B_YSYV19dJ5_1(.din(w_dff_B_pXv33GAe6_1),.dout(w_dff_B_YSYV19dJ5_1),.clk(gclk));
	jdff dff_B_ATGUKbGM5_1(.din(w_dff_B_YSYV19dJ5_1),.dout(w_dff_B_ATGUKbGM5_1),.clk(gclk));
	jdff dff_B_SzUDHR6b7_1(.din(w_dff_B_ATGUKbGM5_1),.dout(w_dff_B_SzUDHR6b7_1),.clk(gclk));
	jdff dff_B_LpWTZVwP6_1(.din(w_dff_B_SzUDHR6b7_1),.dout(w_dff_B_LpWTZVwP6_1),.clk(gclk));
	jdff dff_B_p6Dvi9i21_1(.din(w_dff_B_LpWTZVwP6_1),.dout(w_dff_B_p6Dvi9i21_1),.clk(gclk));
	jdff dff_B_oUEGXJvf0_1(.din(w_dff_B_p6Dvi9i21_1),.dout(w_dff_B_oUEGXJvf0_1),.clk(gclk));
	jdff dff_B_5FxkY6i03_1(.din(w_dff_B_oUEGXJvf0_1),.dout(w_dff_B_5FxkY6i03_1),.clk(gclk));
	jdff dff_B_z5Hs1uc00_1(.din(w_dff_B_5FxkY6i03_1),.dout(w_dff_B_z5Hs1uc00_1),.clk(gclk));
	jdff dff_B_yo79W8XW9_1(.din(w_dff_B_z5Hs1uc00_1),.dout(w_dff_B_yo79W8XW9_1),.clk(gclk));
	jdff dff_A_X8KAt6jb7_0(.dout(w_n715_0[0]),.din(w_dff_A_X8KAt6jb7_0),.clk(gclk));
	jdff dff_A_mNktjaKO5_1(.dout(w_n715_0[1]),.din(w_dff_A_mNktjaKO5_1),.clk(gclk));
	jdff dff_A_lX3g4Itf2_0(.dout(w_n1469_0[0]),.din(w_dff_A_lX3g4Itf2_0),.clk(gclk));
	jdff dff_B_dM42cA8C7_2(.din(n1469),.dout(w_dff_B_dM42cA8C7_2),.clk(gclk));
	jdff dff_B_MJTYYIxQ6_2(.din(w_dff_B_dM42cA8C7_2),.dout(w_dff_B_MJTYYIxQ6_2),.clk(gclk));
	jdff dff_B_GXOXjQLM0_2(.din(w_dff_B_MJTYYIxQ6_2),.dout(w_dff_B_GXOXjQLM0_2),.clk(gclk));
	jdff dff_B_zEDiIaCw9_2(.din(w_dff_B_GXOXjQLM0_2),.dout(w_dff_B_zEDiIaCw9_2),.clk(gclk));
	jdff dff_B_G2n4ifS46_2(.din(w_dff_B_zEDiIaCw9_2),.dout(w_dff_B_G2n4ifS46_2),.clk(gclk));
	jdff dff_B_yjrW8SYW8_2(.din(w_dff_B_G2n4ifS46_2),.dout(w_dff_B_yjrW8SYW8_2),.clk(gclk));
	jdff dff_B_ldsqRPJP1_2(.din(w_dff_B_yjrW8SYW8_2),.dout(w_dff_B_ldsqRPJP1_2),.clk(gclk));
	jdff dff_B_AU69szzi5_2(.din(w_dff_B_ldsqRPJP1_2),.dout(w_dff_B_AU69szzi5_2),.clk(gclk));
	jdff dff_B_R8RVR4Em2_2(.din(w_dff_B_AU69szzi5_2),.dout(w_dff_B_R8RVR4Em2_2),.clk(gclk));
	jdff dff_A_ltbWdfQG3_0(.dout(w_n1470_0[0]),.din(w_dff_A_ltbWdfQG3_0),.clk(gclk));
	jdff dff_B_44HkEJvN5_2(.din(n1470),.dout(w_dff_B_44HkEJvN5_2),.clk(gclk));
	jdff dff_B_Qogw2FEU5_2(.din(w_dff_B_44HkEJvN5_2),.dout(w_dff_B_Qogw2FEU5_2),.clk(gclk));
	jdff dff_B_c373aXyp3_2(.din(w_dff_B_Qogw2FEU5_2),.dout(w_dff_B_c373aXyp3_2),.clk(gclk));
	jdff dff_B_G54LPRDw9_2(.din(w_dff_B_c373aXyp3_2),.dout(w_dff_B_G54LPRDw9_2),.clk(gclk));
	jdff dff_B_XD9VrQfq4_2(.din(w_dff_B_G54LPRDw9_2),.dout(w_dff_B_XD9VrQfq4_2),.clk(gclk));
	jdff dff_B_BBr7EVxo5_2(.din(w_dff_B_XD9VrQfq4_2),.dout(w_dff_B_BBr7EVxo5_2),.clk(gclk));
	jdff dff_B_EsLk7yv80_2(.din(w_dff_B_BBr7EVxo5_2),.dout(w_dff_B_EsLk7yv80_2),.clk(gclk));
	jdff dff_B_t0V9Cd6B6_1(.din(n1500),.dout(w_dff_B_t0V9Cd6B6_1),.clk(gclk));
	jdff dff_B_KUAIJL757_1(.din(w_dff_B_t0V9Cd6B6_1),.dout(w_dff_B_KUAIJL757_1),.clk(gclk));
	jdff dff_B_oFG2qDPi6_1(.din(w_dff_B_KUAIJL757_1),.dout(w_dff_B_oFG2qDPi6_1),.clk(gclk));
	jdff dff_B_qu9AU5DH7_1(.din(w_dff_B_oFG2qDPi6_1),.dout(w_dff_B_qu9AU5DH7_1),.clk(gclk));
	jdff dff_B_e1LrZ9FG8_1(.din(w_dff_B_qu9AU5DH7_1),.dout(w_dff_B_e1LrZ9FG8_1),.clk(gclk));
	jdff dff_B_Kqxsl6xq7_1(.din(w_dff_B_e1LrZ9FG8_1),.dout(w_dff_B_Kqxsl6xq7_1),.clk(gclk));
	jdff dff_B_0BdZoDHv6_1(.din(w_dff_B_Kqxsl6xq7_1),.dout(w_dff_B_0BdZoDHv6_1),.clk(gclk));
	jdff dff_B_HtZdZ1D74_1(.din(w_dff_B_0BdZoDHv6_1),.dout(w_dff_B_HtZdZ1D74_1),.clk(gclk));
	jdff dff_B_iCMngwBU5_1(.din(w_dff_B_HtZdZ1D74_1),.dout(w_dff_B_iCMngwBU5_1),.clk(gclk));
	jdff dff_B_d5fv3hk86_1(.din(w_dff_B_iCMngwBU5_1),.dout(w_dff_B_d5fv3hk86_1),.clk(gclk));
	jdff dff_B_SoWd5YXX4_1(.din(w_dff_B_d5fv3hk86_1),.dout(w_dff_B_SoWd5YXX4_1),.clk(gclk));
	jdff dff_B_ryspUru82_1(.din(w_dff_B_SoWd5YXX4_1),.dout(w_dff_B_ryspUru82_1),.clk(gclk));
	jdff dff_B_aYOpmNQu3_1(.din(w_dff_B_ryspUru82_1),.dout(w_dff_B_aYOpmNQu3_1),.clk(gclk));
	jdff dff_B_9zrF3Isv5_1(.din(w_dff_B_aYOpmNQu3_1),.dout(w_dff_B_9zrF3Isv5_1),.clk(gclk));
	jdff dff_B_U8EmEL2h4_1(.din(w_dff_B_9zrF3Isv5_1),.dout(w_dff_B_U8EmEL2h4_1),.clk(gclk));
	jdff dff_B_LNzOzkYx4_0(.din(n1546),.dout(w_dff_B_LNzOzkYx4_0),.clk(gclk));
	jdff dff_B_gnBCZDhH4_0(.din(w_dff_B_LNzOzkYx4_0),.dout(w_dff_B_gnBCZDhH4_0),.clk(gclk));
	jdff dff_B_J5xJEgnn2_0(.din(n1544),.dout(w_dff_B_J5xJEgnn2_0),.clk(gclk));
	jdff dff_B_QTp7Gtxt6_0(.din(w_dff_B_J5xJEgnn2_0),.dout(w_dff_B_QTp7Gtxt6_0),.clk(gclk));
	jdff dff_B_xR1d7E2a2_1(.din(n1533),.dout(w_dff_B_xR1d7E2a2_1),.clk(gclk));
	jdff dff_B_u3cQHpfZ3_1(.din(w_dff_B_xR1d7E2a2_1),.dout(w_dff_B_u3cQHpfZ3_1),.clk(gclk));
	jdff dff_B_AM7IyKHC6_1(.din(w_dff_B_u3cQHpfZ3_1),.dout(w_dff_B_AM7IyKHC6_1),.clk(gclk));
	jdff dff_B_aI1HuN814_1(.din(w_dff_B_AM7IyKHC6_1),.dout(w_dff_B_aI1HuN814_1),.clk(gclk));
	jdff dff_B_HkRHqI9f6_1(.din(n1534),.dout(w_dff_B_HkRHqI9f6_1),.clk(gclk));
	jdff dff_B_V4RiUXRg5_1(.din(w_dff_B_HkRHqI9f6_1),.dout(w_dff_B_V4RiUXRg5_1),.clk(gclk));
	jdff dff_B_AF1N2f3f8_1(.din(w_dff_B_V4RiUXRg5_1),.dout(w_dff_B_AF1N2f3f8_1),.clk(gclk));
	jdff dff_B_RAz5LPa67_1(.din(w_dff_B_AF1N2f3f8_1),.dout(w_dff_B_RAz5LPa67_1),.clk(gclk));
	jdff dff_B_PSFf9n4w9_1(.din(w_dff_B_RAz5LPa67_1),.dout(w_dff_B_PSFf9n4w9_1),.clk(gclk));
	jdff dff_B_HFTzXLQg0_1(.din(w_dff_B_PSFf9n4w9_1),.dout(w_dff_B_HFTzXLQg0_1),.clk(gclk));
	jdff dff_B_PYhRQtCE6_1(.din(w_dff_B_HFTzXLQg0_1),.dout(w_dff_B_PYhRQtCE6_1),.clk(gclk));
	jdff dff_B_X1okK80g2_1(.din(n1538),.dout(w_dff_B_X1okK80g2_1),.clk(gclk));
	jdff dff_B_aeoxuii34_0(.din(n1540),.dout(w_dff_B_aeoxuii34_0),.clk(gclk));
	jdff dff_B_Nh6WyFZo2_1(.din(n1539),.dout(w_dff_B_Nh6WyFZo2_1),.clk(gclk));
	jdff dff_B_xVxqDQz99_0(.din(n1535),.dout(w_dff_B_xVxqDQz99_0),.clk(gclk));
	jdff dff_A_189A6ZlH4_1(.dout(w_n1414_0[1]),.din(w_dff_A_189A6ZlH4_1),.clk(gclk));
	jdff dff_A_eTuTsUzN9_1(.dout(w_dff_A_189A6ZlH4_1),.din(w_dff_A_eTuTsUzN9_1),.clk(gclk));
	jdff dff_A_YeVLCuEd5_1(.dout(w_dff_A_eTuTsUzN9_1),.din(w_dff_A_YeVLCuEd5_1),.clk(gclk));
	jdff dff_A_7Sb9knEw0_1(.dout(w_dff_A_YeVLCuEd5_1),.din(w_dff_A_7Sb9knEw0_1),.clk(gclk));
	jdff dff_A_sBamll1V9_1(.dout(w_dff_A_7Sb9knEw0_1),.din(w_dff_A_sBamll1V9_1),.clk(gclk));
	jdff dff_A_pWlNBqqc1_1(.dout(w_dff_A_sBamll1V9_1),.din(w_dff_A_pWlNBqqc1_1),.clk(gclk));
	jdff dff_A_HTXHixWY6_1(.dout(w_dff_A_pWlNBqqc1_1),.din(w_dff_A_HTXHixWY6_1),.clk(gclk));
	jdff dff_A_qm6gHRym3_1(.dout(w_dff_A_HTXHixWY6_1),.din(w_dff_A_qm6gHRym3_1),.clk(gclk));
	jdff dff_A_buTZcA207_1(.dout(w_dff_A_qm6gHRym3_1),.din(w_dff_A_buTZcA207_1),.clk(gclk));
	jdff dff_A_gQJETuFf1_1(.dout(w_dff_A_buTZcA207_1),.din(w_dff_A_gQJETuFf1_1),.clk(gclk));
	jdff dff_B_Qst8B18I0_1(.din(n1412),.dout(w_dff_B_Qst8B18I0_1),.clk(gclk));
	jdff dff_A_WVjGtuSH1_1(.dout(w_n1404_0[1]),.din(w_dff_A_WVjGtuSH1_1),.clk(gclk));
	jdff dff_A_mLbPJ5GU7_1(.dout(w_dff_A_WVjGtuSH1_1),.din(w_dff_A_mLbPJ5GU7_1),.clk(gclk));
	jdff dff_A_OEGK5aPO0_1(.dout(w_dff_A_mLbPJ5GU7_1),.din(w_dff_A_OEGK5aPO0_1),.clk(gclk));
	jdff dff_A_cA44UuRA4_1(.dout(w_dff_A_OEGK5aPO0_1),.din(w_dff_A_cA44UuRA4_1),.clk(gclk));
	jdff dff_A_dtyJ8XnP2_1(.dout(w_dff_A_cA44UuRA4_1),.din(w_dff_A_dtyJ8XnP2_1),.clk(gclk));
	jdff dff_A_JTWpSgbv7_1(.dout(w_dff_A_dtyJ8XnP2_1),.din(w_dff_A_JTWpSgbv7_1),.clk(gclk));
	jdff dff_A_TMhhQwq76_1(.dout(w_dff_A_JTWpSgbv7_1),.din(w_dff_A_TMhhQwq76_1),.clk(gclk));
	jdff dff_A_sy9AdmYK5_1(.dout(w_dff_A_TMhhQwq76_1),.din(w_dff_A_sy9AdmYK5_1),.clk(gclk));
	jdff dff_A_SuUZyTFP8_1(.dout(w_dff_A_sy9AdmYK5_1),.din(w_dff_A_SuUZyTFP8_1),.clk(gclk));
	jdff dff_B_KlXKBtaX3_2(.din(n1404),.dout(w_dff_B_KlXKBtaX3_2),.clk(gclk));
	jdff dff_B_cUKLYI2q2_0(.din(n1530),.dout(w_dff_B_cUKLYI2q2_0),.clk(gclk));
	jdff dff_B_LMw4H1BS8_0(.din(w_dff_B_cUKLYI2q2_0),.dout(w_dff_B_LMw4H1BS8_0),.clk(gclk));
	jdff dff_B_nHV2rcZB0_0(.din(w_dff_B_LMw4H1BS8_0),.dout(w_dff_B_nHV2rcZB0_0),.clk(gclk));
	jdff dff_B_3Z2683L62_1(.din(n1524),.dout(w_dff_B_3Z2683L62_1),.clk(gclk));
	jdff dff_B_INRxn0Zf8_1(.din(w_dff_B_3Z2683L62_1),.dout(w_dff_B_INRxn0Zf8_1),.clk(gclk));
	jdff dff_B_qYyCQUq50_0(.din(n1527),.dout(w_dff_B_qYyCQUq50_0),.clk(gclk));
	jdff dff_B_puz4657M8_0(.din(w_dff_B_qYyCQUq50_0),.dout(w_dff_B_puz4657M8_0),.clk(gclk));
	jdff dff_B_h1hNkmOI9_0(.din(w_dff_B_puz4657M8_0),.dout(w_dff_B_h1hNkmOI9_0),.clk(gclk));
	jdff dff_B_WS9Io77u8_1(.din(n1525),.dout(w_dff_B_WS9Io77u8_1),.clk(gclk));
	jdff dff_A_t08G5Bbe2_1(.dout(w_n1401_0[1]),.din(w_dff_A_t08G5Bbe2_1),.clk(gclk));
	jdff dff_A_LJD4TZIk5_1(.dout(w_dff_A_t08G5Bbe2_1),.din(w_dff_A_LJD4TZIk5_1),.clk(gclk));
	jdff dff_A_N9e8tcqr4_1(.dout(w_dff_A_LJD4TZIk5_1),.din(w_dff_A_N9e8tcqr4_1),.clk(gclk));
	jdff dff_A_F0FfSBz80_1(.dout(w_dff_A_N9e8tcqr4_1),.din(w_dff_A_F0FfSBz80_1),.clk(gclk));
	jdff dff_A_B62EhZho3_1(.dout(w_dff_A_F0FfSBz80_1),.din(w_dff_A_B62EhZho3_1),.clk(gclk));
	jdff dff_A_gKREzjCS2_1(.dout(w_dff_A_B62EhZho3_1),.din(w_dff_A_gKREzjCS2_1),.clk(gclk));
	jdff dff_A_iasVbBSK8_1(.dout(w_dff_A_gKREzjCS2_1),.din(w_dff_A_iasVbBSK8_1),.clk(gclk));
	jdff dff_A_zCPEnLGe2_1(.dout(w_dff_A_iasVbBSK8_1),.din(w_dff_A_zCPEnLGe2_1),.clk(gclk));
	jdff dff_A_HnnnsTka4_1(.dout(w_dff_A_zCPEnLGe2_1),.din(w_dff_A_HnnnsTka4_1),.clk(gclk));
	jdff dff_B_kXOVzd9I2_2(.din(n1401),.dout(w_dff_B_kXOVzd9I2_2),.clk(gclk));
	jdff dff_B_HTieYIFO7_2(.din(w_dff_B_kXOVzd9I2_2),.dout(w_dff_B_HTieYIFO7_2),.clk(gclk));
	jdff dff_B_nevWWI0v8_2(.din(w_dff_B_HTieYIFO7_2),.dout(w_dff_B_nevWWI0v8_2),.clk(gclk));
	jdff dff_B_iSRBWQMZ6_2(.din(w_dff_B_nevWWI0v8_2),.dout(w_dff_B_iSRBWQMZ6_2),.clk(gclk));
	jdff dff_B_NIXbY9Ao0_2(.din(w_dff_B_iSRBWQMZ6_2),.dout(w_dff_B_NIXbY9Ao0_2),.clk(gclk));
	jdff dff_B_WUarIzIc6_2(.din(w_dff_B_NIXbY9Ao0_2),.dout(w_dff_B_WUarIzIc6_2),.clk(gclk));
	jdff dff_A_kUmEGgAQ2_1(.dout(w_n1520_0[1]),.din(w_dff_A_kUmEGgAQ2_1),.clk(gclk));
	jdff dff_B_bKnFP9Jd3_0(.din(n1516),.dout(w_dff_B_bKnFP9Jd3_0),.clk(gclk));
	jdff dff_B_majlC20b5_0(.din(w_dff_B_bKnFP9Jd3_0),.dout(w_dff_B_majlC20b5_0),.clk(gclk));
	jdff dff_B_gLo6NdRF1_0(.din(w_dff_B_majlC20b5_0),.dout(w_dff_B_gLo6NdRF1_0),.clk(gclk));
	jdff dff_B_Mm9GiAn24_0(.din(w_dff_B_gLo6NdRF1_0),.dout(w_dff_B_Mm9GiAn24_0),.clk(gclk));
	jdff dff_B_qRoOA2Qd9_0(.din(w_dff_B_Mm9GiAn24_0),.dout(w_dff_B_qRoOA2Qd9_0),.clk(gclk));
	jdff dff_B_UMNJLbhl3_1(.din(n1509),.dout(w_dff_B_UMNJLbhl3_1),.clk(gclk));
	jdff dff_B_4Vp9XJcD5_1(.din(w_dff_B_UMNJLbhl3_1),.dout(w_dff_B_4Vp9XJcD5_1),.clk(gclk));
	jdff dff_B_9THo75lP0_1(.din(w_dff_B_4Vp9XJcD5_1),.dout(w_dff_B_9THo75lP0_1),.clk(gclk));
	jdff dff_B_7Hmehq3E6_1(.din(w_dff_B_9THo75lP0_1),.dout(w_dff_B_7Hmehq3E6_1),.clk(gclk));
	jdff dff_B_r8AFxmE49_1(.din(w_dff_B_7Hmehq3E6_1),.dout(w_dff_B_r8AFxmE49_1),.clk(gclk));
	jdff dff_B_jMIpVqyN4_1(.din(w_dff_B_r8AFxmE49_1),.dout(w_dff_B_jMIpVqyN4_1),.clk(gclk));
	jdff dff_B_WfMAqJW37_0(.din(n1513),.dout(w_dff_B_WfMAqJW37_0),.clk(gclk));
	jdff dff_A_wXk9aqtR3_1(.dout(w_n1445_0[1]),.din(w_dff_A_wXk9aqtR3_1),.clk(gclk));
	jdff dff_A_C957GCgo6_1(.dout(w_dff_A_wXk9aqtR3_1),.din(w_dff_A_C957GCgo6_1),.clk(gclk));
	jdff dff_A_4vVxTJGK5_1(.dout(w_dff_A_C957GCgo6_1),.din(w_dff_A_4vVxTJGK5_1),.clk(gclk));
	jdff dff_A_fBWZPxuy6_1(.dout(w_dff_A_4vVxTJGK5_1),.din(w_dff_A_fBWZPxuy6_1),.clk(gclk));
	jdff dff_A_fTYnZjd86_1(.dout(w_dff_A_fBWZPxuy6_1),.din(w_dff_A_fTYnZjd86_1),.clk(gclk));
	jdff dff_A_twiNsobd1_1(.dout(w_dff_A_fTYnZjd86_1),.din(w_dff_A_twiNsobd1_1),.clk(gclk));
	jdff dff_A_Ad1WD2fp6_1(.dout(w_dff_A_twiNsobd1_1),.din(w_dff_A_Ad1WD2fp6_1),.clk(gclk));
	jdff dff_A_se79etU97_1(.dout(w_dff_A_Ad1WD2fp6_1),.din(w_dff_A_se79etU97_1),.clk(gclk));
	jdff dff_A_pOl1XUOm4_1(.dout(w_dff_A_se79etU97_1),.din(w_dff_A_pOl1XUOm4_1),.clk(gclk));
	jdff dff_A_JL2dJkcJ1_1(.dout(w_dff_A_pOl1XUOm4_1),.din(w_dff_A_JL2dJkcJ1_1),.clk(gclk));
	jdff dff_A_vE50oDBr4_1(.dout(w_dff_A_JL2dJkcJ1_1),.din(w_dff_A_vE50oDBr4_1),.clk(gclk));
	jdff dff_B_UthSIp5O4_2(.din(n1445),.dout(w_dff_B_UthSIp5O4_2),.clk(gclk));
	jdff dff_B_8ozVRkdB5_0(.din(n1507),.dout(w_dff_B_8ozVRkdB5_0),.clk(gclk));
	jdff dff_B_eAaxFN4c8_0(.din(w_dff_B_8ozVRkdB5_0),.dout(w_dff_B_eAaxFN4c8_0),.clk(gclk));
	jdff dff_B_GRpiWZ8t0_0(.din(w_dff_B_eAaxFN4c8_0),.dout(w_dff_B_GRpiWZ8t0_0),.clk(gclk));
	jdff dff_B_sJXleZJV5_0(.din(w_dff_B_GRpiWZ8t0_0),.dout(w_dff_B_sJXleZJV5_0),.clk(gclk));
	jdff dff_B_82qNFKIF8_0(.din(w_dff_B_sJXleZJV5_0),.dout(w_dff_B_82qNFKIF8_0),.clk(gclk));
	jdff dff_B_B5qAVPdK2_0(.din(w_dff_B_82qNFKIF8_0),.dout(w_dff_B_B5qAVPdK2_0),.clk(gclk));
	jdff dff_B_KoHBeDLk7_0(.din(n1503),.dout(w_dff_B_KoHBeDLk7_0),.clk(gclk));
	jdff dff_A_xqicetMq9_0(.dout(w_n1444_0[0]),.din(w_dff_A_xqicetMq9_0),.clk(gclk));
	jdff dff_A_tj41q6wh8_0(.dout(w_dff_A_xqicetMq9_0),.din(w_dff_A_tj41q6wh8_0),.clk(gclk));
	jdff dff_A_E6LFlpmq0_2(.dout(w_n1444_0[2]),.din(w_dff_A_E6LFlpmq0_2),.clk(gclk));
	jdff dff_A_k9KSXCIp0_2(.dout(w_dff_A_E6LFlpmq0_2),.din(w_dff_A_k9KSXCIp0_2),.clk(gclk));
	jdff dff_A_VYR4DypP3_2(.dout(w_dff_A_k9KSXCIp0_2),.din(w_dff_A_VYR4DypP3_2),.clk(gclk));
	jdff dff_A_73fzXHMZ8_2(.dout(w_dff_A_VYR4DypP3_2),.din(w_dff_A_73fzXHMZ8_2),.clk(gclk));
	jdff dff_A_PxD9yZqd5_2(.dout(w_dff_A_73fzXHMZ8_2),.din(w_dff_A_PxD9yZqd5_2),.clk(gclk));
	jdff dff_A_w0Iz6dlr5_2(.dout(w_dff_A_PxD9yZqd5_2),.din(w_dff_A_w0Iz6dlr5_2),.clk(gclk));
	jdff dff_A_XqWRHUXo0_2(.dout(w_dff_A_w0Iz6dlr5_2),.din(w_dff_A_XqWRHUXo0_2),.clk(gclk));
	jdff dff_A_DW5A0erl8_2(.dout(w_dff_A_XqWRHUXo0_2),.din(w_dff_A_DW5A0erl8_2),.clk(gclk));
	jdff dff_A_BwmJgd5x7_2(.dout(w_dff_A_DW5A0erl8_2),.din(w_dff_A_BwmJgd5x7_2),.clk(gclk));
	jdff dff_A_SLMe2BuB5_2(.dout(w_dff_A_BwmJgd5x7_2),.din(w_dff_A_SLMe2BuB5_2),.clk(gclk));
	jdff dff_A_uAmDQLEZ8_2(.dout(w_dff_A_SLMe2BuB5_2),.din(w_dff_A_uAmDQLEZ8_2),.clk(gclk));
	jdff dff_A_NSIIuSUk2_2(.dout(w_dff_A_uAmDQLEZ8_2),.din(w_dff_A_NSIIuSUk2_2),.clk(gclk));
	jdff dff_A_dlooAmvU0_2(.dout(w_dff_A_NSIIuSUk2_2),.din(w_dff_A_dlooAmvU0_2),.clk(gclk));
	jdff dff_B_bRi3SU7w6_3(.din(n1444),.dout(w_dff_B_bRi3SU7w6_3),.clk(gclk));
	jdff dff_B_Mb7QQDlE8_3(.din(w_dff_B_bRi3SU7w6_3),.dout(w_dff_B_Mb7QQDlE8_3),.clk(gclk));
	jdff dff_B_atMmZB8Y1_3(.din(w_dff_B_Mb7QQDlE8_3),.dout(w_dff_B_atMmZB8Y1_3),.clk(gclk));
	jdff dff_B_SI0CUn5e3_3(.din(w_dff_B_atMmZB8Y1_3),.dout(w_dff_B_SI0CUn5e3_3),.clk(gclk));
	jdff dff_A_BIyh4ZNm7_1(.dout(w_n1501_0[1]),.din(w_dff_A_BIyh4ZNm7_1),.clk(gclk));
	jdff dff_A_bU0yKjex8_1(.dout(w_dff_A_BIyh4ZNm7_1),.din(w_dff_A_bU0yKjex8_1),.clk(gclk));
	jdff dff_A_garw6vSx8_1(.dout(w_dff_A_bU0yKjex8_1),.din(w_dff_A_garw6vSx8_1),.clk(gclk));
	jdff dff_A_0bdyKZb81_1(.dout(w_dff_A_garw6vSx8_1),.din(w_dff_A_0bdyKZb81_1),.clk(gclk));
	jdff dff_A_iatti9uZ2_1(.dout(w_dff_A_0bdyKZb81_1),.din(w_dff_A_iatti9uZ2_1),.clk(gclk));
	jdff dff_A_2EEXSPAA6_1(.dout(w_n1454_0[1]),.din(w_dff_A_2EEXSPAA6_1),.clk(gclk));
	jdff dff_A_54ofLsbF8_1(.dout(w_dff_A_2EEXSPAA6_1),.din(w_dff_A_54ofLsbF8_1),.clk(gclk));
	jdff dff_A_7jKDsxoq3_1(.dout(w_dff_A_54ofLsbF8_1),.din(w_dff_A_7jKDsxoq3_1),.clk(gclk));
	jdff dff_A_O2xzF8Dh2_1(.dout(w_dff_A_7jKDsxoq3_1),.din(w_dff_A_O2xzF8Dh2_1),.clk(gclk));
	jdff dff_A_8QDMDMFw1_1(.dout(w_dff_A_O2xzF8Dh2_1),.din(w_dff_A_8QDMDMFw1_1),.clk(gclk));
	jdff dff_A_mvDqumTc6_1(.dout(w_dff_A_8QDMDMFw1_1),.din(w_dff_A_mvDqumTc6_1),.clk(gclk));
	jdff dff_A_uX2DG70z2_1(.dout(w_dff_A_mvDqumTc6_1),.din(w_dff_A_uX2DG70z2_1),.clk(gclk));
	jdff dff_B_jNmrxi3S8_2(.din(n1454),.dout(w_dff_B_jNmrxi3S8_2),.clk(gclk));
	jdff dff_B_cZdZCxDD9_2(.din(w_dff_B_jNmrxi3S8_2),.dout(w_dff_B_cZdZCxDD9_2),.clk(gclk));
	jdff dff_B_Nc8LrthW4_2(.din(w_dff_B_cZdZCxDD9_2),.dout(w_dff_B_Nc8LrthW4_2),.clk(gclk));
	jdff dff_B_sThnjLOW4_2(.din(w_dff_B_Nc8LrthW4_2),.dout(w_dff_B_sThnjLOW4_2),.clk(gclk));
	jdff dff_B_2jMqZwdh5_2(.din(w_dff_B_sThnjLOW4_2),.dout(w_dff_B_2jMqZwdh5_2),.clk(gclk));
	jdff dff_B_kyfv9RBk3_0(.din(n1584),.dout(w_dff_B_kyfv9RBk3_0),.clk(gclk));
	jdff dff_B_qMcc0HEP6_0(.din(w_dff_B_kyfv9RBk3_0),.dout(w_dff_B_qMcc0HEP6_0),.clk(gclk));
	jdff dff_B_YLdHd6tD0_0(.din(w_dff_B_qMcc0HEP6_0),.dout(w_dff_B_YLdHd6tD0_0),.clk(gclk));
	jdff dff_B_9YfKdWK08_1(.din(n1561),.dout(w_dff_B_9YfKdWK08_1),.clk(gclk));
	jdff dff_B_UQKYH9Ol9_1(.din(w_dff_B_9YfKdWK08_1),.dout(w_dff_B_UQKYH9Ol9_1),.clk(gclk));
	jdff dff_B_zccf1NQR1_1(.din(w_dff_B_UQKYH9Ol9_1),.dout(w_dff_B_zccf1NQR1_1),.clk(gclk));
	jdff dff_B_DsDLv6TT5_1(.din(w_dff_B_zccf1NQR1_1),.dout(w_dff_B_DsDLv6TT5_1),.clk(gclk));
	jdff dff_B_Kf49E3wu8_1(.din(w_dff_B_DsDLv6TT5_1),.dout(w_dff_B_Kf49E3wu8_1),.clk(gclk));
	jdff dff_B_XjMt2yO34_1(.din(w_dff_B_Kf49E3wu8_1),.dout(w_dff_B_XjMt2yO34_1),.clk(gclk));
	jdff dff_B_SySFhhGT3_1(.din(w_dff_B_XjMt2yO34_1),.dout(w_dff_B_SySFhhGT3_1),.clk(gclk));
	jdff dff_B_cNLpmMdh9_1(.din(w_dff_B_SySFhhGT3_1),.dout(w_dff_B_cNLpmMdh9_1),.clk(gclk));
	jdff dff_B_MGzbcxmn3_1(.din(w_dff_B_cNLpmMdh9_1),.dout(w_dff_B_MGzbcxmn3_1),.clk(gclk));
	jdff dff_B_JUnEuirv2_1(.din(w_dff_B_MGzbcxmn3_1),.dout(w_dff_B_JUnEuirv2_1),.clk(gclk));
	jdff dff_B_BhTQqvKk4_1(.din(w_dff_B_JUnEuirv2_1),.dout(w_dff_B_BhTQqvKk4_1),.clk(gclk));
	jdff dff_B_OKiIDr9X6_1(.din(w_dff_B_BhTQqvKk4_1),.dout(w_dff_B_OKiIDr9X6_1),.clk(gclk));
	jdff dff_B_2O444AIl1_1(.din(w_dff_B_OKiIDr9X6_1),.dout(w_dff_B_2O444AIl1_1),.clk(gclk));
	jdff dff_B_EsPNKSXH3_1(.din(w_dff_B_2O444AIl1_1),.dout(w_dff_B_EsPNKSXH3_1),.clk(gclk));
	jdff dff_B_p4HONLhX2_1(.din(w_dff_B_EsPNKSXH3_1),.dout(w_dff_B_p4HONLhX2_1),.clk(gclk));
	jdff dff_B_x2kVBAV96_1(.din(w_dff_B_p4HONLhX2_1),.dout(w_dff_B_x2kVBAV96_1),.clk(gclk));
	jdff dff_B_8qb9JnrM6_1(.din(w_dff_B_x2kVBAV96_1),.dout(w_dff_B_8qb9JnrM6_1),.clk(gclk));
	jdff dff_B_bVCbw5jP6_0(.din(n1581),.dout(w_dff_B_bVCbw5jP6_0),.clk(gclk));
	jdff dff_B_7FIOKbKe8_0(.din(w_dff_B_bVCbw5jP6_0),.dout(w_dff_B_7FIOKbKe8_0),.clk(gclk));
	jdff dff_B_9zCOOAxD2_0(.din(n1578),.dout(w_dff_B_9zCOOAxD2_0),.clk(gclk));
	jdff dff_B_92bLwit86_0(.din(w_dff_B_9zCOOAxD2_0),.dout(w_dff_B_92bLwit86_0),.clk(gclk));
	jdff dff_B_1nNq9ubr4_0(.din(w_dff_B_92bLwit86_0),.dout(w_dff_B_1nNq9ubr4_0),.clk(gclk));
	jdff dff_B_WYKqQNdS8_0(.din(w_dff_B_1nNq9ubr4_0),.dout(w_dff_B_WYKqQNdS8_0),.clk(gclk));
	jdff dff_B_jgRtkKpr3_0(.din(w_dff_B_WYKqQNdS8_0),.dout(w_dff_B_jgRtkKpr3_0),.clk(gclk));
	jdff dff_B_E5nqfP4x2_0(.din(w_dff_B_jgRtkKpr3_0),.dout(w_dff_B_E5nqfP4x2_0),.clk(gclk));
	jdff dff_B_F2TP6eVx6_1(.din(n1572),.dout(w_dff_B_F2TP6eVx6_1),.clk(gclk));
	jdff dff_B_cPEWPHhX5_1(.din(w_dff_B_F2TP6eVx6_1),.dout(w_dff_B_cPEWPHhX5_1),.clk(gclk));
	jdff dff_B_AQXSGaOY9_1(.din(w_dff_B_cPEWPHhX5_1),.dout(w_dff_B_AQXSGaOY9_1),.clk(gclk));
	jdff dff_B_Jdd7TguC6_0(.din(n1574),.dout(w_dff_B_Jdd7TguC6_0),.clk(gclk));
	jdff dff_B_AsBXhVOA6_0(.din(n1570),.dout(w_dff_B_AsBXhVOA6_0),.clk(gclk));
	jdff dff_B_gtqeDLaA1_0(.din(w_dff_B_AsBXhVOA6_0),.dout(w_dff_B_gtqeDLaA1_0),.clk(gclk));
	jdff dff_B_qUMsoeRw8_0(.din(n1568),.dout(w_dff_B_qUMsoeRw8_0),.clk(gclk));
	jdff dff_B_54ePHx2p1_0(.din(w_dff_B_qUMsoeRw8_0),.dout(w_dff_B_54ePHx2p1_0),.clk(gclk));
	jdff dff_B_VuDupfmp4_0(.din(w_dff_B_54ePHx2p1_0),.dout(w_dff_B_VuDupfmp4_0),.clk(gclk));
	jdff dff_B_UXMno1W47_0(.din(w_dff_B_VuDupfmp4_0),.dout(w_dff_B_UXMno1W47_0),.clk(gclk));
	jdff dff_B_eqgWUqGr2_0(.din(w_dff_B_UXMno1W47_0),.dout(w_dff_B_eqgWUqGr2_0),.clk(gclk));
	jdff dff_B_d7qp4tb85_0(.din(w_dff_B_eqgWUqGr2_0),.dout(w_dff_B_d7qp4tb85_0),.clk(gclk));
	jdff dff_B_11Q2SXGH8_0(.din(n1567),.dout(w_dff_B_11Q2SXGH8_0),.clk(gclk));
	jdff dff_B_g6FwZoqP4_0(.din(w_dff_B_11Q2SXGH8_0),.dout(w_dff_B_g6FwZoqP4_0),.clk(gclk));
	jdff dff_B_oJAojJul3_0(.din(w_dff_B_g6FwZoqP4_0),.dout(w_dff_B_oJAojJul3_0),.clk(gclk));
	jdff dff_B_7T2CMOVL2_0(.din(w_dff_B_oJAojJul3_0),.dout(w_dff_B_7T2CMOVL2_0),.clk(gclk));
	jdff dff_B_qqXNUt202_0(.din(w_dff_B_7T2CMOVL2_0),.dout(w_dff_B_qqXNUt202_0),.clk(gclk));
	jdff dff_B_ESh5Qf9G8_0(.din(n1566),.dout(w_dff_B_ESh5Qf9G8_0),.clk(gclk));
	jdff dff_B_zxuyijCv3_0(.din(w_dff_B_ESh5Qf9G8_0),.dout(w_dff_B_zxuyijCv3_0),.clk(gclk));
	jdff dff_B_XZZm6ftf0_0(.din(n1562),.dout(w_dff_B_XZZm6ftf0_0),.clk(gclk));
	jdff dff_A_PXGPS2LS4_1(.dout(w_n1420_0[1]),.din(w_dff_A_PXGPS2LS4_1),.clk(gclk));
	jdff dff_A_1W9ogM5S2_1(.dout(w_dff_A_PXGPS2LS4_1),.din(w_dff_A_1W9ogM5S2_1),.clk(gclk));
	jdff dff_A_YAhy02zL6_1(.dout(w_dff_A_1W9ogM5S2_1),.din(w_dff_A_YAhy02zL6_1),.clk(gclk));
	jdff dff_A_hJn7yT7j7_1(.dout(w_dff_A_YAhy02zL6_1),.din(w_dff_A_hJn7yT7j7_1),.clk(gclk));
	jdff dff_A_KuhxwjDN7_2(.dout(w_n1420_0[2]),.din(w_dff_A_KuhxwjDN7_2),.clk(gclk));
	jdff dff_A_9B3hDVd52_2(.dout(w_dff_A_KuhxwjDN7_2),.din(w_dff_A_9B3hDVd52_2),.clk(gclk));
	jdff dff_A_VRs2VgW55_2(.dout(w_dff_A_9B3hDVd52_2),.din(w_dff_A_VRs2VgW55_2),.clk(gclk));
	jdff dff_A_uEyEvH4i8_2(.dout(w_dff_A_VRs2VgW55_2),.din(w_dff_A_uEyEvH4i8_2),.clk(gclk));
	jdff dff_A_mTIZ4Kb78_2(.dout(w_dff_A_uEyEvH4i8_2),.din(w_dff_A_mTIZ4Kb78_2),.clk(gclk));
	jdff dff_A_TwBweXs65_2(.dout(w_dff_A_mTIZ4Kb78_2),.din(w_dff_A_TwBweXs65_2),.clk(gclk));
	jdff dff_A_yFR6T61W9_2(.dout(w_dff_A_TwBweXs65_2),.din(w_dff_A_yFR6T61W9_2),.clk(gclk));
	jdff dff_A_LOyNwaeG2_2(.dout(w_dff_A_yFR6T61W9_2),.din(w_dff_A_LOyNwaeG2_2),.clk(gclk));
	jdff dff_A_0VUNrvOx1_2(.dout(w_dff_A_LOyNwaeG2_2),.din(w_dff_A_0VUNrvOx1_2),.clk(gclk));
	jdff dff_A_K9bwiR2B9_2(.dout(w_dff_A_0VUNrvOx1_2),.din(w_dff_A_K9bwiR2B9_2),.clk(gclk));
	jdff dff_A_o0RjupcQ4_2(.dout(w_dff_A_K9bwiR2B9_2),.din(w_dff_A_o0RjupcQ4_2),.clk(gclk));
	jdff dff_A_5Ppzryr87_2(.dout(w_dff_A_o0RjupcQ4_2),.din(w_dff_A_5Ppzryr87_2),.clk(gclk));
	jdff dff_A_D2lhm79R9_2(.dout(w_dff_A_5Ppzryr87_2),.din(w_dff_A_D2lhm79R9_2),.clk(gclk));
	jdff dff_A_whQeeJ9W9_2(.dout(w_dff_A_D2lhm79R9_2),.din(w_dff_A_whQeeJ9W9_2),.clk(gclk));
	jdff dff_A_LDUmc2re1_2(.dout(w_dff_A_whQeeJ9W9_2),.din(w_dff_A_LDUmc2re1_2),.clk(gclk));
	jdff dff_A_t7v2Foso9_2(.dout(w_dff_A_LDUmc2re1_2),.din(w_dff_A_t7v2Foso9_2),.clk(gclk));
	jdff dff_B_riTkMIhQ1_3(.din(n1420),.dout(w_dff_B_riTkMIhQ1_3),.clk(gclk));
	jdff dff_B_BA6ypliL0_3(.din(w_dff_B_riTkMIhQ1_3),.dout(w_dff_B_BA6ypliL0_3),.clk(gclk));
	jdff dff_B_prn8QpJd1_3(.din(w_dff_B_BA6ypliL0_3),.dout(w_dff_B_prn8QpJd1_3),.clk(gclk));
	jdff dff_B_uP0Es38F6_0(.din(n1559),.dout(w_dff_B_uP0Es38F6_0),.clk(gclk));
	jdff dff_B_ySHsmOrS1_0(.din(w_dff_B_uP0Es38F6_0),.dout(w_dff_B_ySHsmOrS1_0),.clk(gclk));
	jdff dff_B_p8TN8DnC6_0(.din(w_dff_B_ySHsmOrS1_0),.dout(w_dff_B_p8TN8DnC6_0),.clk(gclk));
	jdff dff_B_PI4UAjCe7_0(.din(w_dff_B_p8TN8DnC6_0),.dout(w_dff_B_PI4UAjCe7_0),.clk(gclk));
	jdff dff_B_ULeS2Hdb5_0(.din(n1558),.dout(w_dff_B_ULeS2Hdb5_0),.clk(gclk));
	jdff dff_B_8MufqKta2_0(.din(w_dff_B_ULeS2Hdb5_0),.dout(w_dff_B_8MufqKta2_0),.clk(gclk));
	jdff dff_B_BFXyUr5n4_0(.din(w_dff_B_8MufqKta2_0),.dout(w_dff_B_BFXyUr5n4_0),.clk(gclk));
	jdff dff_B_xS7EoXhY9_0(.din(w_dff_B_BFXyUr5n4_0),.dout(w_dff_B_xS7EoXhY9_0),.clk(gclk));
	jdff dff_B_M7sTA4wo4_0(.din(n1556),.dout(w_dff_B_M7sTA4wo4_0),.clk(gclk));
	jdff dff_B_WMdstgmH6_0(.din(n1554),.dout(w_dff_B_WMdstgmH6_0),.clk(gclk));
	jdff dff_B_dQ2XVzZb1_0(.din(w_dff_B_WMdstgmH6_0),.dout(w_dff_B_dQ2XVzZb1_0),.clk(gclk));
	jdff dff_B_pBDQt7Fm1_0(.din(w_dff_B_dQ2XVzZb1_0),.dout(w_dff_B_pBDQt7Fm1_0),.clk(gclk));
	jdff dff_A_hYRC2GmT0_1(.dout(w_n1464_0[1]),.din(w_dff_A_hYRC2GmT0_1),.clk(gclk));
	jdff dff_A_ETdLGiEY0_1(.dout(w_dff_A_hYRC2GmT0_1),.din(w_dff_A_ETdLGiEY0_1),.clk(gclk));
	jdff dff_A_csLbnYY68_1(.dout(w_dff_A_ETdLGiEY0_1),.din(w_dff_A_csLbnYY68_1),.clk(gclk));
	jdff dff_A_KbhxKYfc1_1(.dout(w_dff_A_csLbnYY68_1),.din(w_dff_A_KbhxKYfc1_1),.clk(gclk));
	jdff dff_A_KIdcbo8U6_1(.dout(w_dff_A_KbhxKYfc1_1),.din(w_dff_A_KIdcbo8U6_1),.clk(gclk));
	jdff dff_A_cIAROaMX8_1(.dout(w_dff_A_KIdcbo8U6_1),.din(w_dff_A_cIAROaMX8_1),.clk(gclk));
	jdff dff_A_ykPomkwX5_1(.dout(w_dff_A_cIAROaMX8_1),.din(w_dff_A_ykPomkwX5_1),.clk(gclk));
	jdff dff_B_wrLotaPu8_2(.din(n1464),.dout(w_dff_B_wrLotaPu8_2),.clk(gclk));
	jdff dff_B_qlpbRo6X8_2(.din(w_dff_B_wrLotaPu8_2),.dout(w_dff_B_qlpbRo6X8_2),.clk(gclk));
	jdff dff_B_OslxSPui1_2(.din(w_dff_B_qlpbRo6X8_2),.dout(w_dff_B_OslxSPui1_2),.clk(gclk));
	jdff dff_B_LMZAH95D2_2(.din(w_dff_B_OslxSPui1_2),.dout(w_dff_B_LMZAH95D2_2),.clk(gclk));
	jdff dff_B_W7sI2l7y4_2(.din(w_dff_B_LMZAH95D2_2),.dout(w_dff_B_W7sI2l7y4_2),.clk(gclk));
	jdff dff_B_jY4d4e6v0_2(.din(w_dff_B_W7sI2l7y4_2),.dout(w_dff_B_jY4d4e6v0_2),.clk(gclk));
	jdff dff_B_xfjsJTi02_2(.din(w_dff_B_jY4d4e6v0_2),.dout(w_dff_B_xfjsJTi02_2),.clk(gclk));
	jdff dff_B_MZyPwBM32_2(.din(w_dff_B_xfjsJTi02_2),.dout(w_dff_B_MZyPwBM32_2),.clk(gclk));
	jdff dff_B_XHc56SKP0_2(.din(w_dff_B_MZyPwBM32_2),.dout(w_dff_B_XHc56SKP0_2),.clk(gclk));
	jdff dff_B_ixzvRv4d5_2(.din(w_dff_B_XHc56SKP0_2),.dout(w_dff_B_ixzvRv4d5_2),.clk(gclk));
	jdff dff_B_Ue1tB1dW8_2(.din(w_dff_B_ixzvRv4d5_2),.dout(w_dff_B_Ue1tB1dW8_2),.clk(gclk));
	jdff dff_B_2rNbrDSn7_2(.din(w_dff_B_Ue1tB1dW8_2),.dout(w_dff_B_2rNbrDSn7_2),.clk(gclk));
	jdff dff_B_HuXvoX1q7_0(.din(n1391),.dout(w_dff_B_HuXvoX1q7_0),.clk(gclk));
	jdff dff_B_wIXhcqSn5_0(.din(w_dff_B_HuXvoX1q7_0),.dout(w_dff_B_wIXhcqSn5_0),.clk(gclk));
	jdff dff_B_AnSrUlyW8_0(.din(w_dff_B_wIXhcqSn5_0),.dout(w_dff_B_AnSrUlyW8_0),.clk(gclk));
	jdff dff_B_oUAMA5Bw9_0(.din(w_dff_B_AnSrUlyW8_0),.dout(w_dff_B_oUAMA5Bw9_0),.clk(gclk));
	jdff dff_B_blBRfFA76_0(.din(w_dff_B_oUAMA5Bw9_0),.dout(w_dff_B_blBRfFA76_0),.clk(gclk));
	jdff dff_B_RVNBsr5A7_0(.din(w_dff_B_blBRfFA76_0),.dout(w_dff_B_RVNBsr5A7_0),.clk(gclk));
	jdff dff_B_Feo5D2xO0_0(.din(w_dff_B_RVNBsr5A7_0),.dout(w_dff_B_Feo5D2xO0_0),.clk(gclk));
	jdff dff_B_vdXXe8U12_0(.din(w_dff_B_Feo5D2xO0_0),.dout(w_dff_B_vdXXe8U12_0),.clk(gclk));
	jdff dff_B_mecUcKPL7_0(.din(n1388),.dout(w_dff_B_mecUcKPL7_0),.clk(gclk));
	jdff dff_B_6JClkLPU5_0(.din(w_dff_B_mecUcKPL7_0),.dout(w_dff_B_6JClkLPU5_0),.clk(gclk));
	jdff dff_B_iot4Zr9i4_0(.din(w_dff_B_6JClkLPU5_0),.dout(w_dff_B_iot4Zr9i4_0),.clk(gclk));
	jdff dff_B_o9eZOgmS1_0(.din(w_dff_B_iot4Zr9i4_0),.dout(w_dff_B_o9eZOgmS1_0),.clk(gclk));
	jdff dff_B_GIOaFgy69_3(.din(n713),.dout(w_dff_B_GIOaFgy69_3),.clk(gclk));
	jdff dff_B_AthcAGN26_3(.din(w_dff_B_GIOaFgy69_3),.dout(w_dff_B_AthcAGN26_3),.clk(gclk));
	jdff dff_B_02lejIxl3_3(.din(w_dff_B_AthcAGN26_3),.dout(w_dff_B_02lejIxl3_3),.clk(gclk));
	jdff dff_B_Xp3YSTii9_3(.din(w_dff_B_02lejIxl3_3),.dout(w_dff_B_Xp3YSTii9_3),.clk(gclk));
	jdff dff_B_WHQ1Ggsp6_3(.din(w_dff_B_Xp3YSTii9_3),.dout(w_dff_B_WHQ1Ggsp6_3),.clk(gclk));
	jdff dff_B_CsnQHbpm0_3(.din(w_dff_B_WHQ1Ggsp6_3),.dout(w_dff_B_CsnQHbpm0_3),.clk(gclk));
	jdff dff_B_lLWNjJ9j3_3(.din(w_dff_B_CsnQHbpm0_3),.dout(w_dff_B_lLWNjJ9j3_3),.clk(gclk));
	jdff dff_B_y3fjucnV8_3(.din(w_dff_B_lLWNjJ9j3_3),.dout(w_dff_B_y3fjucnV8_3),.clk(gclk));
	jdff dff_B_qJra4Pqc5_3(.din(w_dff_B_y3fjucnV8_3),.dout(w_dff_B_qJra4Pqc5_3),.clk(gclk));
	jdff dff_B_l1SLN5z83_3(.din(w_dff_B_qJra4Pqc5_3),.dout(w_dff_B_l1SLN5z83_3),.clk(gclk));
	jdff dff_B_vBcehRgJ4_3(.din(w_dff_B_l1SLN5z83_3),.dout(w_dff_B_vBcehRgJ4_3),.clk(gclk));
	jdff dff_B_syuzaC8i3_3(.din(w_dff_B_vBcehRgJ4_3),.dout(w_dff_B_syuzaC8i3_3),.clk(gclk));
	jdff dff_B_xWHdXOLP2_3(.din(w_dff_B_syuzaC8i3_3),.dout(w_dff_B_xWHdXOLP2_3),.clk(gclk));
	jdff dff_B_fQZma7k94_3(.din(w_dff_B_xWHdXOLP2_3),.dout(w_dff_B_fQZma7k94_3),.clk(gclk));
	jdff dff_B_nKlIzAtF4_3(.din(w_dff_B_fQZma7k94_3),.dout(w_dff_B_nKlIzAtF4_3),.clk(gclk));
	jdff dff_B_fiaUomy91_3(.din(w_dff_B_nKlIzAtF4_3),.dout(w_dff_B_fiaUomy91_3),.clk(gclk));
	jdff dff_B_1rzDFzsj1_3(.din(w_dff_B_fiaUomy91_3),.dout(w_dff_B_1rzDFzsj1_3),.clk(gclk));
	jdff dff_B_wcNfDzhL9_3(.din(w_dff_B_1rzDFzsj1_3),.dout(w_dff_B_wcNfDzhL9_3),.clk(gclk));
	jdff dff_B_FivChyJd2_3(.din(w_dff_B_wcNfDzhL9_3),.dout(w_dff_B_FivChyJd2_3),.clk(gclk));
	jdff dff_A_2pLA6sGi2_0(.dout(w_n712_0[0]),.din(w_dff_A_2pLA6sGi2_0),.clk(gclk));
	jdff dff_A_IScrSnDp4_0(.dout(w_dff_A_2pLA6sGi2_0),.din(w_dff_A_IScrSnDp4_0),.clk(gclk));
	jdff dff_A_RIj09X6r4_0(.dout(w_dff_A_IScrSnDp4_0),.din(w_dff_A_RIj09X6r4_0),.clk(gclk));
	jdff dff_A_5miIlYs52_0(.dout(w_dff_A_RIj09X6r4_0),.din(w_dff_A_5miIlYs52_0),.clk(gclk));
	jdff dff_A_8S2mVXtp5_0(.dout(w_dff_A_5miIlYs52_0),.din(w_dff_A_8S2mVXtp5_0),.clk(gclk));
	jdff dff_A_bVnIap0S4_0(.dout(w_dff_A_8S2mVXtp5_0),.din(w_dff_A_bVnIap0S4_0),.clk(gclk));
	jdff dff_A_RUIAskX05_0(.dout(w_dff_A_bVnIap0S4_0),.din(w_dff_A_RUIAskX05_0),.clk(gclk));
	jdff dff_A_bqr44H7R8_0(.dout(w_dff_A_RUIAskX05_0),.din(w_dff_A_bqr44H7R8_0),.clk(gclk));
	jdff dff_A_s2bnclLQ6_0(.dout(w_dff_A_bqr44H7R8_0),.din(w_dff_A_s2bnclLQ6_0),.clk(gclk));
	jdff dff_A_NKs9K9fI5_0(.dout(w_dff_A_s2bnclLQ6_0),.din(w_dff_A_NKs9K9fI5_0),.clk(gclk));
	jdff dff_A_rVwvjIRN8_0(.dout(w_dff_A_NKs9K9fI5_0),.din(w_dff_A_rVwvjIRN8_0),.clk(gclk));
	jdff dff_A_TEOTdLan2_0(.dout(w_dff_A_rVwvjIRN8_0),.din(w_dff_A_TEOTdLan2_0),.clk(gclk));
	jdff dff_A_4pEt9iRe8_0(.dout(w_dff_A_TEOTdLan2_0),.din(w_dff_A_4pEt9iRe8_0),.clk(gclk));
	jdff dff_A_2fsMJv6Z9_0(.dout(w_dff_A_4pEt9iRe8_0),.din(w_dff_A_2fsMJv6Z9_0),.clk(gclk));
	jdff dff_A_rYs4GucR6_1(.dout(w_n708_0[1]),.din(w_dff_A_rYs4GucR6_1),.clk(gclk));
	jdff dff_A_DSUFAiTB4_1(.dout(w_dff_A_rYs4GucR6_1),.din(w_dff_A_DSUFAiTB4_1),.clk(gclk));
	jdff dff_A_AAIVqFnq0_1(.dout(w_dff_A_DSUFAiTB4_1),.din(w_dff_A_AAIVqFnq0_1),.clk(gclk));
	jdff dff_A_aKdzrLD49_1(.dout(w_dff_A_AAIVqFnq0_1),.din(w_dff_A_aKdzrLD49_1),.clk(gclk));
	jdff dff_A_93P75Fw56_1(.dout(w_dff_A_aKdzrLD49_1),.din(w_dff_A_93P75Fw56_1),.clk(gclk));
	jdff dff_A_63JeO8yX5_1(.dout(w_n707_0[1]),.din(w_dff_A_63JeO8yX5_1),.clk(gclk));
	jdff dff_A_RToS7jYS6_1(.dout(w_dff_A_63JeO8yX5_1),.din(w_dff_A_RToS7jYS6_1),.clk(gclk));
	jdff dff_A_0N8FCyks1_1(.dout(w_dff_A_RToS7jYS6_1),.din(w_dff_A_0N8FCyks1_1),.clk(gclk));
	jdff dff_A_6EiRPQPw6_1(.dout(w_dff_A_0N8FCyks1_1),.din(w_dff_A_6EiRPQPw6_1),.clk(gclk));
	jdff dff_A_DUwVtVMp5_1(.dout(w_dff_A_6EiRPQPw6_1),.din(w_dff_A_DUwVtVMp5_1),.clk(gclk));
	jdff dff_B_5GJbIelO2_1(.din(n684),.dout(w_dff_B_5GJbIelO2_1),.clk(gclk));
	jdff dff_B_6QqI81sW6_1(.din(w_dff_B_5GJbIelO2_1),.dout(w_dff_B_6QqI81sW6_1),.clk(gclk));
	jdff dff_B_31axOZ779_1(.din(w_dff_B_6QqI81sW6_1),.dout(w_dff_B_31axOZ779_1),.clk(gclk));
	jdff dff_B_WcgBQG6L5_1(.din(w_dff_B_31axOZ779_1),.dout(w_dff_B_WcgBQG6L5_1),.clk(gclk));
	jdff dff_B_AW24cn5E4_1(.din(w_dff_B_WcgBQG6L5_1),.dout(w_dff_B_AW24cn5E4_1),.clk(gclk));
	jdff dff_B_98DFixQV3_1(.din(w_dff_B_AW24cn5E4_1),.dout(w_dff_B_98DFixQV3_1),.clk(gclk));
	jdff dff_B_6CyJdoem4_1(.din(w_dff_B_98DFixQV3_1),.dout(w_dff_B_6CyJdoem4_1),.clk(gclk));
	jdff dff_B_j5sFEgj30_1(.din(w_dff_B_6CyJdoem4_1),.dout(w_dff_B_j5sFEgj30_1),.clk(gclk));
	jdff dff_B_nBGwLroT7_1(.din(w_dff_B_j5sFEgj30_1),.dout(w_dff_B_nBGwLroT7_1),.clk(gclk));
	jdff dff_B_dBcfTNrF6_1(.din(w_dff_B_nBGwLroT7_1),.dout(w_dff_B_dBcfTNrF6_1),.clk(gclk));
	jdff dff_B_QSBeyMPl2_1(.din(n685),.dout(w_dff_B_QSBeyMPl2_1),.clk(gclk));
	jdff dff_B_31TRHZrU5_1(.din(w_dff_B_QSBeyMPl2_1),.dout(w_dff_B_31TRHZrU5_1),.clk(gclk));
	jdff dff_B_j117HOou5_1(.din(w_dff_B_31TRHZrU5_1),.dout(w_dff_B_j117HOou5_1),.clk(gclk));
	jdff dff_B_nAACLr1z2_1(.din(w_dff_B_j117HOou5_1),.dout(w_dff_B_nAACLr1z2_1),.clk(gclk));
	jdff dff_B_DQ1EHF7V3_1(.din(w_dff_B_nAACLr1z2_1),.dout(w_dff_B_DQ1EHF7V3_1),.clk(gclk));
	jdff dff_B_xJnr10EK2_1(.din(w_dff_B_DQ1EHF7V3_1),.dout(w_dff_B_xJnr10EK2_1),.clk(gclk));
	jdff dff_B_qnY7mpwh9_1(.din(w_dff_B_xJnr10EK2_1),.dout(w_dff_B_qnY7mpwh9_1),.clk(gclk));
	jdff dff_B_CrkyE9VK5_1(.din(w_dff_B_qnY7mpwh9_1),.dout(w_dff_B_CrkyE9VK5_1),.clk(gclk));
	jdff dff_B_R8R1GegZ9_1(.din(w_dff_B_CrkyE9VK5_1),.dout(w_dff_B_R8R1GegZ9_1),.clk(gclk));
	jdff dff_A_b3NQQGGA8_0(.dout(w_n704_0[0]),.din(w_dff_A_b3NQQGGA8_0),.clk(gclk));
	jdff dff_A_QP6gin3t0_0(.dout(w_dff_A_b3NQQGGA8_0),.din(w_dff_A_QP6gin3t0_0),.clk(gclk));
	jdff dff_A_Cy4gb3jU5_0(.dout(w_dff_A_QP6gin3t0_0),.din(w_dff_A_Cy4gb3jU5_0),.clk(gclk));
	jdff dff_A_XtNZ2cwT4_0(.dout(w_dff_A_Cy4gb3jU5_0),.din(w_dff_A_XtNZ2cwT4_0),.clk(gclk));
	jdff dff_A_uztjHBXS0_0(.dout(w_dff_A_XtNZ2cwT4_0),.din(w_dff_A_uztjHBXS0_0),.clk(gclk));
	jdff dff_A_AFbJ8nJ87_0(.dout(w_dff_A_uztjHBXS0_0),.din(w_dff_A_AFbJ8nJ87_0),.clk(gclk));
	jdff dff_A_F2FgUrfK6_0(.dout(w_dff_A_AFbJ8nJ87_0),.din(w_dff_A_F2FgUrfK6_0),.clk(gclk));
	jdff dff_A_0ehuDGa37_0(.dout(w_dff_A_F2FgUrfK6_0),.din(w_dff_A_0ehuDGa37_0),.clk(gclk));
	jdff dff_A_geo1gBGY6_0(.dout(w_dff_A_0ehuDGa37_0),.din(w_dff_A_geo1gBGY6_0),.clk(gclk));
	jdff dff_A_QVllah6X5_0(.dout(w_dff_A_geo1gBGY6_0),.din(w_dff_A_QVllah6X5_0),.clk(gclk));
	jdff dff_A_W7cqJDbd8_0(.dout(w_dff_A_QVllah6X5_0),.din(w_dff_A_W7cqJDbd8_0),.clk(gclk));
	jdff dff_B_mMspoOhi8_1(.din(n688),.dout(w_dff_B_mMspoOhi8_1),.clk(gclk));
	jdff dff_B_SbXtGPCx1_1(.din(w_dff_B_mMspoOhi8_1),.dout(w_dff_B_SbXtGPCx1_1),.clk(gclk));
	jdff dff_B_3RZrnDtC6_1(.din(w_dff_B_SbXtGPCx1_1),.dout(w_dff_B_3RZrnDtC6_1),.clk(gclk));
	jdff dff_B_k26eojcT9_1(.din(w_dff_B_3RZrnDtC6_1),.dout(w_dff_B_k26eojcT9_1),.clk(gclk));
	jdff dff_B_eirtcAzx3_1(.din(w_dff_B_k26eojcT9_1),.dout(w_dff_B_eirtcAzx3_1),.clk(gclk));
	jdff dff_B_USI1XqZs9_1(.din(n689),.dout(w_dff_B_USI1XqZs9_1),.clk(gclk));
	jdff dff_B_lbDXiSBl2_1(.din(w_dff_B_USI1XqZs9_1),.dout(w_dff_B_lbDXiSBl2_1),.clk(gclk));
	jdff dff_B_c7vP74jz2_1(.din(w_dff_B_lbDXiSBl2_1),.dout(w_dff_B_c7vP74jz2_1),.clk(gclk));
	jdff dff_B_fuS5g3We1_1(.din(w_dff_B_c7vP74jz2_1),.dout(w_dff_B_fuS5g3We1_1),.clk(gclk));
	jdff dff_B_ZrU08K1A0_0(.din(n698),.dout(w_dff_B_ZrU08K1A0_0),.clk(gclk));
	jdff dff_A_pDvDnkNp0_0(.dout(w_n697_0[0]),.din(w_dff_A_pDvDnkNp0_0),.clk(gclk));
	jdff dff_A_VHmyh0658_0(.dout(w_dff_A_pDvDnkNp0_0),.din(w_dff_A_VHmyh0658_0),.clk(gclk));
	jdff dff_A_llREnJMm9_0(.dout(w_dff_A_VHmyh0658_0),.din(w_dff_A_llREnJMm9_0),.clk(gclk));
	jdff dff_A_5plgl53j5_0(.dout(w_dff_A_llREnJMm9_0),.din(w_dff_A_5plgl53j5_0),.clk(gclk));
	jdff dff_A_FUNQwxCo7_0(.dout(w_dff_A_5plgl53j5_0),.din(w_dff_A_FUNQwxCo7_0),.clk(gclk));
	jdff dff_A_rFRXfMHw8_0(.dout(w_dff_A_FUNQwxCo7_0),.din(w_dff_A_rFRXfMHw8_0),.clk(gclk));
	jdff dff_A_Heppkal78_0(.dout(w_dff_A_rFRXfMHw8_0),.din(w_dff_A_Heppkal78_0),.clk(gclk));
	jdff dff_A_S98k5jCQ7_0(.dout(w_dff_A_Heppkal78_0),.din(w_dff_A_S98k5jCQ7_0),.clk(gclk));
	jdff dff_A_yGyzPe4B2_0(.dout(w_dff_A_S98k5jCQ7_0),.din(w_dff_A_yGyzPe4B2_0),.clk(gclk));
	jdff dff_A_7FMjB3Vu6_0(.dout(w_dff_A_yGyzPe4B2_0),.din(w_dff_A_7FMjB3Vu6_0),.clk(gclk));
	jdff dff_A_63wWsD236_0(.dout(w_dff_A_7FMjB3Vu6_0),.din(w_dff_A_63wWsD236_0),.clk(gclk));
	jdff dff_A_VnPbcDzP7_0(.dout(w_dff_A_63wWsD236_0),.din(w_dff_A_VnPbcDzP7_0),.clk(gclk));
	jdff dff_A_u7F2Q8m55_1(.dout(w_n697_0[1]),.din(w_dff_A_u7F2Q8m55_1),.clk(gclk));
	jdff dff_A_OXz8K64H4_1(.dout(w_dff_A_u7F2Q8m55_1),.din(w_dff_A_OXz8K64H4_1),.clk(gclk));
	jdff dff_A_h6WxvGi87_1(.dout(w_dff_A_OXz8K64H4_1),.din(w_dff_A_h6WxvGi87_1),.clk(gclk));
	jdff dff_A_N1hFQIAX4_1(.dout(w_dff_A_h6WxvGi87_1),.din(w_dff_A_N1hFQIAX4_1),.clk(gclk));
	jdff dff_A_kqHA7SEI9_1(.dout(w_dff_A_N1hFQIAX4_1),.din(w_dff_A_kqHA7SEI9_1),.clk(gclk));
	jdff dff_A_OHcH1tg02_1(.dout(w_dff_A_kqHA7SEI9_1),.din(w_dff_A_OHcH1tg02_1),.clk(gclk));
	jdff dff_A_pIWS2X621_1(.dout(w_dff_A_OHcH1tg02_1),.din(w_dff_A_pIWS2X621_1),.clk(gclk));
	jdff dff_A_Cy9aYAbq4_1(.dout(w_dff_A_pIWS2X621_1),.din(w_dff_A_Cy9aYAbq4_1),.clk(gclk));
	jdff dff_A_fSmbRiGw6_1(.dout(w_dff_A_Cy9aYAbq4_1),.din(w_dff_A_fSmbRiGw6_1),.clk(gclk));
	jdff dff_A_ntRiys6G6_1(.dout(w_dff_A_fSmbRiGw6_1),.din(w_dff_A_ntRiys6G6_1),.clk(gclk));
	jdff dff_A_GtSFQ6Iu6_1(.dout(w_dff_A_ntRiys6G6_1),.din(w_dff_A_GtSFQ6Iu6_1),.clk(gclk));
	jdff dff_A_NxWtbGzu4_1(.dout(w_dff_A_GtSFQ6Iu6_1),.din(w_dff_A_NxWtbGzu4_1),.clk(gclk));
	jdff dff_A_h48hVY0p1_1(.dout(w_dff_A_NxWtbGzu4_1),.din(w_dff_A_h48hVY0p1_1),.clk(gclk));
	jdff dff_A_39wYxN6T5_1(.dout(w_dff_A_h48hVY0p1_1),.din(w_dff_A_39wYxN6T5_1),.clk(gclk));
	jdff dff_A_ywic1fHk4_1(.dout(w_dff_A_39wYxN6T5_1),.din(w_dff_A_ywic1fHk4_1),.clk(gclk));
	jdff dff_A_ohcuHZ8E6_1(.dout(w_dff_A_ywic1fHk4_1),.din(w_dff_A_ohcuHZ8E6_1),.clk(gclk));
	jdff dff_A_T8J0NI7b7_1(.dout(w_dff_A_ohcuHZ8E6_1),.din(w_dff_A_T8J0NI7b7_1),.clk(gclk));
	jdff dff_A_N0r6384D1_1(.dout(w_n692_0[1]),.din(w_dff_A_N0r6384D1_1),.clk(gclk));
	jdff dff_A_1IQtyevN2_1(.dout(w_n687_0[1]),.din(w_dff_A_1IQtyevN2_1),.clk(gclk));
	jdff dff_B_3CWIUYUh5_2(.din(n687),.dout(w_dff_B_3CWIUYUh5_2),.clk(gclk));
	jdff dff_B_ZSb2eyue1_2(.din(w_dff_B_3CWIUYUh5_2),.dout(w_dff_B_ZSb2eyue1_2),.clk(gclk));
	jdff dff_B_UEr6zIbv1_2(.din(w_dff_B_ZSb2eyue1_2),.dout(w_dff_B_UEr6zIbv1_2),.clk(gclk));
	jdff dff_B_JqLPROAF1_2(.din(w_dff_B_UEr6zIbv1_2),.dout(w_dff_B_JqLPROAF1_2),.clk(gclk));
	jdff dff_B_FRjIx0s29_2(.din(w_dff_B_JqLPROAF1_2),.dout(w_dff_B_FRjIx0s29_2),.clk(gclk));
	jdff dff_A_0uQLXxFj7_0(.dout(w_n686_0[0]),.din(w_dff_A_0uQLXxFj7_0),.clk(gclk));
	jdff dff_A_se3lgJdO6_0(.dout(w_dff_A_0uQLXxFj7_0),.din(w_dff_A_se3lgJdO6_0),.clk(gclk));
	jdff dff_A_tw1W2qY31_0(.dout(w_dff_A_se3lgJdO6_0),.din(w_dff_A_tw1W2qY31_0),.clk(gclk));
	jdff dff_A_HijjC0fh7_0(.dout(w_dff_A_tw1W2qY31_0),.din(w_dff_A_HijjC0fh7_0),.clk(gclk));
	jdff dff_A_OzFdgeut2_0(.dout(w_dff_A_HijjC0fh7_0),.din(w_dff_A_OzFdgeut2_0),.clk(gclk));
	jdff dff_B_a6vI01Xa7_0(.din(n682),.dout(w_dff_B_a6vI01Xa7_0),.clk(gclk));
	jdff dff_B_PbVZSAaj7_0(.din(w_dff_B_a6vI01Xa7_0),.dout(w_dff_B_PbVZSAaj7_0),.clk(gclk));
	jdff dff_B_zoGqrCsr9_0(.din(w_dff_B_PbVZSAaj7_0),.dout(w_dff_B_zoGqrCsr9_0),.clk(gclk));
	jdff dff_B_8TrRRcVy0_0(.din(w_dff_B_zoGqrCsr9_0),.dout(w_dff_B_8TrRRcVy0_0),.clk(gclk));
	jdff dff_B_UD8zV4Fo8_0(.din(w_dff_B_8TrRRcVy0_0),.dout(w_dff_B_UD8zV4Fo8_0),.clk(gclk));
	jdff dff_B_3vhR5FRd5_0(.din(w_dff_B_UD8zV4Fo8_0),.dout(w_dff_B_3vhR5FRd5_0),.clk(gclk));
	jdff dff_B_egxG1bLp0_0(.din(w_dff_B_3vhR5FRd5_0),.dout(w_dff_B_egxG1bLp0_0),.clk(gclk));
	jdff dff_B_wzsIbGOs3_0(.din(w_dff_B_egxG1bLp0_0),.dout(w_dff_B_wzsIbGOs3_0),.clk(gclk));
	jdff dff_B_M597tXan2_0(.din(w_dff_B_wzsIbGOs3_0),.dout(w_dff_B_M597tXan2_0),.clk(gclk));
	jdff dff_B_oSwk6T4H0_0(.din(w_dff_B_M597tXan2_0),.dout(w_dff_B_oSwk6T4H0_0),.clk(gclk));
	jdff dff_B_lbYoKhjc4_0(.din(w_dff_B_oSwk6T4H0_0),.dout(w_dff_B_lbYoKhjc4_0),.clk(gclk));
	jdff dff_B_v6k1PaaS2_0(.din(w_dff_B_lbYoKhjc4_0),.dout(w_dff_B_v6k1PaaS2_0),.clk(gclk));
	jdff dff_A_nRk0F1yu3_0(.dout(w_n680_0[0]),.din(w_dff_A_nRk0F1yu3_0),.clk(gclk));
	jdff dff_A_9F0lqJYL3_0(.dout(w_dff_A_nRk0F1yu3_0),.din(w_dff_A_9F0lqJYL3_0),.clk(gclk));
	jdff dff_A_ahdHbyKk0_0(.dout(w_dff_A_9F0lqJYL3_0),.din(w_dff_A_ahdHbyKk0_0),.clk(gclk));
	jdff dff_A_BsN9hC1e8_0(.dout(w_dff_A_ahdHbyKk0_0),.din(w_dff_A_BsN9hC1e8_0),.clk(gclk));
	jdff dff_A_bmHVwHPA3_0(.dout(w_dff_A_BsN9hC1e8_0),.din(w_dff_A_bmHVwHPA3_0),.clk(gclk));
	jdff dff_A_8v14q7Rr6_1(.dout(w_n679_0[1]),.din(w_dff_A_8v14q7Rr6_1),.clk(gclk));
	jdff dff_A_bxt3cWg04_1(.dout(w_dff_A_8v14q7Rr6_1),.din(w_dff_A_bxt3cWg04_1),.clk(gclk));
	jdff dff_A_ROvKrg5y1_2(.dout(w_n679_0[2]),.din(w_dff_A_ROvKrg5y1_2),.clk(gclk));
	jdff dff_A_IUaQs51h2_0(.dout(w_n678_0[0]),.din(w_dff_A_IUaQs51h2_0),.clk(gclk));
	jdff dff_A_RQV5umD88_0(.dout(w_dff_A_IUaQs51h2_0),.din(w_dff_A_RQV5umD88_0),.clk(gclk));
	jdff dff_A_DZvNQCFr8_0(.dout(w_dff_A_RQV5umD88_0),.din(w_dff_A_DZvNQCFr8_0),.clk(gclk));
	jdff dff_A_Efe0r4uT8_0(.dout(w_dff_A_DZvNQCFr8_0),.din(w_dff_A_Efe0r4uT8_0),.clk(gclk));
	jdff dff_A_BOeQg6d50_0(.dout(w_dff_A_Efe0r4uT8_0),.din(w_dff_A_BOeQg6d50_0),.clk(gclk));
	jdff dff_A_mcxyT3IL0_0(.dout(w_dff_A_BOeQg6d50_0),.din(w_dff_A_mcxyT3IL0_0),.clk(gclk));
	jdff dff_A_83idBDcV2_0(.dout(w_dff_A_mcxyT3IL0_0),.din(w_dff_A_83idBDcV2_0),.clk(gclk));
	jdff dff_A_1SOOwDKX2_0(.dout(w_dff_A_83idBDcV2_0),.din(w_dff_A_1SOOwDKX2_0),.clk(gclk));
	jdff dff_A_GfgfAQdm0_0(.dout(w_dff_A_1SOOwDKX2_0),.din(w_dff_A_GfgfAQdm0_0),.clk(gclk));
	jdff dff_A_qN9E9QMu1_0(.dout(w_dff_A_GfgfAQdm0_0),.din(w_dff_A_qN9E9QMu1_0),.clk(gclk));
	jdff dff_A_SZwoJk737_0(.dout(w_dff_A_qN9E9QMu1_0),.din(w_dff_A_SZwoJk737_0),.clk(gclk));
	jdff dff_A_FoAN2lGm2_0(.dout(w_dff_A_SZwoJk737_0),.din(w_dff_A_FoAN2lGm2_0),.clk(gclk));
	jdff dff_A_U9khHxe71_0(.dout(w_dff_A_FoAN2lGm2_0),.din(w_dff_A_U9khHxe71_0),.clk(gclk));
	jdff dff_A_LOgY3SDJ6_0(.dout(w_dff_A_U9khHxe71_0),.din(w_dff_A_LOgY3SDJ6_0),.clk(gclk));
	jdff dff_A_24HZQlwX4_0(.dout(w_dff_A_LOgY3SDJ6_0),.din(w_dff_A_24HZQlwX4_0),.clk(gclk));
	jdff dff_A_Hk3heCbt6_0(.dout(w_dff_A_24HZQlwX4_0),.din(w_dff_A_Hk3heCbt6_0),.clk(gclk));
	jdff dff_A_dy8idU0p2_1(.dout(w_n678_0[1]),.din(w_dff_A_dy8idU0p2_1),.clk(gclk));
	jdff dff_A_0k3ywTYN8_1(.dout(w_dff_A_dy8idU0p2_1),.din(w_dff_A_0k3ywTYN8_1),.clk(gclk));
	jdff dff_A_FfUNx92S1_1(.dout(w_dff_A_0k3ywTYN8_1),.din(w_dff_A_FfUNx92S1_1),.clk(gclk));
	jdff dff_A_xeqNNqnp7_1(.dout(w_dff_A_FfUNx92S1_1),.din(w_dff_A_xeqNNqnp7_1),.clk(gclk));
	jdff dff_A_uhzyLWyT7_1(.dout(w_dff_A_xeqNNqnp7_1),.din(w_dff_A_uhzyLWyT7_1),.clk(gclk));
	jdff dff_A_yI1dmKmU2_1(.dout(w_dff_A_uhzyLWyT7_1),.din(w_dff_A_yI1dmKmU2_1),.clk(gclk));
	jdff dff_A_7ed9KzhY5_1(.dout(w_dff_A_yI1dmKmU2_1),.din(w_dff_A_7ed9KzhY5_1),.clk(gclk));
	jdff dff_A_g9dXKNb59_1(.dout(w_dff_A_7ed9KzhY5_1),.din(w_dff_A_g9dXKNb59_1),.clk(gclk));
	jdff dff_A_fivInbil4_1(.dout(w_dff_A_g9dXKNb59_1),.din(w_dff_A_fivInbil4_1),.clk(gclk));
	jdff dff_A_TuC4Q1IY3_1(.dout(w_dff_A_fivInbil4_1),.din(w_dff_A_TuC4Q1IY3_1),.clk(gclk));
	jdff dff_A_zHTplkiB0_1(.dout(w_dff_A_TuC4Q1IY3_1),.din(w_dff_A_zHTplkiB0_1),.clk(gclk));
	jdff dff_A_HCOkP9kF2_1(.dout(w_dff_A_zHTplkiB0_1),.din(w_dff_A_HCOkP9kF2_1),.clk(gclk));
	jdff dff_A_pFcKP18F0_1(.dout(w_dff_A_HCOkP9kF2_1),.din(w_dff_A_pFcKP18F0_1),.clk(gclk));
	jdff dff_A_aQekNMNG6_1(.dout(w_dff_A_pFcKP18F0_1),.din(w_dff_A_aQekNMNG6_1),.clk(gclk));
	jdff dff_A_BrggSZaM2_1(.dout(w_dff_A_aQekNMNG6_1),.din(w_dff_A_BrggSZaM2_1),.clk(gclk));
	jdff dff_A_ksJ7tGhk9_1(.dout(w_dff_A_BrggSZaM2_1),.din(w_dff_A_ksJ7tGhk9_1),.clk(gclk));
	jdff dff_B_ntO3dZxz6_0(.din(G209),.dout(w_dff_B_ntO3dZxz6_0),.clk(gclk));
	jdff dff_B_Eb137lpD7_3(.din(n675),.dout(w_dff_B_Eb137lpD7_3),.clk(gclk));
	jdff dff_B_1b42s4Cf3_3(.din(w_dff_B_Eb137lpD7_3),.dout(w_dff_B_1b42s4Cf3_3),.clk(gclk));
	jdff dff_A_FXzQTZBz9_0(.dout(w_n674_1[0]),.din(w_dff_A_FXzQTZBz9_0),.clk(gclk));
	jdff dff_A_W3wYQSli9_0(.dout(w_dff_A_FXzQTZBz9_0),.din(w_dff_A_W3wYQSli9_0),.clk(gclk));
	jdff dff_A_JXQWSPKi0_0(.dout(w_dff_A_W3wYQSli9_0),.din(w_dff_A_JXQWSPKi0_0),.clk(gclk));
	jdff dff_A_Vtxl6EgM4_0(.dout(w_dff_A_JXQWSPKi0_0),.din(w_dff_A_Vtxl6EgM4_0),.clk(gclk));
	jdff dff_A_IS4t9m6n0_0(.dout(w_dff_A_Vtxl6EgM4_0),.din(w_dff_A_IS4t9m6n0_0),.clk(gclk));
	jdff dff_A_qnmJzlNA5_0(.dout(w_dff_A_IS4t9m6n0_0),.din(w_dff_A_qnmJzlNA5_0),.clk(gclk));
	jdff dff_A_traQn1J99_0(.dout(w_dff_A_qnmJzlNA5_0),.din(w_dff_A_traQn1J99_0),.clk(gclk));
	jdff dff_A_0KY4L7qb6_0(.dout(w_dff_A_traQn1J99_0),.din(w_dff_A_0KY4L7qb6_0),.clk(gclk));
	jdff dff_A_cLN2eEGx0_0(.dout(w_dff_A_0KY4L7qb6_0),.din(w_dff_A_cLN2eEGx0_0),.clk(gclk));
	jdff dff_A_J3qQsUsv8_0(.dout(w_dff_A_cLN2eEGx0_0),.din(w_dff_A_J3qQsUsv8_0),.clk(gclk));
	jdff dff_A_hpwijWbA4_0(.dout(w_dff_A_J3qQsUsv8_0),.din(w_dff_A_hpwijWbA4_0),.clk(gclk));
	jdff dff_A_w8FTFYUL0_0(.dout(w_dff_A_hpwijWbA4_0),.din(w_dff_A_w8FTFYUL0_0),.clk(gclk));
	jdff dff_A_6Hl9xR1E1_0(.dout(w_dff_A_w8FTFYUL0_0),.din(w_dff_A_6Hl9xR1E1_0),.clk(gclk));
	jdff dff_A_jPop937a0_0(.dout(w_dff_A_6Hl9xR1E1_0),.din(w_dff_A_jPop937a0_0),.clk(gclk));
	jdff dff_A_csVXd10E6_0(.dout(w_dff_A_jPop937a0_0),.din(w_dff_A_csVXd10E6_0),.clk(gclk));
	jdff dff_A_m1C0VH770_0(.dout(w_dff_A_csVXd10E6_0),.din(w_dff_A_m1C0VH770_0),.clk(gclk));
	jdff dff_A_CIVjT5VM8_0(.dout(w_dff_A_m1C0VH770_0),.din(w_dff_A_CIVjT5VM8_0),.clk(gclk));
	jdff dff_A_v7RfquDs0_0(.dout(w_dff_A_CIVjT5VM8_0),.din(w_dff_A_v7RfquDs0_0),.clk(gclk));
	jdff dff_A_QUy4eyxe1_1(.dout(w_n674_0[1]),.din(w_dff_A_QUy4eyxe1_1),.clk(gclk));
	jdff dff_A_phBDlMg71_1(.dout(w_dff_A_QUy4eyxe1_1),.din(w_dff_A_phBDlMg71_1),.clk(gclk));
	jdff dff_A_fIC2p0Xx1_1(.dout(w_dff_A_phBDlMg71_1),.din(w_dff_A_fIC2p0Xx1_1),.clk(gclk));
	jdff dff_A_uCNOdBRd7_1(.dout(w_dff_A_fIC2p0Xx1_1),.din(w_dff_A_uCNOdBRd7_1),.clk(gclk));
	jdff dff_A_A0vxmUpU9_1(.dout(w_dff_A_uCNOdBRd7_1),.din(w_dff_A_A0vxmUpU9_1),.clk(gclk));
	jdff dff_A_TxJfzI5u1_1(.dout(w_dff_A_A0vxmUpU9_1),.din(w_dff_A_TxJfzI5u1_1),.clk(gclk));
	jdff dff_A_9Q4iBcA39_1(.dout(w_dff_A_TxJfzI5u1_1),.din(w_dff_A_9Q4iBcA39_1),.clk(gclk));
	jdff dff_A_OKZphSOh1_1(.dout(w_dff_A_9Q4iBcA39_1),.din(w_dff_A_OKZphSOh1_1),.clk(gclk));
	jdff dff_A_pVVPqvYX2_1(.dout(w_dff_A_OKZphSOh1_1),.din(w_dff_A_pVVPqvYX2_1),.clk(gclk));
	jdff dff_A_QZfrvL4I7_1(.dout(w_dff_A_pVVPqvYX2_1),.din(w_dff_A_QZfrvL4I7_1),.clk(gclk));
	jdff dff_A_8O7LrDql9_1(.dout(w_dff_A_QZfrvL4I7_1),.din(w_dff_A_8O7LrDql9_1),.clk(gclk));
	jdff dff_A_FhDUAYYh0_1(.dout(w_dff_A_8O7LrDql9_1),.din(w_dff_A_FhDUAYYh0_1),.clk(gclk));
	jdff dff_A_mzieiADk9_1(.dout(w_dff_A_FhDUAYYh0_1),.din(w_dff_A_mzieiADk9_1),.clk(gclk));
	jdff dff_A_ohXg0I1s7_0(.dout(w_n672_0[0]),.din(w_dff_A_ohXg0I1s7_0),.clk(gclk));
	jdff dff_A_1aqJqf1o2_0(.dout(w_dff_A_ohXg0I1s7_0),.din(w_dff_A_1aqJqf1o2_0),.clk(gclk));
	jdff dff_B_k0FUDk4O7_0(.din(G216),.dout(w_dff_B_k0FUDk4O7_0),.clk(gclk));
	jdff dff_B_UFEOpjR45_2(.din(n671),.dout(w_dff_B_UFEOpjR45_2),.clk(gclk));
	jdff dff_B_xfvM5hH19_2(.din(w_dff_B_UFEOpjR45_2),.dout(w_dff_B_xfvM5hH19_2),.clk(gclk));
	jdff dff_A_D4pDAyua3_0(.dout(w_G1469_1[0]),.din(w_dff_A_D4pDAyua3_0),.clk(gclk));
	jdff dff_A_dA0aAkgi9_0(.dout(w_dff_A_D4pDAyua3_0),.din(w_dff_A_dA0aAkgi9_0),.clk(gclk));
	jdff dff_A_66mRX9688_0(.dout(w_dff_A_dA0aAkgi9_0),.din(w_dff_A_66mRX9688_0),.clk(gclk));
	jdff dff_A_6HCsU9672_0(.dout(w_dff_A_66mRX9688_0),.din(w_dff_A_6HCsU9672_0),.clk(gclk));
	jdff dff_A_iVqUbNYz1_0(.dout(w_n667_0[0]),.din(w_dff_A_iVqUbNYz1_0),.clk(gclk));
	jdff dff_A_Rt6Qggwj7_0(.dout(w_dff_A_iVqUbNYz1_0),.din(w_dff_A_Rt6Qggwj7_0),.clk(gclk));
	jdff dff_B_XHcYUwEC3_0(.din(G215),.dout(w_dff_B_XHcYUwEC3_0),.clk(gclk));
	jdff dff_B_ZdNvDYb41_2(.din(n666),.dout(w_dff_B_ZdNvDYb41_2),.clk(gclk));
	jdff dff_B_xceFMOFW7_2(.din(w_dff_B_ZdNvDYb41_2),.dout(w_dff_B_xceFMOFW7_2),.clk(gclk));
	jdff dff_A_IuovkDfs4_0(.dout(w_G106_1[0]),.din(w_dff_A_IuovkDfs4_0),.clk(gclk));
	jdff dff_A_A3N2WasT5_0(.dout(w_dff_A_IuovkDfs4_0),.din(w_dff_A_A3N2WasT5_0),.clk(gclk));
	jdff dff_A_v0z01ZgM1_0(.dout(w_dff_A_A3N2WasT5_0),.din(w_dff_A_v0z01ZgM1_0),.clk(gclk));
	jdff dff_A_pPlrvx5T9_0(.dout(w_dff_A_v0z01ZgM1_0),.din(w_dff_A_pPlrvx5T9_0),.clk(gclk));
	jdff dff_B_n7oZ3W448_0(.din(G214),.dout(w_dff_B_n7oZ3W448_0),.clk(gclk));
	jdff dff_B_rNlhbg6w2_3(.din(n662),.dout(w_dff_B_rNlhbg6w2_3),.clk(gclk));
	jdff dff_B_pmxFTMoD6_3(.din(w_dff_B_rNlhbg6w2_3),.dout(w_dff_B_pmxFTMoD6_3),.clk(gclk));
	jdff dff_A_N0kDuRwy6_1(.dout(w_n661_0[1]),.din(w_dff_A_N0kDuRwy6_1),.clk(gclk));
	jdff dff_A_Ivn3BrT31_1(.dout(w_dff_A_N0kDuRwy6_1),.din(w_dff_A_Ivn3BrT31_1),.clk(gclk));
	jdff dff_B_tR2LbQ4n4_0(.din(G213),.dout(w_dff_B_tR2LbQ4n4_0),.clk(gclk));
	jdff dff_B_z6Iml3TC6_3(.din(n658),.dout(w_dff_B_z6Iml3TC6_3),.clk(gclk));
	jdff dff_B_VXaHy9Hx2_3(.din(w_dff_B_z6Iml3TC6_3),.dout(w_dff_B_VXaHy9Hx2_3),.clk(gclk));
	jdff dff_A_LhYOVxyI5_1(.dout(w_n656_0[1]),.din(w_dff_A_LhYOVxyI5_1),.clk(gclk));
	jdff dff_A_Ug3mK5NG0_1(.dout(w_dff_A_LhYOVxyI5_1),.din(w_dff_A_Ug3mK5NG0_1),.clk(gclk));
	jdff dff_A_7wd10qIo0_1(.dout(w_dff_A_Ug3mK5NG0_1),.din(w_dff_A_7wd10qIo0_1),.clk(gclk));
	jdff dff_A_EAb3kC1d5_1(.dout(w_dff_A_7wd10qIo0_1),.din(w_dff_A_EAb3kC1d5_1),.clk(gclk));
	jdff dff_A_MAQeO5oo4_1(.dout(w_dff_A_EAb3kC1d5_1),.din(w_dff_A_MAQeO5oo4_1),.clk(gclk));
	jdff dff_A_B6LaQCym1_1(.dout(w_dff_A_MAQeO5oo4_1),.din(w_dff_A_B6LaQCym1_1),.clk(gclk));
	jdff dff_A_mRWBJonj2_1(.dout(w_dff_A_B6LaQCym1_1),.din(w_dff_A_mRWBJonj2_1),.clk(gclk));
	jdff dff_A_15KflhwZ3_1(.dout(w_dff_A_mRWBJonj2_1),.din(w_dff_A_15KflhwZ3_1),.clk(gclk));
	jdff dff_A_HSuaGMv20_1(.dout(w_dff_A_15KflhwZ3_1),.din(w_dff_A_HSuaGMv20_1),.clk(gclk));
	jdff dff_B_fVfsT3JD2_1(.din(n641),.dout(w_dff_B_fVfsT3JD2_1),.clk(gclk));
	jdff dff_B_Mkxo0zjz7_1(.din(w_dff_B_fVfsT3JD2_1),.dout(w_dff_B_Mkxo0zjz7_1),.clk(gclk));
	jdff dff_B_Z7mHQ0hz1_1(.din(w_dff_B_Mkxo0zjz7_1),.dout(w_dff_B_Z7mHQ0hz1_1),.clk(gclk));
	jdff dff_B_M9KreNBI5_1(.din(w_dff_B_Z7mHQ0hz1_1),.dout(w_dff_B_M9KreNBI5_1),.clk(gclk));
	jdff dff_B_hAhFDvod4_0(.din(n654),.dout(w_dff_B_hAhFDvod4_0),.clk(gclk));
	jdff dff_B_QRx72X1R3_0(.din(w_dff_B_hAhFDvod4_0),.dout(w_dff_B_QRx72X1R3_0),.clk(gclk));
	jdff dff_A_nx74sppU0_0(.dout(w_n653_1[0]),.din(w_dff_A_nx74sppU0_0),.clk(gclk));
	jdff dff_A_pLdcDt4v1_0(.dout(w_dff_A_nx74sppU0_0),.din(w_dff_A_pLdcDt4v1_0),.clk(gclk));
	jdff dff_A_UmgNyxXY9_0(.dout(w_dff_A_pLdcDt4v1_0),.din(w_dff_A_UmgNyxXY9_0),.clk(gclk));
	jdff dff_A_whLRc9xJ3_0(.dout(w_dff_A_UmgNyxXY9_0),.din(w_dff_A_whLRc9xJ3_0),.clk(gclk));
	jdff dff_A_mdlHZwOP4_0(.dout(w_dff_A_whLRc9xJ3_0),.din(w_dff_A_mdlHZwOP4_0),.clk(gclk));
	jdff dff_A_1lprh0ls4_0(.dout(w_dff_A_mdlHZwOP4_0),.din(w_dff_A_1lprh0ls4_0),.clk(gclk));
	jdff dff_A_afMyLor28_0(.dout(w_dff_A_1lprh0ls4_0),.din(w_dff_A_afMyLor28_0),.clk(gclk));
	jdff dff_A_vQHn923G0_0(.dout(w_dff_A_afMyLor28_0),.din(w_dff_A_vQHn923G0_0),.clk(gclk));
	jdff dff_A_H5ozfvEf8_0(.dout(w_dff_A_vQHn923G0_0),.din(w_dff_A_H5ozfvEf8_0),.clk(gclk));
	jdff dff_A_Bn4mYZrY0_0(.dout(w_dff_A_H5ozfvEf8_0),.din(w_dff_A_Bn4mYZrY0_0),.clk(gclk));
	jdff dff_A_1fPSTm731_0(.dout(w_dff_A_Bn4mYZrY0_0),.din(w_dff_A_1fPSTm731_0),.clk(gclk));
	jdff dff_A_hPBh4mk55_0(.dout(w_dff_A_1fPSTm731_0),.din(w_dff_A_hPBh4mk55_0),.clk(gclk));
	jdff dff_A_LAnBHev18_0(.dout(w_dff_A_hPBh4mk55_0),.din(w_dff_A_LAnBHev18_0),.clk(gclk));
	jdff dff_A_N85r8T5u6_0(.dout(w_dff_A_LAnBHev18_0),.din(w_dff_A_N85r8T5u6_0),.clk(gclk));
	jdff dff_A_bYH1Yk4w1_0(.dout(w_dff_A_N85r8T5u6_0),.din(w_dff_A_bYH1Yk4w1_0),.clk(gclk));
	jdff dff_A_piWLtxRU3_1(.dout(w_n653_0[1]),.din(w_dff_A_piWLtxRU3_1),.clk(gclk));
	jdff dff_A_wne7cskn8_1(.dout(w_dff_A_piWLtxRU3_1),.din(w_dff_A_wne7cskn8_1),.clk(gclk));
	jdff dff_A_sUtFUMxE0_1(.dout(w_dff_A_wne7cskn8_1),.din(w_dff_A_sUtFUMxE0_1),.clk(gclk));
	jdff dff_A_mni2gDwA4_1(.dout(w_n648_0[1]),.din(w_dff_A_mni2gDwA4_1),.clk(gclk));
	jdff dff_A_9qscZx968_1(.dout(w_dff_A_mni2gDwA4_1),.din(w_dff_A_9qscZx968_1),.clk(gclk));
	jdff dff_A_DOr04mro5_1(.dout(w_dff_A_9qscZx968_1),.din(w_dff_A_DOr04mro5_1),.clk(gclk));
	jdff dff_A_VTSm0hsC0_1(.dout(w_dff_A_DOr04mro5_1),.din(w_dff_A_VTSm0hsC0_1),.clk(gclk));
	jdff dff_A_ZCxDpFtE6_1(.dout(w_dff_A_VTSm0hsC0_1),.din(w_dff_A_ZCxDpFtE6_1),.clk(gclk));
	jdff dff_A_ucRnVag98_1(.dout(w_dff_A_ZCxDpFtE6_1),.din(w_dff_A_ucRnVag98_1),.clk(gclk));
	jdff dff_A_0EK1odHV0_1(.dout(w_dff_A_ucRnVag98_1),.din(w_dff_A_0EK1odHV0_1),.clk(gclk));
	jdff dff_A_PMyYqndW8_1(.dout(w_dff_A_0EK1odHV0_1),.din(w_dff_A_PMyYqndW8_1),.clk(gclk));
	jdff dff_A_DB7tKIUf7_1(.dout(w_dff_A_PMyYqndW8_1),.din(w_dff_A_DB7tKIUf7_1),.clk(gclk));
	jdff dff_A_YR6YSlRF7_1(.dout(w_dff_A_DB7tKIUf7_1),.din(w_dff_A_YR6YSlRF7_1),.clk(gclk));
	jdff dff_A_IpbrTOhL4_1(.dout(w_dff_A_YR6YSlRF7_1),.din(w_dff_A_IpbrTOhL4_1),.clk(gclk));
	jdff dff_A_LnBaAuQd1_1(.dout(w_dff_A_IpbrTOhL4_1),.din(w_dff_A_LnBaAuQd1_1),.clk(gclk));
	jdff dff_B_C4tzDZ6m2_1(.din(n644),.dout(w_dff_B_C4tzDZ6m2_1),.clk(gclk));
	jdff dff_A_NlXmhPtA6_0(.dout(w_n645_0[0]),.din(w_dff_A_NlXmhPtA6_0),.clk(gclk));
	jdff dff_A_qb3jlVHQ1_1(.dout(w_n645_0[1]),.din(w_dff_A_qb3jlVHQ1_1),.clk(gclk));
	jdff dff_A_imvC1xlh9_1(.dout(w_dff_A_qb3jlVHQ1_1),.din(w_dff_A_imvC1xlh9_1),.clk(gclk));
	jdff dff_A_SlLxopcg6_1(.dout(w_dff_A_imvC1xlh9_1),.din(w_dff_A_SlLxopcg6_1),.clk(gclk));
	jdff dff_A_SntQfvgC6_1(.dout(w_dff_A_SlLxopcg6_1),.din(w_dff_A_SntQfvgC6_1),.clk(gclk));
	jdff dff_A_rORgkK0L6_1(.dout(w_dff_A_SntQfvgC6_1),.din(w_dff_A_rORgkK0L6_1),.clk(gclk));
	jdff dff_A_i8Ge2UoJ1_1(.dout(w_dff_A_rORgkK0L6_1),.din(w_dff_A_i8Ge2UoJ1_1),.clk(gclk));
	jdff dff_A_xTDhwCkA7_1(.dout(w_dff_A_i8Ge2UoJ1_1),.din(w_dff_A_xTDhwCkA7_1),.clk(gclk));
	jdff dff_A_u1XntUmo6_1(.dout(w_dff_A_xTDhwCkA7_1),.din(w_dff_A_u1XntUmo6_1),.clk(gclk));
	jdff dff_A_A3w1LbOh4_1(.dout(w_dff_A_u1XntUmo6_1),.din(w_dff_A_A3w1LbOh4_1),.clk(gclk));
	jdff dff_A_hAcYqbdW5_1(.dout(w_dff_A_A3w1LbOh4_1),.din(w_dff_A_hAcYqbdW5_1),.clk(gclk));
	jdff dff_A_URvGaDG78_1(.dout(w_dff_A_hAcYqbdW5_1),.din(w_dff_A_URvGaDG78_1),.clk(gclk));
	jdff dff_A_o77milgf7_1(.dout(w_dff_A_URvGaDG78_1),.din(w_dff_A_o77milgf7_1),.clk(gclk));
	jdff dff_A_UkMHL19G4_1(.dout(w_dff_A_o77milgf7_1),.din(w_dff_A_UkMHL19G4_1),.clk(gclk));
	jdff dff_A_TYce3fmA5_1(.dout(w_dff_A_UkMHL19G4_1),.din(w_dff_A_TYce3fmA5_1),.clk(gclk));
	jdff dff_A_xKhpYeJo3_1(.dout(w_dff_A_TYce3fmA5_1),.din(w_dff_A_xKhpYeJo3_1),.clk(gclk));
	jdff dff_A_TF2dRplP6_0(.dout(w_n643_0[0]),.din(w_dff_A_TF2dRplP6_0),.clk(gclk));
	jdff dff_A_NSQ0FXRP2_0(.dout(w_dff_A_TF2dRplP6_0),.din(w_dff_A_NSQ0FXRP2_0),.clk(gclk));
	jdff dff_A_xjREGCon4_0(.dout(w_dff_A_NSQ0FXRP2_0),.din(w_dff_A_xjREGCon4_0),.clk(gclk));
	jdff dff_A_gTFgY2Nd6_0(.dout(w_dff_A_xjREGCon4_0),.din(w_dff_A_gTFgY2Nd6_0),.clk(gclk));
	jdff dff_A_YdIucaZ67_0(.dout(w_dff_A_gTFgY2Nd6_0),.din(w_dff_A_YdIucaZ67_0),.clk(gclk));
	jdff dff_A_WVB6Expa2_0(.dout(w_dff_A_YdIucaZ67_0),.din(w_dff_A_WVB6Expa2_0),.clk(gclk));
	jdff dff_A_b9qFrL5p4_0(.dout(w_dff_A_WVB6Expa2_0),.din(w_dff_A_b9qFrL5p4_0),.clk(gclk));
	jdff dff_A_kZNUPEa16_0(.dout(w_dff_A_b9qFrL5p4_0),.din(w_dff_A_kZNUPEa16_0),.clk(gclk));
	jdff dff_A_UzbzHfDK9_0(.dout(w_dff_A_kZNUPEa16_0),.din(w_dff_A_UzbzHfDK9_0),.clk(gclk));
	jdff dff_A_bO5DoJI41_0(.dout(w_dff_A_UzbzHfDK9_0),.din(w_dff_A_bO5DoJI41_0),.clk(gclk));
	jdff dff_A_BhdhF3A34_0(.dout(w_dff_A_bO5DoJI41_0),.din(w_dff_A_BhdhF3A34_0),.clk(gclk));
	jdff dff_A_H378nXVf0_0(.dout(w_dff_A_BhdhF3A34_0),.din(w_dff_A_H378nXVf0_0),.clk(gclk));
	jdff dff_A_xApNFDDi8_0(.dout(w_dff_A_H378nXVf0_0),.din(w_dff_A_xApNFDDi8_0),.clk(gclk));
	jdff dff_A_htWSNZ0U3_0(.dout(w_dff_A_xApNFDDi8_0),.din(w_dff_A_htWSNZ0U3_0),.clk(gclk));
	jdff dff_B_8bzvD6Xj6_2(.din(n643),.dout(w_dff_B_8bzvD6Xj6_2),.clk(gclk));
	jdff dff_B_64BnYiHV3_2(.din(w_dff_B_8bzvD6Xj6_2),.dout(w_dff_B_64BnYiHV3_2),.clk(gclk));
	jdff dff_A_kTkwB2Kb6_0(.dout(w_n642_0[0]),.din(w_dff_A_kTkwB2Kb6_0),.clk(gclk));
	jdff dff_A_g5E6Xoil8_0(.dout(w_dff_A_kTkwB2Kb6_0),.din(w_dff_A_g5E6Xoil8_0),.clk(gclk));
	jdff dff_A_PxZd0RBT7_0(.dout(w_dff_A_g5E6Xoil8_0),.din(w_dff_A_PxZd0RBT7_0),.clk(gclk));
	jdff dff_A_e1l956lS8_0(.dout(w_dff_A_PxZd0RBT7_0),.din(w_dff_A_e1l956lS8_0),.clk(gclk));
	jdff dff_A_8nXhsAqp5_0(.dout(w_dff_A_e1l956lS8_0),.din(w_dff_A_8nXhsAqp5_0),.clk(gclk));
	jdff dff_B_ePSTFwxn2_0(.din(n638),.dout(w_dff_B_ePSTFwxn2_0),.clk(gclk));
	jdff dff_B_dZZlInJA2_0(.din(w_dff_B_ePSTFwxn2_0),.dout(w_dff_B_dZZlInJA2_0),.clk(gclk));
	jdff dff_B_5FdAPyX25_0(.din(w_dff_B_dZZlInJA2_0),.dout(w_dff_B_5FdAPyX25_0),.clk(gclk));
	jdff dff_B_yE7AFs3X2_0(.din(w_dff_B_5FdAPyX25_0),.dout(w_dff_B_yE7AFs3X2_0),.clk(gclk));
	jdff dff_B_P4AxfDd10_0(.din(w_dff_B_yE7AFs3X2_0),.dout(w_dff_B_P4AxfDd10_0),.clk(gclk));
	jdff dff_B_2dTI95Ag6_0(.din(w_dff_B_P4AxfDd10_0),.dout(w_dff_B_2dTI95Ag6_0),.clk(gclk));
	jdff dff_B_GJhZjZyj5_0(.din(w_dff_B_2dTI95Ag6_0),.dout(w_dff_B_GJhZjZyj5_0),.clk(gclk));
	jdff dff_B_GF1bxYkC6_0(.din(w_dff_B_GJhZjZyj5_0),.dout(w_dff_B_GF1bxYkC6_0),.clk(gclk));
	jdff dff_B_cDhyUstl7_0(.din(w_dff_B_GF1bxYkC6_0),.dout(w_dff_B_cDhyUstl7_0),.clk(gclk));
	jdff dff_B_hyaXkRZh4_0(.din(w_dff_B_cDhyUstl7_0),.dout(w_dff_B_hyaXkRZh4_0),.clk(gclk));
	jdff dff_B_5bVHzCoB6_0(.din(w_dff_B_hyaXkRZh4_0),.dout(w_dff_B_5bVHzCoB6_0),.clk(gclk));
	jdff dff_A_dI8kEoUQ0_0(.dout(w_n637_0[0]),.din(w_dff_A_dI8kEoUQ0_0),.clk(gclk));
	jdff dff_A_v283yLyc2_0(.dout(w_dff_A_dI8kEoUQ0_0),.din(w_dff_A_v283yLyc2_0),.clk(gclk));
	jdff dff_A_9CzZbaMW0_0(.dout(w_dff_A_v283yLyc2_0),.din(w_dff_A_9CzZbaMW0_0),.clk(gclk));
	jdff dff_A_PTXyHzPb2_0(.dout(w_dff_A_9CzZbaMW0_0),.din(w_dff_A_PTXyHzPb2_0),.clk(gclk));
	jdff dff_A_7yrQxVyh3_0(.dout(w_dff_A_PTXyHzPb2_0),.din(w_dff_A_7yrQxVyh3_0),.clk(gclk));
	jdff dff_A_hXgRrwjt0_0(.dout(w_dff_A_7yrQxVyh3_0),.din(w_dff_A_hXgRrwjt0_0),.clk(gclk));
	jdff dff_A_mQ7JHL7A0_0(.dout(w_dff_A_hXgRrwjt0_0),.din(w_dff_A_mQ7JHL7A0_0),.clk(gclk));
	jdff dff_A_jJWjSZLk1_0(.dout(w_dff_A_mQ7JHL7A0_0),.din(w_dff_A_jJWjSZLk1_0),.clk(gclk));
	jdff dff_A_tGKiAFJ45_0(.dout(w_dff_A_jJWjSZLk1_0),.din(w_dff_A_tGKiAFJ45_0),.clk(gclk));
	jdff dff_A_OAwK0ZCv7_0(.dout(w_dff_A_tGKiAFJ45_0),.din(w_dff_A_OAwK0ZCv7_0),.clk(gclk));
	jdff dff_A_GJ4scgZd6_0(.dout(w_dff_A_OAwK0ZCv7_0),.din(w_dff_A_GJ4scgZd6_0),.clk(gclk));
	jdff dff_A_YBLe62Qq7_0(.dout(w_dff_A_GJ4scgZd6_0),.din(w_dff_A_YBLe62Qq7_0),.clk(gclk));
	jdff dff_A_U3iOSSB60_0(.dout(w_n635_0[0]),.din(w_dff_A_U3iOSSB60_0),.clk(gclk));
	jdff dff_A_BhhxFeUR3_0(.dout(w_n633_0[0]),.din(w_dff_A_BhhxFeUR3_0),.clk(gclk));
	jdff dff_A_z6Z7PJLr0_0(.dout(w_dff_A_BhhxFeUR3_0),.din(w_dff_A_z6Z7PJLr0_0),.clk(gclk));
	jdff dff_B_gmR2tVV00_0(.din(G154),.dout(w_dff_B_gmR2tVV00_0),.clk(gclk));
	jdff dff_B_Wun7VePb7_2(.din(n632),.dout(w_dff_B_Wun7VePb7_2),.clk(gclk));
	jdff dff_B_TLKxVHrz8_2(.din(w_dff_B_Wun7VePb7_2),.dout(w_dff_B_TLKxVHrz8_2),.clk(gclk));
	jdff dff_A_5KOVEoVw7_0(.dout(w_G2253_1[0]),.din(w_dff_A_5KOVEoVw7_0),.clk(gclk));
	jdff dff_A_ZMWNQO8U4_0(.dout(w_dff_A_5KOVEoVw7_0),.din(w_dff_A_ZMWNQO8U4_0),.clk(gclk));
	jdff dff_A_MwA18U3m5_0(.dout(w_dff_A_ZMWNQO8U4_0),.din(w_dff_A_MwA18U3m5_0),.clk(gclk));
	jdff dff_A_9uuk3uJU2_0(.dout(w_dff_A_MwA18U3m5_0),.din(w_dff_A_9uuk3uJU2_0),.clk(gclk));
	jdff dff_A_PlpkORAv3_0(.dout(w_n629_0[0]),.din(w_dff_A_PlpkORAv3_0),.clk(gclk));
	jdff dff_A_EX3ZzQQk9_0(.dout(w_dff_A_PlpkORAv3_0),.din(w_dff_A_EX3ZzQQk9_0),.clk(gclk));
	jdff dff_B_9U7qMuqH0_0(.din(G153),.dout(w_dff_B_9U7qMuqH0_0),.clk(gclk));
	jdff dff_B_wkLN8WmT3_2(.din(n628),.dout(w_dff_B_wkLN8WmT3_2),.clk(gclk));
	jdff dff_B_KqGlf3EU9_2(.din(w_dff_B_wkLN8WmT3_2),.dout(w_dff_B_KqGlf3EU9_2),.clk(gclk));
	jdff dff_A_H4W4do6z0_0(.dout(w_G2256_1[0]),.din(w_dff_A_H4W4do6z0_0),.clk(gclk));
	jdff dff_A_oif6KGoZ0_0(.dout(w_dff_A_H4W4do6z0_0),.din(w_dff_A_oif6KGoZ0_0),.clk(gclk));
	jdff dff_A_8cHYjrwL0_0(.dout(w_dff_A_oif6KGoZ0_0),.din(w_dff_A_8cHYjrwL0_0),.clk(gclk));
	jdff dff_A_Of6m4djP1_0(.dout(w_dff_A_8cHYjrwL0_0),.din(w_dff_A_Of6m4djP1_0),.clk(gclk));
	jdff dff_A_s8YrdGsc3_0(.dout(w_n626_0[0]),.din(w_dff_A_s8YrdGsc3_0),.clk(gclk));
	jdff dff_A_RnCEZq7s6_0(.dout(w_dff_A_s8YrdGsc3_0),.din(w_dff_A_RnCEZq7s6_0),.clk(gclk));
	jdff dff_A_tjQ9oybE9_0(.dout(w_dff_A_RnCEZq7s6_0),.din(w_dff_A_tjQ9oybE9_0),.clk(gclk));
	jdff dff_A_CWdmyTBg6_0(.dout(w_dff_A_tjQ9oybE9_0),.din(w_dff_A_CWdmyTBg6_0),.clk(gclk));
	jdff dff_A_xgzkMFPV2_0(.dout(w_dff_A_CWdmyTBg6_0),.din(w_dff_A_xgzkMFPV2_0),.clk(gclk));
	jdff dff_A_n6EGCexi3_0(.dout(w_dff_A_xgzkMFPV2_0),.din(w_dff_A_n6EGCexi3_0),.clk(gclk));
	jdff dff_A_Lyuesbap7_0(.dout(w_dff_A_n6EGCexi3_0),.din(w_dff_A_Lyuesbap7_0),.clk(gclk));
	jdff dff_A_UaKZasdC2_0(.dout(w_dff_A_Lyuesbap7_0),.din(w_dff_A_UaKZasdC2_0),.clk(gclk));
	jdff dff_A_xVfsRKwD1_0(.dout(w_dff_A_UaKZasdC2_0),.din(w_dff_A_xVfsRKwD1_0),.clk(gclk));
	jdff dff_A_I12FHI8l0_0(.dout(w_dff_A_xVfsRKwD1_0),.din(w_dff_A_I12FHI8l0_0),.clk(gclk));
	jdff dff_A_NRpGR77t6_0(.dout(w_dff_A_I12FHI8l0_0),.din(w_dff_A_NRpGR77t6_0),.clk(gclk));
	jdff dff_A_kOdyl9j68_0(.dout(w_dff_A_NRpGR77t6_0),.din(w_dff_A_kOdyl9j68_0),.clk(gclk));
	jdff dff_A_YcCrtlXV4_0(.dout(w_dff_A_kOdyl9j68_0),.din(w_dff_A_YcCrtlXV4_0),.clk(gclk));
	jdff dff_A_DqfIZIe95_0(.dout(w_dff_A_YcCrtlXV4_0),.din(w_dff_A_DqfIZIe95_0),.clk(gclk));
	jdff dff_A_OnR7F0Ov0_0(.dout(w_n624_0[0]),.din(w_dff_A_OnR7F0Ov0_0),.clk(gclk));
	jdff dff_A_xUWqSw9H1_0(.dout(w_dff_A_OnR7F0Ov0_0),.din(w_dff_A_xUWqSw9H1_0),.clk(gclk));
	jdff dff_B_q90zLv3b6_0(.din(G156),.dout(w_dff_B_q90zLv3b6_0),.clk(gclk));
	jdff dff_A_8IlHPIpi6_1(.dout(w_n623_0[1]),.din(w_dff_A_8IlHPIpi6_1),.clk(gclk));
	jdff dff_A_hhuo9bPa3_1(.dout(w_dff_A_8IlHPIpi6_1),.din(w_dff_A_hhuo9bPa3_1),.clk(gclk));
	jdff dff_A_jOYC5UJN4_2(.dout(w_n623_0[2]),.din(w_dff_A_jOYC5UJN4_2),.clk(gclk));
	jdff dff_A_82enB9Zl4_2(.dout(w_dff_A_jOYC5UJN4_2),.din(w_dff_A_82enB9Zl4_2),.clk(gclk));
	jdff dff_A_K6kRUXt23_1(.dout(w_G2239_0[1]),.din(w_dff_A_K6kRUXt23_1),.clk(gclk));
	jdff dff_A_lzE1Hsi35_1(.dout(w_dff_A_K6kRUXt23_1),.din(w_dff_A_lzE1Hsi35_1),.clk(gclk));
	jdff dff_A_L8NjtLMm4_1(.dout(w_dff_A_lzE1Hsi35_1),.din(w_dff_A_L8NjtLMm4_1),.clk(gclk));
	jdff dff_A_mBJGbxOA3_1(.dout(w_dff_A_L8NjtLMm4_1),.din(w_dff_A_mBJGbxOA3_1),.clk(gclk));
	jdff dff_A_Jx6Nmo0H4_2(.dout(w_n622_0[2]),.din(w_dff_A_Jx6Nmo0H4_2),.clk(gclk));
	jdff dff_A_Inpx9wdH7_2(.dout(w_dff_A_Jx6Nmo0H4_2),.din(w_dff_A_Inpx9wdH7_2),.clk(gclk));
	jdff dff_A_1sTzqk7F1_2(.dout(w_dff_A_Inpx9wdH7_2),.din(w_dff_A_1sTzqk7F1_2),.clk(gclk));
	jdff dff_A_n9sFzddv8_2(.dout(w_dff_A_1sTzqk7F1_2),.din(w_dff_A_n9sFzddv8_2),.clk(gclk));
	jdff dff_A_5hBpT9Dg3_2(.dout(w_dff_A_n9sFzddv8_2),.din(w_dff_A_5hBpT9Dg3_2),.clk(gclk));
	jdff dff_A_H9zOAFHx9_2(.dout(w_dff_A_5hBpT9Dg3_2),.din(w_dff_A_H9zOAFHx9_2),.clk(gclk));
	jdff dff_A_DepeEy322_2(.dout(w_dff_A_H9zOAFHx9_2),.din(w_dff_A_DepeEy322_2),.clk(gclk));
	jdff dff_A_xiHKryJN7_2(.dout(w_dff_A_DepeEy322_2),.din(w_dff_A_xiHKryJN7_2),.clk(gclk));
	jdff dff_A_zCrUtDH90_2(.dout(w_dff_A_xiHKryJN7_2),.din(w_dff_A_zCrUtDH90_2),.clk(gclk));
	jdff dff_A_eN39hUaF2_2(.dout(w_dff_A_zCrUtDH90_2),.din(w_dff_A_eN39hUaF2_2),.clk(gclk));
	jdff dff_A_pLg4OBT42_2(.dout(w_dff_A_eN39hUaF2_2),.din(w_dff_A_pLg4OBT42_2),.clk(gclk));
	jdff dff_A_66N60CTd1_2(.dout(w_dff_A_pLg4OBT42_2),.din(w_dff_A_66N60CTd1_2),.clk(gclk));
	jdff dff_A_famUi9Ow7_2(.dout(w_dff_A_66N60CTd1_2),.din(w_dff_A_famUi9Ow7_2),.clk(gclk));
	jdff dff_A_FlQ3axMt0_2(.dout(w_dff_A_famUi9Ow7_2),.din(w_dff_A_FlQ3axMt0_2),.clk(gclk));
	jdff dff_A_w0z19Z6F8_2(.dout(w_dff_A_FlQ3axMt0_2),.din(w_dff_A_w0z19Z6F8_2),.clk(gclk));
	jdff dff_A_QOjGnQml7_2(.dout(w_dff_A_w0z19Z6F8_2),.din(w_dff_A_QOjGnQml7_2),.clk(gclk));
	jdff dff_A_j7dIH2GR1_0(.dout(w_n620_0[0]),.din(w_dff_A_j7dIH2GR1_0),.clk(gclk));
	jdff dff_A_Kir7Rrku2_0(.dout(w_dff_A_j7dIH2GR1_0),.din(w_dff_A_Kir7Rrku2_0),.clk(gclk));
	jdff dff_B_ushaR9vI3_0(.din(G155),.dout(w_dff_B_ushaR9vI3_0),.clk(gclk));
	jdff dff_B_g6uKnzF50_2(.din(n619),.dout(w_dff_B_g6uKnzF50_2),.clk(gclk));
	jdff dff_B_an6MDwmU2_2(.din(w_dff_B_g6uKnzF50_2),.dout(w_dff_B_an6MDwmU2_2),.clk(gclk));
	jdff dff_A_7hEVAEFb8_1(.dout(w_n617_0[1]),.din(w_dff_A_7hEVAEFb8_1),.clk(gclk));
	jdff dff_A_HWHE1biM3_1(.dout(w_dff_A_7hEVAEFb8_1),.din(w_dff_A_HWHE1biM3_1),.clk(gclk));
	jdff dff_A_prTVDyTp7_1(.dout(w_dff_A_HWHE1biM3_1),.din(w_dff_A_prTVDyTp7_1),.clk(gclk));
	jdff dff_A_8ufHP8OR6_1(.dout(w_dff_A_prTVDyTp7_1),.din(w_dff_A_8ufHP8OR6_1),.clk(gclk));
	jdff dff_A_6arFQ3iJ3_1(.dout(w_dff_A_8ufHP8OR6_1),.din(w_dff_A_6arFQ3iJ3_1),.clk(gclk));
	jdff dff_B_7BmYyDMm7_1(.din(n596),.dout(w_dff_B_7BmYyDMm7_1),.clk(gclk));
	jdff dff_B_SlYEXmrL8_1(.din(w_dff_B_7BmYyDMm7_1),.dout(w_dff_B_SlYEXmrL8_1),.clk(gclk));
	jdff dff_B_xlCfDRVl8_1(.din(w_dff_B_SlYEXmrL8_1),.dout(w_dff_B_xlCfDRVl8_1),.clk(gclk));
	jdff dff_B_LHWRhSg61_1(.din(w_dff_B_xlCfDRVl8_1),.dout(w_dff_B_LHWRhSg61_1),.clk(gclk));
	jdff dff_B_bOwuuzCy2_1(.din(w_dff_B_LHWRhSg61_1),.dout(w_dff_B_bOwuuzCy2_1),.clk(gclk));
	jdff dff_B_9fDOTzUJ0_1(.din(w_dff_B_bOwuuzCy2_1),.dout(w_dff_B_9fDOTzUJ0_1),.clk(gclk));
	jdff dff_B_D5Q2xOZA1_1(.din(n598),.dout(w_dff_B_D5Q2xOZA1_1),.clk(gclk));
	jdff dff_B_yME1aZo34_1(.din(w_dff_B_D5Q2xOZA1_1),.dout(w_dff_B_yME1aZo34_1),.clk(gclk));
	jdff dff_B_rpVKhQ6F6_1(.din(w_dff_B_yME1aZo34_1),.dout(w_dff_B_rpVKhQ6F6_1),.clk(gclk));
	jdff dff_B_l3n405Ep5_1(.din(w_dff_B_rpVKhQ6F6_1),.dout(w_dff_B_l3n405Ep5_1),.clk(gclk));
	jdff dff_B_IFTfh1mX6_1(.din(w_dff_B_l3n405Ep5_1),.dout(w_dff_B_IFTfh1mX6_1),.clk(gclk));
	jdff dff_A_81XBlqvm4_0(.dout(w_n615_1[0]),.din(w_dff_A_81XBlqvm4_0),.clk(gclk));
	jdff dff_A_D1phObl95_0(.dout(w_dff_A_81XBlqvm4_0),.din(w_dff_A_D1phObl95_0),.clk(gclk));
	jdff dff_A_uHmO9OH33_0(.dout(w_dff_A_D1phObl95_0),.din(w_dff_A_uHmO9OH33_0),.clk(gclk));
	jdff dff_A_h3AVsrzd6_0(.dout(w_dff_A_uHmO9OH33_0),.din(w_dff_A_h3AVsrzd6_0),.clk(gclk));
	jdff dff_A_REXG7Zhp7_0(.dout(w_dff_A_h3AVsrzd6_0),.din(w_dff_A_REXG7Zhp7_0),.clk(gclk));
	jdff dff_A_vklsPczg5_0(.dout(w_dff_A_REXG7Zhp7_0),.din(w_dff_A_vklsPczg5_0),.clk(gclk));
	jdff dff_A_4QMJZCK65_0(.dout(w_dff_A_vklsPczg5_0),.din(w_dff_A_4QMJZCK65_0),.clk(gclk));
	jdff dff_A_VsAIbkmZ9_0(.dout(w_dff_A_4QMJZCK65_0),.din(w_dff_A_VsAIbkmZ9_0),.clk(gclk));
	jdff dff_A_KrygBMp55_0(.dout(w_dff_A_VsAIbkmZ9_0),.din(w_dff_A_KrygBMp55_0),.clk(gclk));
	jdff dff_B_6pPOnS6H0_1(.din(n600),.dout(w_dff_B_6pPOnS6H0_1),.clk(gclk));
	jdff dff_B_TlsEcBTW6_1(.din(w_dff_B_6pPOnS6H0_1),.dout(w_dff_B_TlsEcBTW6_1),.clk(gclk));
	jdff dff_B_iTUWS4sz1_1(.din(w_dff_B_TlsEcBTW6_1),.dout(w_dff_B_iTUWS4sz1_1),.clk(gclk));
	jdff dff_B_bO2tCcQc4_1(.din(w_dff_B_iTUWS4sz1_1),.dout(w_dff_B_bO2tCcQc4_1),.clk(gclk));
	jdff dff_B_x1Yl5yVa8_1(.din(n602),.dout(w_dff_B_x1Yl5yVa8_1),.clk(gclk));
	jdff dff_B_wFDA0cag7_1(.din(w_dff_B_x1Yl5yVa8_1),.dout(w_dff_B_wFDA0cag7_1),.clk(gclk));
	jdff dff_B_PSNRXKgT4_1(.din(w_dff_B_wFDA0cag7_1),.dout(w_dff_B_PSNRXKgT4_1),.clk(gclk));
	jdff dff_A_wjUihQaD1_1(.dout(w_n613_0[1]),.din(w_dff_A_wjUihQaD1_1),.clk(gclk));
	jdff dff_A_x70VSDT46_1(.dout(w_dff_A_wjUihQaD1_1),.din(w_dff_A_x70VSDT46_1),.clk(gclk));
	jdff dff_A_KmiCco6I6_1(.dout(w_dff_A_x70VSDT46_1),.din(w_dff_A_KmiCco6I6_1),.clk(gclk));
	jdff dff_A_JyowotkQ5_1(.dout(w_dff_A_KmiCco6I6_1),.din(w_dff_A_JyowotkQ5_1),.clk(gclk));
	jdff dff_A_5jgCpFzy0_1(.dout(w_dff_A_JyowotkQ5_1),.din(w_dff_A_5jgCpFzy0_1),.clk(gclk));
	jdff dff_A_AmXvraAA1_1(.dout(w_dff_A_5jgCpFzy0_1),.din(w_dff_A_AmXvraAA1_1),.clk(gclk));
	jdff dff_A_8UQcol652_1(.dout(w_dff_A_AmXvraAA1_1),.din(w_dff_A_8UQcol652_1),.clk(gclk));
	jdff dff_A_WbBHUvTq9_1(.dout(w_dff_A_8UQcol652_1),.din(w_dff_A_WbBHUvTq9_1),.clk(gclk));
	jdff dff_A_9cezoIdV4_1(.dout(w_dff_A_WbBHUvTq9_1),.din(w_dff_A_9cezoIdV4_1),.clk(gclk));
	jdff dff_A_AeGQcbZC4_1(.dout(w_dff_A_9cezoIdV4_1),.din(w_dff_A_AeGQcbZC4_1),.clk(gclk));
	jdff dff_A_JOD0nreV1_0(.dout(w_n610_0[0]),.din(w_dff_A_JOD0nreV1_0),.clk(gclk));
	jdff dff_A_Nei84SfY4_0(.dout(w_dff_A_JOD0nreV1_0),.din(w_dff_A_Nei84SfY4_0),.clk(gclk));
	jdff dff_A_OyMjnSER3_0(.dout(w_n608_0[0]),.din(w_dff_A_OyMjnSER3_0),.clk(gclk));
	jdff dff_A_nv66cA3z1_0(.dout(w_dff_A_OyMjnSER3_0),.din(w_dff_A_nv66cA3z1_0),.clk(gclk));
	jdff dff_A_PGBKZuMi7_0(.dout(w_n606_1[0]),.din(w_dff_A_PGBKZuMi7_0),.clk(gclk));
	jdff dff_A_D2YnCEkM4_0(.dout(w_dff_A_PGBKZuMi7_0),.din(w_dff_A_D2YnCEkM4_0),.clk(gclk));
	jdff dff_A_FuQ2lwZi3_0(.dout(w_dff_A_D2YnCEkM4_0),.din(w_dff_A_FuQ2lwZi3_0),.clk(gclk));
	jdff dff_A_8CDfmc8z6_0(.dout(w_dff_A_FuQ2lwZi3_0),.din(w_dff_A_8CDfmc8z6_0),.clk(gclk));
	jdff dff_A_gFW2FglF0_1(.dout(w_n606_1[1]),.din(w_dff_A_gFW2FglF0_1),.clk(gclk));
	jdff dff_A_MfH5EZsL5_1(.dout(w_dff_A_gFW2FglF0_1),.din(w_dff_A_MfH5EZsL5_1),.clk(gclk));
	jdff dff_A_OgMELuPM1_1(.dout(w_dff_A_MfH5EZsL5_1),.din(w_dff_A_OgMELuPM1_1),.clk(gclk));
	jdff dff_A_lI0VZls23_1(.dout(w_dff_A_OgMELuPM1_1),.din(w_dff_A_lI0VZls23_1),.clk(gclk));
	jdff dff_A_y36RNCp36_1(.dout(w_dff_A_lI0VZls23_1),.din(w_dff_A_y36RNCp36_1),.clk(gclk));
	jdff dff_A_auSOT7Ez1_1(.dout(w_dff_A_y36RNCp36_1),.din(w_dff_A_auSOT7Ez1_1),.clk(gclk));
	jdff dff_A_07zLDTuy0_1(.dout(w_dff_A_auSOT7Ez1_1),.din(w_dff_A_07zLDTuy0_1),.clk(gclk));
	jdff dff_A_3Gaffbtx8_1(.dout(w_dff_A_07zLDTuy0_1),.din(w_dff_A_3Gaffbtx8_1),.clk(gclk));
	jdff dff_A_Legihi8a8_1(.dout(w_dff_A_3Gaffbtx8_1),.din(w_dff_A_Legihi8a8_1),.clk(gclk));
	jdff dff_A_pRiVCr5C8_1(.dout(w_dff_A_Legihi8a8_1),.din(w_dff_A_pRiVCr5C8_1),.clk(gclk));
	jdff dff_A_nQrK5SOy7_1(.dout(w_dff_A_pRiVCr5C8_1),.din(w_dff_A_nQrK5SOy7_1),.clk(gclk));
	jdff dff_A_90PfBetN6_1(.dout(w_dff_A_nQrK5SOy7_1),.din(w_dff_A_90PfBetN6_1),.clk(gclk));
	jdff dff_A_sIc5B8IA5_1(.dout(w_dff_A_90PfBetN6_1),.din(w_dff_A_sIc5B8IA5_1),.clk(gclk));
	jdff dff_A_bpIZOWyw1_0(.dout(w_n599_0[0]),.din(w_dff_A_bpIZOWyw1_0),.clk(gclk));
	jdff dff_A_gsuy1xhg7_0(.dout(w_dff_A_bpIZOWyw1_0),.din(w_dff_A_gsuy1xhg7_0),.clk(gclk));
	jdff dff_A_NVkVw5Rr0_0(.dout(w_dff_A_gsuy1xhg7_0),.din(w_dff_A_NVkVw5Rr0_0),.clk(gclk));
	jdff dff_A_9kPS5u6Z9_0(.dout(w_dff_A_NVkVw5Rr0_0),.din(w_dff_A_9kPS5u6Z9_0),.clk(gclk));
	jdff dff_A_cOrKHC8r7_0(.dout(w_dff_A_9kPS5u6Z9_0),.din(w_dff_A_cOrKHC8r7_0),.clk(gclk));
	jdff dff_B_ALmpcn5E2_0(.din(n593),.dout(w_dff_B_ALmpcn5E2_0),.clk(gclk));
	jdff dff_B_8DMOOf4i3_0(.din(w_dff_B_ALmpcn5E2_0),.dout(w_dff_B_8DMOOf4i3_0),.clk(gclk));
	jdff dff_B_m293t9WZ8_0(.din(w_dff_B_8DMOOf4i3_0),.dout(w_dff_B_m293t9WZ8_0),.clk(gclk));
	jdff dff_B_gmoTMHaR0_0(.din(w_dff_B_m293t9WZ8_0),.dout(w_dff_B_gmoTMHaR0_0),.clk(gclk));
	jdff dff_B_d5sNZA4I3_0(.din(w_dff_B_gmoTMHaR0_0),.dout(w_dff_B_d5sNZA4I3_0),.clk(gclk));
	jdff dff_B_IDfMCid82_0(.din(w_dff_B_d5sNZA4I3_0),.dout(w_dff_B_IDfMCid82_0),.clk(gclk));
	jdff dff_B_3MDwyOK57_0(.din(w_dff_B_IDfMCid82_0),.dout(w_dff_B_3MDwyOK57_0),.clk(gclk));
	jdff dff_B_fuApnOfa2_0(.din(w_dff_B_3MDwyOK57_0),.dout(w_dff_B_fuApnOfa2_0),.clk(gclk));
	jdff dff_A_zcwsYSNy8_0(.dout(w_n592_0[0]),.din(w_dff_A_zcwsYSNy8_0),.clk(gclk));
	jdff dff_A_lLbhIJXG0_0(.dout(w_dff_A_zcwsYSNy8_0),.din(w_dff_A_lLbhIJXG0_0),.clk(gclk));
	jdff dff_A_pM3KtXqT8_0(.dout(w_dff_A_lLbhIJXG0_0),.din(w_dff_A_pM3KtXqT8_0),.clk(gclk));
	jdff dff_A_ps7QqfkW5_0(.dout(w_dff_A_pM3KtXqT8_0),.din(w_dff_A_ps7QqfkW5_0),.clk(gclk));
	jdff dff_A_z7tTAFy69_0(.dout(w_dff_A_ps7QqfkW5_0),.din(w_dff_A_z7tTAFy69_0),.clk(gclk));
	jdff dff_A_No7cUPur3_0(.dout(w_dff_A_z7tTAFy69_0),.din(w_dff_A_No7cUPur3_0),.clk(gclk));
	jdff dff_A_PTQffy812_0(.dout(w_dff_A_No7cUPur3_0),.din(w_dff_A_PTQffy812_0),.clk(gclk));
	jdff dff_A_6lDzlWRP6_0(.dout(w_dff_A_PTQffy812_0),.din(w_dff_A_6lDzlWRP6_0),.clk(gclk));
	jdff dff_A_LwVKvSsc3_0(.dout(w_dff_A_6lDzlWRP6_0),.din(w_dff_A_LwVKvSsc3_0),.clk(gclk));
	jdff dff_A_VcZ0ObV67_1(.dout(w_n589_0[1]),.din(w_dff_A_VcZ0ObV67_1),.clk(gclk));
	jdff dff_B_DeBhIout9_0(.din(n587),.dout(w_dff_B_DeBhIout9_0),.clk(gclk));
	jdff dff_B_lV3ChrZN8_0(.din(G144),.dout(w_dff_B_lV3ChrZN8_0),.clk(gclk));
	jdff dff_B_xZ08vA4y3_2(.din(n585),.dout(w_dff_B_xZ08vA4y3_2),.clk(gclk));
	jdff dff_B_WDEbrLem7_2(.din(w_dff_B_xZ08vA4y3_2),.dout(w_dff_B_WDEbrLem7_2),.clk(gclk));
	jdff dff_A_fzbjfxrA9_0(.dout(w_G2224_1[0]),.din(w_dff_A_fzbjfxrA9_0),.clk(gclk));
	jdff dff_A_479Mr7cO0_0(.dout(w_dff_A_fzbjfxrA9_0),.din(w_dff_A_479Mr7cO0_0),.clk(gclk));
	jdff dff_A_W3X3aebx9_0(.dout(w_dff_A_479Mr7cO0_0),.din(w_dff_A_W3X3aebx9_0),.clk(gclk));
	jdff dff_A_mm6HwVJP0_0(.dout(w_dff_A_W3X3aebx9_0),.din(w_dff_A_mm6HwVJP0_0),.clk(gclk));
	jdff dff_B_D5js8nOw4_0(.din(n582),.dout(w_dff_B_D5js8nOw4_0),.clk(gclk));
	jdff dff_B_1N5R0yCL3_0(.din(G135),.dout(w_dff_B_1N5R0yCL3_0),.clk(gclk));
	jdff dff_B_0K0C5rfL1_2(.din(n580),.dout(w_dff_B_0K0C5rfL1_2),.clk(gclk));
	jdff dff_B_0BNgGgMg3_2(.din(w_dff_B_0K0C5rfL1_2),.dout(w_dff_B_0BNgGgMg3_2),.clk(gclk));
	jdff dff_A_cm1WQzw24_0(.dout(w_G2230_1[0]),.din(w_dff_A_cm1WQzw24_0),.clk(gclk));
	jdff dff_A_AxAcsGCx7_0(.dout(w_dff_A_cm1WQzw24_0),.din(w_dff_A_AxAcsGCx7_0),.clk(gclk));
	jdff dff_A_UmwWKvEW7_0(.dout(w_dff_A_AxAcsGCx7_0),.din(w_dff_A_UmwWKvEW7_0),.clk(gclk));
	jdff dff_A_1rQxkaMZ6_0(.dout(w_dff_A_UmwWKvEW7_0),.din(w_dff_A_1rQxkaMZ6_0),.clk(gclk));
	jdff dff_A_zXQNcWHq8_0(.dout(w_n578_1[0]),.din(w_dff_A_zXQNcWHq8_0),.clk(gclk));
	jdff dff_A_LZhMNDa49_0(.dout(w_dff_A_zXQNcWHq8_0),.din(w_dff_A_LZhMNDa49_0),.clk(gclk));
	jdff dff_A_IYbuSqnC5_0(.dout(w_dff_A_LZhMNDa49_0),.din(w_dff_A_IYbuSqnC5_0),.clk(gclk));
	jdff dff_A_hTIxALdH9_0(.dout(w_dff_A_IYbuSqnC5_0),.din(w_dff_A_hTIxALdH9_0),.clk(gclk));
	jdff dff_A_MKUfhvux9_0(.dout(w_dff_A_hTIxALdH9_0),.din(w_dff_A_MKUfhvux9_0),.clk(gclk));
	jdff dff_A_2mCGjD1i9_0(.dout(w_dff_A_MKUfhvux9_0),.din(w_dff_A_2mCGjD1i9_0),.clk(gclk));
	jdff dff_A_QL5ApbaD7_0(.dout(w_dff_A_2mCGjD1i9_0),.din(w_dff_A_QL5ApbaD7_0),.clk(gclk));
	jdff dff_A_Gz8E25yi4_0(.dout(w_dff_A_QL5ApbaD7_0),.din(w_dff_A_Gz8E25yi4_0),.clk(gclk));
	jdff dff_A_iuTt8jDK2_0(.dout(w_dff_A_Gz8E25yi4_0),.din(w_dff_A_iuTt8jDK2_0),.clk(gclk));
	jdff dff_A_4Px20A4r9_0(.dout(w_dff_A_iuTt8jDK2_0),.din(w_dff_A_4Px20A4r9_0),.clk(gclk));
	jdff dff_A_iK6pO9725_0(.dout(w_dff_A_4Px20A4r9_0),.din(w_dff_A_iK6pO9725_0),.clk(gclk));
	jdff dff_A_BLNwJD364_0(.dout(w_dff_A_iK6pO9725_0),.din(w_dff_A_BLNwJD364_0),.clk(gclk));
	jdff dff_A_GcFNFohd4_1(.dout(w_n578_0[1]),.din(w_dff_A_GcFNFohd4_1),.clk(gclk));
	jdff dff_A_GipSjDUt4_1(.dout(w_dff_A_GcFNFohd4_1),.din(w_dff_A_GipSjDUt4_1),.clk(gclk));
	jdff dff_A_OP4lTLMV3_1(.dout(w_dff_A_GipSjDUt4_1),.din(w_dff_A_OP4lTLMV3_1),.clk(gclk));
	jdff dff_A_qtJnsGNi4_1(.dout(w_dff_A_OP4lTLMV3_1),.din(w_dff_A_qtJnsGNi4_1),.clk(gclk));
	jdff dff_A_q2fnkuVw8_2(.dout(w_n578_0[2]),.din(w_dff_A_q2fnkuVw8_2),.clk(gclk));
	jdff dff_A_batIeYWG1_2(.dout(w_dff_A_q2fnkuVw8_2),.din(w_dff_A_batIeYWG1_2),.clk(gclk));
	jdff dff_A_OINP2Htl1_2(.dout(w_dff_A_batIeYWG1_2),.din(w_dff_A_OINP2Htl1_2),.clk(gclk));
	jdff dff_A_f7oh9e0H0_2(.dout(w_dff_A_OINP2Htl1_2),.din(w_dff_A_f7oh9e0H0_2),.clk(gclk));
	jdff dff_A_7qcirIbk1_2(.dout(w_dff_A_f7oh9e0H0_2),.din(w_dff_A_7qcirIbk1_2),.clk(gclk));
	jdff dff_A_NZAOmBEF5_2(.dout(w_dff_A_7qcirIbk1_2),.din(w_dff_A_NZAOmBEF5_2),.clk(gclk));
	jdff dff_A_Z41uG3Qb5_2(.dout(w_dff_A_NZAOmBEF5_2),.din(w_dff_A_Z41uG3Qb5_2),.clk(gclk));
	jdff dff_A_dct5lZS76_2(.dout(w_dff_A_Z41uG3Qb5_2),.din(w_dff_A_dct5lZS76_2),.clk(gclk));
	jdff dff_A_6B2059224_2(.dout(w_dff_A_dct5lZS76_2),.din(w_dff_A_6B2059224_2),.clk(gclk));
	jdff dff_A_kTiYQC3z8_2(.dout(w_dff_A_6B2059224_2),.din(w_dff_A_kTiYQC3z8_2),.clk(gclk));
	jdff dff_A_1G46lzN70_2(.dout(w_dff_A_kTiYQC3z8_2),.din(w_dff_A_1G46lzN70_2),.clk(gclk));
	jdff dff_A_AR6PB7eS3_2(.dout(w_dff_A_1G46lzN70_2),.din(w_dff_A_AR6PB7eS3_2),.clk(gclk));
	jdff dff_B_3C2QXZfv3_0(.din(n576),.dout(w_dff_B_3C2QXZfv3_0),.clk(gclk));
	jdff dff_B_rnocEosP8_0(.din(G147),.dout(w_dff_B_rnocEosP8_0),.clk(gclk));
	jdff dff_B_77YsmIWU1_2(.din(n574),.dout(w_dff_B_77YsmIWU1_2),.clk(gclk));
	jdff dff_B_sKxW7ouH5_2(.din(w_dff_B_77YsmIWU1_2),.dout(w_dff_B_sKxW7ouH5_2),.clk(gclk));
	jdff dff_A_wILlbT7T3_2(.dout(w_n573_0[2]),.din(w_dff_A_wILlbT7T3_2),.clk(gclk));
	jdff dff_A_4YWfzSay5_2(.dout(w_dff_A_wILlbT7T3_2),.din(w_dff_A_4YWfzSay5_2),.clk(gclk));
	jdff dff_A_Kne2JWyF3_2(.dout(w_dff_A_4YWfzSay5_2),.din(w_dff_A_Kne2JWyF3_2),.clk(gclk));
	jdff dff_A_6MKETmv02_2(.dout(w_dff_A_Kne2JWyF3_2),.din(w_dff_A_6MKETmv02_2),.clk(gclk));
	jdff dff_A_BFa9jBAm4_2(.dout(w_dff_A_6MKETmv02_2),.din(w_dff_A_BFa9jBAm4_2),.clk(gclk));
	jdff dff_A_UZhSkQ3u9_2(.dout(w_dff_A_BFa9jBAm4_2),.din(w_dff_A_UZhSkQ3u9_2),.clk(gclk));
	jdff dff_A_QcSwRD9w2_2(.dout(w_dff_A_UZhSkQ3u9_2),.din(w_dff_A_QcSwRD9w2_2),.clk(gclk));
	jdff dff_A_zFfFWEtR2_2(.dout(w_dff_A_QcSwRD9w2_2),.din(w_dff_A_zFfFWEtR2_2),.clk(gclk));
	jdff dff_A_yICARhwM9_2(.dout(w_dff_A_zFfFWEtR2_2),.din(w_dff_A_yICARhwM9_2),.clk(gclk));
	jdff dff_A_SW4xabWb7_2(.dout(w_dff_A_yICARhwM9_2),.din(w_dff_A_SW4xabWb7_2),.clk(gclk));
	jdff dff_A_rpso9bRS2_2(.dout(w_dff_A_SW4xabWb7_2),.din(w_dff_A_rpso9bRS2_2),.clk(gclk));
	jdff dff_A_gRtxQXhT5_2(.dout(w_dff_A_rpso9bRS2_2),.din(w_dff_A_gRtxQXhT5_2),.clk(gclk));
	jdff dff_A_txnbFa000_2(.dout(w_dff_A_gRtxQXhT5_2),.din(w_dff_A_txnbFa000_2),.clk(gclk));
	jdff dff_A_xnCWaTuR7_2(.dout(w_dff_A_txnbFa000_2),.din(w_dff_A_xnCWaTuR7_2),.clk(gclk));
	jdff dff_A_Ao79kSAN0_2(.dout(w_n572_0[2]),.din(w_dff_A_Ao79kSAN0_2),.clk(gclk));
	jdff dff_B_KhfQAqlt3_0(.din(n571),.dout(w_dff_B_KhfQAqlt3_0),.clk(gclk));
	jdff dff_B_3uEs4dVE0_0(.din(G138),.dout(w_dff_B_3uEs4dVE0_0),.clk(gclk));
	jdff dff_B_oNNov6Cs0_3(.din(n569),.dout(w_dff_B_oNNov6Cs0_3),.clk(gclk));
	jdff dff_B_syGTL4xv9_3(.din(w_dff_B_oNNov6Cs0_3),.dout(w_dff_B_syGTL4xv9_3),.clk(gclk));
	jdff dff_A_iL4NUDBV5_0(.dout(w_n568_0[0]),.din(w_dff_A_iL4NUDBV5_0),.clk(gclk));
	jdff dff_A_kb6YfBSF5_0(.dout(w_dff_A_iL4NUDBV5_0),.din(w_dff_A_kb6YfBSF5_0),.clk(gclk));
	jdff dff_A_bUkzMEKL9_0(.dout(w_dff_A_kb6YfBSF5_0),.din(w_dff_A_bUkzMEKL9_0),.clk(gclk));
	jdff dff_A_7k2u0Uhk4_0(.dout(w_dff_A_bUkzMEKL9_0),.din(w_dff_A_7k2u0Uhk4_0),.clk(gclk));
	jdff dff_A_mBGChZA09_2(.dout(w_n568_0[2]),.din(w_dff_A_mBGChZA09_2),.clk(gclk));
	jdff dff_A_KB6PSNHp2_2(.dout(w_dff_A_mBGChZA09_2),.din(w_dff_A_KB6PSNHp2_2),.clk(gclk));
	jdff dff_B_gkRoOqZ43_0(.din(G157),.dout(w_dff_B_gkRoOqZ43_0),.clk(gclk));
	jdff dff_A_FdM5IzSU3_0(.dout(w_n564_0[0]),.din(w_dff_A_FdM5IzSU3_0),.clk(gclk));
	jdff dff_A_yGaO7Vih8_0(.dout(w_dff_A_FdM5IzSU3_0),.din(w_dff_A_yGaO7Vih8_0),.clk(gclk));
	jdff dff_A_VMS3oj4g6_0(.dout(w_dff_A_yGaO7Vih8_0),.din(w_dff_A_VMS3oj4g6_0),.clk(gclk));
	jdff dff_A_d8qwEVrX0_1(.dout(w_n564_0[1]),.din(w_dff_A_d8qwEVrX0_1),.clk(gclk));
	jdff dff_B_yVkI5nMr4_2(.din(n563),.dout(w_dff_B_yVkI5nMr4_2),.clk(gclk));
	jdff dff_B_YAXYqcGI0_2(.din(w_dff_B_yVkI5nMr4_2),.dout(w_dff_B_YAXYqcGI0_2),.clk(gclk));
	jdff dff_A_u6ht5Zzm1_0(.dout(w_G2236_1[0]),.din(w_dff_A_u6ht5Zzm1_0),.clk(gclk));
	jdff dff_A_fPsIodG79_0(.dout(w_dff_A_u6ht5Zzm1_0),.din(w_dff_A_fPsIodG79_0),.clk(gclk));
	jdff dff_A_soUu5tBA0_0(.dout(w_dff_A_fPsIodG79_0),.din(w_dff_A_soUu5tBA0_0),.clk(gclk));
	jdff dff_A_j7vDye4R5_0(.dout(w_dff_A_soUu5tBA0_0),.din(w_dff_A_j7vDye4R5_0),.clk(gclk));
	jdff dff_B_6qNqKJ7I7_0(.din(n561),.dout(w_dff_B_6qNqKJ7I7_0),.clk(gclk));
	jdff dff_B_zhQ5zoaN3_0(.din(w_dff_B_6qNqKJ7I7_0),.dout(w_dff_B_zhQ5zoaN3_0),.clk(gclk));
	jdff dff_B_oZxpILHP5_0(.din(w_dff_B_zhQ5zoaN3_0),.dout(w_dff_B_oZxpILHP5_0),.clk(gclk));
	jdff dff_B_eqNB2x3B1_0(.din(w_dff_B_oZxpILHP5_0),.dout(w_dff_B_eqNB2x3B1_0),.clk(gclk));
	jdff dff_A_pf5blDt83_0(.dout(w_n560_0[0]),.din(w_dff_A_pf5blDt83_0),.clk(gclk));
	jdff dff_A_GJmzwBgT8_0(.dout(w_dff_A_pf5blDt83_0),.din(w_dff_A_GJmzwBgT8_0),.clk(gclk));
	jdff dff_A_j8v0MkH30_0(.dout(w_dff_A_GJmzwBgT8_0),.din(w_dff_A_j8v0MkH30_0),.clk(gclk));
	jdff dff_A_ugtOsKZg0_0(.dout(w_dff_A_j8v0MkH30_0),.din(w_dff_A_ugtOsKZg0_0),.clk(gclk));
	jdff dff_A_GOtlVnN46_0(.dout(w_dff_A_ugtOsKZg0_0),.din(w_dff_A_GOtlVnN46_0),.clk(gclk));
	jdff dff_B_j2k8mZZE5_1(.din(n547),.dout(w_dff_B_j2k8mZZE5_1),.clk(gclk));
	jdff dff_B_v4dk76pM1_1(.din(w_dff_B_j2k8mZZE5_1),.dout(w_dff_B_v4dk76pM1_1),.clk(gclk));
	jdff dff_B_INxAodTD2_1(.din(w_dff_B_v4dk76pM1_1),.dout(w_dff_B_INxAodTD2_1),.clk(gclk));
	jdff dff_B_3EeUhV7m3_1(.din(n548),.dout(w_dff_B_3EeUhV7m3_1),.clk(gclk));
	jdff dff_B_4KCJDPpx6_1(.din(w_dff_B_3EeUhV7m3_1),.dout(w_dff_B_4KCJDPpx6_1),.clk(gclk));
	jdff dff_B_YYMfaYUU9_1(.din(w_dff_B_4KCJDPpx6_1),.dout(w_dff_B_YYMfaYUU9_1),.clk(gclk));
	jdff dff_B_bU2JFqUT9_1(.din(w_dff_B_YYMfaYUU9_1),.dout(w_dff_B_bU2JFqUT9_1),.clk(gclk));
	jdff dff_B_DTSOZ4kH2_0(.din(n543),.dout(w_dff_B_DTSOZ4kH2_0),.clk(gclk));
	jdff dff_B_HVTNJEOF6_0(.din(w_dff_B_DTSOZ4kH2_0),.dout(w_dff_B_HVTNJEOF6_0),.clk(gclk));
	jdff dff_B_SnIFAloN7_0(.din(w_dff_B_HVTNJEOF6_0),.dout(w_dff_B_SnIFAloN7_0),.clk(gclk));
	jdff dff_B_6UuhMnFy3_0(.din(w_dff_B_SnIFAloN7_0),.dout(w_dff_B_6UuhMnFy3_0),.clk(gclk));
	jdff dff_B_6h0p151i4_0(.din(w_dff_B_6UuhMnFy3_0),.dout(w_dff_B_6h0p151i4_0),.clk(gclk));
	jdff dff_B_g93XN7Hd9_0(.din(w_dff_B_6h0p151i4_0),.dout(w_dff_B_g93XN7Hd9_0),.clk(gclk));
	jdff dff_B_Cd0jMb9i0_0(.din(w_dff_B_g93XN7Hd9_0),.dout(w_dff_B_Cd0jMb9i0_0),.clk(gclk));
	jdff dff_A_0tNitACA4_0(.dout(w_n542_0[0]),.din(w_dff_A_0tNitACA4_0),.clk(gclk));
	jdff dff_A_NqvdE97N4_0(.dout(w_dff_A_0tNitACA4_0),.din(w_dff_A_NqvdE97N4_0),.clk(gclk));
	jdff dff_A_V0ljnoLg8_0(.dout(w_dff_A_NqvdE97N4_0),.din(w_dff_A_V0ljnoLg8_0),.clk(gclk));
	jdff dff_A_ccNtsWX08_0(.dout(w_dff_A_V0ljnoLg8_0),.din(w_dff_A_ccNtsWX08_0),.clk(gclk));
	jdff dff_A_FIyJsI0G3_0(.dout(w_dff_A_ccNtsWX08_0),.din(w_dff_A_FIyJsI0G3_0),.clk(gclk));
	jdff dff_A_xnYzgbV02_0(.dout(w_dff_A_FIyJsI0G3_0),.din(w_dff_A_xnYzgbV02_0),.clk(gclk));
	jdff dff_A_5Z8h4EPz9_0(.dout(w_dff_A_xnYzgbV02_0),.din(w_dff_A_5Z8h4EPz9_0),.clk(gclk));
	jdff dff_A_DjpXitUl9_0(.dout(w_dff_A_5Z8h4EPz9_0),.din(w_dff_A_DjpXitUl9_0),.clk(gclk));
	jdff dff_A_JovB0lwN3_0(.dout(w_n535_1[0]),.din(w_dff_A_JovB0lwN3_0),.clk(gclk));
	jdff dff_A_E5K7alzc4_0(.dout(w_dff_A_JovB0lwN3_0),.din(w_dff_A_E5K7alzc4_0),.clk(gclk));
	jdff dff_A_KJ3vDEya8_0(.dout(w_dff_A_E5K7alzc4_0),.din(w_dff_A_KJ3vDEya8_0),.clk(gclk));
	jdff dff_A_eheffV112_0(.dout(w_dff_A_KJ3vDEya8_0),.din(w_dff_A_eheffV112_0),.clk(gclk));
	jdff dff_A_joYyMP7n7_0(.dout(w_dff_A_eheffV112_0),.din(w_dff_A_joYyMP7n7_0),.clk(gclk));
	jdff dff_A_KU3rHIqv9_0(.dout(w_dff_A_joYyMP7n7_0),.din(w_dff_A_KU3rHIqv9_0),.clk(gclk));
	jdff dff_A_hB3e9Lal8_0(.dout(w_dff_A_KU3rHIqv9_0),.din(w_dff_A_hB3e9Lal8_0),.clk(gclk));
	jdff dff_A_czRxNlFA7_0(.dout(w_dff_A_hB3e9Lal8_0),.din(w_dff_A_czRxNlFA7_0),.clk(gclk));
	jdff dff_A_xfECxXcF3_0(.dout(w_dff_A_czRxNlFA7_0),.din(w_dff_A_xfECxXcF3_0),.clk(gclk));
	jdff dff_A_PJSjd5ZO0_0(.dout(w_dff_A_xfECxXcF3_0),.din(w_dff_A_PJSjd5ZO0_0),.clk(gclk));
	jdff dff_A_EXpZaSpZ3_0(.dout(w_dff_A_PJSjd5ZO0_0),.din(w_dff_A_EXpZaSpZ3_0),.clk(gclk));
	jdff dff_A_R5aBBOiV2_0(.dout(w_dff_A_EXpZaSpZ3_0),.din(w_dff_A_R5aBBOiV2_0),.clk(gclk));
	jdff dff_A_1GIilQCR3_0(.dout(w_dff_A_R5aBBOiV2_0),.din(w_dff_A_1GIilQCR3_0),.clk(gclk));
	jdff dff_A_px7SGiXE3_0(.dout(w_n530_0[0]),.din(w_dff_A_px7SGiXE3_0),.clk(gclk));
	jdff dff_A_m3rSiGQ31_0(.dout(w_dff_A_px7SGiXE3_0),.din(w_dff_A_m3rSiGQ31_0),.clk(gclk));
	jdff dff_A_suR2No9l5_0(.dout(w_dff_A_m3rSiGQ31_0),.din(w_dff_A_suR2No9l5_0),.clk(gclk));
	jdff dff_A_0NvkXn7P2_0(.dout(w_dff_A_suR2No9l5_0),.din(w_dff_A_0NvkXn7P2_0),.clk(gclk));
	jdff dff_A_Mk4ll8HJ2_0(.dout(w_dff_A_0NvkXn7P2_0),.din(w_dff_A_Mk4ll8HJ2_0),.clk(gclk));
	jdff dff_A_G0ExnXCE7_0(.dout(w_dff_A_Mk4ll8HJ2_0),.din(w_dff_A_G0ExnXCE7_0),.clk(gclk));
	jdff dff_A_niLYAnRN9_0(.dout(w_dff_A_G0ExnXCE7_0),.din(w_dff_A_niLYAnRN9_0),.clk(gclk));
	jdff dff_A_BFIbBuJj1_0(.dout(w_dff_A_niLYAnRN9_0),.din(w_dff_A_BFIbBuJj1_0),.clk(gclk));
	jdff dff_A_CmHLRX2u3_0(.dout(w_dff_A_BFIbBuJj1_0),.din(w_dff_A_CmHLRX2u3_0),.clk(gclk));
	jdff dff_A_CJ2XfhFk2_0(.dout(w_n529_0[0]),.din(w_dff_A_CJ2XfhFk2_0),.clk(gclk));
	jdff dff_A_VCRb9KBz1_0(.dout(w_dff_A_CJ2XfhFk2_0),.din(w_dff_A_VCRb9KBz1_0),.clk(gclk));
	jdff dff_A_wh4rldlH9_0(.dout(w_dff_A_VCRb9KBz1_0),.din(w_dff_A_wh4rldlH9_0),.clk(gclk));
	jdff dff_A_kusIEkBs1_0(.dout(w_dff_A_wh4rldlH9_0),.din(w_dff_A_kusIEkBs1_0),.clk(gclk));
	jdff dff_A_DpbZDXwP0_0(.dout(w_dff_A_kusIEkBs1_0),.din(w_dff_A_DpbZDXwP0_0),.clk(gclk));
	jdff dff_A_lPdV6RPk9_0(.dout(w_dff_A_DpbZDXwP0_0),.din(w_dff_A_lPdV6RPk9_0),.clk(gclk));
	jdff dff_A_dDUxUmdE1_0(.dout(w_dff_A_lPdV6RPk9_0),.din(w_dff_A_dDUxUmdE1_0),.clk(gclk));
	jdff dff_A_mmuEb3QL8_0(.dout(w_dff_A_dDUxUmdE1_0),.din(w_dff_A_mmuEb3QL8_0),.clk(gclk));
	jdff dff_A_AhamDzMV9_0(.dout(w_dff_A_mmuEb3QL8_0),.din(w_dff_A_AhamDzMV9_0),.clk(gclk));
	jdff dff_A_CscisU493_0(.dout(w_dff_A_AhamDzMV9_0),.din(w_dff_A_CscisU493_0),.clk(gclk));
	jdff dff_A_vO6IatWr4_0(.dout(w_n1463_0[0]),.din(w_dff_A_vO6IatWr4_0),.clk(gclk));
	jdff dff_A_rJFI9lK38_0(.dout(w_dff_A_vO6IatWr4_0),.din(w_dff_A_rJFI9lK38_0),.clk(gclk));
	jdff dff_A_qKcgb3jQ7_0(.dout(w_dff_A_rJFI9lK38_0),.din(w_dff_A_qKcgb3jQ7_0),.clk(gclk));
	jdff dff_A_gDjcuU4m7_0(.dout(w_dff_A_qKcgb3jQ7_0),.din(w_dff_A_gDjcuU4m7_0),.clk(gclk));
	jdff dff_A_KfEs8R6r0_0(.dout(w_dff_A_gDjcuU4m7_0),.din(w_dff_A_KfEs8R6r0_0),.clk(gclk));
	jdff dff_A_kRLrKGtV7_0(.dout(w_dff_A_KfEs8R6r0_0),.din(w_dff_A_kRLrKGtV7_0),.clk(gclk));
	jdff dff_A_HiBM4pVC7_0(.dout(w_dff_A_kRLrKGtV7_0),.din(w_dff_A_HiBM4pVC7_0),.clk(gclk));
	jdff dff_A_EGetv3MI1_0(.dout(w_dff_A_HiBM4pVC7_0),.din(w_dff_A_EGetv3MI1_0),.clk(gclk));
	jdff dff_A_cKy94sAX5_0(.dout(w_dff_A_EGetv3MI1_0),.din(w_dff_A_cKy94sAX5_0),.clk(gclk));
	jdff dff_A_tXHQJMnv0_0(.dout(w_dff_A_cKy94sAX5_0),.din(w_dff_A_tXHQJMnv0_0),.clk(gclk));
	jdff dff_A_ZxbK0vmW0_0(.dout(w_dff_A_tXHQJMnv0_0),.din(w_dff_A_ZxbK0vmW0_0),.clk(gclk));
	jdff dff_A_gMf7R9sU2_1(.dout(w_n1463_0[1]),.din(w_dff_A_gMf7R9sU2_1),.clk(gclk));
	jdff dff_A_D5fs9vIB1_1(.dout(w_dff_A_gMf7R9sU2_1),.din(w_dff_A_D5fs9vIB1_1),.clk(gclk));
	jdff dff_A_3K7rC5Qk6_1(.dout(w_dff_A_D5fs9vIB1_1),.din(w_dff_A_3K7rC5Qk6_1),.clk(gclk));
	jdff dff_A_WiNWTh6M3_1(.dout(w_dff_A_3K7rC5Qk6_1),.din(w_dff_A_WiNWTh6M3_1),.clk(gclk));
	jdff dff_A_AZaIBfQd3_1(.dout(w_dff_A_WiNWTh6M3_1),.din(w_dff_A_AZaIBfQd3_1),.clk(gclk));
	jdff dff_A_0gFLWxzC7_1(.dout(w_dff_A_AZaIBfQd3_1),.din(w_dff_A_0gFLWxzC7_1),.clk(gclk));
	jdff dff_A_ranaJklK5_1(.dout(w_dff_A_0gFLWxzC7_1),.din(w_dff_A_ranaJklK5_1),.clk(gclk));
	jdff dff_A_4FRVz7XB5_1(.dout(w_dff_A_ranaJklK5_1),.din(w_dff_A_4FRVz7XB5_1),.clk(gclk));
	jdff dff_A_jEvkwzsX6_1(.dout(w_dff_A_4FRVz7XB5_1),.din(w_dff_A_jEvkwzsX6_1),.clk(gclk));
	jdff dff_A_t6sEAL5Z8_1(.dout(w_dff_A_jEvkwzsX6_1),.din(w_dff_A_t6sEAL5Z8_1),.clk(gclk));
	jdff dff_A_iwIUXNDC4_1(.dout(w_dff_A_t6sEAL5Z8_1),.din(w_dff_A_iwIUXNDC4_1),.clk(gclk));
	jdff dff_A_MbKVSPC10_1(.dout(w_dff_A_iwIUXNDC4_1),.din(w_dff_A_MbKVSPC10_1),.clk(gclk));
	jdff dff_A_hfE9EebZ0_1(.dout(w_dff_A_MbKVSPC10_1),.din(w_dff_A_hfE9EebZ0_1),.clk(gclk));
	jdff dff_A_2LREpPro2_1(.dout(w_dff_A_hfE9EebZ0_1),.din(w_dff_A_2LREpPro2_1),.clk(gclk));
	jdff dff_A_GAxHeVLN5_1(.dout(w_dff_A_2LREpPro2_1),.din(w_dff_A_GAxHeVLN5_1),.clk(gclk));
	jdff dff_A_bvKcreuB4_1(.dout(w_dff_A_GAxHeVLN5_1),.din(w_dff_A_bvKcreuB4_1),.clk(gclk));
	jdff dff_A_hIUtR8a03_1(.dout(w_dff_A_bvKcreuB4_1),.din(w_dff_A_hIUtR8a03_1),.clk(gclk));
	jdff dff_A_PBd0LuDz8_1(.dout(w_dff_A_hIUtR8a03_1),.din(w_dff_A_PBd0LuDz8_1),.clk(gclk));
	jdff dff_A_RGme1VQO3_1(.dout(w_dff_A_PBd0LuDz8_1),.din(w_dff_A_RGme1VQO3_1),.clk(gclk));
	jdff dff_B_uHLU5VDr0_0(.din(n1462),.dout(w_dff_B_uHLU5VDr0_0),.clk(gclk));
	jdff dff_A_eAUesVzk7_1(.dout(w_n365_0[1]),.din(w_dff_A_eAUesVzk7_1),.clk(gclk));
	jdff dff_A_xFztVBjF1_1(.dout(w_dff_A_eAUesVzk7_1),.din(w_dff_A_xFztVBjF1_1),.clk(gclk));
	jdff dff_A_xmevM6pX6_1(.dout(w_dff_A_xFztVBjF1_1),.din(w_dff_A_xmevM6pX6_1),.clk(gclk));
	jdff dff_A_IjN4mPtd6_1(.dout(w_dff_A_xmevM6pX6_1),.din(w_dff_A_IjN4mPtd6_1),.clk(gclk));
	jdff dff_A_5KN7Waln8_1(.dout(w_dff_A_IjN4mPtd6_1),.din(w_dff_A_5KN7Waln8_1),.clk(gclk));
	jdff dff_A_oeUb5HEf1_1(.dout(w_dff_A_5KN7Waln8_1),.din(w_dff_A_oeUb5HEf1_1),.clk(gclk));
	jdff dff_A_WgF7CZ8P1_1(.dout(w_dff_A_oeUb5HEf1_1),.din(w_dff_A_WgF7CZ8P1_1),.clk(gclk));
	jdff dff_A_2VlzlvdJ3_1(.dout(w_dff_A_WgF7CZ8P1_1),.din(w_dff_A_2VlzlvdJ3_1),.clk(gclk));
	jdff dff_A_aeGU1Iix2_1(.dout(w_dff_A_2VlzlvdJ3_1),.din(w_dff_A_aeGU1Iix2_1),.clk(gclk));
	jdff dff_A_t5iGKbeR6_1(.dout(w_dff_A_aeGU1Iix2_1),.din(w_dff_A_t5iGKbeR6_1),.clk(gclk));
	jdff dff_A_gx9i3qNR3_1(.dout(w_dff_A_t5iGKbeR6_1),.din(w_dff_A_gx9i3qNR3_1),.clk(gclk));
	jdff dff_A_6aVfz3u40_1(.dout(w_dff_A_gx9i3qNR3_1),.din(w_dff_A_6aVfz3u40_1),.clk(gclk));
	jdff dff_A_DrolHScC2_1(.dout(w_dff_A_6aVfz3u40_1),.din(w_dff_A_DrolHScC2_1),.clk(gclk));
	jdff dff_A_S4OE00AN7_1(.dout(w_dff_A_DrolHScC2_1),.din(w_dff_A_S4OE00AN7_1),.clk(gclk));
	jdff dff_A_R9H01SW31_1(.dout(w_dff_A_S4OE00AN7_1),.din(w_dff_A_R9H01SW31_1),.clk(gclk));
	jdff dff_A_n78vXkR71_1(.dout(w_dff_A_R9H01SW31_1),.din(w_dff_A_n78vXkR71_1),.clk(gclk));
	jdff dff_A_eagtifbf5_1(.dout(w_dff_A_n78vXkR71_1),.din(w_dff_A_eagtifbf5_1),.clk(gclk));
	jdff dff_A_DInUTTPn0_1(.dout(w_dff_A_eagtifbf5_1),.din(w_dff_A_DInUTTPn0_1),.clk(gclk));
	jdff dff_A_dzkYWVGd4_1(.dout(w_dff_A_DInUTTPn0_1),.din(w_dff_A_dzkYWVGd4_1),.clk(gclk));
	jdff dff_A_EvcAKS2p6_1(.dout(w_dff_A_dzkYWVGd4_1),.din(w_dff_A_EvcAKS2p6_1),.clk(gclk));
	jdff dff_A_9zWEW9xr4_1(.dout(w_dff_A_EvcAKS2p6_1),.din(w_dff_A_9zWEW9xr4_1),.clk(gclk));
	jdff dff_A_FDYHxj9q1_0(.dout(w_G38_1[0]),.din(w_dff_A_FDYHxj9q1_0),.clk(gclk));
	jdff dff_A_YVjUeDoE8_0(.dout(w_dff_A_FDYHxj9q1_0),.din(w_dff_A_YVjUeDoE8_0),.clk(gclk));
	jdff dff_A_5gGa3kNr3_0(.dout(w_dff_A_YVjUeDoE8_0),.din(w_dff_A_5gGa3kNr3_0),.clk(gclk));
	jdff dff_A_VmzUsI6k4_2(.dout(w_G38_1[2]),.din(w_dff_A_VmzUsI6k4_2),.clk(gclk));
	jdff dff_A_WJWqTm6j3_1(.dout(w_G38_0[1]),.din(w_dff_A_WJWqTm6j3_1),.clk(gclk));
	jdff dff_A_GrQxdQNd2_2(.dout(w_G38_0[2]),.din(w_dff_A_GrQxdQNd2_2),.clk(gclk));
	jdff dff_A_DvvVmoVy6_2(.dout(w_dff_A_GrQxdQNd2_2),.din(w_dff_A_DvvVmoVy6_2),.clk(gclk));
	jdff dff_B_H54XB8QL4_1(.din(n1587),.dout(w_dff_B_H54XB8QL4_1),.clk(gclk));
	jdff dff_B_kEK1mXdw5_1(.din(w_dff_B_H54XB8QL4_1),.dout(w_dff_B_kEK1mXdw5_1),.clk(gclk));
	jdff dff_B_5dHBPNPx4_1(.din(w_dff_B_kEK1mXdw5_1),.dout(w_dff_B_5dHBPNPx4_1),.clk(gclk));
	jdff dff_B_mIULG2T30_1(.din(w_dff_B_5dHBPNPx4_1),.dout(w_dff_B_mIULG2T30_1),.clk(gclk));
	jdff dff_B_2zhiKpty8_1(.din(w_dff_B_mIULG2T30_1),.dout(w_dff_B_2zhiKpty8_1),.clk(gclk));
	jdff dff_B_4A3Dnlax8_1(.din(w_dff_B_2zhiKpty8_1),.dout(w_dff_B_4A3Dnlax8_1),.clk(gclk));
	jdff dff_B_pA6yzUWF7_1(.din(w_dff_B_4A3Dnlax8_1),.dout(w_dff_B_pA6yzUWF7_1),.clk(gclk));
	jdff dff_B_60QWl5sd9_1(.din(w_dff_B_pA6yzUWF7_1),.dout(w_dff_B_60QWl5sd9_1),.clk(gclk));
	jdff dff_B_xqiXDl2v5_1(.din(w_dff_B_60QWl5sd9_1),.dout(w_dff_B_xqiXDl2v5_1),.clk(gclk));
	jdff dff_B_ceOtUC3a3_1(.din(w_dff_B_xqiXDl2v5_1),.dout(w_dff_B_ceOtUC3a3_1),.clk(gclk));
	jdff dff_B_WPeyNfHw0_1(.din(w_dff_B_ceOtUC3a3_1),.dout(w_dff_B_WPeyNfHw0_1),.clk(gclk));
	jdff dff_B_ASHbUCWz7_1(.din(w_dff_B_WPeyNfHw0_1),.dout(w_dff_B_ASHbUCWz7_1),.clk(gclk));
	jdff dff_B_OKEBBw1v9_1(.din(n1606),.dout(w_dff_B_OKEBBw1v9_1),.clk(gclk));
	jdff dff_B_xMBW8gtM9_1(.din(w_dff_B_OKEBBw1v9_1),.dout(w_dff_B_xMBW8gtM9_1),.clk(gclk));
	jdff dff_B_ez4oe8O89_1(.din(n1620),.dout(w_dff_B_ez4oe8O89_1),.clk(gclk));
	jdff dff_B_tP5QGGy90_1(.din(w_dff_B_ez4oe8O89_1),.dout(w_dff_B_tP5QGGy90_1),.clk(gclk));
	jdff dff_B_4Gm3sYUt8_1(.din(n1622),.dout(w_dff_B_4Gm3sYUt8_1),.clk(gclk));
	jdff dff_B_FUVbq3kE0_1(.din(w_dff_B_4Gm3sYUt8_1),.dout(w_dff_B_FUVbq3kE0_1),.clk(gclk));
	jdff dff_B_82E0SqC84_1(.din(w_dff_B_FUVbq3kE0_1),.dout(w_dff_B_82E0SqC84_1),.clk(gclk));
	jdff dff_B_H0YLKs2Y6_1(.din(w_dff_B_82E0SqC84_1),.dout(w_dff_B_H0YLKs2Y6_1),.clk(gclk));
	jdff dff_B_AMKVK5VG7_1(.din(w_dff_B_H0YLKs2Y6_1),.dout(w_dff_B_AMKVK5VG7_1),.clk(gclk));
	jdff dff_B_79HMWNLb4_1(.din(w_dff_B_AMKVK5VG7_1),.dout(w_dff_B_79HMWNLb4_1),.clk(gclk));
	jdff dff_B_nw132nbh3_1(.din(n1623),.dout(w_dff_B_nw132nbh3_1),.clk(gclk));
	jdff dff_B_wwJVCGX44_1(.din(w_dff_B_nw132nbh3_1),.dout(w_dff_B_wwJVCGX44_1),.clk(gclk));
	jdff dff_B_MkWhOmse4_1(.din(w_dff_B_wwJVCGX44_1),.dout(w_dff_B_MkWhOmse4_1),.clk(gclk));
	jdff dff_B_MjDQdwRa4_1(.din(w_dff_B_MkWhOmse4_1),.dout(w_dff_B_MjDQdwRa4_1),.clk(gclk));
	jdff dff_B_1UGtU2pP1_1(.din(w_dff_B_MjDQdwRa4_1),.dout(w_dff_B_1UGtU2pP1_1),.clk(gclk));
	jdff dff_B_eYsFY6Dz2_1(.din(w_dff_B_1UGtU2pP1_1),.dout(w_dff_B_eYsFY6Dz2_1),.clk(gclk));
	jdff dff_B_ldlJ2nWL0_1(.din(w_dff_B_eYsFY6Dz2_1),.dout(w_dff_B_ldlJ2nWL0_1),.clk(gclk));
	jdff dff_B_lxx2CanO3_1(.din(w_dff_B_ldlJ2nWL0_1),.dout(w_dff_B_lxx2CanO3_1),.clk(gclk));
	jdff dff_B_tmvJ6XVG7_1(.din(n1626),.dout(w_dff_B_tmvJ6XVG7_1),.clk(gclk));
	jdff dff_B_nGaZYB9h6_1(.din(w_dff_B_tmvJ6XVG7_1),.dout(w_dff_B_nGaZYB9h6_1),.clk(gclk));
	jdff dff_B_9XJZ6PK16_0(.din(n1624),.dout(w_dff_B_9XJZ6PK16_0),.clk(gclk));
	jdff dff_B_4stDTBS90_0(.din(w_dff_B_9XJZ6PK16_0),.dout(w_dff_B_4stDTBS90_0),.clk(gclk));
	jdff dff_A_g0sE4gYu5_1(.dout(w_n1479_0[1]),.din(w_dff_A_g0sE4gYu5_1),.clk(gclk));
	jdff dff_A_WG64xLY17_1(.dout(w_dff_A_g0sE4gYu5_1),.din(w_dff_A_WG64xLY17_1),.clk(gclk));
	jdff dff_A_sjwH9waE9_1(.dout(w_dff_A_WG64xLY17_1),.din(w_dff_A_sjwH9waE9_1),.clk(gclk));
	jdff dff_A_Qzifh2BF2_1(.dout(w_dff_A_sjwH9waE9_1),.din(w_dff_A_Qzifh2BF2_1),.clk(gclk));
	jdff dff_A_XyOJ4ZVF4_1(.dout(w_dff_A_Qzifh2BF2_1),.din(w_dff_A_XyOJ4ZVF4_1),.clk(gclk));
	jdff dff_A_KtsyxYg13_1(.dout(w_dff_A_XyOJ4ZVF4_1),.din(w_dff_A_KtsyxYg13_1),.clk(gclk));
	jdff dff_A_Ed8GysSM6_1(.dout(w_n1471_0[1]),.din(w_dff_A_Ed8GysSM6_1),.clk(gclk));
	jdff dff_A_VkjFpfeo2_1(.dout(w_dff_A_Ed8GysSM6_1),.din(w_dff_A_VkjFpfeo2_1),.clk(gclk));
	jdff dff_A_L9MFRLub6_1(.dout(w_dff_A_VkjFpfeo2_1),.din(w_dff_A_L9MFRLub6_1),.clk(gclk));
	jdff dff_A_t1OorFeT8_1(.dout(w_dff_A_L9MFRLub6_1),.din(w_dff_A_t1OorFeT8_1),.clk(gclk));
	jdff dff_A_pJKJ5JGS9_1(.dout(w_dff_A_t1OorFeT8_1),.din(w_dff_A_pJKJ5JGS9_1),.clk(gclk));
	jdff dff_B_AFVHb2Dm8_1(.din(n1609),.dout(w_dff_B_AFVHb2Dm8_1),.clk(gclk));
	jdff dff_B_VTOZJaWd5_1(.din(w_dff_B_AFVHb2Dm8_1),.dout(w_dff_B_VTOZJaWd5_1),.clk(gclk));
	jdff dff_B_zMT5VBaP1_1(.din(w_dff_B_VTOZJaWd5_1),.dout(w_dff_B_zMT5VBaP1_1),.clk(gclk));
	jdff dff_B_Jmwo1Vpq5_1(.din(w_dff_B_zMT5VBaP1_1),.dout(w_dff_B_Jmwo1Vpq5_1),.clk(gclk));
	jdff dff_B_hIlveP8D7_1(.din(w_dff_B_Jmwo1Vpq5_1),.dout(w_dff_B_hIlveP8D7_1),.clk(gclk));
	jdff dff_B_2yNwb2Rz4_1(.din(w_dff_B_hIlveP8D7_1),.dout(w_dff_B_2yNwb2Rz4_1),.clk(gclk));
	jdff dff_B_XKqHvp1z8_0(.din(n1615),.dout(w_dff_B_XKqHvp1z8_0),.clk(gclk));
	jdff dff_A_KjU7AqUT0_1(.dout(w_n1482_0[1]),.din(w_dff_A_KjU7AqUT0_1),.clk(gclk));
	jdff dff_A_tLo5OXNk5_1(.dout(w_dff_A_KjU7AqUT0_1),.din(w_dff_A_tLo5OXNk5_1),.clk(gclk));
	jdff dff_A_5lvn2ewi5_1(.dout(w_dff_A_tLo5OXNk5_1),.din(w_dff_A_5lvn2ewi5_1),.clk(gclk));
	jdff dff_A_W1Q2ulZp0_1(.dout(w_dff_A_5lvn2ewi5_1),.din(w_dff_A_W1Q2ulZp0_1),.clk(gclk));
	jdff dff_A_iO7mZrfs7_1(.dout(w_dff_A_W1Q2ulZp0_1),.din(w_dff_A_iO7mZrfs7_1),.clk(gclk));
	jdff dff_A_Y5jRghTd6_1(.dout(w_dff_A_iO7mZrfs7_1),.din(w_dff_A_Y5jRghTd6_1),.clk(gclk));
	jdff dff_A_0WAxktpG4_1(.dout(w_dff_A_Y5jRghTd6_1),.din(w_dff_A_0WAxktpG4_1),.clk(gclk));
	jdff dff_A_syDZq2026_1(.dout(w_n1468_0[1]),.din(w_dff_A_syDZq2026_1),.clk(gclk));
	jdff dff_A_F77pSxzR3_1(.dout(w_dff_A_syDZq2026_1),.din(w_dff_A_F77pSxzR3_1),.clk(gclk));
	jdff dff_A_jLvMlcrl4_1(.dout(w_dff_A_F77pSxzR3_1),.din(w_dff_A_jLvMlcrl4_1),.clk(gclk));
	jdff dff_A_JR4JKGp92_1(.dout(w_dff_A_jLvMlcrl4_1),.din(w_dff_A_JR4JKGp92_1),.clk(gclk));
	jdff dff_A_vaUUkInl2_1(.dout(w_dff_A_JR4JKGp92_1),.din(w_dff_A_vaUUkInl2_1),.clk(gclk));
	jdff dff_B_donYkLVC3_2(.din(n1468),.dout(w_dff_B_donYkLVC3_2),.clk(gclk));
	jdff dff_B_mbjCN1LT8_2(.din(w_dff_B_donYkLVC3_2),.dout(w_dff_B_mbjCN1LT8_2),.clk(gclk));
	jdff dff_B_IoS9XBZo6_2(.din(w_dff_B_mbjCN1LT8_2),.dout(w_dff_B_IoS9XBZo6_2),.clk(gclk));
	jdff dff_B_WdTyTBTI2_2(.din(w_dff_B_IoS9XBZo6_2),.dout(w_dff_B_WdTyTBTI2_2),.clk(gclk));
	jdff dff_B_p5naMZBK5_2(.din(w_dff_B_WdTyTBTI2_2),.dout(w_dff_B_p5naMZBK5_2),.clk(gclk));
	jdff dff_B_jllnJNpC9_2(.din(w_dff_B_p5naMZBK5_2),.dout(w_dff_B_jllnJNpC9_2),.clk(gclk));
	jdff dff_B_2ZlPMjFp5_2(.din(n1610),.dout(w_dff_B_2ZlPMjFp5_2),.clk(gclk));
	jdff dff_B_4ORWPjYZ0_1(.din(n1607),.dout(w_dff_B_4ORWPjYZ0_1),.clk(gclk));
	jdff dff_B_IERriCYy9_0(.din(n1604),.dout(w_dff_B_IERriCYy9_0),.clk(gclk));
	jdff dff_B_EjHF14WT6_0(.din(w_dff_B_IERriCYy9_0),.dout(w_dff_B_EjHF14WT6_0),.clk(gclk));
	jdff dff_B_ornnWYyA2_1(.din(n1597),.dout(w_dff_B_ornnWYyA2_1),.clk(gclk));
	jdff dff_B_IDeAhHgO2_1(.din(w_dff_B_ornnWYyA2_1),.dout(w_dff_B_IDeAhHgO2_1),.clk(gclk));
	jdff dff_B_86ioJiNl5_1(.din(w_dff_B_IDeAhHgO2_1),.dout(w_dff_B_86ioJiNl5_1),.clk(gclk));
	jdff dff_B_DpYNnzbp2_1(.din(w_dff_B_86ioJiNl5_1),.dout(w_dff_B_DpYNnzbp2_1),.clk(gclk));
	jdff dff_B_1DOt81Ad4_1(.din(w_dff_B_DpYNnzbp2_1),.dout(w_dff_B_1DOt81Ad4_1),.clk(gclk));
	jdff dff_B_sel0X8RR9_0(.din(n1602),.dout(w_dff_B_sel0X8RR9_0),.clk(gclk));
	jdff dff_A_FnpgA7eZ4_0(.dout(w_n558_0[0]),.din(w_dff_A_FnpgA7eZ4_0),.clk(gclk));
	jdff dff_A_Ng5qy9pI2_1(.dout(w_n558_0[1]),.din(w_dff_A_Ng5qy9pI2_1),.clk(gclk));
	jdff dff_A_kUyaWBU63_1(.dout(w_dff_A_Ng5qy9pI2_1),.din(w_dff_A_kUyaWBU63_1),.clk(gclk));
	jdff dff_A_lRVvlXKr1_1(.dout(w_dff_A_kUyaWBU63_1),.din(w_dff_A_lRVvlXKr1_1),.clk(gclk));
	jdff dff_A_4BSE3NL41_1(.dout(w_dff_A_lRVvlXKr1_1),.din(w_dff_A_4BSE3NL41_1),.clk(gclk));
	jdff dff_A_bHanTw4u7_1(.dout(w_dff_A_4BSE3NL41_1),.din(w_dff_A_bHanTw4u7_1),.clk(gclk));
	jdff dff_A_P3pamEE47_1(.dout(w_dff_A_bHanTw4u7_1),.din(w_dff_A_P3pamEE47_1),.clk(gclk));
	jdff dff_A_5E4wL1zE3_1(.dout(w_dff_A_P3pamEE47_1),.din(w_dff_A_5E4wL1zE3_1),.clk(gclk));
	jdff dff_A_XixEvbBh8_1(.dout(w_dff_A_5E4wL1zE3_1),.din(w_dff_A_XixEvbBh8_1),.clk(gclk));
	jdff dff_A_IynqEskC4_1(.dout(w_n1380_0[1]),.din(w_dff_A_IynqEskC4_1),.clk(gclk));
	jdff dff_A_0gA4mnx75_1(.dout(w_dff_A_IynqEskC4_1),.din(w_dff_A_0gA4mnx75_1),.clk(gclk));
	jdff dff_B_vi9gKCrh7_0(.din(n1377),.dout(w_dff_B_vi9gKCrh7_0),.clk(gclk));
	jdff dff_B_Pr4cRVXm5_0(.din(n1594),.dout(w_dff_B_Pr4cRVXm5_0),.clk(gclk));
	jdff dff_B_Eh2Rk16E7_0(.din(w_dff_B_Pr4cRVXm5_0),.dout(w_dff_B_Eh2Rk16E7_0),.clk(gclk));
	jdff dff_B_VkEavW1t2_0(.din(w_dff_B_Eh2Rk16E7_0),.dout(w_dff_B_VkEavW1t2_0),.clk(gclk));
	jdff dff_B_9ZpuAkHu2_0(.din(n1593),.dout(w_dff_B_9ZpuAkHu2_0),.clk(gclk));
	jdff dff_B_RjQZLPU06_0(.din(w_dff_B_9ZpuAkHu2_0),.dout(w_dff_B_RjQZLPU06_0),.clk(gclk));
	jdff dff_B_XX9PT8uf5_0(.din(w_dff_B_RjQZLPU06_0),.dout(w_dff_B_XX9PT8uf5_0),.clk(gclk));
	jdff dff_A_CMDxxD1q7_2(.dout(w_n1494_0[2]),.din(w_dff_A_CMDxxD1q7_2),.clk(gclk));
	jdff dff_A_CCfkFeBt8_2(.dout(w_dff_A_CMDxxD1q7_2),.din(w_dff_A_CCfkFeBt8_2),.clk(gclk));
	jdff dff_A_4GL5I2FX7_2(.dout(w_dff_A_CCfkFeBt8_2),.din(w_dff_A_4GL5I2FX7_2),.clk(gclk));
	jdff dff_A_9C6nb4KK7_2(.dout(w_dff_A_4GL5I2FX7_2),.din(w_dff_A_9C6nb4KK7_2),.clk(gclk));
	jdff dff_A_CHLv29ha1_2(.dout(w_dff_A_9C6nb4KK7_2),.din(w_dff_A_CHLv29ha1_2),.clk(gclk));
	jdff dff_A_27sUQoDV3_2(.dout(w_dff_A_CHLv29ha1_2),.din(w_dff_A_27sUQoDV3_2),.clk(gclk));
	jdff dff_A_I8542ZhQ6_2(.dout(w_dff_A_27sUQoDV3_2),.din(w_dff_A_I8542ZhQ6_2),.clk(gclk));
	jdff dff_A_IGyUEtNS0_2(.dout(w_dff_A_I8542ZhQ6_2),.din(w_dff_A_IGyUEtNS0_2),.clk(gclk));
	jdff dff_A_opi42OKV6_1(.dout(w_n524_1[1]),.din(w_dff_A_opi42OKV6_1),.clk(gclk));
	jdff dff_A_50Pk9rpa7_1(.dout(w_dff_A_opi42OKV6_1),.din(w_dff_A_50Pk9rpa7_1),.clk(gclk));
	jdff dff_A_h97gtSDy3_2(.dout(w_n524_1[2]),.din(w_dff_A_h97gtSDy3_2),.clk(gclk));
	jdff dff_A_KDwJqF2U7_2(.dout(w_dff_A_h97gtSDy3_2),.din(w_dff_A_KDwJqF2U7_2),.clk(gclk));
	jdff dff_A_nyalX7Vu4_2(.dout(w_dff_A_KDwJqF2U7_2),.din(w_dff_A_nyalX7Vu4_2),.clk(gclk));
	jdff dff_A_EJWBJjO24_2(.dout(w_dff_A_nyalX7Vu4_2),.din(w_dff_A_EJWBJjO24_2),.clk(gclk));
	jdff dff_A_kyC7fiAW9_2(.dout(w_dff_A_EJWBJjO24_2),.din(w_dff_A_kyC7fiAW9_2),.clk(gclk));
	jdff dff_A_gSCgWGLe3_2(.dout(w_dff_A_kyC7fiAW9_2),.din(w_dff_A_gSCgWGLe3_2),.clk(gclk));
	jdff dff_A_UasxrxzM1_2(.dout(w_dff_A_gSCgWGLe3_2),.din(w_dff_A_UasxrxzM1_2),.clk(gclk));
	jdff dff_A_3loQDpa12_2(.dout(w_dff_A_UasxrxzM1_2),.din(w_dff_A_3loQDpa12_2),.clk(gclk));
	jdff dff_A_tJTwwsdY4_2(.dout(w_dff_A_3loQDpa12_2),.din(w_dff_A_tJTwwsdY4_2),.clk(gclk));
	jdff dff_A_RAC4MjRG2_2(.dout(w_dff_A_tJTwwsdY4_2),.din(w_dff_A_RAC4MjRG2_2),.clk(gclk));
	jdff dff_A_ihl4IpdQ5_2(.dout(w_dff_A_RAC4MjRG2_2),.din(w_dff_A_ihl4IpdQ5_2),.clk(gclk));
	jdff dff_A_GMvBdxUO4_2(.dout(w_dff_A_ihl4IpdQ5_2),.din(w_dff_A_GMvBdxUO4_2),.clk(gclk));
	jdff dff_B_OIKxCJxU6_1(.din(n1588),.dout(w_dff_B_OIKxCJxU6_1),.clk(gclk));
	jdff dff_B_GJv8SWDd3_1(.din(w_dff_B_OIKxCJxU6_1),.dout(w_dff_B_GJv8SWDd3_1),.clk(gclk));
	jdff dff_B_xgc1Od2f3_1(.din(w_dff_B_GJv8SWDd3_1),.dout(w_dff_B_xgc1Od2f3_1),.clk(gclk));
	jdff dff_B_mm7fPUEe4_1(.din(w_dff_B_xgc1Od2f3_1),.dout(w_dff_B_mm7fPUEe4_1),.clk(gclk));
	jdff dff_B_2DsdV5O88_0(.din(n1590),.dout(w_dff_B_2DsdV5O88_0),.clk(gclk));
	jdff dff_A_x19YsS0i6_1(.dout(w_n549_0[1]),.din(w_dff_A_x19YsS0i6_1),.clk(gclk));
	jdff dff_B_SAlCeFYl0_2(.din(n549),.dout(w_dff_B_SAlCeFYl0_2),.clk(gclk));
	jdff dff_B_rFAGAFOx4_2(.din(w_dff_B_SAlCeFYl0_2),.dout(w_dff_B_rFAGAFOx4_2),.clk(gclk));
	jdff dff_A_fzKjvWig5_1(.dout(w_n556_0[1]),.din(w_dff_A_fzKjvWig5_1),.clk(gclk));
	jdff dff_A_HtvCpDy58_1(.dout(w_dff_A_fzKjvWig5_1),.din(w_dff_A_HtvCpDy58_1),.clk(gclk));
	jdff dff_A_Ns2WddQp2_1(.dout(w_dff_A_HtvCpDy58_1),.din(w_dff_A_Ns2WddQp2_1),.clk(gclk));
	jdff dff_A_s7orHyME7_1(.dout(w_dff_A_Ns2WddQp2_1),.din(w_dff_A_s7orHyME7_1),.clk(gclk));
	jdff dff_A_9BI1CyFY4_1(.dout(w_dff_A_s7orHyME7_1),.din(w_dff_A_9BI1CyFY4_1),.clk(gclk));
	jdff dff_A_sKP7S97R2_1(.dout(w_dff_A_9BI1CyFY4_1),.din(w_dff_A_sKP7S97R2_1),.clk(gclk));
	jdff dff_A_7MI3tEFm7_1(.dout(w_dff_A_sKP7S97R2_1),.din(w_dff_A_7MI3tEFm7_1),.clk(gclk));
	jdff dff_A_lwZauxQ99_1(.dout(w_dff_A_7MI3tEFm7_1),.din(w_dff_A_lwZauxQ99_1),.clk(gclk));
	jdff dff_A_W9Oe9Irk5_1(.dout(w_dff_A_lwZauxQ99_1),.din(w_dff_A_W9Oe9Irk5_1),.clk(gclk));
	jdff dff_A_nCU9MRR05_1(.dout(w_n554_0[1]),.din(w_dff_A_nCU9MRR05_1),.clk(gclk));
	jdff dff_A_hHJMPfl68_1(.dout(w_dff_A_nCU9MRR05_1),.din(w_dff_A_hHJMPfl68_1),.clk(gclk));
	jdff dff_A_UqO1TnTV9_1(.dout(w_dff_A_hHJMPfl68_1),.din(w_dff_A_UqO1TnTV9_1),.clk(gclk));
	jdff dff_A_iGjyd2mM3_1(.dout(w_dff_A_UqO1TnTV9_1),.din(w_dff_A_iGjyd2mM3_1),.clk(gclk));
	jdff dff_A_fNXRIG3F4_1(.dout(w_dff_A_iGjyd2mM3_1),.din(w_dff_A_fNXRIG3F4_1),.clk(gclk));
	jdff dff_A_6qYis3IZ4_1(.dout(w_dff_A_fNXRIG3F4_1),.din(w_dff_A_6qYis3IZ4_1),.clk(gclk));
	jdff dff_A_GIqro3PQ5_1(.dout(w_dff_A_6qYis3IZ4_1),.din(w_dff_A_GIqro3PQ5_1),.clk(gclk));
	jdff dff_A_pvqZuXdk9_1(.dout(w_dff_A_GIqro3PQ5_1),.din(w_dff_A_pvqZuXdk9_1),.clk(gclk));
	jdff dff_A_TcSk9PEH7_1(.dout(w_dff_A_pvqZuXdk9_1),.din(w_dff_A_TcSk9PEH7_1),.clk(gclk));
	jdff dff_A_fIfmGo6g3_1(.dout(w_dff_A_TcSk9PEH7_1),.din(w_dff_A_fIfmGo6g3_1),.clk(gclk));
	jdff dff_A_ck0iszft9_1(.dout(w_dff_A_fIfmGo6g3_1),.din(w_dff_A_ck0iszft9_1),.clk(gclk));
	jdff dff_B_PcBIj1gP7_1(.din(n526),.dout(w_dff_B_PcBIj1gP7_1),.clk(gclk));
	jdff dff_B_4FoRgvuD6_0(.din(G35),.dout(w_dff_B_4FoRgvuD6_0),.clk(gclk));
	jdff dff_A_AqZSHEOy8_1(.dout(w_n525_0[1]),.din(w_dff_A_AqZSHEOy8_1),.clk(gclk));
	jdff dff_A_4E7K3r0y5_1(.dout(w_dff_A_AqZSHEOy8_1),.din(w_dff_A_4E7K3r0y5_1),.clk(gclk));
	jdff dff_A_EiVtXFOz7_2(.dout(w_n525_0[2]),.din(w_dff_A_EiVtXFOz7_2),.clk(gclk));
	jdff dff_A_JIK2jnnq1_2(.dout(w_dff_A_EiVtXFOz7_2),.din(w_dff_A_JIK2jnnq1_2),.clk(gclk));
	jdff dff_A_lAvt5qLZ3_1(.dout(w_G4420_0[1]),.din(w_dff_A_lAvt5qLZ3_1),.clk(gclk));
	jdff dff_A_KCyLF0xG5_1(.dout(w_dff_A_lAvt5qLZ3_1),.din(w_dff_A_KCyLF0xG5_1),.clk(gclk));
	jdff dff_A_3jSymNVW0_1(.dout(w_dff_A_KCyLF0xG5_1),.din(w_dff_A_3jSymNVW0_1),.clk(gclk));
	jdff dff_A_8eBzixrq7_1(.dout(w_dff_A_3jSymNVW0_1),.din(w_dff_A_8eBzixrq7_1),.clk(gclk));
	jdff dff_A_DgDAJlvf3_2(.dout(w_n524_0[2]),.din(w_dff_A_DgDAJlvf3_2),.clk(gclk));
	jdff dff_A_Iuxr2gKJ8_2(.dout(w_dff_A_DgDAJlvf3_2),.din(w_dff_A_Iuxr2gKJ8_2),.clk(gclk));
	jdff dff_A_pE32UJ6Y0_0(.dout(w_n553_0[0]),.din(w_dff_A_pE32UJ6Y0_0),.clk(gclk));
	jdff dff_A_5dgnjyY68_0(.dout(w_dff_A_pE32UJ6Y0_0),.din(w_dff_A_5dgnjyY68_0),.clk(gclk));
	jdff dff_B_JGSCKHOj3_2(.din(n553),.dout(w_dff_B_JGSCKHOj3_2),.clk(gclk));
	jdff dff_B_fzUH6Gwg3_1(.din(n521),.dout(w_dff_B_fzUH6Gwg3_1),.clk(gclk));
	jdff dff_B_AJSqunPQ4_0(.din(G32),.dout(w_dff_B_AJSqunPQ4_0),.clk(gclk));
	jdff dff_A_EhA8q3zh6_1(.dout(w_n520_0[1]),.din(w_dff_A_EhA8q3zh6_1),.clk(gclk));
	jdff dff_A_rPxpNk2v5_1(.dout(w_dff_A_EhA8q3zh6_1),.din(w_dff_A_rPxpNk2v5_1),.clk(gclk));
	jdff dff_A_6cgcbzJM4_2(.dout(w_n520_0[2]),.din(w_dff_A_6cgcbzJM4_2),.clk(gclk));
	jdff dff_A_t8sJnWpR2_2(.dout(w_dff_A_6cgcbzJM4_2),.din(w_dff_A_t8sJnWpR2_2),.clk(gclk));
	jdff dff_A_fDzA0mv00_0(.dout(w_n552_0[0]),.din(w_dff_A_fDzA0mv00_0),.clk(gclk));
	jdff dff_A_o5zNdw3o6_0(.dout(w_dff_A_fDzA0mv00_0),.din(w_dff_A_o5zNdw3o6_0),.clk(gclk));
	jdff dff_A_Q9lzvkjn7_0(.dout(w_dff_A_o5zNdw3o6_0),.din(w_dff_A_Q9lzvkjn7_0),.clk(gclk));
	jdff dff_A_gCT6V1oP9_0(.dout(w_dff_A_Q9lzvkjn7_0),.din(w_dff_A_gCT6V1oP9_0),.clk(gclk));
	jdff dff_A_o1KJXdOF0_0(.dout(w_dff_A_gCT6V1oP9_0),.din(w_dff_A_o1KJXdOF0_0),.clk(gclk));
	jdff dff_A_DSPztC9M3_0(.dout(w_dff_A_o1KJXdOF0_0),.din(w_dff_A_DSPztC9M3_0),.clk(gclk));
	jdff dff_A_4Jyj9n3U1_0(.dout(w_dff_A_DSPztC9M3_0),.din(w_dff_A_4Jyj9n3U1_0),.clk(gclk));
	jdff dff_A_v7Y8xzsW1_0(.dout(w_dff_A_4Jyj9n3U1_0),.din(w_dff_A_v7Y8xzsW1_0),.clk(gclk));
	jdff dff_A_EZo0lXF13_0(.dout(w_dff_A_v7Y8xzsW1_0),.din(w_dff_A_EZo0lXF13_0),.clk(gclk));
	jdff dff_A_wUx0yTa09_0(.dout(w_n551_0[0]),.din(w_dff_A_wUx0yTa09_0),.clk(gclk));
	jdff dff_A_UzABrpJR6_0(.dout(w_dff_A_wUx0yTa09_0),.din(w_dff_A_UzABrpJR6_0),.clk(gclk));
	jdff dff_A_EYlpZPJq4_0(.dout(w_dff_A_UzABrpJR6_0),.din(w_dff_A_EYlpZPJq4_0),.clk(gclk));
	jdff dff_A_egm8n0ej7_1(.dout(w_n535_0[1]),.din(w_dff_A_egm8n0ej7_1),.clk(gclk));
	jdff dff_B_yAKEZt6k3_1(.din(n532),.dout(w_dff_B_yAKEZt6k3_1),.clk(gclk));
	jdff dff_B_84iRtvq86_0(.din(G66),.dout(w_dff_B_84iRtvq86_0),.clk(gclk));
	jdff dff_A_0iBeJp9B8_1(.dout(w_n531_0[1]),.din(w_dff_A_0iBeJp9B8_1),.clk(gclk));
	jdff dff_A_T9rOa2NS6_1(.dout(w_dff_A_0iBeJp9B8_1),.din(w_dff_A_T9rOa2NS6_1),.clk(gclk));
	jdff dff_A_6gtT0VQr7_2(.dout(w_n531_0[2]),.din(w_dff_A_6gtT0VQr7_2),.clk(gclk));
	jdff dff_A_bcAtzUew4_2(.dout(w_dff_A_6gtT0VQr7_2),.din(w_dff_A_bcAtzUew4_2),.clk(gclk));
	jdff dff_A_XB3GkqvB2_1(.dout(w_G4437_0[1]),.din(w_dff_A_XB3GkqvB2_1),.clk(gclk));
	jdff dff_A_r1Eae4on4_1(.dout(w_dff_A_XB3GkqvB2_1),.din(w_dff_A_r1Eae4on4_1),.clk(gclk));
	jdff dff_A_BKMaKKir6_1(.dout(w_dff_A_r1Eae4on4_1),.din(w_dff_A_BKMaKKir6_1),.clk(gclk));
	jdff dff_A_VgHUHFeN3_1(.dout(w_dff_A_BKMaKKir6_1),.din(w_dff_A_VgHUHFeN3_1),.clk(gclk));
	jdff dff_A_5nLHnB6C4_1(.dout(w_n518_0[1]),.din(w_dff_A_5nLHnB6C4_1),.clk(gclk));
	jdff dff_B_nM3yZrsY8_1(.din(n498),.dout(w_dff_B_nM3yZrsY8_1),.clk(gclk));
	jdff dff_B_lUP2YVfW1_1(.din(w_dff_B_nM3yZrsY8_1),.dout(w_dff_B_lUP2YVfW1_1),.clk(gclk));
	jdff dff_B_B0NN0BAE9_1(.din(w_dff_B_lUP2YVfW1_1),.dout(w_dff_B_B0NN0BAE9_1),.clk(gclk));
	jdff dff_B_FX4kO5pn5_1(.din(w_dff_B_B0NN0BAE9_1),.dout(w_dff_B_FX4kO5pn5_1),.clk(gclk));
	jdff dff_B_G3a7yDBn7_1(.din(w_dff_B_FX4kO5pn5_1),.dout(w_dff_B_G3a7yDBn7_1),.clk(gclk));
	jdff dff_B_ReywKQIc6_1(.din(w_dff_B_G3a7yDBn7_1),.dout(w_dff_B_ReywKQIc6_1),.clk(gclk));
	jdff dff_B_4c1rMKSY1_1(.din(n500),.dout(w_dff_B_4c1rMKSY1_1),.clk(gclk));
	jdff dff_B_kVQlZe7Y6_1(.din(w_dff_B_4c1rMKSY1_1),.dout(w_dff_B_kVQlZe7Y6_1),.clk(gclk));
	jdff dff_B_VV4ipEa63_1(.din(w_dff_B_kVQlZe7Y6_1),.dout(w_dff_B_VV4ipEa63_1),.clk(gclk));
	jdff dff_B_NU9PT9Tc7_1(.din(w_dff_B_VV4ipEa63_1),.dout(w_dff_B_NU9PT9Tc7_1),.clk(gclk));
	jdff dff_B_7bPW3G278_1(.din(w_dff_B_NU9PT9Tc7_1),.dout(w_dff_B_7bPW3G278_1),.clk(gclk));
	jdff dff_A_u77RTt2G0_1(.dout(w_n516_0[1]),.din(w_dff_A_u77RTt2G0_1),.clk(gclk));
	jdff dff_A_qgFMoNKm5_1(.dout(w_dff_A_u77RTt2G0_1),.din(w_dff_A_qgFMoNKm5_1),.clk(gclk));
	jdff dff_A_XTAzeNi84_1(.dout(w_dff_A_qgFMoNKm5_1),.din(w_dff_A_XTAzeNi84_1),.clk(gclk));
	jdff dff_A_0LzmGCC08_1(.dout(w_dff_A_XTAzeNi84_1),.din(w_dff_A_0LzmGCC08_1),.clk(gclk));
	jdff dff_A_5qzCAV2S8_1(.dout(w_dff_A_0LzmGCC08_1),.din(w_dff_A_5qzCAV2S8_1),.clk(gclk));
	jdff dff_B_uW98lKMF6_1(.din(n504),.dout(w_dff_B_uW98lKMF6_1),.clk(gclk));
	jdff dff_B_wJZHFkYc5_1(.din(w_dff_B_uW98lKMF6_1),.dout(w_dff_B_wJZHFkYc5_1),.clk(gclk));
	jdff dff_B_RSpnqIE92_1(.din(w_dff_B_wJZHFkYc5_1),.dout(w_dff_B_RSpnqIE92_1),.clk(gclk));
	jdff dff_A_GsSCDuzU2_1(.dout(w_n514_0[1]),.din(w_dff_A_GsSCDuzU2_1),.clk(gclk));
	jdff dff_A_Lh6XoaEJ7_1(.dout(w_dff_A_GsSCDuzU2_1),.din(w_dff_A_Lh6XoaEJ7_1),.clk(gclk));
	jdff dff_A_vznTILIU3_1(.dout(w_dff_A_Lh6XoaEJ7_1),.din(w_dff_A_vznTILIU3_1),.clk(gclk));
	jdff dff_A_DMkJGa9p8_1(.dout(w_dff_A_vznTILIU3_1),.din(w_dff_A_DMkJGa9p8_1),.clk(gclk));
	jdff dff_A_xvBOGYZI5_1(.dout(w_dff_A_DMkJGa9p8_1),.din(w_dff_A_xvBOGYZI5_1),.clk(gclk));
	jdff dff_A_pH4My2IA7_1(.dout(w_dff_A_xvBOGYZI5_1),.din(w_dff_A_pH4My2IA7_1),.clk(gclk));
	jdff dff_A_NdcOEkCb6_0(.dout(w_n512_0[0]),.din(w_dff_A_NdcOEkCb6_0),.clk(gclk));
	jdff dff_A_6U1UqLW16_0(.dout(w_n510_0[0]),.din(w_dff_A_6U1UqLW16_0),.clk(gclk));
	jdff dff_A_xxOlJ3CW8_0(.dout(w_n509_0[0]),.din(w_dff_A_xxOlJ3CW8_0),.clk(gclk));
	jdff dff_A_U0hXA5h91_0(.dout(w_dff_A_xxOlJ3CW8_0),.din(w_dff_A_U0hXA5h91_0),.clk(gclk));
	jdff dff_A_JE9mLRAe8_2(.dout(w_n507_0[2]),.din(w_dff_A_JE9mLRAe8_2),.clk(gclk));
	jdff dff_A_YOXyXLCP3_2(.dout(w_dff_A_JE9mLRAe8_2),.din(w_dff_A_YOXyXLCP3_2),.clk(gclk));
	jdff dff_A_QXQ9j92N2_2(.dout(w_dff_A_YOXyXLCP3_2),.din(w_dff_A_QXQ9j92N2_2),.clk(gclk));
	jdff dff_A_zIdw6yhx1_2(.dout(w_dff_A_QXQ9j92N2_2),.din(w_dff_A_zIdw6yhx1_2),.clk(gclk));
	jdff dff_A_L8v9zKPK0_1(.dout(w_n505_0[1]),.din(w_dff_A_L8v9zKPK0_1),.clk(gclk));
	jdff dff_B_BpLrxlZp9_2(.din(n505),.dout(w_dff_B_BpLrxlZp9_2),.clk(gclk));
	jdff dff_A_zzibIUZP2_0(.dout(w_n503_0[0]),.din(w_dff_A_zzibIUZP2_0),.clk(gclk));
	jdff dff_A_WeQLK4OR9_0(.dout(w_n502_0[0]),.din(w_dff_A_WeQLK4OR9_0),.clk(gclk));
	jdff dff_B_KV71pfwJ2_2(.din(n502),.dout(w_dff_B_KV71pfwJ2_2),.clk(gclk));
	jdff dff_B_pMrX8p496_2(.din(w_dff_B_KV71pfwJ2_2),.dout(w_dff_B_pMrX8p496_2),.clk(gclk));
	jdff dff_B_EYruc3vf3_2(.din(w_dff_B_pMrX8p496_2),.dout(w_dff_B_EYruc3vf3_2),.clk(gclk));
	jdff dff_B_Kmrt3sfJ7_2(.din(w_dff_B_EYruc3vf3_2),.dout(w_dff_B_Kmrt3sfJ7_2),.clk(gclk));
	jdff dff_B_VVfKKsny1_0(.din(n495),.dout(w_dff_B_VVfKKsny1_0),.clk(gclk));
	jdff dff_B_vqSnrWII8_0(.din(w_dff_B_VVfKKsny1_0),.dout(w_dff_B_vqSnrWII8_0),.clk(gclk));
	jdff dff_B_2GNWMdUI1_0(.din(w_dff_B_vqSnrWII8_0),.dout(w_dff_B_2GNWMdUI1_0),.clk(gclk));
	jdff dff_A_u1xDV8Vf1_0(.dout(w_n494_0[0]),.din(w_dff_A_u1xDV8Vf1_0),.clk(gclk));
	jdff dff_A_iRiUx5rP2_0(.dout(w_dff_A_u1xDV8Vf1_0),.din(w_dff_A_iRiUx5rP2_0),.clk(gclk));
	jdff dff_A_0siaQzSh6_0(.dout(w_dff_A_iRiUx5rP2_0),.din(w_dff_A_0siaQzSh6_0),.clk(gclk));
	jdff dff_A_tOfU8hJU1_0(.dout(w_dff_A_0siaQzSh6_0),.din(w_dff_A_tOfU8hJU1_0),.clk(gclk));
	jdff dff_A_6t7b2Fct8_0(.dout(w_n493_0[0]),.din(w_dff_A_6t7b2Fct8_0),.clk(gclk));
	jdff dff_A_5pYyDCjl1_0(.dout(w_dff_A_6t7b2Fct8_0),.din(w_dff_A_5pYyDCjl1_0),.clk(gclk));
	jdff dff_A_F5L11Xlj2_0(.dout(w_dff_A_5pYyDCjl1_0),.din(w_dff_A_F5L11Xlj2_0),.clk(gclk));
	jdff dff_A_ajUlbdyL5_0(.dout(w_dff_A_F5L11Xlj2_0),.din(w_dff_A_ajUlbdyL5_0),.clk(gclk));
	jdff dff_A_ldFYse3U6_0(.dout(w_n480_1[0]),.din(w_dff_A_ldFYse3U6_0),.clk(gclk));
	jdff dff_A_8uUtDvTF5_0(.dout(w_dff_A_ldFYse3U6_0),.din(w_dff_A_8uUtDvTF5_0),.clk(gclk));
	jdff dff_A_tTHkCHta4_0(.dout(w_dff_A_8uUtDvTF5_0),.din(w_dff_A_tTHkCHta4_0),.clk(gclk));
	jdff dff_A_kwfy8KXb7_0(.dout(w_dff_A_tTHkCHta4_0),.din(w_dff_A_kwfy8KXb7_0),.clk(gclk));
	jdff dff_A_kqH5AU9u5_0(.dout(w_dff_A_kwfy8KXb7_0),.din(w_dff_A_kqH5AU9u5_0),.clk(gclk));
	jdff dff_A_qEgsXavU1_0(.dout(w_dff_A_kqH5AU9u5_0),.din(w_dff_A_qEgsXavU1_0),.clk(gclk));
	jdff dff_A_PXkeGuLe9_0(.dout(w_dff_A_qEgsXavU1_0),.din(w_dff_A_PXkeGuLe9_0),.clk(gclk));
	jdff dff_A_fdpewNTe8_1(.dout(w_n480_0[1]),.din(w_dff_A_fdpewNTe8_1),.clk(gclk));
	jdff dff_A_WvhCOYmd0_1(.dout(w_dff_A_fdpewNTe8_1),.din(w_dff_A_WvhCOYmd0_1),.clk(gclk));
	jdff dff_A_tVXKqJGB9_1(.dout(w_dff_A_WvhCOYmd0_1),.din(w_dff_A_tVXKqJGB9_1),.clk(gclk));
	jdff dff_A_EP0sGnie1_2(.dout(w_n480_0[2]),.din(w_dff_A_EP0sGnie1_2),.clk(gclk));
	jdff dff_A_hKmYyrgv9_2(.dout(w_dff_A_EP0sGnie1_2),.din(w_dff_A_hKmYyrgv9_2),.clk(gclk));
	jdff dff_A_p77vMcCr0_2(.dout(w_dff_A_hKmYyrgv9_2),.din(w_dff_A_p77vMcCr0_2),.clk(gclk));
	jdff dff_A_ojFg92OK0_2(.dout(w_dff_A_p77vMcCr0_2),.din(w_dff_A_ojFg92OK0_2),.clk(gclk));
	jdff dff_A_VvOpbdxn0_2(.dout(w_dff_A_ojFg92OK0_2),.din(w_dff_A_VvOpbdxn0_2),.clk(gclk));
	jdff dff_A_ENMNb7XV9_2(.dout(w_dff_A_VvOpbdxn0_2),.din(w_dff_A_ENMNb7XV9_2),.clk(gclk));
	jdff dff_A_NwdEVlzB8_2(.dout(w_dff_A_ENMNb7XV9_2),.din(w_dff_A_NwdEVlzB8_2),.clk(gclk));
	jdff dff_B_I7HteV6h8_1(.din(n476),.dout(w_dff_B_I7HteV6h8_1),.clk(gclk));
	jdff dff_B_EYX6X5V06_0(.din(G118),.dout(w_dff_B_EYX6X5V06_0),.clk(gclk));
	jdff dff_A_TDelmwbm7_0(.dout(w_G4394_0[0]),.din(w_dff_A_TDelmwbm7_0),.clk(gclk));
	jdff dff_A_okpQ7hcA6_0(.dout(w_dff_A_TDelmwbm7_0),.din(w_dff_A_okpQ7hcA6_0),.clk(gclk));
	jdff dff_A_o0jEiWOW7_0(.dout(w_dff_A_okpQ7hcA6_0),.din(w_dff_A_o0jEiWOW7_0),.clk(gclk));
	jdff dff_A_F6zSoCrM3_0(.dout(w_dff_A_o0jEiWOW7_0),.din(w_dff_A_F6zSoCrM3_0),.clk(gclk));
	jdff dff_A_UMlRGQE61_1(.dout(w_n475_1[1]),.din(w_dff_A_UMlRGQE61_1),.clk(gclk));
	jdff dff_A_Ar2t3l8F8_1(.dout(w_n475_0[1]),.din(w_dff_A_Ar2t3l8F8_1),.clk(gclk));
	jdff dff_A_ZtNUuRnv6_2(.dout(w_n475_0[2]),.din(w_dff_A_ZtNUuRnv6_2),.clk(gclk));
	jdff dff_A_3o7m0Os36_2(.dout(w_dff_A_ZtNUuRnv6_2),.din(w_dff_A_3o7m0Os36_2),.clk(gclk));
	jdff dff_A_k7JJI3cr8_2(.dout(w_dff_A_3o7m0Os36_2),.din(w_dff_A_k7JJI3cr8_2),.clk(gclk));
	jdff dff_A_atQfae210_2(.dout(w_dff_A_k7JJI3cr8_2),.din(w_dff_A_atQfae210_2),.clk(gclk));
	jdff dff_A_1iOGvwmI5_2(.dout(w_dff_A_atQfae210_2),.din(w_dff_A_1iOGvwmI5_2),.clk(gclk));
	jdff dff_A_sdAdEEBW6_2(.dout(w_dff_A_1iOGvwmI5_2),.din(w_dff_A_sdAdEEBW6_2),.clk(gclk));
	jdff dff_A_gk9VVL3Z7_2(.dout(w_dff_A_sdAdEEBW6_2),.din(w_dff_A_gk9VVL3Z7_2),.clk(gclk));
	jdff dff_A_CUvmDf5J0_2(.dout(w_dff_A_gk9VVL3Z7_2),.din(w_dff_A_CUvmDf5J0_2),.clk(gclk));
	jdff dff_A_abvw01o64_2(.dout(w_dff_A_CUvmDf5J0_2),.din(w_dff_A_abvw01o64_2),.clk(gclk));
	jdff dff_A_KGEqSJ7R2_2(.dout(w_dff_A_abvw01o64_2),.din(w_dff_A_KGEqSJ7R2_2),.clk(gclk));
	jdff dff_B_QMTRnMAr5_1(.din(n472),.dout(w_dff_B_QMTRnMAr5_1),.clk(gclk));
	jdff dff_B_Y2u8jKVw1_0(.din(G97),.dout(w_dff_B_Y2u8jKVw1_0),.clk(gclk));
	jdff dff_B_T69QBFzD0_3(.din(n471),.dout(w_dff_B_T69QBFzD0_3),.clk(gclk));
	jdff dff_B_QCLCXMcC4_3(.din(w_dff_B_T69QBFzD0_3),.dout(w_dff_B_QCLCXMcC4_3),.clk(gclk));
	jdff dff_A_TnqZL3N03_0(.dout(w_n470_0[0]),.din(w_dff_A_TnqZL3N03_0),.clk(gclk));
	jdff dff_A_3WBdhEWs9_0(.dout(w_dff_A_TnqZL3N03_0),.din(w_dff_A_3WBdhEWs9_0),.clk(gclk));
	jdff dff_A_vmr5aENK6_0(.dout(w_dff_A_3WBdhEWs9_0),.din(w_dff_A_vmr5aENK6_0),.clk(gclk));
	jdff dff_A_R0cohlg94_0(.dout(w_dff_A_vmr5aENK6_0),.din(w_dff_A_R0cohlg94_0),.clk(gclk));
	jdff dff_A_azehETn11_2(.dout(w_n470_0[2]),.din(w_dff_A_azehETn11_2),.clk(gclk));
	jdff dff_A_sclD5zdd4_2(.dout(w_dff_A_azehETn11_2),.din(w_dff_A_sclD5zdd4_2),.clk(gclk));
	jdff dff_A_Iu8Av3AH3_2(.dout(w_dff_A_sclD5zdd4_2),.din(w_dff_A_Iu8Av3AH3_2),.clk(gclk));
	jdff dff_B_wSeJvHvY2_1(.din(n467),.dout(w_dff_B_wSeJvHvY2_1),.clk(gclk));
	jdff dff_B_Bzm4aaA47_0(.din(G47),.dout(w_dff_B_Bzm4aaA47_0),.clk(gclk));
	jdff dff_B_G4bOJIy79_2(.din(n466),.dout(w_dff_B_G4bOJIy79_2),.clk(gclk));
	jdff dff_B_jr5IL4iN8_2(.din(w_dff_B_G4bOJIy79_2),.dout(w_dff_B_jr5IL4iN8_2),.clk(gclk));
	jdff dff_A_yoOFCVWY1_0(.dout(w_G4415_1[0]),.din(w_dff_A_yoOFCVWY1_0),.clk(gclk));
	jdff dff_A_1ETaXjQF7_0(.dout(w_dff_A_yoOFCVWY1_0),.din(w_dff_A_1ETaXjQF7_0),.clk(gclk));
	jdff dff_A_70SR8ZAK3_0(.dout(w_dff_A_1ETaXjQF7_0),.din(w_dff_A_70SR8ZAK3_0),.clk(gclk));
	jdff dff_A_YppMUfdg6_0(.dout(w_dff_A_70SR8ZAK3_0),.din(w_dff_A_YppMUfdg6_0),.clk(gclk));
	jdff dff_A_4OlQz9K68_0(.dout(w_n465_0[0]),.din(w_dff_A_4OlQz9K68_0),.clk(gclk));
	jdff dff_A_o4THdZ0n0_0(.dout(w_dff_A_4OlQz9K68_0),.din(w_dff_A_o4THdZ0n0_0),.clk(gclk));
	jdff dff_A_plzDQIpw4_0(.dout(w_dff_A_o4THdZ0n0_0),.din(w_dff_A_plzDQIpw4_0),.clk(gclk));
	jdff dff_A_b5VbxXny3_0(.dout(w_dff_A_plzDQIpw4_0),.din(w_dff_A_b5VbxXny3_0),.clk(gclk));
	jdff dff_A_GO7S0n6C9_1(.dout(w_n464_0[1]),.din(w_dff_A_GO7S0n6C9_1),.clk(gclk));
	jdff dff_A_sqp9Njm17_1(.dout(w_n452_0[1]),.din(w_dff_A_sqp9Njm17_1),.clk(gclk));
	jdff dff_A_ayvScaaT2_1(.dout(w_dff_A_sqp9Njm17_1),.din(w_dff_A_ayvScaaT2_1),.clk(gclk));
	jdff dff_A_dfPLcqln1_0(.dout(w_n446_1[0]),.din(w_dff_A_dfPLcqln1_0),.clk(gclk));
	jdff dff_A_kXBd5JXl6_0(.dout(w_dff_A_dfPLcqln1_0),.din(w_dff_A_kXBd5JXl6_0),.clk(gclk));
	jdff dff_A_mjnJcMV75_0(.dout(w_dff_A_kXBd5JXl6_0),.din(w_dff_A_mjnJcMV75_0),.clk(gclk));
	jdff dff_A_ttlRrIgr0_0(.dout(w_dff_A_mjnJcMV75_0),.din(w_dff_A_ttlRrIgr0_0),.clk(gclk));
	jdff dff_A_0szJyxE99_0(.dout(w_dff_A_ttlRrIgr0_0),.din(w_dff_A_0szJyxE99_0),.clk(gclk));
	jdff dff_A_WJQMmuie9_0(.dout(w_dff_A_0szJyxE99_0),.din(w_dff_A_WJQMmuie9_0),.clk(gclk));
	jdff dff_A_NBaBoVcZ7_0(.dout(w_dff_A_WJQMmuie9_0),.din(w_dff_A_NBaBoVcZ7_0),.clk(gclk));
	jdff dff_A_IiN5JI5s8_0(.dout(w_n437_0[0]),.din(w_dff_A_IiN5JI5s8_0),.clk(gclk));
	jdff dff_A_W5tLDX4L7_0(.dout(w_dff_A_IiN5JI5s8_0),.din(w_dff_A_W5tLDX4L7_0),.clk(gclk));
	jdff dff_A_7zf17ZJ46_0(.dout(w_dff_A_W5tLDX4L7_0),.din(w_dff_A_7zf17ZJ46_0),.clk(gclk));
	jdff dff_B_XJUEGaX61_2(.din(n437),.dout(w_dff_B_XJUEGaX61_2),.clk(gclk));
	jdff dff_B_cteXpGLd6_2(.din(w_dff_B_XJUEGaX61_2),.dout(w_dff_B_cteXpGLd6_2),.clk(gclk));
	jdff dff_A_rYZP6bhc0_0(.dout(w_n436_0[0]),.din(w_dff_A_rYZP6bhc0_0),.clk(gclk));
	jdff dff_A_lXbV1seQ8_0(.dout(w_dff_A_rYZP6bhc0_0),.din(w_dff_A_lXbV1seQ8_0),.clk(gclk));
	jdff dff_A_OloIHzAR1_0(.dout(w_dff_A_lXbV1seQ8_0),.din(w_dff_A_OloIHzAR1_0),.clk(gclk));
	jdff dff_A_T2HkbbHv0_0(.dout(w_dff_A_OloIHzAR1_0),.din(w_dff_A_T2HkbbHv0_0),.clk(gclk));
	jdff dff_A_GTbnRU559_0(.dout(w_dff_A_T2HkbbHv0_0),.din(w_dff_A_GTbnRU559_0),.clk(gclk));
	jdff dff_A_mtPxmBZR7_0(.dout(w_dff_A_GTbnRU559_0),.din(w_dff_A_mtPxmBZR7_0),.clk(gclk));
	jdff dff_A_p7UtFTKd6_1(.dout(w_n430_0[1]),.din(w_dff_A_p7UtFTKd6_1),.clk(gclk));
	jdff dff_A_zUKcF8oA4_1(.dout(w_dff_A_p7UtFTKd6_1),.din(w_dff_A_zUKcF8oA4_1),.clk(gclk));
	jdff dff_A_IxiQpLBq7_1(.dout(w_n491_0[1]),.din(w_dff_A_IxiQpLBq7_1),.clk(gclk));
	jdff dff_B_5hU4vHiZ8_1(.din(n487),.dout(w_dff_B_5hU4vHiZ8_1),.clk(gclk));
	jdff dff_B_0QEtDJod2_0(.din(G94),.dout(w_dff_B_0QEtDJod2_0),.clk(gclk));
	jdff dff_A_bIhfmbo90_0(.dout(w_G4405_0[0]),.din(w_dff_A_bIhfmbo90_0),.clk(gclk));
	jdff dff_A_mdiprYfS9_0(.dout(w_dff_A_bIhfmbo90_0),.din(w_dff_A_mdiprYfS9_0),.clk(gclk));
	jdff dff_A_mb7C1QHa8_0(.dout(w_dff_A_mdiprYfS9_0),.din(w_dff_A_mb7C1QHa8_0),.clk(gclk));
	jdff dff_A_J2qPaUXQ6_0(.dout(w_dff_A_mb7C1QHa8_0),.din(w_dff_A_J2qPaUXQ6_0),.clk(gclk));
	jdff dff_A_xdlzvDjW9_0(.dout(w_n486_0[0]),.din(w_dff_A_xdlzvDjW9_0),.clk(gclk));
	jdff dff_A_x71sLdCq3_2(.dout(w_n486_0[2]),.din(w_dff_A_x71sLdCq3_2),.clk(gclk));
	jdff dff_B_JjtPmCHB3_1(.din(n483),.dout(w_dff_B_JjtPmCHB3_1),.clk(gclk));
	jdff dff_B_r7ZZahyA5_0(.din(G121),.dout(w_dff_B_r7ZZahyA5_0),.clk(gclk));
	jdff dff_B_vh3Uguei7_2(.din(n482),.dout(w_dff_B_vh3Uguei7_2),.clk(gclk));
	jdff dff_B_2P58I5eT7_2(.din(w_dff_B_vh3Uguei7_2),.dout(w_dff_B_2P58I5eT7_2),.clk(gclk));
	jdff dff_A_vIvxKYgN7_0(.dout(w_G4410_1[0]),.din(w_dff_A_vIvxKYgN7_0),.clk(gclk));
	jdff dff_A_U9HEbJgo5_0(.dout(w_dff_A_vIvxKYgN7_0),.din(w_dff_A_U9HEbJgo5_0),.clk(gclk));
	jdff dff_A_K48xyCr10_0(.dout(w_dff_A_U9HEbJgo5_0),.din(w_dff_A_K48xyCr10_0),.clk(gclk));
	jdff dff_A_6pxG1Fq52_0(.dout(w_dff_A_K48xyCr10_0),.din(w_dff_A_6pxG1Fq52_0),.clk(gclk));
	jdff dff_A_5EbDisAo9_0(.dout(w_n540_0[0]),.din(w_dff_A_5EbDisAo9_0),.clk(gclk));
	jdff dff_A_IlnJLqiF5_0(.dout(w_dff_A_5EbDisAo9_0),.din(w_dff_A_IlnJLqiF5_0),.clk(gclk));
	jdff dff_A_TzbzIG4M8_1(.dout(w_n540_0[1]),.din(w_dff_A_TzbzIG4M8_1),.clk(gclk));
	jdff dff_A_9LNjiWNT4_1(.dout(w_dff_A_TzbzIG4M8_1),.din(w_dff_A_9LNjiWNT4_1),.clk(gclk));
	jdff dff_A_TO5rHO6z6_1(.dout(w_dff_A_9LNjiWNT4_1),.din(w_dff_A_TO5rHO6z6_1),.clk(gclk));
	jdff dff_A_xb40rgLK8_1(.dout(w_dff_A_TO5rHO6z6_1),.din(w_dff_A_xb40rgLK8_1),.clk(gclk));
	jdff dff_A_3bsSzGkA5_1(.dout(w_dff_A_xb40rgLK8_1),.din(w_dff_A_3bsSzGkA5_1),.clk(gclk));
	jdff dff_A_OL3a0SAZ9_1(.dout(w_dff_A_3bsSzGkA5_1),.din(w_dff_A_OL3a0SAZ9_1),.clk(gclk));
	jdff dff_A_LqKGtasU1_1(.dout(w_dff_A_OL3a0SAZ9_1),.din(w_dff_A_LqKGtasU1_1),.clk(gclk));
	jdff dff_A_NdTm2IRH8_1(.dout(w_dff_A_LqKGtasU1_1),.din(w_dff_A_NdTm2IRH8_1),.clk(gclk));
	jdff dff_A_UIODt7P69_1(.dout(w_dff_A_NdTm2IRH8_1),.din(w_dff_A_UIODt7P69_1),.clk(gclk));
	jdff dff_A_KJ01KZjo3_1(.dout(w_dff_A_UIODt7P69_1),.din(w_dff_A_KJ01KZjo3_1),.clk(gclk));
	jdff dff_A_HpI7Zu6e0_1(.dout(w_dff_A_KJ01KZjo3_1),.din(w_dff_A_HpI7Zu6e0_1),.clk(gclk));
	jdff dff_A_nW4mItQv2_1(.dout(w_dff_A_HpI7Zu6e0_1),.din(w_dff_A_nW4mItQv2_1),.clk(gclk));
	jdff dff_B_Uq25joIQ0_1(.din(n537),.dout(w_dff_B_Uq25joIQ0_1),.clk(gclk));
	jdff dff_B_RbOHchf68_0(.din(G50),.dout(w_dff_B_RbOHchf68_0),.clk(gclk));
	jdff dff_B_Th2dA3IE6_2(.din(n536),.dout(w_dff_B_Th2dA3IE6_2),.clk(gclk));
	jdff dff_B_clWffWiI2_2(.din(w_dff_B_Th2dA3IE6_2),.dout(w_dff_B_clWffWiI2_2),.clk(gclk));
	jdff dff_A_232Wcgk02_0(.dout(w_G4432_1[0]),.din(w_dff_A_232Wcgk02_0),.clk(gclk));
	jdff dff_A_h4ekmAyz2_0(.dout(w_dff_A_232Wcgk02_0),.din(w_dff_A_h4ekmAyz2_0),.clk(gclk));
	jdff dff_A_MAUrdrhs9_0(.dout(w_dff_A_h4ekmAyz2_0),.din(w_dff_A_MAUrdrhs9_0),.clk(gclk));
	jdff dff_A_vK1SaVCu5_0(.dout(w_dff_A_MAUrdrhs9_0),.din(w_dff_A_vK1SaVCu5_0),.clk(gclk));
	jdff dff_B_zr9TvNSk1_1(.din(n1637),.dout(w_dff_B_zr9TvNSk1_1),.clk(gclk));
	jdff dff_B_Wfe7UT0x5_1(.din(w_dff_B_zr9TvNSk1_1),.dout(w_dff_B_Wfe7UT0x5_1),.clk(gclk));
	jdff dff_B_KqnuhGgy5_1(.din(w_dff_B_Wfe7UT0x5_1),.dout(w_dff_B_KqnuhGgy5_1),.clk(gclk));
	jdff dff_B_kmOdv2Jc1_1(.din(w_dff_B_KqnuhGgy5_1),.dout(w_dff_B_kmOdv2Jc1_1),.clk(gclk));
	jdff dff_B_2iXF6qVS1_1(.din(w_dff_B_kmOdv2Jc1_1),.dout(w_dff_B_2iXF6qVS1_1),.clk(gclk));
	jdff dff_B_VR6pvUXp8_1(.din(w_dff_B_2iXF6qVS1_1),.dout(w_dff_B_VR6pvUXp8_1),.clk(gclk));
	jdff dff_B_Z8lwB16C9_1(.din(w_dff_B_VR6pvUXp8_1),.dout(w_dff_B_Z8lwB16C9_1),.clk(gclk));
	jdff dff_B_aMHTsw7C1_1(.din(w_dff_B_Z8lwB16C9_1),.dout(w_dff_B_aMHTsw7C1_1),.clk(gclk));
	jdff dff_B_NpLUcPD67_1(.din(w_dff_B_aMHTsw7C1_1),.dout(w_dff_B_NpLUcPD67_1),.clk(gclk));
	jdff dff_B_KBuj21bs4_1(.din(w_dff_B_NpLUcPD67_1),.dout(w_dff_B_KBuj21bs4_1),.clk(gclk));
	jdff dff_B_VzJehx210_1(.din(w_dff_B_KBuj21bs4_1),.dout(w_dff_B_VzJehx210_1),.clk(gclk));
	jdff dff_B_U7wBcD9C1_1(.din(w_dff_B_VzJehx210_1),.dout(w_dff_B_U7wBcD9C1_1),.clk(gclk));
	jdff dff_B_iXzO8Qrp3_1(.din(w_dff_B_U7wBcD9C1_1),.dout(w_dff_B_iXzO8Qrp3_1),.clk(gclk));
	jdff dff_B_KiFOFoT63_1(.din(w_dff_B_iXzO8Qrp3_1),.dout(w_dff_B_KiFOFoT63_1),.clk(gclk));
	jdff dff_B_3LGbg9YE5_1(.din(w_dff_B_KiFOFoT63_1),.dout(w_dff_B_3LGbg9YE5_1),.clk(gclk));
	jdff dff_B_YN8G514S2_1(.din(n1666),.dout(w_dff_B_YN8G514S2_1),.clk(gclk));
	jdff dff_B_Ot2uxS2b8_1(.din(w_dff_B_YN8G514S2_1),.dout(w_dff_B_Ot2uxS2b8_1),.clk(gclk));
	jdff dff_B_LqYwp0DK4_1(.din(w_dff_B_Ot2uxS2b8_1),.dout(w_dff_B_LqYwp0DK4_1),.clk(gclk));
	jdff dff_B_cC0B5eQI6_0(.din(n1705),.dout(w_dff_B_cC0B5eQI6_0),.clk(gclk));
	jdff dff_B_mHSsPA474_1(.din(n1702),.dout(w_dff_B_mHSsPA474_1),.clk(gclk));
	jdff dff_B_FqaGOYoO0_1(.din(w_dff_B_mHSsPA474_1),.dout(w_dff_B_FqaGOYoO0_1),.clk(gclk));
	jdff dff_B_29kOIiyV1_0(.din(n1698),.dout(w_dff_B_29kOIiyV1_0),.clk(gclk));
	jdff dff_B_AOo5QAEB4_0(.din(w_dff_B_29kOIiyV1_0),.dout(w_dff_B_AOo5QAEB4_0),.clk(gclk));
	jdff dff_B_4WpU1ehT3_0(.din(w_dff_B_AOo5QAEB4_0),.dout(w_dff_B_4WpU1ehT3_0),.clk(gclk));
	jdff dff_B_fvd44txS3_0(.din(w_dff_B_4WpU1ehT3_0),.dout(w_dff_B_fvd44txS3_0),.clk(gclk));
	jdff dff_B_H5omkcwW9_0(.din(w_dff_B_fvd44txS3_0),.dout(w_dff_B_H5omkcwW9_0),.clk(gclk));
	jdff dff_B_ryHRoTbl5_0(.din(w_dff_B_H5omkcwW9_0),.dout(w_dff_B_ryHRoTbl5_0),.clk(gclk));
	jdff dff_B_tUAfxP7n4_0(.din(w_dff_B_ryHRoTbl5_0),.dout(w_dff_B_tUAfxP7n4_0),.clk(gclk));
	jdff dff_B_H0K3lUBb0_1(.din(n1690),.dout(w_dff_B_H0K3lUBb0_1),.clk(gclk));
	jdff dff_B_xleab02x0_1(.din(w_dff_B_H0K3lUBb0_1),.dout(w_dff_B_xleab02x0_1),.clk(gclk));
	jdff dff_B_tuMJqVnd7_1(.din(w_dff_B_xleab02x0_1),.dout(w_dff_B_tuMJqVnd7_1),.clk(gclk));
	jdff dff_B_2bGQ9w4O4_1(.din(w_dff_B_tuMJqVnd7_1),.dout(w_dff_B_2bGQ9w4O4_1),.clk(gclk));
	jdff dff_B_FuQFIgH88_1(.din(w_dff_B_2bGQ9w4O4_1),.dout(w_dff_B_FuQFIgH88_1),.clk(gclk));
	jdff dff_B_CIsA5jLb0_1(.din(n1691),.dout(w_dff_B_CIsA5jLb0_1),.clk(gclk));
	jdff dff_B_hWdk9Lp90_1(.din(w_dff_B_CIsA5jLb0_1),.dout(w_dff_B_hWdk9Lp90_1),.clk(gclk));
	jdff dff_B_v2w6Y5368_1(.din(w_dff_B_hWdk9Lp90_1),.dout(w_dff_B_v2w6Y5368_1),.clk(gclk));
	jdff dff_B_BaY2riKL9_1(.din(w_dff_B_v2w6Y5368_1),.dout(w_dff_B_BaY2riKL9_1),.clk(gclk));
	jdff dff_A_I1cbKSU18_1(.dout(w_n1687_0[1]),.din(w_dff_A_I1cbKSU18_1),.clk(gclk));
	jdff dff_A_qiZJRdEy0_1(.dout(w_dff_A_I1cbKSU18_1),.din(w_dff_A_qiZJRdEy0_1),.clk(gclk));
	jdff dff_A_riHYd6Xt7_1(.dout(w_dff_A_qiZJRdEy0_1),.din(w_dff_A_riHYd6Xt7_1),.clk(gclk));
	jdff dff_A_ybqhCZ7i9_1(.dout(w_dff_A_riHYd6Xt7_1),.din(w_dff_A_ybqhCZ7i9_1),.clk(gclk));
	jdff dff_B_yaGAndz76_1(.din(n1683),.dout(w_dff_B_yaGAndz76_1),.clk(gclk));
	jdff dff_A_qRjD17OP6_0(.dout(w_n1127_0[0]),.din(w_dff_A_qRjD17OP6_0),.clk(gclk));
	jdff dff_A_dTfLmEGw5_0(.dout(w_dff_A_qRjD17OP6_0),.din(w_dff_A_dTfLmEGw5_0),.clk(gclk));
	jdff dff_A_azqyXgUa4_0(.dout(w_dff_A_dTfLmEGw5_0),.din(w_dff_A_azqyXgUa4_0),.clk(gclk));
	jdff dff_B_78qQyTrY1_2(.din(n1127),.dout(w_dff_B_78qQyTrY1_2),.clk(gclk));
	jdff dff_B_zFxoyLqs4_2(.din(w_dff_B_78qQyTrY1_2),.dout(w_dff_B_zFxoyLqs4_2),.clk(gclk));
	jdff dff_B_yKeTjvzk6_2(.din(w_dff_B_zFxoyLqs4_2),.dout(w_dff_B_yKeTjvzk6_2),.clk(gclk));
	jdff dff_B_pfOlVf9R1_2(.din(w_dff_B_yKeTjvzk6_2),.dout(w_dff_B_pfOlVf9R1_2),.clk(gclk));
	jdff dff_A_T06DSO181_1(.dout(w_n1675_0[1]),.din(w_dff_A_T06DSO181_1),.clk(gclk));
	jdff dff_A_bUccLvCp0_1(.dout(w_dff_A_T06DSO181_1),.din(w_dff_A_bUccLvCp0_1),.clk(gclk));
	jdff dff_A_4DWiGXIG0_1(.dout(w_dff_A_bUccLvCp0_1),.din(w_dff_A_4DWiGXIG0_1),.clk(gclk));
	jdff dff_B_OGgUC0wS8_1(.din(n1669),.dout(w_dff_B_OGgUC0wS8_1),.clk(gclk));
	jdff dff_B_REeW9gvT5_1(.din(w_dff_B_OGgUC0wS8_1),.dout(w_dff_B_REeW9gvT5_1),.clk(gclk));
	jdff dff_B_psoXIpxT9_0(.din(n1671),.dout(w_dff_B_psoXIpxT9_0),.clk(gclk));
	jdff dff_B_jxRLmfFY1_0(.din(w_dff_B_psoXIpxT9_0),.dout(w_dff_B_jxRLmfFY1_0),.clk(gclk));
	jdff dff_A_ZJHbP3dP6_0(.dout(w_n1667_0[0]),.din(w_dff_A_ZJHbP3dP6_0),.clk(gclk));
	jdff dff_A_CBVuSnub1_0(.dout(w_dff_A_ZJHbP3dP6_0),.din(w_dff_A_CBVuSnub1_0),.clk(gclk));
	jdff dff_A_ZPEdoOs90_0(.dout(w_dff_A_CBVuSnub1_0),.din(w_dff_A_ZPEdoOs90_0),.clk(gclk));
	jdff dff_A_vpVwBZGG7_1(.dout(w_n1136_0[1]),.din(w_dff_A_vpVwBZGG7_1),.clk(gclk));
	jdff dff_B_rjvqatEd1_1(.din(n1649),.dout(w_dff_B_rjvqatEd1_1),.clk(gclk));
	jdff dff_B_wHCiczz55_1(.din(w_dff_B_rjvqatEd1_1),.dout(w_dff_B_wHCiczz55_1),.clk(gclk));
	jdff dff_B_JRcaNep85_1(.din(w_dff_B_wHCiczz55_1),.dout(w_dff_B_JRcaNep85_1),.clk(gclk));
	jdff dff_B_QUIsBXBh1_1(.din(n1660),.dout(w_dff_B_QUIsBXBh1_1),.clk(gclk));
	jdff dff_B_j4SVgvbl0_1(.din(w_dff_B_QUIsBXBh1_1),.dout(w_dff_B_j4SVgvbl0_1),.clk(gclk));
	jdff dff_B_4Wj5yp2j5_1(.din(n1661),.dout(w_dff_B_4Wj5yp2j5_1),.clk(gclk));
	jdff dff_B_qAlmacbT0_1(.din(w_dff_B_4Wj5yp2j5_1),.dout(w_dff_B_qAlmacbT0_1),.clk(gclk));
	jdff dff_B_Lzk0vi2H7_1(.din(w_dff_B_qAlmacbT0_1),.dout(w_dff_B_Lzk0vi2H7_1),.clk(gclk));
	jdff dff_B_zd0yajDr0_1(.din(w_dff_B_Lzk0vi2H7_1),.dout(w_dff_B_zd0yajDr0_1),.clk(gclk));
	jdff dff_B_lbznyI1u1_1(.din(w_dff_B_zd0yajDr0_1),.dout(w_dff_B_lbznyI1u1_1),.clk(gclk));
	jdff dff_A_9qZgzsNs9_0(.dout(w_n1376_0[0]),.din(w_dff_A_9qZgzsNs9_0),.clk(gclk));
	jdff dff_A_TdBdHRL18_0(.dout(w_dff_A_9qZgzsNs9_0),.din(w_dff_A_TdBdHRL18_0),.clk(gclk));
	jdff dff_A_9yFEB4Tk7_0(.dout(w_dff_A_TdBdHRL18_0),.din(w_dff_A_9yFEB4Tk7_0),.clk(gclk));
	jdff dff_A_6Yzdt3Ak2_0(.dout(w_dff_A_9yFEB4Tk7_0),.din(w_dff_A_6Yzdt3Ak2_0),.clk(gclk));
	jdff dff_B_o9uY41Ac7_1(.din(n1366),.dout(w_dff_B_o9uY41Ac7_1),.clk(gclk));
	jdff dff_A_cV1ghasb7_1(.dout(w_n1361_0[1]),.din(w_dff_A_cV1ghasb7_1),.clk(gclk));
	jdff dff_A_MK79zHne4_0(.dout(w_G3705_1[0]),.din(w_dff_A_MK79zHne4_0),.clk(gclk));
	jdff dff_A_mqnS2Z4X2_0(.dout(w_dff_A_MK79zHne4_0),.din(w_dff_A_mqnS2Z4X2_0),.clk(gclk));
	jdff dff_A_Pbera6bC7_0(.dout(w_dff_A_mqnS2Z4X2_0),.din(w_dff_A_Pbera6bC7_0),.clk(gclk));
	jdff dff_A_MV8HZdIY7_1(.dout(w_G3705_1[1]),.din(w_dff_A_MV8HZdIY7_1),.clk(gclk));
	jdff dff_A_wEcAMxBO0_1(.dout(w_dff_A_MV8HZdIY7_1),.din(w_dff_A_wEcAMxBO0_1),.clk(gclk));
	jdff dff_A_r4uRtzhq8_1(.dout(w_dff_A_wEcAMxBO0_1),.din(w_dff_A_r4uRtzhq8_1),.clk(gclk));
	jdff dff_A_kNbcT2hR0_0(.dout(w_n362_0[0]),.din(w_dff_A_kNbcT2hR0_0),.clk(gclk));
	jdff dff_A_BXHabmH63_0(.dout(w_dff_A_kNbcT2hR0_0),.din(w_dff_A_BXHabmH63_0),.clk(gclk));
	jdff dff_A_CszolQZC5_0(.dout(w_dff_A_BXHabmH63_0),.din(w_dff_A_CszolQZC5_0),.clk(gclk));
	jdff dff_A_7BAqe4RH3_0(.dout(w_dff_A_CszolQZC5_0),.din(w_dff_A_7BAqe4RH3_0),.clk(gclk));
	jdff dff_A_sOHOWnrF9_0(.dout(w_dff_A_7BAqe4RH3_0),.din(w_dff_A_sOHOWnrF9_0),.clk(gclk));
	jdff dff_B_qH8YMZAq3_0(.din(n357),.dout(w_dff_B_qH8YMZAq3_0),.clk(gclk));
	jdff dff_A_zgO2fUiT9_1(.dout(w_n1360_1[1]),.din(w_dff_A_zgO2fUiT9_1),.clk(gclk));
	jdff dff_A_5wPFBUs39_1(.dout(w_dff_A_zgO2fUiT9_1),.din(w_dff_A_5wPFBUs39_1),.clk(gclk));
	jdff dff_A_YU2PxwHh9_1(.dout(w_n1359_0[1]),.din(w_dff_A_YU2PxwHh9_1),.clk(gclk));
	jdff dff_A_u9w86PM44_2(.dout(w_n1359_0[2]),.din(w_dff_A_u9w86PM44_2),.clk(gclk));
	jdff dff_A_1fPZMeRr7_2(.dout(w_dff_A_u9w86PM44_2),.din(w_dff_A_1fPZMeRr7_2),.clk(gclk));
	jdff dff_B_P9QBsc5k9_0(.din(n1358),.dout(w_dff_B_P9QBsc5k9_0),.clk(gclk));
	jdff dff_A_8VN8W2Jp5_0(.dout(w_G3717_1[0]),.din(w_dff_A_8VN8W2Jp5_0),.clk(gclk));
	jdff dff_A_FFoxzIYb8_0(.dout(w_dff_A_8VN8W2Jp5_0),.din(w_dff_A_FFoxzIYb8_0),.clk(gclk));
	jdff dff_A_fUSrVCF72_0(.dout(w_dff_A_FFoxzIYb8_0),.din(w_dff_A_fUSrVCF72_0),.clk(gclk));
	jdff dff_A_UZkBPwWu9_1(.dout(w_G3717_1[1]),.din(w_dff_A_UZkBPwWu9_1),.clk(gclk));
	jdff dff_A_BRbsPw8B7_1(.dout(w_dff_A_UZkBPwWu9_1),.din(w_dff_A_BRbsPw8B7_1),.clk(gclk));
	jdff dff_A_SXnMlaJE4_1(.dout(w_dff_A_BRbsPw8B7_1),.din(w_dff_A_SXnMlaJE4_1),.clk(gclk));
	jdff dff_B_vA4D5r9z7_0(.din(n1658),.dout(w_dff_B_vA4D5r9z7_0),.clk(gclk));
	jdff dff_B_wtTzXQZ68_0(.din(w_dff_B_vA4D5r9z7_0),.dout(w_dff_B_wtTzXQZ68_0),.clk(gclk));
	jdff dff_B_5MKJui9C7_0(.din(w_dff_B_wtTzXQZ68_0),.dout(w_dff_B_5MKJui9C7_0),.clk(gclk));
	jdff dff_B_iWkXe2AJ4_0(.din(w_dff_B_5MKJui9C7_0),.dout(w_dff_B_iWkXe2AJ4_0),.clk(gclk));
	jdff dff_A_BxX42A2O3_1(.dout(w_n1654_0[1]),.din(w_dff_A_BxX42A2O3_1),.clk(gclk));
	jdff dff_A_5gRjoGy61_1(.dout(w_dff_A_BxX42A2O3_1),.din(w_dff_A_5gRjoGy61_1),.clk(gclk));
	jdff dff_A_0WhToFMW5_1(.dout(w_dff_A_5gRjoGy61_1),.din(w_dff_A_0WhToFMW5_1),.clk(gclk));
	jdff dff_A_fDmLV9JP5_1(.dout(w_n462_0[1]),.din(w_dff_A_fDmLV9JP5_1),.clk(gclk));
	jdff dff_A_wWhXJe5g4_1(.dout(w_dff_A_fDmLV9JP5_1),.din(w_dff_A_wWhXJe5g4_1),.clk(gclk));
	jdff dff_A_oqZruxcR8_1(.dout(w_dff_A_wWhXJe5g4_1),.din(w_dff_A_oqZruxcR8_1),.clk(gclk));
	jdff dff_A_PKKRSAtR4_1(.dout(w_dff_A_oqZruxcR8_1),.din(w_dff_A_PKKRSAtR4_1),.clk(gclk));
	jdff dff_A_DOXs29d90_1(.dout(w_n1651_0[1]),.din(w_dff_A_DOXs29d90_1),.clk(gclk));
	jdff dff_A_X1w6X3UH9_1(.dout(w_dff_A_DOXs29d90_1),.din(w_dff_A_X1w6X3UH9_1),.clk(gclk));
	jdff dff_A_oJGc6wik0_1(.dout(w_dff_A_X1w6X3UH9_1),.din(w_dff_A_oJGc6wik0_1),.clk(gclk));
	jdff dff_A_tvCdJFBR8_1(.dout(w_dff_A_oJGc6wik0_1),.din(w_dff_A_tvCdJFBR8_1),.clk(gclk));
	jdff dff_A_bMRYvsgy9_1(.dout(w_dff_A_tvCdJFBR8_1),.din(w_dff_A_bMRYvsgy9_1),.clk(gclk));
	jdff dff_B_KeNprzu58_0(.din(n1650),.dout(w_dff_B_KeNprzu58_0),.clk(gclk));
	jdff dff_A_sTYy0b9H1_1(.dout(w_n422_0[1]),.din(w_dff_A_sTYy0b9H1_1),.clk(gclk));
	jdff dff_A_sBgJxJKt1_1(.dout(w_n419_0[1]),.din(w_dff_A_sBgJxJKt1_1),.clk(gclk));
	jdff dff_B_5GHdNSKJ6_1(.din(n415),.dout(w_dff_B_5GHdNSKJ6_1),.clk(gclk));
	jdff dff_A_Oh3JpdHS7_0(.dout(w_n417_0[0]),.din(w_dff_A_Oh3JpdHS7_0),.clk(gclk));
	jdff dff_A_6M5Ju3np0_0(.dout(w_dff_A_Oh3JpdHS7_0),.din(w_dff_A_6M5Ju3np0_0),.clk(gclk));
	jdff dff_A_5vS2KP6j3_0(.dout(w_dff_A_6M5Ju3np0_0),.din(w_dff_A_5vS2KP6j3_0),.clk(gclk));
	jdff dff_A_uuWTafWp4_0(.dout(w_dff_A_5vS2KP6j3_0),.din(w_dff_A_uuWTafWp4_0),.clk(gclk));
	jdff dff_A_iqDMWr1G8_0(.dout(w_dff_A_uuWTafWp4_0),.din(w_dff_A_iqDMWr1G8_0),.clk(gclk));
	jdff dff_A_2ORK7MJ96_0(.dout(w_dff_A_iqDMWr1G8_0),.din(w_dff_A_2ORK7MJ96_0),.clk(gclk));
	jdff dff_A_ruTERdd65_0(.dout(w_dff_A_2ORK7MJ96_0),.din(w_dff_A_ruTERdd65_0),.clk(gclk));
	jdff dff_A_PFrRtPz72_0(.dout(w_dff_A_ruTERdd65_0),.din(w_dff_A_PFrRtPz72_0),.clk(gclk));
	jdff dff_A_v76VSXqZ6_1(.dout(w_n417_0[1]),.din(w_dff_A_v76VSXqZ6_1),.clk(gclk));
	jdff dff_A_JAoynUOq8_1(.dout(w_dff_A_v76VSXqZ6_1),.din(w_dff_A_JAoynUOq8_1),.clk(gclk));
	jdff dff_A_rShiufyc4_1(.dout(w_dff_A_JAoynUOq8_1),.din(w_dff_A_rShiufyc4_1),.clk(gclk));
	jdff dff_A_u95AvtUA5_1(.dout(w_dff_A_rShiufyc4_1),.din(w_dff_A_u95AvtUA5_1),.clk(gclk));
	jdff dff_A_Mu6B6EbU7_1(.dout(w_dff_A_u95AvtUA5_1),.din(w_dff_A_Mu6B6EbU7_1),.clk(gclk));
	jdff dff_A_8TRro6Rh2_0(.dout(w_n413_1[0]),.din(w_dff_A_8TRro6Rh2_0),.clk(gclk));
	jdff dff_A_74cnW4016_0(.dout(w_n413_0[0]),.din(w_dff_A_74cnW4016_0),.clk(gclk));
	jdff dff_A_qPeJQYRD1_0(.dout(w_n412_0[0]),.din(w_dff_A_qPeJQYRD1_0),.clk(gclk));
	jdff dff_A_9H4knwf08_1(.dout(w_n412_0[1]),.din(w_dff_A_9H4knwf08_1),.clk(gclk));
	jdff dff_A_AIM5S5t53_0(.dout(w_n354_1[0]),.din(w_dff_A_AIM5S5t53_0),.clk(gclk));
	jdff dff_A_5gSkhRnC7_0(.dout(w_dff_A_AIM5S5t53_0),.din(w_dff_A_5gSkhRnC7_0),.clk(gclk));
	jdff dff_A_TbXBDE7v1_2(.dout(w_n354_0[2]),.din(w_dff_A_TbXBDE7v1_2),.clk(gclk));
	jdff dff_A_68KSUdat4_2(.dout(w_dff_A_TbXBDE7v1_2),.din(w_dff_A_68KSUdat4_2),.clk(gclk));
	jdff dff_A_B6Cf6Acw1_2(.dout(w_dff_A_68KSUdat4_2),.din(w_dff_A_B6Cf6Acw1_2),.clk(gclk));
	jdff dff_A_WFaEeLe79_2(.dout(w_dff_A_B6Cf6Acw1_2),.din(w_dff_A_WFaEeLe79_2),.clk(gclk));
	jdff dff_A_8oLxctnW1_2(.dout(w_dff_A_WFaEeLe79_2),.din(w_dff_A_8oLxctnW1_2),.clk(gclk));
	jdff dff_A_G9vcx2wh9_2(.dout(w_dff_A_8oLxctnW1_2),.din(w_dff_A_G9vcx2wh9_2),.clk(gclk));
	jdff dff_A_36dz6SZj6_2(.dout(w_dff_A_G9vcx2wh9_2),.din(w_dff_A_36dz6SZj6_2),.clk(gclk));
	jdff dff_A_PWZDMPJl4_2(.dout(w_dff_A_36dz6SZj6_2),.din(w_dff_A_PWZDMPJl4_2),.clk(gclk));
	jdff dff_A_WWKtgBrA9_2(.dout(w_dff_A_PWZDMPJl4_2),.din(w_dff_A_WWKtgBrA9_2),.clk(gclk));
	jdff dff_A_b2eYmO4R5_2(.dout(w_dff_A_WWKtgBrA9_2),.din(w_dff_A_b2eYmO4R5_2),.clk(gclk));
	jdff dff_B_KidPtzUp6_3(.din(n354),.dout(w_dff_B_KidPtzUp6_3),.clk(gclk));
	jdff dff_A_wN9Pvajd7_2(.dout(w_n407_0[2]),.din(w_dff_A_wN9Pvajd7_2),.clk(gclk));
	jdff dff_A_VW7Yj6298_2(.dout(w_dff_A_wN9Pvajd7_2),.din(w_dff_A_VW7Yj6298_2),.clk(gclk));
	jdff dff_A_DknvD8Cx1_1(.dout(w_n402_1[1]),.din(w_dff_A_DknvD8Cx1_1),.clk(gclk));
	jdff dff_A_hy19a9jk7_1(.dout(w_n402_0[1]),.din(w_dff_A_hy19a9jk7_1),.clk(gclk));
	jdff dff_A_UK6liytN6_1(.dout(w_dff_A_hy19a9jk7_1),.din(w_dff_A_UK6liytN6_1),.clk(gclk));
	jdff dff_A_Y35dsLT03_1(.dout(w_dff_A_UK6liytN6_1),.din(w_dff_A_Y35dsLT03_1),.clk(gclk));
	jdff dff_A_NW0XW22D6_1(.dout(w_dff_A_Y35dsLT03_1),.din(w_dff_A_NW0XW22D6_1),.clk(gclk));
	jdff dff_A_5hMSZaFC4_1(.dout(w_dff_A_NW0XW22D6_1),.din(w_dff_A_5hMSZaFC4_1),.clk(gclk));
	jdff dff_A_JmylGvGX8_1(.dout(w_dff_A_5hMSZaFC4_1),.din(w_dff_A_JmylGvGX8_1),.clk(gclk));
	jdff dff_A_GRIDOSq39_1(.dout(w_dff_A_JmylGvGX8_1),.din(w_dff_A_GRIDOSq39_1),.clk(gclk));
	jdff dff_A_0cOZA6cA9_1(.dout(w_dff_A_GRIDOSq39_1),.din(w_dff_A_0cOZA6cA9_1),.clk(gclk));
	jdff dff_A_7gf8DVbR1_1(.dout(w_dff_A_0cOZA6cA9_1),.din(w_dff_A_7gf8DVbR1_1),.clk(gclk));
	jdff dff_A_fn373POl2_2(.dout(w_n402_0[2]),.din(w_dff_A_fn373POl2_2),.clk(gclk));
	jdff dff_A_Agm25rVm7_2(.dout(w_dff_A_fn373POl2_2),.din(w_dff_A_Agm25rVm7_2),.clk(gclk));
	jdff dff_A_QTlFZtkZ7_2(.dout(w_dff_A_Agm25rVm7_2),.din(w_dff_A_QTlFZtkZ7_2),.clk(gclk));
	jdff dff_B_ijgckosu9_1(.din(n396),.dout(w_dff_B_ijgckosu9_1),.clk(gclk));
	jdff dff_B_sTsRkrCo0_1(.din(w_dff_B_ijgckosu9_1),.dout(w_dff_B_sTsRkrCo0_1),.clk(gclk));
	jdff dff_A_0fReXTFg6_0(.dout(w_G3705_2[0]),.din(w_dff_A_0fReXTFg6_0),.clk(gclk));
	jdff dff_A_kVT3uzCz5_0(.dout(w_dff_A_0fReXTFg6_0),.din(w_dff_A_kVT3uzCz5_0),.clk(gclk));
	jdff dff_A_MeHNMQtc8_0(.dout(w_dff_A_kVT3uzCz5_0),.din(w_dff_A_MeHNMQtc8_0),.clk(gclk));
	jdff dff_A_uSWqszjk6_0(.dout(w_n395_0[0]),.din(w_dff_A_uSWqszjk6_0),.clk(gclk));
	jdff dff_A_sK9IWy2v7_0(.dout(w_n359_0[0]),.din(w_dff_A_sK9IWy2v7_0),.clk(gclk));
	jdff dff_A_MSVHLPQs9_1(.dout(w_G3701_1[1]),.din(w_dff_A_MSVHLPQs9_1),.clk(gclk));
	jdff dff_A_ZxAd4Hdj4_2(.dout(w_n390_0[2]),.din(w_dff_A_ZxAd4Hdj4_2),.clk(gclk));
	jdff dff_A_xb6S6qui0_2(.dout(w_dff_A_ZxAd4Hdj4_2),.din(w_dff_A_xb6S6qui0_2),.clk(gclk));
	jdff dff_A_nMiP9VN05_2(.dout(w_dff_A_xb6S6qui0_2),.din(w_dff_A_nMiP9VN05_2),.clk(gclk));
	jdff dff_A_fNiV9ITl2_2(.dout(w_dff_A_nMiP9VN05_2),.din(w_dff_A_fNiV9ITl2_2),.clk(gclk));
	jdff dff_A_oaivMi756_2(.dout(w_dff_A_fNiV9ITl2_2),.din(w_dff_A_oaivMi756_2),.clk(gclk));
	jdff dff_B_26IBZNyP1_3(.din(n390),.dout(w_dff_B_26IBZNyP1_3),.clk(gclk));
	jdff dff_A_5Sf6yYef6_0(.dout(w_n356_0[0]),.din(w_dff_A_5Sf6yYef6_0),.clk(gclk));
	jdff dff_A_DItjsZtr7_0(.dout(w_G41_0[0]),.din(w_dff_A_DItjsZtr7_0),.clk(gclk));
	jdff dff_A_aE5bhzcy6_0(.dout(w_dff_A_DItjsZtr7_0),.din(w_dff_A_aE5bhzcy6_0),.clk(gclk));
	jdff dff_A_VMwgvIR75_0(.dout(w_dff_A_aE5bhzcy6_0),.din(w_dff_A_VMwgvIR75_0),.clk(gclk));
	jdff dff_A_1JWV0Pyl7_1(.dout(w_G41_0[1]),.din(w_dff_A_1JWV0Pyl7_1),.clk(gclk));
	jdff dff_A_NVapzCBn3_1(.dout(w_n389_0[1]),.din(w_dff_A_NVapzCBn3_1),.clk(gclk));
	jdff dff_A_iUgl4et14_0(.dout(w_G3701_0[0]),.din(w_dff_A_iUgl4et14_0),.clk(gclk));
	jdff dff_A_7xgMrx8f8_0(.dout(w_n388_0[0]),.din(w_dff_A_7xgMrx8f8_0),.clk(gclk));
	jdff dff_A_L8oEP3pi9_0(.dout(w_dff_A_7xgMrx8f8_0),.din(w_dff_A_L8oEP3pi9_0),.clk(gclk));
	jdff dff_A_CM5uF7Q79_0(.dout(w_dff_A_L8oEP3pi9_0),.din(w_dff_A_CM5uF7Q79_0),.clk(gclk));
	jdff dff_A_jQm4POQd1_0(.dout(w_dff_A_CM5uF7Q79_0),.din(w_dff_A_jQm4POQd1_0),.clk(gclk));
	jdff dff_A_ueMveMMH3_0(.dout(w_dff_A_jQm4POQd1_0),.din(w_dff_A_ueMveMMH3_0),.clk(gclk));
	jdff dff_A_7njmmzcU3_0(.dout(w_dff_A_ueMveMMH3_0),.din(w_dff_A_7njmmzcU3_0),.clk(gclk));
	jdff dff_A_JivydptM7_0(.dout(w_dff_A_7njmmzcU3_0),.din(w_dff_A_JivydptM7_0),.clk(gclk));
	jdff dff_A_FHod2HfN7_0(.dout(w_dff_A_JivydptM7_0),.din(w_dff_A_FHod2HfN7_0),.clk(gclk));
	jdff dff_A_n9lY1H8r0_0(.dout(w_dff_A_FHod2HfN7_0),.din(w_dff_A_n9lY1H8r0_0),.clk(gclk));
	jdff dff_A_DsbOikcy1_0(.dout(w_dff_A_n9lY1H8r0_0),.din(w_dff_A_DsbOikcy1_0),.clk(gclk));
	jdff dff_A_QLd0u7Pk2_0(.dout(w_dff_A_DsbOikcy1_0),.din(w_dff_A_QLd0u7Pk2_0),.clk(gclk));
	jdff dff_A_t2vvxLIv2_2(.dout(w_n388_0[2]),.din(w_dff_A_t2vvxLIv2_2),.clk(gclk));
	jdff dff_B_P9oTzFiG0_3(.din(n388),.dout(w_dff_B_P9oTzFiG0_3),.clk(gclk));
	jdff dff_B_pLDP2Vqt9_3(.din(w_dff_B_P9oTzFiG0_3),.dout(w_dff_B_pLDP2Vqt9_3),.clk(gclk));
	jdff dff_B_TBNi1hV02_3(.din(w_dff_B_pLDP2Vqt9_3),.dout(w_dff_B_TBNi1hV02_3),.clk(gclk));
	jdff dff_B_mLOxX17m9_3(.din(w_dff_B_TBNi1hV02_3),.dout(w_dff_B_mLOxX17m9_3),.clk(gclk));
	jdff dff_A_X2hJZbNH9_1(.dout(w_G4526_1[1]),.din(w_dff_A_X2hJZbNH9_1),.clk(gclk));
	jdff dff_A_rTCYYuTb9_1(.dout(w_dff_A_X2hJZbNH9_1),.din(w_dff_A_rTCYYuTb9_1),.clk(gclk));
	jdff dff_A_MJsQ6nGm6_1(.dout(w_dff_A_rTCYYuTb9_1),.din(w_dff_A_MJsQ6nGm6_1),.clk(gclk));
	jdff dff_A_BpQsFthV1_1(.dout(w_dff_A_MJsQ6nGm6_1),.din(w_dff_A_BpQsFthV1_1),.clk(gclk));
	jdff dff_A_ms5Q6tOQ7_1(.dout(w_dff_A_BpQsFthV1_1),.din(w_dff_A_ms5Q6tOQ7_1),.clk(gclk));
	jdff dff_A_9PM9D7hK7_1(.dout(w_G4526_0[1]),.din(w_dff_A_9PM9D7hK7_1),.clk(gclk));
	jdff dff_A_WKlATLgI7_1(.dout(w_dff_A_9PM9D7hK7_1),.din(w_dff_A_WKlATLgI7_1),.clk(gclk));
	jdff dff_A_fy6nSdI54_1(.dout(w_dff_A_WKlATLgI7_1),.din(w_dff_A_fy6nSdI54_1),.clk(gclk));
	jdff dff_A_PgvoQJuA2_1(.dout(w_dff_A_fy6nSdI54_1),.din(w_dff_A_PgvoQJuA2_1),.clk(gclk));
	jdff dff_A_UdbUjPSL4_1(.dout(w_dff_A_PgvoQJuA2_1),.din(w_dff_A_UdbUjPSL4_1),.clk(gclk));
	jdff dff_A_VpOZSvnH0_1(.dout(w_dff_A_UdbUjPSL4_1),.din(w_dff_A_VpOZSvnH0_1),.clk(gclk));
	jdff dff_A_PRsLHwbW7_1(.dout(w_dff_A_VpOZSvnH0_1),.din(w_dff_A_PRsLHwbW7_1),.clk(gclk));
	jdff dff_A_VDwri5zt0_1(.dout(w_dff_A_PRsLHwbW7_1),.din(w_dff_A_VDwri5zt0_1),.clk(gclk));
	jdff dff_A_6LaLYoZz7_1(.dout(w_dff_A_VDwri5zt0_1),.din(w_dff_A_6LaLYoZz7_1),.clk(gclk));
	jdff dff_A_XDKhkYet6_1(.dout(w_dff_A_6LaLYoZz7_1),.din(w_dff_A_XDKhkYet6_1),.clk(gclk));
	jdff dff_A_DLlCpuQU8_1(.dout(w_dff_A_XDKhkYet6_1),.din(w_dff_A_DLlCpuQU8_1),.clk(gclk));
	jdff dff_A_Vvn0hPCn1_1(.dout(w_dff_A_DLlCpuQU8_1),.din(w_dff_A_Vvn0hPCn1_1),.clk(gclk));
	jdff dff_A_YOC4rDdX5_1(.dout(w_dff_A_Vvn0hPCn1_1),.din(w_dff_A_YOC4rDdX5_1),.clk(gclk));
	jdff dff_A_2bAkTEUW4_1(.dout(w_dff_A_YOC4rDdX5_1),.din(w_dff_A_2bAkTEUW4_1),.clk(gclk));
	jdff dff_A_d505jNZO2_1(.dout(w_dff_A_2bAkTEUW4_1),.din(w_dff_A_d505jNZO2_1),.clk(gclk));
	jdff dff_A_9M9WJaAl2_2(.dout(w_G4526_0[2]),.din(w_dff_A_9M9WJaAl2_2),.clk(gclk));
	jdff dff_A_vPudiIHb7_2(.dout(w_dff_A_9M9WJaAl2_2),.din(w_dff_A_vPudiIHb7_2),.clk(gclk));
	jdff dff_A_nuR6vZS55_2(.dout(w_dff_A_vPudiIHb7_2),.din(w_dff_A_nuR6vZS55_2),.clk(gclk));
	jdff dff_A_u6pCXeVY1_2(.dout(w_dff_A_nuR6vZS55_2),.din(w_dff_A_u6pCXeVY1_2),.clk(gclk));
	jdff dff_A_FlXCStQ04_2(.dout(w_dff_A_u6pCXeVY1_2),.din(w_dff_A_FlXCStQ04_2),.clk(gclk));
	jdff dff_A_CGzIPUJQ0_2(.dout(w_dff_A_FlXCStQ04_2),.din(w_dff_A_CGzIPUJQ0_2),.clk(gclk));
	jdff dff_A_fptldo2Z1_1(.dout(w_n387_1[1]),.din(w_dff_A_fptldo2Z1_1),.clk(gclk));
	jdff dff_A_UfqrjIig3_2(.dout(w_n387_1[2]),.din(w_dff_A_UfqrjIig3_2),.clk(gclk));
	jdff dff_A_XjEUdPLg8_2(.dout(w_dff_A_UfqrjIig3_2),.din(w_dff_A_XjEUdPLg8_2),.clk(gclk));
	jdff dff_A_8zOw0JFN9_2(.dout(w_dff_A_XjEUdPLg8_2),.din(w_dff_A_8zOw0JFN9_2),.clk(gclk));
	jdff dff_A_ujmd7dth2_1(.dout(w_n380_0[1]),.din(w_dff_A_ujmd7dth2_1),.clk(gclk));
	jdff dff_A_fxhrM4H85_2(.dout(w_n380_0[2]),.din(w_dff_A_fxhrM4H85_2),.clk(gclk));
	jdff dff_A_QCnVwtnx0_2(.dout(w_dff_A_fxhrM4H85_2),.din(w_dff_A_QCnVwtnx0_2),.clk(gclk));
	jdff dff_A_NsVQY6dY5_0(.dout(w_n379_1[0]),.din(w_dff_A_NsVQY6dY5_0),.clk(gclk));
	jdff dff_A_tlg9K5ml4_0(.dout(w_dff_A_NsVQY6dY5_0),.din(w_dff_A_tlg9K5ml4_0),.clk(gclk));
	jdff dff_A_uFNboZ7w4_0(.dout(w_dff_A_tlg9K5ml4_0),.din(w_dff_A_uFNboZ7w4_0),.clk(gclk));
	jdff dff_A_KIbxWG680_1(.dout(w_n379_0[1]),.din(w_dff_A_KIbxWG680_1),.clk(gclk));
	jdff dff_A_nsY4tZgM7_1(.dout(w_dff_A_KIbxWG680_1),.din(w_dff_A_nsY4tZgM7_1),.clk(gclk));
	jdff dff_A_T4oDNzeA1_1(.dout(w_dff_A_nsY4tZgM7_1),.din(w_dff_A_T4oDNzeA1_1),.clk(gclk));
	jdff dff_A_lAUA7D2V6_1(.dout(w_dff_A_T4oDNzeA1_1),.din(w_dff_A_lAUA7D2V6_1),.clk(gclk));
	jdff dff_A_E1HN2sYi3_1(.dout(w_dff_A_lAUA7D2V6_1),.din(w_dff_A_E1HN2sYi3_1),.clk(gclk));
	jdff dff_A_gi09h5j40_1(.dout(w_dff_A_E1HN2sYi3_1),.din(w_dff_A_gi09h5j40_1),.clk(gclk));
	jdff dff_A_AiXPINR31_1(.dout(w_dff_A_gi09h5j40_1),.din(w_dff_A_AiXPINR31_1),.clk(gclk));
	jdff dff_A_c0J9rYi81_1(.dout(w_dff_A_AiXPINR31_1),.din(w_dff_A_c0J9rYi81_1),.clk(gclk));
	jdff dff_A_wDZaEiJY1_1(.dout(w_dff_A_c0J9rYi81_1),.din(w_dff_A_wDZaEiJY1_1),.clk(gclk));
	jdff dff_A_YFnBr3dz8_1(.dout(w_dff_A_wDZaEiJY1_1),.din(w_dff_A_YFnBr3dz8_1),.clk(gclk));
	jdff dff_A_rLEOKtgO7_1(.dout(w_dff_A_YFnBr3dz8_1),.din(w_dff_A_rLEOKtgO7_1),.clk(gclk));
	jdff dff_A_Y7XVqhIw2_1(.dout(w_dff_A_rLEOKtgO7_1),.din(w_dff_A_Y7XVqhIw2_1),.clk(gclk));
	jdff dff_A_2xgicKFQ5_1(.dout(w_dff_A_Y7XVqhIw2_1),.din(w_dff_A_2xgicKFQ5_1),.clk(gclk));
	jdff dff_A_k9uy9nRV1_1(.dout(w_dff_A_2xgicKFQ5_1),.din(w_dff_A_k9uy9nRV1_1),.clk(gclk));
	jdff dff_A_lxXH7riZ8_2(.dout(w_n379_0[2]),.din(w_dff_A_lxXH7riZ8_2),.clk(gclk));
	jdff dff_A_isE6yyPm5_2(.dout(w_dff_A_lxXH7riZ8_2),.din(w_dff_A_isE6yyPm5_2),.clk(gclk));
	jdff dff_A_yXdKgWiP7_2(.dout(w_dff_A_isE6yyPm5_2),.din(w_dff_A_yXdKgWiP7_2),.clk(gclk));
	jdff dff_A_JeDlUWyh1_2(.dout(w_dff_A_yXdKgWiP7_2),.din(w_dff_A_JeDlUWyh1_2),.clk(gclk));
	jdff dff_A_pzV3NkDf7_2(.dout(w_n377_0[2]),.din(w_dff_A_pzV3NkDf7_2),.clk(gclk));
	jdff dff_A_Y5zX2Jn48_1(.dout(w_G3717_2[1]),.din(w_dff_A_Y5zX2Jn48_1),.clk(gclk));
	jdff dff_A_Awt1ZS5b6_1(.dout(w_G3717_0[1]),.din(w_dff_A_Awt1ZS5b6_1),.clk(gclk));
	jdff dff_A_f4GZOwov5_1(.dout(w_dff_A_Awt1ZS5b6_1),.din(w_dff_A_f4GZOwov5_1),.clk(gclk));
	jdff dff_A_MjfUwtZn7_1(.dout(w_dff_A_f4GZOwov5_1),.din(w_dff_A_MjfUwtZn7_1),.clk(gclk));
	jdff dff_A_QzaHcTNw8_1(.dout(w_n372_1[1]),.din(w_dff_A_QzaHcTNw8_1),.clk(gclk));
	jdff dff_A_xNRUv05R1_1(.dout(w_dff_A_QzaHcTNw8_1),.din(w_dff_A_xNRUv05R1_1),.clk(gclk));
	jdff dff_A_zfdkBFJC6_1(.dout(w_dff_A_xNRUv05R1_1),.din(w_dff_A_zfdkBFJC6_1),.clk(gclk));
	jdff dff_A_qxygZq8W6_1(.dout(w_dff_A_zfdkBFJC6_1),.din(w_dff_A_qxygZq8W6_1),.clk(gclk));
	jdff dff_A_viZejYLv6_1(.dout(w_dff_A_qxygZq8W6_1),.din(w_dff_A_viZejYLv6_1),.clk(gclk));
	jdff dff_A_xBUmBKqi3_1(.dout(w_dff_A_viZejYLv6_1),.din(w_dff_A_xBUmBKqi3_1),.clk(gclk));
	jdff dff_A_aPEOWLYQ7_1(.dout(w_dff_A_xBUmBKqi3_1),.din(w_dff_A_aPEOWLYQ7_1),.clk(gclk));
	jdff dff_A_sCnlMVHi9_2(.dout(w_n372_1[2]),.din(w_dff_A_sCnlMVHi9_2),.clk(gclk));
	jdff dff_A_O1OWSXsT9_1(.dout(w_n372_0[1]),.din(w_dff_A_O1OWSXsT9_1),.clk(gclk));
	jdff dff_A_O09Sv88N4_1(.dout(w_dff_A_O1OWSXsT9_1),.din(w_dff_A_O09Sv88N4_1),.clk(gclk));
	jdff dff_A_myC7Op7m9_1(.dout(w_dff_A_O09Sv88N4_1),.din(w_dff_A_myC7Op7m9_1),.clk(gclk));
	jdff dff_A_lVTS1oef4_1(.dout(w_dff_A_myC7Op7m9_1),.din(w_dff_A_lVTS1oef4_1),.clk(gclk));
	jdff dff_A_1F408bzs9_1(.dout(w_dff_A_lVTS1oef4_1),.din(w_dff_A_1F408bzs9_1),.clk(gclk));
	jdff dff_A_OvmsPZXt0_1(.dout(w_dff_A_1F408bzs9_1),.din(w_dff_A_OvmsPZXt0_1),.clk(gclk));
	jdff dff_A_kGUs8Ygl7_2(.dout(w_n372_0[2]),.din(w_dff_A_kGUs8Ygl7_2),.clk(gclk));
	jdff dff_A_2PKsHjju1_2(.dout(w_dff_A_kGUs8Ygl7_2),.din(w_dff_A_2PKsHjju1_2),.clk(gclk));
	jdff dff_A_O3pZ11if4_2(.dout(w_dff_A_2PKsHjju1_2),.din(w_dff_A_O3pZ11if4_2),.clk(gclk));
	jdff dff_A_G4vODcwN8_2(.dout(w_dff_A_O3pZ11if4_2),.din(w_dff_A_G4vODcwN8_2),.clk(gclk));
	jdff dff_A_BfEahovQ1_2(.dout(w_dff_A_G4vODcwN8_2),.din(w_dff_A_BfEahovQ1_2),.clk(gclk));
	jdff dff_A_IPFhCnFv0_2(.dout(w_dff_A_BfEahovQ1_2),.din(w_dff_A_IPFhCnFv0_2),.clk(gclk));
	jdff dff_A_bUV5ZSHt7_2(.dout(w_dff_A_IPFhCnFv0_2),.din(w_dff_A_bUV5ZSHt7_2),.clk(gclk));
	jdff dff_A_nvfLFF5L2_2(.dout(w_dff_A_bUV5ZSHt7_2),.din(w_dff_A_nvfLFF5L2_2),.clk(gclk));
	jdff dff_A_siTTxv4V7_1(.dout(w_G18_57[1]),.din(w_dff_A_siTTxv4V7_1),.clk(gclk));
	jdff dff_A_7OWMYmKc6_1(.dout(w_n366_0[1]),.din(w_dff_A_7OWMYmKc6_1),.clk(gclk));
	jdff dff_A_rkwUqV5s2_1(.dout(w_dff_A_7OWMYmKc6_1),.din(w_dff_A_rkwUqV5s2_1),.clk(gclk));
	jdff dff_A_A0c8EOMR5_0(.dout(w_G3723_1[0]),.din(w_dff_A_A0c8EOMR5_0),.clk(gclk));
	jdff dff_A_oT3PokxN3_0(.dout(w_dff_A_A0c8EOMR5_0),.din(w_dff_A_oT3PokxN3_0),.clk(gclk));
	jdff dff_A_WhROGiIe9_0(.dout(w_dff_A_oT3PokxN3_0),.din(w_dff_A_WhROGiIe9_0),.clk(gclk));
	jdff dff_A_9SzzS9C42_2(.dout(w_G3723_0[2]),.din(w_dff_A_9SzzS9C42_2),.clk(gclk));
	jdff dff_A_9IeOG2S09_2(.dout(w_dff_A_9SzzS9C42_2),.din(w_dff_A_9IeOG2S09_2),.clk(gclk));
	jdff dff_A_heDmG2sM6_2(.dout(w_dff_A_9IeOG2S09_2),.din(w_dff_A_heDmG2sM6_2),.clk(gclk));
	jdff dff_B_IDWVY7Qp0_0(.din(n1645),.dout(w_dff_B_IDWVY7Qp0_0),.clk(gclk));
	jdff dff_B_HKpF9qpd8_0(.din(w_dff_B_IDWVY7Qp0_0),.dout(w_dff_B_HKpF9qpd8_0),.clk(gclk));
	jdff dff_B_glvbTKBU9_0(.din(w_dff_B_HKpF9qpd8_0),.dout(w_dff_B_glvbTKBU9_0),.clk(gclk));
	jdff dff_B_M0X3wcWY0_0(.din(w_dff_B_glvbTKBU9_0),.dout(w_dff_B_M0X3wcWY0_0),.clk(gclk));
	jdff dff_B_XYYkBOti0_0(.din(w_dff_B_M0X3wcWY0_0),.dout(w_dff_B_XYYkBOti0_0),.clk(gclk));
	jdff dff_A_bxT6hRH78_0(.dout(w_n1644_0[0]),.din(w_dff_A_bxT6hRH78_0),.clk(gclk));
	jdff dff_A_n78Njfyl6_0(.dout(w_dff_A_bxT6hRH78_0),.din(w_dff_A_n78Njfyl6_0),.clk(gclk));
	jdff dff_A_c3nTc5gs1_0(.dout(w_dff_A_n78Njfyl6_0),.din(w_dff_A_c3nTc5gs1_0),.clk(gclk));
	jdff dff_A_J4TEJD776_0(.dout(w_dff_A_c3nTc5gs1_0),.din(w_dff_A_J4TEJD776_0),.clk(gclk));
	jdff dff_A_N99NFegW8_0(.dout(w_dff_A_J4TEJD776_0),.din(w_dff_A_N99NFegW8_0),.clk(gclk));
	jdff dff_A_srNQeTzb1_2(.dout(w_n1148_0[2]),.din(w_dff_A_srNQeTzb1_2),.clk(gclk));
	jdff dff_A_O97I3AvY0_2(.dout(w_dff_A_srNQeTzb1_2),.din(w_dff_A_O97I3AvY0_2),.clk(gclk));
	jdff dff_A_epmZ90cf7_2(.dout(w_dff_A_O97I3AvY0_2),.din(w_dff_A_epmZ90cf7_2),.clk(gclk));
	jdff dff_A_ORIrRChN2_2(.dout(w_dff_A_epmZ90cf7_2),.din(w_dff_A_ORIrRChN2_2),.clk(gclk));
	jdff dff_A_nkNKKBf63_2(.dout(w_dff_A_ORIrRChN2_2),.din(w_dff_A_nkNKKBf63_2),.clk(gclk));
	jdff dff_A_ua17eETB6_2(.dout(w_dff_A_nkNKKBf63_2),.din(w_dff_A_ua17eETB6_2),.clk(gclk));
	jdff dff_A_Z8dSX2lB7_2(.dout(w_n429_1[2]),.din(w_dff_A_Z8dSX2lB7_2),.clk(gclk));
	jdff dff_A_N77G8Ucv9_2(.dout(w_dff_A_Z8dSX2lB7_2),.din(w_dff_A_N77G8Ucv9_2),.clk(gclk));
	jdff dff_A_7gOmAGjr3_2(.dout(w_dff_A_N77G8Ucv9_2),.din(w_dff_A_7gOmAGjr3_2),.clk(gclk));
	jdff dff_A_ZIz1Wk376_2(.dout(w_dff_A_7gOmAGjr3_2),.din(w_dff_A_ZIz1Wk376_2),.clk(gclk));
	jdff dff_A_a9jK7E3F3_2(.dout(w_dff_A_ZIz1Wk376_2),.din(w_dff_A_a9jK7E3F3_2),.clk(gclk));
	jdff dff_A_jj0BgXic4_2(.dout(w_dff_A_a9jK7E3F3_2),.din(w_dff_A_jj0BgXic4_2),.clk(gclk));
	jdff dff_A_M2sNt5aJ0_2(.dout(w_dff_A_jj0BgXic4_2),.din(w_dff_A_M2sNt5aJ0_2),.clk(gclk));
	jdff dff_A_SuogiHgF1_2(.dout(w_dff_A_M2sNt5aJ0_2),.din(w_dff_A_SuogiHgF1_2),.clk(gclk));
	jdff dff_B_8HgM9npp3_1(.din(n1638),.dout(w_dff_B_8HgM9npp3_1),.clk(gclk));
	jdff dff_A_WQ7rGcbR6_1(.dout(w_n455_0[1]),.din(w_dff_A_WQ7rGcbR6_1),.clk(gclk));
	jdff dff_A_7KKGRqGr4_1(.dout(w_dff_A_WQ7rGcbR6_1),.din(w_dff_A_7KKGRqGr4_1),.clk(gclk));
	jdff dff_A_Eo8pjj496_0(.dout(w_n461_0[0]),.din(w_dff_A_Eo8pjj496_0),.clk(gclk));
	jdff dff_A_iiFUvMV99_1(.dout(w_n460_0[1]),.din(w_dff_A_iiFUvMV99_1),.clk(gclk));
	jdff dff_A_e9pqetUX0_1(.dout(w_dff_A_iiFUvMV99_1),.din(w_dff_A_e9pqetUX0_1),.clk(gclk));
	jdff dff_A_BI8gDIYZ4_1(.dout(w_dff_A_e9pqetUX0_1),.din(w_dff_A_BI8gDIYZ4_1),.clk(gclk));
	jdff dff_A_c1RFncXA6_1(.dout(w_dff_A_BI8gDIYZ4_1),.din(w_dff_A_c1RFncXA6_1),.clk(gclk));
	jdff dff_A_UFFdpIeU1_1(.dout(w_dff_A_c1RFncXA6_1),.din(w_dff_A_UFFdpIeU1_1),.clk(gclk));
	jdff dff_A_Ei9lQM4A3_1(.dout(w_n458_0[1]),.din(w_dff_A_Ei9lQM4A3_1),.clk(gclk));
	jdff dff_A_VNLWXNkb2_1(.dout(w_dff_A_Ei9lQM4A3_1),.din(w_dff_A_VNLWXNkb2_1),.clk(gclk));
	jdff dff_A_EnvjuNp65_1(.dout(w_dff_A_VNLWXNkb2_1),.din(w_dff_A_EnvjuNp65_1),.clk(gclk));
	jdff dff_A_UKT2WkAc4_1(.dout(w_dff_A_EnvjuNp65_1),.din(w_dff_A_UKT2WkAc4_1),.clk(gclk));
	jdff dff_A_x11vc7E51_1(.dout(w_dff_A_UKT2WkAc4_1),.din(w_dff_A_x11vc7E51_1),.clk(gclk));
	jdff dff_A_3lQu6qF98_1(.dout(w_dff_A_x11vc7E51_1),.din(w_dff_A_3lQu6qF98_1),.clk(gclk));
	jdff dff_A_v5z2xYqi5_1(.dout(w_dff_A_3lQu6qF98_1),.din(w_dff_A_v5z2xYqi5_1),.clk(gclk));
	jdff dff_A_Pa5T8Khv1_0(.dout(w_G3729_1[0]),.din(w_dff_A_Pa5T8Khv1_0),.clk(gclk));
	jdff dff_A_8LcK8OjW1_0(.dout(w_dff_A_Pa5T8Khv1_0),.din(w_dff_A_8LcK8OjW1_0),.clk(gclk));
	jdff dff_A_FABQIxU61_0(.dout(w_dff_A_8LcK8OjW1_0),.din(w_dff_A_FABQIxU61_0),.clk(gclk));
	jdff dff_A_oU161Ncu3_2(.dout(w_G3729_0[2]),.din(w_dff_A_oU161Ncu3_2),.clk(gclk));
	jdff dff_A_PsQowceb7_2(.dout(w_dff_A_oU161Ncu3_2),.din(w_dff_A_PsQowceb7_2),.clk(gclk));
	jdff dff_A_aF5AZzhG1_2(.dout(w_dff_A_PsQowceb7_2),.din(w_dff_A_aF5AZzhG1_2),.clk(gclk));
	jdff dff_B_h21CaGwJ6_1(.din(n423),.dout(w_dff_B_h21CaGwJ6_1),.clk(gclk));
	jdff dff_B_l6O1nGen5_1(.din(w_dff_B_h21CaGwJ6_1),.dout(w_dff_B_l6O1nGen5_1),.clk(gclk));
	jdff dff_B_aoQ4cO6G4_2(.din(n457),.dout(w_dff_B_aoQ4cO6G4_2),.clk(gclk));
	jdff dff_A_Ez3fDP7O2_0(.dout(w_G18_55[0]),.din(w_dff_A_Ez3fDP7O2_0),.clk(gclk));
	jdff dff_A_LnfPSjCj1_2(.dout(w_G18_55[2]),.din(w_dff_A_LnfPSjCj1_2),.clk(gclk));
	jdff dff_A_5wOY19y38_0(.dout(w_G3737_1[0]),.din(w_dff_A_5wOY19y38_0),.clk(gclk));
	jdff dff_A_TwEkicrX2_0(.dout(w_dff_A_5wOY19y38_0),.din(w_dff_A_TwEkicrX2_0),.clk(gclk));
	jdff dff_A_HfR9wvXH0_0(.dout(w_dff_A_TwEkicrX2_0),.din(w_dff_A_HfR9wvXH0_0),.clk(gclk));
	jdff dff_A_xFFZkzla9_1(.dout(w_n456_0[1]),.din(w_dff_A_xFFZkzla9_1),.clk(gclk));
	jdff dff_A_l1nYXMXi6_1(.dout(w_dff_A_xFFZkzla9_1),.din(w_dff_A_l1nYXMXi6_1),.clk(gclk));
	jdff dff_A_S887kdNf8_1(.dout(w_dff_A_l1nYXMXi6_1),.din(w_dff_A_S887kdNf8_1),.clk(gclk));
	jdff dff_A_ldZ1KY7c8_1(.dout(w_dff_A_S887kdNf8_1),.din(w_dff_A_ldZ1KY7c8_1),.clk(gclk));
	jdff dff_A_YkCQntDW9_1(.dout(w_dff_A_ldZ1KY7c8_1),.din(w_dff_A_YkCQntDW9_1),.clk(gclk));
	jdff dff_A_41bqDbRo2_1(.dout(w_dff_A_YkCQntDW9_1),.din(w_dff_A_41bqDbRo2_1),.clk(gclk));
	jdff dff_A_fSaZrFse3_2(.dout(w_n456_0[2]),.din(w_dff_A_fSaZrFse3_2),.clk(gclk));
	jdff dff_A_zlrFOdIx5_2(.dout(w_n446_0[2]),.din(w_dff_A_zlrFOdIx5_2),.clk(gclk));
	jdff dff_A_Oh7A8BMG5_2(.dout(w_dff_A_zlrFOdIx5_2),.din(w_dff_A_Oh7A8BMG5_2),.clk(gclk));
	jdff dff_A_Mbxmu5IA8_2(.dout(w_dff_A_Oh7A8BMG5_2),.din(w_dff_A_Mbxmu5IA8_2),.clk(gclk));
	jdff dff_A_7nHzeAQE8_0(.dout(w_n445_0[0]),.din(w_dff_A_7nHzeAQE8_0),.clk(gclk));
	jdff dff_A_i8MxtEqX8_0(.dout(w_dff_A_7nHzeAQE8_0),.din(w_dff_A_i8MxtEqX8_0),.clk(gclk));
	jdff dff_A_gJo61eAj1_0(.dout(w_dff_A_i8MxtEqX8_0),.din(w_dff_A_gJo61eAj1_0),.clk(gclk));
	jdff dff_A_jCSaDnGt3_0(.dout(w_dff_A_gJo61eAj1_0),.din(w_dff_A_jCSaDnGt3_0),.clk(gclk));
	jdff dff_B_PlwNksKA7_2(.din(n445),.dout(w_dff_B_PlwNksKA7_2),.clk(gclk));
	jdff dff_A_UiYgcqjj0_0(.dout(w_n443_0[0]),.din(w_dff_A_UiYgcqjj0_0),.clk(gclk));
	jdff dff_A_4K5YfUEq1_0(.dout(w_dff_A_UiYgcqjj0_0),.din(w_dff_A_4K5YfUEq1_0),.clk(gclk));
	jdff dff_A_qYFnchSb5_0(.dout(w_dff_A_4K5YfUEq1_0),.din(w_dff_A_qYFnchSb5_0),.clk(gclk));
	jdff dff_A_qg2u1FFT9_0(.dout(w_dff_A_qYFnchSb5_0),.din(w_dff_A_qg2u1FFT9_0),.clk(gclk));
	jdff dff_A_NME46QeS8_1(.dout(w_G18_54[1]),.din(w_dff_A_NME46QeS8_1),.clk(gclk));
	jdff dff_A_hrTl2yRI2_0(.dout(w_G3749_0[0]),.din(w_dff_A_hrTl2yRI2_0),.clk(gclk));
	jdff dff_A_ZBdNzVag3_0(.dout(w_dff_A_hrTl2yRI2_0),.din(w_dff_A_ZBdNzVag3_0),.clk(gclk));
	jdff dff_A_6QumpSRY2_0(.dout(w_dff_A_ZBdNzVag3_0),.din(w_dff_A_6QumpSRY2_0),.clk(gclk));
	jdff dff_A_zAZyEvqU4_1(.dout(w_n450_0[1]),.din(w_dff_A_zAZyEvqU4_1),.clk(gclk));
	jdff dff_A_S2y8jGwy7_1(.dout(w_dff_A_zAZyEvqU4_1),.din(w_dff_A_S2y8jGwy7_1),.clk(gclk));
	jdff dff_A_eBkTexpT7_1(.dout(w_dff_A_S2y8jGwy7_1),.din(w_dff_A_eBkTexpT7_1),.clk(gclk));
	jdff dff_A_1GyyuEdD3_1(.dout(w_dff_A_eBkTexpT7_1),.din(w_dff_A_1GyyuEdD3_1),.clk(gclk));
	jdff dff_A_7Jc62E2n3_1(.dout(w_dff_A_1GyyuEdD3_1),.din(w_dff_A_7Jc62E2n3_1),.clk(gclk));
	jdff dff_A_Pgbhg1V60_1(.dout(w_dff_A_7Jc62E2n3_1),.din(w_dff_A_Pgbhg1V60_1),.clk(gclk));
	jdff dff_A_yGPNZGOU3_1(.dout(w_dff_A_Pgbhg1V60_1),.din(w_dff_A_yGPNZGOU3_1),.clk(gclk));
	jdff dff_A_DQ9xXhsI5_2(.dout(w_n450_0[2]),.din(w_dff_A_DQ9xXhsI5_2),.clk(gclk));
	jdff dff_B_JFMYzIFG6_3(.din(n450),.dout(w_dff_B_JFMYzIFG6_3),.clk(gclk));
	jdff dff_B_44dd0rRk9_1(.din(n447),.dout(w_dff_B_44dd0rRk9_1),.clk(gclk));
	jdff dff_B_hcyQBnBz9_0(.din(G124),.dout(w_dff_B_hcyQBnBz9_0),.clk(gclk));
	jdff dff_A_JffuGsQJ7_2(.dout(w_G18_58[2]),.din(w_dff_A_JffuGsQJ7_2),.clk(gclk));
	jdff dff_A_cXHyq6OK4_1(.dout(w_G18_6[1]),.din(w_dff_A_cXHyq6OK4_1),.clk(gclk));
	jdff dff_A_984qphLh4_2(.dout(w_G18_6[2]),.din(w_dff_A_984qphLh4_2),.clk(gclk));
	jdff dff_A_n0yhwvps7_2(.dout(w_G18_53[2]),.din(w_dff_A_n0yhwvps7_2),.clk(gclk));
	jdff dff_A_yxDm7fX93_0(.dout(w_G3743_1[0]),.din(w_dff_A_yxDm7fX93_0),.clk(gclk));
	jdff dff_A_j8emn42k0_1(.dout(w_G3743_1[1]),.din(w_dff_A_j8emn42k0_1),.clk(gclk));
	jdff dff_A_Mop6iPGY8_0(.dout(w_G3743_0[0]),.din(w_dff_A_Mop6iPGY8_0),.clk(gclk));
	jdff dff_A_WIVPdZkN8_0(.dout(w_dff_A_Mop6iPGY8_0),.din(w_dff_A_WIVPdZkN8_0),.clk(gclk));
	jdff dff_A_vVahhG232_0(.dout(w_dff_A_WIVPdZkN8_0),.din(w_dff_A_vVahhG232_0),.clk(gclk));
	jdff dff_A_hSoXGY9p8_1(.dout(w_n1360_0[1]),.din(w_dff_A_hSoXGY9p8_1),.clk(gclk));
	jdff dff_A_rsI4cXCp7_2(.dout(w_n387_0[2]),.din(w_dff_A_rsI4cXCp7_2),.clk(gclk));
	jdff dff_A_s7ItAJyX3_2(.dout(w_dff_A_rsI4cXCp7_2),.din(w_dff_A_s7ItAJyX3_2),.clk(gclk));
	jdff dff_A_EagitJIb6_2(.dout(w_dff_A_s7ItAJyX3_2),.din(w_dff_A_EagitJIb6_2),.clk(gclk));
	jdff dff_A_GOOt5XX88_2(.dout(w_dff_A_EagitJIb6_2),.din(w_dff_A_GOOt5XX88_2),.clk(gclk));
	jdff dff_B_8A4vRwvi3_1(.din(n381),.dout(w_dff_B_8A4vRwvi3_1),.clk(gclk));
	jdff dff_B_Lmpe7ff84_1(.din(w_dff_B_8A4vRwvi3_1),.dout(w_dff_B_Lmpe7ff84_1),.clk(gclk));
	jdff dff_A_g8Yd2so27_0(.dout(w_G18_56[0]),.din(w_dff_A_g8Yd2so27_0),.clk(gclk));
	jdff dff_A_e7OVtupO2_2(.dout(w_G18_56[2]),.din(w_dff_A_e7OVtupO2_2),.clk(gclk));
	jdff dff_A_DIwKuMg99_0(.dout(w_G3711_1[0]),.din(w_dff_A_DIwKuMg99_0),.clk(gclk));
	jdff dff_A_7OXfBqVa7_0(.dout(w_dff_A_DIwKuMg99_0),.din(w_dff_A_7OXfBqVa7_0),.clk(gclk));
	jdff dff_A_nDhm2kq96_0(.dout(w_dff_A_7OXfBqVa7_0),.din(w_dff_A_nDhm2kq96_0),.clk(gclk));
	jdff dff_A_Lj9zbcUa6_1(.dout(w_dff_A_ywehXCUa1_0),.din(w_dff_A_Lj9zbcUa6_1),.clk(gclk));
	jdff dff_A_ywehXCUa1_0(.dout(w_dff_A_hpZHBmGS3_0),.din(w_dff_A_ywehXCUa1_0),.clk(gclk));
	jdff dff_A_hpZHBmGS3_0(.dout(w_dff_A_sfSARdCR5_0),.din(w_dff_A_hpZHBmGS3_0),.clk(gclk));
	jdff dff_A_sfSARdCR5_0(.dout(w_dff_A_nBd1YF5H6_0),.din(w_dff_A_sfSARdCR5_0),.clk(gclk));
	jdff dff_A_nBd1YF5H6_0(.dout(w_dff_A_M3jxpyfz4_0),.din(w_dff_A_nBd1YF5H6_0),.clk(gclk));
	jdff dff_A_M3jxpyfz4_0(.dout(w_dff_A_PFYmG4hZ5_0),.din(w_dff_A_M3jxpyfz4_0),.clk(gclk));
	jdff dff_A_PFYmG4hZ5_0(.dout(w_dff_A_eiOEw5107_0),.din(w_dff_A_PFYmG4hZ5_0),.clk(gclk));
	jdff dff_A_eiOEw5107_0(.dout(w_dff_A_YXbuUOnv8_0),.din(w_dff_A_eiOEw5107_0),.clk(gclk));
	jdff dff_A_YXbuUOnv8_0(.dout(w_dff_A_XCVPSGM95_0),.din(w_dff_A_YXbuUOnv8_0),.clk(gclk));
	jdff dff_A_XCVPSGM95_0(.dout(w_dff_A_ZX6fe0lf9_0),.din(w_dff_A_XCVPSGM95_0),.clk(gclk));
	jdff dff_A_ZX6fe0lf9_0(.dout(w_dff_A_uWzz0TLL9_0),.din(w_dff_A_ZX6fe0lf9_0),.clk(gclk));
	jdff dff_A_uWzz0TLL9_0(.dout(w_dff_A_EfuQuOuc9_0),.din(w_dff_A_uWzz0TLL9_0),.clk(gclk));
	jdff dff_A_EfuQuOuc9_0(.dout(w_dff_A_hgvHOupC1_0),.din(w_dff_A_EfuQuOuc9_0),.clk(gclk));
	jdff dff_A_hgvHOupC1_0(.dout(w_dff_A_wtqYKzGc1_0),.din(w_dff_A_hgvHOupC1_0),.clk(gclk));
	jdff dff_A_wtqYKzGc1_0(.dout(w_dff_A_7XduDj1U7_0),.din(w_dff_A_wtqYKzGc1_0),.clk(gclk));
	jdff dff_A_7XduDj1U7_0(.dout(w_dff_A_A7GNF2XS4_0),.din(w_dff_A_7XduDj1U7_0),.clk(gclk));
	jdff dff_A_A7GNF2XS4_0(.dout(w_dff_A_CEmI8Lxr6_0),.din(w_dff_A_A7GNF2XS4_0),.clk(gclk));
	jdff dff_A_CEmI8Lxr6_0(.dout(w_dff_A_5PrQnNSk7_0),.din(w_dff_A_CEmI8Lxr6_0),.clk(gclk));
	jdff dff_A_5PrQnNSk7_0(.dout(w_dff_A_2sPFJEsh9_0),.din(w_dff_A_5PrQnNSk7_0),.clk(gclk));
	jdff dff_A_2sPFJEsh9_0(.dout(w_dff_A_9b6dwdyC6_0),.din(w_dff_A_2sPFJEsh9_0),.clk(gclk));
	jdff dff_A_9b6dwdyC6_0(.dout(w_dff_A_aZWE634o2_0),.din(w_dff_A_9b6dwdyC6_0),.clk(gclk));
	jdff dff_A_aZWE634o2_0(.dout(w_dff_A_BEWgpPnm6_0),.din(w_dff_A_aZWE634o2_0),.clk(gclk));
	jdff dff_A_BEWgpPnm6_0(.dout(w_dff_A_MNU1QNoV9_0),.din(w_dff_A_BEWgpPnm6_0),.clk(gclk));
	jdff dff_A_MNU1QNoV9_0(.dout(w_dff_A_LX11k00f7_0),.din(w_dff_A_MNU1QNoV9_0),.clk(gclk));
	jdff dff_A_LX11k00f7_0(.dout(w_dff_A_iNnnpCsJ0_0),.din(w_dff_A_LX11k00f7_0),.clk(gclk));
	jdff dff_A_iNnnpCsJ0_0(.dout(G2),.din(w_dff_A_iNnnpCsJ0_0),.clk(gclk));
	jdff dff_A_bKUyBodi8_1(.dout(w_dff_A_v285L7xL5_0),.din(w_dff_A_bKUyBodi8_1),.clk(gclk));
	jdff dff_A_v285L7xL5_0(.dout(w_dff_A_rUDYX13a7_0),.din(w_dff_A_v285L7xL5_0),.clk(gclk));
	jdff dff_A_rUDYX13a7_0(.dout(w_dff_A_4tDnO5nJ5_0),.din(w_dff_A_rUDYX13a7_0),.clk(gclk));
	jdff dff_A_4tDnO5nJ5_0(.dout(w_dff_A_h0o3o1xr8_0),.din(w_dff_A_4tDnO5nJ5_0),.clk(gclk));
	jdff dff_A_h0o3o1xr8_0(.dout(w_dff_A_OYeP2yOu7_0),.din(w_dff_A_h0o3o1xr8_0),.clk(gclk));
	jdff dff_A_OYeP2yOu7_0(.dout(w_dff_A_uKTFaQJ35_0),.din(w_dff_A_OYeP2yOu7_0),.clk(gclk));
	jdff dff_A_uKTFaQJ35_0(.dout(w_dff_A_eUrAMSmT5_0),.din(w_dff_A_uKTFaQJ35_0),.clk(gclk));
	jdff dff_A_eUrAMSmT5_0(.dout(w_dff_A_yHDXYlgH7_0),.din(w_dff_A_eUrAMSmT5_0),.clk(gclk));
	jdff dff_A_yHDXYlgH7_0(.dout(w_dff_A_TMxFEqwz9_0),.din(w_dff_A_yHDXYlgH7_0),.clk(gclk));
	jdff dff_A_TMxFEqwz9_0(.dout(w_dff_A_tVliGP8n1_0),.din(w_dff_A_TMxFEqwz9_0),.clk(gclk));
	jdff dff_A_tVliGP8n1_0(.dout(w_dff_A_nt2KtYtx8_0),.din(w_dff_A_tVliGP8n1_0),.clk(gclk));
	jdff dff_A_nt2KtYtx8_0(.dout(w_dff_A_8p4nqR3a8_0),.din(w_dff_A_nt2KtYtx8_0),.clk(gclk));
	jdff dff_A_8p4nqR3a8_0(.dout(w_dff_A_BKsLBISq9_0),.din(w_dff_A_8p4nqR3a8_0),.clk(gclk));
	jdff dff_A_BKsLBISq9_0(.dout(w_dff_A_YZsBBmMq7_0),.din(w_dff_A_BKsLBISq9_0),.clk(gclk));
	jdff dff_A_YZsBBmMq7_0(.dout(w_dff_A_lSdz3bWj1_0),.din(w_dff_A_YZsBBmMq7_0),.clk(gclk));
	jdff dff_A_lSdz3bWj1_0(.dout(w_dff_A_C3PejpNi8_0),.din(w_dff_A_lSdz3bWj1_0),.clk(gclk));
	jdff dff_A_C3PejpNi8_0(.dout(w_dff_A_1tqrNl0d8_0),.din(w_dff_A_C3PejpNi8_0),.clk(gclk));
	jdff dff_A_1tqrNl0d8_0(.dout(w_dff_A_7dJI4oOY1_0),.din(w_dff_A_1tqrNl0d8_0),.clk(gclk));
	jdff dff_A_7dJI4oOY1_0(.dout(w_dff_A_JG1vOCvW3_0),.din(w_dff_A_7dJI4oOY1_0),.clk(gclk));
	jdff dff_A_JG1vOCvW3_0(.dout(w_dff_A_MdcULH4j6_0),.din(w_dff_A_JG1vOCvW3_0),.clk(gclk));
	jdff dff_A_MdcULH4j6_0(.dout(w_dff_A_rnzCGt0E3_0),.din(w_dff_A_MdcULH4j6_0),.clk(gclk));
	jdff dff_A_rnzCGt0E3_0(.dout(w_dff_A_LpNmMvXA5_0),.din(w_dff_A_rnzCGt0E3_0),.clk(gclk));
	jdff dff_A_LpNmMvXA5_0(.dout(w_dff_A_8pPVXDib0_0),.din(w_dff_A_LpNmMvXA5_0),.clk(gclk));
	jdff dff_A_8pPVXDib0_0(.dout(w_dff_A_wOKaWCPZ0_0),.din(w_dff_A_8pPVXDib0_0),.clk(gclk));
	jdff dff_A_wOKaWCPZ0_0(.dout(w_dff_A_4RoSXpPO6_0),.din(w_dff_A_wOKaWCPZ0_0),.clk(gclk));
	jdff dff_A_4RoSXpPO6_0(.dout(G3),.din(w_dff_A_4RoSXpPO6_0),.clk(gclk));
	jdff dff_A_ykkR7BTX5_1(.dout(w_dff_A_EpDTHM1d0_0),.din(w_dff_A_ykkR7BTX5_1),.clk(gclk));
	jdff dff_A_EpDTHM1d0_0(.dout(w_dff_A_brZ3xIhE2_0),.din(w_dff_A_EpDTHM1d0_0),.clk(gclk));
	jdff dff_A_brZ3xIhE2_0(.dout(w_dff_A_mqLJ9KNt3_0),.din(w_dff_A_brZ3xIhE2_0),.clk(gclk));
	jdff dff_A_mqLJ9KNt3_0(.dout(w_dff_A_ToyAXf8w3_0),.din(w_dff_A_mqLJ9KNt3_0),.clk(gclk));
	jdff dff_A_ToyAXf8w3_0(.dout(w_dff_A_LuN51aD65_0),.din(w_dff_A_ToyAXf8w3_0),.clk(gclk));
	jdff dff_A_LuN51aD65_0(.dout(w_dff_A_XH5w1yxR1_0),.din(w_dff_A_LuN51aD65_0),.clk(gclk));
	jdff dff_A_XH5w1yxR1_0(.dout(w_dff_A_3nAWI0la7_0),.din(w_dff_A_XH5w1yxR1_0),.clk(gclk));
	jdff dff_A_3nAWI0la7_0(.dout(w_dff_A_ZRPZAtOX5_0),.din(w_dff_A_3nAWI0la7_0),.clk(gclk));
	jdff dff_A_ZRPZAtOX5_0(.dout(w_dff_A_c7HJVQT50_0),.din(w_dff_A_ZRPZAtOX5_0),.clk(gclk));
	jdff dff_A_c7HJVQT50_0(.dout(w_dff_A_7wrTDaOS1_0),.din(w_dff_A_c7HJVQT50_0),.clk(gclk));
	jdff dff_A_7wrTDaOS1_0(.dout(w_dff_A_VAz7b4Gi5_0),.din(w_dff_A_7wrTDaOS1_0),.clk(gclk));
	jdff dff_A_VAz7b4Gi5_0(.dout(w_dff_A_6SFwqig01_0),.din(w_dff_A_VAz7b4Gi5_0),.clk(gclk));
	jdff dff_A_6SFwqig01_0(.dout(w_dff_A_IOVpHB1G7_0),.din(w_dff_A_6SFwqig01_0),.clk(gclk));
	jdff dff_A_IOVpHB1G7_0(.dout(w_dff_A_RyEOauqP4_0),.din(w_dff_A_IOVpHB1G7_0),.clk(gclk));
	jdff dff_A_RyEOauqP4_0(.dout(w_dff_A_6ZTgUnNV6_0),.din(w_dff_A_RyEOauqP4_0),.clk(gclk));
	jdff dff_A_6ZTgUnNV6_0(.dout(w_dff_A_VThvqpi84_0),.din(w_dff_A_6ZTgUnNV6_0),.clk(gclk));
	jdff dff_A_VThvqpi84_0(.dout(w_dff_A_K5pe7vPB7_0),.din(w_dff_A_VThvqpi84_0),.clk(gclk));
	jdff dff_A_K5pe7vPB7_0(.dout(w_dff_A_K3AtxB7M4_0),.din(w_dff_A_K5pe7vPB7_0),.clk(gclk));
	jdff dff_A_K3AtxB7M4_0(.dout(w_dff_A_A9TpM5qa7_0),.din(w_dff_A_K3AtxB7M4_0),.clk(gclk));
	jdff dff_A_A9TpM5qa7_0(.dout(w_dff_A_jhEdUKFC0_0),.din(w_dff_A_A9TpM5qa7_0),.clk(gclk));
	jdff dff_A_jhEdUKFC0_0(.dout(w_dff_A_Coq6BMl46_0),.din(w_dff_A_jhEdUKFC0_0),.clk(gclk));
	jdff dff_A_Coq6BMl46_0(.dout(w_dff_A_hv1lnQ6D7_0),.din(w_dff_A_Coq6BMl46_0),.clk(gclk));
	jdff dff_A_hv1lnQ6D7_0(.dout(w_dff_A_AVvk53uu6_0),.din(w_dff_A_hv1lnQ6D7_0),.clk(gclk));
	jdff dff_A_AVvk53uu6_0(.dout(w_dff_A_zRW9CPGS3_0),.din(w_dff_A_AVvk53uu6_0),.clk(gclk));
	jdff dff_A_zRW9CPGS3_0(.dout(w_dff_A_teD8M2gk8_0),.din(w_dff_A_zRW9CPGS3_0),.clk(gclk));
	jdff dff_A_teD8M2gk8_0(.dout(G450),.din(w_dff_A_teD8M2gk8_0),.clk(gclk));
	jdff dff_A_5BZl4JPk1_1(.dout(w_dff_A_PIJL7jhG7_0),.din(w_dff_A_5BZl4JPk1_1),.clk(gclk));
	jdff dff_A_PIJL7jhG7_0(.dout(w_dff_A_FnQYp6ul2_0),.din(w_dff_A_PIJL7jhG7_0),.clk(gclk));
	jdff dff_A_FnQYp6ul2_0(.dout(w_dff_A_i4X35nkB3_0),.din(w_dff_A_FnQYp6ul2_0),.clk(gclk));
	jdff dff_A_i4X35nkB3_0(.dout(w_dff_A_X1aQbOx61_0),.din(w_dff_A_i4X35nkB3_0),.clk(gclk));
	jdff dff_A_X1aQbOx61_0(.dout(w_dff_A_Tz9Ll54v1_0),.din(w_dff_A_X1aQbOx61_0),.clk(gclk));
	jdff dff_A_Tz9Ll54v1_0(.dout(w_dff_A_N9m2u4dY9_0),.din(w_dff_A_Tz9Ll54v1_0),.clk(gclk));
	jdff dff_A_N9m2u4dY9_0(.dout(w_dff_A_xSNJ1BTN8_0),.din(w_dff_A_N9m2u4dY9_0),.clk(gclk));
	jdff dff_A_xSNJ1BTN8_0(.dout(w_dff_A_4kKgQLrM4_0),.din(w_dff_A_xSNJ1BTN8_0),.clk(gclk));
	jdff dff_A_4kKgQLrM4_0(.dout(w_dff_A_h1PCNJ8L1_0),.din(w_dff_A_4kKgQLrM4_0),.clk(gclk));
	jdff dff_A_h1PCNJ8L1_0(.dout(w_dff_A_LWfeLkUz3_0),.din(w_dff_A_h1PCNJ8L1_0),.clk(gclk));
	jdff dff_A_LWfeLkUz3_0(.dout(w_dff_A_XFMDUF8M2_0),.din(w_dff_A_LWfeLkUz3_0),.clk(gclk));
	jdff dff_A_XFMDUF8M2_0(.dout(w_dff_A_USC1GW618_0),.din(w_dff_A_XFMDUF8M2_0),.clk(gclk));
	jdff dff_A_USC1GW618_0(.dout(w_dff_A_f0pTPOsW2_0),.din(w_dff_A_USC1GW618_0),.clk(gclk));
	jdff dff_A_f0pTPOsW2_0(.dout(w_dff_A_6dARqQ2a3_0),.din(w_dff_A_f0pTPOsW2_0),.clk(gclk));
	jdff dff_A_6dARqQ2a3_0(.dout(w_dff_A_svgvGrkX3_0),.din(w_dff_A_6dARqQ2a3_0),.clk(gclk));
	jdff dff_A_svgvGrkX3_0(.dout(w_dff_A_qZKJUXgl6_0),.din(w_dff_A_svgvGrkX3_0),.clk(gclk));
	jdff dff_A_qZKJUXgl6_0(.dout(w_dff_A_aw2zk8MI0_0),.din(w_dff_A_qZKJUXgl6_0),.clk(gclk));
	jdff dff_A_aw2zk8MI0_0(.dout(w_dff_A_FnH9o1Tb4_0),.din(w_dff_A_aw2zk8MI0_0),.clk(gclk));
	jdff dff_A_FnH9o1Tb4_0(.dout(w_dff_A_eOlFEr7z1_0),.din(w_dff_A_FnH9o1Tb4_0),.clk(gclk));
	jdff dff_A_eOlFEr7z1_0(.dout(w_dff_A_bVOZMBm67_0),.din(w_dff_A_eOlFEr7z1_0),.clk(gclk));
	jdff dff_A_bVOZMBm67_0(.dout(w_dff_A_14yrAvKb5_0),.din(w_dff_A_bVOZMBm67_0),.clk(gclk));
	jdff dff_A_14yrAvKb5_0(.dout(w_dff_A_lkSNs8He8_0),.din(w_dff_A_14yrAvKb5_0),.clk(gclk));
	jdff dff_A_lkSNs8He8_0(.dout(w_dff_A_vvfK3lCp9_0),.din(w_dff_A_lkSNs8He8_0),.clk(gclk));
	jdff dff_A_vvfK3lCp9_0(.dout(w_dff_A_v2yELCdE9_0),.din(w_dff_A_vvfK3lCp9_0),.clk(gclk));
	jdff dff_A_v2yELCdE9_0(.dout(w_dff_A_3PEnCtBv8_0),.din(w_dff_A_v2yELCdE9_0),.clk(gclk));
	jdff dff_A_3PEnCtBv8_0(.dout(G448),.din(w_dff_A_3PEnCtBv8_0),.clk(gclk));
	jdff dff_A_lpzyHoCB3_1(.dout(w_dff_A_oDbiegJ57_0),.din(w_dff_A_lpzyHoCB3_1),.clk(gclk));
	jdff dff_A_oDbiegJ57_0(.dout(w_dff_A_Hhzsciea1_0),.din(w_dff_A_oDbiegJ57_0),.clk(gclk));
	jdff dff_A_Hhzsciea1_0(.dout(w_dff_A_YwcUCT5Z8_0),.din(w_dff_A_Hhzsciea1_0),.clk(gclk));
	jdff dff_A_YwcUCT5Z8_0(.dout(w_dff_A_n817RTmT7_0),.din(w_dff_A_YwcUCT5Z8_0),.clk(gclk));
	jdff dff_A_n817RTmT7_0(.dout(w_dff_A_nxrsyCh59_0),.din(w_dff_A_n817RTmT7_0),.clk(gclk));
	jdff dff_A_nxrsyCh59_0(.dout(w_dff_A_7voHvPDZ3_0),.din(w_dff_A_nxrsyCh59_0),.clk(gclk));
	jdff dff_A_7voHvPDZ3_0(.dout(w_dff_A_UqJ05x1V3_0),.din(w_dff_A_7voHvPDZ3_0),.clk(gclk));
	jdff dff_A_UqJ05x1V3_0(.dout(w_dff_A_5n1Pyn2d8_0),.din(w_dff_A_UqJ05x1V3_0),.clk(gclk));
	jdff dff_A_5n1Pyn2d8_0(.dout(w_dff_A_u8dNkfQO1_0),.din(w_dff_A_5n1Pyn2d8_0),.clk(gclk));
	jdff dff_A_u8dNkfQO1_0(.dout(w_dff_A_1yUxlyNT3_0),.din(w_dff_A_u8dNkfQO1_0),.clk(gclk));
	jdff dff_A_1yUxlyNT3_0(.dout(w_dff_A_0N75zwGr0_0),.din(w_dff_A_1yUxlyNT3_0),.clk(gclk));
	jdff dff_A_0N75zwGr0_0(.dout(w_dff_A_1rln8GPN5_0),.din(w_dff_A_0N75zwGr0_0),.clk(gclk));
	jdff dff_A_1rln8GPN5_0(.dout(w_dff_A_9yOpdUW36_0),.din(w_dff_A_1rln8GPN5_0),.clk(gclk));
	jdff dff_A_9yOpdUW36_0(.dout(w_dff_A_FdeNCbK17_0),.din(w_dff_A_9yOpdUW36_0),.clk(gclk));
	jdff dff_A_FdeNCbK17_0(.dout(w_dff_A_SWqyt6at7_0),.din(w_dff_A_FdeNCbK17_0),.clk(gclk));
	jdff dff_A_SWqyt6at7_0(.dout(w_dff_A_JZ3Vvpni9_0),.din(w_dff_A_SWqyt6at7_0),.clk(gclk));
	jdff dff_A_JZ3Vvpni9_0(.dout(w_dff_A_i8ZCNfUd9_0),.din(w_dff_A_JZ3Vvpni9_0),.clk(gclk));
	jdff dff_A_i8ZCNfUd9_0(.dout(w_dff_A_0lmWSpFa0_0),.din(w_dff_A_i8ZCNfUd9_0),.clk(gclk));
	jdff dff_A_0lmWSpFa0_0(.dout(w_dff_A_3j3Lnv4x0_0),.din(w_dff_A_0lmWSpFa0_0),.clk(gclk));
	jdff dff_A_3j3Lnv4x0_0(.dout(w_dff_A_fqLPO4jp5_0),.din(w_dff_A_3j3Lnv4x0_0),.clk(gclk));
	jdff dff_A_fqLPO4jp5_0(.dout(w_dff_A_y7pZHwE02_0),.din(w_dff_A_fqLPO4jp5_0),.clk(gclk));
	jdff dff_A_y7pZHwE02_0(.dout(w_dff_A_sUDznM3e7_0),.din(w_dff_A_y7pZHwE02_0),.clk(gclk));
	jdff dff_A_sUDznM3e7_0(.dout(w_dff_A_4KUrw3ax4_0),.din(w_dff_A_sUDznM3e7_0),.clk(gclk));
	jdff dff_A_4KUrw3ax4_0(.dout(w_dff_A_9XzUPOPa3_0),.din(w_dff_A_4KUrw3ax4_0),.clk(gclk));
	jdff dff_A_9XzUPOPa3_0(.dout(w_dff_A_LrxXiihK5_0),.din(w_dff_A_9XzUPOPa3_0),.clk(gclk));
	jdff dff_A_LrxXiihK5_0(.dout(G444),.din(w_dff_A_LrxXiihK5_0),.clk(gclk));
	jdff dff_A_rEh14yc44_1(.dout(w_dff_A_WHwPWy2u7_0),.din(w_dff_A_rEh14yc44_1),.clk(gclk));
	jdff dff_A_WHwPWy2u7_0(.dout(w_dff_A_u3PY3FCf3_0),.din(w_dff_A_WHwPWy2u7_0),.clk(gclk));
	jdff dff_A_u3PY3FCf3_0(.dout(w_dff_A_IAxjzWOd2_0),.din(w_dff_A_u3PY3FCf3_0),.clk(gclk));
	jdff dff_A_IAxjzWOd2_0(.dout(w_dff_A_tkmeiAQe7_0),.din(w_dff_A_IAxjzWOd2_0),.clk(gclk));
	jdff dff_A_tkmeiAQe7_0(.dout(w_dff_A_E7tDs0jO9_0),.din(w_dff_A_tkmeiAQe7_0),.clk(gclk));
	jdff dff_A_E7tDs0jO9_0(.dout(w_dff_A_PvvokCLV7_0),.din(w_dff_A_E7tDs0jO9_0),.clk(gclk));
	jdff dff_A_PvvokCLV7_0(.dout(w_dff_A_UjGj5Ycc8_0),.din(w_dff_A_PvvokCLV7_0),.clk(gclk));
	jdff dff_A_UjGj5Ycc8_0(.dout(w_dff_A_1F61HQYx6_0),.din(w_dff_A_UjGj5Ycc8_0),.clk(gclk));
	jdff dff_A_1F61HQYx6_0(.dout(w_dff_A_ixNBkNpN0_0),.din(w_dff_A_1F61HQYx6_0),.clk(gclk));
	jdff dff_A_ixNBkNpN0_0(.dout(w_dff_A_VrxocDes2_0),.din(w_dff_A_ixNBkNpN0_0),.clk(gclk));
	jdff dff_A_VrxocDes2_0(.dout(w_dff_A_wT6ECk2p1_0),.din(w_dff_A_VrxocDes2_0),.clk(gclk));
	jdff dff_A_wT6ECk2p1_0(.dout(w_dff_A_Oq07xbS00_0),.din(w_dff_A_wT6ECk2p1_0),.clk(gclk));
	jdff dff_A_Oq07xbS00_0(.dout(w_dff_A_2CA241fZ3_0),.din(w_dff_A_Oq07xbS00_0),.clk(gclk));
	jdff dff_A_2CA241fZ3_0(.dout(w_dff_A_nDr6tM732_0),.din(w_dff_A_2CA241fZ3_0),.clk(gclk));
	jdff dff_A_nDr6tM732_0(.dout(w_dff_A_zvMdIWmt8_0),.din(w_dff_A_nDr6tM732_0),.clk(gclk));
	jdff dff_A_zvMdIWmt8_0(.dout(w_dff_A_0BcZrKz53_0),.din(w_dff_A_zvMdIWmt8_0),.clk(gclk));
	jdff dff_A_0BcZrKz53_0(.dout(w_dff_A_XcAMIdEi2_0),.din(w_dff_A_0BcZrKz53_0),.clk(gclk));
	jdff dff_A_XcAMIdEi2_0(.dout(w_dff_A_EK9vnq0r5_0),.din(w_dff_A_XcAMIdEi2_0),.clk(gclk));
	jdff dff_A_EK9vnq0r5_0(.dout(w_dff_A_M64VN9N93_0),.din(w_dff_A_EK9vnq0r5_0),.clk(gclk));
	jdff dff_A_M64VN9N93_0(.dout(w_dff_A_PXIRguxK4_0),.din(w_dff_A_M64VN9N93_0),.clk(gclk));
	jdff dff_A_PXIRguxK4_0(.dout(w_dff_A_1dGvCvkD2_0),.din(w_dff_A_PXIRguxK4_0),.clk(gclk));
	jdff dff_A_1dGvCvkD2_0(.dout(w_dff_A_aGWXHUdU9_0),.din(w_dff_A_1dGvCvkD2_0),.clk(gclk));
	jdff dff_A_aGWXHUdU9_0(.dout(w_dff_A_oKOQuPsj7_0),.din(w_dff_A_aGWXHUdU9_0),.clk(gclk));
	jdff dff_A_oKOQuPsj7_0(.dout(w_dff_A_PMovNCDZ8_0),.din(w_dff_A_oKOQuPsj7_0),.clk(gclk));
	jdff dff_A_PMovNCDZ8_0(.dout(w_dff_A_RUro9E0k3_0),.din(w_dff_A_PMovNCDZ8_0),.clk(gclk));
	jdff dff_A_RUro9E0k3_0(.dout(G442),.din(w_dff_A_RUro9E0k3_0),.clk(gclk));
	jdff dff_A_Qb2jOS5o0_1(.dout(w_dff_A_tIWBtJn27_0),.din(w_dff_A_Qb2jOS5o0_1),.clk(gclk));
	jdff dff_A_tIWBtJn27_0(.dout(w_dff_A_OA0wYm853_0),.din(w_dff_A_tIWBtJn27_0),.clk(gclk));
	jdff dff_A_OA0wYm853_0(.dout(w_dff_A_G3QHnqgV6_0),.din(w_dff_A_OA0wYm853_0),.clk(gclk));
	jdff dff_A_G3QHnqgV6_0(.dout(w_dff_A_gFSGMReh4_0),.din(w_dff_A_G3QHnqgV6_0),.clk(gclk));
	jdff dff_A_gFSGMReh4_0(.dout(w_dff_A_XM9QDtR27_0),.din(w_dff_A_gFSGMReh4_0),.clk(gclk));
	jdff dff_A_XM9QDtR27_0(.dout(w_dff_A_F7xGfi0s8_0),.din(w_dff_A_XM9QDtR27_0),.clk(gclk));
	jdff dff_A_F7xGfi0s8_0(.dout(w_dff_A_OWvvromt7_0),.din(w_dff_A_F7xGfi0s8_0),.clk(gclk));
	jdff dff_A_OWvvromt7_0(.dout(w_dff_A_PX9v89ft9_0),.din(w_dff_A_OWvvromt7_0),.clk(gclk));
	jdff dff_A_PX9v89ft9_0(.dout(w_dff_A_piwCPmhX3_0),.din(w_dff_A_PX9v89ft9_0),.clk(gclk));
	jdff dff_A_piwCPmhX3_0(.dout(w_dff_A_NO5XX01t3_0),.din(w_dff_A_piwCPmhX3_0),.clk(gclk));
	jdff dff_A_NO5XX01t3_0(.dout(w_dff_A_5f7o3nb18_0),.din(w_dff_A_NO5XX01t3_0),.clk(gclk));
	jdff dff_A_5f7o3nb18_0(.dout(w_dff_A_2oEv4P7U4_0),.din(w_dff_A_5f7o3nb18_0),.clk(gclk));
	jdff dff_A_2oEv4P7U4_0(.dout(w_dff_A_SlzhVd5S8_0),.din(w_dff_A_2oEv4P7U4_0),.clk(gclk));
	jdff dff_A_SlzhVd5S8_0(.dout(w_dff_A_cSzB5Gr83_0),.din(w_dff_A_SlzhVd5S8_0),.clk(gclk));
	jdff dff_A_cSzB5Gr83_0(.dout(w_dff_A_t2p3AynC4_0),.din(w_dff_A_cSzB5Gr83_0),.clk(gclk));
	jdff dff_A_t2p3AynC4_0(.dout(w_dff_A_fE6VYTnp9_0),.din(w_dff_A_t2p3AynC4_0),.clk(gclk));
	jdff dff_A_fE6VYTnp9_0(.dout(w_dff_A_KIr9fKK00_0),.din(w_dff_A_fE6VYTnp9_0),.clk(gclk));
	jdff dff_A_KIr9fKK00_0(.dout(w_dff_A_rDeUE6176_0),.din(w_dff_A_KIr9fKK00_0),.clk(gclk));
	jdff dff_A_rDeUE6176_0(.dout(w_dff_A_HaGEhSji1_0),.din(w_dff_A_rDeUE6176_0),.clk(gclk));
	jdff dff_A_HaGEhSji1_0(.dout(w_dff_A_Inbqn0dD7_0),.din(w_dff_A_HaGEhSji1_0),.clk(gclk));
	jdff dff_A_Inbqn0dD7_0(.dout(w_dff_A_3q9vZQW89_0),.din(w_dff_A_Inbqn0dD7_0),.clk(gclk));
	jdff dff_A_3q9vZQW89_0(.dout(w_dff_A_IGygduFJ1_0),.din(w_dff_A_3q9vZQW89_0),.clk(gclk));
	jdff dff_A_IGygduFJ1_0(.dout(w_dff_A_Bv5RYsxJ9_0),.din(w_dff_A_IGygduFJ1_0),.clk(gclk));
	jdff dff_A_Bv5RYsxJ9_0(.dout(w_dff_A_zDxST4zS3_0),.din(w_dff_A_Bv5RYsxJ9_0),.clk(gclk));
	jdff dff_A_zDxST4zS3_0(.dout(w_dff_A_bZbRI6vH5_0),.din(w_dff_A_zDxST4zS3_0),.clk(gclk));
	jdff dff_A_bZbRI6vH5_0(.dout(G440),.din(w_dff_A_bZbRI6vH5_0),.clk(gclk));
	jdff dff_A_lmpG2qDt1_1(.dout(w_dff_A_uNDxEd1U6_0),.din(w_dff_A_lmpG2qDt1_1),.clk(gclk));
	jdff dff_A_uNDxEd1U6_0(.dout(w_dff_A_goDTdAAp2_0),.din(w_dff_A_uNDxEd1U6_0),.clk(gclk));
	jdff dff_A_goDTdAAp2_0(.dout(w_dff_A_XRqvAbIk7_0),.din(w_dff_A_goDTdAAp2_0),.clk(gclk));
	jdff dff_A_XRqvAbIk7_0(.dout(w_dff_A_gsrNM9RN2_0),.din(w_dff_A_XRqvAbIk7_0),.clk(gclk));
	jdff dff_A_gsrNM9RN2_0(.dout(w_dff_A_guYgLIJS6_0),.din(w_dff_A_gsrNM9RN2_0),.clk(gclk));
	jdff dff_A_guYgLIJS6_0(.dout(w_dff_A_9AMwW71b3_0),.din(w_dff_A_guYgLIJS6_0),.clk(gclk));
	jdff dff_A_9AMwW71b3_0(.dout(w_dff_A_ykmvIyn41_0),.din(w_dff_A_9AMwW71b3_0),.clk(gclk));
	jdff dff_A_ykmvIyn41_0(.dout(w_dff_A_xoOlKdZ24_0),.din(w_dff_A_ykmvIyn41_0),.clk(gclk));
	jdff dff_A_xoOlKdZ24_0(.dout(w_dff_A_GburK90B9_0),.din(w_dff_A_xoOlKdZ24_0),.clk(gclk));
	jdff dff_A_GburK90B9_0(.dout(w_dff_A_OeN8qLYi2_0),.din(w_dff_A_GburK90B9_0),.clk(gclk));
	jdff dff_A_OeN8qLYi2_0(.dout(w_dff_A_EvhxFCeK1_0),.din(w_dff_A_OeN8qLYi2_0),.clk(gclk));
	jdff dff_A_EvhxFCeK1_0(.dout(w_dff_A_O203UWHR0_0),.din(w_dff_A_EvhxFCeK1_0),.clk(gclk));
	jdff dff_A_O203UWHR0_0(.dout(w_dff_A_FeU06reW0_0),.din(w_dff_A_O203UWHR0_0),.clk(gclk));
	jdff dff_A_FeU06reW0_0(.dout(w_dff_A_ZBYZw6Ck2_0),.din(w_dff_A_FeU06reW0_0),.clk(gclk));
	jdff dff_A_ZBYZw6Ck2_0(.dout(w_dff_A_KQ5R8WS64_0),.din(w_dff_A_ZBYZw6Ck2_0),.clk(gclk));
	jdff dff_A_KQ5R8WS64_0(.dout(w_dff_A_paOEspV96_0),.din(w_dff_A_KQ5R8WS64_0),.clk(gclk));
	jdff dff_A_paOEspV96_0(.dout(w_dff_A_sjJDN5VP2_0),.din(w_dff_A_paOEspV96_0),.clk(gclk));
	jdff dff_A_sjJDN5VP2_0(.dout(w_dff_A_QS5hikjm0_0),.din(w_dff_A_sjJDN5VP2_0),.clk(gclk));
	jdff dff_A_QS5hikjm0_0(.dout(w_dff_A_pS4Sz9By5_0),.din(w_dff_A_QS5hikjm0_0),.clk(gclk));
	jdff dff_A_pS4Sz9By5_0(.dout(w_dff_A_U3z2FtCz3_0),.din(w_dff_A_pS4Sz9By5_0),.clk(gclk));
	jdff dff_A_U3z2FtCz3_0(.dout(w_dff_A_FrdDRHar5_0),.din(w_dff_A_U3z2FtCz3_0),.clk(gclk));
	jdff dff_A_FrdDRHar5_0(.dout(w_dff_A_r8DucLA32_0),.din(w_dff_A_FrdDRHar5_0),.clk(gclk));
	jdff dff_A_r8DucLA32_0(.dout(w_dff_A_pX4mqxh24_0),.din(w_dff_A_r8DucLA32_0),.clk(gclk));
	jdff dff_A_pX4mqxh24_0(.dout(w_dff_A_0BrYTy6u5_0),.din(w_dff_A_pX4mqxh24_0),.clk(gclk));
	jdff dff_A_0BrYTy6u5_0(.dout(w_dff_A_6BcXm8jQ7_0),.din(w_dff_A_0BrYTy6u5_0),.clk(gclk));
	jdff dff_A_6BcXm8jQ7_0(.dout(G438),.din(w_dff_A_6BcXm8jQ7_0),.clk(gclk));
	jdff dff_A_6XQh2fku4_1(.dout(w_dff_A_refaBZnK1_0),.din(w_dff_A_6XQh2fku4_1),.clk(gclk));
	jdff dff_A_refaBZnK1_0(.dout(w_dff_A_v7pSivbv4_0),.din(w_dff_A_refaBZnK1_0),.clk(gclk));
	jdff dff_A_v7pSivbv4_0(.dout(w_dff_A_5WO8c8WX3_0),.din(w_dff_A_v7pSivbv4_0),.clk(gclk));
	jdff dff_A_5WO8c8WX3_0(.dout(w_dff_A_9ctrAMm45_0),.din(w_dff_A_5WO8c8WX3_0),.clk(gclk));
	jdff dff_A_9ctrAMm45_0(.dout(w_dff_A_XG5Z3lUp0_0),.din(w_dff_A_9ctrAMm45_0),.clk(gclk));
	jdff dff_A_XG5Z3lUp0_0(.dout(w_dff_A_mIdx8PiL0_0),.din(w_dff_A_XG5Z3lUp0_0),.clk(gclk));
	jdff dff_A_mIdx8PiL0_0(.dout(w_dff_A_s97xlK6J4_0),.din(w_dff_A_mIdx8PiL0_0),.clk(gclk));
	jdff dff_A_s97xlK6J4_0(.dout(w_dff_A_MgW2xVXs6_0),.din(w_dff_A_s97xlK6J4_0),.clk(gclk));
	jdff dff_A_MgW2xVXs6_0(.dout(w_dff_A_hYAfsJQT8_0),.din(w_dff_A_MgW2xVXs6_0),.clk(gclk));
	jdff dff_A_hYAfsJQT8_0(.dout(w_dff_A_4HD76SjN7_0),.din(w_dff_A_hYAfsJQT8_0),.clk(gclk));
	jdff dff_A_4HD76SjN7_0(.dout(w_dff_A_lmRroHVc8_0),.din(w_dff_A_4HD76SjN7_0),.clk(gclk));
	jdff dff_A_lmRroHVc8_0(.dout(w_dff_A_Y5QSLk240_0),.din(w_dff_A_lmRroHVc8_0),.clk(gclk));
	jdff dff_A_Y5QSLk240_0(.dout(w_dff_A_850XsCfT5_0),.din(w_dff_A_Y5QSLk240_0),.clk(gclk));
	jdff dff_A_850XsCfT5_0(.dout(w_dff_A_JBpYG9X07_0),.din(w_dff_A_850XsCfT5_0),.clk(gclk));
	jdff dff_A_JBpYG9X07_0(.dout(w_dff_A_WjllqeKO9_0),.din(w_dff_A_JBpYG9X07_0),.clk(gclk));
	jdff dff_A_WjllqeKO9_0(.dout(w_dff_A_i7k7jgCg0_0),.din(w_dff_A_WjllqeKO9_0),.clk(gclk));
	jdff dff_A_i7k7jgCg0_0(.dout(w_dff_A_yloCJqOE0_0),.din(w_dff_A_i7k7jgCg0_0),.clk(gclk));
	jdff dff_A_yloCJqOE0_0(.dout(w_dff_A_0OnIPhgy8_0),.din(w_dff_A_yloCJqOE0_0),.clk(gclk));
	jdff dff_A_0OnIPhgy8_0(.dout(w_dff_A_z8RBLO0Y4_0),.din(w_dff_A_0OnIPhgy8_0),.clk(gclk));
	jdff dff_A_z8RBLO0Y4_0(.dout(w_dff_A_4ecQ7nfB0_0),.din(w_dff_A_z8RBLO0Y4_0),.clk(gclk));
	jdff dff_A_4ecQ7nfB0_0(.dout(w_dff_A_3C99x4QS6_0),.din(w_dff_A_4ecQ7nfB0_0),.clk(gclk));
	jdff dff_A_3C99x4QS6_0(.dout(w_dff_A_FP1CR0gh5_0),.din(w_dff_A_3C99x4QS6_0),.clk(gclk));
	jdff dff_A_FP1CR0gh5_0(.dout(w_dff_A_xSRs55z35_0),.din(w_dff_A_FP1CR0gh5_0),.clk(gclk));
	jdff dff_A_xSRs55z35_0(.dout(w_dff_A_skyWf8pi4_0),.din(w_dff_A_xSRs55z35_0),.clk(gclk));
	jdff dff_A_skyWf8pi4_0(.dout(w_dff_A_9kzeriYN3_0),.din(w_dff_A_skyWf8pi4_0),.clk(gclk));
	jdff dff_A_9kzeriYN3_0(.dout(G496),.din(w_dff_A_9kzeriYN3_0),.clk(gclk));
	jdff dff_A_hlgqtfXa0_1(.dout(w_dff_A_tbOYvf3p0_0),.din(w_dff_A_hlgqtfXa0_1),.clk(gclk));
	jdff dff_A_tbOYvf3p0_0(.dout(w_dff_A_hLJMW56M1_0),.din(w_dff_A_tbOYvf3p0_0),.clk(gclk));
	jdff dff_A_hLJMW56M1_0(.dout(w_dff_A_dejgQg8S3_0),.din(w_dff_A_hLJMW56M1_0),.clk(gclk));
	jdff dff_A_dejgQg8S3_0(.dout(w_dff_A_ps2e0bHv0_0),.din(w_dff_A_dejgQg8S3_0),.clk(gclk));
	jdff dff_A_ps2e0bHv0_0(.dout(w_dff_A_eStmDrLs9_0),.din(w_dff_A_ps2e0bHv0_0),.clk(gclk));
	jdff dff_A_eStmDrLs9_0(.dout(w_dff_A_m7KfGna07_0),.din(w_dff_A_eStmDrLs9_0),.clk(gclk));
	jdff dff_A_m7KfGna07_0(.dout(w_dff_A_3SlH0Ty24_0),.din(w_dff_A_m7KfGna07_0),.clk(gclk));
	jdff dff_A_3SlH0Ty24_0(.dout(w_dff_A_oG9KUfTy3_0),.din(w_dff_A_3SlH0Ty24_0),.clk(gclk));
	jdff dff_A_oG9KUfTy3_0(.dout(w_dff_A_wjNvo2rN9_0),.din(w_dff_A_oG9KUfTy3_0),.clk(gclk));
	jdff dff_A_wjNvo2rN9_0(.dout(w_dff_A_2TqheRFW2_0),.din(w_dff_A_wjNvo2rN9_0),.clk(gclk));
	jdff dff_A_2TqheRFW2_0(.dout(w_dff_A_NoRlpiHW3_0),.din(w_dff_A_2TqheRFW2_0),.clk(gclk));
	jdff dff_A_NoRlpiHW3_0(.dout(w_dff_A_YGEGc6Wu1_0),.din(w_dff_A_NoRlpiHW3_0),.clk(gclk));
	jdff dff_A_YGEGc6Wu1_0(.dout(w_dff_A_4iv8EiES8_0),.din(w_dff_A_YGEGc6Wu1_0),.clk(gclk));
	jdff dff_A_4iv8EiES8_0(.dout(w_dff_A_74ndzxJd2_0),.din(w_dff_A_4iv8EiES8_0),.clk(gclk));
	jdff dff_A_74ndzxJd2_0(.dout(w_dff_A_6UgmVWUd7_0),.din(w_dff_A_74ndzxJd2_0),.clk(gclk));
	jdff dff_A_6UgmVWUd7_0(.dout(w_dff_A_BrI94TK16_0),.din(w_dff_A_6UgmVWUd7_0),.clk(gclk));
	jdff dff_A_BrI94TK16_0(.dout(w_dff_A_UKYlCVZ00_0),.din(w_dff_A_BrI94TK16_0),.clk(gclk));
	jdff dff_A_UKYlCVZ00_0(.dout(w_dff_A_0CxWStX33_0),.din(w_dff_A_UKYlCVZ00_0),.clk(gclk));
	jdff dff_A_0CxWStX33_0(.dout(w_dff_A_1cE0Kbcx5_0),.din(w_dff_A_0CxWStX33_0),.clk(gclk));
	jdff dff_A_1cE0Kbcx5_0(.dout(w_dff_A_Bc9wqrlK4_0),.din(w_dff_A_1cE0Kbcx5_0),.clk(gclk));
	jdff dff_A_Bc9wqrlK4_0(.dout(w_dff_A_pgItJNNg9_0),.din(w_dff_A_Bc9wqrlK4_0),.clk(gclk));
	jdff dff_A_pgItJNNg9_0(.dout(w_dff_A_CTE9SC373_0),.din(w_dff_A_pgItJNNg9_0),.clk(gclk));
	jdff dff_A_CTE9SC373_0(.dout(w_dff_A_0b5GBUFN6_0),.din(w_dff_A_CTE9SC373_0),.clk(gclk));
	jdff dff_A_0b5GBUFN6_0(.dout(w_dff_A_iTnffcDf9_0),.din(w_dff_A_0b5GBUFN6_0),.clk(gclk));
	jdff dff_A_iTnffcDf9_0(.dout(w_dff_A_plhMp4FJ4_0),.din(w_dff_A_iTnffcDf9_0),.clk(gclk));
	jdff dff_A_plhMp4FJ4_0(.dout(G494),.din(w_dff_A_plhMp4FJ4_0),.clk(gclk));
	jdff dff_A_k7VluDx66_1(.dout(w_dff_A_4JCyLnPT8_0),.din(w_dff_A_k7VluDx66_1),.clk(gclk));
	jdff dff_A_4JCyLnPT8_0(.dout(w_dff_A_CqQVVofU5_0),.din(w_dff_A_4JCyLnPT8_0),.clk(gclk));
	jdff dff_A_CqQVVofU5_0(.dout(w_dff_A_0tGO98om5_0),.din(w_dff_A_CqQVVofU5_0),.clk(gclk));
	jdff dff_A_0tGO98om5_0(.dout(w_dff_A_cus2wNyR3_0),.din(w_dff_A_0tGO98om5_0),.clk(gclk));
	jdff dff_A_cus2wNyR3_0(.dout(w_dff_A_ykwg2N3S4_0),.din(w_dff_A_cus2wNyR3_0),.clk(gclk));
	jdff dff_A_ykwg2N3S4_0(.dout(w_dff_A_rHEvjDg05_0),.din(w_dff_A_ykwg2N3S4_0),.clk(gclk));
	jdff dff_A_rHEvjDg05_0(.dout(w_dff_A_Nr2H2tn92_0),.din(w_dff_A_rHEvjDg05_0),.clk(gclk));
	jdff dff_A_Nr2H2tn92_0(.dout(w_dff_A_OWbhJzUE5_0),.din(w_dff_A_Nr2H2tn92_0),.clk(gclk));
	jdff dff_A_OWbhJzUE5_0(.dout(w_dff_A_SyABLrul8_0),.din(w_dff_A_OWbhJzUE5_0),.clk(gclk));
	jdff dff_A_SyABLrul8_0(.dout(w_dff_A_oAEcGWz79_0),.din(w_dff_A_SyABLrul8_0),.clk(gclk));
	jdff dff_A_oAEcGWz79_0(.dout(w_dff_A_1JtRs0mg6_0),.din(w_dff_A_oAEcGWz79_0),.clk(gclk));
	jdff dff_A_1JtRs0mg6_0(.dout(w_dff_A_QvhOosfP7_0),.din(w_dff_A_1JtRs0mg6_0),.clk(gclk));
	jdff dff_A_QvhOosfP7_0(.dout(w_dff_A_cldCjiAI9_0),.din(w_dff_A_QvhOosfP7_0),.clk(gclk));
	jdff dff_A_cldCjiAI9_0(.dout(w_dff_A_2dCumnk10_0),.din(w_dff_A_cldCjiAI9_0),.clk(gclk));
	jdff dff_A_2dCumnk10_0(.dout(w_dff_A_drQEzZcd0_0),.din(w_dff_A_2dCumnk10_0),.clk(gclk));
	jdff dff_A_drQEzZcd0_0(.dout(w_dff_A_6m0xKfwG8_0),.din(w_dff_A_drQEzZcd0_0),.clk(gclk));
	jdff dff_A_6m0xKfwG8_0(.dout(w_dff_A_EMeWYtEd7_0),.din(w_dff_A_6m0xKfwG8_0),.clk(gclk));
	jdff dff_A_EMeWYtEd7_0(.dout(w_dff_A_mq1eryS33_0),.din(w_dff_A_EMeWYtEd7_0),.clk(gclk));
	jdff dff_A_mq1eryS33_0(.dout(w_dff_A_vw7Fow2q3_0),.din(w_dff_A_mq1eryS33_0),.clk(gclk));
	jdff dff_A_vw7Fow2q3_0(.dout(w_dff_A_7X219nVw4_0),.din(w_dff_A_vw7Fow2q3_0),.clk(gclk));
	jdff dff_A_7X219nVw4_0(.dout(w_dff_A_zTqGXTec1_0),.din(w_dff_A_7X219nVw4_0),.clk(gclk));
	jdff dff_A_zTqGXTec1_0(.dout(w_dff_A_SVAf83Wu1_0),.din(w_dff_A_zTqGXTec1_0),.clk(gclk));
	jdff dff_A_SVAf83Wu1_0(.dout(w_dff_A_GYtMXHAg0_0),.din(w_dff_A_SVAf83Wu1_0),.clk(gclk));
	jdff dff_A_GYtMXHAg0_0(.dout(w_dff_A_Lg75cSrF3_0),.din(w_dff_A_GYtMXHAg0_0),.clk(gclk));
	jdff dff_A_Lg75cSrF3_0(.dout(w_dff_A_7Aqi7KFB9_0),.din(w_dff_A_Lg75cSrF3_0),.clk(gclk));
	jdff dff_A_7Aqi7KFB9_0(.dout(G492),.din(w_dff_A_7Aqi7KFB9_0),.clk(gclk));
	jdff dff_A_f0loBwmj7_1(.dout(w_dff_A_UA06XAEd3_0),.din(w_dff_A_f0loBwmj7_1),.clk(gclk));
	jdff dff_A_UA06XAEd3_0(.dout(w_dff_A_KQkcnd6s5_0),.din(w_dff_A_UA06XAEd3_0),.clk(gclk));
	jdff dff_A_KQkcnd6s5_0(.dout(w_dff_A_Xebfgn7k8_0),.din(w_dff_A_KQkcnd6s5_0),.clk(gclk));
	jdff dff_A_Xebfgn7k8_0(.dout(w_dff_A_Kb6DbJdl0_0),.din(w_dff_A_Xebfgn7k8_0),.clk(gclk));
	jdff dff_A_Kb6DbJdl0_0(.dout(w_dff_A_oiQwF4St6_0),.din(w_dff_A_Kb6DbJdl0_0),.clk(gclk));
	jdff dff_A_oiQwF4St6_0(.dout(w_dff_A_7LVfNoyI8_0),.din(w_dff_A_oiQwF4St6_0),.clk(gclk));
	jdff dff_A_7LVfNoyI8_0(.dout(w_dff_A_fbw2mTka4_0),.din(w_dff_A_7LVfNoyI8_0),.clk(gclk));
	jdff dff_A_fbw2mTka4_0(.dout(w_dff_A_sguDky4c4_0),.din(w_dff_A_fbw2mTka4_0),.clk(gclk));
	jdff dff_A_sguDky4c4_0(.dout(w_dff_A_6G8WXdwX6_0),.din(w_dff_A_sguDky4c4_0),.clk(gclk));
	jdff dff_A_6G8WXdwX6_0(.dout(w_dff_A_uVPYL2Fk3_0),.din(w_dff_A_6G8WXdwX6_0),.clk(gclk));
	jdff dff_A_uVPYL2Fk3_0(.dout(w_dff_A_4VR2xzza4_0),.din(w_dff_A_uVPYL2Fk3_0),.clk(gclk));
	jdff dff_A_4VR2xzza4_0(.dout(w_dff_A_3c7hkXfT7_0),.din(w_dff_A_4VR2xzza4_0),.clk(gclk));
	jdff dff_A_3c7hkXfT7_0(.dout(w_dff_A_PLL3p1Ae0_0),.din(w_dff_A_3c7hkXfT7_0),.clk(gclk));
	jdff dff_A_PLL3p1Ae0_0(.dout(w_dff_A_UDPIlZY19_0),.din(w_dff_A_PLL3p1Ae0_0),.clk(gclk));
	jdff dff_A_UDPIlZY19_0(.dout(w_dff_A_gPGJ0XNR6_0),.din(w_dff_A_UDPIlZY19_0),.clk(gclk));
	jdff dff_A_gPGJ0XNR6_0(.dout(w_dff_A_VApq8idV0_0),.din(w_dff_A_gPGJ0XNR6_0),.clk(gclk));
	jdff dff_A_VApq8idV0_0(.dout(w_dff_A_PCnDiEUn8_0),.din(w_dff_A_VApq8idV0_0),.clk(gclk));
	jdff dff_A_PCnDiEUn8_0(.dout(w_dff_A_QcPzhlbh9_0),.din(w_dff_A_PCnDiEUn8_0),.clk(gclk));
	jdff dff_A_QcPzhlbh9_0(.dout(w_dff_A_PErFiEsZ7_0),.din(w_dff_A_QcPzhlbh9_0),.clk(gclk));
	jdff dff_A_PErFiEsZ7_0(.dout(w_dff_A_LPQLaZXx8_0),.din(w_dff_A_PErFiEsZ7_0),.clk(gclk));
	jdff dff_A_LPQLaZXx8_0(.dout(w_dff_A_nU3rmj2L1_0),.din(w_dff_A_LPQLaZXx8_0),.clk(gclk));
	jdff dff_A_nU3rmj2L1_0(.dout(w_dff_A_K9Z7zOhI0_0),.din(w_dff_A_nU3rmj2L1_0),.clk(gclk));
	jdff dff_A_K9Z7zOhI0_0(.dout(w_dff_A_5J3jbhlA4_0),.din(w_dff_A_K9Z7zOhI0_0),.clk(gclk));
	jdff dff_A_5J3jbhlA4_0(.dout(w_dff_A_qfbcGDFo5_0),.din(w_dff_A_5J3jbhlA4_0),.clk(gclk));
	jdff dff_A_qfbcGDFo5_0(.dout(w_dff_A_W040WQg59_0),.din(w_dff_A_qfbcGDFo5_0),.clk(gclk));
	jdff dff_A_W040WQg59_0(.dout(G490),.din(w_dff_A_W040WQg59_0),.clk(gclk));
	jdff dff_A_KZTb2yWC7_1(.dout(w_dff_A_9m7fLkwH1_0),.din(w_dff_A_KZTb2yWC7_1),.clk(gclk));
	jdff dff_A_9m7fLkwH1_0(.dout(w_dff_A_9o66xI0j9_0),.din(w_dff_A_9m7fLkwH1_0),.clk(gclk));
	jdff dff_A_9o66xI0j9_0(.dout(w_dff_A_74RbtHo87_0),.din(w_dff_A_9o66xI0j9_0),.clk(gclk));
	jdff dff_A_74RbtHo87_0(.dout(w_dff_A_SJrsLISZ6_0),.din(w_dff_A_74RbtHo87_0),.clk(gclk));
	jdff dff_A_SJrsLISZ6_0(.dout(w_dff_A_YDCImGTg2_0),.din(w_dff_A_SJrsLISZ6_0),.clk(gclk));
	jdff dff_A_YDCImGTg2_0(.dout(w_dff_A_pKIbaLtX3_0),.din(w_dff_A_YDCImGTg2_0),.clk(gclk));
	jdff dff_A_pKIbaLtX3_0(.dout(w_dff_A_8u03lCP34_0),.din(w_dff_A_pKIbaLtX3_0),.clk(gclk));
	jdff dff_A_8u03lCP34_0(.dout(w_dff_A_XAn5zpBf1_0),.din(w_dff_A_8u03lCP34_0),.clk(gclk));
	jdff dff_A_XAn5zpBf1_0(.dout(w_dff_A_ji7vzwIU7_0),.din(w_dff_A_XAn5zpBf1_0),.clk(gclk));
	jdff dff_A_ji7vzwIU7_0(.dout(w_dff_A_0CFrNTyK3_0),.din(w_dff_A_ji7vzwIU7_0),.clk(gclk));
	jdff dff_A_0CFrNTyK3_0(.dout(w_dff_A_SpUmqvJX4_0),.din(w_dff_A_0CFrNTyK3_0),.clk(gclk));
	jdff dff_A_SpUmqvJX4_0(.dout(w_dff_A_JFCxMApy4_0),.din(w_dff_A_SpUmqvJX4_0),.clk(gclk));
	jdff dff_A_JFCxMApy4_0(.dout(w_dff_A_2o52tIzB6_0),.din(w_dff_A_JFCxMApy4_0),.clk(gclk));
	jdff dff_A_2o52tIzB6_0(.dout(w_dff_A_X0IpWm9L2_0),.din(w_dff_A_2o52tIzB6_0),.clk(gclk));
	jdff dff_A_X0IpWm9L2_0(.dout(w_dff_A_67dkHOgN2_0),.din(w_dff_A_X0IpWm9L2_0),.clk(gclk));
	jdff dff_A_67dkHOgN2_0(.dout(w_dff_A_gC4IHWYU7_0),.din(w_dff_A_67dkHOgN2_0),.clk(gclk));
	jdff dff_A_gC4IHWYU7_0(.dout(w_dff_A_NuZIAZZe1_0),.din(w_dff_A_gC4IHWYU7_0),.clk(gclk));
	jdff dff_A_NuZIAZZe1_0(.dout(w_dff_A_YurapNLy8_0),.din(w_dff_A_NuZIAZZe1_0),.clk(gclk));
	jdff dff_A_YurapNLy8_0(.dout(w_dff_A_BLCgKjbE5_0),.din(w_dff_A_YurapNLy8_0),.clk(gclk));
	jdff dff_A_BLCgKjbE5_0(.dout(w_dff_A_nHtR25q09_0),.din(w_dff_A_BLCgKjbE5_0),.clk(gclk));
	jdff dff_A_nHtR25q09_0(.dout(w_dff_A_5m64xqTj3_0),.din(w_dff_A_nHtR25q09_0),.clk(gclk));
	jdff dff_A_5m64xqTj3_0(.dout(w_dff_A_C39eLG786_0),.din(w_dff_A_5m64xqTj3_0),.clk(gclk));
	jdff dff_A_C39eLG786_0(.dout(w_dff_A_Z5fCVx9H0_0),.din(w_dff_A_C39eLG786_0),.clk(gclk));
	jdff dff_A_Z5fCVx9H0_0(.dout(w_dff_A_Ypbcdhpv7_0),.din(w_dff_A_Z5fCVx9H0_0),.clk(gclk));
	jdff dff_A_Ypbcdhpv7_0(.dout(w_dff_A_Qm1nj8Uz2_0),.din(w_dff_A_Ypbcdhpv7_0),.clk(gclk));
	jdff dff_A_Qm1nj8Uz2_0(.dout(G488),.din(w_dff_A_Qm1nj8Uz2_0),.clk(gclk));
	jdff dff_A_QLfkh51b8_1(.dout(w_dff_A_DUa9HZnC3_0),.din(w_dff_A_QLfkh51b8_1),.clk(gclk));
	jdff dff_A_DUa9HZnC3_0(.dout(w_dff_A_UlCDh2JK1_0),.din(w_dff_A_DUa9HZnC3_0),.clk(gclk));
	jdff dff_A_UlCDh2JK1_0(.dout(w_dff_A_N2V6AKne6_0),.din(w_dff_A_UlCDh2JK1_0),.clk(gclk));
	jdff dff_A_N2V6AKne6_0(.dout(w_dff_A_cG8znGBF0_0),.din(w_dff_A_N2V6AKne6_0),.clk(gclk));
	jdff dff_A_cG8znGBF0_0(.dout(w_dff_A_jU9dvUXv4_0),.din(w_dff_A_cG8znGBF0_0),.clk(gclk));
	jdff dff_A_jU9dvUXv4_0(.dout(w_dff_A_6cpxOmBw2_0),.din(w_dff_A_jU9dvUXv4_0),.clk(gclk));
	jdff dff_A_6cpxOmBw2_0(.dout(w_dff_A_mc0wcpd06_0),.din(w_dff_A_6cpxOmBw2_0),.clk(gclk));
	jdff dff_A_mc0wcpd06_0(.dout(w_dff_A_LHj9tWjm9_0),.din(w_dff_A_mc0wcpd06_0),.clk(gclk));
	jdff dff_A_LHj9tWjm9_0(.dout(w_dff_A_1hts7Ibg8_0),.din(w_dff_A_LHj9tWjm9_0),.clk(gclk));
	jdff dff_A_1hts7Ibg8_0(.dout(w_dff_A_oB5odyPv2_0),.din(w_dff_A_1hts7Ibg8_0),.clk(gclk));
	jdff dff_A_oB5odyPv2_0(.dout(w_dff_A_MKcANnJ04_0),.din(w_dff_A_oB5odyPv2_0),.clk(gclk));
	jdff dff_A_MKcANnJ04_0(.dout(w_dff_A_9CFgohJx4_0),.din(w_dff_A_MKcANnJ04_0),.clk(gclk));
	jdff dff_A_9CFgohJx4_0(.dout(w_dff_A_QwEVE3bG8_0),.din(w_dff_A_9CFgohJx4_0),.clk(gclk));
	jdff dff_A_QwEVE3bG8_0(.dout(w_dff_A_vd3cvdKb9_0),.din(w_dff_A_QwEVE3bG8_0),.clk(gclk));
	jdff dff_A_vd3cvdKb9_0(.dout(w_dff_A_f0Zkd5IP9_0),.din(w_dff_A_vd3cvdKb9_0),.clk(gclk));
	jdff dff_A_f0Zkd5IP9_0(.dout(w_dff_A_W3zNEd0U5_0),.din(w_dff_A_f0Zkd5IP9_0),.clk(gclk));
	jdff dff_A_W3zNEd0U5_0(.dout(w_dff_A_z1aJ5j6L9_0),.din(w_dff_A_W3zNEd0U5_0),.clk(gclk));
	jdff dff_A_z1aJ5j6L9_0(.dout(w_dff_A_FjTypjNG6_0),.din(w_dff_A_z1aJ5j6L9_0),.clk(gclk));
	jdff dff_A_FjTypjNG6_0(.dout(w_dff_A_G7vqqoYa4_0),.din(w_dff_A_FjTypjNG6_0),.clk(gclk));
	jdff dff_A_G7vqqoYa4_0(.dout(w_dff_A_xw6jvl1U5_0),.din(w_dff_A_G7vqqoYa4_0),.clk(gclk));
	jdff dff_A_xw6jvl1U5_0(.dout(w_dff_A_SDEeN8se9_0),.din(w_dff_A_xw6jvl1U5_0),.clk(gclk));
	jdff dff_A_SDEeN8se9_0(.dout(w_dff_A_bIifVykH6_0),.din(w_dff_A_SDEeN8se9_0),.clk(gclk));
	jdff dff_A_bIifVykH6_0(.dout(w_dff_A_CtIWqBnI8_0),.din(w_dff_A_bIifVykH6_0),.clk(gclk));
	jdff dff_A_CtIWqBnI8_0(.dout(w_dff_A_5PdX3Cv19_0),.din(w_dff_A_CtIWqBnI8_0),.clk(gclk));
	jdff dff_A_5PdX3Cv19_0(.dout(w_dff_A_RIUIkOOA8_0),.din(w_dff_A_5PdX3Cv19_0),.clk(gclk));
	jdff dff_A_RIUIkOOA8_0(.dout(G486),.din(w_dff_A_RIUIkOOA8_0),.clk(gclk));
	jdff dff_A_OfURwhBQ4_1(.dout(w_dff_A_ytSQMmZV7_0),.din(w_dff_A_OfURwhBQ4_1),.clk(gclk));
	jdff dff_A_ytSQMmZV7_0(.dout(w_dff_A_yINPCqiF1_0),.din(w_dff_A_ytSQMmZV7_0),.clk(gclk));
	jdff dff_A_yINPCqiF1_0(.dout(w_dff_A_aX0zZrfI5_0),.din(w_dff_A_yINPCqiF1_0),.clk(gclk));
	jdff dff_A_aX0zZrfI5_0(.dout(w_dff_A_Z4owilih7_0),.din(w_dff_A_aX0zZrfI5_0),.clk(gclk));
	jdff dff_A_Z4owilih7_0(.dout(w_dff_A_tA2mEIM04_0),.din(w_dff_A_Z4owilih7_0),.clk(gclk));
	jdff dff_A_tA2mEIM04_0(.dout(w_dff_A_RNvZio891_0),.din(w_dff_A_tA2mEIM04_0),.clk(gclk));
	jdff dff_A_RNvZio891_0(.dout(w_dff_A_7PgBZI536_0),.din(w_dff_A_RNvZio891_0),.clk(gclk));
	jdff dff_A_7PgBZI536_0(.dout(w_dff_A_ZMV5J3RQ6_0),.din(w_dff_A_7PgBZI536_0),.clk(gclk));
	jdff dff_A_ZMV5J3RQ6_0(.dout(w_dff_A_zDAudBa62_0),.din(w_dff_A_ZMV5J3RQ6_0),.clk(gclk));
	jdff dff_A_zDAudBa62_0(.dout(w_dff_A_drX3DFpO8_0),.din(w_dff_A_zDAudBa62_0),.clk(gclk));
	jdff dff_A_drX3DFpO8_0(.dout(w_dff_A_iwCJhtCM6_0),.din(w_dff_A_drX3DFpO8_0),.clk(gclk));
	jdff dff_A_iwCJhtCM6_0(.dout(w_dff_A_VnZKnpWY9_0),.din(w_dff_A_iwCJhtCM6_0),.clk(gclk));
	jdff dff_A_VnZKnpWY9_0(.dout(w_dff_A_uRyf39Wa0_0),.din(w_dff_A_VnZKnpWY9_0),.clk(gclk));
	jdff dff_A_uRyf39Wa0_0(.dout(w_dff_A_XCCaCKBf8_0),.din(w_dff_A_uRyf39Wa0_0),.clk(gclk));
	jdff dff_A_XCCaCKBf8_0(.dout(w_dff_A_0RZ9zW1X4_0),.din(w_dff_A_XCCaCKBf8_0),.clk(gclk));
	jdff dff_A_0RZ9zW1X4_0(.dout(w_dff_A_WfZcjshR7_0),.din(w_dff_A_0RZ9zW1X4_0),.clk(gclk));
	jdff dff_A_WfZcjshR7_0(.dout(w_dff_A_B88VNbXs3_0),.din(w_dff_A_WfZcjshR7_0),.clk(gclk));
	jdff dff_A_B88VNbXs3_0(.dout(w_dff_A_YkKK2TBb4_0),.din(w_dff_A_B88VNbXs3_0),.clk(gclk));
	jdff dff_A_YkKK2TBb4_0(.dout(w_dff_A_3JpGJlkj6_0),.din(w_dff_A_YkKK2TBb4_0),.clk(gclk));
	jdff dff_A_3JpGJlkj6_0(.dout(w_dff_A_aRnGBIFF9_0),.din(w_dff_A_3JpGJlkj6_0),.clk(gclk));
	jdff dff_A_aRnGBIFF9_0(.dout(w_dff_A_9LIutuJ13_0),.din(w_dff_A_aRnGBIFF9_0),.clk(gclk));
	jdff dff_A_9LIutuJ13_0(.dout(w_dff_A_AagqdROk1_0),.din(w_dff_A_9LIutuJ13_0),.clk(gclk));
	jdff dff_A_AagqdROk1_0(.dout(w_dff_A_QmDodXM35_0),.din(w_dff_A_AagqdROk1_0),.clk(gclk));
	jdff dff_A_QmDodXM35_0(.dout(w_dff_A_9HjBWwfe6_0),.din(w_dff_A_QmDodXM35_0),.clk(gclk));
	jdff dff_A_9HjBWwfe6_0(.dout(w_dff_A_980EDFiP5_0),.din(w_dff_A_9HjBWwfe6_0),.clk(gclk));
	jdff dff_A_980EDFiP5_0(.dout(G484),.din(w_dff_A_980EDFiP5_0),.clk(gclk));
	jdff dff_A_fIekaECE3_1(.dout(w_dff_A_bk775PTy5_0),.din(w_dff_A_fIekaECE3_1),.clk(gclk));
	jdff dff_A_bk775PTy5_0(.dout(w_dff_A_IIfDcN731_0),.din(w_dff_A_bk775PTy5_0),.clk(gclk));
	jdff dff_A_IIfDcN731_0(.dout(w_dff_A_5PMu0ONu2_0),.din(w_dff_A_IIfDcN731_0),.clk(gclk));
	jdff dff_A_5PMu0ONu2_0(.dout(w_dff_A_eLol9rpd9_0),.din(w_dff_A_5PMu0ONu2_0),.clk(gclk));
	jdff dff_A_eLol9rpd9_0(.dout(w_dff_A_PLHaiAic9_0),.din(w_dff_A_eLol9rpd9_0),.clk(gclk));
	jdff dff_A_PLHaiAic9_0(.dout(w_dff_A_mZTV7jyz6_0),.din(w_dff_A_PLHaiAic9_0),.clk(gclk));
	jdff dff_A_mZTV7jyz6_0(.dout(w_dff_A_lcJl65Ah2_0),.din(w_dff_A_mZTV7jyz6_0),.clk(gclk));
	jdff dff_A_lcJl65Ah2_0(.dout(w_dff_A_6QXCIqm39_0),.din(w_dff_A_lcJl65Ah2_0),.clk(gclk));
	jdff dff_A_6QXCIqm39_0(.dout(w_dff_A_dSNySXUc9_0),.din(w_dff_A_6QXCIqm39_0),.clk(gclk));
	jdff dff_A_dSNySXUc9_0(.dout(w_dff_A_7l5v8nxi4_0),.din(w_dff_A_dSNySXUc9_0),.clk(gclk));
	jdff dff_A_7l5v8nxi4_0(.dout(w_dff_A_rNrrtCYT4_0),.din(w_dff_A_7l5v8nxi4_0),.clk(gclk));
	jdff dff_A_rNrrtCYT4_0(.dout(w_dff_A_CHI7qLaG5_0),.din(w_dff_A_rNrrtCYT4_0),.clk(gclk));
	jdff dff_A_CHI7qLaG5_0(.dout(w_dff_A_sELod8Nb5_0),.din(w_dff_A_CHI7qLaG5_0),.clk(gclk));
	jdff dff_A_sELod8Nb5_0(.dout(w_dff_A_xf27V03z0_0),.din(w_dff_A_sELod8Nb5_0),.clk(gclk));
	jdff dff_A_xf27V03z0_0(.dout(w_dff_A_7tmE429A8_0),.din(w_dff_A_xf27V03z0_0),.clk(gclk));
	jdff dff_A_7tmE429A8_0(.dout(w_dff_A_MESAuxb88_0),.din(w_dff_A_7tmE429A8_0),.clk(gclk));
	jdff dff_A_MESAuxb88_0(.dout(w_dff_A_vwHscXbt7_0),.din(w_dff_A_MESAuxb88_0),.clk(gclk));
	jdff dff_A_vwHscXbt7_0(.dout(w_dff_A_PLGKFfh65_0),.din(w_dff_A_vwHscXbt7_0),.clk(gclk));
	jdff dff_A_PLGKFfh65_0(.dout(w_dff_A_d75bt1mm2_0),.din(w_dff_A_PLGKFfh65_0),.clk(gclk));
	jdff dff_A_d75bt1mm2_0(.dout(w_dff_A_etmB4GOC4_0),.din(w_dff_A_d75bt1mm2_0),.clk(gclk));
	jdff dff_A_etmB4GOC4_0(.dout(w_dff_A_sBArkJi94_0),.din(w_dff_A_etmB4GOC4_0),.clk(gclk));
	jdff dff_A_sBArkJi94_0(.dout(w_dff_A_Z8MyH8wl9_0),.din(w_dff_A_sBArkJi94_0),.clk(gclk));
	jdff dff_A_Z8MyH8wl9_0(.dout(w_dff_A_Z2kC9TQE6_0),.din(w_dff_A_Z8MyH8wl9_0),.clk(gclk));
	jdff dff_A_Z2kC9TQE6_0(.dout(w_dff_A_nLGhbYri1_0),.din(w_dff_A_Z2kC9TQE6_0),.clk(gclk));
	jdff dff_A_nLGhbYri1_0(.dout(w_dff_A_CCE3pTEC0_0),.din(w_dff_A_nLGhbYri1_0),.clk(gclk));
	jdff dff_A_CCE3pTEC0_0(.dout(G482),.din(w_dff_A_CCE3pTEC0_0),.clk(gclk));
	jdff dff_A_gOv57F6o7_1(.dout(w_dff_A_4ycNk5ue3_0),.din(w_dff_A_gOv57F6o7_1),.clk(gclk));
	jdff dff_A_4ycNk5ue3_0(.dout(w_dff_A_kQb6alwb4_0),.din(w_dff_A_4ycNk5ue3_0),.clk(gclk));
	jdff dff_A_kQb6alwb4_0(.dout(w_dff_A_750YHGfC0_0),.din(w_dff_A_kQb6alwb4_0),.clk(gclk));
	jdff dff_A_750YHGfC0_0(.dout(w_dff_A_1jsP5YW74_0),.din(w_dff_A_750YHGfC0_0),.clk(gclk));
	jdff dff_A_1jsP5YW74_0(.dout(w_dff_A_rQRGYg105_0),.din(w_dff_A_1jsP5YW74_0),.clk(gclk));
	jdff dff_A_rQRGYg105_0(.dout(w_dff_A_pGGC2MO08_0),.din(w_dff_A_rQRGYg105_0),.clk(gclk));
	jdff dff_A_pGGC2MO08_0(.dout(w_dff_A_hz0j8EbO0_0),.din(w_dff_A_pGGC2MO08_0),.clk(gclk));
	jdff dff_A_hz0j8EbO0_0(.dout(w_dff_A_wvPlMp6f5_0),.din(w_dff_A_hz0j8EbO0_0),.clk(gclk));
	jdff dff_A_wvPlMp6f5_0(.dout(w_dff_A_te0lC6vD2_0),.din(w_dff_A_wvPlMp6f5_0),.clk(gclk));
	jdff dff_A_te0lC6vD2_0(.dout(w_dff_A_lTnOwFar8_0),.din(w_dff_A_te0lC6vD2_0),.clk(gclk));
	jdff dff_A_lTnOwFar8_0(.dout(w_dff_A_axSqLTYo9_0),.din(w_dff_A_lTnOwFar8_0),.clk(gclk));
	jdff dff_A_axSqLTYo9_0(.dout(w_dff_A_vVKtUhnG0_0),.din(w_dff_A_axSqLTYo9_0),.clk(gclk));
	jdff dff_A_vVKtUhnG0_0(.dout(w_dff_A_gKwZEhym9_0),.din(w_dff_A_vVKtUhnG0_0),.clk(gclk));
	jdff dff_A_gKwZEhym9_0(.dout(w_dff_A_SQYHVqPZ2_0),.din(w_dff_A_gKwZEhym9_0),.clk(gclk));
	jdff dff_A_SQYHVqPZ2_0(.dout(w_dff_A_GszOT3Ft5_0),.din(w_dff_A_SQYHVqPZ2_0),.clk(gclk));
	jdff dff_A_GszOT3Ft5_0(.dout(w_dff_A_1KIl7Y784_0),.din(w_dff_A_GszOT3Ft5_0),.clk(gclk));
	jdff dff_A_1KIl7Y784_0(.dout(w_dff_A_HGmNnvMP1_0),.din(w_dff_A_1KIl7Y784_0),.clk(gclk));
	jdff dff_A_HGmNnvMP1_0(.dout(w_dff_A_fjvhIx1R6_0),.din(w_dff_A_HGmNnvMP1_0),.clk(gclk));
	jdff dff_A_fjvhIx1R6_0(.dout(w_dff_A_VKCNYq9P8_0),.din(w_dff_A_fjvhIx1R6_0),.clk(gclk));
	jdff dff_A_VKCNYq9P8_0(.dout(w_dff_A_lM8MGmMt3_0),.din(w_dff_A_VKCNYq9P8_0),.clk(gclk));
	jdff dff_A_lM8MGmMt3_0(.dout(w_dff_A_N8yYnooQ6_0),.din(w_dff_A_lM8MGmMt3_0),.clk(gclk));
	jdff dff_A_N8yYnooQ6_0(.dout(w_dff_A_NSmpGyrU1_0),.din(w_dff_A_N8yYnooQ6_0),.clk(gclk));
	jdff dff_A_NSmpGyrU1_0(.dout(w_dff_A_PWWzkdMT3_0),.din(w_dff_A_NSmpGyrU1_0),.clk(gclk));
	jdff dff_A_PWWzkdMT3_0(.dout(w_dff_A_AcKnVu8F1_0),.din(w_dff_A_PWWzkdMT3_0),.clk(gclk));
	jdff dff_A_AcKnVu8F1_0(.dout(w_dff_A_1IMPCMjz6_0),.din(w_dff_A_AcKnVu8F1_0),.clk(gclk));
	jdff dff_A_1IMPCMjz6_0(.dout(G480),.din(w_dff_A_1IMPCMjz6_0),.clk(gclk));
	jdff dff_A_11QQyRH85_1(.dout(w_dff_A_UjXJohJy7_0),.din(w_dff_A_11QQyRH85_1),.clk(gclk));
	jdff dff_A_UjXJohJy7_0(.dout(w_dff_A_ShEUuRJO0_0),.din(w_dff_A_UjXJohJy7_0),.clk(gclk));
	jdff dff_A_ShEUuRJO0_0(.dout(w_dff_A_tg3mlVew4_0),.din(w_dff_A_ShEUuRJO0_0),.clk(gclk));
	jdff dff_A_tg3mlVew4_0(.dout(w_dff_A_4J1i6TzQ3_0),.din(w_dff_A_tg3mlVew4_0),.clk(gclk));
	jdff dff_A_4J1i6TzQ3_0(.dout(w_dff_A_7ZwDlCyW6_0),.din(w_dff_A_4J1i6TzQ3_0),.clk(gclk));
	jdff dff_A_7ZwDlCyW6_0(.dout(w_dff_A_VXPcrupP7_0),.din(w_dff_A_7ZwDlCyW6_0),.clk(gclk));
	jdff dff_A_VXPcrupP7_0(.dout(w_dff_A_Itga5flg1_0),.din(w_dff_A_VXPcrupP7_0),.clk(gclk));
	jdff dff_A_Itga5flg1_0(.dout(w_dff_A_VwnCLoSN9_0),.din(w_dff_A_Itga5flg1_0),.clk(gclk));
	jdff dff_A_VwnCLoSN9_0(.dout(w_dff_A_91dpDgg91_0),.din(w_dff_A_VwnCLoSN9_0),.clk(gclk));
	jdff dff_A_91dpDgg91_0(.dout(w_dff_A_UpWY8KVq9_0),.din(w_dff_A_91dpDgg91_0),.clk(gclk));
	jdff dff_A_UpWY8KVq9_0(.dout(w_dff_A_bAoMvQUp4_0),.din(w_dff_A_UpWY8KVq9_0),.clk(gclk));
	jdff dff_A_bAoMvQUp4_0(.dout(w_dff_A_UgK6i5xj8_0),.din(w_dff_A_bAoMvQUp4_0),.clk(gclk));
	jdff dff_A_UgK6i5xj8_0(.dout(w_dff_A_3H0IbKDz8_0),.din(w_dff_A_UgK6i5xj8_0),.clk(gclk));
	jdff dff_A_3H0IbKDz8_0(.dout(w_dff_A_wbSVtmAL5_0),.din(w_dff_A_3H0IbKDz8_0),.clk(gclk));
	jdff dff_A_wbSVtmAL5_0(.dout(w_dff_A_83nN3jnE0_0),.din(w_dff_A_wbSVtmAL5_0),.clk(gclk));
	jdff dff_A_83nN3jnE0_0(.dout(w_dff_A_52jTadLY9_0),.din(w_dff_A_83nN3jnE0_0),.clk(gclk));
	jdff dff_A_52jTadLY9_0(.dout(w_dff_A_Bt01Oqwz6_0),.din(w_dff_A_52jTadLY9_0),.clk(gclk));
	jdff dff_A_Bt01Oqwz6_0(.dout(w_dff_A_BAh45ch20_0),.din(w_dff_A_Bt01Oqwz6_0),.clk(gclk));
	jdff dff_A_BAh45ch20_0(.dout(w_dff_A_lVSsa0Tp3_0),.din(w_dff_A_BAh45ch20_0),.clk(gclk));
	jdff dff_A_lVSsa0Tp3_0(.dout(w_dff_A_WlWbRkXP1_0),.din(w_dff_A_lVSsa0Tp3_0),.clk(gclk));
	jdff dff_A_WlWbRkXP1_0(.dout(w_dff_A_P2OROSa06_0),.din(w_dff_A_WlWbRkXP1_0),.clk(gclk));
	jdff dff_A_P2OROSa06_0(.dout(w_dff_A_SxaMNOeq4_0),.din(w_dff_A_P2OROSa06_0),.clk(gclk));
	jdff dff_A_SxaMNOeq4_0(.dout(w_dff_A_yA0kOM8s5_0),.din(w_dff_A_SxaMNOeq4_0),.clk(gclk));
	jdff dff_A_yA0kOM8s5_0(.dout(w_dff_A_2QpzgJ2M6_0),.din(w_dff_A_yA0kOM8s5_0),.clk(gclk));
	jdff dff_A_2QpzgJ2M6_0(.dout(w_dff_A_Cnhvxw4A4_0),.din(w_dff_A_2QpzgJ2M6_0),.clk(gclk));
	jdff dff_A_Cnhvxw4A4_0(.dout(G560),.din(w_dff_A_Cnhvxw4A4_0),.clk(gclk));
	jdff dff_A_9okMP1UV2_1(.dout(w_dff_A_W0z5pZCe5_0),.din(w_dff_A_9okMP1UV2_1),.clk(gclk));
	jdff dff_A_W0z5pZCe5_0(.dout(w_dff_A_tqrobSO45_0),.din(w_dff_A_W0z5pZCe5_0),.clk(gclk));
	jdff dff_A_tqrobSO45_0(.dout(w_dff_A_olNmtkdm8_0),.din(w_dff_A_tqrobSO45_0),.clk(gclk));
	jdff dff_A_olNmtkdm8_0(.dout(w_dff_A_vckhYKQb4_0),.din(w_dff_A_olNmtkdm8_0),.clk(gclk));
	jdff dff_A_vckhYKQb4_0(.dout(w_dff_A_kBPXqeMc7_0),.din(w_dff_A_vckhYKQb4_0),.clk(gclk));
	jdff dff_A_kBPXqeMc7_0(.dout(w_dff_A_g3WJ2c3N6_0),.din(w_dff_A_kBPXqeMc7_0),.clk(gclk));
	jdff dff_A_g3WJ2c3N6_0(.dout(w_dff_A_wM3Xz4T23_0),.din(w_dff_A_g3WJ2c3N6_0),.clk(gclk));
	jdff dff_A_wM3Xz4T23_0(.dout(w_dff_A_CCiZ0XNY6_0),.din(w_dff_A_wM3Xz4T23_0),.clk(gclk));
	jdff dff_A_CCiZ0XNY6_0(.dout(w_dff_A_xLCoukH15_0),.din(w_dff_A_CCiZ0XNY6_0),.clk(gclk));
	jdff dff_A_xLCoukH15_0(.dout(w_dff_A_XGY4ms5n3_0),.din(w_dff_A_xLCoukH15_0),.clk(gclk));
	jdff dff_A_XGY4ms5n3_0(.dout(w_dff_A_G41BNQGi2_0),.din(w_dff_A_XGY4ms5n3_0),.clk(gclk));
	jdff dff_A_G41BNQGi2_0(.dout(w_dff_A_FL7zkHKh0_0),.din(w_dff_A_G41BNQGi2_0),.clk(gclk));
	jdff dff_A_FL7zkHKh0_0(.dout(w_dff_A_3HXQdHjF9_0),.din(w_dff_A_FL7zkHKh0_0),.clk(gclk));
	jdff dff_A_3HXQdHjF9_0(.dout(w_dff_A_5gDjCqpK0_0),.din(w_dff_A_3HXQdHjF9_0),.clk(gclk));
	jdff dff_A_5gDjCqpK0_0(.dout(w_dff_A_nOXzo6UW1_0),.din(w_dff_A_5gDjCqpK0_0),.clk(gclk));
	jdff dff_A_nOXzo6UW1_0(.dout(w_dff_A_9zHsPENT5_0),.din(w_dff_A_nOXzo6UW1_0),.clk(gclk));
	jdff dff_A_9zHsPENT5_0(.dout(w_dff_A_SSqTzJ4a8_0),.din(w_dff_A_9zHsPENT5_0),.clk(gclk));
	jdff dff_A_SSqTzJ4a8_0(.dout(w_dff_A_WC0oSFax0_0),.din(w_dff_A_SSqTzJ4a8_0),.clk(gclk));
	jdff dff_A_WC0oSFax0_0(.dout(w_dff_A_Nw7VJFwA3_0),.din(w_dff_A_WC0oSFax0_0),.clk(gclk));
	jdff dff_A_Nw7VJFwA3_0(.dout(w_dff_A_a2kMC4mj5_0),.din(w_dff_A_Nw7VJFwA3_0),.clk(gclk));
	jdff dff_A_a2kMC4mj5_0(.dout(w_dff_A_FMGgHupn6_0),.din(w_dff_A_a2kMC4mj5_0),.clk(gclk));
	jdff dff_A_FMGgHupn6_0(.dout(w_dff_A_F6impo4g7_0),.din(w_dff_A_FMGgHupn6_0),.clk(gclk));
	jdff dff_A_F6impo4g7_0(.dout(w_dff_A_T8b8AyAx1_0),.din(w_dff_A_F6impo4g7_0),.clk(gclk));
	jdff dff_A_T8b8AyAx1_0(.dout(w_dff_A_B7P0jwiJ3_0),.din(w_dff_A_T8b8AyAx1_0),.clk(gclk));
	jdff dff_A_B7P0jwiJ3_0(.dout(w_dff_A_QByHr7ms8_0),.din(w_dff_A_B7P0jwiJ3_0),.clk(gclk));
	jdff dff_A_QByHr7ms8_0(.dout(G542),.din(w_dff_A_QByHr7ms8_0),.clk(gclk));
	jdff dff_A_XMLPmksm8_1(.dout(w_dff_A_nXCBi7Zg4_0),.din(w_dff_A_XMLPmksm8_1),.clk(gclk));
	jdff dff_A_nXCBi7Zg4_0(.dout(w_dff_A_vata1kJy9_0),.din(w_dff_A_nXCBi7Zg4_0),.clk(gclk));
	jdff dff_A_vata1kJy9_0(.dout(w_dff_A_X5xU5kKc2_0),.din(w_dff_A_vata1kJy9_0),.clk(gclk));
	jdff dff_A_X5xU5kKc2_0(.dout(w_dff_A_OcHyEATI4_0),.din(w_dff_A_X5xU5kKc2_0),.clk(gclk));
	jdff dff_A_OcHyEATI4_0(.dout(w_dff_A_xtrwPTaF7_0),.din(w_dff_A_OcHyEATI4_0),.clk(gclk));
	jdff dff_A_xtrwPTaF7_0(.dout(w_dff_A_TuikUtQJ5_0),.din(w_dff_A_xtrwPTaF7_0),.clk(gclk));
	jdff dff_A_TuikUtQJ5_0(.dout(w_dff_A_ScJYNUfR6_0),.din(w_dff_A_TuikUtQJ5_0),.clk(gclk));
	jdff dff_A_ScJYNUfR6_0(.dout(w_dff_A_EFkx2fPr0_0),.din(w_dff_A_ScJYNUfR6_0),.clk(gclk));
	jdff dff_A_EFkx2fPr0_0(.dout(w_dff_A_05fRovvS0_0),.din(w_dff_A_EFkx2fPr0_0),.clk(gclk));
	jdff dff_A_05fRovvS0_0(.dout(w_dff_A_gOoMGAOP1_0),.din(w_dff_A_05fRovvS0_0),.clk(gclk));
	jdff dff_A_gOoMGAOP1_0(.dout(w_dff_A_6CdV0Dx76_0),.din(w_dff_A_gOoMGAOP1_0),.clk(gclk));
	jdff dff_A_6CdV0Dx76_0(.dout(w_dff_A_vhsbPAM43_0),.din(w_dff_A_6CdV0Dx76_0),.clk(gclk));
	jdff dff_A_vhsbPAM43_0(.dout(w_dff_A_U2PW0Nf06_0),.din(w_dff_A_vhsbPAM43_0),.clk(gclk));
	jdff dff_A_U2PW0Nf06_0(.dout(w_dff_A_x6PQxXnG6_0),.din(w_dff_A_U2PW0Nf06_0),.clk(gclk));
	jdff dff_A_x6PQxXnG6_0(.dout(w_dff_A_g1Ki7iYn5_0),.din(w_dff_A_x6PQxXnG6_0),.clk(gclk));
	jdff dff_A_g1Ki7iYn5_0(.dout(w_dff_A_LSN81seR6_0),.din(w_dff_A_g1Ki7iYn5_0),.clk(gclk));
	jdff dff_A_LSN81seR6_0(.dout(w_dff_A_umLDc4e32_0),.din(w_dff_A_LSN81seR6_0),.clk(gclk));
	jdff dff_A_umLDc4e32_0(.dout(w_dff_A_D3Z8w65C0_0),.din(w_dff_A_umLDc4e32_0),.clk(gclk));
	jdff dff_A_D3Z8w65C0_0(.dout(w_dff_A_kZ0VP6MF3_0),.din(w_dff_A_D3Z8w65C0_0),.clk(gclk));
	jdff dff_A_kZ0VP6MF3_0(.dout(w_dff_A_9MQfuMzn7_0),.din(w_dff_A_kZ0VP6MF3_0),.clk(gclk));
	jdff dff_A_9MQfuMzn7_0(.dout(w_dff_A_Q4hBb8IV3_0),.din(w_dff_A_9MQfuMzn7_0),.clk(gclk));
	jdff dff_A_Q4hBb8IV3_0(.dout(w_dff_A_zSXUF6JB8_0),.din(w_dff_A_Q4hBb8IV3_0),.clk(gclk));
	jdff dff_A_zSXUF6JB8_0(.dout(w_dff_A_FxPuHxzq9_0),.din(w_dff_A_zSXUF6JB8_0),.clk(gclk));
	jdff dff_A_FxPuHxzq9_0(.dout(w_dff_A_fIEu4iUG2_0),.din(w_dff_A_FxPuHxzq9_0),.clk(gclk));
	jdff dff_A_fIEu4iUG2_0(.dout(w_dff_A_aSYzNRAE5_0),.din(w_dff_A_fIEu4iUG2_0),.clk(gclk));
	jdff dff_A_aSYzNRAE5_0(.dout(G558),.din(w_dff_A_aSYzNRAE5_0),.clk(gclk));
	jdff dff_A_RwGKFHG76_1(.dout(w_dff_A_pSsJqAGi2_0),.din(w_dff_A_RwGKFHG76_1),.clk(gclk));
	jdff dff_A_pSsJqAGi2_0(.dout(w_dff_A_QTQ3LRou3_0),.din(w_dff_A_pSsJqAGi2_0),.clk(gclk));
	jdff dff_A_QTQ3LRou3_0(.dout(w_dff_A_zHpTy2Ma4_0),.din(w_dff_A_QTQ3LRou3_0),.clk(gclk));
	jdff dff_A_zHpTy2Ma4_0(.dout(w_dff_A_6U9Q47tX8_0),.din(w_dff_A_zHpTy2Ma4_0),.clk(gclk));
	jdff dff_A_6U9Q47tX8_0(.dout(w_dff_A_vQSlVRYl5_0),.din(w_dff_A_6U9Q47tX8_0),.clk(gclk));
	jdff dff_A_vQSlVRYl5_0(.dout(w_dff_A_lqbPE6rA9_0),.din(w_dff_A_vQSlVRYl5_0),.clk(gclk));
	jdff dff_A_lqbPE6rA9_0(.dout(w_dff_A_DhQ8CBJN5_0),.din(w_dff_A_lqbPE6rA9_0),.clk(gclk));
	jdff dff_A_DhQ8CBJN5_0(.dout(w_dff_A_0mmd6iAP6_0),.din(w_dff_A_DhQ8CBJN5_0),.clk(gclk));
	jdff dff_A_0mmd6iAP6_0(.dout(w_dff_A_B4B3iqNi7_0),.din(w_dff_A_0mmd6iAP6_0),.clk(gclk));
	jdff dff_A_B4B3iqNi7_0(.dout(w_dff_A_6V3SgN718_0),.din(w_dff_A_B4B3iqNi7_0),.clk(gclk));
	jdff dff_A_6V3SgN718_0(.dout(w_dff_A_xPzwMw5Y4_0),.din(w_dff_A_6V3SgN718_0),.clk(gclk));
	jdff dff_A_xPzwMw5Y4_0(.dout(w_dff_A_pFhm7M850_0),.din(w_dff_A_xPzwMw5Y4_0),.clk(gclk));
	jdff dff_A_pFhm7M850_0(.dout(w_dff_A_DHgizohK1_0),.din(w_dff_A_pFhm7M850_0),.clk(gclk));
	jdff dff_A_DHgizohK1_0(.dout(w_dff_A_QoKQdfTy8_0),.din(w_dff_A_DHgizohK1_0),.clk(gclk));
	jdff dff_A_QoKQdfTy8_0(.dout(w_dff_A_xdsvHBIa9_0),.din(w_dff_A_QoKQdfTy8_0),.clk(gclk));
	jdff dff_A_xdsvHBIa9_0(.dout(w_dff_A_FqKVM69n1_0),.din(w_dff_A_xdsvHBIa9_0),.clk(gclk));
	jdff dff_A_FqKVM69n1_0(.dout(w_dff_A_z73PWgP01_0),.din(w_dff_A_FqKVM69n1_0),.clk(gclk));
	jdff dff_A_z73PWgP01_0(.dout(w_dff_A_KZNvMPRo8_0),.din(w_dff_A_z73PWgP01_0),.clk(gclk));
	jdff dff_A_KZNvMPRo8_0(.dout(w_dff_A_DDY7NAzT2_0),.din(w_dff_A_KZNvMPRo8_0),.clk(gclk));
	jdff dff_A_DDY7NAzT2_0(.dout(w_dff_A_WmMGUKcV8_0),.din(w_dff_A_DDY7NAzT2_0),.clk(gclk));
	jdff dff_A_WmMGUKcV8_0(.dout(w_dff_A_Eu8t7ZoD2_0),.din(w_dff_A_WmMGUKcV8_0),.clk(gclk));
	jdff dff_A_Eu8t7ZoD2_0(.dout(w_dff_A_Ui7AEILB9_0),.din(w_dff_A_Eu8t7ZoD2_0),.clk(gclk));
	jdff dff_A_Ui7AEILB9_0(.dout(w_dff_A_MXzLsN6d8_0),.din(w_dff_A_Ui7AEILB9_0),.clk(gclk));
	jdff dff_A_MXzLsN6d8_0(.dout(w_dff_A_uaTHpDKo8_0),.din(w_dff_A_MXzLsN6d8_0),.clk(gclk));
	jdff dff_A_uaTHpDKo8_0(.dout(w_dff_A_yI6apG2r3_0),.din(w_dff_A_uaTHpDKo8_0),.clk(gclk));
	jdff dff_A_yI6apG2r3_0(.dout(G556),.din(w_dff_A_yI6apG2r3_0),.clk(gclk));
	jdff dff_A_o7j95bj09_1(.dout(w_dff_A_RCk2tpz64_0),.din(w_dff_A_o7j95bj09_1),.clk(gclk));
	jdff dff_A_RCk2tpz64_0(.dout(w_dff_A_9iGhDWcK7_0),.din(w_dff_A_RCk2tpz64_0),.clk(gclk));
	jdff dff_A_9iGhDWcK7_0(.dout(w_dff_A_dsHEauon1_0),.din(w_dff_A_9iGhDWcK7_0),.clk(gclk));
	jdff dff_A_dsHEauon1_0(.dout(w_dff_A_8AZu8qJD2_0),.din(w_dff_A_dsHEauon1_0),.clk(gclk));
	jdff dff_A_8AZu8qJD2_0(.dout(w_dff_A_7uOv7Jir4_0),.din(w_dff_A_8AZu8qJD2_0),.clk(gclk));
	jdff dff_A_7uOv7Jir4_0(.dout(w_dff_A_0Cliso2d7_0),.din(w_dff_A_7uOv7Jir4_0),.clk(gclk));
	jdff dff_A_0Cliso2d7_0(.dout(w_dff_A_1qFCwSei7_0),.din(w_dff_A_0Cliso2d7_0),.clk(gclk));
	jdff dff_A_1qFCwSei7_0(.dout(w_dff_A_G4vSpu0G5_0),.din(w_dff_A_1qFCwSei7_0),.clk(gclk));
	jdff dff_A_G4vSpu0G5_0(.dout(w_dff_A_wE2z1JIn6_0),.din(w_dff_A_G4vSpu0G5_0),.clk(gclk));
	jdff dff_A_wE2z1JIn6_0(.dout(w_dff_A_bcaSGDxa1_0),.din(w_dff_A_wE2z1JIn6_0),.clk(gclk));
	jdff dff_A_bcaSGDxa1_0(.dout(w_dff_A_JKQi14PJ0_0),.din(w_dff_A_bcaSGDxa1_0),.clk(gclk));
	jdff dff_A_JKQi14PJ0_0(.dout(w_dff_A_C0DiUZfg5_0),.din(w_dff_A_JKQi14PJ0_0),.clk(gclk));
	jdff dff_A_C0DiUZfg5_0(.dout(w_dff_A_XkoFf4qk1_0),.din(w_dff_A_C0DiUZfg5_0),.clk(gclk));
	jdff dff_A_XkoFf4qk1_0(.dout(w_dff_A_Sb6cXqc88_0),.din(w_dff_A_XkoFf4qk1_0),.clk(gclk));
	jdff dff_A_Sb6cXqc88_0(.dout(w_dff_A_HXKwbOBe7_0),.din(w_dff_A_Sb6cXqc88_0),.clk(gclk));
	jdff dff_A_HXKwbOBe7_0(.dout(w_dff_A_SsSbmzrP0_0),.din(w_dff_A_HXKwbOBe7_0),.clk(gclk));
	jdff dff_A_SsSbmzrP0_0(.dout(w_dff_A_fT3hszoY9_0),.din(w_dff_A_SsSbmzrP0_0),.clk(gclk));
	jdff dff_A_fT3hszoY9_0(.dout(w_dff_A_4jYnIGsu8_0),.din(w_dff_A_fT3hszoY9_0),.clk(gclk));
	jdff dff_A_4jYnIGsu8_0(.dout(w_dff_A_mSQhwvnh6_0),.din(w_dff_A_4jYnIGsu8_0),.clk(gclk));
	jdff dff_A_mSQhwvnh6_0(.dout(w_dff_A_R2BG7Hr51_0),.din(w_dff_A_mSQhwvnh6_0),.clk(gclk));
	jdff dff_A_R2BG7Hr51_0(.dout(w_dff_A_qiy3e5fv6_0),.din(w_dff_A_R2BG7Hr51_0),.clk(gclk));
	jdff dff_A_qiy3e5fv6_0(.dout(w_dff_A_v4Qi1qBk1_0),.din(w_dff_A_qiy3e5fv6_0),.clk(gclk));
	jdff dff_A_v4Qi1qBk1_0(.dout(w_dff_A_DZwuPhxq7_0),.din(w_dff_A_v4Qi1qBk1_0),.clk(gclk));
	jdff dff_A_DZwuPhxq7_0(.dout(w_dff_A_gcSvZpbq3_0),.din(w_dff_A_DZwuPhxq7_0),.clk(gclk));
	jdff dff_A_gcSvZpbq3_0(.dout(w_dff_A_h2PKgTfh5_0),.din(w_dff_A_gcSvZpbq3_0),.clk(gclk));
	jdff dff_A_h2PKgTfh5_0(.dout(G554),.din(w_dff_A_h2PKgTfh5_0),.clk(gclk));
	jdff dff_A_SwcSZ5mu2_1(.dout(w_dff_A_I5TtFsPO3_0),.din(w_dff_A_SwcSZ5mu2_1),.clk(gclk));
	jdff dff_A_I5TtFsPO3_0(.dout(w_dff_A_I7sBW1ym7_0),.din(w_dff_A_I5TtFsPO3_0),.clk(gclk));
	jdff dff_A_I7sBW1ym7_0(.dout(w_dff_A_8nuYlqo78_0),.din(w_dff_A_I7sBW1ym7_0),.clk(gclk));
	jdff dff_A_8nuYlqo78_0(.dout(w_dff_A_H1pT0KGG1_0),.din(w_dff_A_8nuYlqo78_0),.clk(gclk));
	jdff dff_A_H1pT0KGG1_0(.dout(w_dff_A_mTgeVoxi5_0),.din(w_dff_A_H1pT0KGG1_0),.clk(gclk));
	jdff dff_A_mTgeVoxi5_0(.dout(w_dff_A_r4j6ACKh3_0),.din(w_dff_A_mTgeVoxi5_0),.clk(gclk));
	jdff dff_A_r4j6ACKh3_0(.dout(w_dff_A_OpoqpKPM1_0),.din(w_dff_A_r4j6ACKh3_0),.clk(gclk));
	jdff dff_A_OpoqpKPM1_0(.dout(w_dff_A_JlLzhrCR7_0),.din(w_dff_A_OpoqpKPM1_0),.clk(gclk));
	jdff dff_A_JlLzhrCR7_0(.dout(w_dff_A_1NKXrdeO7_0),.din(w_dff_A_JlLzhrCR7_0),.clk(gclk));
	jdff dff_A_1NKXrdeO7_0(.dout(w_dff_A_FY8pf0bB7_0),.din(w_dff_A_1NKXrdeO7_0),.clk(gclk));
	jdff dff_A_FY8pf0bB7_0(.dout(w_dff_A_qNhI5oZQ8_0),.din(w_dff_A_FY8pf0bB7_0),.clk(gclk));
	jdff dff_A_qNhI5oZQ8_0(.dout(w_dff_A_ex65tSP45_0),.din(w_dff_A_qNhI5oZQ8_0),.clk(gclk));
	jdff dff_A_ex65tSP45_0(.dout(w_dff_A_LzjMLhai6_0),.din(w_dff_A_ex65tSP45_0),.clk(gclk));
	jdff dff_A_LzjMLhai6_0(.dout(w_dff_A_0s70ksDY3_0),.din(w_dff_A_LzjMLhai6_0),.clk(gclk));
	jdff dff_A_0s70ksDY3_0(.dout(w_dff_A_eahvI2Tw5_0),.din(w_dff_A_0s70ksDY3_0),.clk(gclk));
	jdff dff_A_eahvI2Tw5_0(.dout(w_dff_A_O5ChEaQ90_0),.din(w_dff_A_eahvI2Tw5_0),.clk(gclk));
	jdff dff_A_O5ChEaQ90_0(.dout(w_dff_A_xUzzNqTC1_0),.din(w_dff_A_O5ChEaQ90_0),.clk(gclk));
	jdff dff_A_xUzzNqTC1_0(.dout(w_dff_A_JTDcJUGE2_0),.din(w_dff_A_xUzzNqTC1_0),.clk(gclk));
	jdff dff_A_JTDcJUGE2_0(.dout(w_dff_A_OrQMIMW96_0),.din(w_dff_A_JTDcJUGE2_0),.clk(gclk));
	jdff dff_A_OrQMIMW96_0(.dout(w_dff_A_Z0MWjToV7_0),.din(w_dff_A_OrQMIMW96_0),.clk(gclk));
	jdff dff_A_Z0MWjToV7_0(.dout(w_dff_A_asxkmu0C6_0),.din(w_dff_A_Z0MWjToV7_0),.clk(gclk));
	jdff dff_A_asxkmu0C6_0(.dout(w_dff_A_CnTbIlim7_0),.din(w_dff_A_asxkmu0C6_0),.clk(gclk));
	jdff dff_A_CnTbIlim7_0(.dout(w_dff_A_5eOxR1ck5_0),.din(w_dff_A_CnTbIlim7_0),.clk(gclk));
	jdff dff_A_5eOxR1ck5_0(.dout(w_dff_A_YRco1Ivp7_0),.din(w_dff_A_5eOxR1ck5_0),.clk(gclk));
	jdff dff_A_YRco1Ivp7_0(.dout(w_dff_A_WqGolFye2_0),.din(w_dff_A_YRco1Ivp7_0),.clk(gclk));
	jdff dff_A_WqGolFye2_0(.dout(G552),.din(w_dff_A_WqGolFye2_0),.clk(gclk));
	jdff dff_A_UOFpF7hR0_1(.dout(w_dff_A_DFmfw6vG3_0),.din(w_dff_A_UOFpF7hR0_1),.clk(gclk));
	jdff dff_A_DFmfw6vG3_0(.dout(w_dff_A_ne2TrUOm7_0),.din(w_dff_A_DFmfw6vG3_0),.clk(gclk));
	jdff dff_A_ne2TrUOm7_0(.dout(w_dff_A_HixFBzjI3_0),.din(w_dff_A_ne2TrUOm7_0),.clk(gclk));
	jdff dff_A_HixFBzjI3_0(.dout(w_dff_A_NtJ9bVEG1_0),.din(w_dff_A_HixFBzjI3_0),.clk(gclk));
	jdff dff_A_NtJ9bVEG1_0(.dout(w_dff_A_QP80W6xl8_0),.din(w_dff_A_NtJ9bVEG1_0),.clk(gclk));
	jdff dff_A_QP80W6xl8_0(.dout(w_dff_A_sufIrqeR3_0),.din(w_dff_A_QP80W6xl8_0),.clk(gclk));
	jdff dff_A_sufIrqeR3_0(.dout(w_dff_A_QHxrtEBw3_0),.din(w_dff_A_sufIrqeR3_0),.clk(gclk));
	jdff dff_A_QHxrtEBw3_0(.dout(w_dff_A_RmGhJCkc5_0),.din(w_dff_A_QHxrtEBw3_0),.clk(gclk));
	jdff dff_A_RmGhJCkc5_0(.dout(w_dff_A_gjMK7HsI2_0),.din(w_dff_A_RmGhJCkc5_0),.clk(gclk));
	jdff dff_A_gjMK7HsI2_0(.dout(w_dff_A_63XSR0MP2_0),.din(w_dff_A_gjMK7HsI2_0),.clk(gclk));
	jdff dff_A_63XSR0MP2_0(.dout(w_dff_A_ldZWNcFg1_0),.din(w_dff_A_63XSR0MP2_0),.clk(gclk));
	jdff dff_A_ldZWNcFg1_0(.dout(w_dff_A_sgeEwrXI0_0),.din(w_dff_A_ldZWNcFg1_0),.clk(gclk));
	jdff dff_A_sgeEwrXI0_0(.dout(w_dff_A_T1s58ywb7_0),.din(w_dff_A_sgeEwrXI0_0),.clk(gclk));
	jdff dff_A_T1s58ywb7_0(.dout(w_dff_A_cS2UAUHB4_0),.din(w_dff_A_T1s58ywb7_0),.clk(gclk));
	jdff dff_A_cS2UAUHB4_0(.dout(w_dff_A_hHRRzcPO5_0),.din(w_dff_A_cS2UAUHB4_0),.clk(gclk));
	jdff dff_A_hHRRzcPO5_0(.dout(w_dff_A_GMB2abC96_0),.din(w_dff_A_hHRRzcPO5_0),.clk(gclk));
	jdff dff_A_GMB2abC96_0(.dout(w_dff_A_SUMRqDyo5_0),.din(w_dff_A_GMB2abC96_0),.clk(gclk));
	jdff dff_A_SUMRqDyo5_0(.dout(w_dff_A_bdWj76Op9_0),.din(w_dff_A_SUMRqDyo5_0),.clk(gclk));
	jdff dff_A_bdWj76Op9_0(.dout(w_dff_A_DqUTDiHQ6_0),.din(w_dff_A_bdWj76Op9_0),.clk(gclk));
	jdff dff_A_DqUTDiHQ6_0(.dout(w_dff_A_2reMXbBq1_0),.din(w_dff_A_DqUTDiHQ6_0),.clk(gclk));
	jdff dff_A_2reMXbBq1_0(.dout(w_dff_A_h7KHJgaO4_0),.din(w_dff_A_2reMXbBq1_0),.clk(gclk));
	jdff dff_A_h7KHJgaO4_0(.dout(w_dff_A_dwLIIFPH4_0),.din(w_dff_A_h7KHJgaO4_0),.clk(gclk));
	jdff dff_A_dwLIIFPH4_0(.dout(w_dff_A_1Wbd86ql5_0),.din(w_dff_A_dwLIIFPH4_0),.clk(gclk));
	jdff dff_A_1Wbd86ql5_0(.dout(w_dff_A_E6XSqH0Y5_0),.din(w_dff_A_1Wbd86ql5_0),.clk(gclk));
	jdff dff_A_E6XSqH0Y5_0(.dout(w_dff_A_XzveyaxA5_0),.din(w_dff_A_E6XSqH0Y5_0),.clk(gclk));
	jdff dff_A_XzveyaxA5_0(.dout(G550),.din(w_dff_A_XzveyaxA5_0),.clk(gclk));
	jdff dff_A_3rAom8zd6_1(.dout(w_dff_A_fYXRzNNc1_0),.din(w_dff_A_3rAom8zd6_1),.clk(gclk));
	jdff dff_A_fYXRzNNc1_0(.dout(w_dff_A_Mtc00sxC0_0),.din(w_dff_A_fYXRzNNc1_0),.clk(gclk));
	jdff dff_A_Mtc00sxC0_0(.dout(w_dff_A_t5bc0efI2_0),.din(w_dff_A_Mtc00sxC0_0),.clk(gclk));
	jdff dff_A_t5bc0efI2_0(.dout(w_dff_A_C3oAI2Fi4_0),.din(w_dff_A_t5bc0efI2_0),.clk(gclk));
	jdff dff_A_C3oAI2Fi4_0(.dout(w_dff_A_FH2lil4W1_0),.din(w_dff_A_C3oAI2Fi4_0),.clk(gclk));
	jdff dff_A_FH2lil4W1_0(.dout(w_dff_A_QqZeptEe5_0),.din(w_dff_A_FH2lil4W1_0),.clk(gclk));
	jdff dff_A_QqZeptEe5_0(.dout(w_dff_A_BvkR98yw1_0),.din(w_dff_A_QqZeptEe5_0),.clk(gclk));
	jdff dff_A_BvkR98yw1_0(.dout(w_dff_A_wBytA4eS0_0),.din(w_dff_A_BvkR98yw1_0),.clk(gclk));
	jdff dff_A_wBytA4eS0_0(.dout(w_dff_A_W1Nj9btQ3_0),.din(w_dff_A_wBytA4eS0_0),.clk(gclk));
	jdff dff_A_W1Nj9btQ3_0(.dout(w_dff_A_WIoNprCO3_0),.din(w_dff_A_W1Nj9btQ3_0),.clk(gclk));
	jdff dff_A_WIoNprCO3_0(.dout(w_dff_A_oTH6z8ii4_0),.din(w_dff_A_WIoNprCO3_0),.clk(gclk));
	jdff dff_A_oTH6z8ii4_0(.dout(w_dff_A_iNIdyMhq9_0),.din(w_dff_A_oTH6z8ii4_0),.clk(gclk));
	jdff dff_A_iNIdyMhq9_0(.dout(w_dff_A_wr3GPQIf2_0),.din(w_dff_A_iNIdyMhq9_0),.clk(gclk));
	jdff dff_A_wr3GPQIf2_0(.dout(w_dff_A_RN5oxCKr4_0),.din(w_dff_A_wr3GPQIf2_0),.clk(gclk));
	jdff dff_A_RN5oxCKr4_0(.dout(w_dff_A_GBLQJdzc8_0),.din(w_dff_A_RN5oxCKr4_0),.clk(gclk));
	jdff dff_A_GBLQJdzc8_0(.dout(w_dff_A_6GrH231a8_0),.din(w_dff_A_GBLQJdzc8_0),.clk(gclk));
	jdff dff_A_6GrH231a8_0(.dout(w_dff_A_LzCj4MQa3_0),.din(w_dff_A_6GrH231a8_0),.clk(gclk));
	jdff dff_A_LzCj4MQa3_0(.dout(w_dff_A_YNuIQ53q7_0),.din(w_dff_A_LzCj4MQa3_0),.clk(gclk));
	jdff dff_A_YNuIQ53q7_0(.dout(w_dff_A_Qv19K5je0_0),.din(w_dff_A_YNuIQ53q7_0),.clk(gclk));
	jdff dff_A_Qv19K5je0_0(.dout(w_dff_A_uVgXRt9m1_0),.din(w_dff_A_Qv19K5je0_0),.clk(gclk));
	jdff dff_A_uVgXRt9m1_0(.dout(w_dff_A_0fqMLhtF9_0),.din(w_dff_A_uVgXRt9m1_0),.clk(gclk));
	jdff dff_A_0fqMLhtF9_0(.dout(w_dff_A_IxknPB2B0_0),.din(w_dff_A_0fqMLhtF9_0),.clk(gclk));
	jdff dff_A_IxknPB2B0_0(.dout(w_dff_A_lDRYKVjv0_0),.din(w_dff_A_IxknPB2B0_0),.clk(gclk));
	jdff dff_A_lDRYKVjv0_0(.dout(w_dff_A_rfayoZ0G4_0),.din(w_dff_A_lDRYKVjv0_0),.clk(gclk));
	jdff dff_A_rfayoZ0G4_0(.dout(w_dff_A_HGvALjB69_0),.din(w_dff_A_rfayoZ0G4_0),.clk(gclk));
	jdff dff_A_HGvALjB69_0(.dout(G548),.din(w_dff_A_HGvALjB69_0),.clk(gclk));
	jdff dff_A_jC7At71Q2_1(.dout(w_dff_A_LxBBIU8o3_0),.din(w_dff_A_jC7At71Q2_1),.clk(gclk));
	jdff dff_A_LxBBIU8o3_0(.dout(w_dff_A_r9UDQrDN1_0),.din(w_dff_A_LxBBIU8o3_0),.clk(gclk));
	jdff dff_A_r9UDQrDN1_0(.dout(w_dff_A_FkUvftfL8_0),.din(w_dff_A_r9UDQrDN1_0),.clk(gclk));
	jdff dff_A_FkUvftfL8_0(.dout(w_dff_A_tDVD6uAd0_0),.din(w_dff_A_FkUvftfL8_0),.clk(gclk));
	jdff dff_A_tDVD6uAd0_0(.dout(w_dff_A_ujznNtWB1_0),.din(w_dff_A_tDVD6uAd0_0),.clk(gclk));
	jdff dff_A_ujznNtWB1_0(.dout(w_dff_A_9u2bSJuP0_0),.din(w_dff_A_ujznNtWB1_0),.clk(gclk));
	jdff dff_A_9u2bSJuP0_0(.dout(w_dff_A_6A8laloR9_0),.din(w_dff_A_9u2bSJuP0_0),.clk(gclk));
	jdff dff_A_6A8laloR9_0(.dout(w_dff_A_4bnnsnk34_0),.din(w_dff_A_6A8laloR9_0),.clk(gclk));
	jdff dff_A_4bnnsnk34_0(.dout(w_dff_A_hCILH0XJ5_0),.din(w_dff_A_4bnnsnk34_0),.clk(gclk));
	jdff dff_A_hCILH0XJ5_0(.dout(w_dff_A_8E1PgMP80_0),.din(w_dff_A_hCILH0XJ5_0),.clk(gclk));
	jdff dff_A_8E1PgMP80_0(.dout(w_dff_A_cOc4c2bI7_0),.din(w_dff_A_8E1PgMP80_0),.clk(gclk));
	jdff dff_A_cOc4c2bI7_0(.dout(w_dff_A_it3y7hed1_0),.din(w_dff_A_cOc4c2bI7_0),.clk(gclk));
	jdff dff_A_it3y7hed1_0(.dout(w_dff_A_GhWC7yu38_0),.din(w_dff_A_it3y7hed1_0),.clk(gclk));
	jdff dff_A_GhWC7yu38_0(.dout(w_dff_A_H5skBDB29_0),.din(w_dff_A_GhWC7yu38_0),.clk(gclk));
	jdff dff_A_H5skBDB29_0(.dout(w_dff_A_6obFelOy3_0),.din(w_dff_A_H5skBDB29_0),.clk(gclk));
	jdff dff_A_6obFelOy3_0(.dout(w_dff_A_cJ7KDIQ20_0),.din(w_dff_A_6obFelOy3_0),.clk(gclk));
	jdff dff_A_cJ7KDIQ20_0(.dout(w_dff_A_9qrHKiPs2_0),.din(w_dff_A_cJ7KDIQ20_0),.clk(gclk));
	jdff dff_A_9qrHKiPs2_0(.dout(w_dff_A_yclbE7nM1_0),.din(w_dff_A_9qrHKiPs2_0),.clk(gclk));
	jdff dff_A_yclbE7nM1_0(.dout(w_dff_A_WHkxj6nR7_0),.din(w_dff_A_yclbE7nM1_0),.clk(gclk));
	jdff dff_A_WHkxj6nR7_0(.dout(w_dff_A_ADqu8nAL5_0),.din(w_dff_A_WHkxj6nR7_0),.clk(gclk));
	jdff dff_A_ADqu8nAL5_0(.dout(w_dff_A_wvVlABbh6_0),.din(w_dff_A_ADqu8nAL5_0),.clk(gclk));
	jdff dff_A_wvVlABbh6_0(.dout(w_dff_A_V6m99F9k9_0),.din(w_dff_A_wvVlABbh6_0),.clk(gclk));
	jdff dff_A_V6m99F9k9_0(.dout(w_dff_A_iGzYGW3S4_0),.din(w_dff_A_V6m99F9k9_0),.clk(gclk));
	jdff dff_A_iGzYGW3S4_0(.dout(w_dff_A_L4fSNyRt2_0),.din(w_dff_A_iGzYGW3S4_0),.clk(gclk));
	jdff dff_A_L4fSNyRt2_0(.dout(w_dff_A_Cu3qY5nH9_0),.din(w_dff_A_L4fSNyRt2_0),.clk(gclk));
	jdff dff_A_Cu3qY5nH9_0(.dout(G546),.din(w_dff_A_Cu3qY5nH9_0),.clk(gclk));
	jdff dff_A_O7RMNuf06_1(.dout(w_dff_A_doiTLMWg7_0),.din(w_dff_A_O7RMNuf06_1),.clk(gclk));
	jdff dff_A_doiTLMWg7_0(.dout(w_dff_A_pg5VpNzU3_0),.din(w_dff_A_doiTLMWg7_0),.clk(gclk));
	jdff dff_A_pg5VpNzU3_0(.dout(w_dff_A_uWjlNu2E3_0),.din(w_dff_A_pg5VpNzU3_0),.clk(gclk));
	jdff dff_A_uWjlNu2E3_0(.dout(w_dff_A_ljXNqORV6_0),.din(w_dff_A_uWjlNu2E3_0),.clk(gclk));
	jdff dff_A_ljXNqORV6_0(.dout(w_dff_A_WqFnMp7F1_0),.din(w_dff_A_ljXNqORV6_0),.clk(gclk));
	jdff dff_A_WqFnMp7F1_0(.dout(w_dff_A_yIgB1hws4_0),.din(w_dff_A_WqFnMp7F1_0),.clk(gclk));
	jdff dff_A_yIgB1hws4_0(.dout(w_dff_A_3Mn7T0Mc1_0),.din(w_dff_A_yIgB1hws4_0),.clk(gclk));
	jdff dff_A_3Mn7T0Mc1_0(.dout(w_dff_A_vKDjREg19_0),.din(w_dff_A_3Mn7T0Mc1_0),.clk(gclk));
	jdff dff_A_vKDjREg19_0(.dout(w_dff_A_y6BvsBzb5_0),.din(w_dff_A_vKDjREg19_0),.clk(gclk));
	jdff dff_A_y6BvsBzb5_0(.dout(w_dff_A_JefxyndS9_0),.din(w_dff_A_y6BvsBzb5_0),.clk(gclk));
	jdff dff_A_JefxyndS9_0(.dout(w_dff_A_OWHgQ3gL0_0),.din(w_dff_A_JefxyndS9_0),.clk(gclk));
	jdff dff_A_OWHgQ3gL0_0(.dout(w_dff_A_w8U8XJOq5_0),.din(w_dff_A_OWHgQ3gL0_0),.clk(gclk));
	jdff dff_A_w8U8XJOq5_0(.dout(w_dff_A_QbVkguio0_0),.din(w_dff_A_w8U8XJOq5_0),.clk(gclk));
	jdff dff_A_QbVkguio0_0(.dout(w_dff_A_NT8Dk4SR2_0),.din(w_dff_A_QbVkguio0_0),.clk(gclk));
	jdff dff_A_NT8Dk4SR2_0(.dout(w_dff_A_aRnnqE9j7_0),.din(w_dff_A_NT8Dk4SR2_0),.clk(gclk));
	jdff dff_A_aRnnqE9j7_0(.dout(w_dff_A_jkl0cphT9_0),.din(w_dff_A_aRnnqE9j7_0),.clk(gclk));
	jdff dff_A_jkl0cphT9_0(.dout(w_dff_A_MIVY0kBj5_0),.din(w_dff_A_jkl0cphT9_0),.clk(gclk));
	jdff dff_A_MIVY0kBj5_0(.dout(w_dff_A_I2AoVKde4_0),.din(w_dff_A_MIVY0kBj5_0),.clk(gclk));
	jdff dff_A_I2AoVKde4_0(.dout(w_dff_A_4pytqjya8_0),.din(w_dff_A_I2AoVKde4_0),.clk(gclk));
	jdff dff_A_4pytqjya8_0(.dout(w_dff_A_EP2uysYu8_0),.din(w_dff_A_4pytqjya8_0),.clk(gclk));
	jdff dff_A_EP2uysYu8_0(.dout(w_dff_A_OylISZWJ4_0),.din(w_dff_A_EP2uysYu8_0),.clk(gclk));
	jdff dff_A_OylISZWJ4_0(.dout(w_dff_A_U3RlEzgC0_0),.din(w_dff_A_OylISZWJ4_0),.clk(gclk));
	jdff dff_A_U3RlEzgC0_0(.dout(w_dff_A_SkPYBmGP8_0),.din(w_dff_A_U3RlEzgC0_0),.clk(gclk));
	jdff dff_A_SkPYBmGP8_0(.dout(w_dff_A_fDWQvJ6h5_0),.din(w_dff_A_SkPYBmGP8_0),.clk(gclk));
	jdff dff_A_fDWQvJ6h5_0(.dout(w_dff_A_6MiqYO5M0_0),.din(w_dff_A_fDWQvJ6h5_0),.clk(gclk));
	jdff dff_A_6MiqYO5M0_0(.dout(G544),.din(w_dff_A_6MiqYO5M0_0),.clk(gclk));
	jdff dff_A_cykvuITa8_1(.dout(w_dff_A_770ukYv22_0),.din(w_dff_A_cykvuITa8_1),.clk(gclk));
	jdff dff_A_770ukYv22_0(.dout(w_dff_A_aJRWQdhK0_0),.din(w_dff_A_770ukYv22_0),.clk(gclk));
	jdff dff_A_aJRWQdhK0_0(.dout(w_dff_A_lKFzJtcr0_0),.din(w_dff_A_aJRWQdhK0_0),.clk(gclk));
	jdff dff_A_lKFzJtcr0_0(.dout(w_dff_A_q9bJKAqu5_0),.din(w_dff_A_lKFzJtcr0_0),.clk(gclk));
	jdff dff_A_q9bJKAqu5_0(.dout(w_dff_A_zVZkXWJq6_0),.din(w_dff_A_q9bJKAqu5_0),.clk(gclk));
	jdff dff_A_zVZkXWJq6_0(.dout(w_dff_A_xo0s4Jdx9_0),.din(w_dff_A_zVZkXWJq6_0),.clk(gclk));
	jdff dff_A_xo0s4Jdx9_0(.dout(w_dff_A_qYZ9UaqO6_0),.din(w_dff_A_xo0s4Jdx9_0),.clk(gclk));
	jdff dff_A_qYZ9UaqO6_0(.dout(w_dff_A_zeNUlbEx4_0),.din(w_dff_A_qYZ9UaqO6_0),.clk(gclk));
	jdff dff_A_zeNUlbEx4_0(.dout(w_dff_A_WqjG7eI77_0),.din(w_dff_A_zeNUlbEx4_0),.clk(gclk));
	jdff dff_A_WqjG7eI77_0(.dout(w_dff_A_1Zn3Ue1k8_0),.din(w_dff_A_WqjG7eI77_0),.clk(gclk));
	jdff dff_A_1Zn3Ue1k8_0(.dout(w_dff_A_u1bfDX7C2_0),.din(w_dff_A_1Zn3Ue1k8_0),.clk(gclk));
	jdff dff_A_u1bfDX7C2_0(.dout(w_dff_A_E1CkVYeH5_0),.din(w_dff_A_u1bfDX7C2_0),.clk(gclk));
	jdff dff_A_E1CkVYeH5_0(.dout(w_dff_A_TymXuwcy5_0),.din(w_dff_A_E1CkVYeH5_0),.clk(gclk));
	jdff dff_A_TymXuwcy5_0(.dout(w_dff_A_wG4UJRUV2_0),.din(w_dff_A_TymXuwcy5_0),.clk(gclk));
	jdff dff_A_wG4UJRUV2_0(.dout(w_dff_A_DMadvdJh4_0),.din(w_dff_A_wG4UJRUV2_0),.clk(gclk));
	jdff dff_A_DMadvdJh4_0(.dout(w_dff_A_bM89scTp8_0),.din(w_dff_A_DMadvdJh4_0),.clk(gclk));
	jdff dff_A_bM89scTp8_0(.dout(w_dff_A_jUY7NL5b5_0),.din(w_dff_A_bM89scTp8_0),.clk(gclk));
	jdff dff_A_jUY7NL5b5_0(.dout(w_dff_A_aMmGBlsD6_0),.din(w_dff_A_jUY7NL5b5_0),.clk(gclk));
	jdff dff_A_aMmGBlsD6_0(.dout(w_dff_A_s7grm0hQ4_0),.din(w_dff_A_aMmGBlsD6_0),.clk(gclk));
	jdff dff_A_s7grm0hQ4_0(.dout(w_dff_A_56FFMSOa8_0),.din(w_dff_A_s7grm0hQ4_0),.clk(gclk));
	jdff dff_A_56FFMSOa8_0(.dout(w_dff_A_VhFAjZOL5_0),.din(w_dff_A_56FFMSOa8_0),.clk(gclk));
	jdff dff_A_VhFAjZOL5_0(.dout(w_dff_A_rSbD6nUO1_0),.din(w_dff_A_VhFAjZOL5_0),.clk(gclk));
	jdff dff_A_rSbD6nUO1_0(.dout(w_dff_A_4S3Q3aPN4_0),.din(w_dff_A_rSbD6nUO1_0),.clk(gclk));
	jdff dff_A_4S3Q3aPN4_0(.dout(w_dff_A_f2bmOJli8_0),.din(w_dff_A_4S3Q3aPN4_0),.clk(gclk));
	jdff dff_A_f2bmOJli8_0(.dout(w_dff_A_Ub6SdZnE2_0),.din(w_dff_A_f2bmOJli8_0),.clk(gclk));
	jdff dff_A_Ub6SdZnE2_0(.dout(G540),.din(w_dff_A_Ub6SdZnE2_0),.clk(gclk));
	jdff dff_A_ZmdyHmdd8_1(.dout(w_dff_A_mcWpOpJu8_0),.din(w_dff_A_ZmdyHmdd8_1),.clk(gclk));
	jdff dff_A_mcWpOpJu8_0(.dout(w_dff_A_JAMipuF20_0),.din(w_dff_A_mcWpOpJu8_0),.clk(gclk));
	jdff dff_A_JAMipuF20_0(.dout(w_dff_A_lcdRUCoI8_0),.din(w_dff_A_JAMipuF20_0),.clk(gclk));
	jdff dff_A_lcdRUCoI8_0(.dout(w_dff_A_l0sFi7ci9_0),.din(w_dff_A_lcdRUCoI8_0),.clk(gclk));
	jdff dff_A_l0sFi7ci9_0(.dout(w_dff_A_14pZ2zFV1_0),.din(w_dff_A_l0sFi7ci9_0),.clk(gclk));
	jdff dff_A_14pZ2zFV1_0(.dout(w_dff_A_kM4IefWL3_0),.din(w_dff_A_14pZ2zFV1_0),.clk(gclk));
	jdff dff_A_kM4IefWL3_0(.dout(w_dff_A_3SC9EuCc1_0),.din(w_dff_A_kM4IefWL3_0),.clk(gclk));
	jdff dff_A_3SC9EuCc1_0(.dout(w_dff_A_p9rERASQ0_0),.din(w_dff_A_3SC9EuCc1_0),.clk(gclk));
	jdff dff_A_p9rERASQ0_0(.dout(w_dff_A_w18NPP820_0),.din(w_dff_A_p9rERASQ0_0),.clk(gclk));
	jdff dff_A_w18NPP820_0(.dout(w_dff_A_xQNOfzUB7_0),.din(w_dff_A_w18NPP820_0),.clk(gclk));
	jdff dff_A_xQNOfzUB7_0(.dout(w_dff_A_z1NqDnVO2_0),.din(w_dff_A_xQNOfzUB7_0),.clk(gclk));
	jdff dff_A_z1NqDnVO2_0(.dout(w_dff_A_Pznzn9Fh9_0),.din(w_dff_A_z1NqDnVO2_0),.clk(gclk));
	jdff dff_A_Pznzn9Fh9_0(.dout(w_dff_A_RnIBIxir5_0),.din(w_dff_A_Pznzn9Fh9_0),.clk(gclk));
	jdff dff_A_RnIBIxir5_0(.dout(w_dff_A_bilz34lm8_0),.din(w_dff_A_RnIBIxir5_0),.clk(gclk));
	jdff dff_A_bilz34lm8_0(.dout(w_dff_A_AefvOYKG9_0),.din(w_dff_A_bilz34lm8_0),.clk(gclk));
	jdff dff_A_AefvOYKG9_0(.dout(w_dff_A_DhX6PBLq1_0),.din(w_dff_A_AefvOYKG9_0),.clk(gclk));
	jdff dff_A_DhX6PBLq1_0(.dout(w_dff_A_7kpp6Y2X0_0),.din(w_dff_A_DhX6PBLq1_0),.clk(gclk));
	jdff dff_A_7kpp6Y2X0_0(.dout(w_dff_A_il0yoA8c2_0),.din(w_dff_A_7kpp6Y2X0_0),.clk(gclk));
	jdff dff_A_il0yoA8c2_0(.dout(w_dff_A_VNUV6xRn4_0),.din(w_dff_A_il0yoA8c2_0),.clk(gclk));
	jdff dff_A_VNUV6xRn4_0(.dout(w_dff_A_UsKiHWMT2_0),.din(w_dff_A_VNUV6xRn4_0),.clk(gclk));
	jdff dff_A_UsKiHWMT2_0(.dout(w_dff_A_RhI2wq0z5_0),.din(w_dff_A_UsKiHWMT2_0),.clk(gclk));
	jdff dff_A_RhI2wq0z5_0(.dout(w_dff_A_NTf5VPGD7_0),.din(w_dff_A_RhI2wq0z5_0),.clk(gclk));
	jdff dff_A_NTf5VPGD7_0(.dout(w_dff_A_bTcdFqlR5_0),.din(w_dff_A_NTf5VPGD7_0),.clk(gclk));
	jdff dff_A_bTcdFqlR5_0(.dout(w_dff_A_1E3cOk3U5_0),.din(w_dff_A_bTcdFqlR5_0),.clk(gclk));
	jdff dff_A_1E3cOk3U5_0(.dout(w_dff_A_6latRHez4_0),.din(w_dff_A_1E3cOk3U5_0),.clk(gclk));
	jdff dff_A_6latRHez4_0(.dout(G538),.din(w_dff_A_6latRHez4_0),.clk(gclk));
	jdff dff_A_bVT2Wp258_1(.dout(w_dff_A_TWjxMiy76_0),.din(w_dff_A_bVT2Wp258_1),.clk(gclk));
	jdff dff_A_TWjxMiy76_0(.dout(w_dff_A_ZEcQB5Jl7_0),.din(w_dff_A_TWjxMiy76_0),.clk(gclk));
	jdff dff_A_ZEcQB5Jl7_0(.dout(w_dff_A_DNfbcwZX4_0),.din(w_dff_A_ZEcQB5Jl7_0),.clk(gclk));
	jdff dff_A_DNfbcwZX4_0(.dout(w_dff_A_rt1KetpS8_0),.din(w_dff_A_DNfbcwZX4_0),.clk(gclk));
	jdff dff_A_rt1KetpS8_0(.dout(w_dff_A_d83EbDdg2_0),.din(w_dff_A_rt1KetpS8_0),.clk(gclk));
	jdff dff_A_d83EbDdg2_0(.dout(w_dff_A_3bZAt0Hm5_0),.din(w_dff_A_d83EbDdg2_0),.clk(gclk));
	jdff dff_A_3bZAt0Hm5_0(.dout(w_dff_A_gBrCuvdu4_0),.din(w_dff_A_3bZAt0Hm5_0),.clk(gclk));
	jdff dff_A_gBrCuvdu4_0(.dout(w_dff_A_W5yMHXz95_0),.din(w_dff_A_gBrCuvdu4_0),.clk(gclk));
	jdff dff_A_W5yMHXz95_0(.dout(w_dff_A_ZZ9zmRnp3_0),.din(w_dff_A_W5yMHXz95_0),.clk(gclk));
	jdff dff_A_ZZ9zmRnp3_0(.dout(w_dff_A_31WN9WR89_0),.din(w_dff_A_ZZ9zmRnp3_0),.clk(gclk));
	jdff dff_A_31WN9WR89_0(.dout(w_dff_A_dGioZHas1_0),.din(w_dff_A_31WN9WR89_0),.clk(gclk));
	jdff dff_A_dGioZHas1_0(.dout(w_dff_A_NP4F7CHk5_0),.din(w_dff_A_dGioZHas1_0),.clk(gclk));
	jdff dff_A_NP4F7CHk5_0(.dout(w_dff_A_txfAdmnr5_0),.din(w_dff_A_NP4F7CHk5_0),.clk(gclk));
	jdff dff_A_txfAdmnr5_0(.dout(w_dff_A_dE6GOoFS8_0),.din(w_dff_A_txfAdmnr5_0),.clk(gclk));
	jdff dff_A_dE6GOoFS8_0(.dout(w_dff_A_bL9jkJr21_0),.din(w_dff_A_dE6GOoFS8_0),.clk(gclk));
	jdff dff_A_bL9jkJr21_0(.dout(w_dff_A_PCsnKyw47_0),.din(w_dff_A_bL9jkJr21_0),.clk(gclk));
	jdff dff_A_PCsnKyw47_0(.dout(w_dff_A_WKZ7MFIb3_0),.din(w_dff_A_PCsnKyw47_0),.clk(gclk));
	jdff dff_A_WKZ7MFIb3_0(.dout(w_dff_A_dehq0JxD4_0),.din(w_dff_A_WKZ7MFIb3_0),.clk(gclk));
	jdff dff_A_dehq0JxD4_0(.dout(w_dff_A_PRdaNg3o0_0),.din(w_dff_A_dehq0JxD4_0),.clk(gclk));
	jdff dff_A_PRdaNg3o0_0(.dout(w_dff_A_73lR5fPK3_0),.din(w_dff_A_PRdaNg3o0_0),.clk(gclk));
	jdff dff_A_73lR5fPK3_0(.dout(w_dff_A_BwZ9htRo1_0),.din(w_dff_A_73lR5fPK3_0),.clk(gclk));
	jdff dff_A_BwZ9htRo1_0(.dout(w_dff_A_VUwT3GaX3_0),.din(w_dff_A_BwZ9htRo1_0),.clk(gclk));
	jdff dff_A_VUwT3GaX3_0(.dout(w_dff_A_apxQIS8p5_0),.din(w_dff_A_VUwT3GaX3_0),.clk(gclk));
	jdff dff_A_apxQIS8p5_0(.dout(w_dff_A_CK0UtfAN4_0),.din(w_dff_A_apxQIS8p5_0),.clk(gclk));
	jdff dff_A_CK0UtfAN4_0(.dout(w_dff_A_9vdyOd9n5_0),.din(w_dff_A_CK0UtfAN4_0),.clk(gclk));
	jdff dff_A_9vdyOd9n5_0(.dout(G536),.din(w_dff_A_9vdyOd9n5_0),.clk(gclk));
	jdff dff_A_1ISwIh973_1(.dout(w_dff_A_xxcJnGPc1_0),.din(w_dff_A_1ISwIh973_1),.clk(gclk));
	jdff dff_A_xxcJnGPc1_0(.dout(w_dff_A_1f89aRfw3_0),.din(w_dff_A_xxcJnGPc1_0),.clk(gclk));
	jdff dff_A_1f89aRfw3_0(.dout(w_dff_A_zaiDhMWa6_0),.din(w_dff_A_1f89aRfw3_0),.clk(gclk));
	jdff dff_A_zaiDhMWa6_0(.dout(w_dff_A_xlZk6Hun3_0),.din(w_dff_A_zaiDhMWa6_0),.clk(gclk));
	jdff dff_A_xlZk6Hun3_0(.dout(w_dff_A_IiRPdPLX1_0),.din(w_dff_A_xlZk6Hun3_0),.clk(gclk));
	jdff dff_A_IiRPdPLX1_0(.dout(w_dff_A_AmsLyTTL7_0),.din(w_dff_A_IiRPdPLX1_0),.clk(gclk));
	jdff dff_A_AmsLyTTL7_0(.dout(w_dff_A_UYH5WbYg5_0),.din(w_dff_A_AmsLyTTL7_0),.clk(gclk));
	jdff dff_A_UYH5WbYg5_0(.dout(w_dff_A_xzCKYHee1_0),.din(w_dff_A_UYH5WbYg5_0),.clk(gclk));
	jdff dff_A_xzCKYHee1_0(.dout(w_dff_A_F0ydn2vw7_0),.din(w_dff_A_xzCKYHee1_0),.clk(gclk));
	jdff dff_A_F0ydn2vw7_0(.dout(w_dff_A_lf1zOueQ8_0),.din(w_dff_A_F0ydn2vw7_0),.clk(gclk));
	jdff dff_A_lf1zOueQ8_0(.dout(w_dff_A_mrDtIXis0_0),.din(w_dff_A_lf1zOueQ8_0),.clk(gclk));
	jdff dff_A_mrDtIXis0_0(.dout(w_dff_A_CiyHWuyA4_0),.din(w_dff_A_mrDtIXis0_0),.clk(gclk));
	jdff dff_A_CiyHWuyA4_0(.dout(w_dff_A_5yH4yel01_0),.din(w_dff_A_CiyHWuyA4_0),.clk(gclk));
	jdff dff_A_5yH4yel01_0(.dout(w_dff_A_zLGMLEYs7_0),.din(w_dff_A_5yH4yel01_0),.clk(gclk));
	jdff dff_A_zLGMLEYs7_0(.dout(w_dff_A_V1JJ2rO97_0),.din(w_dff_A_zLGMLEYs7_0),.clk(gclk));
	jdff dff_A_V1JJ2rO97_0(.dout(w_dff_A_4oZSJe060_0),.din(w_dff_A_V1JJ2rO97_0),.clk(gclk));
	jdff dff_A_4oZSJe060_0(.dout(w_dff_A_t118G6i42_0),.din(w_dff_A_4oZSJe060_0),.clk(gclk));
	jdff dff_A_t118G6i42_0(.dout(w_dff_A_Ot5bP7Dg0_0),.din(w_dff_A_t118G6i42_0),.clk(gclk));
	jdff dff_A_Ot5bP7Dg0_0(.dout(w_dff_A_Ty92eDGb9_0),.din(w_dff_A_Ot5bP7Dg0_0),.clk(gclk));
	jdff dff_A_Ty92eDGb9_0(.dout(w_dff_A_qKlU8vAu5_0),.din(w_dff_A_Ty92eDGb9_0),.clk(gclk));
	jdff dff_A_qKlU8vAu5_0(.dout(w_dff_A_qzBzlYFR7_0),.din(w_dff_A_qKlU8vAu5_0),.clk(gclk));
	jdff dff_A_qzBzlYFR7_0(.dout(w_dff_A_qOnaJgEF2_0),.din(w_dff_A_qzBzlYFR7_0),.clk(gclk));
	jdff dff_A_qOnaJgEF2_0(.dout(w_dff_A_rP1B7lWF8_0),.din(w_dff_A_qOnaJgEF2_0),.clk(gclk));
	jdff dff_A_rP1B7lWF8_0(.dout(w_dff_A_qbRmjG5t1_0),.din(w_dff_A_rP1B7lWF8_0),.clk(gclk));
	jdff dff_A_qbRmjG5t1_0(.dout(w_dff_A_CAN7PF2s2_0),.din(w_dff_A_qbRmjG5t1_0),.clk(gclk));
	jdff dff_A_CAN7PF2s2_0(.dout(G534),.din(w_dff_A_CAN7PF2s2_0),.clk(gclk));
	jdff dff_A_uyVV29G02_1(.dout(w_dff_A_YpAS42Pd0_0),.din(w_dff_A_uyVV29G02_1),.clk(gclk));
	jdff dff_A_YpAS42Pd0_0(.dout(w_dff_A_aABiHqDV8_0),.din(w_dff_A_YpAS42Pd0_0),.clk(gclk));
	jdff dff_A_aABiHqDV8_0(.dout(w_dff_A_wUqlU6bb6_0),.din(w_dff_A_aABiHqDV8_0),.clk(gclk));
	jdff dff_A_wUqlU6bb6_0(.dout(w_dff_A_HpeNI6hu8_0),.din(w_dff_A_wUqlU6bb6_0),.clk(gclk));
	jdff dff_A_HpeNI6hu8_0(.dout(w_dff_A_31ifhgLe3_0),.din(w_dff_A_HpeNI6hu8_0),.clk(gclk));
	jdff dff_A_31ifhgLe3_0(.dout(w_dff_A_20LL0kXl3_0),.din(w_dff_A_31ifhgLe3_0),.clk(gclk));
	jdff dff_A_20LL0kXl3_0(.dout(w_dff_A_5frTfrNj9_0),.din(w_dff_A_20LL0kXl3_0),.clk(gclk));
	jdff dff_A_5frTfrNj9_0(.dout(w_dff_A_MnRCGrLU2_0),.din(w_dff_A_5frTfrNj9_0),.clk(gclk));
	jdff dff_A_MnRCGrLU2_0(.dout(w_dff_A_iyKzf2e81_0),.din(w_dff_A_MnRCGrLU2_0),.clk(gclk));
	jdff dff_A_iyKzf2e81_0(.dout(w_dff_A_bHVODOSr4_0),.din(w_dff_A_iyKzf2e81_0),.clk(gclk));
	jdff dff_A_bHVODOSr4_0(.dout(w_dff_A_BgMe5zfd0_0),.din(w_dff_A_bHVODOSr4_0),.clk(gclk));
	jdff dff_A_BgMe5zfd0_0(.dout(w_dff_A_IYQi4gKK1_0),.din(w_dff_A_BgMe5zfd0_0),.clk(gclk));
	jdff dff_A_IYQi4gKK1_0(.dout(w_dff_A_vyipA3Is1_0),.din(w_dff_A_IYQi4gKK1_0),.clk(gclk));
	jdff dff_A_vyipA3Is1_0(.dout(w_dff_A_QQxLPPac5_0),.din(w_dff_A_vyipA3Is1_0),.clk(gclk));
	jdff dff_A_QQxLPPac5_0(.dout(w_dff_A_bYELoScb0_0),.din(w_dff_A_QQxLPPac5_0),.clk(gclk));
	jdff dff_A_bYELoScb0_0(.dout(w_dff_A_zy7vFfa32_0),.din(w_dff_A_bYELoScb0_0),.clk(gclk));
	jdff dff_A_zy7vFfa32_0(.dout(w_dff_A_JDIrwvVA2_0),.din(w_dff_A_zy7vFfa32_0),.clk(gclk));
	jdff dff_A_JDIrwvVA2_0(.dout(w_dff_A_627Yje469_0),.din(w_dff_A_JDIrwvVA2_0),.clk(gclk));
	jdff dff_A_627Yje469_0(.dout(w_dff_A_TMA9OBaf5_0),.din(w_dff_A_627Yje469_0),.clk(gclk));
	jdff dff_A_TMA9OBaf5_0(.dout(w_dff_A_O8OwSJCu5_0),.din(w_dff_A_TMA9OBaf5_0),.clk(gclk));
	jdff dff_A_O8OwSJCu5_0(.dout(w_dff_A_wsyX4SW31_0),.din(w_dff_A_O8OwSJCu5_0),.clk(gclk));
	jdff dff_A_wsyX4SW31_0(.dout(w_dff_A_Y70sezAz6_0),.din(w_dff_A_wsyX4SW31_0),.clk(gclk));
	jdff dff_A_Y70sezAz6_0(.dout(w_dff_A_dc3tr08t9_0),.din(w_dff_A_Y70sezAz6_0),.clk(gclk));
	jdff dff_A_dc3tr08t9_0(.dout(w_dff_A_C1dJ18Gh8_0),.din(w_dff_A_dc3tr08t9_0),.clk(gclk));
	jdff dff_A_C1dJ18Gh8_0(.dout(w_dff_A_XzuygA3z9_0),.din(w_dff_A_C1dJ18Gh8_0),.clk(gclk));
	jdff dff_A_XzuygA3z9_0(.dout(G532),.din(w_dff_A_XzuygA3z9_0),.clk(gclk));
	jdff dff_A_paBQc1dR5_1(.dout(w_dff_A_KrKWbOFh4_0),.din(w_dff_A_paBQc1dR5_1),.clk(gclk));
	jdff dff_A_KrKWbOFh4_0(.dout(w_dff_A_owVCqCIt3_0),.din(w_dff_A_KrKWbOFh4_0),.clk(gclk));
	jdff dff_A_owVCqCIt3_0(.dout(w_dff_A_8tjNKYJW7_0),.din(w_dff_A_owVCqCIt3_0),.clk(gclk));
	jdff dff_A_8tjNKYJW7_0(.dout(w_dff_A_IKRWkruj3_0),.din(w_dff_A_8tjNKYJW7_0),.clk(gclk));
	jdff dff_A_IKRWkruj3_0(.dout(w_dff_A_7ILXqpvi9_0),.din(w_dff_A_IKRWkruj3_0),.clk(gclk));
	jdff dff_A_7ILXqpvi9_0(.dout(w_dff_A_9ssq8esx2_0),.din(w_dff_A_7ILXqpvi9_0),.clk(gclk));
	jdff dff_A_9ssq8esx2_0(.dout(w_dff_A_mz5ZwWi41_0),.din(w_dff_A_9ssq8esx2_0),.clk(gclk));
	jdff dff_A_mz5ZwWi41_0(.dout(w_dff_A_S3H3brTp1_0),.din(w_dff_A_mz5ZwWi41_0),.clk(gclk));
	jdff dff_A_S3H3brTp1_0(.dout(w_dff_A_R3hJPeZ30_0),.din(w_dff_A_S3H3brTp1_0),.clk(gclk));
	jdff dff_A_R3hJPeZ30_0(.dout(w_dff_A_M19Bz4np1_0),.din(w_dff_A_R3hJPeZ30_0),.clk(gclk));
	jdff dff_A_M19Bz4np1_0(.dout(w_dff_A_1xd8j4TM9_0),.din(w_dff_A_M19Bz4np1_0),.clk(gclk));
	jdff dff_A_1xd8j4TM9_0(.dout(w_dff_A_bjysYcGH5_0),.din(w_dff_A_1xd8j4TM9_0),.clk(gclk));
	jdff dff_A_bjysYcGH5_0(.dout(w_dff_A_yFlYAY4Q1_0),.din(w_dff_A_bjysYcGH5_0),.clk(gclk));
	jdff dff_A_yFlYAY4Q1_0(.dout(w_dff_A_Itab8r2P7_0),.din(w_dff_A_yFlYAY4Q1_0),.clk(gclk));
	jdff dff_A_Itab8r2P7_0(.dout(w_dff_A_nxHJwfuq2_0),.din(w_dff_A_Itab8r2P7_0),.clk(gclk));
	jdff dff_A_nxHJwfuq2_0(.dout(w_dff_A_qjpSuRHT0_0),.din(w_dff_A_nxHJwfuq2_0),.clk(gclk));
	jdff dff_A_qjpSuRHT0_0(.dout(w_dff_A_M21h6pYF5_0),.din(w_dff_A_qjpSuRHT0_0),.clk(gclk));
	jdff dff_A_M21h6pYF5_0(.dout(w_dff_A_meqkVuQd2_0),.din(w_dff_A_M21h6pYF5_0),.clk(gclk));
	jdff dff_A_meqkVuQd2_0(.dout(w_dff_A_1SqBkC2z1_0),.din(w_dff_A_meqkVuQd2_0),.clk(gclk));
	jdff dff_A_1SqBkC2z1_0(.dout(w_dff_A_mfmqXWB09_0),.din(w_dff_A_1SqBkC2z1_0),.clk(gclk));
	jdff dff_A_mfmqXWB09_0(.dout(w_dff_A_wkbJbniV5_0),.din(w_dff_A_mfmqXWB09_0),.clk(gclk));
	jdff dff_A_wkbJbniV5_0(.dout(w_dff_A_bDCKCygv0_0),.din(w_dff_A_wkbJbniV5_0),.clk(gclk));
	jdff dff_A_bDCKCygv0_0(.dout(w_dff_A_tRoI4P0z5_0),.din(w_dff_A_bDCKCygv0_0),.clk(gclk));
	jdff dff_A_tRoI4P0z5_0(.dout(w_dff_A_Ulamf9mu4_0),.din(w_dff_A_tRoI4P0z5_0),.clk(gclk));
	jdff dff_A_Ulamf9mu4_0(.dout(w_dff_A_DLzrrKos7_0),.din(w_dff_A_Ulamf9mu4_0),.clk(gclk));
	jdff dff_A_DLzrrKos7_0(.dout(G530),.din(w_dff_A_DLzrrKos7_0),.clk(gclk));
	jdff dff_A_BhtDhst74_1(.dout(w_dff_A_PAVZXrKf0_0),.din(w_dff_A_BhtDhst74_1),.clk(gclk));
	jdff dff_A_PAVZXrKf0_0(.dout(w_dff_A_01cYpg8b6_0),.din(w_dff_A_PAVZXrKf0_0),.clk(gclk));
	jdff dff_A_01cYpg8b6_0(.dout(w_dff_A_fajuVp6Z6_0),.din(w_dff_A_01cYpg8b6_0),.clk(gclk));
	jdff dff_A_fajuVp6Z6_0(.dout(w_dff_A_DJXiWyPe2_0),.din(w_dff_A_fajuVp6Z6_0),.clk(gclk));
	jdff dff_A_DJXiWyPe2_0(.dout(w_dff_A_dlsyUagO4_0),.din(w_dff_A_DJXiWyPe2_0),.clk(gclk));
	jdff dff_A_dlsyUagO4_0(.dout(w_dff_A_vmKx730D5_0),.din(w_dff_A_dlsyUagO4_0),.clk(gclk));
	jdff dff_A_vmKx730D5_0(.dout(w_dff_A_0RmeoFv85_0),.din(w_dff_A_vmKx730D5_0),.clk(gclk));
	jdff dff_A_0RmeoFv85_0(.dout(w_dff_A_IZaZ4JT98_0),.din(w_dff_A_0RmeoFv85_0),.clk(gclk));
	jdff dff_A_IZaZ4JT98_0(.dout(w_dff_A_o7wAR7Kf5_0),.din(w_dff_A_IZaZ4JT98_0),.clk(gclk));
	jdff dff_A_o7wAR7Kf5_0(.dout(w_dff_A_ZWrN8TAT6_0),.din(w_dff_A_o7wAR7Kf5_0),.clk(gclk));
	jdff dff_A_ZWrN8TAT6_0(.dout(w_dff_A_GC1pX1l39_0),.din(w_dff_A_ZWrN8TAT6_0),.clk(gclk));
	jdff dff_A_GC1pX1l39_0(.dout(w_dff_A_DAT3tjR14_0),.din(w_dff_A_GC1pX1l39_0),.clk(gclk));
	jdff dff_A_DAT3tjR14_0(.dout(w_dff_A_Lp3fWjAx2_0),.din(w_dff_A_DAT3tjR14_0),.clk(gclk));
	jdff dff_A_Lp3fWjAx2_0(.dout(w_dff_A_HhyK5uS78_0),.din(w_dff_A_Lp3fWjAx2_0),.clk(gclk));
	jdff dff_A_HhyK5uS78_0(.dout(w_dff_A_I6VdQDZF7_0),.din(w_dff_A_HhyK5uS78_0),.clk(gclk));
	jdff dff_A_I6VdQDZF7_0(.dout(w_dff_A_sBPhlIxo5_0),.din(w_dff_A_I6VdQDZF7_0),.clk(gclk));
	jdff dff_A_sBPhlIxo5_0(.dout(w_dff_A_gZb17gAj1_0),.din(w_dff_A_sBPhlIxo5_0),.clk(gclk));
	jdff dff_A_gZb17gAj1_0(.dout(w_dff_A_3eYdNwvV9_0),.din(w_dff_A_gZb17gAj1_0),.clk(gclk));
	jdff dff_A_3eYdNwvV9_0(.dout(w_dff_A_hKabU6aP9_0),.din(w_dff_A_3eYdNwvV9_0),.clk(gclk));
	jdff dff_A_hKabU6aP9_0(.dout(w_dff_A_GRmOsZCc2_0),.din(w_dff_A_hKabU6aP9_0),.clk(gclk));
	jdff dff_A_GRmOsZCc2_0(.dout(w_dff_A_jOt2u3W90_0),.din(w_dff_A_GRmOsZCc2_0),.clk(gclk));
	jdff dff_A_jOt2u3W90_0(.dout(w_dff_A_2nW35xZC6_0),.din(w_dff_A_jOt2u3W90_0),.clk(gclk));
	jdff dff_A_2nW35xZC6_0(.dout(w_dff_A_pEyMk4PZ2_0),.din(w_dff_A_2nW35xZC6_0),.clk(gclk));
	jdff dff_A_pEyMk4PZ2_0(.dout(w_dff_A_Ef2unXg22_0),.din(w_dff_A_pEyMk4PZ2_0),.clk(gclk));
	jdff dff_A_Ef2unXg22_0(.dout(w_dff_A_f6nhjreC0_0),.din(w_dff_A_Ef2unXg22_0),.clk(gclk));
	jdff dff_A_f6nhjreC0_0(.dout(G528),.din(w_dff_A_f6nhjreC0_0),.clk(gclk));
	jdff dff_A_xoVdo85w5_1(.dout(w_dff_A_5gDDdwws1_0),.din(w_dff_A_xoVdo85w5_1),.clk(gclk));
	jdff dff_A_5gDDdwws1_0(.dout(w_dff_A_tDSURJ8L5_0),.din(w_dff_A_5gDDdwws1_0),.clk(gclk));
	jdff dff_A_tDSURJ8L5_0(.dout(w_dff_A_7T47Z8Ee6_0),.din(w_dff_A_tDSURJ8L5_0),.clk(gclk));
	jdff dff_A_7T47Z8Ee6_0(.dout(w_dff_A_0qzoXbNm6_0),.din(w_dff_A_7T47Z8Ee6_0),.clk(gclk));
	jdff dff_A_0qzoXbNm6_0(.dout(w_dff_A_emAtNjXO1_0),.din(w_dff_A_0qzoXbNm6_0),.clk(gclk));
	jdff dff_A_emAtNjXO1_0(.dout(w_dff_A_Gm5iDwRD3_0),.din(w_dff_A_emAtNjXO1_0),.clk(gclk));
	jdff dff_A_Gm5iDwRD3_0(.dout(w_dff_A_ijIOBYxc4_0),.din(w_dff_A_Gm5iDwRD3_0),.clk(gclk));
	jdff dff_A_ijIOBYxc4_0(.dout(w_dff_A_jFEJhcw94_0),.din(w_dff_A_ijIOBYxc4_0),.clk(gclk));
	jdff dff_A_jFEJhcw94_0(.dout(w_dff_A_JVvijcYU1_0),.din(w_dff_A_jFEJhcw94_0),.clk(gclk));
	jdff dff_A_JVvijcYU1_0(.dout(w_dff_A_yGx7oG0K3_0),.din(w_dff_A_JVvijcYU1_0),.clk(gclk));
	jdff dff_A_yGx7oG0K3_0(.dout(w_dff_A_FHiqnv7H8_0),.din(w_dff_A_yGx7oG0K3_0),.clk(gclk));
	jdff dff_A_FHiqnv7H8_0(.dout(w_dff_A_f0gM1s5W2_0),.din(w_dff_A_FHiqnv7H8_0),.clk(gclk));
	jdff dff_A_f0gM1s5W2_0(.dout(w_dff_A_4iHu8ezz9_0),.din(w_dff_A_f0gM1s5W2_0),.clk(gclk));
	jdff dff_A_4iHu8ezz9_0(.dout(w_dff_A_mJY6w7js8_0),.din(w_dff_A_4iHu8ezz9_0),.clk(gclk));
	jdff dff_A_mJY6w7js8_0(.dout(w_dff_A_LD26rznv4_0),.din(w_dff_A_mJY6w7js8_0),.clk(gclk));
	jdff dff_A_LD26rznv4_0(.dout(w_dff_A_HNHrvkNo8_0),.din(w_dff_A_LD26rznv4_0),.clk(gclk));
	jdff dff_A_HNHrvkNo8_0(.dout(w_dff_A_Qj9BCZR75_0),.din(w_dff_A_HNHrvkNo8_0),.clk(gclk));
	jdff dff_A_Qj9BCZR75_0(.dout(w_dff_A_5czEvGOu2_0),.din(w_dff_A_Qj9BCZR75_0),.clk(gclk));
	jdff dff_A_5czEvGOu2_0(.dout(w_dff_A_nsgSRCgU3_0),.din(w_dff_A_5czEvGOu2_0),.clk(gclk));
	jdff dff_A_nsgSRCgU3_0(.dout(w_dff_A_okbHxb314_0),.din(w_dff_A_nsgSRCgU3_0),.clk(gclk));
	jdff dff_A_okbHxb314_0(.dout(w_dff_A_5ZmMUI1l1_0),.din(w_dff_A_okbHxb314_0),.clk(gclk));
	jdff dff_A_5ZmMUI1l1_0(.dout(w_dff_A_6hMGT60p9_0),.din(w_dff_A_5ZmMUI1l1_0),.clk(gclk));
	jdff dff_A_6hMGT60p9_0(.dout(w_dff_A_HuYc30OT2_0),.din(w_dff_A_6hMGT60p9_0),.clk(gclk));
	jdff dff_A_HuYc30OT2_0(.dout(w_dff_A_NbavnChT7_0),.din(w_dff_A_HuYc30OT2_0),.clk(gclk));
	jdff dff_A_NbavnChT7_0(.dout(w_dff_A_xNJ98UHb0_0),.din(w_dff_A_NbavnChT7_0),.clk(gclk));
	jdff dff_A_xNJ98UHb0_0(.dout(G526),.din(w_dff_A_xNJ98UHb0_0),.clk(gclk));
	jdff dff_A_7CNN2QGj1_1(.dout(w_dff_A_wPADSHmc3_0),.din(w_dff_A_7CNN2QGj1_1),.clk(gclk));
	jdff dff_A_wPADSHmc3_0(.dout(w_dff_A_UfqHfyUg4_0),.din(w_dff_A_wPADSHmc3_0),.clk(gclk));
	jdff dff_A_UfqHfyUg4_0(.dout(w_dff_A_XLoXWYXv6_0),.din(w_dff_A_UfqHfyUg4_0),.clk(gclk));
	jdff dff_A_XLoXWYXv6_0(.dout(w_dff_A_9CZaF95Y6_0),.din(w_dff_A_XLoXWYXv6_0),.clk(gclk));
	jdff dff_A_9CZaF95Y6_0(.dout(w_dff_A_fXX5esH14_0),.din(w_dff_A_9CZaF95Y6_0),.clk(gclk));
	jdff dff_A_fXX5esH14_0(.dout(w_dff_A_H6sED84P5_0),.din(w_dff_A_fXX5esH14_0),.clk(gclk));
	jdff dff_A_H6sED84P5_0(.dout(w_dff_A_ixSHJUKU4_0),.din(w_dff_A_H6sED84P5_0),.clk(gclk));
	jdff dff_A_ixSHJUKU4_0(.dout(w_dff_A_Ax5ViNf71_0),.din(w_dff_A_ixSHJUKU4_0),.clk(gclk));
	jdff dff_A_Ax5ViNf71_0(.dout(w_dff_A_xIk4ZfjZ1_0),.din(w_dff_A_Ax5ViNf71_0),.clk(gclk));
	jdff dff_A_xIk4ZfjZ1_0(.dout(w_dff_A_ww5h3tzY7_0),.din(w_dff_A_xIk4ZfjZ1_0),.clk(gclk));
	jdff dff_A_ww5h3tzY7_0(.dout(w_dff_A_T2WSgOqE8_0),.din(w_dff_A_ww5h3tzY7_0),.clk(gclk));
	jdff dff_A_T2WSgOqE8_0(.dout(w_dff_A_H7KwQJ684_0),.din(w_dff_A_T2WSgOqE8_0),.clk(gclk));
	jdff dff_A_H7KwQJ684_0(.dout(w_dff_A_AB3GZso39_0),.din(w_dff_A_H7KwQJ684_0),.clk(gclk));
	jdff dff_A_AB3GZso39_0(.dout(w_dff_A_tEJ9L1XR0_0),.din(w_dff_A_AB3GZso39_0),.clk(gclk));
	jdff dff_A_tEJ9L1XR0_0(.dout(w_dff_A_XObD0KSJ3_0),.din(w_dff_A_tEJ9L1XR0_0),.clk(gclk));
	jdff dff_A_XObD0KSJ3_0(.dout(w_dff_A_ftVRf9Jn2_0),.din(w_dff_A_XObD0KSJ3_0),.clk(gclk));
	jdff dff_A_ftVRf9Jn2_0(.dout(w_dff_A_VfMZnpqv9_0),.din(w_dff_A_ftVRf9Jn2_0),.clk(gclk));
	jdff dff_A_VfMZnpqv9_0(.dout(w_dff_A_CzQ4pz1a5_0),.din(w_dff_A_VfMZnpqv9_0),.clk(gclk));
	jdff dff_A_CzQ4pz1a5_0(.dout(w_dff_A_OOAtbI1m4_0),.din(w_dff_A_CzQ4pz1a5_0),.clk(gclk));
	jdff dff_A_OOAtbI1m4_0(.dout(w_dff_A_Gsx3K5yd6_0),.din(w_dff_A_OOAtbI1m4_0),.clk(gclk));
	jdff dff_A_Gsx3K5yd6_0(.dout(w_dff_A_FESGzfjc1_0),.din(w_dff_A_Gsx3K5yd6_0),.clk(gclk));
	jdff dff_A_FESGzfjc1_0(.dout(w_dff_A_4E4cdKaC4_0),.din(w_dff_A_FESGzfjc1_0),.clk(gclk));
	jdff dff_A_4E4cdKaC4_0(.dout(w_dff_A_gYgrfdEk4_0),.din(w_dff_A_4E4cdKaC4_0),.clk(gclk));
	jdff dff_A_gYgrfdEk4_0(.dout(w_dff_A_EVpZsa9A0_0),.din(w_dff_A_gYgrfdEk4_0),.clk(gclk));
	jdff dff_A_EVpZsa9A0_0(.dout(w_dff_A_kLXAngYK6_0),.din(w_dff_A_EVpZsa9A0_0),.clk(gclk));
	jdff dff_A_kLXAngYK6_0(.dout(G524),.din(w_dff_A_kLXAngYK6_0),.clk(gclk));
	jdff dff_A_rfiYBFTn8_1(.dout(w_dff_A_KBv17TNX9_0),.din(w_dff_A_rfiYBFTn8_1),.clk(gclk));
	jdff dff_A_KBv17TNX9_0(.dout(w_dff_A_eYF8b48w9_0),.din(w_dff_A_KBv17TNX9_0),.clk(gclk));
	jdff dff_A_eYF8b48w9_0(.dout(w_dff_A_Bws8PJEh4_0),.din(w_dff_A_eYF8b48w9_0),.clk(gclk));
	jdff dff_A_Bws8PJEh4_0(.dout(w_dff_A_3DAFSLe24_0),.din(w_dff_A_Bws8PJEh4_0),.clk(gclk));
	jdff dff_A_3DAFSLe24_0(.dout(w_dff_A_EqiYcGl26_0),.din(w_dff_A_3DAFSLe24_0),.clk(gclk));
	jdff dff_A_EqiYcGl26_0(.dout(w_dff_A_kvlIc9Fz3_0),.din(w_dff_A_EqiYcGl26_0),.clk(gclk));
	jdff dff_A_kvlIc9Fz3_0(.dout(w_dff_A_6Z60N6TK4_0),.din(w_dff_A_kvlIc9Fz3_0),.clk(gclk));
	jdff dff_A_6Z60N6TK4_0(.dout(w_dff_A_6FalZRrc5_0),.din(w_dff_A_6Z60N6TK4_0),.clk(gclk));
	jdff dff_A_6FalZRrc5_0(.dout(w_dff_A_v7Zzebew6_0),.din(w_dff_A_6FalZRrc5_0),.clk(gclk));
	jdff dff_A_v7Zzebew6_0(.dout(w_dff_A_lDTvXDzZ3_0),.din(w_dff_A_v7Zzebew6_0),.clk(gclk));
	jdff dff_A_lDTvXDzZ3_0(.dout(w_dff_A_8yNCk5pb1_0),.din(w_dff_A_lDTvXDzZ3_0),.clk(gclk));
	jdff dff_A_8yNCk5pb1_0(.dout(w_dff_A_HXlHmMDz8_0),.din(w_dff_A_8yNCk5pb1_0),.clk(gclk));
	jdff dff_A_HXlHmMDz8_0(.dout(w_dff_A_YAQm3VGj2_0),.din(w_dff_A_HXlHmMDz8_0),.clk(gclk));
	jdff dff_A_YAQm3VGj2_0(.dout(w_dff_A_TyTEpEEQ6_0),.din(w_dff_A_YAQm3VGj2_0),.clk(gclk));
	jdff dff_A_TyTEpEEQ6_0(.dout(w_dff_A_GnILxcXe2_0),.din(w_dff_A_TyTEpEEQ6_0),.clk(gclk));
	jdff dff_A_GnILxcXe2_0(.dout(w_dff_A_BjlgeGGf3_0),.din(w_dff_A_GnILxcXe2_0),.clk(gclk));
	jdff dff_A_BjlgeGGf3_0(.dout(w_dff_A_LWN4IjBz3_0),.din(w_dff_A_BjlgeGGf3_0),.clk(gclk));
	jdff dff_A_LWN4IjBz3_0(.dout(w_dff_A_7CQEVQDv5_0),.din(w_dff_A_LWN4IjBz3_0),.clk(gclk));
	jdff dff_A_7CQEVQDv5_0(.dout(w_dff_A_Svu2ui5v0_0),.din(w_dff_A_7CQEVQDv5_0),.clk(gclk));
	jdff dff_A_Svu2ui5v0_0(.dout(w_dff_A_5SUASKkG3_0),.din(w_dff_A_Svu2ui5v0_0),.clk(gclk));
	jdff dff_A_5SUASKkG3_0(.dout(w_dff_A_vEzzzN135_0),.din(w_dff_A_5SUASKkG3_0),.clk(gclk));
	jdff dff_A_vEzzzN135_0(.dout(w_dff_A_GvabwsAo3_0),.din(w_dff_A_vEzzzN135_0),.clk(gclk));
	jdff dff_A_GvabwsAo3_0(.dout(w_dff_A_srrWgsu77_0),.din(w_dff_A_GvabwsAo3_0),.clk(gclk));
	jdff dff_A_srrWgsu77_0(.dout(w_dff_A_o1tEZ4r95_0),.din(w_dff_A_srrWgsu77_0),.clk(gclk));
	jdff dff_A_o1tEZ4r95_0(.dout(w_dff_A_NhoOKTcF7_0),.din(w_dff_A_o1tEZ4r95_0),.clk(gclk));
	jdff dff_A_NhoOKTcF7_0(.dout(G279),.din(w_dff_A_NhoOKTcF7_0),.clk(gclk));
	jdff dff_A_vzwKrL7w6_1(.dout(w_dff_A_6JOIMAZh5_0),.din(w_dff_A_vzwKrL7w6_1),.clk(gclk));
	jdff dff_A_6JOIMAZh5_0(.dout(w_dff_A_HXCK9GeG6_0),.din(w_dff_A_6JOIMAZh5_0),.clk(gclk));
	jdff dff_A_HXCK9GeG6_0(.dout(w_dff_A_jnAEY3hC4_0),.din(w_dff_A_HXCK9GeG6_0),.clk(gclk));
	jdff dff_A_jnAEY3hC4_0(.dout(w_dff_A_5T71wfnt9_0),.din(w_dff_A_jnAEY3hC4_0),.clk(gclk));
	jdff dff_A_5T71wfnt9_0(.dout(w_dff_A_RSOKYoRU9_0),.din(w_dff_A_5T71wfnt9_0),.clk(gclk));
	jdff dff_A_RSOKYoRU9_0(.dout(w_dff_A_kMdOAi0x2_0),.din(w_dff_A_RSOKYoRU9_0),.clk(gclk));
	jdff dff_A_kMdOAi0x2_0(.dout(w_dff_A_J3I9FHX88_0),.din(w_dff_A_kMdOAi0x2_0),.clk(gclk));
	jdff dff_A_J3I9FHX88_0(.dout(w_dff_A_zerZj92j0_0),.din(w_dff_A_J3I9FHX88_0),.clk(gclk));
	jdff dff_A_zerZj92j0_0(.dout(w_dff_A_pox6fFuC4_0),.din(w_dff_A_zerZj92j0_0),.clk(gclk));
	jdff dff_A_pox6fFuC4_0(.dout(w_dff_A_Duz2K8qb1_0),.din(w_dff_A_pox6fFuC4_0),.clk(gclk));
	jdff dff_A_Duz2K8qb1_0(.dout(w_dff_A_sCyRjIMc0_0),.din(w_dff_A_Duz2K8qb1_0),.clk(gclk));
	jdff dff_A_sCyRjIMc0_0(.dout(w_dff_A_cq5ftkKE6_0),.din(w_dff_A_sCyRjIMc0_0),.clk(gclk));
	jdff dff_A_cq5ftkKE6_0(.dout(w_dff_A_YLNZXz9w3_0),.din(w_dff_A_cq5ftkKE6_0),.clk(gclk));
	jdff dff_A_YLNZXz9w3_0(.dout(w_dff_A_iEgz1ea65_0),.din(w_dff_A_YLNZXz9w3_0),.clk(gclk));
	jdff dff_A_iEgz1ea65_0(.dout(w_dff_A_cw8y85bi0_0),.din(w_dff_A_iEgz1ea65_0),.clk(gclk));
	jdff dff_A_cw8y85bi0_0(.dout(w_dff_A_Uslt2Quc2_0),.din(w_dff_A_cw8y85bi0_0),.clk(gclk));
	jdff dff_A_Uslt2Quc2_0(.dout(w_dff_A_nczOkbvE2_0),.din(w_dff_A_Uslt2Quc2_0),.clk(gclk));
	jdff dff_A_nczOkbvE2_0(.dout(w_dff_A_LMIHyfFj4_0),.din(w_dff_A_nczOkbvE2_0),.clk(gclk));
	jdff dff_A_LMIHyfFj4_0(.dout(w_dff_A_6chGvKM88_0),.din(w_dff_A_LMIHyfFj4_0),.clk(gclk));
	jdff dff_A_6chGvKM88_0(.dout(w_dff_A_bRBAi5Lb3_0),.din(w_dff_A_6chGvKM88_0),.clk(gclk));
	jdff dff_A_bRBAi5Lb3_0(.dout(w_dff_A_OW8nLXc88_0),.din(w_dff_A_bRBAi5Lb3_0),.clk(gclk));
	jdff dff_A_OW8nLXc88_0(.dout(w_dff_A_3TrrA0Ne9_0),.din(w_dff_A_OW8nLXc88_0),.clk(gclk));
	jdff dff_A_3TrrA0Ne9_0(.dout(w_dff_A_ISuiKvfN8_0),.din(w_dff_A_3TrrA0Ne9_0),.clk(gclk));
	jdff dff_A_ISuiKvfN8_0(.dout(w_dff_A_ctXFwlbt2_0),.din(w_dff_A_ISuiKvfN8_0),.clk(gclk));
	jdff dff_A_ctXFwlbt2_0(.dout(w_dff_A_7eIriKKN8_0),.din(w_dff_A_ctXFwlbt2_0),.clk(gclk));
	jdff dff_A_7eIriKKN8_0(.dout(G436),.din(w_dff_A_7eIriKKN8_0),.clk(gclk));
	jdff dff_A_FaNycJh43_1(.dout(w_dff_A_qGY3H2J69_0),.din(w_dff_A_FaNycJh43_1),.clk(gclk));
	jdff dff_A_qGY3H2J69_0(.dout(w_dff_A_lsSkBHxA3_0),.din(w_dff_A_qGY3H2J69_0),.clk(gclk));
	jdff dff_A_lsSkBHxA3_0(.dout(w_dff_A_GcliZzoZ7_0),.din(w_dff_A_lsSkBHxA3_0),.clk(gclk));
	jdff dff_A_GcliZzoZ7_0(.dout(w_dff_A_vV6ldDxr2_0),.din(w_dff_A_GcliZzoZ7_0),.clk(gclk));
	jdff dff_A_vV6ldDxr2_0(.dout(w_dff_A_YWZF2o7m3_0),.din(w_dff_A_vV6ldDxr2_0),.clk(gclk));
	jdff dff_A_YWZF2o7m3_0(.dout(w_dff_A_ySXUJJNC7_0),.din(w_dff_A_YWZF2o7m3_0),.clk(gclk));
	jdff dff_A_ySXUJJNC7_0(.dout(w_dff_A_HgFrOgpO1_0),.din(w_dff_A_ySXUJJNC7_0),.clk(gclk));
	jdff dff_A_HgFrOgpO1_0(.dout(w_dff_A_MCzTh2bB6_0),.din(w_dff_A_HgFrOgpO1_0),.clk(gclk));
	jdff dff_A_MCzTh2bB6_0(.dout(w_dff_A_KecxzNaP9_0),.din(w_dff_A_MCzTh2bB6_0),.clk(gclk));
	jdff dff_A_KecxzNaP9_0(.dout(w_dff_A_BORnleMq9_0),.din(w_dff_A_KecxzNaP9_0),.clk(gclk));
	jdff dff_A_BORnleMq9_0(.dout(w_dff_A_cssMt9s20_0),.din(w_dff_A_BORnleMq9_0),.clk(gclk));
	jdff dff_A_cssMt9s20_0(.dout(w_dff_A_ZnpVQHlJ1_0),.din(w_dff_A_cssMt9s20_0),.clk(gclk));
	jdff dff_A_ZnpVQHlJ1_0(.dout(w_dff_A_deleM0tD5_0),.din(w_dff_A_ZnpVQHlJ1_0),.clk(gclk));
	jdff dff_A_deleM0tD5_0(.dout(w_dff_A_ErLBn5y45_0),.din(w_dff_A_deleM0tD5_0),.clk(gclk));
	jdff dff_A_ErLBn5y45_0(.dout(w_dff_A_55Q1owVA1_0),.din(w_dff_A_ErLBn5y45_0),.clk(gclk));
	jdff dff_A_55Q1owVA1_0(.dout(w_dff_A_LbLt0Dhv2_0),.din(w_dff_A_55Q1owVA1_0),.clk(gclk));
	jdff dff_A_LbLt0Dhv2_0(.dout(w_dff_A_LstWs4qX6_0),.din(w_dff_A_LbLt0Dhv2_0),.clk(gclk));
	jdff dff_A_LstWs4qX6_0(.dout(w_dff_A_NACdGWnd0_0),.din(w_dff_A_LstWs4qX6_0),.clk(gclk));
	jdff dff_A_NACdGWnd0_0(.dout(w_dff_A_O7Pr7R1k4_0),.din(w_dff_A_NACdGWnd0_0),.clk(gclk));
	jdff dff_A_O7Pr7R1k4_0(.dout(w_dff_A_GjOo3sNm4_0),.din(w_dff_A_O7Pr7R1k4_0),.clk(gclk));
	jdff dff_A_GjOo3sNm4_0(.dout(w_dff_A_K2M5jAHP2_0),.din(w_dff_A_GjOo3sNm4_0),.clk(gclk));
	jdff dff_A_K2M5jAHP2_0(.dout(w_dff_A_MJuuir9n5_0),.din(w_dff_A_K2M5jAHP2_0),.clk(gclk));
	jdff dff_A_MJuuir9n5_0(.dout(w_dff_A_robZoaqS9_0),.din(w_dff_A_MJuuir9n5_0),.clk(gclk));
	jdff dff_A_robZoaqS9_0(.dout(w_dff_A_gAIBCOyk9_0),.din(w_dff_A_robZoaqS9_0),.clk(gclk));
	jdff dff_A_gAIBCOyk9_0(.dout(w_dff_A_AMKGO00a5_0),.din(w_dff_A_gAIBCOyk9_0),.clk(gclk));
	jdff dff_A_AMKGO00a5_0(.dout(G478),.din(w_dff_A_AMKGO00a5_0),.clk(gclk));
	jdff dff_A_brqg9SVn2_1(.dout(w_dff_A_i2nClWBd8_0),.din(w_dff_A_brqg9SVn2_1),.clk(gclk));
	jdff dff_A_i2nClWBd8_0(.dout(w_dff_A_rjGy2gj30_0),.din(w_dff_A_i2nClWBd8_0),.clk(gclk));
	jdff dff_A_rjGy2gj30_0(.dout(w_dff_A_8a2xj6IU7_0),.din(w_dff_A_rjGy2gj30_0),.clk(gclk));
	jdff dff_A_8a2xj6IU7_0(.dout(w_dff_A_SIGElxjj8_0),.din(w_dff_A_8a2xj6IU7_0),.clk(gclk));
	jdff dff_A_SIGElxjj8_0(.dout(w_dff_A_wJTkngWn6_0),.din(w_dff_A_SIGElxjj8_0),.clk(gclk));
	jdff dff_A_wJTkngWn6_0(.dout(w_dff_A_mLbAkSGR0_0),.din(w_dff_A_wJTkngWn6_0),.clk(gclk));
	jdff dff_A_mLbAkSGR0_0(.dout(w_dff_A_klxBYdW41_0),.din(w_dff_A_mLbAkSGR0_0),.clk(gclk));
	jdff dff_A_klxBYdW41_0(.dout(w_dff_A_Xbv4C9a58_0),.din(w_dff_A_klxBYdW41_0),.clk(gclk));
	jdff dff_A_Xbv4C9a58_0(.dout(w_dff_A_aoc4nmTr8_0),.din(w_dff_A_Xbv4C9a58_0),.clk(gclk));
	jdff dff_A_aoc4nmTr8_0(.dout(w_dff_A_ZSaE2QXU7_0),.din(w_dff_A_aoc4nmTr8_0),.clk(gclk));
	jdff dff_A_ZSaE2QXU7_0(.dout(w_dff_A_266lQG9v2_0),.din(w_dff_A_ZSaE2QXU7_0),.clk(gclk));
	jdff dff_A_266lQG9v2_0(.dout(w_dff_A_ACClf9oO2_0),.din(w_dff_A_266lQG9v2_0),.clk(gclk));
	jdff dff_A_ACClf9oO2_0(.dout(w_dff_A_xt4hKMK18_0),.din(w_dff_A_ACClf9oO2_0),.clk(gclk));
	jdff dff_A_xt4hKMK18_0(.dout(w_dff_A_8EV2gJwp6_0),.din(w_dff_A_xt4hKMK18_0),.clk(gclk));
	jdff dff_A_8EV2gJwp6_0(.dout(w_dff_A_0qYkfXI60_0),.din(w_dff_A_8EV2gJwp6_0),.clk(gclk));
	jdff dff_A_0qYkfXI60_0(.dout(w_dff_A_3JpaDPRG0_0),.din(w_dff_A_0qYkfXI60_0),.clk(gclk));
	jdff dff_A_3JpaDPRG0_0(.dout(w_dff_A_29vsu59F3_0),.din(w_dff_A_3JpaDPRG0_0),.clk(gclk));
	jdff dff_A_29vsu59F3_0(.dout(w_dff_A_9K2fRsf20_0),.din(w_dff_A_29vsu59F3_0),.clk(gclk));
	jdff dff_A_9K2fRsf20_0(.dout(w_dff_A_wexf8Kp48_0),.din(w_dff_A_9K2fRsf20_0),.clk(gclk));
	jdff dff_A_wexf8Kp48_0(.dout(w_dff_A_MOslUsCL4_0),.din(w_dff_A_wexf8Kp48_0),.clk(gclk));
	jdff dff_A_MOslUsCL4_0(.dout(w_dff_A_wtQqCkoa2_0),.din(w_dff_A_MOslUsCL4_0),.clk(gclk));
	jdff dff_A_wtQqCkoa2_0(.dout(w_dff_A_JpM7Yh8f2_0),.din(w_dff_A_wtQqCkoa2_0),.clk(gclk));
	jdff dff_A_JpM7Yh8f2_0(.dout(w_dff_A_WozjK2822_0),.din(w_dff_A_JpM7Yh8f2_0),.clk(gclk));
	jdff dff_A_WozjK2822_0(.dout(w_dff_A_oR7RuUwk7_0),.din(w_dff_A_WozjK2822_0),.clk(gclk));
	jdff dff_A_oR7RuUwk7_0(.dout(w_dff_A_UJXTa3yz1_0),.din(w_dff_A_oR7RuUwk7_0),.clk(gclk));
	jdff dff_A_UJXTa3yz1_0(.dout(G522),.din(w_dff_A_UJXTa3yz1_0),.clk(gclk));
	jdff dff_A_ZwI2TXIA4_2(.dout(w_dff_A_sYOBUnNc1_0),.din(w_dff_A_ZwI2TXIA4_2),.clk(gclk));
	jdff dff_A_sYOBUnNc1_0(.dout(w_dff_A_SWDkKvin7_0),.din(w_dff_A_sYOBUnNc1_0),.clk(gclk));
	jdff dff_A_SWDkKvin7_0(.dout(w_dff_A_JjIlIpCG1_0),.din(w_dff_A_SWDkKvin7_0),.clk(gclk));
	jdff dff_A_JjIlIpCG1_0(.dout(w_dff_A_ABN2chsT9_0),.din(w_dff_A_JjIlIpCG1_0),.clk(gclk));
	jdff dff_A_ABN2chsT9_0(.dout(w_dff_A_Btkxkv7A9_0),.din(w_dff_A_ABN2chsT9_0),.clk(gclk));
	jdff dff_A_Btkxkv7A9_0(.dout(w_dff_A_cwgUJgkC7_0),.din(w_dff_A_Btkxkv7A9_0),.clk(gclk));
	jdff dff_A_cwgUJgkC7_0(.dout(w_dff_A_vipA9yt70_0),.din(w_dff_A_cwgUJgkC7_0),.clk(gclk));
	jdff dff_A_vipA9yt70_0(.dout(w_dff_A_OdKV93LJ2_0),.din(w_dff_A_vipA9yt70_0),.clk(gclk));
	jdff dff_A_OdKV93LJ2_0(.dout(w_dff_A_kSn5jDc07_0),.din(w_dff_A_OdKV93LJ2_0),.clk(gclk));
	jdff dff_A_kSn5jDc07_0(.dout(w_dff_A_KNQPhlBV5_0),.din(w_dff_A_kSn5jDc07_0),.clk(gclk));
	jdff dff_A_KNQPhlBV5_0(.dout(w_dff_A_ZrlN9XDj7_0),.din(w_dff_A_KNQPhlBV5_0),.clk(gclk));
	jdff dff_A_ZrlN9XDj7_0(.dout(w_dff_A_qHJFyHS24_0),.din(w_dff_A_ZrlN9XDj7_0),.clk(gclk));
	jdff dff_A_qHJFyHS24_0(.dout(w_dff_A_8CNmKfhf2_0),.din(w_dff_A_qHJFyHS24_0),.clk(gclk));
	jdff dff_A_8CNmKfhf2_0(.dout(w_dff_A_zWxyZbO43_0),.din(w_dff_A_8CNmKfhf2_0),.clk(gclk));
	jdff dff_A_zWxyZbO43_0(.dout(w_dff_A_2c8CazQk6_0),.din(w_dff_A_zWxyZbO43_0),.clk(gclk));
	jdff dff_A_2c8CazQk6_0(.dout(w_dff_A_3Ah7ubNf7_0),.din(w_dff_A_2c8CazQk6_0),.clk(gclk));
	jdff dff_A_3Ah7ubNf7_0(.dout(w_dff_A_m0PycPBr2_0),.din(w_dff_A_3Ah7ubNf7_0),.clk(gclk));
	jdff dff_A_m0PycPBr2_0(.dout(w_dff_A_3errfxBV5_0),.din(w_dff_A_m0PycPBr2_0),.clk(gclk));
	jdff dff_A_3errfxBV5_0(.dout(w_dff_A_4lcwrkSK1_0),.din(w_dff_A_3errfxBV5_0),.clk(gclk));
	jdff dff_A_4lcwrkSK1_0(.dout(w_dff_A_O2j4AT3g2_0),.din(w_dff_A_4lcwrkSK1_0),.clk(gclk));
	jdff dff_A_O2j4AT3g2_0(.dout(w_dff_A_Apx7J8mW7_0),.din(w_dff_A_O2j4AT3g2_0),.clk(gclk));
	jdff dff_A_Apx7J8mW7_0(.dout(w_dff_A_e7RAeC0K0_0),.din(w_dff_A_Apx7J8mW7_0),.clk(gclk));
	jdff dff_A_e7RAeC0K0_0(.dout(w_dff_A_QjToOTvY1_0),.din(w_dff_A_e7RAeC0K0_0),.clk(gclk));
	jdff dff_A_QjToOTvY1_0(.dout(w_dff_A_tVxoQLMN0_0),.din(w_dff_A_QjToOTvY1_0),.clk(gclk));
	jdff dff_A_tVxoQLMN0_0(.dout(w_dff_A_7lcWiGlO9_0),.din(w_dff_A_tVxoQLMN0_0),.clk(gclk));
	jdff dff_A_7lcWiGlO9_0(.dout(G402),.din(w_dff_A_7lcWiGlO9_0),.clk(gclk));
	jdff dff_A_amYEkAj00_1(.dout(w_dff_A_LaqWwdLI9_0),.din(w_dff_A_amYEkAj00_1),.clk(gclk));
	jdff dff_A_LaqWwdLI9_0(.dout(w_dff_A_AKECcuck3_0),.din(w_dff_A_LaqWwdLI9_0),.clk(gclk));
	jdff dff_A_AKECcuck3_0(.dout(w_dff_A_RpsUUWyQ1_0),.din(w_dff_A_AKECcuck3_0),.clk(gclk));
	jdff dff_A_RpsUUWyQ1_0(.dout(w_dff_A_eROdEdx10_0),.din(w_dff_A_RpsUUWyQ1_0),.clk(gclk));
	jdff dff_A_eROdEdx10_0(.dout(w_dff_A_4DHT6LpY4_0),.din(w_dff_A_eROdEdx10_0),.clk(gclk));
	jdff dff_A_4DHT6LpY4_0(.dout(w_dff_A_5mDj9NIa8_0),.din(w_dff_A_4DHT6LpY4_0),.clk(gclk));
	jdff dff_A_5mDj9NIa8_0(.dout(w_dff_A_bw0vr69i8_0),.din(w_dff_A_5mDj9NIa8_0),.clk(gclk));
	jdff dff_A_bw0vr69i8_0(.dout(w_dff_A_dLmmBDjx3_0),.din(w_dff_A_bw0vr69i8_0),.clk(gclk));
	jdff dff_A_dLmmBDjx3_0(.dout(w_dff_A_vPFBJJbJ9_0),.din(w_dff_A_dLmmBDjx3_0),.clk(gclk));
	jdff dff_A_vPFBJJbJ9_0(.dout(w_dff_A_Twal4M3a4_0),.din(w_dff_A_vPFBJJbJ9_0),.clk(gclk));
	jdff dff_A_Twal4M3a4_0(.dout(w_dff_A_oqWc8lh36_0),.din(w_dff_A_Twal4M3a4_0),.clk(gclk));
	jdff dff_A_oqWc8lh36_0(.dout(w_dff_A_U6HvmVBJ8_0),.din(w_dff_A_oqWc8lh36_0),.clk(gclk));
	jdff dff_A_U6HvmVBJ8_0(.dout(w_dff_A_aoOGWk9v8_0),.din(w_dff_A_U6HvmVBJ8_0),.clk(gclk));
	jdff dff_A_aoOGWk9v8_0(.dout(w_dff_A_1Jo9rpXr5_0),.din(w_dff_A_aoOGWk9v8_0),.clk(gclk));
	jdff dff_A_1Jo9rpXr5_0(.dout(w_dff_A_xQ9nMkpX1_0),.din(w_dff_A_1Jo9rpXr5_0),.clk(gclk));
	jdff dff_A_xQ9nMkpX1_0(.dout(w_dff_A_5SbnuXRR1_0),.din(w_dff_A_xQ9nMkpX1_0),.clk(gclk));
	jdff dff_A_5SbnuXRR1_0(.dout(w_dff_A_w3mJGjV52_0),.din(w_dff_A_5SbnuXRR1_0),.clk(gclk));
	jdff dff_A_w3mJGjV52_0(.dout(w_dff_A_7gPHDzAO7_0),.din(w_dff_A_w3mJGjV52_0),.clk(gclk));
	jdff dff_A_7gPHDzAO7_0(.dout(w_dff_A_fUfY2IBG8_0),.din(w_dff_A_7gPHDzAO7_0),.clk(gclk));
	jdff dff_A_fUfY2IBG8_0(.dout(w_dff_A_WkWstzRA6_0),.din(w_dff_A_fUfY2IBG8_0),.clk(gclk));
	jdff dff_A_WkWstzRA6_0(.dout(w_dff_A_8QG85tXQ5_0),.din(w_dff_A_WkWstzRA6_0),.clk(gclk));
	jdff dff_A_8QG85tXQ5_0(.dout(w_dff_A_rPwfwKyQ7_0),.din(w_dff_A_8QG85tXQ5_0),.clk(gclk));
	jdff dff_A_rPwfwKyQ7_0(.dout(w_dff_A_GnEmrQDq6_0),.din(w_dff_A_rPwfwKyQ7_0),.clk(gclk));
	jdff dff_A_GnEmrQDq6_0(.dout(G404),.din(w_dff_A_GnEmrQDq6_0),.clk(gclk));
	jdff dff_A_t6zLtL210_1(.dout(w_dff_A_0GahgdHp1_0),.din(w_dff_A_t6zLtL210_1),.clk(gclk));
	jdff dff_A_0GahgdHp1_0(.dout(w_dff_A_jMA16JGn6_0),.din(w_dff_A_0GahgdHp1_0),.clk(gclk));
	jdff dff_A_jMA16JGn6_0(.dout(w_dff_A_TDTUcUn22_0),.din(w_dff_A_jMA16JGn6_0),.clk(gclk));
	jdff dff_A_TDTUcUn22_0(.dout(w_dff_A_jWjxuwBj5_0),.din(w_dff_A_TDTUcUn22_0),.clk(gclk));
	jdff dff_A_jWjxuwBj5_0(.dout(w_dff_A_lkwW53Hb9_0),.din(w_dff_A_jWjxuwBj5_0),.clk(gclk));
	jdff dff_A_lkwW53Hb9_0(.dout(w_dff_A_WpFj8LLB2_0),.din(w_dff_A_lkwW53Hb9_0),.clk(gclk));
	jdff dff_A_WpFj8LLB2_0(.dout(w_dff_A_aolWF1GW7_0),.din(w_dff_A_WpFj8LLB2_0),.clk(gclk));
	jdff dff_A_aolWF1GW7_0(.dout(w_dff_A_GWLXQRzp2_0),.din(w_dff_A_aolWF1GW7_0),.clk(gclk));
	jdff dff_A_GWLXQRzp2_0(.dout(w_dff_A_qO5YtnWr3_0),.din(w_dff_A_GWLXQRzp2_0),.clk(gclk));
	jdff dff_A_qO5YtnWr3_0(.dout(w_dff_A_BSs8seSw3_0),.din(w_dff_A_qO5YtnWr3_0),.clk(gclk));
	jdff dff_A_BSs8seSw3_0(.dout(w_dff_A_OWT6ucqT4_0),.din(w_dff_A_BSs8seSw3_0),.clk(gclk));
	jdff dff_A_OWT6ucqT4_0(.dout(w_dff_A_z4W6vr4U3_0),.din(w_dff_A_OWT6ucqT4_0),.clk(gclk));
	jdff dff_A_z4W6vr4U3_0(.dout(w_dff_A_E9n4eXgP9_0),.din(w_dff_A_z4W6vr4U3_0),.clk(gclk));
	jdff dff_A_E9n4eXgP9_0(.dout(w_dff_A_w3jBFa2V8_0),.din(w_dff_A_E9n4eXgP9_0),.clk(gclk));
	jdff dff_A_w3jBFa2V8_0(.dout(w_dff_A_OYdpdVrd2_0),.din(w_dff_A_w3jBFa2V8_0),.clk(gclk));
	jdff dff_A_OYdpdVrd2_0(.dout(w_dff_A_7wJGjD7S5_0),.din(w_dff_A_OYdpdVrd2_0),.clk(gclk));
	jdff dff_A_7wJGjD7S5_0(.dout(w_dff_A_8KaPnuhh1_0),.din(w_dff_A_7wJGjD7S5_0),.clk(gclk));
	jdff dff_A_8KaPnuhh1_0(.dout(w_dff_A_eIuhuls23_0),.din(w_dff_A_8KaPnuhh1_0),.clk(gclk));
	jdff dff_A_eIuhuls23_0(.dout(w_dff_A_4UfwIdWz5_0),.din(w_dff_A_eIuhuls23_0),.clk(gclk));
	jdff dff_A_4UfwIdWz5_0(.dout(w_dff_A_6pgKHLx60_0),.din(w_dff_A_4UfwIdWz5_0),.clk(gclk));
	jdff dff_A_6pgKHLx60_0(.dout(w_dff_A_uyafAuev0_0),.din(w_dff_A_6pgKHLx60_0),.clk(gclk));
	jdff dff_A_uyafAuev0_0(.dout(w_dff_A_ZvUt2NIY0_0),.din(w_dff_A_uyafAuev0_0),.clk(gclk));
	jdff dff_A_ZvUt2NIY0_0(.dout(w_dff_A_Chpxamw89_0),.din(w_dff_A_ZvUt2NIY0_0),.clk(gclk));
	jdff dff_A_Chpxamw89_0(.dout(G406),.din(w_dff_A_Chpxamw89_0),.clk(gclk));
	jdff dff_A_08FIgT3x3_1(.dout(w_dff_A_DEWlQHHu2_0),.din(w_dff_A_08FIgT3x3_1),.clk(gclk));
	jdff dff_A_DEWlQHHu2_0(.dout(w_dff_A_NMtfxNaz9_0),.din(w_dff_A_DEWlQHHu2_0),.clk(gclk));
	jdff dff_A_NMtfxNaz9_0(.dout(w_dff_A_QEoySopq9_0),.din(w_dff_A_NMtfxNaz9_0),.clk(gclk));
	jdff dff_A_QEoySopq9_0(.dout(w_dff_A_8Q0uVE093_0),.din(w_dff_A_QEoySopq9_0),.clk(gclk));
	jdff dff_A_8Q0uVE093_0(.dout(w_dff_A_ZFv72X4T8_0),.din(w_dff_A_8Q0uVE093_0),.clk(gclk));
	jdff dff_A_ZFv72X4T8_0(.dout(w_dff_A_CXac6MEm2_0),.din(w_dff_A_ZFv72X4T8_0),.clk(gclk));
	jdff dff_A_CXac6MEm2_0(.dout(w_dff_A_DMK9C7R25_0),.din(w_dff_A_CXac6MEm2_0),.clk(gclk));
	jdff dff_A_DMK9C7R25_0(.dout(w_dff_A_LQkf1OU52_0),.din(w_dff_A_DMK9C7R25_0),.clk(gclk));
	jdff dff_A_LQkf1OU52_0(.dout(w_dff_A_1GojHfPY9_0),.din(w_dff_A_LQkf1OU52_0),.clk(gclk));
	jdff dff_A_1GojHfPY9_0(.dout(w_dff_A_qRdmqRbv7_0),.din(w_dff_A_1GojHfPY9_0),.clk(gclk));
	jdff dff_A_qRdmqRbv7_0(.dout(w_dff_A_K6kgOyaC8_0),.din(w_dff_A_qRdmqRbv7_0),.clk(gclk));
	jdff dff_A_K6kgOyaC8_0(.dout(w_dff_A_z9ssNojK7_0),.din(w_dff_A_K6kgOyaC8_0),.clk(gclk));
	jdff dff_A_z9ssNojK7_0(.dout(w_dff_A_D9iUZg1s9_0),.din(w_dff_A_z9ssNojK7_0),.clk(gclk));
	jdff dff_A_D9iUZg1s9_0(.dout(w_dff_A_d5h4aF7y9_0),.din(w_dff_A_D9iUZg1s9_0),.clk(gclk));
	jdff dff_A_d5h4aF7y9_0(.dout(w_dff_A_p4SBo7ed9_0),.din(w_dff_A_d5h4aF7y9_0),.clk(gclk));
	jdff dff_A_p4SBo7ed9_0(.dout(w_dff_A_OUFQjWLF5_0),.din(w_dff_A_p4SBo7ed9_0),.clk(gclk));
	jdff dff_A_OUFQjWLF5_0(.dout(w_dff_A_GKB4SBDy1_0),.din(w_dff_A_OUFQjWLF5_0),.clk(gclk));
	jdff dff_A_GKB4SBDy1_0(.dout(w_dff_A_pBwVRTGm3_0),.din(w_dff_A_GKB4SBDy1_0),.clk(gclk));
	jdff dff_A_pBwVRTGm3_0(.dout(w_dff_A_Y2ftOXnw3_0),.din(w_dff_A_pBwVRTGm3_0),.clk(gclk));
	jdff dff_A_Y2ftOXnw3_0(.dout(w_dff_A_rycyxBW90_0),.din(w_dff_A_Y2ftOXnw3_0),.clk(gclk));
	jdff dff_A_rycyxBW90_0(.dout(w_dff_A_6Hi7eGz54_0),.din(w_dff_A_rycyxBW90_0),.clk(gclk));
	jdff dff_A_6Hi7eGz54_0(.dout(w_dff_A_cm03bSxK5_0),.din(w_dff_A_6Hi7eGz54_0),.clk(gclk));
	jdff dff_A_cm03bSxK5_0(.dout(w_dff_A_HanoiqVF5_0),.din(w_dff_A_cm03bSxK5_0),.clk(gclk));
	jdff dff_A_HanoiqVF5_0(.dout(G408),.din(w_dff_A_HanoiqVF5_0),.clk(gclk));
	jdff dff_A_OYPAWhe44_1(.dout(w_dff_A_Dp7qLDe60_0),.din(w_dff_A_OYPAWhe44_1),.clk(gclk));
	jdff dff_A_Dp7qLDe60_0(.dout(w_dff_A_RQOGItHR2_0),.din(w_dff_A_Dp7qLDe60_0),.clk(gclk));
	jdff dff_A_RQOGItHR2_0(.dout(w_dff_A_qsVKNdr56_0),.din(w_dff_A_RQOGItHR2_0),.clk(gclk));
	jdff dff_A_qsVKNdr56_0(.dout(w_dff_A_1VrXme1e0_0),.din(w_dff_A_qsVKNdr56_0),.clk(gclk));
	jdff dff_A_1VrXme1e0_0(.dout(w_dff_A_Z7DtqWKy9_0),.din(w_dff_A_1VrXme1e0_0),.clk(gclk));
	jdff dff_A_Z7DtqWKy9_0(.dout(w_dff_A_AyOK5qy39_0),.din(w_dff_A_Z7DtqWKy9_0),.clk(gclk));
	jdff dff_A_AyOK5qy39_0(.dout(w_dff_A_XHSITl1N6_0),.din(w_dff_A_AyOK5qy39_0),.clk(gclk));
	jdff dff_A_XHSITl1N6_0(.dout(w_dff_A_25gz9LWm6_0),.din(w_dff_A_XHSITl1N6_0),.clk(gclk));
	jdff dff_A_25gz9LWm6_0(.dout(w_dff_A_tMyhFtJO9_0),.din(w_dff_A_25gz9LWm6_0),.clk(gclk));
	jdff dff_A_tMyhFtJO9_0(.dout(w_dff_A_CxaKyIIo8_0),.din(w_dff_A_tMyhFtJO9_0),.clk(gclk));
	jdff dff_A_CxaKyIIo8_0(.dout(w_dff_A_CnP9KI3A0_0),.din(w_dff_A_CxaKyIIo8_0),.clk(gclk));
	jdff dff_A_CnP9KI3A0_0(.dout(w_dff_A_zsbHjANn7_0),.din(w_dff_A_CnP9KI3A0_0),.clk(gclk));
	jdff dff_A_zsbHjANn7_0(.dout(w_dff_A_8CoC8X014_0),.din(w_dff_A_zsbHjANn7_0),.clk(gclk));
	jdff dff_A_8CoC8X014_0(.dout(w_dff_A_XhWbLnqH2_0),.din(w_dff_A_8CoC8X014_0),.clk(gclk));
	jdff dff_A_XhWbLnqH2_0(.dout(w_dff_A_T0i8zvlZ5_0),.din(w_dff_A_XhWbLnqH2_0),.clk(gclk));
	jdff dff_A_T0i8zvlZ5_0(.dout(w_dff_A_Gqjgf0B03_0),.din(w_dff_A_T0i8zvlZ5_0),.clk(gclk));
	jdff dff_A_Gqjgf0B03_0(.dout(w_dff_A_vMeWpli98_0),.din(w_dff_A_Gqjgf0B03_0),.clk(gclk));
	jdff dff_A_vMeWpli98_0(.dout(w_dff_A_Uz9TNndU9_0),.din(w_dff_A_vMeWpli98_0),.clk(gclk));
	jdff dff_A_Uz9TNndU9_0(.dout(w_dff_A_XvS0LSSn0_0),.din(w_dff_A_Uz9TNndU9_0),.clk(gclk));
	jdff dff_A_XvS0LSSn0_0(.dout(w_dff_A_PPBrGKr10_0),.din(w_dff_A_XvS0LSSn0_0),.clk(gclk));
	jdff dff_A_PPBrGKr10_0(.dout(w_dff_A_rM2fcNiD2_0),.din(w_dff_A_PPBrGKr10_0),.clk(gclk));
	jdff dff_A_rM2fcNiD2_0(.dout(w_dff_A_OP2oINcU6_0),.din(w_dff_A_rM2fcNiD2_0),.clk(gclk));
	jdff dff_A_OP2oINcU6_0(.dout(w_dff_A_0x6LqtEa7_0),.din(w_dff_A_OP2oINcU6_0),.clk(gclk));
	jdff dff_A_0x6LqtEa7_0(.dout(G410),.din(w_dff_A_0x6LqtEa7_0),.clk(gclk));
	jdff dff_A_72jiinuu9_1(.dout(w_dff_A_9EfaEjWq2_0),.din(w_dff_A_72jiinuu9_1),.clk(gclk));
	jdff dff_A_9EfaEjWq2_0(.dout(w_dff_A_JJ9ymX5w3_0),.din(w_dff_A_9EfaEjWq2_0),.clk(gclk));
	jdff dff_A_JJ9ymX5w3_0(.dout(w_dff_A_oIQSNchm2_0),.din(w_dff_A_JJ9ymX5w3_0),.clk(gclk));
	jdff dff_A_oIQSNchm2_0(.dout(w_dff_A_6GloHEU80_0),.din(w_dff_A_oIQSNchm2_0),.clk(gclk));
	jdff dff_A_6GloHEU80_0(.dout(w_dff_A_dKoQ4bme0_0),.din(w_dff_A_6GloHEU80_0),.clk(gclk));
	jdff dff_A_dKoQ4bme0_0(.dout(w_dff_A_foZ7Xmps6_0),.din(w_dff_A_dKoQ4bme0_0),.clk(gclk));
	jdff dff_A_foZ7Xmps6_0(.dout(w_dff_A_hs7SzKHx5_0),.din(w_dff_A_foZ7Xmps6_0),.clk(gclk));
	jdff dff_A_hs7SzKHx5_0(.dout(w_dff_A_aABwAC8k3_0),.din(w_dff_A_hs7SzKHx5_0),.clk(gclk));
	jdff dff_A_aABwAC8k3_0(.dout(w_dff_A_987uaKlJ6_0),.din(w_dff_A_aABwAC8k3_0),.clk(gclk));
	jdff dff_A_987uaKlJ6_0(.dout(w_dff_A_RIApDNOh1_0),.din(w_dff_A_987uaKlJ6_0),.clk(gclk));
	jdff dff_A_RIApDNOh1_0(.dout(w_dff_A_fFDtMKm58_0),.din(w_dff_A_RIApDNOh1_0),.clk(gclk));
	jdff dff_A_fFDtMKm58_0(.dout(w_dff_A_zvFqjdZP1_0),.din(w_dff_A_fFDtMKm58_0),.clk(gclk));
	jdff dff_A_zvFqjdZP1_0(.dout(w_dff_A_F14rt1un7_0),.din(w_dff_A_zvFqjdZP1_0),.clk(gclk));
	jdff dff_A_F14rt1un7_0(.dout(w_dff_A_1fxqwxrk0_0),.din(w_dff_A_F14rt1un7_0),.clk(gclk));
	jdff dff_A_1fxqwxrk0_0(.dout(w_dff_A_rqv531aD1_0),.din(w_dff_A_1fxqwxrk0_0),.clk(gclk));
	jdff dff_A_rqv531aD1_0(.dout(w_dff_A_M9RJhOXS1_0),.din(w_dff_A_rqv531aD1_0),.clk(gclk));
	jdff dff_A_M9RJhOXS1_0(.dout(w_dff_A_s7dAlhV41_0),.din(w_dff_A_M9RJhOXS1_0),.clk(gclk));
	jdff dff_A_s7dAlhV41_0(.dout(w_dff_A_bZDnzNKi7_0),.din(w_dff_A_s7dAlhV41_0),.clk(gclk));
	jdff dff_A_bZDnzNKi7_0(.dout(w_dff_A_pPf9xNxG2_0),.din(w_dff_A_bZDnzNKi7_0),.clk(gclk));
	jdff dff_A_pPf9xNxG2_0(.dout(w_dff_A_YO1pMBP66_0),.din(w_dff_A_pPf9xNxG2_0),.clk(gclk));
	jdff dff_A_YO1pMBP66_0(.dout(w_dff_A_7F4X4YAc1_0),.din(w_dff_A_YO1pMBP66_0),.clk(gclk));
	jdff dff_A_7F4X4YAc1_0(.dout(w_dff_A_PoAmZBwf0_0),.din(w_dff_A_7F4X4YAc1_0),.clk(gclk));
	jdff dff_A_PoAmZBwf0_0(.dout(w_dff_A_bFsmNfY29_0),.din(w_dff_A_PoAmZBwf0_0),.clk(gclk));
	jdff dff_A_bFsmNfY29_0(.dout(w_dff_A_bLpXWvvb6_0),.din(w_dff_A_bFsmNfY29_0),.clk(gclk));
	jdff dff_A_bLpXWvvb6_0(.dout(w_dff_A_OvPuv0aa0_0),.din(w_dff_A_bLpXWvvb6_0),.clk(gclk));
	jdff dff_A_OvPuv0aa0_0(.dout(G432),.din(w_dff_A_OvPuv0aa0_0),.clk(gclk));
	jdff dff_A_VcYMcl4d4_1(.dout(w_dff_A_Yf6Mekoh8_0),.din(w_dff_A_VcYMcl4d4_1),.clk(gclk));
	jdff dff_A_Yf6Mekoh8_0(.dout(w_dff_A_Yzq3GCri5_0),.din(w_dff_A_Yf6Mekoh8_0),.clk(gclk));
	jdff dff_A_Yzq3GCri5_0(.dout(w_dff_A_FzC9c08i2_0),.din(w_dff_A_Yzq3GCri5_0),.clk(gclk));
	jdff dff_A_FzC9c08i2_0(.dout(w_dff_A_BLjghiPx3_0),.din(w_dff_A_FzC9c08i2_0),.clk(gclk));
	jdff dff_A_BLjghiPx3_0(.dout(w_dff_A_D2MU0aDz7_0),.din(w_dff_A_BLjghiPx3_0),.clk(gclk));
	jdff dff_A_D2MU0aDz7_0(.dout(w_dff_A_mPT6bhaT9_0),.din(w_dff_A_D2MU0aDz7_0),.clk(gclk));
	jdff dff_A_mPT6bhaT9_0(.dout(w_dff_A_yB4gbMmo9_0),.din(w_dff_A_mPT6bhaT9_0),.clk(gclk));
	jdff dff_A_yB4gbMmo9_0(.dout(w_dff_A_tF0P8ENf7_0),.din(w_dff_A_yB4gbMmo9_0),.clk(gclk));
	jdff dff_A_tF0P8ENf7_0(.dout(w_dff_A_jVbVynpX2_0),.din(w_dff_A_tF0P8ENf7_0),.clk(gclk));
	jdff dff_A_jVbVynpX2_0(.dout(w_dff_A_sR8KRVtc9_0),.din(w_dff_A_jVbVynpX2_0),.clk(gclk));
	jdff dff_A_sR8KRVtc9_0(.dout(w_dff_A_zYfAKsO99_0),.din(w_dff_A_sR8KRVtc9_0),.clk(gclk));
	jdff dff_A_zYfAKsO99_0(.dout(w_dff_A_InB5Ribs0_0),.din(w_dff_A_zYfAKsO99_0),.clk(gclk));
	jdff dff_A_InB5Ribs0_0(.dout(w_dff_A_0lDEJ6Vf9_0),.din(w_dff_A_InB5Ribs0_0),.clk(gclk));
	jdff dff_A_0lDEJ6Vf9_0(.dout(w_dff_A_uqtJAVxu4_0),.din(w_dff_A_0lDEJ6Vf9_0),.clk(gclk));
	jdff dff_A_uqtJAVxu4_0(.dout(w_dff_A_lackjnTj4_0),.din(w_dff_A_uqtJAVxu4_0),.clk(gclk));
	jdff dff_A_lackjnTj4_0(.dout(w_dff_A_C3Wea6Qn8_0),.din(w_dff_A_lackjnTj4_0),.clk(gclk));
	jdff dff_A_C3Wea6Qn8_0(.dout(w_dff_A_INP3Vl365_0),.din(w_dff_A_C3Wea6Qn8_0),.clk(gclk));
	jdff dff_A_INP3Vl365_0(.dout(w_dff_A_2h5znEYC7_0),.din(w_dff_A_INP3Vl365_0),.clk(gclk));
	jdff dff_A_2h5znEYC7_0(.dout(w_dff_A_pDkLOFAW9_0),.din(w_dff_A_2h5znEYC7_0),.clk(gclk));
	jdff dff_A_pDkLOFAW9_0(.dout(w_dff_A_Xovkznt48_0),.din(w_dff_A_pDkLOFAW9_0),.clk(gclk));
	jdff dff_A_Xovkznt48_0(.dout(w_dff_A_rR1PNAVS2_0),.din(w_dff_A_Xovkznt48_0),.clk(gclk));
	jdff dff_A_rR1PNAVS2_0(.dout(w_dff_A_KqK4n9an8_0),.din(w_dff_A_rR1PNAVS2_0),.clk(gclk));
	jdff dff_A_KqK4n9an8_0(.dout(w_dff_A_zWXHBiP27_0),.din(w_dff_A_KqK4n9an8_0),.clk(gclk));
	jdff dff_A_zWXHBiP27_0(.dout(w_dff_A_BiNXUr146_0),.din(w_dff_A_zWXHBiP27_0),.clk(gclk));
	jdff dff_A_BiNXUr146_0(.dout(w_dff_A_nbWEwK1h1_0),.din(w_dff_A_BiNXUr146_0),.clk(gclk));
	jdff dff_A_nbWEwK1h1_0(.dout(G446),.din(w_dff_A_nbWEwK1h1_0),.clk(gclk));
	jdff dff_A_g7IbVewx2_2(.dout(w_dff_A_5wY67q0c8_0),.din(w_dff_A_g7IbVewx2_2),.clk(gclk));
	jdff dff_A_5wY67q0c8_0(.dout(w_dff_A_pwJQ3Uk11_0),.din(w_dff_A_5wY67q0c8_0),.clk(gclk));
	jdff dff_A_pwJQ3Uk11_0(.dout(w_dff_A_2KxLRPgB1_0),.din(w_dff_A_pwJQ3Uk11_0),.clk(gclk));
	jdff dff_A_2KxLRPgB1_0(.dout(w_dff_A_c9WI7ptW7_0),.din(w_dff_A_2KxLRPgB1_0),.clk(gclk));
	jdff dff_A_c9WI7ptW7_0(.dout(w_dff_A_l6Mr2j9G6_0),.din(w_dff_A_c9WI7ptW7_0),.clk(gclk));
	jdff dff_A_l6Mr2j9G6_0(.dout(w_dff_A_gg64z5bj4_0),.din(w_dff_A_l6Mr2j9G6_0),.clk(gclk));
	jdff dff_A_gg64z5bj4_0(.dout(w_dff_A_08gqP7Sd4_0),.din(w_dff_A_gg64z5bj4_0),.clk(gclk));
	jdff dff_A_08gqP7Sd4_0(.dout(w_dff_A_BkYoCBqS3_0),.din(w_dff_A_08gqP7Sd4_0),.clk(gclk));
	jdff dff_A_BkYoCBqS3_0(.dout(w_dff_A_4GXBB69u9_0),.din(w_dff_A_BkYoCBqS3_0),.clk(gclk));
	jdff dff_A_4GXBB69u9_0(.dout(w_dff_A_gMYI0Bi43_0),.din(w_dff_A_4GXBB69u9_0),.clk(gclk));
	jdff dff_A_gMYI0Bi43_0(.dout(w_dff_A_nZpA95Uc8_0),.din(w_dff_A_gMYI0Bi43_0),.clk(gclk));
	jdff dff_A_nZpA95Uc8_0(.dout(w_dff_A_xcBzd2uN8_0),.din(w_dff_A_nZpA95Uc8_0),.clk(gclk));
	jdff dff_A_xcBzd2uN8_0(.dout(w_dff_A_ZDQDla7X1_0),.din(w_dff_A_xcBzd2uN8_0),.clk(gclk));
	jdff dff_A_ZDQDla7X1_0(.dout(w_dff_A_JaYtXLZq9_0),.din(w_dff_A_ZDQDla7X1_0),.clk(gclk));
	jdff dff_A_JaYtXLZq9_0(.dout(w_dff_A_ehqFbnaG5_0),.din(w_dff_A_JaYtXLZq9_0),.clk(gclk));
	jdff dff_A_ehqFbnaG5_0(.dout(w_dff_A_B6PFfiDO5_0),.din(w_dff_A_ehqFbnaG5_0),.clk(gclk));
	jdff dff_A_B6PFfiDO5_0(.dout(w_dff_A_bt8591e34_0),.din(w_dff_A_B6PFfiDO5_0),.clk(gclk));
	jdff dff_A_bt8591e34_0(.dout(w_dff_A_wtQeivoA9_0),.din(w_dff_A_bt8591e34_0),.clk(gclk));
	jdff dff_A_wtQeivoA9_0(.dout(w_dff_A_jQaCBwwH6_0),.din(w_dff_A_wtQeivoA9_0),.clk(gclk));
	jdff dff_A_jQaCBwwH6_0(.dout(w_dff_A_JZoykD9o0_0),.din(w_dff_A_jQaCBwwH6_0),.clk(gclk));
	jdff dff_A_JZoykD9o0_0(.dout(w_dff_A_HEctrAiX7_0),.din(w_dff_A_JZoykD9o0_0),.clk(gclk));
	jdff dff_A_HEctrAiX7_0(.dout(w_dff_A_8ky1ZFCm5_0),.din(w_dff_A_HEctrAiX7_0),.clk(gclk));
	jdff dff_A_8ky1ZFCm5_0(.dout(w_dff_A_N445o3Rm9_0),.din(w_dff_A_8ky1ZFCm5_0),.clk(gclk));
	jdff dff_A_N445o3Rm9_0(.dout(w_dff_A_X9VjWtUB8_0),.din(w_dff_A_N445o3Rm9_0),.clk(gclk));
	jdff dff_A_X9VjWtUB8_0(.dout(G284),.din(w_dff_A_X9VjWtUB8_0),.clk(gclk));
	jdff dff_A_X70tw3Lb1_1(.dout(w_dff_A_ivQxTsSS9_0),.din(w_dff_A_X70tw3Lb1_1),.clk(gclk));
	jdff dff_A_ivQxTsSS9_0(.dout(w_dff_A_bbtb0N6U5_0),.din(w_dff_A_ivQxTsSS9_0),.clk(gclk));
	jdff dff_A_bbtb0N6U5_0(.dout(w_dff_A_hPzLgahQ0_0),.din(w_dff_A_bbtb0N6U5_0),.clk(gclk));
	jdff dff_A_hPzLgahQ0_0(.dout(w_dff_A_2Nla7SxG5_0),.din(w_dff_A_hPzLgahQ0_0),.clk(gclk));
	jdff dff_A_2Nla7SxG5_0(.dout(w_dff_A_mVvi4glR3_0),.din(w_dff_A_2Nla7SxG5_0),.clk(gclk));
	jdff dff_A_mVvi4glR3_0(.dout(w_dff_A_Dzv8NsPq9_0),.din(w_dff_A_mVvi4glR3_0),.clk(gclk));
	jdff dff_A_Dzv8NsPq9_0(.dout(w_dff_A_22z3wZQn7_0),.din(w_dff_A_Dzv8NsPq9_0),.clk(gclk));
	jdff dff_A_22z3wZQn7_0(.dout(w_dff_A_s9tWOigg2_0),.din(w_dff_A_22z3wZQn7_0),.clk(gclk));
	jdff dff_A_s9tWOigg2_0(.dout(w_dff_A_H3DCpLJK0_0),.din(w_dff_A_s9tWOigg2_0),.clk(gclk));
	jdff dff_A_H3DCpLJK0_0(.dout(w_dff_A_s43xw4uT1_0),.din(w_dff_A_H3DCpLJK0_0),.clk(gclk));
	jdff dff_A_s43xw4uT1_0(.dout(w_dff_A_pywCpTOG2_0),.din(w_dff_A_s43xw4uT1_0),.clk(gclk));
	jdff dff_A_pywCpTOG2_0(.dout(w_dff_A_fXXipKZO0_0),.din(w_dff_A_pywCpTOG2_0),.clk(gclk));
	jdff dff_A_fXXipKZO0_0(.dout(w_dff_A_1Vhkare43_0),.din(w_dff_A_fXXipKZO0_0),.clk(gclk));
	jdff dff_A_1Vhkare43_0(.dout(w_dff_A_3tbOnTc90_0),.din(w_dff_A_1Vhkare43_0),.clk(gclk));
	jdff dff_A_3tbOnTc90_0(.dout(w_dff_A_IVfxt1M71_0),.din(w_dff_A_3tbOnTc90_0),.clk(gclk));
	jdff dff_A_IVfxt1M71_0(.dout(w_dff_A_SAgrBDqA8_0),.din(w_dff_A_IVfxt1M71_0),.clk(gclk));
	jdff dff_A_SAgrBDqA8_0(.dout(w_dff_A_gruBKQpP1_0),.din(w_dff_A_SAgrBDqA8_0),.clk(gclk));
	jdff dff_A_gruBKQpP1_0(.dout(w_dff_A_QIAjReQU7_0),.din(w_dff_A_gruBKQpP1_0),.clk(gclk));
	jdff dff_A_QIAjReQU7_0(.dout(w_dff_A_jUh98gZM4_0),.din(w_dff_A_QIAjReQU7_0),.clk(gclk));
	jdff dff_A_jUh98gZM4_0(.dout(w_dff_A_YX9ndtTA1_0),.din(w_dff_A_jUh98gZM4_0),.clk(gclk));
	jdff dff_A_YX9ndtTA1_0(.dout(w_dff_A_AMOmrFv77_0),.din(w_dff_A_YX9ndtTA1_0),.clk(gclk));
	jdff dff_A_AMOmrFv77_0(.dout(w_dff_A_vmednM2Z1_0),.din(w_dff_A_AMOmrFv77_0),.clk(gclk));
	jdff dff_A_vmednM2Z1_0(.dout(w_dff_A_9t4FJwtc1_0),.din(w_dff_A_vmednM2Z1_0),.clk(gclk));
	jdff dff_A_9t4FJwtc1_0(.dout(w_dff_A_JqeIkt3S9_0),.din(w_dff_A_9t4FJwtc1_0),.clk(gclk));
	jdff dff_A_JqeIkt3S9_0(.dout(w_dff_A_bJdDKUnI4_0),.din(w_dff_A_JqeIkt3S9_0),.clk(gclk));
	jdff dff_A_bJdDKUnI4_0(.dout(G286),.din(w_dff_A_bJdDKUnI4_0),.clk(gclk));
	jdff dff_A_B1dnqkxZ4_2(.dout(w_dff_A_FjlWCj2b4_0),.din(w_dff_A_B1dnqkxZ4_2),.clk(gclk));
	jdff dff_A_FjlWCj2b4_0(.dout(w_dff_A_Ob68xE3g0_0),.din(w_dff_A_FjlWCj2b4_0),.clk(gclk));
	jdff dff_A_Ob68xE3g0_0(.dout(w_dff_A_SRZrteZt4_0),.din(w_dff_A_Ob68xE3g0_0),.clk(gclk));
	jdff dff_A_SRZrteZt4_0(.dout(w_dff_A_BjoHQKXg5_0),.din(w_dff_A_SRZrteZt4_0),.clk(gclk));
	jdff dff_A_BjoHQKXg5_0(.dout(w_dff_A_Ys4vWhET0_0),.din(w_dff_A_BjoHQKXg5_0),.clk(gclk));
	jdff dff_A_Ys4vWhET0_0(.dout(w_dff_A_9U4sHRSA4_0),.din(w_dff_A_Ys4vWhET0_0),.clk(gclk));
	jdff dff_A_9U4sHRSA4_0(.dout(w_dff_A_RiaeiVOj0_0),.din(w_dff_A_9U4sHRSA4_0),.clk(gclk));
	jdff dff_A_RiaeiVOj0_0(.dout(w_dff_A_tqr91HKx9_0),.din(w_dff_A_RiaeiVOj0_0),.clk(gclk));
	jdff dff_A_tqr91HKx9_0(.dout(w_dff_A_td3SoSxZ4_0),.din(w_dff_A_tqr91HKx9_0),.clk(gclk));
	jdff dff_A_td3SoSxZ4_0(.dout(w_dff_A_B5xA7uuC2_0),.din(w_dff_A_td3SoSxZ4_0),.clk(gclk));
	jdff dff_A_B5xA7uuC2_0(.dout(w_dff_A_7i0u7VnG0_0),.din(w_dff_A_B5xA7uuC2_0),.clk(gclk));
	jdff dff_A_7i0u7VnG0_0(.dout(w_dff_A_uvS5cts93_0),.din(w_dff_A_7i0u7VnG0_0),.clk(gclk));
	jdff dff_A_uvS5cts93_0(.dout(w_dff_A_jtelvk5G4_0),.din(w_dff_A_uvS5cts93_0),.clk(gclk));
	jdff dff_A_jtelvk5G4_0(.dout(w_dff_A_ffF48l0z7_0),.din(w_dff_A_jtelvk5G4_0),.clk(gclk));
	jdff dff_A_ffF48l0z7_0(.dout(w_dff_A_PFBddvsS8_0),.din(w_dff_A_ffF48l0z7_0),.clk(gclk));
	jdff dff_A_PFBddvsS8_0(.dout(w_dff_A_EoD8049A5_0),.din(w_dff_A_PFBddvsS8_0),.clk(gclk));
	jdff dff_A_EoD8049A5_0(.dout(w_dff_A_qO8Kzqhg2_0),.din(w_dff_A_EoD8049A5_0),.clk(gclk));
	jdff dff_A_qO8Kzqhg2_0(.dout(w_dff_A_K8MY7GbE9_0),.din(w_dff_A_qO8Kzqhg2_0),.clk(gclk));
	jdff dff_A_K8MY7GbE9_0(.dout(w_dff_A_RVwgB2Tj4_0),.din(w_dff_A_K8MY7GbE9_0),.clk(gclk));
	jdff dff_A_RVwgB2Tj4_0(.dout(w_dff_A_MQJAntPL9_0),.din(w_dff_A_RVwgB2Tj4_0),.clk(gclk));
	jdff dff_A_MQJAntPL9_0(.dout(w_dff_A_nPVIIYij4_0),.din(w_dff_A_MQJAntPL9_0),.clk(gclk));
	jdff dff_A_nPVIIYij4_0(.dout(w_dff_A_mpA9ibvw3_0),.din(w_dff_A_nPVIIYij4_0),.clk(gclk));
	jdff dff_A_mpA9ibvw3_0(.dout(w_dff_A_r6dNMP9X2_0),.din(w_dff_A_mpA9ibvw3_0),.clk(gclk));
	jdff dff_A_r6dNMP9X2_0(.dout(w_dff_A_jzj3M23R2_0),.din(w_dff_A_r6dNMP9X2_0),.clk(gclk));
	jdff dff_A_jzj3M23R2_0(.dout(G289),.din(w_dff_A_jzj3M23R2_0),.clk(gclk));
	jdff dff_A_Ti7Z5XKL2_2(.dout(w_dff_A_XZJSgp7Q0_0),.din(w_dff_A_Ti7Z5XKL2_2),.clk(gclk));
	jdff dff_A_XZJSgp7Q0_0(.dout(w_dff_A_6uYZIZJe3_0),.din(w_dff_A_XZJSgp7Q0_0),.clk(gclk));
	jdff dff_A_6uYZIZJe3_0(.dout(w_dff_A_kWDoJ2f79_0),.din(w_dff_A_6uYZIZJe3_0),.clk(gclk));
	jdff dff_A_kWDoJ2f79_0(.dout(w_dff_A_HwwT2VBs3_0),.din(w_dff_A_kWDoJ2f79_0),.clk(gclk));
	jdff dff_A_HwwT2VBs3_0(.dout(w_dff_A_0IYeoJO08_0),.din(w_dff_A_HwwT2VBs3_0),.clk(gclk));
	jdff dff_A_0IYeoJO08_0(.dout(w_dff_A_jYew3Hxd8_0),.din(w_dff_A_0IYeoJO08_0),.clk(gclk));
	jdff dff_A_jYew3Hxd8_0(.dout(w_dff_A_3Q53PGQx6_0),.din(w_dff_A_jYew3Hxd8_0),.clk(gclk));
	jdff dff_A_3Q53PGQx6_0(.dout(w_dff_A_DzcVN8oE2_0),.din(w_dff_A_3Q53PGQx6_0),.clk(gclk));
	jdff dff_A_DzcVN8oE2_0(.dout(w_dff_A_atxPUGMS8_0),.din(w_dff_A_DzcVN8oE2_0),.clk(gclk));
	jdff dff_A_atxPUGMS8_0(.dout(w_dff_A_jbFWPGkK0_0),.din(w_dff_A_atxPUGMS8_0),.clk(gclk));
	jdff dff_A_jbFWPGkK0_0(.dout(w_dff_A_uYEAjJdY3_0),.din(w_dff_A_jbFWPGkK0_0),.clk(gclk));
	jdff dff_A_uYEAjJdY3_0(.dout(w_dff_A_WltOxQ4d6_0),.din(w_dff_A_uYEAjJdY3_0),.clk(gclk));
	jdff dff_A_WltOxQ4d6_0(.dout(w_dff_A_yq4ktUSW8_0),.din(w_dff_A_WltOxQ4d6_0),.clk(gclk));
	jdff dff_A_yq4ktUSW8_0(.dout(w_dff_A_Xr7dG80L3_0),.din(w_dff_A_yq4ktUSW8_0),.clk(gclk));
	jdff dff_A_Xr7dG80L3_0(.dout(w_dff_A_3NTHNzxg5_0),.din(w_dff_A_Xr7dG80L3_0),.clk(gclk));
	jdff dff_A_3NTHNzxg5_0(.dout(w_dff_A_eCEWwOLG8_0),.din(w_dff_A_3NTHNzxg5_0),.clk(gclk));
	jdff dff_A_eCEWwOLG8_0(.dout(w_dff_A_BQ2wGKp42_0),.din(w_dff_A_eCEWwOLG8_0),.clk(gclk));
	jdff dff_A_BQ2wGKp42_0(.dout(w_dff_A_uKEtiqzL7_0),.din(w_dff_A_BQ2wGKp42_0),.clk(gclk));
	jdff dff_A_uKEtiqzL7_0(.dout(w_dff_A_WB6mi2477_0),.din(w_dff_A_uKEtiqzL7_0),.clk(gclk));
	jdff dff_A_WB6mi2477_0(.dout(w_dff_A_mTDUt9HN2_0),.din(w_dff_A_WB6mi2477_0),.clk(gclk));
	jdff dff_A_mTDUt9HN2_0(.dout(w_dff_A_4UzhitIC0_0),.din(w_dff_A_mTDUt9HN2_0),.clk(gclk));
	jdff dff_A_4UzhitIC0_0(.dout(w_dff_A_tVeKdouP0_0),.din(w_dff_A_4UzhitIC0_0),.clk(gclk));
	jdff dff_A_tVeKdouP0_0(.dout(w_dff_A_sSTDtCZF9_0),.din(w_dff_A_tVeKdouP0_0),.clk(gclk));
	jdff dff_A_sSTDtCZF9_0(.dout(G292),.din(w_dff_A_sSTDtCZF9_0),.clk(gclk));
	jdff dff_A_w5MdrG526_1(.dout(w_dff_A_ZmDIu1cI5_0),.din(w_dff_A_w5MdrG526_1),.clk(gclk));
	jdff dff_A_ZmDIu1cI5_0(.dout(w_dff_A_RGEZTkao7_0),.din(w_dff_A_ZmDIu1cI5_0),.clk(gclk));
	jdff dff_A_RGEZTkao7_0(.dout(w_dff_A_RowHP7Ov6_0),.din(w_dff_A_RGEZTkao7_0),.clk(gclk));
	jdff dff_A_RowHP7Ov6_0(.dout(w_dff_A_KQ3zL1Bu0_0),.din(w_dff_A_RowHP7Ov6_0),.clk(gclk));
	jdff dff_A_KQ3zL1Bu0_0(.dout(w_dff_A_Z58CL2R31_0),.din(w_dff_A_KQ3zL1Bu0_0),.clk(gclk));
	jdff dff_A_Z58CL2R31_0(.dout(w_dff_A_vL7Wn4443_0),.din(w_dff_A_Z58CL2R31_0),.clk(gclk));
	jdff dff_A_vL7Wn4443_0(.dout(w_dff_A_x2gAadT62_0),.din(w_dff_A_vL7Wn4443_0),.clk(gclk));
	jdff dff_A_x2gAadT62_0(.dout(w_dff_A_frIeChTW7_0),.din(w_dff_A_x2gAadT62_0),.clk(gclk));
	jdff dff_A_frIeChTW7_0(.dout(w_dff_A_Z2Wsc5eu7_0),.din(w_dff_A_frIeChTW7_0),.clk(gclk));
	jdff dff_A_Z2Wsc5eu7_0(.dout(w_dff_A_re6X1cVW3_0),.din(w_dff_A_Z2Wsc5eu7_0),.clk(gclk));
	jdff dff_A_re6X1cVW3_0(.dout(w_dff_A_mwV8252j8_0),.din(w_dff_A_re6X1cVW3_0),.clk(gclk));
	jdff dff_A_mwV8252j8_0(.dout(w_dff_A_oNmloiZZ7_0),.din(w_dff_A_mwV8252j8_0),.clk(gclk));
	jdff dff_A_oNmloiZZ7_0(.dout(w_dff_A_7bf8dao58_0),.din(w_dff_A_oNmloiZZ7_0),.clk(gclk));
	jdff dff_A_7bf8dao58_0(.dout(w_dff_A_I6Pd9k5c6_0),.din(w_dff_A_7bf8dao58_0),.clk(gclk));
	jdff dff_A_I6Pd9k5c6_0(.dout(w_dff_A_VFB3a0un3_0),.din(w_dff_A_I6Pd9k5c6_0),.clk(gclk));
	jdff dff_A_VFB3a0un3_0(.dout(w_dff_A_bnM2uTsC1_0),.din(w_dff_A_VFB3a0un3_0),.clk(gclk));
	jdff dff_A_bnM2uTsC1_0(.dout(w_dff_A_qKiuXRsu4_0),.din(w_dff_A_bnM2uTsC1_0),.clk(gclk));
	jdff dff_A_qKiuXRsu4_0(.dout(w_dff_A_Px8UShAx9_0),.din(w_dff_A_qKiuXRsu4_0),.clk(gclk));
	jdff dff_A_Px8UShAx9_0(.dout(w_dff_A_PDcYMmLt2_0),.din(w_dff_A_Px8UShAx9_0),.clk(gclk));
	jdff dff_A_PDcYMmLt2_0(.dout(w_dff_A_IJyfc8eZ7_0),.din(w_dff_A_PDcYMmLt2_0),.clk(gclk));
	jdff dff_A_IJyfc8eZ7_0(.dout(w_dff_A_Rau2rxJ47_0),.din(w_dff_A_IJyfc8eZ7_0),.clk(gclk));
	jdff dff_A_Rau2rxJ47_0(.dout(w_dff_A_CHKqgrw39_0),.din(w_dff_A_Rau2rxJ47_0),.clk(gclk));
	jdff dff_A_CHKqgrw39_0(.dout(w_dff_A_jJFIApff5_0),.din(w_dff_A_CHKqgrw39_0),.clk(gclk));
	jdff dff_A_jJFIApff5_0(.dout(w_dff_A_TUnYOaP23_0),.din(w_dff_A_jJFIApff5_0),.clk(gclk));
	jdff dff_A_TUnYOaP23_0(.dout(w_dff_A_ypRPQATu8_0),.din(w_dff_A_TUnYOaP23_0),.clk(gclk));
	jdff dff_A_ypRPQATu8_0(.dout(G341),.din(w_dff_A_ypRPQATu8_0),.clk(gclk));
	jdff dff_A_KrEOdKkt7_2(.dout(w_dff_A_mVZ1O6Hg3_0),.din(w_dff_A_KrEOdKkt7_2),.clk(gclk));
	jdff dff_A_mVZ1O6Hg3_0(.dout(w_dff_A_OgrGov5P8_0),.din(w_dff_A_mVZ1O6Hg3_0),.clk(gclk));
	jdff dff_A_OgrGov5P8_0(.dout(w_dff_A_CCfZjVuf9_0),.din(w_dff_A_OgrGov5P8_0),.clk(gclk));
	jdff dff_A_CCfZjVuf9_0(.dout(w_dff_A_JBkwmDO49_0),.din(w_dff_A_CCfZjVuf9_0),.clk(gclk));
	jdff dff_A_JBkwmDO49_0(.dout(w_dff_A_dd5Lt2ZD9_0),.din(w_dff_A_JBkwmDO49_0),.clk(gclk));
	jdff dff_A_dd5Lt2ZD9_0(.dout(w_dff_A_JnR1XVpz2_0),.din(w_dff_A_dd5Lt2ZD9_0),.clk(gclk));
	jdff dff_A_JnR1XVpz2_0(.dout(w_dff_A_mfh1uOZu7_0),.din(w_dff_A_JnR1XVpz2_0),.clk(gclk));
	jdff dff_A_mfh1uOZu7_0(.dout(w_dff_A_qdpVz5IX4_0),.din(w_dff_A_mfh1uOZu7_0),.clk(gclk));
	jdff dff_A_qdpVz5IX4_0(.dout(w_dff_A_CDgFEVpt9_0),.din(w_dff_A_qdpVz5IX4_0),.clk(gclk));
	jdff dff_A_CDgFEVpt9_0(.dout(w_dff_A_aZe4e1ew5_0),.din(w_dff_A_CDgFEVpt9_0),.clk(gclk));
	jdff dff_A_aZe4e1ew5_0(.dout(w_dff_A_TGP3O5wA8_0),.din(w_dff_A_aZe4e1ew5_0),.clk(gclk));
	jdff dff_A_TGP3O5wA8_0(.dout(w_dff_A_1CjAG2pP2_0),.din(w_dff_A_TGP3O5wA8_0),.clk(gclk));
	jdff dff_A_1CjAG2pP2_0(.dout(w_dff_A_euzOGjlo0_0),.din(w_dff_A_1CjAG2pP2_0),.clk(gclk));
	jdff dff_A_euzOGjlo0_0(.dout(w_dff_A_Vf3PdFCW9_0),.din(w_dff_A_euzOGjlo0_0),.clk(gclk));
	jdff dff_A_Vf3PdFCW9_0(.dout(w_dff_A_WuzeQQ1s7_0),.din(w_dff_A_Vf3PdFCW9_0),.clk(gclk));
	jdff dff_A_WuzeQQ1s7_0(.dout(w_dff_A_t8W8UlgB0_0),.din(w_dff_A_WuzeQQ1s7_0),.clk(gclk));
	jdff dff_A_t8W8UlgB0_0(.dout(w_dff_A_LtRtOvmL0_0),.din(w_dff_A_t8W8UlgB0_0),.clk(gclk));
	jdff dff_A_LtRtOvmL0_0(.dout(w_dff_A_ItvX0lT74_0),.din(w_dff_A_LtRtOvmL0_0),.clk(gclk));
	jdff dff_A_ItvX0lT74_0(.dout(w_dff_A_vLeYnClR3_0),.din(w_dff_A_ItvX0lT74_0),.clk(gclk));
	jdff dff_A_vLeYnClR3_0(.dout(w_dff_A_cuKXS15k1_0),.din(w_dff_A_vLeYnClR3_0),.clk(gclk));
	jdff dff_A_cuKXS15k1_0(.dout(w_dff_A_ERkJuYSS5_0),.din(w_dff_A_cuKXS15k1_0),.clk(gclk));
	jdff dff_A_ERkJuYSS5_0(.dout(w_dff_A_JU682vyY6_0),.din(w_dff_A_ERkJuYSS5_0),.clk(gclk));
	jdff dff_A_JU682vyY6_0(.dout(w_dff_A_iq9tyi289_0),.din(w_dff_A_JU682vyY6_0),.clk(gclk));
	jdff dff_A_iq9tyi289_0(.dout(G281),.din(w_dff_A_iq9tyi289_0),.clk(gclk));
	jdff dff_A_WfeN12RN7_1(.dout(w_dff_A_tZyf03n89_0),.din(w_dff_A_WfeN12RN7_1),.clk(gclk));
	jdff dff_A_tZyf03n89_0(.dout(w_dff_A_Gjvg1V2t4_0),.din(w_dff_A_tZyf03n89_0),.clk(gclk));
	jdff dff_A_Gjvg1V2t4_0(.dout(w_dff_A_azWxccFr5_0),.din(w_dff_A_Gjvg1V2t4_0),.clk(gclk));
	jdff dff_A_azWxccFr5_0(.dout(w_dff_A_CtB9QTOK3_0),.din(w_dff_A_azWxccFr5_0),.clk(gclk));
	jdff dff_A_CtB9QTOK3_0(.dout(w_dff_A_8ZxcYVqP1_0),.din(w_dff_A_CtB9QTOK3_0),.clk(gclk));
	jdff dff_A_8ZxcYVqP1_0(.dout(w_dff_A_NtXSZeMD2_0),.din(w_dff_A_8ZxcYVqP1_0),.clk(gclk));
	jdff dff_A_NtXSZeMD2_0(.dout(w_dff_A_IFbVjk4p0_0),.din(w_dff_A_NtXSZeMD2_0),.clk(gclk));
	jdff dff_A_IFbVjk4p0_0(.dout(w_dff_A_tmjihczE0_0),.din(w_dff_A_IFbVjk4p0_0),.clk(gclk));
	jdff dff_A_tmjihczE0_0(.dout(w_dff_A_mJaz4RL47_0),.din(w_dff_A_tmjihczE0_0),.clk(gclk));
	jdff dff_A_mJaz4RL47_0(.dout(w_dff_A_jGsiy5Vs4_0),.din(w_dff_A_mJaz4RL47_0),.clk(gclk));
	jdff dff_A_jGsiy5Vs4_0(.dout(w_dff_A_cWKhQbOq7_0),.din(w_dff_A_jGsiy5Vs4_0),.clk(gclk));
	jdff dff_A_cWKhQbOq7_0(.dout(w_dff_A_l2yFXSXP9_0),.din(w_dff_A_cWKhQbOq7_0),.clk(gclk));
	jdff dff_A_l2yFXSXP9_0(.dout(w_dff_A_4AJOowQ61_0),.din(w_dff_A_l2yFXSXP9_0),.clk(gclk));
	jdff dff_A_4AJOowQ61_0(.dout(w_dff_A_Ggj6PLQA7_0),.din(w_dff_A_4AJOowQ61_0),.clk(gclk));
	jdff dff_A_Ggj6PLQA7_0(.dout(w_dff_A_sCvFeNMs8_0),.din(w_dff_A_Ggj6PLQA7_0),.clk(gclk));
	jdff dff_A_sCvFeNMs8_0(.dout(w_dff_A_Pr7Qdmus9_0),.din(w_dff_A_sCvFeNMs8_0),.clk(gclk));
	jdff dff_A_Pr7Qdmus9_0(.dout(w_dff_A_828TThmF2_0),.din(w_dff_A_Pr7Qdmus9_0),.clk(gclk));
	jdff dff_A_828TThmF2_0(.dout(w_dff_A_kMdQl0sT9_0),.din(w_dff_A_828TThmF2_0),.clk(gclk));
	jdff dff_A_kMdQl0sT9_0(.dout(w_dff_A_rw9JupFW6_0),.din(w_dff_A_kMdQl0sT9_0),.clk(gclk));
	jdff dff_A_rw9JupFW6_0(.dout(w_dff_A_6YDxurMj0_0),.din(w_dff_A_rw9JupFW6_0),.clk(gclk));
	jdff dff_A_6YDxurMj0_0(.dout(w_dff_A_nJBLzrFr4_0),.din(w_dff_A_6YDxurMj0_0),.clk(gclk));
	jdff dff_A_nJBLzrFr4_0(.dout(w_dff_A_jI5PA4cr5_0),.din(w_dff_A_nJBLzrFr4_0),.clk(gclk));
	jdff dff_A_jI5PA4cr5_0(.dout(w_dff_A_8JYjHguq9_0),.din(w_dff_A_jI5PA4cr5_0),.clk(gclk));
	jdff dff_A_8JYjHguq9_0(.dout(w_dff_A_LnjKUAvC2_0),.din(w_dff_A_8JYjHguq9_0),.clk(gclk));
	jdff dff_A_LnjKUAvC2_0(.dout(w_dff_A_ZsdjeHLx7_0),.din(w_dff_A_LnjKUAvC2_0),.clk(gclk));
	jdff dff_A_ZsdjeHLx7_0(.dout(G453),.din(w_dff_A_ZsdjeHLx7_0),.clk(gclk));
	jdff dff_A_NHAxy8Qq4_2(.dout(w_dff_A_Ed2rPu1D0_0),.din(w_dff_A_NHAxy8Qq4_2),.clk(gclk));
	jdff dff_A_Ed2rPu1D0_0(.dout(w_dff_A_5GKxlkRZ6_0),.din(w_dff_A_Ed2rPu1D0_0),.clk(gclk));
	jdff dff_A_5GKxlkRZ6_0(.dout(w_dff_A_12W7fw4g4_0),.din(w_dff_A_5GKxlkRZ6_0),.clk(gclk));
	jdff dff_A_12W7fw4g4_0(.dout(w_dff_A_qnwoH1QE8_0),.din(w_dff_A_12W7fw4g4_0),.clk(gclk));
	jdff dff_A_qnwoH1QE8_0(.dout(w_dff_A_l4jzBRgz9_0),.din(w_dff_A_qnwoH1QE8_0),.clk(gclk));
	jdff dff_A_l4jzBRgz9_0(.dout(w_dff_A_g855YBmC2_0),.din(w_dff_A_l4jzBRgz9_0),.clk(gclk));
	jdff dff_A_g855YBmC2_0(.dout(w_dff_A_9HW4GkQG2_0),.din(w_dff_A_g855YBmC2_0),.clk(gclk));
	jdff dff_A_9HW4GkQG2_0(.dout(w_dff_A_lpZiuo7Q5_0),.din(w_dff_A_9HW4GkQG2_0),.clk(gclk));
	jdff dff_A_lpZiuo7Q5_0(.dout(w_dff_A_Vywao6KF8_0),.din(w_dff_A_lpZiuo7Q5_0),.clk(gclk));
	jdff dff_A_Vywao6KF8_0(.dout(w_dff_A_uB2ThT4B7_0),.din(w_dff_A_Vywao6KF8_0),.clk(gclk));
	jdff dff_A_uB2ThT4B7_0(.dout(w_dff_A_EKIfQgUg4_0),.din(w_dff_A_uB2ThT4B7_0),.clk(gclk));
	jdff dff_A_EKIfQgUg4_0(.dout(w_dff_A_rFhaQCry4_0),.din(w_dff_A_EKIfQgUg4_0),.clk(gclk));
	jdff dff_A_rFhaQCry4_0(.dout(w_dff_A_4lu8Ud9g5_0),.din(w_dff_A_rFhaQCry4_0),.clk(gclk));
	jdff dff_A_4lu8Ud9g5_0(.dout(w_dff_A_NsMAW75Q4_0),.din(w_dff_A_4lu8Ud9g5_0),.clk(gclk));
	jdff dff_A_NsMAW75Q4_0(.dout(w_dff_A_u37X9amP7_0),.din(w_dff_A_NsMAW75Q4_0),.clk(gclk));
	jdff dff_A_u37X9amP7_0(.dout(w_dff_A_hIO7XOSO3_0),.din(w_dff_A_u37X9amP7_0),.clk(gclk));
	jdff dff_A_hIO7XOSO3_0(.dout(w_dff_A_juM6jieX6_0),.din(w_dff_A_hIO7XOSO3_0),.clk(gclk));
	jdff dff_A_juM6jieX6_0(.dout(w_dff_A_Kk3CIjBV7_0),.din(w_dff_A_juM6jieX6_0),.clk(gclk));
	jdff dff_A_Kk3CIjBV7_0(.dout(w_dff_A_FvC1yZEg1_0),.din(w_dff_A_Kk3CIjBV7_0),.clk(gclk));
	jdff dff_A_FvC1yZEg1_0(.dout(w_dff_A_6uv0cKzz0_0),.din(w_dff_A_FvC1yZEg1_0),.clk(gclk));
	jdff dff_A_6uv0cKzz0_0(.dout(w_dff_A_1KH2B4jk1_0),.din(w_dff_A_6uv0cKzz0_0),.clk(gclk));
	jdff dff_A_1KH2B4jk1_0(.dout(w_dff_A_aRdiGPis4_0),.din(w_dff_A_1KH2B4jk1_0),.clk(gclk));
	jdff dff_A_aRdiGPis4_0(.dout(w_dff_A_g3TADX9Q0_0),.din(w_dff_A_aRdiGPis4_0),.clk(gclk));
	jdff dff_A_g3TADX9Q0_0(.dout(w_dff_A_FTt1kzgv0_0),.din(w_dff_A_g3TADX9Q0_0),.clk(gclk));
	jdff dff_A_FTt1kzgv0_0(.dout(w_dff_A_616RzkKH1_0),.din(w_dff_A_FTt1kzgv0_0),.clk(gclk));
	jdff dff_A_616RzkKH1_0(.dout(G278),.din(w_dff_A_616RzkKH1_0),.clk(gclk));
	jdff dff_A_CGluyyLx8_2(.dout(w_dff_A_7g34HPfj9_0),.din(w_dff_A_CGluyyLx8_2),.clk(gclk));
	jdff dff_A_7g34HPfj9_0(.dout(w_dff_A_VHezfZ6H0_0),.din(w_dff_A_7g34HPfj9_0),.clk(gclk));
	jdff dff_A_VHezfZ6H0_0(.dout(w_dff_A_AW4dAvYN2_0),.din(w_dff_A_VHezfZ6H0_0),.clk(gclk));
	jdff dff_A_AW4dAvYN2_0(.dout(w_dff_A_k30oTUpH7_0),.din(w_dff_A_AW4dAvYN2_0),.clk(gclk));
	jdff dff_A_k30oTUpH7_0(.dout(w_dff_A_RViSHWIa6_0),.din(w_dff_A_k30oTUpH7_0),.clk(gclk));
	jdff dff_A_RViSHWIa6_0(.dout(w_dff_A_UkK3hfsn5_0),.din(w_dff_A_RViSHWIa6_0),.clk(gclk));
	jdff dff_A_UkK3hfsn5_0(.dout(w_dff_A_cRyE3iZd2_0),.din(w_dff_A_UkK3hfsn5_0),.clk(gclk));
	jdff dff_A_cRyE3iZd2_0(.dout(w_dff_A_0FfUMgF40_0),.din(w_dff_A_cRyE3iZd2_0),.clk(gclk));
	jdff dff_A_0FfUMgF40_0(.dout(w_dff_A_ffppzAl97_0),.din(w_dff_A_0FfUMgF40_0),.clk(gclk));
	jdff dff_A_ffppzAl97_0(.dout(w_dff_A_7lvWxaUV1_0),.din(w_dff_A_ffppzAl97_0),.clk(gclk));
	jdff dff_A_7lvWxaUV1_0(.dout(w_dff_A_rDQulIv00_0),.din(w_dff_A_7lvWxaUV1_0),.clk(gclk));
	jdff dff_A_rDQulIv00_0(.dout(w_dff_A_2K8I8pYJ2_0),.din(w_dff_A_rDQulIv00_0),.clk(gclk));
	jdff dff_A_2K8I8pYJ2_0(.dout(w_dff_A_duZ6ox7B9_0),.din(w_dff_A_2K8I8pYJ2_0),.clk(gclk));
	jdff dff_A_duZ6ox7B9_0(.dout(w_dff_A_J9CsCj704_0),.din(w_dff_A_duZ6ox7B9_0),.clk(gclk));
	jdff dff_A_J9CsCj704_0(.dout(w_dff_A_IZKCF9bv4_0),.din(w_dff_A_J9CsCj704_0),.clk(gclk));
	jdff dff_A_IZKCF9bv4_0(.dout(w_dff_A_tUg9irBn6_0),.din(w_dff_A_IZKCF9bv4_0),.clk(gclk));
	jdff dff_A_tUg9irBn6_0(.dout(w_dff_A_aOg81CMv9_0),.din(w_dff_A_tUg9irBn6_0),.clk(gclk));
	jdff dff_A_aOg81CMv9_0(.dout(w_dff_A_AOegXKqA3_0),.din(w_dff_A_aOg81CMv9_0),.clk(gclk));
	jdff dff_A_AOegXKqA3_0(.dout(w_dff_A_wt6Hobxm6_0),.din(w_dff_A_AOegXKqA3_0),.clk(gclk));
	jdff dff_A_wt6Hobxm6_0(.dout(w_dff_A_Vdzrohec1_0),.din(w_dff_A_wt6Hobxm6_0),.clk(gclk));
	jdff dff_A_Vdzrohec1_0(.dout(G373),.din(w_dff_A_Vdzrohec1_0),.clk(gclk));
	jdff dff_A_R2YdaLCt7_2(.dout(G246),.din(w_dff_A_R2YdaLCt7_2),.clk(gclk));
	jdff dff_A_Q0JJXQ6q2_2(.dout(w_dff_A_EolVQK7x9_0),.din(w_dff_A_Q0JJXQ6q2_2),.clk(gclk));
	jdff dff_A_EolVQK7x9_0(.dout(w_dff_A_sC8XpTxb0_0),.din(w_dff_A_EolVQK7x9_0),.clk(gclk));
	jdff dff_A_sC8XpTxb0_0(.dout(w_dff_A_mlraThnj5_0),.din(w_dff_A_sC8XpTxb0_0),.clk(gclk));
	jdff dff_A_mlraThnj5_0(.dout(w_dff_A_hqOvNHIe1_0),.din(w_dff_A_mlraThnj5_0),.clk(gclk));
	jdff dff_A_hqOvNHIe1_0(.dout(w_dff_A_xBLn3BnK2_0),.din(w_dff_A_hqOvNHIe1_0),.clk(gclk));
	jdff dff_A_xBLn3BnK2_0(.dout(w_dff_A_VxpAgs9w9_0),.din(w_dff_A_xBLn3BnK2_0),.clk(gclk));
	jdff dff_A_VxpAgs9w9_0(.dout(G258),.din(w_dff_A_VxpAgs9w9_0),.clk(gclk));
	jdff dff_A_A5XS2GlF0_2(.dout(w_dff_A_NfaO50cd0_0),.din(w_dff_A_A5XS2GlF0_2),.clk(gclk));
	jdff dff_A_NfaO50cd0_0(.dout(w_dff_A_WaQ6FwW05_0),.din(w_dff_A_NfaO50cd0_0),.clk(gclk));
	jdff dff_A_WaQ6FwW05_0(.dout(w_dff_A_XCW9JrQp7_0),.din(w_dff_A_WaQ6FwW05_0),.clk(gclk));
	jdff dff_A_XCW9JrQp7_0(.dout(w_dff_A_B7VaiMwO9_0),.din(w_dff_A_XCW9JrQp7_0),.clk(gclk));
	jdff dff_A_B7VaiMwO9_0(.dout(w_dff_A_0qrM3nOe3_0),.din(w_dff_A_B7VaiMwO9_0),.clk(gclk));
	jdff dff_A_0qrM3nOe3_0(.dout(w_dff_A_k292zF0g9_0),.din(w_dff_A_0qrM3nOe3_0),.clk(gclk));
	jdff dff_A_k292zF0g9_0(.dout(G264),.din(w_dff_A_k292zF0g9_0),.clk(gclk));
	jdff dff_A_nl5Rctji5_2(.dout(G270),.din(w_dff_A_nl5Rctji5_2),.clk(gclk));
	jdff dff_A_l9LCgxGv9_2(.dout(w_dff_A_kyTaRLFF9_0),.din(w_dff_A_l9LCgxGv9_2),.clk(gclk));
	jdff dff_A_kyTaRLFF9_0(.dout(w_dff_A_cYIudUaM3_0),.din(w_dff_A_kyTaRLFF9_0),.clk(gclk));
	jdff dff_A_cYIudUaM3_0(.dout(w_dff_A_LfJ9L3gi7_0),.din(w_dff_A_cYIudUaM3_0),.clk(gclk));
	jdff dff_A_LfJ9L3gi7_0(.dout(w_dff_A_DstrArim9_0),.din(w_dff_A_LfJ9L3gi7_0),.clk(gclk));
	jdff dff_A_DstrArim9_0(.dout(w_dff_A_CRC1ax6O2_0),.din(w_dff_A_DstrArim9_0),.clk(gclk));
	jdff dff_A_CRC1ax6O2_0(.dout(w_dff_A_RgXVgALg9_0),.din(w_dff_A_CRC1ax6O2_0),.clk(gclk));
	jdff dff_A_RgXVgALg9_0(.dout(w_dff_A_RL0IalGz4_0),.din(w_dff_A_RgXVgALg9_0),.clk(gclk));
	jdff dff_A_RL0IalGz4_0(.dout(w_dff_A_lfTIEuZs4_0),.din(w_dff_A_RL0IalGz4_0),.clk(gclk));
	jdff dff_A_lfTIEuZs4_0(.dout(w_dff_A_AXXGvaV37_0),.din(w_dff_A_lfTIEuZs4_0),.clk(gclk));
	jdff dff_A_AXXGvaV37_0(.dout(w_dff_A_REsitmqL9_0),.din(w_dff_A_AXXGvaV37_0),.clk(gclk));
	jdff dff_A_REsitmqL9_0(.dout(w_dff_A_PBnnuB6u7_0),.din(w_dff_A_REsitmqL9_0),.clk(gclk));
	jdff dff_A_PBnnuB6u7_0(.dout(w_dff_A_XE6rjJ8Q7_0),.din(w_dff_A_PBnnuB6u7_0),.clk(gclk));
	jdff dff_A_XE6rjJ8Q7_0(.dout(w_dff_A_Uw3YYzYS7_0),.din(w_dff_A_XE6rjJ8Q7_0),.clk(gclk));
	jdff dff_A_Uw3YYzYS7_0(.dout(w_dff_A_iTOYy22w6_0),.din(w_dff_A_Uw3YYzYS7_0),.clk(gclk));
	jdff dff_A_iTOYy22w6_0(.dout(G388),.din(w_dff_A_iTOYy22w6_0),.clk(gclk));
	jdff dff_A_f4MjxiJZ3_2(.dout(w_dff_A_YjJZ0vk19_0),.din(w_dff_A_f4MjxiJZ3_2),.clk(gclk));
	jdff dff_A_YjJZ0vk19_0(.dout(w_dff_A_evzt3vR01_0),.din(w_dff_A_YjJZ0vk19_0),.clk(gclk));
	jdff dff_A_evzt3vR01_0(.dout(w_dff_A_jJkwxnye2_0),.din(w_dff_A_evzt3vR01_0),.clk(gclk));
	jdff dff_A_jJkwxnye2_0(.dout(w_dff_A_nwtmSoKe8_0),.din(w_dff_A_jJkwxnye2_0),.clk(gclk));
	jdff dff_A_nwtmSoKe8_0(.dout(w_dff_A_h9k8PZIV0_0),.din(w_dff_A_nwtmSoKe8_0),.clk(gclk));
	jdff dff_A_h9k8PZIV0_0(.dout(w_dff_A_L7xEiLZH9_0),.din(w_dff_A_h9k8PZIV0_0),.clk(gclk));
	jdff dff_A_L7xEiLZH9_0(.dout(w_dff_A_fOBBr3vE7_0),.din(w_dff_A_L7xEiLZH9_0),.clk(gclk));
	jdff dff_A_fOBBr3vE7_0(.dout(w_dff_A_5Dx3uy0W1_0),.din(w_dff_A_fOBBr3vE7_0),.clk(gclk));
	jdff dff_A_5Dx3uy0W1_0(.dout(w_dff_A_RUKf3Paw2_0),.din(w_dff_A_5Dx3uy0W1_0),.clk(gclk));
	jdff dff_A_RUKf3Paw2_0(.dout(w_dff_A_5OJnOWhJ3_0),.din(w_dff_A_RUKf3Paw2_0),.clk(gclk));
	jdff dff_A_5OJnOWhJ3_0(.dout(w_dff_A_B1GN1IsM6_0),.din(w_dff_A_5OJnOWhJ3_0),.clk(gclk));
	jdff dff_A_B1GN1IsM6_0(.dout(w_dff_A_mRydFenQ2_0),.din(w_dff_A_B1GN1IsM6_0),.clk(gclk));
	jdff dff_A_mRydFenQ2_0(.dout(w_dff_A_bUZ8UM2f2_0),.din(w_dff_A_mRydFenQ2_0),.clk(gclk));
	jdff dff_A_bUZ8UM2f2_0(.dout(w_dff_A_hMRbFHPt0_0),.din(w_dff_A_bUZ8UM2f2_0),.clk(gclk));
	jdff dff_A_hMRbFHPt0_0(.dout(w_dff_A_ahq94RXh2_0),.din(w_dff_A_hMRbFHPt0_0),.clk(gclk));
	jdff dff_A_ahq94RXh2_0(.dout(w_dff_A_xb28ihKw9_0),.din(w_dff_A_ahq94RXh2_0),.clk(gclk));
	jdff dff_A_xb28ihKw9_0(.dout(G391),.din(w_dff_A_xb28ihKw9_0),.clk(gclk));
	jdff dff_A_wd3queQl0_2(.dout(w_dff_A_bGy4FE5o1_0),.din(w_dff_A_wd3queQl0_2),.clk(gclk));
	jdff dff_A_bGy4FE5o1_0(.dout(w_dff_A_JvoLXZv29_0),.din(w_dff_A_bGy4FE5o1_0),.clk(gclk));
	jdff dff_A_JvoLXZv29_0(.dout(w_dff_A_nc2zuewP2_0),.din(w_dff_A_JvoLXZv29_0),.clk(gclk));
	jdff dff_A_nc2zuewP2_0(.dout(w_dff_A_fEJYJaC64_0),.din(w_dff_A_nc2zuewP2_0),.clk(gclk));
	jdff dff_A_fEJYJaC64_0(.dout(w_dff_A_Bqrd55ic6_0),.din(w_dff_A_fEJYJaC64_0),.clk(gclk));
	jdff dff_A_Bqrd55ic6_0(.dout(w_dff_A_6pg4YxwW2_0),.din(w_dff_A_Bqrd55ic6_0),.clk(gclk));
	jdff dff_A_6pg4YxwW2_0(.dout(w_dff_A_JFg8rEiJ6_0),.din(w_dff_A_6pg4YxwW2_0),.clk(gclk));
	jdff dff_A_JFg8rEiJ6_0(.dout(w_dff_A_OcCMQ68y4_0),.din(w_dff_A_JFg8rEiJ6_0),.clk(gclk));
	jdff dff_A_OcCMQ68y4_0(.dout(w_dff_A_pUlb9P5P1_0),.din(w_dff_A_OcCMQ68y4_0),.clk(gclk));
	jdff dff_A_pUlb9P5P1_0(.dout(w_dff_A_wSkeehsm1_0),.din(w_dff_A_pUlb9P5P1_0),.clk(gclk));
	jdff dff_A_wSkeehsm1_0(.dout(w_dff_A_Ly7xUSq95_0),.din(w_dff_A_wSkeehsm1_0),.clk(gclk));
	jdff dff_A_Ly7xUSq95_0(.dout(w_dff_A_r8yX35OL0_0),.din(w_dff_A_Ly7xUSq95_0),.clk(gclk));
	jdff dff_A_r8yX35OL0_0(.dout(w_dff_A_OvuI36Xm3_0),.din(w_dff_A_r8yX35OL0_0),.clk(gclk));
	jdff dff_A_OvuI36Xm3_0(.dout(w_dff_A_b4esieFH2_0),.din(w_dff_A_OvuI36Xm3_0),.clk(gclk));
	jdff dff_A_b4esieFH2_0(.dout(w_dff_A_rGQ9rEbx1_0),.din(w_dff_A_b4esieFH2_0),.clk(gclk));
	jdff dff_A_rGQ9rEbx1_0(.dout(w_dff_A_bA3xXtm41_0),.din(w_dff_A_rGQ9rEbx1_0),.clk(gclk));
	jdff dff_A_bA3xXtm41_0(.dout(w_dff_A_fqNnckpX0_0),.din(w_dff_A_bA3xXtm41_0),.clk(gclk));
	jdff dff_A_fqNnckpX0_0(.dout(G394),.din(w_dff_A_fqNnckpX0_0),.clk(gclk));
	jdff dff_A_vEddeJa75_2(.dout(w_dff_A_vmdaJfph6_0),.din(w_dff_A_vEddeJa75_2),.clk(gclk));
	jdff dff_A_vmdaJfph6_0(.dout(w_dff_A_FMvSAZ0R2_0),.din(w_dff_A_vmdaJfph6_0),.clk(gclk));
	jdff dff_A_FMvSAZ0R2_0(.dout(w_dff_A_iLpUerIY1_0),.din(w_dff_A_FMvSAZ0R2_0),.clk(gclk));
	jdff dff_A_iLpUerIY1_0(.dout(w_dff_A_ZUoOI0BO5_0),.din(w_dff_A_iLpUerIY1_0),.clk(gclk));
	jdff dff_A_ZUoOI0BO5_0(.dout(w_dff_A_VYie8oKZ4_0),.din(w_dff_A_ZUoOI0BO5_0),.clk(gclk));
	jdff dff_A_VYie8oKZ4_0(.dout(w_dff_A_D8skds636_0),.din(w_dff_A_VYie8oKZ4_0),.clk(gclk));
	jdff dff_A_D8skds636_0(.dout(w_dff_A_GNuP6mjp8_0),.din(w_dff_A_D8skds636_0),.clk(gclk));
	jdff dff_A_GNuP6mjp8_0(.dout(w_dff_A_z1gzQNb06_0),.din(w_dff_A_GNuP6mjp8_0),.clk(gclk));
	jdff dff_A_z1gzQNb06_0(.dout(w_dff_A_OSTDsA4W7_0),.din(w_dff_A_z1gzQNb06_0),.clk(gclk));
	jdff dff_A_OSTDsA4W7_0(.dout(w_dff_A_3WbuAF9l4_0),.din(w_dff_A_OSTDsA4W7_0),.clk(gclk));
	jdff dff_A_3WbuAF9l4_0(.dout(w_dff_A_xfZCYeKO1_0),.din(w_dff_A_3WbuAF9l4_0),.clk(gclk));
	jdff dff_A_xfZCYeKO1_0(.dout(w_dff_A_yg8BF1l82_0),.din(w_dff_A_xfZCYeKO1_0),.clk(gclk));
	jdff dff_A_yg8BF1l82_0(.dout(w_dff_A_wXGwjV8M1_0),.din(w_dff_A_yg8BF1l82_0),.clk(gclk));
	jdff dff_A_wXGwjV8M1_0(.dout(w_dff_A_4J9jGk8k2_0),.din(w_dff_A_wXGwjV8M1_0),.clk(gclk));
	jdff dff_A_4J9jGk8k2_0(.dout(w_dff_A_nYIGNC6q8_0),.din(w_dff_A_4J9jGk8k2_0),.clk(gclk));
	jdff dff_A_nYIGNC6q8_0(.dout(w_dff_A_paqg3lvO4_0),.din(w_dff_A_nYIGNC6q8_0),.clk(gclk));
	jdff dff_A_paqg3lvO4_0(.dout(w_dff_A_STpoYxwp4_0),.din(w_dff_A_paqg3lvO4_0),.clk(gclk));
	jdff dff_A_STpoYxwp4_0(.dout(w_dff_A_2FJp0xsN4_0),.din(w_dff_A_STpoYxwp4_0),.clk(gclk));
	jdff dff_A_2FJp0xsN4_0(.dout(G397),.din(w_dff_A_2FJp0xsN4_0),.clk(gclk));
	jdff dff_A_KMCbaGeF1_2(.dout(w_dff_A_q36PlStj3_0),.din(w_dff_A_KMCbaGeF1_2),.clk(gclk));
	jdff dff_A_q36PlStj3_0(.dout(w_dff_A_dBqpDcpe0_0),.din(w_dff_A_q36PlStj3_0),.clk(gclk));
	jdff dff_A_dBqpDcpe0_0(.dout(w_dff_A_hvDXOGaJ2_0),.din(w_dff_A_dBqpDcpe0_0),.clk(gclk));
	jdff dff_A_hvDXOGaJ2_0(.dout(w_dff_A_Qfzya5Ze6_0),.din(w_dff_A_hvDXOGaJ2_0),.clk(gclk));
	jdff dff_A_Qfzya5Ze6_0(.dout(w_dff_A_bv59T8UL8_0),.din(w_dff_A_Qfzya5Ze6_0),.clk(gclk));
	jdff dff_A_bv59T8UL8_0(.dout(w_dff_A_Gd6waxCM1_0),.din(w_dff_A_bv59T8UL8_0),.clk(gclk));
	jdff dff_A_Gd6waxCM1_0(.dout(w_dff_A_hMo2T9ni6_0),.din(w_dff_A_Gd6waxCM1_0),.clk(gclk));
	jdff dff_A_hMo2T9ni6_0(.dout(w_dff_A_IOOoSHDD5_0),.din(w_dff_A_hMo2T9ni6_0),.clk(gclk));
	jdff dff_A_IOOoSHDD5_0(.dout(w_dff_A_MJlkpX5O9_0),.din(w_dff_A_IOOoSHDD5_0),.clk(gclk));
	jdff dff_A_MJlkpX5O9_0(.dout(w_dff_A_MqYYqK3a1_0),.din(w_dff_A_MJlkpX5O9_0),.clk(gclk));
	jdff dff_A_MqYYqK3a1_0(.dout(w_dff_A_RuO7mcqB9_0),.din(w_dff_A_MqYYqK3a1_0),.clk(gclk));
	jdff dff_A_RuO7mcqB9_0(.dout(w_dff_A_dUxt6AWx7_0),.din(w_dff_A_RuO7mcqB9_0),.clk(gclk));
	jdff dff_A_dUxt6AWx7_0(.dout(G376),.din(w_dff_A_dUxt6AWx7_0),.clk(gclk));
	jdff dff_A_8VidLIuF6_2(.dout(w_dff_A_dnP6G8TY7_0),.din(w_dff_A_8VidLIuF6_2),.clk(gclk));
	jdff dff_A_dnP6G8TY7_0(.dout(w_dff_A_FmiXhclr4_0),.din(w_dff_A_dnP6G8TY7_0),.clk(gclk));
	jdff dff_A_FmiXhclr4_0(.dout(w_dff_A_OMstosv94_0),.din(w_dff_A_FmiXhclr4_0),.clk(gclk));
	jdff dff_A_OMstosv94_0(.dout(w_dff_A_vsPVKiou5_0),.din(w_dff_A_OMstosv94_0),.clk(gclk));
	jdff dff_A_vsPVKiou5_0(.dout(w_dff_A_1wUGljjO2_0),.din(w_dff_A_vsPVKiou5_0),.clk(gclk));
	jdff dff_A_1wUGljjO2_0(.dout(w_dff_A_rdtp5aFN2_0),.din(w_dff_A_1wUGljjO2_0),.clk(gclk));
	jdff dff_A_rdtp5aFN2_0(.dout(w_dff_A_p8pYFDhF7_0),.din(w_dff_A_rdtp5aFN2_0),.clk(gclk));
	jdff dff_A_p8pYFDhF7_0(.dout(w_dff_A_aXzsrJp07_0),.din(w_dff_A_p8pYFDhF7_0),.clk(gclk));
	jdff dff_A_aXzsrJp07_0(.dout(w_dff_A_0Bx1f9IE1_0),.din(w_dff_A_aXzsrJp07_0),.clk(gclk));
	jdff dff_A_0Bx1f9IE1_0(.dout(w_dff_A_I4jCtoFc9_0),.din(w_dff_A_0Bx1f9IE1_0),.clk(gclk));
	jdff dff_A_I4jCtoFc9_0(.dout(w_dff_A_57TMX5lc6_0),.din(w_dff_A_I4jCtoFc9_0),.clk(gclk));
	jdff dff_A_57TMX5lc6_0(.dout(w_dff_A_SJ3isSEu3_0),.din(w_dff_A_57TMX5lc6_0),.clk(gclk));
	jdff dff_A_SJ3isSEu3_0(.dout(w_dff_A_M1p3FErj9_0),.din(w_dff_A_SJ3isSEu3_0),.clk(gclk));
	jdff dff_A_M1p3FErj9_0(.dout(G379),.din(w_dff_A_M1p3FErj9_0),.clk(gclk));
	jdff dff_A_f3sHIXSK4_2(.dout(w_dff_A_9WmLhrWF7_0),.din(w_dff_A_f3sHIXSK4_2),.clk(gclk));
	jdff dff_A_9WmLhrWF7_0(.dout(w_dff_A_8nnZTuLO6_0),.din(w_dff_A_9WmLhrWF7_0),.clk(gclk));
	jdff dff_A_8nnZTuLO6_0(.dout(w_dff_A_ao8l4W4i3_0),.din(w_dff_A_8nnZTuLO6_0),.clk(gclk));
	jdff dff_A_ao8l4W4i3_0(.dout(w_dff_A_NdYWOdoP6_0),.din(w_dff_A_ao8l4W4i3_0),.clk(gclk));
	jdff dff_A_NdYWOdoP6_0(.dout(w_dff_A_SeZHf1mh4_0),.din(w_dff_A_NdYWOdoP6_0),.clk(gclk));
	jdff dff_A_SeZHf1mh4_0(.dout(w_dff_A_mVqDdQf03_0),.din(w_dff_A_SeZHf1mh4_0),.clk(gclk));
	jdff dff_A_mVqDdQf03_0(.dout(w_dff_A_Rz8PGoUa2_0),.din(w_dff_A_mVqDdQf03_0),.clk(gclk));
	jdff dff_A_Rz8PGoUa2_0(.dout(w_dff_A_MRYJka3J2_0),.din(w_dff_A_Rz8PGoUa2_0),.clk(gclk));
	jdff dff_A_MRYJka3J2_0(.dout(w_dff_A_Mzv24KvU8_0),.din(w_dff_A_MRYJka3J2_0),.clk(gclk));
	jdff dff_A_Mzv24KvU8_0(.dout(w_dff_A_BbYuBmPy4_0),.din(w_dff_A_Mzv24KvU8_0),.clk(gclk));
	jdff dff_A_BbYuBmPy4_0(.dout(w_dff_A_E0shbqX76_0),.din(w_dff_A_BbYuBmPy4_0),.clk(gclk));
	jdff dff_A_E0shbqX76_0(.dout(w_dff_A_MZeBBfbI7_0),.din(w_dff_A_E0shbqX76_0),.clk(gclk));
	jdff dff_A_MZeBBfbI7_0(.dout(w_dff_A_zOjJnjDn1_0),.din(w_dff_A_MZeBBfbI7_0),.clk(gclk));
	jdff dff_A_zOjJnjDn1_0(.dout(G382),.din(w_dff_A_zOjJnjDn1_0),.clk(gclk));
	jdff dff_A_H03IRAWS8_2(.dout(w_dff_A_NxRbqHJi1_0),.din(w_dff_A_H03IRAWS8_2),.clk(gclk));
	jdff dff_A_NxRbqHJi1_0(.dout(w_dff_A_kn56FF7D5_0),.din(w_dff_A_NxRbqHJi1_0),.clk(gclk));
	jdff dff_A_kn56FF7D5_0(.dout(w_dff_A_Do8OgmES8_0),.din(w_dff_A_kn56FF7D5_0),.clk(gclk));
	jdff dff_A_Do8OgmES8_0(.dout(w_dff_A_507IISw87_0),.din(w_dff_A_Do8OgmES8_0),.clk(gclk));
	jdff dff_A_507IISw87_0(.dout(w_dff_A_19jiPMKQ0_0),.din(w_dff_A_507IISw87_0),.clk(gclk));
	jdff dff_A_19jiPMKQ0_0(.dout(w_dff_A_udbXHxti9_0),.din(w_dff_A_19jiPMKQ0_0),.clk(gclk));
	jdff dff_A_udbXHxti9_0(.dout(w_dff_A_wfrMokYK3_0),.din(w_dff_A_udbXHxti9_0),.clk(gclk));
	jdff dff_A_wfrMokYK3_0(.dout(w_dff_A_3oRT5DHU4_0),.din(w_dff_A_wfrMokYK3_0),.clk(gclk));
	jdff dff_A_3oRT5DHU4_0(.dout(w_dff_A_MmLIGxEI6_0),.din(w_dff_A_3oRT5DHU4_0),.clk(gclk));
	jdff dff_A_MmLIGxEI6_0(.dout(w_dff_A_kT2xvXs51_0),.din(w_dff_A_MmLIGxEI6_0),.clk(gclk));
	jdff dff_A_kT2xvXs51_0(.dout(w_dff_A_bwfAXsGr4_0),.din(w_dff_A_kT2xvXs51_0),.clk(gclk));
	jdff dff_A_bwfAXsGr4_0(.dout(w_dff_A_La0VcisY5_0),.din(w_dff_A_bwfAXsGr4_0),.clk(gclk));
	jdff dff_A_La0VcisY5_0(.dout(w_dff_A_DzVLEwtQ3_0),.din(w_dff_A_La0VcisY5_0),.clk(gclk));
	jdff dff_A_DzVLEwtQ3_0(.dout(w_dff_A_G4xBhRH19_0),.din(w_dff_A_DzVLEwtQ3_0),.clk(gclk));
	jdff dff_A_G4xBhRH19_0(.dout(w_dff_A_Z4ta4T7k2_0),.din(w_dff_A_G4xBhRH19_0),.clk(gclk));
	jdff dff_A_Z4ta4T7k2_0(.dout(G385),.din(w_dff_A_Z4ta4T7k2_0),.clk(gclk));
	jdff dff_A_wykqDbm08_1(.dout(w_dff_A_9zPqFGQz7_0),.din(w_dff_A_wykqDbm08_1),.clk(gclk));
	jdff dff_A_9zPqFGQz7_0(.dout(w_dff_A_wc9ihYAb6_0),.din(w_dff_A_9zPqFGQz7_0),.clk(gclk));
	jdff dff_A_wc9ihYAb6_0(.dout(w_dff_A_KSSYnzCg4_0),.din(w_dff_A_wc9ihYAb6_0),.clk(gclk));
	jdff dff_A_KSSYnzCg4_0(.dout(w_dff_A_JEMkHivD3_0),.din(w_dff_A_KSSYnzCg4_0),.clk(gclk));
	jdff dff_A_JEMkHivD3_0(.dout(w_dff_A_wwXYz9bQ8_0),.din(w_dff_A_JEMkHivD3_0),.clk(gclk));
	jdff dff_A_wwXYz9bQ8_0(.dout(w_dff_A_fJtPq6tq7_0),.din(w_dff_A_wwXYz9bQ8_0),.clk(gclk));
	jdff dff_A_fJtPq6tq7_0(.dout(w_dff_A_1EZv6f307_0),.din(w_dff_A_fJtPq6tq7_0),.clk(gclk));
	jdff dff_A_1EZv6f307_0(.dout(w_dff_A_W2Pe5qtY8_0),.din(w_dff_A_1EZv6f307_0),.clk(gclk));
	jdff dff_A_W2Pe5qtY8_0(.dout(w_dff_A_lpC5Yjxz4_0),.din(w_dff_A_W2Pe5qtY8_0),.clk(gclk));
	jdff dff_A_lpC5Yjxz4_0(.dout(w_dff_A_AXYOX6if8_0),.din(w_dff_A_lpC5Yjxz4_0),.clk(gclk));
	jdff dff_A_AXYOX6if8_0(.dout(w_dff_A_zoXH8DyH0_0),.din(w_dff_A_AXYOX6if8_0),.clk(gclk));
	jdff dff_A_zoXH8DyH0_0(.dout(w_dff_A_AYx6ANXW1_0),.din(w_dff_A_zoXH8DyH0_0),.clk(gclk));
	jdff dff_A_AYx6ANXW1_0(.dout(w_dff_A_bCsRiVss5_0),.din(w_dff_A_AYx6ANXW1_0),.clk(gclk));
	jdff dff_A_bCsRiVss5_0(.dout(w_dff_A_12cptL5E3_0),.din(w_dff_A_bCsRiVss5_0),.clk(gclk));
	jdff dff_A_12cptL5E3_0(.dout(w_dff_A_tgV96mPK7_0),.din(w_dff_A_12cptL5E3_0),.clk(gclk));
	jdff dff_A_tgV96mPK7_0(.dout(G412),.din(w_dff_A_tgV96mPK7_0),.clk(gclk));
	jdff dff_A_nyyEt9jd2_1(.dout(w_dff_A_pkJ0GkZQ3_0),.din(w_dff_A_nyyEt9jd2_1),.clk(gclk));
	jdff dff_A_pkJ0GkZQ3_0(.dout(w_dff_A_trM5DOrX7_0),.din(w_dff_A_pkJ0GkZQ3_0),.clk(gclk));
	jdff dff_A_trM5DOrX7_0(.dout(w_dff_A_ZHXGwIji4_0),.din(w_dff_A_trM5DOrX7_0),.clk(gclk));
	jdff dff_A_ZHXGwIji4_0(.dout(w_dff_A_ydPQZw6P4_0),.din(w_dff_A_ZHXGwIji4_0),.clk(gclk));
	jdff dff_A_ydPQZw6P4_0(.dout(w_dff_A_KZ876fa08_0),.din(w_dff_A_ydPQZw6P4_0),.clk(gclk));
	jdff dff_A_KZ876fa08_0(.dout(w_dff_A_KCQfCrxM3_0),.din(w_dff_A_KZ876fa08_0),.clk(gclk));
	jdff dff_A_KCQfCrxM3_0(.dout(w_dff_A_8I9NFbmK2_0),.din(w_dff_A_KCQfCrxM3_0),.clk(gclk));
	jdff dff_A_8I9NFbmK2_0(.dout(w_dff_A_2VFTo9823_0),.din(w_dff_A_8I9NFbmK2_0),.clk(gclk));
	jdff dff_A_2VFTo9823_0(.dout(w_dff_A_f8kk55bC7_0),.din(w_dff_A_2VFTo9823_0),.clk(gclk));
	jdff dff_A_f8kk55bC7_0(.dout(w_dff_A_E0G0wta24_0),.din(w_dff_A_f8kk55bC7_0),.clk(gclk));
	jdff dff_A_E0G0wta24_0(.dout(w_dff_A_AJCzSzAi8_0),.din(w_dff_A_E0G0wta24_0),.clk(gclk));
	jdff dff_A_AJCzSzAi8_0(.dout(w_dff_A_uu30PPq45_0),.din(w_dff_A_AJCzSzAi8_0),.clk(gclk));
	jdff dff_A_uu30PPq45_0(.dout(w_dff_A_l36IXXuE2_0),.din(w_dff_A_uu30PPq45_0),.clk(gclk));
	jdff dff_A_l36IXXuE2_0(.dout(w_dff_A_7yOlvR0b9_0),.din(w_dff_A_l36IXXuE2_0),.clk(gclk));
	jdff dff_A_7yOlvR0b9_0(.dout(w_dff_A_cJ8tRCMf1_0),.din(w_dff_A_7yOlvR0b9_0),.clk(gclk));
	jdff dff_A_cJ8tRCMf1_0(.dout(G414),.din(w_dff_A_cJ8tRCMf1_0),.clk(gclk));
	jdff dff_A_5Phao2qY9_1(.dout(w_dff_A_SlpxzlWo9_0),.din(w_dff_A_5Phao2qY9_1),.clk(gclk));
	jdff dff_A_SlpxzlWo9_0(.dout(w_dff_A_IPLLeTBj4_0),.din(w_dff_A_SlpxzlWo9_0),.clk(gclk));
	jdff dff_A_IPLLeTBj4_0(.dout(w_dff_A_9HxK52q10_0),.din(w_dff_A_IPLLeTBj4_0),.clk(gclk));
	jdff dff_A_9HxK52q10_0(.dout(w_dff_A_ZIlnqiwe7_0),.din(w_dff_A_9HxK52q10_0),.clk(gclk));
	jdff dff_A_ZIlnqiwe7_0(.dout(w_dff_A_Y6Rgkjl59_0),.din(w_dff_A_ZIlnqiwe7_0),.clk(gclk));
	jdff dff_A_Y6Rgkjl59_0(.dout(w_dff_A_BLZDHSPz7_0),.din(w_dff_A_Y6Rgkjl59_0),.clk(gclk));
	jdff dff_A_BLZDHSPz7_0(.dout(w_dff_A_dtQrnXPr1_0),.din(w_dff_A_BLZDHSPz7_0),.clk(gclk));
	jdff dff_A_dtQrnXPr1_0(.dout(w_dff_A_xtdju5j15_0),.din(w_dff_A_dtQrnXPr1_0),.clk(gclk));
	jdff dff_A_xtdju5j15_0(.dout(w_dff_A_RUF0Bp9h5_0),.din(w_dff_A_xtdju5j15_0),.clk(gclk));
	jdff dff_A_RUF0Bp9h5_0(.dout(w_dff_A_gGKKYrL76_0),.din(w_dff_A_RUF0Bp9h5_0),.clk(gclk));
	jdff dff_A_gGKKYrL76_0(.dout(w_dff_A_eZsSL7no0_0),.din(w_dff_A_gGKKYrL76_0),.clk(gclk));
	jdff dff_A_eZsSL7no0_0(.dout(w_dff_A_JgCU2Fav8_0),.din(w_dff_A_eZsSL7no0_0),.clk(gclk));
	jdff dff_A_JgCU2Fav8_0(.dout(w_dff_A_IFN6ScqP4_0),.din(w_dff_A_JgCU2Fav8_0),.clk(gclk));
	jdff dff_A_IFN6ScqP4_0(.dout(G416),.din(w_dff_A_IFN6ScqP4_0),.clk(gclk));
	jdff dff_A_hMJWlTAb8_2(.dout(w_dff_A_7iyGzNrG8_0),.din(w_dff_A_hMJWlTAb8_2),.clk(gclk));
	jdff dff_A_7iyGzNrG8_0(.dout(w_dff_A_HRHixrIo2_0),.din(w_dff_A_7iyGzNrG8_0),.clk(gclk));
	jdff dff_A_HRHixrIo2_0(.dout(w_dff_A_IShvtZLt9_0),.din(w_dff_A_HRHixrIo2_0),.clk(gclk));
	jdff dff_A_IShvtZLt9_0(.dout(w_dff_A_AACjyD1C0_0),.din(w_dff_A_IShvtZLt9_0),.clk(gclk));
	jdff dff_A_AACjyD1C0_0(.dout(w_dff_A_dz6pocrP5_0),.din(w_dff_A_AACjyD1C0_0),.clk(gclk));
	jdff dff_A_dz6pocrP5_0(.dout(w_dff_A_oXOkdpwq9_0),.din(w_dff_A_dz6pocrP5_0),.clk(gclk));
	jdff dff_A_oXOkdpwq9_0(.dout(G249),.din(w_dff_A_oXOkdpwq9_0),.clk(gclk));
	jdff dff_A_k8fwsG6X8_2(.dout(w_dff_A_GI0MnWIo1_0),.din(w_dff_A_k8fwsG6X8_2),.clk(gclk));
	jdff dff_A_GI0MnWIo1_0(.dout(w_dff_A_Otjvdvdr9_0),.din(w_dff_A_GI0MnWIo1_0),.clk(gclk));
	jdff dff_A_Otjvdvdr9_0(.dout(w_dff_A_EZQyUxsP2_0),.din(w_dff_A_Otjvdvdr9_0),.clk(gclk));
	jdff dff_A_EZQyUxsP2_0(.dout(w_dff_A_e9EVMRV11_0),.din(w_dff_A_EZQyUxsP2_0),.clk(gclk));
	jdff dff_A_e9EVMRV11_0(.dout(w_dff_A_nvdRjiDF3_0),.din(w_dff_A_e9EVMRV11_0),.clk(gclk));
	jdff dff_A_nvdRjiDF3_0(.dout(w_dff_A_kdjx6fiP2_0),.din(w_dff_A_nvdRjiDF3_0),.clk(gclk));
	jdff dff_A_kdjx6fiP2_0(.dout(w_dff_A_r89USscb9_0),.din(w_dff_A_kdjx6fiP2_0),.clk(gclk));
	jdff dff_A_r89USscb9_0(.dout(w_dff_A_6if8DXLV5_0),.din(w_dff_A_r89USscb9_0),.clk(gclk));
	jdff dff_A_6if8DXLV5_0(.dout(w_dff_A_ncsEIN7l2_0),.din(w_dff_A_6if8DXLV5_0),.clk(gclk));
	jdff dff_A_ncsEIN7l2_0(.dout(G295),.din(w_dff_A_ncsEIN7l2_0),.clk(gclk));
	jdff dff_A_ouDDPZkR1_2(.dout(w_dff_A_I97Xg4N51_0),.din(w_dff_A_ouDDPZkR1_2),.clk(gclk));
	jdff dff_A_I97Xg4N51_0(.dout(w_dff_A_zYoIwaxo4_0),.din(w_dff_A_I97Xg4N51_0),.clk(gclk));
	jdff dff_A_zYoIwaxo4_0(.dout(w_dff_A_Cle7SSIO7_0),.din(w_dff_A_zYoIwaxo4_0),.clk(gclk));
	jdff dff_A_Cle7SSIO7_0(.dout(w_dff_A_rf51OD4G6_0),.din(w_dff_A_Cle7SSIO7_0),.clk(gclk));
	jdff dff_A_rf51OD4G6_0(.dout(w_dff_A_6x2DiZCh2_0),.din(w_dff_A_rf51OD4G6_0),.clk(gclk));
	jdff dff_A_6x2DiZCh2_0(.dout(G324),.din(w_dff_A_6x2DiZCh2_0),.clk(gclk));
	jdff dff_A_y1lICjJJ6_2(.dout(w_dff_A_xV6enaR67_0),.din(w_dff_A_y1lICjJJ6_2),.clk(gclk));
	jdff dff_A_xV6enaR67_0(.dout(w_dff_A_aYv5HA7j9_0),.din(w_dff_A_xV6enaR67_0),.clk(gclk));
	jdff dff_A_aYv5HA7j9_0(.dout(w_dff_A_V1Y6LPsY3_0),.din(w_dff_A_aYv5HA7j9_0),.clk(gclk));
	jdff dff_A_V1Y6LPsY3_0(.dout(w_dff_A_Uy4DScXa9_0),.din(w_dff_A_V1Y6LPsY3_0),.clk(gclk));
	jdff dff_A_Uy4DScXa9_0(.dout(w_dff_A_r0NcR0A47_0),.din(w_dff_A_Uy4DScXa9_0),.clk(gclk));
	jdff dff_A_r0NcR0A47_0(.dout(w_dff_A_lgpTcbSX8_0),.din(w_dff_A_r0NcR0A47_0),.clk(gclk));
	jdff dff_A_lgpTcbSX8_0(.dout(w_dff_A_jsap1kaJ3_0),.din(w_dff_A_lgpTcbSX8_0),.clk(gclk));
	jdff dff_A_jsap1kaJ3_0(.dout(w_dff_A_Tsmut07i4_0),.din(w_dff_A_jsap1kaJ3_0),.clk(gclk));
	jdff dff_A_Tsmut07i4_0(.dout(w_dff_A_NfzkrZUl7_0),.din(w_dff_A_Tsmut07i4_0),.clk(gclk));
	jdff dff_A_NfzkrZUl7_0(.dout(G252),.din(w_dff_A_NfzkrZUl7_0),.clk(gclk));
	jdff dff_A_kfLFkw6M5_2(.dout(G276),.din(w_dff_A_kfLFkw6M5_2),.clk(gclk));
	jdff dff_A_ACqslBCv7_2(.dout(w_dff_A_Y4t8sdBm8_0),.din(w_dff_A_ACqslBCv7_2),.clk(gclk));
	jdff dff_A_Y4t8sdBm8_0(.dout(w_dff_A_kifR7LAe6_0),.din(w_dff_A_Y4t8sdBm8_0),.clk(gclk));
	jdff dff_A_kifR7LAe6_0(.dout(w_dff_A_uw9UyzKk2_0),.din(w_dff_A_kifR7LAe6_0),.clk(gclk));
	jdff dff_A_uw9UyzKk2_0(.dout(w_dff_A_Bo9l5qom6_0),.din(w_dff_A_uw9UyzKk2_0),.clk(gclk));
	jdff dff_A_Bo9l5qom6_0(.dout(w_dff_A_pHtuYwCX5_0),.din(w_dff_A_Bo9l5qom6_0),.clk(gclk));
	jdff dff_A_pHtuYwCX5_0(.dout(G310),.din(w_dff_A_pHtuYwCX5_0),.clk(gclk));
	jdff dff_A_u94kLzpL1_2(.dout(w_dff_A_7l6AgJFW3_0),.din(w_dff_A_u94kLzpL1_2),.clk(gclk));
	jdff dff_A_7l6AgJFW3_0(.dout(w_dff_A_ruIjEfsc5_0),.din(w_dff_A_7l6AgJFW3_0),.clk(gclk));
	jdff dff_A_ruIjEfsc5_0(.dout(w_dff_A_eGCBi7UI3_0),.din(w_dff_A_ruIjEfsc5_0),.clk(gclk));
	jdff dff_A_eGCBi7UI3_0(.dout(w_dff_A_IMsKFPMu0_0),.din(w_dff_A_eGCBi7UI3_0),.clk(gclk));
	jdff dff_A_IMsKFPMu0_0(.dout(w_dff_A_BkSUfK953_0),.din(w_dff_A_IMsKFPMu0_0),.clk(gclk));
	jdff dff_A_BkSUfK953_0(.dout(w_dff_A_S7sW2fzJ2_0),.din(w_dff_A_BkSUfK953_0),.clk(gclk));
	jdff dff_A_S7sW2fzJ2_0(.dout(G313),.din(w_dff_A_S7sW2fzJ2_0),.clk(gclk));
	jdff dff_A_iJCHvIYW2_2(.dout(w_dff_A_DwVU4p0z8_0),.din(w_dff_A_iJCHvIYW2_2),.clk(gclk));
	jdff dff_A_DwVU4p0z8_0(.dout(w_dff_A_RxdP6a0E7_0),.din(w_dff_A_DwVU4p0z8_0),.clk(gclk));
	jdff dff_A_RxdP6a0E7_0(.dout(w_dff_A_t5Uihtn31_0),.din(w_dff_A_RxdP6a0E7_0),.clk(gclk));
	jdff dff_A_t5Uihtn31_0(.dout(w_dff_A_THjpltkp3_0),.din(w_dff_A_t5Uihtn31_0),.clk(gclk));
	jdff dff_A_THjpltkp3_0(.dout(w_dff_A_a5BYp71V9_0),.din(w_dff_A_THjpltkp3_0),.clk(gclk));
	jdff dff_A_a5BYp71V9_0(.dout(w_dff_A_eKNM7vN50_0),.din(w_dff_A_a5BYp71V9_0),.clk(gclk));
	jdff dff_A_eKNM7vN50_0(.dout(w_dff_A_7WMxIowz2_0),.din(w_dff_A_eKNM7vN50_0),.clk(gclk));
	jdff dff_A_7WMxIowz2_0(.dout(G316),.din(w_dff_A_7WMxIowz2_0),.clk(gclk));
	jdff dff_A_IhK2kk8i6_2(.dout(w_dff_A_KDAv0QYT0_0),.din(w_dff_A_IhK2kk8i6_2),.clk(gclk));
	jdff dff_A_KDAv0QYT0_0(.dout(w_dff_A_j0C65L6g2_0),.din(w_dff_A_KDAv0QYT0_0),.clk(gclk));
	jdff dff_A_j0C65L6g2_0(.dout(w_dff_A_aVSyyIGQ5_0),.din(w_dff_A_j0C65L6g2_0),.clk(gclk));
	jdff dff_A_aVSyyIGQ5_0(.dout(w_dff_A_4AYGEmap7_0),.din(w_dff_A_aVSyyIGQ5_0),.clk(gclk));
	jdff dff_A_4AYGEmap7_0(.dout(w_dff_A_xI4IW2bo6_0),.din(w_dff_A_4AYGEmap7_0),.clk(gclk));
	jdff dff_A_xI4IW2bo6_0(.dout(w_dff_A_h8Q04HCz0_0),.din(w_dff_A_xI4IW2bo6_0),.clk(gclk));
	jdff dff_A_h8Q04HCz0_0(.dout(w_dff_A_yZTlQUTQ7_0),.din(w_dff_A_h8Q04HCz0_0),.clk(gclk));
	jdff dff_A_yZTlQUTQ7_0(.dout(G319),.din(w_dff_A_yZTlQUTQ7_0),.clk(gclk));
	jdff dff_A_IyoCa8wx8_2(.dout(w_dff_A_NvrgdMKU2_0),.din(w_dff_A_IyoCa8wx8_2),.clk(gclk));
	jdff dff_A_NvrgdMKU2_0(.dout(G327),.din(w_dff_A_NvrgdMKU2_0),.clk(gclk));
	jdff dff_A_HUfgb5F17_2(.dout(w_dff_A_WZFDRTZ02_0),.din(w_dff_A_HUfgb5F17_2),.clk(gclk));
	jdff dff_A_WZFDRTZ02_0(.dout(w_dff_A_UgHHmDTh0_0),.din(w_dff_A_WZFDRTZ02_0),.clk(gclk));
	jdff dff_A_UgHHmDTh0_0(.dout(G330),.din(w_dff_A_UgHHmDTh0_0),.clk(gclk));
	jdff dff_A_56MDtBHq7_2(.dout(w_dff_A_YMbsQHww3_0),.din(w_dff_A_56MDtBHq7_2),.clk(gclk));
	jdff dff_A_YMbsQHww3_0(.dout(w_dff_A_eoKninLD1_0),.din(w_dff_A_YMbsQHww3_0),.clk(gclk));
	jdff dff_A_eoKninLD1_0(.dout(w_dff_A_jVNl1AUr1_0),.din(w_dff_A_eoKninLD1_0),.clk(gclk));
	jdff dff_A_jVNl1AUr1_0(.dout(G333),.din(w_dff_A_jVNl1AUr1_0),.clk(gclk));
	jdff dff_A_bmy2DIyV3_2(.dout(w_dff_A_DmiOXxqU7_0),.din(w_dff_A_bmy2DIyV3_2),.clk(gclk));
	jdff dff_A_DmiOXxqU7_0(.dout(w_dff_A_MrFmcRjM9_0),.din(w_dff_A_DmiOXxqU7_0),.clk(gclk));
	jdff dff_A_MrFmcRjM9_0(.dout(w_dff_A_Faa1tfed9_0),.din(w_dff_A_MrFmcRjM9_0),.clk(gclk));
	jdff dff_A_Faa1tfed9_0(.dout(G336),.din(w_dff_A_Faa1tfed9_0),.clk(gclk));
	jdff dff_A_jhWvCLTd0_2(.dout(w_dff_A_DOhhlZFY7_0),.din(w_dff_A_jhWvCLTd0_2),.clk(gclk));
	jdff dff_A_DOhhlZFY7_0(.dout(w_dff_A_IydLM9Go8_0),.din(w_dff_A_DOhhlZFY7_0),.clk(gclk));
	jdff dff_A_IydLM9Go8_0(.dout(w_dff_A_r7pMVeiv4_0),.din(w_dff_A_IydLM9Go8_0),.clk(gclk));
	jdff dff_A_r7pMVeiv4_0(.dout(w_dff_A_W32TXfhs9_0),.din(w_dff_A_r7pMVeiv4_0),.clk(gclk));
	jdff dff_A_W32TXfhs9_0(.dout(w_dff_A_89CIiKXN0_0),.din(w_dff_A_W32TXfhs9_0),.clk(gclk));
	jdff dff_A_89CIiKXN0_0(.dout(w_dff_A_yTIIXXdG2_0),.din(w_dff_A_89CIiKXN0_0),.clk(gclk));
	jdff dff_A_yTIIXXdG2_0(.dout(w_dff_A_n4QvVDPh2_0),.din(w_dff_A_yTIIXXdG2_0),.clk(gclk));
	jdff dff_A_n4QvVDPh2_0(.dout(w_dff_A_DmSxY9v33_0),.din(w_dff_A_n4QvVDPh2_0),.clk(gclk));
	jdff dff_A_DmSxY9v33_0(.dout(w_dff_A_JZZMLKg54_0),.din(w_dff_A_DmSxY9v33_0),.clk(gclk));
	jdff dff_A_JZZMLKg54_0(.dout(w_dff_A_mmQlEfuy6_0),.din(w_dff_A_JZZMLKg54_0),.clk(gclk));
	jdff dff_A_mmQlEfuy6_0(.dout(w_dff_A_8zlm28G46_0),.din(w_dff_A_mmQlEfuy6_0),.clk(gclk));
	jdff dff_A_8zlm28G46_0(.dout(G418),.din(w_dff_A_8zlm28G46_0),.clk(gclk));
	jdff dff_A_FoWZznBm6_2(.dout(G273),.din(w_dff_A_FoWZznBm6_2),.clk(gclk));
	jdff dff_A_bXHu9UF51_2(.dout(w_dff_A_Yexk4taD4_0),.din(w_dff_A_bXHu9UF51_2),.clk(gclk));
	jdff dff_A_Yexk4taD4_0(.dout(w_dff_A_9IN6LYZ30_0),.din(w_dff_A_Yexk4taD4_0),.clk(gclk));
	jdff dff_A_9IN6LYZ30_0(.dout(w_dff_A_3ubhS1Ve3_0),.din(w_dff_A_9IN6LYZ30_0),.clk(gclk));
	jdff dff_A_3ubhS1Ve3_0(.dout(G298),.din(w_dff_A_3ubhS1Ve3_0),.clk(gclk));
	jdff dff_A_kO1eFYA95_2(.dout(w_dff_A_KvSYlQtB0_0),.din(w_dff_A_kO1eFYA95_2),.clk(gclk));
	jdff dff_A_KvSYlQtB0_0(.dout(w_dff_A_2e7Pzvlt4_0),.din(w_dff_A_KvSYlQtB0_0),.clk(gclk));
	jdff dff_A_2e7Pzvlt4_0(.dout(w_dff_A_wI0jkKM02_0),.din(w_dff_A_2e7Pzvlt4_0),.clk(gclk));
	jdff dff_A_wI0jkKM02_0(.dout(w_dff_A_pq520oT52_0),.din(w_dff_A_wI0jkKM02_0),.clk(gclk));
	jdff dff_A_pq520oT52_0(.dout(w_dff_A_FQeftoZR1_0),.din(w_dff_A_pq520oT52_0),.clk(gclk));
	jdff dff_A_FQeftoZR1_0(.dout(G301),.din(w_dff_A_FQeftoZR1_0),.clk(gclk));
	jdff dff_A_QNPL4Nn99_2(.dout(w_dff_A_eF8HMsmM0_0),.din(w_dff_A_QNPL4Nn99_2),.clk(gclk));
	jdff dff_A_eF8HMsmM0_0(.dout(w_dff_A_nVo2cKWp6_0),.din(w_dff_A_eF8HMsmM0_0),.clk(gclk));
	jdff dff_A_nVo2cKWp6_0(.dout(w_dff_A_wMRy0g015_0),.din(w_dff_A_nVo2cKWp6_0),.clk(gclk));
	jdff dff_A_wMRy0g015_0(.dout(w_dff_A_JqoY9hF47_0),.din(w_dff_A_wMRy0g015_0),.clk(gclk));
	jdff dff_A_JqoY9hF47_0(.dout(w_dff_A_15EPoaaV9_0),.din(w_dff_A_JqoY9hF47_0),.clk(gclk));
	jdff dff_A_15EPoaaV9_0(.dout(G304),.din(w_dff_A_15EPoaaV9_0),.clk(gclk));
	jdff dff_A_GtDw502C2_2(.dout(w_dff_A_idBcVgJA1_0),.din(w_dff_A_GtDw502C2_2),.clk(gclk));
	jdff dff_A_idBcVgJA1_0(.dout(w_dff_A_QW7ti7wh7_0),.din(w_dff_A_idBcVgJA1_0),.clk(gclk));
	jdff dff_A_QW7ti7wh7_0(.dout(w_dff_A_F74uv20G6_0),.din(w_dff_A_QW7ti7wh7_0),.clk(gclk));
	jdff dff_A_F74uv20G6_0(.dout(w_dff_A_4at4GPYc7_0),.din(w_dff_A_F74uv20G6_0),.clk(gclk));
	jdff dff_A_4at4GPYc7_0(.dout(w_dff_A_gmPvQ6Lp0_0),.din(w_dff_A_4at4GPYc7_0),.clk(gclk));
	jdff dff_A_gmPvQ6Lp0_0(.dout(w_dff_A_7tF7lrrX4_0),.din(w_dff_A_gmPvQ6Lp0_0),.clk(gclk));
	jdff dff_A_7tF7lrrX4_0(.dout(w_dff_A_CLY8YUQh0_0),.din(w_dff_A_7tF7lrrX4_0),.clk(gclk));
	jdff dff_A_CLY8YUQh0_0(.dout(G307),.din(w_dff_A_CLY8YUQh0_0),.clk(gclk));
	jdff dff_A_u2VS0eu85_2(.dout(w_dff_A_0WEmXAVP9_0),.din(w_dff_A_u2VS0eu85_2),.clk(gclk));
	jdff dff_A_0WEmXAVP9_0(.dout(w_dff_A_AmHEvaNU2_0),.din(w_dff_A_0WEmXAVP9_0),.clk(gclk));
	jdff dff_A_AmHEvaNU2_0(.dout(w_dff_A_DVNHGDkx9_0),.din(w_dff_A_AmHEvaNU2_0),.clk(gclk));
	jdff dff_A_DVNHGDkx9_0(.dout(w_dff_A_PZYJlCxG8_0),.din(w_dff_A_DVNHGDkx9_0),.clk(gclk));
	jdff dff_A_PZYJlCxG8_0(.dout(w_dff_A_hgG319v29_0),.din(w_dff_A_PZYJlCxG8_0),.clk(gclk));
	jdff dff_A_hgG319v29_0(.dout(w_dff_A_XGIEQCg10_0),.din(w_dff_A_hgG319v29_0),.clk(gclk));
	jdff dff_A_XGIEQCg10_0(.dout(w_dff_A_SpyAcNEH9_0),.din(w_dff_A_XGIEQCg10_0),.clk(gclk));
	jdff dff_A_SpyAcNEH9_0(.dout(w_dff_A_nRWXLRke4_0),.din(w_dff_A_SpyAcNEH9_0),.clk(gclk));
	jdff dff_A_nRWXLRke4_0(.dout(w_dff_A_r2jAo6Mu9_0),.din(w_dff_A_nRWXLRke4_0),.clk(gclk));
	jdff dff_A_r2jAo6Mu9_0(.dout(w_dff_A_vN0bMFAx7_0),.din(w_dff_A_r2jAo6Mu9_0),.clk(gclk));
	jdff dff_A_vN0bMFAx7_0(.dout(w_dff_A_dGxuGP4h3_0),.din(w_dff_A_vN0bMFAx7_0),.clk(gclk));
	jdff dff_A_dGxuGP4h3_0(.dout(w_dff_A_dflpMAFK7_0),.din(w_dff_A_dGxuGP4h3_0),.clk(gclk));
	jdff dff_A_dflpMAFK7_0(.dout(w_dff_A_d63CencI3_0),.din(w_dff_A_dflpMAFK7_0),.clk(gclk));
	jdff dff_A_d63CencI3_0(.dout(G344),.din(w_dff_A_d63CencI3_0),.clk(gclk));
	jdff dff_A_u8189vHk1_2(.dout(G422),.din(w_dff_A_u8189vHk1_2),.clk(gclk));
	jdff dff_A_KJykaV3M0_2(.dout(G469),.din(w_dff_A_KJykaV3M0_2),.clk(gclk));
	jdff dff_A_pN6IxNGh5_2(.dout(w_dff_A_TeChXTMa7_0),.din(w_dff_A_pN6IxNGh5_2),.clk(gclk));
	jdff dff_A_TeChXTMa7_0(.dout(w_dff_A_ikIdkQUw3_0),.din(w_dff_A_TeChXTMa7_0),.clk(gclk));
	jdff dff_A_ikIdkQUw3_0(.dout(w_dff_A_EoeqTSWy8_0),.din(w_dff_A_ikIdkQUw3_0),.clk(gclk));
	jdff dff_A_EoeqTSWy8_0(.dout(G419),.din(w_dff_A_EoeqTSWy8_0),.clk(gclk));
	jdff dff_A_E8jalRTs2_2(.dout(w_dff_A_wfUaDLW66_0),.din(w_dff_A_E8jalRTs2_2),.clk(gclk));
	jdff dff_A_wfUaDLW66_0(.dout(w_dff_A_arKIhtye4_0),.din(w_dff_A_wfUaDLW66_0),.clk(gclk));
	jdff dff_A_arKIhtye4_0(.dout(w_dff_A_QzOwvaFh3_0),.din(w_dff_A_arKIhtye4_0),.clk(gclk));
	jdff dff_A_QzOwvaFh3_0(.dout(G471),.din(w_dff_A_QzOwvaFh3_0),.clk(gclk));
	jdff dff_A_Qutbbi7W3_2(.dout(w_dff_A_j9wtRz0k2_0),.din(w_dff_A_Qutbbi7W3_2),.clk(gclk));
	jdff dff_A_j9wtRz0k2_0(.dout(w_dff_A_zB9ZqTqK2_0),.din(w_dff_A_j9wtRz0k2_0),.clk(gclk));
	jdff dff_A_zB9ZqTqK2_0(.dout(w_dff_A_bwLEuQlq6_0),.din(w_dff_A_zB9ZqTqK2_0),.clk(gclk));
	jdff dff_A_bwLEuQlq6_0(.dout(w_dff_A_U7c5MoiX0_0),.din(w_dff_A_bwLEuQlq6_0),.clk(gclk));
	jdff dff_A_U7c5MoiX0_0(.dout(w_dff_A_gi4w7YCi8_0),.din(w_dff_A_U7c5MoiX0_0),.clk(gclk));
	jdff dff_A_gi4w7YCi8_0(.dout(w_dff_A_J5yOHCRL9_0),.din(w_dff_A_gi4w7YCi8_0),.clk(gclk));
	jdff dff_A_J5yOHCRL9_0(.dout(w_dff_A_i45KJBzy6_0),.din(w_dff_A_J5yOHCRL9_0),.clk(gclk));
	jdff dff_A_i45KJBzy6_0(.dout(w_dff_A_AQx62qQL1_0),.din(w_dff_A_i45KJBzy6_0),.clk(gclk));
	jdff dff_A_AQx62qQL1_0(.dout(w_dff_A_Xe1ad79S1_0),.din(w_dff_A_AQx62qQL1_0),.clk(gclk));
	jdff dff_A_Xe1ad79S1_0(.dout(G359),.din(w_dff_A_Xe1ad79S1_0),.clk(gclk));
	jdff dff_A_QxgVD2QB2_2(.dout(w_dff_A_zgWesmuJ1_0),.din(w_dff_A_QxgVD2QB2_2),.clk(gclk));
	jdff dff_A_zgWesmuJ1_0(.dout(w_dff_A_aaoXjhMP0_0),.din(w_dff_A_zgWesmuJ1_0),.clk(gclk));
	jdff dff_A_aaoXjhMP0_0(.dout(w_dff_A_FiiC9BSW1_0),.din(w_dff_A_aaoXjhMP0_0),.clk(gclk));
	jdff dff_A_FiiC9BSW1_0(.dout(w_dff_A_m5y08wEu6_0),.din(w_dff_A_FiiC9BSW1_0),.clk(gclk));
	jdff dff_A_m5y08wEu6_0(.dout(w_dff_A_5dlFzehl4_0),.din(w_dff_A_m5y08wEu6_0),.clk(gclk));
	jdff dff_A_5dlFzehl4_0(.dout(w_dff_A_HRaAPMWW8_0),.din(w_dff_A_5dlFzehl4_0),.clk(gclk));
	jdff dff_A_HRaAPMWW8_0(.dout(w_dff_A_z4W1hAW05_0),.din(w_dff_A_HRaAPMWW8_0),.clk(gclk));
	jdff dff_A_z4W1hAW05_0(.dout(w_dff_A_SphUPevv8_0),.din(w_dff_A_z4W1hAW05_0),.clk(gclk));
	jdff dff_A_SphUPevv8_0(.dout(w_dff_A_dqPJ984U6_0),.din(w_dff_A_SphUPevv8_0),.clk(gclk));
	jdff dff_A_dqPJ984U6_0(.dout(w_dff_A_6FJsb1lw2_0),.din(w_dff_A_dqPJ984U6_0),.clk(gclk));
	jdff dff_A_6FJsb1lw2_0(.dout(G362),.din(w_dff_A_6FJsb1lw2_0),.clk(gclk));
	jdff dff_A_OEN3E7xB2_2(.dout(w_dff_A_FBPSAZrq3_0),.din(w_dff_A_OEN3E7xB2_2),.clk(gclk));
	jdff dff_A_FBPSAZrq3_0(.dout(w_dff_A_73WPHF0a8_0),.din(w_dff_A_FBPSAZrq3_0),.clk(gclk));
	jdff dff_A_73WPHF0a8_0(.dout(w_dff_A_ugyj3iQ65_0),.din(w_dff_A_73WPHF0a8_0),.clk(gclk));
	jdff dff_A_ugyj3iQ65_0(.dout(w_dff_A_ZZ2Y7ZiW0_0),.din(w_dff_A_ugyj3iQ65_0),.clk(gclk));
	jdff dff_A_ZZ2Y7ZiW0_0(.dout(w_dff_A_EklCC1Fx2_0),.din(w_dff_A_ZZ2Y7ZiW0_0),.clk(gclk));
	jdff dff_A_EklCC1Fx2_0(.dout(w_dff_A_hdHDfOPH7_0),.din(w_dff_A_EklCC1Fx2_0),.clk(gclk));
	jdff dff_A_hdHDfOPH7_0(.dout(w_dff_A_Gb0kjhg59_0),.din(w_dff_A_hdHDfOPH7_0),.clk(gclk));
	jdff dff_A_Gb0kjhg59_0(.dout(w_dff_A_oQuZ9C3o7_0),.din(w_dff_A_Gb0kjhg59_0),.clk(gclk));
	jdff dff_A_oQuZ9C3o7_0(.dout(w_dff_A_HdHLYKd25_0),.din(w_dff_A_oQuZ9C3o7_0),.clk(gclk));
	jdff dff_A_HdHLYKd25_0(.dout(w_dff_A_4YZ7HJAB9_0),.din(w_dff_A_HdHLYKd25_0),.clk(gclk));
	jdff dff_A_4YZ7HJAB9_0(.dout(w_dff_A_LLUDcLli2_0),.din(w_dff_A_4YZ7HJAB9_0),.clk(gclk));
	jdff dff_A_LLUDcLli2_0(.dout(G365),.din(w_dff_A_LLUDcLli2_0),.clk(gclk));
	jdff dff_A_BRr7V1Dd0_2(.dout(w_dff_A_bTLj5nNy8_0),.din(w_dff_A_BRr7V1Dd0_2),.clk(gclk));
	jdff dff_A_bTLj5nNy8_0(.dout(w_dff_A_5waj8wW36_0),.din(w_dff_A_bTLj5nNy8_0),.clk(gclk));
	jdff dff_A_5waj8wW36_0(.dout(w_dff_A_RMkVxy4D8_0),.din(w_dff_A_5waj8wW36_0),.clk(gclk));
	jdff dff_A_RMkVxy4D8_0(.dout(w_dff_A_jVXSzJcQ9_0),.din(w_dff_A_RMkVxy4D8_0),.clk(gclk));
	jdff dff_A_jVXSzJcQ9_0(.dout(w_dff_A_AOsmoC2R4_0),.din(w_dff_A_jVXSzJcQ9_0),.clk(gclk));
	jdff dff_A_AOsmoC2R4_0(.dout(w_dff_A_3e1Lm0s86_0),.din(w_dff_A_AOsmoC2R4_0),.clk(gclk));
	jdff dff_A_3e1Lm0s86_0(.dout(w_dff_A_1HCHJbDg8_0),.din(w_dff_A_3e1Lm0s86_0),.clk(gclk));
	jdff dff_A_1HCHJbDg8_0(.dout(w_dff_A_0T8uOQtH3_0),.din(w_dff_A_1HCHJbDg8_0),.clk(gclk));
	jdff dff_A_0T8uOQtH3_0(.dout(w_dff_A_kJM8BYLq2_0),.din(w_dff_A_0T8uOQtH3_0),.clk(gclk));
	jdff dff_A_kJM8BYLq2_0(.dout(w_dff_A_cHjh7vKg0_0),.din(w_dff_A_kJM8BYLq2_0),.clk(gclk));
	jdff dff_A_cHjh7vKg0_0(.dout(w_dff_A_mPaS6Mha1_0),.din(w_dff_A_cHjh7vKg0_0),.clk(gclk));
	jdff dff_A_mPaS6Mha1_0(.dout(G368),.din(w_dff_A_mPaS6Mha1_0),.clk(gclk));
	jdff dff_A_VimgZs4n3_2(.dout(w_dff_A_3PbZ1Jbq8_0),.din(w_dff_A_VimgZs4n3_2),.clk(gclk));
	jdff dff_A_3PbZ1Jbq8_0(.dout(w_dff_A_zXS4Xfyi0_0),.din(w_dff_A_3PbZ1Jbq8_0),.clk(gclk));
	jdff dff_A_zXS4Xfyi0_0(.dout(w_dff_A_GRpvyfWq5_0),.din(w_dff_A_zXS4Xfyi0_0),.clk(gclk));
	jdff dff_A_GRpvyfWq5_0(.dout(w_dff_A_psKGp7Cq9_0),.din(w_dff_A_GRpvyfWq5_0),.clk(gclk));
	jdff dff_A_psKGp7Cq9_0(.dout(w_dff_A_lxkcQEtM0_0),.din(w_dff_A_psKGp7Cq9_0),.clk(gclk));
	jdff dff_A_lxkcQEtM0_0(.dout(w_dff_A_Q58gQSBR2_0),.din(w_dff_A_lxkcQEtM0_0),.clk(gclk));
	jdff dff_A_Q58gQSBR2_0(.dout(w_dff_A_ekUOwAko3_0),.din(w_dff_A_Q58gQSBR2_0),.clk(gclk));
	jdff dff_A_ekUOwAko3_0(.dout(w_dff_A_dx0HSNzG9_0),.din(w_dff_A_ekUOwAko3_0),.clk(gclk));
	jdff dff_A_dx0HSNzG9_0(.dout(G347),.din(w_dff_A_dx0HSNzG9_0),.clk(gclk));
	jdff dff_A_djG7tKrZ7_2(.dout(w_dff_A_ghteABgK6_0),.din(w_dff_A_djG7tKrZ7_2),.clk(gclk));
	jdff dff_A_ghteABgK6_0(.dout(w_dff_A_Ab0KCW1j2_0),.din(w_dff_A_ghteABgK6_0),.clk(gclk));
	jdff dff_A_Ab0KCW1j2_0(.dout(w_dff_A_pZELC5nk3_0),.din(w_dff_A_Ab0KCW1j2_0),.clk(gclk));
	jdff dff_A_pZELC5nk3_0(.dout(w_dff_A_9iZodpNr8_0),.din(w_dff_A_pZELC5nk3_0),.clk(gclk));
	jdff dff_A_9iZodpNr8_0(.dout(w_dff_A_IVFAHnMD3_0),.din(w_dff_A_9iZodpNr8_0),.clk(gclk));
	jdff dff_A_IVFAHnMD3_0(.dout(w_dff_A_VIktzUjc1_0),.din(w_dff_A_IVFAHnMD3_0),.clk(gclk));
	jdff dff_A_VIktzUjc1_0(.dout(w_dff_A_GjlOPqmp8_0),.din(w_dff_A_VIktzUjc1_0),.clk(gclk));
	jdff dff_A_GjlOPqmp8_0(.dout(w_dff_A_6Y8UhFqg3_0),.din(w_dff_A_GjlOPqmp8_0),.clk(gclk));
	jdff dff_A_6Y8UhFqg3_0(.dout(w_dff_A_CzzP5pjZ0_0),.din(w_dff_A_6Y8UhFqg3_0),.clk(gclk));
	jdff dff_A_CzzP5pjZ0_0(.dout(G350),.din(w_dff_A_CzzP5pjZ0_0),.clk(gclk));
	jdff dff_A_P8hPtzqU4_2(.dout(w_dff_A_9ybG1xG72_0),.din(w_dff_A_P8hPtzqU4_2),.clk(gclk));
	jdff dff_A_9ybG1xG72_0(.dout(w_dff_A_21VOdRlb4_0),.din(w_dff_A_9ybG1xG72_0),.clk(gclk));
	jdff dff_A_21VOdRlb4_0(.dout(w_dff_A_ALy7YhUb2_0),.din(w_dff_A_21VOdRlb4_0),.clk(gclk));
	jdff dff_A_ALy7YhUb2_0(.dout(w_dff_A_WrKJH55W6_0),.din(w_dff_A_ALy7YhUb2_0),.clk(gclk));
	jdff dff_A_WrKJH55W6_0(.dout(w_dff_A_ieoW1bNp6_0),.din(w_dff_A_WrKJH55W6_0),.clk(gclk));
	jdff dff_A_ieoW1bNp6_0(.dout(w_dff_A_ea7jBFts1_0),.din(w_dff_A_ieoW1bNp6_0),.clk(gclk));
	jdff dff_A_ea7jBFts1_0(.dout(w_dff_A_0iF253ta6_0),.din(w_dff_A_ea7jBFts1_0),.clk(gclk));
	jdff dff_A_0iF253ta6_0(.dout(w_dff_A_Z3sOWuaz0_0),.din(w_dff_A_0iF253ta6_0),.clk(gclk));
	jdff dff_A_Z3sOWuaz0_0(.dout(w_dff_A_rw5qINAa0_0),.din(w_dff_A_Z3sOWuaz0_0),.clk(gclk));
	jdff dff_A_rw5qINAa0_0(.dout(G353),.din(w_dff_A_rw5qINAa0_0),.clk(gclk));
	jdff dff_A_ypcAw9sg9_2(.dout(w_dff_A_mOswMUxg3_0),.din(w_dff_A_ypcAw9sg9_2),.clk(gclk));
	jdff dff_A_mOswMUxg3_0(.dout(w_dff_A_tIzFAeLt4_0),.din(w_dff_A_mOswMUxg3_0),.clk(gclk));
	jdff dff_A_tIzFAeLt4_0(.dout(w_dff_A_7BPlkgWi9_0),.din(w_dff_A_tIzFAeLt4_0),.clk(gclk));
	jdff dff_A_7BPlkgWi9_0(.dout(w_dff_A_dAgHZCA45_0),.din(w_dff_A_7BPlkgWi9_0),.clk(gclk));
	jdff dff_A_dAgHZCA45_0(.dout(w_dff_A_QWZOHusX0_0),.din(w_dff_A_dAgHZCA45_0),.clk(gclk));
	jdff dff_A_QWZOHusX0_0(.dout(w_dff_A_E1az6nZ82_0),.din(w_dff_A_QWZOHusX0_0),.clk(gclk));
	jdff dff_A_E1az6nZ82_0(.dout(w_dff_A_XiIHYqRH8_0),.din(w_dff_A_E1az6nZ82_0),.clk(gclk));
	jdff dff_A_XiIHYqRH8_0(.dout(w_dff_A_OsqvV3eo7_0),.din(w_dff_A_XiIHYqRH8_0),.clk(gclk));
	jdff dff_A_OsqvV3eo7_0(.dout(w_dff_A_38FS1zn56_0),.din(w_dff_A_OsqvV3eo7_0),.clk(gclk));
	jdff dff_A_38FS1zn56_0(.dout(w_dff_A_y6MjP8Qb8_0),.din(w_dff_A_38FS1zn56_0),.clk(gclk));
	jdff dff_A_y6MjP8Qb8_0(.dout(w_dff_A_nv0Y42PX8_0),.din(w_dff_A_y6MjP8Qb8_0),.clk(gclk));
	jdff dff_A_nv0Y42PX8_0(.dout(G356),.din(w_dff_A_nv0Y42PX8_0),.clk(gclk));
	jdff dff_A_O0ichDPW1_2(.dout(w_dff_A_PtgjT43b1_0),.din(w_dff_A_O0ichDPW1_2),.clk(gclk));
	jdff dff_A_PtgjT43b1_0(.dout(w_dff_A_IOZH2WS93_0),.din(w_dff_A_PtgjT43b1_0),.clk(gclk));
	jdff dff_A_IOZH2WS93_0(.dout(w_dff_A_jfawbR8f2_0),.din(w_dff_A_IOZH2WS93_0),.clk(gclk));
	jdff dff_A_jfawbR8f2_0(.dout(w_dff_A_LEzamXti6_0),.din(w_dff_A_jfawbR8f2_0),.clk(gclk));
	jdff dff_A_LEzamXti6_0(.dout(G321),.din(w_dff_A_LEzamXti6_0),.clk(gclk));
	jdff dff_A_p7vnaGTp4_2(.dout(w_dff_A_yDtmijmt8_0),.din(w_dff_A_p7vnaGTp4_2),.clk(gclk));
	jdff dff_A_yDtmijmt8_0(.dout(w_dff_A_5B511Ywc8_0),.din(w_dff_A_yDtmijmt8_0),.clk(gclk));
	jdff dff_A_5B511Ywc8_0(.dout(w_dff_A_Y0TP6KzS4_0),.din(w_dff_A_5B511Ywc8_0),.clk(gclk));
	jdff dff_A_Y0TP6KzS4_0(.dout(w_dff_A_8x9IJLGt1_0),.din(w_dff_A_Y0TP6KzS4_0),.clk(gclk));
	jdff dff_A_8x9IJLGt1_0(.dout(w_dff_A_reD76IVv3_0),.din(w_dff_A_8x9IJLGt1_0),.clk(gclk));
	jdff dff_A_reD76IVv3_0(.dout(w_dff_A_T0RPmTc91_0),.din(w_dff_A_reD76IVv3_0),.clk(gclk));
	jdff dff_A_T0RPmTc91_0(.dout(G370),.din(w_dff_A_T0RPmTc91_0),.clk(gclk));
	jdff dff_A_neBD5Ml89_2(.dout(w_dff_A_LeXqoUCC1_0),.din(w_dff_A_neBD5Ml89_2),.clk(gclk));
	jdff dff_A_LeXqoUCC1_0(.dout(w_dff_A_tlVoCh1Z5_0),.din(w_dff_A_LeXqoUCC1_0),.clk(gclk));
	jdff dff_A_tlVoCh1Z5_0(.dout(w_dff_A_uh82oImW5_0),.din(w_dff_A_tlVoCh1Z5_0),.clk(gclk));
	jdff dff_A_uh82oImW5_0(.dout(w_dff_A_BG2uy8SX9_0),.din(w_dff_A_uh82oImW5_0),.clk(gclk));
	jdff dff_A_BG2uy8SX9_0(.dout(G399),.din(w_dff_A_BG2uy8SX9_0),.clk(gclk));
endmodule

