module gf_c1908(G902, G900, G116, G143, G125, G227, G134, G952, G122, G221, G119, G898, G224, G107, G101, G140, G472, G110, G478, G104, G128, G131, G234, G137, G146, G210, G217, G953, G113, G237, G214, G469, G475, G57, G66, G69, G63, G54, G51, G72, G42, G39, G36, G3, G45, G6, G9, G27, G12, G30, G48, G15, G18, G21, G24, G60, G75, G33);
    input G902, G900, G116, G143, G125, G227, G134, G952, G122, G221, G119, G898, G224, G107, G101, G140, G472, G110, G478, G104, G128, G131, G234, G137, G146, G210, G217, G953, G113, G237, G214, G469, G475;
    output G57, G66, G69, G63, G54, G51, G72, G42, G39, G36, G3, G45, G6, G9, G27, G12, G30, G48, G15, G18, G21, G24, G60, G75, G33;
    wire n60;
    wire n63;
    wire n66;
    wire n70;
    wire n74;
    wire n77;
    wire n81;
    wire n85;
    wire n89;
    wire n93;
    wire n97;
    wire n101;
    wire n105;
    wire n109;
    wire n113;
    wire n116;
    wire n120;
    wire n123;
    wire n127;
    wire n131;
    wire n135;
    wire n139;
    wire n143;
    wire n147;
    wire n150;
    wire n154;
    wire n158;
    wire n161;
    wire n165;
    wire n169;
    wire n173;
    wire n177;
    wire n181;
    wire n185;
    wire n189;
    wire n193;
    wire n197;
    wire n201;
    wire n204;
    wire n207;
    wire n211;
    wire n215;
    wire n219;
    wire n223;
    wire n227;
    wire n230;
    wire n234;
    wire n238;
    wire n242;
    wire n246;
    wire n250;
    wire n254;
    wire n258;
    wire n262;
    wire n266;
    wire n269;
    wire n273;
    wire n277;
    wire n281;
    wire n285;
    wire n289;
    wire n293;
    wire n297;
    wire n301;
    wire n305;
    wire n309;
    wire n312;
    wire n316;
    wire n319;
    wire n323;
    wire n327;
    wire n331;
    wire n335;
    wire n339;
    wire n342;
    wire n346;
    wire n350;
    wire n354;
    wire n358;
    wire n362;
    wire n366;
    wire n370;
    wire n374;
    wire n378;
    wire n381;
    wire n385;
    wire n389;
    wire n392;
    wire n396;
    wire n399;
    wire n403;
    wire n407;
    wire n411;
    wire n415;
    wire n419;
    wire n423;
    wire n427;
    wire n431;
    wire n435;
    wire n439;
    wire n443;
    wire n446;
    wire n450;
    wire n454;
    wire n458;
    wire n462;
    wire n466;
    wire n470;
    wire n474;
    wire n478;
    wire n482;
    wire n486;
    wire n490;
    wire n494;
    wire n498;
    wire n502;
    wire n506;
    wire n510;
    wire n514;
    wire n518;
    wire n522;
    wire n526;
    wire n529;
    wire n533;
    wire n537;
    wire n541;
    wire n545;
    wire n549;
    wire n553;
    wire n557;
    wire n561;
    wire n565;
    wire n569;
    wire n573;
    wire n577;
    wire n581;
    wire n584;
    wire n588;
    wire n592;
    wire n596;
    wire n600;
    wire n604;
    wire n608;
    wire n612;
    wire n616;
    wire n620;
    wire n624;
    wire n628;
    wire n632;
    wire n636;
    wire n640;
    wire n644;
    wire n648;
    wire n652;
    wire n656;
    wire n659;
    wire n663;
    wire n667;
    wire n671;
    wire n675;
    wire n679;
    wire n683;
    wire n687;
    wire n691;
    wire n695;
    wire n699;
    wire n703;
    wire n707;
    wire n711;
    wire n715;
    wire n719;
    wire n723;
    wire n727;
    wire n731;
    wire n735;
    wire n739;
    wire n743;
    wire n747;
    wire n751;
    wire n755;
    wire n759;
    wire n763;
    wire n767;
    wire n771;
    wire n775;
    wire n779;
    wire n783;
    wire n787;
    wire n791;
    wire n795;
    wire n799;
    wire n803;
    wire n807;
    wire n811;
    wire n815;
    wire n819;
    wire n823;
    wire n827;
    wire n831;
    wire n835;
    wire n839;
    wire n843;
    wire n847;
    wire n851;
    wire n855;
    wire n859;
    wire n863;
    wire n867;
    wire n871;
    wire n875;
    wire n879;
    wire n887;
    wire n891;
    wire n895;
    wire n903;
    wire n907;
    wire n911;
    wire n914;
    wire n917;
    wire n921;
    wire n925;
    wire n929;
    wire n933;
    wire n937;
    wire n941;
    wire n945;
    wire n949;
    wire n953;
    wire n957;
    wire n960;
    wire n964;
    wire n968;
    wire n972;
    wire n976;
    wire n980;
    wire n984;
    wire n988;
    wire n992;
    wire n996;
    wire n1000;
    wire n1004;
    wire n1008;
    wire n1011;
    wire n1015;
    wire n1019;
    wire n1023;
    wire n1027;
    wire n1031;
    wire n1035;
    wire n1039;
    wire n1043;
    wire n1047;
    wire n1051;
    wire n1055;
    wire n1058;
    wire n1062;
    wire n1066;
    wire n1069;
    wire n1073;
    wire n1077;
    wire n1081;
    wire n1085;
    wire n1089;
    wire n1093;
    wire n1097;
    wire n1101;
    wire n1105;
    wire n1109;
    wire n1113;
    wire n1116;
    wire n1120;
    wire n1124;
    wire n1128;
    wire n1132;
    wire n1136;
    wire n1140;
    wire n1144;
    wire n1148;
    wire n1152;
    wire n1156;
    wire n1160;
    wire n1164;
    wire n1168;
    wire n1171;
    wire n1175;
    wire n1179;
    wire n1183;
    wire n1191;
    wire n1195;
    wire n1199;
    wire n1207;
    wire n1211;
    wire n1215;
    wire n1223;
    wire n1227;
    wire n1231;
    wire n1235;
    wire n1239;
    wire n1243;
    wire n1247;
    wire n1251;
    wire n1255;
    wire n1259;
    wire n1263;
    wire n1267;
    wire n1271;
    wire n1275;
    wire n1279;
    wire n1283;
    wire n1287;
    wire n1949;
    wire n1952;
    wire n1955;
    wire n1958;
    wire n1961;
    wire n1964;
    wire n1967;
    wire n1970;
    wire n1972;
    wire n1975;
    wire n1979;
    wire n1982;
    wire n1985;
    wire n1988;
    wire n1991;
    wire n1994;
    wire n1997;
    wire n2000;
    wire n2003;
    wire n2006;
    wire n2009;
    wire n2012;
    wire n2015;
    wire n2018;
    wire n2021;
    wire n2024;
    wire n2027;
    wire n2030;
    wire n2033;
    wire n2036;
    wire n2039;
    wire n2042;
    wire n2045;
    wire n2048;
    wire n2051;
    wire n2054;
    wire n2057;
    wire n2060;
    wire n2063;
    wire n2066;
    wire n2069;
    wire n2071;
    wire n2074;
    wire n2077;
    wire n2080;
    wire n2083;
    wire n2086;
    wire n2089;
    wire n2092;
    wire n2095;
    wire n2098;
    wire n2101;
    wire n2104;
    wire n2107;
    wire n2110;
    wire n2113;
    wire n2116;
    wire n2119;
    wire n2122;
    wire n2125;
    wire n2128;
    wire n2131;
    wire n2134;
    wire n2137;
    wire n2140;
    wire n2143;
    wire n2146;
    wire n2149;
    wire n2152;
    wire n2155;
    wire n2158;
    wire n2161;
    wire n2164;
    wire n2167;
    wire n2170;
    wire n2173;
    wire n2176;
    wire n2179;
    wire n2182;
    wire n2185;
    wire n2188;
    wire n2191;
    wire n2194;
    wire n2197;
    wire n2200;
    wire n2203;
    wire n2206;
    wire n2209;
    wire n2212;
    wire n2215;
    wire n2218;
    wire n2221;
    wire n2225;
    wire n2228;
    wire n2231;
    wire n2234;
    wire n2237;
    wire n2240;
    wire n2243;
    wire n2246;
    wire n2249;
    wire n2252;
    wire n2255;
    wire n2258;
    wire n2261;
    wire n2264;
    wire n2267;
    wire n2270;
    wire n2273;
    wire n2276;
    wire n2279;
    wire n2282;
    wire n2285;
    wire n2288;
    wire n2291;
    wire n2294;
    wire n2297;
    wire n2300;
    wire n2303;
    wire n2306;
    wire n2309;
    wire n2312;
    wire n2315;
    wire n2317;
    wire n2321;
    wire n2323;
    wire n2326;
    wire n2330;
    wire n2333;
    wire n2336;
    wire n2339;
    wire n2342;
    wire n2345;
    wire n2348;
    wire n2351;
    wire n2354;
    wire n2357;
    wire n2360;
    wire n2363;
    wire n2366;
    wire n2369;
    wire n2372;
    wire n2375;
    wire n2378;
    wire n2381;
    wire n2384;
    wire n2387;
    wire n2390;
    wire n2393;
    wire n2396;
    wire n2399;
    wire n2402;
    wire n2405;
    wire n2408;
    wire n2411;
    wire n2414;
    wire n2417;
    wire n2420;
    wire n2422;
    wire n2425;
    wire n2428;
    wire n2431;
    wire n2434;
    wire n2437;
    wire n2440;
    wire n2443;
    wire n2446;
    wire n2449;
    wire n2452;
    wire n2456;
    wire n2458;
    wire n2461;
    wire n2464;
    wire n2467;
    wire n2471;
    wire n2474;
    wire n2476;
    wire n2479;
    wire n2483;
    wire n2486;
    wire n2489;
    wire n2492;
    wire n2495;
    wire n2498;
    wire n2501;
    wire n2504;
    wire n2507;
    wire n2510;
    wire n2513;
    wire n2516;
    wire n2519;
    wire n2522;
    wire n2525;
    wire n2527;
    wire n2530;
    wire n2533;
    wire n2536;
    wire n2539;
    wire n2542;
    wire n2545;
    wire n2548;
    wire n2551;
    wire n2554;
    wire n2557;
    wire n2560;
    wire n2563;
    wire n2566;
    wire n2569;
    wire n2572;
    wire n2575;
    wire n2578;
    wire n2581;
    wire n2584;
    wire n2587;
    wire n2590;
    wire n2593;
    wire n2596;
    wire n2599;
    wire n2602;
    wire n2605;
    wire n2608;
    wire n2611;
    wire n2614;
    wire n2617;
    wire n2620;
    wire n2623;
    wire n2626;
    wire n2630;
    wire n2633;
    wire n2635;
    wire n2638;
    wire n2641;
    wire n2644;
    wire n2647;
    wire n2651;
    wire n2654;
    wire n2657;
    wire n2659;
    wire n2662;
    wire n2665;
    wire n2668;
    wire n2671;
    wire n2674;
    wire n2677;
    wire n2680;
    wire n2683;
    wire n2686;
    wire n2689;
    wire n2692;
    wire n2695;
    wire n2698;
    wire n2701;
    wire n2704;
    wire n2707;
    wire n2711;
    wire n2713;
    wire n2716;
    wire n2719;
    wire n2723;
    wire n2725;
    wire n2728;
    wire n2731;
    wire n2734;
    wire n2738;
    wire n2741;
    wire n2744;
    wire n2747;
    wire n2750;
    wire n2752;
    wire n2755;
    wire n2758;
    wire n2761;
    wire n2764;
    wire n2767;
    wire n2770;
    wire n2774;
    wire n2777;
    wire n2780;
    wire n2783;
    wire n2786;
    wire n2788;
    wire n2791;
    wire n2794;
    wire n2798;
    wire n2801;
    wire n2804;
    wire n2807;
    wire n2810;
    wire n2812;
    wire n2815;
    wire n2818;
    wire n2821;
    wire n2824;
    wire n2827;
    wire n2830;
    wire n2833;
    wire n2836;
    wire n2839;
    wire n2842;
    wire n2845;
    wire n2848;
    wire n2851;
    wire n2854;
    wire n2857;
    wire n2860;
    wire n2863;
    wire n2866;
    wire n2869;
    wire n2872;
    wire n2875;
    wire n2878;
    wire n2881;
    wire n2884;
    wire n2887;
    wire n2890;
    wire n2893;
    wire n2896;
    wire n2899;
    wire n2902;
    wire n2905;
    wire n2908;
    wire n2911;
    wire n2914;
    wire n2917;
    wire n2920;
    wire n2923;
    wire n2926;
    wire n2929;
    wire n2932;
    wire n2935;
    wire n2938;
    wire n2941;
    wire n2944;
    wire n2947;
    wire n2950;
    wire n2953;
    wire n2956;
    wire n2959;
    wire n2962;
    wire n2965;
    wire n2968;
    wire n2971;
    wire n2974;
    wire n2977;
    wire n2980;
    wire n2983;
    wire n2986;
    wire n2989;
    wire n2992;
    wire n2995;
    wire n2998;
    wire n3002;
    wire n3004;
    wire n3008;
    wire n3011;
    wire n3013;
    wire n3016;
    wire n3019;
    wire n3022;
    wire n3025;
    wire n3029;
    wire n3032;
    wire n3034;
    wire n3037;
    wire n3040;
    wire n3043;
    wire n3046;
    wire n3049;
    wire n3052;
    wire n3055;
    wire n3058;
    wire n3061;
    wire n3064;
    wire n3067;
    wire n3070;
    wire n3073;
    wire n3077;
    wire n3080;
    wire n3083;
    wire n3086;
    wire n3089;
    wire n3092;
    wire n3094;
    wire n3097;
    wire n3100;
    wire n3103;
    wire n3106;
    wire n3109;
    wire n3112;
    wire n3115;
    wire n3118;
    wire n3121;
    wire n3124;
    wire n3127;
    wire n3130;
    wire n3133;
    wire n3136;
    wire n3139;
    wire n3142;
    wire n3145;
    wire n3148;
    wire n3151;
    wire n3154;
    wire n3157;
    wire n3160;
    wire n3163;
    wire n3166;
    wire n3169;
    wire n3172;
    wire n3175;
    wire n3178;
    wire n3181;
    wire n3184;
    wire n3187;
    wire n3190;
    wire n3193;
    wire n3196;
    wire n3199;
    wire n3202;
    wire n3205;
    wire n3208;
    wire n3211;
    wire n3214;
    wire n3217;
    wire n3220;
    wire n3223;
    wire n3226;
    wire n3229;
    wire n3232;
    wire n3235;
    wire n3238;
    wire n3241;
    wire n3244;
    wire n3248;
    wire n3250;
    wire n3253;
    wire n3256;
    wire n3259;
    wire n3262;
    wire n3265;
    wire n3268;
    wire n3271;
    wire n3274;
    wire n3277;
    wire n3280;
    wire n3283;
    wire n3286;
    wire n3289;
    wire n3292;
    wire n3296;
    wire n3299;
    wire n3301;
    wire n3304;
    wire n3307;
    wire n3310;
    wire n3313;
    wire n3316;
    wire n3319;
    wire n3322;
    wire n3325;
    wire n3328;
    wire n3331;
    wire n3335;
    wire n3337;
    wire n3340;
    wire n3343;
    wire n3346;
    wire n3349;
    wire n3352;
    wire n3355;
    wire n3358;
    wire n3361;
    wire n3364;
    wire n3367;
    wire n3370;
    wire n3373;
    wire n3376;
    wire n3379;
    wire n3382;
    wire n3385;
    wire n3388;
    wire n3391;
    wire n3394;
    wire n3397;
    wire n3400;
    wire n3403;
    wire n3407;
    wire n3409;
    wire n3412;
    wire n3415;
    wire n3418;
    wire n3421;
    wire n3424;
    wire n3427;
    wire n3430;
    wire n3433;
    wire n3436;
    wire n3439;
    wire n3442;
    wire n3445;
    wire n3448;
    wire n3451;
    wire n3454;
    wire n3457;
    wire n3460;
    wire n3463;
    wire n3466;
    wire n3469;
    wire n3472;
    wire n3475;
    wire n3478;
    wire n3481;
    wire n3484;
    wire n3487;
    wire n3490;
    wire n3493;
    wire n3496;
    wire n3499;
    wire n3502;
    wire n3505;
    wire n3508;
    wire n3511;
    wire n3514;
    wire n3517;
    wire n3520;
    wire n3523;
    wire n3526;
    wire n3529;
    wire n3532;
    wire n3535;
    wire n3538;
    wire n3541;
    wire n3544;
    wire n3547;
    wire n3550;
    wire n3553;
    wire n3556;
    wire n3560;
    wire n3563;
    wire n3565;
    wire n3568;
    wire n3571;
    wire n3574;
    wire n3577;
    wire n3580;
    wire n3583;
    wire n3586;
    wire n3589;
    wire n3592;
    wire n3595;
    wire n3598;
    wire n3601;
    wire n3604;
    wire n3607;
    wire n3610;
    wire n3613;
    wire n3616;
    wire n3619;
    wire n3622;
    wire n3625;
    wire n3628;
    wire n3631;
    wire n3634;
    wire n3637;
    wire n3640;
    wire n3643;
    wire n3646;
    wire n3649;
    wire n3652;
    wire n3655;
    wire n3658;
    wire n3661;
    wire n3664;
    wire n3667;
    wire n3670;
    wire n3673;
    wire n3676;
    wire n3679;
    wire n3682;
    wire n3685;
    wire n3688;
    wire n3691;
    wire n3694;
    wire n3697;
    wire n3700;
    wire n3703;
    wire n3706;
    wire n3709;
    wire n3712;
    wire n3715;
    wire n3718;
    wire n3722;
    wire n3724;
    wire n3727;
    wire n3730;
    wire n3733;
    wire n3736;
    wire n3739;
    wire n3742;
    wire n3745;
    wire n3748;
    wire n3751;
    wire n3754;
    wire n3757;
    wire n3760;
    wire n3763;
    wire n3766;
    wire n3769;
    wire n3772;
    wire n3775;
    wire n3778;
    wire n3781;
    wire n3784;
    wire n3787;
    wire n3790;
    wire n3793;
    wire n3796;
    wire n3799;
    wire n3802;
    wire n3805;
    wire n3808;
    wire n3811;
    wire n3814;
    wire n3817;
    wire n3820;
    wire n3823;
    wire n3826;
    wire n3829;
    wire n3832;
    wire n3835;
    wire n3838;
    wire n3841;
    wire n3844;
    wire n3847;
    wire n3851;
    wire n3854;
    wire n3857;
    wire n3859;
    wire n3862;
    wire n3865;
    wire n3868;
    wire n3871;
    wire n3874;
    wire n3877;
    wire n3880;
    wire n3883;
    wire n3886;
    wire n3889;
    wire n3892;
    wire n3895;
    wire n3898;
    wire n3901;
    wire n3904;
    wire n3907;
    wire n3910;
    wire n3913;
    wire n3916;
    wire n3919;
    wire n3922;
    wire n3925;
    wire n3928;
    wire n3931;
    wire n3934;
    wire n3937;
    wire n3940;
    wire n3943;
    wire n3946;
    wire n3949;
    wire n3952;
    wire n3955;
    wire n3958;
    wire n3961;
    wire n3964;
    wire n3967;
    wire n3970;
    wire n3973;
    wire n3976;
    wire n3979;
    wire n3982;
    wire n3985;
    wire n3988;
    wire n3991;
    wire n3994;
    wire n3997;
    wire n4000;
    wire n4003;
    wire n4006;
    wire n4009;
    wire n4012;
    wire n4015;
    wire n4019;
    wire n4022;
    wire n4024;
    wire n4027;
    wire n4030;
    wire n4033;
    wire n4036;
    wire n4039;
    wire n4042;
    wire n4045;
    wire n4048;
    wire n4051;
    wire n4054;
    wire n4057;
    wire n4060;
    wire n4063;
    wire n4066;
    wire n4069;
    wire n4072;
    wire n4075;
    wire n4078;
    wire n4081;
    wire n4084;
    wire n4087;
    wire n4090;
    wire n4093;
    wire n4096;
    wire n4099;
    wire n4102;
    wire n4105;
    wire n4108;
    wire n4111;
    wire n4114;
    wire n4117;
    wire n4120;
    wire n4123;
    wire n4126;
    wire n4129;
    wire n4132;
    wire n4135;
    wire n4138;
    wire n4141;
    wire n4144;
    wire n4147;
    wire n4150;
    wire n4153;
    wire n4156;
    wire n4159;
    wire n4162;
    wire n4165;
    wire n4168;
    wire n4171;
    wire n4174;
    wire n4177;
    wire n4180;
    wire n4183;
    wire n4186;
    wire n4189;
    wire n4192;
    wire n4195;
    wire n4198;
    wire n4201;
    wire n4204;
    wire n4207;
    wire n4210;
    wire n4213;
    wire n4216;
    wire n4219;
    wire n4222;
    wire n4225;
    wire n4229;
    wire n4232;
    wire n4235;
    wire n4238;
    wire n4241;
    wire n4244;
    wire n4247;
    wire n4250;
    wire n4253;
    wire n4256;
    wire n4259;
    wire n4262;
    wire n4265;
    wire n4268;
    wire n4271;
    wire n4274;
    wire n4276;
    wire n4279;
    wire n4282;
    wire n4285;
    wire n4288;
    wire n4291;
    wire n4294;
    wire n4297;
    wire n4300;
    wire n4303;
    wire n4306;
    wire n4309;
    wire n4312;
    wire n4315;
    wire n4318;
    wire n4321;
    wire n4324;
    wire n4327;
    wire n4330;
    wire n4333;
    wire n4336;
    wire n4339;
    wire n4342;
    wire n4345;
    wire n4348;
    wire n4351;
    wire n4354;
    wire n4357;
    wire n4360;
    wire n4363;
    wire n4366;
    wire n4369;
    wire n4372;
    wire n4375;
    wire n4378;
    wire n4381;
    wire n4384;
    wire n4387;
    wire n4390;
    wire n4393;
    wire n4396;
    wire n4399;
    wire n4402;
    wire n4405;
    wire n4408;
    wire n4411;
    wire n4414;
    wire n4417;
    wire n4420;
    wire n4423;
    wire n4426;
    wire n4429;
    wire n4432;
    wire n4435;
    wire n4438;
    wire n4441;
    wire n4444;
    wire n4447;
    wire n4450;
    wire n4454;
    wire n4456;
    wire n4459;
    wire n4462;
    wire n4465;
    wire n4468;
    wire n4471;
    wire n4474;
    wire n4480;
    wire n4483;
    wire n4486;
    wire n4489;
    wire n4492;
    wire n4495;
    wire n4498;
    wire n4504;
    wire n4507;
    wire n4510;
    wire n4513;
    wire n4516;
    wire n4519;
    wire n4522;
    wire n4528;
    wire n4531;
    wire n4534;
    wire n4537;
    wire n4540;
    wire n4543;
    wire n4546;
    wire n4552;
    wire n4555;
    wire n4558;
    wire n4561;
    wire n4564;
    wire n4567;
    wire n4570;
    wire n4576;
    wire n4579;
    wire n4582;
    wire n4585;
    wire n4588;
    wire n4591;
    wire n4594;
    wire n4600;
    wire n4603;
    wire n4606;
    wire n4609;
    wire n4612;
    wire n4615;
    wire n4618;
    wire n4624;
    wire n4627;
    wire n4630;
    wire n4633;
    wire n4636;
    wire n4639;
    wire n4642;
    wire n4648;
    wire n4651;
    wire n4654;
    wire n4657;
    wire n4660;
    wire n4663;
    wire n4666;
    wire n4672;
    wire n4675;
    wire n4678;
    wire n4681;
    wire n4684;
    wire n4687;
    wire n4690;
    wire n4696;
    wire n4699;
    wire n4702;
    wire n4705;
    wire n4708;
    wire n4711;
    wire n4717;
    wire n4720;
    wire n4723;
    wire n4726;
    wire n4729;
    wire n4732;
    wire n4735;
    wire n4741;
    wire n4744;
    wire n4747;
    wire n4750;
    wire n4753;
    wire n4756;
    wire n4759;
    wire n4765;
    wire n4768;
    wire n4771;
    wire n4774;
    wire n4777;
    wire n4780;
    wire n4783;
    wire n4789;
    wire n4792;
    wire n4795;
    wire n4798;
    wire n4801;
    wire n4804;
    wire n4807;
    wire n4813;
    wire n4816;
    wire n4819;
    wire n4822;
    wire n4825;
    wire n4828;
    wire n4831;
    wire n4840;
    wire n4846;
    jnot g000(.din(G902), .dout(n60));
    jnot g001(.din(G221), .dout(n63));
    jnot g002(.din(G234), .dout(n66));
    jor g003(.dinb(n66), .dina(n3601), .dout(n70));
    jor g004(.dinb(n3407), .dina(n70), .dout(n74));
    jnot g005(.din(G110), .dout(n77));
    jxor g006(.dinb(n77), .dina(n3370), .dout(n81));
    jxor g007(.dinb(n74), .dina(n3335), .dout(n85));
    jxor g008(.dinb(G125), .dina(G140), .dout(n89));
    jxor g009(.dinb(n3722), .dina(n89), .dout(n93));
    jxor g010(.dinb(G128), .dina(G137), .dout(n97));
    jxor g011(.dinb(n93), .dina(n3299), .dout(n101));
    jxor g012(.dinb(n85), .dina(n3296), .dout(n105));
    jand g013(.dinb(n3433), .dina(n105), .dout(n109));
    jand g014(.dinb(n3409), .dina(n60), .dout(n113));
    jnot g015(.din(n113), .dout(n116));
    jand g016(.dinb(n4015), .dina(n116), .dout(n120));
    jnot g017(.din(n120), .dout(n123));
    jxor g018(.dinb(n109), .dina(n3248), .dout(n127));
    jxor g019(.dinb(G128), .dina(G143), .dout(n131));
    jxor g020(.dinb(n3722), .dina(n131), .dout(n135));
    jxor g021(.dinb(G134), .dina(G137), .dout(n139));
    jxor g022(.dinb(n3598), .dina(n139), .dout(n143));
    jxor g023(.dinb(n135), .dina(n143), .dout(n147));
    jnot g024(.din(G113), .dout(n150));
    jxor g025(.dinb(G116), .dina(G119), .dout(n154));
    jxor g026(.dinb(n150), .dina(n154), .dout(n158));
    jnot g027(.din(G210), .dout(n161));
    jor g028(.dinb(G237), .dina(G953), .dout(n165));
    jor g029(.dinb(n161), .dina(n165), .dout(n169));
    jxor g030(.dinb(n3214), .dina(n169), .dout(n173));
    jxor g031(.dinb(n3220), .dina(n173), .dout(n177));
    jxor g032(.dinb(n3226), .dina(n177), .dout(n181));
    jand g033(.dinb(n3421), .dina(n181), .dout(n185));
    jxor g034(.dinb(n3229), .dina(n185), .dout(n189));
    jand g035(.dinb(n127), .dina(n189), .dout(n193));
    jor g036(.dinb(G237), .dina(G902), .dout(n197));
    jand g037(.dinb(n3604), .dina(n197), .dout(n201));
    jnot g038(.din(n201), .dout(n204));
    jnot g039(.din(G101), .dout(n207));
    jxor g040(.dinb(G104), .dina(G107), .dout(n211));
    jxor g041(.dinb(n207), .dina(n211), .dout(n215));
    jxor g042(.dinb(n158), .dina(n215), .dout(n219));
    jxor g043(.dinb(G110), .dina(G122), .dout(n223));
    jxor g044(.dinb(n219), .dina(n3011), .dout(n227));
    jnot g045(.din(G953), .dout(n230));
    jand g046(.dinb(n3004), .dina(n230), .dout(n234));
    jxor g047(.dinb(n3685), .dina(n135), .dout(n238));
    jxor g048(.dinb(n3002), .dina(n238), .dout(n242));
    jxor g049(.dinb(n227), .dina(n242), .dout(n246));
    jand g050(.dinb(n4129), .dina(n246), .dout(n250));
    jand g051(.dinb(n3178), .dina(n197), .dout(n254));
    jxor g052(.dinb(n250), .dina(n2950), .dout(n258));
    jand g053(.dinb(n3022), .dina(n258), .dout(n262));
    jand g054(.dinb(n3412), .dina(n116), .dout(n266));
    jnot g055(.din(n266), .dout(n269));
    jand g056(.dinb(n2851), .dina(n230), .dout(n273));
    jxor g057(.dinb(n77), .dina(n3649), .dout(n277));
    jxor g058(.dinb(n273), .dina(n277), .dout(n281));
    jxor g059(.dinb(n3013), .dina(n281), .dout(n285));
    jxor g060(.dinb(n3223), .dina(n285), .dout(n289));
    jand g061(.dinb(n4129), .dina(n289), .dout(n293));
    jxor g062(.dinb(n2902), .dina(n293), .dout(n297));
    jand g063(.dinb(n2926), .dina(n297), .dout(n301));
    jand g064(.dinb(n262), .dina(n301), .dout(n305));
    jor g065(.dinb(n3511), .dina(n230), .dout(n309));
    jnot g066(.din(n309), .dout(n312));
    jand g067(.dinb(G234), .dina(G237), .dout(n316));
    jnot g068(.din(n316), .dout(n319));
    jand g069(.dinb(n4153), .dina(n319), .dout(n323));
    jand g070(.dinb(n312), .dina(n323), .dout(n327));
    jand g071(.dinb(n4450), .dina(n319), .dout(n331));
    jand g072(.dinb(n3964), .dina(n331), .dout(n335));
    jor g073(.dinb(n327), .dina(n335), .dout(n339));
    jnot g074(.din(G478), .dout(n342));
    jxor g075(.dinb(n4126), .dina(n131), .dout(n346));
    jand g076(.dinb(n3970), .dina(n230), .dout(n350));
    jand g077(.dinb(n4022), .dina(n350), .dout(n354));
    jxor g078(.dinb(G116), .dina(G122), .dout(n358));
    jxor g079(.dinb(n3961), .dina(n358), .dout(n362));
    jxor g080(.dinb(n354), .dina(n3857), .dout(n366));
    jxor g081(.dinb(n3854), .dina(n366), .dout(n370));
    jand g082(.dinb(n4129), .dina(n370), .dout(n374));
    jxor g083(.dinb(n2786), .dina(n374), .dout(n378));
    jnot g084(.din(G475), .dout(n381));
    jxor g085(.dinb(G113), .dina(G122), .dout(n385));
    jxor g086(.dinb(n3790), .dina(n385), .dout(n389));
    jnot g087(.din(G214), .dout(n392));
    jor g088(.dinb(n392), .dina(n165), .dout(n396));
    jnot g089(.din(G131), .dout(n399));
    jxor g090(.dinb(n399), .dina(n4057), .dout(n403));
    jxor g091(.dinb(n396), .dina(n403), .dout(n407));
    jxor g092(.dinb(n3607), .dina(n407), .dout(n411));
    jxor g093(.dinb(n3563), .dina(n411), .dout(n415));
    jand g094(.dinb(n4141), .dina(n415), .dout(n419));
    jxor g095(.dinb(n2750), .dina(n419), .dout(n423));
    jand g096(.dinb(n378), .dina(n423), .dout(n427));
    jand g097(.dinb(n3445), .dina(n427), .dout(n431));
    jand g098(.dinb(n305), .dina(n431), .dout(n435));
    jand g099(.dinb(n2752), .dina(n435), .dout(n439));
    jxor g100(.dinb(n3181), .dina(n439), .dout(n443));
    jnot g101(.din(G472), .dout(n446));
    jxor g102(.dinb(n3092), .dina(n185), .dout(n450));
    jand g103(.dinb(n127), .dina(n450), .dout(n454));
    jand g104(.dinb(n305), .dina(n3077), .dout(n458));
    jxor g105(.dinb(n3793), .dina(n419), .dout(n462));
    jand g106(.dinb(n378), .dina(n462), .dout(n466));
    jand g107(.dinb(n3445), .dina(n466), .dout(n470));
    jand g108(.dinb(n458), .dina(n2770), .dout(n474));
    jxor g109(.dinb(n3757), .dina(n474), .dout(n478));
    jxor g110(.dinb(n4207), .dina(n374), .dout(n482));
    jand g111(.dinb(n482), .dina(n423), .dout(n486));
    jand g112(.dinb(n3445), .dina(n486), .dout(n490));
    jand g113(.dinb(n458), .dina(n2723), .dout(n494));
    jxor g114(.dinb(n3928), .dina(n494), .dout(n498));
    jxor g115(.dinb(n109), .dina(n3250), .dout(n502));
    jand g116(.dinb(n502), .dina(n450), .dout(n506));
    jand g117(.dinb(n435), .dina(n2707), .dout(n510));
    jxor g118(.dinb(n3373), .dina(n510), .dout(n514));
    jand g119(.dinb(n502), .dina(n189), .dout(n518));
    jand g120(.dinb(n305), .dina(n2701), .dout(n522));
    jor g121(.dinb(n2695), .dina(n230), .dout(n526));
    jnot g122(.din(n526), .dout(n529));
    jand g123(.dinb(n323), .dina(n529), .dout(n533));
    jor g124(.dinb(n335), .dina(n533), .dout(n537));
    jand g125(.dinb(n486), .dina(n2671), .dout(n541));
    jand g126(.dinb(n522), .dina(n2641), .dout(n545));
    jxor g127(.dinb(n4060), .dina(n545), .dout(n549));
    jand g128(.dinb(n482), .dina(n462), .dout(n553));
    jand g129(.dinb(n193), .dina(n553), .dout(n557));
    jand g130(.dinb(n2668), .dina(n557), .dout(n561));
    jand g131(.dinb(n2788), .dina(n561), .dout(n565));
    jxor g132(.dinb(n4024), .dina(n565), .dout(n569));
    jand g133(.dinb(n466), .dina(n2671), .dout(n573));
    jand g134(.dinb(n522), .dina(n2665), .dout(n577));
    jxor g135(.dinb(n3691), .dina(n577), .dout(n581));
    jnot g136(.din(G469), .dout(n584));
    jxor g137(.dinb(n2810), .dina(n293), .dout(n588));
    jand g138(.dinb(n2920), .dina(n588), .dout(n592));
    jand g139(.dinb(n262), .dina(n592), .dout(n596));
    jand g140(.dinb(n2761), .dina(n596), .dout(n600));
    jand g141(.dinb(n2767), .dina(n600), .dout(n604));
    jxor g142(.dinb(n3724), .dina(n604), .dout(n608));
    jand g143(.dinb(n2723), .dina(n600), .dout(n612));
    jxor g144(.dinb(n3895), .dina(n612), .dout(n616));
    jand g145(.dinb(n431), .dina(n2698), .dout(n620));
    jand g146(.dinb(n2719), .dina(n620), .dout(n624));
    jxor g147(.dinb(n3337), .dina(n624), .dout(n628));
    jand g148(.dinb(n3077), .dina(n596), .dout(n632));
    jand g149(.dinb(n3454), .dina(n632), .dout(n636));
    jand g150(.dinb(n3514), .dina(n636), .dout(n640));
    jxor g151(.dinb(n3859), .dina(n640), .dout(n644));
    jand g152(.dinb(n2711), .dina(n573), .dout(n648));
    jand g153(.dinb(n2794), .dina(n648), .dout(n652));
    jxor g154(.dinb(n3652), .dina(n652), .dout(n656));
    jnot g155(.din(n254), .dout(n659));
    jxor g156(.dinb(n250), .dina(n2657), .dout(n663));
    jand g157(.dinb(n3016), .dina(n663), .dout(n667));
    jand g158(.dinb(n301), .dina(n667), .dout(n671));
    jand g159(.dinb(n2758), .dina(n671), .dout(n675));
    jand g160(.dinb(n2662), .dina(n675), .dout(n679));
    jxor g161(.dinb(n3565), .dina(n679), .dout(n683));
    jand g162(.dinb(n2638), .dina(n675), .dout(n687));
    jxor g163(.dinb(n4093), .dina(n687), .dout(n691));
    jand g164(.dinb(n427), .dina(n518), .dout(n695));
    jand g165(.dinb(n2680), .dina(n695), .dout(n699));
    jand g166(.dinb(n2644), .dina(n699), .dout(n703));
    jxor g167(.dinb(n3301), .dina(n703), .dout(n707));
    jand g168(.dinb(n648), .dina(n2647), .dout(n711));
    jxor g169(.dinb(n3616), .dina(n711), .dout(n715));
    jor g170(.dinb(n439), .dina(n494), .dout(n719));
    jor g171(.dinb(n2764), .dina(n719), .dout(n723));
    jor g172(.dinb(n2791), .dina(n723), .dout(n727));
    jor g173(.dinb(n612), .dina(n624), .dout(n731));
    jor g174(.dinb(n2704), .dina(n731), .dout(n735));
    jor g175(.dinb(n2713), .dina(n735), .dout(n739));
    jor g176(.dinb(n727), .dina(n739), .dout(n743));
    jor g177(.dinb(n703), .dina(n711), .dout(n747));
    jor g178(.dinb(n2659), .dina(n747), .dout(n751));
    jor g179(.dinb(n679), .dina(n687), .dout(n755));
    jor g180(.dinb(n565), .dina(n652), .dout(n759));
    jor g181(.dinb(n2635), .dina(n759), .dout(n763));
    jor g182(.dinb(n2633), .dina(n763), .dout(n767));
    jor g183(.dinb(n2630), .dina(n767), .dout(n771));
    jor g184(.dinb(n743), .dina(n771), .dout(n775));
    jand g185(.dinb(n663), .dina(n588), .dout(n779));
    jxor g186(.dinb(n3034), .dina(n266), .dout(n783));
    jand g187(.dinb(n779), .dina(n1991), .dout(n787));
    jor g188(.dinb(n671), .dina(n787), .dout(n791));
    jand g189(.dinb(n3073), .dina(n791), .dout(n795));
    jand g190(.dinb(n3032), .dina(n269), .dout(n799));
    jand g191(.dinb(n779), .dina(n1982), .dout(n803));
    jxor g192(.dinb(n127), .dina(n450), .dout(n807));
    jand g193(.dinb(n803), .dina(n1970), .dout(n811));
    jor g194(.dinb(n632), .dina(n811), .dout(n815));
    jor g195(.dinb(n795), .dina(n815), .dout(n819));
    jand g196(.dinb(n2725), .dina(n819), .dout(n823));
    jand g197(.dinb(n3481), .dina(n823), .dout(n827));
    jor g198(.dinb(n775), .dina(n1967), .dout(n831));
    jand g199(.dinb(n4402), .dina(n831), .dout(n835));
    jor g200(.dinb(n378), .dina(n423), .dout(n839));
    jor g201(.dinb(n3469), .dina(n427), .dout(n843));
    jand g202(.dinb(n2437), .dina(n843), .dout(n847));
    jand g203(.dinb(n3070), .dina(n847), .dout(n851));
    jand g204(.dinb(n1972), .dina(n851), .dout(n855));
    jor g205(.dinb(n4321), .dina(n855), .dout(n859));
    jor g206(.dinb(n835), .dina(n1961), .dout(n863));
    jor g207(.dinb(n4454), .dina(n230), .dout(n867));
    jand g208(.dinb(n3130), .dina(n775), .dout(n871));
    jand g209(.dinb(n2167), .dina(n871), .dout(n875));
    jxor g210(.dinb(n2962), .dina(n875), .dout(n879));
    jand g211(.dinb(n4225), .dina(n879), .dout(G51));
    jand g212(.dinb(n2854), .dina(n775), .dout(n887));
    jand g213(.dinb(n2116), .dina(n887), .dout(n891));
    jxor g214(.dinb(n2812), .dina(n891), .dout(n895));
    jand g215(.dinb(n4225), .dina(n895), .dout(G54));
    jand g216(.dinb(G475), .dina(G902), .dout(n903));
    jand g217(.dinb(n775), .dina(n2071), .dout(n907));
    jor g218(.dinb(n3523), .dina(n907), .dout(n911));
    jnot g219(.din(n415), .dout(n914));
    jnot g220(.din(n339), .dout(n917));
    jor g221(.dinb(n502), .dina(n189), .dout(n921));
    jor g222(.dinb(n3055), .dina(n663), .dout(n925));
    jor g223(.dinb(n2941), .dina(n297), .dout(n929));
    jor g224(.dinb(n925), .dina(n929), .dout(n933));
    jor g225(.dinb(n2321), .dina(n933), .dout(n937));
    jor g226(.dinb(n2323), .dina(n937), .dout(n941));
    jor g227(.dinb(n2428), .dina(n941), .dout(n945));
    jor g228(.dinb(n2932), .dina(n588), .dout(n949));
    jor g229(.dinb(n925), .dina(n949), .dout(n953));
    jor g230(.dinb(n953), .dina(n2321), .dout(n957));
    jnot g231(.din(n470), .dout(n960));
    jor g232(.dinb(n957), .dina(n960), .dout(n964));
    jor g233(.dinb(n502), .dina(n450), .dout(n968));
    jor g234(.dinb(n482), .dina(n462), .dout(n972));
    jor g235(.dinb(n2333), .dina(n972), .dout(n976));
    jor g236(.dinb(n953), .dina(n976), .dout(n980));
    jor g237(.dinb(n2317), .dina(n980), .dout(n984));
    jor g238(.dinb(n378), .dina(n462), .dout(n988));
    jor g239(.dinb(n2333), .dina(n988), .dout(n992));
    jor g240(.dinb(n957), .dina(n2315), .dout(n996));
    jand g241(.dinb(n984), .dina(n996), .dout(n1000));
    jand g242(.dinb(n2312), .dina(n1000), .dout(n1004));
    jand g243(.dinb(n2309), .dina(n1004), .dout(n1008));
    jnot g244(.din(n604), .dout(n1011));
    jor g245(.dinb(n127), .dina(n189), .dout(n1015));
    jor g246(.dinb(n980), .dina(n2452), .dout(n1019));
    jor g247(.dinb(n2443), .dina(n933), .dout(n1023));
    jor g248(.dinb(n2315), .dina(n1023), .dout(n1027));
    jor g249(.dinb(n127), .dina(n450), .dout(n1031));
    jor g250(.dinb(n976), .dina(n2461), .dout(n1035));
    jor g251(.dinb(n2425), .dina(n1035), .dout(n1039));
    jand g252(.dinb(n1027), .dina(n1039), .dout(n1043));
    jand g253(.dinb(n2306), .dina(n1043), .dout(n1047));
    jand g254(.dinb(n2303), .dina(n1047), .dout(n1051));
    jand g255(.dinb(n1008), .dina(n1051), .dout(n1055));
    jnot g256(.din(n577), .dout(n1058));
    jor g257(.dinb(n3040), .dina(n258), .dout(n1062));
    jor g258(.dinb(n949), .dina(n1062), .dout(n1066));
    jnot g259(.din(n537), .dout(n1069));
    jor g260(.dinb(n972), .dina(n1031), .dout(n1073));
    jor g261(.dinb(n2467), .dina(n1073), .dout(n1077));
    jor g262(.dinb(n2479), .dina(n1077), .dout(n1081));
    jor g263(.dinb(n482), .dina(n423), .dout(n1085));
    jor g264(.dinb(n1085), .dina(n2474), .dout(n1089));
    jor g265(.dinb(n2456), .dina(n1089), .dout(n1093));
    jor g266(.dinb(n1093), .dina(n2476), .dout(n1097));
    jand g267(.dinb(n1081), .dina(n1097), .dout(n1101));
    jand g268(.dinb(n1058), .dina(n1101), .dout(n1105));
    jor g269(.dinb(n2446), .dina(n1066), .dout(n1109));
    jor g270(.dinb(n2449), .dina(n1109), .dout(n1113));
    jnot g271(.din(n541), .dout(n1116));
    jor g272(.dinb(n1116), .dina(n1109), .dout(n1120));
    jand g273(.dinb(n1113), .dina(n1120), .dout(n1124));
    jor g274(.dinb(n953), .dina(n2458), .dout(n1128));
    jor g275(.dinb(n1128), .dina(n1116), .dout(n1132));
    jor g276(.dinb(n968), .dina(n839), .dout(n1136));
    jor g277(.dinb(n2464), .dina(n1136), .dout(n1140));
    jor g278(.dinb(n2440), .dina(n1140), .dout(n1144));
    jor g279(.dinb(n2422), .dina(n1093), .dout(n1148));
    jand g280(.dinb(n1144), .dina(n1148), .dout(n1152));
    jand g281(.dinb(n2420), .dina(n1152), .dout(n1156));
    jand g282(.dinb(n2417), .dina(n1156), .dout(n1160));
    jand g283(.dinb(n2414), .dina(n1160), .dout(n1164));
    jand g284(.dinb(n1055), .dina(n1164), .dout(n1168));
    jnot g285(.din(n903), .dout(n1171));
    jor g286(.dinb(n1168), .dina(n2069), .dout(n1175));
    jor g287(.dinb(n2027), .dina(n1175), .dout(n1179));
    jand g288(.dinb(n4274), .dina(n1179), .dout(n1183));
    jand g289(.dinb(n1994), .dina(n1183), .dout(G60));
    jand g290(.dinb(n4159), .dina(n775), .dout(n1191));
    jand g291(.dinb(n2578), .dina(n1191), .dout(n1195));
    jxor g292(.dinb(n3811), .dina(n1195), .dout(n1199));
    jand g293(.dinb(n2221), .dina(n1199), .dout(G63));
    jand g294(.dinb(n3973), .dina(n775), .dout(n1207));
    jand g295(.dinb(n2527), .dina(n1207), .dout(n1211));
    jxor g296(.dinb(n3256), .dina(n1211), .dout(n1215));
    jand g297(.dinb(n2218), .dina(n1215), .dout(G66));
    jor g298(.dinb(n227), .dina(n3508), .dout(n1223));
    jor g299(.dinb(n4276), .dina(n1055), .dout(n1227));
    jand g300(.dinb(G224), .dina(G898), .dout(n1231));
    jor g301(.dinb(n230), .dina(n1231), .dout(n1235));
    jand g302(.dinb(n1227), .dina(n2300), .dout(n1239));
    jxor g303(.dinb(n2258), .dina(n1239), .dout(n1243));
    jor g304(.dinb(n4357), .dina(n1164), .dout(n1247));
    jand g305(.dinb(G227), .dina(G900), .dout(n1251));
    jor g306(.dinb(n230), .dina(n1251), .dout(n1255));
    jand g307(.dinb(n1247), .dina(n2411), .dout(n1259));
    jxor g308(.dinb(n3610), .dina(n147), .dout(n1263));
    jor g309(.dinb(n2692), .dina(n1263), .dout(n1267));
    jxor g310(.dinb(n1259), .dina(n2369), .dout(n1271));
    jand g311(.dinb(G472), .dina(G902), .dout(n1275));
    jand g312(.dinb(n775), .dina(n2525), .dout(n1279));
    jxor g313(.dinb(n3094), .dina(n1279), .dout(n1283));
    jand g314(.dinb(n4274), .dina(n1283), .dout(n1287));
    jdff dff_A_CR8MmAXU9_2(.din(n1287), .dout(G57));
    jdff dff_A_Xaaac5Zg9_0(.din(n4846), .dout(G72));
    jdff dff_A_bfIBpwvT2_2(.din(n1271), .dout(n4846));
    jdff dff_A_FggnYhHZ2_0(.din(n4840), .dout(G69));
    jdff dff_A_jrsgWhlw6_2(.din(n1243), .dout(n4840));
    jdff dff_A_NWXt4Snf1_2(.din(n863), .dout(G75));
    jdff dff_A_ADq0GnWf3_0(.din(n4831), .dout(G42));
    jdff dff_A_tGRE1uAg3_0(.din(n4828), .dout(n4831));
    jdff dff_A_KIFz7CH72_0(.din(n4825), .dout(n4828));
    jdff dff_A_C5lsZQZP3_0(.din(n4822), .dout(n4825));
    jdff dff_A_gAgSSfCd1_0(.din(n4819), .dout(n4822));
    jdff dff_A_gIDHvzis8_0(.din(n4816), .dout(n4819));
    jdff dff_A_vxdStgLY0_0(.din(n4813), .dout(n4816));
    jdff dff_A_K9N8MOyh8_2(.din(n715), .dout(n4813));
    jdff dff_A_qGGumymi0_0(.din(n4807), .dout(G39));
    jdff dff_A_yvSMQFQ96_0(.din(n4804), .dout(n4807));
    jdff dff_A_s3ze39kW7_0(.din(n4801), .dout(n4804));
    jdff dff_A_pQ3YMCOW1_0(.din(n4798), .dout(n4801));
    jdff dff_A_gCTlPJdx7_0(.din(n4795), .dout(n4798));
    jdff dff_A_xevfPlMV8_0(.din(n4792), .dout(n4795));
    jdff dff_A_5Bs10Pmm9_0(.din(n4789), .dout(n4792));
    jdff dff_A_H0wbY1Ub8_2(.din(n707), .dout(n4789));
    jdff dff_A_9S8T0T9S2_0(.din(n4783), .dout(G36));
    jdff dff_A_6hExMG0z6_0(.din(n4780), .dout(n4783));
    jdff dff_A_8KdmLDuJ5_0(.din(n4777), .dout(n4780));
    jdff dff_A_WZS4Vqqr7_0(.din(n4774), .dout(n4777));
    jdff dff_A_HinQTAFs2_0(.din(n4771), .dout(n4774));
    jdff dff_A_S2Tp7smu0_0(.din(n4768), .dout(n4771));
    jdff dff_A_uOSfjerm5_0(.din(n4765), .dout(n4768));
    jdff dff_A_9hMXUQKg7_2(.din(n691), .dout(n4765));
    jdff dff_A_2uHjnuT57_0(.din(n4759), .dout(G33));
    jdff dff_A_iY3FJa145_0(.din(n4756), .dout(n4759));
    jdff dff_A_66F1CsVM0_0(.din(n4753), .dout(n4756));
    jdff dff_A_bnlqfMaz2_0(.din(n4750), .dout(n4753));
    jdff dff_A_cFslUK5m3_0(.din(n4747), .dout(n4750));
    jdff dff_A_4AI7CPcV2_0(.din(n4744), .dout(n4747));
    jdff dff_A_BURVCN1F8_0(.din(n4741), .dout(n4744));
    jdff dff_A_pvSnXxJb3_2(.din(n683), .dout(n4741));
    jdff dff_A_UjaTMIZF1_0(.din(n4735), .dout(G27));
    jdff dff_A_3exUiFpL3_0(.din(n4732), .dout(n4735));
    jdff dff_A_jaUi27hL0_0(.din(n4729), .dout(n4732));
    jdff dff_A_q0ckrtDo0_0(.din(n4726), .dout(n4729));
    jdff dff_A_5WpE3FLY3_0(.din(n4723), .dout(n4726));
    jdff dff_A_hrAlhNAm1_0(.din(n4720), .dout(n4723));
    jdff dff_A_RkFR6puO5_0(.din(n4717), .dout(n4720));
    jdff dff_A_ve0cAdrm6_2(.din(n656), .dout(n4717));
    jdff dff_A_fvL8DYi59_0(.din(n4711), .dout(G24));
    jdff dff_A_65Oxlssu0_0(.din(n4708), .dout(n4711));
    jdff dff_A_O11JJmVx6_0(.din(n4705), .dout(n4708));
    jdff dff_A_KoVzu7q37_0(.din(n4702), .dout(n4705));
    jdff dff_A_FEyCJMKm5_0(.din(n4699), .dout(n4702));
    jdff dff_A_pFBbqCNZ4_0(.din(n4696), .dout(n4699));
    jdff dff_A_48L5gWb59_2(.din(n644), .dout(n4696));
    jdff dff_A_Woh6OdVs2_0(.din(n4690), .dout(G21));
    jdff dff_A_dVTLmbqY8_0(.din(n4687), .dout(n4690));
    jdff dff_A_QfYmXPBM9_0(.din(n4684), .dout(n4687));
    jdff dff_A_z5WKZ6gX1_0(.din(n4681), .dout(n4684));
    jdff dff_A_eJCCopJa8_0(.din(n4678), .dout(n4681));
    jdff dff_A_QqLKm64w6_0(.din(n4675), .dout(n4678));
    jdff dff_A_ZZdXydGm6_0(.din(n4672), .dout(n4675));
    jdff dff_A_s8rXBoX56_2(.din(n628), .dout(n4672));
    jdff dff_A_YLO0uwsg6_0(.din(n4666), .dout(G18));
    jdff dff_A_KptFUmx34_0(.din(n4663), .dout(n4666));
    jdff dff_A_LNaBgbuO0_0(.din(n4660), .dout(n4663));
    jdff dff_A_5a5NmolD0_0(.din(n4657), .dout(n4660));
    jdff dff_A_3gpJ598J6_0(.din(n4654), .dout(n4657));
    jdff dff_A_DzfdTRno5_0(.din(n4651), .dout(n4654));
    jdff dff_A_4MA2UY1h2_0(.din(n4648), .dout(n4651));
    jdff dff_A_YMIk41gS8_2(.din(n616), .dout(n4648));
    jdff dff_A_rSjKCHNd3_0(.din(n4642), .dout(G15));
    jdff dff_A_pXdMvCaZ5_0(.din(n4639), .dout(n4642));
    jdff dff_A_8IxNtXV07_0(.din(n4636), .dout(n4639));
    jdff dff_A_Zuo1Q2Tg7_0(.din(n4633), .dout(n4636));
    jdff dff_A_sjmTYC5l1_0(.din(n4630), .dout(n4633));
    jdff dff_A_jQHsaafC8_0(.din(n4627), .dout(n4630));
    jdff dff_A_sXNTBL0W1_0(.din(n4624), .dout(n4627));
    jdff dff_A_E06fr8vG6_2(.din(n608), .dout(n4624));
    jdff dff_A_B8RMUIgp3_0(.din(n4618), .dout(G48));
    jdff dff_A_rH4t5jcW6_0(.din(n4615), .dout(n4618));
    jdff dff_A_KXNZUKy93_0(.din(n4612), .dout(n4615));
    jdff dff_A_Y4lLNQqh1_0(.din(n4609), .dout(n4612));
    jdff dff_A_duzyz5qb1_0(.din(n4606), .dout(n4609));
    jdff dff_A_r50859xe3_0(.din(n4603), .dout(n4606));
    jdff dff_A_TwZMTknQ6_0(.din(n4600), .dout(n4603));
    jdff dff_A_CDdRnRdY1_2(.din(n581), .dout(n4600));
    jdff dff_A_BhoUwC8V8_0(.din(n4594), .dout(G45));
    jdff dff_A_srCUVw1T3_0(.din(n4591), .dout(n4594));
    jdff dff_A_XCrhnlh61_0(.din(n4588), .dout(n4591));
    jdff dff_A_zV37IviQ9_0(.din(n4585), .dout(n4588));
    jdff dff_A_Z6zVLBMN3_0(.din(n4582), .dout(n4585));
    jdff dff_A_MiuQvP6e8_0(.din(n4579), .dout(n4582));
    jdff dff_A_0CGTH1bS1_0(.din(n4576), .dout(n4579));
    jdff dff_A_R0NrbBNi0_2(.din(n569), .dout(n4576));
    jdff dff_A_APq4wjnn3_0(.din(n4570), .dout(G30));
    jdff dff_A_7jMzdGF19_0(.din(n4567), .dout(n4570));
    jdff dff_A_L0YRChQu4_0(.din(n4564), .dout(n4567));
    jdff dff_A_46LN5FKU6_0(.din(n4561), .dout(n4564));
    jdff dff_A_W1YKKNVp8_0(.din(n4558), .dout(n4561));
    jdff dff_A_FBgM1fRJ7_0(.din(n4555), .dout(n4558));
    jdff dff_A_uHEe57WI6_0(.din(n4552), .dout(n4555));
    jdff dff_A_apRAkZg53_2(.din(n549), .dout(n4552));
    jdff dff_A_q9vckpvG5_0(.din(n4546), .dout(G12));
    jdff dff_A_odBtbIM31_0(.din(n4543), .dout(n4546));
    jdff dff_A_1vEWcUA41_0(.din(n4540), .dout(n4543));
    jdff dff_A_7arxUe0W1_0(.din(n4537), .dout(n4540));
    jdff dff_A_BWrBfszh5_0(.din(n4534), .dout(n4537));
    jdff dff_A_z5QkHR330_0(.din(n4531), .dout(n4534));
    jdff dff_A_HEvIMrhO8_0(.din(n4528), .dout(n4531));
    jdff dff_A_DlpRYtCa6_2(.din(n514), .dout(n4528));
    jdff dff_A_TRxK1wIw3_0(.din(n4522), .dout(G9));
    jdff dff_A_6uNN18sl4_0(.din(n4519), .dout(n4522));
    jdff dff_A_UtqTR2KL3_0(.din(n4516), .dout(n4519));
    jdff dff_A_he6nAg600_0(.din(n4513), .dout(n4516));
    jdff dff_A_e86XZncz6_0(.din(n4510), .dout(n4513));
    jdff dff_A_k0UDo0I42_0(.din(n4507), .dout(n4510));
    jdff dff_A_EiKuOHs69_0(.din(n4504), .dout(n4507));
    jdff dff_A_N02qW1yA7_2(.din(n498), .dout(n4504));
    jdff dff_A_d4RSwXSv6_0(.din(n4498), .dout(G6));
    jdff dff_A_0YMYoiDk5_0(.din(n4495), .dout(n4498));
    jdff dff_A_KyyL9Txj4_0(.din(n4492), .dout(n4495));
    jdff dff_A_Eq74QE4D7_0(.din(n4489), .dout(n4492));
    jdff dff_A_987J6CRB3_0(.din(n4486), .dout(n4489));
    jdff dff_A_8USHUJhp6_0(.din(n4483), .dout(n4486));
    jdff dff_A_XU688eYr5_0(.din(n4480), .dout(n4483));
    jdff dff_A_y0S1Air87_2(.din(n478), .dout(n4480));
    jdff dff_A_bHBPXyAM6_0(.din(n4474), .dout(G3));
    jdff dff_A_ujBRfDho2_0(.din(n4471), .dout(n4474));
    jdff dff_A_GI9QouZV0_0(.din(n4468), .dout(n4471));
    jdff dff_A_dpkeVIAL3_0(.din(n4465), .dout(n4468));
    jdff dff_A_OQIf7Pgw2_0(.din(n4462), .dout(n4465));
    jdff dff_A_fve125FU0_0(.din(n4459), .dout(n4462));
    jdff dff_A_SMnVsTUa9_0(.din(n4456), .dout(n4459));
    jdff dff_A_MwqRsx0w6_2(.din(n443), .dout(n4456));
    jdff dff_B_rfC0uYMu3_3(.din(G952), .dout(n4454));
    jdff dff_A_9rtk9RnC4_2(.din(n4454), .dout(n4450));
    jdff dff_A_fyg1Pvi90_1(.din(n4454), .dout(n4447));
    jdff dff_A_Y3lDFskQ4_1(.din(n4447), .dout(n4444));
    jdff dff_A_xR0wmvLR0_1(.din(n4444), .dout(n4441));
    jdff dff_A_dI8Hm2Kf7_1(.din(n4441), .dout(n4438));
    jdff dff_A_56Wg1G6r6_1(.din(n4438), .dout(n4435));
    jdff dff_A_lqCeg8BL0_1(.din(n4435), .dout(n4432));
    jdff dff_A_DNaSOExD5_1(.din(n4432), .dout(n4429));
    jdff dff_A_PE3lYjSi0_1(.din(n4429), .dout(n4426));
    jdff dff_A_rBR9K8g67_1(.din(n4426), .dout(n4423));
    jdff dff_A_oxWsyVxS3_1(.din(n4423), .dout(n4420));
    jdff dff_A_L04gicix8_1(.din(n4420), .dout(n4417));
    jdff dff_A_Bcs8i3FC8_1(.din(n4417), .dout(n4414));
    jdff dff_A_KbNwem6D8_1(.din(n4414), .dout(n4411));
    jdff dff_A_q5XNO7724_1(.din(n4411), .dout(n4408));
    jdff dff_A_kB4SSVFo8_1(.din(n4408), .dout(n4405));
    jdff dff_A_eJ8WeTly5_1(.din(n4405), .dout(n4402));
    jdff dff_A_TcigiV841_2(.din(G953), .dout(n4399));
    jdff dff_A_BnUQP51w1_2(.din(n4399), .dout(n4396));
    jdff dff_A_lFjUfkaK7_2(.din(n4396), .dout(n4393));
    jdff dff_A_9q7KrHWp5_2(.din(n4393), .dout(n4390));
    jdff dff_A_QKLFT9Vj5_2(.din(n4390), .dout(n4387));
    jdff dff_A_KObVYEQX8_2(.din(n4387), .dout(n4384));
    jdff dff_A_i8Bpewt29_2(.din(n4384), .dout(n4381));
    jdff dff_A_41mZbeXE9_2(.din(n4381), .dout(n4378));
    jdff dff_A_NVQNUgLU8_2(.din(n4378), .dout(n4375));
    jdff dff_A_CtgLOVyt6_2(.din(n4375), .dout(n4372));
    jdff dff_A_lF46ez6K4_2(.din(n4372), .dout(n4369));
    jdff dff_A_6a1B3lW21_2(.din(n4369), .dout(n4366));
    jdff dff_A_BLAfd50W6_2(.din(n4366), .dout(n4363));
    jdff dff_A_bbIVZ2GE6_2(.din(n4363), .dout(n4360));
    jdff dff_A_8MQaLwTx7_2(.din(n4360), .dout(n4357));
    jdff dff_A_6Rsph3Hg4_1(.din(G953), .dout(n4354));
    jdff dff_A_wUT6urke0_1(.din(n4354), .dout(n4351));
    jdff dff_A_BVOeA0sq0_1(.din(n4351), .dout(n4348));
    jdff dff_A_kyiRyx2l1_1(.din(n4348), .dout(n4345));
    jdff dff_A_Bi0O1SEm3_1(.din(n4345), .dout(n4342));
    jdff dff_A_NAHX9de54_1(.din(n4342), .dout(n4339));
    jdff dff_A_TMAstcUh7_1(.din(n4339), .dout(n4336));
    jdff dff_A_essMvL466_1(.din(n4336), .dout(n4333));
    jdff dff_A_boM86YGm1_1(.din(n4333), .dout(n4330));
    jdff dff_A_QPQ4pMGT8_1(.din(n4330), .dout(n4327));
    jdff dff_A_JPs7umaD0_1(.din(n4327), .dout(n4324));
    jdff dff_A_dsLaRl0i4_1(.din(n4324), .dout(n4321));
    jdff dff_A_j20f81iP6_0(.din(G953), .dout(n4318));
    jdff dff_A_3qGi0CTf2_0(.din(n4318), .dout(n4315));
    jdff dff_A_EUiMTc6g9_0(.din(n4315), .dout(n4312));
    jdff dff_A_jZCOVcyN5_0(.din(n4312), .dout(n4309));
    jdff dff_A_U89RAlI01_0(.din(n4309), .dout(n4306));
    jdff dff_A_5uLjN7M02_0(.din(n4306), .dout(n4303));
    jdff dff_A_PTOOPFEP7_0(.din(n4303), .dout(n4300));
    jdff dff_A_cmziJ8rH0_0(.din(n4300), .dout(n4297));
    jdff dff_A_noxCN2xs0_0(.din(n4297), .dout(n4294));
    jdff dff_A_dnb0bL5J6_0(.din(n4294), .dout(n4291));
    jdff dff_A_1JkvPatN8_0(.din(n4291), .dout(n4288));
    jdff dff_A_0iwGuBup5_0(.din(n4288), .dout(n4285));
    jdff dff_A_tPvQ50N17_0(.din(n4285), .dout(n4282));
    jdff dff_B_KUG64qFo9_0(.din(n859), .dout(n1949));
    jdff dff_B_394Fxekk6_0(.din(n1949), .dout(n1952));
    jdff dff_B_alWpnuZ68_0(.din(n1952), .dout(n1955));
    jdff dff_B_flIMqsTO9_0(.din(n1955), .dout(n1958));
    jdff dff_B_X1XwYjW90_0(.din(n1958), .dout(n1961));
    jdff dff_B_oCKmzzRJ2_0(.din(n827), .dout(n1964));
    jdff dff_B_HucuwSJG9_0(.din(n1964), .dout(n1967));
    jdff dff_B_eggdHZDG6_0(.din(n807), .dout(n1970));
    jdff dff_A_IG0CL64y6_0(.din(n1975), .dout(n1972));
    jdff dff_A_v3ni466f3_0(.din(n803), .dout(n1975));
    jdff dff_B_k5gOsM257_0(.din(n799), .dout(n1979));
    jdff dff_B_JBz7l3hc8_0(.din(n1979), .dout(n1982));
    jdff dff_B_hT1JvqQo9_0(.din(n783), .dout(n1985));
    jdff dff_B_QTJGx9Zi8_0(.din(n1985), .dout(n1988));
    jdff dff_B_E3zHyqyO6_0(.din(n1988), .dout(n1991));
    jdff dff_B_8UVV9BKq0_1(.din(n911), .dout(n1994));
    jdff dff_B_Lvpku14t8_1(.din(n914), .dout(n1997));
    jdff dff_B_dvRgyTWL3_1(.din(n1997), .dout(n2000));
    jdff dff_B_f3V5GFWe6_1(.din(n2000), .dout(n2003));
    jdff dff_B_w1ZBE5So9_1(.din(n2003), .dout(n2006));
    jdff dff_B_D6vUSOhQ9_1(.din(n2006), .dout(n2009));
    jdff dff_B_wo1dfjjy0_1(.din(n2009), .dout(n2012));
    jdff dff_B_HxB01BHw8_1(.din(n2012), .dout(n2015));
    jdff dff_B_LP0n0gDD2_1(.din(n2015), .dout(n2018));
    jdff dff_B_j5g1Z4K63_1(.din(n2018), .dout(n2021));
    jdff dff_B_nOi7yzSc6_1(.din(n2021), .dout(n2024));
    jdff dff_B_XY4RlwRU3_1(.din(n2024), .dout(n2027));
    jdff dff_B_oVS34vDx7_0(.din(n1171), .dout(n2030));
    jdff dff_B_s2iS1UZf1_0(.din(n2030), .dout(n2033));
    jdff dff_B_Km60sTcO5_0(.din(n2033), .dout(n2036));
    jdff dff_B_7cITet7p8_0(.din(n2036), .dout(n2039));
    jdff dff_B_aJLU51O03_0(.din(n2039), .dout(n2042));
    jdff dff_B_8yblqgjN8_0(.din(n2042), .dout(n2045));
    jdff dff_B_GPNNfbOx8_0(.din(n2045), .dout(n2048));
    jdff dff_B_h0NNqSV74_0(.din(n2048), .dout(n2051));
    jdff dff_B_FmKeF8Sd9_0(.din(n2051), .dout(n2054));
    jdff dff_B_A9yugYQe2_0(.din(n2054), .dout(n2057));
    jdff dff_B_CNdE24Io0_0(.din(n2057), .dout(n2060));
    jdff dff_B_9UvZ2llQ9_0(.din(n2060), .dout(n2063));
    jdff dff_B_f547bRLo4_0(.din(n2063), .dout(n2066));
    jdff dff_B_U4qzGoUC9_0(.din(n2066), .dout(n2069));
    jdff dff_A_XxGbtZY94_1(.din(n2074), .dout(n2071));
    jdff dff_A_I3PxFMEP5_1(.din(n2077), .dout(n2074));
    jdff dff_A_TGFYP5zS4_1(.din(n2080), .dout(n2077));
    jdff dff_A_2ZW7aQZH7_1(.din(n2083), .dout(n2080));
    jdff dff_A_pLuSHK438_1(.din(n2086), .dout(n2083));
    jdff dff_A_crK3MAGE6_1(.din(n2089), .dout(n2086));
    jdff dff_A_QKwrXAwl5_1(.din(n2092), .dout(n2089));
    jdff dff_A_kmB8DmzN6_1(.din(n2095), .dout(n2092));
    jdff dff_A_X7vahN7m6_1(.din(n2098), .dout(n2095));
    jdff dff_A_aohLhlQ79_1(.din(n2101), .dout(n2098));
    jdff dff_A_RYgo71xN7_1(.din(n2104), .dout(n2101));
    jdff dff_A_DGTpZgc44_1(.din(n2107), .dout(n2104));
    jdff dff_A_k12CDglC2_1(.din(n2110), .dout(n2107));
    jdff dff_A_l53IoIuA6_1(.din(n2113), .dout(n2110));
    jdff dff_A_gLLZy1pU5_1(.din(n903), .dout(n2113));
    jdff dff_A_syXOUwlA2_1(.din(n2119), .dout(n2116));
    jdff dff_A_vuuSfQjb4_1(.din(n2122), .dout(n2119));
    jdff dff_A_z7TEBZSF4_1(.din(n2125), .dout(n2122));
    jdff dff_A_p3pKopkY3_1(.din(n2128), .dout(n2125));
    jdff dff_A_FGhfCPHc4_1(.din(n2131), .dout(n2128));
    jdff dff_A_dp7rQfin0_1(.din(n2134), .dout(n2131));
    jdff dff_A_pHGEWigZ7_1(.din(n2137), .dout(n2134));
    jdff dff_A_A9Mpn6Mo7_1(.din(n2140), .dout(n2137));
    jdff dff_A_vEDHGsRF1_1(.din(n2143), .dout(n2140));
    jdff dff_A_wke8CEi98_1(.din(n2146), .dout(n2143));
    jdff dff_A_Hi8O8vN88_1(.din(n2149), .dout(n2146));
    jdff dff_A_kt91S0nH0_1(.din(n2152), .dout(n2149));
    jdff dff_A_mFka8xG79_1(.din(n2155), .dout(n2152));
    jdff dff_A_GmsY3EdE6_1(.din(n2158), .dout(n2155));
    jdff dff_A_AXsYIj0G3_1(.din(n2161), .dout(n2158));
    jdff dff_A_QVseP5Xn5_1(.din(n2164), .dout(n2161));
    jdff dff_A_TYWhiCcb1_1(.din(G902), .dout(n2164));
    jdff dff_A_iGmSLGYQ0_2(.din(n2170), .dout(n2167));
    jdff dff_A_JNDw6oqa7_2(.din(n2173), .dout(n2170));
    jdff dff_A_F7AUvBLO4_2(.din(n2176), .dout(n2173));
    jdff dff_A_v3Az2e4l6_2(.din(n2179), .dout(n2176));
    jdff dff_A_ShRa6vIr0_2(.din(n2182), .dout(n2179));
    jdff dff_A_7ucS4sL53_2(.din(n2185), .dout(n2182));
    jdff dff_A_YPE5SCWC0_2(.din(n2188), .dout(n2185));
    jdff dff_A_QzBMqiCV4_2(.din(n2191), .dout(n2188));
    jdff dff_A_zOufd4Aa8_2(.din(n2194), .dout(n2191));
    jdff dff_A_T2uI2d8G1_2(.din(n2197), .dout(n2194));
    jdff dff_A_ayxp7PCQ1_2(.din(n2200), .dout(n2197));
    jdff dff_A_2KVwM7VM7_2(.din(n2203), .dout(n2200));
    jdff dff_A_GnsqHrad7_2(.din(n2206), .dout(n2203));
    jdff dff_A_ToUJgmBh8_2(.din(n2209), .dout(n2206));
    jdff dff_A_5YD3cgRK2_2(.din(n2212), .dout(n2209));
    jdff dff_A_mDqaywDU7_2(.din(n2215), .dout(n2212));
    jdff dff_A_WXr3mAOY7_2(.din(G902), .dout(n2215));
    jdff dff_A_fX4U4ovf9_0(.din(n4274), .dout(n2218));
    jdff dff_A_cMFoa89n8_1(.din(n4274), .dout(n2221));
    jdff dff_B_hGOzfkvM9_1(.din(n1223), .dout(n2225));
    jdff dff_B_YURzaCoG9_1(.din(n2225), .dout(n2228));
    jdff dff_B_5LsUcDqb1_1(.din(n2228), .dout(n2231));
    jdff dff_B_lWogwtJi2_1(.din(n2231), .dout(n2234));
    jdff dff_B_8Hz62FqG2_1(.din(n2234), .dout(n2237));
    jdff dff_B_vFUmr7hp3_1(.din(n2237), .dout(n2240));
    jdff dff_B_J5luUa8b5_1(.din(n2240), .dout(n2243));
    jdff dff_B_drqsJAl31_1(.din(n2243), .dout(n2246));
    jdff dff_B_aiC7ouoZ6_1(.din(n2246), .dout(n2249));
    jdff dff_B_WNGVCYfI7_1(.din(n2249), .dout(n2252));
    jdff dff_B_0XerGWij3_1(.din(n2252), .dout(n2255));
    jdff dff_B_8QhtpKir0_1(.din(n2255), .dout(n2258));
    jdff dff_B_UX1OY6Gb2_0(.din(n1235), .dout(n2261));
    jdff dff_B_QpE7LmeA5_0(.din(n2261), .dout(n2264));
    jdff dff_B_FbnBAdS51_0(.din(n2264), .dout(n2267));
    jdff dff_B_w35X5nWO4_0(.din(n2267), .dout(n2270));
    jdff dff_B_w41uq7435_0(.din(n2270), .dout(n2273));
    jdff dff_B_3mQRfDGC9_0(.din(n2273), .dout(n2276));
    jdff dff_B_86QDvtdV9_0(.din(n2276), .dout(n2279));
    jdff dff_B_HeISs4qd9_0(.din(n2279), .dout(n2282));
    jdff dff_B_YxJ0zRfD3_0(.din(n2282), .dout(n2285));
    jdff dff_B_vvhr6LsZ4_0(.din(n2285), .dout(n2288));
    jdff dff_B_240jvMa60_0(.din(n2288), .dout(n2291));
    jdff dff_B_HAqUgjKD2_0(.din(n2291), .dout(n2294));
    jdff dff_B_0o4YFTJ35_0(.din(n2294), .dout(n2297));
    jdff dff_B_uSiNie2K1_0(.din(n2297), .dout(n2300));
    jdff dff_B_xxqWYu090_1(.din(n1011), .dout(n2303));
    jdff dff_B_gJdEHobR1_1(.din(n1019), .dout(n2306));
    jdff dff_B_o1k8CBxA6_1(.din(n945), .dout(n2309));
    jdff dff_B_BvqV64tH2_1(.din(n964), .dout(n2312));
    jdff dff_B_i6qCSWfC6_2(.din(n992), .dout(n2315));
    jdff dff_A_ABtNJUFx6_1(.din(n2443), .dout(n2317));
    jdff dff_B_K6u4Fd705_2(.din(n921), .dout(n2321));
    jdff dff_A_DoAoh6qP1_2(.din(n2326), .dout(n2323));
    jdff dff_A_bGwVcjBD4_2(.din(n2333), .dout(n2326));
    jdff dff_B_OqorBsIl3_3(.din(n917), .dout(n2330));
    jdff dff_B_sb9iZ8bG2_3(.din(n2330), .dout(n2333));
    jdff dff_B_VkBUUOFb5_0(.din(n1267), .dout(n2336));
    jdff dff_B_wIc1UPH12_0(.din(n2336), .dout(n2339));
    jdff dff_B_VQ2fVj6Q2_0(.din(n2339), .dout(n2342));
    jdff dff_B_z823ZQ8i2_0(.din(n2342), .dout(n2345));
    jdff dff_B_CKP56xHB2_0(.din(n2345), .dout(n2348));
    jdff dff_B_Xx7E4TlV7_0(.din(n2348), .dout(n2351));
    jdff dff_B_mHbSeaVo7_0(.din(n2351), .dout(n2354));
    jdff dff_B_PygfWZwp8_0(.din(n2354), .dout(n2357));
    jdff dff_B_eh4kMKeL8_0(.din(n2357), .dout(n2360));
    jdff dff_B_WZiz5vdx3_0(.din(n2360), .dout(n2363));
    jdff dff_B_G6Pc5LI60_0(.din(n2363), .dout(n2366));
    jdff dff_B_WGDz4yIs8_0(.din(n2366), .dout(n2369));
    jdff dff_B_lXOg0ONp7_0(.din(n1255), .dout(n2372));
    jdff dff_B_vBaRG9Ml8_0(.din(n2372), .dout(n2375));
    jdff dff_B_C5LRueNP1_0(.din(n2375), .dout(n2378));
    jdff dff_B_d6aTAMLa3_0(.din(n2378), .dout(n2381));
    jdff dff_B_Jho5Yf9L0_0(.din(n2381), .dout(n2384));
    jdff dff_B_jrfgMv3B0_0(.din(n2384), .dout(n2387));
    jdff dff_B_M7QJVnjF3_0(.din(n2387), .dout(n2390));
    jdff dff_B_rWpQweSu9_0(.din(n2390), .dout(n2393));
    jdff dff_B_9a3Fue1j0_0(.din(n2393), .dout(n2396));
    jdff dff_B_Mklt5Ah61_0(.din(n2396), .dout(n2399));
    jdff dff_B_PuUswaoM0_0(.din(n2399), .dout(n2402));
    jdff dff_B_bHWz2Acr8_0(.din(n2402), .dout(n2405));
    jdff dff_B_WPzS1h6Y7_0(.din(n2405), .dout(n2408));
    jdff dff_B_ai9z8Ib93_0(.din(n2408), .dout(n2411));
    jdff dff_B_l8DfnSgd7_1(.din(n1105), .dout(n2414));
    jdff dff_B_slj6ZFIj6_1(.din(n1124), .dout(n2417));
    jdff dff_B_JQNBt3Tw0_1(.din(n1132), .dout(n2420));
    jdff dff_A_AlG92Tz52_1(.din(n933), .dout(n2422));
    jdff dff_A_WANtlcxU1_2(.din(n933), .dout(n2425));
    jdff dff_A_nJmoAc6P5_1(.din(n2431), .dout(n2428));
    jdff dff_A_Mfurm3pw8_1(.din(n2434), .dout(n2431));
    jdff dff_A_1yr2Fkib6_1(.din(n839), .dout(n2434));
    jdff dff_A_FPGOcCb08_2(.din(n839), .dout(n2437));
    jdff dff_A_82Ol37eH4_1(.din(n953), .dout(n2440));
    jdff dff_A_3sTCNM3y5_0(.din(n968), .dout(n2443));
    jdff dff_A_aVPtgSo02_2(.din(n968), .dout(n2446));
    jdff dff_A_Hp3hdCfF5_0(.din(n1089), .dout(n2449));
    jdff dff_A_lGq66MbF9_1(.din(n2456), .dout(n2452));
    jdff dff_B_hFGawRW00_2(.din(n1015), .dout(n2456));
    jdff dff_A_33pc2Raq6_0(.din(n1031), .dout(n2458));
    jdff dff_A_wTKLKhEd4_2(.din(n1031), .dout(n2461));
    jdff dff_A_gmOYxxun3_0(.din(n2474), .dout(n2464));
    jdff dff_A_WSLk10X92_2(.din(n2474), .dout(n2467));
    jdff dff_B_YpyyUZvx8_3(.din(n1069), .dout(n2471));
    jdff dff_B_6OB8wPMk2_3(.din(n2471), .dout(n2474));
    jdff dff_A_cCQcj4iH3_1(.din(n1066), .dout(n2476));
    jdff dff_A_2sTvlTIs9_2(.din(n1066), .dout(n2479));
    jdff dff_B_9j5Z6XY35_0(.din(n1275), .dout(n2483));
    jdff dff_B_To039hLW4_0(.din(n2483), .dout(n2486));
    jdff dff_B_qS0RVbv06_0(.din(n2486), .dout(n2489));
    jdff dff_B_QMmS2fVF6_0(.din(n2489), .dout(n2492));
    jdff dff_B_XWojwD808_0(.din(n2492), .dout(n2495));
    jdff dff_B_wRxdAre98_0(.din(n2495), .dout(n2498));
    jdff dff_B_1bIDSDbp4_0(.din(n2498), .dout(n2501));
    jdff dff_B_z32MSyet2_0(.din(n2501), .dout(n2504));
    jdff dff_B_toAuobQO5_0(.din(n2504), .dout(n2507));
    jdff dff_B_nTDLVa0Y5_0(.din(n2507), .dout(n2510));
    jdff dff_B_C2Wt8arC7_0(.din(n2510), .dout(n2513));
    jdff dff_B_jPLi9S8P9_0(.din(n2513), .dout(n2516));
    jdff dff_B_jzpWERoA1_0(.din(n2516), .dout(n2519));
    jdff dff_B_o3xNFRU61_0(.din(n2519), .dout(n2522));
    jdff dff_B_GVXrhrtJ9_0(.din(n2522), .dout(n2525));
    jdff dff_A_cxbLVBeD5_1(.din(n2530), .dout(n2527));
    jdff dff_A_HVcZbEPt6_1(.din(n2533), .dout(n2530));
    jdff dff_A_uD3aOx0V1_1(.din(n2536), .dout(n2533));
    jdff dff_A_mOpspPGk4_1(.din(n2539), .dout(n2536));
    jdff dff_A_WqcpWQGw2_1(.din(n2542), .dout(n2539));
    jdff dff_A_10g0eqLL5_1(.din(n2545), .dout(n2542));
    jdff dff_A_mNwDuFKi5_1(.din(n2548), .dout(n2545));
    jdff dff_A_6qXO61xc4_1(.din(n2551), .dout(n2548));
    jdff dff_A_fpPIGJVJ4_1(.din(n2554), .dout(n2551));
    jdff dff_A_ntxM5n5S8_1(.din(n2557), .dout(n2554));
    jdff dff_A_6kRSMX3n4_1(.din(n2560), .dout(n2557));
    jdff dff_A_GShpcJh22_1(.din(n2563), .dout(n2560));
    jdff dff_A_NJQ70hQm1_1(.din(n2566), .dout(n2563));
    jdff dff_A_OgvA04eG7_1(.din(n2569), .dout(n2566));
    jdff dff_A_pQFwUsRx7_1(.din(n2572), .dout(n2569));
    jdff dff_A_9JcezBKN5_1(.din(n2575), .dout(n2572));
    jdff dff_A_eveR7xjG5_1(.din(G902), .dout(n2575));
    jdff dff_A_R0P7A7Oe4_2(.din(n2581), .dout(n2578));
    jdff dff_A_doPstua32_2(.din(n2584), .dout(n2581));
    jdff dff_A_IaklNWCl1_2(.din(n2587), .dout(n2584));
    jdff dff_A_vl8SOYU20_2(.din(n2590), .dout(n2587));
    jdff dff_A_OOXBT9eP7_2(.din(n2593), .dout(n2590));
    jdff dff_A_LSOiE9oF1_2(.din(n2596), .dout(n2593));
    jdff dff_A_0UcrAbvE0_2(.din(n2599), .dout(n2596));
    jdff dff_A_ULUrvKIz6_2(.din(n2602), .dout(n2599));
    jdff dff_A_XUxngNkg4_2(.din(n2605), .dout(n2602));
    jdff dff_A_Sj6X3e9V5_2(.din(n2608), .dout(n2605));
    jdff dff_A_Xg6o16VL7_2(.din(n2611), .dout(n2608));
    jdff dff_A_YDDeoh0r5_2(.din(n2614), .dout(n2611));
    jdff dff_A_VtmdS7t47_2(.din(n2617), .dout(n2614));
    jdff dff_A_fIZEEFDX0_2(.din(n2620), .dout(n2617));
    jdff dff_A_SkIp3MHM6_2(.din(n2623), .dout(n2620));
    jdff dff_A_C32Ed3NP0_2(.din(n2626), .dout(n2623));
    jdff dff_A_9vXg7p2U9_2(.din(G902), .dout(n2626));
    jdff dff_B_RqHLDa1b8_1(.din(n751), .dout(n2630));
    jdff dff_B_JC95DaZ65_1(.din(n755), .dout(n2633));
    jdff dff_A_1VRB2xs14_0(.din(n545), .dout(n2635));
    jdff dff_A_szBFXo8J3_1(.din(n541), .dout(n2638));
    jdff dff_A_BsJ2jOKO4_2(.din(n541), .dout(n2641));
    jdff dff_A_qvlnoTIO5_0(.din(n671), .dout(n2644));
    jdff dff_A_zlZRoQlY1_2(.din(n671), .dout(n2647));
    jdff dff_B_PzhPMEus9_0(.din(n659), .dout(n2651));
    jdff dff_B_dkcwcKti5_0(.din(n2651), .dout(n2654));
    jdff dff_B_2muhCsUb1_0(.din(n2654), .dout(n2657));
    jdff dff_A_ZJtyRA0T1_1(.din(n577), .dout(n2659));
    jdff dff_A_CRco7veP1_0(.din(n573), .dout(n2662));
    jdff dff_A_dKrVgv1U3_2(.din(n573), .dout(n2665));
    jdff dff_A_jElLZGmm8_1(.din(n2671), .dout(n2668));
    jdff dff_A_3CCsnjzW2_0(.din(n2674), .dout(n2671));
    jdff dff_A_19G8xX9t3_0(.din(n2677), .dout(n2674));
    jdff dff_A_EwZWUKIS7_0(.din(n537), .dout(n2677));
    jdff dff_A_pmbcomq20_2(.din(n2683), .dout(n2680));
    jdff dff_A_9S237OTl6_2(.din(n2686), .dout(n2683));
    jdff dff_A_8pmT6EMg5_2(.din(n2689), .dout(n2686));
    jdff dff_A_eHRBrCIQ1_2(.din(n537), .dout(n2689));
    jdff dff_A_Xv4Re0VA8_0(.din(n529), .dout(n2692));
    jdff dff_A_Cpn0gaCa7_1(.din(G900), .dout(n2695));
    jdff dff_A_gPnpAazZ3_1(.din(n518), .dout(n2698));
    jdff dff_A_ZwXfHhEL8_2(.din(n518), .dout(n2701));
    jdff dff_A_WjCKIAiK5_0(.din(n510), .dout(n2704));
    jdff dff_A_DTPDCWCH0_1(.din(n2711), .dout(n2707));
    jdff dff_B_vDF4uLgW4_2(.din(n506), .dout(n2711));
    jdff dff_A_yPVhSkGV2_1(.din(n2716), .dout(n2713));
    jdff dff_A_oqBjpYYL8_1(.din(n604), .dout(n2716));
    jdff dff_A_2ypsFFp70_0(.din(n596), .dout(n2719));
    jdff dff_B_L2sw5HXi6_2(.din(n490), .dout(n2723));
    jdff dff_A_REp22pjD7_2(.din(n2728), .dout(n2725));
    jdff dff_A_zT089Ygc2_2(.din(n2731), .dout(n2728));
    jdff dff_A_3b8lsqOb6_2(.din(n2734), .dout(n2731));
    jdff dff_A_SWInxcw56_2(.din(n427), .dout(n2734));
    jdff dff_B_MRaEe7G13_1(.din(n381), .dout(n2738));
    jdff dff_B_2bzhOtmf4_1(.din(n2738), .dout(n2741));
    jdff dff_B_OZ6XhuiB2_1(.din(n2741), .dout(n2744));
    jdff dff_B_S3yyGRCa6_1(.din(n2744), .dout(n2747));
    jdff dff_B_4GcJj6UK9_1(.din(n2747), .dout(n2750));
    jdff dff_A_jeviynMh1_1(.din(n2755), .dout(n2752));
    jdff dff_A_Goheoi8v6_1(.din(n193), .dout(n2755));
    jdff dff_A_UUI63NDL8_1(.din(n193), .dout(n2758));
    jdff dff_A_Zo59uV6y7_2(.din(n193), .dout(n2761));
    jdff dff_A_dgHihsKT6_0(.din(n474), .dout(n2764));
    jdff dff_A_AE1D2ZU45_1(.din(n470), .dout(n2767));
    jdff dff_A_znOEPE3t7_2(.din(n470), .dout(n2770));
    jdff dff_B_5nsrbSC05_1(.din(n342), .dout(n2774));
    jdff dff_B_OPIO8SGq4_1(.din(n2774), .dout(n2777));
    jdff dff_B_UnXNkBs69_1(.din(n2777), .dout(n2780));
    jdff dff_B_pkG8ZWhz3_1(.din(n2780), .dout(n2783));
    jdff dff_B_kbcpQt2j9_1(.din(n2783), .dout(n2786));
    jdff dff_A_NAtrOi5y4_1(.din(n305), .dout(n2788));
    jdff dff_A_6Mu5TVS08_0(.din(n640), .dout(n2791));
    jdff dff_A_ESbhtxXb4_1(.din(n596), .dout(n2794));
    jdff dff_B_k6APoGJQ8_1(.din(n584), .dout(n2798));
    jdff dff_B_DS7aIEQu2_1(.din(n2798), .dout(n2801));
    jdff dff_B_h9cOKgaC6_1(.din(n2801), .dout(n2804));
    jdff dff_B_xn4tmahP4_1(.din(n2804), .dout(n2807));
    jdff dff_B_NsDCSFXi4_1(.din(n2807), .dout(n2810));
    jdff dff_A_zDABCEQv4_0(.din(n2815), .dout(n2812));
    jdff dff_A_IwDaN4mS1_0(.din(n2818), .dout(n2815));
    jdff dff_A_Ep1bIAFe4_0(.din(n2821), .dout(n2818));
    jdff dff_A_nmWGtdch3_0(.din(n2824), .dout(n2821));
    jdff dff_A_B7fuyqWW3_0(.din(n2827), .dout(n2824));
    jdff dff_A_nUzh37dZ2_0(.din(n2830), .dout(n2827));
    jdff dff_A_EJl3uVnT3_0(.din(n2833), .dout(n2830));
    jdff dff_A_DyOqZUPQ7_0(.din(n2836), .dout(n2833));
    jdff dff_A_4kAObYLq2_0(.din(n2839), .dout(n2836));
    jdff dff_A_1ggNEJ7t1_0(.din(n2842), .dout(n2839));
    jdff dff_A_U73lyVPM5_0(.din(n2845), .dout(n2842));
    jdff dff_A_tQh4oj1H7_0(.din(n2848), .dout(n2845));
    jdff dff_A_tqndhuCu4_0(.din(n289), .dout(n2848));
    jdff dff_A_EQkrYTW60_1(.din(G227), .dout(n2851));
    jdff dff_A_Nep6uVWh4_0(.din(n2857), .dout(n2854));
    jdff dff_A_i7U0X4g38_0(.din(n2860), .dout(n2857));
    jdff dff_A_N29Ib9Xp6_0(.din(n2863), .dout(n2860));
    jdff dff_A_iatluKOH0_0(.din(n2866), .dout(n2863));
    jdff dff_A_nxfbMlCP2_0(.din(n2869), .dout(n2866));
    jdff dff_A_oDForQPh5_0(.din(n2872), .dout(n2869));
    jdff dff_A_Z6J848JK0_0(.din(n2875), .dout(n2872));
    jdff dff_A_fpR1vrs22_0(.din(n2878), .dout(n2875));
    jdff dff_A_jIcyLV9S1_0(.din(n2881), .dout(n2878));
    jdff dff_A_BDCUAhlO5_0(.din(n2884), .dout(n2881));
    jdff dff_A_IP1JPemf0_0(.din(n2887), .dout(n2884));
    jdff dff_A_kDqQp4wh2_0(.din(n2890), .dout(n2887));
    jdff dff_A_zoEEl4xc9_0(.din(n2893), .dout(n2890));
    jdff dff_A_MMQqbunt0_0(.din(n2896), .dout(n2893));
    jdff dff_A_NUweUMAO7_0(.din(n2899), .dout(n2896));
    jdff dff_A_HvlivWmk0_0(.din(G469), .dout(n2899));
    jdff dff_A_r5oBXoY02_2(.din(n2905), .dout(n2902));
    jdff dff_A_Fe6t2XlX6_2(.din(n2908), .dout(n2905));
    jdff dff_A_wWIJ0g4Y4_2(.din(n2911), .dout(n2908));
    jdff dff_A_YmUIaqRu3_2(.din(n2914), .dout(n2911));
    jdff dff_A_hDwbYA1M4_2(.din(n2917), .dout(n2914));
    jdff dff_A_ULtBYnlK8_2(.din(G469), .dout(n2917));
    jdff dff_A_sjWVkpVN1_1(.din(n2923), .dout(n2920));
    jdff dff_A_kHyHxSiA5_1(.din(n269), .dout(n2923));
    jdff dff_A_HtiQBFxH9_2(.din(n2929), .dout(n2926));
    jdff dff_A_wQPGfbPQ3_2(.din(n269), .dout(n2929));
    jdff dff_A_OU8Ehhts9_1(.din(n2935), .dout(n2932));
    jdff dff_A_aYi1miGV4_1(.din(n2938), .dout(n2935));
    jdff dff_A_vI1tui6I2_1(.din(n266), .dout(n2938));
    jdff dff_A_tjuDygRx7_2(.din(n2944), .dout(n2941));
    jdff dff_A_Pe5pLhwT1_2(.din(n2947), .dout(n2944));
    jdff dff_A_zSeAZakS0_2(.din(n266), .dout(n2947));
    jdff dff_A_FLf3qhb67_1(.din(n2953), .dout(n2950));
    jdff dff_A_XnCSF2Rn3_1(.din(n2956), .dout(n2953));
    jdff dff_A_9E2EhCul1_1(.din(n2959), .dout(n2956));
    jdff dff_A_BPSgy5466_1(.din(n254), .dout(n2959));
    jdff dff_A_LYnqv5er8_0(.din(n2965), .dout(n2962));
    jdff dff_A_D7vO2Dl39_0(.din(n2968), .dout(n2965));
    jdff dff_A_v0qq9xQJ7_0(.din(n2971), .dout(n2968));
    jdff dff_A_oyVB0b665_0(.din(n2974), .dout(n2971));
    jdff dff_A_8XfYXIVT6_0(.din(n2977), .dout(n2974));
    jdff dff_A_FmUb1ebN6_0(.din(n2980), .dout(n2977));
    jdff dff_A_bOi4UE0B1_0(.din(n2983), .dout(n2980));
    jdff dff_A_Wj38kN3O5_0(.din(n2986), .dout(n2983));
    jdff dff_A_kCc9f4Ez3_0(.din(n2989), .dout(n2986));
    jdff dff_A_ym2UMXSd0_0(.din(n2992), .dout(n2989));
    jdff dff_A_PkLqv2Px5_0(.din(n2995), .dout(n2992));
    jdff dff_A_iQSMFodB5_0(.din(n2998), .dout(n2995));
    jdff dff_A_ASSNhaad5_0(.din(n246), .dout(n2998));
    jdff dff_B_aFnTQLtg1_1(.din(n234), .dout(n3002));
    jdff dff_A_x4CoadrC8_1(.din(G224), .dout(n3004));
    jdff dff_B_mpwLwhvW6_0(.din(n223), .dout(n3008));
    jdff dff_B_JxaDq2Ff9_0(.din(n3008), .dout(n3011));
    jdff dff_A_9dENtCRg6_0(.din(n215), .dout(n3013));
    jdff dff_A_TXUsMIO52_1(.din(n3019), .dout(n3016));
    jdff dff_A_4iQ5PsFD0_1(.din(n3032), .dout(n3019));
    jdff dff_A_SOb0HfFp1_2(.din(n3025), .dout(n3022));
    jdff dff_A_DyND0V2T2_2(.din(n3032), .dout(n3025));
    jdff dff_B_iZSNUWk79_3(.din(n204), .dout(n3029));
    jdff dff_B_sq9N4pXi0_3(.din(n3029), .dout(n3032));
    jdff dff_A_JQVYE69n0_0(.din(n3037), .dout(n3034));
    jdff dff_A_hZVR3lWF6_0(.din(n201), .dout(n3037));
    jdff dff_A_PIaYCAmj5_1(.din(n3043), .dout(n3040));
    jdff dff_A_wcBhESmt3_1(.din(n3046), .dout(n3043));
    jdff dff_A_m9EiKjWD6_1(.din(n3049), .dout(n3046));
    jdff dff_A_geY3g1Pp7_1(.din(n3052), .dout(n3049));
    jdff dff_A_4hau76MP3_1(.din(n201), .dout(n3052));
    jdff dff_A_ZJ1LG8BS8_2(.din(n3058), .dout(n3055));
    jdff dff_A_Mskq4TCj1_2(.din(n3061), .dout(n3058));
    jdff dff_A_laEriNyn6_2(.din(n3064), .dout(n3061));
    jdff dff_A_GrrdG6wv4_2(.din(n3067), .dout(n3064));
    jdff dff_A_woUgFLQV7_2(.din(n201), .dout(n3067));
    jdff dff_A_bZqGKQsJ5_1(.din(n3077), .dout(n3070));
    jdff dff_A_tUN8qgig9_2(.din(n3077), .dout(n3073));
    jdff dff_B_SmSmmBJM7_3(.din(n454), .dout(n3077));
    jdff dff_B_AYMGgiWa9_1(.din(n446), .dout(n3080));
    jdff dff_B_6H4SbxbY6_1(.din(n3080), .dout(n3083));
    jdff dff_B_yHm5oCLr0_1(.din(n3083), .dout(n3086));
    jdff dff_B_ZOuoeaeS6_1(.din(n3086), .dout(n3089));
    jdff dff_B_P7OwcfVU5_1(.din(n3089), .dout(n3092));
    jdff dff_A_kl9t13r57_0(.din(n3097), .dout(n3094));
    jdff dff_A_TNj0WbIB7_0(.din(n3100), .dout(n3097));
    jdff dff_A_U89xG9Vd2_0(.din(n3103), .dout(n3100));
    jdff dff_A_fuuvUbSH8_0(.din(n3106), .dout(n3103));
    jdff dff_A_slbVTk6q2_0(.din(n3109), .dout(n3106));
    jdff dff_A_G9t4kHd51_0(.din(n3112), .dout(n3109));
    jdff dff_A_2X9bSZv90_0(.din(n3115), .dout(n3112));
    jdff dff_A_NWg9P04g9_0(.din(n3118), .dout(n3115));
    jdff dff_A_clhh5mhz1_0(.din(n3121), .dout(n3118));
    jdff dff_A_qKPCwKQn3_0(.din(n3124), .dout(n3121));
    jdff dff_A_ruJATUgD2_0(.din(n3127), .dout(n3124));
    jdff dff_A_tU0QD92Y8_0(.din(n181), .dout(n3127));
    jdff dff_A_hB3DFJRv7_0(.din(n3133), .dout(n3130));
    jdff dff_A_4xVr9j2f6_0(.din(n3136), .dout(n3133));
    jdff dff_A_mjXoH1J22_0(.din(n3139), .dout(n3136));
    jdff dff_A_k6Pbvkn38_0(.din(n3142), .dout(n3139));
    jdff dff_A_SGzMnbvN2_0(.din(n3145), .dout(n3142));
    jdff dff_A_jwQz4vQy2_0(.din(n3148), .dout(n3145));
    jdff dff_A_AXm7U6Us4_0(.din(n3151), .dout(n3148));
    jdff dff_A_zAgb3OdD2_0(.din(n3154), .dout(n3151));
    jdff dff_A_2V1e7Wgg3_0(.din(n3157), .dout(n3154));
    jdff dff_A_vYQArisC2_0(.din(n3160), .dout(n3157));
    jdff dff_A_4blA1VWQ2_0(.din(n3163), .dout(n3160));
    jdff dff_A_mgyOkLTl1_0(.din(n3166), .dout(n3163));
    jdff dff_A_JB0utwUz8_0(.din(n3169), .dout(n3166));
    jdff dff_A_QrAafOiN1_0(.din(n3172), .dout(n3169));
    jdff dff_A_e7Eaff0f4_0(.din(n3175), .dout(n3172));
    jdff dff_A_VyrqZWlM8_0(.din(G210), .dout(n3175));
    jdff dff_A_2wciar0F4_1(.din(G210), .dout(n3178));
    jdff dff_A_eFk3xNBu3_0(.din(n3184), .dout(n3181));
    jdff dff_A_pXDpby4W7_0(.din(n3187), .dout(n3184));
    jdff dff_A_W2ztJ7SQ4_0(.din(n3190), .dout(n3187));
    jdff dff_A_hvYfNHjT3_0(.din(n3193), .dout(n3190));
    jdff dff_A_5V4Ph5x29_0(.din(n3196), .dout(n3193));
    jdff dff_A_hH17uga58_0(.din(n3199), .dout(n3196));
    jdff dff_A_NwXol6hV0_0(.din(n3202), .dout(n3199));
    jdff dff_A_M5IvXN4M6_0(.din(n3205), .dout(n3202));
    jdff dff_A_DiOHebvu5_0(.din(n3208), .dout(n3205));
    jdff dff_A_nHufrf4W8_0(.din(n3211), .dout(n3208));
    jdff dff_A_tkN9220D2_0(.din(G101), .dout(n3211));
    jdff dff_A_5yz7tMgP9_2(.din(n3217), .dout(n3214));
    jdff dff_A_of9VE2Fz6_2(.din(G101), .dout(n3217));
    jdff dff_A_ok4oxW2C4_1(.din(n158), .dout(n3220));
    jdff dff_A_jm8LVCm13_1(.din(n147), .dout(n3223));
    jdff dff_A_wdagkMWX9_2(.din(n147), .dout(n3226));
    jdff dff_A_HL6lsrHG2_2(.din(n3232), .dout(n3229));
    jdff dff_A_jovm5fYq5_2(.din(n3235), .dout(n3232));
    jdff dff_A_Ty6DqOdE5_2(.din(n3238), .dout(n3235));
    jdff dff_A_ux5drhZs3_2(.din(n3241), .dout(n3238));
    jdff dff_A_7PyvplTS7_2(.din(n3244), .dout(n3241));
    jdff dff_A_6gxqJhLc9_2(.din(G472), .dout(n3244));
    jdff dff_B_4qFwiVGm8_0(.din(n123), .dout(n3248));
    jdff dff_A_atZXIHD73_0(.din(n3253), .dout(n3250));
    jdff dff_A_qpoPMpyG5_0(.din(n120), .dout(n3253));
    jdff dff_A_I9CkvksI5_0(.din(n3259), .dout(n3256));
    jdff dff_A_QHyjIXl35_0(.din(n3262), .dout(n3259));
    jdff dff_A_3YG4nnEL4_0(.din(n3265), .dout(n3262));
    jdff dff_A_ene5vLYs2_0(.din(n3268), .dout(n3265));
    jdff dff_A_GzlSrgQs0_0(.din(n3271), .dout(n3268));
    jdff dff_A_jnLxujRO1_0(.din(n3274), .dout(n3271));
    jdff dff_A_0LJTcGe11_0(.din(n3277), .dout(n3274));
    jdff dff_A_MqlHttQF1_0(.din(n3280), .dout(n3277));
    jdff dff_A_n7J2kp7O1_0(.din(n3283), .dout(n3280));
    jdff dff_A_KailyL7u5_0(.din(n3286), .dout(n3283));
    jdff dff_A_QRFDXzvI1_0(.din(n3289), .dout(n3286));
    jdff dff_A_iDaGQMjD6_0(.din(n3292), .dout(n3289));
    jdff dff_A_12fiUFWN7_0(.din(n105), .dout(n3292));
    jdff dff_B_r8oAmEr11_0(.din(n101), .dout(n3296));
    jdff dff_B_LJSWXHrT7_0(.din(n97), .dout(n3299));
    jdff dff_A_Yx99ZoGm0_0(.din(n3304), .dout(n3301));
    jdff dff_A_1E1OJPCW5_0(.din(n3307), .dout(n3304));
    jdff dff_A_j7AwUOtD4_0(.din(n3310), .dout(n3307));
    jdff dff_A_6A9Lev4r5_0(.din(n3313), .dout(n3310));
    jdff dff_A_v3PehkQg4_0(.din(n3316), .dout(n3313));
    jdff dff_A_Y5XU4Hfp1_0(.din(n3319), .dout(n3316));
    jdff dff_A_LTvMCBkk0_0(.din(n3322), .dout(n3319));
    jdff dff_A_IfLVXqSD8_0(.din(n3325), .dout(n3322));
    jdff dff_A_qJTHVnl13_0(.din(n3328), .dout(n3325));
    jdff dff_A_iF4bgQ0X4_0(.din(n3331), .dout(n3328));
    jdff dff_A_NV5cEZc60_0(.din(G137), .dout(n3331));
    jdff dff_B_XiehfK7Z2_0(.din(n81), .dout(n3335));
    jdff dff_A_pYCeHdjc8_0(.din(n3340), .dout(n3337));
    jdff dff_A_iU8Vv90l2_0(.din(n3343), .dout(n3340));
    jdff dff_A_DDLbsdKx4_0(.din(n3346), .dout(n3343));
    jdff dff_A_MIOm2Y5d6_0(.din(n3349), .dout(n3346));
    jdff dff_A_QOpjK0sa1_0(.din(n3352), .dout(n3349));
    jdff dff_A_SNhItwJm2_0(.din(n3355), .dout(n3352));
    jdff dff_A_m6rWxWNt5_0(.din(n3358), .dout(n3355));
    jdff dff_A_kG3Sw8WA6_0(.din(n3361), .dout(n3358));
    jdff dff_A_tUnhX7UW6_0(.din(n3364), .dout(n3361));
    jdff dff_A_SFbsM8nx7_0(.din(n3367), .dout(n3364));
    jdff dff_A_zQr574PS7_0(.din(G119), .dout(n3367));
    jdff dff_A_pnVt8Qtv5_2(.din(G119), .dout(n3370));
    jdff dff_A_d8mwiH3Y7_0(.din(n3376), .dout(n3373));
    jdff dff_A_NVAp0T9d8_0(.din(n3379), .dout(n3376));
    jdff dff_A_KvebgTYX9_0(.din(n3382), .dout(n3379));
    jdff dff_A_lkrQ8U7C8_0(.din(n3385), .dout(n3382));
    jdff dff_A_zWtAHudD5_0(.din(n3388), .dout(n3385));
    jdff dff_A_kl2sIsMx1_0(.din(n3391), .dout(n3388));
    jdff dff_A_p0tcYRmA8_0(.din(n3394), .dout(n3391));
    jdff dff_A_frApIrAX3_0(.din(n3397), .dout(n3394));
    jdff dff_A_YPTbDuYP4_0(.din(n3400), .dout(n3397));
    jdff dff_A_zwFgS79g3_0(.din(n3403), .dout(n3400));
    jdff dff_A_VJyD25BW2_0(.din(G110), .dout(n3403));
    jdff dff_B_LDZoSPUp5_1(.din(n63), .dout(n3407));
    jdff dff_A_rh5X5q869_0(.din(G234), .dout(n3409));
    jdff dff_A_uC1SOD1I5_0(.din(n3415), .dout(n3412));
    jdff dff_A_8kbSZhd42_0(.din(n3418), .dout(n3415));
    jdff dff_A_UmkrL2Bk1_0(.din(G221), .dout(n3418));
    jdff dff_A_XPV2EKVR7_0(.din(n3424), .dout(n3421));
    jdff dff_A_5HXS80rJ5_0(.din(n3427), .dout(n3424));
    jdff dff_A_9srne13f0_0(.din(n3430), .dout(n3427));
    jdff dff_A_IfPdIVTn7_0(.din(n60), .dout(n3430));
    jdff dff_A_oFeZ3aKP2_2(.din(n3436), .dout(n3433));
    jdff dff_A_51Ifwn6Q6_2(.din(n3439), .dout(n3436));
    jdff dff_A_sdkKZKsZ1_2(.din(n3442), .dout(n3439));
    jdff dff_A_H9Rx8CDR8_2(.din(n60), .dout(n3442));
    jdff dff_A_ksj7tYHN6_0(.din(n3448), .dout(n3445));
    jdff dff_A_Itc80Ea72_0(.din(n3451), .dout(n3448));
    jdff dff_A_M39xwuIo0_0(.din(n339), .dout(n3451));
    jdff dff_A_vjxMacjW1_2(.din(n3457), .dout(n3454));
    jdff dff_A_6kFU2oJx0_2(.din(n3460), .dout(n3457));
    jdff dff_A_I3fxLiWP0_2(.din(n3463), .dout(n3460));
    jdff dff_A_UuNkoUaZ8_2(.din(n3466), .dout(n3463));
    jdff dff_A_kdAG6Xfd1_2(.din(n339), .dout(n3466));
    jdff dff_A_eGqH9LWf9_1(.din(n3472), .dout(n3469));
    jdff dff_A_JxLCtbbS1_1(.din(n3475), .dout(n3472));
    jdff dff_A_lQnAgIGT8_1(.din(n3478), .dout(n3475));
    jdff dff_A_IHjKN1eP7_1(.din(n335), .dout(n3478));
    jdff dff_A_TULZPGgB3_2(.din(n3484), .dout(n3481));
    jdff dff_A_PXokvH883_2(.din(n3487), .dout(n3484));
    jdff dff_A_6O1qeEnr7_2(.din(n3490), .dout(n3487));
    jdff dff_A_ranaXLiv7_2(.din(n3493), .dout(n3490));
    jdff dff_A_B7FQSY6u3_2(.din(n3496), .dout(n3493));
    jdff dff_A_lCVW8TrR0_2(.din(n3499), .dout(n3496));
    jdff dff_A_5UsLVNNZ0_2(.din(n3502), .dout(n3499));
    jdff dff_A_mf0Nb3ry8_2(.din(n3505), .dout(n3502));
    jdff dff_A_oEm0Nfpx8_2(.din(n335), .dout(n3505));
    jdff dff_A_raUcn9Zs3_0(.din(n312), .dout(n3508));
    jdff dff_A_HRi1yhR67_1(.din(G898), .dout(n3511));
    jdff dff_A_SipQVlaa6_0(.din(n3517), .dout(n3514));
    jdff dff_A_lZsDVJ0U6_0(.din(n3520), .dout(n3517));
    jdff dff_A_zbzxFhuo2_0(.din(n553), .dout(n3520));
    jdff dff_A_uI0Twndm0_1(.din(n3526), .dout(n3523));
    jdff dff_A_ZMcwRGWY9_1(.din(n3529), .dout(n3526));
    jdff dff_A_0Q9UZn8v8_1(.din(n3532), .dout(n3529));
    jdff dff_A_tod14Z6Y6_1(.din(n3535), .dout(n3532));
    jdff dff_A_n8swF2ru4_1(.din(n3538), .dout(n3535));
    jdff dff_A_zUrRyy1A7_1(.din(n3541), .dout(n3538));
    jdff dff_A_EAxCJBL25_1(.din(n3544), .dout(n3541));
    jdff dff_A_QKGNkm4x4_1(.din(n3547), .dout(n3544));
    jdff dff_A_ZwthStk77_1(.din(n3550), .dout(n3547));
    jdff dff_A_w9kyeGvU5_1(.din(n3553), .dout(n3550));
    jdff dff_A_pqYUnlPZ3_1(.din(n3556), .dout(n3553));
    jdff dff_A_oAl19vRy1_1(.din(n415), .dout(n3556));
    jdff dff_B_MznmxNAg2_1(.din(n389), .dout(n3560));
    jdff dff_B_Ny6Ilyp92_1(.din(n3560), .dout(n3563));
    jdff dff_A_IU5JvZM81_0(.din(n3568), .dout(n3565));
    jdff dff_A_fUlEsfb87_0(.din(n3571), .dout(n3568));
    jdff dff_A_QoXljbPT5_0(.din(n3574), .dout(n3571));
    jdff dff_A_DZezbzRa5_0(.din(n3577), .dout(n3574));
    jdff dff_A_wGEc2Yr71_0(.din(n3580), .dout(n3577));
    jdff dff_A_QOh7BTgc6_0(.din(n3583), .dout(n3580));
    jdff dff_A_ooAehbF87_0(.din(n3586), .dout(n3583));
    jdff dff_A_D6q22Tbe9_0(.din(n3589), .dout(n3586));
    jdff dff_A_I8DYA9Qv1_0(.din(n3592), .dout(n3589));
    jdff dff_A_evfcDjfb0_0(.din(n3595), .dout(n3592));
    jdff dff_A_ttSlfJ5X7_0(.din(G131), .dout(n3595));
    jdff dff_A_CzsLeHrX3_2(.din(G131), .dout(n3598));
    jdff dff_A_4wyfpWne7_1(.din(G953), .dout(n3601));
    jdff dff_A_1s77Wb1L3_1(.din(G214), .dout(n3604));
    jdff dff_A_Hri4DIpK9_0(.din(n93), .dout(n3607));
    jdff dff_A_i447xYnj1_0(.din(n3613), .dout(n3610));
    jdff dff_A_keIiaf2X8_0(.din(n89), .dout(n3613));
    jdff dff_A_rdWeC6J85_0(.din(n3619), .dout(n3616));
    jdff dff_A_BDE4x2dQ5_0(.din(n3622), .dout(n3619));
    jdff dff_A_h0zXj6WS3_0(.din(n3625), .dout(n3622));
    jdff dff_A_voyEWAbT6_0(.din(n3628), .dout(n3625));
    jdff dff_A_THTWZ5bi7_0(.din(n3631), .dout(n3628));
    jdff dff_A_To3tX07H9_0(.din(n3634), .dout(n3631));
    jdff dff_A_e4q1WrRp3_0(.din(n3637), .dout(n3634));
    jdff dff_A_LpAuHaD96_0(.din(n3640), .dout(n3637));
    jdff dff_A_FVrwDWEu1_0(.din(n3643), .dout(n3640));
    jdff dff_A_tg2iyD9N2_0(.din(n3646), .dout(n3643));
    jdff dff_A_muDEwOhg9_0(.din(G140), .dout(n3646));
    jdff dff_A_ZPd97mhW6_1(.din(G140), .dout(n3649));
    jdff dff_A_cXjJ8Opy8_0(.din(n3655), .dout(n3652));
    jdff dff_A_7ke4v4vb5_0(.din(n3658), .dout(n3655));
    jdff dff_A_rD8LgLhk2_0(.din(n3661), .dout(n3658));
    jdff dff_A_z2yKjB7S3_0(.din(n3664), .dout(n3661));
    jdff dff_A_bx9JhTvo5_0(.din(n3667), .dout(n3664));
    jdff dff_A_tMyZlCyb5_0(.din(n3670), .dout(n3667));
    jdff dff_A_szBWCZSm2_0(.din(n3673), .dout(n3670));
    jdff dff_A_2S0qgKkv2_0(.din(n3676), .dout(n3673));
    jdff dff_A_zZLvdgRX9_0(.din(n3679), .dout(n3676));
    jdff dff_A_LcBNfvQP6_0(.din(n3682), .dout(n3679));
    jdff dff_A_tFgBrtCK8_0(.din(G125), .dout(n3682));
    jdff dff_A_0z7d7R0o8_1(.din(n3688), .dout(n3685));
    jdff dff_A_5e6SVyaf6_1(.din(G125), .dout(n3688));
    jdff dff_A_oSJkky0K2_0(.din(n3694), .dout(n3691));
    jdff dff_A_MigrqXIy2_0(.din(n3697), .dout(n3694));
    jdff dff_A_51TVHLii9_0(.din(n3700), .dout(n3697));
    jdff dff_A_qTNc97ON5_0(.din(n3703), .dout(n3700));
    jdff dff_A_TSwgDWBk9_0(.din(n3706), .dout(n3703));
    jdff dff_A_UmJmSd2S3_0(.din(n3709), .dout(n3706));
    jdff dff_A_ZFmGawyg9_0(.din(n3712), .dout(n3709));
    jdff dff_A_5VP60dUO9_0(.din(n3715), .dout(n3712));
    jdff dff_A_sNAq7mdA3_0(.din(n3718), .dout(n3715));
    jdff dff_A_DX3jurAJ6_0(.din(n3722), .dout(n3718));
    jdff dff_B_QYOxYyQh7_3(.din(G146), .dout(n3722));
    jdff dff_A_q10kKYis6_0(.din(n3727), .dout(n3724));
    jdff dff_A_xIbWc7Ky0_0(.din(n3730), .dout(n3727));
    jdff dff_A_gWk1F5el2_0(.din(n3733), .dout(n3730));
    jdff dff_A_mk8zZIpv4_0(.din(n3736), .dout(n3733));
    jdff dff_A_bpPjve709_0(.din(n3739), .dout(n3736));
    jdff dff_A_HFEBdRvo1_0(.din(n3742), .dout(n3739));
    jdff dff_A_T3f7AEBb4_0(.din(n3745), .dout(n3742));
    jdff dff_A_x38dOZzJ8_0(.din(n3748), .dout(n3745));
    jdff dff_A_QAexxTV21_0(.din(n3751), .dout(n3748));
    jdff dff_A_AYKDvV884_0(.din(n3754), .dout(n3751));
    jdff dff_A_NWJHmVeC7_0(.din(G113), .dout(n3754));
    jdff dff_A_O6x76RM51_0(.din(n3760), .dout(n3757));
    jdff dff_A_b90dULUd8_0(.din(n3763), .dout(n3760));
    jdff dff_A_w4W009VD0_0(.din(n3766), .dout(n3763));
    jdff dff_A_UzgZewKc1_0(.din(n3769), .dout(n3766));
    jdff dff_A_BTydVxyW5_0(.din(n3772), .dout(n3769));
    jdff dff_A_8JAonBZg2_0(.din(n3775), .dout(n3772));
    jdff dff_A_ttCS3nBG4_0(.din(n3778), .dout(n3775));
    jdff dff_A_1mz5hszx0_0(.din(n3781), .dout(n3778));
    jdff dff_A_2FjiCEY75_0(.din(n3784), .dout(n3781));
    jdff dff_A_f6iP0Ym57_0(.din(n3787), .dout(n3784));
    jdff dff_A_FBAHzrOq1_0(.din(G104), .dout(n3787));
    jdff dff_A_eUbbvWIE2_1(.din(G104), .dout(n3790));
    jdff dff_A_gxkjBzf02_1(.din(n3796), .dout(n3793));
    jdff dff_A_ZliZVfE29_1(.din(n3799), .dout(n3796));
    jdff dff_A_RMrCSklw6_1(.din(n3802), .dout(n3799));
    jdff dff_A_RjTJWRhP6_1(.din(n3805), .dout(n3802));
    jdff dff_A_wrzlxhLN1_1(.din(n3808), .dout(n3805));
    jdff dff_A_kUu1Mzls8_1(.din(G475), .dout(n3808));
    jdff dff_A_xUoOSNcT2_0(.din(n3814), .dout(n3811));
    jdff dff_A_mcS7BPxg3_0(.din(n3817), .dout(n3814));
    jdff dff_A_YwwUhA365_0(.din(n3820), .dout(n3817));
    jdff dff_A_Qja3vFFE1_0(.din(n3823), .dout(n3820));
    jdff dff_A_hgcMTnVZ5_0(.din(n3826), .dout(n3823));
    jdff dff_A_oF4bRuhQ9_0(.din(n3829), .dout(n3826));
    jdff dff_A_9PowGjIE1_0(.din(n3832), .dout(n3829));
    jdff dff_A_VvIYXqj79_0(.din(n3835), .dout(n3832));
    jdff dff_A_2vxRWCz35_0(.din(n3838), .dout(n3835));
    jdff dff_A_1xla2iDB4_0(.din(n3841), .dout(n3838));
    jdff dff_A_5YYL5PxY7_0(.din(n3844), .dout(n3841));
    jdff dff_A_6MTAriep6_0(.din(n3847), .dout(n3844));
    jdff dff_A_POImPkBN8_0(.din(n370), .dout(n3847));
    jdff dff_B_rSeBfPmu5_1(.din(n346), .dout(n3851));
    jdff dff_B_CN858ycW5_1(.din(n3851), .dout(n3854));
    jdff dff_B_bm62cSlV3_0(.din(n362), .dout(n3857));
    jdff dff_A_IJjrdxt81_1(.din(n3862), .dout(n3859));
    jdff dff_A_Y3wHbrTA3_1(.din(n3865), .dout(n3862));
    jdff dff_A_MQYJhE4y9_1(.din(n3868), .dout(n3865));
    jdff dff_A_EQX7NdHE4_1(.din(n3871), .dout(n3868));
    jdff dff_A_VBLw9gIW4_1(.din(n3874), .dout(n3871));
    jdff dff_A_uHo0OgwD3_1(.din(n3877), .dout(n3874));
    jdff dff_A_8E6CQeG16_1(.din(n3880), .dout(n3877));
    jdff dff_A_6Z6ifrbO5_1(.din(n3883), .dout(n3880));
    jdff dff_A_dSleeQiT2_1(.din(n3886), .dout(n3883));
    jdff dff_A_MFjApbeP1_1(.din(n3889), .dout(n3886));
    jdff dff_A_i3wbb3jA9_1(.din(n3892), .dout(n3889));
    jdff dff_A_68C1tYLB7_1(.din(G122), .dout(n3892));
    jdff dff_A_nga2Iew62_0(.din(n3898), .dout(n3895));
    jdff dff_A_Prbkge5E7_0(.din(n3901), .dout(n3898));
    jdff dff_A_nyqnGPiK0_0(.din(n3904), .dout(n3901));
    jdff dff_A_g30tdJAs5_0(.din(n3907), .dout(n3904));
    jdff dff_A_57r37bCg9_0(.din(n3910), .dout(n3907));
    jdff dff_A_RnaV8Cpi8_0(.din(n3913), .dout(n3910));
    jdff dff_A_3wMrxpah6_0(.din(n3916), .dout(n3913));
    jdff dff_A_TiER8Ba95_0(.din(n3919), .dout(n3916));
    jdff dff_A_0bVYrvQ19_0(.din(n3922), .dout(n3919));
    jdff dff_A_N5DlPHLb0_0(.din(n3925), .dout(n3922));
    jdff dff_A_NLyaARlw7_0(.din(G116), .dout(n3925));
    jdff dff_A_49YsQQxQ0_0(.din(n3931), .dout(n3928));
    jdff dff_A_8p83rKFq1_0(.din(n3934), .dout(n3931));
    jdff dff_A_iUkqLGaB4_0(.din(n3937), .dout(n3934));
    jdff dff_A_yRgsuM321_0(.din(n3940), .dout(n3937));
    jdff dff_A_vVB9dRLj0_0(.din(n3943), .dout(n3940));
    jdff dff_A_2zdQqUdi1_0(.din(n3946), .dout(n3943));
    jdff dff_A_qtxv1z6j6_0(.din(n3949), .dout(n3946));
    jdff dff_A_9oU8Yl8g4_0(.din(n3952), .dout(n3949));
    jdff dff_A_rh4Mc7Np3_0(.din(n3955), .dout(n3952));
    jdff dff_A_yuS9hSMZ4_0(.din(n3958), .dout(n3955));
    jdff dff_A_CesXBU2u2_0(.din(G107), .dout(n3958));
    jdff dff_A_6FeGUKFN4_1(.din(G107), .dout(n3961));
    jdff dff_A_bly7LfRR9_2(.din(n3967), .dout(n3964));
    jdff dff_A_kfr5z0gz9_2(.din(n230), .dout(n3967));
    jdff dff_A_XAwPxIpV3_1(.din(G234), .dout(n3970));
    jdff dff_A_AaRWqBMq8_0(.din(n3976), .dout(n3973));
    jdff dff_A_9P4CbAt02_0(.din(n3979), .dout(n3976));
    jdff dff_A_dcESeOtO4_0(.din(n3982), .dout(n3979));
    jdff dff_A_pDr1Ffty0_0(.din(n3985), .dout(n3982));
    jdff dff_A_1XeUmfh58_0(.din(n3988), .dout(n3985));
    jdff dff_A_UN32hoSG4_0(.din(n3991), .dout(n3988));
    jdff dff_A_hSTybxa97_0(.din(n3994), .dout(n3991));
    jdff dff_A_gY1PkqQ66_0(.din(n3997), .dout(n3994));
    jdff dff_A_zKFyXN3O9_0(.din(n4000), .dout(n3997));
    jdff dff_A_P0HFjRp93_0(.din(n4003), .dout(n4000));
    jdff dff_A_oTlpMXOD9_0(.din(n4006), .dout(n4003));
    jdff dff_A_AjRwY4x19_0(.din(n4009), .dout(n4006));
    jdff dff_A_sI67HIFr7_0(.din(n4012), .dout(n4009));
    jdff dff_A_mYZjQoQo4_0(.din(n4022), .dout(n4012));
    jdff dff_A_JcBqaPAX3_2(.din(n4022), .dout(n4015));
    jdff dff_B_oh5QZlDJ4_3(.din(G217), .dout(n4019));
    jdff dff_B_M3j6QPic7_3(.din(n4019), .dout(n4022));
    jdff dff_A_DcTb4TUm5_0(.din(n4027), .dout(n4024));
    jdff dff_A_fSoIHhZ60_0(.din(n4030), .dout(n4027));
    jdff dff_A_UFQDDTAz1_0(.din(n4033), .dout(n4030));
    jdff dff_A_tqndewNR1_0(.din(n4036), .dout(n4033));
    jdff dff_A_msk2iWml3_0(.din(n4039), .dout(n4036));
    jdff dff_A_g6NQHAoh9_0(.din(n4042), .dout(n4039));
    jdff dff_A_Q03tJHuo7_0(.din(n4045), .dout(n4042));
    jdff dff_A_zS251Rh04_0(.din(n4048), .dout(n4045));
    jdff dff_A_eAuW7okS4_0(.din(n4051), .dout(n4048));
    jdff dff_A_PAAYFXB99_0(.din(n4054), .dout(n4051));
    jdff dff_A_ryEwEkan5_0(.din(G143), .dout(n4054));
    jdff dff_A_dmHWo8dH3_1(.din(G143), .dout(n4057));
    jdff dff_A_1Zt6HHmR4_0(.din(n4063), .dout(n4060));
    jdff dff_A_2OvaMXge7_0(.din(n4066), .dout(n4063));
    jdff dff_A_hHsEpiOP6_0(.din(n4069), .dout(n4066));
    jdff dff_A_naPrRy4H7_0(.din(n4072), .dout(n4069));
    jdff dff_A_6RwbPwZM9_0(.din(n4075), .dout(n4072));
    jdff dff_A_fnWTvjgw0_0(.din(n4078), .dout(n4075));
    jdff dff_A_oszF1gkS2_0(.din(n4081), .dout(n4078));
    jdff dff_A_lEWY4w7D6_0(.din(n4084), .dout(n4081));
    jdff dff_A_bpc1Pi4f8_0(.din(n4087), .dout(n4084));
    jdff dff_A_4U4Dn5B10_0(.din(n4090), .dout(n4087));
    jdff dff_A_7dghcLrw1_0(.din(G128), .dout(n4090));
    jdff dff_A_4MXdOiW35_0(.din(n4096), .dout(n4093));
    jdff dff_A_699554VJ5_0(.din(n4099), .dout(n4096));
    jdff dff_A_WciAu2Qa8_0(.din(n4102), .dout(n4099));
    jdff dff_A_N7BOy3hJ9_0(.din(n4105), .dout(n4102));
    jdff dff_A_3mtpfrEd9_0(.din(n4108), .dout(n4105));
    jdff dff_A_INH41D6U6_0(.din(n4111), .dout(n4108));
    jdff dff_A_PzPKDana9_0(.din(n4114), .dout(n4111));
    jdff dff_A_ZO63gEjH1_0(.din(n4117), .dout(n4114));
    jdff dff_A_rnKEsWx37_0(.din(n4120), .dout(n4117));
    jdff dff_A_NDNan9j49_0(.din(n4123), .dout(n4120));
    jdff dff_A_7gLeVlQI2_0(.din(G134), .dout(n4123));
    jdff dff_A_XcRayItl7_1(.din(G134), .dout(n4126));
    jdff dff_A_i9Og0RTD8_0(.din(n4132), .dout(n4129));
    jdff dff_A_yEqPEles3_0(.din(n4135), .dout(n4132));
    jdff dff_A_cVYZLGLT9_0(.din(n4138), .dout(n4135));
    jdff dff_A_lPlN46Zi2_0(.din(n60), .dout(n4138));
    jdff dff_A_rA1iVUIV8_2(.din(n4144), .dout(n4141));
    jdff dff_A_lqjD7w6a1_2(.din(n4147), .dout(n4144));
    jdff dff_A_6vZRGKSU4_2(.din(n4150), .dout(n4147));
    jdff dff_A_z0LuLn477_2(.din(n60), .dout(n4150));
    jdff dff_A_1yJTqHgw8_0(.din(n4156), .dout(n4153));
    jdff dff_A_ekZdutAZ2_0(.din(G902), .dout(n4156));
    jdff dff_A_v6I2KH7f2_0(.din(n4162), .dout(n4159));
    jdff dff_A_JzvUZGg29_0(.din(n4165), .dout(n4162));
    jdff dff_A_azIfX3Y38_0(.din(n4168), .dout(n4165));
    jdff dff_A_DmcJJByz4_0(.din(n4171), .dout(n4168));
    jdff dff_A_DQ4NMHGq0_0(.din(n4174), .dout(n4171));
    jdff dff_A_g7pf2V5u6_0(.din(n4177), .dout(n4174));
    jdff dff_A_po0E5KME4_0(.din(n4180), .dout(n4177));
    jdff dff_A_sSABVEBM1_0(.din(n4183), .dout(n4180));
    jdff dff_A_wSa2KBbh5_0(.din(n4186), .dout(n4183));
    jdff dff_A_UwQepUMf0_0(.din(n4189), .dout(n4186));
    jdff dff_A_zjJnu9ml6_0(.din(n4192), .dout(n4189));
    jdff dff_A_53XppaRC8_0(.din(n4195), .dout(n4192));
    jdff dff_A_N1vGFIui8_0(.din(n4198), .dout(n4195));
    jdff dff_A_A3mIpxqX5_0(.din(n4201), .dout(n4198));
    jdff dff_A_Pb6hprQj1_0(.din(n4204), .dout(n4201));
    jdff dff_A_H4EUOxXu5_0(.din(G478), .dout(n4204));
    jdff dff_A_z11SiYkI1_1(.din(n4210), .dout(n4207));
    jdff dff_A_u17sdarp3_1(.din(n4213), .dout(n4210));
    jdff dff_A_uejkKqTt8_1(.din(n4216), .dout(n4213));
    jdff dff_A_ErbHBAEZ7_1(.din(n4219), .dout(n4216));
    jdff dff_A_EBDUmzyk5_1(.din(n4222), .dout(n4219));
    jdff dff_A_bF80AltB1_1(.din(G478), .dout(n4222));
    jdff dff_A_apHLc5GV3_1(.din(n4274), .dout(n4225));
    jdff dff_B_FkmzQT5x0_3(.din(n867), .dout(n4229));
    jdff dff_B_sdL8uqzI8_3(.din(n4229), .dout(n4232));
    jdff dff_B_glo3kX217_3(.din(n4232), .dout(n4235));
    jdff dff_B_jqo5RMfB2_3(.din(n4235), .dout(n4238));
    jdff dff_B_3i79ASGC1_3(.din(n4238), .dout(n4241));
    jdff dff_B_orduQgoF1_3(.din(n4241), .dout(n4244));
    jdff dff_B_mKTavY603_3(.din(n4244), .dout(n4247));
    jdff dff_B_YiyA7Xno4_3(.din(n4247), .dout(n4250));
    jdff dff_B_JwMiTnx43_3(.din(n4250), .dout(n4253));
    jdff dff_B_5oOo1v0z3_3(.din(n4253), .dout(n4256));
    jdff dff_B_JDfv641l3_3(.din(n4256), .dout(n4259));
    jdff dff_B_ZOBIZjc95_3(.din(n4259), .dout(n4262));
    jdff dff_B_aM2RjltO6_3(.din(n4262), .dout(n4265));
    jdff dff_B_QKUuJj6k5_3(.din(n4265), .dout(n4268));
    jdff dff_B_PhKd6gim7_3(.din(n4268), .dout(n4271));
    jdff dff_B_ABthXCsD1_3(.din(n4271), .dout(n4274));
    jdff dff_A_zpocZClW1_0(.din(n4279), .dout(n4276));
    jdff dff_A_kzb2hd9g2_0(.din(n4282), .dout(n4279));
endmodule

