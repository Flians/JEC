/*

c6288:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jdff: 8046
	jand: 664
	jor: 312

Summary:
	jxor: 462
	jspl: 936
	jspl3: 251
	jnot: 321
	jdff: 8046
	jand: 664
	jor: 312
*/

module c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G1gat_1;
	wire[2:0] w_G1gat_2;
	wire[2:0] w_G1gat_3;
	wire[2:0] w_G1gat_4;
	wire[2:0] w_G1gat_5;
	wire[2:0] w_G1gat_6;
	wire[1:0] w_G1gat_7;
	wire[2:0] w_G18gat_0;
	wire[2:0] w_G18gat_1;
	wire[2:0] w_G18gat_2;
	wire[2:0] w_G18gat_3;
	wire[2:0] w_G18gat_4;
	wire[2:0] w_G18gat_5;
	wire[2:0] w_G18gat_6;
	wire[1:0] w_G18gat_7;
	wire[2:0] w_G35gat_0;
	wire[2:0] w_G35gat_1;
	wire[2:0] w_G35gat_2;
	wire[2:0] w_G35gat_3;
	wire[2:0] w_G35gat_4;
	wire[2:0] w_G35gat_5;
	wire[2:0] w_G35gat_6;
	wire[2:0] w_G35gat_7;
	wire[2:0] w_G52gat_0;
	wire[2:0] w_G52gat_1;
	wire[2:0] w_G52gat_2;
	wire[2:0] w_G52gat_3;
	wire[2:0] w_G52gat_4;
	wire[2:0] w_G52gat_5;
	wire[2:0] w_G52gat_6;
	wire[2:0] w_G52gat_7;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G69gat_1;
	wire[2:0] w_G69gat_2;
	wire[2:0] w_G69gat_3;
	wire[2:0] w_G69gat_4;
	wire[2:0] w_G69gat_5;
	wire[2:0] w_G69gat_6;
	wire[1:0] w_G69gat_7;
	wire[2:0] w_G86gat_0;
	wire[2:0] w_G86gat_1;
	wire[2:0] w_G86gat_2;
	wire[2:0] w_G86gat_3;
	wire[2:0] w_G86gat_4;
	wire[2:0] w_G86gat_5;
	wire[2:0] w_G86gat_6;
	wire[1:0] w_G86gat_7;
	wire[2:0] w_G103gat_0;
	wire[2:0] w_G103gat_1;
	wire[2:0] w_G103gat_2;
	wire[2:0] w_G103gat_3;
	wire[2:0] w_G103gat_4;
	wire[2:0] w_G103gat_5;
	wire[2:0] w_G103gat_6;
	wire[1:0] w_G103gat_7;
	wire[2:0] w_G120gat_0;
	wire[2:0] w_G120gat_1;
	wire[2:0] w_G120gat_2;
	wire[2:0] w_G120gat_3;
	wire[2:0] w_G120gat_4;
	wire[2:0] w_G120gat_5;
	wire[2:0] w_G120gat_6;
	wire[1:0] w_G120gat_7;
	wire[2:0] w_G137gat_0;
	wire[2:0] w_G137gat_1;
	wire[2:0] w_G137gat_2;
	wire[2:0] w_G137gat_3;
	wire[2:0] w_G137gat_4;
	wire[2:0] w_G137gat_5;
	wire[2:0] w_G137gat_6;
	wire[1:0] w_G137gat_7;
	wire[2:0] w_G154gat_0;
	wire[2:0] w_G154gat_1;
	wire[2:0] w_G154gat_2;
	wire[2:0] w_G154gat_3;
	wire[2:0] w_G154gat_4;
	wire[2:0] w_G154gat_5;
	wire[2:0] w_G154gat_6;
	wire[1:0] w_G154gat_7;
	wire[2:0] w_G171gat_0;
	wire[2:0] w_G171gat_1;
	wire[2:0] w_G171gat_2;
	wire[2:0] w_G171gat_3;
	wire[2:0] w_G171gat_4;
	wire[2:0] w_G171gat_5;
	wire[2:0] w_G171gat_6;
	wire[1:0] w_G171gat_7;
	wire[2:0] w_G188gat_0;
	wire[2:0] w_G188gat_1;
	wire[2:0] w_G188gat_2;
	wire[2:0] w_G188gat_3;
	wire[2:0] w_G188gat_4;
	wire[2:0] w_G188gat_5;
	wire[2:0] w_G188gat_6;
	wire[1:0] w_G188gat_7;
	wire[2:0] w_G205gat_0;
	wire[2:0] w_G205gat_1;
	wire[2:0] w_G205gat_2;
	wire[2:0] w_G205gat_3;
	wire[2:0] w_G205gat_4;
	wire[2:0] w_G205gat_5;
	wire[2:0] w_G205gat_6;
	wire[1:0] w_G205gat_7;
	wire[2:0] w_G222gat_0;
	wire[2:0] w_G222gat_1;
	wire[2:0] w_G222gat_2;
	wire[2:0] w_G222gat_3;
	wire[2:0] w_G222gat_4;
	wire[2:0] w_G222gat_5;
	wire[2:0] w_G222gat_6;
	wire[1:0] w_G222gat_7;
	wire[2:0] w_G239gat_0;
	wire[2:0] w_G239gat_1;
	wire[2:0] w_G239gat_2;
	wire[2:0] w_G239gat_3;
	wire[2:0] w_G239gat_4;
	wire[2:0] w_G239gat_5;
	wire[2:0] w_G239gat_6;
	wire[1:0] w_G239gat_7;
	wire[2:0] w_G256gat_0;
	wire[2:0] w_G256gat_1;
	wire[2:0] w_G256gat_2;
	wire[2:0] w_G256gat_3;
	wire[2:0] w_G256gat_4;
	wire[2:0] w_G256gat_5;
	wire[2:0] w_G256gat_6;
	wire[1:0] w_G256gat_7;
	wire[2:0] w_G273gat_0;
	wire[2:0] w_G273gat_1;
	wire[2:0] w_G273gat_2;
	wire[2:0] w_G273gat_3;
	wire[2:0] w_G273gat_4;
	wire[2:0] w_G273gat_5;
	wire[2:0] w_G273gat_6;
	wire[1:0] w_G273gat_7;
	wire[2:0] w_G290gat_0;
	wire[2:0] w_G290gat_1;
	wire[2:0] w_G290gat_2;
	wire[2:0] w_G290gat_3;
	wire[2:0] w_G290gat_4;
	wire[2:0] w_G290gat_5;
	wire[2:0] w_G290gat_6;
	wire[2:0] w_G290gat_7;
	wire[2:0] w_G307gat_0;
	wire[2:0] w_G307gat_1;
	wire[2:0] w_G307gat_2;
	wire[2:0] w_G307gat_3;
	wire[2:0] w_G307gat_4;
	wire[2:0] w_G307gat_5;
	wire[2:0] w_G307gat_6;
	wire[1:0] w_G307gat_7;
	wire[2:0] w_G324gat_0;
	wire[2:0] w_G324gat_1;
	wire[2:0] w_G324gat_2;
	wire[2:0] w_G324gat_3;
	wire[2:0] w_G324gat_4;
	wire[2:0] w_G324gat_5;
	wire[2:0] w_G324gat_6;
	wire[1:0] w_G324gat_7;
	wire[2:0] w_G341gat_0;
	wire[2:0] w_G341gat_1;
	wire[2:0] w_G341gat_2;
	wire[2:0] w_G341gat_3;
	wire[2:0] w_G341gat_4;
	wire[2:0] w_G341gat_5;
	wire[2:0] w_G341gat_6;
	wire[1:0] w_G341gat_7;
	wire[2:0] w_G358gat_0;
	wire[2:0] w_G358gat_1;
	wire[2:0] w_G358gat_2;
	wire[2:0] w_G358gat_3;
	wire[2:0] w_G358gat_4;
	wire[2:0] w_G358gat_5;
	wire[2:0] w_G358gat_6;
	wire[1:0] w_G358gat_7;
	wire[2:0] w_G375gat_0;
	wire[2:0] w_G375gat_1;
	wire[2:0] w_G375gat_2;
	wire[2:0] w_G375gat_3;
	wire[2:0] w_G375gat_4;
	wire[2:0] w_G375gat_5;
	wire[2:0] w_G375gat_6;
	wire[1:0] w_G375gat_7;
	wire[2:0] w_G392gat_0;
	wire[2:0] w_G392gat_1;
	wire[2:0] w_G392gat_2;
	wire[2:0] w_G392gat_3;
	wire[2:0] w_G392gat_4;
	wire[2:0] w_G392gat_5;
	wire[2:0] w_G392gat_6;
	wire[1:0] w_G392gat_7;
	wire[2:0] w_G409gat_0;
	wire[2:0] w_G409gat_1;
	wire[2:0] w_G409gat_2;
	wire[2:0] w_G409gat_3;
	wire[2:0] w_G409gat_4;
	wire[2:0] w_G409gat_5;
	wire[2:0] w_G409gat_6;
	wire[1:0] w_G409gat_7;
	wire[2:0] w_G426gat_0;
	wire[2:0] w_G426gat_1;
	wire[2:0] w_G426gat_2;
	wire[2:0] w_G426gat_3;
	wire[2:0] w_G426gat_4;
	wire[2:0] w_G426gat_5;
	wire[2:0] w_G426gat_6;
	wire[1:0] w_G426gat_7;
	wire[2:0] w_G443gat_0;
	wire[2:0] w_G443gat_1;
	wire[2:0] w_G443gat_2;
	wire[2:0] w_G443gat_3;
	wire[2:0] w_G443gat_4;
	wire[2:0] w_G443gat_5;
	wire[2:0] w_G443gat_6;
	wire[1:0] w_G443gat_7;
	wire[2:0] w_G460gat_0;
	wire[2:0] w_G460gat_1;
	wire[2:0] w_G460gat_2;
	wire[2:0] w_G460gat_3;
	wire[2:0] w_G460gat_4;
	wire[2:0] w_G460gat_5;
	wire[2:0] w_G460gat_6;
	wire[1:0] w_G460gat_7;
	wire[2:0] w_G477gat_0;
	wire[2:0] w_G477gat_1;
	wire[2:0] w_G477gat_2;
	wire[2:0] w_G477gat_3;
	wire[2:0] w_G477gat_4;
	wire[2:0] w_G477gat_5;
	wire[2:0] w_G477gat_6;
	wire[1:0] w_G477gat_7;
	wire[2:0] w_G494gat_0;
	wire[2:0] w_G494gat_1;
	wire[2:0] w_G494gat_2;
	wire[2:0] w_G494gat_3;
	wire[2:0] w_G494gat_4;
	wire[2:0] w_G494gat_5;
	wire[2:0] w_G494gat_6;
	wire[1:0] w_G494gat_7;
	wire[2:0] w_G511gat_0;
	wire[2:0] w_G511gat_1;
	wire[2:0] w_G511gat_2;
	wire[2:0] w_G511gat_3;
	wire[2:0] w_G511gat_4;
	wire[2:0] w_G511gat_5;
	wire[2:0] w_G511gat_6;
	wire[1:0] w_G511gat_7;
	wire[2:0] w_G528gat_0;
	wire[2:0] w_G528gat_1;
	wire[2:0] w_G528gat_2;
	wire[2:0] w_G528gat_3;
	wire[2:0] w_G528gat_4;
	wire[2:0] w_G528gat_5;
	wire[2:0] w_G528gat_6;
	wire[1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire[1:0] w_n65_0;
	wire[1:0] w_n66_0;
	wire[1:0] w_n67_0;
	wire[1:0] w_n69_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n75_0;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[2:0] w_n80_0;
	wire[1:0] w_n83_0;
	wire[1:0] w_n84_0;
	wire[1:0] w_n86_0;
	wire[1:0] w_n90_0;
	wire[1:0] w_n91_0;
	wire[1:0] w_n93_0;
	wire[1:0] w_n97_0;
	wire[1:0] w_n99_0;
	wire[2:0] w_n101_0;
	wire[1:0] w_n103_0;
	wire[1:0] w_n104_0;
	wire[1:0] w_n106_0;
	wire[1:0] w_n111_0;
	wire[1:0] w_n112_0;
	wire[2:0] w_n117_0;
	wire[1:0] w_n119_0;
	wire[1:0] w_n120_0;
	wire[1:0] w_n121_0;
	wire[1:0] w_n122_0;
	wire[1:0] w_n123_0;
	wire[1:0] w_n125_0;
	wire[1:0] w_n127_0;
	wire[1:0] w_n128_0;
	wire[1:0] w_n129_0;
	wire[1:0] w_n130_0;
	wire[1:0] w_n132_0;
	wire[1:0] w_n133_0;
	wire[1:0] w_n135_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n141_0;
	wire[2:0] w_n146_0;
	wire[1:0] w_n148_0;
	wire[1:0] w_n152_0;
	wire[1:0] w_n154_0;
	wire[1:0] w_n155_0;
	wire[1:0] w_n156_0;
	wire[1:0] w_n157_0;
	wire[1:0] w_n158_0;
	wire[1:0] w_n160_0;
	wire[1:0] w_n161_0;
	wire[1:0] w_n162_0;
	wire[1:0] w_n163_0;
	wire[1:0] w_n164_0;
	wire[1:0] w_n165_0;
	wire[1:0] w_n167_0;
	wire[1:0] w_n168_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n175_0;
	wire[1:0] w_n176_0;
	wire[2:0] w_n181_0;
	wire[1:0] w_n183_0;
	wire[1:0] w_n186_0;
	wire[1:0] w_n188_0;
	wire[1:0] w_n192_0;
	wire[1:0] w_n194_0;
	wire[1:0] w_n195_0;
	wire[2:0] w_n196_0;
	wire[1:0] w_n198_0;
	wire[1:0] w_n200_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n202_0;
	wire[1:0] w_n203_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n205_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n207_0;
	wire[1:0] w_n209_0;
	wire[1:0] w_n210_0;
	wire[1:0] w_n212_0;
	wire[1:0] w_n217_0;
	wire[1:0] w_n218_0;
	wire[2:0] w_n223_0;
	wire[1:0] w_n225_0;
	wire[1:0] w_n228_0;
	wire[1:0] w_n230_0;
	wire[1:0] w_n233_0;
	wire[1:0] w_n235_0;
	wire[1:0] w_n239_0;
	wire[1:0] w_n241_0;
	wire[1:0] w_n242_0;
	wire[2:0] w_n243_0;
	wire[1:0] w_n245_0;
	wire[1:0] w_n247_0;
	wire[1:0] w_n248_0;
	wire[1:0] w_n249_0;
	wire[1:0] w_n250_0;
	wire[1:0] w_n251_0;
	wire[1:0] w_n252_0;
	wire[1:0] w_n253_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n255_0;
	wire[1:0] w_n256_0;
	wire[1:0] w_n258_0;
	wire[1:0] w_n259_0;
	wire[1:0] w_n261_0;
	wire[1:0] w_n266_0;
	wire[1:0] w_n267_0;
	wire[2:0] w_n272_0;
	wire[1:0] w_n274_0;
	wire[1:0] w_n277_0;
	wire[1:0] w_n279_0;
	wire[1:0] w_n282_0;
	wire[1:0] w_n284_0;
	wire[1:0] w_n287_0;
	wire[1:0] w_n289_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n295_0;
	wire[1:0] w_n296_0;
	wire[2:0] w_n297_0;
	wire[1:0] w_n299_0;
	wire[1:0] w_n301_0;
	wire[1:0] w_n302_0;
	wire[1:0] w_n303_0;
	wire[1:0] w_n304_0;
	wire[1:0] w_n305_0;
	wire[1:0] w_n306_0;
	wire[1:0] w_n307_0;
	wire[1:0] w_n308_0;
	wire[1:0] w_n309_0;
	wire[1:0] w_n310_0;
	wire[1:0] w_n311_0;
	wire[1:0] w_n312_0;
	wire[1:0] w_n314_0;
	wire[1:0] w_n315_0;
	wire[1:0] w_n317_0;
	wire[1:0] w_n322_0;
	wire[1:0] w_n323_0;
	wire[2:0] w_n328_0;
	wire[1:0] w_n330_0;
	wire[1:0] w_n333_0;
	wire[1:0] w_n335_0;
	wire[1:0] w_n338_0;
	wire[1:0] w_n340_0;
	wire[1:0] w_n343_0;
	wire[1:0] w_n345_0;
	wire[1:0] w_n348_0;
	wire[1:0] w_n350_0;
	wire[1:0] w_n354_0;
	wire[1:0] w_n356_0;
	wire[1:0] w_n357_0;
	wire[2:0] w_n358_0;
	wire[1:0] w_n360_0;
	wire[1:0] w_n362_0;
	wire[1:0] w_n363_0;
	wire[1:0] w_n364_0;
	wire[1:0] w_n365_0;
	wire[1:0] w_n366_0;
	wire[1:0] w_n367_0;
	wire[1:0] w_n368_0;
	wire[1:0] w_n369_0;
	wire[1:0] w_n370_0;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n373_0;
	wire[1:0] w_n374_0;
	wire[1:0] w_n375_0;
	wire[1:0] w_n377_0;
	wire[1:0] w_n378_0;
	wire[1:0] w_n380_0;
	wire[1:0] w_n385_0;
	wire[1:0] w_n386_0;
	wire[2:0] w_n391_0;
	wire[1:0] w_n393_0;
	wire[1:0] w_n396_0;
	wire[1:0] w_n398_0;
	wire[1:0] w_n401_0;
	wire[1:0] w_n403_0;
	wire[1:0] w_n406_0;
	wire[1:0] w_n408_0;
	wire[1:0] w_n411_0;
	wire[1:0] w_n413_0;
	wire[1:0] w_n416_0;
	wire[1:0] w_n418_0;
	wire[1:0] w_n423_0;
	wire[1:0] w_n425_0;
	wire[1:0] w_n426_0;
	wire[2:0] w_n427_0;
	wire[1:0] w_n429_0;
	wire[1:0] w_n431_0;
	wire[1:0] w_n432_0;
	wire[1:0] w_n433_0;
	wire[1:0] w_n434_0;
	wire[1:0] w_n435_0;
	wire[1:0] w_n436_0;
	wire[1:0] w_n437_0;
	wire[1:0] w_n438_0;
	wire[1:0] w_n439_0;
	wire[1:0] w_n440_0;
	wire[1:0] w_n441_0;
	wire[1:0] w_n442_0;
	wire[1:0] w_n443_0;
	wire[1:0] w_n444_0;
	wire[1:0] w_n445_0;
	wire[1:0] w_n446_0;
	wire[1:0] w_n448_0;
	wire[1:0] w_n449_0;
	wire[1:0] w_n451_0;
	wire[1:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[2:0] w_n462_0;
	wire[1:0] w_n464_0;
	wire[1:0] w_n467_0;
	wire[1:0] w_n469_0;
	wire[1:0] w_n472_0;
	wire[1:0] w_n474_0;
	wire[1:0] w_n477_0;
	wire[1:0] w_n479_0;
	wire[1:0] w_n482_0;
	wire[1:0] w_n484_0;
	wire[1:0] w_n487_0;
	wire[1:0] w_n489_0;
	wire[1:0] w_n492_0;
	wire[1:0] w_n494_0;
	wire[1:0] w_n499_0;
	wire[1:0] w_n501_0;
	wire[1:0] w_n502_0;
	wire[2:0] w_n503_0;
	wire[1:0] w_n505_0;
	wire[1:0] w_n507_0;
	wire[1:0] w_n508_0;
	wire[1:0] w_n509_0;
	wire[1:0] w_n510_0;
	wire[1:0] w_n511_0;
	wire[1:0] w_n512_0;
	wire[1:0] w_n513_0;
	wire[1:0] w_n514_0;
	wire[1:0] w_n515_0;
	wire[1:0] w_n516_0;
	wire[1:0] w_n517_0;
	wire[1:0] w_n518_0;
	wire[1:0] w_n519_0;
	wire[1:0] w_n520_0;
	wire[1:0] w_n521_0;
	wire[1:0] w_n522_0;
	wire[1:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n526_0;
	wire[1:0] w_n527_0;
	wire[1:0] w_n529_0;
	wire[1:0] w_n534_0;
	wire[1:0] w_n535_0;
	wire[2:0] w_n540_0;
	wire[1:0] w_n542_0;
	wire[1:0] w_n545_0;
	wire[1:0] w_n547_0;
	wire[1:0] w_n550_0;
	wire[1:0] w_n552_0;
	wire[1:0] w_n555_0;
	wire[1:0] w_n557_0;
	wire[1:0] w_n560_0;
	wire[1:0] w_n562_0;
	wire[1:0] w_n565_0;
	wire[1:0] w_n567_0;
	wire[1:0] w_n570_0;
	wire[1:0] w_n572_0;
	wire[1:0] w_n575_0;
	wire[1:0] w_n577_0;
	wire[1:0] w_n582_0;
	wire[1:0] w_n584_0;
	wire[1:0] w_n585_0;
	wire[2:0] w_n586_0;
	wire[1:0] w_n588_0;
	wire[1:0] w_n590_0;
	wire[1:0] w_n591_0;
	wire[1:0] w_n592_0;
	wire[1:0] w_n593_0;
	wire[1:0] w_n594_0;
	wire[1:0] w_n595_0;
	wire[1:0] w_n596_0;
	wire[1:0] w_n597_0;
	wire[1:0] w_n598_0;
	wire[1:0] w_n599_0;
	wire[1:0] w_n600_0;
	wire[1:0] w_n601_0;
	wire[1:0] w_n602_0;
	wire[1:0] w_n603_0;
	wire[1:0] w_n604_0;
	wire[1:0] w_n605_0;
	wire[1:0] w_n606_0;
	wire[1:0] w_n607_0;
	wire[1:0] w_n608_0;
	wire[1:0] w_n609_0;
	wire[1:0] w_n611_0;
	wire[1:0] w_n612_0;
	wire[1:0] w_n614_0;
	wire[1:0] w_n619_0;
	wire[1:0] w_n620_0;
	wire[2:0] w_n625_0;
	wire[1:0] w_n627_0;
	wire[1:0] w_n630_0;
	wire[1:0] w_n632_0;
	wire[1:0] w_n635_0;
	wire[1:0] w_n637_0;
	wire[1:0] w_n640_0;
	wire[1:0] w_n642_0;
	wire[1:0] w_n645_0;
	wire[1:0] w_n647_0;
	wire[1:0] w_n650_0;
	wire[1:0] w_n652_0;
	wire[1:0] w_n655_0;
	wire[1:0] w_n657_0;
	wire[1:0] w_n660_0;
	wire[1:0] w_n662_0;
	wire[1:0] w_n665_0;
	wire[1:0] w_n667_0;
	wire[1:0] w_n672_0;
	wire[1:0] w_n674_0;
	wire[1:0] w_n675_0;
	wire[2:0] w_n676_0;
	wire[1:0] w_n678_0;
	wire[1:0] w_n680_0;
	wire[1:0] w_n681_0;
	wire[1:0] w_n682_0;
	wire[1:0] w_n683_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n685_0;
	wire[1:0] w_n686_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n688_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n691_0;
	wire[1:0] w_n692_0;
	wire[1:0] w_n693_0;
	wire[1:0] w_n694_0;
	wire[1:0] w_n695_0;
	wire[1:0] w_n696_0;
	wire[1:0] w_n697_0;
	wire[1:0] w_n698_0;
	wire[1:0] w_n699_0;
	wire[1:0] w_n700_0;
	wire[1:0] w_n701_0;
	wire[1:0] w_n703_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n706_0;
	wire[1:0] w_n711_0;
	wire[1:0] w_n712_0;
	wire[2:0] w_n717_0;
	wire[1:0] w_n719_0;
	wire[1:0] w_n722_0;
	wire[1:0] w_n724_0;
	wire[1:0] w_n727_0;
	wire[1:0] w_n729_0;
	wire[1:0] w_n732_0;
	wire[1:0] w_n734_0;
	wire[1:0] w_n737_0;
	wire[1:0] w_n739_0;
	wire[1:0] w_n742_0;
	wire[1:0] w_n744_0;
	wire[1:0] w_n747_0;
	wire[1:0] w_n749_0;
	wire[1:0] w_n752_0;
	wire[1:0] w_n754_0;
	wire[1:0] w_n757_0;
	wire[1:0] w_n759_0;
	wire[1:0] w_n762_0;
	wire[1:0] w_n764_0;
	wire[1:0] w_n769_0;
	wire[1:0] w_n771_0;
	wire[1:0] w_n772_0;
	wire[1:0] w_n773_0;
	wire[1:0] w_n774_0;
	wire[1:0] w_n775_0;
	wire[1:0] w_n777_0;
	wire[1:0] w_n778_0;
	wire[1:0] w_n779_0;
	wire[1:0] w_n780_0;
	wire[1:0] w_n781_0;
	wire[1:0] w_n782_0;
	wire[1:0] w_n783_0;
	wire[1:0] w_n784_0;
	wire[1:0] w_n785_0;
	wire[1:0] w_n786_0;
	wire[1:0] w_n787_0;
	wire[1:0] w_n788_0;
	wire[1:0] w_n789_0;
	wire[1:0] w_n790_0;
	wire[1:0] w_n791_0;
	wire[1:0] w_n792_0;
	wire[1:0] w_n793_0;
	wire[1:0] w_n794_0;
	wire[1:0] w_n795_0;
	wire[1:0] w_n796_0;
	wire[1:0] w_n797_0;
	wire[1:0] w_n798_0;
	wire[1:0] w_n799_0;
	wire[1:0] w_n800_0;
	wire[1:0] w_n802_0;
	wire[1:0] w_n803_0;
	wire[1:0] w_n805_0;
	wire[1:0] w_n810_0;
	wire[1:0] w_n811_0;
	wire[1:0] w_n815_0;
	wire[1:0] w_n816_0;
	wire[2:0] w_n820_0;
	wire[1:0] w_n822_0;
	wire[1:0] w_n825_0;
	wire[1:0] w_n827_0;
	wire[1:0] w_n830_0;
	wire[1:0] w_n832_0;
	wire[1:0] w_n835_0;
	wire[1:0] w_n837_0;
	wire[1:0] w_n840_0;
	wire[1:0] w_n842_0;
	wire[1:0] w_n845_0;
	wire[1:0] w_n847_0;
	wire[1:0] w_n850_0;
	wire[1:0] w_n852_0;
	wire[1:0] w_n855_0;
	wire[1:0] w_n857_0;
	wire[1:0] w_n860_0;
	wire[1:0] w_n862_0;
	wire[1:0] w_n865_0;
	wire[1:0] w_n867_0;
	wire[1:0] w_n872_0;
	wire[1:0] w_n874_0;
	wire[1:0] w_n875_0;
	wire[1:0] w_n877_0;
	wire[1:0] w_n879_0;
	wire[1:0] w_n880_0;
	wire[1:0] w_n881_0;
	wire[1:0] w_n882_0;
	wire[1:0] w_n883_0;
	wire[1:0] w_n884_0;
	wire[1:0] w_n885_0;
	wire[1:0] w_n886_0;
	wire[1:0] w_n887_0;
	wire[1:0] w_n888_0;
	wire[1:0] w_n889_0;
	wire[1:0] w_n890_0;
	wire[1:0] w_n891_0;
	wire[1:0] w_n892_0;
	wire[1:0] w_n893_0;
	wire[1:0] w_n894_0;
	wire[1:0] w_n895_0;
	wire[1:0] w_n896_0;
	wire[1:0] w_n897_0;
	wire[1:0] w_n898_0;
	wire[1:0] w_n899_0;
	wire[2:0] w_n900_0;
	wire[1:0] w_n902_0;
	wire[1:0] w_n903_0;
	wire[1:0] w_n904_0;
	wire[1:0] w_n905_0;
	wire[1:0] w_n910_0;
	wire[1:0] w_n911_0;
	wire[2:0] w_n915_0;
	wire[1:0] w_n916_0;
	wire[1:0] w_n922_0;
	wire[1:0] w_n924_0;
	wire[1:0] w_n927_0;
	wire[1:0] w_n929_0;
	wire[1:0] w_n932_0;
	wire[1:0] w_n934_0;
	wire[1:0] w_n937_0;
	wire[1:0] w_n939_0;
	wire[1:0] w_n942_0;
	wire[1:0] w_n944_0;
	wire[1:0] w_n947_0;
	wire[1:0] w_n949_0;
	wire[1:0] w_n952_0;
	wire[1:0] w_n954_0;
	wire[1:0] w_n957_0;
	wire[1:0] w_n959_0;
	wire[1:0] w_n962_0;
	wire[1:0] w_n964_0;
	wire[1:0] w_n967_0;
	wire[1:0] w_n969_0;
	wire[1:0] w_n972_0;
	wire[1:0] w_n974_0;
	wire[1:0] w_n978_0;
	wire[1:0] w_n980_0;
	wire[1:0] w_n982_0;
	wire[1:0] w_n983_0;
	wire[1:0] w_n984_0;
	wire[1:0] w_n985_0;
	wire[1:0] w_n986_0;
	wire[1:0] w_n987_0;
	wire[1:0] w_n988_0;
	wire[1:0] w_n989_0;
	wire[1:0] w_n990_0;
	wire[1:0] w_n991_0;
	wire[1:0] w_n992_0;
	wire[1:0] w_n993_0;
	wire[1:0] w_n994_0;
	wire[1:0] w_n995_0;
	wire[1:0] w_n996_0;
	wire[1:0] w_n997_0;
	wire[1:0] w_n998_0;
	wire[1:0] w_n999_0;
	wire[1:0] w_n1000_0;
	wire[1:0] w_n1001_0;
	wire[1:0] w_n1002_0;
	wire[1:0] w_n1003_0;
	wire[1:0] w_n1004_0;
	wire[1:0] w_n1005_0;
	wire[1:0] w_n1006_0;
	wire[1:0] w_n1007_0;
	wire[1:0] w_n1008_0;
	wire[1:0] w_n1009_0;
	wire[1:0] w_n1011_0;
	wire[1:0] w_n1013_0;
	wire[1:0] w_n1017_0;
	wire[1:0] w_n1018_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1023_0;
	wire[1:0] w_n1026_0;
	wire[1:0] w_n1028_0;
	wire[1:0] w_n1031_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1036_0;
	wire[1:0] w_n1038_0;
	wire[1:0] w_n1041_0;
	wire[1:0] w_n1043_0;
	wire[1:0] w_n1046_0;
	wire[1:0] w_n1048_0;
	wire[1:0] w_n1051_0;
	wire[1:0] w_n1053_0;
	wire[1:0] w_n1056_0;
	wire[1:0] w_n1058_0;
	wire[1:0] w_n1061_0;
	wire[1:0] w_n1063_0;
	wire[1:0] w_n1066_0;
	wire[1:0] w_n1068_0;
	wire[1:0] w_n1071_0;
	wire[1:0] w_n1073_0;
	wire[1:0] w_n1076_0;
	wire[1:0] w_n1077_0;
	wire[1:0] w_n1078_0;
	wire[1:0] w_n1080_0;
	wire[1:0] w_n1082_0;
	wire[1:0] w_n1083_0;
	wire[1:0] w_n1084_0;
	wire[1:0] w_n1085_0;
	wire[1:0] w_n1086_0;
	wire[1:0] w_n1087_0;
	wire[1:0] w_n1088_0;
	wire[1:0] w_n1089_0;
	wire[1:0] w_n1090_0;
	wire[1:0] w_n1091_0;
	wire[1:0] w_n1092_0;
	wire[1:0] w_n1093_0;
	wire[1:0] w_n1094_0;
	wire[1:0] w_n1095_0;
	wire[1:0] w_n1096_0;
	wire[1:0] w_n1097_0;
	wire[1:0] w_n1098_0;
	wire[1:0] w_n1099_0;
	wire[1:0] w_n1100_0;
	wire[1:0] w_n1101_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1103_0;
	wire[1:0] w_n1105_0;
	wire[1:0] w_n1106_0;
	wire[1:0] w_n1107_0;
	wire[1:0] w_n1108_0;
	wire[1:0] w_n1109_0;
	wire[1:0] w_n1115_0;
	wire[1:0] w_n1119_0;
	wire[1:0] w_n1120_0;
	wire[1:0] w_n1124_0;
	wire[1:0] w_n1126_0;
	wire[1:0] w_n1129_0;
	wire[1:0] w_n1131_0;
	wire[1:0] w_n1134_0;
	wire[1:0] w_n1136_0;
	wire[1:0] w_n1139_0;
	wire[1:0] w_n1141_0;
	wire[1:0] w_n1144_0;
	wire[1:0] w_n1146_0;
	wire[1:0] w_n1149_0;
	wire[1:0] w_n1151_0;
	wire[1:0] w_n1154_0;
	wire[1:0] w_n1156_0;
	wire[1:0] w_n1159_0;
	wire[1:0] w_n1161_0;
	wire[1:0] w_n1164_0;
	wire[1:0] w_n1166_0;
	wire[1:0] w_n1169_0;
	wire[1:0] w_n1171_0;
	wire[1:0] w_n1174_0;
	wire[1:0] w_n1175_0;
	wire[1:0] w_n1176_0;
	wire[1:0] w_n1179_0;
	wire[1:0] w_n1181_0;
	wire[1:0] w_n1182_0;
	wire[1:0] w_n1183_0;
	wire[1:0] w_n1184_0;
	wire[1:0] w_n1185_0;
	wire[1:0] w_n1186_0;
	wire[1:0] w_n1187_0;
	wire[1:0] w_n1188_0;
	wire[1:0] w_n1189_0;
	wire[1:0] w_n1190_0;
	wire[1:0] w_n1191_0;
	wire[1:0] w_n1192_0;
	wire[1:0] w_n1193_0;
	wire[1:0] w_n1194_0;
	wire[1:0] w_n1195_0;
	wire[1:0] w_n1196_0;
	wire[1:0] w_n1197_0;
	wire[1:0] w_n1198_0;
	wire[1:0] w_n1199_0;
	wire[1:0] w_n1200_0;
	wire[1:0] w_n1201_0;
	wire[1:0] w_n1203_0;
	wire[1:0] w_n1205_0;
	wire[1:0] w_n1206_0;
	wire[1:0] w_n1207_0;
	wire[1:0] w_n1213_0;
	wire[1:0] w_n1216_0;
	wire[1:0] w_n1217_0;
	wire[1:0] w_n1220_0;
	wire[1:0] w_n1222_0;
	wire[1:0] w_n1225_0;
	wire[1:0] w_n1227_0;
	wire[1:0] w_n1230_0;
	wire[1:0] w_n1232_0;
	wire[1:0] w_n1235_0;
	wire[1:0] w_n1237_0;
	wire[1:0] w_n1240_0;
	wire[1:0] w_n1242_0;
	wire[1:0] w_n1245_0;
	wire[1:0] w_n1247_0;
	wire[1:0] w_n1250_0;
	wire[1:0] w_n1252_0;
	wire[1:0] w_n1255_0;
	wire[1:0] w_n1257_0;
	wire[1:0] w_n1260_0;
	wire[1:0] w_n1262_0;
	wire[1:0] w_n1265_0;
	wire[1:0] w_n1266_0;
	wire[1:0] w_n1267_0;
	wire[1:0] w_n1270_0;
	wire[1:0] w_n1272_0;
	wire[1:0] w_n1273_0;
	wire[1:0] w_n1274_0;
	wire[1:0] w_n1275_0;
	wire[1:0] w_n1276_0;
	wire[1:0] w_n1277_0;
	wire[1:0] w_n1278_0;
	wire[1:0] w_n1279_0;
	wire[1:0] w_n1280_0;
	wire[1:0] w_n1281_0;
	wire[1:0] w_n1282_0;
	wire[1:0] w_n1283_0;
	wire[1:0] w_n1284_0;
	wire[1:0] w_n1285_0;
	wire[1:0] w_n1286_0;
	wire[1:0] w_n1287_0;
	wire[1:0] w_n1288_0;
	wire[1:0] w_n1289_0;
	wire[1:0] w_n1290_0;
	wire[1:0] w_n1291_0;
	wire[1:0] w_n1293_0;
	wire[1:0] w_n1294_0;
	wire[1:0] w_n1295_0;
	wire[1:0] w_n1301_0;
	wire[1:0] w_n1306_0;
	wire[1:0] w_n1307_0;
	wire[1:0] w_n1310_0;
	wire[1:0] w_n1312_0;
	wire[1:0] w_n1315_0;
	wire[1:0] w_n1317_0;
	wire[1:0] w_n1320_0;
	wire[1:0] w_n1322_0;
	wire[1:0] w_n1325_0;
	wire[1:0] w_n1327_0;
	wire[1:0] w_n1330_0;
	wire[1:0] w_n1332_0;
	wire[1:0] w_n1335_0;
	wire[1:0] w_n1337_0;
	wire[1:0] w_n1340_0;
	wire[1:0] w_n1342_0;
	wire[1:0] w_n1345_0;
	wire[1:0] w_n1347_0;
	wire[1:0] w_n1350_0;
	wire[1:0] w_n1351_0;
	wire[1:0] w_n1352_0;
	wire[1:0] w_n1355_0;
	wire[1:0] w_n1357_0;
	wire[1:0] w_n1358_0;
	wire[1:0] w_n1359_0;
	wire[1:0] w_n1360_0;
	wire[1:0] w_n1361_0;
	wire[1:0] w_n1362_0;
	wire[1:0] w_n1363_0;
	wire[1:0] w_n1364_0;
	wire[1:0] w_n1365_0;
	wire[1:0] w_n1366_0;
	wire[1:0] w_n1367_0;
	wire[1:0] w_n1368_0;
	wire[1:0] w_n1369_0;
	wire[1:0] w_n1370_0;
	wire[1:0] w_n1371_0;
	wire[1:0] w_n1372_0;
	wire[1:0] w_n1373_0;
	wire[1:0] w_n1374_0;
	wire[1:0] w_n1376_0;
	wire[1:0] w_n1378_0;
	wire[1:0] w_n1379_0;
	wire[1:0] w_n1384_0;
	wire[1:0] w_n1389_0;
	wire[1:0] w_n1390_0;
	wire[1:0] w_n1393_0;
	wire[1:0] w_n1395_0;
	wire[1:0] w_n1398_0;
	wire[1:0] w_n1400_0;
	wire[1:0] w_n1403_0;
	wire[1:0] w_n1405_0;
	wire[1:0] w_n1408_0;
	wire[1:0] w_n1410_0;
	wire[1:0] w_n1413_0;
	wire[1:0] w_n1415_0;
	wire[1:0] w_n1418_0;
	wire[1:0] w_n1420_0;
	wire[1:0] w_n1423_0;
	wire[1:0] w_n1425_0;
	wire[1:0] w_n1428_0;
	wire[1:0] w_n1429_0;
	wire[1:0] w_n1430_0;
	wire[1:0] w_n1433_0;
	wire[1:0] w_n1435_0;
	wire[1:0] w_n1436_0;
	wire[1:0] w_n1437_0;
	wire[1:0] w_n1438_0;
	wire[1:0] w_n1439_0;
	wire[1:0] w_n1440_0;
	wire[1:0] w_n1441_0;
	wire[1:0] w_n1442_0;
	wire[1:0] w_n1443_0;
	wire[1:0] w_n1444_0;
	wire[1:0] w_n1445_0;
	wire[1:0] w_n1446_0;
	wire[1:0] w_n1447_0;
	wire[1:0] w_n1448_0;
	wire[1:0] w_n1449_0;
	wire[1:0] w_n1450_0;
	wire[1:0] w_n1452_0;
	wire[1:0] w_n1454_0;
	wire[1:0] w_n1455_0;
	wire[1:0] w_n1460_0;
	wire[1:0] w_n1465_0;
	wire[1:0] w_n1466_0;
	wire[1:0] w_n1469_0;
	wire[1:0] w_n1471_0;
	wire[1:0] w_n1474_0;
	wire[1:0] w_n1476_0;
	wire[1:0] w_n1479_0;
	wire[1:0] w_n1481_0;
	wire[1:0] w_n1484_0;
	wire[1:0] w_n1486_0;
	wire[1:0] w_n1489_0;
	wire[1:0] w_n1491_0;
	wire[1:0] w_n1494_0;
	wire[1:0] w_n1496_0;
	wire[1:0] w_n1499_0;
	wire[1:0] w_n1500_0;
	wire[1:0] w_n1501_0;
	wire[1:0] w_n1504_0;
	wire[1:0] w_n1506_0;
	wire[1:0] w_n1507_0;
	wire[1:0] w_n1508_0;
	wire[1:0] w_n1509_0;
	wire[1:0] w_n1510_0;
	wire[1:0] w_n1511_0;
	wire[1:0] w_n1512_0;
	wire[1:0] w_n1513_0;
	wire[1:0] w_n1514_0;
	wire[1:0] w_n1515_0;
	wire[1:0] w_n1516_0;
	wire[1:0] w_n1517_0;
	wire[1:0] w_n1518_0;
	wire[1:0] w_n1519_0;
	wire[1:0] w_n1521_0;
	wire[1:0] w_n1523_0;
	wire[1:0] w_n1524_0;
	wire[1:0] w_n1529_0;
	wire[1:0] w_n1534_0;
	wire[1:0] w_n1535_0;
	wire[1:0] w_n1538_0;
	wire[1:0] w_n1540_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1545_0;
	wire[1:0] w_n1548_0;
	wire[1:0] w_n1550_0;
	wire[1:0] w_n1553_0;
	wire[1:0] w_n1555_0;
	wire[1:0] w_n1558_0;
	wire[1:0] w_n1560_0;
	wire[1:0] w_n1563_0;
	wire[1:0] w_n1564_0;
	wire[1:0] w_n1565_0;
	wire[1:0] w_n1568_0;
	wire[1:0] w_n1570_0;
	wire[1:0] w_n1571_0;
	wire[1:0] w_n1572_0;
	wire[1:0] w_n1573_0;
	wire[1:0] w_n1574_0;
	wire[1:0] w_n1575_0;
	wire[1:0] w_n1576_0;
	wire[1:0] w_n1577_0;
	wire[1:0] w_n1578_0;
	wire[1:0] w_n1579_0;
	wire[1:0] w_n1580_0;
	wire[1:0] w_n1581_0;
	wire[1:0] w_n1583_0;
	wire[1:0] w_n1585_0;
	wire[1:0] w_n1586_0;
	wire[1:0] w_n1591_0;
	wire[1:0] w_n1596_0;
	wire[1:0] w_n1597_0;
	wire[1:0] w_n1600_0;
	wire[1:0] w_n1602_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1607_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1612_0;
	wire[1:0] w_n1615_0;
	wire[1:0] w_n1617_0;
	wire[1:0] w_n1620_0;
	wire[1:0] w_n1621_0;
	wire[1:0] w_n1622_0;
	wire[1:0] w_n1625_0;
	wire[1:0] w_n1627_0;
	wire[1:0] w_n1628_0;
	wire[1:0] w_n1629_0;
	wire[1:0] w_n1630_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1632_0;
	wire[1:0] w_n1633_0;
	wire[1:0] w_n1634_0;
	wire[1:0] w_n1635_0;
	wire[1:0] w_n1636_0;
	wire[1:0] w_n1638_0;
	wire[1:0] w_n1640_0;
	wire[1:0] w_n1641_0;
	wire[1:0] w_n1646_0;
	wire[1:0] w_n1651_0;
	wire[1:0] w_n1653_0;
	wire[1:0] w_n1656_0;
	wire[1:0] w_n1658_0;
	wire[1:0] w_n1661_0;
	wire[1:0] w_n1663_0;
	wire[1:0] w_n1666_0;
	wire[1:0] w_n1668_0;
	wire[1:0] w_n1671_0;
	wire[1:0] w_n1672_0;
	wire[1:0] w_n1673_0;
	wire[1:0] w_n1676_0;
	wire[1:0] w_n1678_0;
	wire[1:0] w_n1679_0;
	wire[1:0] w_n1680_0;
	wire[1:0] w_n1681_0;
	wire[1:0] w_n1682_0;
	wire[1:0] w_n1683_0;
	wire[1:0] w_n1684_0;
	wire[1:0] w_n1685_0;
	wire[1:0] w_n1686_0;
	wire[1:0] w_n1688_0;
	wire[1:0] w_n1689_0;
	wire[1:0] w_n1694_0;
	wire[1:0] w_n1697_0;
	wire[1:0] w_n1699_0;
	wire[1:0] w_n1702_0;
	wire[1:0] w_n1704_0;
	wire[1:0] w_n1707_0;
	wire[1:0] w_n1709_0;
	wire[1:0] w_n1712_0;
	wire[1:0] w_n1713_0;
	wire[1:0] w_n1714_0;
	wire[1:0] w_n1717_0;
	wire[1:0] w_n1719_0;
	wire[1:0] w_n1720_0;
	wire[1:0] w_n1721_0;
	wire[1:0] w_n1722_0;
	wire[1:0] w_n1723_0;
	wire[1:0] w_n1724_0;
	wire[1:0] w_n1725_0;
	wire[1:0] w_n1726_0;
	wire[1:0] w_n1727_0;
	wire[1:0] w_n1734_0;
	wire[1:0] w_n1737_0;
	wire[1:0] w_n1739_0;
	wire[1:0] w_n1742_0;
	wire[1:0] w_n1744_0;
	wire[1:0] w_n1747_0;
	wire[1:0] w_n1748_0;
	wire[1:0] w_n1749_0;
	wire[1:0] w_n1752_0;
	wire[1:0] w_n1754_0;
	wire[1:0] w_n1755_0;
	wire[1:0] w_n1756_0;
	wire[1:0] w_n1757_0;
	wire[1:0] w_n1758_0;
	wire[1:0] w_n1759_0;
	wire[1:0] w_n1760_0;
	wire[1:0] w_n1767_0;
	wire[1:0] w_n1770_0;
	wire[1:0] w_n1772_0;
	wire[1:0] w_n1775_0;
	wire[1:0] w_n1776_0;
	wire[1:0] w_n1777_0;
	wire[1:0] w_n1780_0;
	wire[1:0] w_n1782_0;
	wire[1:0] w_n1783_0;
	wire[1:0] w_n1784_0;
	wire[1:0] w_n1785_0;
	wire[1:0] w_n1786_0;
	wire[1:0] w_n1793_0;
	wire[1:0] w_n1796_0;
	wire[1:0] w_n1797_0;
	wire[1:0] w_n1798_0;
	wire[1:0] w_n1801_0;
	wire[1:0] w_n1803_0;
	wire[1:0] w_n1804_0;
	wire[1:0] w_n1805_0;
	wire[1:0] w_n1807_0;
	wire[1:0] w_n1810_0;
	wire[1:0] w_n1817_0;
	wire[1:0] w_n1818_0;
	wire w_dff_B_6EbCXpH77_0;
	wire w_dff_B_xtZmTHUA1_0;
	wire w_dff_B_8eVh8Wnb7_1;
	wire w_dff_B_4JcfhAzb9_1;
	wire w_dff_B_c1j5Gyez3_1;
	wire w_dff_B_PVNT4aGx9_1;
	wire w_dff_B_JaUmz1Va5_1;
	wire w_dff_B_S7dPF5m53_1;
	wire w_dff_B_s7M86MFT7_1;
	wire w_dff_B_1KvYvi7e1_1;
	wire w_dff_B_TnLU4N4R5_1;
	wire w_dff_B_FS2Gflch8_1;
	wire w_dff_B_bTw3ySpl4_1;
	wire w_dff_B_fKN0GiF25_1;
	wire w_dff_B_NvRmulmG2_1;
	wire w_dff_B_FEOzBdld7_1;
	wire w_dff_B_GtpBJpdl5_1;
	wire w_dff_B_trBLxzOo0_1;
	wire w_dff_B_TuXcG4bf5_1;
	wire w_dff_B_2bca4tz20_1;
	wire w_dff_B_fY7JYVwV5_1;
	wire w_dff_B_f80I4H8v9_1;
	wire w_dff_B_n56lUK196_1;
	wire w_dff_B_EfJA0pmZ5_1;
	wire w_dff_B_i89h6el13_1;
	wire w_dff_B_9opOCRek1_1;
	wire w_dff_B_uAw445A47_1;
	wire w_dff_B_6SLWFlgP9_1;
	wire w_dff_B_SoefDKPz1_1;
	wire w_dff_B_WDui7EWV9_1;
	wire w_dff_B_UqUZaCXs4_1;
	wire w_dff_B_M3AxJSlC9_1;
	wire w_dff_B_LFYlq8cZ0_1;
	wire w_dff_B_VKDa8BD95_1;
	wire w_dff_B_B9rGcLtU8_1;
	wire w_dff_B_hTuES3dj1_1;
	wire w_dff_B_v9F38lDU3_1;
	wire w_dff_B_Hx7aAZiW0_1;
	wire w_dff_B_tN1jq0LE5_1;
	wire w_dff_B_KvRtTdHc6_1;
	wire w_dff_B_jrQjBfkc6_1;
	wire w_dff_B_ob4NYxlA0_1;
	wire w_dff_B_N65PrVWl8_1;
	wire w_dff_B_eSr03Dgt7_1;
	wire w_dff_B_daeICTUl4_1;
	wire w_dff_B_J8n7Q3YB3_1;
	wire w_dff_B_DOxgFj537_1;
	wire w_dff_B_StChmr9P4_1;
	wire w_dff_B_YMTpwJuY0_1;
	wire w_dff_B_tmoHPFN09_1;
	wire w_dff_B_yCjB3KRH9_1;
	wire w_dff_B_YZCWiTtL4_1;
	wire w_dff_B_VWRvGCNO2_1;
	wire w_dff_B_uVSwz0Lu1_1;
	wire w_dff_B_cTW4zgFp8_1;
	wire w_dff_B_SGk1TWIE0_1;
	wire w_dff_B_zVogGwtN2_1;
	wire w_dff_B_uOGSDFNo5_1;
	wire w_dff_B_RGfjPcz20_1;
	wire w_dff_B_MTuAQUhG6_1;
	wire w_dff_B_igP4oBDl2_1;
	wire w_dff_B_mi7TkSlU3_1;
	wire w_dff_B_P7CtA1N89_1;
	wire w_dff_B_4pcr0ilK7_1;
	wire w_dff_B_DtxLqxqv7_1;
	wire w_dff_B_SgOCHxAj6_1;
	wire w_dff_B_O3FUU1Ss4_1;
	wire w_dff_B_cyUrzFXY2_1;
	wire w_dff_B_ylPbca7d0_1;
	wire w_dff_B_TezgXW8k5_1;
	wire w_dff_B_chzPvfiq8_1;
	wire w_dff_B_8FA1HqLd1_1;
	wire w_dff_B_9HKf2dSi8_1;
	wire w_dff_B_WbfZrgI67_1;
	wire w_dff_B_3gWwstnp9_1;
	wire w_dff_B_L9SJeKrO7_1;
	wire w_dff_B_LrxxM1bT3_1;
	wire w_dff_B_Cb1wrOak1_1;
	wire w_dff_B_SgKKyl412_1;
	wire w_dff_B_eRwawQsp9_1;
	wire w_dff_B_teDoWhVc9_1;
	wire w_dff_B_xEctTbmu9_1;
	wire w_dff_B_xDzWTUSH9_1;
	wire w_dff_B_XI4hWen59_1;
	wire w_dff_B_dxTOxvBm1_1;
	wire w_dff_B_8TdGlqOt4_1;
	wire w_dff_B_xCe6rYqH2_1;
	wire w_dff_B_rCfwRgoe0_1;
	wire w_dff_B_7xNDPKNx3_1;
	wire w_dff_B_rraDYe3f2_1;
	wire w_dff_B_OZGA47qO8_1;
	wire w_dff_B_cXrSdBwG7_1;
	wire w_dff_B_24VQ7H7T1_1;
	wire w_dff_B_vgfrHnC17_1;
	wire w_dff_B_lwok5KC89_1;
	wire w_dff_B_SiyGT3On8_1;
	wire w_dff_B_Zmoc0Eb75_1;
	wire w_dff_B_67vY2LXH8_1;
	wire w_dff_B_XtFc66aC5_1;
	wire w_dff_B_nX6DvFbs7_1;
	wire w_dff_B_kwkp0b7E2_1;
	wire w_dff_B_zbV1xpA51_1;
	wire w_dff_B_0aJaneqd6_1;
	wire w_dff_B_QwSxNmHY6_1;
	wire w_dff_B_wcTbZlve2_1;
	wire w_dff_B_mf6fPMF03_1;
	wire w_dff_B_l1VaZjya2_1;
	wire w_dff_B_h6EyVqVB2_1;
	wire w_dff_B_WhgrDOYv4_1;
	wire w_dff_B_KsiC9Zr79_1;
	wire w_dff_B_w2Qpxdxx9_1;
	wire w_dff_B_Zog4Q74K6_1;
	wire w_dff_B_0WgXiZAG4_1;
	wire w_dff_B_KJF7FvIw6_1;
	wire w_dff_B_qSq7upvm6_1;
	wire w_dff_B_AoCZsmiq2_1;
	wire w_dff_B_TrGx3jis2_1;
	wire w_dff_B_bJzNGOuL6_1;
	wire w_dff_B_rZeSt5sL0_1;
	wire w_dff_B_DI6sVi8z2_1;
	wire w_dff_B_rR0d9lqD3_1;
	wire w_dff_B_UnQyhgqA3_1;
	wire w_dff_B_vVH6eMGy7_1;
	wire w_dff_B_UHLQIkvA8_1;
	wire w_dff_B_33uwKasO8_1;
	wire w_dff_B_wRKtgU1X9_1;
	wire w_dff_B_6JIsAdm45_1;
	wire w_dff_B_9jo6SD158_1;
	wire w_dff_B_zRaMeYca5_1;
	wire w_dff_B_rpHuyIUg3_1;
	wire w_dff_B_HbSSAAja9_1;
	wire w_dff_B_0znk2DEo2_1;
	wire w_dff_B_uHQTjcxB3_1;
	wire w_dff_B_5SPzbTGA3_1;
	wire w_dff_B_j8pjpo9R2_1;
	wire w_dff_B_kpQP77Kr2_1;
	wire w_dff_B_IFgWrum80_1;
	wire w_dff_B_hL3LG6ve1_1;
	wire w_dff_B_MLkfyhYU5_1;
	wire w_dff_B_BaIaZgFE3_1;
	wire w_dff_B_75WEGCHR1_1;
	wire w_dff_B_1uv7rtZ97_1;
	wire w_dff_B_tT19Tmhp3_1;
	wire w_dff_B_OFGr9D4e7_1;
	wire w_dff_B_zQ3WILTG6_1;
	wire w_dff_B_rPoMADEC8_1;
	wire w_dff_B_WY1oUXNV4_1;
	wire w_dff_B_4JHhzcGh9_1;
	wire w_dff_B_B5oNP1057_1;
	wire w_dff_B_3gks9b4i8_1;
	wire w_dff_B_1ckkkLVM2_1;
	wire w_dff_B_7JVYq7Mk8_1;
	wire w_dff_B_ObFOKFSt2_1;
	wire w_dff_B_N9xsphSB1_1;
	wire w_dff_B_Fs67pSzw2_1;
	wire w_dff_B_TdIJWCCK2_1;
	wire w_dff_B_34XUerzc0_1;
	wire w_dff_B_HQdnTf2A0_1;
	wire w_dff_B_HuzeMcf21_1;
	wire w_dff_B_1YffoFRi6_1;
	wire w_dff_B_7yiP9aLU6_1;
	wire w_dff_B_uEJ6x5EK0_1;
	wire w_dff_B_3Kb2MUQu2_1;
	wire w_dff_B_gSd35X2k7_1;
	wire w_dff_B_agLT5Mwy1_1;
	wire w_dff_B_xIMHMpsd0_1;
	wire w_dff_B_EX4MsRm61_1;
	wire w_dff_B_3p8ppx9t4_1;
	wire w_dff_B_fxhoKKHk4_1;
	wire w_dff_B_zDZM7NoD7_1;
	wire w_dff_B_Rp9MfLq09_1;
	wire w_dff_B_R9PHrWSQ6_1;
	wire w_dff_B_4kLT5PFC5_1;
	wire w_dff_B_O5TH56fR5_1;
	wire w_dff_B_vfzUTUFM7_1;
	wire w_dff_B_zvgPJBZK6_1;
	wire w_dff_B_nkxQ0gpm5_1;
	wire w_dff_B_EBR7MLPw5_1;
	wire w_dff_B_srhPxAMg8_1;
	wire w_dff_B_WSXMOyrr6_1;
	wire w_dff_B_ojdXWzes0_1;
	wire w_dff_B_nYSBzpuP9_1;
	wire w_dff_B_ZmSne4aQ9_1;
	wire w_dff_B_tNebJp1A7_1;
	wire w_dff_B_M3dJ2zW73_1;
	wire w_dff_B_K7wUEF2I0_1;
	wire w_dff_B_0AoavkzU9_1;
	wire w_dff_B_fCzMoOLC1_1;
	wire w_dff_B_0UaRtaB64_1;
	wire w_dff_B_2NxIlVfb1_1;
	wire w_dff_B_mSUjF4GK0_1;
	wire w_dff_B_b53IuW9w5_1;
	wire w_dff_B_29gJcb3l1_1;
	wire w_dff_B_cLYYZ00k1_1;
	wire w_dff_B_JIXTNkLI7_1;
	wire w_dff_B_UW2U5ROp9_1;
	wire w_dff_B_frlRyrlY4_1;
	wire w_dff_B_9Mjys5ry7_1;
	wire w_dff_B_idv9ebLc1_1;
	wire w_dff_B_pnCMdMee4_1;
	wire w_dff_B_ddCYsK5h7_1;
	wire w_dff_B_4z9tfpSV2_1;
	wire w_dff_B_8Onkcvdh3_1;
	wire w_dff_B_mtf9P8PM2_1;
	wire w_dff_B_nBpGjsSK1_1;
	wire w_dff_B_BfZGTwG56_1;
	wire w_dff_B_tNJjdQ0I7_1;
	wire w_dff_B_zs2J7dza5_1;
	wire w_dff_B_1OXU5V3c8_1;
	wire w_dff_B_Vn73s0514_1;
	wire w_dff_B_7wbDTtQ59_1;
	wire w_dff_B_73Dquhxd4_1;
	wire w_dff_B_i95YsMrf5_1;
	wire w_dff_B_iA3P04ht0_1;
	wire w_dff_B_D8gh3Ruy1_1;
	wire w_dff_B_yky5UjuC0_1;
	wire w_dff_B_2kNdDtiR9_1;
	wire w_dff_B_iV5peYyX9_1;
	wire w_dff_B_bsa4ROoh9_1;
	wire w_dff_B_x0GZNjDs1_1;
	wire w_dff_B_SmWZzYXj4_1;
	wire w_dff_B_XV0VQKRM7_1;
	wire w_dff_B_yhEWxIyq7_1;
	wire w_dff_B_RrWDctnL6_1;
	wire w_dff_B_PluXWITn0_1;
	wire w_dff_B_8wW7V9P29_1;
	wire w_dff_B_1ouMGPOL5_1;
	wire w_dff_B_j8SJs5rv6_1;
	wire w_dff_B_MWqaKIe18_1;
	wire w_dff_B_YDf0bTE60_1;
	wire w_dff_B_t31VFgcK7_1;
	wire w_dff_B_q5vUMTHS7_1;
	wire w_dff_B_TBpCQkxo8_1;
	wire w_dff_B_Fq5TI8J04_1;
	wire w_dff_B_vSmBcOzN5_1;
	wire w_dff_B_55BBytC33_1;
	wire w_dff_B_9I11JogR9_1;
	wire w_dff_B_AczLivBM5_1;
	wire w_dff_B_6UpP73mP7_1;
	wire w_dff_B_qqD2Z0GD4_1;
	wire w_dff_B_aKmwxaI15_1;
	wire w_dff_B_QWwkQPb75_1;
	wire w_dff_B_0X2NQNbV7_1;
	wire w_dff_B_jn8UXZli3_1;
	wire w_dff_B_c1wNrggv4_1;
	wire w_dff_B_MITQI8gI8_1;
	wire w_dff_B_ObkCXsxe1_1;
	wire w_dff_B_SWQIp7Rq1_1;
	wire w_dff_B_roRCwGpq1_1;
	wire w_dff_B_PRyxs9Dj8_1;
	wire w_dff_B_iBKZ7qDt8_1;
	wire w_dff_B_K23hHub09_1;
	wire w_dff_B_P2U5OV9H9_1;
	wire w_dff_B_eueJfIIM9_1;
	wire w_dff_B_kot1wLEQ6_1;
	wire w_dff_B_2yBF3vGT2_1;
	wire w_dff_B_2MrJYv3v0_1;
	wire w_dff_B_gzHQXFjs7_1;
	wire w_dff_B_6lrXfArB8_1;
	wire w_dff_B_WgenlHKS4_1;
	wire w_dff_B_ogke7o653_1;
	wire w_dff_B_AKE6WBgO2_1;
	wire w_dff_B_6JcvkoBn3_1;
	wire w_dff_B_qjWchHdH6_1;
	wire w_dff_B_MOYeTtWB8_1;
	wire w_dff_B_Y08ZnuLG5_1;
	wire w_dff_B_71asyolI3_1;
	wire w_dff_B_D3qyxekF7_1;
	wire w_dff_B_aG0sMuV34_1;
	wire w_dff_B_B5hEKQXo3_1;
	wire w_dff_B_GG58iKfq2_1;
	wire w_dff_B_Xzqg8oJW5_1;
	wire w_dff_B_wga2OkXR9_1;
	wire w_dff_B_cZs1tC6j0_1;
	wire w_dff_B_9PkQ9nLG0_1;
	wire w_dff_B_UOySr02X9_1;
	wire w_dff_B_xGqX2sE21_1;
	wire w_dff_B_hIGWddNj8_1;
	wire w_dff_B_tBfiJ1sl4_1;
	wire w_dff_B_zzDAoTbl5_1;
	wire w_dff_B_gHVAWJCW3_1;
	wire w_dff_B_WJFtzMZc2_1;
	wire w_dff_B_xwIMkggk6_1;
	wire w_dff_B_QSLkstkU3_1;
	wire w_dff_B_T1fAoUum7_1;
	wire w_dff_B_dmQa6sMh3_1;
	wire w_dff_B_vr3m0T0t7_1;
	wire w_dff_B_vGHD0Xx13_1;
	wire w_dff_B_W1TAUOEO5_1;
	wire w_dff_B_7WD94D5C1_1;
	wire w_dff_B_yN4pr8wP4_1;
	wire w_dff_B_nTaNbPTO9_1;
	wire w_dff_B_Wcuhr3UH6_1;
	wire w_dff_B_1XCLyNpe8_1;
	wire w_dff_B_lFU5vpFS0_1;
	wire w_dff_B_GJR6hA603_1;
	wire w_dff_B_bY96qWr99_1;
	wire w_dff_B_kuFOyRvF2_1;
	wire w_dff_B_5njfu8GU9_1;
	wire w_dff_B_XhcR2aI06_1;
	wire w_dff_B_PYlWTWKm4_1;
	wire w_dff_B_czH6LOmf5_1;
	wire w_dff_B_q6H1cXHd1_1;
	wire w_dff_B_GxMtINvE2_1;
	wire w_dff_B_M3T1LsCC7_1;
	wire w_dff_B_K47AOfHv3_1;
	wire w_dff_B_xiPhMNUX8_1;
	wire w_dff_B_P7WUDUBO1_1;
	wire w_dff_B_pUbvCtGT7_1;
	wire w_dff_B_ca9BPqXR7_1;
	wire w_dff_B_KBceVWwJ8_1;
	wire w_dff_B_XNQTM6Mn1_1;
	wire w_dff_B_yMcaZczD9_1;
	wire w_dff_B_s4E0WcHW3_1;
	wire w_dff_B_dUWNQoQB4_1;
	wire w_dff_B_kwbDSW4F8_1;
	wire w_dff_B_mW8Cwltp4_1;
	wire w_dff_B_7zYdlvs98_0;
	wire w_dff_B_7EpvMSVl5_1;
	wire w_dff_B_T6QCaNef3_1;
	wire w_dff_B_3XDMxnoE8_1;
	wire w_dff_B_kPASAC0t9_1;
	wire w_dff_B_bjPfQZns6_1;
	wire w_dff_B_nKcYsWBE6_1;
	wire w_dff_B_SksbWreh9_1;
	wire w_dff_B_Ya9DTWMv0_1;
	wire w_dff_B_mtOLx1JO5_1;
	wire w_dff_B_3zryJO885_1;
	wire w_dff_B_FPGRGM5T4_1;
	wire w_dff_B_A6LMD9Hy5_1;
	wire w_dff_B_eSTj5NJB6_1;
	wire w_dff_B_yjNaL4ch6_1;
	wire w_dff_B_phOQFaYs1_1;
	wire w_dff_B_sKBpYG7w6_0;
	wire w_dff_B_c7PyV10g3_0;
	wire w_dff_B_zlCXqYP15_0;
	wire w_dff_B_1m7bE9rQ8_0;
	wire w_dff_B_xobmftXj2_0;
	wire w_dff_B_PIwlu7vU0_0;
	wire w_dff_B_Jfgx368K5_0;
	wire w_dff_B_R9dJDjgQ8_0;
	wire w_dff_B_OSBjIakL5_0;
	wire w_dff_B_nsM6fSXT6_0;
	wire w_dff_B_Y2HbigHG2_0;
	wire w_dff_B_QYDhjXC85_0;
	wire w_dff_B_u8BV5SUB4_0;
	wire w_dff_A_OGLZbC4T0_0;
	wire w_dff_A_fZtf3Zqj6_0;
	wire w_dff_A_Hmu1dZPq4_0;
	wire w_dff_A_2BJdVJ2X9_0;
	wire w_dff_A_FVkfFLj19_0;
	wire w_dff_A_olTvgeWK7_0;
	wire w_dff_A_Dxu63sbT3_0;
	wire w_dff_A_H1MmSlWn2_0;
	wire w_dff_A_u0HMtG4L4_0;
	wire w_dff_A_Yk6WJghu5_0;
	wire w_dff_A_oURrr8Qc5_0;
	wire w_dff_A_5J9vILk98_0;
	wire w_dff_A_aLp7Z5QE0_0;
	wire w_dff_A_5WGFEFAr1_0;
	wire w_dff_B_d36Qvtmv9_1;
	wire w_dff_B_ZdHPZkjT0_1;
	wire w_dff_B_pbjukx3p3_2;
	wire w_dff_B_BnpMevp12_2;
	wire w_dff_B_BgibgsJp5_2;
	wire w_dff_B_FgbljkLo3_2;
	wire w_dff_B_RuJO5MXl4_2;
	wire w_dff_B_aAH60p9E8_2;
	wire w_dff_B_wZ6Naiyz7_2;
	wire w_dff_B_3irCt1cS4_2;
	wire w_dff_B_r2CbHWer7_2;
	wire w_dff_B_FEZZN7fx9_2;
	wire w_dff_B_dOxPNwOr3_2;
	wire w_dff_B_bcl5B0Ji2_2;
	wire w_dff_B_g5nXW3zj7_2;
	wire w_dff_B_LsPfb9yV0_2;
	wire w_dff_B_37eVJ1G91_2;
	wire w_dff_B_JSDHdnHv4_2;
	wire w_dff_B_89sVl6iy5_2;
	wire w_dff_B_7jTaEjpM3_2;
	wire w_dff_B_wrrgvrQ67_2;
	wire w_dff_B_NCl24oB17_2;
	wire w_dff_B_49jATq0G1_2;
	wire w_dff_B_Qq1c6G4n8_2;
	wire w_dff_B_2yg5L7XW3_2;
	wire w_dff_B_afq3mQ3G2_2;
	wire w_dff_B_xPiheAAy0_2;
	wire w_dff_B_eW3s00fe8_2;
	wire w_dff_B_1pw1a6SK8_2;
	wire w_dff_B_8rfYcsID7_2;
	wire w_dff_B_rQvKxmFw5_2;
	wire w_dff_B_famZFcKB5_2;
	wire w_dff_B_tbFlF8UB1_2;
	wire w_dff_B_qMdlOkgv7_2;
	wire w_dff_B_3RX2ORUq0_2;
	wire w_dff_B_mv831Y7I2_2;
	wire w_dff_B_tBPOmc2m2_2;
	wire w_dff_B_OtSpjFUH6_2;
	wire w_dff_B_n30ZIvjc2_2;
	wire w_dff_B_VGVCOS1k9_2;
	wire w_dff_B_JIQOLr3L4_2;
	wire w_dff_B_VjmxtvCP9_2;
	wire w_dff_B_uJsCxzc15_2;
	wire w_dff_B_2wuuOQNM6_2;
	wire w_dff_B_ea6nszm69_2;
	wire w_dff_B_zHSg5EZA8_2;
	wire w_dff_B_5o2CEteu9_2;
	wire w_dff_B_AdjPIj2j3_2;
	wire w_dff_B_1KKQIqhO4_2;
	wire w_dff_B_GuUGSFkC1_2;
	wire w_dff_B_7QK4NaCx4_2;
	wire w_dff_B_LzPIU7lD6_2;
	wire w_dff_B_MAsQbvKE2_2;
	wire w_dff_B_G9WrQf9w3_2;
	wire w_dff_B_EIQDCpFu4_2;
	wire w_dff_B_244B1Wex5_2;
	wire w_dff_B_1FS8p3sa6_2;
	wire w_dff_B_5XV3zr7M5_2;
	wire w_dff_B_U2lBJJDX5_2;
	wire w_dff_B_Bix3zfp38_1;
	wire w_dff_B_HUKiIKo39_1;
	wire w_dff_B_X7tXwIFQ1_1;
	wire w_dff_B_jupwEDHS3_1;
	wire w_dff_B_HxGId1660_1;
	wire w_dff_B_3UXBHJQS2_1;
	wire w_dff_B_Jvmy94ni8_1;
	wire w_dff_B_0sWA1UK89_1;
	wire w_dff_B_0ZwEKrgK9_1;
	wire w_dff_B_11YPltti4_1;
	wire w_dff_B_OSoyy2EH8_1;
	wire w_dff_B_YPELLd6n6_1;
	wire w_dff_B_Qw1tMa5V8_1;
	wire w_dff_B_3lOqtsjK5_0;
	wire w_dff_B_FJJJ8L2U5_0;
	wire w_dff_B_DC7NPE3h0_0;
	wire w_dff_B_yC3cHug76_0;
	wire w_dff_B_RwwjpeXH2_0;
	wire w_dff_B_nc4HFfsQ2_0;
	wire w_dff_B_Qfijb8HS2_0;
	wire w_dff_B_Qc9AZV7I7_0;
	wire w_dff_B_WksdNB8K3_0;
	wire w_dff_B_IjTrR2oE5_0;
	wire w_dff_B_Xfrab0YJ1_0;
	wire w_dff_B_0VGTcHsx1_0;
	wire w_dff_A_pTqzBYu31_1;
	wire w_dff_A_4FePtVCr2_1;
	wire w_dff_A_5F7kZV4w2_1;
	wire w_dff_A_kvi5W9hh3_1;
	wire w_dff_A_OkshN4R91_1;
	wire w_dff_A_yYiUzrlC1_1;
	wire w_dff_A_RMdtxuCP6_1;
	wire w_dff_A_a1q6uYAC1_1;
	wire w_dff_A_WQMxp8Gs8_1;
	wire w_dff_A_7ZYaLpCK1_1;
	wire w_dff_A_bYfNsD6v3_1;
	wire w_dff_A_FhOaXYDI7_1;
	wire w_dff_A_U4LD1zzq3_1;
	wire w_dff_B_8v3WQY2V7_1;
	wire w_dff_B_eKIm7TT43_1;
	wire w_dff_B_qDpLUSQJ5_1;
	wire w_dff_B_SG9rV6eE5_1;
	wire w_dff_B_TDhwSEQc4_1;
	wire w_dff_B_LotP9No29_1;
	wire w_dff_B_WE1PAy2l5_1;
	wire w_dff_B_rLXX39jf1_1;
	wire w_dff_B_sBibyQ3Y8_1;
	wire w_dff_B_GDYGvwbl7_1;
	wire w_dff_B_xhSQ2eNV9_1;
	wire w_dff_B_dMx9PzRk5_1;
	wire w_dff_B_riXXVnAg6_1;
	wire w_dff_B_jNxbnMLI3_0;
	wire w_dff_B_GwVkRXTt3_0;
	wire w_dff_B_MLG8SSbY3_0;
	wire w_dff_B_2jeVg1IQ7_0;
	wire w_dff_B_Jp3TWmxC8_0;
	wire w_dff_B_p58vol1v2_0;
	wire w_dff_B_jerW2Aff7_0;
	wire w_dff_B_15y0Hs482_0;
	wire w_dff_B_PWWwDA3Q3_0;
	wire w_dff_B_ZRk8IG8r4_0;
	wire w_dff_B_zLU5isVA4_0;
	wire w_dff_B_wTDV2G8q2_0;
	wire w_dff_A_pBhS1Xgx7_1;
	wire w_dff_A_kiFRoxr33_1;
	wire w_dff_A_YuBI7OAj3_1;
	wire w_dff_A_FcpZtgMN4_1;
	wire w_dff_A_2y1Mngn19_1;
	wire w_dff_A_OK9QNA8d5_1;
	wire w_dff_A_QgzdG5GI1_1;
	wire w_dff_A_yNYEbi4V6_1;
	wire w_dff_A_M27VZ3eY9_1;
	wire w_dff_A_9xyC4LpG8_1;
	wire w_dff_A_LgJ6lgWz5_1;
	wire w_dff_A_BYSrS0wx7_1;
	wire w_dff_A_X2uFtJnt5_1;
	wire w_dff_B_pFoFlUWE0_1;
	wire w_dff_B_r1PrxLTi4_1;
	wire w_dff_B_BPO2fSng8_1;
	wire w_dff_B_m6704ISZ0_1;
	wire w_dff_B_hiHOPFuQ5_1;
	wire w_dff_B_BzHZeDtJ7_1;
	wire w_dff_B_NbJYKeo75_1;
	wire w_dff_B_bqk360Sm5_1;
	wire w_dff_B_73g31No99_1;
	wire w_dff_B_8EcVF8Sf7_1;
	wire w_dff_B_S398jecD7_1;
	wire w_dff_B_DYBrGr1S5_1;
	wire w_dff_B_LvUM34K53_1;
	wire w_dff_B_SkGD4B6a3_0;
	wire w_dff_B_7WXAFeFZ0_0;
	wire w_dff_B_J5P78yHT3_0;
	wire w_dff_B_qHzjWNrt1_0;
	wire w_dff_B_sIxquQj50_0;
	wire w_dff_B_wgGR5Igf0_0;
	wire w_dff_B_QQZ6U9yX8_0;
	wire w_dff_B_S5Lu6qdr7_0;
	wire w_dff_B_7rWqxsCi8_0;
	wire w_dff_B_w4wAMyPH7_0;
	wire w_dff_B_WOOYhY1H8_0;
	wire w_dff_B_rmZtcw0A2_0;
	wire w_dff_A_uNAV6jyP9_1;
	wire w_dff_A_rsdn4Fvf6_1;
	wire w_dff_A_ec2cygHW9_1;
	wire w_dff_A_wP6v6v4l9_1;
	wire w_dff_A_SKlKZQ3q4_1;
	wire w_dff_A_9RjWiZKk4_1;
	wire w_dff_A_OKriZr6j2_1;
	wire w_dff_A_sSHIpeJ62_1;
	wire w_dff_A_N6W14orn8_1;
	wire w_dff_A_wnKCvNYV1_1;
	wire w_dff_A_qstbFSmp5_1;
	wire w_dff_A_R8FXLjzr9_1;
	wire w_dff_A_vJw6EZhk6_1;
	wire w_dff_B_N9wQQJg86_1;
	wire w_dff_B_SsnF83O28_1;
	wire w_dff_B_KW544CsX5_1;
	wire w_dff_B_TJcVgsp28_1;
	wire w_dff_B_B5jq7bo63_1;
	wire w_dff_B_5bljzWBo5_1;
	wire w_dff_B_76f0BGGX8_1;
	wire w_dff_B_2bpPxMxK3_1;
	wire w_dff_B_fxymJWAO4_1;
	wire w_dff_B_m8Zv5k4W2_1;
	wire w_dff_B_QoVLrXGO4_1;
	wire w_dff_B_y1tpFsAq0_1;
	wire w_dff_B_uDp8zjvm9_1;
	wire w_dff_B_E8Jt4ML90_0;
	wire w_dff_B_XoPospA31_0;
	wire w_dff_B_0alDVRbt3_0;
	wire w_dff_B_hYJZTyWJ0_0;
	wire w_dff_B_786EVvBB0_0;
	wire w_dff_B_4OKTCQay7_0;
	wire w_dff_B_rd3A1EDw4_0;
	wire w_dff_B_Hb7hgK8W9_0;
	wire w_dff_B_f4jijjLA5_0;
	wire w_dff_B_QawrM9Qr4_0;
	wire w_dff_B_eN3dMciJ8_0;
	wire w_dff_B_DXgxM1M27_0;
	wire w_dff_A_hjV3lOHx4_1;
	wire w_dff_A_NDdoCHAe9_1;
	wire w_dff_A_HW0ZDJ4t6_1;
	wire w_dff_A_btICl05A6_1;
	wire w_dff_A_q2F8XsFO5_1;
	wire w_dff_A_kbqibt0p1_1;
	wire w_dff_A_eO1PjrBI2_1;
	wire w_dff_A_czwSC3EB8_1;
	wire w_dff_A_OYzVL8BR8_1;
	wire w_dff_A_rOFx621m8_1;
	wire w_dff_A_u950MIbr0_1;
	wire w_dff_A_mbm2HHbT3_1;
	wire w_dff_A_Sd21jNyI9_1;
	wire w_dff_B_30yM5xKK6_1;
	wire w_dff_B_CGYZkYwP2_1;
	wire w_dff_B_zr07N4Pr6_1;
	wire w_dff_B_6nE8ZbBL8_1;
	wire w_dff_B_LGnK3gLv0_1;
	wire w_dff_B_b31vDNQL9_1;
	wire w_dff_B_weeQiOkW2_1;
	wire w_dff_B_cTuRbi5Y2_1;
	wire w_dff_B_H6VExGyq5_1;
	wire w_dff_B_7cOPp9976_1;
	wire w_dff_B_lvc6ILmI6_1;
	wire w_dff_B_D8PRoUg86_1;
	wire w_dff_B_DNx9ayef5_1;
	wire w_dff_B_0BLcdcqw7_0;
	wire w_dff_B_jQCGwjLa3_0;
	wire w_dff_B_wyZRcVP01_0;
	wire w_dff_B_gV5MsEzD1_0;
	wire w_dff_B_DRUHyAs93_0;
	wire w_dff_B_INf212I59_0;
	wire w_dff_B_rsOKGopn9_0;
	wire w_dff_B_j9P400kM3_0;
	wire w_dff_B_DZNoLCJ52_0;
	wire w_dff_B_ucRAZtgc5_0;
	wire w_dff_B_F08mUVaJ1_0;
	wire w_dff_A_tvreZN8X1_1;
	wire w_dff_A_Cn7XDjv57_1;
	wire w_dff_A_4rZDInLo4_1;
	wire w_dff_A_BAAoP9jH6_1;
	wire w_dff_A_UWVFC1Ic5_1;
	wire w_dff_A_79AkB2Do4_1;
	wire w_dff_A_sOjATV497_1;
	wire w_dff_A_Cat8Zylc3_1;
	wire w_dff_A_lzvz1v0d6_1;
	wire w_dff_A_ZdZNELKh4_1;
	wire w_dff_A_7yapfgYL4_1;
	wire w_dff_A_cIRgkc145_1;
	wire w_dff_B_uWlBIvLo8_1;
	wire w_dff_B_MgA73bY22_1;
	wire w_dff_B_xmXztxwm5_1;
	wire w_dff_B_HlF8PbBy0_1;
	wire w_dff_B_8W7M111H4_1;
	wire w_dff_B_Mdq1B7827_1;
	wire w_dff_B_IwJzkcoX3_1;
	wire w_dff_B_QvlTnmCB9_1;
	wire w_dff_B_2KfT1hEF4_1;
	wire w_dff_B_0cJZaRno9_1;
	wire w_dff_B_oYoAC6kM4_1;
	wire w_dff_B_s5QX8V1B0_1;
	wire w_dff_B_obngi1Mw6_0;
	wire w_dff_B_sZS5H6QN1_0;
	wire w_dff_B_eILZSG073_0;
	wire w_dff_B_7CsJF2TN9_0;
	wire w_dff_B_sIpz9hmA9_0;
	wire w_dff_B_HrfV0fS35_0;
	wire w_dff_B_CkOM9qdK4_0;
	wire w_dff_B_WKxyQKDn9_0;
	wire w_dff_B_Cn15YGIz2_0;
	wire w_dff_B_0kya3YlB7_0;
	wire w_dff_A_PZpdhY025_1;
	wire w_dff_A_2Aeeomrf3_1;
	wire w_dff_A_6ms3FofL1_1;
	wire w_dff_A_MgxkmANA7_1;
	wire w_dff_A_ZnEhY6lB5_1;
	wire w_dff_A_y7GSRsIN9_1;
	wire w_dff_A_0v9Gkyz79_1;
	wire w_dff_A_fxWq5Bfg5_1;
	wire w_dff_A_XVYOy3fL1_1;
	wire w_dff_A_yrIOqe3D5_1;
	wire w_dff_A_TtZdaZ396_1;
	wire w_dff_B_4uJ8Bepp5_1;
	wire w_dff_B_AUzhealC0_1;
	wire w_dff_B_S77Q3T2F2_1;
	wire w_dff_B_a952ppHb0_1;
	wire w_dff_B_PjT0Dn9s2_1;
	wire w_dff_B_ijEFmXS61_1;
	wire w_dff_B_gW7xaS6U3_1;
	wire w_dff_B_O2AeDvK69_1;
	wire w_dff_B_8dCHLFDH7_1;
	wire w_dff_B_YA4uxX2x2_1;
	wire w_dff_B_4vE1JtrY5_0;
	wire w_dff_B_49ivluk90_0;
	wire w_dff_B_75L79S3Z0_0;
	wire w_dff_B_Boao5wH08_0;
	wire w_dff_B_eifM8ikB7_0;
	wire w_dff_B_AeNyD6i78_0;
	wire w_dff_B_57bKYgkk5_0;
	wire w_dff_B_kMbvP8Ys0_0;
	wire w_dff_A_A4IqpdUQ5_1;
	wire w_dff_A_8fL4RIXD2_1;
	wire w_dff_A_eajauNj64_1;
	wire w_dff_A_wspUXdpS9_1;
	wire w_dff_A_myeZBikA5_1;
	wire w_dff_A_v4dCg3kJ4_1;
	wire w_dff_A_1H3sC3Dl2_1;
	wire w_dff_A_eQICZcG63_1;
	wire w_dff_A_UV68AmjS3_1;
	wire w_dff_B_XdGCmkl78_1;
	wire w_dff_B_K8uoeSnC5_1;
	wire w_dff_B_aN7ZBlDt2_1;
	wire w_dff_B_wr3vF4hx2_1;
	wire w_dff_B_Q11UU1Bz4_1;
	wire w_dff_B_PSO2yEQ62_1;
	wire w_dff_B_22LA1uYP2_1;
	wire w_dff_B_tnRGkghO1_1;
	wire w_dff_B_IBPxuKjS9_0;
	wire w_dff_B_qCi3aASs1_0;
	wire w_dff_B_eIQi7tKb4_0;
	wire w_dff_B_bQsmDhh81_0;
	wire w_dff_B_MwJ1wSbg8_0;
	wire w_dff_B_tlSTntkM6_0;
	wire w_dff_A_3JhYv0GU8_1;
	wire w_dff_A_SxywY5UB2_1;
	wire w_dff_A_f48muEoQ5_1;
	wire w_dff_A_XUOQDGnf4_1;
	wire w_dff_A_SD3ES31H9_1;
	wire w_dff_A_aYOi67Ny6_1;
	wire w_dff_A_wCShQUCq8_1;
	wire w_dff_B_Vufxfh1h0_1;
	wire w_dff_B_wkuxKIox2_1;
	wire w_dff_B_24U2AcJ98_1;
	wire w_dff_B_otp3howQ8_1;
	wire w_dff_B_O1mc53Ql2_1;
	wire w_dff_B_yRWGmAue1_1;
	wire w_dff_B_Jum1WBO27_1;
	wire w_dff_B_ZwOkEQIq9_0;
	wire w_dff_B_HqaMKhrT9_0;
	wire w_dff_B_7APDhqe42_0;
	wire w_dff_B_IOOsdPOc2_0;
	wire w_dff_B_BjqKJUgd6_0;
	wire w_dff_A_stdT9izj0_1;
	wire w_dff_A_vDhqPUTt0_1;
	wire w_dff_A_oN0MRBMf9_1;
	wire w_dff_A_6l2COR606_1;
	wire w_dff_A_eoffVhJJ4_1;
	wire w_dff_A_CpR4vvnb3_1;
	wire w_dff_B_DRhGq0Jx3_1;
	wire w_dff_B_f2CfR5yF8_1;
	wire w_dff_B_oWG9Onrk0_1;
	wire w_dff_B_SDVvdd771_1;
	wire w_dff_B_ZJhdyy6G9_1;
	wire w_dff_B_wlGQ1Lsq0_1;
	wire w_dff_B_TgsEjimH4_0;
	wire w_dff_B_qTNqAT652_0;
	wire w_dff_B_4CJJYbYo5_0;
	wire w_dff_B_hVTh9bVH3_0;
	wire w_dff_A_oEnI9cUc0_1;
	wire w_dff_A_ThfkHn2S2_1;
	wire w_dff_A_y6icyVYp4_1;
	wire w_dff_A_95HQoU8P0_1;
	wire w_dff_A_QwUZQSPN3_1;
	wire w_dff_B_JYF0L2XJ8_1;
	wire w_dff_B_510lIA7N8_1;
	wire w_dff_B_jS3TSOxf8_1;
	wire w_dff_A_oxewnWqe5_0;
	wire w_dff_A_d5qDWqJV6_0;
	wire w_dff_B_z5MYaKAx6_1;
	wire w_dff_A_fRkJO1mJ1_0;
	wire w_dff_B_Uj7K2SEj3_1;
	wire w_dff_A_4Ncw3g6H8_1;
	wire w_dff_B_gC9Kk4D31_2;
	wire w_dff_B_kLvZqWp66_1;
	wire w_dff_A_Seyk8gfb3_0;
	wire w_dff_A_1yImg40o4_0;
	wire w_dff_A_ozNheDmb8_0;
	wire w_dff_A_8Oqfx7Y42_0;
	wire w_dff_A_s8vQXMGD9_0;
	wire w_dff_A_L3jATuxM0_0;
	wire w_dff_A_u3AT2OHP4_0;
	wire w_dff_A_MfSNh8Kt5_0;
	wire w_dff_A_1ShWz5oI9_0;
	wire w_dff_A_gzcDSFxN4_0;
	wire w_dff_A_UKl2naQv9_0;
	wire w_dff_A_AmdVlZ4t3_0;
	wire w_dff_A_WYQRrI7A1_0;
	wire w_dff_A_r2uzzCPy2_0;
	wire w_dff_A_OufKW71A1_0;
	wire w_dff_A_PVQkZhej7_0;
	wire w_dff_A_pauUSEtX0_0;
	wire w_dff_A_aN4i3XGp4_0;
	wire w_dff_A_43nPrk3u9_0;
	wire w_dff_A_mK81VH2X9_0;
	wire w_dff_A_6Zg4E4Qp6_0;
	wire w_dff_A_yXbS2Gw17_0;
	wire w_dff_A_mlMGkp182_0;
	wire w_dff_A_58KKJxIu0_0;
	wire w_dff_A_lqpqhx4x1_0;
	wire w_dff_A_ou0a32tw9_0;
	wire w_dff_A_GixbuAfL0_0;
	wire w_dff_A_drcFrAzD4_0;
	wire w_dff_A_f69hM5O12_0;
	wire w_dff_A_NWrmpPhQ9_0;
	wire w_dff_A_65twvrJE0_0;
	wire w_dff_A_4foDo0V27_0;
	wire w_dff_A_VxeqP4YA0_0;
	wire w_dff_A_XU7sFgWb9_0;
	wire w_dff_A_3khLpKQS0_0;
	wire w_dff_A_iXCDGnMZ8_0;
	wire w_dff_A_B1PvtdqP9_0;
	wire w_dff_A_LPCfYOc87_0;
	wire w_dff_A_WCJlgciS9_0;
	wire w_dff_A_PfgyymiN4_0;
	wire w_dff_A_nBHD5X532_0;
	wire w_dff_A_uRpohZrb7_0;
	wire w_dff_A_gsQw3Cox5_0;
	wire w_dff_A_MK0VuhU15_1;
	wire w_dff_B_q0XPWQFi0_1;
	wire w_dff_A_WuTLqNa22_0;
	wire w_dff_A_KfoPNO1Y4_0;
	wire w_dff_A_XSSvmQtG1_0;
	wire w_dff_A_ZlsGnQqO7_0;
	wire w_dff_A_Aa1DoKfs2_0;
	wire w_dff_A_mqjpVsZq5_0;
	wire w_dff_A_5MJeBqd60_0;
	wire w_dff_A_6pmYOGOO3_0;
	wire w_dff_A_ZHU9wbMW3_0;
	wire w_dff_A_Z6vGYTU80_0;
	wire w_dff_A_sOObR9hA0_0;
	wire w_dff_A_0ejioA165_0;
	wire w_dff_A_LffEP1fF1_0;
	wire w_dff_A_Qjav21df6_0;
	wire w_dff_A_xQbIpreV1_0;
	wire w_dff_A_C64Ma2ar9_0;
	wire w_dff_A_fOUgoNZH3_0;
	wire w_dff_A_fskyirpJ7_0;
	wire w_dff_A_N75iOreL9_0;
	wire w_dff_A_UfKbiXcp2_0;
	wire w_dff_A_NAZcYdOt2_0;
	wire w_dff_A_fzlEcLXi8_0;
	wire w_dff_A_xZHh3vOq4_0;
	wire w_dff_A_diknPS3S5_0;
	wire w_dff_A_jVfL5Aub8_0;
	wire w_dff_A_JLn3havl0_0;
	wire w_dff_A_ewHWcpLv0_0;
	wire w_dff_A_pAaIwZXZ5_0;
	wire w_dff_A_xqcYvUh81_0;
	wire w_dff_A_hKojmLny7_0;
	wire w_dff_A_gcK08Eqn0_0;
	wire w_dff_A_MbsevW2o7_0;
	wire w_dff_A_SOwVyMfj0_0;
	wire w_dff_A_sPhTPns42_0;
	wire w_dff_A_dW4RF2Ft7_0;
	wire w_dff_A_ARoe1L8O8_0;
	wire w_dff_A_kXhHpDur1_0;
	wire w_dff_A_YxS1Ph414_0;
	wire w_dff_A_hm4ZlzOA6_0;
	wire w_dff_A_JDpPRqDB1_0;
	wire w_dff_A_7y1XPP7Z4_1;
	wire w_dff_B_g43RiTyq0_1;
	wire w_dff_B_ZxMqnISu0_1;
	wire w_dff_B_Hc8L1sT89_1;
	wire w_dff_B_vrKF4epo2_1;
	wire w_dff_B_8Kww9MzI0_1;
	wire w_dff_B_8x8i6mlF1_1;
	wire w_dff_B_ZjZj9Aby5_1;
	wire w_dff_B_D2oBz4Wa0_1;
	wire w_dff_B_hN8VyDGI1_1;
	wire w_dff_B_DxRVVLY88_1;
	wire w_dff_B_Kn1YLFL86_1;
	wire w_dff_B_eR9WagRX5_1;
	wire w_dff_B_EfijYsn78_1;
	wire w_dff_B_ozXFAZpm0_1;
	wire w_dff_B_84dE1AQn9_1;
	wire w_dff_B_C7Xn6Wbq5_1;
	wire w_dff_B_XF7vc1FB3_1;
	wire w_dff_B_yYPWjdDE5_1;
	wire w_dff_B_5f7EaXK75_1;
	wire w_dff_B_kjvJJgtf9_1;
	wire w_dff_B_taz7nMrq5_1;
	wire w_dff_B_Gie3gtTv3_1;
	wire w_dff_B_DWUFKs3E6_1;
	wire w_dff_B_NKoGWVHk5_1;
	wire w_dff_B_XoeCgNQU5_1;
	wire w_dff_B_mfcqjjRG6_1;
	wire w_dff_B_N1oXcL675_1;
	wire w_dff_B_P73yMuXu2_1;
	wire w_dff_B_4Db8brQB2_1;
	wire w_dff_B_CjtE1QT35_1;
	wire w_dff_B_H7YH7Gy75_1;
	wire w_dff_B_XdewGD5u9_1;
	wire w_dff_B_XEl1n5fU1_1;
	wire w_dff_B_VALSnHhf5_1;
	wire w_dff_B_sdmMjafT8_1;
	wire w_dff_B_Z79BEmHT1_1;
	wire w_dff_B_IwWgFsJp8_1;
	wire w_dff_A_Oa1vXFiX9_0;
	wire w_dff_A_R3bKBnDr9_0;
	wire w_dff_A_ZlLm64wL1_0;
	wire w_dff_A_e4Gtb3Os3_0;
	wire w_dff_A_FN9YtOfB1_0;
	wire w_dff_A_rOPYlOn38_0;
	wire w_dff_A_1WFxNLzI3_0;
	wire w_dff_A_2FslWfwU4_0;
	wire w_dff_A_EtzSNt0L2_0;
	wire w_dff_A_iMLREl8e8_0;
	wire w_dff_A_rxPOp8wx7_0;
	wire w_dff_A_g43Bb1ol8_0;
	wire w_dff_A_ye5rD1Ej7_0;
	wire w_dff_A_HxmDsr3t0_0;
	wire w_dff_A_RbQ6QcXS9_0;
	wire w_dff_A_xFf4yazO4_0;
	wire w_dff_A_Eeg6ZSa59_0;
	wire w_dff_A_R0Y8OcgE7_0;
	wire w_dff_A_iSz0WDy75_0;
	wire w_dff_A_QClbv4NU9_0;
	wire w_dff_A_tjoCZtvS8_0;
	wire w_dff_A_4VcbBO8I7_0;
	wire w_dff_A_6GwuDmAY2_0;
	wire w_dff_A_m0epqztM4_0;
	wire w_dff_A_WWpoYzIe3_0;
	wire w_dff_A_UCCVHBbM7_0;
	wire w_dff_A_Wfq2MU012_0;
	wire w_dff_A_rbpxN1Rn4_0;
	wire w_dff_A_btalWeFR7_0;
	wire w_dff_A_Ii5XlZRL2_0;
	wire w_dff_A_Fes7awqC7_0;
	wire w_dff_A_fMZKtSET8_0;
	wire w_dff_A_0JnkHxpi7_0;
	wire w_dff_A_2hTJTysR2_0;
	wire w_dff_A_y00YJ24C4_0;
	wire w_dff_A_AXw7sj3V1_0;
	wire w_dff_A_kXtpBZXi8_0;
	wire w_dff_A_CSAuEfHm7_1;
	wire w_dff_B_cR2gTOZ97_1;
	wire w_dff_B_54i5Q0MS7_1;
	wire w_dff_B_wtrumuQx4_1;
	wire w_dff_B_6tv5O8MX8_1;
	wire w_dff_B_85mHSmjY2_1;
	wire w_dff_B_olxTzOCY3_1;
	wire w_dff_B_3CPHOMdp8_1;
	wire w_dff_B_QHFoXO5q9_1;
	wire w_dff_B_rB099p4a1_1;
	wire w_dff_B_3aDHaYDp7_1;
	wire w_dff_B_LoZhRq1q7_1;
	wire w_dff_B_yWnOi33b5_1;
	wire w_dff_B_aahxRXEg0_1;
	wire w_dff_B_fz2WoD0H2_1;
	wire w_dff_B_QCOziseq7_1;
	wire w_dff_B_90Tn0qPk1_1;
	wire w_dff_B_2jyAQP1L0_1;
	wire w_dff_B_JEloTsq18_1;
	wire w_dff_B_00823XVm1_1;
	wire w_dff_B_aBqK1NJg7_1;
	wire w_dff_B_V66xwiMO0_1;
	wire w_dff_B_PvkSu1sO1_1;
	wire w_dff_B_bNzryRVm1_1;
	wire w_dff_B_Q3flWllZ2_1;
	wire w_dff_B_ndvr2KGu4_1;
	wire w_dff_B_IiO0KRMc8_1;
	wire w_dff_B_ABYYUiQK7_1;
	wire w_dff_B_TZpxFUax0_1;
	wire w_dff_B_W5ZNOVpY5_1;
	wire w_dff_B_WOYym9X45_1;
	wire w_dff_B_bNIxA3FX7_1;
	wire w_dff_B_4NHOyic36_1;
	wire w_dff_B_XbI8uxyG4_1;
	wire w_dff_B_MJFHgnav4_1;
	wire w_dff_A_p9jKWYMW0_0;
	wire w_dff_A_jsd4sH1j8_0;
	wire w_dff_A_P6ZXIqrC9_0;
	wire w_dff_A_xrVvMFLv8_0;
	wire w_dff_A_NYDw1c584_0;
	wire w_dff_A_dYmh04vC5_0;
	wire w_dff_A_02DZLLnu9_0;
	wire w_dff_A_SNNw2z1M2_0;
	wire w_dff_A_dKJK6svR5_0;
	wire w_dff_A_fOjQaHos0_0;
	wire w_dff_A_uvCSk85k2_0;
	wire w_dff_A_jKvttLj64_0;
	wire w_dff_A_hb2IhXrr6_0;
	wire w_dff_A_PM6uz7Rv9_0;
	wire w_dff_A_bJp0c96x2_0;
	wire w_dff_A_FuGseIGv1_0;
	wire w_dff_A_3QTqhoPC7_0;
	wire w_dff_A_jG9FYM2V2_0;
	wire w_dff_A_3n4B5e6L4_0;
	wire w_dff_A_6frpnqbJ6_0;
	wire w_dff_A_WZh8TLRI9_0;
	wire w_dff_A_iJKnNzY76_0;
	wire w_dff_A_CQiqHLOa7_0;
	wire w_dff_A_56n11hGU8_0;
	wire w_dff_A_zRGzsltV2_0;
	wire w_dff_A_fdUGG1xu6_0;
	wire w_dff_A_ZB7d8JM58_0;
	wire w_dff_A_VoCT5toY1_0;
	wire w_dff_A_DEaZWes05_0;
	wire w_dff_A_d7h3sCZh3_0;
	wire w_dff_A_3yDKZYX31_0;
	wire w_dff_A_n0Z7vuAQ5_0;
	wire w_dff_A_h5FTBKqR0_0;
	wire w_dff_A_8FMft7rY4_0;
	wire w_dff_A_VCBWiqrM6_1;
	wire w_dff_B_VXUxXE5i2_1;
	wire w_dff_B_0NqgOcbr6_1;
	wire w_dff_B_a7UIAezb6_1;
	wire w_dff_B_WoLv6GGD0_1;
	wire w_dff_B_z394AiBi7_1;
	wire w_dff_B_vWoIU1SC6_1;
	wire w_dff_B_2y5u0C9w4_1;
	wire w_dff_B_8Wgyh1953_1;
	wire w_dff_B_JXdJOFc00_1;
	wire w_dff_B_HA7BnoSR1_1;
	wire w_dff_B_vGm4ksid7_1;
	wire w_dff_B_9CEbEvHy7_1;
	wire w_dff_B_0pCRhHbD2_1;
	wire w_dff_B_l1S9vmLL9_1;
	wire w_dff_B_quMxuRZH4_1;
	wire w_dff_B_xpHvWSF86_1;
	wire w_dff_B_xHMh5C4h8_1;
	wire w_dff_B_1IOTEWeh1_1;
	wire w_dff_B_0W4bQnwp0_1;
	wire w_dff_B_6HD1SHxH2_1;
	wire w_dff_B_CEoCruuK5_1;
	wire w_dff_B_wH5rwERM2_1;
	wire w_dff_B_pGf1PXjf4_1;
	wire w_dff_B_VYyTK3eA4_1;
	wire w_dff_B_cZTF5xol6_1;
	wire w_dff_B_4pzDosNZ2_1;
	wire w_dff_B_6EVOQlFo0_1;
	wire w_dff_B_9XwNGk0U2_1;
	wire w_dff_B_eWEe3ipL1_1;
	wire w_dff_B_3mtpIpHT8_1;
	wire w_dff_B_os8dMX4n3_1;
	wire w_dff_A_zojWS9US5_0;
	wire w_dff_A_YAVei9ND7_0;
	wire w_dff_A_5FLD68tZ1_0;
	wire w_dff_A_EzTdPr8q3_0;
	wire w_dff_A_gCIHjZCT1_0;
	wire w_dff_A_Zbd9pH166_0;
	wire w_dff_A_6GruaOuZ0_0;
	wire w_dff_A_GveBnI4F0_0;
	wire w_dff_A_nJUsncYO4_0;
	wire w_dff_A_Emad5PsB9_0;
	wire w_dff_A_pTE7WaHH6_0;
	wire w_dff_A_8asdnRH69_0;
	wire w_dff_A_GVwV9WVe4_0;
	wire w_dff_A_KfDO0agX3_0;
	wire w_dff_A_XuhxZ9mO5_0;
	wire w_dff_A_yK8srXoQ9_0;
	wire w_dff_A_WmY2WDt34_0;
	wire w_dff_A_0K8KwNXu9_0;
	wire w_dff_A_nYsKGQUc6_0;
	wire w_dff_A_9vqx9Qht4_0;
	wire w_dff_A_LOf30NvJ6_0;
	wire w_dff_A_prvmZykS0_0;
	wire w_dff_A_R5x4RGFX9_0;
	wire w_dff_A_qgGvadVp9_0;
	wire w_dff_A_lqobwI2Z9_0;
	wire w_dff_A_LlAoWolS7_0;
	wire w_dff_A_OQDWOHiI4_0;
	wire w_dff_A_pFZ61ev29_0;
	wire w_dff_A_S0iNfoEu0_0;
	wire w_dff_A_TzYCBMEP7_0;
	wire w_dff_A_KESIRdKO2_0;
	wire w_dff_A_lHvD8GlN0_1;
	wire w_dff_B_aSADHQTu3_1;
	wire w_dff_B_3ZdcsKJH9_1;
	wire w_dff_B_ZqWefski7_1;
	wire w_dff_B_hizDrtCA7_1;
	wire w_dff_B_ptBNrwE36_1;
	wire w_dff_B_VwBMDQx89_1;
	wire w_dff_B_8tDafc114_1;
	wire w_dff_B_twfHxHMw7_1;
	wire w_dff_B_a575eMHI3_1;
	wire w_dff_B_swQw10Ym0_1;
	wire w_dff_B_2XznyWvl3_1;
	wire w_dff_B_x7kgNVEF7_1;
	wire w_dff_B_ZCco6TX03_1;
	wire w_dff_B_Vd35OrAI7_1;
	wire w_dff_B_twy1WSuR0_1;
	wire w_dff_B_fFBtw0bh2_1;
	wire w_dff_B_KfambDLf9_1;
	wire w_dff_B_uT46plvO4_1;
	wire w_dff_B_IUZBAAxX6_1;
	wire w_dff_B_8giSlLJ91_1;
	wire w_dff_B_EQX30hvF5_1;
	wire w_dff_B_sBLF6frq1_1;
	wire w_dff_B_bqc2mA7v5_1;
	wire w_dff_B_qIBiK0BQ4_1;
	wire w_dff_B_BYMeohTD0_1;
	wire w_dff_B_NAwfn8bf0_1;
	wire w_dff_B_SB9jIKZE4_1;
	wire w_dff_B_V2FILeAh0_1;
	wire w_dff_A_VuO3Iqgm2_0;
	wire w_dff_A_AtrwzAHS5_0;
	wire w_dff_A_fouVqPd42_0;
	wire w_dff_A_NAIU3vfv8_0;
	wire w_dff_A_vRutJaBF8_0;
	wire w_dff_A_yZEnEJJ37_0;
	wire w_dff_A_nVAERRRU4_0;
	wire w_dff_A_MiKfNUtT0_0;
	wire w_dff_A_lri4jbPY3_0;
	wire w_dff_A_om0DWTBR4_0;
	wire w_dff_A_Cb03oVk69_0;
	wire w_dff_A_TJTBq4iX4_0;
	wire w_dff_A_Dhw3wSJZ4_0;
	wire w_dff_A_4fat33Bv6_0;
	wire w_dff_A_muSacNYn5_0;
	wire w_dff_A_R7n0p3s09_0;
	wire w_dff_A_IaSfGTGT3_0;
	wire w_dff_A_RhBN7Wl41_0;
	wire w_dff_A_QgX6Xu133_0;
	wire w_dff_A_xGh3H45m1_0;
	wire w_dff_A_tcfaNK5u1_0;
	wire w_dff_A_DGJ9JMi79_0;
	wire w_dff_A_ouQ01lMY7_0;
	wire w_dff_A_D0KXoUpF1_0;
	wire w_dff_A_fRLdcCCO6_0;
	wire w_dff_A_qF7n0lNR0_0;
	wire w_dff_A_QAZ1OWo78_0;
	wire w_dff_A_8REIYbrZ2_0;
	wire w_dff_A_DkEdws1O4_1;
	wire w_dff_B_1Hwnia6y5_1;
	wire w_dff_B_7eRMdeHJ6_1;
	wire w_dff_B_XP15YOmj4_1;
	wire w_dff_B_lw6qK0rJ5_1;
	wire w_dff_B_zUPspc0Q0_1;
	wire w_dff_B_Htv7EuUU9_1;
	wire w_dff_B_5b2Rgo8m0_1;
	wire w_dff_B_OkrF5aAh4_1;
	wire w_dff_B_2uVSew0n9_1;
	wire w_dff_B_mJIZdswJ0_1;
	wire w_dff_B_2rXngZl52_1;
	wire w_dff_B_3MwG9N8o0_1;
	wire w_dff_B_iHT480Tn6_1;
	wire w_dff_B_yEywQHVs1_1;
	wire w_dff_B_Rzwsub104_1;
	wire w_dff_B_xRfHIyoQ7_1;
	wire w_dff_B_N5u7Y69e2_1;
	wire w_dff_B_o1Wyqwih8_1;
	wire w_dff_B_0PoCoKpS5_1;
	wire w_dff_B_abBCvjBt5_1;
	wire w_dff_B_zdkpLGdc5_1;
	wire w_dff_B_JoeoQYl15_1;
	wire w_dff_B_ywdPvI0A7_1;
	wire w_dff_B_gBOEeCXE2_1;
	wire w_dff_B_kGQLwCQb2_1;
	wire w_dff_A_lOmWAwmn7_0;
	wire w_dff_A_C8MyfKbz3_0;
	wire w_dff_A_bN5Kgzky8_0;
	wire w_dff_A_6FNsbAd11_0;
	wire w_dff_A_A3eZGUtg0_0;
	wire w_dff_A_60rmtUnQ1_0;
	wire w_dff_A_c4GuJAhG9_0;
	wire w_dff_A_PlPOWuLG1_0;
	wire w_dff_A_si98wfdP8_0;
	wire w_dff_A_kQXNzgLG6_0;
	wire w_dff_A_V6uivRY26_0;
	wire w_dff_A_OcrFrRTl0_0;
	wire w_dff_A_AhyO9wxh9_0;
	wire w_dff_A_0tAqT7jG1_0;
	wire w_dff_A_nAKTEXvw9_0;
	wire w_dff_A_XWLuz7rt9_0;
	wire w_dff_A_jK0aNFSy9_0;
	wire w_dff_A_ynk5SylS1_0;
	wire w_dff_A_koF0IBwu4_0;
	wire w_dff_A_2IZZW4I74_0;
	wire w_dff_A_XaSxk0By8_0;
	wire w_dff_A_pHBec1sl8_0;
	wire w_dff_A_t5WXf41F4_0;
	wire w_dff_A_Blq0YXyK8_0;
	wire w_dff_A_9otDpVqf0_0;
	wire w_dff_A_RVsGh9gK2_1;
	wire w_dff_B_ho3VH9op0_1;
	wire w_dff_B_Fz5biCnP3_1;
	wire w_dff_B_aoBeiQaW0_1;
	wire w_dff_B_zXm3zxue6_1;
	wire w_dff_B_Js4dWb0A8_1;
	wire w_dff_B_XtgDgxAH8_1;
	wire w_dff_B_iFkoXCaA1_1;
	wire w_dff_B_MapPrYeL5_1;
	wire w_dff_B_dYwt28XJ1_1;
	wire w_dff_B_IcoHR6Jl6_1;
	wire w_dff_B_4zcNiNTF9_1;
	wire w_dff_B_ekmokFYU8_1;
	wire w_dff_B_BU0okkuW7_1;
	wire w_dff_B_D2HUPqIi1_1;
	wire w_dff_B_foJYmLVh5_1;
	wire w_dff_B_luqDlp972_1;
	wire w_dff_B_woYQI3Xo1_1;
	wire w_dff_B_DWYYMhFN1_1;
	wire w_dff_B_2KBAuhsx4_1;
	wire w_dff_B_svZT3w2m4_1;
	wire w_dff_B_eZQ8FN4T1_1;
	wire w_dff_B_KXgzlV1M9_1;
	wire w_dff_A_J7WOjswY8_0;
	wire w_dff_A_uL7sbdPp1_0;
	wire w_dff_A_u2OnqcI40_0;
	wire w_dff_A_3HCtycP24_0;
	wire w_dff_A_Asf8COAB8_0;
	wire w_dff_A_d6buk1457_0;
	wire w_dff_A_KHgypmyQ1_0;
	wire w_dff_A_miRXi02Y2_0;
	wire w_dff_A_9uKv9i878_0;
	wire w_dff_A_5gmCLYxM3_0;
	wire w_dff_A_vnXmfF1G1_0;
	wire w_dff_A_zlElvV4I0_0;
	wire w_dff_A_5URrfS203_0;
	wire w_dff_A_e1pVPcMY9_0;
	wire w_dff_A_e9IMCj5g1_0;
	wire w_dff_A_RxNTvOhv2_0;
	wire w_dff_A_GvO1V44g7_0;
	wire w_dff_A_E4SLNtuM0_0;
	wire w_dff_A_cqj1vMHG2_0;
	wire w_dff_A_TWxyknpV1_0;
	wire w_dff_A_N65SNwsB3_0;
	wire w_dff_A_gM2LXppr0_0;
	wire w_dff_A_E2AfKQGi1_1;
	wire w_dff_B_LkzXASl69_1;
	wire w_dff_B_QBY03YW21_1;
	wire w_dff_B_znxiZW4c3_1;
	wire w_dff_B_00jPaK7g9_1;
	wire w_dff_B_r5P06Tk20_1;
	wire w_dff_B_VwUw66dR5_1;
	wire w_dff_B_JVNXc6vS4_1;
	wire w_dff_B_cByGxDKc2_1;
	wire w_dff_B_5ugC1HHl1_1;
	wire w_dff_B_I1qL3ToX2_1;
	wire w_dff_B_cuYa9qI68_1;
	wire w_dff_B_HdWi1d3R2_1;
	wire w_dff_B_f6gA8plr8_1;
	wire w_dff_B_ydGDNvnU7_1;
	wire w_dff_B_Xh79EhiN2_1;
	wire w_dff_B_1YaZ1wIn0_1;
	wire w_dff_B_X3u6fkyO1_1;
	wire w_dff_B_NwoMSljy8_1;
	wire w_dff_B_yHoAoE6P4_1;
	wire w_dff_A_F6HOCl9Z1_0;
	wire w_dff_A_NLMVx5xN4_0;
	wire w_dff_A_SdbbVui39_0;
	wire w_dff_A_ibJZI8Pz8_0;
	wire w_dff_A_NEDW3c189_0;
	wire w_dff_A_DiDbtBgY6_0;
	wire w_dff_A_d9g259gG9_0;
	wire w_dff_A_CVfikeBg8_0;
	wire w_dff_A_nOrqZHBH0_0;
	wire w_dff_A_2b7vdG0w9_0;
	wire w_dff_A_m0njP2kO6_0;
	wire w_dff_A_q0Nn6ixV0_0;
	wire w_dff_A_lMZKy4LX9_0;
	wire w_dff_A_GQIVikUo5_0;
	wire w_dff_A_uVIXtaQe2_0;
	wire w_dff_A_SFM34Hx82_0;
	wire w_dff_A_MgZ8Tsoj1_0;
	wire w_dff_A_uOxkyAHE4_0;
	wire w_dff_A_nXyfF5ZW7_0;
	wire w_dff_A_ujIduFVv2_1;
	wire w_dff_B_uQa7je7J4_1;
	wire w_dff_B_0dXH419U3_1;
	wire w_dff_B_uVc8stqu4_1;
	wire w_dff_B_vTTMyKL42_1;
	wire w_dff_B_IkNeszDg4_1;
	wire w_dff_B_QEH6NRHJ8_1;
	wire w_dff_B_9HLorpzB3_1;
	wire w_dff_B_REtC54pC2_1;
	wire w_dff_B_7Cz5Z4Kr4_1;
	wire w_dff_B_RcFjeqnT6_1;
	wire w_dff_B_VmXVDCV31_1;
	wire w_dff_B_HUFtEnqY0_1;
	wire w_dff_B_HEx40znw5_1;
	wire w_dff_B_NFEyZqW68_1;
	wire w_dff_B_d8EbkTxD8_1;
	wire w_dff_B_4IAinCvK4_1;
	wire w_dff_A_sIr3t28d7_0;
	wire w_dff_A_9iyz4Pte6_0;
	wire w_dff_A_R4Oz2l9q0_0;
	wire w_dff_A_FjSEhMfU8_0;
	wire w_dff_A_j1Xv7zmb2_0;
	wire w_dff_A_L382okfo6_0;
	wire w_dff_A_l9nhwDHr8_0;
	wire w_dff_A_OOlRk1Ny8_0;
	wire w_dff_A_gUhkwX6k5_0;
	wire w_dff_A_938kOzp87_0;
	wire w_dff_A_BeJ7GYUl7_0;
	wire w_dff_A_4YMDY7en1_0;
	wire w_dff_A_rjLEFNFV8_0;
	wire w_dff_A_vUPAaQ5i2_0;
	wire w_dff_A_gs5bTWi95_0;
	wire w_dff_A_3paX2inR4_0;
	wire w_dff_A_2h6ak3GK4_1;
	wire w_dff_B_O1nL2Eme5_1;
	wire w_dff_B_4Dq2Ul1G2_1;
	wire w_dff_B_wXjGVgAc2_1;
	wire w_dff_B_sTcbt0Xc1_1;
	wire w_dff_B_8ludC52q6_1;
	wire w_dff_B_7MFV8VOy2_1;
	wire w_dff_B_b2JeRQLK7_1;
	wire w_dff_B_6qA0x1Dt3_1;
	wire w_dff_B_cgCwIWBN1_1;
	wire w_dff_B_9Ckz7EOK7_1;
	wire w_dff_B_aJJ7xfrT9_1;
	wire w_dff_B_wDNz3IFj5_1;
	wire w_dff_B_e5SXL19y3_1;
	wire w_dff_A_yOPOHtc53_0;
	wire w_dff_A_hBEkpYuJ6_0;
	wire w_dff_A_bUeLdpSR5_0;
	wire w_dff_A_cH1xxg165_0;
	wire w_dff_A_d1p6rDNR2_0;
	wire w_dff_A_DmIQjyM20_0;
	wire w_dff_A_d74gFXDP1_0;
	wire w_dff_A_xTEMoy1Y5_0;
	wire w_dff_A_HnoeuEKP9_0;
	wire w_dff_A_BT1MZ7Sz0_0;
	wire w_dff_A_aHaSUFTv5_0;
	wire w_dff_A_8WGJXl8K4_0;
	wire w_dff_A_9WrAOST24_0;
	wire w_dff_A_RKyRjln93_1;
	wire w_dff_B_l7CIwixh9_1;
	wire w_dff_B_I462lvCz2_1;
	wire w_dff_B_58oxfOiv9_1;
	wire w_dff_B_fSed0ote5_1;
	wire w_dff_B_7ga4towO6_1;
	wire w_dff_B_HHOcYcgn9_1;
	wire w_dff_B_D2ySSSay6_1;
	wire w_dff_B_CsC0BIYR3_1;
	wire w_dff_B_41TCNUGG3_1;
	wire w_dff_B_ZBGSYhqQ2_1;
	wire w_dff_A_I9I1WVz00_0;
	wire w_dff_A_Kwk6TNJB8_0;
	wire w_dff_A_5uHSAbGh7_0;
	wire w_dff_A_adtHeypL6_0;
	wire w_dff_A_Dlr3XBF36_0;
	wire w_dff_A_E1i8Mt5B3_0;
	wire w_dff_A_QAldSDto2_0;
	wire w_dff_A_KPirdrdm9_0;
	wire w_dff_A_QHbmduf29_0;
	wire w_dff_A_qdcJQ49M1_0;
	wire w_dff_A_hivLiakV5_1;
	wire w_dff_B_vznmlZVm5_1;
	wire w_dff_B_1XKIj6og3_1;
	wire w_dff_B_jLPMgnHZ4_1;
	wire w_dff_B_yhm7Gakg5_1;
	wire w_dff_B_8CmJTX035_1;
	wire w_dff_B_gzcghbfG9_1;
	wire w_dff_B_MwfEWbpP9_1;
	wire w_dff_A_DecIt21K5_0;
	wire w_dff_A_a9AaLAWx9_0;
	wire w_dff_A_1c9raQmS9_0;
	wire w_dff_A_gVIRcJBG4_0;
	wire w_dff_A_ioR6XyE70_0;
	wire w_dff_A_o4KfhgMK0_0;
	wire w_dff_A_d8DAIhbV2_0;
	wire w_dff_A_MSEJUAI97_1;
	wire w_dff_B_6M5aIzqv6_1;
	wire w_dff_B_ifezlAmu9_1;
	wire w_dff_B_VxStCGKZ2_1;
	wire w_dff_B_UGGTIAOT5_1;
	wire w_dff_B_DaDNKJQD9_2;
	wire w_dff_A_VvcuaMFH7_0;
	wire w_dff_A_mKL79bUP7_0;
	wire w_dff_A_HiWWr8kQ9_0;
	wire w_dff_A_QnJKV9jW3_0;
	wire w_dff_B_4AVndoHp8_0;
	wire w_dff_A_sICFtYLJ6_0;
	wire w_dff_A_7PsyB8RX7_0;
	wire w_dff_A_g7Cqca0B3_1;
	wire w_dff_B_kUX2dQoU1_1;
	wire w_dff_B_uh08qkyA8_2;
	wire w_dff_B_67SyN4BX0_2;
	wire w_dff_B_3n1TvbgO3_2;
	wire w_dff_B_E23RCO5t0_2;
	wire w_dff_B_kmhO2PBp8_2;
	wire w_dff_B_wpKlsJpS2_2;
	wire w_dff_B_uJhi3PER3_2;
	wire w_dff_B_Rl3aCQEo4_2;
	wire w_dff_B_lXBkLMC50_2;
	wire w_dff_B_rRhLN53z2_2;
	wire w_dff_B_fpVYwdWF7_2;
	wire w_dff_B_D7IdrbQv4_2;
	wire w_dff_B_u9ZhCgMi0_2;
	wire w_dff_B_oceqJu7P4_2;
	wire w_dff_B_JFQ8KwRR2_2;
	wire w_dff_B_jYYsO1in3_2;
	wire w_dff_B_2OWlbafw5_2;
	wire w_dff_B_WcVNyhwX7_2;
	wire w_dff_B_u4pT78iO2_2;
	wire w_dff_B_bjv4PFRx5_2;
	wire w_dff_B_sduVcZIW5_2;
	wire w_dff_B_NGW36fhR9_2;
	wire w_dff_B_r3j6jYjK6_2;
	wire w_dff_B_bBDHLzPL3_2;
	wire w_dff_B_TofsPsMb4_2;
	wire w_dff_B_udEqYqW39_2;
	wire w_dff_B_yGZWIbEw3_2;
	wire w_dff_B_4jdMOdpI9_2;
	wire w_dff_B_i5nC3PJ59_2;
	wire w_dff_B_cpC5Ctxy3_2;
	wire w_dff_B_6uAyAGD86_2;
	wire w_dff_B_Eep8acM41_2;
	wire w_dff_B_HK7RbBR77_2;
	wire w_dff_B_bnjkz5Xs0_2;
	wire w_dff_B_c5oPvu1p9_2;
	wire w_dff_B_ErOjuLIh3_2;
	wire w_dff_B_H4vF8Jzv3_2;
	wire w_dff_B_2dg9xcRF3_2;
	wire w_dff_B_3C3MC2xr3_2;
	wire w_dff_B_xjjOOBCW3_2;
	wire w_dff_B_0HIzmumo0_2;
	wire w_dff_B_YVxJX7bK8_2;
	wire w_dff_B_npU4dBmU0_2;
	wire w_dff_A_4srhdI5f7_0;
	wire w_dff_B_7ZqNEE1X2_1;
	wire w_dff_B_MyRF88Ho1_2;
	wire w_dff_B_vs2i8CRr4_2;
	wire w_dff_B_HxjixdtX4_2;
	wire w_dff_B_2schdg8b4_2;
	wire w_dff_B_X0AEB7865_2;
	wire w_dff_B_wSinLOER6_2;
	wire w_dff_B_ZbenMmdJ3_2;
	wire w_dff_B_w4pjXUgY0_2;
	wire w_dff_B_zixU73o69_2;
	wire w_dff_B_Hg8CQCUM2_2;
	wire w_dff_B_t875ONQ45_2;
	wire w_dff_B_JOVkWgXp1_2;
	wire w_dff_B_P0PgcrjQ4_2;
	wire w_dff_B_oervyHLH9_2;
	wire w_dff_B_JbZSDcwQ1_2;
	wire w_dff_B_yTmfgBJe2_2;
	wire w_dff_B_20aD1xrL6_2;
	wire w_dff_B_Zv2aVvHy0_2;
	wire w_dff_B_2RQgefhu4_2;
	wire w_dff_B_AOMSN1Mt7_2;
	wire w_dff_B_Oj94We1D8_2;
	wire w_dff_B_lA1NGeNw4_2;
	wire w_dff_B_DL1JyQv69_2;
	wire w_dff_B_YpF83VGD4_2;
	wire w_dff_B_sobBcY7u5_2;
	wire w_dff_B_H928jWCT5_2;
	wire w_dff_B_Pdn3zpCf7_2;
	wire w_dff_B_EuvBYWQp7_2;
	wire w_dff_B_88g5pI1W8_2;
	wire w_dff_B_usMhhRpj6_2;
	wire w_dff_B_sKOj6k0h7_2;
	wire w_dff_B_Nf4BGIkL3_2;
	wire w_dff_B_U8VFAW3G6_2;
	wire w_dff_B_6eUkt3ob1_2;
	wire w_dff_B_F96ZW9ZA5_2;
	wire w_dff_B_Yev0Ya1m6_2;
	wire w_dff_B_ofK5VT0q6_2;
	wire w_dff_B_BQyzyyjB3_2;
	wire w_dff_B_nEkoHJJ30_2;
	wire w_dff_B_GjiEG68z4_2;
	wire w_dff_A_pk5fm7722_1;
	wire w_dff_B_mH3YQC8G2_1;
	wire w_dff_B_mi78tRPC4_1;
	wire w_dff_B_CuSZhulK4_1;
	wire w_dff_B_POOwfaAm1_1;
	wire w_dff_B_bUBtQcxz5_1;
	wire w_dff_B_RaTCpOwE7_1;
	wire w_dff_B_79dFNKNP5_1;
	wire w_dff_B_fmMxAAbW0_1;
	wire w_dff_B_OekLfmFc3_1;
	wire w_dff_B_6Zr66Qik3_1;
	wire w_dff_B_9Avhm6r94_1;
	wire w_dff_B_zxje7ffB9_1;
	wire w_dff_B_BBDmSs0x4_1;
	wire w_dff_B_gA4B9JWh8_1;
	wire w_dff_B_uXHsKQAB2_1;
	wire w_dff_B_g3lXLIwq1_1;
	wire w_dff_B_lCZmjHv13_1;
	wire w_dff_B_82cERNsd2_1;
	wire w_dff_B_r8jcfOAp4_1;
	wire w_dff_B_5dn8vxyq0_1;
	wire w_dff_B_eQCeMJtD9_1;
	wire w_dff_B_VBj5hVN94_1;
	wire w_dff_B_yx5b9oMt1_1;
	wire w_dff_B_TP95Tceu1_1;
	wire w_dff_B_NTd7QoBg8_1;
	wire w_dff_B_JpcRq0sr7_1;
	wire w_dff_B_8MWQTBhw6_1;
	wire w_dff_B_ukRNl2yb2_1;
	wire w_dff_B_dXQkpcAo9_1;
	wire w_dff_B_fP1syjHV2_1;
	wire w_dff_B_edtvXeBF9_1;
	wire w_dff_B_ZRecMDAO6_1;
	wire w_dff_B_wazNxPDQ7_1;
	wire w_dff_B_4KHvnmWF6_1;
	wire w_dff_B_ubCutBrC6_1;
	wire w_dff_B_IauIUggA0_1;
	wire w_dff_B_e90BrRBC1_1;
	wire w_dff_A_4cCVeIPs0_0;
	wire w_dff_A_Puj7Y3jZ5_0;
	wire w_dff_A_XM7PygpP9_0;
	wire w_dff_A_7flPWa5f8_0;
	wire w_dff_A_ktjG7CB24_0;
	wire w_dff_A_F4tBUn2w1_0;
	wire w_dff_A_GVQjSI4K8_0;
	wire w_dff_A_9B2KPkSK3_0;
	wire w_dff_A_99fWzCkJ8_0;
	wire w_dff_A_JsBJ9IlF9_0;
	wire w_dff_A_u9Y17Nz70_0;
	wire w_dff_A_zaZuvExN7_0;
	wire w_dff_A_vR9gCxSH4_0;
	wire w_dff_A_o4YK45B50_0;
	wire w_dff_A_vC464gJA6_0;
	wire w_dff_A_SzwDyVug4_0;
	wire w_dff_A_nsS9aEr48_0;
	wire w_dff_A_Zt5QNNE91_0;
	wire w_dff_A_qhJqJTnu3_0;
	wire w_dff_A_m0dD5oNw2_0;
	wire w_dff_A_OUkrUA4s7_0;
	wire w_dff_A_7hkTAzJD5_0;
	wire w_dff_A_NDMZ93ru7_0;
	wire w_dff_A_fnpmKFz18_0;
	wire w_dff_A_dXcqFxTP9_0;
	wire w_dff_A_OFTxbFi85_0;
	wire w_dff_A_rFHXN8Fe6_0;
	wire w_dff_A_y4KpsBnx8_0;
	wire w_dff_A_ex8Vjarn0_0;
	wire w_dff_A_m8PoQSv38_0;
	wire w_dff_A_jp9BR9eU5_0;
	wire w_dff_A_Y5rzik6T1_0;
	wire w_dff_A_EZ16Ww6f0_0;
	wire w_dff_A_UThHCoHP4_0;
	wire w_dff_A_ICtdikRJ5_0;
	wire w_dff_A_SfWTCEAE1_0;
	wire w_dff_A_MZQj5o8y5_0;
	wire w_dff_A_ZPHxKH3L7_0;
	wire w_dff_B_TcMWfGUl2_1;
	wire w_dff_A_yep8Mkb95_0;
	wire w_dff_A_Ml3cU1p46_0;
	wire w_dff_A_cUhWZDR51_0;
	wire w_dff_A_VsJ9vFWg0_0;
	wire w_dff_A_kdsM8Nuk2_0;
	wire w_dff_A_m5FNblAF6_0;
	wire w_dff_A_8o5GQI4n3_0;
	wire w_dff_A_vZQmsyke1_0;
	wire w_dff_A_xqneDfm06_0;
	wire w_dff_A_zqb877gu3_0;
	wire w_dff_A_yZD8demx9_0;
	wire w_dff_A_hfNXxVHy4_0;
	wire w_dff_A_OcUc42Uf2_0;
	wire w_dff_A_nE2Pm5Zp5_0;
	wire w_dff_A_b4DvnkBd7_0;
	wire w_dff_A_Gq0Zcrfz6_0;
	wire w_dff_A_TdTx8Vid6_0;
	wire w_dff_A_by2xzjeB0_0;
	wire w_dff_A_6ePQ0IMP4_0;
	wire w_dff_A_TezrQHhD4_0;
	wire w_dff_A_YYTYTgYW8_0;
	wire w_dff_A_hlOgDtrn2_0;
	wire w_dff_A_RgcRg5WZ4_0;
	wire w_dff_A_srhpZvbs1_0;
	wire w_dff_A_8pZMFplZ5_0;
	wire w_dff_A_dVLxC8g57_0;
	wire w_dff_A_UFUxdAPV2_0;
	wire w_dff_A_09L0zUaT4_0;
	wire w_dff_A_gDRNrXgf6_0;
	wire w_dff_A_18hIphsv7_0;
	wire w_dff_A_XCvrLZwF6_0;
	wire w_dff_A_jYUIfQ6Y2_0;
	wire w_dff_A_SmcgCxUj2_0;
	wire w_dff_A_KIQ1Xrxm6_0;
	wire w_dff_A_D4J8BljM6_0;
	wire w_dff_B_3ol2YPqu2_1;
	wire w_dff_A_i1JM5dwV8_0;
	wire w_dff_A_WOZggPKq5_0;
	wire w_dff_A_6GtOBhRn8_0;
	wire w_dff_A_noy1VxbO8_0;
	wire w_dff_A_qsasqbgO9_0;
	wire w_dff_A_5tDBfrqP1_0;
	wire w_dff_A_q0O0cgm53_0;
	wire w_dff_A_Va48axrL4_0;
	wire w_dff_A_qtWnJQZR8_0;
	wire w_dff_A_WTKJSQpe7_0;
	wire w_dff_A_1Wb5c5Hi8_0;
	wire w_dff_A_G061ckVS1_0;
	wire w_dff_A_hqnuUQHr9_0;
	wire w_dff_A_Tt1tlz4D8_0;
	wire w_dff_A_shqwgRBP3_0;
	wire w_dff_A_LboxpIG64_0;
	wire w_dff_A_2Ks4Js8K2_0;
	wire w_dff_A_TArPpHmr3_0;
	wire w_dff_A_Jqtgd0Un3_0;
	wire w_dff_A_XTw8XSQ82_0;
	wire w_dff_A_q59joT0v6_0;
	wire w_dff_A_H0QPgv0Z4_0;
	wire w_dff_A_ggsxK3ad0_0;
	wire w_dff_A_JvHzqgkK6_0;
	wire w_dff_A_3hDHtTTp4_0;
	wire w_dff_A_Vh4Xs31y1_0;
	wire w_dff_A_s5ABN5T91_0;
	wire w_dff_A_I83dDIWl2_0;
	wire w_dff_A_yBAJ2YQw2_0;
	wire w_dff_A_BQ4RT4cZ8_0;
	wire w_dff_A_QnXpZbch3_0;
	wire w_dff_A_YThLcJGt7_0;
	wire w_dff_B_Wx8gVA3f4_1;
	wire w_dff_A_Dp6pYkgg5_0;
	wire w_dff_A_kLiuxRIq5_0;
	wire w_dff_A_k9SGnOS40_0;
	wire w_dff_A_UxINHyAF6_0;
	wire w_dff_A_yX94VMgY2_0;
	wire w_dff_A_LZASZojU4_0;
	wire w_dff_A_WUL0oOaN2_0;
	wire w_dff_A_OQt0ht2d9_0;
	wire w_dff_A_Qn2YoWTQ8_0;
	wire w_dff_A_wQsDb4ik3_0;
	wire w_dff_A_qorG1gqc8_0;
	wire w_dff_A_RjXcQ55b2_0;
	wire w_dff_A_54zR3vse1_0;
	wire w_dff_A_AkOGVlTY6_0;
	wire w_dff_A_sHm8lLFr8_0;
	wire w_dff_A_6zqJZpsy7_0;
	wire w_dff_A_86V7Tos08_0;
	wire w_dff_A_9jgUymra0_0;
	wire w_dff_A_43oKsjpy8_0;
	wire w_dff_A_oOjK5N8O8_0;
	wire w_dff_A_Q1KcbHFn1_0;
	wire w_dff_A_kibVlbmf0_0;
	wire w_dff_A_6KfgduoD1_0;
	wire w_dff_A_uvKssEkd3_0;
	wire w_dff_A_6hOg0Fg01_0;
	wire w_dff_A_TR5dnRrm7_0;
	wire w_dff_A_xzNnXzgm5_0;
	wire w_dff_A_yRb039tD0_0;
	wire w_dff_A_TVcECwO33_0;
	wire w_dff_B_4nstmJjP9_1;
	wire w_dff_A_GMKIGBu49_0;
	wire w_dff_A_BfaZkGg15_0;
	wire w_dff_A_rVzu2cTz0_0;
	wire w_dff_A_rIusyq2v3_0;
	wire w_dff_A_JXQFsXgi1_0;
	wire w_dff_A_0I8RhK9w5_0;
	wire w_dff_A_OkX2pUTe8_0;
	wire w_dff_A_26MB3cam6_0;
	wire w_dff_A_jkixgHNI8_0;
	wire w_dff_A_dPIAWrUa4_0;
	wire w_dff_A_nJvHBlKN9_0;
	wire w_dff_A_HkOiRcYj8_0;
	wire w_dff_A_TvJWAPnU4_0;
	wire w_dff_A_p2u4AGtI7_0;
	wire w_dff_A_qIVvVm9z7_0;
	wire w_dff_A_tKAoNEmu9_0;
	wire w_dff_A_qpmAS6uv8_0;
	wire w_dff_A_Zu5gOBWU7_0;
	wire w_dff_A_7u2lWCTo1_0;
	wire w_dff_A_Tlfzrtja8_0;
	wire w_dff_A_KULErXji4_0;
	wire w_dff_A_ZjU4JL573_0;
	wire w_dff_A_sEM64owF5_0;
	wire w_dff_A_v6J7VqWj2_0;
	wire w_dff_A_b6WhIoFW7_0;
	wire w_dff_A_ssjJfwfn8_0;
	wire w_dff_B_mGfMoIar4_1;
	wire w_dff_A_TVF0ZkmO6_0;
	wire w_dff_A_WLXBINEZ5_0;
	wire w_dff_A_KZakzYWl0_0;
	wire w_dff_A_U4637zoq2_0;
	wire w_dff_A_kzE1S2iG5_0;
	wire w_dff_A_XNmO402k2_0;
	wire w_dff_A_xst5G28g4_0;
	wire w_dff_A_4RW4rLWP5_0;
	wire w_dff_A_FaRc3B7l3_0;
	wire w_dff_A_XPKGPep44_0;
	wire w_dff_A_kIObjICQ4_0;
	wire w_dff_A_siITKYo55_0;
	wire w_dff_A_lbGDJ6Dz9_0;
	wire w_dff_A_dNwyM5om1_0;
	wire w_dff_A_ro56wlhL7_0;
	wire w_dff_A_nUlHRz308_0;
	wire w_dff_A_hXXeUypV3_0;
	wire w_dff_A_fYfhTmPz2_0;
	wire w_dff_A_581ICQAM8_0;
	wire w_dff_A_CxufCeoR3_0;
	wire w_dff_A_t8Y7zL9k1_0;
	wire w_dff_A_6pazhalA8_0;
	wire w_dff_A_GwuSQdzy9_0;
	wire w_dff_B_GGzwUl4x8_1;
	wire w_dff_A_DmmuvWkU1_0;
	wire w_dff_A_hKOdt0Qq9_0;
	wire w_dff_A_a27edCMS9_0;
	wire w_dff_A_GJuj7Haa8_0;
	wire w_dff_A_vwBnq14B0_0;
	wire w_dff_A_G4vo3dq36_0;
	wire w_dff_A_Yyua2LYt9_0;
	wire w_dff_A_QNaXWpn77_0;
	wire w_dff_A_uW9KqhCg7_0;
	wire w_dff_A_MdginEWG5_0;
	wire w_dff_A_APVKPNtx4_0;
	wire w_dff_A_sE3bSTJf9_0;
	wire w_dff_A_eReiMeQq5_0;
	wire w_dff_A_gpito29p2_0;
	wire w_dff_A_4n0Etl6P1_0;
	wire w_dff_A_RJJcbE8U5_0;
	wire w_dff_A_CafySYUU0_0;
	wire w_dff_A_qgPtQnLD1_0;
	wire w_dff_A_8jxZBe6x3_0;
	wire w_dff_A_Fuhz5ZBN3_0;
	wire w_dff_B_Q4fCHPlP0_1;
	wire w_dff_A_XZpB9fif1_0;
	wire w_dff_A_yKxOAacz9_0;
	wire w_dff_A_N0GyQVKT9_0;
	wire w_dff_A_Xasm4Db38_0;
	wire w_dff_A_pJasGj7f2_0;
	wire w_dff_A_X31MRqSb3_0;
	wire w_dff_A_FihyutwB7_0;
	wire w_dff_A_qpSdDf7k8_0;
	wire w_dff_A_PgChPnc70_0;
	wire w_dff_A_AjcRSVMr6_0;
	wire w_dff_A_IWZFFSnZ2_0;
	wire w_dff_A_E2i69n038_0;
	wire w_dff_A_Ylc8IzWN7_0;
	wire w_dff_A_mPMefKtX8_0;
	wire w_dff_A_YTZMBscv6_0;
	wire w_dff_A_XSkiOj6b1_0;
	wire w_dff_A_ZTA4c5vr1_0;
	wire w_dff_B_Ij7RFoTe0_1;
	wire w_dff_A_54yzyJ4a4_0;
	wire w_dff_A_Lj13HK1f7_0;
	wire w_dff_A_OAC4kflL1_0;
	wire w_dff_A_aVS7udP02_0;
	wire w_dff_A_QTcRTf0u6_0;
	wire w_dff_A_jNqAMyIU6_0;
	wire w_dff_A_j7fXsmhR1_0;
	wire w_dff_A_uSIBpSpI9_0;
	wire w_dff_A_j73k00YD8_0;
	wire w_dff_A_gxnswvGT5_0;
	wire w_dff_A_hc74l10N9_0;
	wire w_dff_A_UIFjVK8s3_0;
	wire w_dff_A_rnaNxX3p0_0;
	wire w_dff_A_l1YxZAyV9_0;
	wire w_dff_B_aBtWMcoy6_1;
	wire w_dff_A_sXPX3wjW9_0;
	wire w_dff_A_UQmalzHI7_0;
	wire w_dff_A_l6yAl2QV8_0;
	wire w_dff_A_UXk6t5Dm4_0;
	wire w_dff_A_svhuoTIV4_0;
	wire w_dff_A_qzcvBLxm7_0;
	wire w_dff_A_urmjdxk04_0;
	wire w_dff_A_wnkYSCaX8_0;
	wire w_dff_A_35krV8GY5_0;
	wire w_dff_A_qETlHZLX2_0;
	wire w_dff_A_dgaDtayp4_0;
	wire w_dff_B_DPmtQp9y6_1;
	wire w_dff_A_dWN7is6d5_0;
	wire w_dff_A_QjWMs8ti8_0;
	wire w_dff_A_TD3fKKkG5_0;
	wire w_dff_A_DCJyXSFZ2_0;
	wire w_dff_A_b8ajZ0vy2_0;
	wire w_dff_A_V0PunVvf7_0;
	wire w_dff_A_sLao2UcO5_0;
	wire w_dff_A_iQhZsTBv4_0;
	wire w_dff_B_665wR8I06_1;
	wire w_dff_A_uNlohcFg2_0;
	wire w_dff_A_GbQgXPnf5_0;
	wire w_dff_A_UEeEy5Yb0_0;
	wire w_dff_A_ekScY5O94_0;
	wire w_dff_B_lUl1Ec815_0;
	wire w_dff_A_Xm4Ois8X2_0;
	wire w_dff_A_MTFXj9jv8_0;
	wire w_dff_B_TE7IUzHw6_2;
	wire w_dff_B_m2D92t4A6_2;
	wire w_dff_B_KvJmMPCZ2_2;
	wire w_dff_B_TUmgFBeP4_2;
	wire w_dff_B_zfbUrtA34_2;
	wire w_dff_B_RJeRf19S1_2;
	wire w_dff_B_y99PNr7M2_2;
	wire w_dff_B_NdhpUcr03_2;
	wire w_dff_B_Ofo8b89l6_2;
	wire w_dff_B_TzIJma0E4_2;
	wire w_dff_B_TPKlGYzw5_2;
	wire w_dff_B_YeQLhzxq8_2;
	wire w_dff_B_jcEzTYw38_2;
	wire w_dff_B_5GsClUeS8_2;
	wire w_dff_B_wNpxeUlw1_2;
	wire w_dff_B_5mnpL7rk9_2;
	wire w_dff_B_iLMfAYs48_2;
	wire w_dff_B_6JYjTF0m1_2;
	wire w_dff_B_GiFFH6du6_2;
	wire w_dff_B_xaPCS9GA0_2;
	wire w_dff_B_QupNyiK51_2;
	wire w_dff_B_zfECBIgh9_2;
	wire w_dff_B_tZqpdtqD4_2;
	wire w_dff_B_cb9E4iQu3_2;
	wire w_dff_B_lIxqaB019_2;
	wire w_dff_B_rebp5DpQ9_2;
	wire w_dff_B_qockIgX34_2;
	wire w_dff_B_H1ZRfpr80_2;
	wire w_dff_B_L9MWqCdD2_2;
	wire w_dff_B_MwCkCbO47_2;
	wire w_dff_B_Tnvf8DVQ3_2;
	wire w_dff_B_RDWDIazy7_2;
	wire w_dff_B_ulTm7mSm4_2;
	wire w_dff_B_7oVIdcJM4_2;
	wire w_dff_B_3dgdwS6e4_2;
	wire w_dff_B_McpLEPzu8_2;
	wire w_dff_B_IcRXRP7O7_2;
	wire w_dff_B_K7d4hIjO0_2;
	wire w_dff_B_GK5aTa5s1_2;
	wire w_dff_B_OfZUHjtI3_2;
	wire w_dff_B_MJKSD1ir7_2;
	wire w_dff_B_omBAHzXb1_2;
	wire w_dff_B_cvsacRiZ6_2;
	wire w_dff_B_5NNsqtcs0_2;
	wire w_dff_A_jtq9VIji0_0;
	wire w_dff_B_L4bM11W03_1;
	wire w_dff_B_NXpybWVb0_2;
	wire w_dff_B_SNfaZxqY4_2;
	wire w_dff_B_unmECFzh3_2;
	wire w_dff_B_lzeeD1D73_2;
	wire w_dff_B_pV981ygm7_2;
	wire w_dff_B_US0csvFV5_2;
	wire w_dff_B_gjQBVSZT0_2;
	wire w_dff_B_7XS5vAmo3_2;
	wire w_dff_B_y7jSaYIm2_2;
	wire w_dff_B_7X16aKI65_2;
	wire w_dff_B_dYzLpyIv9_2;
	wire w_dff_B_DEqnNIst6_2;
	wire w_dff_B_ttTgWAgs7_2;
	wire w_dff_B_aQr5yUPV7_2;
	wire w_dff_B_tkqZrdFq3_2;
	wire w_dff_B_UtvbkyQV0_2;
	wire w_dff_B_YYmzVbct7_2;
	wire w_dff_B_yg1oDqeG3_2;
	wire w_dff_B_QN6STyxv3_2;
	wire w_dff_B_saMXTMqk2_2;
	wire w_dff_B_qO0D7mff5_2;
	wire w_dff_B_aNSdxiyd0_2;
	wire w_dff_B_uM4KoRwI5_2;
	wire w_dff_B_eutStpg04_2;
	wire w_dff_B_Fpge5zU09_2;
	wire w_dff_B_UDRrIOuF2_2;
	wire w_dff_B_2M7o3Xm55_2;
	wire w_dff_B_NMt9eYEZ2_2;
	wire w_dff_B_M8PEl6yE4_2;
	wire w_dff_B_F8UOjfwp2_2;
	wire w_dff_B_BF8davyZ9_2;
	wire w_dff_B_nH9dYGtR9_2;
	wire w_dff_B_sVIqy5wP8_2;
	wire w_dff_B_Magq2tLW1_2;
	wire w_dff_B_42odInzz4_2;
	wire w_dff_B_5JqZnrUw2_2;
	wire w_dff_B_ySZqLxuy4_2;
	wire w_dff_B_E5urkzbu4_2;
	wire w_dff_B_Gp3sfWDO7_2;
	wire w_dff_B_GiPGGvU81_2;
	wire w_dff_A_hYbFF23a1_1;
	wire w_dff_A_UvLQDDSv5_0;
	wire w_dff_A_kstmPLp70_0;
	wire w_dff_A_wFyE6uTZ6_0;
	wire w_dff_A_nSRMrK0O5_0;
	wire w_dff_A_MC0Qs3eK4_0;
	wire w_dff_A_Bnu8nZuB0_0;
	wire w_dff_A_ljA7cAPy1_0;
	wire w_dff_A_vFuPo2Il1_0;
	wire w_dff_A_RlpAuLPe3_0;
	wire w_dff_A_nXICAeIO3_0;
	wire w_dff_A_BdIuxJW48_0;
	wire w_dff_A_iIRk5VLh5_0;
	wire w_dff_A_ezUAFxHZ1_0;
	wire w_dff_A_PeIArAzX7_0;
	wire w_dff_A_1zWLdJ3N7_0;
	wire w_dff_A_kB0tQKH79_0;
	wire w_dff_A_73wH3RgH5_0;
	wire w_dff_A_twPON9eS6_0;
	wire w_dff_A_9O3gJxRv3_0;
	wire w_dff_A_7lk4NUJ14_0;
	wire w_dff_A_HKw6jIgO9_0;
	wire w_dff_A_U2qgJ6413_0;
	wire w_dff_A_VQsAhFVy1_0;
	wire w_dff_A_XdrIhCRw8_0;
	wire w_dff_A_HEXadBW79_0;
	wire w_dff_A_3PsCWxAH3_0;
	wire w_dff_A_KEHKnKex5_0;
	wire w_dff_A_iodJtMTu7_0;
	wire w_dff_A_FWLtlRdZ9_0;
	wire w_dff_A_oQaM2Mvm7_0;
	wire w_dff_A_v3G458jc4_0;
	wire w_dff_A_mFXfWBcB2_0;
	wire w_dff_A_ZB7ACmPt8_0;
	wire w_dff_A_LcHzCn9O8_0;
	wire w_dff_A_kOMYAdAY8_0;
	wire w_dff_A_H8PJtw943_0;
	wire w_dff_A_B8itLeCq2_0;
	wire w_dff_A_Pt0afR317_1;
	wire w_dff_A_0aocDaWj8_2;
	wire w_dff_B_dNQi9PLH0_1;
	wire w_dff_B_P5kqbM7h2_2;
	wire w_dff_B_PPyj4RN67_2;
	wire w_dff_B_FTZvdhQU1_2;
	wire w_dff_B_I5b0sp8H6_2;
	wire w_dff_B_ihd7apOB8_2;
	wire w_dff_B_iNmPesNL5_2;
	wire w_dff_B_idfNLey56_2;
	wire w_dff_B_Eyv94Qvs4_2;
	wire w_dff_B_OMl5hO618_2;
	wire w_dff_B_QO7kxPFe6_2;
	wire w_dff_B_vT1oA9iS5_2;
	wire w_dff_B_raYfew9D8_2;
	wire w_dff_B_tOGUTWXH3_2;
	wire w_dff_B_p2kaPQWR6_2;
	wire w_dff_B_UoFZvXiB8_2;
	wire w_dff_B_zT0Yk9Hi4_2;
	wire w_dff_B_rNqmNcCx6_2;
	wire w_dff_B_lv1SRQXi1_2;
	wire w_dff_B_MdZkpYz10_2;
	wire w_dff_B_bZRHx9if7_2;
	wire w_dff_B_PY2wD7eq7_2;
	wire w_dff_B_b8D34B625_2;
	wire w_dff_B_fAxKGH039_2;
	wire w_dff_B_3n01StlD6_2;
	wire w_dff_B_8AXscg2M5_2;
	wire w_dff_B_stLbKPUz1_2;
	wire w_dff_B_4JcNNLnI1_2;
	wire w_dff_B_KcbvCYKb7_2;
	wire w_dff_B_A5OQRGhH1_2;
	wire w_dff_B_E1rZKPON0_2;
	wire w_dff_B_ErlpDTqi1_2;
	wire w_dff_B_NJuq3n8J9_2;
	wire w_dff_B_LMMTeiyX9_2;
	wire w_dff_B_ah10LIvS1_2;
	wire w_dff_B_Dlogfoix6_1;
	wire w_dff_B_I5qByQ2b0_2;
	wire w_dff_B_AM9CuuDy7_2;
	wire w_dff_B_Ltm5NdKr8_2;
	wire w_dff_B_F5yvn08P8_2;
	wire w_dff_B_2v9bMgNf8_2;
	wire w_dff_B_7wzU8vK20_2;
	wire w_dff_B_tb8bruCo5_2;
	wire w_dff_B_VS5c4Ex44_2;
	wire w_dff_B_gPlquzEW3_2;
	wire w_dff_B_kBc74Hlf1_2;
	wire w_dff_B_9hlGbQcB1_2;
	wire w_dff_B_JKc2WJVm2_2;
	wire w_dff_B_DMgHGdz74_2;
	wire w_dff_B_GjsClQzy5_2;
	wire w_dff_B_Y6EvD0z66_2;
	wire w_dff_B_MOibOGLg5_2;
	wire w_dff_B_Tp1Yx1iJ6_2;
	wire w_dff_B_5susflEF9_2;
	wire w_dff_B_p2w1ZfdA3_2;
	wire w_dff_B_hycbdnRu4_2;
	wire w_dff_B_0qEocB764_2;
	wire w_dff_B_E1EsZ7Zp7_2;
	wire w_dff_B_fTpHpzeg2_2;
	wire w_dff_B_S4CnyiCq6_2;
	wire w_dff_B_vZTI7Q4v9_2;
	wire w_dff_B_PYZxaz5r4_2;
	wire w_dff_B_Oazy7wZj8_2;
	wire w_dff_B_Xg8h8zKW0_2;
	wire w_dff_B_KwQq9Pvw0_2;
	wire w_dff_B_uCo2WFDQ7_2;
	wire w_dff_B_BpsdmnhP5_2;
	wire w_dff_B_VlAwclpH3_1;
	wire w_dff_B_frsO1YE89_2;
	wire w_dff_B_q2OIXh6o9_2;
	wire w_dff_B_AOPQ8Cgv5_2;
	wire w_dff_B_3tgNZQ2M5_2;
	wire w_dff_B_3tOvUodx0_2;
	wire w_dff_B_Qf7Ol6hQ5_2;
	wire w_dff_B_gvOhazXT0_2;
	wire w_dff_B_VHcLtPYa1_2;
	wire w_dff_B_KjcNmx9n4_2;
	wire w_dff_B_OdAHMk085_2;
	wire w_dff_B_M08TkCT50_2;
	wire w_dff_B_KudcsrTK9_2;
	wire w_dff_B_oYaIClRT9_2;
	wire w_dff_B_0yQqW5rK6_2;
	wire w_dff_B_4NfDJ9Do6_2;
	wire w_dff_B_21AlTdPx9_2;
	wire w_dff_B_9R50SdT34_2;
	wire w_dff_B_fNBn6mQi5_2;
	wire w_dff_B_eyd7J8PN4_2;
	wire w_dff_B_mQ9i8Y283_2;
	wire w_dff_B_Pe5S1Bua7_2;
	wire w_dff_B_8GmyEVhh7_2;
	wire w_dff_B_KzNRgZlN9_2;
	wire w_dff_B_debyNz7m6_2;
	wire w_dff_B_71sD4LkC3_2;
	wire w_dff_B_OKLa9Y4w5_2;
	wire w_dff_B_vAR6gnbU2_2;
	wire w_dff_B_SQ2UFCHO7_2;
	wire w_dff_B_L2nPKQmm2_1;
	wire w_dff_B_c4sq8zqR5_2;
	wire w_dff_B_mOoYf1Jb9_2;
	wire w_dff_B_yCZhBPxp8_2;
	wire w_dff_B_Mul37upJ9_2;
	wire w_dff_B_Vr2Pzmrc5_2;
	wire w_dff_B_qo8HQgrj5_2;
	wire w_dff_B_K3DD2AXb5_2;
	wire w_dff_B_HZkZjAfV5_2;
	wire w_dff_B_FH92ztJZ4_2;
	wire w_dff_B_w8i5aEmS3_2;
	wire w_dff_B_cjp2gP3k2_2;
	wire w_dff_B_Z5u0LZ2M7_2;
	wire w_dff_B_XiHaLHLS6_2;
	wire w_dff_B_IXsfg1ad6_2;
	wire w_dff_B_WaX5XqFb4_2;
	wire w_dff_B_7Ze0OYxt3_2;
	wire w_dff_B_WTlshVem5_2;
	wire w_dff_B_d9wXloB33_2;
	wire w_dff_B_RSoPvPgy5_2;
	wire w_dff_B_Xya5hZUY2_2;
	wire w_dff_B_zqATVwVs3_2;
	wire w_dff_B_Xi5AxfYo5_2;
	wire w_dff_B_8Nz5cBEq1_2;
	wire w_dff_B_qarWrr7Y9_2;
	wire w_dff_B_4CbSZ5vX4_2;
	wire w_dff_B_X5omvm2U0_1;
	wire w_dff_B_FL4oPBb72_2;
	wire w_dff_B_LvPyXXkq7_2;
	wire w_dff_B_2bilZ0N25_2;
	wire w_dff_B_ENdoiEJq4_2;
	wire w_dff_B_vese2wvk4_2;
	wire w_dff_B_WM4BWJ4s8_2;
	wire w_dff_B_jNlVsGzh4_2;
	wire w_dff_B_q0eth2wE1_2;
	wire w_dff_B_WG9DLVO93_2;
	wire w_dff_B_FP48xxx35_2;
	wire w_dff_B_WcOaV3KZ7_2;
	wire w_dff_B_u5k8TSn71_2;
	wire w_dff_B_c4e9w2VA4_2;
	wire w_dff_B_jXUeBYB18_2;
	wire w_dff_B_hjc6npKu3_2;
	wire w_dff_B_TfLbHHsW6_2;
	wire w_dff_B_r5XncUOe1_2;
	wire w_dff_B_byJXfhuc8_2;
	wire w_dff_B_j3iwvC752_2;
	wire w_dff_B_JfxA9DbI9_2;
	wire w_dff_B_ym3Zhri70_2;
	wire w_dff_B_zx4XBNOA8_2;
	wire w_dff_B_Bs4DgqRc7_1;
	wire w_dff_B_eVoHHgMh1_2;
	wire w_dff_B_ifv1llP13_2;
	wire w_dff_B_pncGDIyb2_2;
	wire w_dff_B_dpQYugbH5_2;
	wire w_dff_B_sv95vB819_2;
	wire w_dff_B_u2QHBXNp3_2;
	wire w_dff_B_6xU8DAjM9_2;
	wire w_dff_B_rVOc4Pvu7_2;
	wire w_dff_B_Y867QQsv3_2;
	wire w_dff_B_IABYL4ue1_2;
	wire w_dff_B_aKZmd10S1_2;
	wire w_dff_B_P3GWNgdy4_2;
	wire w_dff_B_ptWp9URN8_2;
	wire w_dff_B_Pw44QFse8_2;
	wire w_dff_B_nJAi9NUS2_2;
	wire w_dff_B_xgBntN4U4_2;
	wire w_dff_B_UBMDuBur1_2;
	wire w_dff_B_GcmFsTjW1_2;
	wire w_dff_B_hTY2G8Qz6_2;
	wire w_dff_B_XaXDB1un7_1;
	wire w_dff_B_3AYx6PUb7_2;
	wire w_dff_B_LQ3iHkdQ4_2;
	wire w_dff_B_H27fDRbF5_2;
	wire w_dff_B_nKPtcQ663_2;
	wire w_dff_B_TEIh8Wse9_2;
	wire w_dff_B_ktNZMjEI5_2;
	wire w_dff_B_BeC7EHWL6_2;
	wire w_dff_B_qJimZa2S7_2;
	wire w_dff_B_Qu8p78dQ7_2;
	wire w_dff_B_p96mk8IX7_2;
	wire w_dff_B_VZOo691w6_2;
	wire w_dff_B_D0bKMrlm2_2;
	wire w_dff_B_YHb5QV8n9_2;
	wire w_dff_B_2eL7hIAR7_2;
	wire w_dff_B_n0acGMyX6_2;
	wire w_dff_B_MdHYQ9QH5_2;
	wire w_dff_B_2zdPCp3j5_1;
	wire w_dff_B_fBUYFPWv9_2;
	wire w_dff_B_nLXPnEUn5_2;
	wire w_dff_B_Lb1EoDNV4_2;
	wire w_dff_B_e5TTvIDn2_2;
	wire w_dff_B_8xb3SKbj7_2;
	wire w_dff_B_8pmgmrqv9_2;
	wire w_dff_B_UUxAbdPb9_2;
	wire w_dff_B_tH1kPjGu9_2;
	wire w_dff_B_xiCsUoNt2_2;
	wire w_dff_B_CzKDmZqK4_2;
	wire w_dff_B_o71D0EqK8_2;
	wire w_dff_B_lpY4cnop9_2;
	wire w_dff_B_u8z9iEiN3_2;
	wire w_dff_B_y8neqvKc3_1;
	wire w_dff_B_kyr9crAz3_2;
	wire w_dff_B_a1diWAbW8_2;
	wire w_dff_B_vWOEN5Am9_2;
	wire w_dff_B_qTCT4rn00_2;
	wire w_dff_B_OV1Rcg7f1_2;
	wire w_dff_B_jYusxhKz8_2;
	wire w_dff_B_OOlb4gtb7_2;
	wire w_dff_B_p6zTNLbH6_2;
	wire w_dff_B_RQbxMgue5_2;
	wire w_dff_B_YSaWgmih5_2;
	wire w_dff_B_Ahgr0w2R0_1;
	wire w_dff_B_f3hDQk3h4_2;
	wire w_dff_B_zeCKEgXy2_2;
	wire w_dff_B_ds9YZXoq9_2;
	wire w_dff_B_aeIqsUPX2_2;
	wire w_dff_B_b74r9Gi62_2;
	wire w_dff_B_GKEotS8a1_2;
	wire w_dff_B_3qcV8KCs4_2;
	wire w_dff_B_aPUqMr1Q7_2;
	wire w_dff_B_RrCKCGtT2_2;
	wire w_dff_B_SKjCMl7v6_2;
	wire w_dff_B_Vp1e94050_0;
	wire w_dff_B_eXsPARqE7_0;
	wire w_dff_A_DlOdnnnI0_1;
	wire w_dff_A_SO1P2mKd0_1;
	wire w_dff_B_P9F6kZrV9_1;
	wire w_dff_B_oqfRcZfn8_1;
	wire w_dff_B_EVVFRqZg9_2;
	wire w_dff_B_awF2P6AN6_2;
	wire w_dff_B_8EQXT19O0_2;
	wire w_dff_B_DfazqAdr5_2;
	wire w_dff_B_e4opkjwI4_2;
	wire w_dff_B_2am6qQWW5_2;
	wire w_dff_B_ADZmoE0x3_2;
	wire w_dff_B_rRFl05J20_2;
	wire w_dff_B_Etxsq8lX1_2;
	wire w_dff_B_bdHEFPg50_2;
	wire w_dff_B_WkyDX7Ym8_2;
	wire w_dff_B_VxLzf2U09_2;
	wire w_dff_B_0Op7r6oD3_2;
	wire w_dff_B_aOsRYIrX9_2;
	wire w_dff_B_QkMcCj3B1_2;
	wire w_dff_B_43t4PVte6_2;
	wire w_dff_B_OT7JCWRn5_2;
	wire w_dff_B_YDaXchOg2_2;
	wire w_dff_B_wgCOrgMY7_2;
	wire w_dff_B_RhUz6OvF2_2;
	wire w_dff_B_2MlIBitM5_2;
	wire w_dff_B_2VF38Yei9_2;
	wire w_dff_B_RgLwhXgw5_2;
	wire w_dff_B_WjSiQqSf8_2;
	wire w_dff_B_2TAtEa473_2;
	wire w_dff_B_TsjUJFQZ1_2;
	wire w_dff_B_D0KO3jPT7_2;
	wire w_dff_B_Gm9f3XRR9_2;
	wire w_dff_B_293qiK9z6_2;
	wire w_dff_B_mvUxN0mq1_2;
	wire w_dff_B_SOCLBoWa4_2;
	wire w_dff_B_oKEjuQty0_2;
	wire w_dff_B_ayF3F6j89_2;
	wire w_dff_B_fpGvMBxt1_2;
	wire w_dff_B_NX1yYp398_2;
	wire w_dff_B_u3FVPYPI5_2;
	wire w_dff_B_Y5CJJox81_2;
	wire w_dff_B_8eo7xoXf6_2;
	wire w_dff_B_qISSE5J91_2;
	wire w_dff_B_LEndyedm0_2;
	wire w_dff_B_oyWtLiPE7_2;
	wire w_dff_B_fiNWfDKF5_2;
	wire w_dff_B_6HkBwK4T1_2;
	wire w_dff_B_nzO81hGf5_2;
	wire w_dff_B_k6qpMpUd0_2;
	wire w_dff_B_5rgbaAfY4_2;
	wire w_dff_B_2agerOhh0_1;
	wire w_dff_B_plRlcrQy1_2;
	wire w_dff_B_XHyuMrUU8_2;
	wire w_dff_B_xRCoA3tL9_2;
	wire w_dff_B_bgdDR2Tq7_2;
	wire w_dff_B_o8xBbSY07_2;
	wire w_dff_B_BppLBu097_2;
	wire w_dff_B_w7DjH2Zj6_2;
	wire w_dff_B_GwUYymFD8_2;
	wire w_dff_B_NLaVXcXC1_2;
	wire w_dff_B_CvXsLa9q4_2;
	wire w_dff_B_aWKAKEWC6_2;
	wire w_dff_B_PCkpH6ki9_2;
	wire w_dff_B_IjzZGE777_2;
	wire w_dff_B_vwlhKaln2_2;
	wire w_dff_B_4r9cV33p6_2;
	wire w_dff_B_bcFjwpJ61_2;
	wire w_dff_B_g1QVrJ7F6_2;
	wire w_dff_B_UqJogqPs6_2;
	wire w_dff_B_mqTMNk6f9_2;
	wire w_dff_B_WRGjUugp9_2;
	wire w_dff_B_R0w3avMd0_2;
	wire w_dff_B_NpBR11xX4_2;
	wire w_dff_B_VUN5HsKF1_2;
	wire w_dff_B_HFrn3sbE3_2;
	wire w_dff_B_xXFSDG067_2;
	wire w_dff_B_sypxpxNa8_2;
	wire w_dff_B_SVqo9Ppz3_2;
	wire w_dff_B_YnURCieT3_2;
	wire w_dff_B_CZqbhFpD0_2;
	wire w_dff_B_3qa0X0CI2_2;
	wire w_dff_B_xjHt7fKf4_2;
	wire w_dff_B_BQP1rre78_2;
	wire w_dff_B_l59G6I9D3_2;
	wire w_dff_B_bKRVCC3o7_2;
	wire w_dff_B_pey6Gaoz4_2;
	wire w_dff_B_XvTtMi7d7_2;
	wire w_dff_B_R1QsuEeq6_2;
	wire w_dff_B_9Mpx2Jkw4_2;
	wire w_dff_B_X7HNuwVK1_2;
	wire w_dff_B_osmQoWUC6_2;
	wire w_dff_B_zeGKJ73x9_2;
	wire w_dff_B_SP7NRKBw2_2;
	wire w_dff_B_JZOAAh0m7_1;
	wire w_dff_B_SfGCj1NX8_2;
	wire w_dff_B_BKn5tQhV2_2;
	wire w_dff_B_z8sYq6UD6_2;
	wire w_dff_B_K5y0Uywy1_2;
	wire w_dff_B_yEYlMSue0_2;
	wire w_dff_B_Y37g2gjH6_2;
	wire w_dff_B_kbGAFFd82_2;
	wire w_dff_B_jV8hqtSE5_2;
	wire w_dff_B_qmC5z9LQ6_2;
	wire w_dff_B_VXvuDzya9_2;
	wire w_dff_B_aYTOhepd7_2;
	wire w_dff_B_eFbGPJ9D4_2;
	wire w_dff_B_xJpviDem3_2;
	wire w_dff_B_FsBFaBbz5_2;
	wire w_dff_B_3emKv7rM0_2;
	wire w_dff_B_XC3gfv0r1_2;
	wire w_dff_B_rMrBkCUc2_2;
	wire w_dff_B_BtrmtMzp4_2;
	wire w_dff_B_B1JvIKgZ8_2;
	wire w_dff_B_UxY7OPnX1_2;
	wire w_dff_B_pPFbDXp40_2;
	wire w_dff_B_3UVQFIHO7_2;
	wire w_dff_B_4Zi5bA0R3_2;
	wire w_dff_B_xJY3JMIk0_2;
	wire w_dff_B_o4TAkCq11_2;
	wire w_dff_B_nBtW83Wj8_2;
	wire w_dff_B_yrFlx6x65_2;
	wire w_dff_B_odXFmtme4_2;
	wire w_dff_B_xkzBdazl2_2;
	wire w_dff_B_Uv6GYbcM8_2;
	wire w_dff_B_CHfjPQzu2_2;
	wire w_dff_B_abwMh0ZC7_2;
	wire w_dff_B_2NZmxyyc6_2;
	wire w_dff_B_tnnsRXoL7_2;
	wire w_dff_B_NeNp9QR70_2;
	wire w_dff_B_tA00dRxH2_2;
	wire w_dff_B_zPu8CIsz0_2;
	wire w_dff_B_tWfpopR90_1;
	wire w_dff_B_5xmqKnFL5_2;
	wire w_dff_B_ZZbxtirt1_2;
	wire w_dff_B_9R46VbSd3_2;
	wire w_dff_B_4qQeQjl38_2;
	wire w_dff_B_idy0wPN87_2;
	wire w_dff_B_1m2z7O3Y4_2;
	wire w_dff_B_OUWuT4dg8_2;
	wire w_dff_B_Tmf8wHcL6_2;
	wire w_dff_B_fOpeZru06_2;
	wire w_dff_B_95d57tZi2_2;
	wire w_dff_B_CdyXRYiv6_2;
	wire w_dff_B_2a3lZlvX8_2;
	wire w_dff_B_UCKJ8daa0_2;
	wire w_dff_B_k40dRXGm8_2;
	wire w_dff_B_5G0zsCcN3_2;
	wire w_dff_B_o4Hb9KNs8_2;
	wire w_dff_B_m9ajCnLM7_2;
	wire w_dff_B_o2RQk1c75_2;
	wire w_dff_B_jWFOf66m4_2;
	wire w_dff_B_CZszh0S51_2;
	wire w_dff_B_RgbMZKsJ8_2;
	wire w_dff_B_sOV6mkJm6_2;
	wire w_dff_B_ZxU2XHPK0_2;
	wire w_dff_B_izXJIk7T0_2;
	wire w_dff_B_YAhRNZkW1_2;
	wire w_dff_B_Ct9c1h916_2;
	wire w_dff_B_JxsqKyAW5_2;
	wire w_dff_B_t1XGfg2G0_2;
	wire w_dff_B_FDFs0Ajd6_2;
	wire w_dff_B_diqJhKW81_2;
	wire w_dff_B_bb24lChW1_2;
	wire w_dff_B_nbpakffp1_2;
	wire w_dff_B_3JPXeLls3_2;
	wire w_dff_B_8iCog5Rp9_2;
	wire w_dff_B_BysUlr9y6_1;
	wire w_dff_B_qz2j93Cu9_2;
	wire w_dff_B_pzVR9Z3b0_2;
	wire w_dff_B_RFuSuZLs4_2;
	wire w_dff_B_VPhVP4Xt9_2;
	wire w_dff_B_MxhLVDQj8_2;
	wire w_dff_B_2LXPNHTf1_2;
	wire w_dff_B_yXpl13D91_2;
	wire w_dff_B_cX3mh0TA6_2;
	wire w_dff_B_HcaSunOj6_2;
	wire w_dff_B_iS1G2Wt26_2;
	wire w_dff_B_OuvjgAH26_2;
	wire w_dff_B_gJfVkYUi5_2;
	wire w_dff_B_w3JLBf8L0_2;
	wire w_dff_B_uvdapXKf3_2;
	wire w_dff_B_mB0mnk9N8_2;
	wire w_dff_B_XObe7jZ28_2;
	wire w_dff_B_VzGhWh159_2;
	wire w_dff_B_dSok3YC12_2;
	wire w_dff_B_ZOD1UMvF8_2;
	wire w_dff_B_uIlMGlyK7_2;
	wire w_dff_B_q5hiiK7n0_2;
	wire w_dff_B_1rXs8uF41_2;
	wire w_dff_B_QItZIc6D2_2;
	wire w_dff_B_DrbFUlg39_2;
	wire w_dff_B_ScDjIgIN3_2;
	wire w_dff_B_SDXyv6ay4_2;
	wire w_dff_B_BEQgbryD0_2;
	wire w_dff_B_UImHBzLF6_2;
	wire w_dff_B_KwO1WfyY5_2;
	wire w_dff_B_2FHoCyLs4_2;
	wire w_dff_B_9RmJStxt8_2;
	wire w_dff_B_bl7gv11g3_1;
	wire w_dff_B_sgctC2ms6_2;
	wire w_dff_B_QDlLT5Dg2_2;
	wire w_dff_B_5PJko8JB2_2;
	wire w_dff_B_xg0tMxRL1_2;
	wire w_dff_B_I9VxXEZz3_2;
	wire w_dff_B_tL0DKbUx6_2;
	wire w_dff_B_QuV1SDT26_2;
	wire w_dff_B_BV28o4XO2_2;
	wire w_dff_B_70khY1v44_2;
	wire w_dff_B_6F2iZ29O1_2;
	wire w_dff_B_jgAw1G9q7_2;
	wire w_dff_B_sOofq8fZ9_2;
	wire w_dff_B_mDwnVTuZ6_2;
	wire w_dff_B_h4Szrg7x8_2;
	wire w_dff_B_gEc78X3u3_2;
	wire w_dff_B_FOoxqQW81_2;
	wire w_dff_B_zFZf0V4C5_2;
	wire w_dff_B_ccihcXOc7_2;
	wire w_dff_B_BYTy5ETk6_2;
	wire w_dff_B_dgjtkW2T1_2;
	wire w_dff_B_h6GEwEum3_2;
	wire w_dff_B_x0NX5xOp9_2;
	wire w_dff_B_KKb1EUnh2_2;
	wire w_dff_B_lAiRSUL17_2;
	wire w_dff_B_ZtL614pE9_2;
	wire w_dff_B_nJVDWohz7_2;
	wire w_dff_B_VjjXjdD76_2;
	wire w_dff_B_aBR7h1Hy2_2;
	wire w_dff_B_aD7x3mA87_1;
	wire w_dff_B_THAfjzzN6_2;
	wire w_dff_B_fpMykrte6_2;
	wire w_dff_B_i5MGwZqR6_2;
	wire w_dff_B_wrL4KYTs4_2;
	wire w_dff_B_up88BSOY2_2;
	wire w_dff_B_JXgeXzgy7_2;
	wire w_dff_B_S2FjTR3z9_2;
	wire w_dff_B_NE2Htc2V6_2;
	wire w_dff_B_ZDuH2iOY1_2;
	wire w_dff_B_a2saWzPG6_2;
	wire w_dff_B_Ru4ExJ7l9_2;
	wire w_dff_B_p4PIKxPn9_2;
	wire w_dff_B_IYBh4PKs9_2;
	wire w_dff_B_gn1RbeKP9_2;
	wire w_dff_B_JobxkEj82_2;
	wire w_dff_B_eyyG0nGG4_2;
	wire w_dff_B_SMrOrYep3_2;
	wire w_dff_B_wQB0DR4o7_2;
	wire w_dff_B_SnnuDMwd1_2;
	wire w_dff_B_yA9eEGGP0_2;
	wire w_dff_B_2AykSPL21_2;
	wire w_dff_B_F7yXKers5_2;
	wire w_dff_B_li0uOzq46_2;
	wire w_dff_B_0cTUdrvL2_2;
	wire w_dff_B_zTSUf4yg2_2;
	wire w_dff_B_JMosQLe99_1;
	wire w_dff_B_evkuoxgF7_2;
	wire w_dff_B_vmepfc7l6_2;
	wire w_dff_B_Uv072pIe8_2;
	wire w_dff_B_WiOPty1Y5_2;
	wire w_dff_B_COZ8HxcW5_2;
	wire w_dff_B_pkToUIgK6_2;
	wire w_dff_B_SHoS1vMN9_2;
	wire w_dff_B_tuZ4q8mk1_2;
	wire w_dff_B_adbh6YNe3_2;
	wire w_dff_B_PicBMPJH2_2;
	wire w_dff_B_5lGIudHz2_2;
	wire w_dff_B_kVmSAe5U9_2;
	wire w_dff_B_0EcuB2rK7_2;
	wire w_dff_B_xUEFUTM94_2;
	wire w_dff_B_Yb3MFoWe3_2;
	wire w_dff_B_V3ysKATD7_2;
	wire w_dff_B_lki6xDrr8_2;
	wire w_dff_B_DgVIYWTG7_2;
	wire w_dff_B_zB03IuIx7_2;
	wire w_dff_B_xAiTgPQE0_2;
	wire w_dff_B_VqpNoIgB5_2;
	wire w_dff_B_zFtsBFuG7_2;
	wire w_dff_B_U0htOr0J6_1;
	wire w_dff_B_KUgqZjEE7_2;
	wire w_dff_B_wxUNL26q6_2;
	wire w_dff_B_xiJ0v6c28_2;
	wire w_dff_B_vQplVdSV2_2;
	wire w_dff_B_Cl9pVdzs3_2;
	wire w_dff_B_KlkEIGIx6_2;
	wire w_dff_B_FBu0J2Su7_2;
	wire w_dff_B_w6KgQCQM0_2;
	wire w_dff_B_i4Dilrae4_2;
	wire w_dff_B_3KyqIZti9_2;
	wire w_dff_B_LwtuXjcv0_2;
	wire w_dff_B_8fQ49QiS7_2;
	wire w_dff_B_fEVbJMi30_2;
	wire w_dff_B_juLqisgc0_2;
	wire w_dff_B_wfezRKVB2_2;
	wire w_dff_B_GbsgmZ433_2;
	wire w_dff_B_iPrzVBwB6_2;
	wire w_dff_B_mLPwvyRw6_2;
	wire w_dff_B_XQlWpnvd2_2;
	wire w_dff_B_Iyryb7Ag3_1;
	wire w_dff_B_L0df6ITD8_2;
	wire w_dff_B_aOQyFdbY0_2;
	wire w_dff_B_znBRIrXq5_2;
	wire w_dff_B_gN9lqP0x1_2;
	wire w_dff_B_ktn6rVR98_2;
	wire w_dff_B_a7BAjz0B0_2;
	wire w_dff_B_WXQdLsEp9_2;
	wire w_dff_B_IZ0zSYvF3_2;
	wire w_dff_B_ttIhVM3d9_2;
	wire w_dff_B_ye0jgQYT3_2;
	wire w_dff_B_BW6TAmCM6_2;
	wire w_dff_B_0g5TJARm0_2;
	wire w_dff_B_y88AwWPC6_2;
	wire w_dff_B_NSpNPeqM5_2;
	wire w_dff_B_ZMuS2v2G9_2;
	wire w_dff_B_6WoNTM9e2_2;
	wire w_dff_B_3fp6Nyge0_1;
	wire w_dff_B_HOEKbKf41_2;
	wire w_dff_B_vuuZnh450_2;
	wire w_dff_B_Zjcsl5wP6_2;
	wire w_dff_B_nUi9cYoc0_2;
	wire w_dff_B_NYBsgyeo4_2;
	wire w_dff_B_ZaJKuGs42_2;
	wire w_dff_B_5cZYg6TB4_2;
	wire w_dff_B_r93McewT1_2;
	wire w_dff_B_P3Fm3UB04_2;
	wire w_dff_B_2p6Rr5Ra2_2;
	wire w_dff_B_X7aUmSwt2_2;
	wire w_dff_B_lBNBFkrK6_2;
	wire w_dff_B_LAmdmyhz3_2;
	wire w_dff_B_yNEAHrJk0_1;
	wire w_dff_B_n9ZaYF507_2;
	wire w_dff_B_02VdiIyv7_2;
	wire w_dff_B_gcgRUa4g5_2;
	wire w_dff_B_pUFMYXEQ9_2;
	wire w_dff_B_7KSL262Q3_2;
	wire w_dff_B_XhUVsXSg9_2;
	wire w_dff_B_XXTPQTv89_2;
	wire w_dff_B_5DEFtKar6_2;
	wire w_dff_B_B1atzNu17_2;
	wire w_dff_B_nxiq51Ud2_2;
	wire w_dff_B_bmAOyLyk1_1;
	wire w_dff_B_0iZdEHEx9_2;
	wire w_dff_B_o53S9IqX2_2;
	wire w_dff_B_lcyoUKLj0_2;
	wire w_dff_B_SOX6ZN0Z6_2;
	wire w_dff_B_cxulTZoH0_2;
	wire w_dff_B_8W3jZQuq6_2;
	wire w_dff_B_iUG0sUcw6_2;
	wire w_dff_B_JuzekZtg4_2;
	wire w_dff_B_xb9va1oA8_2;
	wire w_dff_B_xEacR6If5_2;
	wire w_dff_B_r3s5Qos04_0;
	wire w_dff_A_3QQsrz8h0_0;
	wire w_dff_A_tqDlP7NW9_0;
	wire w_dff_A_qChiSjTT1_0;
	wire w_dff_A_9ki8toQ61_0;
	wire w_dff_B_0Tq9flrP8_1;
	wire w_dff_B_RC3DzLJi9_2;
	wire w_dff_B_41vVKmW97_2;
	wire w_dff_B_Vy2zL9cD0_2;
	wire w_dff_B_xvNydhBx9_2;
	wire w_dff_B_yYeXScd81_2;
	wire w_dff_B_xe1jJSAf0_2;
	wire w_dff_B_FMKqSaua2_2;
	wire w_dff_B_H9R5l9Ci5_2;
	wire w_dff_B_RJ6utOV02_2;
	wire w_dff_B_CqkL9ZQR2_2;
	wire w_dff_B_8xhQzuQ41_2;
	wire w_dff_B_qXaQoU6P6_2;
	wire w_dff_B_vOouALVs6_2;
	wire w_dff_B_4TpawNZv0_2;
	wire w_dff_B_HkU3zgBf5_2;
	wire w_dff_B_506aG5TU7_2;
	wire w_dff_B_iMfTyXVX4_2;
	wire w_dff_B_Psn9Xlde3_2;
	wire w_dff_B_MdIewARP2_2;
	wire w_dff_B_PyGevuDR5_2;
	wire w_dff_B_vjyZ07B55_2;
	wire w_dff_B_yMMg5mFA0_2;
	wire w_dff_B_p3mljQqH1_2;
	wire w_dff_B_ga7XhXMp3_2;
	wire w_dff_B_50FIKzDS2_2;
	wire w_dff_B_gp9e7UAL7_2;
	wire w_dff_B_8ZNOG0zT5_2;
	wire w_dff_B_bTM5Vijz5_2;
	wire w_dff_B_ghHWn50z7_2;
	wire w_dff_B_MKu59GoH2_2;
	wire w_dff_B_UP3upJe72_2;
	wire w_dff_B_Gt73K3dY1_2;
	wire w_dff_B_nmZshGw77_2;
	wire w_dff_B_TdlP5mEs6_2;
	wire w_dff_B_RCtarpdH5_2;
	wire w_dff_B_TBChotMj6_2;
	wire w_dff_B_admalDvB7_2;
	wire w_dff_B_dVmmNH8Q3_2;
	wire w_dff_B_LgFQUSNZ4_2;
	wire w_dff_B_yPxKtyo95_2;
	wire w_dff_B_1UWqrAzI4_2;
	wire w_dff_B_ViywdTj95_2;
	wire w_dff_B_RnfD60v84_2;
	wire w_dff_B_8NRw3rHp5_2;
	wire w_dff_B_DIbn7qAF3_0;
	wire w_dff_A_lYf27aFO6_1;
	wire w_dff_B_5b7MHFLe9_1;
	wire w_dff_B_vbDbSqNB6_2;
	wire w_dff_B_OSMIUIRZ4_2;
	wire w_dff_B_LwqzFRSM7_2;
	wire w_dff_B_UWrPxdzc7_2;
	wire w_dff_B_KnFwu6QV4_2;
	wire w_dff_B_qRFYBKY82_2;
	wire w_dff_B_cZtzH5tg7_2;
	wire w_dff_B_KRrw8Jvd2_2;
	wire w_dff_B_ex9EOPU21_2;
	wire w_dff_B_O0tfZ5s76_2;
	wire w_dff_B_4ilJbEqV7_2;
	wire w_dff_B_Z7PfLtWP3_2;
	wire w_dff_B_ejOFnKkv3_2;
	wire w_dff_B_CDZaLuLw8_2;
	wire w_dff_B_YKGkE7RC2_2;
	wire w_dff_B_VdZKIYkh7_2;
	wire w_dff_B_roL2bsNd8_2;
	wire w_dff_B_B5cJly2x4_2;
	wire w_dff_B_WJc95NuN1_2;
	wire w_dff_B_9WeYMuTj5_2;
	wire w_dff_B_lyxoAaqq6_2;
	wire w_dff_B_xaBHL6Jf8_2;
	wire w_dff_B_237AxNRa0_2;
	wire w_dff_B_zjWZUXKu3_2;
	wire w_dff_B_Totrr1c28_2;
	wire w_dff_B_yHnZ6pZd3_2;
	wire w_dff_B_CaqJxvK11_2;
	wire w_dff_B_buvGEhHE4_2;
	wire w_dff_B_21VvH6B65_2;
	wire w_dff_B_C1ONkMfs3_2;
	wire w_dff_B_MMXkNZlI3_2;
	wire w_dff_B_g2Wjjm5N4_2;
	wire w_dff_B_v3Ri2d5g7_2;
	wire w_dff_B_mTtG2pcZ8_2;
	wire w_dff_B_sLrCaugh6_2;
	wire w_dff_B_WTcQIfv96_2;
	wire w_dff_B_qjvsO5PI5_2;
	wire w_dff_B_2Z3H3mR92_2;
	wire w_dff_B_e1hx0Z8G3_2;
	wire w_dff_B_xyI3tAO59_2;
	wire w_dff_B_ALbNq03a9_1;
	wire w_dff_B_v2dMiSA64_2;
	wire w_dff_B_bUR6Jbse2_2;
	wire w_dff_B_LQiljXHt6_2;
	wire w_dff_B_G0NB0KcF0_2;
	wire w_dff_B_sXUbyWm39_2;
	wire w_dff_B_PF3v1WVF3_2;
	wire w_dff_B_vEeFK2NN9_2;
	wire w_dff_B_CTHnz4QK6_2;
	wire w_dff_B_KzRjYztY3_2;
	wire w_dff_B_6YWGK0mB3_2;
	wire w_dff_B_Ne9oEF0r1_2;
	wire w_dff_B_kPvIBqUA6_2;
	wire w_dff_B_DNHDwCFR7_2;
	wire w_dff_B_7h5yKv5G1_2;
	wire w_dff_B_vGzsnYHc3_2;
	wire w_dff_B_dSx3LZEv9_2;
	wire w_dff_B_D0yM60QO6_2;
	wire w_dff_B_LlfVOZ4Y4_2;
	wire w_dff_B_1ia5lneo8_2;
	wire w_dff_B_fNdXa7x81_2;
	wire w_dff_B_mnScxryE3_2;
	wire w_dff_B_mJ0XS2XH3_2;
	wire w_dff_B_0LJkCJNO9_2;
	wire w_dff_B_TYxXuLLp1_2;
	wire w_dff_B_NzfBssT10_2;
	wire w_dff_B_xqc7mgcY6_2;
	wire w_dff_B_NkXm7E5v4_2;
	wire w_dff_B_ki8dsgDd2_2;
	wire w_dff_B_KXl0rC2Y9_2;
	wire w_dff_B_Olt5ViON0_2;
	wire w_dff_B_YPMijV1J2_2;
	wire w_dff_B_FWhOfQcU2_2;
	wire w_dff_B_8DdjDPLX7_2;
	wire w_dff_B_daAklES03_2;
	wire w_dff_B_dTa0L80u3_2;
	wire w_dff_B_DZtWG4YR4_2;
	wire w_dff_B_b33kYsUA6_2;
	wire w_dff_B_tM9aG5Ne4_1;
	wire w_dff_B_X33akk7n2_2;
	wire w_dff_B_DtUVPjlF1_2;
	wire w_dff_B_rd3KiYXc9_2;
	wire w_dff_B_uCXfeUfO7_2;
	wire w_dff_B_1qA0kXFD1_2;
	wire w_dff_B_CALulnsx6_2;
	wire w_dff_B_KXVeKuOc5_2;
	wire w_dff_B_ZDdd0oX22_2;
	wire w_dff_B_qpVt4v6H0_2;
	wire w_dff_B_hhudREVW2_2;
	wire w_dff_B_cEVre46x1_2;
	wire w_dff_B_lBT0qaRG0_2;
	wire w_dff_B_uoSgA8na3_2;
	wire w_dff_B_6ioeJRdx1_2;
	wire w_dff_B_ohYpvn1y2_2;
	wire w_dff_B_mh1Qfucu0_2;
	wire w_dff_B_Km0WM7KA6_2;
	wire w_dff_B_yNq2aYil7_2;
	wire w_dff_B_AsRD1YKj7_2;
	wire w_dff_B_qH8dJJgq0_2;
	wire w_dff_B_oaSuyjv46_2;
	wire w_dff_B_bl5Iuqq96_2;
	wire w_dff_B_kxAFGSW07_2;
	wire w_dff_B_FYRkc7Ru9_2;
	wire w_dff_B_yg0LnYqi5_2;
	wire w_dff_B_I9GAGc4b3_2;
	wire w_dff_B_12DvJwqp2_2;
	wire w_dff_B_3eo30jx80_2;
	wire w_dff_B_uscUeEHA5_2;
	wire w_dff_B_ULinil997_2;
	wire w_dff_B_T2cedTRv7_2;
	wire w_dff_B_GomBGRAp5_2;
	wire w_dff_B_UrvDxQ9U4_2;
	wire w_dff_B_WAhhwlNj0_2;
	wire w_dff_B_ES8A9qFY2_1;
	wire w_dff_B_4OKM4cKp7_2;
	wire w_dff_B_GdG1bUWr0_2;
	wire w_dff_B_McEmyvUX2_2;
	wire w_dff_B_a60qLhFd6_2;
	wire w_dff_B_YzeipnX85_2;
	wire w_dff_B_lR4kSvH20_2;
	wire w_dff_B_ndTj5aDB8_2;
	wire w_dff_B_PAyzfLUT1_2;
	wire w_dff_B_g7jmvIFk6_2;
	wire w_dff_B_zoISVPjS2_2;
	wire w_dff_B_PTJKGiy70_2;
	wire w_dff_B_Dp89tbBr2_2;
	wire w_dff_B_u3fV66GJ7_2;
	wire w_dff_B_9H44FkjQ5_2;
	wire w_dff_B_b8HlkuWd3_2;
	wire w_dff_B_7sLHKdh51_2;
	wire w_dff_B_XBBSYOyr6_2;
	wire w_dff_B_AUNKYcOn9_2;
	wire w_dff_B_wAtPlfI39_2;
	wire w_dff_B_25t42bdX4_2;
	wire w_dff_B_gKD0Gxe66_2;
	wire w_dff_B_jFZoaqyw7_2;
	wire w_dff_B_HWCxjJ2i0_2;
	wire w_dff_B_HvlRzSII5_2;
	wire w_dff_B_Eq8k8tt39_2;
	wire w_dff_B_25aefGon7_2;
	wire w_dff_B_UqxYYvQe9_2;
	wire w_dff_B_psQDKeQz4_2;
	wire w_dff_B_zpf0RMsl6_2;
	wire w_dff_B_QxodiXm21_2;
	wire w_dff_B_J1SboDT76_2;
	wire w_dff_B_BEvijuvY2_1;
	wire w_dff_B_GQ3QdFvL0_2;
	wire w_dff_B_HFHh5zsi0_2;
	wire w_dff_B_aF7loKUi6_2;
	wire w_dff_B_yefhpsUQ8_2;
	wire w_dff_B_AetPeZ4R5_2;
	wire w_dff_B_XXOV84DU6_2;
	wire w_dff_B_B9Vgeurz8_2;
	wire w_dff_B_cFhCzb1c5_2;
	wire w_dff_B_bHTPZ83v2_2;
	wire w_dff_B_7V3YVRwD4_2;
	wire w_dff_B_jrhUNSGX5_2;
	wire w_dff_B_HhUXOQlg9_2;
	wire w_dff_B_BcdhCkD81_2;
	wire w_dff_B_NzrZNvWT0_2;
	wire w_dff_B_V5hvzjcu8_2;
	wire w_dff_B_U0ueuIPn1_2;
	wire w_dff_B_kW9adihj2_2;
	wire w_dff_B_obvdkl5p8_2;
	wire w_dff_B_a42tlBsV7_2;
	wire w_dff_B_nJmuKdlf0_2;
	wire w_dff_B_IRynea0h1_2;
	wire w_dff_B_KwqeBfpv8_2;
	wire w_dff_B_8FlsdvU64_2;
	wire w_dff_B_rfX2w4o63_2;
	wire w_dff_B_7jqHOznN0_2;
	wire w_dff_B_UtuN7ZTW3_2;
	wire w_dff_B_hrcXJnDK9_2;
	wire w_dff_B_svrYkw6u9_2;
	wire w_dff_B_FXe6CwUR4_1;
	wire w_dff_B_t1XBVJht3_2;
	wire w_dff_B_rSySyf5D7_2;
	wire w_dff_B_iks8NdLb4_2;
	wire w_dff_B_ViliiN2U3_2;
	wire w_dff_B_gEyCpVS98_2;
	wire w_dff_B_qozLjBPJ2_2;
	wire w_dff_B_61jcc8J72_2;
	wire w_dff_B_wcCzGFN59_2;
	wire w_dff_B_RUamuXrZ0_2;
	wire w_dff_B_X7mtnsEN2_2;
	wire w_dff_B_sEaYM43W3_2;
	wire w_dff_B_JpJF7PRE8_2;
	wire w_dff_B_xdYxnhQO8_2;
	wire w_dff_B_nRnL4E6W4_2;
	wire w_dff_B_lSIZ6eIi9_2;
	wire w_dff_B_zlKdYJbH3_2;
	wire w_dff_B_m1YmdJ9t1_2;
	wire w_dff_B_0MKCJrkr1_2;
	wire w_dff_B_jLR83C9x0_2;
	wire w_dff_B_Qn3XVrj43_2;
	wire w_dff_B_5EVpO9IP8_2;
	wire w_dff_B_6p0ufAyi4_2;
	wire w_dff_B_c3qKAM3p1_2;
	wire w_dff_B_96dG2lku2_2;
	wire w_dff_B_uPSobetU8_2;
	wire w_dff_B_1euSCDwy0_1;
	wire w_dff_B_jdaWrV129_2;
	wire w_dff_B_Ws6j2AqG6_2;
	wire w_dff_B_JEHKea2e6_2;
	wire w_dff_B_46kIN4dJ8_2;
	wire w_dff_B_tEth13KY7_2;
	wire w_dff_B_BlB4pSDy7_2;
	wire w_dff_B_aomaS7Ha4_2;
	wire w_dff_B_opUpP3oK8_2;
	wire w_dff_B_r8wvA1h25_2;
	wire w_dff_B_P0oLKxNr5_2;
	wire w_dff_B_yTXSK4yW0_2;
	wire w_dff_B_2UHkJSm74_2;
	wire w_dff_B_nzMkGFDw9_2;
	wire w_dff_B_QyOBWDvR4_2;
	wire w_dff_B_PvIhAwNA1_2;
	wire w_dff_B_6f40NG5z5_2;
	wire w_dff_B_b5xwAwts8_2;
	wire w_dff_B_mu7wUGIp4_2;
	wire w_dff_B_OmTfFvBC3_2;
	wire w_dff_B_se3F7SJA5_2;
	wire w_dff_B_QQcdNQza5_2;
	wire w_dff_B_lgr9fuJH8_2;
	wire w_dff_B_uy2SawVe8_1;
	wire w_dff_B_vzemtAjL1_2;
	wire w_dff_B_yFFYn2TD0_2;
	wire w_dff_B_snmph6z98_2;
	wire w_dff_B_sy3F2kV40_2;
	wire w_dff_B_qUdlNRve4_2;
	wire w_dff_B_hSyDXdHs6_2;
	wire w_dff_B_zCYVFSva2_2;
	wire w_dff_B_ovYZAF3U1_2;
	wire w_dff_B_k47Nm3CI9_2;
	wire w_dff_B_iVMjVeeL9_2;
	wire w_dff_B_CfPIXJVu3_2;
	wire w_dff_B_77beoL2m7_2;
	wire w_dff_B_DSJn62HN1_2;
	wire w_dff_B_laxTxQlK7_2;
	wire w_dff_B_V24fdcLu1_2;
	wire w_dff_B_5HOpSRCc4_2;
	wire w_dff_B_k32OGgPv5_2;
	wire w_dff_B_oIoefvFy9_2;
	wire w_dff_B_nZJmTAnu1_2;
	wire w_dff_B_GXqD2o435_1;
	wire w_dff_B_yQWoVcq78_2;
	wire w_dff_B_OzxQIpyc3_2;
	wire w_dff_B_bwWGxP5g0_2;
	wire w_dff_B_b5ciOZUC7_2;
	wire w_dff_B_jFdfFPbR8_2;
	wire w_dff_B_yj84MG5C4_2;
	wire w_dff_B_ZnmMV5Gk3_2;
	wire w_dff_B_BVD23hxG1_2;
	wire w_dff_B_9ZRrLiv72_2;
	wire w_dff_B_MtSGdIjF2_2;
	wire w_dff_B_IKjg6YUZ9_2;
	wire w_dff_B_HRceJayX3_2;
	wire w_dff_B_IVbcteM63_2;
	wire w_dff_B_SsTK8xTm0_2;
	wire w_dff_B_xobzKttg0_2;
	wire w_dff_B_Ef1UaLVG5_2;
	wire w_dff_B_hSfTyuhW6_1;
	wire w_dff_B_PWQJ2Vnu3_2;
	wire w_dff_B_6B2YF9Ay1_2;
	wire w_dff_B_y9ktx8Jb5_2;
	wire w_dff_B_rjQWH52K2_2;
	wire w_dff_B_KQm4MA0M9_2;
	wire w_dff_B_gxsauXrw9_2;
	wire w_dff_B_AjTY6Lo33_2;
	wire w_dff_B_r84F0BXi2_2;
	wire w_dff_B_BVhpNlmg8_2;
	wire w_dff_B_1ZNcWDTJ4_2;
	wire w_dff_B_U1GybGGG9_2;
	wire w_dff_B_b8fAa6Jb0_2;
	wire w_dff_B_IE4fTbbZ3_2;
	wire w_dff_B_TBd7wztu5_1;
	wire w_dff_B_nNKdS2049_2;
	wire w_dff_B_NURwZw7z5_2;
	wire w_dff_B_zQUzFn1p0_2;
	wire w_dff_B_7SibxeSs7_2;
	wire w_dff_B_m9aJIOKE2_2;
	wire w_dff_B_a0Se4UDH4_2;
	wire w_dff_B_V96D4y7W9_2;
	wire w_dff_B_Y6VQH7IZ4_2;
	wire w_dff_B_CbvTIG0O8_2;
	wire w_dff_B_n3Z6e0v41_2;
	wire w_dff_B_YoDQV3J86_1;
	wire w_dff_B_GbOS7NLd1_2;
	wire w_dff_B_WQnTFrOB2_2;
	wire w_dff_B_Wors72lZ0_2;
	wire w_dff_B_X0ggv1W10_2;
	wire w_dff_B_GkuqroHq8_2;
	wire w_dff_B_7mP3ZrFy4_2;
	wire w_dff_B_6moYWDCl8_2;
	wire w_dff_B_tLxctWia2_2;
	wire w_dff_B_epZiYMrb5_2;
	wire w_dff_B_5j9PqDcD1_2;
	wire w_dff_B_vi41Mh5Q9_0;
	wire w_dff_A_T32BztU16_0;
	wire w_dff_A_Rg6AGHtF7_0;
	wire w_dff_A_5EX1W2hZ4_0;
	wire w_dff_A_nGqydeaL0_0;
	wire w_dff_B_HsitQwma1_2;
	wire w_dff_B_3Elpi5LQ4_1;
	wire w_dff_B_DRYQFlrp3_2;
	wire w_dff_B_Gl0SiJCf0_2;
	wire w_dff_B_SVeeDJSP8_2;
	wire w_dff_B_C6iZAuX13_2;
	wire w_dff_B_3IYusue31_2;
	wire w_dff_B_dEEzoEfp9_2;
	wire w_dff_B_jrBR3hNx5_2;
	wire w_dff_B_TD39RoJ25_2;
	wire w_dff_B_xE9dR0lx5_2;
	wire w_dff_B_EgN0PYJT6_2;
	wire w_dff_B_zAIScBcD5_2;
	wire w_dff_B_KgskRtnN4_2;
	wire w_dff_B_fsM45eLY9_2;
	wire w_dff_B_fbwW3KCr9_2;
	wire w_dff_B_GiWfCGXA7_2;
	wire w_dff_B_hHjCLsR01_2;
	wire w_dff_B_cJtUaC1u5_2;
	wire w_dff_B_dgkr1E9x4_2;
	wire w_dff_B_VBvgpe0w2_2;
	wire w_dff_B_K0Mn1GUF2_2;
	wire w_dff_B_TgK9lkI00_2;
	wire w_dff_B_D3UkFlhV2_2;
	wire w_dff_B_X8FVcDj51_2;
	wire w_dff_B_elgSfL0S3_2;
	wire w_dff_B_IR3vG3Zu1_2;
	wire w_dff_B_aWCy2cF89_2;
	wire w_dff_B_SoLQ3Xav9_2;
	wire w_dff_B_ezl1TwEr2_2;
	wire w_dff_B_You15Nnr4_2;
	wire w_dff_B_Vl6gXDkl3_2;
	wire w_dff_B_w4nqc8XN4_2;
	wire w_dff_B_rIxlfcrw2_2;
	wire w_dff_B_YEzMr56n5_2;
	wire w_dff_B_Kwqoe2np4_2;
	wire w_dff_B_XzqoWY2q4_2;
	wire w_dff_B_N2nn0n0g0_2;
	wire w_dff_B_oybLVK4D8_2;
	wire w_dff_B_izwdhGDY8_2;
	wire w_dff_B_LFpGHjxF6_2;
	wire w_dff_B_MxUou9Hc5_2;
	wire w_dff_B_xvJ6aTvz4_2;
	wire w_dff_B_JRknODPh7_2;
	wire w_dff_B_t7ZsAJgh2_2;
	wire w_dff_B_Lo8FIWC53_2;
	wire w_dff_B_k8XlVUA97_1;
	wire w_dff_B_fAgyJvSN6_2;
	wire w_dff_B_mwyaLb3v2_2;
	wire w_dff_B_tJPE0WFp3_2;
	wire w_dff_B_68CUfuxP7_2;
	wire w_dff_B_zlNpVvvW0_2;
	wire w_dff_B_OPM4i01Q4_2;
	wire w_dff_B_fpKwXHvc4_2;
	wire w_dff_B_poSb7Tcn7_2;
	wire w_dff_B_aoMWe0xT4_2;
	wire w_dff_B_rDrlEccx5_2;
	wire w_dff_B_3FbUVB1E7_2;
	wire w_dff_B_nnpi5Kj04_2;
	wire w_dff_B_wray5jyJ6_2;
	wire w_dff_B_yJ6ZsH4o8_2;
	wire w_dff_B_jXAZaE1N3_2;
	wire w_dff_B_iYXLo5l90_2;
	wire w_dff_B_5FOah2fI3_2;
	wire w_dff_B_mnKdMAz65_2;
	wire w_dff_B_vo7eoJt71_2;
	wire w_dff_B_nEYU0SN60_2;
	wire w_dff_B_uSNmt1l58_2;
	wire w_dff_B_d5vHjC0C0_2;
	wire w_dff_B_y0Oo2BPK8_2;
	wire w_dff_B_yNKXbDM99_2;
	wire w_dff_B_m6cRa4Jl3_2;
	wire w_dff_B_DwibTo361_2;
	wire w_dff_B_hg03bV8v8_2;
	wire w_dff_B_RnFolPgg2_2;
	wire w_dff_B_CdCj96At8_2;
	wire w_dff_B_arwfT5Ft4_2;
	wire w_dff_B_tYntJP816_2;
	wire w_dff_B_jg6mtGK87_2;
	wire w_dff_B_O9ILECp82_2;
	wire w_dff_B_swlrL67e4_2;
	wire w_dff_B_A66EmYzY5_2;
	wire w_dff_B_VhcX5Szs4_2;
	wire w_dff_B_D7wBaV4Z1_2;
	wire w_dff_B_N1AHSpAn2_2;
	wire w_dff_B_39RFgBUm3_2;
	wire w_dff_B_fiwM2wYC8_1;
	wire w_dff_B_tKDdBQqd8_2;
	wire w_dff_B_qNEzsbKg7_2;
	wire w_dff_B_vUOUi9cH3_2;
	wire w_dff_B_lP8AAloD7_2;
	wire w_dff_B_W0DFx3Zh8_2;
	wire w_dff_B_ONs93hSM2_2;
	wire w_dff_B_ShxoNOvX9_2;
	wire w_dff_B_01LndCTO5_2;
	wire w_dff_B_aUKBCvj80_2;
	wire w_dff_B_eCkCW5nx3_2;
	wire w_dff_B_lqT8ZVYz1_2;
	wire w_dff_B_o8jYEeQb0_2;
	wire w_dff_B_mnKFgr1B9_2;
	wire w_dff_B_p60nv3tk8_2;
	wire w_dff_B_0BZbX3UZ5_2;
	wire w_dff_B_I14t2u4i9_2;
	wire w_dff_B_x4KC1XaE7_2;
	wire w_dff_B_t5gKtYkM3_2;
	wire w_dff_B_7k9cYEWR5_2;
	wire w_dff_B_35gFl6HC6_2;
	wire w_dff_B_DvyTw6HX9_2;
	wire w_dff_B_aRmcyMxX6_2;
	wire w_dff_B_qVlpD0Ka4_2;
	wire w_dff_B_OsW73hAU7_2;
	wire w_dff_B_gxQu3uKK3_2;
	wire w_dff_B_Ckf0V3sk5_2;
	wire w_dff_B_TFONE8Ha0_2;
	wire w_dff_B_WDDXFCA29_2;
	wire w_dff_B_kUMuguP50_2;
	wire w_dff_B_NakSXBwn8_2;
	wire w_dff_B_qRjbkKcV6_2;
	wire w_dff_B_n9cBxznM3_2;
	wire w_dff_B_ijHw9koU1_2;
	wire w_dff_B_TUI4EmhO3_2;
	wire w_dff_B_1vHsV6SF0_2;
	wire w_dff_B_J3NOWJQd2_2;
	wire w_dff_B_HfWrQ1Ho7_1;
	wire w_dff_B_KODIlDmX1_2;
	wire w_dff_B_csCOtoNU4_2;
	wire w_dff_B_9wGhnw8x6_2;
	wire w_dff_B_CMWpwJBe2_2;
	wire w_dff_B_5y4qAQ0k8_2;
	wire w_dff_B_O1yL9swT8_2;
	wire w_dff_B_K2dzaRKH4_2;
	wire w_dff_B_92z9Qms06_2;
	wire w_dff_B_cWxRY6Ya0_2;
	wire w_dff_B_pPMpScHQ3_2;
	wire w_dff_B_TYUblta39_2;
	wire w_dff_B_XIiO30kZ4_2;
	wire w_dff_B_dfNUeEuS9_2;
	wire w_dff_B_7uOR295C2_2;
	wire w_dff_B_hXbwctaK6_2;
	wire w_dff_B_gtQMHRbk1_2;
	wire w_dff_B_uzVLRekc5_2;
	wire w_dff_B_CARo65hi7_2;
	wire w_dff_B_FDTDgNN44_2;
	wire w_dff_B_YZ4VpJSX8_2;
	wire w_dff_B_OK4Ukae05_2;
	wire w_dff_B_AMWiKE6O4_2;
	wire w_dff_B_TigrChrE8_2;
	wire w_dff_B_lJhJMmwD4_2;
	wire w_dff_B_TZa3XLot5_2;
	wire w_dff_B_Ac4cxLrh2_2;
	wire w_dff_B_zROXxUve7_2;
	wire w_dff_B_UsFytzGm9_2;
	wire w_dff_B_S6HvVgXo8_2;
	wire w_dff_B_DshDVSHv6_2;
	wire w_dff_B_N5EhLutR4_2;
	wire w_dff_B_rxpvaiXx5_2;
	wire w_dff_B_lQyCJl4Y6_2;
	wire w_dff_B_RhSaeNsr6_1;
	wire w_dff_B_W1mFT3IN0_2;
	wire w_dff_B_uTZGI3sU8_2;
	wire w_dff_B_6hRcDbyc0_2;
	wire w_dff_B_fAL3bVqH2_2;
	wire w_dff_B_reVJgRRt1_2;
	wire w_dff_B_iwxoP96i4_2;
	wire w_dff_B_92Jd6xJe0_2;
	wire w_dff_B_1lN2lGqZ9_2;
	wire w_dff_B_bk9xbFrT0_2;
	wire w_dff_B_omEZxyTQ5_2;
	wire w_dff_B_BPrLBHMV3_2;
	wire w_dff_B_ZUwYEeX83_2;
	wire w_dff_B_K4w2dVa61_2;
	wire w_dff_B_tIM5N5Zq1_2;
	wire w_dff_B_hGxe35nt6_2;
	wire w_dff_B_TIjSAsJ70_2;
	wire w_dff_B_nGrFAuFj2_2;
	wire w_dff_B_CwTMXs6S7_2;
	wire w_dff_B_nlxyfOhE6_2;
	wire w_dff_B_ponracsk3_2;
	wire w_dff_B_A3eNbX6Y6_2;
	wire w_dff_B_8iMnrbZi7_2;
	wire w_dff_B_G91A9Xx24_2;
	wire w_dff_B_vlQPEQfi2_2;
	wire w_dff_B_dQVHuCkX2_2;
	wire w_dff_B_WQd0TssQ8_2;
	wire w_dff_B_Di5fBYKC8_2;
	wire w_dff_B_TpaGXncm5_2;
	wire w_dff_B_rRbimV570_2;
	wire w_dff_B_8BHbKbWp9_2;
	wire w_dff_B_QJ7JBseb2_1;
	wire w_dff_B_OHTtpgJ00_2;
	wire w_dff_B_AnhGii639_2;
	wire w_dff_B_rrnvr8jj2_2;
	wire w_dff_B_NnPK0t1N6_2;
	wire w_dff_B_hNpaOvIQ3_2;
	wire w_dff_B_FTw4nQhW1_2;
	wire w_dff_B_cXiKRgxT2_2;
	wire w_dff_B_VbYUTTOn2_2;
	wire w_dff_B_IKda24pJ4_2;
	wire w_dff_B_QpfYUdSV3_2;
	wire w_dff_B_4GN8XVSh0_2;
	wire w_dff_B_BPYizo1R5_2;
	wire w_dff_B_Zi2Esws10_2;
	wire w_dff_B_DzL6x2KE2_2;
	wire w_dff_B_W828Mu7m0_2;
	wire w_dff_B_faAN3UCE9_2;
	wire w_dff_B_Y2TeiGFM2_2;
	wire w_dff_B_D1Mgrz1W5_2;
	wire w_dff_B_cWLBa6684_2;
	wire w_dff_B_LA41AzYl7_2;
	wire w_dff_B_hnH68s2H6_2;
	wire w_dff_B_kAYKam8T5_2;
	wire w_dff_B_ZxOyhqWS8_2;
	wire w_dff_B_XcjG0ExS7_2;
	wire w_dff_B_1kkDEOlE6_2;
	wire w_dff_B_Hiw2Z4ik1_2;
	wire w_dff_B_0jYhmeDR2_2;
	wire w_dff_B_aKoY2FFS5_1;
	wire w_dff_B_7MdYhEU40_2;
	wire w_dff_B_bYsAvfoF0_2;
	wire w_dff_B_8SEpU9cv1_2;
	wire w_dff_B_IxA3BBVu1_2;
	wire w_dff_B_4VHLFzQw3_2;
	wire w_dff_B_jBQ4GdPP9_2;
	wire w_dff_B_LPjKVJF13_2;
	wire w_dff_B_MOmlbwMm4_2;
	wire w_dff_B_cr8VTA2l6_2;
	wire w_dff_B_qlilAu5e1_2;
	wire w_dff_B_nqOWRDfA9_2;
	wire w_dff_B_c95FA0pp0_2;
	wire w_dff_B_7wpSharB5_2;
	wire w_dff_B_iAoUph6s3_2;
	wire w_dff_B_10zKxQgf3_2;
	wire w_dff_B_ebOEtC5u9_2;
	wire w_dff_B_33YMv3sj6_2;
	wire w_dff_B_oOUXpSxl3_2;
	wire w_dff_B_nwcT9UN73_2;
	wire w_dff_B_3u7FlmR44_2;
	wire w_dff_B_Db3Odp5g5_2;
	wire w_dff_B_QywCoaMc4_2;
	wire w_dff_B_aWxI0aVn1_2;
	wire w_dff_B_oRp3NQyX5_2;
	wire w_dff_B_dKuj7UIM9_1;
	wire w_dff_B_q3QMKSYf2_2;
	wire w_dff_B_Aph4nQxB0_2;
	wire w_dff_B_cgHpw67p6_2;
	wire w_dff_B_sl3PHFQe5_2;
	wire w_dff_B_75yho7qO7_2;
	wire w_dff_B_oOhw1uEk5_2;
	wire w_dff_B_8eyCW8ID0_2;
	wire w_dff_B_0z2WCI0I5_2;
	wire w_dff_B_0iTd3ZHM4_2;
	wire w_dff_B_ckLG8WYz6_2;
	wire w_dff_B_FlSiSvfJ8_2;
	wire w_dff_B_KSHntsTn6_2;
	wire w_dff_B_XbMv8Vz49_2;
	wire w_dff_B_4CPKUTPl6_2;
	wire w_dff_B_RXc1X9gg8_2;
	wire w_dff_B_SrOlL3PA3_2;
	wire w_dff_B_boADKgOE7_2;
	wire w_dff_B_hG7l2ONS5_2;
	wire w_dff_B_V92Sy3Sx9_2;
	wire w_dff_B_TuM6Ewv20_2;
	wire w_dff_B_5qY27qCF0_2;
	wire w_dff_B_aQcRGXAd3_1;
	wire w_dff_B_zf7qMEU36_2;
	wire w_dff_B_H0CaMaGA1_2;
	wire w_dff_B_oot3Kj9n4_2;
	wire w_dff_B_r4T12Dzd2_2;
	wire w_dff_B_0ge5Pz5b8_2;
	wire w_dff_B_G5cskc422_2;
	wire w_dff_B_JxoS9pvz3_2;
	wire w_dff_B_heZSkhma0_2;
	wire w_dff_B_wfBTfFld2_2;
	wire w_dff_B_FXD2ZjPd2_2;
	wire w_dff_B_XJ9TIffT4_2;
	wire w_dff_B_mQTIjlwR0_2;
	wire w_dff_B_E0WKH84L1_2;
	wire w_dff_B_C7I1qSDs0_2;
	wire w_dff_B_fssYfKpV7_2;
	wire w_dff_B_Sdh0qhQX6_2;
	wire w_dff_B_fPtc7Jlv2_2;
	wire w_dff_B_5g0nQWiE2_2;
	wire w_dff_B_P1aw5ykX6_1;
	wire w_dff_B_NXFFFSE95_2;
	wire w_dff_B_qUFF4Dlu1_2;
	wire w_dff_B_PmlSuEvl6_2;
	wire w_dff_B_9BnGul3M6_2;
	wire w_dff_B_sIjyY2IA6_2;
	wire w_dff_B_wNgmwsv64_2;
	wire w_dff_B_8kIr1eeO8_2;
	wire w_dff_B_JY2n58mY7_2;
	wire w_dff_B_x1U1S38Z9_2;
	wire w_dff_B_ZXqKzxfj4_2;
	wire w_dff_B_hpZCRbIk6_2;
	wire w_dff_B_3GJtlzYM1_2;
	wire w_dff_B_zgg8Tj2w8_2;
	wire w_dff_B_4w8tkCCg1_2;
	wire w_dff_B_L4ZbzIDi7_2;
	wire w_dff_B_6HH7rVy35_1;
	wire w_dff_B_gVsqYsu18_2;
	wire w_dff_B_ytMNg9Lb1_2;
	wire w_dff_B_6WZRlhWR4_2;
	wire w_dff_B_h0LQLSH50_2;
	wire w_dff_B_I3EjWxr31_2;
	wire w_dff_B_SlXB7Bt70_2;
	wire w_dff_B_HPsLlWeB0_2;
	wire w_dff_B_ulNJqK5x1_2;
	wire w_dff_B_vy5M9ujs3_2;
	wire w_dff_B_3FelmzPf6_2;
	wire w_dff_B_I2vQsKeF9_2;
	wire w_dff_B_hhHb4CZS5_2;
	wire w_dff_B_YL95S5n31_1;
	wire w_dff_B_87uMtoxF9_2;
	wire w_dff_B_HJqRWbSf9_2;
	wire w_dff_B_8yUtVIQm2_2;
	wire w_dff_B_L2En0x2s0_2;
	wire w_dff_B_G4hiu4kD4_2;
	wire w_dff_B_sceqQ9rB1_2;
	wire w_dff_B_Qh4mReII3_2;
	wire w_dff_B_IZ53g2WM5_2;
	wire w_dff_B_9RkqwVp20_2;
	wire w_dff_B_D35Bkf912_2;
	wire w_dff_B_ir1ZwmwY5_1;
	wire w_dff_B_EfvDEuPI7_2;
	wire w_dff_B_SFqcnKhA5_2;
	wire w_dff_B_OVN1Mg9T4_2;
	wire w_dff_B_6kAhJTRB4_2;
	wire w_dff_B_MKnRdFyu1_2;
	wire w_dff_B_EZJuavUv4_2;
	wire w_dff_B_KrkZHRZ11_2;
	wire w_dff_B_HOBApmeT6_2;
	wire w_dff_B_yNro1q3L6_2;
	wire w_dff_B_DPQAd0JT2_2;
	wire w_dff_B_dFtM3qTM2_0;
	wire w_dff_A_ltPdOqju8_0;
	wire w_dff_A_JUhNNVgm0_0;
	wire w_dff_A_Kt85JJ044_1;
	wire w_dff_A_ZLkAxtuN9_1;
	wire w_dff_B_8w74N4ai7_2;
	wire w_dff_B_tyeEbBLJ7_1;
	wire w_dff_B_fVuhJmVK5_2;
	wire w_dff_B_ZJenFmRo7_2;
	wire w_dff_B_HPTKlO0P7_2;
	wire w_dff_B_QutrbreA6_2;
	wire w_dff_B_nk9i37RL3_2;
	wire w_dff_B_Y8DcatZY5_2;
	wire w_dff_B_daMRik372_2;
	wire w_dff_B_TuZLNalW6_2;
	wire w_dff_B_cJyEoYtY8_2;
	wire w_dff_B_uPwcfmdA8_2;
	wire w_dff_B_FdUkVYnb0_2;
	wire w_dff_B_M7U83DY40_2;
	wire w_dff_B_qhWFS2cL0_2;
	wire w_dff_B_jcnHWUJX7_2;
	wire w_dff_B_v5yd2RQ81_2;
	wire w_dff_B_IICoYyHR3_2;
	wire w_dff_B_pmRUkfVb4_2;
	wire w_dff_B_mh4S1d5X4_2;
	wire w_dff_B_S5gXFcqx8_2;
	wire w_dff_B_UdVJUrad3_2;
	wire w_dff_B_CuWwkZcY5_2;
	wire w_dff_B_w0cZCKHO9_2;
	wire w_dff_B_6Z3bVJ5f8_2;
	wire w_dff_B_yzFAqiAR7_2;
	wire w_dff_B_7iYX3Mei0_2;
	wire w_dff_B_6pPTLiTa6_2;
	wire w_dff_B_IoZO6PAx8_2;
	wire w_dff_B_yAXuRTv26_2;
	wire w_dff_B_VNPO8uiN9_2;
	wire w_dff_B_B79uhzjP3_2;
	wire w_dff_B_BlxmijrU6_2;
	wire w_dff_B_58QYTuvJ5_2;
	wire w_dff_B_QTjHgQ1H1_2;
	wire w_dff_B_pbLRlp6D9_2;
	wire w_dff_B_fGObqosS0_2;
	wire w_dff_B_ebXtDkaj5_2;
	wire w_dff_B_2y2RXh0P5_2;
	wire w_dff_B_frlZztg88_2;
	wire w_dff_B_AzscMRNQ4_2;
	wire w_dff_B_bWQfYQug0_2;
	wire w_dff_B_IMR3K2bM4_2;
	wire w_dff_B_wosXpw0K0_2;
	wire w_dff_B_hpoS111w6_2;
	wire w_dff_B_Sr0ExSmE5_2;
	wire w_dff_B_RlCGGr5Y0_2;
	wire w_dff_B_NdHYw2Ji4_1;
	wire w_dff_B_U6Ubw3pp7_2;
	wire w_dff_B_8y31KhAG1_2;
	wire w_dff_B_WDuo4Wx99_2;
	wire w_dff_B_wbsBZ0wh1_2;
	wire w_dff_B_XQBzbO711_2;
	wire w_dff_B_POkTLrYn1_2;
	wire w_dff_B_3Z2dZ2y55_2;
	wire w_dff_B_5C0cvymz5_2;
	wire w_dff_B_KISb0sGm6_2;
	wire w_dff_B_fFfPC3k22_2;
	wire w_dff_B_UG0yZ99Q3_2;
	wire w_dff_B_SLXdx0D89_2;
	wire w_dff_B_oX0d8D2Y1_2;
	wire w_dff_B_Mxmc4wt85_2;
	wire w_dff_B_mrGCGhk83_2;
	wire w_dff_B_LAW0QPg33_2;
	wire w_dff_B_OQrWFPAw2_2;
	wire w_dff_B_gzs3GLYf8_2;
	wire w_dff_B_D9EZcvwU9_2;
	wire w_dff_B_kn0MMw319_2;
	wire w_dff_B_xyfehsFM1_2;
	wire w_dff_B_4OmD33P44_2;
	wire w_dff_B_ONgPNZhT5_2;
	wire w_dff_B_hAyWX5ki0_2;
	wire w_dff_B_29g9LcSI1_2;
	wire w_dff_B_yi1YVyiv9_2;
	wire w_dff_B_MqMIe5CU8_2;
	wire w_dff_B_MJpMMPUn9_2;
	wire w_dff_B_WQ9ZA4Bg5_2;
	wire w_dff_B_T6gQ6IyL3_2;
	wire w_dff_B_z4YkEEGY1_2;
	wire w_dff_B_YDMz8jpm1_2;
	wire w_dff_B_S8lu1yTv5_2;
	wire w_dff_B_EOfLXsNi3_2;
	wire w_dff_B_DVaSfitn6_2;
	wire w_dff_B_oc45YKuR1_2;
	wire w_dff_B_TpuK3uk54_2;
	wire w_dff_B_47ENbsaX8_2;
	wire w_dff_B_kyZA73wn3_2;
	wire w_dff_B_GTCAo03K0_2;
	wire w_dff_B_0H3Hy2HC2_1;
	wire w_dff_B_WaCNSFAD9_2;
	wire w_dff_B_MmTj9uej6_2;
	wire w_dff_B_iSPwaqOV4_2;
	wire w_dff_B_IqpecuSu4_2;
	wire w_dff_B_kboR52OL5_2;
	wire w_dff_B_K1SfeoQm6_2;
	wire w_dff_B_UZ6rPx319_2;
	wire w_dff_B_jldKp3rJ3_2;
	wire w_dff_B_VMT8lu7f3_2;
	wire w_dff_B_koqA6MUA1_2;
	wire w_dff_B_EKJKSklJ0_2;
	wire w_dff_B_Tadc9CTp4_2;
	wire w_dff_B_9U5ceWEf9_2;
	wire w_dff_B_bdaHPO2g3_2;
	wire w_dff_B_5SFXbCKm4_2;
	wire w_dff_B_vjaOVjhX4_2;
	wire w_dff_B_tndIYSkn6_2;
	wire w_dff_B_eYQBbDY71_2;
	wire w_dff_B_KfRiBqqk7_2;
	wire w_dff_B_sVUntn618_2;
	wire w_dff_B_5E0S7Mk61_2;
	wire w_dff_B_AkPqbWMS6_2;
	wire w_dff_B_T29OzGGi0_2;
	wire w_dff_B_dbHMGxAf7_2;
	wire w_dff_B_VYi3cu8q2_2;
	wire w_dff_B_og7Gg05P5_2;
	wire w_dff_B_nxteRPeU9_2;
	wire w_dff_B_2Q601fps1_2;
	wire w_dff_B_LKcnht060_2;
	wire w_dff_B_mp4znJFi8_2;
	wire w_dff_B_2TX2MUxa8_2;
	wire w_dff_B_ybZWlAH97_2;
	wire w_dff_B_mHMSWxFA9_2;
	wire w_dff_B_o7MXoDFr3_2;
	wire w_dff_B_khC0GNDL1_2;
	wire w_dff_B_fQN4zX1Q9_2;
	wire w_dff_B_d8wm2tPJ1_2;
	wire w_dff_B_mv68vdNy4_1;
	wire w_dff_B_N19jddEL1_2;
	wire w_dff_B_zCSAdxRo9_2;
	wire w_dff_B_k7UHKrmN5_2;
	wire w_dff_B_QO4Wi0rH7_2;
	wire w_dff_B_dlYknYU47_2;
	wire w_dff_B_lf8cTiQT3_2;
	wire w_dff_B_jQKFDVaN3_2;
	wire w_dff_B_819MoxBQ6_2;
	wire w_dff_B_ITXowIf06_2;
	wire w_dff_B_9KJNCrAw7_2;
	wire w_dff_B_ghQBMAJ50_2;
	wire w_dff_B_crOhpl8S4_2;
	wire w_dff_B_DBwlyrH25_2;
	wire w_dff_B_na5gIAp41_2;
	wire w_dff_B_kvE4x7du9_2;
	wire w_dff_B_RrvAzQYm0_2;
	wire w_dff_B_1zxwHV1P6_2;
	wire w_dff_B_C2CwjGL09_2;
	wire w_dff_B_omL9CEEb8_2;
	wire w_dff_B_Wv9QBvxG9_2;
	wire w_dff_B_86qSjaqv5_2;
	wire w_dff_B_a2EivDk55_2;
	wire w_dff_B_2wwv2AWA8_2;
	wire w_dff_B_zgBzSHyD9_2;
	wire w_dff_B_OmoqOIOh3_2;
	wire w_dff_B_aVGXOIuJ0_2;
	wire w_dff_B_mn1lX62U7_2;
	wire w_dff_B_3Yt60LoN1_2;
	wire w_dff_B_zSuTzn4U3_2;
	wire w_dff_B_7qrznLfw0_2;
	wire w_dff_B_803htx507_2;
	wire w_dff_B_rVW0ikC74_2;
	wire w_dff_B_Yl3UZDtS0_2;
	wire w_dff_B_mhXbmUcO0_2;
	wire w_dff_B_RZrP3vIZ0_1;
	wire w_dff_B_emabwrZH3_2;
	wire w_dff_B_ih9tL02v4_2;
	wire w_dff_B_8LfxJpnY3_2;
	wire w_dff_B_UnvWLgoe4_2;
	wire w_dff_B_sXLHwsOj3_2;
	wire w_dff_B_fJ4Ys15I5_2;
	wire w_dff_B_4E0A09X87_2;
	wire w_dff_B_mEMRNyYs0_2;
	wire w_dff_B_nX6BpL9K7_2;
	wire w_dff_B_kU34mXxB5_2;
	wire w_dff_B_CHH1R1PH1_2;
	wire w_dff_B_Z9Krbvwn0_2;
	wire w_dff_B_6D06yrvc2_2;
	wire w_dff_B_evHTy8lh5_2;
	wire w_dff_B_tzBsdoiJ9_2;
	wire w_dff_B_8R8pBGxB7_2;
	wire w_dff_B_PJHzxGPt8_2;
	wire w_dff_B_nkJlaTvE7_2;
	wire w_dff_B_Dqj2ac0W8_2;
	wire w_dff_B_beOFBzPl8_2;
	wire w_dff_B_PfCkoZLF5_2;
	wire w_dff_B_0vEl2Oyo4_2;
	wire w_dff_B_CXTPmEgr7_2;
	wire w_dff_B_5xyxvJKs0_2;
	wire w_dff_B_rvrh4gJu6_2;
	wire w_dff_B_jIP2ZTtx8_2;
	wire w_dff_B_0MXe75ZF6_2;
	wire w_dff_B_konae6BJ4_2;
	wire w_dff_B_byl4MSlQ5_2;
	wire w_dff_B_0BUPneNN4_2;
	wire w_dff_B_rid0auL54_2;
	wire w_dff_B_CB0sktN81_1;
	wire w_dff_B_ZuPv0UCP1_2;
	wire w_dff_B_2PhOPdVE6_2;
	wire w_dff_B_eF68Gr4u9_2;
	wire w_dff_B_OgHyAR9h0_2;
	wire w_dff_B_ntxEm7ok8_2;
	wire w_dff_B_Y1pRCgYT7_2;
	wire w_dff_B_RQtvvaoB6_2;
	wire w_dff_B_FWC5jXQF2_2;
	wire w_dff_B_CURFQNWl5_2;
	wire w_dff_B_Zfz6R5ip9_2;
	wire w_dff_B_cI1z6C6B9_2;
	wire w_dff_B_WdR5ugpk1_2;
	wire w_dff_B_5GxzGWHf3_2;
	wire w_dff_B_ioAtN6GD9_2;
	wire w_dff_B_NYbpLxkt9_2;
	wire w_dff_B_vYX7WNda7_2;
	wire w_dff_B_yy1t4VSv5_2;
	wire w_dff_B_BejsI9Wk5_2;
	wire w_dff_B_7JrZ1iPz7_2;
	wire w_dff_B_O86Yp4628_2;
	wire w_dff_B_FBoc3Kks4_2;
	wire w_dff_B_UzydEc451_2;
	wire w_dff_B_790z7C9M9_2;
	wire w_dff_B_4prvWc2y5_2;
	wire w_dff_B_Mgx47BCv9_2;
	wire w_dff_B_otfWY0iH9_2;
	wire w_dff_B_PgAFMw7M5_2;
	wire w_dff_B_guKhFquV9_2;
	wire w_dff_B_euu1EETl5_1;
	wire w_dff_B_140oDg3y9_2;
	wire w_dff_B_IYsYkObq8_2;
	wire w_dff_B_foP3H1gP0_2;
	wire w_dff_B_u7Z2H9ci5_2;
	wire w_dff_B_RznP0vOC0_2;
	wire w_dff_B_IBCdzPW32_2;
	wire w_dff_B_KB20gC9q5_2;
	wire w_dff_B_S5VAJ7gx7_2;
	wire w_dff_B_6ftHPquV8_2;
	wire w_dff_B_Uhkxv0Ek3_2;
	wire w_dff_B_GI15IjLD1_2;
	wire w_dff_B_lIWNvGbD4_2;
	wire w_dff_B_NWq41bgg1_2;
	wire w_dff_B_8yRuhjn20_2;
	wire w_dff_B_Gh9Yabwx6_2;
	wire w_dff_B_PcXjcuxO7_2;
	wire w_dff_B_zjBU6wvI0_2;
	wire w_dff_B_4wCIEq9L2_2;
	wire w_dff_B_OeccjMiK7_2;
	wire w_dff_B_BpxqhOfG3_2;
	wire w_dff_B_UVP3n2FV6_2;
	wire w_dff_B_MHLEkW565_2;
	wire w_dff_B_nxEQdo8F8_2;
	wire w_dff_B_Xeegg63e1_2;
	wire w_dff_B_M7snh6mM0_2;
	wire w_dff_B_80NBw8E22_1;
	wire w_dff_B_gaHa6Ttn8_2;
	wire w_dff_B_2qIe3AW63_2;
	wire w_dff_B_7fImEcFy5_2;
	wire w_dff_B_fUmlFteO5_2;
	wire w_dff_B_Vi6yQiHF6_2;
	wire w_dff_B_2rJ3BzyP8_2;
	wire w_dff_B_QfAQvCrZ5_2;
	wire w_dff_B_HbDuMGaU3_2;
	wire w_dff_B_b6UI1FgC3_2;
	wire w_dff_B_2d1ULuW58_2;
	wire w_dff_B_AAan1nW28_2;
	wire w_dff_B_nEnGV00g8_2;
	wire w_dff_B_XTBEhzw57_2;
	wire w_dff_B_jQLgfyHJ8_2;
	wire w_dff_B_4PbDtGpy8_2;
	wire w_dff_B_61uNtf058_2;
	wire w_dff_B_mV8Jujk52_2;
	wire w_dff_B_VYrb5c288_2;
	wire w_dff_B_dwunB3z69_2;
	wire w_dff_B_WfLAAADk9_2;
	wire w_dff_B_a8fZlPKO3_2;
	wire w_dff_B_cBGvdRqR1_2;
	wire w_dff_B_hEuuqHdi4_1;
	wire w_dff_B_fbvPWilt2_2;
	wire w_dff_B_I5wSJXMr1_2;
	wire w_dff_B_FvnetU492_2;
	wire w_dff_B_vyl0QTHK9_2;
	wire w_dff_B_LfhKWCDh7_2;
	wire w_dff_B_ROchpxLD1_2;
	wire w_dff_B_LJiSSg278_2;
	wire w_dff_B_ZIoIHeRj5_2;
	wire w_dff_B_8uFlPPON6_2;
	wire w_dff_B_OJGwLr494_2;
	wire w_dff_B_ZDhRUGph2_2;
	wire w_dff_B_gN3O8cuC7_2;
	wire w_dff_B_1jTV0hhF5_2;
	wire w_dff_B_8zK6q8DU3_2;
	wire w_dff_B_s2CgjbII3_2;
	wire w_dff_B_9yvpeUFL7_2;
	wire w_dff_B_0OlITHCw5_2;
	wire w_dff_B_DetLcREn6_2;
	wire w_dff_B_i37JVgK58_2;
	wire w_dff_B_X2riWvgE7_1;
	wire w_dff_B_RY9wnxnK4_2;
	wire w_dff_B_Pfpbnudr5_2;
	wire w_dff_B_jQwzLbSu8_2;
	wire w_dff_B_EN54tcqP5_2;
	wire w_dff_B_JLwThOEh0_2;
	wire w_dff_B_OG9oEXUv6_2;
	wire w_dff_B_URsgLQtx1_2;
	wire w_dff_B_nyXakjjf5_2;
	wire w_dff_B_yNLoLpNb1_2;
	wire w_dff_B_BzRJ3EN29_2;
	wire w_dff_B_a9tNjHic7_2;
	wire w_dff_B_bb5Pwi2E8_2;
	wire w_dff_B_eVeuy8Od2_2;
	wire w_dff_B_ZofbYMf14_2;
	wire w_dff_B_ouWBy32k7_2;
	wire w_dff_B_HmOy9gdZ6_2;
	wire w_dff_B_npGZULCR8_1;
	wire w_dff_B_tP8yLYmi3_2;
	wire w_dff_B_KlMpgy0L5_2;
	wire w_dff_B_J4eLG92o3_2;
	wire w_dff_B_eNBPa2Nn4_2;
	wire w_dff_B_CT5KwJnv4_2;
	wire w_dff_B_sXqHW34T9_2;
	wire w_dff_B_cWlML1WQ6_2;
	wire w_dff_B_HcahgT2a9_2;
	wire w_dff_B_u1HP4UEW7_2;
	wire w_dff_B_IKWzQX9x2_2;
	wire w_dff_B_5SQtOB3W8_2;
	wire w_dff_B_eQOmFkzZ5_2;
	wire w_dff_B_fkV0tacZ9_2;
	wire w_dff_B_MhBtpbU40_1;
	wire w_dff_B_AlzyFC0d4_2;
	wire w_dff_B_cAUyq2nS0_2;
	wire w_dff_B_nT4RwkNr1_2;
	wire w_dff_B_4aIHD7BG6_2;
	wire w_dff_B_kkV6g1UX2_2;
	wire w_dff_B_0VdfSvSY1_2;
	wire w_dff_B_D34umgtn8_2;
	wire w_dff_B_CDsU8MiW5_2;
	wire w_dff_B_3jElJUyu7_2;
	wire w_dff_B_s9XxNWqf5_2;
	wire w_dff_B_L38jzCHb3_2;
	wire w_dff_B_hvejbr7D5_1;
	wire w_dff_B_sKjMvSKJ5_2;
	wire w_dff_B_F3xIrhsK2_2;
	wire w_dff_B_JQ8vV1Ct7_2;
	wire w_dff_B_mV2s5AHh3_2;
	wire w_dff_B_JJN7KISF6_2;
	wire w_dff_B_lM87nnUQ3_2;
	wire w_dff_B_yrwF1j462_2;
	wire w_dff_B_8DhbLyL88_2;
	wire w_dff_B_h6T7WqZy2_2;
	wire w_dff_B_muOGxhGJ0_2;
	wire w_dff_B_KO48WI7V7_0;
	wire w_dff_A_xjlCJ5fH0_0;
	wire w_dff_A_HYTriE2r8_0;
	wire w_dff_A_X4THlejH0_1;
	wire w_dff_A_y8ecDZvJ4_1;
	wire w_dff_B_ro5cP48Y3_1;
	wire w_dff_B_e9hx0nUu3_2;
	wire w_dff_B_rxRlKeHn5_2;
	wire w_dff_B_m3tKkT4H1_2;
	wire w_dff_B_eojPBsxJ9_2;
	wire w_dff_B_Aw5oXyTs3_2;
	wire w_dff_B_XKXNnmcC7_2;
	wire w_dff_B_Qnxulk1J9_2;
	wire w_dff_B_azXO8WOf0_2;
	wire w_dff_B_x3FjfZDu1_2;
	wire w_dff_B_cHwPmx7o9_2;
	wire w_dff_B_AunaTG8D8_2;
	wire w_dff_B_IqUEvn7s6_2;
	wire w_dff_B_E2NKaZ5a1_2;
	wire w_dff_B_8fH1qxUN0_2;
	wire w_dff_B_AXLrF5O73_2;
	wire w_dff_B_Oi2AIzEE4_2;
	wire w_dff_B_iIs3XRv60_2;
	wire w_dff_B_Tu1j5mQB1_2;
	wire w_dff_B_tnlgnleI5_2;
	wire w_dff_B_XQHYbaeu4_2;
	wire w_dff_B_BLFWJ7ha6_2;
	wire w_dff_B_64pBxwNZ7_2;
	wire w_dff_B_myrIGuL12_2;
	wire w_dff_B_nGXbkOdq6_2;
	wire w_dff_B_oe1UKJlG4_2;
	wire w_dff_B_EF9vJNIh7_2;
	wire w_dff_B_LPAoNBBK6_2;
	wire w_dff_B_HTfnSY413_2;
	wire w_dff_B_xlbU1lKx0_2;
	wire w_dff_B_dGee7S2H7_2;
	wire w_dff_B_hekHXXVp8_2;
	wire w_dff_B_rLR9XlKF9_2;
	wire w_dff_B_vBX8i7zp2_2;
	wire w_dff_B_tf1dHzvh9_2;
	wire w_dff_B_9LZ5ya752_2;
	wire w_dff_B_062t9TBY1_2;
	wire w_dff_B_vdsF2kNk9_2;
	wire w_dff_B_Xc4cmSKZ7_2;
	wire w_dff_B_TUAjzaQc5_2;
	wire w_dff_B_M1cXpTH12_2;
	wire w_dff_B_9ZJrYBGp7_2;
	wire w_dff_B_eP63CA6Z8_2;
	wire w_dff_B_XbFSq7fE1_2;
	wire w_dff_B_IESZAlaq7_2;
	wire w_dff_B_lfyc2Dh14_2;
	wire w_dff_B_KmYUFH5k9_2;
	wire w_dff_B_Ed9BH3408_0;
	wire w_dff_A_zDIQNUSH4_1;
	wire w_dff_B_SwruDX775_1;
	wire w_dff_B_ZFLKPJdI7_2;
	wire w_dff_B_5YUTvlny2_2;
	wire w_dff_B_fVq5IO5Z8_2;
	wire w_dff_B_UFTdSGGb8_2;
	wire w_dff_B_F961kvvd6_2;
	wire w_dff_B_2tsZpQrR7_2;
	wire w_dff_B_3FqGXqHb6_2;
	wire w_dff_B_ukePDoKZ0_2;
	wire w_dff_B_43K46HWJ1_2;
	wire w_dff_B_choCfG798_2;
	wire w_dff_B_HB2ovhRj3_2;
	wire w_dff_B_v5Wb0iHJ4_2;
	wire w_dff_B_tV1mwPZ21_2;
	wire w_dff_B_OqHRrrz13_2;
	wire w_dff_B_9znQpidB3_2;
	wire w_dff_B_8ohYwqSV2_2;
	wire w_dff_B_Bf3ow6S36_2;
	wire w_dff_B_oF1ZgOQ17_2;
	wire w_dff_B_UDrsoCEv9_2;
	wire w_dff_B_7uFdHyHj5_2;
	wire w_dff_B_sSDQfO7u7_2;
	wire w_dff_B_rpZfSjZL3_2;
	wire w_dff_B_BYMxRWhV9_2;
	wire w_dff_B_hQpLa3C88_2;
	wire w_dff_B_eOTUKhrR2_2;
	wire w_dff_B_blWOgusu2_2;
	wire w_dff_B_aTiybGHH9_2;
	wire w_dff_B_FZ0vuZHe8_2;
	wire w_dff_B_igVgbz570_2;
	wire w_dff_B_6tRHFwrC0_2;
	wire w_dff_B_2QzioibU2_2;
	wire w_dff_B_7Lal1JNS0_2;
	wire w_dff_B_cxwcPxIW9_2;
	wire w_dff_B_UQiUkEWc3_2;
	wire w_dff_B_jKip5CG98_2;
	wire w_dff_B_LYtwX1wa1_2;
	wire w_dff_B_EjwOCjkJ8_2;
	wire w_dff_B_P0Z487Ck5_2;
	wire w_dff_B_lCGCcQDY8_2;
	wire w_dff_B_Nzm1NpCa4_2;
	wire w_dff_B_jTp396Bm6_2;
	wire w_dff_B_jfnSrci08_2;
	wire w_dff_B_72didT1E7_1;
	wire w_dff_B_koLmQBVx9_2;
	wire w_dff_B_2NeL1kKh4_2;
	wire w_dff_B_RJ8OZ77n7_2;
	wire w_dff_B_f3WxRuip5_2;
	wire w_dff_B_zUN74IGU2_2;
	wire w_dff_B_Ysqbm8bS8_2;
	wire w_dff_B_91ITMEux7_2;
	wire w_dff_B_sjKZHQDI0_2;
	wire w_dff_B_MxphXzJP0_2;
	wire w_dff_B_AarvnL5V8_2;
	wire w_dff_B_ICokY8lt5_2;
	wire w_dff_B_6Q24a3Lb8_2;
	wire w_dff_B_HZYMmhHe6_2;
	wire w_dff_B_pkwZdyEq5_2;
	wire w_dff_B_xIGQhoHB5_2;
	wire w_dff_B_DZdqauXq5_2;
	wire w_dff_B_CaLWwJJC1_2;
	wire w_dff_B_Wbxpflml8_2;
	wire w_dff_B_WltMCCl04_2;
	wire w_dff_B_YADgxmS45_2;
	wire w_dff_B_AjzUHZIG9_2;
	wire w_dff_B_MD0dnGNm8_2;
	wire w_dff_B_3dZI2tTN6_2;
	wire w_dff_B_ftYZnWzI9_2;
	wire w_dff_B_xd2ONGLZ8_2;
	wire w_dff_B_iZCDyWct0_2;
	wire w_dff_B_1K44OmuI2_2;
	wire w_dff_B_gc9JE6wK9_2;
	wire w_dff_B_XNKZBaDe0_2;
	wire w_dff_B_mJ7nhXEv2_2;
	wire w_dff_B_Avu5dUl02_2;
	wire w_dff_B_eZ9ABUN80_2;
	wire w_dff_B_OlrDENrr0_2;
	wire w_dff_B_PJyKYYJK4_2;
	wire w_dff_B_7vwcqmpR6_2;
	wire w_dff_B_AY4AJOQO3_2;
	wire w_dff_B_b5ywJgcS4_2;
	wire w_dff_B_2Kdu6SYs4_2;
	wire w_dff_B_SkmqDCMx4_2;
	wire w_dff_B_m5BQ8Cor6_1;
	wire w_dff_B_ZFv2DbFa6_2;
	wire w_dff_B_Rgsdhu8z9_2;
	wire w_dff_B_4loedHyv2_2;
	wire w_dff_B_1irYhlm43_2;
	wire w_dff_B_pKp2z2pW6_2;
	wire w_dff_B_4vPUwsJy7_2;
	wire w_dff_B_yW9mvhdH5_2;
	wire w_dff_B_qppZnRYI5_2;
	wire w_dff_B_eFho2Ocr0_2;
	wire w_dff_B_w6IdzP6c3_2;
	wire w_dff_B_eDyzI75j0_2;
	wire w_dff_B_7x8o2d7b2_2;
	wire w_dff_B_FsVR2xqC3_2;
	wire w_dff_B_zdSw8gB36_2;
	wire w_dff_B_x75q6FaY7_2;
	wire w_dff_B_WmuiCPUb9_2;
	wire w_dff_B_dMHStHUJ0_2;
	wire w_dff_B_RF6Zny4U8_2;
	wire w_dff_B_OWYIk00z9_2;
	wire w_dff_B_DKJTnKOe5_2;
	wire w_dff_B_CJJwGijn9_2;
	wire w_dff_B_rkI5szww7_2;
	wire w_dff_B_y0d4yNIv7_2;
	wire w_dff_B_s6rwE94m2_2;
	wire w_dff_B_mSthmGMl1_2;
	wire w_dff_B_dp4bfbII8_2;
	wire w_dff_B_BaRpYuK41_2;
	wire w_dff_B_b6dAJ7fh2_2;
	wire w_dff_B_ppyBh3EC0_2;
	wire w_dff_B_ZUFVAfxQ6_2;
	wire w_dff_B_pHgVYMsK1_2;
	wire w_dff_B_eDzazIj67_2;
	wire w_dff_B_fEp8Xi859_2;
	wire w_dff_B_bhke1jhb5_2;
	wire w_dff_B_Gs5q38Ow6_2;
	wire w_dff_B_Fhg9wTZk4_2;
	wire w_dff_B_uK9k6vOp8_1;
	wire w_dff_B_YT3Oav0l2_2;
	wire w_dff_B_n7VUH4rp0_2;
	wire w_dff_B_tR6z7l7b3_2;
	wire w_dff_B_gRCHUCka2_2;
	wire w_dff_B_kLCdBYPu0_2;
	wire w_dff_B_LLvt2ApK3_2;
	wire w_dff_B_1QCdPEgW0_2;
	wire w_dff_B_EYsZsjDO7_2;
	wire w_dff_B_YuQ7oVd31_2;
	wire w_dff_B_m9rjNFu97_2;
	wire w_dff_B_cUt6OpAC0_2;
	wire w_dff_B_h8geLlOu5_2;
	wire w_dff_B_PHxDSOKU6_2;
	wire w_dff_B_7I1OUmOt6_2;
	wire w_dff_B_LHxuTWIV8_2;
	wire w_dff_B_iyQbVhyw3_2;
	wire w_dff_B_cQcIEMFr0_2;
	wire w_dff_B_hxj5GZfK8_2;
	wire w_dff_B_RuBPVcm53_2;
	wire w_dff_B_n5h6j43O1_2;
	wire w_dff_B_7uNnuhgy3_2;
	wire w_dff_B_vT9CQ6Jv2_2;
	wire w_dff_B_dW60OF9P0_2;
	wire w_dff_B_W35zB9hd0_2;
	wire w_dff_B_QnuR2BcK0_2;
	wire w_dff_B_W7CSpw3n6_2;
	wire w_dff_B_yzpa4i1u6_2;
	wire w_dff_B_mHYYZmXZ5_2;
	wire w_dff_B_w1W6beGH7_2;
	wire w_dff_B_QxvQZhVJ9_2;
	wire w_dff_B_K6alEr3G9_2;
	wire w_dff_B_YzDpsTeH8_2;
	wire w_dff_B_mToJob0I8_2;
	wire w_dff_B_1LktRM5K5_1;
	wire w_dff_B_J6WTWbRu9_2;
	wire w_dff_B_6ZHoQYwV3_2;
	wire w_dff_B_W1xHsh0Y7_2;
	wire w_dff_B_N8Nrvvdr8_2;
	wire w_dff_B_ZgW69Ha32_2;
	wire w_dff_B_966qRKTz0_2;
	wire w_dff_B_yxCLSotg3_2;
	wire w_dff_B_eBvW2OIU5_2;
	wire w_dff_B_fIOEa8zb1_2;
	wire w_dff_B_bWQjhRvE6_2;
	wire w_dff_B_Q2f95jkD5_2;
	wire w_dff_B_AYwitsEW3_2;
	wire w_dff_B_jEKa6cXH1_2;
	wire w_dff_B_TRTSBtWP8_2;
	wire w_dff_B_GXwVtD863_2;
	wire w_dff_B_7606xbX21_2;
	wire w_dff_B_9jlg54Nl8_2;
	wire w_dff_B_7ejpO0pr5_2;
	wire w_dff_B_izIltxwd8_2;
	wire w_dff_B_A6yHRtyG0_2;
	wire w_dff_B_D0Mjjkng0_2;
	wire w_dff_B_IN1IzNOB8_2;
	wire w_dff_B_qhIPU2ky0_2;
	wire w_dff_B_3oXBbsWI7_2;
	wire w_dff_B_YiHYoCaW1_2;
	wire w_dff_B_GsTU2seh5_2;
	wire w_dff_B_UyWPELAZ8_2;
	wire w_dff_B_miABNWeP6_2;
	wire w_dff_B_Y4ySdTZE1_2;
	wire w_dff_B_Y6GAW0cI0_2;
	wire w_dff_B_sCOjvpwk7_1;
	wire w_dff_B_s8t8Y6jC0_2;
	wire w_dff_B_Fjg59sQk4_2;
	wire w_dff_B_NIVnNRD34_2;
	wire w_dff_B_cPctDPIu9_2;
	wire w_dff_B_ZDsRNgsI3_2;
	wire w_dff_B_2kZISSSF4_2;
	wire w_dff_B_GT4L85wp8_2;
	wire w_dff_B_fXI8qcWG4_2;
	wire w_dff_B_3WbCNHrf9_2;
	wire w_dff_B_3a4zULMd1_2;
	wire w_dff_B_SOBtObaT2_2;
	wire w_dff_B_cb9BPlpi5_2;
	wire w_dff_B_mUR7WmDM7_2;
	wire w_dff_B_85fNOHrM6_2;
	wire w_dff_B_d2lSzW5Z7_2;
	wire w_dff_B_XyPOo3FA9_2;
	wire w_dff_B_iW40ZDY95_2;
	wire w_dff_B_OaECFVQW8_2;
	wire w_dff_B_xAsIWQLc4_2;
	wire w_dff_B_68NWWaE34_2;
	wire w_dff_B_c5F9Q2IR2_2;
	wire w_dff_B_9TfUHFVB1_2;
	wire w_dff_B_qaIPyx9p7_2;
	wire w_dff_B_3KuNxgML2_2;
	wire w_dff_B_LBV9gPn63_2;
	wire w_dff_B_YADlhlg21_2;
	wire w_dff_B_hc93bl1r7_2;
	wire w_dff_B_6kM8FJQY9_1;
	wire w_dff_B_ZyzgSRoN8_2;
	wire w_dff_B_OUeqsrJM9_2;
	wire w_dff_B_jkVpC7Dy5_2;
	wire w_dff_B_gkCR23mv0_2;
	wire w_dff_B_WrIzNfP32_2;
	wire w_dff_B_nkJYK7ve5_2;
	wire w_dff_B_hThd8Uot6_2;
	wire w_dff_B_vfo2Y41P6_2;
	wire w_dff_B_qmqbmAq66_2;
	wire w_dff_B_FynjsJbm4_2;
	wire w_dff_B_bsGDJrYI3_2;
	wire w_dff_B_zBBQ3SDi4_2;
	wire w_dff_B_FyKHuwoQ6_2;
	wire w_dff_B_l2R6oesL6_2;
	wire w_dff_B_GoeeFxNv9_2;
	wire w_dff_B_zYinyuAT5_2;
	wire w_dff_B_ZZD9bShk4_2;
	wire w_dff_B_tUCneVk78_2;
	wire w_dff_B_4x9OCzuh4_2;
	wire w_dff_B_wXYqPP6c4_2;
	wire w_dff_B_LCmPTTOE9_2;
	wire w_dff_B_VgGuNdZS4_2;
	wire w_dff_B_WtYEZnw26_2;
	wire w_dff_B_DI2KDhzz3_2;
	wire w_dff_B_i5rvOa3p3_1;
	wire w_dff_B_FGOo59EC6_2;
	wire w_dff_B_0BzU38913_2;
	wire w_dff_B_A9EtvMiB6_2;
	wire w_dff_B_NB5SXZe11_2;
	wire w_dff_B_PxuWLaUL7_2;
	wire w_dff_B_eAv1dQOL5_2;
	wire w_dff_B_R8wxR1fV5_2;
	wire w_dff_B_wlcobMyC5_2;
	wire w_dff_B_DjF9SevS9_2;
	wire w_dff_B_gH3e6Los9_2;
	wire w_dff_B_3MImr5rk7_2;
	wire w_dff_B_niBvErOj2_2;
	wire w_dff_B_uOWDBK3b1_2;
	wire w_dff_B_tEm9qimH6_2;
	wire w_dff_B_0lvyRvPs7_2;
	wire w_dff_B_4nU3qPdF6_2;
	wire w_dff_B_pV06f9Cc4_2;
	wire w_dff_B_YysPbcvA7_2;
	wire w_dff_B_FuojEz9c7_2;
	wire w_dff_B_YF5CjkL67_2;
	wire w_dff_B_XofydX4J3_2;
	wire w_dff_B_cxqTMeGw6_1;
	wire w_dff_B_OYpVKsSp0_2;
	wire w_dff_B_oicXX7277_2;
	wire w_dff_B_r1U5wM4T0_2;
	wire w_dff_B_1dXnuMea1_2;
	wire w_dff_B_CW7tpbTA8_2;
	wire w_dff_B_qay6GDby2_2;
	wire w_dff_B_S5AWkLQn4_2;
	wire w_dff_B_4KoGR2c12_2;
	wire w_dff_B_KtLuIGYF7_2;
	wire w_dff_B_SVOeVH5J3_2;
	wire w_dff_B_RoFIz7MI8_2;
	wire w_dff_B_TvaTr2md3_2;
	wire w_dff_B_lsZc9F6t0_2;
	wire w_dff_B_IxLePcrZ7_2;
	wire w_dff_B_CxQRB3R63_2;
	wire w_dff_B_I7nGwSX22_2;
	wire w_dff_B_1HcQjVsl8_2;
	wire w_dff_B_aKw7mzUM2_2;
	wire w_dff_B_iYHSkoAI3_1;
	wire w_dff_B_Mgft5F382_2;
	wire w_dff_B_G47GsENl3_2;
	wire w_dff_B_VRctDRZy4_2;
	wire w_dff_B_VdiWadEt1_2;
	wire w_dff_B_j5PSWXcg0_2;
	wire w_dff_B_Czwk7QF38_2;
	wire w_dff_B_5hQbSskh1_2;
	wire w_dff_B_f8ff7PKS8_2;
	wire w_dff_B_NvncKvTK9_2;
	wire w_dff_B_OLSWtFCH0_2;
	wire w_dff_B_ECyh6JfX5_2;
	wire w_dff_B_0gSdxCt41_2;
	wire w_dff_B_7UplmbCD0_2;
	wire w_dff_B_MuPLUmnB9_2;
	wire w_dff_B_8FZDh62H1_2;
	wire w_dff_B_LYvvcZlp2_1;
	wire w_dff_B_NHzErvfo8_2;
	wire w_dff_B_Wh6ejkyV2_2;
	wire w_dff_B_e3MUNzrD9_2;
	wire w_dff_B_zEGRgbGm4_2;
	wire w_dff_B_INOngRA77_2;
	wire w_dff_B_KBYuhoZD1_2;
	wire w_dff_B_hPmpx0wQ8_2;
	wire w_dff_B_qT4cfSNC8_2;
	wire w_dff_B_Be6lNEUY1_2;
	wire w_dff_B_G90Oi5jn9_2;
	wire w_dff_B_T7hkcrGP2_2;
	wire w_dff_B_KbVs6OG40_2;
	wire w_dff_B_1Eksn2Zn3_1;
	wire w_dff_B_O5gyWS1I6_2;
	wire w_dff_B_GvOStkZh7_2;
	wire w_dff_B_QsIJ3ucJ6_2;
	wire w_dff_B_4xyshxkA5_2;
	wire w_dff_B_KmlJ57ou0_2;
	wire w_dff_B_n4fHl4XQ7_2;
	wire w_dff_B_V9mFu0RL1_2;
	wire w_dff_B_3M5uY5Tr9_2;
	wire w_dff_B_ZaWpwy740_2;
	wire w_dff_B_RFwDKia83_2;
	wire w_dff_B_mS9zbmyi8_2;
	wire w_dff_B_VbOJDbnY3_1;
	wire w_dff_B_9n09owlS0_1;
	wire w_dff_B_zQnT7X9Y1_2;
	wire w_dff_B_DGmkYPqP0_2;
	wire w_dff_B_E4u52Zoz7_2;
	wire w_dff_B_x2mpqGpk1_0;
	wire w_dff_A_hG4Qr7px8_0;
	wire w_dff_A_nqIjHJqT2_0;
	wire w_dff_A_nHEdJLsC4_1;
	wire w_dff_A_g1Mpap7a6_1;
	wire w_dff_B_9t040d6f3_1;
	wire w_dff_B_Mev7A2tR5_2;
	wire w_dff_B_EeKtMkSW3_2;
	wire w_dff_B_4jql7c3u4_2;
	wire w_dff_B_hntGXt5R9_2;
	wire w_dff_B_CfNg9dQo8_2;
	wire w_dff_B_6jojmauz7_2;
	wire w_dff_B_yxoYTJqx3_2;
	wire w_dff_B_p2NofYur5_2;
	wire w_dff_B_bAzpiuRG6_2;
	wire w_dff_B_5BKnZWRv1_2;
	wire w_dff_B_r05j243Y0_2;
	wire w_dff_B_kobXswfi0_2;
	wire w_dff_B_RSMXxXds7_2;
	wire w_dff_B_YGSifZPw2_2;
	wire w_dff_B_YNwOSMAk9_2;
	wire w_dff_B_NMYcZaMZ6_2;
	wire w_dff_B_l5mBzfNd7_2;
	wire w_dff_B_fu7N1rfx6_2;
	wire w_dff_B_mBDhIcze4_2;
	wire w_dff_B_ISmq8vt38_2;
	wire w_dff_B_uMziZcN20_2;
	wire w_dff_B_HWjKfqSf5_2;
	wire w_dff_B_63Qul5YC3_2;
	wire w_dff_B_vCqWrtgW6_2;
	wire w_dff_B_E1YEEBaE3_2;
	wire w_dff_B_jx82Vfhe2_2;
	wire w_dff_B_2pLYcsUD1_2;
	wire w_dff_B_x2wMZitc2_2;
	wire w_dff_B_X6Ml1W8V8_2;
	wire w_dff_B_MxeULBOb2_2;
	wire w_dff_B_vzCeqZdo9_2;
	wire w_dff_B_j8gJeYrE7_2;
	wire w_dff_B_uNiqXae08_2;
	wire w_dff_B_lgATJXxJ1_2;
	wire w_dff_B_EAoBZrwA9_2;
	wire w_dff_B_TMgvlIA79_2;
	wire w_dff_B_RrR9zis70_2;
	wire w_dff_B_GmA4Vr5K0_2;
	wire w_dff_B_jz4ORJk21_2;
	wire w_dff_B_MO59b8JA7_2;
	wire w_dff_B_skBfKhuI0_2;
	wire w_dff_B_lTImN72h1_2;
	wire w_dff_B_PND3Uvmr6_2;
	wire w_dff_B_KUj90Kln8_2;
	wire w_dff_B_TiBUXKJU4_2;
	wire w_dff_B_JtkMUbzs3_2;
	wire w_dff_B_wztV4xSX0_0;
	wire w_dff_A_s2XrVx6R2_1;
	wire w_dff_B_mwxOl5mb9_1;
	wire w_dff_B_wXRiHMXH9_2;
	wire w_dff_B_a0W6LTZY3_2;
	wire w_dff_B_gnTokJbh4_2;
	wire w_dff_B_buhPrzya7_2;
	wire w_dff_B_qmGOzqXB2_2;
	wire w_dff_B_2Rwtgp866_2;
	wire w_dff_B_oB3l6RXp6_2;
	wire w_dff_B_6TPLTBmE4_2;
	wire w_dff_B_iijzvRKa6_2;
	wire w_dff_B_CDmkz72u0_2;
	wire w_dff_B_L1abFwff6_2;
	wire w_dff_B_jpUODlBj1_2;
	wire w_dff_B_MlXYdS4E5_2;
	wire w_dff_B_zVo3CANZ2_2;
	wire w_dff_B_Y86smOFu3_2;
	wire w_dff_B_1nIuf5JA9_2;
	wire w_dff_B_F8T7Bx9u6_2;
	wire w_dff_B_PBxRXUcp8_2;
	wire w_dff_B_HEp7zFMA7_2;
	wire w_dff_B_dHRQ70XL4_2;
	wire w_dff_B_sxbtVEAB0_2;
	wire w_dff_B_lkfgfxll7_2;
	wire w_dff_B_jEj45JqO5_2;
	wire w_dff_B_twt6vKDL5_2;
	wire w_dff_B_r17X3Flb5_2;
	wire w_dff_B_qpDD8kv18_2;
	wire w_dff_B_5kpM8K1R9_2;
	wire w_dff_B_J7dseuea3_2;
	wire w_dff_B_6DoHxmma1_2;
	wire w_dff_B_1RVTBdNJ0_2;
	wire w_dff_B_JE9RxYM24_2;
	wire w_dff_B_dmxwLxfi2_2;
	wire w_dff_B_V5VCLTH43_2;
	wire w_dff_B_a4osvAmc2_2;
	wire w_dff_B_N6AHXkbF5_2;
	wire w_dff_B_O0JhIPw07_2;
	wire w_dff_B_DQHEeKIw4_2;
	wire w_dff_B_kcsrwiPU6_2;
	wire w_dff_B_L6Rp2KA26_2;
	wire w_dff_B_npZRYyU75_2;
	wire w_dff_B_tdWHgp7n9_2;
	wire w_dff_B_wuiWfaLW9_2;
	wire w_dff_B_zcHUBgZ90_1;
	wire w_dff_B_8LFVjVyH9_2;
	wire w_dff_B_DpDWqd1R9_2;
	wire w_dff_B_FUWQD5aA9_2;
	wire w_dff_B_CMDEz6jy6_2;
	wire w_dff_B_o4Qq07tr2_2;
	wire w_dff_B_pXFwTl3J0_2;
	wire w_dff_B_SMUDMK8o4_2;
	wire w_dff_B_tYZcWdYQ0_2;
	wire w_dff_B_gcYlqGOP8_2;
	wire w_dff_B_rZoHJuAq7_2;
	wire w_dff_B_GdxRIVTI6_2;
	wire w_dff_B_wXGjJxQu8_2;
	wire w_dff_B_Z2TGY7Zb5_2;
	wire w_dff_B_dQJOBsL50_2;
	wire w_dff_B_Hwl65rLE5_2;
	wire w_dff_B_iDhMGPT26_2;
	wire w_dff_B_TH1ZTvff4_2;
	wire w_dff_B_MIcxA2Vq0_2;
	wire w_dff_B_1gE1HjZl2_2;
	wire w_dff_B_Cynb3zst0_2;
	wire w_dff_B_YIwcJRkS7_2;
	wire w_dff_B_gzp6AcP23_2;
	wire w_dff_B_GyGQnDmy6_2;
	wire w_dff_B_Cpaa194s9_2;
	wire w_dff_B_Vscg8Jay6_2;
	wire w_dff_B_vZUcsHqd7_2;
	wire w_dff_B_4PeIBbgi5_2;
	wire w_dff_B_a4f51BJZ3_2;
	wire w_dff_B_EJUCWQe28_2;
	wire w_dff_B_0e1C559U2_2;
	wire w_dff_B_AdZfayq25_2;
	wire w_dff_B_tfuUpwKE0_2;
	wire w_dff_B_2vbQGTsJ6_2;
	wire w_dff_B_VZssfK2X6_2;
	wire w_dff_B_R6LeE3Ft7_2;
	wire w_dff_B_bljc86PX1_2;
	wire w_dff_B_K8JRXiRX2_2;
	wire w_dff_B_lW0kk8354_2;
	wire w_dff_B_mbhr9m1M1_2;
	wire w_dff_B_lqFfUgs60_1;
	wire w_dff_B_KBeKWEJB4_2;
	wire w_dff_B_JyfXNeKL5_2;
	wire w_dff_B_qEnCukdO6_2;
	wire w_dff_B_W2Rurbls0_2;
	wire w_dff_B_cjfsOv1y8_2;
	wire w_dff_B_qV1g9Prs5_2;
	wire w_dff_B_ONi6J01R7_2;
	wire w_dff_B_HniIYiJL6_2;
	wire w_dff_B_Jmj5DSi88_2;
	wire w_dff_B_dHbY1vWt0_2;
	wire w_dff_B_wl19Ld9m2_2;
	wire w_dff_B_85UvMXL87_2;
	wire w_dff_B_k3iX4E0i5_2;
	wire w_dff_B_Caezq4bY2_2;
	wire w_dff_B_YQrebjQp4_2;
	wire w_dff_B_QuE9XNyK1_2;
	wire w_dff_B_I6lkS5e53_2;
	wire w_dff_B_AWynAbvu6_2;
	wire w_dff_B_hgs86rlD8_2;
	wire w_dff_B_vgPhUIB04_2;
	wire w_dff_B_riKux56G7_2;
	wire w_dff_B_bUr5vGjO8_2;
	wire w_dff_B_M86Ho1Bm1_2;
	wire w_dff_B_m5GmsNR90_2;
	wire w_dff_B_bL3vy8Vl6_2;
	wire w_dff_B_m2sC1NEV4_2;
	wire w_dff_B_1jNKTHhZ1_2;
	wire w_dff_B_llysxnyL1_2;
	wire w_dff_B_Lq9rmOH56_2;
	wire w_dff_B_W4zzFZB87_2;
	wire w_dff_B_AFp6Rvfp9_2;
	wire w_dff_B_sJztinWD0_2;
	wire w_dff_B_HKctigfB6_2;
	wire w_dff_B_GTtQcLjM1_2;
	wire w_dff_B_1yz24uV28_2;
	wire w_dff_B_FRdNxege6_2;
	wire w_dff_B_1MmuV6Vb7_1;
	wire w_dff_B_2qajahL00_2;
	wire w_dff_B_zx5zGZ3z5_2;
	wire w_dff_B_qkXnfkjC3_2;
	wire w_dff_B_QW1dHc2r4_2;
	wire w_dff_B_qXvLha4E2_2;
	wire w_dff_B_VeBiJPly0_2;
	wire w_dff_B_QhKmzk4d2_2;
	wire w_dff_B_xf8nfrmz8_2;
	wire w_dff_B_Amj9SR2e0_2;
	wire w_dff_B_yQXeHfFn3_2;
	wire w_dff_B_3YCtFFb71_2;
	wire w_dff_B_4i5y2rlA0_2;
	wire w_dff_B_FzeFKLdv1_2;
	wire w_dff_B_9fHz8tE97_2;
	wire w_dff_B_kmk8lekL2_2;
	wire w_dff_B_3SClmbQ98_2;
	wire w_dff_B_xAnIGToR2_2;
	wire w_dff_B_Qlcq6qvH2_2;
	wire w_dff_B_s477KKrP8_2;
	wire w_dff_B_qKTptbSZ1_2;
	wire w_dff_B_WlarPdLD0_2;
	wire w_dff_B_45KLFwQS7_2;
	wire w_dff_B_TUyAwlTn3_2;
	wire w_dff_B_b5ylFTOj4_2;
	wire w_dff_B_l91dVKwJ7_2;
	wire w_dff_B_96RTggfs1_2;
	wire w_dff_B_0qOC2W1v2_2;
	wire w_dff_B_NuO0l4nZ5_2;
	wire w_dff_B_TBfQyYoT1_2;
	wire w_dff_B_39pfXZz19_2;
	wire w_dff_B_8bu60b5c9_2;
	wire w_dff_B_61PhXr827_2;
	wire w_dff_B_gQfjdZlo5_2;
	wire w_dff_B_Gsa8nd0s8_1;
	wire w_dff_B_afuhBzha9_2;
	wire w_dff_B_WtZzsr5W8_2;
	wire w_dff_B_Wwc8q2Rw4_2;
	wire w_dff_B_q5QB4lUo2_2;
	wire w_dff_B_swaUDdSF0_2;
	wire w_dff_B_qDYt7nbd2_2;
	wire w_dff_B_2qTqRvlW3_2;
	wire w_dff_B_vRuBQgIE4_2;
	wire w_dff_B_C6nCEh9i5_2;
	wire w_dff_B_pMm4pkmh7_2;
	wire w_dff_B_5I2ou4L92_2;
	wire w_dff_B_dUH4GDyX4_2;
	wire w_dff_B_kTw7f4GD7_2;
	wire w_dff_B_mdN2fhrM6_2;
	wire w_dff_B_mYzYfili8_2;
	wire w_dff_B_CfP76dGT1_2;
	wire w_dff_B_EYDedzUd4_2;
	wire w_dff_B_PSKzpbiE1_2;
	wire w_dff_B_z7sC5bZP5_2;
	wire w_dff_B_UEuPTdyw1_2;
	wire w_dff_B_fwIPDdqK3_2;
	wire w_dff_B_UnrrENxU3_2;
	wire w_dff_B_wzpjEvUe5_2;
	wire w_dff_B_SqVhbY4B1_2;
	wire w_dff_B_KhvejIkn0_2;
	wire w_dff_B_rWSS7VCu7_2;
	wire w_dff_B_RNsonPTE1_2;
	wire w_dff_B_hs2zLa393_2;
	wire w_dff_B_kzrcoXMJ4_2;
	wire w_dff_B_agDZGcgb0_2;
	wire w_dff_B_KmONAJPs5_1;
	wire w_dff_B_9C3wDcnH7_2;
	wire w_dff_B_aYjU6GZ77_2;
	wire w_dff_B_dAQ4DXwb0_2;
	wire w_dff_B_GXnwgz5D6_2;
	wire w_dff_B_wSezUTmB8_2;
	wire w_dff_B_A9Q1NYPP4_2;
	wire w_dff_B_xn9GcnWh8_2;
	wire w_dff_B_9j13FQdz2_2;
	wire w_dff_B_7t34lPtK3_2;
	wire w_dff_B_Kagtc9w50_2;
	wire w_dff_B_H29SMceJ4_2;
	wire w_dff_B_QuDqRJX72_2;
	wire w_dff_B_FKa6rfTr3_2;
	wire w_dff_B_gM8mhMaM2_2;
	wire w_dff_B_D6if3GDK8_2;
	wire w_dff_B_k2LfXZY65_2;
	wire w_dff_B_ff1Wecaz5_2;
	wire w_dff_B_BHTOasWb7_2;
	wire w_dff_B_wdD4OTvt7_2;
	wire w_dff_B_3AAbsJM04_2;
	wire w_dff_B_IklaTZij1_2;
	wire w_dff_B_wtlmhCxI6_2;
	wire w_dff_B_mwhgo5Sm6_2;
	wire w_dff_B_0BakiQWU6_2;
	wire w_dff_B_QJHueJYm9_2;
	wire w_dff_B_bqaJiNvs7_2;
	wire w_dff_B_X5KODBcQ8_2;
	wire w_dff_B_Fm64XX5H4_1;
	wire w_dff_B_oOHcAjoA9_2;
	wire w_dff_B_esaunbSb6_2;
	wire w_dff_B_UC16XmCD7_2;
	wire w_dff_B_GPgHBzW92_2;
	wire w_dff_B_QC8QxRYn7_2;
	wire w_dff_B_7PczbEzD1_2;
	wire w_dff_B_KjjvChe66_2;
	wire w_dff_B_qy9ut7mM2_2;
	wire w_dff_B_pVfqf9br4_2;
	wire w_dff_B_Olcqf9OU1_2;
	wire w_dff_B_wxZsCW0Z7_2;
	wire w_dff_B_Tem6Ds3i6_2;
	wire w_dff_B_JpKp5glT1_2;
	wire w_dff_B_CXmYz1ss1_2;
	wire w_dff_B_yOXM7FSi1_2;
	wire w_dff_B_fyk4inXr3_2;
	wire w_dff_B_uUhqt12A2_2;
	wire w_dff_B_l6TdmEOG4_2;
	wire w_dff_B_ipyvXdGK8_2;
	wire w_dff_B_FtuwAEjf2_2;
	wire w_dff_B_a9QQZFrk2_2;
	wire w_dff_B_3dB2SyH27_2;
	wire w_dff_B_ezzIuTk95_2;
	wire w_dff_B_5zjqFYag2_2;
	wire w_dff_B_8U4bRvfp3_1;
	wire w_dff_B_2KzRaxmx7_2;
	wire w_dff_B_9DUP62Jz3_2;
	wire w_dff_B_D9gNovTs7_2;
	wire w_dff_B_OdEG0UGN2_2;
	wire w_dff_B_XXCYUZkq1_2;
	wire w_dff_B_AiygU9vh8_2;
	wire w_dff_B_dxEzX2fk8_2;
	wire w_dff_B_fpa3Njoi2_2;
	wire w_dff_B_A3IYaeHX9_2;
	wire w_dff_B_AY4zyO7d9_2;
	wire w_dff_B_EjldRlN04_2;
	wire w_dff_B_O1AGV8Mj5_2;
	wire w_dff_B_01r305D21_2;
	wire w_dff_B_z4b6ezLd9_2;
	wire w_dff_B_O6uKpGyC9_2;
	wire w_dff_B_lJItwmgE8_2;
	wire w_dff_B_mQKObdEv8_2;
	wire w_dff_B_s691kwsS4_2;
	wire w_dff_B_ZaMaxq0z2_2;
	wire w_dff_B_Az5yo4cW8_2;
	wire w_dff_B_kPyJZvli6_2;
	wire w_dff_B_GuYSHLCf0_1;
	wire w_dff_B_mUclxpru7_2;
	wire w_dff_B_UqD2P0ku7_2;
	wire w_dff_B_jYBafdmq0_2;
	wire w_dff_B_Bqc89Xmn6_2;
	wire w_dff_B_velkgLsM1_2;
	wire w_dff_B_RKygZ9z57_2;
	wire w_dff_B_jRMC4n5K0_2;
	wire w_dff_B_j4n2Vfjf3_2;
	wire w_dff_B_KEqbxZAs4_2;
	wire w_dff_B_ThCaaDeO8_2;
	wire w_dff_B_2mKLQ3yo5_2;
	wire w_dff_B_vFPDQEYe6_2;
	wire w_dff_B_wHyZ3VmD0_2;
	wire w_dff_B_59OiT60s9_2;
	wire w_dff_B_o5MepG8Q6_2;
	wire w_dff_B_fiHQYdtG8_2;
	wire w_dff_B_e8OA1mjm3_2;
	wire w_dff_B_1fONnGMT0_2;
	wire w_dff_B_TyaiXiWX8_1;
	wire w_dff_B_kSAGYTcu8_2;
	wire w_dff_B_l915hsfN1_2;
	wire w_dff_B_7iAyFHPN8_2;
	wire w_dff_B_jVYgW8v39_2;
	wire w_dff_B_PkLk4g3a4_2;
	wire w_dff_B_r7RM0ham1_2;
	wire w_dff_B_hW1pG5ih6_2;
	wire w_dff_B_lK6Ho6Lu3_2;
	wire w_dff_B_69YT2YFB1_2;
	wire w_dff_B_uJdAzTQq5_2;
	wire w_dff_B_dwCyvl3u9_2;
	wire w_dff_B_puXUq43Z6_2;
	wire w_dff_B_VdZ7G18k2_2;
	wire w_dff_B_cutxkZDZ0_2;
	wire w_dff_B_1OLi2jHj4_2;
	wire w_dff_B_HLJpNWGj5_1;
	wire w_dff_B_mHi4H4Ha4_2;
	wire w_dff_B_oaIatHEk3_2;
	wire w_dff_B_A3pP1mEA4_2;
	wire w_dff_B_wb9IMQ4a4_2;
	wire w_dff_B_7wzD5FRp2_2;
	wire w_dff_B_e1HZEEES3_2;
	wire w_dff_B_GK9OsL6K1_2;
	wire w_dff_B_9NE4ZEbF7_2;
	wire w_dff_B_RYKPiDi66_2;
	wire w_dff_B_NtiND1tn5_2;
	wire w_dff_B_CtZDk9d71_2;
	wire w_dff_B_uXYkKBb94_2;
	wire w_dff_B_sfcCpwer7_1;
	wire w_dff_B_cwChgFb36_2;
	wire w_dff_B_2jW0S4wf9_2;
	wire w_dff_B_4KFNpsED5_2;
	wire w_dff_B_2THOlbMO2_2;
	wire w_dff_B_C8F8gtl95_2;
	wire w_dff_B_LMTNzjtw9_2;
	wire w_dff_B_XpVCeBoh5_2;
	wire w_dff_B_JDMQXHZZ1_2;
	wire w_dff_B_Q5RmVBP66_2;
	wire w_dff_B_jSyAlbkI4_2;
	wire w_dff_B_CHBlmuDm5_2;
	wire w_dff_B_3wmnwqtf4_1;
	wire w_dff_B_jCZ6uKDN9_1;
	wire w_dff_B_vIMy7gBQ4_2;
	wire w_dff_B_kJvLCQcI9_2;
	wire w_dff_B_zDriRcux5_2;
	wire w_dff_B_pnrgftmm8_0;
	wire w_dff_A_YpcDgDI45_0;
	wire w_dff_A_DeY9akHJ1_0;
	wire w_dff_A_6dRNXfir4_1;
	wire w_dff_A_ae8Leg8q5_1;
	wire w_dff_B_5UjToAl94_2;
	wire w_dff_B_SP1HpvoC3_1;
	wire w_dff_B_71cK37nZ6_2;
	wire w_dff_B_YK0SbFRt6_2;
	wire w_dff_B_l9SbmwhF0_2;
	wire w_dff_B_jRxX2vNX1_2;
	wire w_dff_B_TXHHwfc74_2;
	wire w_dff_B_VPUXu7tS8_2;
	wire w_dff_B_P3CeeXQm7_2;
	wire w_dff_B_o9V35KRA9_2;
	wire w_dff_B_nh9s3tTn1_2;
	wire w_dff_B_vSbYCo453_2;
	wire w_dff_B_e9QocAal7_2;
	wire w_dff_B_wgWsdMIV8_2;
	wire w_dff_B_DAbkcINL6_2;
	wire w_dff_B_8x9jV9B98_2;
	wire w_dff_B_G5xoHGjX5_2;
	wire w_dff_B_mjikOwLC7_2;
	wire w_dff_B_u8zQrG3z9_2;
	wire w_dff_B_ZggIJJAC3_2;
	wire w_dff_B_WvfaBn5O1_2;
	wire w_dff_B_zqQtchwe3_2;
	wire w_dff_B_IXOXLDQa0_2;
	wire w_dff_B_R41Ituzw7_2;
	wire w_dff_B_e92hMknu6_2;
	wire w_dff_B_0ZkeI9lZ3_2;
	wire w_dff_B_tuLgRq3u5_2;
	wire w_dff_B_EM5gG7WT6_2;
	wire w_dff_B_2bCPBpfY4_2;
	wire w_dff_B_rFemxtgI9_2;
	wire w_dff_B_TE82Mu566_2;
	wire w_dff_B_YNoogsYC9_2;
	wire w_dff_B_DEJEUtwu3_2;
	wire w_dff_B_Qnw7XuIt0_2;
	wire w_dff_B_Djj2TcPL3_2;
	wire w_dff_B_bKHsVbBg8_2;
	wire w_dff_B_NV0MGv9q6_2;
	wire w_dff_B_kDOhS67u4_2;
	wire w_dff_B_TLj0vM5f8_2;
	wire w_dff_B_dWYwdqNx2_2;
	wire w_dff_B_lljg9htH9_2;
	wire w_dff_B_few84Wq91_2;
	wire w_dff_B_0eo0p8Kg9_2;
	wire w_dff_B_MI4lqtHn0_2;
	wire w_dff_B_ykau3p4K6_2;
	wire w_dff_B_Mk0TUSzN9_2;
	wire w_dff_B_zOpO2JFm7_2;
	wire w_dff_B_sg5RzDjZ8_2;
	wire w_dff_B_ZnchbZUI3_1;
	wire w_dff_B_wdAMPoaF0_2;
	wire w_dff_B_5URAdbae0_2;
	wire w_dff_B_2wvz0KpW4_2;
	wire w_dff_B_BClbjmIh3_2;
	wire w_dff_B_3RZ21tG67_2;
	wire w_dff_B_wRwX9GTn0_2;
	wire w_dff_B_CeA2Fwuc8_2;
	wire w_dff_B_wQ4XOuxH8_2;
	wire w_dff_B_MgCTk6jI1_2;
	wire w_dff_B_w5cP2fYv4_2;
	wire w_dff_B_UDIBngJ91_2;
	wire w_dff_B_bqyMLTma7_2;
	wire w_dff_B_AdknMspm5_2;
	wire w_dff_B_1tY35QHh3_2;
	wire w_dff_B_oxchOEEt4_2;
	wire w_dff_B_64Cmum3t4_2;
	wire w_dff_B_fzBkggOH7_2;
	wire w_dff_B_aHIko8rw1_2;
	wire w_dff_B_cSpqfCL07_2;
	wire w_dff_B_Kd4jgXSm8_2;
	wire w_dff_B_moHWxap25_2;
	wire w_dff_B_RRltPjFi3_2;
	wire w_dff_B_5wKUrzf65_2;
	wire w_dff_B_dGSAcWoX4_2;
	wire w_dff_B_jsmUPEP30_2;
	wire w_dff_B_fv9hfoGt9_2;
	wire w_dff_B_5FZSmRek4_2;
	wire w_dff_B_mjx9Eo4e7_2;
	wire w_dff_B_rUwZoaS78_2;
	wire w_dff_B_D0lFcWPB5_2;
	wire w_dff_B_NjQMJKnR7_2;
	wire w_dff_B_X9DVy4Qx8_2;
	wire w_dff_B_0XLoYU5T4_2;
	wire w_dff_B_Vp3ifSjy0_2;
	wire w_dff_B_okLpPXzQ2_2;
	wire w_dff_B_xCEpiB3p3_2;
	wire w_dff_B_hH3DvJTQ0_2;
	wire w_dff_B_umnE4FMY2_2;
	wire w_dff_B_dmCv4WHx8_2;
	wire w_dff_B_45YYGLI79_2;
	wire w_dff_B_qf6KaGu87_2;
	wire w_dff_B_f5jzpFwY9_2;
	wire w_dff_B_CrfapjXi1_1;
	wire w_dff_B_V69YQsqG4_2;
	wire w_dff_B_6UawjIrV5_2;
	wire w_dff_B_EDDUXb4S1_2;
	wire w_dff_B_ud80M0vy1_2;
	wire w_dff_B_mXgA2FpI4_2;
	wire w_dff_B_09ygmIav2_2;
	wire w_dff_B_Auv3TVh96_2;
	wire w_dff_B_Xi8lea3v9_2;
	wire w_dff_B_BGrSYvj22_2;
	wire w_dff_B_F8gJViX73_2;
	wire w_dff_B_dMF2Ni9S0_2;
	wire w_dff_B_2HGrpTvm3_2;
	wire w_dff_B_Z94lnMzP8_2;
	wire w_dff_B_CGHP00si3_2;
	wire w_dff_B_4raPXYEk1_2;
	wire w_dff_B_RJ5hshh29_2;
	wire w_dff_B_vtNaouEg7_2;
	wire w_dff_B_28g9tOFh2_2;
	wire w_dff_B_FKJ3wFMO7_2;
	wire w_dff_B_prSK7DWw7_2;
	wire w_dff_B_BCAdCdye2_2;
	wire w_dff_B_Q8ulPfxt9_2;
	wire w_dff_B_bHpKbI9B6_2;
	wire w_dff_B_K5ju37lr5_2;
	wire w_dff_B_229QCfxt9_2;
	wire w_dff_B_7v78ovQT2_2;
	wire w_dff_B_JsVFV5wz2_2;
	wire w_dff_B_SdNBurqI6_2;
	wire w_dff_B_pODrh9r59_2;
	wire w_dff_B_7zxmP5Zr7_2;
	wire w_dff_B_x2Z4l0kg9_2;
	wire w_dff_B_jLFTsBHk6_2;
	wire w_dff_B_9D1WOhjy7_2;
	wire w_dff_B_WFLJ8JVs3_2;
	wire w_dff_B_z7olk5Sa9_2;
	wire w_dff_B_pGQqjV7U0_2;
	wire w_dff_B_0hNEUiv10_2;
	wire w_dff_B_ooaUOpmP9_2;
	wire w_dff_B_y0v4w9nr6_2;
	wire w_dff_B_m02Mw1jm9_1;
	wire w_dff_B_cxFXrJTS5_2;
	wire w_dff_B_kqS5ULAi3_2;
	wire w_dff_B_2yRIJCt79_2;
	wire w_dff_B_2zxAJRTr3_2;
	wire w_dff_B_WwHnwgwd0_2;
	wire w_dff_B_SuE322iB6_2;
	wire w_dff_B_9dmu7QGB2_2;
	wire w_dff_B_mLpTjJZh3_2;
	wire w_dff_B_w0Tf9ODh6_2;
	wire w_dff_B_UFDaTRqW1_2;
	wire w_dff_B_UYGEtdvl5_2;
	wire w_dff_B_x2XSTL6S0_2;
	wire w_dff_B_QiZuaDGp4_2;
	wire w_dff_B_3UsTOzIP5_2;
	wire w_dff_B_5P9KJta54_2;
	wire w_dff_B_v9sYggrd1_2;
	wire w_dff_B_Ssl33oJn0_2;
	wire w_dff_B_U1WXKmK53_2;
	wire w_dff_B_wuZPX3pd1_2;
	wire w_dff_B_HGWXxLhB5_2;
	wire w_dff_B_paDfDDmw0_2;
	wire w_dff_B_6GFn8D1V1_2;
	wire w_dff_B_tL76Uq5V2_2;
	wire w_dff_B_cGjkux6G4_2;
	wire w_dff_B_mi4VUHIQ2_2;
	wire w_dff_B_ZMfxlqyd3_2;
	wire w_dff_B_iYhExfym0_2;
	wire w_dff_B_wiwxmdGk2_2;
	wire w_dff_B_2WCuw5mT3_2;
	wire w_dff_B_Tb1vvtYi2_2;
	wire w_dff_B_Ixm0xFCO7_2;
	wire w_dff_B_GR8kSYNR7_2;
	wire w_dff_B_5Vy1W1Gf9_2;
	wire w_dff_B_6uS1MzVD9_2;
	wire w_dff_B_FlcmKFLv6_2;
	wire w_dff_B_9zXT8tMX6_2;
	wire w_dff_B_g8XKJVFw3_1;
	wire w_dff_B_79xcPeQN5_2;
	wire w_dff_B_NVgzO3NF1_2;
	wire w_dff_B_XFdAogwm4_2;
	wire w_dff_B_FtAlXc7k3_2;
	wire w_dff_B_3wdPJEmg0_2;
	wire w_dff_B_dcIfVtK90_2;
	wire w_dff_B_Zuw9jU3M8_2;
	wire w_dff_B_AmqrlRJz0_2;
	wire w_dff_B_3ZkWtzQX2_2;
	wire w_dff_B_Kx9IwpM71_2;
	wire w_dff_B_HUmgC5bV4_2;
	wire w_dff_B_8zupik028_2;
	wire w_dff_B_lKR91fiW8_2;
	wire w_dff_B_gmCZ4vL74_2;
	wire w_dff_B_jd2WnOjq9_2;
	wire w_dff_B_ZiTPcUyT7_2;
	wire w_dff_B_UsvavLb55_2;
	wire w_dff_B_63O8CR9r1_2;
	wire w_dff_B_iNrKj0ju9_2;
	wire w_dff_B_rwpmIUYj5_2;
	wire w_dff_B_ak1xBx2U8_2;
	wire w_dff_B_xA4YWT8C0_2;
	wire w_dff_B_K77LXZyO8_2;
	wire w_dff_B_o72rBbEI4_2;
	wire w_dff_B_Mymlih731_2;
	wire w_dff_B_t1oPpmXf2_2;
	wire w_dff_B_vSj4aknc2_2;
	wire w_dff_B_lluLUQWV3_2;
	wire w_dff_B_AKMhD39Q0_2;
	wire w_dff_B_Yp1yWMb26_2;
	wire w_dff_B_5Zfa1MZy7_2;
	wire w_dff_B_DoOjH9fV8_2;
	wire w_dff_B_krZPfOzy8_2;
	wire w_dff_B_DgelcY9s0_1;
	wire w_dff_B_n2wlbCTp3_2;
	wire w_dff_B_iV9qx05D7_2;
	wire w_dff_B_va4LksZJ6_2;
	wire w_dff_B_wLd8OlM61_2;
	wire w_dff_B_8Tk36hCG3_2;
	wire w_dff_B_WSdfvYBY5_2;
	wire w_dff_B_m0ZDxtK81_2;
	wire w_dff_B_lkPEqwj77_2;
	wire w_dff_B_KC6Jr47j8_2;
	wire w_dff_B_lwgW2GI17_2;
	wire w_dff_B_I0V4xDrm2_2;
	wire w_dff_B_IetvA6Mi8_2;
	wire w_dff_B_Iwr3XN9U5_2;
	wire w_dff_B_6RMFK7qw7_2;
	wire w_dff_B_iVQFYlep3_2;
	wire w_dff_B_vmfQfqnN2_2;
	wire w_dff_B_Icnrj4Bo2_2;
	wire w_dff_B_johYvclZ3_2;
	wire w_dff_B_s4nzUCk26_2;
	wire w_dff_B_od5SsdDx4_2;
	wire w_dff_B_ok7elgaY6_2;
	wire w_dff_B_fB6TQAIy2_2;
	wire w_dff_B_IVfJyvYH3_2;
	wire w_dff_B_KFP4rjqn8_2;
	wire w_dff_B_VvkALyYG6_2;
	wire w_dff_B_4nNpd3uk5_2;
	wire w_dff_B_3p8Vyoyk6_2;
	wire w_dff_B_ixf2x6Qq0_2;
	wire w_dff_B_udHESU6A9_2;
	wire w_dff_B_wqiKM8GG9_2;
	wire w_dff_B_gdrGJvfb5_1;
	wire w_dff_B_6LAxITUM1_2;
	wire w_dff_B_wqR3q3tK0_2;
	wire w_dff_B_x46Z4r6u8_2;
	wire w_dff_B_bZT47peb1_2;
	wire w_dff_B_bRNfpkxY2_2;
	wire w_dff_B_2IO2lG6n8_2;
	wire w_dff_B_holTAT613_2;
	wire w_dff_B_mhZVSbhS8_2;
	wire w_dff_B_EL0OK4th6_2;
	wire w_dff_B_wZD3fL640_2;
	wire w_dff_B_OA5ufeU86_2;
	wire w_dff_B_6XBoNMvw5_2;
	wire w_dff_B_GNbxkuDy3_2;
	wire w_dff_B_aHllh0UQ8_2;
	wire w_dff_B_ORPEDbGn2_2;
	wire w_dff_B_0LQUf4Ah5_2;
	wire w_dff_B_6JmgZ9PH7_2;
	wire w_dff_B_He58tmNP8_2;
	wire w_dff_B_PrL1D6tf4_2;
	wire w_dff_B_aZCe5bF60_2;
	wire w_dff_B_Ueu599mm7_2;
	wire w_dff_B_RHUtLhne3_2;
	wire w_dff_B_M4GdUuWq6_2;
	wire w_dff_B_VZqh0cDT6_2;
	wire w_dff_B_IhLGXj228_2;
	wire w_dff_B_lGtpcAJp7_2;
	wire w_dff_B_03qnLCe22_2;
	wire w_dff_B_hbAs9MRE7_1;
	wire w_dff_B_7YSbfqLc6_2;
	wire w_dff_B_br1dIeQV4_2;
	wire w_dff_B_KpEuoHQc7_2;
	wire w_dff_B_nH6yqGFt7_2;
	wire w_dff_B_k7FErPul7_2;
	wire w_dff_B_n9aGapcV5_2;
	wire w_dff_B_NVE8bpjW7_2;
	wire w_dff_B_bK2InPNT6_2;
	wire w_dff_B_oWdkY0Gi6_2;
	wire w_dff_B_rfjTdLWg6_2;
	wire w_dff_B_6OlVESxY9_2;
	wire w_dff_B_uqLgkRFO9_2;
	wire w_dff_B_Lnio3Zql7_2;
	wire w_dff_B_z4nlAwtf6_2;
	wire w_dff_B_DvKdE5fy1_2;
	wire w_dff_B_ZFyPLXeB2_2;
	wire w_dff_B_PXKTojbK7_2;
	wire w_dff_B_qxRhpnAz0_2;
	wire w_dff_B_OsCNhheQ6_2;
	wire w_dff_B_Z02BIdNg0_2;
	wire w_dff_B_Ebr1VH9l9_2;
	wire w_dff_B_pVJGLeRL7_2;
	wire w_dff_B_ao91obDv1_2;
	wire w_dff_B_4xpjW6mv9_2;
	wire w_dff_B_LAVnKpcM7_1;
	wire w_dff_B_3BT3or5H8_2;
	wire w_dff_B_Z4EtcHTU7_2;
	wire w_dff_B_HU98oJWt6_2;
	wire w_dff_B_Z1xelDDy1_2;
	wire w_dff_B_trYHmvBe8_2;
	wire w_dff_B_4gKp8EFT8_2;
	wire w_dff_B_AF0608h03_2;
	wire w_dff_B_YtbohqzK5_2;
	wire w_dff_B_OkgsXH552_2;
	wire w_dff_B_H5s0HGV35_2;
	wire w_dff_B_frD7O9NK8_2;
	wire w_dff_B_1m8GGWQI6_2;
	wire w_dff_B_CR7uknkT1_2;
	wire w_dff_B_rq8TM1ly0_2;
	wire w_dff_B_yZ2DPA2L6_2;
	wire w_dff_B_qPRdAYD37_2;
	wire w_dff_B_kYnLVwGx9_2;
	wire w_dff_B_ADDWrBKg7_2;
	wire w_dff_B_zNLnX71z2_2;
	wire w_dff_B_d4nEiHRz9_2;
	wire w_dff_B_aoIjgNAi7_2;
	wire w_dff_B_RYkSGtmM3_1;
	wire w_dff_B_YUD9nspG2_2;
	wire w_dff_B_UUqmA8X71_2;
	wire w_dff_B_aubJzKXX8_2;
	wire w_dff_B_qhmQ3wqw2_2;
	wire w_dff_B_JRoSQOaS8_2;
	wire w_dff_B_48cd8Bc66_2;
	wire w_dff_B_EG6g5fEI9_2;
	wire w_dff_B_n5FdlT3x7_2;
	wire w_dff_B_1ZaeDNct5_2;
	wire w_dff_B_bgmMBiAu4_2;
	wire w_dff_B_oJ3U0Udn5_2;
	wire w_dff_B_6WqpbwZZ0_2;
	wire w_dff_B_EFo5p8J57_2;
	wire w_dff_B_J8iXcCjd8_2;
	wire w_dff_B_AqMfvCMo8_2;
	wire w_dff_B_8C8LvwYj9_2;
	wire w_dff_B_atvicVez0_2;
	wire w_dff_B_q9E9E1EZ5_2;
	wire w_dff_B_pky1lf7R0_1;
	wire w_dff_B_cop3KlzS0_2;
	wire w_dff_B_7Pfajhzu8_2;
	wire w_dff_B_Qa3fqE9G6_2;
	wire w_dff_B_WL7rJb5t8_2;
	wire w_dff_B_81MAUXDq3_2;
	wire w_dff_B_bI8U3JD88_2;
	wire w_dff_B_SOrQUK9g3_2;
	wire w_dff_B_bn8T6aC32_2;
	wire w_dff_B_MxMY04SY1_2;
	wire w_dff_B_hoD6JlkO7_2;
	wire w_dff_B_QCN9vbEl6_2;
	wire w_dff_B_XkTyAUcG1_2;
	wire w_dff_B_CkImynzt0_2;
	wire w_dff_B_vtGoz9zg2_2;
	wire w_dff_B_GvEQLVg08_2;
	wire w_dff_B_QHE2z7Ie5_1;
	wire w_dff_B_bLxyMb3P9_2;
	wire w_dff_B_cvBs6jAA5_2;
	wire w_dff_B_Kg8QyU639_2;
	wire w_dff_B_WKoQoKNC6_2;
	wire w_dff_B_IBDF3cDn0_2;
	wire w_dff_B_tzQdXW0o1_2;
	wire w_dff_B_9JWlaWHN3_2;
	wire w_dff_B_kYa6cxna7_2;
	wire w_dff_B_PhvJ10wD4_2;
	wire w_dff_B_z02FG4Ot5_2;
	wire w_dff_B_kjssqN031_2;
	wire w_dff_B_R87REC4W0_2;
	wire w_dff_B_YlGTExVH1_1;
	wire w_dff_B_ePkst0b07_2;
	wire w_dff_B_087CWndQ4_2;
	wire w_dff_B_UsXfUvZq6_2;
	wire w_dff_B_87JjQ5LB2_2;
	wire w_dff_B_hfEbtF9y3_2;
	wire w_dff_B_wIRjB66Y0_2;
	wire w_dff_B_va1fvv802_2;
	wire w_dff_B_fFbYDQIW4_2;
	wire w_dff_B_S4QVlaXz1_2;
	wire w_dff_B_VvMOypjG3_2;
	wire w_dff_B_nCxF0Fs43_2;
	wire w_dff_B_HWfi7Esq8_1;
	wire w_dff_B_6q58Zi7A0_1;
	wire w_dff_B_ATyUjume4_2;
	wire w_dff_B_HjpMqqJB6_2;
	wire w_dff_B_wPhdDcjg4_2;
	wire w_dff_B_JIdhCC2w7_0;
	wire w_dff_A_kmoZ7gjB8_0;
	wire w_dff_A_qgqYeQLl3_0;
	wire w_dff_A_hGhDz4u86_1;
	wire w_dff_A_qSqHHLZm1_1;
	wire w_dff_B_RNmKnxNj1_1;
	wire w_dff_A_kB4EvvLH8_1;
	wire w_dff_B_EjhvP3lH5_1;
	wire w_dff_B_86NpWNeW8_2;
	wire w_dff_B_MHrQKCMV5_2;
	wire w_dff_B_2YxjOSjQ7_2;
	wire w_dff_B_DxQyfBfM7_2;
	wire w_dff_B_1ZJYhFPx1_2;
	wire w_dff_B_ZGAvkeWZ3_2;
	wire w_dff_B_wY2YYS6D7_2;
	wire w_dff_B_nwQcUs8N8_2;
	wire w_dff_B_rRVXfMNa0_2;
	wire w_dff_B_oYbLJG688_2;
	wire w_dff_B_I4PYwhX82_2;
	wire w_dff_B_e4Ss7TB39_2;
	wire w_dff_B_9US6O8uT3_2;
	wire w_dff_B_swadolk93_2;
	wire w_dff_B_HS4oMSVO2_2;
	wire w_dff_B_4TPCzsBT0_2;
	wire w_dff_B_PUCIrwSb8_2;
	wire w_dff_B_iS7dKMz94_2;
	wire w_dff_B_ud2SorNx9_2;
	wire w_dff_B_44ClnKSg6_2;
	wire w_dff_B_AmEBpAcH4_2;
	wire w_dff_B_D1n7xwRJ6_2;
	wire w_dff_B_uga1Kz5B5_2;
	wire w_dff_B_VFfhgVS75_2;
	wire w_dff_B_HmIja5Vp0_2;
	wire w_dff_B_C9x4hNgZ1_2;
	wire w_dff_B_tkL76kbB1_2;
	wire w_dff_B_oG3I6i9v9_2;
	wire w_dff_B_ab25Dm6h1_2;
	wire w_dff_B_bhFxR8fG6_2;
	wire w_dff_B_0ecvAmry6_2;
	wire w_dff_B_A0HQTnRS5_2;
	wire w_dff_B_1Ji9BOsi7_2;
	wire w_dff_B_LaJRO3fp4_2;
	wire w_dff_B_FV0XBqGk8_2;
	wire w_dff_B_NjCPu9Mz0_2;
	wire w_dff_B_I0iEEkOt3_2;
	wire w_dff_B_Lt0jMCye4_2;
	wire w_dff_B_GGFHYT3U8_2;
	wire w_dff_B_tkUk5iCJ8_2;
	wire w_dff_B_kpk8K8ZK8_2;
	wire w_dff_B_VzYXxpMT1_2;
	wire w_dff_B_jRGarOmj8_2;
	wire w_dff_B_vwd53Nsd6_2;
	wire w_dff_B_ogga8Sqf7_2;
	wire w_dff_B_pE3RY6EJ3_2;
	wire w_dff_B_sNHG63tc4_2;
	wire w_dff_B_Hda611ca5_1;
	wire w_dff_B_zXXELH222_2;
	wire w_dff_B_Q5Wo0zzI6_2;
	wire w_dff_B_hFCgGp9V9_2;
	wire w_dff_B_ZIWHJBJw3_2;
	wire w_dff_B_aIgN8ii19_2;
	wire w_dff_B_YZOVsGuE4_2;
	wire w_dff_B_MGVTiXsw6_2;
	wire w_dff_B_78Qz7F2r8_2;
	wire w_dff_B_sfvx99TZ5_2;
	wire w_dff_B_0PMYyms69_2;
	wire w_dff_B_sOnGZSRu0_2;
	wire w_dff_B_jZsMk6Zv9_2;
	wire w_dff_B_JmUourcI3_2;
	wire w_dff_B_27738wuW2_2;
	wire w_dff_B_C1SmVTst8_2;
	wire w_dff_B_QNWiyBi36_2;
	wire w_dff_B_xdFx4idk7_2;
	wire w_dff_B_cHjPVH1P8_2;
	wire w_dff_B_J99FYGp43_2;
	wire w_dff_B_JP3qFZba7_2;
	wire w_dff_B_3oMdCaRj7_2;
	wire w_dff_B_QFVFKalo4_2;
	wire w_dff_B_8T1GbwaS4_2;
	wire w_dff_B_KPiNWqn23_2;
	wire w_dff_B_lmoQQE0S4_2;
	wire w_dff_B_gXzfq2pK9_2;
	wire w_dff_B_yVuYxYSV7_2;
	wire w_dff_B_5fYUDq1q6_2;
	wire w_dff_B_2WKPpk5e7_2;
	wire w_dff_B_zPGj7Znh0_2;
	wire w_dff_B_GML0Fae86_2;
	wire w_dff_B_pJOJ8wix4_2;
	wire w_dff_B_xemwHUVc7_2;
	wire w_dff_B_ttnCY9od6_2;
	wire w_dff_B_E8XeTHSK4_2;
	wire w_dff_B_SfNyBD0v8_2;
	wire w_dff_B_vZKQ6Mfu5_2;
	wire w_dff_B_w5g9bPqK3_2;
	wire w_dff_B_QoEsyjak3_2;
	wire w_dff_B_CYpQHWUI5_2;
	wire w_dff_B_7qTU7lys5_2;
	wire w_dff_B_RQf5jV8H4_2;
	wire w_dff_B_8O6FL66n5_2;
	wire w_dff_B_PWGUw7d86_1;
	wire w_dff_B_UjtCsIq95_2;
	wire w_dff_B_2FBFf7nb9_2;
	wire w_dff_B_A3hZxBXW2_2;
	wire w_dff_B_IxevdxLc8_2;
	wire w_dff_B_xQ3h8aY55_2;
	wire w_dff_B_DkOgFsMV8_2;
	wire w_dff_B_fJBcM0qM6_2;
	wire w_dff_B_L7sjh2oX9_2;
	wire w_dff_B_IyDywO801_2;
	wire w_dff_B_gE8xoJnz6_2;
	wire w_dff_B_0TEbxsic0_2;
	wire w_dff_B_o6TRXdeQ0_2;
	wire w_dff_B_p7CqJLlQ0_2;
	wire w_dff_B_ZneqRuYq6_2;
	wire w_dff_B_45jqCXTn0_2;
	wire w_dff_B_Qq7vmDBE6_2;
	wire w_dff_B_eA3vTREJ7_2;
	wire w_dff_B_KcisPGXK9_2;
	wire w_dff_B_WEDuEVWN1_2;
	wire w_dff_B_plOaHfpE7_2;
	wire w_dff_B_emkmWjAt8_2;
	wire w_dff_B_qvuQ9Hzb7_2;
	wire w_dff_B_5Fzxgran2_2;
	wire w_dff_B_dP9OO4NJ2_2;
	wire w_dff_B_1CLlZGws5_2;
	wire w_dff_B_bq2q6p1G5_2;
	wire w_dff_B_pr619eye4_2;
	wire w_dff_B_Hpxyhvh51_2;
	wire w_dff_B_gbTO50EO7_2;
	wire w_dff_B_jIfg9ag48_2;
	wire w_dff_B_NCdnn3Yy6_2;
	wire w_dff_B_yQ8ZbIFE5_2;
	wire w_dff_B_KQnXlsq47_2;
	wire w_dff_B_VYo8NXq32_2;
	wire w_dff_B_jetdDKut5_2;
	wire w_dff_B_hodL1qM27_2;
	wire w_dff_B_weh610iE4_2;
	wire w_dff_B_ryjsFclc7_2;
	wire w_dff_B_TkxqROVW5_1;
	wire w_dff_B_ILYBq7oC4_2;
	wire w_dff_B_FhiqZvdu7_2;
	wire w_dff_B_jRvyvnNH2_2;
	wire w_dff_B_8SniH8HP9_2;
	wire w_dff_B_7a3dHNp73_2;
	wire w_dff_B_qOPBmmdJ9_2;
	wire w_dff_B_hqkURLnP4_2;
	wire w_dff_B_dYMx2zw50_2;
	wire w_dff_B_e8kVhg791_2;
	wire w_dff_B_F7tCiPu11_2;
	wire w_dff_B_SjbfP5Z02_2;
	wire w_dff_B_xX9DT0jS3_2;
	wire w_dff_B_pU3K24Qg8_2;
	wire w_dff_B_97WXnysl8_2;
	wire w_dff_B_wsh8o2237_2;
	wire w_dff_B_E3vO13B00_2;
	wire w_dff_B_BwToRSrO5_2;
	wire w_dff_B_ta7y8tgH6_2;
	wire w_dff_B_4dE50Gwp8_2;
	wire w_dff_B_4466LlwD0_2;
	wire w_dff_B_MXoQ7O9y8_2;
	wire w_dff_B_D2wU16SM2_2;
	wire w_dff_B_TRmMkrUB4_2;
	wire w_dff_B_wJ2AoZmT2_2;
	wire w_dff_B_rJkbEKeZ2_2;
	wire w_dff_B_QiWiEkcq3_2;
	wire w_dff_B_nz7xI0Ml6_2;
	wire w_dff_B_PO2f7dKZ3_2;
	wire w_dff_B_cg2pk6Qf3_2;
	wire w_dff_B_7VfQK97E2_2;
	wire w_dff_B_0x1OAe0j3_2;
	wire w_dff_B_77bUs3HG7_2;
	wire w_dff_B_BikqO5xy9_2;
	wire w_dff_B_FUvRPWGM6_2;
	wire w_dff_B_7kyonYWH5_2;
	wire w_dff_B_Lxj1A7jA7_2;
	wire w_dff_B_hpSnetn01_1;
	wire w_dff_B_WHa8wRvB1_2;
	wire w_dff_B_49e0OhMy7_2;
	wire w_dff_B_OhDGhI9z1_2;
	wire w_dff_B_HnJpM4PZ3_2;
	wire w_dff_B_y9xdCoen3_2;
	wire w_dff_B_TxxhFT373_2;
	wire w_dff_B_FqhYvdZG8_2;
	wire w_dff_B_fRqZcGXX4_2;
	wire w_dff_B_iNo8s8U23_2;
	wire w_dff_B_tikmd1Ny1_2;
	wire w_dff_B_ikuEt39o1_2;
	wire w_dff_B_O9CkpP3U1_2;
	wire w_dff_B_r82IGXdZ6_2;
	wire w_dff_B_3grm17AD7_2;
	wire w_dff_B_xyafewkp7_2;
	wire w_dff_B_e4RXbdMU0_2;
	wire w_dff_B_I5hyxxs73_2;
	wire w_dff_B_wqi8rNtI1_2;
	wire w_dff_B_G2C80Fdd2_2;
	wire w_dff_B_oD2Hcv5r4_2;
	wire w_dff_B_fog9XP5O2_2;
	wire w_dff_B_5HXJhtaF3_2;
	wire w_dff_B_0NoRYcOp6_2;
	wire w_dff_B_btDNh6wR3_2;
	wire w_dff_B_d87YSAsi0_2;
	wire w_dff_B_DGq3LQSS9_2;
	wire w_dff_B_8mcX23te9_2;
	wire w_dff_B_FrAHjZAT7_2;
	wire w_dff_B_f3ceJS240_2;
	wire w_dff_B_nPrlUkPQ9_2;
	wire w_dff_B_YkPAgCZk6_2;
	wire w_dff_B_Hlxo0DKL6_2;
	wire w_dff_B_tqh4Egzt0_2;
	wire w_dff_B_AGOGhga26_1;
	wire w_dff_B_iKkpZuvh2_2;
	wire w_dff_B_d2JHRYAE6_2;
	wire w_dff_B_dQVzrfqs2_2;
	wire w_dff_B_Y2i3sSXZ1_2;
	wire w_dff_B_hoj4EpN59_2;
	wire w_dff_B_itmNrREO9_2;
	wire w_dff_B_f8KWNAef2_2;
	wire w_dff_B_JUkqhfsD7_2;
	wire w_dff_B_W1exKHoF5_2;
	wire w_dff_B_dnQuA9eV7_2;
	wire w_dff_B_OYrOFMKU8_2;
	wire w_dff_B_ru2tzxYP9_2;
	wire w_dff_B_q2WK9FCg1_2;
	wire w_dff_B_TRrY3cb73_2;
	wire w_dff_B_L2hbt7Qv3_2;
	wire w_dff_B_bomolWtn5_2;
	wire w_dff_B_ExVtAqnd6_2;
	wire w_dff_B_K8NCccEu6_2;
	wire w_dff_B_eZaVu03u2_2;
	wire w_dff_B_WWe23Agw5_2;
	wire w_dff_B_6UxDvB6k9_2;
	wire w_dff_B_9Cqae6962_2;
	wire w_dff_B_atxFZfKO9_2;
	wire w_dff_B_BTNP1cHa8_2;
	wire w_dff_B_JuGvrBSW0_2;
	wire w_dff_B_rj9OZnPs9_2;
	wire w_dff_B_Rwy09Gx62_2;
	wire w_dff_B_35y5uoGK4_2;
	wire w_dff_B_efYzMPz54_2;
	wire w_dff_B_SkDVNICh2_2;
	wire w_dff_B_aLxXaBkb0_1;
	wire w_dff_B_9vvyijU41_2;
	wire w_dff_B_Jc3wGxe92_2;
	wire w_dff_B_uQ6ZivpW7_2;
	wire w_dff_B_PDOuhlgu0_2;
	wire w_dff_B_NZfyBnrl7_2;
	wire w_dff_B_58NyR2xG8_2;
	wire w_dff_B_QEhTsO0T2_2;
	wire w_dff_B_iLLBdhIE1_2;
	wire w_dff_B_2ziVN1Cx5_2;
	wire w_dff_B_XGkMAYdB5_2;
	wire w_dff_B_AORQPlV59_2;
	wire w_dff_B_dzu6utUz2_2;
	wire w_dff_B_9ObBPCfB6_2;
	wire w_dff_B_kVeQ6qku3_2;
	wire w_dff_B_6coCRPyg8_2;
	wire w_dff_B_dAI4pKjT4_2;
	wire w_dff_B_J4mpgpSg0_2;
	wire w_dff_B_PDNZTc5s5_2;
	wire w_dff_B_zAeVcSGl7_2;
	wire w_dff_B_3hbZyOdU6_2;
	wire w_dff_B_CUOsoGQR6_2;
	wire w_dff_B_RPwjE7CU8_2;
	wire w_dff_B_aNEZFJig2_2;
	wire w_dff_B_nnEA6jhf4_2;
	wire w_dff_B_2FugCIN58_2;
	wire w_dff_B_Z2H3KzTz3_2;
	wire w_dff_B_c3ouuaHN5_2;
	wire w_dff_B_C3FFnonp9_1;
	wire w_dff_B_NMSto3Mm2_2;
	wire w_dff_B_I1LkqqKz2_2;
	wire w_dff_B_GxBhb5m90_2;
	wire w_dff_B_LkBNXGK29_2;
	wire w_dff_B_sLmW6l7F5_2;
	wire w_dff_B_CF4SF6d23_2;
	wire w_dff_B_RRYrR1jQ7_2;
	wire w_dff_B_DHizh3n91_2;
	wire w_dff_B_9q7jPIU23_2;
	wire w_dff_B_smlRYZrp1_2;
	wire w_dff_B_jKewHi7F5_2;
	wire w_dff_B_Zx0BdT2J9_2;
	wire w_dff_B_GwqkwY8C5_2;
	wire w_dff_B_qMg2IR714_2;
	wire w_dff_B_8gFIau1v5_2;
	wire w_dff_B_0RWu5RWr2_2;
	wire w_dff_B_6YTeBN2C2_2;
	wire w_dff_B_VDewpwzq9_2;
	wire w_dff_B_qqZ9UZjH3_2;
	wire w_dff_B_1bpYPDPy7_2;
	wire w_dff_B_mbKxSyET4_2;
	wire w_dff_B_zPTss1mL8_2;
	wire w_dff_B_fFzEiE7X7_2;
	wire w_dff_B_gVfB6OuJ0_2;
	wire w_dff_B_6uAOIO527_1;
	wire w_dff_B_Og1E3fEo7_2;
	wire w_dff_B_p1K4nSmB2_2;
	wire w_dff_B_VtvaCsJW8_2;
	wire w_dff_B_GdcaahH54_2;
	wire w_dff_B_cNYtdx9M4_2;
	wire w_dff_B_lTAmXAox1_2;
	wire w_dff_B_MrIi5FUd4_2;
	wire w_dff_B_shbaHQVl7_2;
	wire w_dff_B_kbqHaiSe3_2;
	wire w_dff_B_UAKDsih58_2;
	wire w_dff_B_XPrKZe582_2;
	wire w_dff_B_XTgMDWXg5_2;
	wire w_dff_B_EBQ3XWoe6_2;
	wire w_dff_B_ufxvtP217_2;
	wire w_dff_B_zMjPcx6u5_2;
	wire w_dff_B_kFRRaUWn9_2;
	wire w_dff_B_QCFiVIu31_2;
	wire w_dff_B_UkwlhGwZ4_2;
	wire w_dff_B_4ijmjSmD2_2;
	wire w_dff_B_aeK2CoD29_2;
	wire w_dff_B_642m3ZPH9_2;
	wire w_dff_B_V7jV1Ext4_1;
	wire w_dff_B_H0eY1vCP7_2;
	wire w_dff_B_kGDEyA688_2;
	wire w_dff_B_7midFWKD9_2;
	wire w_dff_B_7RTBT8P87_2;
	wire w_dff_B_O192w7cy9_2;
	wire w_dff_B_MfCgHR8F5_2;
	wire w_dff_B_5xHweeaR5_2;
	wire w_dff_B_UWykl13E0_2;
	wire w_dff_B_S25beSWm8_2;
	wire w_dff_B_2ATTapyC3_2;
	wire w_dff_B_vwNcG6CI9_2;
	wire w_dff_B_fBp0edJv9_2;
	wire w_dff_B_Zp6cFr067_2;
	wire w_dff_B_jIB7rih82_2;
	wire w_dff_B_JEI8yRGU7_2;
	wire w_dff_B_Z4HN1GRr4_2;
	wire w_dff_B_d7RAo6mC7_2;
	wire w_dff_B_6ZVNhIwl0_2;
	wire w_dff_B_hXdk3x3M0_1;
	wire w_dff_B_XJQ9mYHf9_2;
	wire w_dff_B_nnmoNH6T1_2;
	wire w_dff_B_qwE0HqvV7_2;
	wire w_dff_B_Vzqqvx1Y6_2;
	wire w_dff_B_ny6Xgr5Z5_2;
	wire w_dff_B_nKpA752d8_2;
	wire w_dff_B_Pq9P0IlF6_2;
	wire w_dff_B_CijSerZ83_2;
	wire w_dff_B_BY284Atr3_2;
	wire w_dff_B_MfOHYXdU4_2;
	wire w_dff_B_akuff64K9_2;
	wire w_dff_B_0LkS7Hcw8_2;
	wire w_dff_B_cCZloNXb6_2;
	wire w_dff_B_FZkZf7sr3_2;
	wire w_dff_B_KTLbZe9Y4_2;
	wire w_dff_B_rEp1xRQD0_1;
	wire w_dff_B_P969pCJR7_2;
	wire w_dff_B_xE7UWh4n0_2;
	wire w_dff_B_nAKMsubZ1_2;
	wire w_dff_B_QdT3Hk797_2;
	wire w_dff_B_NWTacWc16_2;
	wire w_dff_B_0pBkhihE4_2;
	wire w_dff_B_045Z5u9l8_2;
	wire w_dff_B_JI6TOvjV8_2;
	wire w_dff_B_j6TlcuSh7_2;
	wire w_dff_B_1qYIf7LQ4_2;
	wire w_dff_B_kkq1ZYEO4_2;
	wire w_dff_B_lqGQoYfm1_2;
	wire w_dff_B_vcmnjSc07_1;
	wire w_dff_B_OQTaVFbh9_2;
	wire w_dff_B_WiQUQgJW6_2;
	wire w_dff_B_5Xp2TDOR3_2;
	wire w_dff_B_GD8msEAh0_2;
	wire w_dff_B_vL374RAq1_2;
	wire w_dff_B_jfRUn2a51_2;
	wire w_dff_B_hW8sr8e47_2;
	wire w_dff_B_an79LytC2_2;
	wire w_dff_B_Tu7fwmsW0_2;
	wire w_dff_B_C45puVrB0_2;
	wire w_dff_B_TtyaOiSh6_2;
	wire w_dff_B_FFb2oKXS3_1;
	wire w_dff_B_bX1BMdYa4_1;
	wire w_dff_B_HaImst948_2;
	wire w_dff_B_viGk7c4i9_2;
	wire w_dff_B_neDSvnNh6_2;
	wire w_dff_B_SDciChy19_0;
	wire w_dff_A_CknfTZA03_0;
	wire w_dff_A_W0GH72gf8_0;
	wire w_dff_A_FaAUVDb87_1;
	wire w_dff_A_7j3bc8678_1;
	wire w_dff_B_v8v4A7LS1_1;
	wire w_dff_A_NtY58GGi5_1;
	wire w_dff_B_xxwiKctb7_1;
	wire w_dff_B_LcJA5Bqi7_2;
	wire w_dff_B_UfNDRm7f6_2;
	wire w_dff_B_GY7K8U8i0_2;
	wire w_dff_B_RrKfvWFU5_2;
	wire w_dff_B_OEJT5zoy2_2;
	wire w_dff_B_rLCi2IIq2_2;
	wire w_dff_B_Yu4juAjS4_2;
	wire w_dff_B_8btXofuv6_2;
	wire w_dff_B_y0ga9Pip0_2;
	wire w_dff_B_tMhWONbk2_2;
	wire w_dff_B_fksUxnGO4_2;
	wire w_dff_B_cfaU7hET9_2;
	wire w_dff_B_Mc80C5zE7_2;
	wire w_dff_B_d9Gem43W8_2;
	wire w_dff_B_8SSLVOf56_2;
	wire w_dff_B_XAQOilhm9_2;
	wire w_dff_B_t5VqixS82_2;
	wire w_dff_B_UWdIDvmW0_2;
	wire w_dff_B_GzsXwmeC3_2;
	wire w_dff_B_exzaH3Wo0_2;
	wire w_dff_B_9DKXb4LL4_2;
	wire w_dff_B_dBANWLne5_2;
	wire w_dff_B_mDhSZInk3_2;
	wire w_dff_B_ftViZq3V6_2;
	wire w_dff_B_q92XC5u46_2;
	wire w_dff_B_07zvVMdD3_2;
	wire w_dff_B_eGdnURNa3_2;
	wire w_dff_B_fg9cwdkh9_2;
	wire w_dff_B_jhWfGbIB8_2;
	wire w_dff_B_EcHovQZ33_2;
	wire w_dff_B_wROgSLxf1_2;
	wire w_dff_B_A1qacFVr2_2;
	wire w_dff_B_Oyk20svl8_2;
	wire w_dff_B_UqmthsR98_2;
	wire w_dff_B_YTU2SVhg0_2;
	wire w_dff_B_2KmRIrEo7_2;
	wire w_dff_B_MVrdaGf84_2;
	wire w_dff_B_fxFJaqLv6_2;
	wire w_dff_B_cLlliuTa4_2;
	wire w_dff_B_S9w9TuCP7_2;
	wire w_dff_B_hBCZ7gpB9_2;
	wire w_dff_B_qoc6ogO33_2;
	wire w_dff_B_Xhm2qsxB3_2;
	wire w_dff_B_VJj0m1Do2_2;
	wire w_dff_B_70PEJUXi4_2;
	wire w_dff_B_13gBd8gh5_2;
	wire w_dff_B_i4eIiAC04_2;
	wire w_dff_B_6OjCEdhs7_2;
	wire w_dff_B_JpN0rZj48_2;
	wire w_dff_B_nqvQXrCN6_1;
	wire w_dff_B_xVGKKs8u1_2;
	wire w_dff_B_71oxvSmr9_2;
	wire w_dff_B_VDWJjfHx8_2;
	wire w_dff_B_Xf5vl8hx4_2;
	wire w_dff_B_irXO5eZF6_2;
	wire w_dff_B_PdQXvMXa8_2;
	wire w_dff_B_sv9CjH9b1_2;
	wire w_dff_B_DU2dZiy92_2;
	wire w_dff_B_AWhWqrac2_2;
	wire w_dff_B_3O9FsM545_2;
	wire w_dff_B_RklGZo928_2;
	wire w_dff_B_2RJ4PmOO0_2;
	wire w_dff_B_EsLEBkm56_2;
	wire w_dff_B_4dIAflDz6_2;
	wire w_dff_B_HGAKkdYK3_2;
	wire w_dff_B_HNQ9b8yK1_2;
	wire w_dff_B_R1W7SSfX6_2;
	wire w_dff_B_rmX5oKrJ3_2;
	wire w_dff_B_ua7b4t665_2;
	wire w_dff_B_14X4e4YK8_2;
	wire w_dff_B_rjQagSH03_2;
	wire w_dff_B_tEFkfzHf9_2;
	wire w_dff_B_TKVOVmoL9_2;
	wire w_dff_B_wttPaOG69_2;
	wire w_dff_B_lqo5lrpD9_2;
	wire w_dff_B_fPe0kNB17_2;
	wire w_dff_B_93UqPvIe5_2;
	wire w_dff_B_TyfrnoXd9_2;
	wire w_dff_B_paY5ipUC3_2;
	wire w_dff_B_GvR4kVTr4_2;
	wire w_dff_B_qG3iUPF92_2;
	wire w_dff_B_nZJLRNkM6_2;
	wire w_dff_B_O8zeAHm31_2;
	wire w_dff_B_s43PEsiD1_2;
	wire w_dff_B_k418u75v3_2;
	wire w_dff_B_gvo1yXTy3_2;
	wire w_dff_B_tfm2uLff8_2;
	wire w_dff_B_WnD1Q5Is7_2;
	wire w_dff_B_uoSSnGrC7_2;
	wire w_dff_B_D2DtCYLZ9_2;
	wire w_dff_B_PNkfvJ2l3_2;
	wire w_dff_B_DU0dxzrJ1_2;
	wire w_dff_B_gXL6O2rA7_2;
	wire w_dff_B_XKc9uIkO5_2;
	wire w_dff_B_5O1Mhl5G7_2;
	wire w_dff_B_tJimsX8j4_1;
	wire w_dff_B_frIaj2RI6_2;
	wire w_dff_B_9GUPOc4G3_2;
	wire w_dff_B_GyDejqQZ6_2;
	wire w_dff_B_iE8ZleQ34_2;
	wire w_dff_B_eDtJpeUn1_2;
	wire w_dff_B_HFfVIqOH7_2;
	wire w_dff_B_4dmr9fh66_2;
	wire w_dff_B_cf7s3GCB7_2;
	wire w_dff_B_BCl9MYeo6_2;
	wire w_dff_B_MSz9wcsF6_2;
	wire w_dff_B_El6EXcGj8_2;
	wire w_dff_B_Z7TBncL22_2;
	wire w_dff_B_UQOTd3cL0_2;
	wire w_dff_B_98lTtZWW4_2;
	wire w_dff_B_BCGqecOT6_2;
	wire w_dff_B_VRL736xT1_2;
	wire w_dff_B_xxQ2KoaD6_2;
	wire w_dff_B_pNqlZkVh7_2;
	wire w_dff_B_iNPiKcZZ0_2;
	wire w_dff_B_71H4NSuf0_2;
	wire w_dff_B_Ne9kFWUv8_2;
	wire w_dff_B_CVGfMbPx2_2;
	wire w_dff_B_uOr5SNYT5_2;
	wire w_dff_B_VFBjNAp29_2;
	wire w_dff_B_79WfRfcl2_2;
	wire w_dff_B_9MKOUFEs4_2;
	wire w_dff_B_gpppMwAA8_2;
	wire w_dff_B_yGXQaSIF9_2;
	wire w_dff_B_dIFafHB12_2;
	wire w_dff_B_NAyzPjTs6_2;
	wire w_dff_B_vdgNYJ4J5_2;
	wire w_dff_B_i2HGev2t7_2;
	wire w_dff_B_P98oAzxN1_2;
	wire w_dff_B_acRU4ZJT8_2;
	wire w_dff_B_Gaj7Yz0v5_2;
	wire w_dff_B_ygTh3g6T2_2;
	wire w_dff_B_1UjozB693_2;
	wire w_dff_B_OhDQm7O98_2;
	wire w_dff_B_FcU1j5sf0_2;
	wire w_dff_B_ak5udAVA0_2;
	wire w_dff_B_Ft9mJuO39_2;
	wire w_dff_B_Jm8IZ2yX3_1;
	wire w_dff_B_TLMwKooz6_2;
	wire w_dff_B_NMoIyqNe9_2;
	wire w_dff_B_3LDtzcG92_2;
	wire w_dff_B_hsZxwD3n0_2;
	wire w_dff_B_ho1mJ0n92_2;
	wire w_dff_B_tPMLtXZC4_2;
	wire w_dff_B_jxTAML3I4_2;
	wire w_dff_B_TbalT7X48_2;
	wire w_dff_B_wi6yv5YD4_2;
	wire w_dff_B_9ZMoTj7O2_2;
	wire w_dff_B_XhlUlpmN9_2;
	wire w_dff_B_0Cy7ds3L9_2;
	wire w_dff_B_JEGO43Gh0_2;
	wire w_dff_B_tlA6hnOO0_2;
	wire w_dff_B_zK57mf7V5_2;
	wire w_dff_B_FVjx6qJ20_2;
	wire w_dff_B_FvOmMJRH7_2;
	wire w_dff_B_ZGkvIe3P5_2;
	wire w_dff_B_Ga7PixhE1_2;
	wire w_dff_B_rQxouyCF0_2;
	wire w_dff_B_DDpThMtg6_2;
	wire w_dff_B_XT9cGpH54_2;
	wire w_dff_B_G4qlP3tX2_2;
	wire w_dff_B_o9Ov8vg08_2;
	wire w_dff_B_Gssfd7i91_2;
	wire w_dff_B_gJP2y6Lp0_2;
	wire w_dff_B_LjADZ1Q38_2;
	wire w_dff_B_KqkiHu1Y1_2;
	wire w_dff_B_glA7izOQ6_2;
	wire w_dff_B_fdEBLbDe0_2;
	wire w_dff_B_PiUtUxb49_2;
	wire w_dff_B_2LgUiKan6_2;
	wire w_dff_B_GTlewXVx6_2;
	wire w_dff_B_fAhIAaFB0_2;
	wire w_dff_B_dJfnV5gX4_2;
	wire w_dff_B_74fhHmmo4_2;
	wire w_dff_B_zJmFRF1S3_2;
	wire w_dff_B_Va8VTkjZ2_1;
	wire w_dff_B_evoA3u0e5_2;
	wire w_dff_B_9fjy1hcf7_2;
	wire w_dff_B_jBbS5RuG5_2;
	wire w_dff_B_FMWHfMZr3_2;
	wire w_dff_B_DXSiYJu52_2;
	wire w_dff_B_JpNzzsqb0_2;
	wire w_dff_B_18VsRlV54_2;
	wire w_dff_B_s0Lwa2JG5_2;
	wire w_dff_B_0ohXihXH0_2;
	wire w_dff_B_xE5GTrDl4_2;
	wire w_dff_B_AJjxi0RM7_2;
	wire w_dff_B_kujdne955_2;
	wire w_dff_B_Z4LdgwLL5_2;
	wire w_dff_B_bng3TENJ8_2;
	wire w_dff_B_Wt50lZFc8_2;
	wire w_dff_B_BP5LinwD5_2;
	wire w_dff_B_df3C4cg64_2;
	wire w_dff_B_o6Oc50zP4_2;
	wire w_dff_B_sYraskPq2_2;
	wire w_dff_B_zdGGUdN12_2;
	wire w_dff_B_Cy6oI1Cd3_2;
	wire w_dff_B_eFwuzjGV8_2;
	wire w_dff_B_25Q8x9Lc6_2;
	wire w_dff_B_B7XcN1c74_2;
	wire w_dff_B_kPP1PRpe4_2;
	wire w_dff_B_LvV2Wnea5_2;
	wire w_dff_B_LDa4iBRi6_2;
	wire w_dff_B_9Sb2e7uA3_2;
	wire w_dff_B_iaf79csc3_2;
	wire w_dff_B_Jmpy6PLJ5_2;
	wire w_dff_B_2cvUCt7I8_2;
	wire w_dff_B_vgDz7HGl0_2;
	wire w_dff_B_NOMqsQbb7_1;
	wire w_dff_B_rzAh5RcK6_2;
	wire w_dff_B_TL3k3i9w3_2;
	wire w_dff_B_BdC1pYdW0_2;
	wire w_dff_B_vHZ2E8h42_2;
	wire w_dff_B_KDPvP8p84_2;
	wire w_dff_B_EJm5QPb62_2;
	wire w_dff_B_js9r2Jih3_2;
	wire w_dff_B_lZryZs087_2;
	wire w_dff_B_KVTqR6m77_2;
	wire w_dff_B_ZrHoH6s26_2;
	wire w_dff_B_iEursiol9_2;
	wire w_dff_B_E0Pr9wZX7_2;
	wire w_dff_B_hwMIAubV0_2;
	wire w_dff_B_A8KORzvp6_2;
	wire w_dff_B_B1JptVA97_2;
	wire w_dff_B_DruRNvMn3_2;
	wire w_dff_B_wrziWZtS7_2;
	wire w_dff_B_qATlgHj86_2;
	wire w_dff_B_oB2yIpW74_2;
	wire w_dff_B_XqrWpKwt9_2;
	wire w_dff_B_UuOQwWzo9_2;
	wire w_dff_B_df8D3KrU1_2;
	wire w_dff_B_b4AD2SLo8_2;
	wire w_dff_B_DNJKM7Bh8_2;
	wire w_dff_B_mhtO42R30_2;
	wire w_dff_B_ljmbFGL86_2;
	wire w_dff_B_5KP6FtA28_2;
	wire w_dff_B_ztnEy9jo6_2;
	wire w_dff_B_XmFqVPUy1_2;
	wire w_dff_B_uFhzbbnU0_2;
	wire w_dff_B_JDhLY78t9_1;
	wire w_dff_B_5M1pZYK88_2;
	wire w_dff_B_riturfmM2_2;
	wire w_dff_B_7TW9ku0j0_2;
	wire w_dff_B_c9TestuX8_2;
	wire w_dff_B_cahsJowi9_2;
	wire w_dff_B_nmQWsTmW6_2;
	wire w_dff_B_PXQIHeDt4_2;
	wire w_dff_B_I7y39cJ69_2;
	wire w_dff_B_7f4shHJb2_2;
	wire w_dff_B_9p19iKxK6_2;
	wire w_dff_B_mv4b9fhm6_2;
	wire w_dff_B_LRfPGIup0_2;
	wire w_dff_B_PJk8RI6r2_2;
	wire w_dff_B_O5bwz0rN8_2;
	wire w_dff_B_tFx8tzA56_2;
	wire w_dff_B_sYCDs1rW4_2;
	wire w_dff_B_2sZRzt4m7_2;
	wire w_dff_B_UYh72TEh3_2;
	wire w_dff_B_Q97c5wcB6_2;
	wire w_dff_B_VnPZuiPs2_2;
	wire w_dff_B_wXh85ooP8_2;
	wire w_dff_B_WKA8rCtM8_2;
	wire w_dff_B_60Sy6Wjk2_2;
	wire w_dff_B_2x0X6PHW1_2;
	wire w_dff_B_LCZc02rR6_2;
	wire w_dff_B_YqVPXIAC4_2;
	wire w_dff_B_R2EcHsrg1_2;
	wire w_dff_B_c1etSVAc6_1;
	wire w_dff_B_M8gCdQYB7_2;
	wire w_dff_B_MA7wPNC92_2;
	wire w_dff_B_eMDarAP04_2;
	wire w_dff_B_9RpXHOHZ2_2;
	wire w_dff_B_8JK15M254_2;
	wire w_dff_B_JLmJrbDQ5_2;
	wire w_dff_B_EIoeWHHn1_2;
	wire w_dff_B_49I5weLS8_2;
	wire w_dff_B_Z5jZu9IV5_2;
	wire w_dff_B_8mrcuC5s8_2;
	wire w_dff_B_AGxnscc05_2;
	wire w_dff_B_pN9nYxDw0_2;
	wire w_dff_B_tTQiORyZ9_2;
	wire w_dff_B_C7gKbrz84_2;
	wire w_dff_B_fCFaMa1U8_2;
	wire w_dff_B_nu8UxruK7_2;
	wire w_dff_B_N1dwY88e5_2;
	wire w_dff_B_ntFrNRJQ9_2;
	wire w_dff_B_ZYJtKi7w4_2;
	wire w_dff_B_3COP6sPn6_2;
	wire w_dff_B_jZOdiYwE2_2;
	wire w_dff_B_Fnt90ml08_2;
	wire w_dff_B_im5OGiDU0_2;
	wire w_dff_B_N8V3kiDx4_2;
	wire w_dff_B_QSeZHBz11_1;
	wire w_dff_B_P98EKWL35_2;
	wire w_dff_B_EGITGzLL9_2;
	wire w_dff_B_mZgwUsGu9_2;
	wire w_dff_B_cA0kpSps9_2;
	wire w_dff_B_goHPfu9Y0_2;
	wire w_dff_B_Mb85K9bQ3_2;
	wire w_dff_B_IXgUMDHr0_2;
	wire w_dff_B_Cp5W3Rwi1_2;
	wire w_dff_B_IgGP0blm0_2;
	wire w_dff_B_cGgvSC5R9_2;
	wire w_dff_B_iWfOXjoi9_2;
	wire w_dff_B_N0bKsjRq7_2;
	wire w_dff_B_QI8I4yxY7_2;
	wire w_dff_B_4valJuJS9_2;
	wire w_dff_B_LeXv3NRD9_2;
	wire w_dff_B_7suEemPV6_2;
	wire w_dff_B_A2H9Q2iP2_2;
	wire w_dff_B_vAKrdrEp2_2;
	wire w_dff_B_YVbkSeii8_2;
	wire w_dff_B_KiwMMxOK1_2;
	wire w_dff_B_0SMno3DD3_2;
	wire w_dff_B_BuVg0Fal8_1;
	wire w_dff_B_uRZnHjlG6_2;
	wire w_dff_B_8JTEWFuK7_2;
	wire w_dff_B_puOSgXYT4_2;
	wire w_dff_B_VJZf9ttj0_2;
	wire w_dff_B_7XAjTZvt0_2;
	wire w_dff_B_4ySnrHkG9_2;
	wire w_dff_B_gutEjDEN5_2;
	wire w_dff_B_jOfjCySS2_2;
	wire w_dff_B_4mPQlNFP8_2;
	wire w_dff_B_uubFtQX79_2;
	wire w_dff_B_yOc8uIUD3_2;
	wire w_dff_B_YMadiFVo3_2;
	wire w_dff_B_KaYKnkPc7_2;
	wire w_dff_B_mmk0al6M9_2;
	wire w_dff_B_ZDLXlVxL8_2;
	wire w_dff_B_b6mkOZUi2_2;
	wire w_dff_B_lyy5Ss3G8_2;
	wire w_dff_B_werfbEQm9_2;
	wire w_dff_B_KfPZcrTp9_1;
	wire w_dff_B_F9p8MiAC1_2;
	wire w_dff_B_RecbO2QY7_2;
	wire w_dff_B_vAQcqUzf8_2;
	wire w_dff_B_Jx2yanIf7_2;
	wire w_dff_B_PcsyNyJa7_2;
	wire w_dff_B_824f8WqV7_2;
	wire w_dff_B_7PsSyqiD1_2;
	wire w_dff_B_xsfhwwj28_2;
	wire w_dff_B_ixAxE6Rj1_2;
	wire w_dff_B_ke8KQ10q4_2;
	wire w_dff_B_aAbtQ7CG6_2;
	wire w_dff_B_xwT7C5Bk9_2;
	wire w_dff_B_h4GS01EF2_2;
	wire w_dff_B_UUS9ub6Q8_2;
	wire w_dff_B_HTmzlJ4h1_2;
	wire w_dff_B_9T1eoiix9_1;
	wire w_dff_B_25xqsulN2_2;
	wire w_dff_B_uZE0YxWa2_2;
	wire w_dff_B_p22cGFRo2_2;
	wire w_dff_B_gIUcLDhp8_2;
	wire w_dff_B_APbCrZMR1_2;
	wire w_dff_B_0Z5tLtuI7_2;
	wire w_dff_B_N2Yi987I9_2;
	wire w_dff_B_NijsNKhx4_2;
	wire w_dff_B_4SJ33FUb7_2;
	wire w_dff_B_8Ky5uIpk2_2;
	wire w_dff_B_5scgfOcd7_2;
	wire w_dff_B_uELAWVEd5_2;
	wire w_dff_B_DhUnkwK37_1;
	wire w_dff_B_ozPk56Ju1_2;
	wire w_dff_B_P8dCb00Q8_2;
	wire w_dff_B_VeOTDZB43_2;
	wire w_dff_B_fqXulsCF2_2;
	wire w_dff_B_UT9xhlH88_2;
	wire w_dff_B_ZXbv9itt5_2;
	wire w_dff_B_NfygFl5U8_2;
	wire w_dff_B_mnqJR6yD3_2;
	wire w_dff_B_SMblcq3r0_2;
	wire w_dff_B_bkF6reiD2_2;
	wire w_dff_B_Ol1vyf5o2_2;
	wire w_dff_B_fnPsljRX7_1;
	wire w_dff_B_728XF6378_1;
	wire w_dff_B_ti08sdLI4_2;
	wire w_dff_B_c9BN89Rz8_2;
	wire w_dff_B_nKqnNbB13_2;
	wire w_dff_B_HZOk2ILt2_0;
	wire w_dff_A_j9vhROl75_0;
	wire w_dff_A_jYzDXLF64_0;
	wire w_dff_A_Inffjh1N0_1;
	wire w_dff_A_Px009JHl6_1;
	wire w_dff_B_ETaZKDi58_1;
	wire w_dff_A_bbY4ozxq3_1;
	wire w_dff_B_FpK85Rv57_1;
	wire w_dff_B_0J7Gc0SF7_2;
	wire w_dff_B_RItlMF0x6_2;
	wire w_dff_B_4MaYUbDN9_2;
	wire w_dff_B_jlak0FYh3_2;
	wire w_dff_B_aHf5LmA61_2;
	wire w_dff_B_akiJMh763_2;
	wire w_dff_B_ZOVKDJZA3_2;
	wire w_dff_B_IZZAaECC8_2;
	wire w_dff_B_Jxu8CMxU9_2;
	wire w_dff_B_5001brXV3_2;
	wire w_dff_B_dXcM6R285_2;
	wire w_dff_B_Zaz86RKs9_2;
	wire w_dff_B_vkoTzYjQ7_2;
	wire w_dff_B_UtflPp6t4_2;
	wire w_dff_B_aXq7BneS8_2;
	wire w_dff_B_lucdm2r45_2;
	wire w_dff_B_cA9cdT9m0_2;
	wire w_dff_B_FTlwbQ8F2_2;
	wire w_dff_B_IcLyjPpy4_2;
	wire w_dff_B_vqs514OL9_2;
	wire w_dff_B_o7AcsVXJ5_2;
	wire w_dff_B_SHJbi5ee7_2;
	wire w_dff_B_ninwYxOX8_2;
	wire w_dff_B_kYsFLzp61_2;
	wire w_dff_B_VxEM1pZE0_2;
	wire w_dff_B_h1enl7NK4_2;
	wire w_dff_B_B2evrgU36_2;
	wire w_dff_B_AB64OUGE6_2;
	wire w_dff_B_m2iV2cTa9_2;
	wire w_dff_B_eiv1bLO56_2;
	wire w_dff_B_ERwakILn1_2;
	wire w_dff_B_3tSAaoF18_2;
	wire w_dff_B_XNXOuQKM1_2;
	wire w_dff_B_tEtmH9Uw5_2;
	wire w_dff_B_ySQWxMvM9_2;
	wire w_dff_B_2MHDgYqP0_2;
	wire w_dff_B_EibVGkX51_2;
	wire w_dff_B_hYSdxW9Z8_2;
	wire w_dff_B_XTovOF3k0_2;
	wire w_dff_B_bLrhwQwU1_2;
	wire w_dff_B_FB5yVCJj2_2;
	wire w_dff_B_ynNgCZhF8_2;
	wire w_dff_B_wfrMVCi33_2;
	wire w_dff_B_9YhcK1cV7_2;
	wire w_dff_B_3KexhzEF3_2;
	wire w_dff_B_OOwgU4En3_2;
	wire w_dff_B_FkR01uEE7_2;
	wire w_dff_B_IXyeuhBa9_2;
	wire w_dff_B_2ARDXNAx6_2;
	wire w_dff_B_LKZsNJGw4_2;
	wire w_dff_B_fNHkhFqF1_2;
	wire w_dff_B_Fwtz0GBI3_1;
	wire w_dff_B_c3RRbHhk2_2;
	wire w_dff_B_Lk9HF94M1_2;
	wire w_dff_B_rxSKNL5Y5_2;
	wire w_dff_B_Y7U2s3x88_2;
	wire w_dff_B_V6mELiII3_2;
	wire w_dff_B_ekMijgTn3_2;
	wire w_dff_B_1ior7ngO6_2;
	wire w_dff_B_QLK2MV150_2;
	wire w_dff_B_hHqeOXhU4_2;
	wire w_dff_B_gJrM9ugt1_2;
	wire w_dff_B_3Cucg19M1_2;
	wire w_dff_B_ygluhhKe9_2;
	wire w_dff_B_pde6lBDY9_2;
	wire w_dff_B_JoOifMwG6_2;
	wire w_dff_B_mRU9JJE20_2;
	wire w_dff_B_pyQmTLtt9_2;
	wire w_dff_B_56Cfhd2K9_2;
	wire w_dff_B_Mr5GeYhh2_2;
	wire w_dff_B_WZBDpkOC1_2;
	wire w_dff_B_m5k2qyLm4_2;
	wire w_dff_B_weMayPOr5_2;
	wire w_dff_B_vOTxNLKD4_2;
	wire w_dff_B_QKR0Eo2v2_2;
	wire w_dff_B_X0qbQzhS3_2;
	wire w_dff_B_RBpoRr485_2;
	wire w_dff_B_nOXV2j3n2_2;
	wire w_dff_B_695sRdqD8_2;
	wire w_dff_B_VcDi0xUx4_2;
	wire w_dff_B_FcldosAC6_2;
	wire w_dff_B_4a77vzdv1_2;
	wire w_dff_B_8aF2ljsM5_2;
	wire w_dff_B_lMk6uqgL8_2;
	wire w_dff_B_e2CVeWme4_2;
	wire w_dff_B_w9DTsEyy9_2;
	wire w_dff_B_kQjwzu7a3_2;
	wire w_dff_B_T1G30gkP9_2;
	wire w_dff_B_1ORF6B2k3_2;
	wire w_dff_B_ycRTIGjs3_2;
	wire w_dff_B_aAyhudJG6_2;
	wire w_dff_B_oAdVFYEh6_2;
	wire w_dff_B_J0HjeCu54_2;
	wire w_dff_B_WgN7AWFO4_2;
	wire w_dff_B_gzyMYr3q3_2;
	wire w_dff_B_tUHatfsD4_2;
	wire w_dff_B_50REtMdL3_2;
	wire w_dff_B_99nspnyh2_2;
	wire w_dff_B_9eIiVIDf5_2;
	wire w_dff_B_bKvMIyeU2_1;
	wire w_dff_B_yyktrpNm2_2;
	wire w_dff_B_bu44eu1B6_2;
	wire w_dff_B_Csz3AXj83_2;
	wire w_dff_B_5CIQqlsm6_2;
	wire w_dff_B_ZDKXoh2w4_2;
	wire w_dff_B_jsKNAhOB9_2;
	wire w_dff_B_JAVoLa977_2;
	wire w_dff_B_HEN85mpg4_2;
	wire w_dff_B_nbzo6lFV1_2;
	wire w_dff_B_m8i7scyu2_2;
	wire w_dff_B_jYT64vM47_2;
	wire w_dff_B_4CLFUP2v3_2;
	wire w_dff_B_mATS5brh5_2;
	wire w_dff_B_YbI7v3Ie3_2;
	wire w_dff_B_DlVDXHU01_2;
	wire w_dff_B_x8TSpmYQ5_2;
	wire w_dff_B_0jjHzCaj3_2;
	wire w_dff_B_BzmtM4pE5_2;
	wire w_dff_B_8EGmo8Zb9_2;
	wire w_dff_B_NBkEa6QD6_2;
	wire w_dff_B_pBSoxbIG2_2;
	wire w_dff_B_6Pc5XPYD7_2;
	wire w_dff_B_POEtoDlq7_2;
	wire w_dff_B_PPwdF0Rf0_2;
	wire w_dff_B_b4gHzTWo4_2;
	wire w_dff_B_VXDnRktu9_2;
	wire w_dff_B_I0Jg6Rsa1_2;
	wire w_dff_B_JSnNrEa39_2;
	wire w_dff_B_f3wVelXf8_2;
	wire w_dff_B_b6Qfe2ap6_2;
	wire w_dff_B_MmGvxAvq5_2;
	wire w_dff_B_6IKtcY6Q6_2;
	wire w_dff_B_eCb2YjhA9_2;
	wire w_dff_B_JodLjeCh7_2;
	wire w_dff_B_cbvCIZhe2_2;
	wire w_dff_B_KCwQgi8Y7_2;
	wire w_dff_B_vmF7H9uT4_2;
	wire w_dff_B_tNCXlTSp5_2;
	wire w_dff_B_vik4YCF04_2;
	wire w_dff_B_hX7Hdih84_2;
	wire w_dff_B_6lFIrJ2u2_2;
	wire w_dff_B_YReXbETt0_2;
	wire w_dff_B_AIRwaqk58_2;
	wire w_dff_B_uWD0VSwd7_1;
	wire w_dff_B_9EP9codA9_2;
	wire w_dff_B_FUCf8NxE5_2;
	wire w_dff_B_NtOVCewy8_2;
	wire w_dff_B_AAmU4A087_2;
	wire w_dff_B_SbpVYm8w6_2;
	wire w_dff_B_ARybbmoo7_2;
	wire w_dff_B_E7QsuqFe9_2;
	wire w_dff_B_UY1f4PDI3_2;
	wire w_dff_B_Fva5N2Ee8_2;
	wire w_dff_B_eO7YgJXN7_2;
	wire w_dff_B_JswO11cn4_2;
	wire w_dff_B_fQ3JW1hU4_2;
	wire w_dff_B_CdvN1CaH5_2;
	wire w_dff_B_mIEG6yNy3_2;
	wire w_dff_B_51WJwNha8_2;
	wire w_dff_B_to2EVpos1_2;
	wire w_dff_B_pC4Hs9Zd0_2;
	wire w_dff_B_o3dLxQRK3_2;
	wire w_dff_B_t0hWqOuN2_2;
	wire w_dff_B_G3E3fsmW4_2;
	wire w_dff_B_g4wAVB2x1_2;
	wire w_dff_B_7k9fO9Rr3_2;
	wire w_dff_B_OJA1FgMG0_2;
	wire w_dff_B_sdiTLzAQ9_2;
	wire w_dff_B_D6jVjiLH7_2;
	wire w_dff_B_MNHBAXIj2_2;
	wire w_dff_B_FmG2Xsxj6_2;
	wire w_dff_B_k7thOBWJ9_2;
	wire w_dff_B_tOKQBhwO5_2;
	wire w_dff_B_gXboCuKn2_2;
	wire w_dff_B_LY9pV0b29_2;
	wire w_dff_B_M1NuotcH0_2;
	wire w_dff_B_bPbudhif3_2;
	wire w_dff_B_fXlLPqGG9_2;
	wire w_dff_B_Tz7bpof40_2;
	wire w_dff_B_5pdr62VP2_2;
	wire w_dff_B_pD8rLnxO2_2;
	wire w_dff_B_NU2VaBpl9_2;
	wire w_dff_B_eSWBskYx7_2;
	wire w_dff_B_td0WxbKe1_1;
	wire w_dff_B_lR1OHnT79_2;
	wire w_dff_B_xExEMAf12_2;
	wire w_dff_B_VeUPoq5F9_2;
	wire w_dff_B_KrF5GXoG2_2;
	wire w_dff_B_aLsi9sQW2_2;
	wire w_dff_B_OGRPt5W52_2;
	wire w_dff_B_QeMouNEn3_2;
	wire w_dff_B_oWAms1w90_2;
	wire w_dff_B_1DjPtBAV0_2;
	wire w_dff_B_DVvfyar48_2;
	wire w_dff_B_SwY7dVbT8_2;
	wire w_dff_B_80SXZOAi3_2;
	wire w_dff_B_cZWOhMBL1_2;
	wire w_dff_B_QmLWvtGn2_2;
	wire w_dff_B_wvOn5yyw2_2;
	wire w_dff_B_d7pYEh2H7_2;
	wire w_dff_B_tUBTESTP5_2;
	wire w_dff_B_u2ewzUzZ6_2;
	wire w_dff_B_fp0m2A314_2;
	wire w_dff_B_Ob11gPZD2_2;
	wire w_dff_B_oB4Rfb6C3_2;
	wire w_dff_B_kMjtllTd1_2;
	wire w_dff_B_ws5sLlAW8_2;
	wire w_dff_B_L3Alvh2Z4_2;
	wire w_dff_B_n0fR6AjL1_2;
	wire w_dff_B_R92hkvZX9_2;
	wire w_dff_B_woDCuFZ14_2;
	wire w_dff_B_sDLU0lsD2_2;
	wire w_dff_B_BCpNfPXZ6_2;
	wire w_dff_B_2HS8vD7d7_2;
	wire w_dff_B_8ujHI00n8_2;
	wire w_dff_B_NzcSzjJV8_2;
	wire w_dff_B_4owFNBrb9_2;
	wire w_dff_B_hVjhuHCc7_2;
	wire w_dff_B_wI1VmqpV6_2;
	wire w_dff_B_XibNqeFm6_1;
	wire w_dff_B_5pNB9v7M9_2;
	wire w_dff_B_UcyDdDiE6_2;
	wire w_dff_B_NUu40z0f2_2;
	wire w_dff_B_WepBRDtN2_2;
	wire w_dff_B_AZ0movJs3_2;
	wire w_dff_B_cYCPIotE5_2;
	wire w_dff_B_GbiYccTs0_2;
	wire w_dff_B_xJjZIcJk9_2;
	wire w_dff_B_jZwxBOn14_2;
	wire w_dff_B_qVWqC9VF1_2;
	wire w_dff_B_KMZ0YBCs6_2;
	wire w_dff_B_s8RtqUdJ7_2;
	wire w_dff_B_nIWwlrBD2_2;
	wire w_dff_B_GMfgLclG6_2;
	wire w_dff_B_0ZKYV8au2_2;
	wire w_dff_B_BlNw9jrD4_2;
	wire w_dff_B_ouJldoFm3_2;
	wire w_dff_B_NCxsBkjw6_2;
	wire w_dff_B_6pBiAHQg1_2;
	wire w_dff_B_JepAfnws1_2;
	wire w_dff_B_A0zD2iT57_2;
	wire w_dff_B_panCBQgy1_2;
	wire w_dff_B_Tg96JtO59_2;
	wire w_dff_B_JLp5wwiB9_2;
	wire w_dff_B_VJ36D2oQ1_2;
	wire w_dff_B_jpKFKqBO4_2;
	wire w_dff_B_Z354jVBY8_2;
	wire w_dff_B_3JIOsrOB6_2;
	wire w_dff_B_6o2KRl8z8_2;
	wire w_dff_B_9zzKoBVo7_2;
	wire w_dff_B_Z5aK2Mqf8_2;
	wire w_dff_B_1lgDSPcO0_1;
	wire w_dff_B_lsal0nxM1_2;
	wire w_dff_B_4cOYH2Bv9_2;
	wire w_dff_B_tfd2igIn3_2;
	wire w_dff_B_6gupaslH9_2;
	wire w_dff_B_sU53PKXp3_2;
	wire w_dff_B_e6AALpjn5_2;
	wire w_dff_B_IR7MDgCE1_2;
	wire w_dff_B_b3GhAzpq8_2;
	wire w_dff_B_PCdLxVcJ4_2;
	wire w_dff_B_O2Kwrf1q8_2;
	wire w_dff_B_CRz5nzIH8_2;
	wire w_dff_B_N0dTfSQ35_2;
	wire w_dff_B_lBy6FCxs8_2;
	wire w_dff_B_mpU0aF9C6_2;
	wire w_dff_B_s1C4YxQa4_2;
	wire w_dff_B_pz1SME7d8_2;
	wire w_dff_B_SGkNHoRI2_2;
	wire w_dff_B_oZc2EKs89_2;
	wire w_dff_B_L5MuNCV12_2;
	wire w_dff_B_7ljeYh7z9_2;
	wire w_dff_B_KrP08cMV3_2;
	wire w_dff_B_be7HGxfU7_2;
	wire w_dff_B_XSatfJ2t5_2;
	wire w_dff_B_Kha9fibu0_2;
	wire w_dff_B_Do3CHlZJ4_2;
	wire w_dff_B_e40zLt7F6_2;
	wire w_dff_B_n19aq9WK1_1;
	wire w_dff_B_ocY5mxKI8_2;
	wire w_dff_B_cxtn1Egs2_2;
	wire w_dff_B_1W71HvGN9_2;
	wire w_dff_B_BD4TXV0W6_2;
	wire w_dff_B_dGnguKrX3_2;
	wire w_dff_B_9hSTjei00_2;
	wire w_dff_B_tiimYwi14_2;
	wire w_dff_B_Hxj5JbAl9_2;
	wire w_dff_B_jGtmp9vK8_2;
	wire w_dff_B_JaunJOqk6_2;
	wire w_dff_B_mKJ5yvwJ9_2;
	wire w_dff_B_KHG8SNb73_2;
	wire w_dff_B_5FD3ET3e4_2;
	wire w_dff_B_7tHAWO2m6_2;
	wire w_dff_B_Rv9qCRPw6_2;
	wire w_dff_B_ZJ6g7wCM7_2;
	wire w_dff_B_YKz3RTM64_2;
	wire w_dff_B_qrh9tmJJ1_2;
	wire w_dff_B_aafwFHd19_2;
	wire w_dff_B_DZkDxv8R1_2;
	wire w_dff_B_ffShLiOs1_2;
	wire w_dff_B_lHCWwTcy0_2;
	wire w_dff_B_MxE3o1cU9_2;
	wire w_dff_B_9iqGyKXP9_2;
	wire w_dff_B_hdB6e6E61_1;
	wire w_dff_B_M8Ag9vRB1_2;
	wire w_dff_B_Fcx6PIzr0_2;
	wire w_dff_B_CJ1gukER8_2;
	wire w_dff_B_6XjSYidV3_2;
	wire w_dff_B_UsYIXMgo5_2;
	wire w_dff_B_UYI1MK2r4_2;
	wire w_dff_B_1cF1h3Hw3_2;
	wire w_dff_B_bC9exOXa0_2;
	wire w_dff_B_1otDCR9r1_2;
	wire w_dff_B_FmaWGmFY1_2;
	wire w_dff_B_6waAWmvV4_2;
	wire w_dff_B_3EcrslVx7_2;
	wire w_dff_B_pEUeYrei9_2;
	wire w_dff_B_t3pldeuE7_2;
	wire w_dff_B_WppsMTJk8_2;
	wire w_dff_B_9DC59lOa2_2;
	wire w_dff_B_qh3rdMGx4_2;
	wire w_dff_B_9aVeab610_2;
	wire w_dff_B_hZIvGtRx0_2;
	wire w_dff_B_bV6shDjr6_2;
	wire w_dff_B_xxLYShRk6_2;
	wire w_dff_B_mjBQCs7h3_1;
	wire w_dff_B_fRNpdsny8_2;
	wire w_dff_B_afn9dtFl0_2;
	wire w_dff_B_wtD52uC91_2;
	wire w_dff_B_r4uCN1Ci0_2;
	wire w_dff_B_j4ddA7yP4_2;
	wire w_dff_B_yrUthAg95_2;
	wire w_dff_B_CMldEojj1_2;
	wire w_dff_B_xllfnvYM3_2;
	wire w_dff_B_7s3mM2d98_2;
	wire w_dff_B_QyqQjF4b8_2;
	wire w_dff_B_2RLERi4D3_2;
	wire w_dff_B_hsEK8ghl4_2;
	wire w_dff_B_VbBFQejO1_2;
	wire w_dff_B_NeAIDJ7I6_2;
	wire w_dff_B_AXWu38c30_2;
	wire w_dff_B_mSEpAkhb3_2;
	wire w_dff_B_AdX8cphv6_2;
	wire w_dff_B_pDsZakwK6_2;
	wire w_dff_B_s9KZOleJ3_1;
	wire w_dff_B_lnZdkdhu8_2;
	wire w_dff_B_3uOXyjC45_2;
	wire w_dff_B_XSQuYT9H0_2;
	wire w_dff_B_1IHjAhvv0_2;
	wire w_dff_B_rJYqr7oy9_2;
	wire w_dff_B_YUxIifb32_2;
	wire w_dff_B_NcDSgTR24_2;
	wire w_dff_B_21N4drx09_2;
	wire w_dff_B_kFATyO175_2;
	wire w_dff_B_zUtO91ct9_2;
	wire w_dff_B_BcBRBhx66_2;
	wire w_dff_B_96nKsbR15_2;
	wire w_dff_B_axJgrRFr3_2;
	wire w_dff_B_PrtgEQao9_2;
	wire w_dff_B_4OQ3Tr7o3_2;
	wire w_dff_B_JEKq79lb7_1;
	wire w_dff_B_7qVTZSt23_2;
	wire w_dff_B_x4LXLFhz1_2;
	wire w_dff_B_vkMs8pXZ9_2;
	wire w_dff_B_YP3WyDY45_2;
	wire w_dff_B_5dYUpLsq5_2;
	wire w_dff_B_1Kun2Lk55_2;
	wire w_dff_B_FOpswNle6_2;
	wire w_dff_B_19sugaSe5_2;
	wire w_dff_B_YZjIsvaf6_2;
	wire w_dff_B_1zRM0Uim6_2;
	wire w_dff_B_jri7Ub2C6_2;
	wire w_dff_B_KpAjid0A5_2;
	wire w_dff_B_XDYSzb834_1;
	wire w_dff_B_zpKd6K8c6_2;
	wire w_dff_B_pHrcQcCv0_2;
	wire w_dff_B_lUwl4kVV6_2;
	wire w_dff_B_MvZZh7PX7_2;
	wire w_dff_B_DbUaWsD48_2;
	wire w_dff_B_qniCvI2i3_2;
	wire w_dff_B_Acp5b3Kh4_2;
	wire w_dff_B_EXMcD6pc9_2;
	wire w_dff_B_xP5YrImD0_2;
	wire w_dff_B_XTmIjNuN8_2;
	wire w_dff_B_5wJlXDlD9_2;
	wire w_dff_B_et0YoBfi1_1;
	wire w_dff_B_Rx5fQxCb1_1;
	wire w_dff_B_3tgqI8hW8_2;
	wire w_dff_B_7TqT456q7_2;
	wire w_dff_B_wYrutqXZ8_2;
	wire w_dff_B_scAyxHrg4_0;
	wire w_dff_A_Ehqss91C2_0;
	wire w_dff_A_96WjFtJZ9_0;
	wire w_dff_A_vxfMr52P9_1;
	wire w_dff_A_z1Kp4bwm6_1;
	wire w_dff_B_jsicA2br8_1;
	wire w_dff_B_EqsQe0zZ2_1;
	wire w_dff_B_SQb1nkqy3_1;
	wire w_dff_B_0ZC1Rhkb4_2;
	wire w_dff_B_b9bKABFx3_2;
	wire w_dff_B_v16KuXGp9_2;
	wire w_dff_B_wAqBbolL7_2;
	wire w_dff_B_Mq6sI9D28_2;
	wire w_dff_B_HfCZ0BMs4_2;
	wire w_dff_B_T9QlhBoH0_2;
	wire w_dff_B_5bFb3YYt0_2;
	wire w_dff_B_CHTigQ4K6_2;
	wire w_dff_B_E1mwLwzD3_2;
	wire w_dff_B_KBkld3fv6_2;
	wire w_dff_B_eyyxhrH93_2;
	wire w_dff_B_ViIgY6qx5_2;
	wire w_dff_B_PSjB8nIS1_2;
	wire w_dff_B_BRTnTT3k5_2;
	wire w_dff_B_orq0XXey8_2;
	wire w_dff_B_w5otUtWB7_2;
	wire w_dff_B_WvWMk6WC9_2;
	wire w_dff_B_dKREafO36_2;
	wire w_dff_B_1gzraluq6_2;
	wire w_dff_B_AJVUYrpd2_2;
	wire w_dff_B_U6GHPRTR5_2;
	wire w_dff_B_ljxAg85k1_2;
	wire w_dff_B_vELiSrbG3_2;
	wire w_dff_B_N6RIcCje6_2;
	wire w_dff_B_0AYq1ozq9_2;
	wire w_dff_B_DhlcXIkj0_2;
	wire w_dff_B_rK11GMSa2_2;
	wire w_dff_B_PZ38W6Yx2_2;
	wire w_dff_B_yjgVH1fF0_2;
	wire w_dff_B_Au7sQFSe9_2;
	wire w_dff_B_IQtbwsbQ9_2;
	wire w_dff_B_ZnVnleM24_2;
	wire w_dff_B_FhLgab0R5_2;
	wire w_dff_B_RmOZQAAW1_2;
	wire w_dff_B_mcoHI9228_2;
	wire w_dff_B_nu9yuFi28_2;
	wire w_dff_B_57nUGVQH7_2;
	wire w_dff_B_WZVjoAz74_2;
	wire w_dff_B_Dj8wHJUw3_2;
	wire w_dff_B_CxuOwJ9T4_2;
	wire w_dff_B_YE5usB9l5_2;
	wire w_dff_B_MaLZ22Bi4_2;
	wire w_dff_B_0vlqLkWt1_2;
	wire w_dff_B_yF9Xkmon8_2;
	wire w_dff_B_oQREDpah4_2;
	wire w_dff_B_3bykjGzj4_2;
	wire w_dff_B_olshoiTp9_2;
	wire w_dff_B_HKO57Efn9_2;
	wire w_dff_B_ngOwxPRj8_2;
	wire w_dff_B_ez7O8DKz6_2;
	wire w_dff_B_CJrNqhDw9_2;
	wire w_dff_B_Yqe5obyU9_2;
	wire w_dff_B_MUkFS5jG6_2;
	wire w_dff_B_OGwC6Rvn1_2;
	wire w_dff_B_gUFxVDau1_2;
	wire w_dff_B_YCYUCBC63_2;
	wire w_dff_B_MDn3ANsS2_2;
	wire w_dff_B_KJ8cCYY08_2;
	wire w_dff_B_TKVh6Ytz4_2;
	wire w_dff_B_4liTS6k20_2;
	wire w_dff_B_eOR086B22_2;
	wire w_dff_B_Hvgmn9CN1_2;
	wire w_dff_B_gQPX1R127_2;
	wire w_dff_B_bAiX3mxd1_2;
	wire w_dff_B_9QjRRC6G0_2;
	wire w_dff_B_iYUtJfo63_2;
	wire w_dff_B_BEjzN3Tk8_2;
	wire w_dff_B_oPkqVb122_2;
	wire w_dff_B_ybM8yBJc6_2;
	wire w_dff_B_AwW3Li6B4_2;
	wire w_dff_B_wDiSjjVo0_2;
	wire w_dff_B_IDfo7be52_2;
	wire w_dff_B_v6NPQO604_2;
	wire w_dff_B_oM8ZydWC4_2;
	wire w_dff_B_7gmdIUcN3_2;
	wire w_dff_B_VJn4hN5I0_2;
	wire w_dff_B_ywgb2ue65_2;
	wire w_dff_B_AhWO7RTD7_2;
	wire w_dff_B_dee6IbdF6_2;
	wire w_dff_B_0sTGuZlx4_2;
	wire w_dff_B_U15bZJxy9_2;
	wire w_dff_B_CBzR9XnT5_2;
	wire w_dff_B_hjGEk3FN1_2;
	wire w_dff_B_UwDtDREG3_2;
	wire w_dff_B_eo8weaP44_2;
	wire w_dff_B_kugiXiML7_2;
	wire w_dff_B_XGFTtA0G2_2;
	wire w_dff_B_KI8OEpS27_2;
	wire w_dff_B_YM4G7ZiF1_2;
	wire w_dff_B_zwpbgDYE5_2;
	wire w_dff_B_XtfTWcjP3_2;
	wire w_dff_B_czZGDbNt3_2;
	wire w_dff_B_UsjuP7vh9_2;
	wire w_dff_B_dVmPfubU1_2;
	wire w_dff_B_4QP4v6QC2_2;
	wire w_dff_B_u7vexqQJ7_2;
	wire w_dff_B_vwqbKnIa1_2;
	wire w_dff_B_hbIAKUDn3_2;
	wire w_dff_B_9xf7aOe23_2;
	wire w_dff_B_Lh8zPf0H3_2;
	wire w_dff_B_z7Oi3qKz3_2;
	wire w_dff_B_mJTxB75M7_2;
	wire w_dff_B_GiZa1NzW1_2;
	wire w_dff_B_dTjgFn7P7_2;
	wire w_dff_B_lMh2uqU83_2;
	wire w_dff_B_bQhuycTN1_2;
	wire w_dff_B_hAmTZHFN2_2;
	wire w_dff_A_WUTJTKWd2_1;
	wire w_dff_B_wGgdgUrc1_1;
	wire w_dff_B_sCeb9wVt9_2;
	wire w_dff_B_ylhITx530_2;
	wire w_dff_B_WjBnJe5F8_2;
	wire w_dff_B_Gg7w9Nh92_2;
	wire w_dff_B_Tvph5wDM4_2;
	wire w_dff_B_dPZPOFDB6_2;
	wire w_dff_B_vnzkRU5m8_2;
	wire w_dff_B_9c3FrUCK4_2;
	wire w_dff_B_C2GU6Yls0_2;
	wire w_dff_B_Lu3HTxUo6_2;
	wire w_dff_B_j23Qzexu3_2;
	wire w_dff_B_1wzHLvu67_2;
	wire w_dff_B_kyItvtrt4_2;
	wire w_dff_B_SvUP6WzU9_2;
	wire w_dff_B_nEcOhYSY9_2;
	wire w_dff_B_VGjiVPLY7_2;
	wire w_dff_B_KQWCpyzV0_2;
	wire w_dff_B_LB2brG6O6_2;
	wire w_dff_B_mI1Zg0cW1_2;
	wire w_dff_B_OXIrjBbR2_2;
	wire w_dff_B_g7im5osU3_2;
	wire w_dff_B_BHDgTPr90_2;
	wire w_dff_B_J8HDxvDj5_2;
	wire w_dff_B_DRquSYQP2_2;
	wire w_dff_B_UFQstv0P5_2;
	wire w_dff_B_NiRYfbKi4_2;
	wire w_dff_B_071mX1x89_2;
	wire w_dff_B_7yCmUlGK8_2;
	wire w_dff_B_3ZGp1siw2_2;
	wire w_dff_B_cuQKHB7k7_2;
	wire w_dff_B_FZ78vUyu4_2;
	wire w_dff_B_70P1lBrn5_2;
	wire w_dff_B_wlbwh8KZ7_2;
	wire w_dff_B_iBMZxMjk1_2;
	wire w_dff_B_mr4jFSFb6_2;
	wire w_dff_B_ui9HzCMJ7_2;
	wire w_dff_B_t5Kw2i9u2_2;
	wire w_dff_B_NSouHv6q5_2;
	wire w_dff_B_gXo3zGkQ7_2;
	wire w_dff_B_Ynzsrzsp4_2;
	wire w_dff_B_3cnBLrxN6_2;
	wire w_dff_B_VLdoh07G5_2;
	wire w_dff_B_ZHJi1bYo6_2;
	wire w_dff_B_SXcydJgu3_2;
	wire w_dff_B_tWmGSrej7_2;
	wire w_dff_B_2lda7fOH1_2;
	wire w_dff_B_e867UfEX2_2;
	wire w_dff_B_0cqTYGmW5_2;
	wire w_dff_B_CLZacbvV3_2;
	wire w_dff_B_ygypAn457_2;
	wire w_dff_B_hWcQC6fp4_2;
	wire w_dff_B_85nnEfjK5_2;
	wire w_dff_B_W6rnKeD31_1;
	wire w_dff_B_RZnj8RYO2_1;
	wire w_dff_B_2J865Ohu3_2;
	wire w_dff_B_HVZ3fHA36_2;
	wire w_dff_B_TqHM9f793_2;
	wire w_dff_B_K8tauUjq6_2;
	wire w_dff_B_7O5ZcEF10_2;
	wire w_dff_B_4O5C7DOo9_2;
	wire w_dff_B_MbmSYfdq3_2;
	wire w_dff_B_8ZHRrLpp7_2;
	wire w_dff_B_nth6Zzm01_2;
	wire w_dff_B_ZBCUt1NI2_2;
	wire w_dff_B_8FaVY4zQ0_2;
	wire w_dff_B_KFce92R43_2;
	wire w_dff_B_qgVSkdWw7_2;
	wire w_dff_B_MfUfDEm14_2;
	wire w_dff_B_SWgQFbfC1_2;
	wire w_dff_B_WY7lLxqQ4_2;
	wire w_dff_B_OoDwh6u38_2;
	wire w_dff_B_XyZwpfnq1_2;
	wire w_dff_B_GULrO4eb3_2;
	wire w_dff_B_6rEcWJbo5_2;
	wire w_dff_B_dh9tn2rf4_2;
	wire w_dff_B_WXktlnfk4_2;
	wire w_dff_B_BScdIvYp7_2;
	wire w_dff_B_fCJsykjG5_2;
	wire w_dff_B_13rVuZoF7_2;
	wire w_dff_B_8q6t7x9G8_2;
	wire w_dff_B_UVZGFrqb4_2;
	wire w_dff_B_Thh2GDD83_2;
	wire w_dff_B_qSWBQnpy2_2;
	wire w_dff_B_jYR6UxKH7_2;
	wire w_dff_B_DbNIh9ig4_2;
	wire w_dff_B_GsJrEfF28_2;
	wire w_dff_B_lDy8tTWb4_2;
	wire w_dff_B_84DxAPml2_2;
	wire w_dff_B_qwVJrxPE7_2;
	wire w_dff_B_7y3vtOru1_2;
	wire w_dff_B_jz9gIu8r3_2;
	wire w_dff_B_0MtxO2Sz1_2;
	wire w_dff_B_XyLSfHrD3_2;
	wire w_dff_B_57i03B9h9_2;
	wire w_dff_B_adTaDt612_2;
	wire w_dff_B_DaLsLcXI6_2;
	wire w_dff_B_3kIobVxA7_2;
	wire w_dff_B_oBF2lXrS3_2;
	wire w_dff_B_sBWxF3Ru3_2;
	wire w_dff_B_5jJWr6HJ8_2;
	wire w_dff_B_BKRyAMPI2_2;
	wire w_dff_B_z22qLd3X2_2;
	wire w_dff_B_Z6YhwrNl1_2;
	wire w_dff_B_BVZmH9Fj5_2;
	wire w_dff_B_7JXgpsbT1_2;
	wire w_dff_B_zL97k3z71_2;
	wire w_dff_B_pqGf6b2E9_2;
	wire w_dff_B_q7YYC9048_2;
	wire w_dff_B_fs7uiKUb7_2;
	wire w_dff_B_lfjrS0234_2;
	wire w_dff_B_WsdavIZf1_2;
	wire w_dff_B_C6gMaQTZ2_2;
	wire w_dff_B_qwozOQVE0_2;
	wire w_dff_B_nhX3f3B65_2;
	wire w_dff_B_hKYoVlqY9_2;
	wire w_dff_B_12yvBWWU6_2;
	wire w_dff_B_XiavbY4o8_2;
	wire w_dff_B_Tc3xqEJy7_2;
	wire w_dff_B_93kJDd5I0_2;
	wire w_dff_B_UrLgxFgP5_2;
	wire w_dff_B_Q8DmjmFR8_2;
	wire w_dff_B_aSdGkBWq0_2;
	wire w_dff_B_6VEaBnXq3_2;
	wire w_dff_B_23Xr9Jzk4_2;
	wire w_dff_B_onEYiaQZ5_2;
	wire w_dff_B_k0aWeSkx5_2;
	wire w_dff_B_Qjb1zy3w3_2;
	wire w_dff_B_cZke7L2V5_2;
	wire w_dff_B_bOhgOz0n7_2;
	wire w_dff_B_lKP4KhVR3_2;
	wire w_dff_B_4cmNqf2c6_2;
	wire w_dff_B_hRg4920O2_2;
	wire w_dff_B_0nGkvphh9_2;
	wire w_dff_B_c0oPyYeU3_2;
	wire w_dff_B_5nOaUjMi0_2;
	wire w_dff_B_zstZZFWV7_2;
	wire w_dff_B_bruJMJFn8_2;
	wire w_dff_B_qM5vG8ip3_2;
	wire w_dff_B_Z2E20n928_2;
	wire w_dff_B_vdWqJbFJ6_2;
	wire w_dff_B_CmabRUo87_2;
	wire w_dff_B_KsfOcV4e3_2;
	wire w_dff_B_n5E5HmvU4_2;
	wire w_dff_B_GzRa2q4H0_2;
	wire w_dff_B_staIUWfV4_2;
	wire w_dff_B_CG8DoOEK9_2;
	wire w_dff_B_o3yT1ZIc1_2;
	wire w_dff_B_qHfqmhz79_2;
	wire w_dff_B_4g1I6MsN8_2;
	wire w_dff_B_dmRd39eB5_2;
	wire w_dff_B_gsq2MKZ29_2;
	wire w_dff_B_8057qEsG4_2;
	wire w_dff_B_QULvV8V88_2;
	wire w_dff_B_BMwC0cpx0_2;
	wire w_dff_B_xwJvQPur6_2;
	wire w_dff_B_7dpaZHxq8_1;
	wire w_dff_B_av0Z4jtR1_2;
	wire w_dff_B_6qEj3pS98_2;
	wire w_dff_B_i9tYDqdD2_2;
	wire w_dff_B_4syNUP6B8_2;
	wire w_dff_B_TyzTntKf3_2;
	wire w_dff_B_yy1RzfvQ4_2;
	wire w_dff_B_gCtZIFNU9_2;
	wire w_dff_B_RGmZhSRa0_2;
	wire w_dff_B_Y2dCptr67_2;
	wire w_dff_B_pnUedo9w9_2;
	wire w_dff_B_nxtiiZGi9_2;
	wire w_dff_B_WsO6rbGz8_2;
	wire w_dff_B_t2pv4I0G9_2;
	wire w_dff_B_dM1QLNk81_2;
	wire w_dff_B_cPgayzv85_2;
	wire w_dff_B_eZhtcYPL1_2;
	wire w_dff_B_UVmh4zAv5_2;
	wire w_dff_B_KSttIiVW9_2;
	wire w_dff_B_NuZYHMkO0_2;
	wire w_dff_B_su2KVq545_2;
	wire w_dff_B_2P1inuRz5_2;
	wire w_dff_B_yY6onhTI9_2;
	wire w_dff_B_xoGKECVJ9_2;
	wire w_dff_B_UVaiboU92_2;
	wire w_dff_B_ICW8Ev2L5_2;
	wire w_dff_B_Nf6GLSV29_2;
	wire w_dff_B_VrN9zv2U0_2;
	wire w_dff_B_ddmjZsiA7_2;
	wire w_dff_B_I6WMBrAw8_2;
	wire w_dff_B_VSHuEfxU0_2;
	wire w_dff_B_uDkSno7C4_2;
	wire w_dff_B_PnF0CkH76_2;
	wire w_dff_B_hnNILBVt1_2;
	wire w_dff_B_t62sOwyR2_2;
	wire w_dff_B_dlcYo8dZ8_2;
	wire w_dff_B_5ZtZWLSG3_2;
	wire w_dff_B_iSX1nsKp7_2;
	wire w_dff_B_Dkg3i56c5_2;
	wire w_dff_B_uhQ1kuob9_2;
	wire w_dff_B_1ivoFxOM5_2;
	wire w_dff_B_v0im1tBe6_2;
	wire w_dff_B_9IkQZ6dB1_2;
	wire w_dff_B_daRRA12K6_2;
	wire w_dff_B_DDDeFEzQ2_2;
	wire w_dff_B_WXeeu8oa4_2;
	wire w_dff_B_9Wo1o3nk9_2;
	wire w_dff_B_piTGDidU7_2;
	wire w_dff_B_J8pEQWx43_2;
	wire w_dff_B_xOGJrbx65_1;
	wire w_dff_B_Eb1e4zv05_1;
	wire w_dff_B_QTUrXhTB7_2;
	wire w_dff_B_bDexCrgx5_2;
	wire w_dff_B_Avs9lNBp1_2;
	wire w_dff_B_2SVGwvrh9_2;
	wire w_dff_B_tlsCTcUM0_2;
	wire w_dff_B_N0zI1NNW1_2;
	wire w_dff_B_E3L3xIaM1_2;
	wire w_dff_B_DTvsiQKD0_2;
	wire w_dff_B_QaZTbXsw8_2;
	wire w_dff_B_QzNICzxk3_2;
	wire w_dff_B_mjeW80UN4_2;
	wire w_dff_B_7kYzLfl41_2;
	wire w_dff_B_dQqgCHMh2_2;
	wire w_dff_B_RMPISNWG4_2;
	wire w_dff_B_8T9FbkBe1_2;
	wire w_dff_B_x1xgvqI17_2;
	wire w_dff_B_3aj5npzq6_2;
	wire w_dff_B_ZKXZdRes4_2;
	wire w_dff_B_OOne1VRC8_2;
	wire w_dff_B_cq6H0Ksa1_2;
	wire w_dff_B_TbOS0GcV4_2;
	wire w_dff_B_TE7dmQcq4_2;
	wire w_dff_B_zPEcD1dR1_2;
	wire w_dff_B_OTgWJMc69_2;
	wire w_dff_B_S0dumocq8_2;
	wire w_dff_B_jgvt7n2v2_2;
	wire w_dff_B_nRTinHS83_2;
	wire w_dff_B_AAvTchCT3_2;
	wire w_dff_B_Y6jvpiLY7_2;
	wire w_dff_B_PYTlLPgU2_2;
	wire w_dff_B_g4p8XUGx3_2;
	wire w_dff_B_4Vgkvirh1_2;
	wire w_dff_B_sGD4DW2H3_2;
	wire w_dff_B_sozmydQQ7_2;
	wire w_dff_B_J3qRzl3k4_2;
	wire w_dff_B_aIvhg7WE1_2;
	wire w_dff_B_VOQUcd8l4_2;
	wire w_dff_B_LTv6hB2J8_2;
	wire w_dff_B_0FfXaU3J1_2;
	wire w_dff_B_hfjAzmzM9_2;
	wire w_dff_B_rM7khkJN1_2;
	wire w_dff_B_OrhBpZSr5_2;
	wire w_dff_B_RTdvRxML0_2;
	wire w_dff_B_LtRtLIKV1_2;
	wire w_dff_B_GdviRPqa7_2;
	wire w_dff_B_s0ChG4Md8_2;
	wire w_dff_B_zp14U6pT5_2;
	wire w_dff_B_USgDcLoi1_2;
	wire w_dff_B_A1zY5Kij0_2;
	wire w_dff_B_rFOK6I2c3_2;
	wire w_dff_B_wHKvree92_2;
	wire w_dff_B_ypwBiEOp5_2;
	wire w_dff_B_aVDZ4jek4_2;
	wire w_dff_B_gGL9Nctf8_2;
	wire w_dff_B_2dwFD92M6_2;
	wire w_dff_B_dTB2xocl2_2;
	wire w_dff_B_WTI3i5HF6_2;
	wire w_dff_B_BIaSBGVc9_2;
	wire w_dff_B_bCYW4vfu7_2;
	wire w_dff_B_doOVltAs6_2;
	wire w_dff_B_SNRvUApd2_2;
	wire w_dff_B_il0aZ23A7_2;
	wire w_dff_B_oOKMVDjz3_2;
	wire w_dff_B_6nf6vUhG4_2;
	wire w_dff_B_KU0hY5iM2_2;
	wire w_dff_B_ku4WOzi16_2;
	wire w_dff_B_Q90A9N5n7_2;
	wire w_dff_B_qTNOXtMI8_2;
	wire w_dff_B_Af15cCWq9_2;
	wire w_dff_B_ZaVDupB09_2;
	wire w_dff_B_a79sutxU0_2;
	wire w_dff_B_wPlm9PoA1_2;
	wire w_dff_B_3RIUMySV6_2;
	wire w_dff_B_5VXRJeTX5_2;
	wire w_dff_B_10E7R6jW3_2;
	wire w_dff_B_4wxEo3nc5_2;
	wire w_dff_B_kz4ZAxxS3_2;
	wire w_dff_B_PJxYP14y4_2;
	wire w_dff_B_U8dQpLzK1_2;
	wire w_dff_B_OMk2KzHJ8_2;
	wire w_dff_B_eKIOurO45_2;
	wire w_dff_B_zRAUS7gg5_2;
	wire w_dff_B_OqyqSyrB2_2;
	wire w_dff_B_l0R9GduR1_2;
	wire w_dff_B_srBtELsK7_2;
	wire w_dff_B_U0i14xFa9_2;
	wire w_dff_B_wDQ379xY9_2;
	wire w_dff_B_fmd4f86b2_2;
	wire w_dff_B_ERW3I19F4_2;
	wire w_dff_B_DqXazg6O0_2;
	wire w_dff_B_xvv2OEut9_2;
	wire w_dff_B_sbxCKHqq8_2;
	wire w_dff_B_pFri1iHH0_2;
	wire w_dff_B_8w4XTPpi9_1;
	wire w_dff_B_4ZmHRJrV1_2;
	wire w_dff_B_9DNKNgt53_2;
	wire w_dff_B_FdlhnPA41_2;
	wire w_dff_B_vZU7n0tT8_2;
	wire w_dff_B_3S5Vq60G4_2;
	wire w_dff_B_L96CCz5K7_2;
	wire w_dff_B_SaIBBEzU0_2;
	wire w_dff_B_Ayo4m5VA7_2;
	wire w_dff_B_pcvehPN78_2;
	wire w_dff_B_YOG5Umbu8_2;
	wire w_dff_B_pgx7HPXs2_2;
	wire w_dff_B_h9LwHkWn0_2;
	wire w_dff_B_5XRL5acR6_2;
	wire w_dff_B_fkDkQe9K9_2;
	wire w_dff_B_d0mRO7T62_2;
	wire w_dff_B_LhW3JaGi3_2;
	wire w_dff_B_A4c859rS3_2;
	wire w_dff_B_4HXw9Oxz5_2;
	wire w_dff_B_BAH15Enk3_2;
	wire w_dff_B_AxzJNU8C1_2;
	wire w_dff_B_y7VGyiwD9_2;
	wire w_dff_B_zS9rBlHi4_2;
	wire w_dff_B_z3DVdtej0_2;
	wire w_dff_B_G6J0wWIt7_2;
	wire w_dff_B_2oLprXB86_2;
	wire w_dff_B_WmSjZBjW8_2;
	wire w_dff_B_jTcoAEOm8_2;
	wire w_dff_B_ZzX2JLmr1_2;
	wire w_dff_B_6VDsy6lD4_2;
	wire w_dff_B_2moIeQY85_2;
	wire w_dff_B_Dsjxsjoh1_2;
	wire w_dff_B_0z0GZMjg5_2;
	wire w_dff_B_AWfUhAC55_2;
	wire w_dff_B_EM9w7JRr1_2;
	wire w_dff_B_ARSC4Ftf7_2;
	wire w_dff_B_7WG6CZLr4_2;
	wire w_dff_B_rBbTmy2f3_2;
	wire w_dff_B_1pfvS0JA0_2;
	wire w_dff_B_cBzBdBST9_2;
	wire w_dff_B_q7Gqt4ro1_2;
	wire w_dff_B_M4eqRp689_2;
	wire w_dff_B_e1L6mD2V7_2;
	wire w_dff_B_VmSCkBYu1_2;
	wire w_dff_B_RXpiju8U5_2;
	wire w_dff_B_CqtpbViC8_1;
	wire w_dff_B_ongJG3EE9_1;
	wire w_dff_B_2CyJdK8Z7_2;
	wire w_dff_B_ncZPwi679_2;
	wire w_dff_B_xop6ylVZ1_2;
	wire w_dff_B_DazW0yQB0_2;
	wire w_dff_B_t9qFKXAZ4_2;
	wire w_dff_B_RnAt7tCc0_2;
	wire w_dff_B_c4jEV9eq6_2;
	wire w_dff_B_8YgfvItd4_2;
	wire w_dff_B_N7oLL6FB0_2;
	wire w_dff_B_7U0dit3X6_2;
	wire w_dff_B_49HGPpv23_2;
	wire w_dff_B_nWfFf0ch5_2;
	wire w_dff_B_wK5urF5u2_2;
	wire w_dff_B_HDQRt5lp3_2;
	wire w_dff_B_b37Hy5GF2_2;
	wire w_dff_B_YyrSW5Ct5_2;
	wire w_dff_B_EsY9RjQV9_2;
	wire w_dff_B_QwVvic7U2_2;
	wire w_dff_B_m5itEPoM5_2;
	wire w_dff_B_u3HUYTPv7_2;
	wire w_dff_B_ghN2Zun31_2;
	wire w_dff_B_7Ru9YPn77_2;
	wire w_dff_B_nqV95iwg0_2;
	wire w_dff_B_s5Q5PXGk8_2;
	wire w_dff_B_0gbvO4OC2_2;
	wire w_dff_B_MJTELs1G5_2;
	wire w_dff_B_YqQifkcW1_2;
	wire w_dff_B_vfPaTgFh9_2;
	wire w_dff_B_N86eqlBb5_2;
	wire w_dff_B_7z0q1ZVd8_2;
	wire w_dff_B_j1TY1evc6_2;
	wire w_dff_B_OUtOs0oT9_2;
	wire w_dff_B_XBVwhZ5j4_2;
	wire w_dff_B_EZrCr98L4_2;
	wire w_dff_B_TMTsCZeM5_2;
	wire w_dff_B_KBGpHGoT8_2;
	wire w_dff_B_VUniCjIM8_2;
	wire w_dff_B_QQSf4ZWy6_2;
	wire w_dff_B_3AcoKcs97_2;
	wire w_dff_B_9hxYjqaB7_2;
	wire w_dff_B_c3ReEHRB7_2;
	wire w_dff_B_R6dPuvtn1_2;
	wire w_dff_B_4IjTNubv8_2;
	wire w_dff_B_KDL99OvQ5_2;
	wire w_dff_B_z4YZp4Du2_2;
	wire w_dff_B_3RgO0TWM3_2;
	wire w_dff_B_eZXbr0V54_2;
	wire w_dff_B_hVJTkY7K6_2;
	wire w_dff_B_bUAIVfIs6_2;
	wire w_dff_B_BILmwwex7_2;
	wire w_dff_B_G7rGZoZ10_2;
	wire w_dff_B_TeLTNiLL3_2;
	wire w_dff_B_rCG0LvIx7_2;
	wire w_dff_B_DBn2FbCR2_2;
	wire w_dff_B_b1lEewrK5_2;
	wire w_dff_B_xK1ZFrHW9_2;
	wire w_dff_B_VcdB7Ems5_2;
	wire w_dff_B_FXNntc2K9_2;
	wire w_dff_B_mYwqHzcf8_2;
	wire w_dff_B_atQJYgGv5_2;
	wire w_dff_B_1NwKVTvC7_2;
	wire w_dff_B_h0WYMxQh4_2;
	wire w_dff_B_xgZmrLAf0_2;
	wire w_dff_B_S2YyZGEL4_2;
	wire w_dff_B_E1c6ZsQY3_2;
	wire w_dff_B_lYb19zPu5_2;
	wire w_dff_B_hCE862NY2_2;
	wire w_dff_B_3uhZAm128_2;
	wire w_dff_B_ppVyT4Hw5_2;
	wire w_dff_B_KZxWwOwg2_2;
	wire w_dff_B_eEqE2GBI5_2;
	wire w_dff_B_f1YAp7Xu1_2;
	wire w_dff_B_yudoXnwW9_2;
	wire w_dff_B_icYVq9Sk3_2;
	wire w_dff_B_06cP4HMr5_2;
	wire w_dff_B_eSa1ax943_2;
	wire w_dff_B_NLyXDzBG8_2;
	wire w_dff_B_hXHlc8EP3_2;
	wire w_dff_B_Mc8N4V6c1_2;
	wire w_dff_B_vcIT8ORZ9_2;
	wire w_dff_B_MmA9o2Px5_2;
	wire w_dff_B_U9sq9dXx5_2;
	wire w_dff_B_fjff3wPx7_2;
	wire w_dff_B_VE9RbqXC4_2;
	wire w_dff_B_tXWfrrrp7_2;
	wire w_dff_B_RYVMzpN97_1;
	wire w_dff_B_x9c3PDcI7_2;
	wire w_dff_B_BnFDsRGs0_2;
	wire w_dff_B_K2L8qRO92_2;
	wire w_dff_B_5xNigKaC1_2;
	wire w_dff_B_GqmQDBGx2_2;
	wire w_dff_B_0QCbbunV0_2;
	wire w_dff_B_qUWE1KkA6_2;
	wire w_dff_B_sj9Xg9yW2_2;
	wire w_dff_B_TRHFsr1R0_2;
	wire w_dff_B_LXdu0AkO8_2;
	wire w_dff_B_AKixe2ru9_2;
	wire w_dff_B_30HM3AC04_2;
	wire w_dff_B_N6nEW1yV9_2;
	wire w_dff_B_KKSF2tfy0_2;
	wire w_dff_B_ZwrOPPdG9_2;
	wire w_dff_B_R15dqJNn9_2;
	wire w_dff_B_xii39iJq9_2;
	wire w_dff_B_YKI5l6Hs2_2;
	wire w_dff_B_aIPBVgCe1_2;
	wire w_dff_B_5O9epzDr1_2;
	wire w_dff_B_tzDgVItv0_2;
	wire w_dff_B_iA10L69m2_2;
	wire w_dff_B_2oWl4rML9_2;
	wire w_dff_B_13pGjisS0_2;
	wire w_dff_B_C2Wc6Wvw6_2;
	wire w_dff_B_s78V3ezX4_2;
	wire w_dff_B_Tv2e50Nm6_2;
	wire w_dff_B_V729JHOL8_2;
	wire w_dff_B_ECinXe1W0_2;
	wire w_dff_B_T98C3kRf7_2;
	wire w_dff_B_Ve65sJdP7_2;
	wire w_dff_B_2NtWCb7J9_2;
	wire w_dff_B_ESrSLO466_2;
	wire w_dff_B_ffJ3eKLO3_2;
	wire w_dff_B_sYSEjoPj5_2;
	wire w_dff_B_cvo0OhbJ5_2;
	wire w_dff_B_NBaznYtg5_2;
	wire w_dff_B_D9nY5kld8_2;
	wire w_dff_B_nxNT8YVZ2_2;
	wire w_dff_B_d19QqC920_2;
	wire w_dff_B_qFz2i5bZ3_1;
	wire w_dff_B_BS5jlJis8_1;
	wire w_dff_B_BCHZwWHr9_2;
	wire w_dff_B_3NkGgqFD3_2;
	wire w_dff_B_iOzz3uqc4_2;
	wire w_dff_B_PeJBjRHi5_2;
	wire w_dff_B_R2pf6reC5_2;
	wire w_dff_B_xrSvcZms1_2;
	wire w_dff_B_A4JIWXhJ2_2;
	wire w_dff_B_iJLRGmSm9_2;
	wire w_dff_B_9wXZ4drW7_2;
	wire w_dff_B_H6k7qUr83_2;
	wire w_dff_B_rnR2EMVn3_2;
	wire w_dff_B_cyYKyTcW9_2;
	wire w_dff_B_LG6HglGr7_2;
	wire w_dff_B_4dF0UD2E1_2;
	wire w_dff_B_7sVx1Bbz7_2;
	wire w_dff_B_Yk6VcBVx3_2;
	wire w_dff_B_SvkAqVdf6_2;
	wire w_dff_B_eTpezwir6_2;
	wire w_dff_B_Fv2vJcsU0_2;
	wire w_dff_B_yw91nAdB1_2;
	wire w_dff_B_nt4QY3Pc6_2;
	wire w_dff_B_OCJ0P7RE3_2;
	wire w_dff_B_TPbdEi4f0_2;
	wire w_dff_B_hmxQUuYV9_2;
	wire w_dff_B_OVrobNsX7_2;
	wire w_dff_B_QtWt3vGn0_2;
	wire w_dff_B_EizkcA7N0_2;
	wire w_dff_B_7iGNFEju4_2;
	wire w_dff_B_qDCwc2Dl8_2;
	wire w_dff_B_UhItJk2c3_2;
	wire w_dff_B_YRbCoiYw2_2;
	wire w_dff_B_cDJB2DsX7_2;
	wire w_dff_B_sWYheQJS9_2;
	wire w_dff_B_pq2DPpZI7_2;
	wire w_dff_B_1vPSXQt52_2;
	wire w_dff_B_MWLO8jro5_2;
	wire w_dff_B_uCOPYHHr4_2;
	wire w_dff_B_cMaruJZQ5_2;
	wire w_dff_B_uYUlhEFw7_2;
	wire w_dff_B_8IVAGVyn6_2;
	wire w_dff_B_DQwNWSSj5_2;
	wire w_dff_B_yVi6PexV2_2;
	wire w_dff_B_2smYxZgT2_2;
	wire w_dff_B_Pi5g5RIl7_2;
	wire w_dff_B_HClIwoj19_2;
	wire w_dff_B_FnMWYGRF4_2;
	wire w_dff_B_W6lJyYdW8_2;
	wire w_dff_B_e8CvEH3I0_2;
	wire w_dff_B_NGhIjFql9_2;
	wire w_dff_B_IF2z2di74_2;
	wire w_dff_B_JPAaHdeJ3_2;
	wire w_dff_B_1Nh4SGeK5_2;
	wire w_dff_B_q1FL87Rh1_2;
	wire w_dff_B_HsRMh7uS3_2;
	wire w_dff_B_sf0OTIXx8_2;
	wire w_dff_B_SvxVQAP35_2;
	wire w_dff_B_NKRMDZ1O4_2;
	wire w_dff_B_XgX7ehYZ6_2;
	wire w_dff_B_HkMirg7a2_2;
	wire w_dff_B_M7ywZa7k3_2;
	wire w_dff_B_cP0VlKjz8_2;
	wire w_dff_B_eA3Yygsi4_2;
	wire w_dff_B_S3H5TUMo6_2;
	wire w_dff_B_gtNkzfLy2_2;
	wire w_dff_B_T2vebjFV1_2;
	wire w_dff_B_HX5HcSot8_2;
	wire w_dff_B_WLbUSyTF1_2;
	wire w_dff_B_RCKDo9C86_2;
	wire w_dff_B_cSOKipbt9_2;
	wire w_dff_B_OqUJ9lt96_2;
	wire w_dff_B_4knkifYT9_2;
	wire w_dff_B_Y81BF20X9_2;
	wire w_dff_B_E0W5cjBN1_2;
	wire w_dff_B_tJ9cO7eA7_2;
	wire w_dff_B_jDunCeCm0_2;
	wire w_dff_B_qm4Xdjn60_2;
	wire w_dff_B_KI6zkGY98_2;
	wire w_dff_B_ntwO1BtR6_1;
	wire w_dff_B_YMrTLbXo8_2;
	wire w_dff_B_Dj5C2tG87_2;
	wire w_dff_B_B9Q1NcNt9_2;
	wire w_dff_B_LJcV8DAo4_2;
	wire w_dff_B_yU9GDdmy5_2;
	wire w_dff_B_oj6I1fhT7_2;
	wire w_dff_B_p1friQVX9_2;
	wire w_dff_B_EPbDH7YQ4_2;
	wire w_dff_B_MAqHVTY94_2;
	wire w_dff_B_P2H9yM5T1_2;
	wire w_dff_B_DC05vVfq0_2;
	wire w_dff_B_CA1fzLZ38_2;
	wire w_dff_B_RHvCyUSp5_2;
	wire w_dff_B_jqEfmEm42_2;
	wire w_dff_B_WrKoJqVN5_2;
	wire w_dff_B_mtWdbZf87_2;
	wire w_dff_B_Cl1VHnoQ1_2;
	wire w_dff_B_8nwFrqKH8_2;
	wire w_dff_B_7xNJ6RWm7_2;
	wire w_dff_B_DuCTP03u4_2;
	wire w_dff_B_irzoq4BI7_2;
	wire w_dff_B_GPPHDsy27_2;
	wire w_dff_B_wCPdB5n86_2;
	wire w_dff_B_H55aBVAt2_2;
	wire w_dff_B_3qhzTdwb9_2;
	wire w_dff_B_DTuG6Slf4_2;
	wire w_dff_B_wwpDl90J9_2;
	wire w_dff_B_fjSPGuSj6_2;
	wire w_dff_B_KmBnLnlX7_2;
	wire w_dff_B_mmDMY6Gu5_2;
	wire w_dff_B_au2uUdBm4_2;
	wire w_dff_B_wB5uG7jW4_2;
	wire w_dff_B_SK2KFuYW8_2;
	wire w_dff_B_RLTDLljs4_2;
	wire w_dff_B_a3whaK1s3_2;
	wire w_dff_B_tYEo24vg1_2;
	wire w_dff_B_jL5LBRT13_1;
	wire w_dff_B_CDUyJ6Ha0_1;
	wire w_dff_B_lu2c9jbA0_2;
	wire w_dff_B_MLfHG4xb3_2;
	wire w_dff_B_cQ1pxbYt1_2;
	wire w_dff_B_2U6o0fJL7_2;
	wire w_dff_B_3F2oAwlg3_2;
	wire w_dff_B_xJSs3pD08_2;
	wire w_dff_B_b2iPkQUb6_2;
	wire w_dff_B_wt3HlLd44_2;
	wire w_dff_B_uGAakRTN8_2;
	wire w_dff_B_rdEeYATn5_2;
	wire w_dff_B_60CvUXGm4_2;
	wire w_dff_B_p2OyUcxS9_2;
	wire w_dff_B_9CfXGiuI0_2;
	wire w_dff_B_OvTsoxPy4_2;
	wire w_dff_B_rTQelcBA9_2;
	wire w_dff_B_8D96CdCl9_2;
	wire w_dff_B_OVG0goZC9_2;
	wire w_dff_B_acOnO6Zc4_2;
	wire w_dff_B_9J3eSEQu2_2;
	wire w_dff_B_35gb3vVg5_2;
	wire w_dff_B_2SA6zfzj1_2;
	wire w_dff_B_jd3EjMk98_2;
	wire w_dff_B_6OpeuCrB2_2;
	wire w_dff_B_aGn6E8B36_2;
	wire w_dff_B_v1pevEXP2_2;
	wire w_dff_B_D4ssf82m6_2;
	wire w_dff_B_y1v2CbCH9_2;
	wire w_dff_B_sYk5t9Lx0_2;
	wire w_dff_B_AKirHMAn0_2;
	wire w_dff_B_8N6yDly67_2;
	wire w_dff_B_DvTfPtjn5_2;
	wire w_dff_B_sQNQuede2_2;
	wire w_dff_B_Xpc4Xt2r4_2;
	wire w_dff_B_9sAn7Fcb6_2;
	wire w_dff_B_hFlYIM527_2;
	wire w_dff_B_lsNPF1TA8_2;
	wire w_dff_B_j0qBV0LY6_2;
	wire w_dff_B_gCtvqu4I2_2;
	wire w_dff_B_RidqMonS5_2;
	wire w_dff_B_nYS2B4yV8_2;
	wire w_dff_B_mchIiVzc1_2;
	wire w_dff_B_sNEh0Q967_2;
	wire w_dff_B_VCfgkNlf1_2;
	wire w_dff_B_k1xKFdHo2_2;
	wire w_dff_B_mQq6qvaZ3_2;
	wire w_dff_B_KYdAZ0ES2_2;
	wire w_dff_B_C8c0Fvhr1_2;
	wire w_dff_B_SSKgi54W2_2;
	wire w_dff_B_j8oz2q7E1_2;
	wire w_dff_B_7tgUzNhT3_2;
	wire w_dff_B_kTTGrVnz1_2;
	wire w_dff_B_frKsoiuy9_2;
	wire w_dff_B_hfd3emXe7_2;
	wire w_dff_B_jccaAOYS8_2;
	wire w_dff_B_rkUXDS3V5_2;
	wire w_dff_B_wSPNl7ez7_2;
	wire w_dff_B_P0WkqwtZ3_2;
	wire w_dff_B_Zk9YvXF85_2;
	wire w_dff_B_G1TmgyV26_2;
	wire w_dff_B_IeFKOpvN1_2;
	wire w_dff_B_IigCEz2c6_2;
	wire w_dff_B_L8vOQTb50_2;
	wire w_dff_B_bd73EToM2_2;
	wire w_dff_B_oWdZxOkF7_2;
	wire w_dff_B_wMxHba9J7_2;
	wire w_dff_B_PCX08hoM6_2;
	wire w_dff_B_3Ec1X0q09_2;
	wire w_dff_B_fUIKiS5m0_2;
	wire w_dff_B_RXKSSsqR2_2;
	wire w_dff_B_lVfrHDpd8_1;
	wire w_dff_B_Tbwpf6xt9_2;
	wire w_dff_B_4p6H30yu9_2;
	wire w_dff_B_NCV5bwJ41_2;
	wire w_dff_B_K5lzGnLK5_2;
	wire w_dff_B_bx0cJ6n45_2;
	wire w_dff_B_YIAzdPWe5_2;
	wire w_dff_B_nfE1RCyW4_2;
	wire w_dff_B_mRxCSs2z4_2;
	wire w_dff_B_XE5Bi9jw8_2;
	wire w_dff_B_jUhfG1Wo0_2;
	wire w_dff_B_a345NiQz9_2;
	wire w_dff_B_axaNYMEY7_2;
	wire w_dff_B_VGkCPCOe3_2;
	wire w_dff_B_v6XLbMiq2_2;
	wire w_dff_B_oZ5UZ9j75_2;
	wire w_dff_B_tvbVsxWb7_2;
	wire w_dff_B_HYtGl2de5_2;
	wire w_dff_B_oJ8eMsRB8_2;
	wire w_dff_B_xNXjctV55_2;
	wire w_dff_B_yn6Jz8C52_2;
	wire w_dff_B_gjSxjEzl5_2;
	wire w_dff_B_tpO9zrKX3_2;
	wire w_dff_B_7o4EZgzI3_2;
	wire w_dff_B_pBitbiE92_2;
	wire w_dff_B_7th584bH8_2;
	wire w_dff_B_IL1auyot5_2;
	wire w_dff_B_Kvf7tkbt7_2;
	wire w_dff_B_ul3IkykT6_2;
	wire w_dff_B_8jLUi6t41_2;
	wire w_dff_B_Q8QnPVam5_2;
	wire w_dff_B_dGEwiIKs9_2;
	wire w_dff_B_NCLO9bGl6_2;
	wire w_dff_B_JqBDnx6C6_1;
	wire w_dff_B_akoQDKb85_1;
	wire w_dff_B_80egostb8_2;
	wire w_dff_B_gcHEIEyP4_2;
	wire w_dff_B_Knq085FN6_2;
	wire w_dff_B_xVBIBO344_2;
	wire w_dff_B_9fHuaslc8_2;
	wire w_dff_B_mnsJi2EB1_2;
	wire w_dff_B_SMHASyAu4_2;
	wire w_dff_B_7IqK6qEg9_2;
	wire w_dff_B_G8JdxIRP1_2;
	wire w_dff_B_R4DsbbLR1_2;
	wire w_dff_B_P472hPn29_2;
	wire w_dff_B_lIDlEYAf0_2;
	wire w_dff_B_dzRvG1Lu5_2;
	wire w_dff_B_9EzyEBcd5_2;
	wire w_dff_B_FD3a6GpS4_2;
	wire w_dff_B_CtD1V4Bz7_2;
	wire w_dff_B_aIZ82vB52_2;
	wire w_dff_B_JQSAppdZ4_2;
	wire w_dff_B_zKhtu69H4_2;
	wire w_dff_B_buyjAk7I1_2;
	wire w_dff_B_Bb1KFwxw0_2;
	wire w_dff_B_geQLz2po7_2;
	wire w_dff_B_hU03qZzE1_2;
	wire w_dff_B_O0DEJEvc6_2;
	wire w_dff_B_eQ3Uy3G08_2;
	wire w_dff_B_yh7kAaU98_2;
	wire w_dff_B_h74D9eKU0_2;
	wire w_dff_B_f6waqcye3_2;
	wire w_dff_B_q34FxeZk2_2;
	wire w_dff_B_Bf9YOSqe2_2;
	wire w_dff_B_7nlPZ1h67_2;
	wire w_dff_B_XTMmf55n7_2;
	wire w_dff_B_0wG04RyC6_2;
	wire w_dff_B_lsRLi1j21_2;
	wire w_dff_B_6ZCo8SuC1_2;
	wire w_dff_B_g0yROJRG7_2;
	wire w_dff_B_KvTcEe1y7_2;
	wire w_dff_B_V56bjvL51_2;
	wire w_dff_B_O3GCq6kZ7_2;
	wire w_dff_B_ihzPeJjK7_2;
	wire w_dff_B_mYM5gCoF7_2;
	wire w_dff_B_1yDYon1F2_2;
	wire w_dff_B_k8xZ3v2D6_2;
	wire w_dff_B_UDeZe4N71_2;
	wire w_dff_B_wQN9B2v33_2;
	wire w_dff_B_IgagyY0E8_2;
	wire w_dff_B_HrTCHcvK7_2;
	wire w_dff_B_JEOpD9dL1_2;
	wire w_dff_B_wXmlrgGV1_2;
	wire w_dff_B_WvqBDI8O0_2;
	wire w_dff_B_vzhlZg3w8_2;
	wire w_dff_B_NRMato3z0_2;
	wire w_dff_B_ns0dDKnN3_2;
	wire w_dff_B_eLhoSjZo1_2;
	wire w_dff_B_nnGcM5Q27_2;
	wire w_dff_B_bbUPCRWi9_2;
	wire w_dff_B_CbRoJI7X7_2;
	wire w_dff_B_5o1gj5FO1_2;
	wire w_dff_B_3xWtFiSr9_2;
	wire w_dff_B_AtA3bWf96_2;
	wire w_dff_B_Lc401koj9_2;
	wire w_dff_B_yLu2oWlL0_1;
	wire w_dff_B_BKTdhDnF2_2;
	wire w_dff_B_LzXR7G6t2_2;
	wire w_dff_B_0YeTcVzn2_2;
	wire w_dff_B_E5IgPBqR5_2;
	wire w_dff_B_Mn1sDoBt9_2;
	wire w_dff_B_NiGSt4u23_2;
	wire w_dff_B_tLyMQgIP1_2;
	wire w_dff_B_s48nmVZq0_2;
	wire w_dff_B_eC59fv107_2;
	wire w_dff_B_zE3yWCua2_2;
	wire w_dff_B_dVd6AblZ6_2;
	wire w_dff_B_B8bFEOKm6_2;
	wire w_dff_B_CGsZb66e7_2;
	wire w_dff_B_WPMMIjTt1_2;
	wire w_dff_B_FsH3WjZB3_2;
	wire w_dff_B_ibr7ghrX1_2;
	wire w_dff_B_PnAfyQpd1_2;
	wire w_dff_B_rUVhrAsh8_2;
	wire w_dff_B_zUVLmAQs5_2;
	wire w_dff_B_Ka83XLPu8_2;
	wire w_dff_B_nqQDGSgw0_2;
	wire w_dff_B_6Hq6EAjJ8_2;
	wire w_dff_B_fMHUahLR0_2;
	wire w_dff_B_Gzq7vYFc0_2;
	wire w_dff_B_eLFM84gq6_2;
	wire w_dff_B_37kdYW5B6_2;
	wire w_dff_B_ivKCltzi8_2;
	wire w_dff_B_xOdbxLaE6_2;
	wire w_dff_B_pHyen3Vw5_1;
	wire w_dff_B_O4pQZRa68_1;
	wire w_dff_B_VfOPYxpv2_2;
	wire w_dff_B_sjij758H7_2;
	wire w_dff_B_Yr8CD6EF9_2;
	wire w_dff_B_hdpzD2fa8_2;
	wire w_dff_B_WJPSR8797_2;
	wire w_dff_B_Nbpw8GSc4_2;
	wire w_dff_B_ddQWk0ub5_2;
	wire w_dff_B_SGmKyeeq2_2;
	wire w_dff_B_eAeMZbFl5_2;
	wire w_dff_B_ClXnvXk25_2;
	wire w_dff_B_CbyZSHUz2_2;
	wire w_dff_B_tsmT14vq1_2;
	wire w_dff_B_crN3jRC43_2;
	wire w_dff_B_48Iods5x4_2;
	wire w_dff_B_VQxXYS8l8_2;
	wire w_dff_B_RSIiPJIW6_2;
	wire w_dff_B_ow2pnKit8_2;
	wire w_dff_B_oyZ706BL6_2;
	wire w_dff_B_E5yecxaX6_2;
	wire w_dff_B_TpjybKn51_2;
	wire w_dff_B_3zbxahj84_2;
	wire w_dff_B_1CDqRsBU4_2;
	wire w_dff_B_iz3mqyXT3_2;
	wire w_dff_B_Q3bdpMSd8_2;
	wire w_dff_B_YQMQaZxU4_2;
	wire w_dff_B_2Gvn7DMy9_2;
	wire w_dff_B_cbBRVvAf0_2;
	wire w_dff_B_AS76nUfd4_2;
	wire w_dff_B_DFaZJEyd8_2;
	wire w_dff_B_J24kzodN2_2;
	wire w_dff_B_zwzp4V0h1_2;
	wire w_dff_B_5qoBdjaB4_2;
	wire w_dff_B_cKip2Vh62_2;
	wire w_dff_B_PwhUEkCO8_2;
	wire w_dff_B_8Os835gu0_2;
	wire w_dff_B_qtYUzJo82_2;
	wire w_dff_B_MkqOsuV71_2;
	wire w_dff_B_4lpmtRRx0_2;
	wire w_dff_B_0TZ1s0dd0_2;
	wire w_dff_B_Mu6pU7tz2_2;
	wire w_dff_B_D8GY4yPm3_2;
	wire w_dff_B_l4ulICik2_2;
	wire w_dff_B_yNtCmOZx2_2;
	wire w_dff_B_hHLtnYpG6_2;
	wire w_dff_B_CVVMM4nl2_2;
	wire w_dff_B_iN4KO8l51_2;
	wire w_dff_B_nv21DhVX8_2;
	wire w_dff_B_hMGg3jI35_2;
	wire w_dff_B_Gvxw6GEQ6_2;
	wire w_dff_B_ObiDmNgP1_2;
	wire w_dff_B_kiGupozr8_2;
	wire w_dff_B_sF8K7eJt7_2;
	wire w_dff_B_63ITM0IV8_2;
	wire w_dff_B_Nxts0IYw7_1;
	wire w_dff_B_OqXGtk0r7_2;
	wire w_dff_B_Cvja5RD80_2;
	wire w_dff_B_NY42Quuc6_2;
	wire w_dff_B_M7SOeoaH5_2;
	wire w_dff_B_jpgXIRCc1_2;
	wire w_dff_B_tNWJ3hDc2_2;
	wire w_dff_B_eivDyMDw4_2;
	wire w_dff_B_jFIeS7iS5_2;
	wire w_dff_B_tE7sWGt58_2;
	wire w_dff_B_Blo8dg376_2;
	wire w_dff_B_ZAa6HCIe9_2;
	wire w_dff_B_eGeEOhDo8_2;
	wire w_dff_B_c3LSE7Jp7_2;
	wire w_dff_B_7y4iZ9Np2_2;
	wire w_dff_B_2F2XMy2d5_2;
	wire w_dff_B_368IqZiA5_2;
	wire w_dff_B_SB2h7UB99_2;
	wire w_dff_B_cWwLyUxA9_2;
	wire w_dff_B_AvTLrOPv5_2;
	wire w_dff_B_ZUAe7bqy3_2;
	wire w_dff_B_HOAfO1VV0_2;
	wire w_dff_B_0hpV2Lgu2_2;
	wire w_dff_B_iDM6MtEK6_2;
	wire w_dff_B_cW7nfghM3_2;
	wire w_dff_B_PSOlWlRS9_1;
	wire w_dff_B_kUPrBYtM2_1;
	wire w_dff_B_nYbFUOK69_2;
	wire w_dff_B_ArXbxpJ25_2;
	wire w_dff_B_KTvJJh0v9_2;
	wire w_dff_B_MarX1VX68_2;
	wire w_dff_B_8RpZfeWw6_2;
	wire w_dff_B_F31DFCFA2_2;
	wire w_dff_B_w9m4zXIC9_2;
	wire w_dff_B_wDvJF5NS0_2;
	wire w_dff_B_BBLwHwkQ8_2;
	wire w_dff_B_UuwrVsM92_2;
	wire w_dff_B_EpoIowCu8_2;
	wire w_dff_B_ia5N8OXy8_2;
	wire w_dff_B_Pn8Pv91D0_2;
	wire w_dff_B_svcJVEXU4_2;
	wire w_dff_B_bdYi72WB1_2;
	wire w_dff_B_3TUxJHuE5_2;
	wire w_dff_B_2eJcINEF6_2;
	wire w_dff_B_uV5GGtDX8_2;
	wire w_dff_B_vUkUamBW4_2;
	wire w_dff_B_nDOtVjXs8_2;
	wire w_dff_B_y2SyWNyp8_2;
	wire w_dff_B_OAWrp7nW6_2;
	wire w_dff_B_cc8BGGwY9_2;
	wire w_dff_B_Gx5uZHb87_2;
	wire w_dff_B_XDhq4FBF6_2;
	wire w_dff_B_OfWoQqJH2_2;
	wire w_dff_B_BR4Tjjvr4_2;
	wire w_dff_B_ZaHkSOZg9_2;
	wire w_dff_B_w5vKRf4Z8_2;
	wire w_dff_B_iKbfZKgF7_2;
	wire w_dff_B_Q9IKnMa38_2;
	wire w_dff_B_CQX2jHmG3_2;
	wire w_dff_B_f63iPIcQ4_2;
	wire w_dff_B_38x8kn8X4_2;
	wire w_dff_B_C0vKHX3G1_2;
	wire w_dff_B_hIz0nFUS3_2;
	wire w_dff_B_geBw50nT9_2;
	wire w_dff_B_lKA6DX5k0_2;
	wire w_dff_B_YsxI9lXF3_2;
	wire w_dff_B_vNTh4RgE6_2;
	wire w_dff_B_kEIsEVAr4_2;
	wire w_dff_B_8wSfaBW14_2;
	wire w_dff_B_fNZgH5Ia3_2;
	wire w_dff_B_gF9ti5EF3_2;
	wire w_dff_B_1XAPDj0M1_2;
	wire w_dff_B_0bFHJie74_1;
	wire w_dff_B_4UY19m043_2;
	wire w_dff_B_d9XBYaqX8_2;
	wire w_dff_B_YVabvJQa1_2;
	wire w_dff_B_eC30aI6f6_2;
	wire w_dff_B_CPXcp7ny7_2;
	wire w_dff_B_6dNqTBbT2_2;
	wire w_dff_B_Q5O0HqW16_2;
	wire w_dff_B_efNjonfQ7_2;
	wire w_dff_B_iDnnnMfs1_2;
	wire w_dff_B_fYOrmObb1_2;
	wire w_dff_B_jYhlo0RK9_2;
	wire w_dff_B_o96tmtMv2_2;
	wire w_dff_B_tggmTTTF3_2;
	wire w_dff_B_IbjrAGqq9_2;
	wire w_dff_B_u5zh3mSe2_2;
	wire w_dff_B_MjBcxu072_2;
	wire w_dff_B_eUTUXKbM1_2;
	wire w_dff_B_Ffqu1yuv3_2;
	wire w_dff_B_3qWJqvg82_2;
	wire w_dff_B_jfnFqI8W0_2;
	wire w_dff_B_IUJTneI48_1;
	wire w_dff_B_O9rLtxNu0_1;
	wire w_dff_B_Yo4NJgHU9_2;
	wire w_dff_B_nAYduoFH1_2;
	wire w_dff_B_uASePRO83_2;
	wire w_dff_B_4faQDMdp3_2;
	wire w_dff_B_CPE5SUUB5_2;
	wire w_dff_B_IM3GGFyb2_2;
	wire w_dff_B_BbHgMiGc9_2;
	wire w_dff_B_uY2zE2uQ1_2;
	wire w_dff_B_bCKBVgiw5_2;
	wire w_dff_B_OUade5p45_2;
	wire w_dff_B_urKKBo6M9_2;
	wire w_dff_B_4o4OIB594_2;
	wire w_dff_B_6WX05CD52_2;
	wire w_dff_B_xw50NHlM0_2;
	wire w_dff_B_dmkToIFs6_2;
	wire w_dff_B_7eMuuLbb2_2;
	wire w_dff_B_id4ZkbFR2_2;
	wire w_dff_B_vnMnEEWT2_2;
	wire w_dff_B_sbjTJYux0_2;
	wire w_dff_B_BVFSdiRn2_2;
	wire w_dff_B_O2Pq2xS98_2;
	wire w_dff_B_yWAG5Exw1_2;
	wire w_dff_B_7ON9MR2A7_2;
	wire w_dff_B_hRAbzofl0_2;
	wire w_dff_B_vAjlP61A0_2;
	wire w_dff_B_GUiXVbHH3_2;
	wire w_dff_B_2pkieY3j1_2;
	wire w_dff_B_6MkznyUo3_2;
	wire w_dff_B_TJrw2N5p9_2;
	wire w_dff_B_2kvg4Fv99_2;
	wire w_dff_B_nVoxdnes2_2;
	wire w_dff_B_D5utOWhA6_2;
	wire w_dff_B_jF5xRy7D9_2;
	wire w_dff_B_Kmmi47nv6_2;
	wire w_dff_B_LC3BOYRO6_2;
	wire w_dff_B_R1ismnub3_2;
	wire w_dff_B_3mVv4DRR9_1;
	wire w_dff_B_IWHhk4Ln3_2;
	wire w_dff_B_leddj2aF4_2;
	wire w_dff_B_8rkaynPQ6_2;
	wire w_dff_B_sijKPjN28_2;
	wire w_dff_B_K5YNOlXo8_2;
	wire w_dff_B_M3BiYllW4_2;
	wire w_dff_B_QSITtQkT5_2;
	wire w_dff_B_R0G6dGWk8_2;
	wire w_dff_B_378IHsSa2_2;
	wire w_dff_B_ZG6YCjww7_2;
	wire w_dff_B_tOv6AX2j9_2;
	wire w_dff_B_K0hzm4e26_2;
	wire w_dff_B_I5UfBLWq2_2;
	wire w_dff_B_m2EJuf2V9_2;
	wire w_dff_B_2gu2iADJ0_2;
	wire w_dff_B_elEvupHo3_2;
	wire w_dff_B_AteBDex17_2;
	wire w_dff_B_PKQSLXiP0_2;
	wire w_dff_B_z3lkp7JR6_1;
	wire w_dff_B_CSsJu4ca9_1;
	wire w_dff_B_Xo2BpnRW5_2;
	wire w_dff_B_5XQ0nrF35_2;
	wire w_dff_B_qEXWvxh97_2;
	wire w_dff_B_ZQJPXZFV5_2;
	wire w_dff_B_5IxobdZq5_2;
	wire w_dff_B_Jcy3oZuD4_2;
	wire w_dff_B_sYLgovAu7_2;
	wire w_dff_B_IZ6bZz6v2_2;
	wire w_dff_B_zrOP94kH2_2;
	wire w_dff_B_zompo2d58_2;
	wire w_dff_B_7lUNFWuT8_2;
	wire w_dff_B_usv94h986_2;
	wire w_dff_B_W5C7l31p9_2;
	wire w_dff_B_qEfu1ZfZ0_2;
	wire w_dff_B_ZkRmFNuL2_2;
	wire w_dff_B_VeaPsWuT4_2;
	wire w_dff_B_3lEBNQst8_2;
	wire w_dff_B_wcFO4hM45_2;
	wire w_dff_B_WJpZxDEC1_2;
	wire w_dff_B_E037uTcI2_2;
	wire w_dff_B_Jhkh5mMR1_2;
	wire w_dff_B_UK9mqZU10_2;
	wire w_dff_B_avWyTI751_2;
	wire w_dff_B_GC9wIpFz2_2;
	wire w_dff_B_EIgSh8By8_2;
	wire w_dff_B_tysjgboV3_2;
	wire w_dff_B_0d5u6kvY2_2;
	wire w_dff_B_E3ivLrTe7_2;
	wire w_dff_B_zd2kEF9W7_1;
	wire w_dff_B_uDJOOt0d7_2;
	wire w_dff_B_0nOHOJjq5_2;
	wire w_dff_B_IDCpIKvz6_2;
	wire w_dff_B_74qhtc2l4_2;
	wire w_dff_B_lyUkxFj24_2;
	wire w_dff_B_ezwYcDka4_2;
	wire w_dff_B_ikgVUA8i4_2;
	wire w_dff_B_D1X70OjW9_2;
	wire w_dff_B_tVvhSEI03_2;
	wire w_dff_B_FaPaHFCc3_2;
	wire w_dff_B_q11e93fA8_2;
	wire w_dff_B_CHQM5nyO9_2;
	wire w_dff_B_yAJlfnKR7_2;
	wire w_dff_B_7AgCoNZE4_2;
	wire w_dff_B_XS4WX4E57_2;
	wire w_dff_B_RkzEbBhT9_2;
	wire w_dff_B_bIQlvcg20_1;
	wire w_dff_B_Gjt8d74j1_1;
	wire w_dff_B_LXYLAeB95_2;
	wire w_dff_B_0n2a2h1X1_2;
	wire w_dff_B_wFXnMAqk6_2;
	wire w_dff_B_CXqwzez22_2;
	wire w_dff_B_f59dO4s58_2;
	wire w_dff_B_AVFPRMmi6_2;
	wire w_dff_B_w8A3RxER3_2;
	wire w_dff_B_l1bbskJE9_2;
	wire w_dff_B_Wjv0KT8C0_2;
	wire w_dff_B_WhlOOeS69_2;
	wire w_dff_B_IVbFDPnX4_2;
	wire w_dff_B_bXLmwg2S1_2;
	wire w_dff_B_ERRyIOcK5_2;
	wire w_dff_B_7GO5bWIN1_2;
	wire w_dff_B_Lz2fwbes8_2;
	wire w_dff_B_ZCvR93kx6_2;
	wire w_dff_B_xz6pQ6NE1_2;
	wire w_dff_B_bUScqbrk2_2;
	wire w_dff_B_4HW70j5j1_2;
	wire w_dff_B_WfUqXEjd0_2;
	wire w_dff_B_Ufyikq8N9_1;
	wire w_dff_B_UveMoWF14_2;
	wire w_dff_B_ulyTI7Oq7_2;
	wire w_dff_B_OnKaUG1J7_2;
	wire w_dff_B_hNzvNxiS0_2;
	wire w_dff_B_3vonbvKI4_2;
	wire w_dff_B_2PgK952V4_2;
	wire w_dff_B_bF404Jso3_2;
	wire w_dff_B_9Lzn0eOn5_2;
	wire w_dff_B_SsUnkEGl2_2;
	wire w_dff_B_ScpWsRMN6_2;
	wire w_dff_B_REPYmE8F0_2;
	wire w_dff_B_SuelSZ3s7_2;
	wire w_dff_B_4160zYfZ2_2;
	wire w_dff_B_VcfgjPsI0_2;
	wire w_dff_B_GlaY8Bbk6_2;
	wire w_dff_B_T3ULk5nn6_2;
	wire w_dff_B_mcsrWnJK6_2;
	wire w_dff_B_NbWDpy8r7_2;
	wire w_dff_B_XKFgzDIA2_2;
	wire w_dff_B_eBmO4flu4_2;
	wire w_dff_B_6YAPjww34_2;
	wire w_dff_B_eadTlS2A1_2;
	wire w_dff_B_H8eNOtfX5_2;
	wire w_dff_B_TZmvMU6P3_2;
	wire w_dff_B_91W0zb4V7_2;
	wire w_dff_B_WKGtY2ml4_2;
	wire w_dff_B_vjml4cqS8_1;
	wire w_dff_B_KpVUuAJN5_2;
	wire w_dff_B_w9jauQoR8_2;
	wire w_dff_B_EaHDlXP45_2;
	wire w_dff_B_m8IARHne9_2;
	wire w_dff_B_SJ9DI1s79_2;
	wire w_dff_B_8CrwbxYA8_2;
	wire w_dff_B_Ttx1IJNK3_2;
	wire w_dff_B_mRin9tCy3_2;
	wire w_dff_B_tDITpW1u6_2;
	wire w_dff_B_3e9rjiZe8_2;
	wire w_dff_B_cLrWZABO6_2;
	wire w_dff_B_GaJSvwO06_2;
	wire w_dff_B_gMd2PrvX8_2;
	wire w_dff_B_kc3LZIYa9_2;
	wire w_dff_B_gOT3hRON5_2;
	wire w_dff_A_mBmYYDfz3_0;
	wire w_dff_A_9NCxbHb42_0;
	wire w_dff_A_UX8pD6aF4_0;
	wire w_dff_B_mbQs6htz1_2;
	wire w_dff_A_Y79VpmHU5_0;
	wire w_dff_A_7r8RQZfT3_0;
	wire w_dff_A_cs9E2wFq9_0;
	wire w_dff_B_2jQ3RK4d0_2;
	wire w_dff_A_XBZdRkvs1_0;
	wire w_dff_A_BkdLtBcM6_0;
	wire w_dff_B_lXjMKyo05_2;
	wire w_dff_B_JasEiltx4_2;
	wire w_dff_B_Q2iIP7Qg7_2;
	wire w_dff_A_ooBIzX3Q9_1;
	wire w_dff_A_ooalAoq50_0;
	wire w_dff_A_DSr6ENMU4_0;
	wire w_dff_A_wNznkkHX1_0;
	wire w_dff_A_FrQBhmAr8_0;
	wire w_dff_A_Hhbenz899_0;
	wire w_dff_A_NxH2jbQk7_0;
	wire w_dff_A_TLX1PWnh2_0;
	wire w_dff_A_sN2TyrCa8_0;
	wire w_dff_A_K0FvvkJp9_0;
	wire w_dff_A_LifDZLrE0_0;
	wire w_dff_A_N06ojCkr9_0;
	wire w_dff_A_PY0KxP1a2_0;
	wire w_dff_A_wJFNUXW48_0;
	wire w_dff_A_5iBuQOlB0_0;
	wire w_dff_A_BlHXVJON3_0;
	wire w_dff_A_cnCqwNHi6_0;
	wire w_dff_A_GzQiZkhL6_0;
	wire w_dff_A_Wwvneifu8_0;
	wire w_dff_A_KkzAZReB7_0;
	wire w_dff_A_p1jrxzGC0_0;
	wire w_dff_A_qwlMhPvA7_0;
	wire w_dff_A_zhrHWjME2_0;
	wire w_dff_A_KNVu0Ji99_0;
	wire w_dff_A_JmNUEczm9_0;
	wire w_dff_A_m0nE4OuU7_0;
	wire w_dff_A_BxmNwcYk5_0;
	wire w_dff_A_3k6zDv6d1_0;
	wire w_dff_A_URc29qnp7_0;
	wire w_dff_A_3hSDRLeS9_0;
	wire w_dff_A_fV559tTN4_0;
	wire w_dff_A_471LQcjL6_0;
	wire w_dff_A_j16ILcqv7_0;
	wire w_dff_A_xQF2nmdq4_0;
	wire w_dff_A_9JTXxx1I4_0;
	wire w_dff_A_ZxzDFWJl7_0;
	wire w_dff_A_ChmJP1dU7_0;
	wire w_dff_A_Xr4LdzK80_0;
	wire w_dff_A_JccgSi2u0_0;
	wire w_dff_A_8OcIxksp1_0;
	wire w_dff_A_QuCUHEMZ8_0;
	wire w_dff_A_fdOsw1VI3_0;
	wire w_dff_A_SdXJdlXV0_0;
	wire w_dff_A_cb5J6VfX0_0;
	wire w_dff_A_oDRamxAK6_0;
	wire w_dff_A_HxYkZiuK6_0;
	wire w_dff_A_eeamE3s85_0;
	wire w_dff_A_rVm0TM4c4_0;
	wire w_dff_A_XY5LdrhZ4_0;
	wire w_dff_A_dTmWJk0V3_0;
	wire w_dff_A_tbuDP5oc9_0;
	wire w_dff_A_pFkx1aAh1_0;
	wire w_dff_A_rYeUySUg9_0;
	wire w_dff_A_YfJtFXKK6_0;
	wire w_dff_A_7EWBmJsn3_0;
	wire w_dff_A_hRb4Uy4R2_0;
	wire w_dff_A_1MBESbvS7_0;
	wire w_dff_A_4iKiaaya0_0;
	wire w_dff_A_tPAHFVZ62_0;
	wire w_dff_A_fyTdke9w0_0;
	wire w_dff_A_sPx8JKZc8_0;
	wire w_dff_A_BefKe4R87_0;
	wire w_dff_A_F2E10s9i9_0;
	wire w_dff_A_gXzTkQsB0_0;
	wire w_dff_A_KV3yWYH62_0;
	wire w_dff_A_b4sTED5r7_0;
	wire w_dff_A_kEVgXev02_0;
	wire w_dff_A_wOJOhcwG3_0;
	wire w_dff_A_twS3z4Md7_0;
	wire w_dff_A_c6JWTf9y6_0;
	wire w_dff_A_BEn3V9Gl9_0;
	wire w_dff_A_YYHzYWnv7_0;
	wire w_dff_A_xsrUDg8Q4_0;
	wire w_dff_A_d5AloKRx0_0;
	wire w_dff_A_ERwqQcch6_2;
	wire w_dff_A_n9GB75JS3_0;
	wire w_dff_A_hHvtGTlQ8_0;
	wire w_dff_A_AnFkQSy58_0;
	wire w_dff_A_alQvqies3_0;
	wire w_dff_A_NTsj793Y3_0;
	wire w_dff_A_UdfStCmJ6_0;
	wire w_dff_A_M5Gc7Mn44_0;
	wire w_dff_A_ZoPEDEal0_0;
	wire w_dff_A_MmoN4ZXN2_0;
	wire w_dff_A_GvgcWzc66_0;
	wire w_dff_A_CopCHs636_0;
	wire w_dff_A_j2VkvqY69_0;
	wire w_dff_A_hSgVIXjW7_0;
	wire w_dff_A_j2ztsuy43_0;
	wire w_dff_A_v62F2IWC7_0;
	wire w_dff_A_6mpWp5Zf8_0;
	wire w_dff_A_tdtMLX1A3_0;
	wire w_dff_A_2bhDzNnD9_0;
	wire w_dff_A_HBngTINL3_0;
	wire w_dff_A_44ZYftsj8_0;
	wire w_dff_A_1T0wmQ9Q7_0;
	wire w_dff_A_uwwWCaAN5_0;
	wire w_dff_A_OOVUengi4_0;
	wire w_dff_A_RiNYpsUZ4_0;
	wire w_dff_A_pAz4n5Ij9_0;
	wire w_dff_A_2OUaKl2z8_0;
	wire w_dff_A_ji4ZwdNe3_0;
	wire w_dff_A_LEi7ziF49_0;
	wire w_dff_A_hHqfrAqe9_0;
	wire w_dff_A_iafQQNhc1_0;
	wire w_dff_A_qqEazY6k9_0;
	wire w_dff_A_Zjv5WxxK8_0;
	wire w_dff_A_QStrNx3z2_0;
	wire w_dff_A_iWUXfyjK0_0;
	wire w_dff_A_QHqd1eQe9_0;
	wire w_dff_A_s5bR2fBA6_0;
	wire w_dff_A_7CjraK4O8_0;
	wire w_dff_A_sra1MCyW3_0;
	wire w_dff_A_NqVRCeBe6_0;
	wire w_dff_A_gewLgLH49_0;
	wire w_dff_A_yeUuBgYH3_0;
	wire w_dff_A_e5RL9Fr17_0;
	wire w_dff_A_vkcrJACS5_0;
	wire w_dff_A_FvGyzLDv6_0;
	wire w_dff_A_ynJToruf2_0;
	wire w_dff_A_ibkW8z117_0;
	wire w_dff_A_xQSrxj0P4_0;
	wire w_dff_A_us00chUJ7_0;
	wire w_dff_A_v1nt2IXZ5_0;
	wire w_dff_A_B2YdVD7m5_0;
	wire w_dff_A_fBkfM7Dk9_0;
	wire w_dff_A_T9ce9Asc0_0;
	wire w_dff_A_yLpw7GaN3_0;
	wire w_dff_A_Zr3ERBvI4_0;
	wire w_dff_A_xcp2VARa5_0;
	wire w_dff_A_zVbkba7S3_0;
	wire w_dff_A_sepVj1Tp8_0;
	wire w_dff_A_22FGuTkW5_0;
	wire w_dff_A_sVhuT3xV8_0;
	wire w_dff_A_e975MbsB1_0;
	wire w_dff_A_l2UfLZWH9_0;
	wire w_dff_A_KRDcwiQT3_0;
	wire w_dff_A_U8omtxaO8_0;
	wire w_dff_A_5AqRMy096_0;
	wire w_dff_A_cnOOCoKZ5_0;
	wire w_dff_A_TBTHLLdM3_0;
	wire w_dff_A_cZdjRu643_0;
	wire w_dff_A_8e6dsy809_0;
	wire w_dff_A_v9hUv4tu3_0;
	wire w_dff_A_JVhOTcac7_2;
	wire w_dff_A_NT76UVWY5_0;
	wire w_dff_A_824KkLKS4_0;
	wire w_dff_A_fMtPH8fD4_0;
	wire w_dff_A_VJyafekE9_0;
	wire w_dff_A_ID3HfpM18_0;
	wire w_dff_A_Xa9r3keL2_0;
	wire w_dff_A_fGqx4EVW3_0;
	wire w_dff_A_u5QbZPUF0_0;
	wire w_dff_A_e9Mq2UPP9_0;
	wire w_dff_A_HhxrEXQQ2_0;
	wire w_dff_A_Gnnlkr3h1_0;
	wire w_dff_A_pUiflOiD1_0;
	wire w_dff_A_2lKeuyZs8_0;
	wire w_dff_A_NFITlDAY8_0;
	wire w_dff_A_hNdIgJyg0_0;
	wire w_dff_A_7CtlbZyX5_0;
	wire w_dff_A_8hqeXyt36_0;
	wire w_dff_A_133QnD3y4_0;
	wire w_dff_A_tGlBxxaP5_0;
	wire w_dff_A_D0bWv7nh6_0;
	wire w_dff_A_KBQxncBm3_0;
	wire w_dff_A_07Znfa8p1_0;
	wire w_dff_A_UhdnXtKU9_0;
	wire w_dff_A_WmTEDsOs8_0;
	wire w_dff_A_1xzJKcZs7_0;
	wire w_dff_A_QTjy2HHt2_0;
	wire w_dff_A_ngxFGTSy8_0;
	wire w_dff_A_Kwl2yqEI4_0;
	wire w_dff_A_fqgXS9d36_0;
	wire w_dff_A_97CxQrb70_0;
	wire w_dff_A_tYGfJabt2_0;
	wire w_dff_A_wkMNkgim6_0;
	wire w_dff_A_xNUMPrWg3_0;
	wire w_dff_A_0RGdBZxN3_0;
	wire w_dff_A_kFROo3MS8_0;
	wire w_dff_A_WdROrC0j6_0;
	wire w_dff_A_Ej6knU7C6_0;
	wire w_dff_A_68COWNWm6_0;
	wire w_dff_A_Fs6yXC0n1_0;
	wire w_dff_A_FcdE4FeK9_0;
	wire w_dff_A_8UgCSxG51_0;
	wire w_dff_A_sXMumqT44_0;
	wire w_dff_A_0HM10aIA2_0;
	wire w_dff_A_8FeN6LaS6_0;
	wire w_dff_A_x1E0F7KP0_0;
	wire w_dff_A_YjWzstNl3_0;
	wire w_dff_A_ZXNeWPsI9_0;
	wire w_dff_A_C4jqsiD09_0;
	wire w_dff_A_aiXV3y6k9_0;
	wire w_dff_A_PiXCjjyt8_0;
	wire w_dff_A_FIhdjpn42_0;
	wire w_dff_A_psrtXOYz5_0;
	wire w_dff_A_Inpql7wC1_0;
	wire w_dff_A_uqk1M2Gx6_0;
	wire w_dff_A_Q2CUbeza0_0;
	wire w_dff_A_g0oU4rgc8_0;
	wire w_dff_A_gDlYcnpp3_0;
	wire w_dff_A_p0MP5Sde4_0;
	wire w_dff_A_Q8nhhH208_0;
	wire w_dff_A_9LIkbH8r7_0;
	wire w_dff_A_xOmjsfo56_0;
	wire w_dff_A_fpXNrvut3_0;
	wire w_dff_A_yEu7myOq6_0;
	wire w_dff_A_I7iEgpZ91_0;
	wire w_dff_A_TFyM6XWr9_0;
	wire w_dff_A_170TZJca6_0;
	wire w_dff_A_omAAnoaQ4_0;
	wire w_dff_A_Ipkfrq3U1_0;
	wire w_dff_A_1yMaWZic3_2;
	wire w_dff_A_8X9du1RG9_0;
	wire w_dff_A_rFVpRbud2_0;
	wire w_dff_A_ErdpTLjR2_0;
	wire w_dff_A_s05MepAb6_0;
	wire w_dff_A_TWufy2BV1_0;
	wire w_dff_A_x4kecnmA0_0;
	wire w_dff_A_KyKEaOsH1_0;
	wire w_dff_A_PrEVD5yV7_0;
	wire w_dff_A_b0TfVYAn0_0;
	wire w_dff_A_IbuQTzem8_0;
	wire w_dff_A_R8NDF07a2_0;
	wire w_dff_A_JElYusPA3_0;
	wire w_dff_A_CFpjbw0M6_0;
	wire w_dff_A_jENwXvRN6_0;
	wire w_dff_A_Re96E3ou3_0;
	wire w_dff_A_Yvw7I55z3_0;
	wire w_dff_A_SY9Td5QQ8_0;
	wire w_dff_A_cjVJyWL80_0;
	wire w_dff_A_xY6YpDOM2_0;
	wire w_dff_A_wzuAUU8H2_0;
	wire w_dff_A_8JLkeZUI0_0;
	wire w_dff_A_uheqYr9h6_0;
	wire w_dff_A_iVzxobba6_0;
	wire w_dff_A_GMDtooMm0_0;
	wire w_dff_A_8gG22on23_0;
	wire w_dff_A_igzkPXVb7_0;
	wire w_dff_A_RMxLWcNl9_0;
	wire w_dff_A_vIpiASBy9_0;
	wire w_dff_A_WV4kVZTz5_0;
	wire w_dff_A_oAmK9mjk3_0;
	wire w_dff_A_Ar1CFKkr3_0;
	wire w_dff_A_gAgW4Gp38_0;
	wire w_dff_A_L782zogU6_0;
	wire w_dff_A_q47g306l8_0;
	wire w_dff_A_vcwRjrh79_0;
	wire w_dff_A_PHocqwJc6_0;
	wire w_dff_A_xBN6Utg09_0;
	wire w_dff_A_sggvOKUn2_0;
	wire w_dff_A_4AZEIa1j1_0;
	wire w_dff_A_j2Rwxy2r9_0;
	wire w_dff_A_TKYfrazv0_0;
	wire w_dff_A_77NnLVCI7_0;
	wire w_dff_A_BeqkVDrE2_0;
	wire w_dff_A_ZPJpWdwx2_0;
	wire w_dff_A_X2SBdZSj6_0;
	wire w_dff_A_uUOBhka81_0;
	wire w_dff_A_iRgeIgQo3_0;
	wire w_dff_A_KcS4N9bR1_0;
	wire w_dff_A_VwK39ooS6_0;
	wire w_dff_A_16XwVVWG5_0;
	wire w_dff_A_wbdI8snT1_0;
	wire w_dff_A_irtJAX4c7_0;
	wire w_dff_A_Yr0yTxxK8_0;
	wire w_dff_A_JkE0mIGb2_0;
	wire w_dff_A_vtt15bAz7_0;
	wire w_dff_A_Lusgj4m97_0;
	wire w_dff_A_PNV4wddq2_0;
	wire w_dff_A_ViDl5Bzk1_0;
	wire w_dff_A_IMNEaPK70_0;
	wire w_dff_A_udqJLdeb9_0;
	wire w_dff_A_ryLHRJvm6_0;
	wire w_dff_A_lLEhQVjI2_0;
	wire w_dff_A_CxReM8mW6_0;
	wire w_dff_A_0FjEIobv2_0;
	wire w_dff_A_lY17I36C2_0;
	wire w_dff_A_THDtcXMv5_2;
	wire w_dff_A_ODbkMDGw9_0;
	wire w_dff_A_yzRjjQb78_0;
	wire w_dff_A_nx7lV8ZY8_0;
	wire w_dff_A_6GBtMk3S7_0;
	wire w_dff_A_t4n3Vxnp3_0;
	wire w_dff_A_gnWkttWm2_0;
	wire w_dff_A_Ws57iV842_0;
	wire w_dff_A_IyKUKQ4n2_0;
	wire w_dff_A_mcq8eNv20_0;
	wire w_dff_A_XRGRVtm78_0;
	wire w_dff_A_qXiDv2w52_0;
	wire w_dff_A_MUAd3p4d7_0;
	wire w_dff_A_EAaQ7z5e5_0;
	wire w_dff_A_BpGXNOAY0_0;
	wire w_dff_A_g7OYbm2x0_0;
	wire w_dff_A_xHo15xPE7_0;
	wire w_dff_A_gpvHEGao3_0;
	wire w_dff_A_aUF0kOJh8_0;
	wire w_dff_A_Kj8vqFVc2_0;
	wire w_dff_A_BKloISGC6_0;
	wire w_dff_A_Zvmu7Wwi2_0;
	wire w_dff_A_fyaRnmnx2_0;
	wire w_dff_A_Ay3fC7ts7_0;
	wire w_dff_A_hCAdJnNv5_0;
	wire w_dff_A_pPlhb8708_0;
	wire w_dff_A_WbSZbNhz6_0;
	wire w_dff_A_oWvcKqrA4_0;
	wire w_dff_A_WW2TlCyv3_0;
	wire w_dff_A_f8uAFxet7_0;
	wire w_dff_A_1pdyoYeS8_0;
	wire w_dff_A_QD0p07Am6_0;
	wire w_dff_A_d8P6ylwF7_0;
	wire w_dff_A_Lgm8zHoN0_0;
	wire w_dff_A_6t3link02_0;
	wire w_dff_A_8d8p2Gyi8_0;
	wire w_dff_A_hoTGXh7o0_0;
	wire w_dff_A_AB0CsfNW1_0;
	wire w_dff_A_seXohdPi0_0;
	wire w_dff_A_mTmIwOWB9_0;
	wire w_dff_A_Po82cIcz8_0;
	wire w_dff_A_NFQrKPGr7_0;
	wire w_dff_A_x1aK2mS70_0;
	wire w_dff_A_2eaFZj3w8_0;
	wire w_dff_A_zFNlT83p8_0;
	wire w_dff_A_tqjlsVox0_0;
	wire w_dff_A_yIwuicAw7_0;
	wire w_dff_A_0x4CTKnf7_0;
	wire w_dff_A_0rSnzzPj4_0;
	wire w_dff_A_a2LNhgPD4_0;
	wire w_dff_A_dqVEAAbu3_0;
	wire w_dff_A_DCuBdoDz4_0;
	wire w_dff_A_7Pu2h7lu1_0;
	wire w_dff_A_qQnBUnhz3_0;
	wire w_dff_A_4O8ace7l1_0;
	wire w_dff_A_gyS4asOc8_0;
	wire w_dff_A_MJqVFwi67_0;
	wire w_dff_A_fFFvfhWN2_0;
	wire w_dff_A_xie6wb2G0_0;
	wire w_dff_A_TLjKRVch2_0;
	wire w_dff_A_pNp79i8V9_0;
	wire w_dff_A_wXRBSrFY6_0;
	wire w_dff_A_3sQIG0Ov2_0;
	wire w_dff_A_w3mHM9Py5_2;
	wire w_dff_A_JakqqeV08_0;
	wire w_dff_A_SesUIdQv5_0;
	wire w_dff_A_4E6N3AQ14_0;
	wire w_dff_A_zxi2NWyo2_0;
	wire w_dff_A_7xLM1DEP4_0;
	wire w_dff_A_5m0orVSO7_0;
	wire w_dff_A_yIZrjeEn3_0;
	wire w_dff_A_Vpdpc3n28_0;
	wire w_dff_A_42hxcsI41_0;
	wire w_dff_A_b867YtuE9_0;
	wire w_dff_A_S0yvhFAL4_0;
	wire w_dff_A_S5gYA1oS1_0;
	wire w_dff_A_IZl7vllN8_0;
	wire w_dff_A_GnplEB9y1_0;
	wire w_dff_A_6t176Plu5_0;
	wire w_dff_A_uPyWJ8VS5_0;
	wire w_dff_A_gwWJWCzu0_0;
	wire w_dff_A_pfsJhVjh9_0;
	wire w_dff_A_OEn9XMKV7_0;
	wire w_dff_A_hByr6STF4_0;
	wire w_dff_A_n4IIHgRg9_0;
	wire w_dff_A_XVww6zG93_0;
	wire w_dff_A_15Khhkqz1_0;
	wire w_dff_A_pkr9Ey5o5_0;
	wire w_dff_A_8oemvZsB0_0;
	wire w_dff_A_tHo5P9X98_0;
	wire w_dff_A_1itXeHyd3_0;
	wire w_dff_A_B8cJIMHg6_0;
	wire w_dff_A_c5FiU9ow1_0;
	wire w_dff_A_W3nfsRFu4_0;
	wire w_dff_A_EutsRKl33_0;
	wire w_dff_A_HqVcCpro5_0;
	wire w_dff_A_p5cCwLaK2_0;
	wire w_dff_A_TwB8fXxc6_0;
	wire w_dff_A_oe575g4w7_0;
	wire w_dff_A_B5eLN9NM1_0;
	wire w_dff_A_65Yafg4d4_0;
	wire w_dff_A_DqSOxroJ5_0;
	wire w_dff_A_iE3Vw3Mv5_0;
	wire w_dff_A_V0pYOB5p6_0;
	wire w_dff_A_ioLgQfr38_0;
	wire w_dff_A_vE0OYVYI0_0;
	wire w_dff_A_PTniF9K56_0;
	wire w_dff_A_Sw2QX1vV9_0;
	wire w_dff_A_YMOXujyN8_0;
	wire w_dff_A_2xejjWoa4_0;
	wire w_dff_A_xISFREAK2_0;
	wire w_dff_A_RiW9sP6b9_0;
	wire w_dff_A_Iz342MBE6_0;
	wire w_dff_A_QaB235Zq1_0;
	wire w_dff_A_x2WhwkiH1_0;
	wire w_dff_A_RAtZtlxT2_0;
	wire w_dff_A_16GcYN2g3_0;
	wire w_dff_A_6FrJqOY24_0;
	wire w_dff_A_wNfL901z5_0;
	wire w_dff_A_B1di4oAW9_0;
	wire w_dff_A_tg7uLbtY4_0;
	wire w_dff_A_f5r53jkt1_0;
	wire w_dff_A_pDzvdEB44_0;
	wire w_dff_A_QxM6dCu23_2;
	wire w_dff_A_e01wDhmm2_0;
	wire w_dff_A_71V0GWoh3_0;
	wire w_dff_A_QP9mgEJw6_0;
	wire w_dff_A_q9ky4FRJ8_0;
	wire w_dff_A_34nH5grt4_0;
	wire w_dff_A_3YMOdVJu1_0;
	wire w_dff_A_QsP3bsdy1_0;
	wire w_dff_A_imBaBLJ17_0;
	wire w_dff_A_5mat9fLD2_0;
	wire w_dff_A_Txf3lufu9_0;
	wire w_dff_A_IFFby4vZ6_0;
	wire w_dff_A_cxD9eBeh3_0;
	wire w_dff_A_6yLmLBFt0_0;
	wire w_dff_A_0Idnk2Po7_0;
	wire w_dff_A_qgxjHXtH5_0;
	wire w_dff_A_u9Cu1s053_0;
	wire w_dff_A_2KA2uSxb2_0;
	wire w_dff_A_eMHFlnZR8_0;
	wire w_dff_A_KwjGTL4p3_0;
	wire w_dff_A_LAPk2opK5_0;
	wire w_dff_A_ihZeLB9x2_0;
	wire w_dff_A_HjWGw5N04_0;
	wire w_dff_A_ZOF2eZb34_0;
	wire w_dff_A_NpPYNAmR8_0;
	wire w_dff_A_Jp2DZEsI4_0;
	wire w_dff_A_ALE353iQ5_0;
	wire w_dff_A_W5LgvVxC7_0;
	wire w_dff_A_KXqU0ZAF2_0;
	wire w_dff_A_tK7Da9dN1_0;
	wire w_dff_A_BKfJM7F47_0;
	wire w_dff_A_Gt0mGzhN3_0;
	wire w_dff_A_JnAzQUn49_0;
	wire w_dff_A_i90H7wnC5_0;
	wire w_dff_A_txonvOJh0_0;
	wire w_dff_A_h0Np84wX3_0;
	wire w_dff_A_5b33Sm3G3_0;
	wire w_dff_A_zsL0Qf338_0;
	wire w_dff_A_ZLXs3Jm23_0;
	wire w_dff_A_b4ZMHgzr0_0;
	wire w_dff_A_6UvraaLu0_0;
	wire w_dff_A_x5mWSqiO5_0;
	wire w_dff_A_YsUpNSSN9_0;
	wire w_dff_A_uempqmzs8_0;
	wire w_dff_A_S6X3TZmz0_0;
	wire w_dff_A_gYSrY5SC0_0;
	wire w_dff_A_zMZZJ41B4_0;
	wire w_dff_A_mYWVpp0j7_0;
	wire w_dff_A_XmsPwX095_0;
	wire w_dff_A_C4p2jBQJ3_0;
	wire w_dff_A_eFZQk3Eh1_0;
	wire w_dff_A_zM5vnYCu7_0;
	wire w_dff_A_9Nsn4WGU2_0;
	wire w_dff_A_EeliMwh14_0;
	wire w_dff_A_TGvP4lDF0_0;
	wire w_dff_A_ERuSPKMK5_0;
	wire w_dff_A_vYRT9OcE8_0;
	wire w_dff_A_0JP3jwNj8_2;
	wire w_dff_A_9y7nuPwr7_0;
	wire w_dff_A_rwDIbwDH8_0;
	wire w_dff_A_EC2jM1kI2_0;
	wire w_dff_A_sFFvZO1G5_0;
	wire w_dff_A_o69ULqdI8_0;
	wire w_dff_A_vnvzQmvE8_0;
	wire w_dff_A_vPYQKSFe7_0;
	wire w_dff_A_Q3xFXEYr9_0;
	wire w_dff_A_2p1SoVej6_0;
	wire w_dff_A_gICOUGPW3_0;
	wire w_dff_A_wrJOAbeg2_0;
	wire w_dff_A_OZNbhE6V0_0;
	wire w_dff_A_dXbCAxYc2_0;
	wire w_dff_A_DWCE28Yg2_0;
	wire w_dff_A_ZW80NjQM6_0;
	wire w_dff_A_S5US0VGX6_0;
	wire w_dff_A_dD5cbYH40_0;
	wire w_dff_A_8Tbz3cTc1_0;
	wire w_dff_A_gAAIlYDy1_0;
	wire w_dff_A_aVN2lUok7_0;
	wire w_dff_A_EZkZivps6_0;
	wire w_dff_A_Z6qNvanW8_0;
	wire w_dff_A_YosXUhTH6_0;
	wire w_dff_A_SCZnhn4U6_0;
	wire w_dff_A_QCZh84Pu6_0;
	wire w_dff_A_tmlCZHY94_0;
	wire w_dff_A_UIsUUhaR9_0;
	wire w_dff_A_N9aQ43IP4_0;
	wire w_dff_A_wU9Lxyep3_0;
	wire w_dff_A_c0efwtBe5_0;
	wire w_dff_A_8SbIfut79_0;
	wire w_dff_A_tr4GEd7E8_0;
	wire w_dff_A_x9Ksuv9a4_0;
	wire w_dff_A_fKGrflfG7_0;
	wire w_dff_A_2FXSAPhw0_0;
	wire w_dff_A_8fEcePn13_0;
	wire w_dff_A_dZ2Or8Zg3_0;
	wire w_dff_A_PicvuRuG1_0;
	wire w_dff_A_8kdxz9Ch5_0;
	wire w_dff_A_JTlG9CDe6_0;
	wire w_dff_A_nuB0GE4r1_0;
	wire w_dff_A_MR2XgASb7_0;
	wire w_dff_A_tFWlQKnh6_0;
	wire w_dff_A_bhnfYepS4_0;
	wire w_dff_A_S9bBKKld1_0;
	wire w_dff_A_cHdYMAfi8_0;
	wire w_dff_A_r9Nlqm7i4_0;
	wire w_dff_A_XkHpznFV3_0;
	wire w_dff_A_CyXriHxa6_0;
	wire w_dff_A_GmIQqCmU1_0;
	wire w_dff_A_W06CTYbN9_0;
	wire w_dff_A_S5MkaSO17_0;
	wire w_dff_A_l4fMSMGb2_0;
	wire w_dff_A_tDHTbtHD9_2;
	wire w_dff_A_q8aFmGwZ4_0;
	wire w_dff_A_A0jCiuli4_0;
	wire w_dff_A_h6HUAdhD6_0;
	wire w_dff_A_yNxj5BwM7_0;
	wire w_dff_A_p7RJdatl3_0;
	wire w_dff_A_CiDFMdkw8_0;
	wire w_dff_A_ofCcrgmp4_0;
	wire w_dff_A_Xo7ZIekS3_0;
	wire w_dff_A_RpFuB8Qn1_0;
	wire w_dff_A_14TbbzkY5_0;
	wire w_dff_A_uXxcj9tz7_0;
	wire w_dff_A_BHFk1Yzt1_0;
	wire w_dff_A_50bpTB1X7_0;
	wire w_dff_A_dIi3DsUF7_0;
	wire w_dff_A_upeYc7wD8_0;
	wire w_dff_A_5Ld78PMj9_0;
	wire w_dff_A_SSt2Kutn2_0;
	wire w_dff_A_gDbYxs4x9_0;
	wire w_dff_A_uYgVlVl84_0;
	wire w_dff_A_j2ctZomr5_0;
	wire w_dff_A_ZxJillTQ5_0;
	wire w_dff_A_QJVAZTCR0_0;
	wire w_dff_A_tvh4sAEC5_0;
	wire w_dff_A_bKZ7AmGt4_0;
	wire w_dff_A_U9GbU6Fx4_0;
	wire w_dff_A_GbUPDE3q6_0;
	wire w_dff_A_QiHzXXPs8_0;
	wire w_dff_A_noWrcSJX8_0;
	wire w_dff_A_3XzaxxNv0_0;
	wire w_dff_A_3uePTLzI7_0;
	wire w_dff_A_rzlm0Y8B9_0;
	wire w_dff_A_SdU8bPRz6_0;
	wire w_dff_A_9gdr0Xiz7_0;
	wire w_dff_A_R08VmBP44_0;
	wire w_dff_A_Ik9SmEod2_0;
	wire w_dff_A_rUGlc7xG3_0;
	wire w_dff_A_NE0Xxvtv7_0;
	wire w_dff_A_agiBJQfc9_0;
	wire w_dff_A_5OTMzzmz6_0;
	wire w_dff_A_Pj0pm2Lm9_0;
	wire w_dff_A_3VPgA6oT7_0;
	wire w_dff_A_UU2TEuBj0_0;
	wire w_dff_A_P125C3pf9_0;
	wire w_dff_A_XFrQZNcg6_0;
	wire w_dff_A_emcMfYOC1_0;
	wire w_dff_A_eq14Vo006_0;
	wire w_dff_A_nGM6iWhg4_0;
	wire w_dff_A_0Tuq0Iiq2_0;
	wire w_dff_A_FDDth7LC2_0;
	wire w_dff_A_YVygEv5j9_0;
	wire w_dff_A_yY8yxN6c1_2;
	wire w_dff_A_0b1wWLal0_0;
	wire w_dff_A_9v1dS7BS6_0;
	wire w_dff_A_vM9hfPwR7_0;
	wire w_dff_A_vwnSNPbd6_0;
	wire w_dff_A_t7Nr2H954_0;
	wire w_dff_A_PRPqvJq75_0;
	wire w_dff_A_P8lKd5Ei4_0;
	wire w_dff_A_nClFaeR25_0;
	wire w_dff_A_7OdD3DtH2_0;
	wire w_dff_A_i96Tcl8H9_0;
	wire w_dff_A_z53VELXU9_0;
	wire w_dff_A_JG4tHwD50_0;
	wire w_dff_A_TB75Yj5y7_0;
	wire w_dff_A_fCfZubvv1_0;
	wire w_dff_A_1Sdie3if2_0;
	wire w_dff_A_lkQwCQPJ1_0;
	wire w_dff_A_j3Ohi46O8_0;
	wire w_dff_A_UIP0i0cf1_0;
	wire w_dff_A_fmR0BYtz3_0;
	wire w_dff_A_of14nbZc5_0;
	wire w_dff_A_gAnzB6kQ3_0;
	wire w_dff_A_brmmQzJT5_0;
	wire w_dff_A_NkbS25FG6_0;
	wire w_dff_A_rw3kTQKb0_0;
	wire w_dff_A_40WdcH1w2_0;
	wire w_dff_A_7BYduC8C8_0;
	wire w_dff_A_NeIWGPHg2_0;
	wire w_dff_A_u7aqd18z4_0;
	wire w_dff_A_G4ZC9E6f8_0;
	wire w_dff_A_9k9HSoWQ7_0;
	wire w_dff_A_1XGm5JsJ0_0;
	wire w_dff_A_EJ1X0jFs0_0;
	wire w_dff_A_YJ7iCCNq3_0;
	wire w_dff_A_gLNRFF4J1_0;
	wire w_dff_A_mPZgSX809_0;
	wire w_dff_A_NnglkXpB4_0;
	wire w_dff_A_B8fArUQK7_0;
	wire w_dff_A_CVW4O55p7_0;
	wire w_dff_A_RCwCBnkA9_0;
	wire w_dff_A_E33sluXJ1_0;
	wire w_dff_A_FnVM3lPo6_0;
	wire w_dff_A_1J2KOAl32_0;
	wire w_dff_A_R6MIg0XX3_0;
	wire w_dff_A_aL2jgIDE2_0;
	wire w_dff_A_i1Q5XMKk5_0;
	wire w_dff_A_Q36wvf1V6_0;
	wire w_dff_A_BsgY16DA7_0;
	wire w_dff_A_fbgsIzQB8_2;
	wire w_dff_A_qNCNU8F57_0;
	wire w_dff_A_rfKRqyHU1_0;
	wire w_dff_A_ovHxfjTD4_0;
	wire w_dff_A_OX1r2rZU1_0;
	wire w_dff_A_L5drJ2ae2_0;
	wire w_dff_A_bARdbM5a4_0;
	wire w_dff_A_AuZTwuwb0_0;
	wire w_dff_A_VA6UYDbr0_0;
	wire w_dff_A_nb2VvcMG1_0;
	wire w_dff_A_MePFNjtP3_0;
	wire w_dff_A_ZiV2sNfm9_0;
	wire w_dff_A_q45HJ2GB2_0;
	wire w_dff_A_CZP3qcSt4_0;
	wire w_dff_A_DS6MY5VM5_0;
	wire w_dff_A_DdPtjZeI8_0;
	wire w_dff_A_pFyblxKc4_0;
	wire w_dff_A_f9CFv9jU8_0;
	wire w_dff_A_asFNwthJ7_0;
	wire w_dff_A_W6Apw8iQ4_0;
	wire w_dff_A_oFLy3QE49_0;
	wire w_dff_A_9HvlsRXd7_0;
	wire w_dff_A_fYfG2ma35_0;
	wire w_dff_A_SelniTRZ8_0;
	wire w_dff_A_rV80BmMk3_0;
	wire w_dff_A_qLroIxiw2_0;
	wire w_dff_A_a85xfeTt2_0;
	wire w_dff_A_jGDSUmUd3_0;
	wire w_dff_A_eOOedJWz2_0;
	wire w_dff_A_uDRtnHPv0_0;
	wire w_dff_A_oxMhZN4T2_0;
	wire w_dff_A_ESxJ4YV42_0;
	wire w_dff_A_paPIw30Y4_0;
	wire w_dff_A_qLEpEyQN5_0;
	wire w_dff_A_qVyleftZ2_0;
	wire w_dff_A_4foWbfZS4_0;
	wire w_dff_A_xKh5cuOz4_0;
	wire w_dff_A_RmSzaXQB6_0;
	wire w_dff_A_0MObwkrQ2_0;
	wire w_dff_A_fgKlhONG3_0;
	wire w_dff_A_7V7YIKOI2_0;
	wire w_dff_A_bswxh8ik4_0;
	wire w_dff_A_6frSAAOX8_0;
	wire w_dff_A_T8XkDwd88_0;
	wire w_dff_A_8pOYho5g0_0;
	wire w_dff_A_DQUJXFRm8_2;
	wire w_dff_A_JFTtzcUb4_0;
	wire w_dff_A_HFjeRtC20_0;
	wire w_dff_A_wD8F8hqE4_0;
	wire w_dff_A_wVjVJ9ib8_0;
	wire w_dff_A_7GWRsU4V5_0;
	wire w_dff_A_beufR2cX8_0;
	wire w_dff_A_9gbRHc2e8_0;
	wire w_dff_A_M5tnwTok7_0;
	wire w_dff_A_dysjJHkp7_0;
	wire w_dff_A_5lTRNEKv6_0;
	wire w_dff_A_fkkSoLPu0_0;
	wire w_dff_A_VTBh2ZbQ4_0;
	wire w_dff_A_61uc9PD59_0;
	wire w_dff_A_bWdrDN9S0_0;
	wire w_dff_A_F3zsr08B1_0;
	wire w_dff_A_UjKGELjN8_0;
	wire w_dff_A_M23keRjl5_0;
	wire w_dff_A_H2Ro9ix14_0;
	wire w_dff_A_WAHmXhtO6_0;
	wire w_dff_A_QKKsJc3r3_0;
	wire w_dff_A_hF66G8km0_0;
	wire w_dff_A_Wlx5e4gI1_0;
	wire w_dff_A_L8ZrONbv7_0;
	wire w_dff_A_cBCe8gcX8_0;
	wire w_dff_A_dH9tmkyX1_0;
	wire w_dff_A_imBoMl9G9_0;
	wire w_dff_A_W1mS41bH9_0;
	wire w_dff_A_ACIeM6bW5_0;
	wire w_dff_A_644sRsx45_0;
	wire w_dff_A_LJUwWryI9_0;
	wire w_dff_A_bX0adZO72_0;
	wire w_dff_A_TtQPRtxi8_0;
	wire w_dff_A_ZvkeB0Gf4_0;
	wire w_dff_A_ZYE6agFO2_0;
	wire w_dff_A_JTmjFYKV3_0;
	wire w_dff_A_HzLv7mXe8_0;
	wire w_dff_A_4jUeqfUz6_0;
	wire w_dff_A_YM0Fr3Pz8_0;
	wire w_dff_A_IRmNQcGl4_0;
	wire w_dff_A_hpYCYBbp1_0;
	wire w_dff_A_xdIs2me35_0;
	wire w_dff_A_8ScMJPuv8_2;
	wire w_dff_A_1sXjWFsi8_0;
	wire w_dff_A_vTjFl9Rn3_0;
	wire w_dff_A_NMYpmCh04_0;
	wire w_dff_A_XyPynqNI2_0;
	wire w_dff_A_CmQ5euX20_0;
	wire w_dff_A_kWoSzfOi0_0;
	wire w_dff_A_7c1wBPh17_0;
	wire w_dff_A_pbz9b6dE0_0;
	wire w_dff_A_g1d3kRWY8_0;
	wire w_dff_A_cU7By3wf1_0;
	wire w_dff_A_GsWeOOmM5_0;
	wire w_dff_A_5ApPesxj5_0;
	wire w_dff_A_kDEVRP9n3_0;
	wire w_dff_A_g3OrA6nu4_0;
	wire w_dff_A_icC5L8Iv9_0;
	wire w_dff_A_w2HZqHfQ1_0;
	wire w_dff_A_x3qiTCHS1_0;
	wire w_dff_A_7ZqXSU3f2_0;
	wire w_dff_A_lTpGPtBB9_0;
	wire w_dff_A_eMUjKrFr8_0;
	wire w_dff_A_EEYxIu5s7_0;
	wire w_dff_A_4ZKLbhg75_0;
	wire w_dff_A_CZdMZ5Cv1_0;
	wire w_dff_A_UunUEequ1_0;
	wire w_dff_A_HyF0T5Xn1_0;
	wire w_dff_A_soyjrbM79_0;
	wire w_dff_A_t6fhRwBl7_0;
	wire w_dff_A_ZCBCQ7Wy8_0;
	wire w_dff_A_4bwfYfC41_0;
	wire w_dff_A_wPQlhMFN9_0;
	wire w_dff_A_CvB16kXw1_0;
	wire w_dff_A_EFMkvWW48_0;
	wire w_dff_A_B5lzMnH01_0;
	wire w_dff_A_foGIT7xW2_0;
	wire w_dff_A_7aqBwVGZ2_0;
	wire w_dff_A_vP8nQb8o3_0;
	wire w_dff_A_ogiUPDms9_0;
	wire w_dff_A_mVvJiUQc0_0;
	wire w_dff_A_rUJAEsv64_2;
	wire w_dff_A_JYqPvBDT0_0;
	wire w_dff_A_VYAN729f8_0;
	wire w_dff_A_qtCHvmpF5_0;
	wire w_dff_A_SrxwfNOz6_0;
	wire w_dff_A_BXNLoJpd5_0;
	wire w_dff_A_QhYkGcty4_0;
	wire w_dff_A_t12lW47r2_0;
	wire w_dff_A_hSiAqwwP3_0;
	wire w_dff_A_GwI3OZQm6_0;
	wire w_dff_A_r2Trua028_0;
	wire w_dff_A_Fi9ds2FE8_0;
	wire w_dff_A_clqbhO766_0;
	wire w_dff_A_eCqlIYJn5_0;
	wire w_dff_A_WJqIf4YB2_0;
	wire w_dff_A_fPTxrkDm3_0;
	wire w_dff_A_a2vJftVL1_0;
	wire w_dff_A_x2fm1VxS0_0;
	wire w_dff_A_OEf8OgmG6_0;
	wire w_dff_A_QCqVLBS73_0;
	wire w_dff_A_nZiHrkMA3_0;
	wire w_dff_A_vE1RCgDa7_0;
	wire w_dff_A_G56Oklg13_0;
	wire w_dff_A_CSodMM0w7_0;
	wire w_dff_A_zcaXJL5A1_0;
	wire w_dff_A_YWyc4epU3_0;
	wire w_dff_A_Pjvj8V4g0_0;
	wire w_dff_A_Z0MHmglx6_0;
	wire w_dff_A_ECyjikka2_0;
	wire w_dff_A_yYyqOtGw9_0;
	wire w_dff_A_tH8tLAvU3_0;
	wire w_dff_A_SSE78vj12_0;
	wire w_dff_A_TorGxQLr8_0;
	wire w_dff_A_uww9Xvi05_0;
	wire w_dff_A_RyQFf0FN1_0;
	wire w_dff_A_YBcaU1TX9_0;
	wire w_dff_A_84xyMY4Y3_2;
	wire w_dff_A_XTJhTSGg9_0;
	wire w_dff_A_sXhMawUE8_0;
	wire w_dff_A_sN2E6JPZ3_0;
	wire w_dff_A_b5ZxHcPc0_0;
	wire w_dff_A_FZyfrE312_0;
	wire w_dff_A_QDPN4ozZ1_0;
	wire w_dff_A_OY5geCES6_0;
	wire w_dff_A_ZSWMtmIt5_0;
	wire w_dff_A_MNDivmGy2_0;
	wire w_dff_A_lz1MYfga9_0;
	wire w_dff_A_s4EZuP6e6_0;
	wire w_dff_A_afiW7GTk6_0;
	wire w_dff_A_wQ7vsfjB9_0;
	wire w_dff_A_K8JOOwg21_0;
	wire w_dff_A_kr6VHYWe5_0;
	wire w_dff_A_dEIxKwy43_0;
	wire w_dff_A_nerKESo28_0;
	wire w_dff_A_wPxiTZLp4_0;
	wire w_dff_A_YLDbwvF19_0;
	wire w_dff_A_OdnUEPO55_0;
	wire w_dff_A_P9sAmqPJ3_0;
	wire w_dff_A_dFpb3NUm9_0;
	wire w_dff_A_JLc2T2nW7_0;
	wire w_dff_A_fsLSZjJc9_0;
	wire w_dff_A_PO2quGnb2_0;
	wire w_dff_A_d323YXze7_0;
	wire w_dff_A_gbjPXZff0_0;
	wire w_dff_A_gVATgN0m7_0;
	wire w_dff_A_L4cqZF7I6_0;
	wire w_dff_A_bpGAAgeE1_0;
	wire w_dff_A_xB0BdyQL4_0;
	wire w_dff_A_hRShA0ed5_0;
	wire w_dff_A_1raJBPiI7_2;
	wire w_dff_A_b0A700nA8_0;
	wire w_dff_A_EtbUJt987_0;
	wire w_dff_A_0swVoc0V3_0;
	wire w_dff_A_CHqs3Bxe6_0;
	wire w_dff_A_FyJscuXk5_0;
	wire w_dff_A_DgTOnl1P9_0;
	wire w_dff_A_Ax5KdSXQ6_0;
	wire w_dff_A_mQf30PIE5_0;
	wire w_dff_A_tbPuAVsh2_0;
	wire w_dff_A_LP01NtDK9_0;
	wire w_dff_A_21FkTXyp3_0;
	wire w_dff_A_qIWPi15m5_0;
	wire w_dff_A_lQbnPwvX5_0;
	wire w_dff_A_NtDgGHN10_0;
	wire w_dff_A_uYrhRVcn8_0;
	wire w_dff_A_iF8emuVV5_0;
	wire w_dff_A_S7Rt2u0W1_0;
	wire w_dff_A_T447om4z0_0;
	wire w_dff_A_VVqMdkWK7_0;
	wire w_dff_A_AhsZsNcg0_0;
	wire w_dff_A_1B0OHMJC9_0;
	wire w_dff_A_XWSbTKbY2_0;
	wire w_dff_A_1lvipsKF1_0;
	wire w_dff_A_2lzSU0s65_0;
	wire w_dff_A_KPlMCcWP0_0;
	wire w_dff_A_YKhpwTBF5_0;
	wire w_dff_A_1lOkirMM1_0;
	wire w_dff_A_NgKhnMyS0_0;
	wire w_dff_A_4ZOHlOK03_0;
	wire w_dff_A_y2Cx0Ugv4_2;
	wire w_dff_A_IM9zw3ip2_0;
	wire w_dff_A_GuG5kwK45_0;
	wire w_dff_A_HQDaexNy9_0;
	wire w_dff_A_XFlsTBiF8_0;
	wire w_dff_A_tLsJc26L9_0;
	wire w_dff_A_YPpQaonI8_0;
	wire w_dff_A_JD7hAYLi4_0;
	wire w_dff_A_iyCJsjJN7_0;
	wire w_dff_A_rR3kr6zM4_0;
	wire w_dff_A_sG66h2zR4_0;
	wire w_dff_A_7VOJ2J6Z1_0;
	wire w_dff_A_W3vTYauk0_0;
	wire w_dff_A_NM2eYEB24_0;
	wire w_dff_A_8YuQDSsh2_0;
	wire w_dff_A_T6skV5jX5_0;
	wire w_dff_A_Vt2bouFW6_0;
	wire w_dff_A_H0Wn6B0I3_0;
	wire w_dff_A_1PG892WP2_0;
	wire w_dff_A_agF66L0e9_0;
	wire w_dff_A_JACyKZqv6_0;
	wire w_dff_A_YgNyNfM41_0;
	wire w_dff_A_hrW6acbg0_0;
	wire w_dff_A_WcMAmwaU7_0;
	wire w_dff_A_6SV7dqQK4_0;
	wire w_dff_A_8apvyxvv6_0;
	wire w_dff_A_gd8vqqrV6_0;
	wire w_dff_A_SUNrvR1n8_0;
	wire w_dff_A_SvwK5EUw5_2;
	wire w_dff_A_bjd83Vxj5_0;
	wire w_dff_A_x9BftWh56_0;
	wire w_dff_A_bwo486E10_0;
	wire w_dff_A_xkMMLt5c7_0;
	wire w_dff_A_ruSffF2E4_0;
	wire w_dff_A_u83didJi9_0;
	wire w_dff_A_SX9Eezw61_0;
	wire w_dff_A_VywakCAI0_0;
	wire w_dff_A_HHhOAcAy8_0;
	wire w_dff_A_RGovoSLq4_0;
	wire w_dff_A_c6mK9v437_0;
	wire w_dff_A_Mdxt7XPY9_0;
	wire w_dff_A_5Jr7QOea1_0;
	wire w_dff_A_hoZveZIZ4_0;
	wire w_dff_A_HVlW4p3D1_0;
	wire w_dff_A_nKuLprAn3_0;
	wire w_dff_A_ofZYTtmx6_0;
	wire w_dff_A_DiCHfkEQ6_0;
	wire w_dff_A_x0CBrwWu5_0;
	wire w_dff_A_u5hkAvVI5_0;
	wire w_dff_A_CiM46Hfy3_0;
	wire w_dff_A_H4TnNXJI2_0;
	wire w_dff_A_KLkNfKOu4_0;
	wire w_dff_A_4oFE5pXi0_0;
	wire w_dff_A_s39hK2rb3_0;
	wire w_dff_A_EELcdX9T0_2;
	wire w_dff_A_gufvd4Sv1_0;
	wire w_dff_A_EHNCK4Ft7_0;
	wire w_dff_A_SZNA8S4J5_0;
	wire w_dff_A_UP180uH48_0;
	wire w_dff_A_7tOsaqMl7_0;
	wire w_dff_A_EqdzPePq4_0;
	wire w_dff_A_BFf5iGPR9_0;
	wire w_dff_A_hSUBVtHL8_0;
	wire w_dff_A_gfs4PPv88_0;
	wire w_dff_A_lEIKIGiG4_0;
	wire w_dff_A_NJddlC4g2_0;
	wire w_dff_A_omlpZSum4_0;
	wire w_dff_A_qHPpO4G22_0;
	wire w_dff_A_fYwezJSA2_0;
	wire w_dff_A_Xq5Ii9hC4_0;
	wire w_dff_A_RkjQx0pg0_0;
	wire w_dff_A_posI18bm7_0;
	wire w_dff_A_TsSkDL2w4_0;
	wire w_dff_A_5DnQ9DTu6_0;
	wire w_dff_A_jF8lu5fj3_0;
	wire w_dff_A_Eb4STl0r7_0;
	wire w_dff_A_hW0BFO5Z8_0;
	wire w_dff_A_L1grFQ8m3_0;
	wire w_dff_A_nA71Rspl2_0;
	wire w_dff_A_RRpqyqj39_2;
	wire w_dff_A_W05T6Vtq2_0;
	wire w_dff_A_iB45JsjX3_0;
	wire w_dff_A_WJcSqkwi3_0;
	wire w_dff_A_23r1uK1y2_0;
	wire w_dff_A_r2igO0z46_0;
	wire w_dff_A_aJnIeCz43_0;
	wire w_dff_A_oK8tOAyr2_0;
	wire w_dff_A_OeqywrbW2_0;
	wire w_dff_A_EROGwThe8_0;
	wire w_dff_A_YvPWHAVr6_0;
	wire w_dff_A_AQ2TWwBn4_0;
	wire w_dff_A_SjyFdkBI1_0;
	wire w_dff_A_fYnjaFlm9_0;
	wire w_dff_A_R8zPP88j0_0;
	wire w_dff_A_ZQQzkbON9_0;
	wire w_dff_A_R9C4OhDh2_0;
	wire w_dff_A_ZruFFfjo8_0;
	wire w_dff_A_34NIgfUP0_0;
	wire w_dff_A_hEit6H518_0;
	wire w_dff_A_iNBAwf6Y9_0;
	wire w_dff_A_eS1NZCvx0_0;
	wire w_dff_A_D9cfx2J05_0;
	wire w_dff_A_qnZGkGXX4_2;
	wire w_dff_A_MrUqgbmz4_0;
	wire w_dff_A_YzHzUYsy2_0;
	wire w_dff_A_BQpyPue48_0;
	wire w_dff_A_ToE0Uzaa1_0;
	wire w_dff_A_GTcSazS79_0;
	wire w_dff_A_e1O9BePz0_0;
	wire w_dff_A_L34fsglg0_0;
	wire w_dff_A_5SBShVGD5_0;
	wire w_dff_A_Cac4DcrY6_0;
	wire w_dff_A_dbFnQviG9_0;
	wire w_dff_A_dxRFwI2D7_0;
	wire w_dff_A_IKDAjMqW5_0;
	wire w_dff_A_3b0H7rvu6_0;
	wire w_dff_A_SdRXAC8i4_0;
	wire w_dff_A_CmQM7OPJ6_0;
	wire w_dff_A_Xl1H6DCG8_0;
	wire w_dff_A_pXI6Kagq6_0;
	wire w_dff_A_ijoNJwum0_0;
	wire w_dff_A_WVQpKK2N9_0;
	wire w_dff_A_Xo1pRnTM3_0;
	wire w_dff_A_WXOrmoWW8_2;
	wire w_dff_A_YD9nUo5Y2_0;
	wire w_dff_A_6222Yix48_0;
	wire w_dff_A_VLK1D3XO4_0;
	wire w_dff_A_qqwnvcOY4_0;
	wire w_dff_A_HhTak8JX4_0;
	wire w_dff_A_XeoNVGQX0_0;
	wire w_dff_A_L9N8ivgX5_0;
	wire w_dff_A_UwsvkvX28_0;
	wire w_dff_A_f94bDBZ40_0;
	wire w_dff_A_ugLDeNNj6_0;
	wire w_dff_A_9EmocGAs7_0;
	wire w_dff_A_XOfhhKrZ3_0;
	wire w_dff_A_EA5B83wV8_0;
	wire w_dff_A_292ORCPw0_0;
	wire w_dff_A_scfpyQbO1_0;
	wire w_dff_A_7aiN5HCM8_0;
	wire w_dff_A_eLb1kdS36_0;
	wire w_dff_A_0C9Oi0wz7_0;
	wire w_dff_A_zBf6HHia3_2;
	wire w_dff_A_Cu2Gj7gW1_0;
	wire w_dff_A_mbzG29En6_0;
	wire w_dff_A_1lPBvm1B0_0;
	wire w_dff_A_0oyWFeur6_0;
	wire w_dff_A_QbFecoML7_0;
	wire w_dff_A_YuUqoDk83_0;
	wire w_dff_A_6B1ZG7hd4_0;
	wire w_dff_A_RGKk3GKA7_0;
	wire w_dff_A_Y2WspOBJ8_0;
	wire w_dff_A_2FOAFc9a3_0;
	wire w_dff_A_gbxlx1kB9_0;
	wire w_dff_A_ygU1NomP4_0;
	wire w_dff_A_D51HS72s5_0;
	wire w_dff_A_3SlxXx1b3_0;
	wire w_dff_A_PNUJ3g586_0;
	wire w_dff_A_vkEGzOEX2_0;
	wire w_dff_A_VdYZ4TDy2_2;
	wire w_dff_A_QqM89tHL5_0;
	wire w_dff_A_bQEtXRSJ5_0;
	wire w_dff_A_Xqh191pB3_0;
	wire w_dff_A_MNYBlyGd7_0;
	wire w_dff_A_QEuc27FI9_0;
	wire w_dff_A_3Q6eYBmT0_0;
	wire w_dff_A_HwoLkaH27_0;
	wire w_dff_A_JWFBjUrt6_0;
	wire w_dff_A_TnUyeyoj9_0;
	wire w_dff_A_mBhYgjfA1_0;
	wire w_dff_A_26BAZ0Yn0_0;
	wire w_dff_A_jbabzuMu4_0;
	wire w_dff_A_vc4KjUy91_0;
	wire w_dff_A_rdeBYawA9_0;
	wire w_dff_A_AlZA3pCn3_2;
	wire w_dff_A_IjYaULZR8_0;
	wire w_dff_A_TbbjLwsR9_0;
	wire w_dff_A_CC1v8XDI2_0;
	wire w_dff_A_WuSmD3gK6_0;
	wire w_dff_A_HXNWaxWZ9_0;
	wire w_dff_A_f5cnWkfv1_0;
	wire w_dff_A_kuvEhMcr4_0;
	wire w_dff_A_hnGk9Q8V0_0;
	wire w_dff_A_UeqvxuhD3_0;
	wire w_dff_A_h6LR23uM8_0;
	wire w_dff_A_4yqZ4Pre6_0;
	wire w_dff_A_VzHzPI6Y7_0;
	wire w_dff_A_x9YO84OD2_2;
	wire w_dff_A_q9IerLkm3_0;
	wire w_dff_A_EVgzEf1Q6_0;
	wire w_dff_A_sl9KLPig2_0;
	wire w_dff_A_yxgyofFe1_0;
	wire w_dff_A_5rflpenG1_0;
	wire w_dff_A_WzzfEBtd4_0;
	wire w_dff_A_iKVcCPPa2_0;
	wire w_dff_A_MREacc6p1_0;
	wire w_dff_A_AcLskXXc1_0;
	wire w_dff_A_1g6mJbci7_0;
	wire w_dff_A_YgTyAIea9_2;
	wire w_dff_A_FdapSK7r3_0;
	wire w_dff_A_OQPZteuG2_0;
	wire w_dff_A_iKWHgDRZ0_0;
	wire w_dff_A_TtcaAFp44_0;
	wire w_dff_A_pWpLbvuA9_0;
	wire w_dff_A_N5GSayY97_0;
	wire w_dff_A_LIox8mrh5_0;
	wire w_dff_A_CjxTm4vc0_0;
	wire w_dff_A_1aNiPV9I1_2;
	wire w_dff_A_yw6ZvmmJ6_0;
	wire w_dff_A_RUHFp4pu4_0;
	wire w_dff_A_QqBqEDwE9_0;
	wire w_dff_A_V0roDClD2_0;
	wire w_dff_A_4dMcpDyQ8_0;
	wire w_dff_A_FBcr8KZO8_0;
	wire w_dff_A_xYpvdcGX7_2;
	wire w_dff_A_boGHSrLK5_0;
	wire w_dff_A_setKgQZu2_0;
	wire w_dff_A_pB90dIRx5_0;
	wire w_dff_A_7SeyXxwC1_0;
	wire w_dff_A_oBPVQzMN0_2;
	wire w_dff_A_XdEtSXX40_0;
	wire w_dff_A_JZUSrm1M4_0;
	wire w_dff_A_i6yb8BNW4_2;
	jand g0000(.dina(w_G273gat_7[1]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G290gat_7[2]),.dinb(w_G18gat_7[1]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_n65_0[1]),.dinb(w_G545gat_0),.dout(n66),.clk(gclk));
	jnot g0003(.din(w_n66_0[1]),.dout(n67),.clk(gclk));
	jnot g0004(.din(w_G18gat_7[0]),.dout(n68),.clk(gclk));
	jnot g0005(.din(w_G273gat_7[0]),.dout(n69),.clk(gclk));
	jor g0006(.dina(w_n69_0[1]),.dinb(n68),.dout(n70),.clk(gclk));
	jnot g0007(.din(w_n70_0[1]),.dout(n71),.clk(gclk));
	jand g0008(.dina(w_G290gat_7[1]),.dinb(w_G1gat_7[0]),.dout(n72),.clk(gclk));
	jor g0009(.dina(w_dff_B_xtZmTHUA1_0),.dinb(n71),.dout(n73),.clk(gclk));
	jand g0010(.dina(n73),.dinb(w_n67_0[1]),.dout(w_dff_A_ERwqQcch6_2),.clk(gclk));
	jand g0011(.dina(w_G307gat_7[1]),.dinb(w_G1gat_6[2]),.dout(n75),.clk(gclk));
	jnot g0012(.din(w_n75_0[1]),.dout(n76),.clk(gclk));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G290gat_7[0]),.dout(n78),.clk(gclk));
	jor g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79),.clk(gclk));
	jor g0016(.dina(n79),.dinb(w_n70_0[0]),.dout(n80),.clk(gclk));
	jand g0017(.dina(w_G273gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jor g0018(.dina(n81),.dinb(w_n65_0[0]),.dout(n82),.clk(gclk));
	jand g0019(.dina(w_dff_B_4AVndoHp8_0),.dinb(w_n80_0[2]),.dout(n83),.clk(gclk));
	jxor g0020(.dina(w_n83_0[1]),.dinb(w_n67_0[0]),.dout(n84),.clk(gclk));
	jxor g0021(.dina(w_n84_0[1]),.dinb(w_dff_B_c1j5Gyez3_1),.dout(w_dff_A_JVhOTcac7_2),.clk(gclk));
	jand g0022(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n86),.clk(gclk));
	jnot g0023(.din(w_n86_0[1]),.dout(n87),.clk(gclk));
	jor g0024(.dina(w_n83_0[0]),.dinb(w_n66_0[0]),.dout(n88),.clk(gclk));
	jor g0025(.dina(w_n84_0[0]),.dinb(w_n75_0[0]),.dout(n89),.clk(gclk));
	jand g0026(.dina(n89),.dinb(w_dff_B_UGGTIAOT5_1),.dout(n90),.clk(gclk));
	jand g0027(.dina(w_G307gat_7[0]),.dinb(w_G18gat_6[2]),.dout(n91),.clk(gclk));
	jnot g0028(.din(w_n91_0[1]),.dout(n92),.clk(gclk));
	jnot g0029(.din(w_n80_0[1]),.dout(n93),.clk(gclk));
	jor g0030(.dina(w_n69_0[0]),.dinb(w_n77_0[0]),.dout(n94),.clk(gclk));
	jnot g0031(.din(w_G52gat_7[2]),.dout(n95),.clk(gclk));
	jor g0032(.dina(w_n78_0[0]),.dinb(n95),.dout(n96),.clk(gclk));
	jor g0033(.dina(n96),.dinb(n94),.dout(n97),.clk(gclk));
	jand g0034(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G273gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jor g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100),.clk(gclk));
	jand g0037(.dina(w_dff_B_lUl1Ec815_0),.dinb(w_n97_0[1]),.dout(n101),.clk(gclk));
	jxor g0038(.dina(w_n101_0[2]),.dinb(w_n93_0[1]),.dout(n102),.clk(gclk));
	jxor g0039(.dina(n102),.dinb(w_dff_B_VxStCGKZ2_1),.dout(n103),.clk(gclk));
	jxor g0040(.dina(w_n103_0[1]),.dinb(w_n90_0[1]),.dout(n104),.clk(gclk));
	jxor g0041(.dina(w_n104_0[1]),.dinb(w_dff_B_TnLU4N4R5_1),.dout(w_dff_A_1yMaWZic3_2),.clk(gclk));
	jand g0042(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n106),.clk(gclk));
	jnot g0043(.din(w_n106_0[1]),.dout(n107),.clk(gclk));
	jnot g0044(.din(w_n103_0[0]),.dout(n108),.clk(gclk));
	jor g0045(.dina(n108),.dinb(w_n90_0[0]),.dout(n109),.clk(gclk));
	jor g0046(.dina(w_n104_0[0]),.dinb(w_n86_0[0]),.dout(n110),.clk(gclk));
	jand g0047(.dina(n110),.dinb(w_dff_B_MwfEWbpP9_1),.dout(n111),.clk(gclk));
	jand g0048(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n112),.clk(gclk));
	jnot g0049(.din(w_n112_0[1]),.dout(n113),.clk(gclk));
	jor g0050(.dina(w_n101_0[1]),.dinb(w_n93_0[0]),.dout(n114),.clk(gclk));
	jxor g0051(.dina(w_n101_0[0]),.dinb(w_n80_0[0]),.dout(n115),.clk(gclk));
	jor g0052(.dina(n115),.dinb(w_n91_0[0]),.dout(n116),.clk(gclk));
	jand g0053(.dina(n116),.dinb(w_dff_B_665wR8I06_1),.dout(n117),.clk(gclk));
	jand g0054(.dina(w_G307gat_6[2]),.dinb(w_G35gat_6[2]),.dout(n118),.clk(gclk));
	jnot g0055(.din(n118),.dout(n119),.clk(gclk));
	jnot g0056(.din(w_n97_0[0]),.dout(n120),.clk(gclk));
	jand g0057(.dina(w_G290gat_6[1]),.dinb(w_G69gat_7[1]),.dout(n121),.clk(gclk));
	jand g0058(.dina(w_n121_0[1]),.dinb(w_n99_0[0]),.dout(n122),.clk(gclk));
	jnot g0059(.din(w_n122_0[1]),.dout(n123),.clk(gclk));
	jand g0060(.dina(w_G290gat_6[0]),.dinb(w_G52gat_7[0]),.dout(n124),.clk(gclk));
	jand g0061(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n125),.clk(gclk));
	jor g0062(.dina(w_n125_0[1]),.dinb(n124),.dout(n126),.clk(gclk));
	jand g0063(.dina(w_dff_B_Vp1e94050_0),.dinb(w_n123_0[1]),.dout(n127),.clk(gclk));
	jxor g0064(.dina(w_n127_0[1]),.dinb(w_n120_0[1]),.dout(n128),.clk(gclk));
	jxor g0065(.dina(w_n128_0[1]),.dinb(w_n119_0[1]),.dout(n129),.clk(gclk));
	jnot g0066(.din(w_n129_0[1]),.dout(n130),.clk(gclk));
	jxor g0067(.dina(w_n130_0[1]),.dinb(w_n117_0[2]),.dout(n131),.clk(gclk));
	jxor g0068(.dina(n131),.dinb(w_dff_B_gzcghbfG9_1),.dout(n132),.clk(gclk));
	jxor g0069(.dina(w_n132_0[1]),.dinb(w_n111_0[1]),.dout(n133),.clk(gclk));
	jxor g0070(.dina(w_n133_0[1]),.dinb(w_dff_B_2bca4tz20_1),.dout(w_dff_A_THDtcXMv5_2),.clk(gclk));
	jand g0071(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n135),.clk(gclk));
	jnot g0072(.din(w_n135_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(w_n132_0[0]),.dout(n137),.clk(gclk));
	jor g0074(.dina(n137),.dinb(w_n111_0[0]),.dout(n138),.clk(gclk));
	jor g0075(.dina(w_n133_0[0]),.dinb(w_n106_0[0]),.dout(n139),.clk(gclk));
	jand g0076(.dina(n139),.dinb(w_dff_B_ZBGSYhqQ2_1),.dout(n140),.clk(gclk));
	jand g0077(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n141),.clk(gclk));
	jnot g0078(.din(w_n141_0[1]),.dout(n142),.clk(gclk));
	jor g0079(.dina(w_n130_0[0]),.dinb(w_n117_0[1]),.dout(n143),.clk(gclk));
	jxor g0080(.dina(w_n129_0[0]),.dinb(w_n117_0[0]),.dout(n144),.clk(gclk));
	jor g0081(.dina(n144),.dinb(w_n112_0[0]),.dout(n145),.clk(gclk));
	jand g0082(.dina(n145),.dinb(w_dff_B_DPmtQp9y6_1),.dout(n146),.clk(gclk));
	jand g0083(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n147),.clk(gclk));
	jnot g0084(.din(n147),.dout(n148),.clk(gclk));
	jor g0085(.dina(w_n127_0[0]),.dinb(w_n120_0[0]),.dout(n149),.clk(gclk));
	jnot g0086(.din(n149),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_n128_0[0]),.dinb(w_n119_0[0]),.dout(n151),.clk(gclk));
	jor g0088(.dina(n151),.dinb(n150),.dout(n152),.clk(gclk));
	jand g0089(.dina(w_G307gat_6[1]),.dinb(w_G52gat_6[2]),.dout(n153),.clk(gclk));
	jnot g0090(.din(n153),.dout(n154),.clk(gclk));
	jand g0091(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n155),.clk(gclk));
	jand g0092(.dina(w_n155_0[1]),.dinb(w_n125_0[0]),.dout(n156),.clk(gclk));
	jnot g0093(.din(w_n156_0[1]),.dout(n157),.clk(gclk));
	jand g0094(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n158),.clk(gclk));
	jor g0095(.dina(w_n158_0[1]),.dinb(w_n121_0[0]),.dout(n159),.clk(gclk));
	jand g0096(.dina(w_dff_B_r3s5Qos04_0),.dinb(w_n157_0[1]),.dout(n160),.clk(gclk));
	jxor g0097(.dina(w_n160_0[1]),.dinb(w_n122_0[0]),.dout(n161),.clk(gclk));
	jxor g0098(.dina(w_n161_0[1]),.dinb(w_n154_0[1]),.dout(n162),.clk(gclk));
	jxor g0099(.dina(w_n162_0[1]),.dinb(w_n152_0[1]),.dout(n163),.clk(gclk));
	jxor g0100(.dina(w_n163_0[1]),.dinb(w_n148_0[1]),.dout(n164),.clk(gclk));
	jnot g0101(.din(w_n164_0[1]),.dout(n165),.clk(gclk));
	jxor g0102(.dina(w_n165_0[1]),.dinb(w_n146_0[2]),.dout(n166),.clk(gclk));
	jxor g0103(.dina(n166),.dinb(w_dff_B_41TCNUGG3_1),.dout(n167),.clk(gclk));
	jxor g0104(.dina(w_n167_0[1]),.dinb(w_n140_0[1]),.dout(n168),.clk(gclk));
	jxor g0105(.dina(w_n168_0[1]),.dinb(w_dff_B_M3AxJSlC9_1),.dout(w_dff_A_w3mHM9Py5_2),.clk(gclk));
	jand g0106(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n170),.clk(gclk));
	jnot g0107(.din(w_n170_0[1]),.dout(n171),.clk(gclk));
	jnot g0108(.din(w_n167_0[0]),.dout(n172),.clk(gclk));
	jor g0109(.dina(n172),.dinb(w_n140_0[0]),.dout(n173),.clk(gclk));
	jor g0110(.dina(w_n168_0[0]),.dinb(w_n135_0[0]),.dout(n174),.clk(gclk));
	jand g0111(.dina(n174),.dinb(w_dff_B_e5SXL19y3_1),.dout(n175),.clk(gclk));
	jand g0112(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n176),.clk(gclk));
	jnot g0113(.din(w_n176_0[1]),.dout(n177),.clk(gclk));
	jor g0114(.dina(w_n165_0[0]),.dinb(w_n146_0[1]),.dout(n178),.clk(gclk));
	jxor g0115(.dina(w_n164_0[0]),.dinb(w_n146_0[0]),.dout(n179),.clk(gclk));
	jor g0116(.dina(n179),.dinb(w_n141_0[0]),.dout(n180),.clk(gclk));
	jand g0117(.dina(n180),.dinb(w_dff_B_aBtWMcoy6_1),.dout(n181),.clk(gclk));
	jand g0118(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n182),.clk(gclk));
	jnot g0119(.din(n182),.dout(n183),.clk(gclk));
	jand g0120(.dina(w_n162_0[0]),.dinb(w_n152_0[0]),.dout(n184),.clk(gclk));
	jand g0121(.dina(w_n163_0[0]),.dinb(w_n148_0[0]),.dout(n185),.clk(gclk));
	jor g0122(.dina(n185),.dinb(w_dff_B_Ahgr0w2R0_1),.dout(n186),.clk(gclk));
	jand g0123(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n187),.clk(gclk));
	jnot g0124(.din(n187),.dout(n188),.clk(gclk));
	jnot g0125(.din(w_n160_0[0]),.dout(n189),.clk(gclk));
	jand g0126(.dina(n189),.dinb(w_n123_0[0]),.dout(n190),.clk(gclk));
	jand g0127(.dina(w_n161_0[0]),.dinb(w_n154_0[0]),.dout(n191),.clk(gclk));
	jor g0128(.dina(n191),.dinb(n190),.dout(n192),.clk(gclk));
	jand g0129(.dina(w_G307gat_6[0]),.dinb(w_G69gat_6[2]),.dout(n193),.clk(gclk));
	jnot g0130(.din(n193),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n195),.clk(gclk));
	jand g0132(.dina(w_n195_0[1]),.dinb(w_n158_0[0]),.dout(n196),.clk(gclk));
	jnot g0133(.din(w_n196_0[2]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n198),.clk(gclk));
	jor g0135(.dina(w_n198_0[1]),.dinb(w_n155_0[0]),.dout(n199),.clk(gclk));
	jand g0136(.dina(w_dff_B_vi41Mh5Q9_0),.dinb(n197),.dout(n200),.clk(gclk));
	jxor g0137(.dina(w_n200_0[1]),.dinb(w_n156_0[0]),.dout(n201),.clk(gclk));
	jxor g0138(.dina(w_n201_0[1]),.dinb(w_n194_0[1]),.dout(n202),.clk(gclk));
	jxor g0139(.dina(w_n202_0[1]),.dinb(w_n192_0[1]),.dout(n203),.clk(gclk));
	jxor g0140(.dina(w_n203_0[1]),.dinb(w_n188_0[1]),.dout(n204),.clk(gclk));
	jxor g0141(.dina(w_n204_0[1]),.dinb(w_n186_0[1]),.dout(n205),.clk(gclk));
	jxor g0142(.dina(w_n205_0[1]),.dinb(w_n183_0[1]),.dout(n206),.clk(gclk));
	jnot g0143(.din(w_n206_0[1]),.dout(n207),.clk(gclk));
	jxor g0144(.dina(w_n207_0[1]),.dinb(w_n181_0[2]),.dout(n208),.clk(gclk));
	jxor g0145(.dina(n208),.dinb(w_dff_B_wDNz3IFj5_1),.dout(n209),.clk(gclk));
	jxor g0146(.dina(w_n209_0[1]),.dinb(w_n175_0[1]),.dout(n210),.clk(gclk));
	jxor g0147(.dina(w_n210_0[1]),.dinb(w_dff_B_DOxgFj537_1),.dout(w_dff_A_QxM6dCu23_2),.clk(gclk));
	jand g0148(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n212),.clk(gclk));
	jnot g0149(.din(w_n212_0[1]),.dout(n213),.clk(gclk));
	jnot g0150(.din(w_n209_0[0]),.dout(n214),.clk(gclk));
	jor g0151(.dina(n214),.dinb(w_n175_0[0]),.dout(n215),.clk(gclk));
	jor g0152(.dina(w_n210_0[0]),.dinb(w_n170_0[0]),.dout(n216),.clk(gclk));
	jand g0153(.dina(n216),.dinb(w_dff_B_4IAinCvK4_1),.dout(n217),.clk(gclk));
	jand g0154(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n218),.clk(gclk));
	jnot g0155(.din(w_n218_0[1]),.dout(n219),.clk(gclk));
	jor g0156(.dina(w_n207_0[0]),.dinb(w_n181_0[1]),.dout(n220),.clk(gclk));
	jxor g0157(.dina(w_n206_0[0]),.dinb(w_n181_0[0]),.dout(n221),.clk(gclk));
	jor g0158(.dina(n221),.dinb(w_n176_0[0]),.dout(n222),.clk(gclk));
	jand g0159(.dina(n222),.dinb(w_dff_B_Ij7RFoTe0_1),.dout(n223),.clk(gclk));
	jand g0160(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n224),.clk(gclk));
	jnot g0161(.din(n224),.dout(n225),.clk(gclk));
	jand g0162(.dina(w_n204_0[0]),.dinb(w_n186_0[0]),.dout(n226),.clk(gclk));
	jand g0163(.dina(w_n205_0[0]),.dinb(w_n183_0[0]),.dout(n227),.clk(gclk));
	jor g0164(.dina(n227),.dinb(w_dff_B_y8neqvKc3_1),.dout(n228),.clk(gclk));
	jand g0165(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n229),.clk(gclk));
	jnot g0166(.din(n229),.dout(n230),.clk(gclk));
	jand g0167(.dina(w_n202_0[0]),.dinb(w_n192_0[0]),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_n203_0[0]),.dinb(w_n188_0[0]),.dout(n232),.clk(gclk));
	jor g0169(.dina(n232),.dinb(w_dff_B_bmAOyLyk1_1),.dout(n233),.clk(gclk));
	jand g0170(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n234),.clk(gclk));
	jnot g0171(.din(n234),.dout(n235),.clk(gclk));
	jnot g0172(.din(w_n200_0[0]),.dout(n236),.clk(gclk));
	jand g0173(.dina(n236),.dinb(w_n157_0[0]),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_n201_0[0]),.dinb(w_n194_0[0]),.dout(n238),.clk(gclk));
	jor g0175(.dina(n238),.dinb(n237),.dout(n239),.clk(gclk));
	jand g0176(.dina(w_G307gat_5[2]),.dinb(w_G86gat_6[2]),.dout(n240),.clk(gclk));
	jnot g0177(.din(n240),.dout(n241),.clk(gclk));
	jand g0178(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n242),.clk(gclk));
	jand g0179(.dina(w_n242_0[1]),.dinb(w_n198_0[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(w_n243_0[2]),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n245),.clk(gclk));
	jor g0182(.dina(w_n245_0[1]),.dinb(w_n195_0[0]),.dout(n246),.clk(gclk));
	jand g0183(.dina(w_dff_B_dFtM3qTM2_0),.dinb(n244),.dout(n247),.clk(gclk));
	jxor g0184(.dina(w_n247_0[1]),.dinb(w_n196_0[1]),.dout(n248),.clk(gclk));
	jxor g0185(.dina(w_n248_0[1]),.dinb(w_n241_0[1]),.dout(n249),.clk(gclk));
	jxor g0186(.dina(w_n249_0[1]),.dinb(w_n239_0[1]),.dout(n250),.clk(gclk));
	jxor g0187(.dina(w_n250_0[1]),.dinb(w_n235_0[1]),.dout(n251),.clk(gclk));
	jxor g0188(.dina(w_n251_0[1]),.dinb(w_n233_0[1]),.dout(n252),.clk(gclk));
	jxor g0189(.dina(w_n252_0[1]),.dinb(w_n230_0[1]),.dout(n253),.clk(gclk));
	jxor g0190(.dina(w_n253_0[1]),.dinb(w_n228_0[1]),.dout(n254),.clk(gclk));
	jxor g0191(.dina(w_n254_0[1]),.dinb(w_n225_0[1]),.dout(n255),.clk(gclk));
	jnot g0192(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jxor g0193(.dina(w_n256_0[1]),.dinb(w_n223_0[2]),.dout(n257),.clk(gclk));
	jxor g0194(.dina(n257),.dinb(w_dff_B_d8EbkTxD8_1),.dout(n258),.clk(gclk));
	jxor g0195(.dina(w_n258_0[1]),.dinb(w_n217_0[1]),.dout(n259),.clk(gclk));
	jxor g0196(.dina(w_n259_0[1]),.dinb(w_dff_B_DtxLqxqv7_1),.dout(w_dff_A_0JP3jwNj8_2),.clk(gclk));
	jand g0197(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n261),.clk(gclk));
	jnot g0198(.din(w_n261_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(w_n258_0[0]),.dout(n263),.clk(gclk));
	jor g0200(.dina(n263),.dinb(w_n217_0[0]),.dout(n264),.clk(gclk));
	jor g0201(.dina(w_n259_0[0]),.dinb(w_n212_0[0]),.dout(n265),.clk(gclk));
	jand g0202(.dina(n265),.dinb(w_dff_B_yHoAoE6P4_1),.dout(n266),.clk(gclk));
	jand g0203(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n267),.clk(gclk));
	jnot g0204(.din(w_n267_0[1]),.dout(n268),.clk(gclk));
	jor g0205(.dina(w_n256_0[0]),.dinb(w_n223_0[1]),.dout(n269),.clk(gclk));
	jxor g0206(.dina(w_n255_0[0]),.dinb(w_n223_0[0]),.dout(n270),.clk(gclk));
	jor g0207(.dina(n270),.dinb(w_n218_0[0]),.dout(n271),.clk(gclk));
	jand g0208(.dina(n271),.dinb(w_dff_B_Q4fCHPlP0_1),.dout(n272),.clk(gclk));
	jand g0209(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n273),.clk(gclk));
	jnot g0210(.din(n273),.dout(n274),.clk(gclk));
	jand g0211(.dina(w_n253_0[0]),.dinb(w_n228_0[0]),.dout(n275),.clk(gclk));
	jand g0212(.dina(w_n254_0[0]),.dinb(w_n225_0[0]),.dout(n276),.clk(gclk));
	jor g0213(.dina(n276),.dinb(w_dff_B_2zdPCp3j5_1),.dout(n277),.clk(gclk));
	jand g0214(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n278),.clk(gclk));
	jnot g0215(.din(n278),.dout(n279),.clk(gclk));
	jand g0216(.dina(w_n251_0[0]),.dinb(w_n233_0[0]),.dout(n280),.clk(gclk));
	jand g0217(.dina(w_n252_0[0]),.dinb(w_n230_0[0]),.dout(n281),.clk(gclk));
	jor g0218(.dina(n281),.dinb(w_dff_B_yNEAHrJk0_1),.dout(n282),.clk(gclk));
	jand g0219(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(n283),.dout(n284),.clk(gclk));
	jand g0221(.dina(w_n249_0[0]),.dinb(w_n239_0[0]),.dout(n285),.clk(gclk));
	jand g0222(.dina(w_n250_0[0]),.dinb(w_n235_0[0]),.dout(n286),.clk(gclk));
	jor g0223(.dina(n286),.dinb(w_dff_B_YoDQV3J86_1),.dout(n287),.clk(gclk));
	jand g0224(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n288),.clk(gclk));
	jnot g0225(.din(n288),.dout(n289),.clk(gclk));
	jor g0226(.dina(w_n247_0[0]),.dinb(w_n196_0[0]),.dout(n290),.clk(gclk));
	jnot g0227(.din(n290),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n248_0[0]),.dinb(w_n241_0[0]),.dout(n292),.clk(gclk));
	jor g0229(.dina(n292),.dinb(n291),.dout(n293),.clk(gclk));
	jand g0230(.dina(w_G307gat_5[1]),.dinb(w_G103gat_6[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n296_0[1]),.dinb(w_n245_0[0]),.dout(n297),.clk(gclk));
	jnot g0234(.din(w_n297_0[2]),.dout(n298),.clk(gclk));
	jand g0235(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n299),.clk(gclk));
	jor g0236(.dina(w_n299_0[1]),.dinb(w_n242_0[0]),.dout(n300),.clk(gclk));
	jand g0237(.dina(w_dff_B_KO48WI7V7_0),.dinb(n298),.dout(n301),.clk(gclk));
	jxor g0238(.dina(w_n301_0[1]),.dinb(w_n243_0[1]),.dout(n302),.clk(gclk));
	jxor g0239(.dina(w_n302_0[1]),.dinb(w_n295_0[1]),.dout(n303),.clk(gclk));
	jxor g0240(.dina(w_n303_0[1]),.dinb(w_n293_0[1]),.dout(n304),.clk(gclk));
	jxor g0241(.dina(w_n304_0[1]),.dinb(w_n289_0[1]),.dout(n305),.clk(gclk));
	jxor g0242(.dina(w_n305_0[1]),.dinb(w_n287_0[1]),.dout(n306),.clk(gclk));
	jxor g0243(.dina(w_n306_0[1]),.dinb(w_n284_0[1]),.dout(n307),.clk(gclk));
	jxor g0244(.dina(w_n307_0[1]),.dinb(w_n282_0[1]),.dout(n308),.clk(gclk));
	jxor g0245(.dina(w_n308_0[1]),.dinb(w_n279_0[1]),.dout(n309),.clk(gclk));
	jxor g0246(.dina(w_n309_0[1]),.dinb(w_n277_0[1]),.dout(n310),.clk(gclk));
	jxor g0247(.dina(w_n310_0[1]),.dinb(w_n274_0[1]),.dout(n311),.clk(gclk));
	jnot g0248(.din(w_n311_0[1]),.dout(n312),.clk(gclk));
	jxor g0249(.dina(w_n312_0[1]),.dinb(w_n272_0[2]),.dout(n313),.clk(gclk));
	jxor g0250(.dina(n313),.dinb(w_dff_B_NwoMSljy8_1),.dout(n314),.clk(gclk));
	jxor g0251(.dina(w_n314_0[1]),.dinb(w_n266_0[1]),.dout(n315),.clk(gclk));
	jxor g0252(.dina(w_n315_0[1]),.dinb(w_dff_B_8TdGlqOt4_1),.dout(w_dff_A_tDHTbtHD9_2),.clk(gclk));
	jand g0253(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n317),.clk(gclk));
	jnot g0254(.din(w_n317_0[1]),.dout(n318),.clk(gclk));
	jnot g0255(.din(w_n314_0[0]),.dout(n319),.clk(gclk));
	jor g0256(.dina(n319),.dinb(w_n266_0[0]),.dout(n320),.clk(gclk));
	jor g0257(.dina(w_n315_0[0]),.dinb(w_n261_0[0]),.dout(n321),.clk(gclk));
	jand g0258(.dina(n321),.dinb(w_dff_B_KXgzlV1M9_1),.dout(n322),.clk(gclk));
	jand g0259(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n323),.clk(gclk));
	jnot g0260(.din(w_n323_0[1]),.dout(n324),.clk(gclk));
	jor g0261(.dina(w_n312_0[0]),.dinb(w_n272_0[1]),.dout(n325),.clk(gclk));
	jxor g0262(.dina(w_n311_0[0]),.dinb(w_n272_0[0]),.dout(n326),.clk(gclk));
	jor g0263(.dina(n326),.dinb(w_n267_0[0]),.dout(n327),.clk(gclk));
	jand g0264(.dina(n327),.dinb(w_dff_B_GGzwUl4x8_1),.dout(n328),.clk(gclk));
	jand g0265(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n329),.clk(gclk));
	jnot g0266(.din(n329),.dout(n330),.clk(gclk));
	jand g0267(.dina(w_n309_0[0]),.dinb(w_n277_0[0]),.dout(n331),.clk(gclk));
	jand g0268(.dina(w_n310_0[0]),.dinb(w_n274_0[0]),.dout(n332),.clk(gclk));
	jor g0269(.dina(n332),.dinb(w_dff_B_XaXDB1un7_1),.dout(n333),.clk(gclk));
	jand g0270(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n334),.clk(gclk));
	jnot g0271(.din(n334),.dout(n335),.clk(gclk));
	jand g0272(.dina(w_n307_0[0]),.dinb(w_n282_0[0]),.dout(n336),.clk(gclk));
	jand g0273(.dina(w_n308_0[0]),.dinb(w_n279_0[0]),.dout(n337),.clk(gclk));
	jor g0274(.dina(n337),.dinb(w_dff_B_3fp6Nyge0_1),.dout(n338),.clk(gclk));
	jand g0275(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n339),.clk(gclk));
	jnot g0276(.din(n339),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_n305_0[0]),.dinb(w_n287_0[0]),.dout(n341),.clk(gclk));
	jand g0278(.dina(w_n306_0[0]),.dinb(w_n284_0[0]),.dout(n342),.clk(gclk));
	jor g0279(.dina(n342),.dinb(w_dff_B_TBd7wztu5_1),.dout(n343),.clk(gclk));
	jand g0280(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n344),.clk(gclk));
	jnot g0281(.din(n344),.dout(n345),.clk(gclk));
	jand g0282(.dina(w_n303_0[0]),.dinb(w_n293_0[0]),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_n304_0[0]),.dinb(w_n289_0[0]),.dout(n347),.clk(gclk));
	jor g0284(.dina(n347),.dinb(w_dff_B_ir1ZwmwY5_1),.dout(n348),.clk(gclk));
	jand g0285(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n349),.clk(gclk));
	jnot g0286(.din(n349),.dout(n350),.clk(gclk));
	jor g0287(.dina(w_n301_0[0]),.dinb(w_n243_0[0]),.dout(n351),.clk(gclk));
	jnot g0288(.din(n351),.dout(n352),.clk(gclk));
	jand g0289(.dina(w_n302_0[0]),.dinb(w_n295_0[0]),.dout(n353),.clk(gclk));
	jor g0290(.dina(n353),.dinb(n352),.dout(n354),.clk(gclk));
	jand g0291(.dina(w_G307gat_5[0]),.dinb(w_G120gat_6[2]),.dout(n355),.clk(gclk));
	jnot g0292(.din(n355),.dout(n356),.clk(gclk));
	jand g0293(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n357),.clk(gclk));
	jand g0294(.dina(w_n357_0[1]),.dinb(w_n299_0[0]),.dout(n358),.clk(gclk));
	jnot g0295(.din(w_n358_0[2]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n360),.clk(gclk));
	jor g0297(.dina(w_n360_0[1]),.dinb(w_n296_0[0]),.dout(n361),.clk(gclk));
	jand g0298(.dina(w_dff_B_x2mpqGpk1_0),.dinb(n359),.dout(n362),.clk(gclk));
	jxor g0299(.dina(w_n362_0[1]),.dinb(w_n297_0[1]),.dout(n363),.clk(gclk));
	jxor g0300(.dina(w_n363_0[1]),.dinb(w_n356_0[1]),.dout(n364),.clk(gclk));
	jxor g0301(.dina(w_n364_0[1]),.dinb(w_n354_0[1]),.dout(n365),.clk(gclk));
	jxor g0302(.dina(w_n365_0[1]),.dinb(w_n350_0[1]),.dout(n366),.clk(gclk));
	jxor g0303(.dina(w_n366_0[1]),.dinb(w_n348_0[1]),.dout(n367),.clk(gclk));
	jxor g0304(.dina(w_n367_0[1]),.dinb(w_n345_0[1]),.dout(n368),.clk(gclk));
	jxor g0305(.dina(w_n368_0[1]),.dinb(w_n343_0[1]),.dout(n369),.clk(gclk));
	jxor g0306(.dina(w_n369_0[1]),.dinb(w_n340_0[1]),.dout(n370),.clk(gclk));
	jxor g0307(.dina(w_n370_0[1]),.dinb(w_n338_0[1]),.dout(n371),.clk(gclk));
	jxor g0308(.dina(w_n371_0[1]),.dinb(w_n335_0[1]),.dout(n372),.clk(gclk));
	jxor g0309(.dina(w_n372_0[1]),.dinb(w_n333_0[1]),.dout(n373),.clk(gclk));
	jxor g0310(.dina(w_n373_0[1]),.dinb(w_n330_0[1]),.dout(n374),.clk(gclk));
	jnot g0311(.din(w_n374_0[1]),.dout(n375),.clk(gclk));
	jxor g0312(.dina(w_n375_0[1]),.dinb(w_n328_0[2]),.dout(n376),.clk(gclk));
	jxor g0313(.dina(n376),.dinb(w_dff_B_eZQ8FN4T1_1),.dout(n377),.clk(gclk));
	jxor g0314(.dina(w_n377_0[1]),.dinb(w_n322_0[1]),.dout(n378),.clk(gclk));
	jxor g0315(.dina(w_n378_0[1]),.dinb(w_dff_B_KsiC9Zr79_1),.dout(w_dff_A_yY8yxN6c1_2),.clk(gclk));
	jand g0316(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n380),.clk(gclk));
	jnot g0317(.din(w_n380_0[1]),.dout(n381),.clk(gclk));
	jnot g0318(.din(w_n377_0[0]),.dout(n382),.clk(gclk));
	jor g0319(.dina(n382),.dinb(w_n322_0[0]),.dout(n383),.clk(gclk));
	jor g0320(.dina(w_n378_0[0]),.dinb(w_n317_0[0]),.dout(n384),.clk(gclk));
	jand g0321(.dina(n384),.dinb(w_dff_B_kGQLwCQb2_1),.dout(n385),.clk(gclk));
	jand g0322(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n386),.clk(gclk));
	jnot g0323(.din(w_n386_0[1]),.dout(n387),.clk(gclk));
	jor g0324(.dina(w_n375_0[0]),.dinb(w_n328_0[1]),.dout(n388),.clk(gclk));
	jxor g0325(.dina(w_n374_0[0]),.dinb(w_n328_0[0]),.dout(n389),.clk(gclk));
	jor g0326(.dina(n389),.dinb(w_n323_0[0]),.dout(n390),.clk(gclk));
	jand g0327(.dina(n390),.dinb(w_dff_B_mGfMoIar4_1),.dout(n391),.clk(gclk));
	jand g0328(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n392),.clk(gclk));
	jnot g0329(.din(n392),.dout(n393),.clk(gclk));
	jand g0330(.dina(w_n372_0[0]),.dinb(w_n333_0[0]),.dout(n394),.clk(gclk));
	jand g0331(.dina(w_n373_0[0]),.dinb(w_n330_0[0]),.dout(n395),.clk(gclk));
	jor g0332(.dina(n395),.dinb(w_dff_B_Bs4DgqRc7_1),.dout(n396),.clk(gclk));
	jand g0333(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n397),.clk(gclk));
	jnot g0334(.din(n397),.dout(n398),.clk(gclk));
	jand g0335(.dina(w_n370_0[0]),.dinb(w_n338_0[0]),.dout(n399),.clk(gclk));
	jand g0336(.dina(w_n371_0[0]),.dinb(w_n335_0[0]),.dout(n400),.clk(gclk));
	jor g0337(.dina(n400),.dinb(w_dff_B_Iyryb7Ag3_1),.dout(n401),.clk(gclk));
	jand g0338(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n402),.clk(gclk));
	jnot g0339(.din(n402),.dout(n403),.clk(gclk));
	jand g0340(.dina(w_n368_0[0]),.dinb(w_n343_0[0]),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_n369_0[0]),.dinb(w_n340_0[0]),.dout(n405),.clk(gclk));
	jor g0342(.dina(n405),.dinb(w_dff_B_hSfTyuhW6_1),.dout(n406),.clk(gclk));
	jand g0343(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n407),.clk(gclk));
	jnot g0344(.din(n407),.dout(n408),.clk(gclk));
	jand g0345(.dina(w_n366_0[0]),.dinb(w_n348_0[0]),.dout(n409),.clk(gclk));
	jand g0346(.dina(w_n367_0[0]),.dinb(w_n345_0[0]),.dout(n410),.clk(gclk));
	jor g0347(.dina(n410),.dinb(w_dff_B_YL95S5n31_1),.dout(n411),.clk(gclk));
	jand g0348(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n412),.clk(gclk));
	jnot g0349(.din(n412),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n364_0[0]),.dinb(w_n354_0[0]),.dout(n414),.clk(gclk));
	jand g0351(.dina(w_n365_0[0]),.dinb(w_n350_0[0]),.dout(n415),.clk(gclk));
	jor g0352(.dina(n415),.dinb(w_dff_B_hvejbr7D5_1),.dout(n416),.clk(gclk));
	jand g0353(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n417),.clk(gclk));
	jnot g0354(.din(n417),.dout(n418),.clk(gclk));
	jor g0355(.dina(w_n362_0[0]),.dinb(w_n297_0[0]),.dout(n419),.clk(gclk));
	jand g0356(.dina(w_n363_0[0]),.dinb(w_n356_0[0]),.dout(n420),.clk(gclk));
	jnot g0357(.din(n420),.dout(n421),.clk(gclk));
	jand g0358(.dina(n421),.dinb(w_dff_B_9n09owlS0_1),.dout(n422),.clk(gclk));
	jnot g0359(.din(n422),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_G307gat_4[2]),.dinb(w_G137gat_6[2]),.dout(n424),.clk(gclk));
	jnot g0361(.din(n424),.dout(n425),.clk(gclk));
	jand g0362(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n426),.clk(gclk));
	jand g0363(.dina(w_n426_0[1]),.dinb(w_n360_0[0]),.dout(n427),.clk(gclk));
	jnot g0364(.din(w_n427_0[2]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n429),.clk(gclk));
	jor g0366(.dina(w_n429_0[1]),.dinb(w_n357_0[0]),.dout(n430),.clk(gclk));
	jand g0367(.dina(w_dff_B_pnrgftmm8_0),.dinb(n428),.dout(n431),.clk(gclk));
	jxor g0368(.dina(w_n431_0[1]),.dinb(w_n358_0[1]),.dout(n432),.clk(gclk));
	jxor g0369(.dina(w_n432_0[1]),.dinb(w_n425_0[1]),.dout(n433),.clk(gclk));
	jxor g0370(.dina(w_n433_0[1]),.dinb(w_n423_0[1]),.dout(n434),.clk(gclk));
	jxor g0371(.dina(w_n434_0[1]),.dinb(w_n418_0[1]),.dout(n435),.clk(gclk));
	jxor g0372(.dina(w_n435_0[1]),.dinb(w_n416_0[1]),.dout(n436),.clk(gclk));
	jxor g0373(.dina(w_n436_0[1]),.dinb(w_n413_0[1]),.dout(n437),.clk(gclk));
	jxor g0374(.dina(w_n437_0[1]),.dinb(w_n411_0[1]),.dout(n438),.clk(gclk));
	jxor g0375(.dina(w_n438_0[1]),.dinb(w_n408_0[1]),.dout(n439),.clk(gclk));
	jxor g0376(.dina(w_n439_0[1]),.dinb(w_n406_0[1]),.dout(n440),.clk(gclk));
	jxor g0377(.dina(w_n440_0[1]),.dinb(w_n403_0[1]),.dout(n441),.clk(gclk));
	jxor g0378(.dina(w_n441_0[1]),.dinb(w_n401_0[1]),.dout(n442),.clk(gclk));
	jxor g0379(.dina(w_n442_0[1]),.dinb(w_n398_0[1]),.dout(n443),.clk(gclk));
	jxor g0380(.dina(w_n443_0[1]),.dinb(w_n396_0[1]),.dout(n444),.clk(gclk));
	jxor g0381(.dina(w_n444_0[1]),.dinb(w_n393_0[1]),.dout(n445),.clk(gclk));
	jnot g0382(.din(w_n445_0[1]),.dout(n446),.clk(gclk));
	jxor g0383(.dina(w_n446_0[1]),.dinb(w_n391_0[2]),.dout(n447),.clk(gclk));
	jxor g0384(.dina(n447),.dinb(w_dff_B_gBOEeCXE2_1),.dout(n448),.clk(gclk));
	jxor g0385(.dina(w_n448_0[1]),.dinb(w_n385_0[1]),.dout(n449),.clk(gclk));
	jxor g0386(.dina(w_n449_0[1]),.dinb(w_dff_B_IFgWrum80_1),.dout(w_dff_A_fbgsIzQB8_2),.clk(gclk));
	jand g0387(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n451),.clk(gclk));
	jnot g0388(.din(w_n451_0[1]),.dout(n452),.clk(gclk));
	jnot g0389(.din(w_n448_0[0]),.dout(n453),.clk(gclk));
	jor g0390(.dina(n453),.dinb(w_n385_0[0]),.dout(n454),.clk(gclk));
	jor g0391(.dina(w_n449_0[0]),.dinb(w_n380_0[0]),.dout(n455),.clk(gclk));
	jand g0392(.dina(n455),.dinb(w_dff_B_V2FILeAh0_1),.dout(n456),.clk(gclk));
	jand g0393(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n457),.clk(gclk));
	jnot g0394(.din(w_n457_0[1]),.dout(n458),.clk(gclk));
	jor g0395(.dina(w_n446_0[0]),.dinb(w_n391_0[1]),.dout(n459),.clk(gclk));
	jxor g0396(.dina(w_n445_0[0]),.dinb(w_n391_0[0]),.dout(n460),.clk(gclk));
	jor g0397(.dina(n460),.dinb(w_n386_0[0]),.dout(n461),.clk(gclk));
	jand g0398(.dina(n461),.dinb(w_dff_B_4nstmJjP9_1),.dout(n462),.clk(gclk));
	jand g0399(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n463),.clk(gclk));
	jnot g0400(.din(n463),.dout(n464),.clk(gclk));
	jand g0401(.dina(w_n443_0[0]),.dinb(w_n396_0[0]),.dout(n465),.clk(gclk));
	jand g0402(.dina(w_n444_0[0]),.dinb(w_n393_0[0]),.dout(n466),.clk(gclk));
	jor g0403(.dina(n466),.dinb(w_dff_B_X5omvm2U0_1),.dout(n467),.clk(gclk));
	jand g0404(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n468),.clk(gclk));
	jnot g0405(.din(n468),.dout(n469),.clk(gclk));
	jand g0406(.dina(w_n441_0[0]),.dinb(w_n401_0[0]),.dout(n470),.clk(gclk));
	jand g0407(.dina(w_n442_0[0]),.dinb(w_n398_0[0]),.dout(n471),.clk(gclk));
	jor g0408(.dina(n471),.dinb(w_dff_B_U0htOr0J6_1),.dout(n472),.clk(gclk));
	jand g0409(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n473),.clk(gclk));
	jnot g0410(.din(n473),.dout(n474),.clk(gclk));
	jand g0411(.dina(w_n439_0[0]),.dinb(w_n406_0[0]),.dout(n475),.clk(gclk));
	jand g0412(.dina(w_n440_0[0]),.dinb(w_n403_0[0]),.dout(n476),.clk(gclk));
	jor g0413(.dina(n476),.dinb(w_dff_B_GXqD2o435_1),.dout(n477),.clk(gclk));
	jand g0414(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n478),.clk(gclk));
	jnot g0415(.din(n478),.dout(n479),.clk(gclk));
	jand g0416(.dina(w_n437_0[0]),.dinb(w_n411_0[0]),.dout(n480),.clk(gclk));
	jand g0417(.dina(w_n438_0[0]),.dinb(w_n408_0[0]),.dout(n481),.clk(gclk));
	jor g0418(.dina(n481),.dinb(w_dff_B_6HH7rVy35_1),.dout(n482),.clk(gclk));
	jand g0419(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n435_0[0]),.dinb(w_n416_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n436_0[0]),.dinb(w_n413_0[0]),.dout(n486),.clk(gclk));
	jor g0423(.dina(n486),.dinb(w_dff_B_MhBtpbU40_1),.dout(n487),.clk(gclk));
	jand g0424(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n433_0[0]),.dinb(w_n423_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n434_0[0]),.dinb(w_n418_0[0]),.dout(n491),.clk(gclk));
	jor g0428(.dina(n491),.dinb(w_dff_B_1Eksn2Zn3_1),.dout(n492),.clk(gclk));
	jand g0429(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jor g0431(.dina(w_n431_0[0]),.dinb(w_n358_0[0]),.dout(n495),.clk(gclk));
	jand g0432(.dina(w_n432_0[0]),.dinb(w_n425_0[0]),.dout(n496),.clk(gclk));
	jnot g0433(.din(n496),.dout(n497),.clk(gclk));
	jand g0434(.dina(n497),.dinb(w_dff_B_jCZ6uKDN9_1),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_G307gat_4[1]),.dinb(w_G154gat_6[2]),.dout(n500),.clk(gclk));
	jnot g0437(.din(n500),.dout(n501),.clk(gclk));
	jand g0438(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n502),.clk(gclk));
	jand g0439(.dina(w_n502_0[1]),.dinb(w_n429_0[0]),.dout(n503),.clk(gclk));
	jnot g0440(.din(w_n503_0[2]),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n505),.clk(gclk));
	jor g0442(.dina(w_n505_0[1]),.dinb(w_n426_0[0]),.dout(n506),.clk(gclk));
	jand g0443(.dina(w_dff_B_JIdhCC2w7_0),.dinb(n504),.dout(n507),.clk(gclk));
	jxor g0444(.dina(w_n507_0[1]),.dinb(w_n427_0[1]),.dout(n508),.clk(gclk));
	jxor g0445(.dina(w_n508_0[1]),.dinb(w_n501_0[1]),.dout(n509),.clk(gclk));
	jxor g0446(.dina(w_n509_0[1]),.dinb(w_n499_0[1]),.dout(n510),.clk(gclk));
	jxor g0447(.dina(w_n510_0[1]),.dinb(w_n494_0[1]),.dout(n511),.clk(gclk));
	jxor g0448(.dina(w_n511_0[1]),.dinb(w_n492_0[1]),.dout(n512),.clk(gclk));
	jxor g0449(.dina(w_n512_0[1]),.dinb(w_n489_0[1]),.dout(n513),.clk(gclk));
	jxor g0450(.dina(w_n513_0[1]),.dinb(w_n487_0[1]),.dout(n514),.clk(gclk));
	jxor g0451(.dina(w_n514_0[1]),.dinb(w_n484_0[1]),.dout(n515),.clk(gclk));
	jxor g0452(.dina(w_n515_0[1]),.dinb(w_n482_0[1]),.dout(n516),.clk(gclk));
	jxor g0453(.dina(w_n516_0[1]),.dinb(w_n479_0[1]),.dout(n517),.clk(gclk));
	jxor g0454(.dina(w_n517_0[1]),.dinb(w_n477_0[1]),.dout(n518),.clk(gclk));
	jxor g0455(.dina(w_n518_0[1]),.dinb(w_n474_0[1]),.dout(n519),.clk(gclk));
	jxor g0456(.dina(w_n519_0[1]),.dinb(w_n472_0[1]),.dout(n520),.clk(gclk));
	jxor g0457(.dina(w_n520_0[1]),.dinb(w_n469_0[1]),.dout(n521),.clk(gclk));
	jxor g0458(.dina(w_n521_0[1]),.dinb(w_n467_0[1]),.dout(n522),.clk(gclk));
	jxor g0459(.dina(w_n522_0[1]),.dinb(w_n464_0[1]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[1]),.dout(n524),.clk(gclk));
	jxor g0461(.dina(w_n524_0[1]),.dinb(w_n462_0[2]),.dout(n525),.clk(gclk));
	jxor g0462(.dina(n525),.dinb(w_dff_B_SB9jIKZE4_1),.dout(n526),.clk(gclk));
	jxor g0463(.dina(w_n526_0[1]),.dinb(w_n456_0[1]),.dout(n527),.clk(gclk));
	jxor g0464(.dina(w_n527_0[1]),.dinb(w_dff_B_EX4MsRm61_1),.dout(w_dff_A_DQUJXFRm8_2),.clk(gclk));
	jand g0465(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n529),.clk(gclk));
	jnot g0466(.din(w_n529_0[1]),.dout(n530),.clk(gclk));
	jnot g0467(.din(w_n526_0[0]),.dout(n531),.clk(gclk));
	jor g0468(.dina(n531),.dinb(w_n456_0[0]),.dout(n532),.clk(gclk));
	jor g0469(.dina(w_n527_0[0]),.dinb(w_n451_0[0]),.dout(n533),.clk(gclk));
	jand g0470(.dina(n533),.dinb(w_dff_B_os8dMX4n3_1),.dout(n534),.clk(gclk));
	jand g0471(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n535),.clk(gclk));
	jnot g0472(.din(w_n535_0[1]),.dout(n536),.clk(gclk));
	jor g0473(.dina(w_n524_0[0]),.dinb(w_n462_0[1]),.dout(n537),.clk(gclk));
	jxor g0474(.dina(w_n523_0[0]),.dinb(w_n462_0[0]),.dout(n538),.clk(gclk));
	jor g0475(.dina(n538),.dinb(w_n457_0[0]),.dout(n539),.clk(gclk));
	jand g0476(.dina(n539),.dinb(w_dff_B_Wx8gVA3f4_1),.dout(n540),.clk(gclk));
	jand g0477(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n541),.clk(gclk));
	jnot g0478(.din(n541),.dout(n542),.clk(gclk));
	jand g0479(.dina(w_n521_0[0]),.dinb(w_n467_0[0]),.dout(n543),.clk(gclk));
	jand g0480(.dina(w_n522_0[0]),.dinb(w_n464_0[0]),.dout(n544),.clk(gclk));
	jor g0481(.dina(n544),.dinb(w_dff_B_L2nPKQmm2_1),.dout(n545),.clk(gclk));
	jand g0482(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n546),.clk(gclk));
	jnot g0483(.din(n546),.dout(n547),.clk(gclk));
	jand g0484(.dina(w_n519_0[0]),.dinb(w_n472_0[0]),.dout(n548),.clk(gclk));
	jand g0485(.dina(w_n520_0[0]),.dinb(w_n469_0[0]),.dout(n549),.clk(gclk));
	jor g0486(.dina(n549),.dinb(w_dff_B_JMosQLe99_1),.dout(n550),.clk(gclk));
	jand g0487(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n551),.clk(gclk));
	jnot g0488(.din(n551),.dout(n552),.clk(gclk));
	jand g0489(.dina(w_n517_0[0]),.dinb(w_n477_0[0]),.dout(n553),.clk(gclk));
	jand g0490(.dina(w_n518_0[0]),.dinb(w_n474_0[0]),.dout(n554),.clk(gclk));
	jor g0491(.dina(n554),.dinb(w_dff_B_uy2SawVe8_1),.dout(n555),.clk(gclk));
	jand g0492(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n556),.clk(gclk));
	jnot g0493(.din(n556),.dout(n557),.clk(gclk));
	jand g0494(.dina(w_n515_0[0]),.dinb(w_n482_0[0]),.dout(n558),.clk(gclk));
	jand g0495(.dina(w_n516_0[0]),.dinb(w_n479_0[0]),.dout(n559),.clk(gclk));
	jor g0496(.dina(n559),.dinb(w_dff_B_P1aw5ykX6_1),.dout(n560),.clk(gclk));
	jand g0497(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n561),.clk(gclk));
	jnot g0498(.din(n561),.dout(n562),.clk(gclk));
	jand g0499(.dina(w_n513_0[0]),.dinb(w_n487_0[0]),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n514_0[0]),.dinb(w_n484_0[0]),.dout(n564),.clk(gclk));
	jor g0501(.dina(n564),.dinb(w_dff_B_npGZULCR8_1),.dout(n565),.clk(gclk));
	jand g0502(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n566),.clk(gclk));
	jnot g0503(.din(n566),.dout(n567),.clk(gclk));
	jand g0504(.dina(w_n511_0[0]),.dinb(w_n492_0[0]),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n512_0[0]),.dinb(w_n489_0[0]),.dout(n569),.clk(gclk));
	jor g0506(.dina(n569),.dinb(w_dff_B_LYvvcZlp2_1),.dout(n570),.clk(gclk));
	jand g0507(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n571),.clk(gclk));
	jnot g0508(.din(n571),.dout(n572),.clk(gclk));
	jand g0509(.dina(w_n509_0[0]),.dinb(w_n499_0[0]),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n510_0[0]),.dinb(w_n494_0[0]),.dout(n574),.clk(gclk));
	jor g0511(.dina(n574),.dinb(w_dff_B_sfcCpwer7_1),.dout(n575),.clk(gclk));
	jand g0512(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n576),.clk(gclk));
	jnot g0513(.din(n576),.dout(n577),.clk(gclk));
	jor g0514(.dina(w_n507_0[0]),.dinb(w_n427_0[0]),.dout(n578),.clk(gclk));
	jand g0515(.dina(w_n508_0[0]),.dinb(w_n501_0[0]),.dout(n579),.clk(gclk));
	jnot g0516(.din(n579),.dout(n580),.clk(gclk));
	jand g0517(.dina(n580),.dinb(w_dff_B_6q58Zi7A0_1),.dout(n581),.clk(gclk));
	jnot g0518(.din(n581),.dout(n582),.clk(gclk));
	jand g0519(.dina(w_G307gat_4[0]),.dinb(w_G171gat_6[2]),.dout(n583),.clk(gclk));
	jnot g0520(.din(n583),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n585),.clk(gclk));
	jand g0522(.dina(w_n585_0[1]),.dinb(w_n505_0[0]),.dout(n586),.clk(gclk));
	jnot g0523(.din(w_n586_0[2]),.dout(n587),.clk(gclk));
	jand g0524(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n588),.clk(gclk));
	jor g0525(.dina(w_n588_0[1]),.dinb(w_n502_0[0]),.dout(n589),.clk(gclk));
	jand g0526(.dina(w_dff_B_SDciChy19_0),.dinb(n587),.dout(n590),.clk(gclk));
	jxor g0527(.dina(w_n590_0[1]),.dinb(w_n503_0[1]),.dout(n591),.clk(gclk));
	jxor g0528(.dina(w_n591_0[1]),.dinb(w_n584_0[1]),.dout(n592),.clk(gclk));
	jxor g0529(.dina(w_n592_0[1]),.dinb(w_n582_0[1]),.dout(n593),.clk(gclk));
	jxor g0530(.dina(w_n593_0[1]),.dinb(w_n577_0[1]),.dout(n594),.clk(gclk));
	jxor g0531(.dina(w_n594_0[1]),.dinb(w_n575_0[1]),.dout(n595),.clk(gclk));
	jxor g0532(.dina(w_n595_0[1]),.dinb(w_n572_0[1]),.dout(n596),.clk(gclk));
	jxor g0533(.dina(w_n596_0[1]),.dinb(w_n570_0[1]),.dout(n597),.clk(gclk));
	jxor g0534(.dina(w_n597_0[1]),.dinb(w_n567_0[1]),.dout(n598),.clk(gclk));
	jxor g0535(.dina(w_n598_0[1]),.dinb(w_n565_0[1]),.dout(n599),.clk(gclk));
	jxor g0536(.dina(w_n599_0[1]),.dinb(w_n562_0[1]),.dout(n600),.clk(gclk));
	jxor g0537(.dina(w_n600_0[1]),.dinb(w_n560_0[1]),.dout(n601),.clk(gclk));
	jxor g0538(.dina(w_n601_0[1]),.dinb(w_n557_0[1]),.dout(n602),.clk(gclk));
	jxor g0539(.dina(w_n602_0[1]),.dinb(w_n555_0[1]),.dout(n603),.clk(gclk));
	jxor g0540(.dina(w_n603_0[1]),.dinb(w_n552_0[1]),.dout(n604),.clk(gclk));
	jxor g0541(.dina(w_n604_0[1]),.dinb(w_n550_0[1]),.dout(n605),.clk(gclk));
	jxor g0542(.dina(w_n605_0[1]),.dinb(w_n547_0[1]),.dout(n606),.clk(gclk));
	jxor g0543(.dina(w_n606_0[1]),.dinb(w_n545_0[1]),.dout(n607),.clk(gclk));
	jxor g0544(.dina(w_n607_0[1]),.dinb(w_n542_0[1]),.dout(n608),.clk(gclk));
	jnot g0545(.din(w_n608_0[1]),.dout(n609),.clk(gclk));
	jxor g0546(.dina(w_n609_0[1]),.dinb(w_n540_0[2]),.dout(n610),.clk(gclk));
	jxor g0547(.dina(n610),.dinb(w_dff_B_3mtpIpHT8_1),.dout(n611),.clk(gclk));
	jxor g0548(.dina(w_n611_0[1]),.dinb(w_n534_0[1]),.dout(n612),.clk(gclk));
	jxor g0549(.dina(w_n612_0[1]),.dinb(w_dff_B_pnCMdMee4_1),.dout(w_dff_A_8ScMJPuv8_2),.clk(gclk));
	jand g0550(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n614),.clk(gclk));
	jnot g0551(.din(w_n614_0[1]),.dout(n615),.clk(gclk));
	jnot g0552(.din(w_n611_0[0]),.dout(n616),.clk(gclk));
	jor g0553(.dina(n616),.dinb(w_n534_0[0]),.dout(n617),.clk(gclk));
	jor g0554(.dina(w_n612_0[0]),.dinb(w_n529_0[0]),.dout(n618),.clk(gclk));
	jand g0555(.dina(n618),.dinb(w_dff_B_MJFHgnav4_1),.dout(n619),.clk(gclk));
	jand g0556(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n620),.clk(gclk));
	jnot g0557(.din(w_n620_0[1]),.dout(n621),.clk(gclk));
	jor g0558(.dina(w_n609_0[0]),.dinb(w_n540_0[1]),.dout(n622),.clk(gclk));
	jxor g0559(.dina(w_n608_0[0]),.dinb(w_n540_0[0]),.dout(n623),.clk(gclk));
	jor g0560(.dina(n623),.dinb(w_n535_0[0]),.dout(n624),.clk(gclk));
	jand g0561(.dina(n624),.dinb(w_dff_B_3ol2YPqu2_1),.dout(n625),.clk(gclk));
	jand g0562(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n626),.clk(gclk));
	jnot g0563(.din(n626),.dout(n627),.clk(gclk));
	jand g0564(.dina(w_n606_0[0]),.dinb(w_n545_0[0]),.dout(n628),.clk(gclk));
	jand g0565(.dina(w_n607_0[0]),.dinb(w_n542_0[0]),.dout(n629),.clk(gclk));
	jor g0566(.dina(n629),.dinb(w_dff_B_VlAwclpH3_1),.dout(n630),.clk(gclk));
	jand g0567(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n631),.clk(gclk));
	jnot g0568(.din(n631),.dout(n632),.clk(gclk));
	jand g0569(.dina(w_n604_0[0]),.dinb(w_n550_0[0]),.dout(n633),.clk(gclk));
	jand g0570(.dina(w_n605_0[0]),.dinb(w_n547_0[0]),.dout(n634),.clk(gclk));
	jor g0571(.dina(n634),.dinb(w_dff_B_aD7x3mA87_1),.dout(n635),.clk(gclk));
	jand g0572(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n636),.clk(gclk));
	jnot g0573(.din(n636),.dout(n637),.clk(gclk));
	jand g0574(.dina(w_n602_0[0]),.dinb(w_n555_0[0]),.dout(n638),.clk(gclk));
	jand g0575(.dina(w_n603_0[0]),.dinb(w_n552_0[0]),.dout(n639),.clk(gclk));
	jor g0576(.dina(n639),.dinb(w_dff_B_1euSCDwy0_1),.dout(n640),.clk(gclk));
	jand g0577(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n641),.clk(gclk));
	jnot g0578(.din(n641),.dout(n642),.clk(gclk));
	jand g0579(.dina(w_n600_0[0]),.dinb(w_n560_0[0]),.dout(n643),.clk(gclk));
	jand g0580(.dina(w_n601_0[0]),.dinb(w_n557_0[0]),.dout(n644),.clk(gclk));
	jor g0581(.dina(n644),.dinb(w_dff_B_aQcRGXAd3_1),.dout(n645),.clk(gclk));
	jand g0582(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n646),.clk(gclk));
	jnot g0583(.din(n646),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_n598_0[0]),.dinb(w_n565_0[0]),.dout(n648),.clk(gclk));
	jand g0585(.dina(w_n599_0[0]),.dinb(w_n562_0[0]),.dout(n649),.clk(gclk));
	jor g0586(.dina(n649),.dinb(w_dff_B_X2riWvgE7_1),.dout(n650),.clk(gclk));
	jand g0587(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n651),.clk(gclk));
	jnot g0588(.din(n651),.dout(n652),.clk(gclk));
	jand g0589(.dina(w_n596_0[0]),.dinb(w_n570_0[0]),.dout(n653),.clk(gclk));
	jand g0590(.dina(w_n597_0[0]),.dinb(w_n567_0[0]),.dout(n654),.clk(gclk));
	jor g0591(.dina(n654),.dinb(w_dff_B_iYHSkoAI3_1),.dout(n655),.clk(gclk));
	jand g0592(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n656),.clk(gclk));
	jnot g0593(.din(n656),.dout(n657),.clk(gclk));
	jand g0594(.dina(w_n594_0[0]),.dinb(w_n575_0[0]),.dout(n658),.clk(gclk));
	jand g0595(.dina(w_n595_0[0]),.dinb(w_n572_0[0]),.dout(n659),.clk(gclk));
	jor g0596(.dina(n659),.dinb(w_dff_B_HLJpNWGj5_1),.dout(n660),.clk(gclk));
	jand g0597(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n661),.clk(gclk));
	jnot g0598(.din(n661),.dout(n662),.clk(gclk));
	jand g0599(.dina(w_n592_0[0]),.dinb(w_n582_0[0]),.dout(n663),.clk(gclk));
	jand g0600(.dina(w_n593_0[0]),.dinb(w_n577_0[0]),.dout(n664),.clk(gclk));
	jor g0601(.dina(n664),.dinb(w_dff_B_YlGTExVH1_1),.dout(n665),.clk(gclk));
	jand g0602(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n666),.clk(gclk));
	jnot g0603(.din(n666),.dout(n667),.clk(gclk));
	jor g0604(.dina(w_n590_0[0]),.dinb(w_n503_0[0]),.dout(n668),.clk(gclk));
	jand g0605(.dina(w_n591_0[0]),.dinb(w_n584_0[0]),.dout(n669),.clk(gclk));
	jnot g0606(.din(n669),.dout(n670),.clk(gclk));
	jand g0607(.dina(n670),.dinb(w_dff_B_bX1BMdYa4_1),.dout(n671),.clk(gclk));
	jnot g0608(.din(n671),.dout(n672),.clk(gclk));
	jand g0609(.dina(w_G307gat_3[2]),.dinb(w_G188gat_6[2]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n675_0[1]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jnot g0613(.din(w_n676_0[2]),.dout(n677),.clk(gclk));
	jand g0614(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n678),.clk(gclk));
	jor g0615(.dina(w_n678_0[1]),.dinb(w_n585_0[0]),.dout(n679),.clk(gclk));
	jand g0616(.dina(w_dff_B_HZOk2ILt2_0),.dinb(n677),.dout(n680),.clk(gclk));
	jxor g0617(.dina(w_n680_0[1]),.dinb(w_n586_0[1]),.dout(n681),.clk(gclk));
	jxor g0618(.dina(w_n681_0[1]),.dinb(w_n674_0[1]),.dout(n682),.clk(gclk));
	jxor g0619(.dina(w_n682_0[1]),.dinb(w_n672_0[1]),.dout(n683),.clk(gclk));
	jxor g0620(.dina(w_n683_0[1]),.dinb(w_n667_0[1]),.dout(n684),.clk(gclk));
	jxor g0621(.dina(w_n684_0[1]),.dinb(w_n665_0[1]),.dout(n685),.clk(gclk));
	jxor g0622(.dina(w_n685_0[1]),.dinb(w_n662_0[1]),.dout(n686),.clk(gclk));
	jxor g0623(.dina(w_n686_0[1]),.dinb(w_n660_0[1]),.dout(n687),.clk(gclk));
	jxor g0624(.dina(w_n687_0[1]),.dinb(w_n657_0[1]),.dout(n688),.clk(gclk));
	jxor g0625(.dina(w_n688_0[1]),.dinb(w_n655_0[1]),.dout(n689),.clk(gclk));
	jxor g0626(.dina(w_n689_0[1]),.dinb(w_n652_0[1]),.dout(n690),.clk(gclk));
	jxor g0627(.dina(w_n690_0[1]),.dinb(w_n650_0[1]),.dout(n691),.clk(gclk));
	jxor g0628(.dina(w_n691_0[1]),.dinb(w_n647_0[1]),.dout(n692),.clk(gclk));
	jxor g0629(.dina(w_n692_0[1]),.dinb(w_n645_0[1]),.dout(n693),.clk(gclk));
	jxor g0630(.dina(w_n693_0[1]),.dinb(w_n642_0[1]),.dout(n694),.clk(gclk));
	jxor g0631(.dina(w_n694_0[1]),.dinb(w_n640_0[1]),.dout(n695),.clk(gclk));
	jxor g0632(.dina(w_n695_0[1]),.dinb(w_n637_0[1]),.dout(n696),.clk(gclk));
	jxor g0633(.dina(w_n696_0[1]),.dinb(w_n635_0[1]),.dout(n697),.clk(gclk));
	jxor g0634(.dina(w_n697_0[1]),.dinb(w_n632_0[1]),.dout(n698),.clk(gclk));
	jxor g0635(.dina(w_n698_0[1]),.dinb(w_n630_0[1]),.dout(n699),.clk(gclk));
	jxor g0636(.dina(w_n699_0[1]),.dinb(w_n627_0[1]),.dout(n700),.clk(gclk));
	jnot g0637(.din(w_n700_0[1]),.dout(n701),.clk(gclk));
	jxor g0638(.dina(w_n701_0[1]),.dinb(w_n625_0[2]),.dout(n702),.clk(gclk));
	jxor g0639(.dina(n702),.dinb(w_dff_B_XbI8uxyG4_1),.dout(n703),.clk(gclk));
	jxor g0640(.dina(w_n703_0[1]),.dinb(w_n619_0[1]),.dout(n704),.clk(gclk));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_dff_B_55BBytC33_1),.dout(w_dff_A_rUJAEsv64_2),.clk(gclk));
	jand g0642(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n706),.clk(gclk));
	jnot g0643(.din(w_n706_0[1]),.dout(n707),.clk(gclk));
	jnot g0644(.din(w_n703_0[0]),.dout(n708),.clk(gclk));
	jor g0645(.dina(n708),.dinb(w_n619_0[0]),.dout(n709),.clk(gclk));
	jor g0646(.dina(w_n704_0[0]),.dinb(w_n614_0[0]),.dout(n710),.clk(gclk));
	jand g0647(.dina(n710),.dinb(w_dff_B_IwWgFsJp8_1),.dout(n711),.clk(gclk));
	jand g0648(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n712),.clk(gclk));
	jnot g0649(.din(w_n712_0[1]),.dout(n713),.clk(gclk));
	jor g0650(.dina(w_n701_0[0]),.dinb(w_n625_0[1]),.dout(n714),.clk(gclk));
	jxor g0651(.dina(w_n700_0[0]),.dinb(w_n625_0[0]),.dout(n715),.clk(gclk));
	jor g0652(.dina(n715),.dinb(w_n620_0[0]),.dout(n716),.clk(gclk));
	jand g0653(.dina(n716),.dinb(w_dff_B_TcMWfGUl2_1),.dout(n717),.clk(gclk));
	jand g0654(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n718),.clk(gclk));
	jnot g0655(.din(n718),.dout(n719),.clk(gclk));
	jand g0656(.dina(w_n698_0[0]),.dinb(w_n630_0[0]),.dout(n720),.clk(gclk));
	jand g0657(.dina(w_n699_0[0]),.dinb(w_n627_0[0]),.dout(n721),.clk(gclk));
	jor g0658(.dina(n721),.dinb(w_dff_B_Dlogfoix6_1),.dout(n722),.clk(gclk));
	jand g0659(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n723),.clk(gclk));
	jnot g0660(.din(n723),.dout(n724),.clk(gclk));
	jand g0661(.dina(w_n696_0[0]),.dinb(w_n635_0[0]),.dout(n725),.clk(gclk));
	jand g0662(.dina(w_n697_0[0]),.dinb(w_n632_0[0]),.dout(n726),.clk(gclk));
	jor g0663(.dina(n726),.dinb(w_dff_B_bl7gv11g3_1),.dout(n727),.clk(gclk));
	jand g0664(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n728),.clk(gclk));
	jnot g0665(.din(n728),.dout(n729),.clk(gclk));
	jand g0666(.dina(w_n694_0[0]),.dinb(w_n640_0[0]),.dout(n730),.clk(gclk));
	jand g0667(.dina(w_n695_0[0]),.dinb(w_n637_0[0]),.dout(n731),.clk(gclk));
	jor g0668(.dina(n731),.dinb(w_dff_B_FXe6CwUR4_1),.dout(n732),.clk(gclk));
	jand g0669(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n733),.clk(gclk));
	jnot g0670(.din(n733),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_n692_0[0]),.dinb(w_n645_0[0]),.dout(n735),.clk(gclk));
	jand g0672(.dina(w_n693_0[0]),.dinb(w_n642_0[0]),.dout(n736),.clk(gclk));
	jor g0673(.dina(n736),.dinb(w_dff_B_dKuj7UIM9_1),.dout(n737),.clk(gclk));
	jand g0674(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n738),.clk(gclk));
	jnot g0675(.din(n738),.dout(n739),.clk(gclk));
	jand g0676(.dina(w_n690_0[0]),.dinb(w_n650_0[0]),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_n691_0[0]),.dinb(w_n647_0[0]),.dout(n741),.clk(gclk));
	jor g0678(.dina(n741),.dinb(w_dff_B_hEuuqHdi4_1),.dout(n742),.clk(gclk));
	jand g0679(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n743),.clk(gclk));
	jnot g0680(.din(n743),.dout(n744),.clk(gclk));
	jand g0681(.dina(w_n688_0[0]),.dinb(w_n655_0[0]),.dout(n745),.clk(gclk));
	jand g0682(.dina(w_n689_0[0]),.dinb(w_n652_0[0]),.dout(n746),.clk(gclk));
	jor g0683(.dina(n746),.dinb(w_dff_B_cxqTMeGw6_1),.dout(n747),.clk(gclk));
	jand g0684(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n748),.clk(gclk));
	jnot g0685(.din(n748),.dout(n749),.clk(gclk));
	jand g0686(.dina(w_n686_0[0]),.dinb(w_n660_0[0]),.dout(n750),.clk(gclk));
	jand g0687(.dina(w_n687_0[0]),.dinb(w_n657_0[0]),.dout(n751),.clk(gclk));
	jor g0688(.dina(n751),.dinb(w_dff_B_TyaiXiWX8_1),.dout(n752),.clk(gclk));
	jand g0689(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n753),.clk(gclk));
	jnot g0690(.din(n753),.dout(n754),.clk(gclk));
	jand g0691(.dina(w_n684_0[0]),.dinb(w_n665_0[0]),.dout(n755),.clk(gclk));
	jand g0692(.dina(w_n685_0[0]),.dinb(w_n662_0[0]),.dout(n756),.clk(gclk));
	jor g0693(.dina(n756),.dinb(w_dff_B_QHE2z7Ie5_1),.dout(n757),.clk(gclk));
	jand g0694(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n758),.clk(gclk));
	jnot g0695(.din(n758),.dout(n759),.clk(gclk));
	jand g0696(.dina(w_n682_0[0]),.dinb(w_n672_0[0]),.dout(n760),.clk(gclk));
	jand g0697(.dina(w_n683_0[0]),.dinb(w_n667_0[0]),.dout(n761),.clk(gclk));
	jor g0698(.dina(n761),.dinb(w_dff_B_vcmnjSc07_1),.dout(n762),.clk(gclk));
	jand g0699(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n763),.clk(gclk));
	jnot g0700(.din(n763),.dout(n764),.clk(gclk));
	jor g0701(.dina(w_n680_0[0]),.dinb(w_n586_0[0]),.dout(n765),.clk(gclk));
	jand g0702(.dina(w_n681_0[0]),.dinb(w_n674_0[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(n767),.dinb(w_dff_B_728XF6378_1),.dout(n768),.clk(gclk));
	jnot g0705(.din(n768),.dout(n769),.clk(gclk));
	jand g0706(.dina(w_G307gat_3[1]),.dinb(w_G205gat_6[2]),.dout(n770),.clk(gclk));
	jnot g0707(.din(n770),.dout(n771),.clk(gclk));
	jand g0708(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n772_0[1]),.dinb(w_n678_0[0]),.dout(n773),.clk(gclk));
	jnot g0710(.din(w_n773_0[1]),.dout(n774),.clk(gclk));
	jand g0711(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n775),.clk(gclk));
	jor g0712(.dina(w_n775_0[1]),.dinb(w_n675_0[0]),.dout(n776),.clk(gclk));
	jand g0713(.dina(w_dff_B_scAyxHrg4_0),.dinb(w_n774_0[1]),.dout(n777),.clk(gclk));
	jxor g0714(.dina(w_n777_0[1]),.dinb(w_n676_0[1]),.dout(n778),.clk(gclk));
	jxor g0715(.dina(w_n778_0[1]),.dinb(w_n771_0[1]),.dout(n779),.clk(gclk));
	jxor g0716(.dina(w_n779_0[1]),.dinb(w_n769_0[1]),.dout(n780),.clk(gclk));
	jxor g0717(.dina(w_n780_0[1]),.dinb(w_n764_0[1]),.dout(n781),.clk(gclk));
	jxor g0718(.dina(w_n781_0[1]),.dinb(w_n762_0[1]),.dout(n782),.clk(gclk));
	jxor g0719(.dina(w_n782_0[1]),.dinb(w_n759_0[1]),.dout(n783),.clk(gclk));
	jxor g0720(.dina(w_n783_0[1]),.dinb(w_n757_0[1]),.dout(n784),.clk(gclk));
	jxor g0721(.dina(w_n784_0[1]),.dinb(w_n754_0[1]),.dout(n785),.clk(gclk));
	jxor g0722(.dina(w_n785_0[1]),.dinb(w_n752_0[1]),.dout(n786),.clk(gclk));
	jxor g0723(.dina(w_n786_0[1]),.dinb(w_n749_0[1]),.dout(n787),.clk(gclk));
	jxor g0724(.dina(w_n787_0[1]),.dinb(w_n747_0[1]),.dout(n788),.clk(gclk));
	jxor g0725(.dina(w_n788_0[1]),.dinb(w_n744_0[1]),.dout(n789),.clk(gclk));
	jxor g0726(.dina(w_n789_0[1]),.dinb(w_n742_0[1]),.dout(n790),.clk(gclk));
	jxor g0727(.dina(w_n790_0[1]),.dinb(w_n739_0[1]),.dout(n791),.clk(gclk));
	jxor g0728(.dina(w_n791_0[1]),.dinb(w_n737_0[1]),.dout(n792),.clk(gclk));
	jxor g0729(.dina(w_n792_0[1]),.dinb(w_n734_0[1]),.dout(n793),.clk(gclk));
	jxor g0730(.dina(w_n793_0[1]),.dinb(w_n732_0[1]),.dout(n794),.clk(gclk));
	jxor g0731(.dina(w_n794_0[1]),.dinb(w_n729_0[1]),.dout(n795),.clk(gclk));
	jxor g0732(.dina(w_n795_0[1]),.dinb(w_n727_0[1]),.dout(n796),.clk(gclk));
	jxor g0733(.dina(w_n796_0[1]),.dinb(w_n724_0[1]),.dout(n797),.clk(gclk));
	jxor g0734(.dina(w_n797_0[1]),.dinb(w_n722_0[1]),.dout(n798),.clk(gclk));
	jxor g0735(.dina(w_n798_0[1]),.dinb(w_n719_0[1]),.dout(n799),.clk(gclk));
	jnot g0736(.din(w_n799_0[1]),.dout(n800),.clk(gclk));
	jxor g0737(.dina(w_n800_0[1]),.dinb(w_n717_0[2]),.dout(n801),.clk(gclk));
	jxor g0738(.dina(n801),.dinb(w_dff_B_Z79BEmHT1_1),.dout(n802),.clk(gclk));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n711_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_dff_B_9PkQ9nLG0_1),.dout(w_dff_A_84xyMY4Y3_2),.clk(gclk));
	jand g0741(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n805),.clk(gclk));
	jnot g0742(.din(w_n805_0[1]),.dout(n806),.clk(gclk));
	jnot g0743(.din(w_n802_0[0]),.dout(n807),.clk(gclk));
	jor g0744(.dina(n807),.dinb(w_n711_0[0]),.dout(n808),.clk(gclk));
	jor g0745(.dina(w_n803_0[0]),.dinb(w_n706_0[0]),.dout(n809),.clk(gclk));
	jand g0746(.dina(n809),.dinb(w_dff_B_q0XPWQFi0_1),.dout(n810),.clk(gclk));
	jand g0747(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n811),.clk(gclk));
	jor g0748(.dina(w_n800_0[0]),.dinb(w_n717_0[1]),.dout(n812),.clk(gclk));
	jxor g0749(.dina(w_n799_0[0]),.dinb(w_n717_0[0]),.dout(n813),.clk(gclk));
	jor g0750(.dina(n813),.dinb(w_n712_0[0]),.dout(n814),.clk(gclk));
	jand g0751(.dina(n814),.dinb(w_dff_B_e90BrRBC1_1),.dout(n815),.clk(gclk));
	jand g0752(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n816),.clk(gclk));
	jnot g0753(.din(w_n816_0[1]),.dout(n817),.clk(gclk));
	jand g0754(.dina(w_n797_0[0]),.dinb(w_n722_0[0]),.dout(n818),.clk(gclk));
	jand g0755(.dina(w_n798_0[0]),.dinb(w_n719_0[0]),.dout(n819),.clk(gclk));
	jor g0756(.dina(n819),.dinb(w_dff_B_dNQi9PLH0_1),.dout(n820),.clk(gclk));
	jand g0757(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n821),.clk(gclk));
	jnot g0758(.din(n821),.dout(n822),.clk(gclk));
	jand g0759(.dina(w_n795_0[0]),.dinb(w_n727_0[0]),.dout(n823),.clk(gclk));
	jand g0760(.dina(w_n796_0[0]),.dinb(w_n724_0[0]),.dout(n824),.clk(gclk));
	jor g0761(.dina(n824),.dinb(w_dff_B_BysUlr9y6_1),.dout(n825),.clk(gclk));
	jand g0762(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n826),.clk(gclk));
	jnot g0763(.din(n826),.dout(n827),.clk(gclk));
	jand g0764(.dina(w_n793_0[0]),.dinb(w_n732_0[0]),.dout(n828),.clk(gclk));
	jand g0765(.dina(w_n794_0[0]),.dinb(w_n729_0[0]),.dout(n829),.clk(gclk));
	jor g0766(.dina(n829),.dinb(w_dff_B_BEvijuvY2_1),.dout(n830),.clk(gclk));
	jand g0767(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n831),.clk(gclk));
	jnot g0768(.din(n831),.dout(n832),.clk(gclk));
	jand g0769(.dina(w_n791_0[0]),.dinb(w_n737_0[0]),.dout(n833),.clk(gclk));
	jand g0770(.dina(w_n792_0[0]),.dinb(w_n734_0[0]),.dout(n834),.clk(gclk));
	jor g0771(.dina(n834),.dinb(w_dff_B_aKoY2FFS5_1),.dout(n835),.clk(gclk));
	jand g0772(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n836),.clk(gclk));
	jnot g0773(.din(n836),.dout(n837),.clk(gclk));
	jand g0774(.dina(w_n789_0[0]),.dinb(w_n742_0[0]),.dout(n838),.clk(gclk));
	jand g0775(.dina(w_n790_0[0]),.dinb(w_n739_0[0]),.dout(n839),.clk(gclk));
	jor g0776(.dina(n839),.dinb(w_dff_B_80NBw8E22_1),.dout(n840),.clk(gclk));
	jand g0777(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n841),.clk(gclk));
	jnot g0778(.din(n841),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n787_0[0]),.dinb(w_n747_0[0]),.dout(n843),.clk(gclk));
	jand g0780(.dina(w_n788_0[0]),.dinb(w_n744_0[0]),.dout(n844),.clk(gclk));
	jor g0781(.dina(n844),.dinb(w_dff_B_i5rvOa3p3_1),.dout(n845),.clk(gclk));
	jand g0782(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n846),.clk(gclk));
	jnot g0783(.din(n846),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n785_0[0]),.dinb(w_n752_0[0]),.dout(n848),.clk(gclk));
	jand g0785(.dina(w_n786_0[0]),.dinb(w_n749_0[0]),.dout(n849),.clk(gclk));
	jor g0786(.dina(n849),.dinb(w_dff_B_GuYSHLCf0_1),.dout(n850),.clk(gclk));
	jand g0787(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n851),.clk(gclk));
	jnot g0788(.din(n851),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n783_0[0]),.dinb(w_n757_0[0]),.dout(n853),.clk(gclk));
	jand g0790(.dina(w_n784_0[0]),.dinb(w_n754_0[0]),.dout(n854),.clk(gclk));
	jor g0791(.dina(n854),.dinb(w_dff_B_pky1lf7R0_1),.dout(n855),.clk(gclk));
	jand g0792(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n856),.clk(gclk));
	jnot g0793(.din(n856),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n781_0[0]),.dinb(w_n762_0[0]),.dout(n858),.clk(gclk));
	jand g0795(.dina(w_n782_0[0]),.dinb(w_n759_0[0]),.dout(n859),.clk(gclk));
	jor g0796(.dina(n859),.dinb(w_dff_B_rEp1xRQD0_1),.dout(n860),.clk(gclk));
	jand g0797(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n861),.clk(gclk));
	jnot g0798(.din(n861),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n779_0[0]),.dinb(w_n769_0[0]),.dout(n863),.clk(gclk));
	jand g0800(.dina(w_n780_0[0]),.dinb(w_n764_0[0]),.dout(n864),.clk(gclk));
	jor g0801(.dina(n864),.dinb(w_dff_B_DhUnkwK37_1),.dout(n865),.clk(gclk));
	jand g0802(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n866),.clk(gclk));
	jnot g0803(.din(n866),.dout(n867),.clk(gclk));
	jor g0804(.dina(w_n777_0[0]),.dinb(w_n676_0[0]),.dout(n868),.clk(gclk));
	jand g0805(.dina(w_n778_0[0]),.dinb(w_n771_0[0]),.dout(n869),.clk(gclk));
	jnot g0806(.din(n869),.dout(n870),.clk(gclk));
	jand g0807(.dina(n870),.dinb(w_dff_B_Rx5fQxCb1_1),.dout(n871),.clk(gclk));
	jnot g0808(.din(n871),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_G307gat_3[0]),.dinb(w_G222gat_6[2]),.dout(n873),.clk(gclk));
	jnot g0810(.din(n873),.dout(n874),.clk(gclk));
	jand g0811(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n875),.clk(gclk));
	jxor g0812(.dina(w_n875_0[1]),.dinb(w_n772_0[0]),.dout(n876),.clk(gclk));
	jor g0813(.dina(n876),.dinb(w_n773_0[0]),.dout(n877),.clk(gclk));
	jor g0814(.dina(w_n875_0[0]),.dinb(w_n774_0[0]),.dout(n878),.clk(gclk));
	jand g0815(.dina(n878),.dinb(w_n877_0[1]),.dout(n879),.clk(gclk));
	jxor g0816(.dina(w_n879_0[1]),.dinb(w_n874_0[1]),.dout(n880),.clk(gclk));
	jxor g0817(.dina(w_n880_0[1]),.dinb(w_n872_0[1]),.dout(n881),.clk(gclk));
	jxor g0818(.dina(w_n881_0[1]),.dinb(w_n867_0[1]),.dout(n882),.clk(gclk));
	jxor g0819(.dina(w_n882_0[1]),.dinb(w_n865_0[1]),.dout(n883),.clk(gclk));
	jxor g0820(.dina(w_n883_0[1]),.dinb(w_n862_0[1]),.dout(n884),.clk(gclk));
	jxor g0821(.dina(w_n884_0[1]),.dinb(w_n860_0[1]),.dout(n885),.clk(gclk));
	jxor g0822(.dina(w_n885_0[1]),.dinb(w_n857_0[1]),.dout(n886),.clk(gclk));
	jxor g0823(.dina(w_n886_0[1]),.dinb(w_n855_0[1]),.dout(n887),.clk(gclk));
	jxor g0824(.dina(w_n887_0[1]),.dinb(w_n852_0[1]),.dout(n888),.clk(gclk));
	jxor g0825(.dina(w_n888_0[1]),.dinb(w_n850_0[1]),.dout(n889),.clk(gclk));
	jxor g0826(.dina(w_n889_0[1]),.dinb(w_n847_0[1]),.dout(n890),.clk(gclk));
	jxor g0827(.dina(w_n890_0[1]),.dinb(w_n845_0[1]),.dout(n891),.clk(gclk));
	jxor g0828(.dina(w_n891_0[1]),.dinb(w_n842_0[1]),.dout(n892),.clk(gclk));
	jxor g0829(.dina(w_n892_0[1]),.dinb(w_n840_0[1]),.dout(n893),.clk(gclk));
	jxor g0830(.dina(w_n893_0[1]),.dinb(w_n837_0[1]),.dout(n894),.clk(gclk));
	jxor g0831(.dina(w_n894_0[1]),.dinb(w_n835_0[1]),.dout(n895),.clk(gclk));
	jxor g0832(.dina(w_n895_0[1]),.dinb(w_n832_0[1]),.dout(n896),.clk(gclk));
	jxor g0833(.dina(w_n896_0[1]),.dinb(w_n830_0[1]),.dout(n897),.clk(gclk));
	jxor g0834(.dina(w_n897_0[1]),.dinb(w_n827_0[1]),.dout(n898),.clk(gclk));
	jxor g0835(.dina(w_n898_0[1]),.dinb(w_n825_0[1]),.dout(n899),.clk(gclk));
	jxor g0836(.dina(w_n899_0[1]),.dinb(w_n822_0[1]),.dout(n900),.clk(gclk));
	jxor g0837(.dina(w_n900_0[2]),.dinb(w_n820_0[2]),.dout(n901),.clk(gclk));
	jxor g0838(.dina(n901),.dinb(w_dff_B_IauIUggA0_1),.dout(n902),.clk(gclk));
	jxor g0839(.dina(w_n902_0[1]),.dinb(w_n815_0[1]),.dout(n903),.clk(gclk));
	jxor g0840(.dina(w_n903_0[1]),.dinb(w_n811_0[1]),.dout(n904),.clk(gclk));
	jxor g0841(.dina(w_n904_0[1]),.dinb(w_n810_0[1]),.dout(n905),.clk(gclk));
	jxor g0842(.dina(w_n905_0[1]),.dinb(w_dff_B_mW8Cwltp4_1),.dout(w_dff_A_1raJBPiI7_2),.clk(gclk));
	jnot g0843(.din(w_n904_0[0]),.dout(n907),.clk(gclk));
	jor g0844(.dina(n907),.dinb(w_n810_0[0]),.dout(n908),.clk(gclk));
	jor g0845(.dina(w_n905_0[0]),.dinb(w_n805_0[0]),.dout(n909),.clk(gclk));
	jand g0846(.dina(n909),.dinb(w_dff_B_kLvZqWp66_1),.dout(n910),.clk(gclk));
	jand g0847(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n911),.clk(gclk));
	jnot g0848(.din(w_n902_0[0]),.dout(n912),.clk(gclk));
	jor g0849(.dina(n912),.dinb(w_n815_0[0]),.dout(n913),.clk(gclk));
	jor g0850(.dina(w_n903_0[0]),.dinb(w_n811_0[0]),.dout(n914),.clk(gclk));
	jand g0851(.dina(n914),.dinb(w_dff_B_7ZqNEE1X2_1),.dout(n915),.clk(gclk));
	jand g0852(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n916),.clk(gclk));
	jand g0853(.dina(w_n900_0[1]),.dinb(w_n820_0[1]),.dout(n917),.clk(gclk));
	jnot g0854(.din(n917),.dout(n918),.clk(gclk));
	jnot g0855(.din(w_n900_0[0]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(n919),.dinb(w_n820_0[0]),.dout(n920),.clk(gclk));
	jor g0857(.dina(n920),.dinb(w_n816_0[0]),.dout(n921),.clk(gclk));
	jand g0858(.dina(n921),.dinb(n918),.dout(n922),.clk(gclk));
	jand g0859(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n923),.clk(gclk));
	jnot g0860(.din(n923),.dout(n924),.clk(gclk));
	jand g0861(.dina(w_n898_0[0]),.dinb(w_n825_0[0]),.dout(n925),.clk(gclk));
	jand g0862(.dina(w_n899_0[0]),.dinb(w_n822_0[0]),.dout(n926),.clk(gclk));
	jor g0863(.dina(n926),.dinb(w_dff_B_tWfpopR90_1),.dout(n927),.clk(gclk));
	jand g0864(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n928),.clk(gclk));
	jnot g0865(.din(n928),.dout(n929),.clk(gclk));
	jand g0866(.dina(w_n896_0[0]),.dinb(w_n830_0[0]),.dout(n930),.clk(gclk));
	jand g0867(.dina(w_n897_0[0]),.dinb(w_n827_0[0]),.dout(n931),.clk(gclk));
	jor g0868(.dina(n931),.dinb(w_dff_B_ES8A9qFY2_1),.dout(n932),.clk(gclk));
	jand g0869(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n933),.clk(gclk));
	jnot g0870(.din(n933),.dout(n934),.clk(gclk));
	jand g0871(.dina(w_n894_0[0]),.dinb(w_n835_0[0]),.dout(n935),.clk(gclk));
	jand g0872(.dina(w_n895_0[0]),.dinb(w_n832_0[0]),.dout(n936),.clk(gclk));
	jor g0873(.dina(n936),.dinb(w_dff_B_QJ7JBseb2_1),.dout(n937),.clk(gclk));
	jand g0874(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n938),.clk(gclk));
	jnot g0875(.din(n938),.dout(n939),.clk(gclk));
	jand g0876(.dina(w_n892_0[0]),.dinb(w_n840_0[0]),.dout(n940),.clk(gclk));
	jand g0877(.dina(w_n893_0[0]),.dinb(w_n837_0[0]),.dout(n941),.clk(gclk));
	jor g0878(.dina(n941),.dinb(w_dff_B_euu1EETl5_1),.dout(n942),.clk(gclk));
	jand g0879(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n943),.clk(gclk));
	jnot g0880(.din(n943),.dout(n944),.clk(gclk));
	jand g0881(.dina(w_n890_0[0]),.dinb(w_n845_0[0]),.dout(n945),.clk(gclk));
	jand g0882(.dina(w_n891_0[0]),.dinb(w_n842_0[0]),.dout(n946),.clk(gclk));
	jor g0883(.dina(n946),.dinb(w_dff_B_6kM8FJQY9_1),.dout(n947),.clk(gclk));
	jand g0884(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n948),.clk(gclk));
	jnot g0885(.din(n948),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_n888_0[0]),.dinb(w_n850_0[0]),.dout(n950),.clk(gclk));
	jand g0887(.dina(w_n889_0[0]),.dinb(w_n847_0[0]),.dout(n951),.clk(gclk));
	jor g0888(.dina(n951),.dinb(w_dff_B_8U4bRvfp3_1),.dout(n952),.clk(gclk));
	jand g0889(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n953),.clk(gclk));
	jnot g0890(.din(n953),.dout(n954),.clk(gclk));
	jand g0891(.dina(w_n886_0[0]),.dinb(w_n855_0[0]),.dout(n955),.clk(gclk));
	jand g0892(.dina(w_n887_0[0]),.dinb(w_n852_0[0]),.dout(n956),.clk(gclk));
	jor g0893(.dina(n956),.dinb(w_dff_B_RYkSGtmM3_1),.dout(n957),.clk(gclk));
	jand g0894(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n958),.clk(gclk));
	jnot g0895(.din(n958),.dout(n959),.clk(gclk));
	jand g0896(.dina(w_n884_0[0]),.dinb(w_n860_0[0]),.dout(n960),.clk(gclk));
	jand g0897(.dina(w_n885_0[0]),.dinb(w_n857_0[0]),.dout(n961),.clk(gclk));
	jor g0898(.dina(n961),.dinb(w_dff_B_hXdk3x3M0_1),.dout(n962),.clk(gclk));
	jand g0899(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n963),.clk(gclk));
	jnot g0900(.din(n963),.dout(n964),.clk(gclk));
	jand g0901(.dina(w_n882_0[0]),.dinb(w_n865_0[0]),.dout(n965),.clk(gclk));
	jand g0902(.dina(w_n883_0[0]),.dinb(w_n862_0[0]),.dout(n966),.clk(gclk));
	jor g0903(.dina(n966),.dinb(w_dff_B_9T1eoiix9_1),.dout(n967),.clk(gclk));
	jand g0904(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n968),.clk(gclk));
	jnot g0905(.din(n968),.dout(n969),.clk(gclk));
	jand g0906(.dina(w_n880_0[0]),.dinb(w_n872_0[0]),.dout(n970),.clk(gclk));
	jand g0907(.dina(w_n881_0[0]),.dinb(w_n867_0[0]),.dout(n971),.clk(gclk));
	jor g0908(.dina(n971),.dinb(w_dff_B_XDYSzb834_1),.dout(n972),.clk(gclk));
	jand g0909(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n973),.clk(gclk));
	jnot g0910(.din(n973),.dout(n974),.clk(gclk));
	jand g0911(.dina(w_n879_0[0]),.dinb(w_n874_0[0]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(n976),.dinb(w_n877_0[0]),.dout(n977),.clk(gclk));
	jnot g0914(.din(n977),.dout(n978),.clk(gclk));
	jnot g0915(.din(w_n775_0[0]),.dout(n979),.clk(gclk));
	jand g0916(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n980),.clk(gclk));
	jand g0917(.dina(w_n980_0[1]),.dinb(n979),.dout(n981),.clk(gclk));
	jnot g0918(.din(n981),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_G307gat_2[2]),.dinb(w_G239gat_6[2]),.dout(n983),.clk(gclk));
	jxor g0920(.dina(w_n983_0[1]),.dinb(w_n982_0[1]),.dout(n984),.clk(gclk));
	jxor g0921(.dina(w_n984_0[1]),.dinb(w_n978_0[1]),.dout(n985),.clk(gclk));
	jxor g0922(.dina(w_n985_0[1]),.dinb(w_n974_0[1]),.dout(n986),.clk(gclk));
	jxor g0923(.dina(w_n986_0[1]),.dinb(w_n972_0[1]),.dout(n987),.clk(gclk));
	jxor g0924(.dina(w_n987_0[1]),.dinb(w_n969_0[1]),.dout(n988),.clk(gclk));
	jxor g0925(.dina(w_n988_0[1]),.dinb(w_n967_0[1]),.dout(n989),.clk(gclk));
	jxor g0926(.dina(w_n989_0[1]),.dinb(w_n964_0[1]),.dout(n990),.clk(gclk));
	jxor g0927(.dina(w_n990_0[1]),.dinb(w_n962_0[1]),.dout(n991),.clk(gclk));
	jxor g0928(.dina(w_n991_0[1]),.dinb(w_n959_0[1]),.dout(n992),.clk(gclk));
	jxor g0929(.dina(w_n992_0[1]),.dinb(w_n957_0[1]),.dout(n993),.clk(gclk));
	jxor g0930(.dina(w_n993_0[1]),.dinb(w_n954_0[1]),.dout(n994),.clk(gclk));
	jxor g0931(.dina(w_n994_0[1]),.dinb(w_n952_0[1]),.dout(n995),.clk(gclk));
	jxor g0932(.dina(w_n995_0[1]),.dinb(w_n949_0[1]),.dout(n996),.clk(gclk));
	jxor g0933(.dina(w_n996_0[1]),.dinb(w_n947_0[1]),.dout(n997),.clk(gclk));
	jxor g0934(.dina(w_n997_0[1]),.dinb(w_n944_0[1]),.dout(n998),.clk(gclk));
	jxor g0935(.dina(w_n998_0[1]),.dinb(w_n942_0[1]),.dout(n999),.clk(gclk));
	jxor g0936(.dina(w_n999_0[1]),.dinb(w_n939_0[1]),.dout(n1000),.clk(gclk));
	jxor g0937(.dina(w_n1000_0[1]),.dinb(w_n937_0[1]),.dout(n1001),.clk(gclk));
	jxor g0938(.dina(w_n1001_0[1]),.dinb(w_n934_0[1]),.dout(n1002),.clk(gclk));
	jxor g0939(.dina(w_n1002_0[1]),.dinb(w_n932_0[1]),.dout(n1003),.clk(gclk));
	jxor g0940(.dina(w_n1003_0[1]),.dinb(w_n929_0[1]),.dout(n1004),.clk(gclk));
	jxor g0941(.dina(w_n1004_0[1]),.dinb(w_n927_0[1]),.dout(n1005),.clk(gclk));
	jxor g0942(.dina(w_n1005_0[1]),.dinb(w_n924_0[1]),.dout(n1006),.clk(gclk));
	jxor g0943(.dina(w_n1006_0[1]),.dinb(w_n922_0[1]),.dout(n1007),.clk(gclk));
	jxor g0944(.dina(w_n1007_0[1]),.dinb(w_n916_0[1]),.dout(n1008),.clk(gclk));
	jnot g0945(.din(w_n1008_0[1]),.dout(n1009),.clk(gclk));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n915_0[2]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(n1010),.dinb(w_n911_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n910_0[1]),.dout(w_dff_A_y2Cx0Ugv4_2),.clk(gclk));
	jand g0949(.dina(w_n1011_0[0]),.dinb(w_n910_0[0]),.dout(n1013),.clk(gclk));
	jor g0950(.dina(w_n1009_0[0]),.dinb(w_n915_0[1]),.dout(n1014),.clk(gclk));
	jxor g0951(.dina(w_n1008_0[0]),.dinb(w_n915_0[0]),.dout(n1015),.clk(gclk));
	jor g0952(.dina(n1015),.dinb(w_n911_0[0]),.dout(n1016),.clk(gclk));
	jand g0953(.dina(n1016),.dinb(w_dff_B_kUX2dQoU1_1),.dout(n1017),.clk(gclk));
	jand g0954(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1018),.clk(gclk));
	jnot g0955(.din(w_n1006_0[0]),.dout(n1019),.clk(gclk));
	jor g0956(.dina(n1019),.dinb(w_n922_0[0]),.dout(n1020),.clk(gclk));
	jor g0957(.dina(w_n1007_0[0]),.dinb(w_n916_0[0]),.dout(n1021),.clk(gclk));
	jand g0958(.dina(n1021),.dinb(w_dff_B_L4bM11W03_1),.dout(n1022),.clk(gclk));
	jand g0959(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1023),.clk(gclk));
	jand g0960(.dina(w_n1004_0[0]),.dinb(w_n927_0[0]),.dout(n1024),.clk(gclk));
	jand g0961(.dina(w_n1005_0[0]),.dinb(w_n924_0[0]),.dout(n1025),.clk(gclk));
	jor g0962(.dina(n1025),.dinb(w_dff_B_JZOAAh0m7_1),.dout(n1026),.clk(gclk));
	jand g0963(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1027),.clk(gclk));
	jnot g0964(.din(n1027),.dout(n1028),.clk(gclk));
	jand g0965(.dina(w_n1002_0[0]),.dinb(w_n932_0[0]),.dout(n1029),.clk(gclk));
	jand g0966(.dina(w_n1003_0[0]),.dinb(w_n929_0[0]),.dout(n1030),.clk(gclk));
	jor g0967(.dina(n1030),.dinb(w_dff_B_tM9aG5Ne4_1),.dout(n1031),.clk(gclk));
	jand g0968(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1032),.clk(gclk));
	jnot g0969(.din(n1032),.dout(n1033),.clk(gclk));
	jand g0970(.dina(w_n1000_0[0]),.dinb(w_n937_0[0]),.dout(n1034),.clk(gclk));
	jand g0971(.dina(w_n1001_0[0]),.dinb(w_n934_0[0]),.dout(n1035),.clk(gclk));
	jor g0972(.dina(n1035),.dinb(w_dff_B_RhSaeNsr6_1),.dout(n1036),.clk(gclk));
	jand g0973(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1037),.clk(gclk));
	jnot g0974(.din(n1037),.dout(n1038),.clk(gclk));
	jand g0975(.dina(w_n998_0[0]),.dinb(w_n942_0[0]),.dout(n1039),.clk(gclk));
	jand g0976(.dina(w_n999_0[0]),.dinb(w_n939_0[0]),.dout(n1040),.clk(gclk));
	jor g0977(.dina(n1040),.dinb(w_dff_B_CB0sktN81_1),.dout(n1041),.clk(gclk));
	jand g0978(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1042),.clk(gclk));
	jnot g0979(.din(n1042),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_n996_0[0]),.dinb(w_n947_0[0]),.dout(n1044),.clk(gclk));
	jand g0981(.dina(w_n997_0[0]),.dinb(w_n944_0[0]),.dout(n1045),.clk(gclk));
	jor g0982(.dina(n1045),.dinb(w_dff_B_sCOjvpwk7_1),.dout(n1046),.clk(gclk));
	jand g0983(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1047),.clk(gclk));
	jnot g0984(.din(n1047),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_n994_0[0]),.dinb(w_n952_0[0]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n995_0[0]),.dinb(w_n949_0[0]),.dout(n1050),.clk(gclk));
	jor g0987(.dina(n1050),.dinb(w_dff_B_Fm64XX5H4_1),.dout(n1051),.clk(gclk));
	jand g0988(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1052),.clk(gclk));
	jnot g0989(.din(n1052),.dout(n1053),.clk(gclk));
	jand g0990(.dina(w_n992_0[0]),.dinb(w_n957_0[0]),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n993_0[0]),.dinb(w_n954_0[0]),.dout(n1055),.clk(gclk));
	jor g0992(.dina(n1055),.dinb(w_dff_B_LAVnKpcM7_1),.dout(n1056),.clk(gclk));
	jand g0993(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1057),.clk(gclk));
	jnot g0994(.din(n1057),.dout(n1058),.clk(gclk));
	jand g0995(.dina(w_n990_0[0]),.dinb(w_n962_0[0]),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n991_0[0]),.dinb(w_n959_0[0]),.dout(n1060),.clk(gclk));
	jor g0997(.dina(n1060),.dinb(w_dff_B_V7jV1Ext4_1),.dout(n1061),.clk(gclk));
	jand g0998(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1062),.clk(gclk));
	jnot g0999(.din(n1062),.dout(n1063),.clk(gclk));
	jand g1000(.dina(w_n988_0[0]),.dinb(w_n967_0[0]),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n989_0[0]),.dinb(w_n964_0[0]),.dout(n1065),.clk(gclk));
	jor g1002(.dina(n1065),.dinb(w_dff_B_KfPZcrTp9_1),.dout(n1066),.clk(gclk));
	jand g1003(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1067),.clk(gclk));
	jnot g1004(.din(n1067),.dout(n1068),.clk(gclk));
	jand g1005(.dina(w_n986_0[0]),.dinb(w_n972_0[0]),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n987_0[0]),.dinb(w_n969_0[0]),.dout(n1070),.clk(gclk));
	jor g1007(.dina(n1070),.dinb(w_dff_B_JEKq79lb7_1),.dout(n1071),.clk(gclk));
	jand g1008(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1072),.clk(gclk));
	jnot g1009(.din(n1072),.dout(n1073),.clk(gclk));
	jand g1010(.dina(w_n984_0[0]),.dinb(w_n978_0[0]),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n985_0[0]),.dinb(w_n974_0[0]),.dout(n1075),.clk(gclk));
	jor g1012(.dina(n1075),.dinb(w_dff_B_vjml4cqS8_1),.dout(n1076),.clk(gclk));
	jand g1013(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1077),.clk(gclk));
	jand g1014(.dina(w_G307gat_2[1]),.dinb(w_G256gat_6[2]),.dout(n1078),.clk(gclk));
	jor g1015(.dina(w_n983_0[0]),.dinb(w_n982_0[0]),.dout(n1079),.clk(gclk));
	jand g1016(.dina(n1079),.dinb(w_n980_0[0]),.dout(n1080),.clk(gclk));
	jxor g1017(.dina(w_n1080_0[1]),.dinb(w_n1078_0[1]),.dout(n1081),.clk(gclk));
	jnot g1018(.din(n1081),.dout(n1082),.clk(gclk));
	jxor g1019(.dina(w_n1082_0[1]),.dinb(w_n1077_0[1]),.dout(n1083),.clk(gclk));
	jxor g1020(.dina(w_n1083_0[1]),.dinb(w_n1076_0[1]),.dout(n1084),.clk(gclk));
	jxor g1021(.dina(w_n1084_0[1]),.dinb(w_n1073_0[1]),.dout(n1085),.clk(gclk));
	jxor g1022(.dina(w_n1085_0[1]),.dinb(w_n1071_0[1]),.dout(n1086),.clk(gclk));
	jxor g1023(.dina(w_n1086_0[1]),.dinb(w_n1068_0[1]),.dout(n1087),.clk(gclk));
	jxor g1024(.dina(w_n1087_0[1]),.dinb(w_n1066_0[1]),.dout(n1088),.clk(gclk));
	jxor g1025(.dina(w_n1088_0[1]),.dinb(w_n1063_0[1]),.dout(n1089),.clk(gclk));
	jxor g1026(.dina(w_n1089_0[1]),.dinb(w_n1061_0[1]),.dout(n1090),.clk(gclk));
	jxor g1027(.dina(w_n1090_0[1]),.dinb(w_n1058_0[1]),.dout(n1091),.clk(gclk));
	jxor g1028(.dina(w_n1091_0[1]),.dinb(w_n1056_0[1]),.dout(n1092),.clk(gclk));
	jxor g1029(.dina(w_n1092_0[1]),.dinb(w_n1053_0[1]),.dout(n1093),.clk(gclk));
	jxor g1030(.dina(w_n1093_0[1]),.dinb(w_n1051_0[1]),.dout(n1094),.clk(gclk));
	jxor g1031(.dina(w_n1094_0[1]),.dinb(w_n1048_0[1]),.dout(n1095),.clk(gclk));
	jxor g1032(.dina(w_n1095_0[1]),.dinb(w_n1046_0[1]),.dout(n1096),.clk(gclk));
	jxor g1033(.dina(w_n1096_0[1]),.dinb(w_n1043_0[1]),.dout(n1097),.clk(gclk));
	jxor g1034(.dina(w_n1097_0[1]),.dinb(w_n1041_0[1]),.dout(n1098),.clk(gclk));
	jxor g1035(.dina(w_n1098_0[1]),.dinb(w_n1038_0[1]),.dout(n1099),.clk(gclk));
	jxor g1036(.dina(w_n1099_0[1]),.dinb(w_n1036_0[1]),.dout(n1100),.clk(gclk));
	jxor g1037(.dina(w_n1100_0[1]),.dinb(w_n1033_0[1]),.dout(n1101),.clk(gclk));
	jxor g1038(.dina(w_n1101_0[1]),.dinb(w_n1031_0[1]),.dout(n1102),.clk(gclk));
	jxor g1039(.dina(w_n1102_0[1]),.dinb(w_n1028_0[1]),.dout(n1103),.clk(gclk));
	jxor g1040(.dina(w_n1103_0[1]),.dinb(w_n1026_0[1]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(n1104),.dout(n1105),.clk(gclk));
	jxor g1042(.dina(w_n1105_0[1]),.dinb(w_n1023_0[1]),.dout(n1106),.clk(gclk));
	jxor g1043(.dina(w_n1106_0[1]),.dinb(w_n1022_0[1]),.dout(n1107),.clk(gclk));
	jxor g1044(.dina(w_n1107_0[1]),.dinb(w_n1018_0[1]),.dout(n1108),.clk(gclk));
	jxor g1045(.dina(w_n1108_0[1]),.dinb(w_n1017_0[1]),.dout(n1109),.clk(gclk));
	jnot g1046(.din(w_n1109_0[1]),.dout(n1110),.clk(gclk));
	jxor g1047(.dina(n1110),.dinb(w_n1013_0[1]),.dout(w_dff_A_SvwK5EUw5_2),.clk(gclk));
	jnot g1048(.din(w_n1108_0[0]),.dout(n1112),.clk(gclk));
	jor g1049(.dina(n1112),.dinb(w_n1017_0[0]),.dout(n1113),.clk(gclk));
	jor g1050(.dina(w_n1109_0[0]),.dinb(w_n1013_0[0]),.dout(n1114),.clk(gclk));
	jand g1051(.dina(n1114),.dinb(w_dff_B_Uj7K2SEj3_1),.dout(n1115),.clk(gclk));
	jnot g1052(.din(w_n1106_0[0]),.dout(n1116),.clk(gclk));
	jor g1053(.dina(n1116),.dinb(w_n1022_0[0]),.dout(n1117),.clk(gclk));
	jor g1054(.dina(w_n1107_0[0]),.dinb(w_n1018_0[0]),.dout(n1118),.clk(gclk));
	jand g1055(.dina(n1118),.dinb(n1117),.dout(n1119),.clk(gclk));
	jand g1056(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1120),.clk(gclk));
	jand g1057(.dina(w_n1103_0[0]),.dinb(w_n1026_0[0]),.dout(n1121),.clk(gclk));
	jnot g1058(.din(n1121),.dout(n1122),.clk(gclk));
	jor g1059(.dina(w_n1105_0[0]),.dinb(w_n1023_0[0]),.dout(n1123),.clk(gclk));
	jand g1060(.dina(n1123),.dinb(w_dff_B_2agerOhh0_1),.dout(n1124),.clk(gclk));
	jand g1061(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1125),.clk(gclk));
	jnot g1062(.din(n1125),.dout(n1126),.clk(gclk));
	jand g1063(.dina(w_n1101_0[0]),.dinb(w_n1031_0[0]),.dout(n1127),.clk(gclk));
	jand g1064(.dina(w_n1102_0[0]),.dinb(w_n1028_0[0]),.dout(n1128),.clk(gclk));
	jor g1065(.dina(n1128),.dinb(w_dff_B_ALbNq03a9_1),.dout(n1129),.clk(gclk));
	jand g1066(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1130),.clk(gclk));
	jnot g1067(.din(n1130),.dout(n1131),.clk(gclk));
	jand g1068(.dina(w_n1099_0[0]),.dinb(w_n1036_0[0]),.dout(n1132),.clk(gclk));
	jand g1069(.dina(w_n1100_0[0]),.dinb(w_n1033_0[0]),.dout(n1133),.clk(gclk));
	jor g1070(.dina(n1133),.dinb(w_dff_B_HfWrQ1Ho7_1),.dout(n1134),.clk(gclk));
	jand g1071(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1135),.clk(gclk));
	jnot g1072(.din(n1135),.dout(n1136),.clk(gclk));
	jand g1073(.dina(w_n1097_0[0]),.dinb(w_n1041_0[0]),.dout(n1137),.clk(gclk));
	jand g1074(.dina(w_n1098_0[0]),.dinb(w_n1038_0[0]),.dout(n1138),.clk(gclk));
	jor g1075(.dina(n1138),.dinb(w_dff_B_RZrP3vIZ0_1),.dout(n1139),.clk(gclk));
	jand g1076(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1140),.clk(gclk));
	jnot g1077(.din(n1140),.dout(n1141),.clk(gclk));
	jand g1078(.dina(w_n1095_0[0]),.dinb(w_n1046_0[0]),.dout(n1142),.clk(gclk));
	jand g1079(.dina(w_n1096_0[0]),.dinb(w_n1043_0[0]),.dout(n1143),.clk(gclk));
	jor g1080(.dina(n1143),.dinb(w_dff_B_1LktRM5K5_1),.dout(n1144),.clk(gclk));
	jand g1081(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1145),.clk(gclk));
	jnot g1082(.din(n1145),.dout(n1146),.clk(gclk));
	jand g1083(.dina(w_n1093_0[0]),.dinb(w_n1051_0[0]),.dout(n1147),.clk(gclk));
	jand g1084(.dina(w_n1094_0[0]),.dinb(w_n1048_0[0]),.dout(n1148),.clk(gclk));
	jor g1085(.dina(n1148),.dinb(w_dff_B_KmONAJPs5_1),.dout(n1149),.clk(gclk));
	jand g1086(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1150),.clk(gclk));
	jnot g1087(.din(n1150),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_n1091_0[0]),.dinb(w_n1056_0[0]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1092_0[0]),.dinb(w_n1053_0[0]),.dout(n1153),.clk(gclk));
	jor g1090(.dina(n1153),.dinb(w_dff_B_hbAs9MRE7_1),.dout(n1154),.clk(gclk));
	jand g1091(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1155),.clk(gclk));
	jnot g1092(.din(n1155),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_n1089_0[0]),.dinb(w_n1061_0[0]),.dout(n1157),.clk(gclk));
	jand g1094(.dina(w_n1090_0[0]),.dinb(w_n1058_0[0]),.dout(n1158),.clk(gclk));
	jor g1095(.dina(n1158),.dinb(w_dff_B_6uAOIO527_1),.dout(n1159),.clk(gclk));
	jand g1096(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1160),.clk(gclk));
	jnot g1097(.din(n1160),.dout(n1161),.clk(gclk));
	jand g1098(.dina(w_n1087_0[0]),.dinb(w_n1066_0[0]),.dout(n1162),.clk(gclk));
	jand g1099(.dina(w_n1088_0[0]),.dinb(w_n1063_0[0]),.dout(n1163),.clk(gclk));
	jor g1100(.dina(n1163),.dinb(w_dff_B_BuVg0Fal8_1),.dout(n1164),.clk(gclk));
	jand g1101(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1165),.clk(gclk));
	jnot g1102(.din(n1165),.dout(n1166),.clk(gclk));
	jand g1103(.dina(w_n1085_0[0]),.dinb(w_n1071_0[0]),.dout(n1167),.clk(gclk));
	jand g1104(.dina(w_n1086_0[0]),.dinb(w_n1068_0[0]),.dout(n1168),.clk(gclk));
	jor g1105(.dina(n1168),.dinb(w_dff_B_s9KZOleJ3_1),.dout(n1169),.clk(gclk));
	jand g1106(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1170),.clk(gclk));
	jnot g1107(.din(n1170),.dout(n1171),.clk(gclk));
	jand g1108(.dina(w_n1083_0[0]),.dinb(w_n1076_0[0]),.dout(n1172),.clk(gclk));
	jand g1109(.dina(w_n1084_0[0]),.dinb(w_n1073_0[0]),.dout(n1173),.clk(gclk));
	jor g1110(.dina(n1173),.dinb(w_dff_B_Ufyikq8N9_1),.dout(n1174),.clk(gclk));
	jand g1111(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1175),.clk(gclk));
	jand g1112(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1176),.clk(gclk));
	jor g1113(.dina(w_n1080_0[0]),.dinb(w_n1078_0[0]),.dout(n1177),.clk(gclk));
	jor g1114(.dina(w_n1082_0[0]),.dinb(w_n1077_0[0]),.dout(n1178),.clk(gclk));
	jand g1115(.dina(n1178),.dinb(w_dff_B_Gjt8d74j1_1),.dout(n1179),.clk(gclk));
	jxor g1116(.dina(w_n1179_0[1]),.dinb(w_n1176_0[1]),.dout(n1180),.clk(gclk));
	jnot g1117(.din(n1180),.dout(n1181),.clk(gclk));
	jxor g1118(.dina(w_n1181_0[1]),.dinb(w_n1175_0[1]),.dout(n1182),.clk(gclk));
	jxor g1119(.dina(w_n1182_0[1]),.dinb(w_n1174_0[1]),.dout(n1183),.clk(gclk));
	jxor g1120(.dina(w_n1183_0[1]),.dinb(w_n1171_0[1]),.dout(n1184),.clk(gclk));
	jxor g1121(.dina(w_n1184_0[1]),.dinb(w_n1169_0[1]),.dout(n1185),.clk(gclk));
	jxor g1122(.dina(w_n1185_0[1]),.dinb(w_n1166_0[1]),.dout(n1186),.clk(gclk));
	jxor g1123(.dina(w_n1186_0[1]),.dinb(w_n1164_0[1]),.dout(n1187),.clk(gclk));
	jxor g1124(.dina(w_n1187_0[1]),.dinb(w_n1161_0[1]),.dout(n1188),.clk(gclk));
	jxor g1125(.dina(w_n1188_0[1]),.dinb(w_n1159_0[1]),.dout(n1189),.clk(gclk));
	jxor g1126(.dina(w_n1189_0[1]),.dinb(w_n1156_0[1]),.dout(n1190),.clk(gclk));
	jxor g1127(.dina(w_n1190_0[1]),.dinb(w_n1154_0[1]),.dout(n1191),.clk(gclk));
	jxor g1128(.dina(w_n1191_0[1]),.dinb(w_n1151_0[1]),.dout(n1192),.clk(gclk));
	jxor g1129(.dina(w_n1192_0[1]),.dinb(w_n1149_0[1]),.dout(n1193),.clk(gclk));
	jxor g1130(.dina(w_n1193_0[1]),.dinb(w_n1146_0[1]),.dout(n1194),.clk(gclk));
	jxor g1131(.dina(w_n1194_0[1]),.dinb(w_n1144_0[1]),.dout(n1195),.clk(gclk));
	jxor g1132(.dina(w_n1195_0[1]),.dinb(w_n1141_0[1]),.dout(n1196),.clk(gclk));
	jxor g1133(.dina(w_n1196_0[1]),.dinb(w_n1139_0[1]),.dout(n1197),.clk(gclk));
	jxor g1134(.dina(w_n1197_0[1]),.dinb(w_n1136_0[1]),.dout(n1198),.clk(gclk));
	jxor g1135(.dina(w_n1198_0[1]),.dinb(w_n1134_0[1]),.dout(n1199),.clk(gclk));
	jxor g1136(.dina(w_n1199_0[1]),.dinb(w_n1131_0[1]),.dout(n1200),.clk(gclk));
	jxor g1137(.dina(w_n1200_0[1]),.dinb(w_n1129_0[1]),.dout(n1201),.clk(gclk));
	jxor g1138(.dina(w_n1201_0[1]),.dinb(w_n1126_0[1]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jxor g1140(.dina(w_n1203_0[1]),.dinb(w_n1124_0[1]),.dout(n1204),.clk(gclk));
	jnot g1141(.din(n1204),.dout(n1205),.clk(gclk));
	jxor g1142(.dina(w_n1205_0[1]),.dinb(w_n1120_0[1]),.dout(n1206),.clk(gclk));
	jxor g1143(.dina(w_n1206_0[1]),.dinb(w_n1119_0[1]),.dout(n1207),.clk(gclk));
	jnot g1144(.din(w_n1207_0[1]),.dout(n1208),.clk(gclk));
	jxor g1145(.dina(n1208),.dinb(w_n1115_0[1]),.dout(w_dff_A_EELcdX9T0_2),.clk(gclk));
	jnot g1146(.din(w_n1206_0[0]),.dout(n1210),.clk(gclk));
	jor g1147(.dina(n1210),.dinb(w_n1119_0[0]),.dout(n1211),.clk(gclk));
	jor g1148(.dina(w_n1207_0[0]),.dinb(w_n1115_0[0]),.dout(n1212),.clk(gclk));
	jand g1149(.dina(n1212),.dinb(w_dff_B_z5MYaKAx6_1),.dout(n1213),.clk(gclk));
	jor g1150(.dina(w_n1203_0[0]),.dinb(w_n1124_0[0]),.dout(n1214),.clk(gclk));
	jor g1151(.dina(w_n1205_0[0]),.dinb(w_n1120_0[0]),.dout(n1215),.clk(gclk));
	jand g1152(.dina(n1215),.dinb(w_dff_B_oqfRcZfn8_1),.dout(n1216),.clk(gclk));
	jand g1153(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1217),.clk(gclk));
	jand g1154(.dina(w_n1200_0[0]),.dinb(w_n1129_0[0]),.dout(n1218),.clk(gclk));
	jand g1155(.dina(w_n1201_0[0]),.dinb(w_n1126_0[0]),.dout(n1219),.clk(gclk));
	jor g1156(.dina(n1219),.dinb(w_dff_B_5b7MHFLe9_1),.dout(n1220),.clk(gclk));
	jand g1157(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1221),.clk(gclk));
	jnot g1158(.din(n1221),.dout(n1222),.clk(gclk));
	jand g1159(.dina(w_n1198_0[0]),.dinb(w_n1134_0[0]),.dout(n1223),.clk(gclk));
	jand g1160(.dina(w_n1199_0[0]),.dinb(w_n1131_0[0]),.dout(n1224),.clk(gclk));
	jor g1161(.dina(n1224),.dinb(w_dff_B_fiwM2wYC8_1),.dout(n1225),.clk(gclk));
	jand g1162(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1226),.clk(gclk));
	jnot g1163(.din(n1226),.dout(n1227),.clk(gclk));
	jand g1164(.dina(w_n1196_0[0]),.dinb(w_n1139_0[0]),.dout(n1228),.clk(gclk));
	jand g1165(.dina(w_n1197_0[0]),.dinb(w_n1136_0[0]),.dout(n1229),.clk(gclk));
	jor g1166(.dina(n1229),.dinb(w_dff_B_mv68vdNy4_1),.dout(n1230),.clk(gclk));
	jand g1167(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1231),.clk(gclk));
	jnot g1168(.din(n1231),.dout(n1232),.clk(gclk));
	jand g1169(.dina(w_n1194_0[0]),.dinb(w_n1144_0[0]),.dout(n1233),.clk(gclk));
	jand g1170(.dina(w_n1195_0[0]),.dinb(w_n1141_0[0]),.dout(n1234),.clk(gclk));
	jor g1171(.dina(n1234),.dinb(w_dff_B_uK9k6vOp8_1),.dout(n1235),.clk(gclk));
	jand g1172(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1236),.clk(gclk));
	jnot g1173(.din(n1236),.dout(n1237),.clk(gclk));
	jand g1174(.dina(w_n1192_0[0]),.dinb(w_n1149_0[0]),.dout(n1238),.clk(gclk));
	jand g1175(.dina(w_n1193_0[0]),.dinb(w_n1146_0[0]),.dout(n1239),.clk(gclk));
	jor g1176(.dina(n1239),.dinb(w_dff_B_Gsa8nd0s8_1),.dout(n1240),.clk(gclk));
	jand g1177(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1241),.clk(gclk));
	jnot g1178(.din(n1241),.dout(n1242),.clk(gclk));
	jand g1179(.dina(w_n1190_0[0]),.dinb(w_n1154_0[0]),.dout(n1243),.clk(gclk));
	jand g1180(.dina(w_n1191_0[0]),.dinb(w_n1151_0[0]),.dout(n1244),.clk(gclk));
	jor g1181(.dina(n1244),.dinb(w_dff_B_gdrGJvfb5_1),.dout(n1245),.clk(gclk));
	jand g1182(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1246),.clk(gclk));
	jnot g1183(.din(n1246),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_n1188_0[0]),.dinb(w_n1159_0[0]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1189_0[0]),.dinb(w_n1156_0[0]),.dout(n1249),.clk(gclk));
	jor g1186(.dina(n1249),.dinb(w_dff_B_C3FFnonp9_1),.dout(n1250),.clk(gclk));
	jand g1187(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1251),.clk(gclk));
	jnot g1188(.din(n1251),.dout(n1252),.clk(gclk));
	jand g1189(.dina(w_n1186_0[0]),.dinb(w_n1164_0[0]),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1187_0[0]),.dinb(w_n1161_0[0]),.dout(n1254),.clk(gclk));
	jor g1191(.dina(n1254),.dinb(w_dff_B_QSeZHBz11_1),.dout(n1255),.clk(gclk));
	jand g1192(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1256),.clk(gclk));
	jnot g1193(.din(n1256),.dout(n1257),.clk(gclk));
	jand g1194(.dina(w_n1184_0[0]),.dinb(w_n1169_0[0]),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1185_0[0]),.dinb(w_n1166_0[0]),.dout(n1259),.clk(gclk));
	jor g1196(.dina(n1259),.dinb(w_dff_B_mjBQCs7h3_1),.dout(n1260),.clk(gclk));
	jand g1197(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1261),.clk(gclk));
	jnot g1198(.din(n1261),.dout(n1262),.clk(gclk));
	jand g1199(.dina(w_n1182_0[0]),.dinb(w_n1174_0[0]),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1183_0[0]),.dinb(w_n1171_0[0]),.dout(n1264),.clk(gclk));
	jor g1201(.dina(n1264),.dinb(w_dff_B_zd2kEF9W7_1),.dout(n1265),.clk(gclk));
	jand g1202(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1266),.clk(gclk));
	jand g1203(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1267),.clk(gclk));
	jor g1204(.dina(w_n1179_0[0]),.dinb(w_n1176_0[0]),.dout(n1268),.clk(gclk));
	jor g1205(.dina(w_n1181_0[0]),.dinb(w_n1175_0[0]),.dout(n1269),.clk(gclk));
	jand g1206(.dina(n1269),.dinb(w_dff_B_CSsJu4ca9_1),.dout(n1270),.clk(gclk));
	jxor g1207(.dina(w_n1270_0[1]),.dinb(w_n1267_0[1]),.dout(n1271),.clk(gclk));
	jnot g1208(.din(n1271),.dout(n1272),.clk(gclk));
	jxor g1209(.dina(w_n1272_0[1]),.dinb(w_n1266_0[1]),.dout(n1273),.clk(gclk));
	jxor g1210(.dina(w_n1273_0[1]),.dinb(w_n1265_0[1]),.dout(n1274),.clk(gclk));
	jxor g1211(.dina(w_n1274_0[1]),.dinb(w_n1262_0[1]),.dout(n1275),.clk(gclk));
	jxor g1212(.dina(w_n1275_0[1]),.dinb(w_n1260_0[1]),.dout(n1276),.clk(gclk));
	jxor g1213(.dina(w_n1276_0[1]),.dinb(w_n1257_0[1]),.dout(n1277),.clk(gclk));
	jxor g1214(.dina(w_n1277_0[1]),.dinb(w_n1255_0[1]),.dout(n1278),.clk(gclk));
	jxor g1215(.dina(w_n1278_0[1]),.dinb(w_n1252_0[1]),.dout(n1279),.clk(gclk));
	jxor g1216(.dina(w_n1279_0[1]),.dinb(w_n1250_0[1]),.dout(n1280),.clk(gclk));
	jxor g1217(.dina(w_n1280_0[1]),.dinb(w_n1247_0[1]),.dout(n1281),.clk(gclk));
	jxor g1218(.dina(w_n1281_0[1]),.dinb(w_n1245_0[1]),.dout(n1282),.clk(gclk));
	jxor g1219(.dina(w_n1282_0[1]),.dinb(w_n1242_0[1]),.dout(n1283),.clk(gclk));
	jxor g1220(.dina(w_n1283_0[1]),.dinb(w_n1240_0[1]),.dout(n1284),.clk(gclk));
	jxor g1221(.dina(w_n1284_0[1]),.dinb(w_n1237_0[1]),.dout(n1285),.clk(gclk));
	jxor g1222(.dina(w_n1285_0[1]),.dinb(w_n1235_0[1]),.dout(n1286),.clk(gclk));
	jxor g1223(.dina(w_n1286_0[1]),.dinb(w_n1232_0[1]),.dout(n1287),.clk(gclk));
	jxor g1224(.dina(w_n1287_0[1]),.dinb(w_n1230_0[1]),.dout(n1288),.clk(gclk));
	jxor g1225(.dina(w_n1288_0[1]),.dinb(w_n1227_0[1]),.dout(n1289),.clk(gclk));
	jxor g1226(.dina(w_n1289_0[1]),.dinb(w_n1225_0[1]),.dout(n1290),.clk(gclk));
	jxor g1227(.dina(w_n1290_0[1]),.dinb(w_n1222_0[1]),.dout(n1291),.clk(gclk));
	jxor g1228(.dina(w_n1291_0[1]),.dinb(w_n1220_0[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jxor g1230(.dina(w_n1293_0[1]),.dinb(w_n1217_0[1]),.dout(n1294),.clk(gclk));
	jxor g1231(.dina(w_n1294_0[1]),.dinb(w_n1216_0[1]),.dout(n1295),.clk(gclk));
	jnot g1232(.din(w_n1295_0[1]),.dout(n1296),.clk(gclk));
	jxor g1233(.dina(w_dff_B_7zYdlvs98_0),.dinb(w_n1213_0[1]),.dout(w_dff_A_RRpqyqj39_2),.clk(gclk));
	jnot g1234(.din(w_n1294_0[0]),.dout(n1298),.clk(gclk));
	jor g1235(.dina(w_dff_B_eXsPARqE7_0),.dinb(w_n1216_0[0]),.dout(n1299),.clk(gclk));
	jor g1236(.dina(w_n1295_0[0]),.dinb(w_n1213_0[0]),.dout(n1300),.clk(gclk));
	jand g1237(.dina(n1300),.dinb(w_dff_B_jS3TSOxf8_1),.dout(n1301),.clk(gclk));
	jnot g1238(.din(w_n1220_0[0]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(w_n1291_0[0]),.dout(n1303),.clk(gclk));
	jor g1240(.dina(w_dff_B_DIbn7qAF3_0),.dinb(n1302),.dout(n1304),.clk(gclk));
	jor g1241(.dina(w_n1293_0[0]),.dinb(w_n1217_0[0]),.dout(n1305),.clk(gclk));
	jand g1242(.dina(n1305),.dinb(w_dff_B_0Tq9flrP8_1),.dout(n1306),.clk(gclk));
	jand g1243(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1307),.clk(gclk));
	jand g1244(.dina(w_n1289_0[0]),.dinb(w_n1225_0[0]),.dout(n1308),.clk(gclk));
	jand g1245(.dina(w_n1290_0[0]),.dinb(w_n1222_0[0]),.dout(n1309),.clk(gclk));
	jor g1246(.dina(n1309),.dinb(w_dff_B_k8XlVUA97_1),.dout(n1310),.clk(gclk));
	jand g1247(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1311),.clk(gclk));
	jnot g1248(.din(n1311),.dout(n1312),.clk(gclk));
	jand g1249(.dina(w_n1287_0[0]),.dinb(w_n1230_0[0]),.dout(n1313),.clk(gclk));
	jand g1250(.dina(w_n1288_0[0]),.dinb(w_n1227_0[0]),.dout(n1314),.clk(gclk));
	jor g1251(.dina(n1314),.dinb(w_dff_B_0H3Hy2HC2_1),.dout(n1315),.clk(gclk));
	jand g1252(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1316),.clk(gclk));
	jnot g1253(.din(n1316),.dout(n1317),.clk(gclk));
	jand g1254(.dina(w_n1285_0[0]),.dinb(w_n1235_0[0]),.dout(n1318),.clk(gclk));
	jand g1255(.dina(w_n1286_0[0]),.dinb(w_n1232_0[0]),.dout(n1319),.clk(gclk));
	jor g1256(.dina(n1319),.dinb(w_dff_B_m5BQ8Cor6_1),.dout(n1320),.clk(gclk));
	jand g1257(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1321),.clk(gclk));
	jnot g1258(.din(n1321),.dout(n1322),.clk(gclk));
	jand g1259(.dina(w_n1283_0[0]),.dinb(w_n1240_0[0]),.dout(n1323),.clk(gclk));
	jand g1260(.dina(w_n1284_0[0]),.dinb(w_n1237_0[0]),.dout(n1324),.clk(gclk));
	jor g1261(.dina(n1324),.dinb(w_dff_B_1MmuV6Vb7_1),.dout(n1325),.clk(gclk));
	jand g1262(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(n1326),.dout(n1327),.clk(gclk));
	jand g1264(.dina(w_n1281_0[0]),.dinb(w_n1245_0[0]),.dout(n1328),.clk(gclk));
	jand g1265(.dina(w_n1282_0[0]),.dinb(w_n1242_0[0]),.dout(n1329),.clk(gclk));
	jor g1266(.dina(n1329),.dinb(w_dff_B_DgelcY9s0_1),.dout(n1330),.clk(gclk));
	jand g1267(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1331),.clk(gclk));
	jnot g1268(.din(n1331),.dout(n1332),.clk(gclk));
	jand g1269(.dina(w_n1279_0[0]),.dinb(w_n1250_0[0]),.dout(n1333),.clk(gclk));
	jand g1270(.dina(w_n1280_0[0]),.dinb(w_n1247_0[0]),.dout(n1334),.clk(gclk));
	jor g1271(.dina(n1334),.dinb(w_dff_B_aLxXaBkb0_1),.dout(n1335),.clk(gclk));
	jand g1272(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1336),.clk(gclk));
	jnot g1273(.din(n1336),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_n1277_0[0]),.dinb(w_n1255_0[0]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1278_0[0]),.dinb(w_n1252_0[0]),.dout(n1339),.clk(gclk));
	jor g1276(.dina(n1339),.dinb(w_dff_B_c1etSVAc6_1),.dout(n1340),.clk(gclk));
	jand g1277(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1341),.clk(gclk));
	jnot g1278(.din(n1341),.dout(n1342),.clk(gclk));
	jand g1279(.dina(w_n1275_0[0]),.dinb(w_n1260_0[0]),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1276_0[0]),.dinb(w_n1257_0[0]),.dout(n1344),.clk(gclk));
	jor g1281(.dina(n1344),.dinb(w_dff_B_hdB6e6E61_1),.dout(n1345),.clk(gclk));
	jand g1282(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1346),.clk(gclk));
	jnot g1283(.din(n1346),.dout(n1347),.clk(gclk));
	jand g1284(.dina(w_n1273_0[0]),.dinb(w_n1265_0[0]),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1274_0[0]),.dinb(w_n1262_0[0]),.dout(n1349),.clk(gclk));
	jor g1286(.dina(n1349),.dinb(w_dff_B_3mVv4DRR9_1),.dout(n1350),.clk(gclk));
	jand g1287(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1351),.clk(gclk));
	jand g1288(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1352),.clk(gclk));
	jor g1289(.dina(w_n1270_0[0]),.dinb(w_n1267_0[0]),.dout(n1353),.clk(gclk));
	jor g1290(.dina(w_n1272_0[0]),.dinb(w_n1266_0[0]),.dout(n1354),.clk(gclk));
	jand g1291(.dina(n1354),.dinb(w_dff_B_O9rLtxNu0_1),.dout(n1355),.clk(gclk));
	jxor g1292(.dina(w_n1355_0[1]),.dinb(w_n1352_0[1]),.dout(n1356),.clk(gclk));
	jnot g1293(.din(n1356),.dout(n1357),.clk(gclk));
	jxor g1294(.dina(w_n1357_0[1]),.dinb(w_n1351_0[1]),.dout(n1358),.clk(gclk));
	jxor g1295(.dina(w_n1358_0[1]),.dinb(w_n1350_0[1]),.dout(n1359),.clk(gclk));
	jxor g1296(.dina(w_n1359_0[1]),.dinb(w_n1347_0[1]),.dout(n1360),.clk(gclk));
	jxor g1297(.dina(w_n1360_0[1]),.dinb(w_n1345_0[1]),.dout(n1361),.clk(gclk));
	jxor g1298(.dina(w_n1361_0[1]),.dinb(w_n1342_0[1]),.dout(n1362),.clk(gclk));
	jxor g1299(.dina(w_n1362_0[1]),.dinb(w_n1340_0[1]),.dout(n1363),.clk(gclk));
	jxor g1300(.dina(w_n1363_0[1]),.dinb(w_n1337_0[1]),.dout(n1364),.clk(gclk));
	jxor g1301(.dina(w_n1364_0[1]),.dinb(w_n1335_0[1]),.dout(n1365),.clk(gclk));
	jxor g1302(.dina(w_n1365_0[1]),.dinb(w_n1332_0[1]),.dout(n1366),.clk(gclk));
	jxor g1303(.dina(w_n1366_0[1]),.dinb(w_n1330_0[1]),.dout(n1367),.clk(gclk));
	jxor g1304(.dina(w_n1367_0[1]),.dinb(w_n1327_0[1]),.dout(n1368),.clk(gclk));
	jxor g1305(.dina(w_n1368_0[1]),.dinb(w_n1325_0[1]),.dout(n1369),.clk(gclk));
	jxor g1306(.dina(w_n1369_0[1]),.dinb(w_n1322_0[1]),.dout(n1370),.clk(gclk));
	jxor g1307(.dina(w_n1370_0[1]),.dinb(w_n1320_0[1]),.dout(n1371),.clk(gclk));
	jxor g1308(.dina(w_n1371_0[1]),.dinb(w_n1317_0[1]),.dout(n1372),.clk(gclk));
	jxor g1309(.dina(w_n1372_0[1]),.dinb(w_n1315_0[1]),.dout(n1373),.clk(gclk));
	jxor g1310(.dina(w_n1373_0[1]),.dinb(w_n1312_0[1]),.dout(n1374),.clk(gclk));
	jxor g1311(.dina(w_n1374_0[1]),.dinb(w_n1310_0[1]),.dout(n1375),.clk(gclk));
	jnot g1312(.din(n1375),.dout(n1376),.clk(gclk));
	jxor g1313(.dina(w_n1376_0[1]),.dinb(w_n1307_0[1]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jxor g1315(.dina(w_n1378_0[1]),.dinb(w_n1306_0[1]),.dout(n1379),.clk(gclk));
	jxor g1316(.dina(w_n1379_0[1]),.dinb(w_n1301_0[1]),.dout(w_dff_A_qnZGkGXX4_2),.clk(gclk));
	jor g1317(.dina(w_n1378_0[0]),.dinb(w_n1306_0[0]),.dout(n1381),.clk(gclk));
	jnot g1318(.din(w_n1379_0[0]),.dout(n1382),.clk(gclk));
	jor g1319(.dina(w_dff_B_hVTh9bVH3_0),.dinb(w_n1301_0[0]),.dout(n1383),.clk(gclk));
	jand g1320(.dina(n1383),.dinb(w_dff_B_wlGQ1Lsq0_1),.dout(n1384),.clk(gclk));
	jnot g1321(.din(w_n1310_0[0]),.dout(n1385),.clk(gclk));
	jnot g1322(.din(w_n1374_0[0]),.dout(n1386),.clk(gclk));
	jor g1323(.dina(n1386),.dinb(n1385),.dout(n1387),.clk(gclk));
	jor g1324(.dina(w_n1376_0[0]),.dinb(w_n1307_0[0]),.dout(n1388),.clk(gclk));
	jand g1325(.dina(n1388),.dinb(w_dff_B_3Elpi5LQ4_1),.dout(n1389),.clk(gclk));
	jand g1326(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1390),.clk(gclk));
	jand g1327(.dina(w_n1372_0[0]),.dinb(w_n1315_0[0]),.dout(n1391),.clk(gclk));
	jand g1328(.dina(w_n1373_0[0]),.dinb(w_n1312_0[0]),.dout(n1392),.clk(gclk));
	jor g1329(.dina(n1392),.dinb(w_dff_B_NdHYw2Ji4_1),.dout(n1393),.clk(gclk));
	jand g1330(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1394),.clk(gclk));
	jnot g1331(.din(n1394),.dout(n1395),.clk(gclk));
	jand g1332(.dina(w_n1370_0[0]),.dinb(w_n1320_0[0]),.dout(n1396),.clk(gclk));
	jand g1333(.dina(w_n1371_0[0]),.dinb(w_n1317_0[0]),.dout(n1397),.clk(gclk));
	jor g1334(.dina(n1397),.dinb(w_dff_B_72didT1E7_1),.dout(n1398),.clk(gclk));
	jand g1335(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1399),.clk(gclk));
	jnot g1336(.din(n1399),.dout(n1400),.clk(gclk));
	jand g1337(.dina(w_n1368_0[0]),.dinb(w_n1325_0[0]),.dout(n1401),.clk(gclk));
	jand g1338(.dina(w_n1369_0[0]),.dinb(w_n1322_0[0]),.dout(n1402),.clk(gclk));
	jor g1339(.dina(n1402),.dinb(w_dff_B_lqFfUgs60_1),.dout(n1403),.clk(gclk));
	jand g1340(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1404),.clk(gclk));
	jnot g1341(.din(n1404),.dout(n1405),.clk(gclk));
	jand g1342(.dina(w_n1366_0[0]),.dinb(w_n1330_0[0]),.dout(n1406),.clk(gclk));
	jand g1343(.dina(w_n1367_0[0]),.dinb(w_n1327_0[0]),.dout(n1407),.clk(gclk));
	jor g1344(.dina(n1407),.dinb(w_dff_B_g8XKJVFw3_1),.dout(n1408),.clk(gclk));
	jand g1345(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1409),.clk(gclk));
	jnot g1346(.din(n1409),.dout(n1410),.clk(gclk));
	jand g1347(.dina(w_n1364_0[0]),.dinb(w_n1335_0[0]),.dout(n1411),.clk(gclk));
	jand g1348(.dina(w_n1365_0[0]),.dinb(w_n1332_0[0]),.dout(n1412),.clk(gclk));
	jor g1349(.dina(n1412),.dinb(w_dff_B_AGOGhga26_1),.dout(n1413),.clk(gclk));
	jand g1350(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1414),.clk(gclk));
	jnot g1351(.din(n1414),.dout(n1415),.clk(gclk));
	jand g1352(.dina(w_n1362_0[0]),.dinb(w_n1340_0[0]),.dout(n1416),.clk(gclk));
	jand g1353(.dina(w_n1363_0[0]),.dinb(w_n1337_0[0]),.dout(n1417),.clk(gclk));
	jor g1354(.dina(n1417),.dinb(w_dff_B_JDhLY78t9_1),.dout(n1418),.clk(gclk));
	jand g1355(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1419),.clk(gclk));
	jnot g1356(.din(n1419),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_n1360_0[0]),.dinb(w_n1345_0[0]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1361_0[0]),.dinb(w_n1342_0[0]),.dout(n1422),.clk(gclk));
	jor g1359(.dina(n1422),.dinb(w_dff_B_n19aq9WK1_1),.dout(n1423),.clk(gclk));
	jand g1360(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1424),.clk(gclk));
	jnot g1361(.din(n1424),.dout(n1425),.clk(gclk));
	jand g1362(.dina(w_n1358_0[0]),.dinb(w_n1350_0[0]),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1359_0[0]),.dinb(w_n1347_0[0]),.dout(n1427),.clk(gclk));
	jor g1364(.dina(n1427),.dinb(w_dff_B_0bFHJie74_1),.dout(n1428),.clk(gclk));
	jand g1365(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1429),.clk(gclk));
	jand g1366(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1430),.clk(gclk));
	jor g1367(.dina(w_n1355_0[0]),.dinb(w_n1352_0[0]),.dout(n1431),.clk(gclk));
	jor g1368(.dina(w_n1357_0[0]),.dinb(w_n1351_0[0]),.dout(n1432),.clk(gclk));
	jand g1369(.dina(n1432),.dinb(w_dff_B_kUPrBYtM2_1),.dout(n1433),.clk(gclk));
	jxor g1370(.dina(w_n1433_0[1]),.dinb(w_n1430_0[1]),.dout(n1434),.clk(gclk));
	jnot g1371(.din(n1434),.dout(n1435),.clk(gclk));
	jxor g1372(.dina(w_n1435_0[1]),.dinb(w_n1429_0[1]),.dout(n1436),.clk(gclk));
	jxor g1373(.dina(w_n1436_0[1]),.dinb(w_n1428_0[1]),.dout(n1437),.clk(gclk));
	jxor g1374(.dina(w_n1437_0[1]),.dinb(w_n1425_0[1]),.dout(n1438),.clk(gclk));
	jxor g1375(.dina(w_n1438_0[1]),.dinb(w_n1423_0[1]),.dout(n1439),.clk(gclk));
	jxor g1376(.dina(w_n1439_0[1]),.dinb(w_n1420_0[1]),.dout(n1440),.clk(gclk));
	jxor g1377(.dina(w_n1440_0[1]),.dinb(w_n1418_0[1]),.dout(n1441),.clk(gclk));
	jxor g1378(.dina(w_n1441_0[1]),.dinb(w_n1415_0[1]),.dout(n1442),.clk(gclk));
	jxor g1379(.dina(w_n1442_0[1]),.dinb(w_n1413_0[1]),.dout(n1443),.clk(gclk));
	jxor g1380(.dina(w_n1443_0[1]),.dinb(w_n1410_0[1]),.dout(n1444),.clk(gclk));
	jxor g1381(.dina(w_n1444_0[1]),.dinb(w_n1408_0[1]),.dout(n1445),.clk(gclk));
	jxor g1382(.dina(w_n1445_0[1]),.dinb(w_n1405_0[1]),.dout(n1446),.clk(gclk));
	jxor g1383(.dina(w_n1446_0[1]),.dinb(w_n1403_0[1]),.dout(n1447),.clk(gclk));
	jxor g1384(.dina(w_n1447_0[1]),.dinb(w_n1400_0[1]),.dout(n1448),.clk(gclk));
	jxor g1385(.dina(w_n1448_0[1]),.dinb(w_n1398_0[1]),.dout(n1449),.clk(gclk));
	jxor g1386(.dina(w_n1449_0[1]),.dinb(w_n1395_0[1]),.dout(n1450),.clk(gclk));
	jxor g1387(.dina(w_n1450_0[1]),.dinb(w_n1393_0[1]),.dout(n1451),.clk(gclk));
	jnot g1388(.din(n1451),.dout(n1452),.clk(gclk));
	jxor g1389(.dina(w_n1452_0[1]),.dinb(w_n1390_0[1]),.dout(n1453),.clk(gclk));
	jnot g1390(.din(n1453),.dout(n1454),.clk(gclk));
	jxor g1391(.dina(w_n1454_0[1]),.dinb(w_n1389_0[1]),.dout(n1455),.clk(gclk));
	jxor g1392(.dina(w_n1455_0[1]),.dinb(w_n1384_0[1]),.dout(w_dff_A_WXOrmoWW8_2),.clk(gclk));
	jor g1393(.dina(w_n1454_0[0]),.dinb(w_n1389_0[0]),.dout(n1457),.clk(gclk));
	jnot g1394(.din(w_n1455_0[0]),.dout(n1458),.clk(gclk));
	jor g1395(.dina(w_dff_B_BjqKJUgd6_0),.dinb(w_n1384_0[0]),.dout(n1459),.clk(gclk));
	jand g1396(.dina(n1459),.dinb(w_dff_B_Jum1WBO27_1),.dout(n1460),.clk(gclk));
	jnot g1397(.din(w_n1393_0[0]),.dout(n1461),.clk(gclk));
	jnot g1398(.din(w_n1450_0[0]),.dout(n1462),.clk(gclk));
	jor g1399(.dina(n1462),.dinb(n1461),.dout(n1463),.clk(gclk));
	jor g1400(.dina(w_n1452_0[0]),.dinb(w_n1390_0[0]),.dout(n1464),.clk(gclk));
	jand g1401(.dina(n1464),.dinb(w_dff_B_tyeEbBLJ7_1),.dout(n1465),.clk(gclk));
	jand g1402(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1466),.clk(gclk));
	jand g1403(.dina(w_n1448_0[0]),.dinb(w_n1398_0[0]),.dout(n1467),.clk(gclk));
	jand g1404(.dina(w_n1449_0[0]),.dinb(w_n1395_0[0]),.dout(n1468),.clk(gclk));
	jor g1405(.dina(n1468),.dinb(w_dff_B_SwruDX775_1),.dout(n1469),.clk(gclk));
	jand g1406(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1470),.clk(gclk));
	jnot g1407(.din(n1470),.dout(n1471),.clk(gclk));
	jand g1408(.dina(w_n1446_0[0]),.dinb(w_n1403_0[0]),.dout(n1472),.clk(gclk));
	jand g1409(.dina(w_n1447_0[0]),.dinb(w_n1400_0[0]),.dout(n1473),.clk(gclk));
	jor g1410(.dina(n1473),.dinb(w_dff_B_zcHUBgZ90_1),.dout(n1474),.clk(gclk));
	jand g1411(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1475),.clk(gclk));
	jnot g1412(.din(n1475),.dout(n1476),.clk(gclk));
	jand g1413(.dina(w_n1444_0[0]),.dinb(w_n1408_0[0]),.dout(n1477),.clk(gclk));
	jand g1414(.dina(w_n1445_0[0]),.dinb(w_n1405_0[0]),.dout(n1478),.clk(gclk));
	jor g1415(.dina(n1478),.dinb(w_dff_B_m02Mw1jm9_1),.dout(n1479),.clk(gclk));
	jand g1416(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1480),.clk(gclk));
	jnot g1417(.din(n1480),.dout(n1481),.clk(gclk));
	jand g1418(.dina(w_n1442_0[0]),.dinb(w_n1413_0[0]),.dout(n1482),.clk(gclk));
	jand g1419(.dina(w_n1443_0[0]),.dinb(w_n1410_0[0]),.dout(n1483),.clk(gclk));
	jor g1420(.dina(n1483),.dinb(w_dff_B_hpSnetn01_1),.dout(n1484),.clk(gclk));
	jand g1421(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1485),.clk(gclk));
	jnot g1422(.din(n1485),.dout(n1486),.clk(gclk));
	jand g1423(.dina(w_n1440_0[0]),.dinb(w_n1418_0[0]),.dout(n1487),.clk(gclk));
	jand g1424(.dina(w_n1441_0[0]),.dinb(w_n1415_0[0]),.dout(n1488),.clk(gclk));
	jor g1425(.dina(n1488),.dinb(w_dff_B_NOMqsQbb7_1),.dout(n1489),.clk(gclk));
	jand g1426(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1490),.clk(gclk));
	jnot g1427(.din(n1490),.dout(n1491),.clk(gclk));
	jand g1428(.dina(w_n1438_0[0]),.dinb(w_n1423_0[0]),.dout(n1492),.clk(gclk));
	jand g1429(.dina(w_n1439_0[0]),.dinb(w_n1420_0[0]),.dout(n1493),.clk(gclk));
	jor g1430(.dina(n1493),.dinb(w_dff_B_1lgDSPcO0_1),.dout(n1494),.clk(gclk));
	jand g1431(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1495),.clk(gclk));
	jnot g1432(.din(n1495),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_n1436_0[0]),.dinb(w_n1428_0[0]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1437_0[0]),.dinb(w_n1425_0[0]),.dout(n1498),.clk(gclk));
	jor g1435(.dina(n1498),.dinb(w_dff_B_Nxts0IYw7_1),.dout(n1499),.clk(gclk));
	jand g1436(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1500),.clk(gclk));
	jand g1437(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1501),.clk(gclk));
	jor g1438(.dina(w_n1433_0[0]),.dinb(w_n1430_0[0]),.dout(n1502),.clk(gclk));
	jor g1439(.dina(w_n1435_0[0]),.dinb(w_n1429_0[0]),.dout(n1503),.clk(gclk));
	jand g1440(.dina(n1503),.dinb(w_dff_B_O4pQZRa68_1),.dout(n1504),.clk(gclk));
	jxor g1441(.dina(w_n1504_0[1]),.dinb(w_n1501_0[1]),.dout(n1505),.clk(gclk));
	jnot g1442(.din(n1505),.dout(n1506),.clk(gclk));
	jxor g1443(.dina(w_n1506_0[1]),.dinb(w_n1500_0[1]),.dout(n1507),.clk(gclk));
	jxor g1444(.dina(w_n1507_0[1]),.dinb(w_n1499_0[1]),.dout(n1508),.clk(gclk));
	jxor g1445(.dina(w_n1508_0[1]),.dinb(w_n1496_0[1]),.dout(n1509),.clk(gclk));
	jxor g1446(.dina(w_n1509_0[1]),.dinb(w_n1494_0[1]),.dout(n1510),.clk(gclk));
	jxor g1447(.dina(w_n1510_0[1]),.dinb(w_n1491_0[1]),.dout(n1511),.clk(gclk));
	jxor g1448(.dina(w_n1511_0[1]),.dinb(w_n1489_0[1]),.dout(n1512),.clk(gclk));
	jxor g1449(.dina(w_n1512_0[1]),.dinb(w_n1486_0[1]),.dout(n1513),.clk(gclk));
	jxor g1450(.dina(w_n1513_0[1]),.dinb(w_n1484_0[1]),.dout(n1514),.clk(gclk));
	jxor g1451(.dina(w_n1514_0[1]),.dinb(w_n1481_0[1]),.dout(n1515),.clk(gclk));
	jxor g1452(.dina(w_n1515_0[1]),.dinb(w_n1479_0[1]),.dout(n1516),.clk(gclk));
	jxor g1453(.dina(w_n1516_0[1]),.dinb(w_n1476_0[1]),.dout(n1517),.clk(gclk));
	jxor g1454(.dina(w_n1517_0[1]),.dinb(w_n1474_0[1]),.dout(n1518),.clk(gclk));
	jxor g1455(.dina(w_n1518_0[1]),.dinb(w_n1471_0[1]),.dout(n1519),.clk(gclk));
	jxor g1456(.dina(w_n1519_0[1]),.dinb(w_n1469_0[1]),.dout(n1520),.clk(gclk));
	jnot g1457(.din(n1520),.dout(n1521),.clk(gclk));
	jxor g1458(.dina(w_n1521_0[1]),.dinb(w_n1466_0[1]),.dout(n1522),.clk(gclk));
	jnot g1459(.din(n1522),.dout(n1523),.clk(gclk));
	jxor g1460(.dina(w_n1523_0[1]),.dinb(w_n1465_0[1]),.dout(n1524),.clk(gclk));
	jxor g1461(.dina(w_n1524_0[1]),.dinb(w_n1460_0[1]),.dout(w_dff_A_zBf6HHia3_2),.clk(gclk));
	jor g1462(.dina(w_n1523_0[0]),.dinb(w_n1465_0[0]),.dout(n1526),.clk(gclk));
	jnot g1463(.din(w_n1524_0[0]),.dout(n1527),.clk(gclk));
	jor g1464(.dina(w_dff_B_tlSTntkM6_0),.dinb(w_n1460_0[0]),.dout(n1528),.clk(gclk));
	jand g1465(.dina(n1528),.dinb(w_dff_B_tnRGkghO1_1),.dout(n1529),.clk(gclk));
	jnot g1466(.din(w_n1469_0[0]),.dout(n1530),.clk(gclk));
	jnot g1467(.din(w_n1519_0[0]),.dout(n1531),.clk(gclk));
	jor g1468(.dina(w_dff_B_Ed9BH3408_0),.dinb(n1530),.dout(n1532),.clk(gclk));
	jor g1469(.dina(w_n1521_0[0]),.dinb(w_n1466_0[0]),.dout(n1533),.clk(gclk));
	jand g1470(.dina(n1533),.dinb(w_dff_B_ro5cP48Y3_1),.dout(n1534),.clk(gclk));
	jand g1471(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1535),.clk(gclk));
	jand g1472(.dina(w_n1517_0[0]),.dinb(w_n1474_0[0]),.dout(n1536),.clk(gclk));
	jand g1473(.dina(w_n1518_0[0]),.dinb(w_n1471_0[0]),.dout(n1537),.clk(gclk));
	jor g1474(.dina(n1537),.dinb(w_dff_B_mwxOl5mb9_1),.dout(n1538),.clk(gclk));
	jand g1475(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1539),.clk(gclk));
	jnot g1476(.din(n1539),.dout(n1540),.clk(gclk));
	jand g1477(.dina(w_n1515_0[0]),.dinb(w_n1479_0[0]),.dout(n1541),.clk(gclk));
	jand g1478(.dina(w_n1516_0[0]),.dinb(w_n1476_0[0]),.dout(n1542),.clk(gclk));
	jor g1479(.dina(n1542),.dinb(w_dff_B_CrfapjXi1_1),.dout(n1543),.clk(gclk));
	jand g1480(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1544),.clk(gclk));
	jnot g1481(.din(n1544),.dout(n1545),.clk(gclk));
	jand g1482(.dina(w_n1513_0[0]),.dinb(w_n1484_0[0]),.dout(n1546),.clk(gclk));
	jand g1483(.dina(w_n1514_0[0]),.dinb(w_n1481_0[0]),.dout(n1547),.clk(gclk));
	jor g1484(.dina(n1547),.dinb(w_dff_B_TkxqROVW5_1),.dout(n1548),.clk(gclk));
	jand g1485(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1549),.clk(gclk));
	jnot g1486(.din(n1549),.dout(n1550),.clk(gclk));
	jand g1487(.dina(w_n1511_0[0]),.dinb(w_n1489_0[0]),.dout(n1551),.clk(gclk));
	jand g1488(.dina(w_n1512_0[0]),.dinb(w_n1486_0[0]),.dout(n1552),.clk(gclk));
	jor g1489(.dina(n1552),.dinb(w_dff_B_Va8VTkjZ2_1),.dout(n1553),.clk(gclk));
	jand g1490(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1554),.clk(gclk));
	jnot g1491(.din(n1554),.dout(n1555),.clk(gclk));
	jand g1492(.dina(w_n1509_0[0]),.dinb(w_n1494_0[0]),.dout(n1556),.clk(gclk));
	jand g1493(.dina(w_n1510_0[0]),.dinb(w_n1491_0[0]),.dout(n1557),.clk(gclk));
	jor g1494(.dina(n1557),.dinb(w_dff_B_XibNqeFm6_1),.dout(n1558),.clk(gclk));
	jand g1495(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1559),.clk(gclk));
	jnot g1496(.din(n1559),.dout(n1560),.clk(gclk));
	jand g1497(.dina(w_n1507_0[0]),.dinb(w_n1499_0[0]),.dout(n1561),.clk(gclk));
	jand g1498(.dina(w_n1508_0[0]),.dinb(w_n1496_0[0]),.dout(n1562),.clk(gclk));
	jor g1499(.dina(n1562),.dinb(w_dff_B_yLu2oWlL0_1),.dout(n1563),.clk(gclk));
	jand g1500(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1564),.clk(gclk));
	jand g1501(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1565),.clk(gclk));
	jor g1502(.dina(w_n1504_0[0]),.dinb(w_n1501_0[0]),.dout(n1566),.clk(gclk));
	jor g1503(.dina(w_n1506_0[0]),.dinb(w_n1500_0[0]),.dout(n1567),.clk(gclk));
	jand g1504(.dina(n1567),.dinb(w_dff_B_akoQDKb85_1),.dout(n1568),.clk(gclk));
	jxor g1505(.dina(w_n1568_0[1]),.dinb(w_n1565_0[1]),.dout(n1569),.clk(gclk));
	jnot g1506(.din(n1569),.dout(n1570),.clk(gclk));
	jxor g1507(.dina(w_n1570_0[1]),.dinb(w_n1564_0[1]),.dout(n1571),.clk(gclk));
	jxor g1508(.dina(w_n1571_0[1]),.dinb(w_n1563_0[1]),.dout(n1572),.clk(gclk));
	jxor g1509(.dina(w_n1572_0[1]),.dinb(w_n1560_0[1]),.dout(n1573),.clk(gclk));
	jxor g1510(.dina(w_n1573_0[1]),.dinb(w_n1558_0[1]),.dout(n1574),.clk(gclk));
	jxor g1511(.dina(w_n1574_0[1]),.dinb(w_n1555_0[1]),.dout(n1575),.clk(gclk));
	jxor g1512(.dina(w_n1575_0[1]),.dinb(w_n1553_0[1]),.dout(n1576),.clk(gclk));
	jxor g1513(.dina(w_n1576_0[1]),.dinb(w_n1550_0[1]),.dout(n1577),.clk(gclk));
	jxor g1514(.dina(w_n1577_0[1]),.dinb(w_n1548_0[1]),.dout(n1578),.clk(gclk));
	jxor g1515(.dina(w_n1578_0[1]),.dinb(w_n1545_0[1]),.dout(n1579),.clk(gclk));
	jxor g1516(.dina(w_n1579_0[1]),.dinb(w_n1543_0[1]),.dout(n1580),.clk(gclk));
	jxor g1517(.dina(w_n1580_0[1]),.dinb(w_n1540_0[1]),.dout(n1581),.clk(gclk));
	jxor g1518(.dina(w_n1581_0[1]),.dinb(w_n1538_0[1]),.dout(n1582),.clk(gclk));
	jnot g1519(.din(n1582),.dout(n1583),.clk(gclk));
	jxor g1520(.dina(w_n1583_0[1]),.dinb(w_n1535_0[1]),.dout(n1584),.clk(gclk));
	jnot g1521(.din(n1584),.dout(n1585),.clk(gclk));
	jxor g1522(.dina(w_n1585_0[1]),.dinb(w_n1534_0[1]),.dout(n1586),.clk(gclk));
	jxor g1523(.dina(w_n1586_0[1]),.dinb(w_n1529_0[1]),.dout(w_dff_A_VdYZ4TDy2_2),.clk(gclk));
	jor g1524(.dina(w_n1585_0[0]),.dinb(w_n1534_0[0]),.dout(n1588),.clk(gclk));
	jnot g1525(.din(w_n1586_0[0]),.dout(n1589),.clk(gclk));
	jor g1526(.dina(w_dff_B_kMbvP8Ys0_0),.dinb(w_n1529_0[0]),.dout(n1590),.clk(gclk));
	jand g1527(.dina(n1590),.dinb(w_dff_B_YA4uxX2x2_1),.dout(n1591),.clk(gclk));
	jnot g1528(.din(w_n1538_0[0]),.dout(n1592),.clk(gclk));
	jnot g1529(.din(w_n1581_0[0]),.dout(n1593),.clk(gclk));
	jor g1530(.dina(w_dff_B_wztV4xSX0_0),.dinb(n1592),.dout(n1594),.clk(gclk));
	jor g1531(.dina(w_n1583_0[0]),.dinb(w_n1535_0[0]),.dout(n1595),.clk(gclk));
	jand g1532(.dina(n1595),.dinb(w_dff_B_9t040d6f3_1),.dout(n1596),.clk(gclk));
	jand g1533(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1597),.clk(gclk));
	jand g1534(.dina(w_n1579_0[0]),.dinb(w_n1543_0[0]),.dout(n1598),.clk(gclk));
	jand g1535(.dina(w_n1580_0[0]),.dinb(w_n1540_0[0]),.dout(n1599),.clk(gclk));
	jor g1536(.dina(n1599),.dinb(w_dff_B_ZnchbZUI3_1),.dout(n1600),.clk(gclk));
	jand g1537(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1601),.clk(gclk));
	jnot g1538(.din(n1601),.dout(n1602),.clk(gclk));
	jand g1539(.dina(w_n1577_0[0]),.dinb(w_n1548_0[0]),.dout(n1603),.clk(gclk));
	jand g1540(.dina(w_n1578_0[0]),.dinb(w_n1545_0[0]),.dout(n1604),.clk(gclk));
	jor g1541(.dina(n1604),.dinb(w_dff_B_PWGUw7d86_1),.dout(n1605),.clk(gclk));
	jand g1542(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1606),.clk(gclk));
	jnot g1543(.din(n1606),.dout(n1607),.clk(gclk));
	jand g1544(.dina(w_n1575_0[0]),.dinb(w_n1553_0[0]),.dout(n1608),.clk(gclk));
	jand g1545(.dina(w_n1576_0[0]),.dinb(w_n1550_0[0]),.dout(n1609),.clk(gclk));
	jor g1546(.dina(n1609),.dinb(w_dff_B_Jm8IZ2yX3_1),.dout(n1610),.clk(gclk));
	jand g1547(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1611),.clk(gclk));
	jnot g1548(.din(n1611),.dout(n1612),.clk(gclk));
	jand g1549(.dina(w_n1573_0[0]),.dinb(w_n1558_0[0]),.dout(n1613),.clk(gclk));
	jand g1550(.dina(w_n1574_0[0]),.dinb(w_n1555_0[0]),.dout(n1614),.clk(gclk));
	jor g1551(.dina(n1614),.dinb(w_dff_B_td0WxbKe1_1),.dout(n1615),.clk(gclk));
	jand g1552(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1616),.clk(gclk));
	jnot g1553(.din(n1616),.dout(n1617),.clk(gclk));
	jand g1554(.dina(w_n1571_0[0]),.dinb(w_n1563_0[0]),.dout(n1618),.clk(gclk));
	jand g1555(.dina(w_n1572_0[0]),.dinb(w_n1560_0[0]),.dout(n1619),.clk(gclk));
	jor g1556(.dina(n1619),.dinb(w_dff_B_lVfrHDpd8_1),.dout(n1620),.clk(gclk));
	jand g1557(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1621),.clk(gclk));
	jand g1558(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1622),.clk(gclk));
	jor g1559(.dina(w_n1568_0[0]),.dinb(w_n1565_0[0]),.dout(n1623),.clk(gclk));
	jor g1560(.dina(w_n1570_0[0]),.dinb(w_n1564_0[0]),.dout(n1624),.clk(gclk));
	jand g1561(.dina(n1624),.dinb(w_dff_B_CDUyJ6Ha0_1),.dout(n1625),.clk(gclk));
	jxor g1562(.dina(w_n1625_0[1]),.dinb(w_n1622_0[1]),.dout(n1626),.clk(gclk));
	jnot g1563(.din(n1626),.dout(n1627),.clk(gclk));
	jxor g1564(.dina(w_n1627_0[1]),.dinb(w_n1621_0[1]),.dout(n1628),.clk(gclk));
	jxor g1565(.dina(w_n1628_0[1]),.dinb(w_n1620_0[1]),.dout(n1629),.clk(gclk));
	jxor g1566(.dina(w_n1629_0[1]),.dinb(w_n1617_0[1]),.dout(n1630),.clk(gclk));
	jxor g1567(.dina(w_n1630_0[1]),.dinb(w_n1615_0[1]),.dout(n1631),.clk(gclk));
	jxor g1568(.dina(w_n1631_0[1]),.dinb(w_n1612_0[1]),.dout(n1632),.clk(gclk));
	jxor g1569(.dina(w_n1632_0[1]),.dinb(w_n1610_0[1]),.dout(n1633),.clk(gclk));
	jxor g1570(.dina(w_n1633_0[1]),.dinb(w_n1607_0[1]),.dout(n1634),.clk(gclk));
	jxor g1571(.dina(w_n1634_0[1]),.dinb(w_n1605_0[1]),.dout(n1635),.clk(gclk));
	jxor g1572(.dina(w_n1635_0[1]),.dinb(w_n1602_0[1]),.dout(n1636),.clk(gclk));
	jxor g1573(.dina(w_n1636_0[1]),.dinb(w_n1600_0[1]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jxor g1575(.dina(w_n1638_0[1]),.dinb(w_n1597_0[1]),.dout(n1639),.clk(gclk));
	jnot g1576(.din(n1639),.dout(n1640),.clk(gclk));
	jxor g1577(.dina(w_n1640_0[1]),.dinb(w_n1596_0[1]),.dout(n1641),.clk(gclk));
	jxor g1578(.dina(w_n1641_0[1]),.dinb(w_n1591_0[1]),.dout(w_dff_A_AlZA3pCn3_2),.clk(gclk));
	jor g1579(.dina(w_n1640_0[0]),.dinb(w_n1596_0[0]),.dout(n1643),.clk(gclk));
	jnot g1580(.din(w_n1641_0[0]),.dout(n1644),.clk(gclk));
	jor g1581(.dina(w_dff_B_0kya3YlB7_0),.dinb(w_n1591_0[0]),.dout(n1645),.clk(gclk));
	jand g1582(.dina(n1645),.dinb(w_dff_B_s5QX8V1B0_1),.dout(n1646),.clk(gclk));
	jnot g1583(.din(w_n1600_0[0]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(w_n1636_0[0]),.dout(n1648),.clk(gclk));
	jor g1585(.dina(n1648),.dinb(n1647),.dout(n1649),.clk(gclk));
	jor g1586(.dina(w_n1638_0[0]),.dinb(w_n1597_0[0]),.dout(n1650),.clk(gclk));
	jand g1587(.dina(n1650),.dinb(w_dff_B_SP1HpvoC3_1),.dout(n1651),.clk(gclk));
	jand g1588(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1652),.clk(gclk));
	jnot g1589(.din(n1652),.dout(n1653),.clk(gclk));
	jand g1590(.dina(w_n1634_0[0]),.dinb(w_n1605_0[0]),.dout(n1654),.clk(gclk));
	jand g1591(.dina(w_n1635_0[0]),.dinb(w_n1602_0[0]),.dout(n1655),.clk(gclk));
	jor g1592(.dina(n1655),.dinb(w_dff_B_Hda611ca5_1),.dout(n1656),.clk(gclk));
	jand g1593(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jand g1595(.dina(w_n1632_0[0]),.dinb(w_n1610_0[0]),.dout(n1659),.clk(gclk));
	jand g1596(.dina(w_n1633_0[0]),.dinb(w_n1607_0[0]),.dout(n1660),.clk(gclk));
	jor g1597(.dina(n1660),.dinb(w_dff_B_tJimsX8j4_1),.dout(n1661),.clk(gclk));
	jand g1598(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1662),.clk(gclk));
	jnot g1599(.din(n1662),.dout(n1663),.clk(gclk));
	jand g1600(.dina(w_n1630_0[0]),.dinb(w_n1615_0[0]),.dout(n1664),.clk(gclk));
	jand g1601(.dina(w_n1631_0[0]),.dinb(w_n1612_0[0]),.dout(n1665),.clk(gclk));
	jor g1602(.dina(n1665),.dinb(w_dff_B_uWD0VSwd7_1),.dout(n1666),.clk(gclk));
	jand g1603(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1667),.clk(gclk));
	jnot g1604(.din(n1667),.dout(n1668),.clk(gclk));
	jand g1605(.dina(w_n1628_0[0]),.dinb(w_n1620_0[0]),.dout(n1669),.clk(gclk));
	jand g1606(.dina(w_n1629_0[0]),.dinb(w_n1617_0[0]),.dout(n1670),.clk(gclk));
	jor g1607(.dina(n1670),.dinb(w_dff_B_ntwO1BtR6_1),.dout(n1671),.clk(gclk));
	jand g1608(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1672),.clk(gclk));
	jand g1609(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1673),.clk(gclk));
	jor g1610(.dina(w_n1625_0[0]),.dinb(w_n1622_0[0]),.dout(n1674),.clk(gclk));
	jor g1611(.dina(w_n1627_0[0]),.dinb(w_n1621_0[0]),.dout(n1675),.clk(gclk));
	jand g1612(.dina(n1675),.dinb(w_dff_B_BS5jlJis8_1),.dout(n1676),.clk(gclk));
	jxor g1613(.dina(w_n1676_0[1]),.dinb(w_n1673_0[1]),.dout(n1677),.clk(gclk));
	jnot g1614(.din(n1677),.dout(n1678),.clk(gclk));
	jxor g1615(.dina(w_n1678_0[1]),.dinb(w_n1672_0[1]),.dout(n1679),.clk(gclk));
	jxor g1616(.dina(w_n1679_0[1]),.dinb(w_n1671_0[1]),.dout(n1680),.clk(gclk));
	jxor g1617(.dina(w_n1680_0[1]),.dinb(w_n1668_0[1]),.dout(n1681),.clk(gclk));
	jxor g1618(.dina(w_n1681_0[1]),.dinb(w_n1666_0[1]),.dout(n1682),.clk(gclk));
	jxor g1619(.dina(w_n1682_0[1]),.dinb(w_n1663_0[1]),.dout(n1683),.clk(gclk));
	jxor g1620(.dina(w_n1683_0[1]),.dinb(w_n1661_0[1]),.dout(n1684),.clk(gclk));
	jxor g1621(.dina(w_n1684_0[1]),.dinb(w_n1658_0[1]),.dout(n1685),.clk(gclk));
	jxor g1622(.dina(w_n1685_0[1]),.dinb(w_n1656_0[1]),.dout(n1686),.clk(gclk));
	jxor g1623(.dina(w_n1686_0[1]),.dinb(w_n1653_0[1]),.dout(n1687),.clk(gclk));
	jnot g1624(.din(n1687),.dout(n1688),.clk(gclk));
	jxor g1625(.dina(w_n1688_0[1]),.dinb(w_n1651_0[1]),.dout(n1689),.clk(gclk));
	jxor g1626(.dina(w_n1689_0[1]),.dinb(w_n1646_0[1]),.dout(w_dff_A_x9YO84OD2_2),.clk(gclk));
	jor g1627(.dina(w_n1688_0[0]),.dinb(w_n1651_0[0]),.dout(n1691),.clk(gclk));
	jnot g1628(.din(w_n1689_0[0]),.dout(n1692),.clk(gclk));
	jor g1629(.dina(w_dff_B_F08mUVaJ1_0),.dinb(w_n1646_0[0]),.dout(n1693),.clk(gclk));
	jand g1630(.dina(n1693),.dinb(w_dff_B_DNx9ayef5_1),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1685_0[0]),.dinb(w_n1656_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1686_0[0]),.dinb(w_n1653_0[0]),.dout(n1696),.clk(gclk));
	jor g1633(.dina(n1696),.dinb(w_dff_B_EjhvP3lH5_1),.dout(n1697),.clk(gclk));
	jand g1634(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1683_0[0]),.dinb(w_n1661_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1684_0[0]),.dinb(w_n1658_0[0]),.dout(n1701),.clk(gclk));
	jor g1638(.dina(n1701),.dinb(w_dff_B_nqvQXrCN6_1),.dout(n1702),.clk(gclk));
	jand g1639(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1703),.clk(gclk));
	jnot g1640(.din(n1703),.dout(n1704),.clk(gclk));
	jand g1641(.dina(w_n1681_0[0]),.dinb(w_n1666_0[0]),.dout(n1705),.clk(gclk));
	jand g1642(.dina(w_n1682_0[0]),.dinb(w_n1663_0[0]),.dout(n1706),.clk(gclk));
	jor g1643(.dina(n1706),.dinb(w_dff_B_bKvMIyeU2_1),.dout(n1707),.clk(gclk));
	jand g1644(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jand g1646(.dina(w_n1679_0[0]),.dinb(w_n1671_0[0]),.dout(n1710),.clk(gclk));
	jand g1647(.dina(w_n1680_0[0]),.dinb(w_n1668_0[0]),.dout(n1711),.clk(gclk));
	jor g1648(.dina(n1711),.dinb(w_dff_B_RYVMzpN97_1),.dout(n1712),.clk(gclk));
	jand g1649(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1713),.clk(gclk));
	jand g1650(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1714),.clk(gclk));
	jor g1651(.dina(w_n1676_0[0]),.dinb(w_n1673_0[0]),.dout(n1715),.clk(gclk));
	jor g1652(.dina(w_n1678_0[0]),.dinb(w_n1672_0[0]),.dout(n1716),.clk(gclk));
	jand g1653(.dina(n1716),.dinb(w_dff_B_ongJG3EE9_1),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1714_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1713_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1712_0[1]),.dout(n1721),.clk(gclk));
	jxor g1658(.dina(w_n1721_0[1]),.dinb(w_n1709_0[1]),.dout(n1722),.clk(gclk));
	jxor g1659(.dina(w_n1722_0[1]),.dinb(w_n1707_0[1]),.dout(n1723),.clk(gclk));
	jxor g1660(.dina(w_n1723_0[1]),.dinb(w_n1704_0[1]),.dout(n1724),.clk(gclk));
	jxor g1661(.dina(w_n1724_0[1]),.dinb(w_n1702_0[1]),.dout(n1725),.clk(gclk));
	jxor g1662(.dina(w_n1725_0[1]),.dinb(w_n1699_0[1]),.dout(n1726),.clk(gclk));
	jxor g1663(.dina(w_n1726_0[1]),.dinb(w_n1697_0[1]),.dout(n1727),.clk(gclk));
	jxor g1664(.dina(w_n1727_0[1]),.dinb(w_n1694_0[1]),.dout(w_dff_A_YgTyAIea9_2),.clk(gclk));
	jnot g1665(.din(w_n1697_0[0]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(w_n1726_0[0]),.dout(n1730),.clk(gclk));
	jor g1667(.dina(n1730),.dinb(w_dff_B_RNmKnxNj1_1),.dout(n1731),.clk(gclk));
	jnot g1668(.din(w_n1727_0[0]),.dout(n1732),.clk(gclk));
	jor g1669(.dina(w_dff_B_DXgxM1M27_0),.dinb(w_n1694_0[0]),.dout(n1733),.clk(gclk));
	jand g1670(.dina(n1733),.dinb(w_dff_B_uDp8zjvm9_1),.dout(n1734),.clk(gclk));
	jand g1671(.dina(w_n1724_0[0]),.dinb(w_n1702_0[0]),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1725_0[0]),.dinb(w_n1699_0[0]),.dout(n1736),.clk(gclk));
	jor g1673(.dina(n1736),.dinb(w_dff_B_xxwiKctb7_1),.dout(n1737),.clk(gclk));
	jand g1674(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1738),.clk(gclk));
	jnot g1675(.din(n1738),.dout(n1739),.clk(gclk));
	jand g1676(.dina(w_n1722_0[0]),.dinb(w_n1707_0[0]),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1723_0[0]),.dinb(w_n1704_0[0]),.dout(n1741),.clk(gclk));
	jor g1678(.dina(n1741),.dinb(w_dff_B_Fwtz0GBI3_1),.dout(n1742),.clk(gclk));
	jand g1679(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1743),.clk(gclk));
	jnot g1680(.din(n1743),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_n1720_0[0]),.dinb(w_n1712_0[0]),.dout(n1745),.clk(gclk));
	jand g1682(.dina(w_n1721_0[0]),.dinb(w_n1709_0[0]),.dout(n1746),.clk(gclk));
	jor g1683(.dina(n1746),.dinb(w_dff_B_8w4XTPpi9_1),.dout(n1747),.clk(gclk));
	jand g1684(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1748),.clk(gclk));
	jand g1685(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1749),.clk(gclk));
	jor g1686(.dina(w_n1717_0[0]),.dinb(w_n1714_0[0]),.dout(n1750),.clk(gclk));
	jor g1687(.dina(w_n1719_0[0]),.dinb(w_n1713_0[0]),.dout(n1751),.clk(gclk));
	jand g1688(.dina(n1751),.dinb(w_dff_B_Eb1e4zv05_1),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1749_0[1]),.dout(n1753),.clk(gclk));
	jnot g1690(.din(n1753),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1748_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1747_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1744_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1742_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1739_0[1]),.dout(n1759),.clk(gclk));
	jxor g1696(.dina(w_n1759_0[1]),.dinb(w_n1737_0[1]),.dout(n1760),.clk(gclk));
	jxor g1697(.dina(w_n1760_0[1]),.dinb(w_n1734_0[1]),.dout(w_dff_A_1aNiPV9I1_2),.clk(gclk));
	jnot g1698(.din(w_n1737_0[0]),.dout(n1762),.clk(gclk));
	jnot g1699(.din(w_n1759_0[0]),.dout(n1763),.clk(gclk));
	jor g1700(.dina(n1763),.dinb(w_dff_B_v8v4A7LS1_1),.dout(n1764),.clk(gclk));
	jnot g1701(.din(w_n1760_0[0]),.dout(n1765),.clk(gclk));
	jor g1702(.dina(w_dff_B_rmZtcw0A2_0),.dinb(w_n1734_0[0]),.dout(n1766),.clk(gclk));
	jand g1703(.dina(n1766),.dinb(w_dff_B_LvUM34K53_1),.dout(n1767),.clk(gclk));
	jand g1704(.dina(w_n1757_0[0]),.dinb(w_n1742_0[0]),.dout(n1768),.clk(gclk));
	jand g1705(.dina(w_n1758_0[0]),.dinb(w_n1739_0[0]),.dout(n1769),.clk(gclk));
	jor g1706(.dina(n1769),.dinb(w_dff_B_FpK85Rv57_1),.dout(n1770),.clk(gclk));
	jand g1707(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1771),.clk(gclk));
	jnot g1708(.din(n1771),.dout(n1772),.clk(gclk));
	jand g1709(.dina(w_n1755_0[0]),.dinb(w_n1747_0[0]),.dout(n1773),.clk(gclk));
	jand g1710(.dina(w_n1756_0[0]),.dinb(w_n1744_0[0]),.dout(n1774),.clk(gclk));
	jor g1711(.dina(n1774),.dinb(w_dff_B_7dpaZHxq8_1),.dout(n1775),.clk(gclk));
	jand g1712(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1777),.clk(gclk));
	jor g1714(.dina(w_n1752_0[0]),.dinb(w_n1749_0[0]),.dout(n1778),.clk(gclk));
	jor g1715(.dina(w_n1754_0[0]),.dinb(w_n1748_0[0]),.dout(n1779),.clk(gclk));
	jand g1716(.dina(n1779),.dinb(w_dff_B_RZnj8RYO2_1),.dout(n1780),.clk(gclk));
	jxor g1717(.dina(w_n1780_0[1]),.dinb(w_n1777_0[1]),.dout(n1781),.clk(gclk));
	jnot g1718(.din(n1781),.dout(n1782),.clk(gclk));
	jxor g1719(.dina(w_n1782_0[1]),.dinb(w_n1776_0[1]),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1775_0[1]),.dout(n1784),.clk(gclk));
	jxor g1721(.dina(w_n1784_0[1]),.dinb(w_n1772_0[1]),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1770_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1767_0[1]),.dout(w_dff_A_xYpvdcGX7_2),.clk(gclk));
	jnot g1724(.din(w_n1770_0[0]),.dout(n1788),.clk(gclk));
	jnot g1725(.din(w_n1785_0[0]),.dout(n1789),.clk(gclk));
	jor g1726(.dina(n1789),.dinb(w_dff_B_ETaZKDi58_1),.dout(n1790),.clk(gclk));
	jnot g1727(.din(w_n1786_0[0]),.dout(n1791),.clk(gclk));
	jor g1728(.dina(w_dff_B_wTDV2G8q2_0),.dinb(w_n1767_0[0]),.dout(n1792),.clk(gclk));
	jand g1729(.dina(n1792),.dinb(w_dff_B_riXXVnAg6_1),.dout(n1793),.clk(gclk));
	jand g1730(.dina(w_n1783_0[0]),.dinb(w_n1775_0[0]),.dout(n1794),.clk(gclk));
	jand g1731(.dina(w_n1784_0[0]),.dinb(w_n1772_0[0]),.dout(n1795),.clk(gclk));
	jor g1732(.dina(n1795),.dinb(w_dff_B_wGgdgUrc1_1),.dout(n1796),.clk(gclk));
	jand g1733(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1797),.clk(gclk));
	jand g1734(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1798),.clk(gclk));
	jor g1735(.dina(w_n1780_0[0]),.dinb(w_n1777_0[0]),.dout(n1799),.clk(gclk));
	jor g1736(.dina(w_n1782_0[0]),.dinb(w_n1776_0[0]),.dout(n1800),.clk(gclk));
	jand g1737(.dina(n1800),.dinb(w_dff_B_SQb1nkqy3_1),.dout(n1801),.clk(gclk));
	jxor g1738(.dina(w_n1801_0[1]),.dinb(w_n1798_0[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jxor g1740(.dina(w_n1803_0[1]),.dinb(w_n1797_0[1]),.dout(n1804),.clk(gclk));
	jxor g1741(.dina(w_n1804_0[1]),.dinb(w_n1796_0[1]),.dout(n1805),.clk(gclk));
	jxor g1742(.dina(w_n1805_0[1]),.dinb(w_n1793_0[1]),.dout(w_dff_A_oBPVQzMN0_2),.clk(gclk));
	jand g1743(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1807),.clk(gclk));
	jor g1744(.dina(w_n1801_0[0]),.dinb(w_n1798_0[0]),.dout(n1808),.clk(gclk));
	jor g1745(.dina(w_n1803_0[0]),.dinb(w_n1797_0[0]),.dout(n1809),.clk(gclk));
	jand g1746(.dina(n1809),.dinb(w_dff_B_ZdHPZkjT0_1),.dout(n1810),.clk(gclk));
	jor g1747(.dina(w_n1810_0[1]),.dinb(w_n1807_0[1]),.dout(n1811),.clk(gclk));
	jnot g1748(.din(w_n1796_0[0]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(w_n1804_0[0]),.dout(n1813),.clk(gclk));
	jor g1750(.dina(n1813),.dinb(w_dff_B_jsicA2br8_1),.dout(n1814),.clk(gclk));
	jnot g1751(.din(w_n1805_0[0]),.dout(n1815),.clk(gclk));
	jor g1752(.dina(w_dff_B_0VGTcHsx1_0),.dinb(w_n1793_0[0]),.dout(n1816),.clk(gclk));
	jand g1753(.dina(n1816),.dinb(w_dff_B_Qw1tMa5V8_1),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1810_0[0]),.dinb(w_n1807_0[0]),.dout(n1818),.clk(gclk));
	jnot g1755(.din(w_n1818_0[1]),.dout(n1819),.clk(gclk));
	jor g1756(.dina(w_dff_B_u8BV5SUB4_0),.dinb(w_n1817_0[1]),.dout(n1820),.clk(gclk));
	jand g1757(.dina(n1820),.dinb(w_dff_B_phOQFaYs1_1),.dout(G6287gat),.clk(gclk));
	jxor g1758(.dina(w_n1818_0[0]),.dinb(w_n1817_0[0]),.dout(w_dff_A_i6yb8BNW4_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl jspl_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl jspl_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_G307gat_2[1]),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl jspl_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(w_dff_A_ooBIzX3Q9_1),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n66_0(.douta(w_dff_A_7PsyB8RX7_0),.doutb(w_n66_0[1]),.din(n66));
	jspl jspl_w_n67_0(.douta(w_n67_0[0]),.doutb(w_n67_0[1]),.din(w_dff_B_DaDNKJQD9_2));
	jspl jspl_w_n69_0(.douta(w_n69_0[0]),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n75_0(.douta(w_dff_A_QnJKV9jW3_0),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl3 jspl3_w_n80_0(.douta(w_dff_A_Xm4Ois8X2_0),.doutb(w_n80_0[1]),.doutc(w_n80_0[2]),.din(n80));
	jspl jspl_w_n83_0(.douta(w_n83_0[0]),.doutb(w_n83_0[1]),.din(n83));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n86_0(.douta(w_dff_A_d8DAIhbV2_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n90_0(.douta(w_n90_0[0]),.doutb(w_n90_0[1]),.din(n90));
	jspl jspl_w_n91_0(.douta(w_dff_A_ekScY5O94_0),.doutb(w_n91_0[1]),.din(n91));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_MSEJUAI97_1),.din(n103));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n106_0(.douta(w_dff_A_qdcJQ49M1_0),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl jspl_w_n112_0(.douta(w_dff_A_sLao2UcO5_0),.doutb(w_n112_0[1]),.din(n112));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_n117_0[1]),.doutc(w_n117_0[2]),.din(n117));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(w_dff_B_SKjCMl7v6_2));
	jspl jspl_w_n120_0(.douta(w_n120_0[0]),.doutb(w_n120_0[1]),.din(n120));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n122_0(.douta(w_dff_A_9ki8toQ61_0),.doutb(w_n122_0[1]),.din(n122));
	jspl jspl_w_n123_0(.douta(w_dff_A_tqDlP7NW9_0),.doutb(w_n123_0[1]),.din(n123));
	jspl jspl_w_n125_0(.douta(w_n125_0[0]),.doutb(w_n125_0[1]),.din(n125));
	jspl jspl_w_n127_0(.douta(w_n127_0[0]),.doutb(w_n127_0[1]),.din(n127));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(n128));
	jspl jspl_w_n129_0(.douta(w_dff_A_iQhZsTBv4_0),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.din(n130));
	jspl jspl_w_n132_0(.douta(w_n132_0[0]),.doutb(w_dff_A_hivLiakV5_1),.din(n132));
	jspl jspl_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.din(n133));
	jspl jspl_w_n135_0(.douta(w_dff_A_9WrAOST24_0),.doutb(w_n135_0[1]),.din(n135));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n141_0(.douta(w_dff_A_qETlHZLX2_0),.doutb(w_n141_0[1]),.din(n141));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.doutc(w_n146_0[2]),.din(n146));
	jspl jspl_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.din(w_dff_B_GKEotS8a1_2));
	jspl jspl_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(w_dff_B_xEacR6If5_2));
	jspl jspl_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.din(n155));
	jspl jspl_w_n156_0(.douta(w_dff_A_nGqydeaL0_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n157_0(.douta(w_dff_A_Rg6AGHtF7_0),.doutb(w_n157_0[1]),.din(n157));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(n158));
	jspl jspl_w_n160_0(.douta(w_n160_0[0]),.doutb(w_n160_0[1]),.din(n160));
	jspl jspl_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.din(n161));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(w_dff_B_3qcV8KCs4_2));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n164_0(.douta(w_dff_A_dgaDtayp4_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(n165));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_dff_A_RKyRjln93_1),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl jspl_w_n170_0(.douta(w_dff_A_3paX2inR4_0),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(n175));
	jspl jspl_w_n176_0(.douta(w_dff_A_rnaNxX3p0_0),.doutb(w_n176_0[1]),.din(n176));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl jspl_w_n183_0(.douta(w_n183_0[0]),.doutb(w_n183_0[1]),.din(w_dff_B_RQbxMgue5_2));
	jspl jspl_w_n186_0(.douta(w_n186_0[0]),.doutb(w_n186_0[1]),.din(n186));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(w_dff_B_8W3jZQuq6_2));
	jspl jspl_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.din(n192));
	jspl jspl_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.din(w_dff_B_5j9PqDcD1_2));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_dff_A_JUhNNVgm0_0),.doutb(w_dff_A_ZLkAxtuN9_1),.doutc(w_n196_0[2]),.din(n196));
	jspl jspl_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.din(w_dff_B_iUG0sUcw6_2));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(n203));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(w_dff_B_YSaWgmih5_2));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(n205));
	jspl jspl_w_n206_0(.douta(w_dff_A_l1YxZAyV9_0),.doutb(w_n206_0[1]),.din(n206));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_dff_A_2h6ak3GK4_1),.din(n209));
	jspl jspl_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.din(n210));
	jspl jspl_w_n212_0(.douta(w_dff_A_nXyfF5ZW7_0),.doutb(w_n212_0[1]),.din(n212));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_dff_A_XSkiOj6b1_0),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.doutc(w_n223_0[2]),.din(n223));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(w_dff_B_lpY4cnop9_2));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.din(w_dff_B_B1atzNu17_2));
	jspl jspl_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.din(n233));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_n235_0[1]),.din(w_dff_B_7mP3ZrFy4_2));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(n239));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(w_dff_B_DPQAd0JT2_2));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_dff_A_HYTriE2r8_0),.doutb(w_dff_A_y8ecDZvJ4_1),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n248_0(.douta(w_n248_0[0]),.doutb(w_n248_0[1]),.din(n248));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_6moYWDCl8_2));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl jspl_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.din(w_dff_B_nxiq51Ud2_2));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl jspl_w_n253_0(.douta(w_n253_0[0]),.doutb(w_n253_0[1]),.din(w_dff_B_u8z9iEiN3_2));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n255_0(.douta(w_dff_A_ZTA4c5vr1_0),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n256_0(.douta(w_n256_0[0]),.doutb(w_n256_0[1]),.din(n256));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_dff_A_ujIduFVv2_1),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_dff_A_gM2LXppr0_0),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_dff_A_8jxZBe6x3_0),.doutb(w_n267_0[1]),.din(n267));
	jspl3 jspl3_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.doutc(w_n272_0[2]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(w_dff_B_n0acGMyX6_2));
	jspl jspl_w_n277_0(.douta(w_n277_0[0]),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(w_dff_B_lBNBFkrK6_2));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n284_0(.douta(w_n284_0[0]),.doutb(w_n284_0[1]),.din(w_dff_B_CbvTIG0O8_2));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl jspl_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.din(w_dff_B_EZJuavUv4_2));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(w_dff_B_muOGxhGJ0_2));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl3 jspl3_w_n297_0(.douta(w_dff_A_nqIjHJqT2_0),.doutb(w_dff_A_g1Mpap7a6_1),.doutc(w_n297_0[2]),.din(n297));
	jspl jspl_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.din(n299));
	jspl jspl_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.din(n301));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_n302_0[1]),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(w_dff_B_KrkZHRZ11_2));
	jspl jspl_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.din(n304));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(w_dff_B_n3Z6e0v41_2));
	jspl jspl_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.din(n306));
	jspl jspl_w_n307_0(.douta(w_n307_0[0]),.doutb(w_n307_0[1]),.din(w_dff_B_LAmdmyhz3_2));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(w_dff_B_MdHYQ9QH5_2));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(n310));
	jspl jspl_w_n311_0(.douta(w_dff_A_Fuhz5ZBN3_0),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.din(n312));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_dff_A_E2AfKQGi1_1),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_dff_A_9otDpVqf0_0),.doutb(w_n317_0[1]),.din(n317));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_dff_A_6pazhalA8_0),.doutb(w_n323_0[1]),.din(n323));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(w_dff_B_GcmFsTjW1_2));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.din(w_dff_B_ZMuS2v2G9_2));
	jspl jspl_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.din(n338));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(w_dff_B_b8fAa6Jb0_2));
	jspl jspl_w_n343_0(.douta(w_n343_0[0]),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(w_dff_B_9RkqwVp20_2));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(w_dff_B_lM87nnUQ3_2));
	jspl jspl_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.din(n354));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(w_dff_B_E4u52Zoz7_2));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl3 jspl3_w_n358_0(.douta(w_dff_A_DeY9akHJ1_0),.doutb(w_dff_A_ae8Leg8q5_1),.doutc(w_n358_0[2]),.din(n358));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(n363));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(w_dff_B_yrwF1j462_2));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_n365_0[1]),.din(n365));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(w_dff_B_D35Bkf912_2));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(w_dff_B_IE4fTbbZ3_2));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(w_dff_B_6WoNTM9e2_2));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(w_dff_B_hTY2G8Qz6_2));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n374_0(.douta(w_dff_A_GwuSQdzy9_0),.doutb(w_n374_0[1]),.din(n374));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_dff_A_RVsGh9gK2_1),.din(n377));
	jspl jspl_w_n378_0(.douta(w_n378_0[0]),.doutb(w_n378_0[1]),.din(n378));
	jspl jspl_w_n380_0(.douta(w_dff_A_8REIYbrZ2_0),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl jspl_w_n386_0(.douta(w_dff_A_b6WhIoFW7_0),.doutb(w_n386_0[1]),.din(n386));
	jspl3 jspl3_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.doutc(w_n391_0[2]),.din(n391));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(w_dff_B_ym3Zhri70_2));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.din(n396));
	jspl jspl_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.din(w_dff_B_mLPwvyRw6_2));
	jspl jspl_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.din(n401));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(w_dff_B_xobzKttg0_2));
	jspl jspl_w_n406_0(.douta(w_n406_0[0]),.doutb(w_n406_0[1]),.din(n406));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(w_dff_B_hhHb4CZS5_2));
	jspl jspl_w_n411_0(.douta(w_n411_0[0]),.doutb(w_n411_0[1]),.din(n411));
	jspl jspl_w_n413_0(.douta(w_n413_0[0]),.doutb(w_n413_0[1]),.din(w_dff_B_s9XxNWqf5_2));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(w_dff_B_L38jzCHb3_2));
	jspl jspl_w_n418_0(.douta(w_n418_0[0]),.doutb(w_n418_0[1]),.din(w_dff_B_3M5uY5Tr9_2));
	jspl jspl_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.din(n423));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(w_dff_B_zDriRcux5_2));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl3 jspl3_w_n427_0(.douta(w_dff_A_qgqYeQLl3_0),.doutb(w_dff_A_qSqHHLZm1_1),.doutc(w_n427_0[2]),.din(n427));
	jspl jspl_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.din(n429));
	jspl jspl_w_n431_0(.douta(w_n431_0[0]),.doutb(w_n431_0[1]),.din(n431));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(n432));
	jspl jspl_w_n433_0(.douta(w_n433_0[0]),.doutb(w_n433_0[1]),.din(w_dff_B_mS9zbmyi8_2));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl jspl_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.din(n436));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(n437));
	jspl jspl_w_n438_0(.douta(w_n438_0[0]),.doutb(w_n438_0[1]),.din(n438));
	jspl jspl_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.din(w_dff_B_Ef1UaLVG5_2));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(w_dff_B_XQlWpnvd2_2));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_n442_0[1]),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(w_dff_B_zx4XBNOA8_2));
	jspl jspl_w_n444_0(.douta(w_n444_0[0]),.doutb(w_n444_0[1]),.din(n444));
	jspl jspl_w_n445_0(.douta(w_dff_A_ssjJfwfn8_0),.doutb(w_n445_0[1]),.din(n445));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_dff_A_DkEdws1O4_1),.din(n448));
	jspl jspl_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.din(n449));
	jspl jspl_w_n451_0(.douta(w_dff_A_KESIRdKO2_0),.doutb(w_n451_0[1]),.din(n451));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_dff_A_yRb039tD0_0),.doutb(w_n457_0[1]),.din(n457));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(w_dff_B_qarWrr7Y9_2));
	jspl jspl_w_n467_0(.douta(w_n467_0[0]),.doutb(w_n467_0[1]),.din(n467));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(w_dff_B_VqpNoIgB5_2));
	jspl jspl_w_n472_0(.douta(w_n472_0[0]),.doutb(w_n472_0[1]),.din(n472));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(w_dff_B_oIoefvFy9_2));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(w_dff_B_L4ZbzIDi7_2));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(w_dff_B_fkV0tacZ9_2));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(w_dff_B_T7hkcrGP2_2));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(w_dff_B_JDMQXHZZ1_2));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(n499));
	jspl jspl_w_n501_0(.douta(w_n501_0[0]),.doutb(w_n501_0[1]),.din(w_dff_B_wPhdDcjg4_2));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl3 jspl3_w_n503_0(.douta(w_dff_A_W0GH72gf8_0),.doutb(w_dff_A_7j3bc8678_1),.doutc(w_n503_0[2]),.din(n503));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_CHBlmuDm5_2));
	jspl jspl_w_n510_0(.douta(w_n510_0[0]),.doutb(w_n510_0[1]),.din(n510));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(w_dff_B_KbVs6OG40_2));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n513_0(.douta(w_n513_0[0]),.doutb(w_n513_0[1]),.din(n513));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(n514));
	jspl jspl_w_n515_0(.douta(w_n515_0[0]),.doutb(w_n515_0[1]),.din(n515));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(w_dff_B_nZJmTAnu1_2));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(w_dff_B_zFtsBFuG7_2));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n521_0(.douta(w_n521_0[0]),.doutb(w_n521_0[1]),.din(w_dff_B_4CbSZ5vX4_2));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl jspl_w_n523_0(.douta(w_dff_A_TVcECwO33_0),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n526_0(.douta(w_n526_0[0]),.doutb(w_dff_A_lHvD8GlN0_1),.din(n526));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_dff_A_8FMft7rY4_0),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_dff_A_QnXpZbch3_0),.doutb(w_n535_0[1]),.din(n535));
	jspl3 jspl3_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.doutc(w_n540_0[2]),.din(n540));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(w_dff_B_vAR6gnbU2_2));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(w_dff_B_0cTUdrvL2_2));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.din(w_dff_B_QQcdNQza5_2));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(w_dff_B_5g0nQWiE2_2));
	jspl jspl_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.din(n560));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(w_dff_B_HmOy9gdZ6_2));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(w_dff_B_MuPLUmnB9_2));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl jspl_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.din(w_dff_B_CtZDk9d71_2));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(w_dff_B_fFbYDQIW4_2));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(w_dff_B_neDSvnNh6_2));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n586_0(.douta(w_dff_A_jYzDXLF64_0),.doutb(w_dff_A_Px009JHl6_1),.doutc(w_n586_0[2]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(n588));
	jspl jspl_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.din(n590));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(w_dff_B_nCxF0Fs43_2));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl jspl_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.din(w_dff_B_uXYkKBb94_2));
	jspl jspl_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.din(n595));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(w_dff_B_8FZDh62H1_2));
	jspl jspl_w_n597_0(.douta(w_n597_0[0]),.doutb(w_n597_0[1]),.din(n597));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl jspl_w_n599_0(.douta(w_n599_0[0]),.doutb(w_n599_0[1]),.din(n599));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(n600));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(w_dff_B_lgr9fuJH8_2));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(w_dff_B_zTSUf4yg2_2));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(w_dff_B_SQ2UFCHO7_2));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_dff_A_YThLcJGt7_0),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.din(n609));
	jspl jspl_w_n611_0(.douta(w_n611_0[0]),.doutb(w_dff_A_VCBWiqrM6_1),.din(n611));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl jspl_w_n614_0(.douta(w_dff_A_kXtpBZXi8_0),.doutb(w_n614_0[1]),.din(n614));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_dff_A_KIQ1Xrxm6_0),.doutb(w_n620_0[1]),.din(n620));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(w_dff_B_uCo2WFDQ7_2));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(w_dff_B_VjjXjdD76_2));
	jspl jspl_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.din(n635));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(w_dff_B_96dG2lku2_2));
	jspl jspl_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.din(n640));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(w_dff_B_5qY27qCF0_2));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(w_dff_B_i37JVgK58_2));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(w_dff_B_1HcQjVsl8_2));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(w_dff_B_cutxkZDZ0_2));
	jspl jspl_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.din(n660));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(w_dff_B_kjssqN031_2));
	jspl jspl_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.din(n665));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(w_dff_B_an79LytC2_2));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(w_dff_B_nKqnNbB13_2));
	jspl jspl_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.din(n675));
	jspl3 jspl3_w_n676_0(.douta(w_dff_A_96WjFtJZ9_0),.doutb(w_dff_A_z1Kp4bwm6_1),.doutc(w_n676_0[2]),.din(n676));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl jspl_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.din(n681));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(w_dff_B_TtyaOiSh6_2));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(w_dff_B_R87REC4W0_2));
	jspl jspl_w_n685_0(.douta(w_n685_0[0]),.doutb(w_n685_0[1]),.din(n685));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(w_dff_B_1OLi2jHj4_2));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n688_0(.douta(w_n688_0[0]),.doutb(w_n688_0[1]),.din(w_dff_B_aKw7mzUM2_2));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n691_0(.douta(w_n691_0[0]),.doutb(w_n691_0[1]),.din(n691));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.din(n692));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_n694_0[1]),.din(w_dff_B_uPSobetU8_2));
	jspl jspl_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.din(n695));
	jspl jspl_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.din(w_dff_B_aBR7h1Hy2_2));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(w_dff_B_BpsdmnhP5_2));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n700_0(.douta(w_dff_A_D4J8BljM6_0),.doutb(w_n700_0[1]),.din(n700));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_dff_A_CSAuEfHm7_1),.din(n703));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n706_0(.douta(w_dff_A_JDpPRqDB1_0),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_dff_A_MZQj5o8y5_0),.doutb(w_n712_0[1]),.din(n712));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.doutc(w_n717_0[2]),.din(n717));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(w_dff_B_LMMTeiyX9_2));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(w_dff_B_2FHoCyLs4_2));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.din(w_dff_B_hrcXJnDK9_2));
	jspl jspl_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.din(n732));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(w_dff_B_oRp3NQyX5_2));
	jspl jspl_w_n737_0(.douta(w_n737_0[0]),.doutb(w_n737_0[1]),.din(n737));
	jspl jspl_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.din(w_dff_B_cBGvdRqR1_2));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl jspl_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.din(w_dff_B_YF5CjkL67_2));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(n747));
	jspl jspl_w_n749_0(.douta(w_n749_0[0]),.doutb(w_n749_0[1]),.din(w_dff_B_e8OA1mjm3_2));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(w_dff_B_vtGoz9zg2_2));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(w_dff_B_kkq1ZYEO4_2));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(n762));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(w_dff_B_mnqJR6yD3_2));
	jspl jspl_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.din(n769));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(w_dff_B_wYrutqXZ8_2));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl jspl_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.din(n774));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(n777));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.din(w_dff_B_Ol1vyf5o2_2));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.din(w_dff_B_lqGQoYfm1_2));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl jspl_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.din(w_dff_B_GvEQLVg08_2));
	jspl jspl_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.din(n784));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(w_dff_B_1fONnGMT0_2));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_XofydX4J3_2));
	jspl jspl_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.din(n788));
	jspl jspl_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.din(n789));
	jspl jspl_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.din(n790));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl jspl_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.din(w_dff_B_svrYkw6u9_2));
	jspl jspl_w_n794_0(.douta(w_n794_0[0]),.doutb(w_n794_0[1]),.din(n794));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(w_dff_B_9RmJStxt8_2));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl jspl_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.din(w_dff_B_ah10LIvS1_2));
	jspl jspl_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.din(n798));
	jspl jspl_w_n799_0(.douta(w_dff_A_ZPHxKH3L7_0),.doutb(w_n799_0[1]),.din(n799));
	jspl jspl_w_n800_0(.douta(w_n800_0[0]),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_dff_A_7y1XPP7Z4_1),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(n803));
	jspl jspl_w_n805_0(.douta(w_dff_A_gsQw3Cox5_0),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(w_dff_B_GjiEG68z4_2));
	jspl jspl_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_dff_A_B8itLeCq2_0),.doutb(w_n816_0[1]),.din(n816));
	jspl3 jspl3_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.doutc(w_n820_0[2]),.din(n820));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(w_dff_B_3JPXeLls3_2));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(w_dff_B_QxodiXm21_2));
	jspl jspl_w_n830_0(.douta(w_n830_0[0]),.doutb(w_n830_0[1]),.din(n830));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(w_dff_B_0jYhmeDR2_2));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(n835));
	jspl jspl_w_n837_0(.douta(w_n837_0[0]),.doutb(w_n837_0[1]),.din(w_dff_B_M7snh6mM0_2));
	jspl jspl_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.din(n840));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(w_dff_B_WtYEZnw26_2));
	jspl jspl_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.din(n845));
	jspl jspl_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.din(w_dff_B_Az5yo4cW8_2));
	jspl jspl_w_n850_0(.douta(w_n850_0[0]),.doutb(w_n850_0[1]),.din(n850));
	jspl jspl_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.din(w_dff_B_atvicVez0_2));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(w_dff_B_FZkZf7sr3_2));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(w_dff_B_5scgfOcd7_2));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.din(n865));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(w_dff_B_EXMcD6pc9_2));
	jspl jspl_w_n872_0(.douta(w_n872_0[0]),.doutb(w_n872_0[1]),.din(n872));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(w_dff_B_Q2iIP7Qg7_2));
	jspl jspl_w_n875_0(.douta(w_dff_A_BkdLtBcM6_0),.doutb(w_n875_0[1]),.din(n875));
	jspl jspl_w_n877_0(.douta(w_dff_A_cs9E2wFq9_0),.doutb(w_n877_0[1]),.din(w_dff_B_2jQ3RK4d0_2));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n880_0(.douta(w_n880_0[0]),.doutb(w_n880_0[1]),.din(w_dff_B_5wJlXDlD9_2));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n882_0(.douta(w_n882_0[0]),.doutb(w_n882_0[1]),.din(w_dff_B_uELAWVEd5_2));
	jspl jspl_w_n883_0(.douta(w_n883_0[0]),.doutb(w_n883_0[1]),.din(n883));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(w_dff_B_KTLbZe9Y4_2));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(w_dff_B_q9E9E1EZ5_2));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.din(n887));
	jspl jspl_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.din(w_dff_B_kPyJZvli6_2));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n890_0(.douta(w_n890_0[0]),.doutb(w_n890_0[1]),.din(w_dff_B_DI2KDhzz3_2));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(n891));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n893_0(.douta(w_n893_0[0]),.doutb(w_n893_0[1]),.din(n893));
	jspl jspl_w_n894_0(.douta(w_n894_0[0]),.doutb(w_n894_0[1]),.din(n894));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(w_dff_B_J1SboDT76_2));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(w_dff_B_8iCog5Rp9_2));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.din(n899));
	jspl3 jspl3_w_n900_0(.douta(w_n900_0[0]),.doutb(w_dff_A_Pt0afR317_1),.doutc(w_dff_A_0aocDaWj8_2),.din(n900));
	jspl jspl_w_n902_0(.douta(w_n902_0[0]),.doutb(w_dff_A_pk5fm7722_1),.din(n902));
	jspl jspl_w_n903_0(.douta(w_n903_0[0]),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n904_0(.douta(w_n904_0[0]),.doutb(w_dff_A_MK0VuhU15_1),.din(n904));
	jspl jspl_w_n905_0(.douta(w_n905_0[0]),.doutb(w_n905_0[1]),.din(n905));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(n910));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(w_dff_B_npU4dBmU0_2));
	jspl3 jspl3_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.doutc(w_n915_0[2]),.din(n915));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(w_dff_B_GiPGGvU81_2));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(w_dff_B_tA00dRxH2_2));
	jspl jspl_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(w_dff_B_UrvDxQ9U4_2));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n934_0(.douta(w_n934_0[0]),.doutb(w_n934_0[1]),.din(w_dff_B_8BHbKbWp9_2));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n939_0(.douta(w_n939_0[0]),.doutb(w_n939_0[1]),.din(w_dff_B_guKhFquV9_2));
	jspl jspl_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.din(n942));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_n944_0[1]),.din(w_dff_B_YADlhlg21_2));
	jspl jspl_w_n947_0(.douta(w_n947_0[0]),.doutb(w_n947_0[1]),.din(n947));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(w_dff_B_ezzIuTk95_2));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(w_dff_B_d4nEiHRz9_2));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(w_dff_B_d7RAo6mC7_2));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(w_dff_B_UUS9ub6Q8_2));
	jspl jspl_w_n967_0(.douta(w_n967_0[0]),.doutb(w_n967_0[1]),.din(n967));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(w_dff_B_jri7Ub2C6_2));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(w_dff_B_mRin9tCy3_2));
	jspl jspl_w_n978_0(.douta(w_n978_0[0]),.doutb(w_n978_0[1]),.din(n978));
	jspl jspl_w_n980_0(.douta(w_dff_A_UX8pD6aF4_0),.doutb(w_n980_0[1]),.din(w_dff_B_mbQs6htz1_2));
	jspl jspl_w_n982_0(.douta(w_n982_0[0]),.doutb(w_n982_0[1]),.din(n982));
	jspl jspl_w_n983_0(.douta(w_n983_0[0]),.doutb(w_n983_0[1]),.din(w_dff_B_gOT3hRON5_2));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(w_dff_B_GaJSvwO06_2));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(w_dff_B_KpAjid0A5_2));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl jspl_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.din(w_dff_B_HTmzlJ4h1_2));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.din(w_dff_B_6ZVNhIwl0_2));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(w_dff_B_aoIjgNAi7_2));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(w_dff_B_5zjqFYag2_2));
	jspl jspl_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.din(n995));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(w_dff_B_hc93bl1r7_2));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl jspl_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_n1002_0[1]),.din(w_dff_B_WAhhwlNj0_2));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.din(w_dff_B_zPu8CIsz0_2));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_dff_A_hYbFF23a1_1),.din(n1006));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_dff_A_4srhdI5f7_0),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(w_dff_B_gC9Kk4D31_2));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_dff_A_4Ncw3g6H8_1),.din(n1013));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(w_dff_B_5NNsqtcs0_2));
	jspl jspl_w_n1022_0(.douta(w_dff_A_jtq9VIji0_0),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(w_dff_B_zeGKJ73x9_2));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(w_dff_B_DZtWG4YR4_2));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(w_dff_B_lQyCJl4Y6_2));
	jspl jspl_w_n1036_0(.douta(w_n1036_0[0]),.doutb(w_n1036_0[1]),.din(n1036));
	jspl jspl_w_n1038_0(.douta(w_n1038_0[0]),.doutb(w_n1038_0[1]),.din(w_dff_B_rid0auL54_2));
	jspl jspl_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.din(n1041));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(w_dff_B_Y4ySdTZE1_2));
	jspl jspl_w_n1046_0(.douta(w_n1046_0[0]),.doutb(w_n1046_0[1]),.din(n1046));
	jspl jspl_w_n1048_0(.douta(w_n1048_0[0]),.doutb(w_n1048_0[1]),.din(w_dff_B_bqaJiNvs7_2));
	jspl jspl_w_n1051_0(.douta(w_n1051_0[0]),.doutb(w_n1051_0[1]),.din(n1051));
	jspl jspl_w_n1053_0(.douta(w_n1053_0[0]),.doutb(w_n1053_0[1]),.din(w_dff_B_ao91obDv1_2));
	jspl jspl_w_n1056_0(.douta(w_n1056_0[0]),.doutb(w_n1056_0[1]),.din(n1056));
	jspl jspl_w_n1058_0(.douta(w_n1058_0[0]),.doutb(w_n1058_0[1]),.din(w_dff_B_aeK2CoD29_2));
	jspl jspl_w_n1061_0(.douta(w_n1061_0[0]),.doutb(w_n1061_0[1]),.din(n1061));
	jspl jspl_w_n1063_0(.douta(w_n1063_0[0]),.doutb(w_n1063_0[1]),.din(w_dff_B_lyy5Ss3G8_2));
	jspl jspl_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.din(n1066));
	jspl jspl_w_n1068_0(.douta(w_n1068_0[0]),.doutb(w_n1068_0[1]),.din(w_dff_B_PrtgEQao9_2));
	jspl jspl_w_n1071_0(.douta(w_n1071_0[0]),.doutb(w_n1071_0[1]),.din(n1071));
	jspl jspl_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.din(w_dff_B_REPYmE8F0_2));
	jspl jspl_w_n1076_0(.douta(w_n1076_0[0]),.doutb(w_n1076_0[1]),.din(n1076));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(w_dff_B_WKGtY2ml4_2));
	jspl jspl_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.din(w_dff_B_XKFgzDIA2_2));
	jspl jspl_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.din(n1080));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl jspl_w_n1083_0(.douta(w_n1083_0[0]),.doutb(w_n1083_0[1]),.din(w_dff_B_VcfgjPsI0_2));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(n1084));
	jspl jspl_w_n1085_0(.douta(w_n1085_0[0]),.doutb(w_n1085_0[1]),.din(w_dff_B_4OQ3Tr7o3_2));
	jspl jspl_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.din(n1086));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(w_dff_B_werfbEQm9_2));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(w_dff_B_642m3ZPH9_2));
	jspl jspl_w_n1090_0(.douta(w_n1090_0[0]),.doutb(w_n1090_0[1]),.din(n1090));
	jspl jspl_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.din(w_dff_B_4xpjW6mv9_2));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1093_0(.douta(w_n1093_0[0]),.doutb(w_n1093_0[1]),.din(w_dff_B_X5KODBcQ8_2));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(n1094));
	jspl jspl_w_n1095_0(.douta(w_n1095_0[0]),.doutb(w_n1095_0[1]),.din(w_dff_B_Y6GAW0cI0_2));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1098_0(.douta(w_n1098_0[0]),.doutb(w_n1098_0[1]),.din(n1098));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(n1099));
	jspl jspl_w_n1100_0(.douta(w_n1100_0[0]),.doutb(w_n1100_0[1]),.din(n1100));
	jspl jspl_w_n1101_0(.douta(w_n1101_0[0]),.doutb(w_n1101_0[1]),.din(w_dff_B_b33kYsUA6_2));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(w_dff_B_SP7NRKBw2_2));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.din(n1105));
	jspl jspl_w_n1106_0(.douta(w_n1106_0[0]),.doutb(w_n1106_0[1]),.din(n1106));
	jspl jspl_w_n1107_0(.douta(w_n1107_0[0]),.doutb(w_n1107_0[1]),.din(n1107));
	jspl jspl_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_dff_A_g7Cqca0B3_1),.din(n1108));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1119_0(.douta(w_dff_A_MTFXj9jv8_0),.doutb(w_n1119_0[1]),.din(w_dff_B_TE7IUzHw6_2));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(w_dff_B_k6qpMpUd0_2));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(w_dff_B_e1hx0Z8G3_2));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(w_dff_B_J3NOWJQd2_2));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1136_0(.douta(w_n1136_0[0]),.doutb(w_n1136_0[1]),.din(w_dff_B_mhXbmUcO0_2));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(w_dff_B_YzDpsTeH8_2));
	jspl jspl_w_n1144_0(.douta(w_n1144_0[0]),.doutb(w_n1144_0[1]),.din(n1144));
	jspl jspl_w_n1146_0(.douta(w_n1146_0[0]),.doutb(w_n1146_0[1]),.din(w_dff_B_kzrcoXMJ4_2));
	jspl jspl_w_n1149_0(.douta(w_n1149_0[0]),.doutb(w_n1149_0[1]),.din(n1149));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(w_dff_B_lGtpcAJp7_2));
	jspl jspl_w_n1154_0(.douta(w_n1154_0[0]),.doutb(w_n1154_0[1]),.din(n1154));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(w_dff_B_fFzEiE7X7_2));
	jspl jspl_w_n1159_0(.douta(w_n1159_0[0]),.doutb(w_n1159_0[1]),.din(n1159));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(w_dff_B_KiwMMxOK1_2));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_n1164_0[1]),.din(n1164));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(w_dff_B_AdX8cphv6_2));
	jspl jspl_w_n1169_0(.douta(w_n1169_0[0]),.doutb(w_n1169_0[1]),.din(n1169));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(w_dff_B_7AgCoNZE4_2));
	jspl jspl_w_n1174_0(.douta(w_n1174_0[0]),.doutb(w_n1174_0[1]),.din(n1174));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_n1175_0[1]),.din(w_dff_B_WfUqXEjd0_2));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(w_dff_B_Wjv0KT8C0_2));
	jspl jspl_w_n1179_0(.douta(w_n1179_0[0]),.doutb(w_n1179_0[1]),.din(n1179));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1182_0(.douta(w_n1182_0[0]),.doutb(w_n1182_0[1]),.din(w_dff_B_RkzEbBhT9_2));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_n1184_0[0]),.doutb(w_n1184_0[1]),.din(w_dff_B_pDsZakwK6_2));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(w_dff_B_0SMno3DD3_2));
	jspl jspl_w_n1187_0(.douta(w_n1187_0[0]),.doutb(w_n1187_0[1]),.din(n1187));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(w_dff_B_gVfB6OuJ0_2));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1190_0(.douta(w_n1190_0[0]),.doutb(w_n1190_0[1]),.din(w_dff_B_03qnLCe22_2));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(n1191));
	jspl jspl_w_n1192_0(.douta(w_n1192_0[0]),.doutb(w_n1192_0[1]),.din(w_dff_B_agDZGcgb0_2));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(n1193));
	jspl jspl_w_n1194_0(.douta(w_n1194_0[0]),.doutb(w_n1194_0[1]),.din(w_dff_B_mToJob0I8_2));
	jspl jspl_w_n1195_0(.douta(w_n1195_0[0]),.doutb(w_n1195_0[1]),.din(n1195));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.din(n1197));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(n1198));
	jspl jspl_w_n1199_0(.douta(w_n1199_0[0]),.doutb(w_n1199_0[1]),.din(n1199));
	jspl jspl_w_n1200_0(.douta(w_n1200_0[0]),.doutb(w_n1200_0[1]),.din(w_dff_B_xyI3tAO59_2));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(w_dff_B_5rgbaAfY4_2));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(n1206));
	jspl jspl_w_n1207_0(.douta(w_dff_A_fRkJO1mJ1_0),.doutb(w_n1207_0[1]),.din(n1207));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(w_dff_B_8NRw3rHp5_2));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(w_dff_B_39RFgBUm3_2));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(n1225));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(w_dff_B_d8wm2tPJ1_2));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(w_dff_B_Gs5q38Ow6_2));
	jspl jspl_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.din(n1235));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(w_dff_B_61PhXr827_2));
	jspl jspl_w_n1240_0(.douta(w_n1240_0[0]),.doutb(w_n1240_0[1]),.din(n1240));
	jspl jspl_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.din(w_dff_B_udHESU6A9_2));
	jspl jspl_w_n1245_0(.douta(w_n1245_0[0]),.doutb(w_n1245_0[1]),.din(n1245));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(w_dff_B_Z2H3KzTz3_2));
	jspl jspl_w_n1250_0(.douta(w_n1250_0[0]),.doutb(w_n1250_0[1]),.din(n1250));
	jspl jspl_w_n1252_0(.douta(w_n1252_0[0]),.doutb(w_n1252_0[1]),.din(w_dff_B_im5OGiDU0_2));
	jspl jspl_w_n1255_0(.douta(w_n1255_0[0]),.doutb(w_n1255_0[1]),.din(n1255));
	jspl jspl_w_n1257_0(.douta(w_n1257_0[0]),.doutb(w_n1257_0[1]),.din(w_dff_B_bV6shDjr6_2));
	jspl jspl_w_n1260_0(.douta(w_n1260_0[0]),.doutb(w_n1260_0[1]),.din(n1260));
	jspl jspl_w_n1262_0(.douta(w_n1262_0[0]),.doutb(w_n1262_0[1]),.din(w_dff_B_AteBDex17_2));
	jspl jspl_w_n1265_0(.douta(w_n1265_0[0]),.doutb(w_n1265_0[1]),.din(n1265));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(w_dff_B_E3ivLrTe7_2));
	jspl jspl_w_n1267_0(.douta(w_n1267_0[0]),.doutb(w_n1267_0[1]),.din(w_dff_B_W5C7l31p9_2));
	jspl jspl_w_n1270_0(.douta(w_n1270_0[0]),.doutb(w_n1270_0[1]),.din(n1270));
	jspl jspl_w_n1272_0(.douta(w_n1272_0[0]),.doutb(w_n1272_0[1]),.din(n1272));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(w_dff_B_PKQSLXiP0_2));
	jspl jspl_w_n1274_0(.douta(w_n1274_0[0]),.doutb(w_n1274_0[1]),.din(n1274));
	jspl jspl_w_n1275_0(.douta(w_n1275_0[0]),.doutb(w_n1275_0[1]),.din(w_dff_B_xxLYShRk6_2));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(n1276));
	jspl jspl_w_n1277_0(.douta(w_n1277_0[0]),.doutb(w_n1277_0[1]),.din(w_dff_B_N8V3kiDx4_2));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(n1278));
	jspl jspl_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.din(w_dff_B_c3ouuaHN5_2));
	jspl jspl_w_n1280_0(.douta(w_n1280_0[0]),.doutb(w_n1280_0[1]),.din(n1280));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(w_dff_B_wqiKM8GG9_2));
	jspl jspl_w_n1282_0(.douta(w_n1282_0[0]),.doutb(w_n1282_0[1]),.din(n1282));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(w_dff_B_gQfjdZlo5_2));
	jspl jspl_w_n1284_0(.douta(w_n1284_0[0]),.doutb(w_n1284_0[1]),.din(n1284));
	jspl jspl_w_n1285_0(.douta(w_n1285_0[0]),.doutb(w_n1285_0[1]),.din(w_dff_B_Fhg9wTZk4_2));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(n1286));
	jspl jspl_w_n1287_0(.douta(w_n1287_0[0]),.doutb(w_n1287_0[1]),.din(n1287));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(n1288));
	jspl jspl_w_n1289_0(.douta(w_n1289_0[0]),.doutb(w_n1289_0[1]),.din(n1289));
	jspl jspl_w_n1290_0(.douta(w_n1290_0[0]),.doutb(w_n1290_0[1]),.din(n1290));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_dff_A_lYf27aFO6_1),.din(n1291));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(n1293));
	jspl jspl_w_n1294_0(.douta(w_n1294_0[0]),.doutb(w_dff_A_SO1P2mKd0_1),.din(n1294));
	jspl jspl_w_n1295_0(.douta(w_dff_A_d5qDWqJV6_0),.doutb(w_n1295_0[1]),.din(n1295));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(w_dff_B_Lo8FIWC53_2));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(w_dff_B_GTCAo03K0_2));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(w_dff_B_2Kdu6SYs4_2));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.din(w_dff_B_1yz24uV28_2));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl jspl_w_n1327_0(.douta(w_n1327_0[0]),.doutb(w_n1327_0[1]),.din(w_dff_B_DoOjH9fV8_2));
	jspl jspl_w_n1330_0(.douta(w_n1330_0[0]),.doutb(w_n1330_0[1]),.din(n1330));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(w_dff_B_efYzMPz54_2));
	jspl jspl_w_n1335_0(.douta(w_n1335_0[0]),.doutb(w_n1335_0[1]),.din(n1335));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(w_dff_B_YqVPXIAC4_2));
	jspl jspl_w_n1340_0(.douta(w_n1340_0[0]),.doutb(w_n1340_0[1]),.din(n1340));
	jspl jspl_w_n1342_0(.douta(w_n1342_0[0]),.doutb(w_n1342_0[1]),.din(w_dff_B_MxE3o1cU9_2));
	jspl jspl_w_n1345_0(.douta(w_n1345_0[0]),.doutb(w_n1345_0[1]),.din(n1345));
	jspl jspl_w_n1347_0(.douta(w_n1347_0[0]),.doutb(w_n1347_0[1]),.din(w_dff_B_jfnFqI8W0_2));
	jspl jspl_w_n1350_0(.douta(w_n1350_0[0]),.doutb(w_n1350_0[1]),.din(n1350));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(w_dff_B_R1ismnub3_2));
	jspl jspl_w_n1352_0(.douta(w_n1352_0[0]),.doutb(w_n1352_0[1]),.din(w_dff_B_id4ZkbFR2_2));
	jspl jspl_w_n1355_0(.douta(w_n1355_0[0]),.doutb(w_n1355_0[1]),.din(n1355));
	jspl jspl_w_n1357_0(.douta(w_n1357_0[0]),.doutb(w_n1357_0[1]),.din(n1357));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_n1359_0[1]),.din(n1359));
	jspl jspl_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.din(w_dff_B_9iqGyKXP9_2));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1362_0(.douta(w_n1362_0[0]),.doutb(w_n1362_0[1]),.din(w_dff_B_R2EcHsrg1_2));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(n1363));
	jspl jspl_w_n1364_0(.douta(w_n1364_0[0]),.doutb(w_n1364_0[1]),.din(w_dff_B_SkDVNICh2_2));
	jspl jspl_w_n1365_0(.douta(w_n1365_0[0]),.doutb(w_n1365_0[1]),.din(n1365));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(w_dff_B_krZPfOzy8_2));
	jspl jspl_w_n1367_0(.douta(w_n1367_0[0]),.doutb(w_n1367_0[1]),.din(n1367));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(w_dff_B_FRdNxege6_2));
	jspl jspl_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.din(n1369));
	jspl jspl_w_n1370_0(.douta(w_n1370_0[0]),.doutb(w_n1370_0[1]),.din(w_dff_B_SkmqDCMx4_2));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.din(n1372));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(n1373));
	jspl jspl_w_n1374_0(.douta(w_n1374_0[0]),.doutb(w_n1374_0[1]),.din(n1374));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(n1376));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(n1378));
	jspl jspl_w_n1379_0(.douta(w_n1379_0[0]),.doutb(w_dff_A_QwUZQSPN3_1),.din(n1379));
	jspl jspl_w_n1384_0(.douta(w_n1384_0[0]),.doutb(w_n1384_0[1]),.din(n1384));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(w_dff_B_HsitQwma1_2));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(w_dff_B_RlCGGr5Y0_2));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(w_dff_B_jTp396Bm6_2));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(w_dff_B_lW0kk8354_2));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(w_dff_B_FlcmKFLv6_2));
	jspl jspl_w_n1408_0(.douta(w_n1408_0[0]),.doutb(w_n1408_0[1]),.din(n1408));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(w_dff_B_Hlxo0DKL6_2));
	jspl jspl_w_n1413_0(.douta(w_n1413_0[0]),.doutb(w_n1413_0[1]),.din(n1413));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(w_dff_B_XmFqVPUy1_2));
	jspl jspl_w_n1418_0(.douta(w_n1418_0[0]),.doutb(w_n1418_0[1]),.din(n1418));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(w_dff_B_e40zLt7F6_2));
	jspl jspl_w_n1423_0(.douta(w_n1423_0[0]),.doutb(w_n1423_0[1]),.din(n1423));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(w_dff_B_cW7nfghM3_2));
	jspl jspl_w_n1428_0(.douta(w_n1428_0[0]),.doutb(w_n1428_0[1]),.din(w_dff_B_1XAPDj0M1_2));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(w_dff_B_gF9ti5EF3_2));
	jspl jspl_w_n1430_0(.douta(w_n1430_0[0]),.doutb(w_n1430_0[1]),.din(w_dff_B_y2SyWNyp8_2));
	jspl jspl_w_n1433_0(.douta(w_n1433_0[0]),.doutb(w_n1433_0[1]),.din(n1433));
	jspl jspl_w_n1435_0(.douta(w_n1435_0[0]),.doutb(w_n1435_0[1]),.din(n1435));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(n1436));
	jspl jspl_w_n1437_0(.douta(w_n1437_0[0]),.doutb(w_n1437_0[1]),.din(n1437));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_n1438_0[1]),.din(n1438));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.din(w_dff_B_uFhzbbnU0_2));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl jspl_w_n1442_0(.douta(w_n1442_0[0]),.doutb(w_n1442_0[1]),.din(w_dff_B_tqh4Egzt0_2));
	jspl jspl_w_n1443_0(.douta(w_n1443_0[0]),.doutb(w_n1443_0[1]),.din(n1443));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(w_dff_B_9zXT8tMX6_2));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(w_dff_B_mbhr9m1M1_2));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1448_0(.douta(w_n1448_0[0]),.doutb(w_n1448_0[1]),.din(w_dff_B_jfnSrci08_2));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(n1449));
	jspl jspl_w_n1450_0(.douta(w_n1450_0[0]),.doutb(w_n1450_0[1]),.din(n1450));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(n1454));
	jspl jspl_w_n1455_0(.douta(w_n1455_0[0]),.doutb(w_dff_A_CpR4vvnb3_1),.din(n1455));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(n1460));
	jspl jspl_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.din(w_dff_B_8w74N4ai7_2));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(w_dff_B_KmYUFH5k9_2));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(w_dff_B_tdWHgp7n9_2));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(n1474));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(w_dff_B_ooaUOpmP9_2));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(n1479));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(w_dff_B_7kyonYWH5_2));
	jspl jspl_w_n1484_0(.douta(w_n1484_0[0]),.doutb(w_n1484_0[1]),.din(n1484));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(w_dff_B_vgDz7HGl0_2));
	jspl jspl_w_n1489_0(.douta(w_n1489_0[0]),.doutb(w_n1489_0[1]),.din(n1489));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(w_dff_B_9zzKoBVo7_2));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(w_dff_B_Z5aK2Mqf8_2));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(w_dff_B_xOdbxLaE6_2));
	jspl jspl_w_n1499_0(.douta(w_n1499_0[0]),.doutb(w_n1499_0[1]),.din(w_dff_B_63ITM0IV8_2));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(w_dff_B_sF8K7eJt7_2));
	jspl jspl_w_n1501_0(.douta(w_n1501_0[0]),.doutb(w_n1501_0[1]),.din(w_dff_B_YQMQaZxU4_2));
	jspl jspl_w_n1504_0(.douta(w_n1504_0[0]),.doutb(w_n1504_0[1]),.din(n1504));
	jspl jspl_w_n1506_0(.douta(w_n1506_0[0]),.doutb(w_n1506_0[1]),.din(n1506));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(n1507));
	jspl jspl_w_n1508_0(.douta(w_n1508_0[0]),.doutb(w_n1508_0[1]),.din(n1508));
	jspl jspl_w_n1509_0(.douta(w_n1509_0[0]),.doutb(w_n1509_0[1]),.din(n1509));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1511_0(.douta(w_n1511_0[0]),.doutb(w_n1511_0[1]),.din(n1511));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(n1512));
	jspl jspl_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.din(w_dff_B_Lxj1A7jA7_2));
	jspl jspl_w_n1514_0(.douta(w_n1514_0[0]),.doutb(w_n1514_0[1]),.din(n1514));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(w_dff_B_y0v4w9nr6_2));
	jspl jspl_w_n1516_0(.douta(w_n1516_0[0]),.doutb(w_n1516_0[1]),.din(n1516));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(w_dff_B_wuiWfaLW9_2));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl jspl_w_n1519_0(.douta(w_n1519_0[0]),.doutb(w_dff_A_zDIQNUSH4_1),.din(n1519));
	jspl jspl_w_n1521_0(.douta(w_n1521_0[0]),.doutb(w_n1521_0[1]),.din(n1521));
	jspl jspl_w_n1523_0(.douta(w_n1523_0[0]),.doutb(w_n1523_0[1]),.din(n1523));
	jspl jspl_w_n1524_0(.douta(w_n1524_0[0]),.doutb(w_dff_A_wCShQUCq8_1),.din(n1524));
	jspl jspl_w_n1529_0(.douta(w_n1529_0[0]),.doutb(w_n1529_0[1]),.din(n1529));
	jspl jspl_w_n1534_0(.douta(w_n1534_0[0]),.doutb(w_n1534_0[1]),.din(n1534));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(w_dff_B_JtkMUbzs3_2));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(w_dff_B_qf6KaGu87_2));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(w_dff_B_ryjsFclc7_2));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(n1548));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_n1550_0[1]),.din(w_dff_B_74fhHmmo4_2));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(w_dff_B_zJmFRF1S3_2));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(w_dff_B_hVjhuHCc7_2));
	jspl jspl_w_n1558_0(.douta(w_n1558_0[0]),.doutb(w_n1558_0[1]),.din(w_dff_B_wI1VmqpV6_2));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(w_dff_B_NCLO9bGl6_2));
	jspl jspl_w_n1563_0(.douta(w_n1563_0[0]),.doutb(w_n1563_0[1]),.din(w_dff_B_Lc401koj9_2));
	jspl jspl_w_n1564_0(.douta(w_n1564_0[0]),.doutb(w_n1564_0[1]),.din(w_dff_B_AtA3bWf96_2));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(w_dff_B_q34FxeZk2_2));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_n1568_0[1]),.din(n1568));
	jspl jspl_w_n1570_0(.douta(w_n1570_0[0]),.doutb(w_n1570_0[1]),.din(n1570));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(n1571));
	jspl jspl_w_n1572_0(.douta(w_n1572_0[0]),.doutb(w_n1572_0[1]),.din(n1572));
	jspl jspl_w_n1573_0(.douta(w_n1573_0[0]),.doutb(w_n1573_0[1]),.din(n1573));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(n1574));
	jspl jspl_w_n1575_0(.douta(w_n1575_0[0]),.doutb(w_n1575_0[1]),.din(n1575));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(n1576));
	jspl jspl_w_n1577_0(.douta(w_n1577_0[0]),.doutb(w_n1577_0[1]),.din(n1577));
	jspl jspl_w_n1578_0(.douta(w_n1578_0[0]),.doutb(w_n1578_0[1]),.din(n1578));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(w_dff_B_f5jzpFwY9_2));
	jspl jspl_w_n1580_0(.douta(w_n1580_0[0]),.doutb(w_n1580_0[1]),.din(n1580));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_dff_A_s2XrVx6R2_1),.din(n1581));
	jspl jspl_w_n1583_0(.douta(w_n1583_0[0]),.doutb(w_n1583_0[1]),.din(n1583));
	jspl jspl_w_n1585_0(.douta(w_n1585_0[0]),.doutb(w_n1585_0[1]),.din(n1585));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_dff_A_UV68AmjS3_1),.din(n1586));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(n1596));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(w_dff_B_sg5RzDjZ8_2));
	jspl jspl_w_n1600_0(.douta(w_n1600_0[0]),.doutb(w_n1600_0[1]),.din(n1600));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(w_dff_B_RQf5jV8H4_2));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(w_dff_B_8O6FL66n5_2));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(w_dff_B_ak5udAVA0_2));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(w_dff_B_Ft9mJuO39_2));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(w_dff_B_NU2VaBpl9_2));
	jspl jspl_w_n1615_0(.douta(w_n1615_0[0]),.doutb(w_n1615_0[1]),.din(w_dff_B_eSWBskYx7_2));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_n1617_0[1]),.din(w_dff_B_tYEo24vg1_2));
	jspl jspl_w_n1620_0(.douta(w_n1620_0[0]),.doutb(w_n1620_0[1]),.din(w_dff_B_RXKSSsqR2_2));
	jspl jspl_w_n1621_0(.douta(w_n1621_0[0]),.doutb(w_n1621_0[1]),.din(w_dff_B_fUIKiS5m0_2));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(w_dff_B_Xpc4Xt2r4_2));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(n1628));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1630_0(.douta(w_n1630_0[0]),.doutb(w_n1630_0[1]),.din(n1630));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(n1631));
	jspl jspl_w_n1632_0(.douta(w_n1632_0[0]),.doutb(w_n1632_0[1]),.din(n1632));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(n1633));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(n1634));
	jspl jspl_w_n1635_0(.douta(w_n1635_0[0]),.doutb(w_n1635_0[1]),.din(n1635));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(n1636));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(n1638));
	jspl jspl_w_n1640_0(.douta(w_n1640_0[0]),.doutb(w_n1640_0[1]),.din(n1640));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_dff_A_TtZdaZ396_1),.din(n1641));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(n1646));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(w_dff_B_5UjToAl94_2));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(w_dff_B_pE3RY6EJ3_2));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(w_dff_B_sNHG63tc4_2));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(w_dff_B_XKc9uIkO5_2));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(w_dff_B_5O1Mhl5G7_2));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(w_dff_B_YReXbETt0_2));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(w_dff_B_AIRwaqk58_2));
	jspl jspl_w_n1668_0(.douta(w_n1668_0[0]),.doutb(w_n1668_0[1]),.din(w_dff_B_d19QqC920_2));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(w_dff_B_KI6zkGY98_2));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(w_dff_B_qm4Xdjn60_2));
	jspl jspl_w_n1673_0(.douta(w_n1673_0[0]),.doutb(w_n1673_0[1]),.din(w_dff_B_uCOPYHHr4_2));
	jspl jspl_w_n1676_0(.douta(w_n1676_0[0]),.doutb(w_n1676_0[1]),.din(n1676));
	jspl jspl_w_n1678_0(.douta(w_n1678_0[0]),.doutb(w_n1678_0[1]),.din(n1678));
	jspl jspl_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.din(n1679));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1681_0(.douta(w_n1681_0[0]),.doutb(w_n1681_0[1]),.din(n1681));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(n1682));
	jspl jspl_w_n1683_0(.douta(w_n1683_0[0]),.doutb(w_n1683_0[1]),.din(n1683));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(n1684));
	jspl jspl_w_n1685_0(.douta(w_n1685_0[0]),.doutb(w_n1685_0[1]),.din(n1685));
	jspl jspl_w_n1686_0(.douta(w_n1686_0[0]),.doutb(w_n1686_0[1]),.din(n1686));
	jspl jspl_w_n1688_0(.douta(w_n1688_0[0]),.doutb(w_n1688_0[1]),.din(n1688));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_dff_A_cIRgkc145_1),.din(n1689));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(n1694));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_dff_A_kB4EvvLH8_1),.din(n1697));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(w_dff_B_6OjCEdhs7_2));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(w_dff_B_JpN0rZj48_2));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(w_dff_B_99nspnyh2_2));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(w_dff_B_9eIiVIDf5_2));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(w_dff_B_RXpiju8U5_2));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(w_dff_B_tXWfrrrp7_2));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(w_dff_B_VE9RbqXC4_2));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(w_dff_B_c3ReEHRB7_2));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_n1720_0[1]),.din(n1720));
	jspl jspl_w_n1721_0(.douta(w_n1721_0[0]),.doutb(w_n1721_0[1]),.din(n1721));
	jspl jspl_w_n1722_0(.douta(w_n1722_0[0]),.doutb(w_n1722_0[1]),.din(n1722));
	jspl jspl_w_n1723_0(.douta(w_n1723_0[0]),.doutb(w_n1723_0[1]),.din(n1723));
	jspl jspl_w_n1724_0(.douta(w_n1724_0[0]),.doutb(w_n1724_0[1]),.din(n1724));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1726_0(.douta(w_n1726_0[0]),.doutb(w_n1726_0[1]),.din(n1726));
	jspl jspl_w_n1727_0(.douta(w_n1727_0[0]),.doutb(w_dff_A_Sd21jNyI9_1),.din(n1727));
	jspl jspl_w_n1734_0(.douta(w_n1734_0[0]),.doutb(w_n1734_0[1]),.din(n1734));
	jspl jspl_w_n1737_0(.douta(w_n1737_0[0]),.doutb(w_dff_A_NtY58GGi5_1),.din(n1737));
	jspl jspl_w_n1739_0(.douta(w_n1739_0[0]),.doutb(w_n1739_0[1]),.din(w_dff_B_LKZsNJGw4_2));
	jspl jspl_w_n1742_0(.douta(w_n1742_0[0]),.doutb(w_n1742_0[1]),.din(w_dff_B_fNHkhFqF1_2));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(w_dff_B_J8pEQWx43_2));
	jspl jspl_w_n1747_0(.douta(w_n1747_0[0]),.doutb(w_n1747_0[1]),.din(w_dff_B_pFri1iHH0_2));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(w_dff_B_sbxCKHqq8_2));
	jspl jspl_w_n1749_0(.douta(w_n1749_0[0]),.doutb(w_n1749_0[1]),.din(w_dff_B_GdviRPqa7_2));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_n1758_0[1]),.din(n1758));
	jspl jspl_w_n1759_0(.douta(w_n1759_0[0]),.doutb(w_n1759_0[1]),.din(n1759));
	jspl jspl_w_n1760_0(.douta(w_n1760_0[0]),.doutb(w_dff_A_vJw6EZhk6_1),.din(n1760));
	jspl jspl_w_n1767_0(.douta(w_n1767_0[0]),.doutb(w_n1767_0[1]),.din(n1767));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_dff_A_bbY4ozxq3_1),.din(n1770));
	jspl jspl_w_n1772_0(.douta(w_n1772_0[0]),.doutb(w_n1772_0[1]),.din(w_dff_B_85nnEfjK5_2));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(w_dff_B_xwJvQPur6_2));
	jspl jspl_w_n1776_0(.douta(w_n1776_0[0]),.doutb(w_n1776_0[1]),.din(w_dff_B_BMwC0cpx0_2));
	jspl jspl_w_n1777_0(.douta(w_n1777_0[0]),.doutb(w_n1777_0[1]),.din(w_dff_B_Z6YhwrNl1_2));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(n1780));
	jspl jspl_w_n1782_0(.douta(w_n1782_0[0]),.doutb(w_n1782_0[1]),.din(n1782));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1784_0(.douta(w_n1784_0[0]),.doutb(w_n1784_0[1]),.din(n1784));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_dff_A_X2uFtJnt5_1),.din(n1786));
	jspl jspl_w_n1793_0(.douta(w_n1793_0[0]),.doutb(w_n1793_0[1]),.din(n1793));
	jspl jspl_w_n1796_0(.douta(w_n1796_0[0]),.doutb(w_dff_A_WUTJTKWd2_1),.din(n1796));
	jspl jspl_w_n1797_0(.douta(w_n1797_0[0]),.doutb(w_n1797_0[1]),.din(w_dff_B_hAmTZHFN2_2));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(w_dff_B_Yqe5obyU9_2));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_n1801_0[1]),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(n1803));
	jspl jspl_w_n1804_0(.douta(w_n1804_0[0]),.doutb(w_n1804_0[1]),.din(n1804));
	jspl jspl_w_n1805_0(.douta(w_n1805_0[0]),.doutb(w_dff_A_U4LD1zzq3_1),.din(n1805));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(w_dff_B_U2lBJJDX5_2));
	jspl jspl_w_n1810_0(.douta(w_n1810_0[0]),.doutb(w_n1810_0[1]),.din(n1810));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_n1817_0[1]),.din(n1817));
	jspl jspl_w_n1818_0(.douta(w_dff_A_5WGFEFAr1_0),.doutb(w_n1818_0[1]),.din(n1818));
	jdff dff_B_6EbCXpH77_0(.din(n72),.dout(w_dff_B_6EbCXpH77_0),.clk(gclk));
	jdff dff_B_xtZmTHUA1_0(.din(w_dff_B_6EbCXpH77_0),.dout(w_dff_B_xtZmTHUA1_0),.clk(gclk));
	jdff dff_B_8eVh8Wnb7_1(.din(n76),.dout(w_dff_B_8eVh8Wnb7_1),.clk(gclk));
	jdff dff_B_4JcfhAzb9_1(.din(w_dff_B_8eVh8Wnb7_1),.dout(w_dff_B_4JcfhAzb9_1),.clk(gclk));
	jdff dff_B_c1j5Gyez3_1(.din(w_dff_B_4JcfhAzb9_1),.dout(w_dff_B_c1j5Gyez3_1),.clk(gclk));
	jdff dff_B_PVNT4aGx9_1(.din(n87),.dout(w_dff_B_PVNT4aGx9_1),.clk(gclk));
	jdff dff_B_JaUmz1Va5_1(.din(w_dff_B_PVNT4aGx9_1),.dout(w_dff_B_JaUmz1Va5_1),.clk(gclk));
	jdff dff_B_S7dPF5m53_1(.din(w_dff_B_JaUmz1Va5_1),.dout(w_dff_B_S7dPF5m53_1),.clk(gclk));
	jdff dff_B_s7M86MFT7_1(.din(w_dff_B_S7dPF5m53_1),.dout(w_dff_B_s7M86MFT7_1),.clk(gclk));
	jdff dff_B_1KvYvi7e1_1(.din(w_dff_B_s7M86MFT7_1),.dout(w_dff_B_1KvYvi7e1_1),.clk(gclk));
	jdff dff_B_TnLU4N4R5_1(.din(w_dff_B_1KvYvi7e1_1),.dout(w_dff_B_TnLU4N4R5_1),.clk(gclk));
	jdff dff_B_FS2Gflch8_1(.din(n107),.dout(w_dff_B_FS2Gflch8_1),.clk(gclk));
	jdff dff_B_bTw3ySpl4_1(.din(w_dff_B_FS2Gflch8_1),.dout(w_dff_B_bTw3ySpl4_1),.clk(gclk));
	jdff dff_B_fKN0GiF25_1(.din(w_dff_B_bTw3ySpl4_1),.dout(w_dff_B_fKN0GiF25_1),.clk(gclk));
	jdff dff_B_NvRmulmG2_1(.din(w_dff_B_fKN0GiF25_1),.dout(w_dff_B_NvRmulmG2_1),.clk(gclk));
	jdff dff_B_FEOzBdld7_1(.din(w_dff_B_NvRmulmG2_1),.dout(w_dff_B_FEOzBdld7_1),.clk(gclk));
	jdff dff_B_GtpBJpdl5_1(.din(w_dff_B_FEOzBdld7_1),.dout(w_dff_B_GtpBJpdl5_1),.clk(gclk));
	jdff dff_B_trBLxzOo0_1(.din(w_dff_B_GtpBJpdl5_1),.dout(w_dff_B_trBLxzOo0_1),.clk(gclk));
	jdff dff_B_TuXcG4bf5_1(.din(w_dff_B_trBLxzOo0_1),.dout(w_dff_B_TuXcG4bf5_1),.clk(gclk));
	jdff dff_B_2bca4tz20_1(.din(w_dff_B_TuXcG4bf5_1),.dout(w_dff_B_2bca4tz20_1),.clk(gclk));
	jdff dff_B_fY7JYVwV5_1(.din(n136),.dout(w_dff_B_fY7JYVwV5_1),.clk(gclk));
	jdff dff_B_f80I4H8v9_1(.din(w_dff_B_fY7JYVwV5_1),.dout(w_dff_B_f80I4H8v9_1),.clk(gclk));
	jdff dff_B_n56lUK196_1(.din(w_dff_B_f80I4H8v9_1),.dout(w_dff_B_n56lUK196_1),.clk(gclk));
	jdff dff_B_EfJA0pmZ5_1(.din(w_dff_B_n56lUK196_1),.dout(w_dff_B_EfJA0pmZ5_1),.clk(gclk));
	jdff dff_B_i89h6el13_1(.din(w_dff_B_EfJA0pmZ5_1),.dout(w_dff_B_i89h6el13_1),.clk(gclk));
	jdff dff_B_9opOCRek1_1(.din(w_dff_B_i89h6el13_1),.dout(w_dff_B_9opOCRek1_1),.clk(gclk));
	jdff dff_B_uAw445A47_1(.din(w_dff_B_9opOCRek1_1),.dout(w_dff_B_uAw445A47_1),.clk(gclk));
	jdff dff_B_6SLWFlgP9_1(.din(w_dff_B_uAw445A47_1),.dout(w_dff_B_6SLWFlgP9_1),.clk(gclk));
	jdff dff_B_SoefDKPz1_1(.din(w_dff_B_6SLWFlgP9_1),.dout(w_dff_B_SoefDKPz1_1),.clk(gclk));
	jdff dff_B_WDui7EWV9_1(.din(w_dff_B_SoefDKPz1_1),.dout(w_dff_B_WDui7EWV9_1),.clk(gclk));
	jdff dff_B_UqUZaCXs4_1(.din(w_dff_B_WDui7EWV9_1),.dout(w_dff_B_UqUZaCXs4_1),.clk(gclk));
	jdff dff_B_M3AxJSlC9_1(.din(w_dff_B_UqUZaCXs4_1),.dout(w_dff_B_M3AxJSlC9_1),.clk(gclk));
	jdff dff_B_LFYlq8cZ0_1(.din(n171),.dout(w_dff_B_LFYlq8cZ0_1),.clk(gclk));
	jdff dff_B_VKDa8BD95_1(.din(w_dff_B_LFYlq8cZ0_1),.dout(w_dff_B_VKDa8BD95_1),.clk(gclk));
	jdff dff_B_B9rGcLtU8_1(.din(w_dff_B_VKDa8BD95_1),.dout(w_dff_B_B9rGcLtU8_1),.clk(gclk));
	jdff dff_B_hTuES3dj1_1(.din(w_dff_B_B9rGcLtU8_1),.dout(w_dff_B_hTuES3dj1_1),.clk(gclk));
	jdff dff_B_v9F38lDU3_1(.din(w_dff_B_hTuES3dj1_1),.dout(w_dff_B_v9F38lDU3_1),.clk(gclk));
	jdff dff_B_Hx7aAZiW0_1(.din(w_dff_B_v9F38lDU3_1),.dout(w_dff_B_Hx7aAZiW0_1),.clk(gclk));
	jdff dff_B_tN1jq0LE5_1(.din(w_dff_B_Hx7aAZiW0_1),.dout(w_dff_B_tN1jq0LE5_1),.clk(gclk));
	jdff dff_B_KvRtTdHc6_1(.din(w_dff_B_tN1jq0LE5_1),.dout(w_dff_B_KvRtTdHc6_1),.clk(gclk));
	jdff dff_B_jrQjBfkc6_1(.din(w_dff_B_KvRtTdHc6_1),.dout(w_dff_B_jrQjBfkc6_1),.clk(gclk));
	jdff dff_B_ob4NYxlA0_1(.din(w_dff_B_jrQjBfkc6_1),.dout(w_dff_B_ob4NYxlA0_1),.clk(gclk));
	jdff dff_B_N65PrVWl8_1(.din(w_dff_B_ob4NYxlA0_1),.dout(w_dff_B_N65PrVWl8_1),.clk(gclk));
	jdff dff_B_eSr03Dgt7_1(.din(w_dff_B_N65PrVWl8_1),.dout(w_dff_B_eSr03Dgt7_1),.clk(gclk));
	jdff dff_B_daeICTUl4_1(.din(w_dff_B_eSr03Dgt7_1),.dout(w_dff_B_daeICTUl4_1),.clk(gclk));
	jdff dff_B_J8n7Q3YB3_1(.din(w_dff_B_daeICTUl4_1),.dout(w_dff_B_J8n7Q3YB3_1),.clk(gclk));
	jdff dff_B_DOxgFj537_1(.din(w_dff_B_J8n7Q3YB3_1),.dout(w_dff_B_DOxgFj537_1),.clk(gclk));
	jdff dff_B_StChmr9P4_1(.din(n213),.dout(w_dff_B_StChmr9P4_1),.clk(gclk));
	jdff dff_B_YMTpwJuY0_1(.din(w_dff_B_StChmr9P4_1),.dout(w_dff_B_YMTpwJuY0_1),.clk(gclk));
	jdff dff_B_tmoHPFN09_1(.din(w_dff_B_YMTpwJuY0_1),.dout(w_dff_B_tmoHPFN09_1),.clk(gclk));
	jdff dff_B_yCjB3KRH9_1(.din(w_dff_B_tmoHPFN09_1),.dout(w_dff_B_yCjB3KRH9_1),.clk(gclk));
	jdff dff_B_YZCWiTtL4_1(.din(w_dff_B_yCjB3KRH9_1),.dout(w_dff_B_YZCWiTtL4_1),.clk(gclk));
	jdff dff_B_VWRvGCNO2_1(.din(w_dff_B_YZCWiTtL4_1),.dout(w_dff_B_VWRvGCNO2_1),.clk(gclk));
	jdff dff_B_uVSwz0Lu1_1(.din(w_dff_B_VWRvGCNO2_1),.dout(w_dff_B_uVSwz0Lu1_1),.clk(gclk));
	jdff dff_B_cTW4zgFp8_1(.din(w_dff_B_uVSwz0Lu1_1),.dout(w_dff_B_cTW4zgFp8_1),.clk(gclk));
	jdff dff_B_SGk1TWIE0_1(.din(w_dff_B_cTW4zgFp8_1),.dout(w_dff_B_SGk1TWIE0_1),.clk(gclk));
	jdff dff_B_zVogGwtN2_1(.din(w_dff_B_SGk1TWIE0_1),.dout(w_dff_B_zVogGwtN2_1),.clk(gclk));
	jdff dff_B_uOGSDFNo5_1(.din(w_dff_B_zVogGwtN2_1),.dout(w_dff_B_uOGSDFNo5_1),.clk(gclk));
	jdff dff_B_RGfjPcz20_1(.din(w_dff_B_uOGSDFNo5_1),.dout(w_dff_B_RGfjPcz20_1),.clk(gclk));
	jdff dff_B_MTuAQUhG6_1(.din(w_dff_B_RGfjPcz20_1),.dout(w_dff_B_MTuAQUhG6_1),.clk(gclk));
	jdff dff_B_igP4oBDl2_1(.din(w_dff_B_MTuAQUhG6_1),.dout(w_dff_B_igP4oBDl2_1),.clk(gclk));
	jdff dff_B_mi7TkSlU3_1(.din(w_dff_B_igP4oBDl2_1),.dout(w_dff_B_mi7TkSlU3_1),.clk(gclk));
	jdff dff_B_P7CtA1N89_1(.din(w_dff_B_mi7TkSlU3_1),.dout(w_dff_B_P7CtA1N89_1),.clk(gclk));
	jdff dff_B_4pcr0ilK7_1(.din(w_dff_B_P7CtA1N89_1),.dout(w_dff_B_4pcr0ilK7_1),.clk(gclk));
	jdff dff_B_DtxLqxqv7_1(.din(w_dff_B_4pcr0ilK7_1),.dout(w_dff_B_DtxLqxqv7_1),.clk(gclk));
	jdff dff_B_SgOCHxAj6_1(.din(n262),.dout(w_dff_B_SgOCHxAj6_1),.clk(gclk));
	jdff dff_B_O3FUU1Ss4_1(.din(w_dff_B_SgOCHxAj6_1),.dout(w_dff_B_O3FUU1Ss4_1),.clk(gclk));
	jdff dff_B_cyUrzFXY2_1(.din(w_dff_B_O3FUU1Ss4_1),.dout(w_dff_B_cyUrzFXY2_1),.clk(gclk));
	jdff dff_B_ylPbca7d0_1(.din(w_dff_B_cyUrzFXY2_1),.dout(w_dff_B_ylPbca7d0_1),.clk(gclk));
	jdff dff_B_TezgXW8k5_1(.din(w_dff_B_ylPbca7d0_1),.dout(w_dff_B_TezgXW8k5_1),.clk(gclk));
	jdff dff_B_chzPvfiq8_1(.din(w_dff_B_TezgXW8k5_1),.dout(w_dff_B_chzPvfiq8_1),.clk(gclk));
	jdff dff_B_8FA1HqLd1_1(.din(w_dff_B_chzPvfiq8_1),.dout(w_dff_B_8FA1HqLd1_1),.clk(gclk));
	jdff dff_B_9HKf2dSi8_1(.din(w_dff_B_8FA1HqLd1_1),.dout(w_dff_B_9HKf2dSi8_1),.clk(gclk));
	jdff dff_B_WbfZrgI67_1(.din(w_dff_B_9HKf2dSi8_1),.dout(w_dff_B_WbfZrgI67_1),.clk(gclk));
	jdff dff_B_3gWwstnp9_1(.din(w_dff_B_WbfZrgI67_1),.dout(w_dff_B_3gWwstnp9_1),.clk(gclk));
	jdff dff_B_L9SJeKrO7_1(.din(w_dff_B_3gWwstnp9_1),.dout(w_dff_B_L9SJeKrO7_1),.clk(gclk));
	jdff dff_B_LrxxM1bT3_1(.din(w_dff_B_L9SJeKrO7_1),.dout(w_dff_B_LrxxM1bT3_1),.clk(gclk));
	jdff dff_B_Cb1wrOak1_1(.din(w_dff_B_LrxxM1bT3_1),.dout(w_dff_B_Cb1wrOak1_1),.clk(gclk));
	jdff dff_B_SgKKyl412_1(.din(w_dff_B_Cb1wrOak1_1),.dout(w_dff_B_SgKKyl412_1),.clk(gclk));
	jdff dff_B_eRwawQsp9_1(.din(w_dff_B_SgKKyl412_1),.dout(w_dff_B_eRwawQsp9_1),.clk(gclk));
	jdff dff_B_teDoWhVc9_1(.din(w_dff_B_eRwawQsp9_1),.dout(w_dff_B_teDoWhVc9_1),.clk(gclk));
	jdff dff_B_xEctTbmu9_1(.din(w_dff_B_teDoWhVc9_1),.dout(w_dff_B_xEctTbmu9_1),.clk(gclk));
	jdff dff_B_xDzWTUSH9_1(.din(w_dff_B_xEctTbmu9_1),.dout(w_dff_B_xDzWTUSH9_1),.clk(gclk));
	jdff dff_B_XI4hWen59_1(.din(w_dff_B_xDzWTUSH9_1),.dout(w_dff_B_XI4hWen59_1),.clk(gclk));
	jdff dff_B_dxTOxvBm1_1(.din(w_dff_B_XI4hWen59_1),.dout(w_dff_B_dxTOxvBm1_1),.clk(gclk));
	jdff dff_B_8TdGlqOt4_1(.din(w_dff_B_dxTOxvBm1_1),.dout(w_dff_B_8TdGlqOt4_1),.clk(gclk));
	jdff dff_B_xCe6rYqH2_1(.din(n318),.dout(w_dff_B_xCe6rYqH2_1),.clk(gclk));
	jdff dff_B_rCfwRgoe0_1(.din(w_dff_B_xCe6rYqH2_1),.dout(w_dff_B_rCfwRgoe0_1),.clk(gclk));
	jdff dff_B_7xNDPKNx3_1(.din(w_dff_B_rCfwRgoe0_1),.dout(w_dff_B_7xNDPKNx3_1),.clk(gclk));
	jdff dff_B_rraDYe3f2_1(.din(w_dff_B_7xNDPKNx3_1),.dout(w_dff_B_rraDYe3f2_1),.clk(gclk));
	jdff dff_B_OZGA47qO8_1(.din(w_dff_B_rraDYe3f2_1),.dout(w_dff_B_OZGA47qO8_1),.clk(gclk));
	jdff dff_B_cXrSdBwG7_1(.din(w_dff_B_OZGA47qO8_1),.dout(w_dff_B_cXrSdBwG7_1),.clk(gclk));
	jdff dff_B_24VQ7H7T1_1(.din(w_dff_B_cXrSdBwG7_1),.dout(w_dff_B_24VQ7H7T1_1),.clk(gclk));
	jdff dff_B_vgfrHnC17_1(.din(w_dff_B_24VQ7H7T1_1),.dout(w_dff_B_vgfrHnC17_1),.clk(gclk));
	jdff dff_B_lwok5KC89_1(.din(w_dff_B_vgfrHnC17_1),.dout(w_dff_B_lwok5KC89_1),.clk(gclk));
	jdff dff_B_SiyGT3On8_1(.din(w_dff_B_lwok5KC89_1),.dout(w_dff_B_SiyGT3On8_1),.clk(gclk));
	jdff dff_B_Zmoc0Eb75_1(.din(w_dff_B_SiyGT3On8_1),.dout(w_dff_B_Zmoc0Eb75_1),.clk(gclk));
	jdff dff_B_67vY2LXH8_1(.din(w_dff_B_Zmoc0Eb75_1),.dout(w_dff_B_67vY2LXH8_1),.clk(gclk));
	jdff dff_B_XtFc66aC5_1(.din(w_dff_B_67vY2LXH8_1),.dout(w_dff_B_XtFc66aC5_1),.clk(gclk));
	jdff dff_B_nX6DvFbs7_1(.din(w_dff_B_XtFc66aC5_1),.dout(w_dff_B_nX6DvFbs7_1),.clk(gclk));
	jdff dff_B_kwkp0b7E2_1(.din(w_dff_B_nX6DvFbs7_1),.dout(w_dff_B_kwkp0b7E2_1),.clk(gclk));
	jdff dff_B_zbV1xpA51_1(.din(w_dff_B_kwkp0b7E2_1),.dout(w_dff_B_zbV1xpA51_1),.clk(gclk));
	jdff dff_B_0aJaneqd6_1(.din(w_dff_B_zbV1xpA51_1),.dout(w_dff_B_0aJaneqd6_1),.clk(gclk));
	jdff dff_B_QwSxNmHY6_1(.din(w_dff_B_0aJaneqd6_1),.dout(w_dff_B_QwSxNmHY6_1),.clk(gclk));
	jdff dff_B_wcTbZlve2_1(.din(w_dff_B_QwSxNmHY6_1),.dout(w_dff_B_wcTbZlve2_1),.clk(gclk));
	jdff dff_B_mf6fPMF03_1(.din(w_dff_B_wcTbZlve2_1),.dout(w_dff_B_mf6fPMF03_1),.clk(gclk));
	jdff dff_B_l1VaZjya2_1(.din(w_dff_B_mf6fPMF03_1),.dout(w_dff_B_l1VaZjya2_1),.clk(gclk));
	jdff dff_B_h6EyVqVB2_1(.din(w_dff_B_l1VaZjya2_1),.dout(w_dff_B_h6EyVqVB2_1),.clk(gclk));
	jdff dff_B_WhgrDOYv4_1(.din(w_dff_B_h6EyVqVB2_1),.dout(w_dff_B_WhgrDOYv4_1),.clk(gclk));
	jdff dff_B_KsiC9Zr79_1(.din(w_dff_B_WhgrDOYv4_1),.dout(w_dff_B_KsiC9Zr79_1),.clk(gclk));
	jdff dff_B_w2Qpxdxx9_1(.din(n381),.dout(w_dff_B_w2Qpxdxx9_1),.clk(gclk));
	jdff dff_B_Zog4Q74K6_1(.din(w_dff_B_w2Qpxdxx9_1),.dout(w_dff_B_Zog4Q74K6_1),.clk(gclk));
	jdff dff_B_0WgXiZAG4_1(.din(w_dff_B_Zog4Q74K6_1),.dout(w_dff_B_0WgXiZAG4_1),.clk(gclk));
	jdff dff_B_KJF7FvIw6_1(.din(w_dff_B_0WgXiZAG4_1),.dout(w_dff_B_KJF7FvIw6_1),.clk(gclk));
	jdff dff_B_qSq7upvm6_1(.din(w_dff_B_KJF7FvIw6_1),.dout(w_dff_B_qSq7upvm6_1),.clk(gclk));
	jdff dff_B_AoCZsmiq2_1(.din(w_dff_B_qSq7upvm6_1),.dout(w_dff_B_AoCZsmiq2_1),.clk(gclk));
	jdff dff_B_TrGx3jis2_1(.din(w_dff_B_AoCZsmiq2_1),.dout(w_dff_B_TrGx3jis2_1),.clk(gclk));
	jdff dff_B_bJzNGOuL6_1(.din(w_dff_B_TrGx3jis2_1),.dout(w_dff_B_bJzNGOuL6_1),.clk(gclk));
	jdff dff_B_rZeSt5sL0_1(.din(w_dff_B_bJzNGOuL6_1),.dout(w_dff_B_rZeSt5sL0_1),.clk(gclk));
	jdff dff_B_DI6sVi8z2_1(.din(w_dff_B_rZeSt5sL0_1),.dout(w_dff_B_DI6sVi8z2_1),.clk(gclk));
	jdff dff_B_rR0d9lqD3_1(.din(w_dff_B_DI6sVi8z2_1),.dout(w_dff_B_rR0d9lqD3_1),.clk(gclk));
	jdff dff_B_UnQyhgqA3_1(.din(w_dff_B_rR0d9lqD3_1),.dout(w_dff_B_UnQyhgqA3_1),.clk(gclk));
	jdff dff_B_vVH6eMGy7_1(.din(w_dff_B_UnQyhgqA3_1),.dout(w_dff_B_vVH6eMGy7_1),.clk(gclk));
	jdff dff_B_UHLQIkvA8_1(.din(w_dff_B_vVH6eMGy7_1),.dout(w_dff_B_UHLQIkvA8_1),.clk(gclk));
	jdff dff_B_33uwKasO8_1(.din(w_dff_B_UHLQIkvA8_1),.dout(w_dff_B_33uwKasO8_1),.clk(gclk));
	jdff dff_B_wRKtgU1X9_1(.din(w_dff_B_33uwKasO8_1),.dout(w_dff_B_wRKtgU1X9_1),.clk(gclk));
	jdff dff_B_6JIsAdm45_1(.din(w_dff_B_wRKtgU1X9_1),.dout(w_dff_B_6JIsAdm45_1),.clk(gclk));
	jdff dff_B_9jo6SD158_1(.din(w_dff_B_6JIsAdm45_1),.dout(w_dff_B_9jo6SD158_1),.clk(gclk));
	jdff dff_B_zRaMeYca5_1(.din(w_dff_B_9jo6SD158_1),.dout(w_dff_B_zRaMeYca5_1),.clk(gclk));
	jdff dff_B_rpHuyIUg3_1(.din(w_dff_B_zRaMeYca5_1),.dout(w_dff_B_rpHuyIUg3_1),.clk(gclk));
	jdff dff_B_HbSSAAja9_1(.din(w_dff_B_rpHuyIUg3_1),.dout(w_dff_B_HbSSAAja9_1),.clk(gclk));
	jdff dff_B_0znk2DEo2_1(.din(w_dff_B_HbSSAAja9_1),.dout(w_dff_B_0znk2DEo2_1),.clk(gclk));
	jdff dff_B_uHQTjcxB3_1(.din(w_dff_B_0znk2DEo2_1),.dout(w_dff_B_uHQTjcxB3_1),.clk(gclk));
	jdff dff_B_5SPzbTGA3_1(.din(w_dff_B_uHQTjcxB3_1),.dout(w_dff_B_5SPzbTGA3_1),.clk(gclk));
	jdff dff_B_j8pjpo9R2_1(.din(w_dff_B_5SPzbTGA3_1),.dout(w_dff_B_j8pjpo9R2_1),.clk(gclk));
	jdff dff_B_kpQP77Kr2_1(.din(w_dff_B_j8pjpo9R2_1),.dout(w_dff_B_kpQP77Kr2_1),.clk(gclk));
	jdff dff_B_IFgWrum80_1(.din(w_dff_B_kpQP77Kr2_1),.dout(w_dff_B_IFgWrum80_1),.clk(gclk));
	jdff dff_B_hL3LG6ve1_1(.din(n452),.dout(w_dff_B_hL3LG6ve1_1),.clk(gclk));
	jdff dff_B_MLkfyhYU5_1(.din(w_dff_B_hL3LG6ve1_1),.dout(w_dff_B_MLkfyhYU5_1),.clk(gclk));
	jdff dff_B_BaIaZgFE3_1(.din(w_dff_B_MLkfyhYU5_1),.dout(w_dff_B_BaIaZgFE3_1),.clk(gclk));
	jdff dff_B_75WEGCHR1_1(.din(w_dff_B_BaIaZgFE3_1),.dout(w_dff_B_75WEGCHR1_1),.clk(gclk));
	jdff dff_B_1uv7rtZ97_1(.din(w_dff_B_75WEGCHR1_1),.dout(w_dff_B_1uv7rtZ97_1),.clk(gclk));
	jdff dff_B_tT19Tmhp3_1(.din(w_dff_B_1uv7rtZ97_1),.dout(w_dff_B_tT19Tmhp3_1),.clk(gclk));
	jdff dff_B_OFGr9D4e7_1(.din(w_dff_B_tT19Tmhp3_1),.dout(w_dff_B_OFGr9D4e7_1),.clk(gclk));
	jdff dff_B_zQ3WILTG6_1(.din(w_dff_B_OFGr9D4e7_1),.dout(w_dff_B_zQ3WILTG6_1),.clk(gclk));
	jdff dff_B_rPoMADEC8_1(.din(w_dff_B_zQ3WILTG6_1),.dout(w_dff_B_rPoMADEC8_1),.clk(gclk));
	jdff dff_B_WY1oUXNV4_1(.din(w_dff_B_rPoMADEC8_1),.dout(w_dff_B_WY1oUXNV4_1),.clk(gclk));
	jdff dff_B_4JHhzcGh9_1(.din(w_dff_B_WY1oUXNV4_1),.dout(w_dff_B_4JHhzcGh9_1),.clk(gclk));
	jdff dff_B_B5oNP1057_1(.din(w_dff_B_4JHhzcGh9_1),.dout(w_dff_B_B5oNP1057_1),.clk(gclk));
	jdff dff_B_3gks9b4i8_1(.din(w_dff_B_B5oNP1057_1),.dout(w_dff_B_3gks9b4i8_1),.clk(gclk));
	jdff dff_B_1ckkkLVM2_1(.din(w_dff_B_3gks9b4i8_1),.dout(w_dff_B_1ckkkLVM2_1),.clk(gclk));
	jdff dff_B_7JVYq7Mk8_1(.din(w_dff_B_1ckkkLVM2_1),.dout(w_dff_B_7JVYq7Mk8_1),.clk(gclk));
	jdff dff_B_ObFOKFSt2_1(.din(w_dff_B_7JVYq7Mk8_1),.dout(w_dff_B_ObFOKFSt2_1),.clk(gclk));
	jdff dff_B_N9xsphSB1_1(.din(w_dff_B_ObFOKFSt2_1),.dout(w_dff_B_N9xsphSB1_1),.clk(gclk));
	jdff dff_B_Fs67pSzw2_1(.din(w_dff_B_N9xsphSB1_1),.dout(w_dff_B_Fs67pSzw2_1),.clk(gclk));
	jdff dff_B_TdIJWCCK2_1(.din(w_dff_B_Fs67pSzw2_1),.dout(w_dff_B_TdIJWCCK2_1),.clk(gclk));
	jdff dff_B_34XUerzc0_1(.din(w_dff_B_TdIJWCCK2_1),.dout(w_dff_B_34XUerzc0_1),.clk(gclk));
	jdff dff_B_HQdnTf2A0_1(.din(w_dff_B_34XUerzc0_1),.dout(w_dff_B_HQdnTf2A0_1),.clk(gclk));
	jdff dff_B_HuzeMcf21_1(.din(w_dff_B_HQdnTf2A0_1),.dout(w_dff_B_HuzeMcf21_1),.clk(gclk));
	jdff dff_B_1YffoFRi6_1(.din(w_dff_B_HuzeMcf21_1),.dout(w_dff_B_1YffoFRi6_1),.clk(gclk));
	jdff dff_B_7yiP9aLU6_1(.din(w_dff_B_1YffoFRi6_1),.dout(w_dff_B_7yiP9aLU6_1),.clk(gclk));
	jdff dff_B_uEJ6x5EK0_1(.din(w_dff_B_7yiP9aLU6_1),.dout(w_dff_B_uEJ6x5EK0_1),.clk(gclk));
	jdff dff_B_3Kb2MUQu2_1(.din(w_dff_B_uEJ6x5EK0_1),.dout(w_dff_B_3Kb2MUQu2_1),.clk(gclk));
	jdff dff_B_gSd35X2k7_1(.din(w_dff_B_3Kb2MUQu2_1),.dout(w_dff_B_gSd35X2k7_1),.clk(gclk));
	jdff dff_B_agLT5Mwy1_1(.din(w_dff_B_gSd35X2k7_1),.dout(w_dff_B_agLT5Mwy1_1),.clk(gclk));
	jdff dff_B_xIMHMpsd0_1(.din(w_dff_B_agLT5Mwy1_1),.dout(w_dff_B_xIMHMpsd0_1),.clk(gclk));
	jdff dff_B_EX4MsRm61_1(.din(w_dff_B_xIMHMpsd0_1),.dout(w_dff_B_EX4MsRm61_1),.clk(gclk));
	jdff dff_B_3p8ppx9t4_1(.din(n530),.dout(w_dff_B_3p8ppx9t4_1),.clk(gclk));
	jdff dff_B_fxhoKKHk4_1(.din(w_dff_B_3p8ppx9t4_1),.dout(w_dff_B_fxhoKKHk4_1),.clk(gclk));
	jdff dff_B_zDZM7NoD7_1(.din(w_dff_B_fxhoKKHk4_1),.dout(w_dff_B_zDZM7NoD7_1),.clk(gclk));
	jdff dff_B_Rp9MfLq09_1(.din(w_dff_B_zDZM7NoD7_1),.dout(w_dff_B_Rp9MfLq09_1),.clk(gclk));
	jdff dff_B_R9PHrWSQ6_1(.din(w_dff_B_Rp9MfLq09_1),.dout(w_dff_B_R9PHrWSQ6_1),.clk(gclk));
	jdff dff_B_4kLT5PFC5_1(.din(w_dff_B_R9PHrWSQ6_1),.dout(w_dff_B_4kLT5PFC5_1),.clk(gclk));
	jdff dff_B_O5TH56fR5_1(.din(w_dff_B_4kLT5PFC5_1),.dout(w_dff_B_O5TH56fR5_1),.clk(gclk));
	jdff dff_B_vfzUTUFM7_1(.din(w_dff_B_O5TH56fR5_1),.dout(w_dff_B_vfzUTUFM7_1),.clk(gclk));
	jdff dff_B_zvgPJBZK6_1(.din(w_dff_B_vfzUTUFM7_1),.dout(w_dff_B_zvgPJBZK6_1),.clk(gclk));
	jdff dff_B_nkxQ0gpm5_1(.din(w_dff_B_zvgPJBZK6_1),.dout(w_dff_B_nkxQ0gpm5_1),.clk(gclk));
	jdff dff_B_EBR7MLPw5_1(.din(w_dff_B_nkxQ0gpm5_1),.dout(w_dff_B_EBR7MLPw5_1),.clk(gclk));
	jdff dff_B_srhPxAMg8_1(.din(w_dff_B_EBR7MLPw5_1),.dout(w_dff_B_srhPxAMg8_1),.clk(gclk));
	jdff dff_B_WSXMOyrr6_1(.din(w_dff_B_srhPxAMg8_1),.dout(w_dff_B_WSXMOyrr6_1),.clk(gclk));
	jdff dff_B_ojdXWzes0_1(.din(w_dff_B_WSXMOyrr6_1),.dout(w_dff_B_ojdXWzes0_1),.clk(gclk));
	jdff dff_B_nYSBzpuP9_1(.din(w_dff_B_ojdXWzes0_1),.dout(w_dff_B_nYSBzpuP9_1),.clk(gclk));
	jdff dff_B_ZmSne4aQ9_1(.din(w_dff_B_nYSBzpuP9_1),.dout(w_dff_B_ZmSne4aQ9_1),.clk(gclk));
	jdff dff_B_tNebJp1A7_1(.din(w_dff_B_ZmSne4aQ9_1),.dout(w_dff_B_tNebJp1A7_1),.clk(gclk));
	jdff dff_B_M3dJ2zW73_1(.din(w_dff_B_tNebJp1A7_1),.dout(w_dff_B_M3dJ2zW73_1),.clk(gclk));
	jdff dff_B_K7wUEF2I0_1(.din(w_dff_B_M3dJ2zW73_1),.dout(w_dff_B_K7wUEF2I0_1),.clk(gclk));
	jdff dff_B_0AoavkzU9_1(.din(w_dff_B_K7wUEF2I0_1),.dout(w_dff_B_0AoavkzU9_1),.clk(gclk));
	jdff dff_B_fCzMoOLC1_1(.din(w_dff_B_0AoavkzU9_1),.dout(w_dff_B_fCzMoOLC1_1),.clk(gclk));
	jdff dff_B_0UaRtaB64_1(.din(w_dff_B_fCzMoOLC1_1),.dout(w_dff_B_0UaRtaB64_1),.clk(gclk));
	jdff dff_B_2NxIlVfb1_1(.din(w_dff_B_0UaRtaB64_1),.dout(w_dff_B_2NxIlVfb1_1),.clk(gclk));
	jdff dff_B_mSUjF4GK0_1(.din(w_dff_B_2NxIlVfb1_1),.dout(w_dff_B_mSUjF4GK0_1),.clk(gclk));
	jdff dff_B_b53IuW9w5_1(.din(w_dff_B_mSUjF4GK0_1),.dout(w_dff_B_b53IuW9w5_1),.clk(gclk));
	jdff dff_B_29gJcb3l1_1(.din(w_dff_B_b53IuW9w5_1),.dout(w_dff_B_29gJcb3l1_1),.clk(gclk));
	jdff dff_B_cLYYZ00k1_1(.din(w_dff_B_29gJcb3l1_1),.dout(w_dff_B_cLYYZ00k1_1),.clk(gclk));
	jdff dff_B_JIXTNkLI7_1(.din(w_dff_B_cLYYZ00k1_1),.dout(w_dff_B_JIXTNkLI7_1),.clk(gclk));
	jdff dff_B_UW2U5ROp9_1(.din(w_dff_B_JIXTNkLI7_1),.dout(w_dff_B_UW2U5ROp9_1),.clk(gclk));
	jdff dff_B_frlRyrlY4_1(.din(w_dff_B_UW2U5ROp9_1),.dout(w_dff_B_frlRyrlY4_1),.clk(gclk));
	jdff dff_B_9Mjys5ry7_1(.din(w_dff_B_frlRyrlY4_1),.dout(w_dff_B_9Mjys5ry7_1),.clk(gclk));
	jdff dff_B_idv9ebLc1_1(.din(w_dff_B_9Mjys5ry7_1),.dout(w_dff_B_idv9ebLc1_1),.clk(gclk));
	jdff dff_B_pnCMdMee4_1(.din(w_dff_B_idv9ebLc1_1),.dout(w_dff_B_pnCMdMee4_1),.clk(gclk));
	jdff dff_B_ddCYsK5h7_1(.din(n615),.dout(w_dff_B_ddCYsK5h7_1),.clk(gclk));
	jdff dff_B_4z9tfpSV2_1(.din(w_dff_B_ddCYsK5h7_1),.dout(w_dff_B_4z9tfpSV2_1),.clk(gclk));
	jdff dff_B_8Onkcvdh3_1(.din(w_dff_B_4z9tfpSV2_1),.dout(w_dff_B_8Onkcvdh3_1),.clk(gclk));
	jdff dff_B_mtf9P8PM2_1(.din(w_dff_B_8Onkcvdh3_1),.dout(w_dff_B_mtf9P8PM2_1),.clk(gclk));
	jdff dff_B_nBpGjsSK1_1(.din(w_dff_B_mtf9P8PM2_1),.dout(w_dff_B_nBpGjsSK1_1),.clk(gclk));
	jdff dff_B_BfZGTwG56_1(.din(w_dff_B_nBpGjsSK1_1),.dout(w_dff_B_BfZGTwG56_1),.clk(gclk));
	jdff dff_B_tNJjdQ0I7_1(.din(w_dff_B_BfZGTwG56_1),.dout(w_dff_B_tNJjdQ0I7_1),.clk(gclk));
	jdff dff_B_zs2J7dza5_1(.din(w_dff_B_tNJjdQ0I7_1),.dout(w_dff_B_zs2J7dza5_1),.clk(gclk));
	jdff dff_B_1OXU5V3c8_1(.din(w_dff_B_zs2J7dza5_1),.dout(w_dff_B_1OXU5V3c8_1),.clk(gclk));
	jdff dff_B_Vn73s0514_1(.din(w_dff_B_1OXU5V3c8_1),.dout(w_dff_B_Vn73s0514_1),.clk(gclk));
	jdff dff_B_7wbDTtQ59_1(.din(w_dff_B_Vn73s0514_1),.dout(w_dff_B_7wbDTtQ59_1),.clk(gclk));
	jdff dff_B_73Dquhxd4_1(.din(w_dff_B_7wbDTtQ59_1),.dout(w_dff_B_73Dquhxd4_1),.clk(gclk));
	jdff dff_B_i95YsMrf5_1(.din(w_dff_B_73Dquhxd4_1),.dout(w_dff_B_i95YsMrf5_1),.clk(gclk));
	jdff dff_B_iA3P04ht0_1(.din(w_dff_B_i95YsMrf5_1),.dout(w_dff_B_iA3P04ht0_1),.clk(gclk));
	jdff dff_B_D8gh3Ruy1_1(.din(w_dff_B_iA3P04ht0_1),.dout(w_dff_B_D8gh3Ruy1_1),.clk(gclk));
	jdff dff_B_yky5UjuC0_1(.din(w_dff_B_D8gh3Ruy1_1),.dout(w_dff_B_yky5UjuC0_1),.clk(gclk));
	jdff dff_B_2kNdDtiR9_1(.din(w_dff_B_yky5UjuC0_1),.dout(w_dff_B_2kNdDtiR9_1),.clk(gclk));
	jdff dff_B_iV5peYyX9_1(.din(w_dff_B_2kNdDtiR9_1),.dout(w_dff_B_iV5peYyX9_1),.clk(gclk));
	jdff dff_B_bsa4ROoh9_1(.din(w_dff_B_iV5peYyX9_1),.dout(w_dff_B_bsa4ROoh9_1),.clk(gclk));
	jdff dff_B_x0GZNjDs1_1(.din(w_dff_B_bsa4ROoh9_1),.dout(w_dff_B_x0GZNjDs1_1),.clk(gclk));
	jdff dff_B_SmWZzYXj4_1(.din(w_dff_B_x0GZNjDs1_1),.dout(w_dff_B_SmWZzYXj4_1),.clk(gclk));
	jdff dff_B_XV0VQKRM7_1(.din(w_dff_B_SmWZzYXj4_1),.dout(w_dff_B_XV0VQKRM7_1),.clk(gclk));
	jdff dff_B_yhEWxIyq7_1(.din(w_dff_B_XV0VQKRM7_1),.dout(w_dff_B_yhEWxIyq7_1),.clk(gclk));
	jdff dff_B_RrWDctnL6_1(.din(w_dff_B_yhEWxIyq7_1),.dout(w_dff_B_RrWDctnL6_1),.clk(gclk));
	jdff dff_B_PluXWITn0_1(.din(w_dff_B_RrWDctnL6_1),.dout(w_dff_B_PluXWITn0_1),.clk(gclk));
	jdff dff_B_8wW7V9P29_1(.din(w_dff_B_PluXWITn0_1),.dout(w_dff_B_8wW7V9P29_1),.clk(gclk));
	jdff dff_B_1ouMGPOL5_1(.din(w_dff_B_8wW7V9P29_1),.dout(w_dff_B_1ouMGPOL5_1),.clk(gclk));
	jdff dff_B_j8SJs5rv6_1(.din(w_dff_B_1ouMGPOL5_1),.dout(w_dff_B_j8SJs5rv6_1),.clk(gclk));
	jdff dff_B_MWqaKIe18_1(.din(w_dff_B_j8SJs5rv6_1),.dout(w_dff_B_MWqaKIe18_1),.clk(gclk));
	jdff dff_B_YDf0bTE60_1(.din(w_dff_B_MWqaKIe18_1),.dout(w_dff_B_YDf0bTE60_1),.clk(gclk));
	jdff dff_B_t31VFgcK7_1(.din(w_dff_B_YDf0bTE60_1),.dout(w_dff_B_t31VFgcK7_1),.clk(gclk));
	jdff dff_B_q5vUMTHS7_1(.din(w_dff_B_t31VFgcK7_1),.dout(w_dff_B_q5vUMTHS7_1),.clk(gclk));
	jdff dff_B_TBpCQkxo8_1(.din(w_dff_B_q5vUMTHS7_1),.dout(w_dff_B_TBpCQkxo8_1),.clk(gclk));
	jdff dff_B_Fq5TI8J04_1(.din(w_dff_B_TBpCQkxo8_1),.dout(w_dff_B_Fq5TI8J04_1),.clk(gclk));
	jdff dff_B_vSmBcOzN5_1(.din(w_dff_B_Fq5TI8J04_1),.dout(w_dff_B_vSmBcOzN5_1),.clk(gclk));
	jdff dff_B_55BBytC33_1(.din(w_dff_B_vSmBcOzN5_1),.dout(w_dff_B_55BBytC33_1),.clk(gclk));
	jdff dff_B_9I11JogR9_1(.din(n707),.dout(w_dff_B_9I11JogR9_1),.clk(gclk));
	jdff dff_B_AczLivBM5_1(.din(w_dff_B_9I11JogR9_1),.dout(w_dff_B_AczLivBM5_1),.clk(gclk));
	jdff dff_B_6UpP73mP7_1(.din(w_dff_B_AczLivBM5_1),.dout(w_dff_B_6UpP73mP7_1),.clk(gclk));
	jdff dff_B_qqD2Z0GD4_1(.din(w_dff_B_6UpP73mP7_1),.dout(w_dff_B_qqD2Z0GD4_1),.clk(gclk));
	jdff dff_B_aKmwxaI15_1(.din(w_dff_B_qqD2Z0GD4_1),.dout(w_dff_B_aKmwxaI15_1),.clk(gclk));
	jdff dff_B_QWwkQPb75_1(.din(w_dff_B_aKmwxaI15_1),.dout(w_dff_B_QWwkQPb75_1),.clk(gclk));
	jdff dff_B_0X2NQNbV7_1(.din(w_dff_B_QWwkQPb75_1),.dout(w_dff_B_0X2NQNbV7_1),.clk(gclk));
	jdff dff_B_jn8UXZli3_1(.din(w_dff_B_0X2NQNbV7_1),.dout(w_dff_B_jn8UXZli3_1),.clk(gclk));
	jdff dff_B_c1wNrggv4_1(.din(w_dff_B_jn8UXZli3_1),.dout(w_dff_B_c1wNrggv4_1),.clk(gclk));
	jdff dff_B_MITQI8gI8_1(.din(w_dff_B_c1wNrggv4_1),.dout(w_dff_B_MITQI8gI8_1),.clk(gclk));
	jdff dff_B_ObkCXsxe1_1(.din(w_dff_B_MITQI8gI8_1),.dout(w_dff_B_ObkCXsxe1_1),.clk(gclk));
	jdff dff_B_SWQIp7Rq1_1(.din(w_dff_B_ObkCXsxe1_1),.dout(w_dff_B_SWQIp7Rq1_1),.clk(gclk));
	jdff dff_B_roRCwGpq1_1(.din(w_dff_B_SWQIp7Rq1_1),.dout(w_dff_B_roRCwGpq1_1),.clk(gclk));
	jdff dff_B_PRyxs9Dj8_1(.din(w_dff_B_roRCwGpq1_1),.dout(w_dff_B_PRyxs9Dj8_1),.clk(gclk));
	jdff dff_B_iBKZ7qDt8_1(.din(w_dff_B_PRyxs9Dj8_1),.dout(w_dff_B_iBKZ7qDt8_1),.clk(gclk));
	jdff dff_B_K23hHub09_1(.din(w_dff_B_iBKZ7qDt8_1),.dout(w_dff_B_K23hHub09_1),.clk(gclk));
	jdff dff_B_P2U5OV9H9_1(.din(w_dff_B_K23hHub09_1),.dout(w_dff_B_P2U5OV9H9_1),.clk(gclk));
	jdff dff_B_eueJfIIM9_1(.din(w_dff_B_P2U5OV9H9_1),.dout(w_dff_B_eueJfIIM9_1),.clk(gclk));
	jdff dff_B_kot1wLEQ6_1(.din(w_dff_B_eueJfIIM9_1),.dout(w_dff_B_kot1wLEQ6_1),.clk(gclk));
	jdff dff_B_2yBF3vGT2_1(.din(w_dff_B_kot1wLEQ6_1),.dout(w_dff_B_2yBF3vGT2_1),.clk(gclk));
	jdff dff_B_2MrJYv3v0_1(.din(w_dff_B_2yBF3vGT2_1),.dout(w_dff_B_2MrJYv3v0_1),.clk(gclk));
	jdff dff_B_gzHQXFjs7_1(.din(w_dff_B_2MrJYv3v0_1),.dout(w_dff_B_gzHQXFjs7_1),.clk(gclk));
	jdff dff_B_6lrXfArB8_1(.din(w_dff_B_gzHQXFjs7_1),.dout(w_dff_B_6lrXfArB8_1),.clk(gclk));
	jdff dff_B_WgenlHKS4_1(.din(w_dff_B_6lrXfArB8_1),.dout(w_dff_B_WgenlHKS4_1),.clk(gclk));
	jdff dff_B_ogke7o653_1(.din(w_dff_B_WgenlHKS4_1),.dout(w_dff_B_ogke7o653_1),.clk(gclk));
	jdff dff_B_AKE6WBgO2_1(.din(w_dff_B_ogke7o653_1),.dout(w_dff_B_AKE6WBgO2_1),.clk(gclk));
	jdff dff_B_6JcvkoBn3_1(.din(w_dff_B_AKE6WBgO2_1),.dout(w_dff_B_6JcvkoBn3_1),.clk(gclk));
	jdff dff_B_qjWchHdH6_1(.din(w_dff_B_6JcvkoBn3_1),.dout(w_dff_B_qjWchHdH6_1),.clk(gclk));
	jdff dff_B_MOYeTtWB8_1(.din(w_dff_B_qjWchHdH6_1),.dout(w_dff_B_MOYeTtWB8_1),.clk(gclk));
	jdff dff_B_Y08ZnuLG5_1(.din(w_dff_B_MOYeTtWB8_1),.dout(w_dff_B_Y08ZnuLG5_1),.clk(gclk));
	jdff dff_B_71asyolI3_1(.din(w_dff_B_Y08ZnuLG5_1),.dout(w_dff_B_71asyolI3_1),.clk(gclk));
	jdff dff_B_D3qyxekF7_1(.din(w_dff_B_71asyolI3_1),.dout(w_dff_B_D3qyxekF7_1),.clk(gclk));
	jdff dff_B_aG0sMuV34_1(.din(w_dff_B_D3qyxekF7_1),.dout(w_dff_B_aG0sMuV34_1),.clk(gclk));
	jdff dff_B_B5hEKQXo3_1(.din(w_dff_B_aG0sMuV34_1),.dout(w_dff_B_B5hEKQXo3_1),.clk(gclk));
	jdff dff_B_GG58iKfq2_1(.din(w_dff_B_B5hEKQXo3_1),.dout(w_dff_B_GG58iKfq2_1),.clk(gclk));
	jdff dff_B_Xzqg8oJW5_1(.din(w_dff_B_GG58iKfq2_1),.dout(w_dff_B_Xzqg8oJW5_1),.clk(gclk));
	jdff dff_B_wga2OkXR9_1(.din(w_dff_B_Xzqg8oJW5_1),.dout(w_dff_B_wga2OkXR9_1),.clk(gclk));
	jdff dff_B_cZs1tC6j0_1(.din(w_dff_B_wga2OkXR9_1),.dout(w_dff_B_cZs1tC6j0_1),.clk(gclk));
	jdff dff_B_9PkQ9nLG0_1(.din(w_dff_B_cZs1tC6j0_1),.dout(w_dff_B_9PkQ9nLG0_1),.clk(gclk));
	jdff dff_B_UOySr02X9_1(.din(n806),.dout(w_dff_B_UOySr02X9_1),.clk(gclk));
	jdff dff_B_xGqX2sE21_1(.din(w_dff_B_UOySr02X9_1),.dout(w_dff_B_xGqX2sE21_1),.clk(gclk));
	jdff dff_B_hIGWddNj8_1(.din(w_dff_B_xGqX2sE21_1),.dout(w_dff_B_hIGWddNj8_1),.clk(gclk));
	jdff dff_B_tBfiJ1sl4_1(.din(w_dff_B_hIGWddNj8_1),.dout(w_dff_B_tBfiJ1sl4_1),.clk(gclk));
	jdff dff_B_zzDAoTbl5_1(.din(w_dff_B_tBfiJ1sl4_1),.dout(w_dff_B_zzDAoTbl5_1),.clk(gclk));
	jdff dff_B_gHVAWJCW3_1(.din(w_dff_B_zzDAoTbl5_1),.dout(w_dff_B_gHVAWJCW3_1),.clk(gclk));
	jdff dff_B_WJFtzMZc2_1(.din(w_dff_B_gHVAWJCW3_1),.dout(w_dff_B_WJFtzMZc2_1),.clk(gclk));
	jdff dff_B_xwIMkggk6_1(.din(w_dff_B_WJFtzMZc2_1),.dout(w_dff_B_xwIMkggk6_1),.clk(gclk));
	jdff dff_B_QSLkstkU3_1(.din(w_dff_B_xwIMkggk6_1),.dout(w_dff_B_QSLkstkU3_1),.clk(gclk));
	jdff dff_B_T1fAoUum7_1(.din(w_dff_B_QSLkstkU3_1),.dout(w_dff_B_T1fAoUum7_1),.clk(gclk));
	jdff dff_B_dmQa6sMh3_1(.din(w_dff_B_T1fAoUum7_1),.dout(w_dff_B_dmQa6sMh3_1),.clk(gclk));
	jdff dff_B_vr3m0T0t7_1(.din(w_dff_B_dmQa6sMh3_1),.dout(w_dff_B_vr3m0T0t7_1),.clk(gclk));
	jdff dff_B_vGHD0Xx13_1(.din(w_dff_B_vr3m0T0t7_1),.dout(w_dff_B_vGHD0Xx13_1),.clk(gclk));
	jdff dff_B_W1TAUOEO5_1(.din(w_dff_B_vGHD0Xx13_1),.dout(w_dff_B_W1TAUOEO5_1),.clk(gclk));
	jdff dff_B_7WD94D5C1_1(.din(w_dff_B_W1TAUOEO5_1),.dout(w_dff_B_7WD94D5C1_1),.clk(gclk));
	jdff dff_B_yN4pr8wP4_1(.din(w_dff_B_7WD94D5C1_1),.dout(w_dff_B_yN4pr8wP4_1),.clk(gclk));
	jdff dff_B_nTaNbPTO9_1(.din(w_dff_B_yN4pr8wP4_1),.dout(w_dff_B_nTaNbPTO9_1),.clk(gclk));
	jdff dff_B_Wcuhr3UH6_1(.din(w_dff_B_nTaNbPTO9_1),.dout(w_dff_B_Wcuhr3UH6_1),.clk(gclk));
	jdff dff_B_1XCLyNpe8_1(.din(w_dff_B_Wcuhr3UH6_1),.dout(w_dff_B_1XCLyNpe8_1),.clk(gclk));
	jdff dff_B_lFU5vpFS0_1(.din(w_dff_B_1XCLyNpe8_1),.dout(w_dff_B_lFU5vpFS0_1),.clk(gclk));
	jdff dff_B_GJR6hA603_1(.din(w_dff_B_lFU5vpFS0_1),.dout(w_dff_B_GJR6hA603_1),.clk(gclk));
	jdff dff_B_bY96qWr99_1(.din(w_dff_B_GJR6hA603_1),.dout(w_dff_B_bY96qWr99_1),.clk(gclk));
	jdff dff_B_kuFOyRvF2_1(.din(w_dff_B_bY96qWr99_1),.dout(w_dff_B_kuFOyRvF2_1),.clk(gclk));
	jdff dff_B_5njfu8GU9_1(.din(w_dff_B_kuFOyRvF2_1),.dout(w_dff_B_5njfu8GU9_1),.clk(gclk));
	jdff dff_B_XhcR2aI06_1(.din(w_dff_B_5njfu8GU9_1),.dout(w_dff_B_XhcR2aI06_1),.clk(gclk));
	jdff dff_B_PYlWTWKm4_1(.din(w_dff_B_XhcR2aI06_1),.dout(w_dff_B_PYlWTWKm4_1),.clk(gclk));
	jdff dff_B_czH6LOmf5_1(.din(w_dff_B_PYlWTWKm4_1),.dout(w_dff_B_czH6LOmf5_1),.clk(gclk));
	jdff dff_B_q6H1cXHd1_1(.din(w_dff_B_czH6LOmf5_1),.dout(w_dff_B_q6H1cXHd1_1),.clk(gclk));
	jdff dff_B_GxMtINvE2_1(.din(w_dff_B_q6H1cXHd1_1),.dout(w_dff_B_GxMtINvE2_1),.clk(gclk));
	jdff dff_B_M3T1LsCC7_1(.din(w_dff_B_GxMtINvE2_1),.dout(w_dff_B_M3T1LsCC7_1),.clk(gclk));
	jdff dff_B_K47AOfHv3_1(.din(w_dff_B_M3T1LsCC7_1),.dout(w_dff_B_K47AOfHv3_1),.clk(gclk));
	jdff dff_B_xiPhMNUX8_1(.din(w_dff_B_K47AOfHv3_1),.dout(w_dff_B_xiPhMNUX8_1),.clk(gclk));
	jdff dff_B_P7WUDUBO1_1(.din(w_dff_B_xiPhMNUX8_1),.dout(w_dff_B_P7WUDUBO1_1),.clk(gclk));
	jdff dff_B_pUbvCtGT7_1(.din(w_dff_B_P7WUDUBO1_1),.dout(w_dff_B_pUbvCtGT7_1),.clk(gclk));
	jdff dff_B_ca9BPqXR7_1(.din(w_dff_B_pUbvCtGT7_1),.dout(w_dff_B_ca9BPqXR7_1),.clk(gclk));
	jdff dff_B_KBceVWwJ8_1(.din(w_dff_B_ca9BPqXR7_1),.dout(w_dff_B_KBceVWwJ8_1),.clk(gclk));
	jdff dff_B_XNQTM6Mn1_1(.din(w_dff_B_KBceVWwJ8_1),.dout(w_dff_B_XNQTM6Mn1_1),.clk(gclk));
	jdff dff_B_yMcaZczD9_1(.din(w_dff_B_XNQTM6Mn1_1),.dout(w_dff_B_yMcaZczD9_1),.clk(gclk));
	jdff dff_B_s4E0WcHW3_1(.din(w_dff_B_yMcaZczD9_1),.dout(w_dff_B_s4E0WcHW3_1),.clk(gclk));
	jdff dff_B_dUWNQoQB4_1(.din(w_dff_B_s4E0WcHW3_1),.dout(w_dff_B_dUWNQoQB4_1),.clk(gclk));
	jdff dff_B_kwbDSW4F8_1(.din(w_dff_B_dUWNQoQB4_1),.dout(w_dff_B_kwbDSW4F8_1),.clk(gclk));
	jdff dff_B_mW8Cwltp4_1(.din(w_dff_B_kwbDSW4F8_1),.dout(w_dff_B_mW8Cwltp4_1),.clk(gclk));
	jdff dff_B_7zYdlvs98_0(.din(n1296),.dout(w_dff_B_7zYdlvs98_0),.clk(gclk));
	jdff dff_B_7EpvMSVl5_1(.din(n1811),.dout(w_dff_B_7EpvMSVl5_1),.clk(gclk));
	jdff dff_B_T6QCaNef3_1(.din(w_dff_B_7EpvMSVl5_1),.dout(w_dff_B_T6QCaNef3_1),.clk(gclk));
	jdff dff_B_3XDMxnoE8_1(.din(w_dff_B_T6QCaNef3_1),.dout(w_dff_B_3XDMxnoE8_1),.clk(gclk));
	jdff dff_B_kPASAC0t9_1(.din(w_dff_B_3XDMxnoE8_1),.dout(w_dff_B_kPASAC0t9_1),.clk(gclk));
	jdff dff_B_bjPfQZns6_1(.din(w_dff_B_kPASAC0t9_1),.dout(w_dff_B_bjPfQZns6_1),.clk(gclk));
	jdff dff_B_nKcYsWBE6_1(.din(w_dff_B_bjPfQZns6_1),.dout(w_dff_B_nKcYsWBE6_1),.clk(gclk));
	jdff dff_B_SksbWreh9_1(.din(w_dff_B_nKcYsWBE6_1),.dout(w_dff_B_SksbWreh9_1),.clk(gclk));
	jdff dff_B_Ya9DTWMv0_1(.din(w_dff_B_SksbWreh9_1),.dout(w_dff_B_Ya9DTWMv0_1),.clk(gclk));
	jdff dff_B_mtOLx1JO5_1(.din(w_dff_B_Ya9DTWMv0_1),.dout(w_dff_B_mtOLx1JO5_1),.clk(gclk));
	jdff dff_B_3zryJO885_1(.din(w_dff_B_mtOLx1JO5_1),.dout(w_dff_B_3zryJO885_1),.clk(gclk));
	jdff dff_B_FPGRGM5T4_1(.din(w_dff_B_3zryJO885_1),.dout(w_dff_B_FPGRGM5T4_1),.clk(gclk));
	jdff dff_B_A6LMD9Hy5_1(.din(w_dff_B_FPGRGM5T4_1),.dout(w_dff_B_A6LMD9Hy5_1),.clk(gclk));
	jdff dff_B_eSTj5NJB6_1(.din(w_dff_B_A6LMD9Hy5_1),.dout(w_dff_B_eSTj5NJB6_1),.clk(gclk));
	jdff dff_B_yjNaL4ch6_1(.din(w_dff_B_eSTj5NJB6_1),.dout(w_dff_B_yjNaL4ch6_1),.clk(gclk));
	jdff dff_B_phOQFaYs1_1(.din(w_dff_B_yjNaL4ch6_1),.dout(w_dff_B_phOQFaYs1_1),.clk(gclk));
	jdff dff_B_sKBpYG7w6_0(.din(n1819),.dout(w_dff_B_sKBpYG7w6_0),.clk(gclk));
	jdff dff_B_c7PyV10g3_0(.din(w_dff_B_sKBpYG7w6_0),.dout(w_dff_B_c7PyV10g3_0),.clk(gclk));
	jdff dff_B_zlCXqYP15_0(.din(w_dff_B_c7PyV10g3_0),.dout(w_dff_B_zlCXqYP15_0),.clk(gclk));
	jdff dff_B_1m7bE9rQ8_0(.din(w_dff_B_zlCXqYP15_0),.dout(w_dff_B_1m7bE9rQ8_0),.clk(gclk));
	jdff dff_B_xobmftXj2_0(.din(w_dff_B_1m7bE9rQ8_0),.dout(w_dff_B_xobmftXj2_0),.clk(gclk));
	jdff dff_B_PIwlu7vU0_0(.din(w_dff_B_xobmftXj2_0),.dout(w_dff_B_PIwlu7vU0_0),.clk(gclk));
	jdff dff_B_Jfgx368K5_0(.din(w_dff_B_PIwlu7vU0_0),.dout(w_dff_B_Jfgx368K5_0),.clk(gclk));
	jdff dff_B_R9dJDjgQ8_0(.din(w_dff_B_Jfgx368K5_0),.dout(w_dff_B_R9dJDjgQ8_0),.clk(gclk));
	jdff dff_B_OSBjIakL5_0(.din(w_dff_B_R9dJDjgQ8_0),.dout(w_dff_B_OSBjIakL5_0),.clk(gclk));
	jdff dff_B_nsM6fSXT6_0(.din(w_dff_B_OSBjIakL5_0),.dout(w_dff_B_nsM6fSXT6_0),.clk(gclk));
	jdff dff_B_Y2HbigHG2_0(.din(w_dff_B_nsM6fSXT6_0),.dout(w_dff_B_Y2HbigHG2_0),.clk(gclk));
	jdff dff_B_QYDhjXC85_0(.din(w_dff_B_Y2HbigHG2_0),.dout(w_dff_B_QYDhjXC85_0),.clk(gclk));
	jdff dff_B_u8BV5SUB4_0(.din(w_dff_B_QYDhjXC85_0),.dout(w_dff_B_u8BV5SUB4_0),.clk(gclk));
	jdff dff_A_OGLZbC4T0_0(.dout(w_n1818_0[0]),.din(w_dff_A_OGLZbC4T0_0),.clk(gclk));
	jdff dff_A_fZtf3Zqj6_0(.dout(w_dff_A_OGLZbC4T0_0),.din(w_dff_A_fZtf3Zqj6_0),.clk(gclk));
	jdff dff_A_Hmu1dZPq4_0(.dout(w_dff_A_fZtf3Zqj6_0),.din(w_dff_A_Hmu1dZPq4_0),.clk(gclk));
	jdff dff_A_2BJdVJ2X9_0(.dout(w_dff_A_Hmu1dZPq4_0),.din(w_dff_A_2BJdVJ2X9_0),.clk(gclk));
	jdff dff_A_FVkfFLj19_0(.dout(w_dff_A_2BJdVJ2X9_0),.din(w_dff_A_FVkfFLj19_0),.clk(gclk));
	jdff dff_A_olTvgeWK7_0(.dout(w_dff_A_FVkfFLj19_0),.din(w_dff_A_olTvgeWK7_0),.clk(gclk));
	jdff dff_A_Dxu63sbT3_0(.dout(w_dff_A_olTvgeWK7_0),.din(w_dff_A_Dxu63sbT3_0),.clk(gclk));
	jdff dff_A_H1MmSlWn2_0(.dout(w_dff_A_Dxu63sbT3_0),.din(w_dff_A_H1MmSlWn2_0),.clk(gclk));
	jdff dff_A_u0HMtG4L4_0(.dout(w_dff_A_H1MmSlWn2_0),.din(w_dff_A_u0HMtG4L4_0),.clk(gclk));
	jdff dff_A_Yk6WJghu5_0(.dout(w_dff_A_u0HMtG4L4_0),.din(w_dff_A_Yk6WJghu5_0),.clk(gclk));
	jdff dff_A_oURrr8Qc5_0(.dout(w_dff_A_Yk6WJghu5_0),.din(w_dff_A_oURrr8Qc5_0),.clk(gclk));
	jdff dff_A_5J9vILk98_0(.dout(w_dff_A_oURrr8Qc5_0),.din(w_dff_A_5J9vILk98_0),.clk(gclk));
	jdff dff_A_aLp7Z5QE0_0(.dout(w_dff_A_5J9vILk98_0),.din(w_dff_A_aLp7Z5QE0_0),.clk(gclk));
	jdff dff_A_5WGFEFAr1_0(.dout(w_dff_A_aLp7Z5QE0_0),.din(w_dff_A_5WGFEFAr1_0),.clk(gclk));
	jdff dff_B_d36Qvtmv9_1(.din(n1808),.dout(w_dff_B_d36Qvtmv9_1),.clk(gclk));
	jdff dff_B_ZdHPZkjT0_1(.din(w_dff_B_d36Qvtmv9_1),.dout(w_dff_B_ZdHPZkjT0_1),.clk(gclk));
	jdff dff_B_pbjukx3p3_2(.din(n1807),.dout(w_dff_B_pbjukx3p3_2),.clk(gclk));
	jdff dff_B_BnpMevp12_2(.din(w_dff_B_pbjukx3p3_2),.dout(w_dff_B_BnpMevp12_2),.clk(gclk));
	jdff dff_B_BgibgsJp5_2(.din(w_dff_B_BnpMevp12_2),.dout(w_dff_B_BgibgsJp5_2),.clk(gclk));
	jdff dff_B_FgbljkLo3_2(.din(w_dff_B_BgibgsJp5_2),.dout(w_dff_B_FgbljkLo3_2),.clk(gclk));
	jdff dff_B_RuJO5MXl4_2(.din(w_dff_B_FgbljkLo3_2),.dout(w_dff_B_RuJO5MXl4_2),.clk(gclk));
	jdff dff_B_aAH60p9E8_2(.din(w_dff_B_RuJO5MXl4_2),.dout(w_dff_B_aAH60p9E8_2),.clk(gclk));
	jdff dff_B_wZ6Naiyz7_2(.din(w_dff_B_aAH60p9E8_2),.dout(w_dff_B_wZ6Naiyz7_2),.clk(gclk));
	jdff dff_B_3irCt1cS4_2(.din(w_dff_B_wZ6Naiyz7_2),.dout(w_dff_B_3irCt1cS4_2),.clk(gclk));
	jdff dff_B_r2CbHWer7_2(.din(w_dff_B_3irCt1cS4_2),.dout(w_dff_B_r2CbHWer7_2),.clk(gclk));
	jdff dff_B_FEZZN7fx9_2(.din(w_dff_B_r2CbHWer7_2),.dout(w_dff_B_FEZZN7fx9_2),.clk(gclk));
	jdff dff_B_dOxPNwOr3_2(.din(w_dff_B_FEZZN7fx9_2),.dout(w_dff_B_dOxPNwOr3_2),.clk(gclk));
	jdff dff_B_bcl5B0Ji2_2(.din(w_dff_B_dOxPNwOr3_2),.dout(w_dff_B_bcl5B0Ji2_2),.clk(gclk));
	jdff dff_B_g5nXW3zj7_2(.din(w_dff_B_bcl5B0Ji2_2),.dout(w_dff_B_g5nXW3zj7_2),.clk(gclk));
	jdff dff_B_LsPfb9yV0_2(.din(w_dff_B_g5nXW3zj7_2),.dout(w_dff_B_LsPfb9yV0_2),.clk(gclk));
	jdff dff_B_37eVJ1G91_2(.din(w_dff_B_LsPfb9yV0_2),.dout(w_dff_B_37eVJ1G91_2),.clk(gclk));
	jdff dff_B_JSDHdnHv4_2(.din(w_dff_B_37eVJ1G91_2),.dout(w_dff_B_JSDHdnHv4_2),.clk(gclk));
	jdff dff_B_89sVl6iy5_2(.din(w_dff_B_JSDHdnHv4_2),.dout(w_dff_B_89sVl6iy5_2),.clk(gclk));
	jdff dff_B_7jTaEjpM3_2(.din(w_dff_B_89sVl6iy5_2),.dout(w_dff_B_7jTaEjpM3_2),.clk(gclk));
	jdff dff_B_wrrgvrQ67_2(.din(w_dff_B_7jTaEjpM3_2),.dout(w_dff_B_wrrgvrQ67_2),.clk(gclk));
	jdff dff_B_NCl24oB17_2(.din(w_dff_B_wrrgvrQ67_2),.dout(w_dff_B_NCl24oB17_2),.clk(gclk));
	jdff dff_B_49jATq0G1_2(.din(w_dff_B_NCl24oB17_2),.dout(w_dff_B_49jATq0G1_2),.clk(gclk));
	jdff dff_B_Qq1c6G4n8_2(.din(w_dff_B_49jATq0G1_2),.dout(w_dff_B_Qq1c6G4n8_2),.clk(gclk));
	jdff dff_B_2yg5L7XW3_2(.din(w_dff_B_Qq1c6G4n8_2),.dout(w_dff_B_2yg5L7XW3_2),.clk(gclk));
	jdff dff_B_afq3mQ3G2_2(.din(w_dff_B_2yg5L7XW3_2),.dout(w_dff_B_afq3mQ3G2_2),.clk(gclk));
	jdff dff_B_xPiheAAy0_2(.din(w_dff_B_afq3mQ3G2_2),.dout(w_dff_B_xPiheAAy0_2),.clk(gclk));
	jdff dff_B_eW3s00fe8_2(.din(w_dff_B_xPiheAAy0_2),.dout(w_dff_B_eW3s00fe8_2),.clk(gclk));
	jdff dff_B_1pw1a6SK8_2(.din(w_dff_B_eW3s00fe8_2),.dout(w_dff_B_1pw1a6SK8_2),.clk(gclk));
	jdff dff_B_8rfYcsID7_2(.din(w_dff_B_1pw1a6SK8_2),.dout(w_dff_B_8rfYcsID7_2),.clk(gclk));
	jdff dff_B_rQvKxmFw5_2(.din(w_dff_B_8rfYcsID7_2),.dout(w_dff_B_rQvKxmFw5_2),.clk(gclk));
	jdff dff_B_famZFcKB5_2(.din(w_dff_B_rQvKxmFw5_2),.dout(w_dff_B_famZFcKB5_2),.clk(gclk));
	jdff dff_B_tbFlF8UB1_2(.din(w_dff_B_famZFcKB5_2),.dout(w_dff_B_tbFlF8UB1_2),.clk(gclk));
	jdff dff_B_qMdlOkgv7_2(.din(w_dff_B_tbFlF8UB1_2),.dout(w_dff_B_qMdlOkgv7_2),.clk(gclk));
	jdff dff_B_3RX2ORUq0_2(.din(w_dff_B_qMdlOkgv7_2),.dout(w_dff_B_3RX2ORUq0_2),.clk(gclk));
	jdff dff_B_mv831Y7I2_2(.din(w_dff_B_3RX2ORUq0_2),.dout(w_dff_B_mv831Y7I2_2),.clk(gclk));
	jdff dff_B_tBPOmc2m2_2(.din(w_dff_B_mv831Y7I2_2),.dout(w_dff_B_tBPOmc2m2_2),.clk(gclk));
	jdff dff_B_OtSpjFUH6_2(.din(w_dff_B_tBPOmc2m2_2),.dout(w_dff_B_OtSpjFUH6_2),.clk(gclk));
	jdff dff_B_n30ZIvjc2_2(.din(w_dff_B_OtSpjFUH6_2),.dout(w_dff_B_n30ZIvjc2_2),.clk(gclk));
	jdff dff_B_VGVCOS1k9_2(.din(w_dff_B_n30ZIvjc2_2),.dout(w_dff_B_VGVCOS1k9_2),.clk(gclk));
	jdff dff_B_JIQOLr3L4_2(.din(w_dff_B_VGVCOS1k9_2),.dout(w_dff_B_JIQOLr3L4_2),.clk(gclk));
	jdff dff_B_VjmxtvCP9_2(.din(w_dff_B_JIQOLr3L4_2),.dout(w_dff_B_VjmxtvCP9_2),.clk(gclk));
	jdff dff_B_uJsCxzc15_2(.din(w_dff_B_VjmxtvCP9_2),.dout(w_dff_B_uJsCxzc15_2),.clk(gclk));
	jdff dff_B_2wuuOQNM6_2(.din(w_dff_B_uJsCxzc15_2),.dout(w_dff_B_2wuuOQNM6_2),.clk(gclk));
	jdff dff_B_ea6nszm69_2(.din(w_dff_B_2wuuOQNM6_2),.dout(w_dff_B_ea6nszm69_2),.clk(gclk));
	jdff dff_B_zHSg5EZA8_2(.din(w_dff_B_ea6nszm69_2),.dout(w_dff_B_zHSg5EZA8_2),.clk(gclk));
	jdff dff_B_5o2CEteu9_2(.din(w_dff_B_zHSg5EZA8_2),.dout(w_dff_B_5o2CEteu9_2),.clk(gclk));
	jdff dff_B_AdjPIj2j3_2(.din(w_dff_B_5o2CEteu9_2),.dout(w_dff_B_AdjPIj2j3_2),.clk(gclk));
	jdff dff_B_1KKQIqhO4_2(.din(w_dff_B_AdjPIj2j3_2),.dout(w_dff_B_1KKQIqhO4_2),.clk(gclk));
	jdff dff_B_GuUGSFkC1_2(.din(w_dff_B_1KKQIqhO4_2),.dout(w_dff_B_GuUGSFkC1_2),.clk(gclk));
	jdff dff_B_7QK4NaCx4_2(.din(w_dff_B_GuUGSFkC1_2),.dout(w_dff_B_7QK4NaCx4_2),.clk(gclk));
	jdff dff_B_LzPIU7lD6_2(.din(w_dff_B_7QK4NaCx4_2),.dout(w_dff_B_LzPIU7lD6_2),.clk(gclk));
	jdff dff_B_MAsQbvKE2_2(.din(w_dff_B_LzPIU7lD6_2),.dout(w_dff_B_MAsQbvKE2_2),.clk(gclk));
	jdff dff_B_G9WrQf9w3_2(.din(w_dff_B_MAsQbvKE2_2),.dout(w_dff_B_G9WrQf9w3_2),.clk(gclk));
	jdff dff_B_EIQDCpFu4_2(.din(w_dff_B_G9WrQf9w3_2),.dout(w_dff_B_EIQDCpFu4_2),.clk(gclk));
	jdff dff_B_244B1Wex5_2(.din(w_dff_B_EIQDCpFu4_2),.dout(w_dff_B_244B1Wex5_2),.clk(gclk));
	jdff dff_B_1FS8p3sa6_2(.din(w_dff_B_244B1Wex5_2),.dout(w_dff_B_1FS8p3sa6_2),.clk(gclk));
	jdff dff_B_5XV3zr7M5_2(.din(w_dff_B_1FS8p3sa6_2),.dout(w_dff_B_5XV3zr7M5_2),.clk(gclk));
	jdff dff_B_U2lBJJDX5_2(.din(w_dff_B_5XV3zr7M5_2),.dout(w_dff_B_U2lBJJDX5_2),.clk(gclk));
	jdff dff_B_Bix3zfp38_1(.din(n1814),.dout(w_dff_B_Bix3zfp38_1),.clk(gclk));
	jdff dff_B_HUKiIKo39_1(.din(w_dff_B_Bix3zfp38_1),.dout(w_dff_B_HUKiIKo39_1),.clk(gclk));
	jdff dff_B_X7tXwIFQ1_1(.din(w_dff_B_HUKiIKo39_1),.dout(w_dff_B_X7tXwIFQ1_1),.clk(gclk));
	jdff dff_B_jupwEDHS3_1(.din(w_dff_B_X7tXwIFQ1_1),.dout(w_dff_B_jupwEDHS3_1),.clk(gclk));
	jdff dff_B_HxGId1660_1(.din(w_dff_B_jupwEDHS3_1),.dout(w_dff_B_HxGId1660_1),.clk(gclk));
	jdff dff_B_3UXBHJQS2_1(.din(w_dff_B_HxGId1660_1),.dout(w_dff_B_3UXBHJQS2_1),.clk(gclk));
	jdff dff_B_Jvmy94ni8_1(.din(w_dff_B_3UXBHJQS2_1),.dout(w_dff_B_Jvmy94ni8_1),.clk(gclk));
	jdff dff_B_0sWA1UK89_1(.din(w_dff_B_Jvmy94ni8_1),.dout(w_dff_B_0sWA1UK89_1),.clk(gclk));
	jdff dff_B_0ZwEKrgK9_1(.din(w_dff_B_0sWA1UK89_1),.dout(w_dff_B_0ZwEKrgK9_1),.clk(gclk));
	jdff dff_B_11YPltti4_1(.din(w_dff_B_0ZwEKrgK9_1),.dout(w_dff_B_11YPltti4_1),.clk(gclk));
	jdff dff_B_OSoyy2EH8_1(.din(w_dff_B_11YPltti4_1),.dout(w_dff_B_OSoyy2EH8_1),.clk(gclk));
	jdff dff_B_YPELLd6n6_1(.din(w_dff_B_OSoyy2EH8_1),.dout(w_dff_B_YPELLd6n6_1),.clk(gclk));
	jdff dff_B_Qw1tMa5V8_1(.din(w_dff_B_YPELLd6n6_1),.dout(w_dff_B_Qw1tMa5V8_1),.clk(gclk));
	jdff dff_B_3lOqtsjK5_0(.din(n1815),.dout(w_dff_B_3lOqtsjK5_0),.clk(gclk));
	jdff dff_B_FJJJ8L2U5_0(.din(w_dff_B_3lOqtsjK5_0),.dout(w_dff_B_FJJJ8L2U5_0),.clk(gclk));
	jdff dff_B_DC7NPE3h0_0(.din(w_dff_B_FJJJ8L2U5_0),.dout(w_dff_B_DC7NPE3h0_0),.clk(gclk));
	jdff dff_B_yC3cHug76_0(.din(w_dff_B_DC7NPE3h0_0),.dout(w_dff_B_yC3cHug76_0),.clk(gclk));
	jdff dff_B_RwwjpeXH2_0(.din(w_dff_B_yC3cHug76_0),.dout(w_dff_B_RwwjpeXH2_0),.clk(gclk));
	jdff dff_B_nc4HFfsQ2_0(.din(w_dff_B_RwwjpeXH2_0),.dout(w_dff_B_nc4HFfsQ2_0),.clk(gclk));
	jdff dff_B_Qfijb8HS2_0(.din(w_dff_B_nc4HFfsQ2_0),.dout(w_dff_B_Qfijb8HS2_0),.clk(gclk));
	jdff dff_B_Qc9AZV7I7_0(.din(w_dff_B_Qfijb8HS2_0),.dout(w_dff_B_Qc9AZV7I7_0),.clk(gclk));
	jdff dff_B_WksdNB8K3_0(.din(w_dff_B_Qc9AZV7I7_0),.dout(w_dff_B_WksdNB8K3_0),.clk(gclk));
	jdff dff_B_IjTrR2oE5_0(.din(w_dff_B_WksdNB8K3_0),.dout(w_dff_B_IjTrR2oE5_0),.clk(gclk));
	jdff dff_B_Xfrab0YJ1_0(.din(w_dff_B_IjTrR2oE5_0),.dout(w_dff_B_Xfrab0YJ1_0),.clk(gclk));
	jdff dff_B_0VGTcHsx1_0(.din(w_dff_B_Xfrab0YJ1_0),.dout(w_dff_B_0VGTcHsx1_0),.clk(gclk));
	jdff dff_A_pTqzBYu31_1(.dout(w_n1805_0[1]),.din(w_dff_A_pTqzBYu31_1),.clk(gclk));
	jdff dff_A_4FePtVCr2_1(.dout(w_dff_A_pTqzBYu31_1),.din(w_dff_A_4FePtVCr2_1),.clk(gclk));
	jdff dff_A_5F7kZV4w2_1(.dout(w_dff_A_4FePtVCr2_1),.din(w_dff_A_5F7kZV4w2_1),.clk(gclk));
	jdff dff_A_kvi5W9hh3_1(.dout(w_dff_A_5F7kZV4w2_1),.din(w_dff_A_kvi5W9hh3_1),.clk(gclk));
	jdff dff_A_OkshN4R91_1(.dout(w_dff_A_kvi5W9hh3_1),.din(w_dff_A_OkshN4R91_1),.clk(gclk));
	jdff dff_A_yYiUzrlC1_1(.dout(w_dff_A_OkshN4R91_1),.din(w_dff_A_yYiUzrlC1_1),.clk(gclk));
	jdff dff_A_RMdtxuCP6_1(.dout(w_dff_A_yYiUzrlC1_1),.din(w_dff_A_RMdtxuCP6_1),.clk(gclk));
	jdff dff_A_a1q6uYAC1_1(.dout(w_dff_A_RMdtxuCP6_1),.din(w_dff_A_a1q6uYAC1_1),.clk(gclk));
	jdff dff_A_WQMxp8Gs8_1(.dout(w_dff_A_a1q6uYAC1_1),.din(w_dff_A_WQMxp8Gs8_1),.clk(gclk));
	jdff dff_A_7ZYaLpCK1_1(.dout(w_dff_A_WQMxp8Gs8_1),.din(w_dff_A_7ZYaLpCK1_1),.clk(gclk));
	jdff dff_A_bYfNsD6v3_1(.dout(w_dff_A_7ZYaLpCK1_1),.din(w_dff_A_bYfNsD6v3_1),.clk(gclk));
	jdff dff_A_FhOaXYDI7_1(.dout(w_dff_A_bYfNsD6v3_1),.din(w_dff_A_FhOaXYDI7_1),.clk(gclk));
	jdff dff_A_U4LD1zzq3_1(.dout(w_dff_A_FhOaXYDI7_1),.din(w_dff_A_U4LD1zzq3_1),.clk(gclk));
	jdff dff_B_8v3WQY2V7_1(.din(n1790),.dout(w_dff_B_8v3WQY2V7_1),.clk(gclk));
	jdff dff_B_eKIm7TT43_1(.din(w_dff_B_8v3WQY2V7_1),.dout(w_dff_B_eKIm7TT43_1),.clk(gclk));
	jdff dff_B_qDpLUSQJ5_1(.din(w_dff_B_eKIm7TT43_1),.dout(w_dff_B_qDpLUSQJ5_1),.clk(gclk));
	jdff dff_B_SG9rV6eE5_1(.din(w_dff_B_qDpLUSQJ5_1),.dout(w_dff_B_SG9rV6eE5_1),.clk(gclk));
	jdff dff_B_TDhwSEQc4_1(.din(w_dff_B_SG9rV6eE5_1),.dout(w_dff_B_TDhwSEQc4_1),.clk(gclk));
	jdff dff_B_LotP9No29_1(.din(w_dff_B_TDhwSEQc4_1),.dout(w_dff_B_LotP9No29_1),.clk(gclk));
	jdff dff_B_WE1PAy2l5_1(.din(w_dff_B_LotP9No29_1),.dout(w_dff_B_WE1PAy2l5_1),.clk(gclk));
	jdff dff_B_rLXX39jf1_1(.din(w_dff_B_WE1PAy2l5_1),.dout(w_dff_B_rLXX39jf1_1),.clk(gclk));
	jdff dff_B_sBibyQ3Y8_1(.din(w_dff_B_rLXX39jf1_1),.dout(w_dff_B_sBibyQ3Y8_1),.clk(gclk));
	jdff dff_B_GDYGvwbl7_1(.din(w_dff_B_sBibyQ3Y8_1),.dout(w_dff_B_GDYGvwbl7_1),.clk(gclk));
	jdff dff_B_xhSQ2eNV9_1(.din(w_dff_B_GDYGvwbl7_1),.dout(w_dff_B_xhSQ2eNV9_1),.clk(gclk));
	jdff dff_B_dMx9PzRk5_1(.din(w_dff_B_xhSQ2eNV9_1),.dout(w_dff_B_dMx9PzRk5_1),.clk(gclk));
	jdff dff_B_riXXVnAg6_1(.din(w_dff_B_dMx9PzRk5_1),.dout(w_dff_B_riXXVnAg6_1),.clk(gclk));
	jdff dff_B_jNxbnMLI3_0(.din(n1791),.dout(w_dff_B_jNxbnMLI3_0),.clk(gclk));
	jdff dff_B_GwVkRXTt3_0(.din(w_dff_B_jNxbnMLI3_0),.dout(w_dff_B_GwVkRXTt3_0),.clk(gclk));
	jdff dff_B_MLG8SSbY3_0(.din(w_dff_B_GwVkRXTt3_0),.dout(w_dff_B_MLG8SSbY3_0),.clk(gclk));
	jdff dff_B_2jeVg1IQ7_0(.din(w_dff_B_MLG8SSbY3_0),.dout(w_dff_B_2jeVg1IQ7_0),.clk(gclk));
	jdff dff_B_Jp3TWmxC8_0(.din(w_dff_B_2jeVg1IQ7_0),.dout(w_dff_B_Jp3TWmxC8_0),.clk(gclk));
	jdff dff_B_p58vol1v2_0(.din(w_dff_B_Jp3TWmxC8_0),.dout(w_dff_B_p58vol1v2_0),.clk(gclk));
	jdff dff_B_jerW2Aff7_0(.din(w_dff_B_p58vol1v2_0),.dout(w_dff_B_jerW2Aff7_0),.clk(gclk));
	jdff dff_B_15y0Hs482_0(.din(w_dff_B_jerW2Aff7_0),.dout(w_dff_B_15y0Hs482_0),.clk(gclk));
	jdff dff_B_PWWwDA3Q3_0(.din(w_dff_B_15y0Hs482_0),.dout(w_dff_B_PWWwDA3Q3_0),.clk(gclk));
	jdff dff_B_ZRk8IG8r4_0(.din(w_dff_B_PWWwDA3Q3_0),.dout(w_dff_B_ZRk8IG8r4_0),.clk(gclk));
	jdff dff_B_zLU5isVA4_0(.din(w_dff_B_ZRk8IG8r4_0),.dout(w_dff_B_zLU5isVA4_0),.clk(gclk));
	jdff dff_B_wTDV2G8q2_0(.din(w_dff_B_zLU5isVA4_0),.dout(w_dff_B_wTDV2G8q2_0),.clk(gclk));
	jdff dff_A_pBhS1Xgx7_1(.dout(w_n1786_0[1]),.din(w_dff_A_pBhS1Xgx7_1),.clk(gclk));
	jdff dff_A_kiFRoxr33_1(.dout(w_dff_A_pBhS1Xgx7_1),.din(w_dff_A_kiFRoxr33_1),.clk(gclk));
	jdff dff_A_YuBI7OAj3_1(.dout(w_dff_A_kiFRoxr33_1),.din(w_dff_A_YuBI7OAj3_1),.clk(gclk));
	jdff dff_A_FcpZtgMN4_1(.dout(w_dff_A_YuBI7OAj3_1),.din(w_dff_A_FcpZtgMN4_1),.clk(gclk));
	jdff dff_A_2y1Mngn19_1(.dout(w_dff_A_FcpZtgMN4_1),.din(w_dff_A_2y1Mngn19_1),.clk(gclk));
	jdff dff_A_OK9QNA8d5_1(.dout(w_dff_A_2y1Mngn19_1),.din(w_dff_A_OK9QNA8d5_1),.clk(gclk));
	jdff dff_A_QgzdG5GI1_1(.dout(w_dff_A_OK9QNA8d5_1),.din(w_dff_A_QgzdG5GI1_1),.clk(gclk));
	jdff dff_A_yNYEbi4V6_1(.dout(w_dff_A_QgzdG5GI1_1),.din(w_dff_A_yNYEbi4V6_1),.clk(gclk));
	jdff dff_A_M27VZ3eY9_1(.dout(w_dff_A_yNYEbi4V6_1),.din(w_dff_A_M27VZ3eY9_1),.clk(gclk));
	jdff dff_A_9xyC4LpG8_1(.dout(w_dff_A_M27VZ3eY9_1),.din(w_dff_A_9xyC4LpG8_1),.clk(gclk));
	jdff dff_A_LgJ6lgWz5_1(.dout(w_dff_A_9xyC4LpG8_1),.din(w_dff_A_LgJ6lgWz5_1),.clk(gclk));
	jdff dff_A_BYSrS0wx7_1(.dout(w_dff_A_LgJ6lgWz5_1),.din(w_dff_A_BYSrS0wx7_1),.clk(gclk));
	jdff dff_A_X2uFtJnt5_1(.dout(w_dff_A_BYSrS0wx7_1),.din(w_dff_A_X2uFtJnt5_1),.clk(gclk));
	jdff dff_B_pFoFlUWE0_1(.din(n1764),.dout(w_dff_B_pFoFlUWE0_1),.clk(gclk));
	jdff dff_B_r1PrxLTi4_1(.din(w_dff_B_pFoFlUWE0_1),.dout(w_dff_B_r1PrxLTi4_1),.clk(gclk));
	jdff dff_B_BPO2fSng8_1(.din(w_dff_B_r1PrxLTi4_1),.dout(w_dff_B_BPO2fSng8_1),.clk(gclk));
	jdff dff_B_m6704ISZ0_1(.din(w_dff_B_BPO2fSng8_1),.dout(w_dff_B_m6704ISZ0_1),.clk(gclk));
	jdff dff_B_hiHOPFuQ5_1(.din(w_dff_B_m6704ISZ0_1),.dout(w_dff_B_hiHOPFuQ5_1),.clk(gclk));
	jdff dff_B_BzHZeDtJ7_1(.din(w_dff_B_hiHOPFuQ5_1),.dout(w_dff_B_BzHZeDtJ7_1),.clk(gclk));
	jdff dff_B_NbJYKeo75_1(.din(w_dff_B_BzHZeDtJ7_1),.dout(w_dff_B_NbJYKeo75_1),.clk(gclk));
	jdff dff_B_bqk360Sm5_1(.din(w_dff_B_NbJYKeo75_1),.dout(w_dff_B_bqk360Sm5_1),.clk(gclk));
	jdff dff_B_73g31No99_1(.din(w_dff_B_bqk360Sm5_1),.dout(w_dff_B_73g31No99_1),.clk(gclk));
	jdff dff_B_8EcVF8Sf7_1(.din(w_dff_B_73g31No99_1),.dout(w_dff_B_8EcVF8Sf7_1),.clk(gclk));
	jdff dff_B_S398jecD7_1(.din(w_dff_B_8EcVF8Sf7_1),.dout(w_dff_B_S398jecD7_1),.clk(gclk));
	jdff dff_B_DYBrGr1S5_1(.din(w_dff_B_S398jecD7_1),.dout(w_dff_B_DYBrGr1S5_1),.clk(gclk));
	jdff dff_B_LvUM34K53_1(.din(w_dff_B_DYBrGr1S5_1),.dout(w_dff_B_LvUM34K53_1),.clk(gclk));
	jdff dff_B_SkGD4B6a3_0(.din(n1765),.dout(w_dff_B_SkGD4B6a3_0),.clk(gclk));
	jdff dff_B_7WXAFeFZ0_0(.din(w_dff_B_SkGD4B6a3_0),.dout(w_dff_B_7WXAFeFZ0_0),.clk(gclk));
	jdff dff_B_J5P78yHT3_0(.din(w_dff_B_7WXAFeFZ0_0),.dout(w_dff_B_J5P78yHT3_0),.clk(gclk));
	jdff dff_B_qHzjWNrt1_0(.din(w_dff_B_J5P78yHT3_0),.dout(w_dff_B_qHzjWNrt1_0),.clk(gclk));
	jdff dff_B_sIxquQj50_0(.din(w_dff_B_qHzjWNrt1_0),.dout(w_dff_B_sIxquQj50_0),.clk(gclk));
	jdff dff_B_wgGR5Igf0_0(.din(w_dff_B_sIxquQj50_0),.dout(w_dff_B_wgGR5Igf0_0),.clk(gclk));
	jdff dff_B_QQZ6U9yX8_0(.din(w_dff_B_wgGR5Igf0_0),.dout(w_dff_B_QQZ6U9yX8_0),.clk(gclk));
	jdff dff_B_S5Lu6qdr7_0(.din(w_dff_B_QQZ6U9yX8_0),.dout(w_dff_B_S5Lu6qdr7_0),.clk(gclk));
	jdff dff_B_7rWqxsCi8_0(.din(w_dff_B_S5Lu6qdr7_0),.dout(w_dff_B_7rWqxsCi8_0),.clk(gclk));
	jdff dff_B_w4wAMyPH7_0(.din(w_dff_B_7rWqxsCi8_0),.dout(w_dff_B_w4wAMyPH7_0),.clk(gclk));
	jdff dff_B_WOOYhY1H8_0(.din(w_dff_B_w4wAMyPH7_0),.dout(w_dff_B_WOOYhY1H8_0),.clk(gclk));
	jdff dff_B_rmZtcw0A2_0(.din(w_dff_B_WOOYhY1H8_0),.dout(w_dff_B_rmZtcw0A2_0),.clk(gclk));
	jdff dff_A_uNAV6jyP9_1(.dout(w_n1760_0[1]),.din(w_dff_A_uNAV6jyP9_1),.clk(gclk));
	jdff dff_A_rsdn4Fvf6_1(.dout(w_dff_A_uNAV6jyP9_1),.din(w_dff_A_rsdn4Fvf6_1),.clk(gclk));
	jdff dff_A_ec2cygHW9_1(.dout(w_dff_A_rsdn4Fvf6_1),.din(w_dff_A_ec2cygHW9_1),.clk(gclk));
	jdff dff_A_wP6v6v4l9_1(.dout(w_dff_A_ec2cygHW9_1),.din(w_dff_A_wP6v6v4l9_1),.clk(gclk));
	jdff dff_A_SKlKZQ3q4_1(.dout(w_dff_A_wP6v6v4l9_1),.din(w_dff_A_SKlKZQ3q4_1),.clk(gclk));
	jdff dff_A_9RjWiZKk4_1(.dout(w_dff_A_SKlKZQ3q4_1),.din(w_dff_A_9RjWiZKk4_1),.clk(gclk));
	jdff dff_A_OKriZr6j2_1(.dout(w_dff_A_9RjWiZKk4_1),.din(w_dff_A_OKriZr6j2_1),.clk(gclk));
	jdff dff_A_sSHIpeJ62_1(.dout(w_dff_A_OKriZr6j2_1),.din(w_dff_A_sSHIpeJ62_1),.clk(gclk));
	jdff dff_A_N6W14orn8_1(.dout(w_dff_A_sSHIpeJ62_1),.din(w_dff_A_N6W14orn8_1),.clk(gclk));
	jdff dff_A_wnKCvNYV1_1(.dout(w_dff_A_N6W14orn8_1),.din(w_dff_A_wnKCvNYV1_1),.clk(gclk));
	jdff dff_A_qstbFSmp5_1(.dout(w_dff_A_wnKCvNYV1_1),.din(w_dff_A_qstbFSmp5_1),.clk(gclk));
	jdff dff_A_R8FXLjzr9_1(.dout(w_dff_A_qstbFSmp5_1),.din(w_dff_A_R8FXLjzr9_1),.clk(gclk));
	jdff dff_A_vJw6EZhk6_1(.dout(w_dff_A_R8FXLjzr9_1),.din(w_dff_A_vJw6EZhk6_1),.clk(gclk));
	jdff dff_B_N9wQQJg86_1(.din(n1731),.dout(w_dff_B_N9wQQJg86_1),.clk(gclk));
	jdff dff_B_SsnF83O28_1(.din(w_dff_B_N9wQQJg86_1),.dout(w_dff_B_SsnF83O28_1),.clk(gclk));
	jdff dff_B_KW544CsX5_1(.din(w_dff_B_SsnF83O28_1),.dout(w_dff_B_KW544CsX5_1),.clk(gclk));
	jdff dff_B_TJcVgsp28_1(.din(w_dff_B_KW544CsX5_1),.dout(w_dff_B_TJcVgsp28_1),.clk(gclk));
	jdff dff_B_B5jq7bo63_1(.din(w_dff_B_TJcVgsp28_1),.dout(w_dff_B_B5jq7bo63_1),.clk(gclk));
	jdff dff_B_5bljzWBo5_1(.din(w_dff_B_B5jq7bo63_1),.dout(w_dff_B_5bljzWBo5_1),.clk(gclk));
	jdff dff_B_76f0BGGX8_1(.din(w_dff_B_5bljzWBo5_1),.dout(w_dff_B_76f0BGGX8_1),.clk(gclk));
	jdff dff_B_2bpPxMxK3_1(.din(w_dff_B_76f0BGGX8_1),.dout(w_dff_B_2bpPxMxK3_1),.clk(gclk));
	jdff dff_B_fxymJWAO4_1(.din(w_dff_B_2bpPxMxK3_1),.dout(w_dff_B_fxymJWAO4_1),.clk(gclk));
	jdff dff_B_m8Zv5k4W2_1(.din(w_dff_B_fxymJWAO4_1),.dout(w_dff_B_m8Zv5k4W2_1),.clk(gclk));
	jdff dff_B_QoVLrXGO4_1(.din(w_dff_B_m8Zv5k4W2_1),.dout(w_dff_B_QoVLrXGO4_1),.clk(gclk));
	jdff dff_B_y1tpFsAq0_1(.din(w_dff_B_QoVLrXGO4_1),.dout(w_dff_B_y1tpFsAq0_1),.clk(gclk));
	jdff dff_B_uDp8zjvm9_1(.din(w_dff_B_y1tpFsAq0_1),.dout(w_dff_B_uDp8zjvm9_1),.clk(gclk));
	jdff dff_B_E8Jt4ML90_0(.din(n1732),.dout(w_dff_B_E8Jt4ML90_0),.clk(gclk));
	jdff dff_B_XoPospA31_0(.din(w_dff_B_E8Jt4ML90_0),.dout(w_dff_B_XoPospA31_0),.clk(gclk));
	jdff dff_B_0alDVRbt3_0(.din(w_dff_B_XoPospA31_0),.dout(w_dff_B_0alDVRbt3_0),.clk(gclk));
	jdff dff_B_hYJZTyWJ0_0(.din(w_dff_B_0alDVRbt3_0),.dout(w_dff_B_hYJZTyWJ0_0),.clk(gclk));
	jdff dff_B_786EVvBB0_0(.din(w_dff_B_hYJZTyWJ0_0),.dout(w_dff_B_786EVvBB0_0),.clk(gclk));
	jdff dff_B_4OKTCQay7_0(.din(w_dff_B_786EVvBB0_0),.dout(w_dff_B_4OKTCQay7_0),.clk(gclk));
	jdff dff_B_rd3A1EDw4_0(.din(w_dff_B_4OKTCQay7_0),.dout(w_dff_B_rd3A1EDw4_0),.clk(gclk));
	jdff dff_B_Hb7hgK8W9_0(.din(w_dff_B_rd3A1EDw4_0),.dout(w_dff_B_Hb7hgK8W9_0),.clk(gclk));
	jdff dff_B_f4jijjLA5_0(.din(w_dff_B_Hb7hgK8W9_0),.dout(w_dff_B_f4jijjLA5_0),.clk(gclk));
	jdff dff_B_QawrM9Qr4_0(.din(w_dff_B_f4jijjLA5_0),.dout(w_dff_B_QawrM9Qr4_0),.clk(gclk));
	jdff dff_B_eN3dMciJ8_0(.din(w_dff_B_QawrM9Qr4_0),.dout(w_dff_B_eN3dMciJ8_0),.clk(gclk));
	jdff dff_B_DXgxM1M27_0(.din(w_dff_B_eN3dMciJ8_0),.dout(w_dff_B_DXgxM1M27_0),.clk(gclk));
	jdff dff_A_hjV3lOHx4_1(.dout(w_n1727_0[1]),.din(w_dff_A_hjV3lOHx4_1),.clk(gclk));
	jdff dff_A_NDdoCHAe9_1(.dout(w_dff_A_hjV3lOHx4_1),.din(w_dff_A_NDdoCHAe9_1),.clk(gclk));
	jdff dff_A_HW0ZDJ4t6_1(.dout(w_dff_A_NDdoCHAe9_1),.din(w_dff_A_HW0ZDJ4t6_1),.clk(gclk));
	jdff dff_A_btICl05A6_1(.dout(w_dff_A_HW0ZDJ4t6_1),.din(w_dff_A_btICl05A6_1),.clk(gclk));
	jdff dff_A_q2F8XsFO5_1(.dout(w_dff_A_btICl05A6_1),.din(w_dff_A_q2F8XsFO5_1),.clk(gclk));
	jdff dff_A_kbqibt0p1_1(.dout(w_dff_A_q2F8XsFO5_1),.din(w_dff_A_kbqibt0p1_1),.clk(gclk));
	jdff dff_A_eO1PjrBI2_1(.dout(w_dff_A_kbqibt0p1_1),.din(w_dff_A_eO1PjrBI2_1),.clk(gclk));
	jdff dff_A_czwSC3EB8_1(.dout(w_dff_A_eO1PjrBI2_1),.din(w_dff_A_czwSC3EB8_1),.clk(gclk));
	jdff dff_A_OYzVL8BR8_1(.dout(w_dff_A_czwSC3EB8_1),.din(w_dff_A_OYzVL8BR8_1),.clk(gclk));
	jdff dff_A_rOFx621m8_1(.dout(w_dff_A_OYzVL8BR8_1),.din(w_dff_A_rOFx621m8_1),.clk(gclk));
	jdff dff_A_u950MIbr0_1(.dout(w_dff_A_rOFx621m8_1),.din(w_dff_A_u950MIbr0_1),.clk(gclk));
	jdff dff_A_mbm2HHbT3_1(.dout(w_dff_A_u950MIbr0_1),.din(w_dff_A_mbm2HHbT3_1),.clk(gclk));
	jdff dff_A_Sd21jNyI9_1(.dout(w_dff_A_mbm2HHbT3_1),.din(w_dff_A_Sd21jNyI9_1),.clk(gclk));
	jdff dff_B_30yM5xKK6_1(.din(n1691),.dout(w_dff_B_30yM5xKK6_1),.clk(gclk));
	jdff dff_B_CGYZkYwP2_1(.din(w_dff_B_30yM5xKK6_1),.dout(w_dff_B_CGYZkYwP2_1),.clk(gclk));
	jdff dff_B_zr07N4Pr6_1(.din(w_dff_B_CGYZkYwP2_1),.dout(w_dff_B_zr07N4Pr6_1),.clk(gclk));
	jdff dff_B_6nE8ZbBL8_1(.din(w_dff_B_zr07N4Pr6_1),.dout(w_dff_B_6nE8ZbBL8_1),.clk(gclk));
	jdff dff_B_LGnK3gLv0_1(.din(w_dff_B_6nE8ZbBL8_1),.dout(w_dff_B_LGnK3gLv0_1),.clk(gclk));
	jdff dff_B_b31vDNQL9_1(.din(w_dff_B_LGnK3gLv0_1),.dout(w_dff_B_b31vDNQL9_1),.clk(gclk));
	jdff dff_B_weeQiOkW2_1(.din(w_dff_B_b31vDNQL9_1),.dout(w_dff_B_weeQiOkW2_1),.clk(gclk));
	jdff dff_B_cTuRbi5Y2_1(.din(w_dff_B_weeQiOkW2_1),.dout(w_dff_B_cTuRbi5Y2_1),.clk(gclk));
	jdff dff_B_H6VExGyq5_1(.din(w_dff_B_cTuRbi5Y2_1),.dout(w_dff_B_H6VExGyq5_1),.clk(gclk));
	jdff dff_B_7cOPp9976_1(.din(w_dff_B_H6VExGyq5_1),.dout(w_dff_B_7cOPp9976_1),.clk(gclk));
	jdff dff_B_lvc6ILmI6_1(.din(w_dff_B_7cOPp9976_1),.dout(w_dff_B_lvc6ILmI6_1),.clk(gclk));
	jdff dff_B_D8PRoUg86_1(.din(w_dff_B_lvc6ILmI6_1),.dout(w_dff_B_D8PRoUg86_1),.clk(gclk));
	jdff dff_B_DNx9ayef5_1(.din(w_dff_B_D8PRoUg86_1),.dout(w_dff_B_DNx9ayef5_1),.clk(gclk));
	jdff dff_B_0BLcdcqw7_0(.din(n1692),.dout(w_dff_B_0BLcdcqw7_0),.clk(gclk));
	jdff dff_B_jQCGwjLa3_0(.din(w_dff_B_0BLcdcqw7_0),.dout(w_dff_B_jQCGwjLa3_0),.clk(gclk));
	jdff dff_B_wyZRcVP01_0(.din(w_dff_B_jQCGwjLa3_0),.dout(w_dff_B_wyZRcVP01_0),.clk(gclk));
	jdff dff_B_gV5MsEzD1_0(.din(w_dff_B_wyZRcVP01_0),.dout(w_dff_B_gV5MsEzD1_0),.clk(gclk));
	jdff dff_B_DRUHyAs93_0(.din(w_dff_B_gV5MsEzD1_0),.dout(w_dff_B_DRUHyAs93_0),.clk(gclk));
	jdff dff_B_INf212I59_0(.din(w_dff_B_DRUHyAs93_0),.dout(w_dff_B_INf212I59_0),.clk(gclk));
	jdff dff_B_rsOKGopn9_0(.din(w_dff_B_INf212I59_0),.dout(w_dff_B_rsOKGopn9_0),.clk(gclk));
	jdff dff_B_j9P400kM3_0(.din(w_dff_B_rsOKGopn9_0),.dout(w_dff_B_j9P400kM3_0),.clk(gclk));
	jdff dff_B_DZNoLCJ52_0(.din(w_dff_B_j9P400kM3_0),.dout(w_dff_B_DZNoLCJ52_0),.clk(gclk));
	jdff dff_B_ucRAZtgc5_0(.din(w_dff_B_DZNoLCJ52_0),.dout(w_dff_B_ucRAZtgc5_0),.clk(gclk));
	jdff dff_B_F08mUVaJ1_0(.din(w_dff_B_ucRAZtgc5_0),.dout(w_dff_B_F08mUVaJ1_0),.clk(gclk));
	jdff dff_A_tvreZN8X1_1(.dout(w_n1689_0[1]),.din(w_dff_A_tvreZN8X1_1),.clk(gclk));
	jdff dff_A_Cn7XDjv57_1(.dout(w_dff_A_tvreZN8X1_1),.din(w_dff_A_Cn7XDjv57_1),.clk(gclk));
	jdff dff_A_4rZDInLo4_1(.dout(w_dff_A_Cn7XDjv57_1),.din(w_dff_A_4rZDInLo4_1),.clk(gclk));
	jdff dff_A_BAAoP9jH6_1(.dout(w_dff_A_4rZDInLo4_1),.din(w_dff_A_BAAoP9jH6_1),.clk(gclk));
	jdff dff_A_UWVFC1Ic5_1(.dout(w_dff_A_BAAoP9jH6_1),.din(w_dff_A_UWVFC1Ic5_1),.clk(gclk));
	jdff dff_A_79AkB2Do4_1(.dout(w_dff_A_UWVFC1Ic5_1),.din(w_dff_A_79AkB2Do4_1),.clk(gclk));
	jdff dff_A_sOjATV497_1(.dout(w_dff_A_79AkB2Do4_1),.din(w_dff_A_sOjATV497_1),.clk(gclk));
	jdff dff_A_Cat8Zylc3_1(.dout(w_dff_A_sOjATV497_1),.din(w_dff_A_Cat8Zylc3_1),.clk(gclk));
	jdff dff_A_lzvz1v0d6_1(.dout(w_dff_A_Cat8Zylc3_1),.din(w_dff_A_lzvz1v0d6_1),.clk(gclk));
	jdff dff_A_ZdZNELKh4_1(.dout(w_dff_A_lzvz1v0d6_1),.din(w_dff_A_ZdZNELKh4_1),.clk(gclk));
	jdff dff_A_7yapfgYL4_1(.dout(w_dff_A_ZdZNELKh4_1),.din(w_dff_A_7yapfgYL4_1),.clk(gclk));
	jdff dff_A_cIRgkc145_1(.dout(w_dff_A_7yapfgYL4_1),.din(w_dff_A_cIRgkc145_1),.clk(gclk));
	jdff dff_B_uWlBIvLo8_1(.din(n1643),.dout(w_dff_B_uWlBIvLo8_1),.clk(gclk));
	jdff dff_B_MgA73bY22_1(.din(w_dff_B_uWlBIvLo8_1),.dout(w_dff_B_MgA73bY22_1),.clk(gclk));
	jdff dff_B_xmXztxwm5_1(.din(w_dff_B_MgA73bY22_1),.dout(w_dff_B_xmXztxwm5_1),.clk(gclk));
	jdff dff_B_HlF8PbBy0_1(.din(w_dff_B_xmXztxwm5_1),.dout(w_dff_B_HlF8PbBy0_1),.clk(gclk));
	jdff dff_B_8W7M111H4_1(.din(w_dff_B_HlF8PbBy0_1),.dout(w_dff_B_8W7M111H4_1),.clk(gclk));
	jdff dff_B_Mdq1B7827_1(.din(w_dff_B_8W7M111H4_1),.dout(w_dff_B_Mdq1B7827_1),.clk(gclk));
	jdff dff_B_IwJzkcoX3_1(.din(w_dff_B_Mdq1B7827_1),.dout(w_dff_B_IwJzkcoX3_1),.clk(gclk));
	jdff dff_B_QvlTnmCB9_1(.din(w_dff_B_IwJzkcoX3_1),.dout(w_dff_B_QvlTnmCB9_1),.clk(gclk));
	jdff dff_B_2KfT1hEF4_1(.din(w_dff_B_QvlTnmCB9_1),.dout(w_dff_B_2KfT1hEF4_1),.clk(gclk));
	jdff dff_B_0cJZaRno9_1(.din(w_dff_B_2KfT1hEF4_1),.dout(w_dff_B_0cJZaRno9_1),.clk(gclk));
	jdff dff_B_oYoAC6kM4_1(.din(w_dff_B_0cJZaRno9_1),.dout(w_dff_B_oYoAC6kM4_1),.clk(gclk));
	jdff dff_B_s5QX8V1B0_1(.din(w_dff_B_oYoAC6kM4_1),.dout(w_dff_B_s5QX8V1B0_1),.clk(gclk));
	jdff dff_B_obngi1Mw6_0(.din(n1644),.dout(w_dff_B_obngi1Mw6_0),.clk(gclk));
	jdff dff_B_sZS5H6QN1_0(.din(w_dff_B_obngi1Mw6_0),.dout(w_dff_B_sZS5H6QN1_0),.clk(gclk));
	jdff dff_B_eILZSG073_0(.din(w_dff_B_sZS5H6QN1_0),.dout(w_dff_B_eILZSG073_0),.clk(gclk));
	jdff dff_B_7CsJF2TN9_0(.din(w_dff_B_eILZSG073_0),.dout(w_dff_B_7CsJF2TN9_0),.clk(gclk));
	jdff dff_B_sIpz9hmA9_0(.din(w_dff_B_7CsJF2TN9_0),.dout(w_dff_B_sIpz9hmA9_0),.clk(gclk));
	jdff dff_B_HrfV0fS35_0(.din(w_dff_B_sIpz9hmA9_0),.dout(w_dff_B_HrfV0fS35_0),.clk(gclk));
	jdff dff_B_CkOM9qdK4_0(.din(w_dff_B_HrfV0fS35_0),.dout(w_dff_B_CkOM9qdK4_0),.clk(gclk));
	jdff dff_B_WKxyQKDn9_0(.din(w_dff_B_CkOM9qdK4_0),.dout(w_dff_B_WKxyQKDn9_0),.clk(gclk));
	jdff dff_B_Cn15YGIz2_0(.din(w_dff_B_WKxyQKDn9_0),.dout(w_dff_B_Cn15YGIz2_0),.clk(gclk));
	jdff dff_B_0kya3YlB7_0(.din(w_dff_B_Cn15YGIz2_0),.dout(w_dff_B_0kya3YlB7_0),.clk(gclk));
	jdff dff_A_PZpdhY025_1(.dout(w_n1641_0[1]),.din(w_dff_A_PZpdhY025_1),.clk(gclk));
	jdff dff_A_2Aeeomrf3_1(.dout(w_dff_A_PZpdhY025_1),.din(w_dff_A_2Aeeomrf3_1),.clk(gclk));
	jdff dff_A_6ms3FofL1_1(.dout(w_dff_A_2Aeeomrf3_1),.din(w_dff_A_6ms3FofL1_1),.clk(gclk));
	jdff dff_A_MgxkmANA7_1(.dout(w_dff_A_6ms3FofL1_1),.din(w_dff_A_MgxkmANA7_1),.clk(gclk));
	jdff dff_A_ZnEhY6lB5_1(.dout(w_dff_A_MgxkmANA7_1),.din(w_dff_A_ZnEhY6lB5_1),.clk(gclk));
	jdff dff_A_y7GSRsIN9_1(.dout(w_dff_A_ZnEhY6lB5_1),.din(w_dff_A_y7GSRsIN9_1),.clk(gclk));
	jdff dff_A_0v9Gkyz79_1(.dout(w_dff_A_y7GSRsIN9_1),.din(w_dff_A_0v9Gkyz79_1),.clk(gclk));
	jdff dff_A_fxWq5Bfg5_1(.dout(w_dff_A_0v9Gkyz79_1),.din(w_dff_A_fxWq5Bfg5_1),.clk(gclk));
	jdff dff_A_XVYOy3fL1_1(.dout(w_dff_A_fxWq5Bfg5_1),.din(w_dff_A_XVYOy3fL1_1),.clk(gclk));
	jdff dff_A_yrIOqe3D5_1(.dout(w_dff_A_XVYOy3fL1_1),.din(w_dff_A_yrIOqe3D5_1),.clk(gclk));
	jdff dff_A_TtZdaZ396_1(.dout(w_dff_A_yrIOqe3D5_1),.din(w_dff_A_TtZdaZ396_1),.clk(gclk));
	jdff dff_B_4uJ8Bepp5_1(.din(n1588),.dout(w_dff_B_4uJ8Bepp5_1),.clk(gclk));
	jdff dff_B_AUzhealC0_1(.din(w_dff_B_4uJ8Bepp5_1),.dout(w_dff_B_AUzhealC0_1),.clk(gclk));
	jdff dff_B_S77Q3T2F2_1(.din(w_dff_B_AUzhealC0_1),.dout(w_dff_B_S77Q3T2F2_1),.clk(gclk));
	jdff dff_B_a952ppHb0_1(.din(w_dff_B_S77Q3T2F2_1),.dout(w_dff_B_a952ppHb0_1),.clk(gclk));
	jdff dff_B_PjT0Dn9s2_1(.din(w_dff_B_a952ppHb0_1),.dout(w_dff_B_PjT0Dn9s2_1),.clk(gclk));
	jdff dff_B_ijEFmXS61_1(.din(w_dff_B_PjT0Dn9s2_1),.dout(w_dff_B_ijEFmXS61_1),.clk(gclk));
	jdff dff_B_gW7xaS6U3_1(.din(w_dff_B_ijEFmXS61_1),.dout(w_dff_B_gW7xaS6U3_1),.clk(gclk));
	jdff dff_B_O2AeDvK69_1(.din(w_dff_B_gW7xaS6U3_1),.dout(w_dff_B_O2AeDvK69_1),.clk(gclk));
	jdff dff_B_8dCHLFDH7_1(.din(w_dff_B_O2AeDvK69_1),.dout(w_dff_B_8dCHLFDH7_1),.clk(gclk));
	jdff dff_B_YA4uxX2x2_1(.din(w_dff_B_8dCHLFDH7_1),.dout(w_dff_B_YA4uxX2x2_1),.clk(gclk));
	jdff dff_B_4vE1JtrY5_0(.din(n1589),.dout(w_dff_B_4vE1JtrY5_0),.clk(gclk));
	jdff dff_B_49ivluk90_0(.din(w_dff_B_4vE1JtrY5_0),.dout(w_dff_B_49ivluk90_0),.clk(gclk));
	jdff dff_B_75L79S3Z0_0(.din(w_dff_B_49ivluk90_0),.dout(w_dff_B_75L79S3Z0_0),.clk(gclk));
	jdff dff_B_Boao5wH08_0(.din(w_dff_B_75L79S3Z0_0),.dout(w_dff_B_Boao5wH08_0),.clk(gclk));
	jdff dff_B_eifM8ikB7_0(.din(w_dff_B_Boao5wH08_0),.dout(w_dff_B_eifM8ikB7_0),.clk(gclk));
	jdff dff_B_AeNyD6i78_0(.din(w_dff_B_eifM8ikB7_0),.dout(w_dff_B_AeNyD6i78_0),.clk(gclk));
	jdff dff_B_57bKYgkk5_0(.din(w_dff_B_AeNyD6i78_0),.dout(w_dff_B_57bKYgkk5_0),.clk(gclk));
	jdff dff_B_kMbvP8Ys0_0(.din(w_dff_B_57bKYgkk5_0),.dout(w_dff_B_kMbvP8Ys0_0),.clk(gclk));
	jdff dff_A_A4IqpdUQ5_1(.dout(w_n1586_0[1]),.din(w_dff_A_A4IqpdUQ5_1),.clk(gclk));
	jdff dff_A_8fL4RIXD2_1(.dout(w_dff_A_A4IqpdUQ5_1),.din(w_dff_A_8fL4RIXD2_1),.clk(gclk));
	jdff dff_A_eajauNj64_1(.dout(w_dff_A_8fL4RIXD2_1),.din(w_dff_A_eajauNj64_1),.clk(gclk));
	jdff dff_A_wspUXdpS9_1(.dout(w_dff_A_eajauNj64_1),.din(w_dff_A_wspUXdpS9_1),.clk(gclk));
	jdff dff_A_myeZBikA5_1(.dout(w_dff_A_wspUXdpS9_1),.din(w_dff_A_myeZBikA5_1),.clk(gclk));
	jdff dff_A_v4dCg3kJ4_1(.dout(w_dff_A_myeZBikA5_1),.din(w_dff_A_v4dCg3kJ4_1),.clk(gclk));
	jdff dff_A_1H3sC3Dl2_1(.dout(w_dff_A_v4dCg3kJ4_1),.din(w_dff_A_1H3sC3Dl2_1),.clk(gclk));
	jdff dff_A_eQICZcG63_1(.dout(w_dff_A_1H3sC3Dl2_1),.din(w_dff_A_eQICZcG63_1),.clk(gclk));
	jdff dff_A_UV68AmjS3_1(.dout(w_dff_A_eQICZcG63_1),.din(w_dff_A_UV68AmjS3_1),.clk(gclk));
	jdff dff_B_XdGCmkl78_1(.din(n1526),.dout(w_dff_B_XdGCmkl78_1),.clk(gclk));
	jdff dff_B_K8uoeSnC5_1(.din(w_dff_B_XdGCmkl78_1),.dout(w_dff_B_K8uoeSnC5_1),.clk(gclk));
	jdff dff_B_aN7ZBlDt2_1(.din(w_dff_B_K8uoeSnC5_1),.dout(w_dff_B_aN7ZBlDt2_1),.clk(gclk));
	jdff dff_B_wr3vF4hx2_1(.din(w_dff_B_aN7ZBlDt2_1),.dout(w_dff_B_wr3vF4hx2_1),.clk(gclk));
	jdff dff_B_Q11UU1Bz4_1(.din(w_dff_B_wr3vF4hx2_1),.dout(w_dff_B_Q11UU1Bz4_1),.clk(gclk));
	jdff dff_B_PSO2yEQ62_1(.din(w_dff_B_Q11UU1Bz4_1),.dout(w_dff_B_PSO2yEQ62_1),.clk(gclk));
	jdff dff_B_22LA1uYP2_1(.din(w_dff_B_PSO2yEQ62_1),.dout(w_dff_B_22LA1uYP2_1),.clk(gclk));
	jdff dff_B_tnRGkghO1_1(.din(w_dff_B_22LA1uYP2_1),.dout(w_dff_B_tnRGkghO1_1),.clk(gclk));
	jdff dff_B_IBPxuKjS9_0(.din(n1527),.dout(w_dff_B_IBPxuKjS9_0),.clk(gclk));
	jdff dff_B_qCi3aASs1_0(.din(w_dff_B_IBPxuKjS9_0),.dout(w_dff_B_qCi3aASs1_0),.clk(gclk));
	jdff dff_B_eIQi7tKb4_0(.din(w_dff_B_qCi3aASs1_0),.dout(w_dff_B_eIQi7tKb4_0),.clk(gclk));
	jdff dff_B_bQsmDhh81_0(.din(w_dff_B_eIQi7tKb4_0),.dout(w_dff_B_bQsmDhh81_0),.clk(gclk));
	jdff dff_B_MwJ1wSbg8_0(.din(w_dff_B_bQsmDhh81_0),.dout(w_dff_B_MwJ1wSbg8_0),.clk(gclk));
	jdff dff_B_tlSTntkM6_0(.din(w_dff_B_MwJ1wSbg8_0),.dout(w_dff_B_tlSTntkM6_0),.clk(gclk));
	jdff dff_A_3JhYv0GU8_1(.dout(w_n1524_0[1]),.din(w_dff_A_3JhYv0GU8_1),.clk(gclk));
	jdff dff_A_SxywY5UB2_1(.dout(w_dff_A_3JhYv0GU8_1),.din(w_dff_A_SxywY5UB2_1),.clk(gclk));
	jdff dff_A_f48muEoQ5_1(.dout(w_dff_A_SxywY5UB2_1),.din(w_dff_A_f48muEoQ5_1),.clk(gclk));
	jdff dff_A_XUOQDGnf4_1(.dout(w_dff_A_f48muEoQ5_1),.din(w_dff_A_XUOQDGnf4_1),.clk(gclk));
	jdff dff_A_SD3ES31H9_1(.dout(w_dff_A_XUOQDGnf4_1),.din(w_dff_A_SD3ES31H9_1),.clk(gclk));
	jdff dff_A_aYOi67Ny6_1(.dout(w_dff_A_SD3ES31H9_1),.din(w_dff_A_aYOi67Ny6_1),.clk(gclk));
	jdff dff_A_wCShQUCq8_1(.dout(w_dff_A_aYOi67Ny6_1),.din(w_dff_A_wCShQUCq8_1),.clk(gclk));
	jdff dff_B_Vufxfh1h0_1(.din(n1457),.dout(w_dff_B_Vufxfh1h0_1),.clk(gclk));
	jdff dff_B_wkuxKIox2_1(.din(w_dff_B_Vufxfh1h0_1),.dout(w_dff_B_wkuxKIox2_1),.clk(gclk));
	jdff dff_B_24U2AcJ98_1(.din(w_dff_B_wkuxKIox2_1),.dout(w_dff_B_24U2AcJ98_1),.clk(gclk));
	jdff dff_B_otp3howQ8_1(.din(w_dff_B_24U2AcJ98_1),.dout(w_dff_B_otp3howQ8_1),.clk(gclk));
	jdff dff_B_O1mc53Ql2_1(.din(w_dff_B_otp3howQ8_1),.dout(w_dff_B_O1mc53Ql2_1),.clk(gclk));
	jdff dff_B_yRWGmAue1_1(.din(w_dff_B_O1mc53Ql2_1),.dout(w_dff_B_yRWGmAue1_1),.clk(gclk));
	jdff dff_B_Jum1WBO27_1(.din(w_dff_B_yRWGmAue1_1),.dout(w_dff_B_Jum1WBO27_1),.clk(gclk));
	jdff dff_B_ZwOkEQIq9_0(.din(n1458),.dout(w_dff_B_ZwOkEQIq9_0),.clk(gclk));
	jdff dff_B_HqaMKhrT9_0(.din(w_dff_B_ZwOkEQIq9_0),.dout(w_dff_B_HqaMKhrT9_0),.clk(gclk));
	jdff dff_B_7APDhqe42_0(.din(w_dff_B_HqaMKhrT9_0),.dout(w_dff_B_7APDhqe42_0),.clk(gclk));
	jdff dff_B_IOOsdPOc2_0(.din(w_dff_B_7APDhqe42_0),.dout(w_dff_B_IOOsdPOc2_0),.clk(gclk));
	jdff dff_B_BjqKJUgd6_0(.din(w_dff_B_IOOsdPOc2_0),.dout(w_dff_B_BjqKJUgd6_0),.clk(gclk));
	jdff dff_A_stdT9izj0_1(.dout(w_n1455_0[1]),.din(w_dff_A_stdT9izj0_1),.clk(gclk));
	jdff dff_A_vDhqPUTt0_1(.dout(w_dff_A_stdT9izj0_1),.din(w_dff_A_vDhqPUTt0_1),.clk(gclk));
	jdff dff_A_oN0MRBMf9_1(.dout(w_dff_A_vDhqPUTt0_1),.din(w_dff_A_oN0MRBMf9_1),.clk(gclk));
	jdff dff_A_6l2COR606_1(.dout(w_dff_A_oN0MRBMf9_1),.din(w_dff_A_6l2COR606_1),.clk(gclk));
	jdff dff_A_eoffVhJJ4_1(.dout(w_dff_A_6l2COR606_1),.din(w_dff_A_eoffVhJJ4_1),.clk(gclk));
	jdff dff_A_CpR4vvnb3_1(.dout(w_dff_A_eoffVhJJ4_1),.din(w_dff_A_CpR4vvnb3_1),.clk(gclk));
	jdff dff_B_DRhGq0Jx3_1(.din(n1381),.dout(w_dff_B_DRhGq0Jx3_1),.clk(gclk));
	jdff dff_B_f2CfR5yF8_1(.din(w_dff_B_DRhGq0Jx3_1),.dout(w_dff_B_f2CfR5yF8_1),.clk(gclk));
	jdff dff_B_oWG9Onrk0_1(.din(w_dff_B_f2CfR5yF8_1),.dout(w_dff_B_oWG9Onrk0_1),.clk(gclk));
	jdff dff_B_SDVvdd771_1(.din(w_dff_B_oWG9Onrk0_1),.dout(w_dff_B_SDVvdd771_1),.clk(gclk));
	jdff dff_B_ZJhdyy6G9_1(.din(w_dff_B_SDVvdd771_1),.dout(w_dff_B_ZJhdyy6G9_1),.clk(gclk));
	jdff dff_B_wlGQ1Lsq0_1(.din(w_dff_B_ZJhdyy6G9_1),.dout(w_dff_B_wlGQ1Lsq0_1),.clk(gclk));
	jdff dff_B_TgsEjimH4_0(.din(n1382),.dout(w_dff_B_TgsEjimH4_0),.clk(gclk));
	jdff dff_B_qTNqAT652_0(.din(w_dff_B_TgsEjimH4_0),.dout(w_dff_B_qTNqAT652_0),.clk(gclk));
	jdff dff_B_4CJJYbYo5_0(.din(w_dff_B_qTNqAT652_0),.dout(w_dff_B_4CJJYbYo5_0),.clk(gclk));
	jdff dff_B_hVTh9bVH3_0(.din(w_dff_B_4CJJYbYo5_0),.dout(w_dff_B_hVTh9bVH3_0),.clk(gclk));
	jdff dff_A_oEnI9cUc0_1(.dout(w_n1379_0[1]),.din(w_dff_A_oEnI9cUc0_1),.clk(gclk));
	jdff dff_A_ThfkHn2S2_1(.dout(w_dff_A_oEnI9cUc0_1),.din(w_dff_A_ThfkHn2S2_1),.clk(gclk));
	jdff dff_A_y6icyVYp4_1(.dout(w_dff_A_ThfkHn2S2_1),.din(w_dff_A_y6icyVYp4_1),.clk(gclk));
	jdff dff_A_95HQoU8P0_1(.dout(w_dff_A_y6icyVYp4_1),.din(w_dff_A_95HQoU8P0_1),.clk(gclk));
	jdff dff_A_QwUZQSPN3_1(.dout(w_dff_A_95HQoU8P0_1),.din(w_dff_A_QwUZQSPN3_1),.clk(gclk));
	jdff dff_B_JYF0L2XJ8_1(.din(n1299),.dout(w_dff_B_JYF0L2XJ8_1),.clk(gclk));
	jdff dff_B_510lIA7N8_1(.din(w_dff_B_JYF0L2XJ8_1),.dout(w_dff_B_510lIA7N8_1),.clk(gclk));
	jdff dff_B_jS3TSOxf8_1(.din(w_dff_B_510lIA7N8_1),.dout(w_dff_B_jS3TSOxf8_1),.clk(gclk));
	jdff dff_A_oxewnWqe5_0(.dout(w_n1295_0[0]),.din(w_dff_A_oxewnWqe5_0),.clk(gclk));
	jdff dff_A_d5qDWqJV6_0(.dout(w_dff_A_oxewnWqe5_0),.din(w_dff_A_d5qDWqJV6_0),.clk(gclk));
	jdff dff_B_z5MYaKAx6_1(.din(n1211),.dout(w_dff_B_z5MYaKAx6_1),.clk(gclk));
	jdff dff_A_fRkJO1mJ1_0(.dout(w_n1207_0[0]),.din(w_dff_A_fRkJO1mJ1_0),.clk(gclk));
	jdff dff_B_Uj7K2SEj3_1(.din(n1113),.dout(w_dff_B_Uj7K2SEj3_1),.clk(gclk));
	jdff dff_A_4Ncw3g6H8_1(.dout(w_n1013_0[1]),.din(w_dff_A_4Ncw3g6H8_1),.clk(gclk));
	jdff dff_B_gC9Kk4D31_2(.din(n1011),.dout(w_dff_B_gC9Kk4D31_2),.clk(gclk));
	jdff dff_B_kLvZqWp66_1(.din(n908),.dout(w_dff_B_kLvZqWp66_1),.clk(gclk));
	jdff dff_A_Seyk8gfb3_0(.dout(w_n805_0[0]),.din(w_dff_A_Seyk8gfb3_0),.clk(gclk));
	jdff dff_A_1yImg40o4_0(.dout(w_dff_A_Seyk8gfb3_0),.din(w_dff_A_1yImg40o4_0),.clk(gclk));
	jdff dff_A_ozNheDmb8_0(.dout(w_dff_A_1yImg40o4_0),.din(w_dff_A_ozNheDmb8_0),.clk(gclk));
	jdff dff_A_8Oqfx7Y42_0(.dout(w_dff_A_ozNheDmb8_0),.din(w_dff_A_8Oqfx7Y42_0),.clk(gclk));
	jdff dff_A_s8vQXMGD9_0(.dout(w_dff_A_8Oqfx7Y42_0),.din(w_dff_A_s8vQXMGD9_0),.clk(gclk));
	jdff dff_A_L3jATuxM0_0(.dout(w_dff_A_s8vQXMGD9_0),.din(w_dff_A_L3jATuxM0_0),.clk(gclk));
	jdff dff_A_u3AT2OHP4_0(.dout(w_dff_A_L3jATuxM0_0),.din(w_dff_A_u3AT2OHP4_0),.clk(gclk));
	jdff dff_A_MfSNh8Kt5_0(.dout(w_dff_A_u3AT2OHP4_0),.din(w_dff_A_MfSNh8Kt5_0),.clk(gclk));
	jdff dff_A_1ShWz5oI9_0(.dout(w_dff_A_MfSNh8Kt5_0),.din(w_dff_A_1ShWz5oI9_0),.clk(gclk));
	jdff dff_A_gzcDSFxN4_0(.dout(w_dff_A_1ShWz5oI9_0),.din(w_dff_A_gzcDSFxN4_0),.clk(gclk));
	jdff dff_A_UKl2naQv9_0(.dout(w_dff_A_gzcDSFxN4_0),.din(w_dff_A_UKl2naQv9_0),.clk(gclk));
	jdff dff_A_AmdVlZ4t3_0(.dout(w_dff_A_UKl2naQv9_0),.din(w_dff_A_AmdVlZ4t3_0),.clk(gclk));
	jdff dff_A_WYQRrI7A1_0(.dout(w_dff_A_AmdVlZ4t3_0),.din(w_dff_A_WYQRrI7A1_0),.clk(gclk));
	jdff dff_A_r2uzzCPy2_0(.dout(w_dff_A_WYQRrI7A1_0),.din(w_dff_A_r2uzzCPy2_0),.clk(gclk));
	jdff dff_A_OufKW71A1_0(.dout(w_dff_A_r2uzzCPy2_0),.din(w_dff_A_OufKW71A1_0),.clk(gclk));
	jdff dff_A_PVQkZhej7_0(.dout(w_dff_A_OufKW71A1_0),.din(w_dff_A_PVQkZhej7_0),.clk(gclk));
	jdff dff_A_pauUSEtX0_0(.dout(w_dff_A_PVQkZhej7_0),.din(w_dff_A_pauUSEtX0_0),.clk(gclk));
	jdff dff_A_aN4i3XGp4_0(.dout(w_dff_A_pauUSEtX0_0),.din(w_dff_A_aN4i3XGp4_0),.clk(gclk));
	jdff dff_A_43nPrk3u9_0(.dout(w_dff_A_aN4i3XGp4_0),.din(w_dff_A_43nPrk3u9_0),.clk(gclk));
	jdff dff_A_mK81VH2X9_0(.dout(w_dff_A_43nPrk3u9_0),.din(w_dff_A_mK81VH2X9_0),.clk(gclk));
	jdff dff_A_6Zg4E4Qp6_0(.dout(w_dff_A_mK81VH2X9_0),.din(w_dff_A_6Zg4E4Qp6_0),.clk(gclk));
	jdff dff_A_yXbS2Gw17_0(.dout(w_dff_A_6Zg4E4Qp6_0),.din(w_dff_A_yXbS2Gw17_0),.clk(gclk));
	jdff dff_A_mlMGkp182_0(.dout(w_dff_A_yXbS2Gw17_0),.din(w_dff_A_mlMGkp182_0),.clk(gclk));
	jdff dff_A_58KKJxIu0_0(.dout(w_dff_A_mlMGkp182_0),.din(w_dff_A_58KKJxIu0_0),.clk(gclk));
	jdff dff_A_lqpqhx4x1_0(.dout(w_dff_A_58KKJxIu0_0),.din(w_dff_A_lqpqhx4x1_0),.clk(gclk));
	jdff dff_A_ou0a32tw9_0(.dout(w_dff_A_lqpqhx4x1_0),.din(w_dff_A_ou0a32tw9_0),.clk(gclk));
	jdff dff_A_GixbuAfL0_0(.dout(w_dff_A_ou0a32tw9_0),.din(w_dff_A_GixbuAfL0_0),.clk(gclk));
	jdff dff_A_drcFrAzD4_0(.dout(w_dff_A_GixbuAfL0_0),.din(w_dff_A_drcFrAzD4_0),.clk(gclk));
	jdff dff_A_f69hM5O12_0(.dout(w_dff_A_drcFrAzD4_0),.din(w_dff_A_f69hM5O12_0),.clk(gclk));
	jdff dff_A_NWrmpPhQ9_0(.dout(w_dff_A_f69hM5O12_0),.din(w_dff_A_NWrmpPhQ9_0),.clk(gclk));
	jdff dff_A_65twvrJE0_0(.dout(w_dff_A_NWrmpPhQ9_0),.din(w_dff_A_65twvrJE0_0),.clk(gclk));
	jdff dff_A_4foDo0V27_0(.dout(w_dff_A_65twvrJE0_0),.din(w_dff_A_4foDo0V27_0),.clk(gclk));
	jdff dff_A_VxeqP4YA0_0(.dout(w_dff_A_4foDo0V27_0),.din(w_dff_A_VxeqP4YA0_0),.clk(gclk));
	jdff dff_A_XU7sFgWb9_0(.dout(w_dff_A_VxeqP4YA0_0),.din(w_dff_A_XU7sFgWb9_0),.clk(gclk));
	jdff dff_A_3khLpKQS0_0(.dout(w_dff_A_XU7sFgWb9_0),.din(w_dff_A_3khLpKQS0_0),.clk(gclk));
	jdff dff_A_iXCDGnMZ8_0(.dout(w_dff_A_3khLpKQS0_0),.din(w_dff_A_iXCDGnMZ8_0),.clk(gclk));
	jdff dff_A_B1PvtdqP9_0(.dout(w_dff_A_iXCDGnMZ8_0),.din(w_dff_A_B1PvtdqP9_0),.clk(gclk));
	jdff dff_A_LPCfYOc87_0(.dout(w_dff_A_B1PvtdqP9_0),.din(w_dff_A_LPCfYOc87_0),.clk(gclk));
	jdff dff_A_WCJlgciS9_0(.dout(w_dff_A_LPCfYOc87_0),.din(w_dff_A_WCJlgciS9_0),.clk(gclk));
	jdff dff_A_PfgyymiN4_0(.dout(w_dff_A_WCJlgciS9_0),.din(w_dff_A_PfgyymiN4_0),.clk(gclk));
	jdff dff_A_nBHD5X532_0(.dout(w_dff_A_PfgyymiN4_0),.din(w_dff_A_nBHD5X532_0),.clk(gclk));
	jdff dff_A_uRpohZrb7_0(.dout(w_dff_A_nBHD5X532_0),.din(w_dff_A_uRpohZrb7_0),.clk(gclk));
	jdff dff_A_gsQw3Cox5_0(.dout(w_dff_A_uRpohZrb7_0),.din(w_dff_A_gsQw3Cox5_0),.clk(gclk));
	jdff dff_A_MK0VuhU15_1(.dout(w_n904_0[1]),.din(w_dff_A_MK0VuhU15_1),.clk(gclk));
	jdff dff_B_q0XPWQFi0_1(.din(n808),.dout(w_dff_B_q0XPWQFi0_1),.clk(gclk));
	jdff dff_A_WuTLqNa22_0(.dout(w_n706_0[0]),.din(w_dff_A_WuTLqNa22_0),.clk(gclk));
	jdff dff_A_KfoPNO1Y4_0(.dout(w_dff_A_WuTLqNa22_0),.din(w_dff_A_KfoPNO1Y4_0),.clk(gclk));
	jdff dff_A_XSSvmQtG1_0(.dout(w_dff_A_KfoPNO1Y4_0),.din(w_dff_A_XSSvmQtG1_0),.clk(gclk));
	jdff dff_A_ZlsGnQqO7_0(.dout(w_dff_A_XSSvmQtG1_0),.din(w_dff_A_ZlsGnQqO7_0),.clk(gclk));
	jdff dff_A_Aa1DoKfs2_0(.dout(w_dff_A_ZlsGnQqO7_0),.din(w_dff_A_Aa1DoKfs2_0),.clk(gclk));
	jdff dff_A_mqjpVsZq5_0(.dout(w_dff_A_Aa1DoKfs2_0),.din(w_dff_A_mqjpVsZq5_0),.clk(gclk));
	jdff dff_A_5MJeBqd60_0(.dout(w_dff_A_mqjpVsZq5_0),.din(w_dff_A_5MJeBqd60_0),.clk(gclk));
	jdff dff_A_6pmYOGOO3_0(.dout(w_dff_A_5MJeBqd60_0),.din(w_dff_A_6pmYOGOO3_0),.clk(gclk));
	jdff dff_A_ZHU9wbMW3_0(.dout(w_dff_A_6pmYOGOO3_0),.din(w_dff_A_ZHU9wbMW3_0),.clk(gclk));
	jdff dff_A_Z6vGYTU80_0(.dout(w_dff_A_ZHU9wbMW3_0),.din(w_dff_A_Z6vGYTU80_0),.clk(gclk));
	jdff dff_A_sOObR9hA0_0(.dout(w_dff_A_Z6vGYTU80_0),.din(w_dff_A_sOObR9hA0_0),.clk(gclk));
	jdff dff_A_0ejioA165_0(.dout(w_dff_A_sOObR9hA0_0),.din(w_dff_A_0ejioA165_0),.clk(gclk));
	jdff dff_A_LffEP1fF1_0(.dout(w_dff_A_0ejioA165_0),.din(w_dff_A_LffEP1fF1_0),.clk(gclk));
	jdff dff_A_Qjav21df6_0(.dout(w_dff_A_LffEP1fF1_0),.din(w_dff_A_Qjav21df6_0),.clk(gclk));
	jdff dff_A_xQbIpreV1_0(.dout(w_dff_A_Qjav21df6_0),.din(w_dff_A_xQbIpreV1_0),.clk(gclk));
	jdff dff_A_C64Ma2ar9_0(.dout(w_dff_A_xQbIpreV1_0),.din(w_dff_A_C64Ma2ar9_0),.clk(gclk));
	jdff dff_A_fOUgoNZH3_0(.dout(w_dff_A_C64Ma2ar9_0),.din(w_dff_A_fOUgoNZH3_0),.clk(gclk));
	jdff dff_A_fskyirpJ7_0(.dout(w_dff_A_fOUgoNZH3_0),.din(w_dff_A_fskyirpJ7_0),.clk(gclk));
	jdff dff_A_N75iOreL9_0(.dout(w_dff_A_fskyirpJ7_0),.din(w_dff_A_N75iOreL9_0),.clk(gclk));
	jdff dff_A_UfKbiXcp2_0(.dout(w_dff_A_N75iOreL9_0),.din(w_dff_A_UfKbiXcp2_0),.clk(gclk));
	jdff dff_A_NAZcYdOt2_0(.dout(w_dff_A_UfKbiXcp2_0),.din(w_dff_A_NAZcYdOt2_0),.clk(gclk));
	jdff dff_A_fzlEcLXi8_0(.dout(w_dff_A_NAZcYdOt2_0),.din(w_dff_A_fzlEcLXi8_0),.clk(gclk));
	jdff dff_A_xZHh3vOq4_0(.dout(w_dff_A_fzlEcLXi8_0),.din(w_dff_A_xZHh3vOq4_0),.clk(gclk));
	jdff dff_A_diknPS3S5_0(.dout(w_dff_A_xZHh3vOq4_0),.din(w_dff_A_diknPS3S5_0),.clk(gclk));
	jdff dff_A_jVfL5Aub8_0(.dout(w_dff_A_diknPS3S5_0),.din(w_dff_A_jVfL5Aub8_0),.clk(gclk));
	jdff dff_A_JLn3havl0_0(.dout(w_dff_A_jVfL5Aub8_0),.din(w_dff_A_JLn3havl0_0),.clk(gclk));
	jdff dff_A_ewHWcpLv0_0(.dout(w_dff_A_JLn3havl0_0),.din(w_dff_A_ewHWcpLv0_0),.clk(gclk));
	jdff dff_A_pAaIwZXZ5_0(.dout(w_dff_A_ewHWcpLv0_0),.din(w_dff_A_pAaIwZXZ5_0),.clk(gclk));
	jdff dff_A_xqcYvUh81_0(.dout(w_dff_A_pAaIwZXZ5_0),.din(w_dff_A_xqcYvUh81_0),.clk(gclk));
	jdff dff_A_hKojmLny7_0(.dout(w_dff_A_xqcYvUh81_0),.din(w_dff_A_hKojmLny7_0),.clk(gclk));
	jdff dff_A_gcK08Eqn0_0(.dout(w_dff_A_hKojmLny7_0),.din(w_dff_A_gcK08Eqn0_0),.clk(gclk));
	jdff dff_A_MbsevW2o7_0(.dout(w_dff_A_gcK08Eqn0_0),.din(w_dff_A_MbsevW2o7_0),.clk(gclk));
	jdff dff_A_SOwVyMfj0_0(.dout(w_dff_A_MbsevW2o7_0),.din(w_dff_A_SOwVyMfj0_0),.clk(gclk));
	jdff dff_A_sPhTPns42_0(.dout(w_dff_A_SOwVyMfj0_0),.din(w_dff_A_sPhTPns42_0),.clk(gclk));
	jdff dff_A_dW4RF2Ft7_0(.dout(w_dff_A_sPhTPns42_0),.din(w_dff_A_dW4RF2Ft7_0),.clk(gclk));
	jdff dff_A_ARoe1L8O8_0(.dout(w_dff_A_dW4RF2Ft7_0),.din(w_dff_A_ARoe1L8O8_0),.clk(gclk));
	jdff dff_A_kXhHpDur1_0(.dout(w_dff_A_ARoe1L8O8_0),.din(w_dff_A_kXhHpDur1_0),.clk(gclk));
	jdff dff_A_YxS1Ph414_0(.dout(w_dff_A_kXhHpDur1_0),.din(w_dff_A_YxS1Ph414_0),.clk(gclk));
	jdff dff_A_hm4ZlzOA6_0(.dout(w_dff_A_YxS1Ph414_0),.din(w_dff_A_hm4ZlzOA6_0),.clk(gclk));
	jdff dff_A_JDpPRqDB1_0(.dout(w_dff_A_hm4ZlzOA6_0),.din(w_dff_A_JDpPRqDB1_0),.clk(gclk));
	jdff dff_A_7y1XPP7Z4_1(.dout(w_n802_0[1]),.din(w_dff_A_7y1XPP7Z4_1),.clk(gclk));
	jdff dff_B_g43RiTyq0_1(.din(n713),.dout(w_dff_B_g43RiTyq0_1),.clk(gclk));
	jdff dff_B_ZxMqnISu0_1(.din(w_dff_B_g43RiTyq0_1),.dout(w_dff_B_ZxMqnISu0_1),.clk(gclk));
	jdff dff_B_Hc8L1sT89_1(.din(w_dff_B_ZxMqnISu0_1),.dout(w_dff_B_Hc8L1sT89_1),.clk(gclk));
	jdff dff_B_vrKF4epo2_1(.din(w_dff_B_Hc8L1sT89_1),.dout(w_dff_B_vrKF4epo2_1),.clk(gclk));
	jdff dff_B_8Kww9MzI0_1(.din(w_dff_B_vrKF4epo2_1),.dout(w_dff_B_8Kww9MzI0_1),.clk(gclk));
	jdff dff_B_8x8i6mlF1_1(.din(w_dff_B_8Kww9MzI0_1),.dout(w_dff_B_8x8i6mlF1_1),.clk(gclk));
	jdff dff_B_ZjZj9Aby5_1(.din(w_dff_B_8x8i6mlF1_1),.dout(w_dff_B_ZjZj9Aby5_1),.clk(gclk));
	jdff dff_B_D2oBz4Wa0_1(.din(w_dff_B_ZjZj9Aby5_1),.dout(w_dff_B_D2oBz4Wa0_1),.clk(gclk));
	jdff dff_B_hN8VyDGI1_1(.din(w_dff_B_D2oBz4Wa0_1),.dout(w_dff_B_hN8VyDGI1_1),.clk(gclk));
	jdff dff_B_DxRVVLY88_1(.din(w_dff_B_hN8VyDGI1_1),.dout(w_dff_B_DxRVVLY88_1),.clk(gclk));
	jdff dff_B_Kn1YLFL86_1(.din(w_dff_B_DxRVVLY88_1),.dout(w_dff_B_Kn1YLFL86_1),.clk(gclk));
	jdff dff_B_eR9WagRX5_1(.din(w_dff_B_Kn1YLFL86_1),.dout(w_dff_B_eR9WagRX5_1),.clk(gclk));
	jdff dff_B_EfijYsn78_1(.din(w_dff_B_eR9WagRX5_1),.dout(w_dff_B_EfijYsn78_1),.clk(gclk));
	jdff dff_B_ozXFAZpm0_1(.din(w_dff_B_EfijYsn78_1),.dout(w_dff_B_ozXFAZpm0_1),.clk(gclk));
	jdff dff_B_84dE1AQn9_1(.din(w_dff_B_ozXFAZpm0_1),.dout(w_dff_B_84dE1AQn9_1),.clk(gclk));
	jdff dff_B_C7Xn6Wbq5_1(.din(w_dff_B_84dE1AQn9_1),.dout(w_dff_B_C7Xn6Wbq5_1),.clk(gclk));
	jdff dff_B_XF7vc1FB3_1(.din(w_dff_B_C7Xn6Wbq5_1),.dout(w_dff_B_XF7vc1FB3_1),.clk(gclk));
	jdff dff_B_yYPWjdDE5_1(.din(w_dff_B_XF7vc1FB3_1),.dout(w_dff_B_yYPWjdDE5_1),.clk(gclk));
	jdff dff_B_5f7EaXK75_1(.din(w_dff_B_yYPWjdDE5_1),.dout(w_dff_B_5f7EaXK75_1),.clk(gclk));
	jdff dff_B_kjvJJgtf9_1(.din(w_dff_B_5f7EaXK75_1),.dout(w_dff_B_kjvJJgtf9_1),.clk(gclk));
	jdff dff_B_taz7nMrq5_1(.din(w_dff_B_kjvJJgtf9_1),.dout(w_dff_B_taz7nMrq5_1),.clk(gclk));
	jdff dff_B_Gie3gtTv3_1(.din(w_dff_B_taz7nMrq5_1),.dout(w_dff_B_Gie3gtTv3_1),.clk(gclk));
	jdff dff_B_DWUFKs3E6_1(.din(w_dff_B_Gie3gtTv3_1),.dout(w_dff_B_DWUFKs3E6_1),.clk(gclk));
	jdff dff_B_NKoGWVHk5_1(.din(w_dff_B_DWUFKs3E6_1),.dout(w_dff_B_NKoGWVHk5_1),.clk(gclk));
	jdff dff_B_XoeCgNQU5_1(.din(w_dff_B_NKoGWVHk5_1),.dout(w_dff_B_XoeCgNQU5_1),.clk(gclk));
	jdff dff_B_mfcqjjRG6_1(.din(w_dff_B_XoeCgNQU5_1),.dout(w_dff_B_mfcqjjRG6_1),.clk(gclk));
	jdff dff_B_N1oXcL675_1(.din(w_dff_B_mfcqjjRG6_1),.dout(w_dff_B_N1oXcL675_1),.clk(gclk));
	jdff dff_B_P73yMuXu2_1(.din(w_dff_B_N1oXcL675_1),.dout(w_dff_B_P73yMuXu2_1),.clk(gclk));
	jdff dff_B_4Db8brQB2_1(.din(w_dff_B_P73yMuXu2_1),.dout(w_dff_B_4Db8brQB2_1),.clk(gclk));
	jdff dff_B_CjtE1QT35_1(.din(w_dff_B_4Db8brQB2_1),.dout(w_dff_B_CjtE1QT35_1),.clk(gclk));
	jdff dff_B_H7YH7Gy75_1(.din(w_dff_B_CjtE1QT35_1),.dout(w_dff_B_H7YH7Gy75_1),.clk(gclk));
	jdff dff_B_XdewGD5u9_1(.din(w_dff_B_H7YH7Gy75_1),.dout(w_dff_B_XdewGD5u9_1),.clk(gclk));
	jdff dff_B_XEl1n5fU1_1(.din(w_dff_B_XdewGD5u9_1),.dout(w_dff_B_XEl1n5fU1_1),.clk(gclk));
	jdff dff_B_VALSnHhf5_1(.din(w_dff_B_XEl1n5fU1_1),.dout(w_dff_B_VALSnHhf5_1),.clk(gclk));
	jdff dff_B_sdmMjafT8_1(.din(w_dff_B_VALSnHhf5_1),.dout(w_dff_B_sdmMjafT8_1),.clk(gclk));
	jdff dff_B_Z79BEmHT1_1(.din(w_dff_B_sdmMjafT8_1),.dout(w_dff_B_Z79BEmHT1_1),.clk(gclk));
	jdff dff_B_IwWgFsJp8_1(.din(n709),.dout(w_dff_B_IwWgFsJp8_1),.clk(gclk));
	jdff dff_A_Oa1vXFiX9_0(.dout(w_n614_0[0]),.din(w_dff_A_Oa1vXFiX9_0),.clk(gclk));
	jdff dff_A_R3bKBnDr9_0(.dout(w_dff_A_Oa1vXFiX9_0),.din(w_dff_A_R3bKBnDr9_0),.clk(gclk));
	jdff dff_A_ZlLm64wL1_0(.dout(w_dff_A_R3bKBnDr9_0),.din(w_dff_A_ZlLm64wL1_0),.clk(gclk));
	jdff dff_A_e4Gtb3Os3_0(.dout(w_dff_A_ZlLm64wL1_0),.din(w_dff_A_e4Gtb3Os3_0),.clk(gclk));
	jdff dff_A_FN9YtOfB1_0(.dout(w_dff_A_e4Gtb3Os3_0),.din(w_dff_A_FN9YtOfB1_0),.clk(gclk));
	jdff dff_A_rOPYlOn38_0(.dout(w_dff_A_FN9YtOfB1_0),.din(w_dff_A_rOPYlOn38_0),.clk(gclk));
	jdff dff_A_1WFxNLzI3_0(.dout(w_dff_A_rOPYlOn38_0),.din(w_dff_A_1WFxNLzI3_0),.clk(gclk));
	jdff dff_A_2FslWfwU4_0(.dout(w_dff_A_1WFxNLzI3_0),.din(w_dff_A_2FslWfwU4_0),.clk(gclk));
	jdff dff_A_EtzSNt0L2_0(.dout(w_dff_A_2FslWfwU4_0),.din(w_dff_A_EtzSNt0L2_0),.clk(gclk));
	jdff dff_A_iMLREl8e8_0(.dout(w_dff_A_EtzSNt0L2_0),.din(w_dff_A_iMLREl8e8_0),.clk(gclk));
	jdff dff_A_rxPOp8wx7_0(.dout(w_dff_A_iMLREl8e8_0),.din(w_dff_A_rxPOp8wx7_0),.clk(gclk));
	jdff dff_A_g43Bb1ol8_0(.dout(w_dff_A_rxPOp8wx7_0),.din(w_dff_A_g43Bb1ol8_0),.clk(gclk));
	jdff dff_A_ye5rD1Ej7_0(.dout(w_dff_A_g43Bb1ol8_0),.din(w_dff_A_ye5rD1Ej7_0),.clk(gclk));
	jdff dff_A_HxmDsr3t0_0(.dout(w_dff_A_ye5rD1Ej7_0),.din(w_dff_A_HxmDsr3t0_0),.clk(gclk));
	jdff dff_A_RbQ6QcXS9_0(.dout(w_dff_A_HxmDsr3t0_0),.din(w_dff_A_RbQ6QcXS9_0),.clk(gclk));
	jdff dff_A_xFf4yazO4_0(.dout(w_dff_A_RbQ6QcXS9_0),.din(w_dff_A_xFf4yazO4_0),.clk(gclk));
	jdff dff_A_Eeg6ZSa59_0(.dout(w_dff_A_xFf4yazO4_0),.din(w_dff_A_Eeg6ZSa59_0),.clk(gclk));
	jdff dff_A_R0Y8OcgE7_0(.dout(w_dff_A_Eeg6ZSa59_0),.din(w_dff_A_R0Y8OcgE7_0),.clk(gclk));
	jdff dff_A_iSz0WDy75_0(.dout(w_dff_A_R0Y8OcgE7_0),.din(w_dff_A_iSz0WDy75_0),.clk(gclk));
	jdff dff_A_QClbv4NU9_0(.dout(w_dff_A_iSz0WDy75_0),.din(w_dff_A_QClbv4NU9_0),.clk(gclk));
	jdff dff_A_tjoCZtvS8_0(.dout(w_dff_A_QClbv4NU9_0),.din(w_dff_A_tjoCZtvS8_0),.clk(gclk));
	jdff dff_A_4VcbBO8I7_0(.dout(w_dff_A_tjoCZtvS8_0),.din(w_dff_A_4VcbBO8I7_0),.clk(gclk));
	jdff dff_A_6GwuDmAY2_0(.dout(w_dff_A_4VcbBO8I7_0),.din(w_dff_A_6GwuDmAY2_0),.clk(gclk));
	jdff dff_A_m0epqztM4_0(.dout(w_dff_A_6GwuDmAY2_0),.din(w_dff_A_m0epqztM4_0),.clk(gclk));
	jdff dff_A_WWpoYzIe3_0(.dout(w_dff_A_m0epqztM4_0),.din(w_dff_A_WWpoYzIe3_0),.clk(gclk));
	jdff dff_A_UCCVHBbM7_0(.dout(w_dff_A_WWpoYzIe3_0),.din(w_dff_A_UCCVHBbM7_0),.clk(gclk));
	jdff dff_A_Wfq2MU012_0(.dout(w_dff_A_UCCVHBbM7_0),.din(w_dff_A_Wfq2MU012_0),.clk(gclk));
	jdff dff_A_rbpxN1Rn4_0(.dout(w_dff_A_Wfq2MU012_0),.din(w_dff_A_rbpxN1Rn4_0),.clk(gclk));
	jdff dff_A_btalWeFR7_0(.dout(w_dff_A_rbpxN1Rn4_0),.din(w_dff_A_btalWeFR7_0),.clk(gclk));
	jdff dff_A_Ii5XlZRL2_0(.dout(w_dff_A_btalWeFR7_0),.din(w_dff_A_Ii5XlZRL2_0),.clk(gclk));
	jdff dff_A_Fes7awqC7_0(.dout(w_dff_A_Ii5XlZRL2_0),.din(w_dff_A_Fes7awqC7_0),.clk(gclk));
	jdff dff_A_fMZKtSET8_0(.dout(w_dff_A_Fes7awqC7_0),.din(w_dff_A_fMZKtSET8_0),.clk(gclk));
	jdff dff_A_0JnkHxpi7_0(.dout(w_dff_A_fMZKtSET8_0),.din(w_dff_A_0JnkHxpi7_0),.clk(gclk));
	jdff dff_A_2hTJTysR2_0(.dout(w_dff_A_0JnkHxpi7_0),.din(w_dff_A_2hTJTysR2_0),.clk(gclk));
	jdff dff_A_y00YJ24C4_0(.dout(w_dff_A_2hTJTysR2_0),.din(w_dff_A_y00YJ24C4_0),.clk(gclk));
	jdff dff_A_AXw7sj3V1_0(.dout(w_dff_A_y00YJ24C4_0),.din(w_dff_A_AXw7sj3V1_0),.clk(gclk));
	jdff dff_A_kXtpBZXi8_0(.dout(w_dff_A_AXw7sj3V1_0),.din(w_dff_A_kXtpBZXi8_0),.clk(gclk));
	jdff dff_A_CSAuEfHm7_1(.dout(w_n703_0[1]),.din(w_dff_A_CSAuEfHm7_1),.clk(gclk));
	jdff dff_B_cR2gTOZ97_1(.din(n621),.dout(w_dff_B_cR2gTOZ97_1),.clk(gclk));
	jdff dff_B_54i5Q0MS7_1(.din(w_dff_B_cR2gTOZ97_1),.dout(w_dff_B_54i5Q0MS7_1),.clk(gclk));
	jdff dff_B_wtrumuQx4_1(.din(w_dff_B_54i5Q0MS7_1),.dout(w_dff_B_wtrumuQx4_1),.clk(gclk));
	jdff dff_B_6tv5O8MX8_1(.din(w_dff_B_wtrumuQx4_1),.dout(w_dff_B_6tv5O8MX8_1),.clk(gclk));
	jdff dff_B_85mHSmjY2_1(.din(w_dff_B_6tv5O8MX8_1),.dout(w_dff_B_85mHSmjY2_1),.clk(gclk));
	jdff dff_B_olxTzOCY3_1(.din(w_dff_B_85mHSmjY2_1),.dout(w_dff_B_olxTzOCY3_1),.clk(gclk));
	jdff dff_B_3CPHOMdp8_1(.din(w_dff_B_olxTzOCY3_1),.dout(w_dff_B_3CPHOMdp8_1),.clk(gclk));
	jdff dff_B_QHFoXO5q9_1(.din(w_dff_B_3CPHOMdp8_1),.dout(w_dff_B_QHFoXO5q9_1),.clk(gclk));
	jdff dff_B_rB099p4a1_1(.din(w_dff_B_QHFoXO5q9_1),.dout(w_dff_B_rB099p4a1_1),.clk(gclk));
	jdff dff_B_3aDHaYDp7_1(.din(w_dff_B_rB099p4a1_1),.dout(w_dff_B_3aDHaYDp7_1),.clk(gclk));
	jdff dff_B_LoZhRq1q7_1(.din(w_dff_B_3aDHaYDp7_1),.dout(w_dff_B_LoZhRq1q7_1),.clk(gclk));
	jdff dff_B_yWnOi33b5_1(.din(w_dff_B_LoZhRq1q7_1),.dout(w_dff_B_yWnOi33b5_1),.clk(gclk));
	jdff dff_B_aahxRXEg0_1(.din(w_dff_B_yWnOi33b5_1),.dout(w_dff_B_aahxRXEg0_1),.clk(gclk));
	jdff dff_B_fz2WoD0H2_1(.din(w_dff_B_aahxRXEg0_1),.dout(w_dff_B_fz2WoD0H2_1),.clk(gclk));
	jdff dff_B_QCOziseq7_1(.din(w_dff_B_fz2WoD0H2_1),.dout(w_dff_B_QCOziseq7_1),.clk(gclk));
	jdff dff_B_90Tn0qPk1_1(.din(w_dff_B_QCOziseq7_1),.dout(w_dff_B_90Tn0qPk1_1),.clk(gclk));
	jdff dff_B_2jyAQP1L0_1(.din(w_dff_B_90Tn0qPk1_1),.dout(w_dff_B_2jyAQP1L0_1),.clk(gclk));
	jdff dff_B_JEloTsq18_1(.din(w_dff_B_2jyAQP1L0_1),.dout(w_dff_B_JEloTsq18_1),.clk(gclk));
	jdff dff_B_00823XVm1_1(.din(w_dff_B_JEloTsq18_1),.dout(w_dff_B_00823XVm1_1),.clk(gclk));
	jdff dff_B_aBqK1NJg7_1(.din(w_dff_B_00823XVm1_1),.dout(w_dff_B_aBqK1NJg7_1),.clk(gclk));
	jdff dff_B_V66xwiMO0_1(.din(w_dff_B_aBqK1NJg7_1),.dout(w_dff_B_V66xwiMO0_1),.clk(gclk));
	jdff dff_B_PvkSu1sO1_1(.din(w_dff_B_V66xwiMO0_1),.dout(w_dff_B_PvkSu1sO1_1),.clk(gclk));
	jdff dff_B_bNzryRVm1_1(.din(w_dff_B_PvkSu1sO1_1),.dout(w_dff_B_bNzryRVm1_1),.clk(gclk));
	jdff dff_B_Q3flWllZ2_1(.din(w_dff_B_bNzryRVm1_1),.dout(w_dff_B_Q3flWllZ2_1),.clk(gclk));
	jdff dff_B_ndvr2KGu4_1(.din(w_dff_B_Q3flWllZ2_1),.dout(w_dff_B_ndvr2KGu4_1),.clk(gclk));
	jdff dff_B_IiO0KRMc8_1(.din(w_dff_B_ndvr2KGu4_1),.dout(w_dff_B_IiO0KRMc8_1),.clk(gclk));
	jdff dff_B_ABYYUiQK7_1(.din(w_dff_B_IiO0KRMc8_1),.dout(w_dff_B_ABYYUiQK7_1),.clk(gclk));
	jdff dff_B_TZpxFUax0_1(.din(w_dff_B_ABYYUiQK7_1),.dout(w_dff_B_TZpxFUax0_1),.clk(gclk));
	jdff dff_B_W5ZNOVpY5_1(.din(w_dff_B_TZpxFUax0_1),.dout(w_dff_B_W5ZNOVpY5_1),.clk(gclk));
	jdff dff_B_WOYym9X45_1(.din(w_dff_B_W5ZNOVpY5_1),.dout(w_dff_B_WOYym9X45_1),.clk(gclk));
	jdff dff_B_bNIxA3FX7_1(.din(w_dff_B_WOYym9X45_1),.dout(w_dff_B_bNIxA3FX7_1),.clk(gclk));
	jdff dff_B_4NHOyic36_1(.din(w_dff_B_bNIxA3FX7_1),.dout(w_dff_B_4NHOyic36_1),.clk(gclk));
	jdff dff_B_XbI8uxyG4_1(.din(w_dff_B_4NHOyic36_1),.dout(w_dff_B_XbI8uxyG4_1),.clk(gclk));
	jdff dff_B_MJFHgnav4_1(.din(n617),.dout(w_dff_B_MJFHgnav4_1),.clk(gclk));
	jdff dff_A_p9jKWYMW0_0(.dout(w_n529_0[0]),.din(w_dff_A_p9jKWYMW0_0),.clk(gclk));
	jdff dff_A_jsd4sH1j8_0(.dout(w_dff_A_p9jKWYMW0_0),.din(w_dff_A_jsd4sH1j8_0),.clk(gclk));
	jdff dff_A_P6ZXIqrC9_0(.dout(w_dff_A_jsd4sH1j8_0),.din(w_dff_A_P6ZXIqrC9_0),.clk(gclk));
	jdff dff_A_xrVvMFLv8_0(.dout(w_dff_A_P6ZXIqrC9_0),.din(w_dff_A_xrVvMFLv8_0),.clk(gclk));
	jdff dff_A_NYDw1c584_0(.dout(w_dff_A_xrVvMFLv8_0),.din(w_dff_A_NYDw1c584_0),.clk(gclk));
	jdff dff_A_dYmh04vC5_0(.dout(w_dff_A_NYDw1c584_0),.din(w_dff_A_dYmh04vC5_0),.clk(gclk));
	jdff dff_A_02DZLLnu9_0(.dout(w_dff_A_dYmh04vC5_0),.din(w_dff_A_02DZLLnu9_0),.clk(gclk));
	jdff dff_A_SNNw2z1M2_0(.dout(w_dff_A_02DZLLnu9_0),.din(w_dff_A_SNNw2z1M2_0),.clk(gclk));
	jdff dff_A_dKJK6svR5_0(.dout(w_dff_A_SNNw2z1M2_0),.din(w_dff_A_dKJK6svR5_0),.clk(gclk));
	jdff dff_A_fOjQaHos0_0(.dout(w_dff_A_dKJK6svR5_0),.din(w_dff_A_fOjQaHos0_0),.clk(gclk));
	jdff dff_A_uvCSk85k2_0(.dout(w_dff_A_fOjQaHos0_0),.din(w_dff_A_uvCSk85k2_0),.clk(gclk));
	jdff dff_A_jKvttLj64_0(.dout(w_dff_A_uvCSk85k2_0),.din(w_dff_A_jKvttLj64_0),.clk(gclk));
	jdff dff_A_hb2IhXrr6_0(.dout(w_dff_A_jKvttLj64_0),.din(w_dff_A_hb2IhXrr6_0),.clk(gclk));
	jdff dff_A_PM6uz7Rv9_0(.dout(w_dff_A_hb2IhXrr6_0),.din(w_dff_A_PM6uz7Rv9_0),.clk(gclk));
	jdff dff_A_bJp0c96x2_0(.dout(w_dff_A_PM6uz7Rv9_0),.din(w_dff_A_bJp0c96x2_0),.clk(gclk));
	jdff dff_A_FuGseIGv1_0(.dout(w_dff_A_bJp0c96x2_0),.din(w_dff_A_FuGseIGv1_0),.clk(gclk));
	jdff dff_A_3QTqhoPC7_0(.dout(w_dff_A_FuGseIGv1_0),.din(w_dff_A_3QTqhoPC7_0),.clk(gclk));
	jdff dff_A_jG9FYM2V2_0(.dout(w_dff_A_3QTqhoPC7_0),.din(w_dff_A_jG9FYM2V2_0),.clk(gclk));
	jdff dff_A_3n4B5e6L4_0(.dout(w_dff_A_jG9FYM2V2_0),.din(w_dff_A_3n4B5e6L4_0),.clk(gclk));
	jdff dff_A_6frpnqbJ6_0(.dout(w_dff_A_3n4B5e6L4_0),.din(w_dff_A_6frpnqbJ6_0),.clk(gclk));
	jdff dff_A_WZh8TLRI9_0(.dout(w_dff_A_6frpnqbJ6_0),.din(w_dff_A_WZh8TLRI9_0),.clk(gclk));
	jdff dff_A_iJKnNzY76_0(.dout(w_dff_A_WZh8TLRI9_0),.din(w_dff_A_iJKnNzY76_0),.clk(gclk));
	jdff dff_A_CQiqHLOa7_0(.dout(w_dff_A_iJKnNzY76_0),.din(w_dff_A_CQiqHLOa7_0),.clk(gclk));
	jdff dff_A_56n11hGU8_0(.dout(w_dff_A_CQiqHLOa7_0),.din(w_dff_A_56n11hGU8_0),.clk(gclk));
	jdff dff_A_zRGzsltV2_0(.dout(w_dff_A_56n11hGU8_0),.din(w_dff_A_zRGzsltV2_0),.clk(gclk));
	jdff dff_A_fdUGG1xu6_0(.dout(w_dff_A_zRGzsltV2_0),.din(w_dff_A_fdUGG1xu6_0),.clk(gclk));
	jdff dff_A_ZB7d8JM58_0(.dout(w_dff_A_fdUGG1xu6_0),.din(w_dff_A_ZB7d8JM58_0),.clk(gclk));
	jdff dff_A_VoCT5toY1_0(.dout(w_dff_A_ZB7d8JM58_0),.din(w_dff_A_VoCT5toY1_0),.clk(gclk));
	jdff dff_A_DEaZWes05_0(.dout(w_dff_A_VoCT5toY1_0),.din(w_dff_A_DEaZWes05_0),.clk(gclk));
	jdff dff_A_d7h3sCZh3_0(.dout(w_dff_A_DEaZWes05_0),.din(w_dff_A_d7h3sCZh3_0),.clk(gclk));
	jdff dff_A_3yDKZYX31_0(.dout(w_dff_A_d7h3sCZh3_0),.din(w_dff_A_3yDKZYX31_0),.clk(gclk));
	jdff dff_A_n0Z7vuAQ5_0(.dout(w_dff_A_3yDKZYX31_0),.din(w_dff_A_n0Z7vuAQ5_0),.clk(gclk));
	jdff dff_A_h5FTBKqR0_0(.dout(w_dff_A_n0Z7vuAQ5_0),.din(w_dff_A_h5FTBKqR0_0),.clk(gclk));
	jdff dff_A_8FMft7rY4_0(.dout(w_dff_A_h5FTBKqR0_0),.din(w_dff_A_8FMft7rY4_0),.clk(gclk));
	jdff dff_A_VCBWiqrM6_1(.dout(w_n611_0[1]),.din(w_dff_A_VCBWiqrM6_1),.clk(gclk));
	jdff dff_B_VXUxXE5i2_1(.din(n536),.dout(w_dff_B_VXUxXE5i2_1),.clk(gclk));
	jdff dff_B_0NqgOcbr6_1(.din(w_dff_B_VXUxXE5i2_1),.dout(w_dff_B_0NqgOcbr6_1),.clk(gclk));
	jdff dff_B_a7UIAezb6_1(.din(w_dff_B_0NqgOcbr6_1),.dout(w_dff_B_a7UIAezb6_1),.clk(gclk));
	jdff dff_B_WoLv6GGD0_1(.din(w_dff_B_a7UIAezb6_1),.dout(w_dff_B_WoLv6GGD0_1),.clk(gclk));
	jdff dff_B_z394AiBi7_1(.din(w_dff_B_WoLv6GGD0_1),.dout(w_dff_B_z394AiBi7_1),.clk(gclk));
	jdff dff_B_vWoIU1SC6_1(.din(w_dff_B_z394AiBi7_1),.dout(w_dff_B_vWoIU1SC6_1),.clk(gclk));
	jdff dff_B_2y5u0C9w4_1(.din(w_dff_B_vWoIU1SC6_1),.dout(w_dff_B_2y5u0C9w4_1),.clk(gclk));
	jdff dff_B_8Wgyh1953_1(.din(w_dff_B_2y5u0C9w4_1),.dout(w_dff_B_8Wgyh1953_1),.clk(gclk));
	jdff dff_B_JXdJOFc00_1(.din(w_dff_B_8Wgyh1953_1),.dout(w_dff_B_JXdJOFc00_1),.clk(gclk));
	jdff dff_B_HA7BnoSR1_1(.din(w_dff_B_JXdJOFc00_1),.dout(w_dff_B_HA7BnoSR1_1),.clk(gclk));
	jdff dff_B_vGm4ksid7_1(.din(w_dff_B_HA7BnoSR1_1),.dout(w_dff_B_vGm4ksid7_1),.clk(gclk));
	jdff dff_B_9CEbEvHy7_1(.din(w_dff_B_vGm4ksid7_1),.dout(w_dff_B_9CEbEvHy7_1),.clk(gclk));
	jdff dff_B_0pCRhHbD2_1(.din(w_dff_B_9CEbEvHy7_1),.dout(w_dff_B_0pCRhHbD2_1),.clk(gclk));
	jdff dff_B_l1S9vmLL9_1(.din(w_dff_B_0pCRhHbD2_1),.dout(w_dff_B_l1S9vmLL9_1),.clk(gclk));
	jdff dff_B_quMxuRZH4_1(.din(w_dff_B_l1S9vmLL9_1),.dout(w_dff_B_quMxuRZH4_1),.clk(gclk));
	jdff dff_B_xpHvWSF86_1(.din(w_dff_B_quMxuRZH4_1),.dout(w_dff_B_xpHvWSF86_1),.clk(gclk));
	jdff dff_B_xHMh5C4h8_1(.din(w_dff_B_xpHvWSF86_1),.dout(w_dff_B_xHMh5C4h8_1),.clk(gclk));
	jdff dff_B_1IOTEWeh1_1(.din(w_dff_B_xHMh5C4h8_1),.dout(w_dff_B_1IOTEWeh1_1),.clk(gclk));
	jdff dff_B_0W4bQnwp0_1(.din(w_dff_B_1IOTEWeh1_1),.dout(w_dff_B_0W4bQnwp0_1),.clk(gclk));
	jdff dff_B_6HD1SHxH2_1(.din(w_dff_B_0W4bQnwp0_1),.dout(w_dff_B_6HD1SHxH2_1),.clk(gclk));
	jdff dff_B_CEoCruuK5_1(.din(w_dff_B_6HD1SHxH2_1),.dout(w_dff_B_CEoCruuK5_1),.clk(gclk));
	jdff dff_B_wH5rwERM2_1(.din(w_dff_B_CEoCruuK5_1),.dout(w_dff_B_wH5rwERM2_1),.clk(gclk));
	jdff dff_B_pGf1PXjf4_1(.din(w_dff_B_wH5rwERM2_1),.dout(w_dff_B_pGf1PXjf4_1),.clk(gclk));
	jdff dff_B_VYyTK3eA4_1(.din(w_dff_B_pGf1PXjf4_1),.dout(w_dff_B_VYyTK3eA4_1),.clk(gclk));
	jdff dff_B_cZTF5xol6_1(.din(w_dff_B_VYyTK3eA4_1),.dout(w_dff_B_cZTF5xol6_1),.clk(gclk));
	jdff dff_B_4pzDosNZ2_1(.din(w_dff_B_cZTF5xol6_1),.dout(w_dff_B_4pzDosNZ2_1),.clk(gclk));
	jdff dff_B_6EVOQlFo0_1(.din(w_dff_B_4pzDosNZ2_1),.dout(w_dff_B_6EVOQlFo0_1),.clk(gclk));
	jdff dff_B_9XwNGk0U2_1(.din(w_dff_B_6EVOQlFo0_1),.dout(w_dff_B_9XwNGk0U2_1),.clk(gclk));
	jdff dff_B_eWEe3ipL1_1(.din(w_dff_B_9XwNGk0U2_1),.dout(w_dff_B_eWEe3ipL1_1),.clk(gclk));
	jdff dff_B_3mtpIpHT8_1(.din(w_dff_B_eWEe3ipL1_1),.dout(w_dff_B_3mtpIpHT8_1),.clk(gclk));
	jdff dff_B_os8dMX4n3_1(.din(n532),.dout(w_dff_B_os8dMX4n3_1),.clk(gclk));
	jdff dff_A_zojWS9US5_0(.dout(w_n451_0[0]),.din(w_dff_A_zojWS9US5_0),.clk(gclk));
	jdff dff_A_YAVei9ND7_0(.dout(w_dff_A_zojWS9US5_0),.din(w_dff_A_YAVei9ND7_0),.clk(gclk));
	jdff dff_A_5FLD68tZ1_0(.dout(w_dff_A_YAVei9ND7_0),.din(w_dff_A_5FLD68tZ1_0),.clk(gclk));
	jdff dff_A_EzTdPr8q3_0(.dout(w_dff_A_5FLD68tZ1_0),.din(w_dff_A_EzTdPr8q3_0),.clk(gclk));
	jdff dff_A_gCIHjZCT1_0(.dout(w_dff_A_EzTdPr8q3_0),.din(w_dff_A_gCIHjZCT1_0),.clk(gclk));
	jdff dff_A_Zbd9pH166_0(.dout(w_dff_A_gCIHjZCT1_0),.din(w_dff_A_Zbd9pH166_0),.clk(gclk));
	jdff dff_A_6GruaOuZ0_0(.dout(w_dff_A_Zbd9pH166_0),.din(w_dff_A_6GruaOuZ0_0),.clk(gclk));
	jdff dff_A_GveBnI4F0_0(.dout(w_dff_A_6GruaOuZ0_0),.din(w_dff_A_GveBnI4F0_0),.clk(gclk));
	jdff dff_A_nJUsncYO4_0(.dout(w_dff_A_GveBnI4F0_0),.din(w_dff_A_nJUsncYO4_0),.clk(gclk));
	jdff dff_A_Emad5PsB9_0(.dout(w_dff_A_nJUsncYO4_0),.din(w_dff_A_Emad5PsB9_0),.clk(gclk));
	jdff dff_A_pTE7WaHH6_0(.dout(w_dff_A_Emad5PsB9_0),.din(w_dff_A_pTE7WaHH6_0),.clk(gclk));
	jdff dff_A_8asdnRH69_0(.dout(w_dff_A_pTE7WaHH6_0),.din(w_dff_A_8asdnRH69_0),.clk(gclk));
	jdff dff_A_GVwV9WVe4_0(.dout(w_dff_A_8asdnRH69_0),.din(w_dff_A_GVwV9WVe4_0),.clk(gclk));
	jdff dff_A_KfDO0agX3_0(.dout(w_dff_A_GVwV9WVe4_0),.din(w_dff_A_KfDO0agX3_0),.clk(gclk));
	jdff dff_A_XuhxZ9mO5_0(.dout(w_dff_A_KfDO0agX3_0),.din(w_dff_A_XuhxZ9mO5_0),.clk(gclk));
	jdff dff_A_yK8srXoQ9_0(.dout(w_dff_A_XuhxZ9mO5_0),.din(w_dff_A_yK8srXoQ9_0),.clk(gclk));
	jdff dff_A_WmY2WDt34_0(.dout(w_dff_A_yK8srXoQ9_0),.din(w_dff_A_WmY2WDt34_0),.clk(gclk));
	jdff dff_A_0K8KwNXu9_0(.dout(w_dff_A_WmY2WDt34_0),.din(w_dff_A_0K8KwNXu9_0),.clk(gclk));
	jdff dff_A_nYsKGQUc6_0(.dout(w_dff_A_0K8KwNXu9_0),.din(w_dff_A_nYsKGQUc6_0),.clk(gclk));
	jdff dff_A_9vqx9Qht4_0(.dout(w_dff_A_nYsKGQUc6_0),.din(w_dff_A_9vqx9Qht4_0),.clk(gclk));
	jdff dff_A_LOf30NvJ6_0(.dout(w_dff_A_9vqx9Qht4_0),.din(w_dff_A_LOf30NvJ6_0),.clk(gclk));
	jdff dff_A_prvmZykS0_0(.dout(w_dff_A_LOf30NvJ6_0),.din(w_dff_A_prvmZykS0_0),.clk(gclk));
	jdff dff_A_R5x4RGFX9_0(.dout(w_dff_A_prvmZykS0_0),.din(w_dff_A_R5x4RGFX9_0),.clk(gclk));
	jdff dff_A_qgGvadVp9_0(.dout(w_dff_A_R5x4RGFX9_0),.din(w_dff_A_qgGvadVp9_0),.clk(gclk));
	jdff dff_A_lqobwI2Z9_0(.dout(w_dff_A_qgGvadVp9_0),.din(w_dff_A_lqobwI2Z9_0),.clk(gclk));
	jdff dff_A_LlAoWolS7_0(.dout(w_dff_A_lqobwI2Z9_0),.din(w_dff_A_LlAoWolS7_0),.clk(gclk));
	jdff dff_A_OQDWOHiI4_0(.dout(w_dff_A_LlAoWolS7_0),.din(w_dff_A_OQDWOHiI4_0),.clk(gclk));
	jdff dff_A_pFZ61ev29_0(.dout(w_dff_A_OQDWOHiI4_0),.din(w_dff_A_pFZ61ev29_0),.clk(gclk));
	jdff dff_A_S0iNfoEu0_0(.dout(w_dff_A_pFZ61ev29_0),.din(w_dff_A_S0iNfoEu0_0),.clk(gclk));
	jdff dff_A_TzYCBMEP7_0(.dout(w_dff_A_S0iNfoEu0_0),.din(w_dff_A_TzYCBMEP7_0),.clk(gclk));
	jdff dff_A_KESIRdKO2_0(.dout(w_dff_A_TzYCBMEP7_0),.din(w_dff_A_KESIRdKO2_0),.clk(gclk));
	jdff dff_A_lHvD8GlN0_1(.dout(w_n526_0[1]),.din(w_dff_A_lHvD8GlN0_1),.clk(gclk));
	jdff dff_B_aSADHQTu3_1(.din(n458),.dout(w_dff_B_aSADHQTu3_1),.clk(gclk));
	jdff dff_B_3ZdcsKJH9_1(.din(w_dff_B_aSADHQTu3_1),.dout(w_dff_B_3ZdcsKJH9_1),.clk(gclk));
	jdff dff_B_ZqWefski7_1(.din(w_dff_B_3ZdcsKJH9_1),.dout(w_dff_B_ZqWefski7_1),.clk(gclk));
	jdff dff_B_hizDrtCA7_1(.din(w_dff_B_ZqWefski7_1),.dout(w_dff_B_hizDrtCA7_1),.clk(gclk));
	jdff dff_B_ptBNrwE36_1(.din(w_dff_B_hizDrtCA7_1),.dout(w_dff_B_ptBNrwE36_1),.clk(gclk));
	jdff dff_B_VwBMDQx89_1(.din(w_dff_B_ptBNrwE36_1),.dout(w_dff_B_VwBMDQx89_1),.clk(gclk));
	jdff dff_B_8tDafc114_1(.din(w_dff_B_VwBMDQx89_1),.dout(w_dff_B_8tDafc114_1),.clk(gclk));
	jdff dff_B_twfHxHMw7_1(.din(w_dff_B_8tDafc114_1),.dout(w_dff_B_twfHxHMw7_1),.clk(gclk));
	jdff dff_B_a575eMHI3_1(.din(w_dff_B_twfHxHMw7_1),.dout(w_dff_B_a575eMHI3_1),.clk(gclk));
	jdff dff_B_swQw10Ym0_1(.din(w_dff_B_a575eMHI3_1),.dout(w_dff_B_swQw10Ym0_1),.clk(gclk));
	jdff dff_B_2XznyWvl3_1(.din(w_dff_B_swQw10Ym0_1),.dout(w_dff_B_2XznyWvl3_1),.clk(gclk));
	jdff dff_B_x7kgNVEF7_1(.din(w_dff_B_2XznyWvl3_1),.dout(w_dff_B_x7kgNVEF7_1),.clk(gclk));
	jdff dff_B_ZCco6TX03_1(.din(w_dff_B_x7kgNVEF7_1),.dout(w_dff_B_ZCco6TX03_1),.clk(gclk));
	jdff dff_B_Vd35OrAI7_1(.din(w_dff_B_ZCco6TX03_1),.dout(w_dff_B_Vd35OrAI7_1),.clk(gclk));
	jdff dff_B_twy1WSuR0_1(.din(w_dff_B_Vd35OrAI7_1),.dout(w_dff_B_twy1WSuR0_1),.clk(gclk));
	jdff dff_B_fFBtw0bh2_1(.din(w_dff_B_twy1WSuR0_1),.dout(w_dff_B_fFBtw0bh2_1),.clk(gclk));
	jdff dff_B_KfambDLf9_1(.din(w_dff_B_fFBtw0bh2_1),.dout(w_dff_B_KfambDLf9_1),.clk(gclk));
	jdff dff_B_uT46plvO4_1(.din(w_dff_B_KfambDLf9_1),.dout(w_dff_B_uT46plvO4_1),.clk(gclk));
	jdff dff_B_IUZBAAxX6_1(.din(w_dff_B_uT46plvO4_1),.dout(w_dff_B_IUZBAAxX6_1),.clk(gclk));
	jdff dff_B_8giSlLJ91_1(.din(w_dff_B_IUZBAAxX6_1),.dout(w_dff_B_8giSlLJ91_1),.clk(gclk));
	jdff dff_B_EQX30hvF5_1(.din(w_dff_B_8giSlLJ91_1),.dout(w_dff_B_EQX30hvF5_1),.clk(gclk));
	jdff dff_B_sBLF6frq1_1(.din(w_dff_B_EQX30hvF5_1),.dout(w_dff_B_sBLF6frq1_1),.clk(gclk));
	jdff dff_B_bqc2mA7v5_1(.din(w_dff_B_sBLF6frq1_1),.dout(w_dff_B_bqc2mA7v5_1),.clk(gclk));
	jdff dff_B_qIBiK0BQ4_1(.din(w_dff_B_bqc2mA7v5_1),.dout(w_dff_B_qIBiK0BQ4_1),.clk(gclk));
	jdff dff_B_BYMeohTD0_1(.din(w_dff_B_qIBiK0BQ4_1),.dout(w_dff_B_BYMeohTD0_1),.clk(gclk));
	jdff dff_B_NAwfn8bf0_1(.din(w_dff_B_BYMeohTD0_1),.dout(w_dff_B_NAwfn8bf0_1),.clk(gclk));
	jdff dff_B_SB9jIKZE4_1(.din(w_dff_B_NAwfn8bf0_1),.dout(w_dff_B_SB9jIKZE4_1),.clk(gclk));
	jdff dff_B_V2FILeAh0_1(.din(n454),.dout(w_dff_B_V2FILeAh0_1),.clk(gclk));
	jdff dff_A_VuO3Iqgm2_0(.dout(w_n380_0[0]),.din(w_dff_A_VuO3Iqgm2_0),.clk(gclk));
	jdff dff_A_AtrwzAHS5_0(.dout(w_dff_A_VuO3Iqgm2_0),.din(w_dff_A_AtrwzAHS5_0),.clk(gclk));
	jdff dff_A_fouVqPd42_0(.dout(w_dff_A_AtrwzAHS5_0),.din(w_dff_A_fouVqPd42_0),.clk(gclk));
	jdff dff_A_NAIU3vfv8_0(.dout(w_dff_A_fouVqPd42_0),.din(w_dff_A_NAIU3vfv8_0),.clk(gclk));
	jdff dff_A_vRutJaBF8_0(.dout(w_dff_A_NAIU3vfv8_0),.din(w_dff_A_vRutJaBF8_0),.clk(gclk));
	jdff dff_A_yZEnEJJ37_0(.dout(w_dff_A_vRutJaBF8_0),.din(w_dff_A_yZEnEJJ37_0),.clk(gclk));
	jdff dff_A_nVAERRRU4_0(.dout(w_dff_A_yZEnEJJ37_0),.din(w_dff_A_nVAERRRU4_0),.clk(gclk));
	jdff dff_A_MiKfNUtT0_0(.dout(w_dff_A_nVAERRRU4_0),.din(w_dff_A_MiKfNUtT0_0),.clk(gclk));
	jdff dff_A_lri4jbPY3_0(.dout(w_dff_A_MiKfNUtT0_0),.din(w_dff_A_lri4jbPY3_0),.clk(gclk));
	jdff dff_A_om0DWTBR4_0(.dout(w_dff_A_lri4jbPY3_0),.din(w_dff_A_om0DWTBR4_0),.clk(gclk));
	jdff dff_A_Cb03oVk69_0(.dout(w_dff_A_om0DWTBR4_0),.din(w_dff_A_Cb03oVk69_0),.clk(gclk));
	jdff dff_A_TJTBq4iX4_0(.dout(w_dff_A_Cb03oVk69_0),.din(w_dff_A_TJTBq4iX4_0),.clk(gclk));
	jdff dff_A_Dhw3wSJZ4_0(.dout(w_dff_A_TJTBq4iX4_0),.din(w_dff_A_Dhw3wSJZ4_0),.clk(gclk));
	jdff dff_A_4fat33Bv6_0(.dout(w_dff_A_Dhw3wSJZ4_0),.din(w_dff_A_4fat33Bv6_0),.clk(gclk));
	jdff dff_A_muSacNYn5_0(.dout(w_dff_A_4fat33Bv6_0),.din(w_dff_A_muSacNYn5_0),.clk(gclk));
	jdff dff_A_R7n0p3s09_0(.dout(w_dff_A_muSacNYn5_0),.din(w_dff_A_R7n0p3s09_0),.clk(gclk));
	jdff dff_A_IaSfGTGT3_0(.dout(w_dff_A_R7n0p3s09_0),.din(w_dff_A_IaSfGTGT3_0),.clk(gclk));
	jdff dff_A_RhBN7Wl41_0(.dout(w_dff_A_IaSfGTGT3_0),.din(w_dff_A_RhBN7Wl41_0),.clk(gclk));
	jdff dff_A_QgX6Xu133_0(.dout(w_dff_A_RhBN7Wl41_0),.din(w_dff_A_QgX6Xu133_0),.clk(gclk));
	jdff dff_A_xGh3H45m1_0(.dout(w_dff_A_QgX6Xu133_0),.din(w_dff_A_xGh3H45m1_0),.clk(gclk));
	jdff dff_A_tcfaNK5u1_0(.dout(w_dff_A_xGh3H45m1_0),.din(w_dff_A_tcfaNK5u1_0),.clk(gclk));
	jdff dff_A_DGJ9JMi79_0(.dout(w_dff_A_tcfaNK5u1_0),.din(w_dff_A_DGJ9JMi79_0),.clk(gclk));
	jdff dff_A_ouQ01lMY7_0(.dout(w_dff_A_DGJ9JMi79_0),.din(w_dff_A_ouQ01lMY7_0),.clk(gclk));
	jdff dff_A_D0KXoUpF1_0(.dout(w_dff_A_ouQ01lMY7_0),.din(w_dff_A_D0KXoUpF1_0),.clk(gclk));
	jdff dff_A_fRLdcCCO6_0(.dout(w_dff_A_D0KXoUpF1_0),.din(w_dff_A_fRLdcCCO6_0),.clk(gclk));
	jdff dff_A_qF7n0lNR0_0(.dout(w_dff_A_fRLdcCCO6_0),.din(w_dff_A_qF7n0lNR0_0),.clk(gclk));
	jdff dff_A_QAZ1OWo78_0(.dout(w_dff_A_qF7n0lNR0_0),.din(w_dff_A_QAZ1OWo78_0),.clk(gclk));
	jdff dff_A_8REIYbrZ2_0(.dout(w_dff_A_QAZ1OWo78_0),.din(w_dff_A_8REIYbrZ2_0),.clk(gclk));
	jdff dff_A_DkEdws1O4_1(.dout(w_n448_0[1]),.din(w_dff_A_DkEdws1O4_1),.clk(gclk));
	jdff dff_B_1Hwnia6y5_1(.din(n387),.dout(w_dff_B_1Hwnia6y5_1),.clk(gclk));
	jdff dff_B_7eRMdeHJ6_1(.din(w_dff_B_1Hwnia6y5_1),.dout(w_dff_B_7eRMdeHJ6_1),.clk(gclk));
	jdff dff_B_XP15YOmj4_1(.din(w_dff_B_7eRMdeHJ6_1),.dout(w_dff_B_XP15YOmj4_1),.clk(gclk));
	jdff dff_B_lw6qK0rJ5_1(.din(w_dff_B_XP15YOmj4_1),.dout(w_dff_B_lw6qK0rJ5_1),.clk(gclk));
	jdff dff_B_zUPspc0Q0_1(.din(w_dff_B_lw6qK0rJ5_1),.dout(w_dff_B_zUPspc0Q0_1),.clk(gclk));
	jdff dff_B_Htv7EuUU9_1(.din(w_dff_B_zUPspc0Q0_1),.dout(w_dff_B_Htv7EuUU9_1),.clk(gclk));
	jdff dff_B_5b2Rgo8m0_1(.din(w_dff_B_Htv7EuUU9_1),.dout(w_dff_B_5b2Rgo8m0_1),.clk(gclk));
	jdff dff_B_OkrF5aAh4_1(.din(w_dff_B_5b2Rgo8m0_1),.dout(w_dff_B_OkrF5aAh4_1),.clk(gclk));
	jdff dff_B_2uVSew0n9_1(.din(w_dff_B_OkrF5aAh4_1),.dout(w_dff_B_2uVSew0n9_1),.clk(gclk));
	jdff dff_B_mJIZdswJ0_1(.din(w_dff_B_2uVSew0n9_1),.dout(w_dff_B_mJIZdswJ0_1),.clk(gclk));
	jdff dff_B_2rXngZl52_1(.din(w_dff_B_mJIZdswJ0_1),.dout(w_dff_B_2rXngZl52_1),.clk(gclk));
	jdff dff_B_3MwG9N8o0_1(.din(w_dff_B_2rXngZl52_1),.dout(w_dff_B_3MwG9N8o0_1),.clk(gclk));
	jdff dff_B_iHT480Tn6_1(.din(w_dff_B_3MwG9N8o0_1),.dout(w_dff_B_iHT480Tn6_1),.clk(gclk));
	jdff dff_B_yEywQHVs1_1(.din(w_dff_B_iHT480Tn6_1),.dout(w_dff_B_yEywQHVs1_1),.clk(gclk));
	jdff dff_B_Rzwsub104_1(.din(w_dff_B_yEywQHVs1_1),.dout(w_dff_B_Rzwsub104_1),.clk(gclk));
	jdff dff_B_xRfHIyoQ7_1(.din(w_dff_B_Rzwsub104_1),.dout(w_dff_B_xRfHIyoQ7_1),.clk(gclk));
	jdff dff_B_N5u7Y69e2_1(.din(w_dff_B_xRfHIyoQ7_1),.dout(w_dff_B_N5u7Y69e2_1),.clk(gclk));
	jdff dff_B_o1Wyqwih8_1(.din(w_dff_B_N5u7Y69e2_1),.dout(w_dff_B_o1Wyqwih8_1),.clk(gclk));
	jdff dff_B_0PoCoKpS5_1(.din(w_dff_B_o1Wyqwih8_1),.dout(w_dff_B_0PoCoKpS5_1),.clk(gclk));
	jdff dff_B_abBCvjBt5_1(.din(w_dff_B_0PoCoKpS5_1),.dout(w_dff_B_abBCvjBt5_1),.clk(gclk));
	jdff dff_B_zdkpLGdc5_1(.din(w_dff_B_abBCvjBt5_1),.dout(w_dff_B_zdkpLGdc5_1),.clk(gclk));
	jdff dff_B_JoeoQYl15_1(.din(w_dff_B_zdkpLGdc5_1),.dout(w_dff_B_JoeoQYl15_1),.clk(gclk));
	jdff dff_B_ywdPvI0A7_1(.din(w_dff_B_JoeoQYl15_1),.dout(w_dff_B_ywdPvI0A7_1),.clk(gclk));
	jdff dff_B_gBOEeCXE2_1(.din(w_dff_B_ywdPvI0A7_1),.dout(w_dff_B_gBOEeCXE2_1),.clk(gclk));
	jdff dff_B_kGQLwCQb2_1(.din(n383),.dout(w_dff_B_kGQLwCQb2_1),.clk(gclk));
	jdff dff_A_lOmWAwmn7_0(.dout(w_n317_0[0]),.din(w_dff_A_lOmWAwmn7_0),.clk(gclk));
	jdff dff_A_C8MyfKbz3_0(.dout(w_dff_A_lOmWAwmn7_0),.din(w_dff_A_C8MyfKbz3_0),.clk(gclk));
	jdff dff_A_bN5Kgzky8_0(.dout(w_dff_A_C8MyfKbz3_0),.din(w_dff_A_bN5Kgzky8_0),.clk(gclk));
	jdff dff_A_6FNsbAd11_0(.dout(w_dff_A_bN5Kgzky8_0),.din(w_dff_A_6FNsbAd11_0),.clk(gclk));
	jdff dff_A_A3eZGUtg0_0(.dout(w_dff_A_6FNsbAd11_0),.din(w_dff_A_A3eZGUtg0_0),.clk(gclk));
	jdff dff_A_60rmtUnQ1_0(.dout(w_dff_A_A3eZGUtg0_0),.din(w_dff_A_60rmtUnQ1_0),.clk(gclk));
	jdff dff_A_c4GuJAhG9_0(.dout(w_dff_A_60rmtUnQ1_0),.din(w_dff_A_c4GuJAhG9_0),.clk(gclk));
	jdff dff_A_PlPOWuLG1_0(.dout(w_dff_A_c4GuJAhG9_0),.din(w_dff_A_PlPOWuLG1_0),.clk(gclk));
	jdff dff_A_si98wfdP8_0(.dout(w_dff_A_PlPOWuLG1_0),.din(w_dff_A_si98wfdP8_0),.clk(gclk));
	jdff dff_A_kQXNzgLG6_0(.dout(w_dff_A_si98wfdP8_0),.din(w_dff_A_kQXNzgLG6_0),.clk(gclk));
	jdff dff_A_V6uivRY26_0(.dout(w_dff_A_kQXNzgLG6_0),.din(w_dff_A_V6uivRY26_0),.clk(gclk));
	jdff dff_A_OcrFrRTl0_0(.dout(w_dff_A_V6uivRY26_0),.din(w_dff_A_OcrFrRTl0_0),.clk(gclk));
	jdff dff_A_AhyO9wxh9_0(.dout(w_dff_A_OcrFrRTl0_0),.din(w_dff_A_AhyO9wxh9_0),.clk(gclk));
	jdff dff_A_0tAqT7jG1_0(.dout(w_dff_A_AhyO9wxh9_0),.din(w_dff_A_0tAqT7jG1_0),.clk(gclk));
	jdff dff_A_nAKTEXvw9_0(.dout(w_dff_A_0tAqT7jG1_0),.din(w_dff_A_nAKTEXvw9_0),.clk(gclk));
	jdff dff_A_XWLuz7rt9_0(.dout(w_dff_A_nAKTEXvw9_0),.din(w_dff_A_XWLuz7rt9_0),.clk(gclk));
	jdff dff_A_jK0aNFSy9_0(.dout(w_dff_A_XWLuz7rt9_0),.din(w_dff_A_jK0aNFSy9_0),.clk(gclk));
	jdff dff_A_ynk5SylS1_0(.dout(w_dff_A_jK0aNFSy9_0),.din(w_dff_A_ynk5SylS1_0),.clk(gclk));
	jdff dff_A_koF0IBwu4_0(.dout(w_dff_A_ynk5SylS1_0),.din(w_dff_A_koF0IBwu4_0),.clk(gclk));
	jdff dff_A_2IZZW4I74_0(.dout(w_dff_A_koF0IBwu4_0),.din(w_dff_A_2IZZW4I74_0),.clk(gclk));
	jdff dff_A_XaSxk0By8_0(.dout(w_dff_A_2IZZW4I74_0),.din(w_dff_A_XaSxk0By8_0),.clk(gclk));
	jdff dff_A_pHBec1sl8_0(.dout(w_dff_A_XaSxk0By8_0),.din(w_dff_A_pHBec1sl8_0),.clk(gclk));
	jdff dff_A_t5WXf41F4_0(.dout(w_dff_A_pHBec1sl8_0),.din(w_dff_A_t5WXf41F4_0),.clk(gclk));
	jdff dff_A_Blq0YXyK8_0(.dout(w_dff_A_t5WXf41F4_0),.din(w_dff_A_Blq0YXyK8_0),.clk(gclk));
	jdff dff_A_9otDpVqf0_0(.dout(w_dff_A_Blq0YXyK8_0),.din(w_dff_A_9otDpVqf0_0),.clk(gclk));
	jdff dff_A_RVsGh9gK2_1(.dout(w_n377_0[1]),.din(w_dff_A_RVsGh9gK2_1),.clk(gclk));
	jdff dff_B_ho3VH9op0_1(.din(n324),.dout(w_dff_B_ho3VH9op0_1),.clk(gclk));
	jdff dff_B_Fz5biCnP3_1(.din(w_dff_B_ho3VH9op0_1),.dout(w_dff_B_Fz5biCnP3_1),.clk(gclk));
	jdff dff_B_aoBeiQaW0_1(.din(w_dff_B_Fz5biCnP3_1),.dout(w_dff_B_aoBeiQaW0_1),.clk(gclk));
	jdff dff_B_zXm3zxue6_1(.din(w_dff_B_aoBeiQaW0_1),.dout(w_dff_B_zXm3zxue6_1),.clk(gclk));
	jdff dff_B_Js4dWb0A8_1(.din(w_dff_B_zXm3zxue6_1),.dout(w_dff_B_Js4dWb0A8_1),.clk(gclk));
	jdff dff_B_XtgDgxAH8_1(.din(w_dff_B_Js4dWb0A8_1),.dout(w_dff_B_XtgDgxAH8_1),.clk(gclk));
	jdff dff_B_iFkoXCaA1_1(.din(w_dff_B_XtgDgxAH8_1),.dout(w_dff_B_iFkoXCaA1_1),.clk(gclk));
	jdff dff_B_MapPrYeL5_1(.din(w_dff_B_iFkoXCaA1_1),.dout(w_dff_B_MapPrYeL5_1),.clk(gclk));
	jdff dff_B_dYwt28XJ1_1(.din(w_dff_B_MapPrYeL5_1),.dout(w_dff_B_dYwt28XJ1_1),.clk(gclk));
	jdff dff_B_IcoHR6Jl6_1(.din(w_dff_B_dYwt28XJ1_1),.dout(w_dff_B_IcoHR6Jl6_1),.clk(gclk));
	jdff dff_B_4zcNiNTF9_1(.din(w_dff_B_IcoHR6Jl6_1),.dout(w_dff_B_4zcNiNTF9_1),.clk(gclk));
	jdff dff_B_ekmokFYU8_1(.din(w_dff_B_4zcNiNTF9_1),.dout(w_dff_B_ekmokFYU8_1),.clk(gclk));
	jdff dff_B_BU0okkuW7_1(.din(w_dff_B_ekmokFYU8_1),.dout(w_dff_B_BU0okkuW7_1),.clk(gclk));
	jdff dff_B_D2HUPqIi1_1(.din(w_dff_B_BU0okkuW7_1),.dout(w_dff_B_D2HUPqIi1_1),.clk(gclk));
	jdff dff_B_foJYmLVh5_1(.din(w_dff_B_D2HUPqIi1_1),.dout(w_dff_B_foJYmLVh5_1),.clk(gclk));
	jdff dff_B_luqDlp972_1(.din(w_dff_B_foJYmLVh5_1),.dout(w_dff_B_luqDlp972_1),.clk(gclk));
	jdff dff_B_woYQI3Xo1_1(.din(w_dff_B_luqDlp972_1),.dout(w_dff_B_woYQI3Xo1_1),.clk(gclk));
	jdff dff_B_DWYYMhFN1_1(.din(w_dff_B_woYQI3Xo1_1),.dout(w_dff_B_DWYYMhFN1_1),.clk(gclk));
	jdff dff_B_2KBAuhsx4_1(.din(w_dff_B_DWYYMhFN1_1),.dout(w_dff_B_2KBAuhsx4_1),.clk(gclk));
	jdff dff_B_svZT3w2m4_1(.din(w_dff_B_2KBAuhsx4_1),.dout(w_dff_B_svZT3w2m4_1),.clk(gclk));
	jdff dff_B_eZQ8FN4T1_1(.din(w_dff_B_svZT3w2m4_1),.dout(w_dff_B_eZQ8FN4T1_1),.clk(gclk));
	jdff dff_B_KXgzlV1M9_1(.din(n320),.dout(w_dff_B_KXgzlV1M9_1),.clk(gclk));
	jdff dff_A_J7WOjswY8_0(.dout(w_n261_0[0]),.din(w_dff_A_J7WOjswY8_0),.clk(gclk));
	jdff dff_A_uL7sbdPp1_0(.dout(w_dff_A_J7WOjswY8_0),.din(w_dff_A_uL7sbdPp1_0),.clk(gclk));
	jdff dff_A_u2OnqcI40_0(.dout(w_dff_A_uL7sbdPp1_0),.din(w_dff_A_u2OnqcI40_0),.clk(gclk));
	jdff dff_A_3HCtycP24_0(.dout(w_dff_A_u2OnqcI40_0),.din(w_dff_A_3HCtycP24_0),.clk(gclk));
	jdff dff_A_Asf8COAB8_0(.dout(w_dff_A_3HCtycP24_0),.din(w_dff_A_Asf8COAB8_0),.clk(gclk));
	jdff dff_A_d6buk1457_0(.dout(w_dff_A_Asf8COAB8_0),.din(w_dff_A_d6buk1457_0),.clk(gclk));
	jdff dff_A_KHgypmyQ1_0(.dout(w_dff_A_d6buk1457_0),.din(w_dff_A_KHgypmyQ1_0),.clk(gclk));
	jdff dff_A_miRXi02Y2_0(.dout(w_dff_A_KHgypmyQ1_0),.din(w_dff_A_miRXi02Y2_0),.clk(gclk));
	jdff dff_A_9uKv9i878_0(.dout(w_dff_A_miRXi02Y2_0),.din(w_dff_A_9uKv9i878_0),.clk(gclk));
	jdff dff_A_5gmCLYxM3_0(.dout(w_dff_A_9uKv9i878_0),.din(w_dff_A_5gmCLYxM3_0),.clk(gclk));
	jdff dff_A_vnXmfF1G1_0(.dout(w_dff_A_5gmCLYxM3_0),.din(w_dff_A_vnXmfF1G1_0),.clk(gclk));
	jdff dff_A_zlElvV4I0_0(.dout(w_dff_A_vnXmfF1G1_0),.din(w_dff_A_zlElvV4I0_0),.clk(gclk));
	jdff dff_A_5URrfS203_0(.dout(w_dff_A_zlElvV4I0_0),.din(w_dff_A_5URrfS203_0),.clk(gclk));
	jdff dff_A_e1pVPcMY9_0(.dout(w_dff_A_5URrfS203_0),.din(w_dff_A_e1pVPcMY9_0),.clk(gclk));
	jdff dff_A_e9IMCj5g1_0(.dout(w_dff_A_e1pVPcMY9_0),.din(w_dff_A_e9IMCj5g1_0),.clk(gclk));
	jdff dff_A_RxNTvOhv2_0(.dout(w_dff_A_e9IMCj5g1_0),.din(w_dff_A_RxNTvOhv2_0),.clk(gclk));
	jdff dff_A_GvO1V44g7_0(.dout(w_dff_A_RxNTvOhv2_0),.din(w_dff_A_GvO1V44g7_0),.clk(gclk));
	jdff dff_A_E4SLNtuM0_0(.dout(w_dff_A_GvO1V44g7_0),.din(w_dff_A_E4SLNtuM0_0),.clk(gclk));
	jdff dff_A_cqj1vMHG2_0(.dout(w_dff_A_E4SLNtuM0_0),.din(w_dff_A_cqj1vMHG2_0),.clk(gclk));
	jdff dff_A_TWxyknpV1_0(.dout(w_dff_A_cqj1vMHG2_0),.din(w_dff_A_TWxyknpV1_0),.clk(gclk));
	jdff dff_A_N65SNwsB3_0(.dout(w_dff_A_TWxyknpV1_0),.din(w_dff_A_N65SNwsB3_0),.clk(gclk));
	jdff dff_A_gM2LXppr0_0(.dout(w_dff_A_N65SNwsB3_0),.din(w_dff_A_gM2LXppr0_0),.clk(gclk));
	jdff dff_A_E2AfKQGi1_1(.dout(w_n314_0[1]),.din(w_dff_A_E2AfKQGi1_1),.clk(gclk));
	jdff dff_B_LkzXASl69_1(.din(n268),.dout(w_dff_B_LkzXASl69_1),.clk(gclk));
	jdff dff_B_QBY03YW21_1(.din(w_dff_B_LkzXASl69_1),.dout(w_dff_B_QBY03YW21_1),.clk(gclk));
	jdff dff_B_znxiZW4c3_1(.din(w_dff_B_QBY03YW21_1),.dout(w_dff_B_znxiZW4c3_1),.clk(gclk));
	jdff dff_B_00jPaK7g9_1(.din(w_dff_B_znxiZW4c3_1),.dout(w_dff_B_00jPaK7g9_1),.clk(gclk));
	jdff dff_B_r5P06Tk20_1(.din(w_dff_B_00jPaK7g9_1),.dout(w_dff_B_r5P06Tk20_1),.clk(gclk));
	jdff dff_B_VwUw66dR5_1(.din(w_dff_B_r5P06Tk20_1),.dout(w_dff_B_VwUw66dR5_1),.clk(gclk));
	jdff dff_B_JVNXc6vS4_1(.din(w_dff_B_VwUw66dR5_1),.dout(w_dff_B_JVNXc6vS4_1),.clk(gclk));
	jdff dff_B_cByGxDKc2_1(.din(w_dff_B_JVNXc6vS4_1),.dout(w_dff_B_cByGxDKc2_1),.clk(gclk));
	jdff dff_B_5ugC1HHl1_1(.din(w_dff_B_cByGxDKc2_1),.dout(w_dff_B_5ugC1HHl1_1),.clk(gclk));
	jdff dff_B_I1qL3ToX2_1(.din(w_dff_B_5ugC1HHl1_1),.dout(w_dff_B_I1qL3ToX2_1),.clk(gclk));
	jdff dff_B_cuYa9qI68_1(.din(w_dff_B_I1qL3ToX2_1),.dout(w_dff_B_cuYa9qI68_1),.clk(gclk));
	jdff dff_B_HdWi1d3R2_1(.din(w_dff_B_cuYa9qI68_1),.dout(w_dff_B_HdWi1d3R2_1),.clk(gclk));
	jdff dff_B_f6gA8plr8_1(.din(w_dff_B_HdWi1d3R2_1),.dout(w_dff_B_f6gA8plr8_1),.clk(gclk));
	jdff dff_B_ydGDNvnU7_1(.din(w_dff_B_f6gA8plr8_1),.dout(w_dff_B_ydGDNvnU7_1),.clk(gclk));
	jdff dff_B_Xh79EhiN2_1(.din(w_dff_B_ydGDNvnU7_1),.dout(w_dff_B_Xh79EhiN2_1),.clk(gclk));
	jdff dff_B_1YaZ1wIn0_1(.din(w_dff_B_Xh79EhiN2_1),.dout(w_dff_B_1YaZ1wIn0_1),.clk(gclk));
	jdff dff_B_X3u6fkyO1_1(.din(w_dff_B_1YaZ1wIn0_1),.dout(w_dff_B_X3u6fkyO1_1),.clk(gclk));
	jdff dff_B_NwoMSljy8_1(.din(w_dff_B_X3u6fkyO1_1),.dout(w_dff_B_NwoMSljy8_1),.clk(gclk));
	jdff dff_B_yHoAoE6P4_1(.din(n264),.dout(w_dff_B_yHoAoE6P4_1),.clk(gclk));
	jdff dff_A_F6HOCl9Z1_0(.dout(w_n212_0[0]),.din(w_dff_A_F6HOCl9Z1_0),.clk(gclk));
	jdff dff_A_NLMVx5xN4_0(.dout(w_dff_A_F6HOCl9Z1_0),.din(w_dff_A_NLMVx5xN4_0),.clk(gclk));
	jdff dff_A_SdbbVui39_0(.dout(w_dff_A_NLMVx5xN4_0),.din(w_dff_A_SdbbVui39_0),.clk(gclk));
	jdff dff_A_ibJZI8Pz8_0(.dout(w_dff_A_SdbbVui39_0),.din(w_dff_A_ibJZI8Pz8_0),.clk(gclk));
	jdff dff_A_NEDW3c189_0(.dout(w_dff_A_ibJZI8Pz8_0),.din(w_dff_A_NEDW3c189_0),.clk(gclk));
	jdff dff_A_DiDbtBgY6_0(.dout(w_dff_A_NEDW3c189_0),.din(w_dff_A_DiDbtBgY6_0),.clk(gclk));
	jdff dff_A_d9g259gG9_0(.dout(w_dff_A_DiDbtBgY6_0),.din(w_dff_A_d9g259gG9_0),.clk(gclk));
	jdff dff_A_CVfikeBg8_0(.dout(w_dff_A_d9g259gG9_0),.din(w_dff_A_CVfikeBg8_0),.clk(gclk));
	jdff dff_A_nOrqZHBH0_0(.dout(w_dff_A_CVfikeBg8_0),.din(w_dff_A_nOrqZHBH0_0),.clk(gclk));
	jdff dff_A_2b7vdG0w9_0(.dout(w_dff_A_nOrqZHBH0_0),.din(w_dff_A_2b7vdG0w9_0),.clk(gclk));
	jdff dff_A_m0njP2kO6_0(.dout(w_dff_A_2b7vdG0w9_0),.din(w_dff_A_m0njP2kO6_0),.clk(gclk));
	jdff dff_A_q0Nn6ixV0_0(.dout(w_dff_A_m0njP2kO6_0),.din(w_dff_A_q0Nn6ixV0_0),.clk(gclk));
	jdff dff_A_lMZKy4LX9_0(.dout(w_dff_A_q0Nn6ixV0_0),.din(w_dff_A_lMZKy4LX9_0),.clk(gclk));
	jdff dff_A_GQIVikUo5_0(.dout(w_dff_A_lMZKy4LX9_0),.din(w_dff_A_GQIVikUo5_0),.clk(gclk));
	jdff dff_A_uVIXtaQe2_0(.dout(w_dff_A_GQIVikUo5_0),.din(w_dff_A_uVIXtaQe2_0),.clk(gclk));
	jdff dff_A_SFM34Hx82_0(.dout(w_dff_A_uVIXtaQe2_0),.din(w_dff_A_SFM34Hx82_0),.clk(gclk));
	jdff dff_A_MgZ8Tsoj1_0(.dout(w_dff_A_SFM34Hx82_0),.din(w_dff_A_MgZ8Tsoj1_0),.clk(gclk));
	jdff dff_A_uOxkyAHE4_0(.dout(w_dff_A_MgZ8Tsoj1_0),.din(w_dff_A_uOxkyAHE4_0),.clk(gclk));
	jdff dff_A_nXyfF5ZW7_0(.dout(w_dff_A_uOxkyAHE4_0),.din(w_dff_A_nXyfF5ZW7_0),.clk(gclk));
	jdff dff_A_ujIduFVv2_1(.dout(w_n258_0[1]),.din(w_dff_A_ujIduFVv2_1),.clk(gclk));
	jdff dff_B_uQa7je7J4_1(.din(n219),.dout(w_dff_B_uQa7je7J4_1),.clk(gclk));
	jdff dff_B_0dXH419U3_1(.din(w_dff_B_uQa7je7J4_1),.dout(w_dff_B_0dXH419U3_1),.clk(gclk));
	jdff dff_B_uVc8stqu4_1(.din(w_dff_B_0dXH419U3_1),.dout(w_dff_B_uVc8stqu4_1),.clk(gclk));
	jdff dff_B_vTTMyKL42_1(.din(w_dff_B_uVc8stqu4_1),.dout(w_dff_B_vTTMyKL42_1),.clk(gclk));
	jdff dff_B_IkNeszDg4_1(.din(w_dff_B_vTTMyKL42_1),.dout(w_dff_B_IkNeszDg4_1),.clk(gclk));
	jdff dff_B_QEH6NRHJ8_1(.din(w_dff_B_IkNeszDg4_1),.dout(w_dff_B_QEH6NRHJ8_1),.clk(gclk));
	jdff dff_B_9HLorpzB3_1(.din(w_dff_B_QEH6NRHJ8_1),.dout(w_dff_B_9HLorpzB3_1),.clk(gclk));
	jdff dff_B_REtC54pC2_1(.din(w_dff_B_9HLorpzB3_1),.dout(w_dff_B_REtC54pC2_1),.clk(gclk));
	jdff dff_B_7Cz5Z4Kr4_1(.din(w_dff_B_REtC54pC2_1),.dout(w_dff_B_7Cz5Z4Kr4_1),.clk(gclk));
	jdff dff_B_RcFjeqnT6_1(.din(w_dff_B_7Cz5Z4Kr4_1),.dout(w_dff_B_RcFjeqnT6_1),.clk(gclk));
	jdff dff_B_VmXVDCV31_1(.din(w_dff_B_RcFjeqnT6_1),.dout(w_dff_B_VmXVDCV31_1),.clk(gclk));
	jdff dff_B_HUFtEnqY0_1(.din(w_dff_B_VmXVDCV31_1),.dout(w_dff_B_HUFtEnqY0_1),.clk(gclk));
	jdff dff_B_HEx40znw5_1(.din(w_dff_B_HUFtEnqY0_1),.dout(w_dff_B_HEx40znw5_1),.clk(gclk));
	jdff dff_B_NFEyZqW68_1(.din(w_dff_B_HEx40znw5_1),.dout(w_dff_B_NFEyZqW68_1),.clk(gclk));
	jdff dff_B_d8EbkTxD8_1(.din(w_dff_B_NFEyZqW68_1),.dout(w_dff_B_d8EbkTxD8_1),.clk(gclk));
	jdff dff_B_4IAinCvK4_1(.din(n215),.dout(w_dff_B_4IAinCvK4_1),.clk(gclk));
	jdff dff_A_sIr3t28d7_0(.dout(w_n170_0[0]),.din(w_dff_A_sIr3t28d7_0),.clk(gclk));
	jdff dff_A_9iyz4Pte6_0(.dout(w_dff_A_sIr3t28d7_0),.din(w_dff_A_9iyz4Pte6_0),.clk(gclk));
	jdff dff_A_R4Oz2l9q0_0(.dout(w_dff_A_9iyz4Pte6_0),.din(w_dff_A_R4Oz2l9q0_0),.clk(gclk));
	jdff dff_A_FjSEhMfU8_0(.dout(w_dff_A_R4Oz2l9q0_0),.din(w_dff_A_FjSEhMfU8_0),.clk(gclk));
	jdff dff_A_j1Xv7zmb2_0(.dout(w_dff_A_FjSEhMfU8_0),.din(w_dff_A_j1Xv7zmb2_0),.clk(gclk));
	jdff dff_A_L382okfo6_0(.dout(w_dff_A_j1Xv7zmb2_0),.din(w_dff_A_L382okfo6_0),.clk(gclk));
	jdff dff_A_l9nhwDHr8_0(.dout(w_dff_A_L382okfo6_0),.din(w_dff_A_l9nhwDHr8_0),.clk(gclk));
	jdff dff_A_OOlRk1Ny8_0(.dout(w_dff_A_l9nhwDHr8_0),.din(w_dff_A_OOlRk1Ny8_0),.clk(gclk));
	jdff dff_A_gUhkwX6k5_0(.dout(w_dff_A_OOlRk1Ny8_0),.din(w_dff_A_gUhkwX6k5_0),.clk(gclk));
	jdff dff_A_938kOzp87_0(.dout(w_dff_A_gUhkwX6k5_0),.din(w_dff_A_938kOzp87_0),.clk(gclk));
	jdff dff_A_BeJ7GYUl7_0(.dout(w_dff_A_938kOzp87_0),.din(w_dff_A_BeJ7GYUl7_0),.clk(gclk));
	jdff dff_A_4YMDY7en1_0(.dout(w_dff_A_BeJ7GYUl7_0),.din(w_dff_A_4YMDY7en1_0),.clk(gclk));
	jdff dff_A_rjLEFNFV8_0(.dout(w_dff_A_4YMDY7en1_0),.din(w_dff_A_rjLEFNFV8_0),.clk(gclk));
	jdff dff_A_vUPAaQ5i2_0(.dout(w_dff_A_rjLEFNFV8_0),.din(w_dff_A_vUPAaQ5i2_0),.clk(gclk));
	jdff dff_A_gs5bTWi95_0(.dout(w_dff_A_vUPAaQ5i2_0),.din(w_dff_A_gs5bTWi95_0),.clk(gclk));
	jdff dff_A_3paX2inR4_0(.dout(w_dff_A_gs5bTWi95_0),.din(w_dff_A_3paX2inR4_0),.clk(gclk));
	jdff dff_A_2h6ak3GK4_1(.dout(w_n209_0[1]),.din(w_dff_A_2h6ak3GK4_1),.clk(gclk));
	jdff dff_B_O1nL2Eme5_1(.din(n177),.dout(w_dff_B_O1nL2Eme5_1),.clk(gclk));
	jdff dff_B_4Dq2Ul1G2_1(.din(w_dff_B_O1nL2Eme5_1),.dout(w_dff_B_4Dq2Ul1G2_1),.clk(gclk));
	jdff dff_B_wXjGVgAc2_1(.din(w_dff_B_4Dq2Ul1G2_1),.dout(w_dff_B_wXjGVgAc2_1),.clk(gclk));
	jdff dff_B_sTcbt0Xc1_1(.din(w_dff_B_wXjGVgAc2_1),.dout(w_dff_B_sTcbt0Xc1_1),.clk(gclk));
	jdff dff_B_8ludC52q6_1(.din(w_dff_B_sTcbt0Xc1_1),.dout(w_dff_B_8ludC52q6_1),.clk(gclk));
	jdff dff_B_7MFV8VOy2_1(.din(w_dff_B_8ludC52q6_1),.dout(w_dff_B_7MFV8VOy2_1),.clk(gclk));
	jdff dff_B_b2JeRQLK7_1(.din(w_dff_B_7MFV8VOy2_1),.dout(w_dff_B_b2JeRQLK7_1),.clk(gclk));
	jdff dff_B_6qA0x1Dt3_1(.din(w_dff_B_b2JeRQLK7_1),.dout(w_dff_B_6qA0x1Dt3_1),.clk(gclk));
	jdff dff_B_cgCwIWBN1_1(.din(w_dff_B_6qA0x1Dt3_1),.dout(w_dff_B_cgCwIWBN1_1),.clk(gclk));
	jdff dff_B_9Ckz7EOK7_1(.din(w_dff_B_cgCwIWBN1_1),.dout(w_dff_B_9Ckz7EOK7_1),.clk(gclk));
	jdff dff_B_aJJ7xfrT9_1(.din(w_dff_B_9Ckz7EOK7_1),.dout(w_dff_B_aJJ7xfrT9_1),.clk(gclk));
	jdff dff_B_wDNz3IFj5_1(.din(w_dff_B_aJJ7xfrT9_1),.dout(w_dff_B_wDNz3IFj5_1),.clk(gclk));
	jdff dff_B_e5SXL19y3_1(.din(n173),.dout(w_dff_B_e5SXL19y3_1),.clk(gclk));
	jdff dff_A_yOPOHtc53_0(.dout(w_n135_0[0]),.din(w_dff_A_yOPOHtc53_0),.clk(gclk));
	jdff dff_A_hBEkpYuJ6_0(.dout(w_dff_A_yOPOHtc53_0),.din(w_dff_A_hBEkpYuJ6_0),.clk(gclk));
	jdff dff_A_bUeLdpSR5_0(.dout(w_dff_A_hBEkpYuJ6_0),.din(w_dff_A_bUeLdpSR5_0),.clk(gclk));
	jdff dff_A_cH1xxg165_0(.dout(w_dff_A_bUeLdpSR5_0),.din(w_dff_A_cH1xxg165_0),.clk(gclk));
	jdff dff_A_d1p6rDNR2_0(.dout(w_dff_A_cH1xxg165_0),.din(w_dff_A_d1p6rDNR2_0),.clk(gclk));
	jdff dff_A_DmIQjyM20_0(.dout(w_dff_A_d1p6rDNR2_0),.din(w_dff_A_DmIQjyM20_0),.clk(gclk));
	jdff dff_A_d74gFXDP1_0(.dout(w_dff_A_DmIQjyM20_0),.din(w_dff_A_d74gFXDP1_0),.clk(gclk));
	jdff dff_A_xTEMoy1Y5_0(.dout(w_dff_A_d74gFXDP1_0),.din(w_dff_A_xTEMoy1Y5_0),.clk(gclk));
	jdff dff_A_HnoeuEKP9_0(.dout(w_dff_A_xTEMoy1Y5_0),.din(w_dff_A_HnoeuEKP9_0),.clk(gclk));
	jdff dff_A_BT1MZ7Sz0_0(.dout(w_dff_A_HnoeuEKP9_0),.din(w_dff_A_BT1MZ7Sz0_0),.clk(gclk));
	jdff dff_A_aHaSUFTv5_0(.dout(w_dff_A_BT1MZ7Sz0_0),.din(w_dff_A_aHaSUFTv5_0),.clk(gclk));
	jdff dff_A_8WGJXl8K4_0(.dout(w_dff_A_aHaSUFTv5_0),.din(w_dff_A_8WGJXl8K4_0),.clk(gclk));
	jdff dff_A_9WrAOST24_0(.dout(w_dff_A_8WGJXl8K4_0),.din(w_dff_A_9WrAOST24_0),.clk(gclk));
	jdff dff_A_RKyRjln93_1(.dout(w_n167_0[1]),.din(w_dff_A_RKyRjln93_1),.clk(gclk));
	jdff dff_B_l7CIwixh9_1(.din(n142),.dout(w_dff_B_l7CIwixh9_1),.clk(gclk));
	jdff dff_B_I462lvCz2_1(.din(w_dff_B_l7CIwixh9_1),.dout(w_dff_B_I462lvCz2_1),.clk(gclk));
	jdff dff_B_58oxfOiv9_1(.din(w_dff_B_I462lvCz2_1),.dout(w_dff_B_58oxfOiv9_1),.clk(gclk));
	jdff dff_B_fSed0ote5_1(.din(w_dff_B_58oxfOiv9_1),.dout(w_dff_B_fSed0ote5_1),.clk(gclk));
	jdff dff_B_7ga4towO6_1(.din(w_dff_B_fSed0ote5_1),.dout(w_dff_B_7ga4towO6_1),.clk(gclk));
	jdff dff_B_HHOcYcgn9_1(.din(w_dff_B_7ga4towO6_1),.dout(w_dff_B_HHOcYcgn9_1),.clk(gclk));
	jdff dff_B_D2ySSSay6_1(.din(w_dff_B_HHOcYcgn9_1),.dout(w_dff_B_D2ySSSay6_1),.clk(gclk));
	jdff dff_B_CsC0BIYR3_1(.din(w_dff_B_D2ySSSay6_1),.dout(w_dff_B_CsC0BIYR3_1),.clk(gclk));
	jdff dff_B_41TCNUGG3_1(.din(w_dff_B_CsC0BIYR3_1),.dout(w_dff_B_41TCNUGG3_1),.clk(gclk));
	jdff dff_B_ZBGSYhqQ2_1(.din(n138),.dout(w_dff_B_ZBGSYhqQ2_1),.clk(gclk));
	jdff dff_A_I9I1WVz00_0(.dout(w_n106_0[0]),.din(w_dff_A_I9I1WVz00_0),.clk(gclk));
	jdff dff_A_Kwk6TNJB8_0(.dout(w_dff_A_I9I1WVz00_0),.din(w_dff_A_Kwk6TNJB8_0),.clk(gclk));
	jdff dff_A_5uHSAbGh7_0(.dout(w_dff_A_Kwk6TNJB8_0),.din(w_dff_A_5uHSAbGh7_0),.clk(gclk));
	jdff dff_A_adtHeypL6_0(.dout(w_dff_A_5uHSAbGh7_0),.din(w_dff_A_adtHeypL6_0),.clk(gclk));
	jdff dff_A_Dlr3XBF36_0(.dout(w_dff_A_adtHeypL6_0),.din(w_dff_A_Dlr3XBF36_0),.clk(gclk));
	jdff dff_A_E1i8Mt5B3_0(.dout(w_dff_A_Dlr3XBF36_0),.din(w_dff_A_E1i8Mt5B3_0),.clk(gclk));
	jdff dff_A_QAldSDto2_0(.dout(w_dff_A_E1i8Mt5B3_0),.din(w_dff_A_QAldSDto2_0),.clk(gclk));
	jdff dff_A_KPirdrdm9_0(.dout(w_dff_A_QAldSDto2_0),.din(w_dff_A_KPirdrdm9_0),.clk(gclk));
	jdff dff_A_QHbmduf29_0(.dout(w_dff_A_KPirdrdm9_0),.din(w_dff_A_QHbmduf29_0),.clk(gclk));
	jdff dff_A_qdcJQ49M1_0(.dout(w_dff_A_QHbmduf29_0),.din(w_dff_A_qdcJQ49M1_0),.clk(gclk));
	jdff dff_A_hivLiakV5_1(.dout(w_n132_0[1]),.din(w_dff_A_hivLiakV5_1),.clk(gclk));
	jdff dff_B_vznmlZVm5_1(.din(n113),.dout(w_dff_B_vznmlZVm5_1),.clk(gclk));
	jdff dff_B_1XKIj6og3_1(.din(w_dff_B_vznmlZVm5_1),.dout(w_dff_B_1XKIj6og3_1),.clk(gclk));
	jdff dff_B_jLPMgnHZ4_1(.din(w_dff_B_1XKIj6og3_1),.dout(w_dff_B_jLPMgnHZ4_1),.clk(gclk));
	jdff dff_B_yhm7Gakg5_1(.din(w_dff_B_jLPMgnHZ4_1),.dout(w_dff_B_yhm7Gakg5_1),.clk(gclk));
	jdff dff_B_8CmJTX035_1(.din(w_dff_B_yhm7Gakg5_1),.dout(w_dff_B_8CmJTX035_1),.clk(gclk));
	jdff dff_B_gzcghbfG9_1(.din(w_dff_B_8CmJTX035_1),.dout(w_dff_B_gzcghbfG9_1),.clk(gclk));
	jdff dff_B_MwfEWbpP9_1(.din(n109),.dout(w_dff_B_MwfEWbpP9_1),.clk(gclk));
	jdff dff_A_DecIt21K5_0(.dout(w_n86_0[0]),.din(w_dff_A_DecIt21K5_0),.clk(gclk));
	jdff dff_A_a9AaLAWx9_0(.dout(w_dff_A_DecIt21K5_0),.din(w_dff_A_a9AaLAWx9_0),.clk(gclk));
	jdff dff_A_1c9raQmS9_0(.dout(w_dff_A_a9AaLAWx9_0),.din(w_dff_A_1c9raQmS9_0),.clk(gclk));
	jdff dff_A_gVIRcJBG4_0(.dout(w_dff_A_1c9raQmS9_0),.din(w_dff_A_gVIRcJBG4_0),.clk(gclk));
	jdff dff_A_ioR6XyE70_0(.dout(w_dff_A_gVIRcJBG4_0),.din(w_dff_A_ioR6XyE70_0),.clk(gclk));
	jdff dff_A_o4KfhgMK0_0(.dout(w_dff_A_ioR6XyE70_0),.din(w_dff_A_o4KfhgMK0_0),.clk(gclk));
	jdff dff_A_d8DAIhbV2_0(.dout(w_dff_A_o4KfhgMK0_0),.din(w_dff_A_d8DAIhbV2_0),.clk(gclk));
	jdff dff_A_MSEJUAI97_1(.dout(w_n103_0[1]),.din(w_dff_A_MSEJUAI97_1),.clk(gclk));
	jdff dff_B_6M5aIzqv6_1(.din(n92),.dout(w_dff_B_6M5aIzqv6_1),.clk(gclk));
	jdff dff_B_ifezlAmu9_1(.din(w_dff_B_6M5aIzqv6_1),.dout(w_dff_B_ifezlAmu9_1),.clk(gclk));
	jdff dff_B_VxStCGKZ2_1(.din(w_dff_B_ifezlAmu9_1),.dout(w_dff_B_VxStCGKZ2_1),.clk(gclk));
	jdff dff_B_UGGTIAOT5_1(.din(n88),.dout(w_dff_B_UGGTIAOT5_1),.clk(gclk));
	jdff dff_B_DaDNKJQD9_2(.din(n67),.dout(w_dff_B_DaDNKJQD9_2),.clk(gclk));
	jdff dff_A_VvcuaMFH7_0(.dout(w_n75_0[0]),.din(w_dff_A_VvcuaMFH7_0),.clk(gclk));
	jdff dff_A_mKL79bUP7_0(.dout(w_dff_A_VvcuaMFH7_0),.din(w_dff_A_mKL79bUP7_0),.clk(gclk));
	jdff dff_A_HiWWr8kQ9_0(.dout(w_dff_A_mKL79bUP7_0),.din(w_dff_A_HiWWr8kQ9_0),.clk(gclk));
	jdff dff_A_QnJKV9jW3_0(.dout(w_dff_A_HiWWr8kQ9_0),.din(w_dff_A_QnJKV9jW3_0),.clk(gclk));
	jdff dff_B_4AVndoHp8_0(.din(n82),.dout(w_dff_B_4AVndoHp8_0),.clk(gclk));
	jdff dff_A_sICFtYLJ6_0(.dout(w_n66_0[0]),.din(w_dff_A_sICFtYLJ6_0),.clk(gclk));
	jdff dff_A_7PsyB8RX7_0(.dout(w_dff_A_sICFtYLJ6_0),.din(w_dff_A_7PsyB8RX7_0),.clk(gclk));
	jdff dff_A_g7Cqca0B3_1(.dout(w_n1108_0[1]),.din(w_dff_A_g7Cqca0B3_1),.clk(gclk));
	jdff dff_B_kUX2dQoU1_1(.din(n1014),.dout(w_dff_B_kUX2dQoU1_1),.clk(gclk));
	jdff dff_B_uh08qkyA8_2(.din(n911),.dout(w_dff_B_uh08qkyA8_2),.clk(gclk));
	jdff dff_B_67SyN4BX0_2(.din(w_dff_B_uh08qkyA8_2),.dout(w_dff_B_67SyN4BX0_2),.clk(gclk));
	jdff dff_B_3n1TvbgO3_2(.din(w_dff_B_67SyN4BX0_2),.dout(w_dff_B_3n1TvbgO3_2),.clk(gclk));
	jdff dff_B_E23RCO5t0_2(.din(w_dff_B_3n1TvbgO3_2),.dout(w_dff_B_E23RCO5t0_2),.clk(gclk));
	jdff dff_B_kmhO2PBp8_2(.din(w_dff_B_E23RCO5t0_2),.dout(w_dff_B_kmhO2PBp8_2),.clk(gclk));
	jdff dff_B_wpKlsJpS2_2(.din(w_dff_B_kmhO2PBp8_2),.dout(w_dff_B_wpKlsJpS2_2),.clk(gclk));
	jdff dff_B_uJhi3PER3_2(.din(w_dff_B_wpKlsJpS2_2),.dout(w_dff_B_uJhi3PER3_2),.clk(gclk));
	jdff dff_B_Rl3aCQEo4_2(.din(w_dff_B_uJhi3PER3_2),.dout(w_dff_B_Rl3aCQEo4_2),.clk(gclk));
	jdff dff_B_lXBkLMC50_2(.din(w_dff_B_Rl3aCQEo4_2),.dout(w_dff_B_lXBkLMC50_2),.clk(gclk));
	jdff dff_B_rRhLN53z2_2(.din(w_dff_B_lXBkLMC50_2),.dout(w_dff_B_rRhLN53z2_2),.clk(gclk));
	jdff dff_B_fpVYwdWF7_2(.din(w_dff_B_rRhLN53z2_2),.dout(w_dff_B_fpVYwdWF7_2),.clk(gclk));
	jdff dff_B_D7IdrbQv4_2(.din(w_dff_B_fpVYwdWF7_2),.dout(w_dff_B_D7IdrbQv4_2),.clk(gclk));
	jdff dff_B_u9ZhCgMi0_2(.din(w_dff_B_D7IdrbQv4_2),.dout(w_dff_B_u9ZhCgMi0_2),.clk(gclk));
	jdff dff_B_oceqJu7P4_2(.din(w_dff_B_u9ZhCgMi0_2),.dout(w_dff_B_oceqJu7P4_2),.clk(gclk));
	jdff dff_B_JFQ8KwRR2_2(.din(w_dff_B_oceqJu7P4_2),.dout(w_dff_B_JFQ8KwRR2_2),.clk(gclk));
	jdff dff_B_jYYsO1in3_2(.din(w_dff_B_JFQ8KwRR2_2),.dout(w_dff_B_jYYsO1in3_2),.clk(gclk));
	jdff dff_B_2OWlbafw5_2(.din(w_dff_B_jYYsO1in3_2),.dout(w_dff_B_2OWlbafw5_2),.clk(gclk));
	jdff dff_B_WcVNyhwX7_2(.din(w_dff_B_2OWlbafw5_2),.dout(w_dff_B_WcVNyhwX7_2),.clk(gclk));
	jdff dff_B_u4pT78iO2_2(.din(w_dff_B_WcVNyhwX7_2),.dout(w_dff_B_u4pT78iO2_2),.clk(gclk));
	jdff dff_B_bjv4PFRx5_2(.din(w_dff_B_u4pT78iO2_2),.dout(w_dff_B_bjv4PFRx5_2),.clk(gclk));
	jdff dff_B_sduVcZIW5_2(.din(w_dff_B_bjv4PFRx5_2),.dout(w_dff_B_sduVcZIW5_2),.clk(gclk));
	jdff dff_B_NGW36fhR9_2(.din(w_dff_B_sduVcZIW5_2),.dout(w_dff_B_NGW36fhR9_2),.clk(gclk));
	jdff dff_B_r3j6jYjK6_2(.din(w_dff_B_NGW36fhR9_2),.dout(w_dff_B_r3j6jYjK6_2),.clk(gclk));
	jdff dff_B_bBDHLzPL3_2(.din(w_dff_B_r3j6jYjK6_2),.dout(w_dff_B_bBDHLzPL3_2),.clk(gclk));
	jdff dff_B_TofsPsMb4_2(.din(w_dff_B_bBDHLzPL3_2),.dout(w_dff_B_TofsPsMb4_2),.clk(gclk));
	jdff dff_B_udEqYqW39_2(.din(w_dff_B_TofsPsMb4_2),.dout(w_dff_B_udEqYqW39_2),.clk(gclk));
	jdff dff_B_yGZWIbEw3_2(.din(w_dff_B_udEqYqW39_2),.dout(w_dff_B_yGZWIbEw3_2),.clk(gclk));
	jdff dff_B_4jdMOdpI9_2(.din(w_dff_B_yGZWIbEw3_2),.dout(w_dff_B_4jdMOdpI9_2),.clk(gclk));
	jdff dff_B_i5nC3PJ59_2(.din(w_dff_B_4jdMOdpI9_2),.dout(w_dff_B_i5nC3PJ59_2),.clk(gclk));
	jdff dff_B_cpC5Ctxy3_2(.din(w_dff_B_i5nC3PJ59_2),.dout(w_dff_B_cpC5Ctxy3_2),.clk(gclk));
	jdff dff_B_6uAyAGD86_2(.din(w_dff_B_cpC5Ctxy3_2),.dout(w_dff_B_6uAyAGD86_2),.clk(gclk));
	jdff dff_B_Eep8acM41_2(.din(w_dff_B_6uAyAGD86_2),.dout(w_dff_B_Eep8acM41_2),.clk(gclk));
	jdff dff_B_HK7RbBR77_2(.din(w_dff_B_Eep8acM41_2),.dout(w_dff_B_HK7RbBR77_2),.clk(gclk));
	jdff dff_B_bnjkz5Xs0_2(.din(w_dff_B_HK7RbBR77_2),.dout(w_dff_B_bnjkz5Xs0_2),.clk(gclk));
	jdff dff_B_c5oPvu1p9_2(.din(w_dff_B_bnjkz5Xs0_2),.dout(w_dff_B_c5oPvu1p9_2),.clk(gclk));
	jdff dff_B_ErOjuLIh3_2(.din(w_dff_B_c5oPvu1p9_2),.dout(w_dff_B_ErOjuLIh3_2),.clk(gclk));
	jdff dff_B_H4vF8Jzv3_2(.din(w_dff_B_ErOjuLIh3_2),.dout(w_dff_B_H4vF8Jzv3_2),.clk(gclk));
	jdff dff_B_2dg9xcRF3_2(.din(w_dff_B_H4vF8Jzv3_2),.dout(w_dff_B_2dg9xcRF3_2),.clk(gclk));
	jdff dff_B_3C3MC2xr3_2(.din(w_dff_B_2dg9xcRF3_2),.dout(w_dff_B_3C3MC2xr3_2),.clk(gclk));
	jdff dff_B_xjjOOBCW3_2(.din(w_dff_B_3C3MC2xr3_2),.dout(w_dff_B_xjjOOBCW3_2),.clk(gclk));
	jdff dff_B_0HIzmumo0_2(.din(w_dff_B_xjjOOBCW3_2),.dout(w_dff_B_0HIzmumo0_2),.clk(gclk));
	jdff dff_B_YVxJX7bK8_2(.din(w_dff_B_0HIzmumo0_2),.dout(w_dff_B_YVxJX7bK8_2),.clk(gclk));
	jdff dff_B_npU4dBmU0_2(.din(w_dff_B_YVxJX7bK8_2),.dout(w_dff_B_npU4dBmU0_2),.clk(gclk));
	jdff dff_A_4srhdI5f7_0(.dout(w_n1008_0[0]),.din(w_dff_A_4srhdI5f7_0),.clk(gclk));
	jdff dff_B_7ZqNEE1X2_1(.din(n913),.dout(w_dff_B_7ZqNEE1X2_1),.clk(gclk));
	jdff dff_B_MyRF88Ho1_2(.din(n811),.dout(w_dff_B_MyRF88Ho1_2),.clk(gclk));
	jdff dff_B_vs2i8CRr4_2(.din(w_dff_B_MyRF88Ho1_2),.dout(w_dff_B_vs2i8CRr4_2),.clk(gclk));
	jdff dff_B_HxjixdtX4_2(.din(w_dff_B_vs2i8CRr4_2),.dout(w_dff_B_HxjixdtX4_2),.clk(gclk));
	jdff dff_B_2schdg8b4_2(.din(w_dff_B_HxjixdtX4_2),.dout(w_dff_B_2schdg8b4_2),.clk(gclk));
	jdff dff_B_X0AEB7865_2(.din(w_dff_B_2schdg8b4_2),.dout(w_dff_B_X0AEB7865_2),.clk(gclk));
	jdff dff_B_wSinLOER6_2(.din(w_dff_B_X0AEB7865_2),.dout(w_dff_B_wSinLOER6_2),.clk(gclk));
	jdff dff_B_ZbenMmdJ3_2(.din(w_dff_B_wSinLOER6_2),.dout(w_dff_B_ZbenMmdJ3_2),.clk(gclk));
	jdff dff_B_w4pjXUgY0_2(.din(w_dff_B_ZbenMmdJ3_2),.dout(w_dff_B_w4pjXUgY0_2),.clk(gclk));
	jdff dff_B_zixU73o69_2(.din(w_dff_B_w4pjXUgY0_2),.dout(w_dff_B_zixU73o69_2),.clk(gclk));
	jdff dff_B_Hg8CQCUM2_2(.din(w_dff_B_zixU73o69_2),.dout(w_dff_B_Hg8CQCUM2_2),.clk(gclk));
	jdff dff_B_t875ONQ45_2(.din(w_dff_B_Hg8CQCUM2_2),.dout(w_dff_B_t875ONQ45_2),.clk(gclk));
	jdff dff_B_JOVkWgXp1_2(.din(w_dff_B_t875ONQ45_2),.dout(w_dff_B_JOVkWgXp1_2),.clk(gclk));
	jdff dff_B_P0PgcrjQ4_2(.din(w_dff_B_JOVkWgXp1_2),.dout(w_dff_B_P0PgcrjQ4_2),.clk(gclk));
	jdff dff_B_oervyHLH9_2(.din(w_dff_B_P0PgcrjQ4_2),.dout(w_dff_B_oervyHLH9_2),.clk(gclk));
	jdff dff_B_JbZSDcwQ1_2(.din(w_dff_B_oervyHLH9_2),.dout(w_dff_B_JbZSDcwQ1_2),.clk(gclk));
	jdff dff_B_yTmfgBJe2_2(.din(w_dff_B_JbZSDcwQ1_2),.dout(w_dff_B_yTmfgBJe2_2),.clk(gclk));
	jdff dff_B_20aD1xrL6_2(.din(w_dff_B_yTmfgBJe2_2),.dout(w_dff_B_20aD1xrL6_2),.clk(gclk));
	jdff dff_B_Zv2aVvHy0_2(.din(w_dff_B_20aD1xrL6_2),.dout(w_dff_B_Zv2aVvHy0_2),.clk(gclk));
	jdff dff_B_2RQgefhu4_2(.din(w_dff_B_Zv2aVvHy0_2),.dout(w_dff_B_2RQgefhu4_2),.clk(gclk));
	jdff dff_B_AOMSN1Mt7_2(.din(w_dff_B_2RQgefhu4_2),.dout(w_dff_B_AOMSN1Mt7_2),.clk(gclk));
	jdff dff_B_Oj94We1D8_2(.din(w_dff_B_AOMSN1Mt7_2),.dout(w_dff_B_Oj94We1D8_2),.clk(gclk));
	jdff dff_B_lA1NGeNw4_2(.din(w_dff_B_Oj94We1D8_2),.dout(w_dff_B_lA1NGeNw4_2),.clk(gclk));
	jdff dff_B_DL1JyQv69_2(.din(w_dff_B_lA1NGeNw4_2),.dout(w_dff_B_DL1JyQv69_2),.clk(gclk));
	jdff dff_B_YpF83VGD4_2(.din(w_dff_B_DL1JyQv69_2),.dout(w_dff_B_YpF83VGD4_2),.clk(gclk));
	jdff dff_B_sobBcY7u5_2(.din(w_dff_B_YpF83VGD4_2),.dout(w_dff_B_sobBcY7u5_2),.clk(gclk));
	jdff dff_B_H928jWCT5_2(.din(w_dff_B_sobBcY7u5_2),.dout(w_dff_B_H928jWCT5_2),.clk(gclk));
	jdff dff_B_Pdn3zpCf7_2(.din(w_dff_B_H928jWCT5_2),.dout(w_dff_B_Pdn3zpCf7_2),.clk(gclk));
	jdff dff_B_EuvBYWQp7_2(.din(w_dff_B_Pdn3zpCf7_2),.dout(w_dff_B_EuvBYWQp7_2),.clk(gclk));
	jdff dff_B_88g5pI1W8_2(.din(w_dff_B_EuvBYWQp7_2),.dout(w_dff_B_88g5pI1W8_2),.clk(gclk));
	jdff dff_B_usMhhRpj6_2(.din(w_dff_B_88g5pI1W8_2),.dout(w_dff_B_usMhhRpj6_2),.clk(gclk));
	jdff dff_B_sKOj6k0h7_2(.din(w_dff_B_usMhhRpj6_2),.dout(w_dff_B_sKOj6k0h7_2),.clk(gclk));
	jdff dff_B_Nf4BGIkL3_2(.din(w_dff_B_sKOj6k0h7_2),.dout(w_dff_B_Nf4BGIkL3_2),.clk(gclk));
	jdff dff_B_U8VFAW3G6_2(.din(w_dff_B_Nf4BGIkL3_2),.dout(w_dff_B_U8VFAW3G6_2),.clk(gclk));
	jdff dff_B_6eUkt3ob1_2(.din(w_dff_B_U8VFAW3G6_2),.dout(w_dff_B_6eUkt3ob1_2),.clk(gclk));
	jdff dff_B_F96ZW9ZA5_2(.din(w_dff_B_6eUkt3ob1_2),.dout(w_dff_B_F96ZW9ZA5_2),.clk(gclk));
	jdff dff_B_Yev0Ya1m6_2(.din(w_dff_B_F96ZW9ZA5_2),.dout(w_dff_B_Yev0Ya1m6_2),.clk(gclk));
	jdff dff_B_ofK5VT0q6_2(.din(w_dff_B_Yev0Ya1m6_2),.dout(w_dff_B_ofK5VT0q6_2),.clk(gclk));
	jdff dff_B_BQyzyyjB3_2(.din(w_dff_B_ofK5VT0q6_2),.dout(w_dff_B_BQyzyyjB3_2),.clk(gclk));
	jdff dff_B_nEkoHJJ30_2(.din(w_dff_B_BQyzyyjB3_2),.dout(w_dff_B_nEkoHJJ30_2),.clk(gclk));
	jdff dff_B_GjiEG68z4_2(.din(w_dff_B_nEkoHJJ30_2),.dout(w_dff_B_GjiEG68z4_2),.clk(gclk));
	jdff dff_A_pk5fm7722_1(.dout(w_n902_0[1]),.din(w_dff_A_pk5fm7722_1),.clk(gclk));
	jdff dff_B_mH3YQC8G2_1(.din(n817),.dout(w_dff_B_mH3YQC8G2_1),.clk(gclk));
	jdff dff_B_mi78tRPC4_1(.din(w_dff_B_mH3YQC8G2_1),.dout(w_dff_B_mi78tRPC4_1),.clk(gclk));
	jdff dff_B_CuSZhulK4_1(.din(w_dff_B_mi78tRPC4_1),.dout(w_dff_B_CuSZhulK4_1),.clk(gclk));
	jdff dff_B_POOwfaAm1_1(.din(w_dff_B_CuSZhulK4_1),.dout(w_dff_B_POOwfaAm1_1),.clk(gclk));
	jdff dff_B_bUBtQcxz5_1(.din(w_dff_B_POOwfaAm1_1),.dout(w_dff_B_bUBtQcxz5_1),.clk(gclk));
	jdff dff_B_RaTCpOwE7_1(.din(w_dff_B_bUBtQcxz5_1),.dout(w_dff_B_RaTCpOwE7_1),.clk(gclk));
	jdff dff_B_79dFNKNP5_1(.din(w_dff_B_RaTCpOwE7_1),.dout(w_dff_B_79dFNKNP5_1),.clk(gclk));
	jdff dff_B_fmMxAAbW0_1(.din(w_dff_B_79dFNKNP5_1),.dout(w_dff_B_fmMxAAbW0_1),.clk(gclk));
	jdff dff_B_OekLfmFc3_1(.din(w_dff_B_fmMxAAbW0_1),.dout(w_dff_B_OekLfmFc3_1),.clk(gclk));
	jdff dff_B_6Zr66Qik3_1(.din(w_dff_B_OekLfmFc3_1),.dout(w_dff_B_6Zr66Qik3_1),.clk(gclk));
	jdff dff_B_9Avhm6r94_1(.din(w_dff_B_6Zr66Qik3_1),.dout(w_dff_B_9Avhm6r94_1),.clk(gclk));
	jdff dff_B_zxje7ffB9_1(.din(w_dff_B_9Avhm6r94_1),.dout(w_dff_B_zxje7ffB9_1),.clk(gclk));
	jdff dff_B_BBDmSs0x4_1(.din(w_dff_B_zxje7ffB9_1),.dout(w_dff_B_BBDmSs0x4_1),.clk(gclk));
	jdff dff_B_gA4B9JWh8_1(.din(w_dff_B_BBDmSs0x4_1),.dout(w_dff_B_gA4B9JWh8_1),.clk(gclk));
	jdff dff_B_uXHsKQAB2_1(.din(w_dff_B_gA4B9JWh8_1),.dout(w_dff_B_uXHsKQAB2_1),.clk(gclk));
	jdff dff_B_g3lXLIwq1_1(.din(w_dff_B_uXHsKQAB2_1),.dout(w_dff_B_g3lXLIwq1_1),.clk(gclk));
	jdff dff_B_lCZmjHv13_1(.din(w_dff_B_g3lXLIwq1_1),.dout(w_dff_B_lCZmjHv13_1),.clk(gclk));
	jdff dff_B_82cERNsd2_1(.din(w_dff_B_lCZmjHv13_1),.dout(w_dff_B_82cERNsd2_1),.clk(gclk));
	jdff dff_B_r8jcfOAp4_1(.din(w_dff_B_82cERNsd2_1),.dout(w_dff_B_r8jcfOAp4_1),.clk(gclk));
	jdff dff_B_5dn8vxyq0_1(.din(w_dff_B_r8jcfOAp4_1),.dout(w_dff_B_5dn8vxyq0_1),.clk(gclk));
	jdff dff_B_eQCeMJtD9_1(.din(w_dff_B_5dn8vxyq0_1),.dout(w_dff_B_eQCeMJtD9_1),.clk(gclk));
	jdff dff_B_VBj5hVN94_1(.din(w_dff_B_eQCeMJtD9_1),.dout(w_dff_B_VBj5hVN94_1),.clk(gclk));
	jdff dff_B_yx5b9oMt1_1(.din(w_dff_B_VBj5hVN94_1),.dout(w_dff_B_yx5b9oMt1_1),.clk(gclk));
	jdff dff_B_TP95Tceu1_1(.din(w_dff_B_yx5b9oMt1_1),.dout(w_dff_B_TP95Tceu1_1),.clk(gclk));
	jdff dff_B_NTd7QoBg8_1(.din(w_dff_B_TP95Tceu1_1),.dout(w_dff_B_NTd7QoBg8_1),.clk(gclk));
	jdff dff_B_JpcRq0sr7_1(.din(w_dff_B_NTd7QoBg8_1),.dout(w_dff_B_JpcRq0sr7_1),.clk(gclk));
	jdff dff_B_8MWQTBhw6_1(.din(w_dff_B_JpcRq0sr7_1),.dout(w_dff_B_8MWQTBhw6_1),.clk(gclk));
	jdff dff_B_ukRNl2yb2_1(.din(w_dff_B_8MWQTBhw6_1),.dout(w_dff_B_ukRNl2yb2_1),.clk(gclk));
	jdff dff_B_dXQkpcAo9_1(.din(w_dff_B_ukRNl2yb2_1),.dout(w_dff_B_dXQkpcAo9_1),.clk(gclk));
	jdff dff_B_fP1syjHV2_1(.din(w_dff_B_dXQkpcAo9_1),.dout(w_dff_B_fP1syjHV2_1),.clk(gclk));
	jdff dff_B_edtvXeBF9_1(.din(w_dff_B_fP1syjHV2_1),.dout(w_dff_B_edtvXeBF9_1),.clk(gclk));
	jdff dff_B_ZRecMDAO6_1(.din(w_dff_B_edtvXeBF9_1),.dout(w_dff_B_ZRecMDAO6_1),.clk(gclk));
	jdff dff_B_wazNxPDQ7_1(.din(w_dff_B_ZRecMDAO6_1),.dout(w_dff_B_wazNxPDQ7_1),.clk(gclk));
	jdff dff_B_4KHvnmWF6_1(.din(w_dff_B_wazNxPDQ7_1),.dout(w_dff_B_4KHvnmWF6_1),.clk(gclk));
	jdff dff_B_ubCutBrC6_1(.din(w_dff_B_4KHvnmWF6_1),.dout(w_dff_B_ubCutBrC6_1),.clk(gclk));
	jdff dff_B_IauIUggA0_1(.din(w_dff_B_ubCutBrC6_1),.dout(w_dff_B_IauIUggA0_1),.clk(gclk));
	jdff dff_B_e90BrRBC1_1(.din(n812),.dout(w_dff_B_e90BrRBC1_1),.clk(gclk));
	jdff dff_A_4cCVeIPs0_0(.dout(w_n712_0[0]),.din(w_dff_A_4cCVeIPs0_0),.clk(gclk));
	jdff dff_A_Puj7Y3jZ5_0(.dout(w_dff_A_4cCVeIPs0_0),.din(w_dff_A_Puj7Y3jZ5_0),.clk(gclk));
	jdff dff_A_XM7PygpP9_0(.dout(w_dff_A_Puj7Y3jZ5_0),.din(w_dff_A_XM7PygpP9_0),.clk(gclk));
	jdff dff_A_7flPWa5f8_0(.dout(w_dff_A_XM7PygpP9_0),.din(w_dff_A_7flPWa5f8_0),.clk(gclk));
	jdff dff_A_ktjG7CB24_0(.dout(w_dff_A_7flPWa5f8_0),.din(w_dff_A_ktjG7CB24_0),.clk(gclk));
	jdff dff_A_F4tBUn2w1_0(.dout(w_dff_A_ktjG7CB24_0),.din(w_dff_A_F4tBUn2w1_0),.clk(gclk));
	jdff dff_A_GVQjSI4K8_0(.dout(w_dff_A_F4tBUn2w1_0),.din(w_dff_A_GVQjSI4K8_0),.clk(gclk));
	jdff dff_A_9B2KPkSK3_0(.dout(w_dff_A_GVQjSI4K8_0),.din(w_dff_A_9B2KPkSK3_0),.clk(gclk));
	jdff dff_A_99fWzCkJ8_0(.dout(w_dff_A_9B2KPkSK3_0),.din(w_dff_A_99fWzCkJ8_0),.clk(gclk));
	jdff dff_A_JsBJ9IlF9_0(.dout(w_dff_A_99fWzCkJ8_0),.din(w_dff_A_JsBJ9IlF9_0),.clk(gclk));
	jdff dff_A_u9Y17Nz70_0(.dout(w_dff_A_JsBJ9IlF9_0),.din(w_dff_A_u9Y17Nz70_0),.clk(gclk));
	jdff dff_A_zaZuvExN7_0(.dout(w_dff_A_u9Y17Nz70_0),.din(w_dff_A_zaZuvExN7_0),.clk(gclk));
	jdff dff_A_vR9gCxSH4_0(.dout(w_dff_A_zaZuvExN7_0),.din(w_dff_A_vR9gCxSH4_0),.clk(gclk));
	jdff dff_A_o4YK45B50_0(.dout(w_dff_A_vR9gCxSH4_0),.din(w_dff_A_o4YK45B50_0),.clk(gclk));
	jdff dff_A_vC464gJA6_0(.dout(w_dff_A_o4YK45B50_0),.din(w_dff_A_vC464gJA6_0),.clk(gclk));
	jdff dff_A_SzwDyVug4_0(.dout(w_dff_A_vC464gJA6_0),.din(w_dff_A_SzwDyVug4_0),.clk(gclk));
	jdff dff_A_nsS9aEr48_0(.dout(w_dff_A_SzwDyVug4_0),.din(w_dff_A_nsS9aEr48_0),.clk(gclk));
	jdff dff_A_Zt5QNNE91_0(.dout(w_dff_A_nsS9aEr48_0),.din(w_dff_A_Zt5QNNE91_0),.clk(gclk));
	jdff dff_A_qhJqJTnu3_0(.dout(w_dff_A_Zt5QNNE91_0),.din(w_dff_A_qhJqJTnu3_0),.clk(gclk));
	jdff dff_A_m0dD5oNw2_0(.dout(w_dff_A_qhJqJTnu3_0),.din(w_dff_A_m0dD5oNw2_0),.clk(gclk));
	jdff dff_A_OUkrUA4s7_0(.dout(w_dff_A_m0dD5oNw2_0),.din(w_dff_A_OUkrUA4s7_0),.clk(gclk));
	jdff dff_A_7hkTAzJD5_0(.dout(w_dff_A_OUkrUA4s7_0),.din(w_dff_A_7hkTAzJD5_0),.clk(gclk));
	jdff dff_A_NDMZ93ru7_0(.dout(w_dff_A_7hkTAzJD5_0),.din(w_dff_A_NDMZ93ru7_0),.clk(gclk));
	jdff dff_A_fnpmKFz18_0(.dout(w_dff_A_NDMZ93ru7_0),.din(w_dff_A_fnpmKFz18_0),.clk(gclk));
	jdff dff_A_dXcqFxTP9_0(.dout(w_dff_A_fnpmKFz18_0),.din(w_dff_A_dXcqFxTP9_0),.clk(gclk));
	jdff dff_A_OFTxbFi85_0(.dout(w_dff_A_dXcqFxTP9_0),.din(w_dff_A_OFTxbFi85_0),.clk(gclk));
	jdff dff_A_rFHXN8Fe6_0(.dout(w_dff_A_OFTxbFi85_0),.din(w_dff_A_rFHXN8Fe6_0),.clk(gclk));
	jdff dff_A_y4KpsBnx8_0(.dout(w_dff_A_rFHXN8Fe6_0),.din(w_dff_A_y4KpsBnx8_0),.clk(gclk));
	jdff dff_A_ex8Vjarn0_0(.dout(w_dff_A_y4KpsBnx8_0),.din(w_dff_A_ex8Vjarn0_0),.clk(gclk));
	jdff dff_A_m8PoQSv38_0(.dout(w_dff_A_ex8Vjarn0_0),.din(w_dff_A_m8PoQSv38_0),.clk(gclk));
	jdff dff_A_jp9BR9eU5_0(.dout(w_dff_A_m8PoQSv38_0),.din(w_dff_A_jp9BR9eU5_0),.clk(gclk));
	jdff dff_A_Y5rzik6T1_0(.dout(w_dff_A_jp9BR9eU5_0),.din(w_dff_A_Y5rzik6T1_0),.clk(gclk));
	jdff dff_A_EZ16Ww6f0_0(.dout(w_dff_A_Y5rzik6T1_0),.din(w_dff_A_EZ16Ww6f0_0),.clk(gclk));
	jdff dff_A_UThHCoHP4_0(.dout(w_dff_A_EZ16Ww6f0_0),.din(w_dff_A_UThHCoHP4_0),.clk(gclk));
	jdff dff_A_ICtdikRJ5_0(.dout(w_dff_A_UThHCoHP4_0),.din(w_dff_A_ICtdikRJ5_0),.clk(gclk));
	jdff dff_A_SfWTCEAE1_0(.dout(w_dff_A_ICtdikRJ5_0),.din(w_dff_A_SfWTCEAE1_0),.clk(gclk));
	jdff dff_A_MZQj5o8y5_0(.dout(w_dff_A_SfWTCEAE1_0),.din(w_dff_A_MZQj5o8y5_0),.clk(gclk));
	jdff dff_A_ZPHxKH3L7_0(.dout(w_n799_0[0]),.din(w_dff_A_ZPHxKH3L7_0),.clk(gclk));
	jdff dff_B_TcMWfGUl2_1(.din(n714),.dout(w_dff_B_TcMWfGUl2_1),.clk(gclk));
	jdff dff_A_yep8Mkb95_0(.dout(w_n620_0[0]),.din(w_dff_A_yep8Mkb95_0),.clk(gclk));
	jdff dff_A_Ml3cU1p46_0(.dout(w_dff_A_yep8Mkb95_0),.din(w_dff_A_Ml3cU1p46_0),.clk(gclk));
	jdff dff_A_cUhWZDR51_0(.dout(w_dff_A_Ml3cU1p46_0),.din(w_dff_A_cUhWZDR51_0),.clk(gclk));
	jdff dff_A_VsJ9vFWg0_0(.dout(w_dff_A_cUhWZDR51_0),.din(w_dff_A_VsJ9vFWg0_0),.clk(gclk));
	jdff dff_A_kdsM8Nuk2_0(.dout(w_dff_A_VsJ9vFWg0_0),.din(w_dff_A_kdsM8Nuk2_0),.clk(gclk));
	jdff dff_A_m5FNblAF6_0(.dout(w_dff_A_kdsM8Nuk2_0),.din(w_dff_A_m5FNblAF6_0),.clk(gclk));
	jdff dff_A_8o5GQI4n3_0(.dout(w_dff_A_m5FNblAF6_0),.din(w_dff_A_8o5GQI4n3_0),.clk(gclk));
	jdff dff_A_vZQmsyke1_0(.dout(w_dff_A_8o5GQI4n3_0),.din(w_dff_A_vZQmsyke1_0),.clk(gclk));
	jdff dff_A_xqneDfm06_0(.dout(w_dff_A_vZQmsyke1_0),.din(w_dff_A_xqneDfm06_0),.clk(gclk));
	jdff dff_A_zqb877gu3_0(.dout(w_dff_A_xqneDfm06_0),.din(w_dff_A_zqb877gu3_0),.clk(gclk));
	jdff dff_A_yZD8demx9_0(.dout(w_dff_A_zqb877gu3_0),.din(w_dff_A_yZD8demx9_0),.clk(gclk));
	jdff dff_A_hfNXxVHy4_0(.dout(w_dff_A_yZD8demx9_0),.din(w_dff_A_hfNXxVHy4_0),.clk(gclk));
	jdff dff_A_OcUc42Uf2_0(.dout(w_dff_A_hfNXxVHy4_0),.din(w_dff_A_OcUc42Uf2_0),.clk(gclk));
	jdff dff_A_nE2Pm5Zp5_0(.dout(w_dff_A_OcUc42Uf2_0),.din(w_dff_A_nE2Pm5Zp5_0),.clk(gclk));
	jdff dff_A_b4DvnkBd7_0(.dout(w_dff_A_nE2Pm5Zp5_0),.din(w_dff_A_b4DvnkBd7_0),.clk(gclk));
	jdff dff_A_Gq0Zcrfz6_0(.dout(w_dff_A_b4DvnkBd7_0),.din(w_dff_A_Gq0Zcrfz6_0),.clk(gclk));
	jdff dff_A_TdTx8Vid6_0(.dout(w_dff_A_Gq0Zcrfz6_0),.din(w_dff_A_TdTx8Vid6_0),.clk(gclk));
	jdff dff_A_by2xzjeB0_0(.dout(w_dff_A_TdTx8Vid6_0),.din(w_dff_A_by2xzjeB0_0),.clk(gclk));
	jdff dff_A_6ePQ0IMP4_0(.dout(w_dff_A_by2xzjeB0_0),.din(w_dff_A_6ePQ0IMP4_0),.clk(gclk));
	jdff dff_A_TezrQHhD4_0(.dout(w_dff_A_6ePQ0IMP4_0),.din(w_dff_A_TezrQHhD4_0),.clk(gclk));
	jdff dff_A_YYTYTgYW8_0(.dout(w_dff_A_TezrQHhD4_0),.din(w_dff_A_YYTYTgYW8_0),.clk(gclk));
	jdff dff_A_hlOgDtrn2_0(.dout(w_dff_A_YYTYTgYW8_0),.din(w_dff_A_hlOgDtrn2_0),.clk(gclk));
	jdff dff_A_RgcRg5WZ4_0(.dout(w_dff_A_hlOgDtrn2_0),.din(w_dff_A_RgcRg5WZ4_0),.clk(gclk));
	jdff dff_A_srhpZvbs1_0(.dout(w_dff_A_RgcRg5WZ4_0),.din(w_dff_A_srhpZvbs1_0),.clk(gclk));
	jdff dff_A_8pZMFplZ5_0(.dout(w_dff_A_srhpZvbs1_0),.din(w_dff_A_8pZMFplZ5_0),.clk(gclk));
	jdff dff_A_dVLxC8g57_0(.dout(w_dff_A_8pZMFplZ5_0),.din(w_dff_A_dVLxC8g57_0),.clk(gclk));
	jdff dff_A_UFUxdAPV2_0(.dout(w_dff_A_dVLxC8g57_0),.din(w_dff_A_UFUxdAPV2_0),.clk(gclk));
	jdff dff_A_09L0zUaT4_0(.dout(w_dff_A_UFUxdAPV2_0),.din(w_dff_A_09L0zUaT4_0),.clk(gclk));
	jdff dff_A_gDRNrXgf6_0(.dout(w_dff_A_09L0zUaT4_0),.din(w_dff_A_gDRNrXgf6_0),.clk(gclk));
	jdff dff_A_18hIphsv7_0(.dout(w_dff_A_gDRNrXgf6_0),.din(w_dff_A_18hIphsv7_0),.clk(gclk));
	jdff dff_A_XCvrLZwF6_0(.dout(w_dff_A_18hIphsv7_0),.din(w_dff_A_XCvrLZwF6_0),.clk(gclk));
	jdff dff_A_jYUIfQ6Y2_0(.dout(w_dff_A_XCvrLZwF6_0),.din(w_dff_A_jYUIfQ6Y2_0),.clk(gclk));
	jdff dff_A_SmcgCxUj2_0(.dout(w_dff_A_jYUIfQ6Y2_0),.din(w_dff_A_SmcgCxUj2_0),.clk(gclk));
	jdff dff_A_KIQ1Xrxm6_0(.dout(w_dff_A_SmcgCxUj2_0),.din(w_dff_A_KIQ1Xrxm6_0),.clk(gclk));
	jdff dff_A_D4J8BljM6_0(.dout(w_n700_0[0]),.din(w_dff_A_D4J8BljM6_0),.clk(gclk));
	jdff dff_B_3ol2YPqu2_1(.din(n622),.dout(w_dff_B_3ol2YPqu2_1),.clk(gclk));
	jdff dff_A_i1JM5dwV8_0(.dout(w_n535_0[0]),.din(w_dff_A_i1JM5dwV8_0),.clk(gclk));
	jdff dff_A_WOZggPKq5_0(.dout(w_dff_A_i1JM5dwV8_0),.din(w_dff_A_WOZggPKq5_0),.clk(gclk));
	jdff dff_A_6GtOBhRn8_0(.dout(w_dff_A_WOZggPKq5_0),.din(w_dff_A_6GtOBhRn8_0),.clk(gclk));
	jdff dff_A_noy1VxbO8_0(.dout(w_dff_A_6GtOBhRn8_0),.din(w_dff_A_noy1VxbO8_0),.clk(gclk));
	jdff dff_A_qsasqbgO9_0(.dout(w_dff_A_noy1VxbO8_0),.din(w_dff_A_qsasqbgO9_0),.clk(gclk));
	jdff dff_A_5tDBfrqP1_0(.dout(w_dff_A_qsasqbgO9_0),.din(w_dff_A_5tDBfrqP1_0),.clk(gclk));
	jdff dff_A_q0O0cgm53_0(.dout(w_dff_A_5tDBfrqP1_0),.din(w_dff_A_q0O0cgm53_0),.clk(gclk));
	jdff dff_A_Va48axrL4_0(.dout(w_dff_A_q0O0cgm53_0),.din(w_dff_A_Va48axrL4_0),.clk(gclk));
	jdff dff_A_qtWnJQZR8_0(.dout(w_dff_A_Va48axrL4_0),.din(w_dff_A_qtWnJQZR8_0),.clk(gclk));
	jdff dff_A_WTKJSQpe7_0(.dout(w_dff_A_qtWnJQZR8_0),.din(w_dff_A_WTKJSQpe7_0),.clk(gclk));
	jdff dff_A_1Wb5c5Hi8_0(.dout(w_dff_A_WTKJSQpe7_0),.din(w_dff_A_1Wb5c5Hi8_0),.clk(gclk));
	jdff dff_A_G061ckVS1_0(.dout(w_dff_A_1Wb5c5Hi8_0),.din(w_dff_A_G061ckVS1_0),.clk(gclk));
	jdff dff_A_hqnuUQHr9_0(.dout(w_dff_A_G061ckVS1_0),.din(w_dff_A_hqnuUQHr9_0),.clk(gclk));
	jdff dff_A_Tt1tlz4D8_0(.dout(w_dff_A_hqnuUQHr9_0),.din(w_dff_A_Tt1tlz4D8_0),.clk(gclk));
	jdff dff_A_shqwgRBP3_0(.dout(w_dff_A_Tt1tlz4D8_0),.din(w_dff_A_shqwgRBP3_0),.clk(gclk));
	jdff dff_A_LboxpIG64_0(.dout(w_dff_A_shqwgRBP3_0),.din(w_dff_A_LboxpIG64_0),.clk(gclk));
	jdff dff_A_2Ks4Js8K2_0(.dout(w_dff_A_LboxpIG64_0),.din(w_dff_A_2Ks4Js8K2_0),.clk(gclk));
	jdff dff_A_TArPpHmr3_0(.dout(w_dff_A_2Ks4Js8K2_0),.din(w_dff_A_TArPpHmr3_0),.clk(gclk));
	jdff dff_A_Jqtgd0Un3_0(.dout(w_dff_A_TArPpHmr3_0),.din(w_dff_A_Jqtgd0Un3_0),.clk(gclk));
	jdff dff_A_XTw8XSQ82_0(.dout(w_dff_A_Jqtgd0Un3_0),.din(w_dff_A_XTw8XSQ82_0),.clk(gclk));
	jdff dff_A_q59joT0v6_0(.dout(w_dff_A_XTw8XSQ82_0),.din(w_dff_A_q59joT0v6_0),.clk(gclk));
	jdff dff_A_H0QPgv0Z4_0(.dout(w_dff_A_q59joT0v6_0),.din(w_dff_A_H0QPgv0Z4_0),.clk(gclk));
	jdff dff_A_ggsxK3ad0_0(.dout(w_dff_A_H0QPgv0Z4_0),.din(w_dff_A_ggsxK3ad0_0),.clk(gclk));
	jdff dff_A_JvHzqgkK6_0(.dout(w_dff_A_ggsxK3ad0_0),.din(w_dff_A_JvHzqgkK6_0),.clk(gclk));
	jdff dff_A_3hDHtTTp4_0(.dout(w_dff_A_JvHzqgkK6_0),.din(w_dff_A_3hDHtTTp4_0),.clk(gclk));
	jdff dff_A_Vh4Xs31y1_0(.dout(w_dff_A_3hDHtTTp4_0),.din(w_dff_A_Vh4Xs31y1_0),.clk(gclk));
	jdff dff_A_s5ABN5T91_0(.dout(w_dff_A_Vh4Xs31y1_0),.din(w_dff_A_s5ABN5T91_0),.clk(gclk));
	jdff dff_A_I83dDIWl2_0(.dout(w_dff_A_s5ABN5T91_0),.din(w_dff_A_I83dDIWl2_0),.clk(gclk));
	jdff dff_A_yBAJ2YQw2_0(.dout(w_dff_A_I83dDIWl2_0),.din(w_dff_A_yBAJ2YQw2_0),.clk(gclk));
	jdff dff_A_BQ4RT4cZ8_0(.dout(w_dff_A_yBAJ2YQw2_0),.din(w_dff_A_BQ4RT4cZ8_0),.clk(gclk));
	jdff dff_A_QnXpZbch3_0(.dout(w_dff_A_BQ4RT4cZ8_0),.din(w_dff_A_QnXpZbch3_0),.clk(gclk));
	jdff dff_A_YThLcJGt7_0(.dout(w_n608_0[0]),.din(w_dff_A_YThLcJGt7_0),.clk(gclk));
	jdff dff_B_Wx8gVA3f4_1(.din(n537),.dout(w_dff_B_Wx8gVA3f4_1),.clk(gclk));
	jdff dff_A_Dp6pYkgg5_0(.dout(w_n457_0[0]),.din(w_dff_A_Dp6pYkgg5_0),.clk(gclk));
	jdff dff_A_kLiuxRIq5_0(.dout(w_dff_A_Dp6pYkgg5_0),.din(w_dff_A_kLiuxRIq5_0),.clk(gclk));
	jdff dff_A_k9SGnOS40_0(.dout(w_dff_A_kLiuxRIq5_0),.din(w_dff_A_k9SGnOS40_0),.clk(gclk));
	jdff dff_A_UxINHyAF6_0(.dout(w_dff_A_k9SGnOS40_0),.din(w_dff_A_UxINHyAF6_0),.clk(gclk));
	jdff dff_A_yX94VMgY2_0(.dout(w_dff_A_UxINHyAF6_0),.din(w_dff_A_yX94VMgY2_0),.clk(gclk));
	jdff dff_A_LZASZojU4_0(.dout(w_dff_A_yX94VMgY2_0),.din(w_dff_A_LZASZojU4_0),.clk(gclk));
	jdff dff_A_WUL0oOaN2_0(.dout(w_dff_A_LZASZojU4_0),.din(w_dff_A_WUL0oOaN2_0),.clk(gclk));
	jdff dff_A_OQt0ht2d9_0(.dout(w_dff_A_WUL0oOaN2_0),.din(w_dff_A_OQt0ht2d9_0),.clk(gclk));
	jdff dff_A_Qn2YoWTQ8_0(.dout(w_dff_A_OQt0ht2d9_0),.din(w_dff_A_Qn2YoWTQ8_0),.clk(gclk));
	jdff dff_A_wQsDb4ik3_0(.dout(w_dff_A_Qn2YoWTQ8_0),.din(w_dff_A_wQsDb4ik3_0),.clk(gclk));
	jdff dff_A_qorG1gqc8_0(.dout(w_dff_A_wQsDb4ik3_0),.din(w_dff_A_qorG1gqc8_0),.clk(gclk));
	jdff dff_A_RjXcQ55b2_0(.dout(w_dff_A_qorG1gqc8_0),.din(w_dff_A_RjXcQ55b2_0),.clk(gclk));
	jdff dff_A_54zR3vse1_0(.dout(w_dff_A_RjXcQ55b2_0),.din(w_dff_A_54zR3vse1_0),.clk(gclk));
	jdff dff_A_AkOGVlTY6_0(.dout(w_dff_A_54zR3vse1_0),.din(w_dff_A_AkOGVlTY6_0),.clk(gclk));
	jdff dff_A_sHm8lLFr8_0(.dout(w_dff_A_AkOGVlTY6_0),.din(w_dff_A_sHm8lLFr8_0),.clk(gclk));
	jdff dff_A_6zqJZpsy7_0(.dout(w_dff_A_sHm8lLFr8_0),.din(w_dff_A_6zqJZpsy7_0),.clk(gclk));
	jdff dff_A_86V7Tos08_0(.dout(w_dff_A_6zqJZpsy7_0),.din(w_dff_A_86V7Tos08_0),.clk(gclk));
	jdff dff_A_9jgUymra0_0(.dout(w_dff_A_86V7Tos08_0),.din(w_dff_A_9jgUymra0_0),.clk(gclk));
	jdff dff_A_43oKsjpy8_0(.dout(w_dff_A_9jgUymra0_0),.din(w_dff_A_43oKsjpy8_0),.clk(gclk));
	jdff dff_A_oOjK5N8O8_0(.dout(w_dff_A_43oKsjpy8_0),.din(w_dff_A_oOjK5N8O8_0),.clk(gclk));
	jdff dff_A_Q1KcbHFn1_0(.dout(w_dff_A_oOjK5N8O8_0),.din(w_dff_A_Q1KcbHFn1_0),.clk(gclk));
	jdff dff_A_kibVlbmf0_0(.dout(w_dff_A_Q1KcbHFn1_0),.din(w_dff_A_kibVlbmf0_0),.clk(gclk));
	jdff dff_A_6KfgduoD1_0(.dout(w_dff_A_kibVlbmf0_0),.din(w_dff_A_6KfgduoD1_0),.clk(gclk));
	jdff dff_A_uvKssEkd3_0(.dout(w_dff_A_6KfgduoD1_0),.din(w_dff_A_uvKssEkd3_0),.clk(gclk));
	jdff dff_A_6hOg0Fg01_0(.dout(w_dff_A_uvKssEkd3_0),.din(w_dff_A_6hOg0Fg01_0),.clk(gclk));
	jdff dff_A_TR5dnRrm7_0(.dout(w_dff_A_6hOg0Fg01_0),.din(w_dff_A_TR5dnRrm7_0),.clk(gclk));
	jdff dff_A_xzNnXzgm5_0(.dout(w_dff_A_TR5dnRrm7_0),.din(w_dff_A_xzNnXzgm5_0),.clk(gclk));
	jdff dff_A_yRb039tD0_0(.dout(w_dff_A_xzNnXzgm5_0),.din(w_dff_A_yRb039tD0_0),.clk(gclk));
	jdff dff_A_TVcECwO33_0(.dout(w_n523_0[0]),.din(w_dff_A_TVcECwO33_0),.clk(gclk));
	jdff dff_B_4nstmJjP9_1(.din(n459),.dout(w_dff_B_4nstmJjP9_1),.clk(gclk));
	jdff dff_A_GMKIGBu49_0(.dout(w_n386_0[0]),.din(w_dff_A_GMKIGBu49_0),.clk(gclk));
	jdff dff_A_BfaZkGg15_0(.dout(w_dff_A_GMKIGBu49_0),.din(w_dff_A_BfaZkGg15_0),.clk(gclk));
	jdff dff_A_rVzu2cTz0_0(.dout(w_dff_A_BfaZkGg15_0),.din(w_dff_A_rVzu2cTz0_0),.clk(gclk));
	jdff dff_A_rIusyq2v3_0(.dout(w_dff_A_rVzu2cTz0_0),.din(w_dff_A_rIusyq2v3_0),.clk(gclk));
	jdff dff_A_JXQFsXgi1_0(.dout(w_dff_A_rIusyq2v3_0),.din(w_dff_A_JXQFsXgi1_0),.clk(gclk));
	jdff dff_A_0I8RhK9w5_0(.dout(w_dff_A_JXQFsXgi1_0),.din(w_dff_A_0I8RhK9w5_0),.clk(gclk));
	jdff dff_A_OkX2pUTe8_0(.dout(w_dff_A_0I8RhK9w5_0),.din(w_dff_A_OkX2pUTe8_0),.clk(gclk));
	jdff dff_A_26MB3cam6_0(.dout(w_dff_A_OkX2pUTe8_0),.din(w_dff_A_26MB3cam6_0),.clk(gclk));
	jdff dff_A_jkixgHNI8_0(.dout(w_dff_A_26MB3cam6_0),.din(w_dff_A_jkixgHNI8_0),.clk(gclk));
	jdff dff_A_dPIAWrUa4_0(.dout(w_dff_A_jkixgHNI8_0),.din(w_dff_A_dPIAWrUa4_0),.clk(gclk));
	jdff dff_A_nJvHBlKN9_0(.dout(w_dff_A_dPIAWrUa4_0),.din(w_dff_A_nJvHBlKN9_0),.clk(gclk));
	jdff dff_A_HkOiRcYj8_0(.dout(w_dff_A_nJvHBlKN9_0),.din(w_dff_A_HkOiRcYj8_0),.clk(gclk));
	jdff dff_A_TvJWAPnU4_0(.dout(w_dff_A_HkOiRcYj8_0),.din(w_dff_A_TvJWAPnU4_0),.clk(gclk));
	jdff dff_A_p2u4AGtI7_0(.dout(w_dff_A_TvJWAPnU4_0),.din(w_dff_A_p2u4AGtI7_0),.clk(gclk));
	jdff dff_A_qIVvVm9z7_0(.dout(w_dff_A_p2u4AGtI7_0),.din(w_dff_A_qIVvVm9z7_0),.clk(gclk));
	jdff dff_A_tKAoNEmu9_0(.dout(w_dff_A_qIVvVm9z7_0),.din(w_dff_A_tKAoNEmu9_0),.clk(gclk));
	jdff dff_A_qpmAS6uv8_0(.dout(w_dff_A_tKAoNEmu9_0),.din(w_dff_A_qpmAS6uv8_0),.clk(gclk));
	jdff dff_A_Zu5gOBWU7_0(.dout(w_dff_A_qpmAS6uv8_0),.din(w_dff_A_Zu5gOBWU7_0),.clk(gclk));
	jdff dff_A_7u2lWCTo1_0(.dout(w_dff_A_Zu5gOBWU7_0),.din(w_dff_A_7u2lWCTo1_0),.clk(gclk));
	jdff dff_A_Tlfzrtja8_0(.dout(w_dff_A_7u2lWCTo1_0),.din(w_dff_A_Tlfzrtja8_0),.clk(gclk));
	jdff dff_A_KULErXji4_0(.dout(w_dff_A_Tlfzrtja8_0),.din(w_dff_A_KULErXji4_0),.clk(gclk));
	jdff dff_A_ZjU4JL573_0(.dout(w_dff_A_KULErXji4_0),.din(w_dff_A_ZjU4JL573_0),.clk(gclk));
	jdff dff_A_sEM64owF5_0(.dout(w_dff_A_ZjU4JL573_0),.din(w_dff_A_sEM64owF5_0),.clk(gclk));
	jdff dff_A_v6J7VqWj2_0(.dout(w_dff_A_sEM64owF5_0),.din(w_dff_A_v6J7VqWj2_0),.clk(gclk));
	jdff dff_A_b6WhIoFW7_0(.dout(w_dff_A_v6J7VqWj2_0),.din(w_dff_A_b6WhIoFW7_0),.clk(gclk));
	jdff dff_A_ssjJfwfn8_0(.dout(w_n445_0[0]),.din(w_dff_A_ssjJfwfn8_0),.clk(gclk));
	jdff dff_B_mGfMoIar4_1(.din(n388),.dout(w_dff_B_mGfMoIar4_1),.clk(gclk));
	jdff dff_A_TVF0ZkmO6_0(.dout(w_n323_0[0]),.din(w_dff_A_TVF0ZkmO6_0),.clk(gclk));
	jdff dff_A_WLXBINEZ5_0(.dout(w_dff_A_TVF0ZkmO6_0),.din(w_dff_A_WLXBINEZ5_0),.clk(gclk));
	jdff dff_A_KZakzYWl0_0(.dout(w_dff_A_WLXBINEZ5_0),.din(w_dff_A_KZakzYWl0_0),.clk(gclk));
	jdff dff_A_U4637zoq2_0(.dout(w_dff_A_KZakzYWl0_0),.din(w_dff_A_U4637zoq2_0),.clk(gclk));
	jdff dff_A_kzE1S2iG5_0(.dout(w_dff_A_U4637zoq2_0),.din(w_dff_A_kzE1S2iG5_0),.clk(gclk));
	jdff dff_A_XNmO402k2_0(.dout(w_dff_A_kzE1S2iG5_0),.din(w_dff_A_XNmO402k2_0),.clk(gclk));
	jdff dff_A_xst5G28g4_0(.dout(w_dff_A_XNmO402k2_0),.din(w_dff_A_xst5G28g4_0),.clk(gclk));
	jdff dff_A_4RW4rLWP5_0(.dout(w_dff_A_xst5G28g4_0),.din(w_dff_A_4RW4rLWP5_0),.clk(gclk));
	jdff dff_A_FaRc3B7l3_0(.dout(w_dff_A_4RW4rLWP5_0),.din(w_dff_A_FaRc3B7l3_0),.clk(gclk));
	jdff dff_A_XPKGPep44_0(.dout(w_dff_A_FaRc3B7l3_0),.din(w_dff_A_XPKGPep44_0),.clk(gclk));
	jdff dff_A_kIObjICQ4_0(.dout(w_dff_A_XPKGPep44_0),.din(w_dff_A_kIObjICQ4_0),.clk(gclk));
	jdff dff_A_siITKYo55_0(.dout(w_dff_A_kIObjICQ4_0),.din(w_dff_A_siITKYo55_0),.clk(gclk));
	jdff dff_A_lbGDJ6Dz9_0(.dout(w_dff_A_siITKYo55_0),.din(w_dff_A_lbGDJ6Dz9_0),.clk(gclk));
	jdff dff_A_dNwyM5om1_0(.dout(w_dff_A_lbGDJ6Dz9_0),.din(w_dff_A_dNwyM5om1_0),.clk(gclk));
	jdff dff_A_ro56wlhL7_0(.dout(w_dff_A_dNwyM5om1_0),.din(w_dff_A_ro56wlhL7_0),.clk(gclk));
	jdff dff_A_nUlHRz308_0(.dout(w_dff_A_ro56wlhL7_0),.din(w_dff_A_nUlHRz308_0),.clk(gclk));
	jdff dff_A_hXXeUypV3_0(.dout(w_dff_A_nUlHRz308_0),.din(w_dff_A_hXXeUypV3_0),.clk(gclk));
	jdff dff_A_fYfhTmPz2_0(.dout(w_dff_A_hXXeUypV3_0),.din(w_dff_A_fYfhTmPz2_0),.clk(gclk));
	jdff dff_A_581ICQAM8_0(.dout(w_dff_A_fYfhTmPz2_0),.din(w_dff_A_581ICQAM8_0),.clk(gclk));
	jdff dff_A_CxufCeoR3_0(.dout(w_dff_A_581ICQAM8_0),.din(w_dff_A_CxufCeoR3_0),.clk(gclk));
	jdff dff_A_t8Y7zL9k1_0(.dout(w_dff_A_CxufCeoR3_0),.din(w_dff_A_t8Y7zL9k1_0),.clk(gclk));
	jdff dff_A_6pazhalA8_0(.dout(w_dff_A_t8Y7zL9k1_0),.din(w_dff_A_6pazhalA8_0),.clk(gclk));
	jdff dff_A_GwuSQdzy9_0(.dout(w_n374_0[0]),.din(w_dff_A_GwuSQdzy9_0),.clk(gclk));
	jdff dff_B_GGzwUl4x8_1(.din(n325),.dout(w_dff_B_GGzwUl4x8_1),.clk(gclk));
	jdff dff_A_DmmuvWkU1_0(.dout(w_n267_0[0]),.din(w_dff_A_DmmuvWkU1_0),.clk(gclk));
	jdff dff_A_hKOdt0Qq9_0(.dout(w_dff_A_DmmuvWkU1_0),.din(w_dff_A_hKOdt0Qq9_0),.clk(gclk));
	jdff dff_A_a27edCMS9_0(.dout(w_dff_A_hKOdt0Qq9_0),.din(w_dff_A_a27edCMS9_0),.clk(gclk));
	jdff dff_A_GJuj7Haa8_0(.dout(w_dff_A_a27edCMS9_0),.din(w_dff_A_GJuj7Haa8_0),.clk(gclk));
	jdff dff_A_vwBnq14B0_0(.dout(w_dff_A_GJuj7Haa8_0),.din(w_dff_A_vwBnq14B0_0),.clk(gclk));
	jdff dff_A_G4vo3dq36_0(.dout(w_dff_A_vwBnq14B0_0),.din(w_dff_A_G4vo3dq36_0),.clk(gclk));
	jdff dff_A_Yyua2LYt9_0(.dout(w_dff_A_G4vo3dq36_0),.din(w_dff_A_Yyua2LYt9_0),.clk(gclk));
	jdff dff_A_QNaXWpn77_0(.dout(w_dff_A_Yyua2LYt9_0),.din(w_dff_A_QNaXWpn77_0),.clk(gclk));
	jdff dff_A_uW9KqhCg7_0(.dout(w_dff_A_QNaXWpn77_0),.din(w_dff_A_uW9KqhCg7_0),.clk(gclk));
	jdff dff_A_MdginEWG5_0(.dout(w_dff_A_uW9KqhCg7_0),.din(w_dff_A_MdginEWG5_0),.clk(gclk));
	jdff dff_A_APVKPNtx4_0(.dout(w_dff_A_MdginEWG5_0),.din(w_dff_A_APVKPNtx4_0),.clk(gclk));
	jdff dff_A_sE3bSTJf9_0(.dout(w_dff_A_APVKPNtx4_0),.din(w_dff_A_sE3bSTJf9_0),.clk(gclk));
	jdff dff_A_eReiMeQq5_0(.dout(w_dff_A_sE3bSTJf9_0),.din(w_dff_A_eReiMeQq5_0),.clk(gclk));
	jdff dff_A_gpito29p2_0(.dout(w_dff_A_eReiMeQq5_0),.din(w_dff_A_gpito29p2_0),.clk(gclk));
	jdff dff_A_4n0Etl6P1_0(.dout(w_dff_A_gpito29p2_0),.din(w_dff_A_4n0Etl6P1_0),.clk(gclk));
	jdff dff_A_RJJcbE8U5_0(.dout(w_dff_A_4n0Etl6P1_0),.din(w_dff_A_RJJcbE8U5_0),.clk(gclk));
	jdff dff_A_CafySYUU0_0(.dout(w_dff_A_RJJcbE8U5_0),.din(w_dff_A_CafySYUU0_0),.clk(gclk));
	jdff dff_A_qgPtQnLD1_0(.dout(w_dff_A_CafySYUU0_0),.din(w_dff_A_qgPtQnLD1_0),.clk(gclk));
	jdff dff_A_8jxZBe6x3_0(.dout(w_dff_A_qgPtQnLD1_0),.din(w_dff_A_8jxZBe6x3_0),.clk(gclk));
	jdff dff_A_Fuhz5ZBN3_0(.dout(w_n311_0[0]),.din(w_dff_A_Fuhz5ZBN3_0),.clk(gclk));
	jdff dff_B_Q4fCHPlP0_1(.din(n269),.dout(w_dff_B_Q4fCHPlP0_1),.clk(gclk));
	jdff dff_A_XZpB9fif1_0(.dout(w_n218_0[0]),.din(w_dff_A_XZpB9fif1_0),.clk(gclk));
	jdff dff_A_yKxOAacz9_0(.dout(w_dff_A_XZpB9fif1_0),.din(w_dff_A_yKxOAacz9_0),.clk(gclk));
	jdff dff_A_N0GyQVKT9_0(.dout(w_dff_A_yKxOAacz9_0),.din(w_dff_A_N0GyQVKT9_0),.clk(gclk));
	jdff dff_A_Xasm4Db38_0(.dout(w_dff_A_N0GyQVKT9_0),.din(w_dff_A_Xasm4Db38_0),.clk(gclk));
	jdff dff_A_pJasGj7f2_0(.dout(w_dff_A_Xasm4Db38_0),.din(w_dff_A_pJasGj7f2_0),.clk(gclk));
	jdff dff_A_X31MRqSb3_0(.dout(w_dff_A_pJasGj7f2_0),.din(w_dff_A_X31MRqSb3_0),.clk(gclk));
	jdff dff_A_FihyutwB7_0(.dout(w_dff_A_X31MRqSb3_0),.din(w_dff_A_FihyutwB7_0),.clk(gclk));
	jdff dff_A_qpSdDf7k8_0(.dout(w_dff_A_FihyutwB7_0),.din(w_dff_A_qpSdDf7k8_0),.clk(gclk));
	jdff dff_A_PgChPnc70_0(.dout(w_dff_A_qpSdDf7k8_0),.din(w_dff_A_PgChPnc70_0),.clk(gclk));
	jdff dff_A_AjcRSVMr6_0(.dout(w_dff_A_PgChPnc70_0),.din(w_dff_A_AjcRSVMr6_0),.clk(gclk));
	jdff dff_A_IWZFFSnZ2_0(.dout(w_dff_A_AjcRSVMr6_0),.din(w_dff_A_IWZFFSnZ2_0),.clk(gclk));
	jdff dff_A_E2i69n038_0(.dout(w_dff_A_IWZFFSnZ2_0),.din(w_dff_A_E2i69n038_0),.clk(gclk));
	jdff dff_A_Ylc8IzWN7_0(.dout(w_dff_A_E2i69n038_0),.din(w_dff_A_Ylc8IzWN7_0),.clk(gclk));
	jdff dff_A_mPMefKtX8_0(.dout(w_dff_A_Ylc8IzWN7_0),.din(w_dff_A_mPMefKtX8_0),.clk(gclk));
	jdff dff_A_YTZMBscv6_0(.dout(w_dff_A_mPMefKtX8_0),.din(w_dff_A_YTZMBscv6_0),.clk(gclk));
	jdff dff_A_XSkiOj6b1_0(.dout(w_dff_A_YTZMBscv6_0),.din(w_dff_A_XSkiOj6b1_0),.clk(gclk));
	jdff dff_A_ZTA4c5vr1_0(.dout(w_n255_0[0]),.din(w_dff_A_ZTA4c5vr1_0),.clk(gclk));
	jdff dff_B_Ij7RFoTe0_1(.din(n220),.dout(w_dff_B_Ij7RFoTe0_1),.clk(gclk));
	jdff dff_A_54yzyJ4a4_0(.dout(w_n176_0[0]),.din(w_dff_A_54yzyJ4a4_0),.clk(gclk));
	jdff dff_A_Lj13HK1f7_0(.dout(w_dff_A_54yzyJ4a4_0),.din(w_dff_A_Lj13HK1f7_0),.clk(gclk));
	jdff dff_A_OAC4kflL1_0(.dout(w_dff_A_Lj13HK1f7_0),.din(w_dff_A_OAC4kflL1_0),.clk(gclk));
	jdff dff_A_aVS7udP02_0(.dout(w_dff_A_OAC4kflL1_0),.din(w_dff_A_aVS7udP02_0),.clk(gclk));
	jdff dff_A_QTcRTf0u6_0(.dout(w_dff_A_aVS7udP02_0),.din(w_dff_A_QTcRTf0u6_0),.clk(gclk));
	jdff dff_A_jNqAMyIU6_0(.dout(w_dff_A_QTcRTf0u6_0),.din(w_dff_A_jNqAMyIU6_0),.clk(gclk));
	jdff dff_A_j7fXsmhR1_0(.dout(w_dff_A_jNqAMyIU6_0),.din(w_dff_A_j7fXsmhR1_0),.clk(gclk));
	jdff dff_A_uSIBpSpI9_0(.dout(w_dff_A_j7fXsmhR1_0),.din(w_dff_A_uSIBpSpI9_0),.clk(gclk));
	jdff dff_A_j73k00YD8_0(.dout(w_dff_A_uSIBpSpI9_0),.din(w_dff_A_j73k00YD8_0),.clk(gclk));
	jdff dff_A_gxnswvGT5_0(.dout(w_dff_A_j73k00YD8_0),.din(w_dff_A_gxnswvGT5_0),.clk(gclk));
	jdff dff_A_hc74l10N9_0(.dout(w_dff_A_gxnswvGT5_0),.din(w_dff_A_hc74l10N9_0),.clk(gclk));
	jdff dff_A_UIFjVK8s3_0(.dout(w_dff_A_hc74l10N9_0),.din(w_dff_A_UIFjVK8s3_0),.clk(gclk));
	jdff dff_A_rnaNxX3p0_0(.dout(w_dff_A_UIFjVK8s3_0),.din(w_dff_A_rnaNxX3p0_0),.clk(gclk));
	jdff dff_A_l1YxZAyV9_0(.dout(w_n206_0[0]),.din(w_dff_A_l1YxZAyV9_0),.clk(gclk));
	jdff dff_B_aBtWMcoy6_1(.din(n178),.dout(w_dff_B_aBtWMcoy6_1),.clk(gclk));
	jdff dff_A_sXPX3wjW9_0(.dout(w_n141_0[0]),.din(w_dff_A_sXPX3wjW9_0),.clk(gclk));
	jdff dff_A_UQmalzHI7_0(.dout(w_dff_A_sXPX3wjW9_0),.din(w_dff_A_UQmalzHI7_0),.clk(gclk));
	jdff dff_A_l6yAl2QV8_0(.dout(w_dff_A_UQmalzHI7_0),.din(w_dff_A_l6yAl2QV8_0),.clk(gclk));
	jdff dff_A_UXk6t5Dm4_0(.dout(w_dff_A_l6yAl2QV8_0),.din(w_dff_A_UXk6t5Dm4_0),.clk(gclk));
	jdff dff_A_svhuoTIV4_0(.dout(w_dff_A_UXk6t5Dm4_0),.din(w_dff_A_svhuoTIV4_0),.clk(gclk));
	jdff dff_A_qzcvBLxm7_0(.dout(w_dff_A_svhuoTIV4_0),.din(w_dff_A_qzcvBLxm7_0),.clk(gclk));
	jdff dff_A_urmjdxk04_0(.dout(w_dff_A_qzcvBLxm7_0),.din(w_dff_A_urmjdxk04_0),.clk(gclk));
	jdff dff_A_wnkYSCaX8_0(.dout(w_dff_A_urmjdxk04_0),.din(w_dff_A_wnkYSCaX8_0),.clk(gclk));
	jdff dff_A_35krV8GY5_0(.dout(w_dff_A_wnkYSCaX8_0),.din(w_dff_A_35krV8GY5_0),.clk(gclk));
	jdff dff_A_qETlHZLX2_0(.dout(w_dff_A_35krV8GY5_0),.din(w_dff_A_qETlHZLX2_0),.clk(gclk));
	jdff dff_A_dgaDtayp4_0(.dout(w_n164_0[0]),.din(w_dff_A_dgaDtayp4_0),.clk(gclk));
	jdff dff_B_DPmtQp9y6_1(.din(n143),.dout(w_dff_B_DPmtQp9y6_1),.clk(gclk));
	jdff dff_A_dWN7is6d5_0(.dout(w_n112_0[0]),.din(w_dff_A_dWN7is6d5_0),.clk(gclk));
	jdff dff_A_QjWMs8ti8_0(.dout(w_dff_A_dWN7is6d5_0),.din(w_dff_A_QjWMs8ti8_0),.clk(gclk));
	jdff dff_A_TD3fKKkG5_0(.dout(w_dff_A_QjWMs8ti8_0),.din(w_dff_A_TD3fKKkG5_0),.clk(gclk));
	jdff dff_A_DCJyXSFZ2_0(.dout(w_dff_A_TD3fKKkG5_0),.din(w_dff_A_DCJyXSFZ2_0),.clk(gclk));
	jdff dff_A_b8ajZ0vy2_0(.dout(w_dff_A_DCJyXSFZ2_0),.din(w_dff_A_b8ajZ0vy2_0),.clk(gclk));
	jdff dff_A_V0PunVvf7_0(.dout(w_dff_A_b8ajZ0vy2_0),.din(w_dff_A_V0PunVvf7_0),.clk(gclk));
	jdff dff_A_sLao2UcO5_0(.dout(w_dff_A_V0PunVvf7_0),.din(w_dff_A_sLao2UcO5_0),.clk(gclk));
	jdff dff_A_iQhZsTBv4_0(.dout(w_n129_0[0]),.din(w_dff_A_iQhZsTBv4_0),.clk(gclk));
	jdff dff_B_665wR8I06_1(.din(n114),.dout(w_dff_B_665wR8I06_1),.clk(gclk));
	jdff dff_A_uNlohcFg2_0(.dout(w_n91_0[0]),.din(w_dff_A_uNlohcFg2_0),.clk(gclk));
	jdff dff_A_GbQgXPnf5_0(.dout(w_dff_A_uNlohcFg2_0),.din(w_dff_A_GbQgXPnf5_0),.clk(gclk));
	jdff dff_A_UEeEy5Yb0_0(.dout(w_dff_A_GbQgXPnf5_0),.din(w_dff_A_UEeEy5Yb0_0),.clk(gclk));
	jdff dff_A_ekScY5O94_0(.dout(w_dff_A_UEeEy5Yb0_0),.din(w_dff_A_ekScY5O94_0),.clk(gclk));
	jdff dff_B_lUl1Ec815_0(.din(n100),.dout(w_dff_B_lUl1Ec815_0),.clk(gclk));
	jdff dff_A_Xm4Ois8X2_0(.dout(w_n80_0[0]),.din(w_dff_A_Xm4Ois8X2_0),.clk(gclk));
	jdff dff_A_MTFXj9jv8_0(.dout(w_n1119_0[0]),.din(w_dff_A_MTFXj9jv8_0),.clk(gclk));
	jdff dff_B_TE7IUzHw6_2(.din(n1119),.dout(w_dff_B_TE7IUzHw6_2),.clk(gclk));
	jdff dff_B_m2D92t4A6_2(.din(n1018),.dout(w_dff_B_m2D92t4A6_2),.clk(gclk));
	jdff dff_B_KvJmMPCZ2_2(.din(w_dff_B_m2D92t4A6_2),.dout(w_dff_B_KvJmMPCZ2_2),.clk(gclk));
	jdff dff_B_TUmgFBeP4_2(.din(w_dff_B_KvJmMPCZ2_2),.dout(w_dff_B_TUmgFBeP4_2),.clk(gclk));
	jdff dff_B_zfbUrtA34_2(.din(w_dff_B_TUmgFBeP4_2),.dout(w_dff_B_zfbUrtA34_2),.clk(gclk));
	jdff dff_B_RJeRf19S1_2(.din(w_dff_B_zfbUrtA34_2),.dout(w_dff_B_RJeRf19S1_2),.clk(gclk));
	jdff dff_B_y99PNr7M2_2(.din(w_dff_B_RJeRf19S1_2),.dout(w_dff_B_y99PNr7M2_2),.clk(gclk));
	jdff dff_B_NdhpUcr03_2(.din(w_dff_B_y99PNr7M2_2),.dout(w_dff_B_NdhpUcr03_2),.clk(gclk));
	jdff dff_B_Ofo8b89l6_2(.din(w_dff_B_NdhpUcr03_2),.dout(w_dff_B_Ofo8b89l6_2),.clk(gclk));
	jdff dff_B_TzIJma0E4_2(.din(w_dff_B_Ofo8b89l6_2),.dout(w_dff_B_TzIJma0E4_2),.clk(gclk));
	jdff dff_B_TPKlGYzw5_2(.din(w_dff_B_TzIJma0E4_2),.dout(w_dff_B_TPKlGYzw5_2),.clk(gclk));
	jdff dff_B_YeQLhzxq8_2(.din(w_dff_B_TPKlGYzw5_2),.dout(w_dff_B_YeQLhzxq8_2),.clk(gclk));
	jdff dff_B_jcEzTYw38_2(.din(w_dff_B_YeQLhzxq8_2),.dout(w_dff_B_jcEzTYw38_2),.clk(gclk));
	jdff dff_B_5GsClUeS8_2(.din(w_dff_B_jcEzTYw38_2),.dout(w_dff_B_5GsClUeS8_2),.clk(gclk));
	jdff dff_B_wNpxeUlw1_2(.din(w_dff_B_5GsClUeS8_2),.dout(w_dff_B_wNpxeUlw1_2),.clk(gclk));
	jdff dff_B_5mnpL7rk9_2(.din(w_dff_B_wNpxeUlw1_2),.dout(w_dff_B_5mnpL7rk9_2),.clk(gclk));
	jdff dff_B_iLMfAYs48_2(.din(w_dff_B_5mnpL7rk9_2),.dout(w_dff_B_iLMfAYs48_2),.clk(gclk));
	jdff dff_B_6JYjTF0m1_2(.din(w_dff_B_iLMfAYs48_2),.dout(w_dff_B_6JYjTF0m1_2),.clk(gclk));
	jdff dff_B_GiFFH6du6_2(.din(w_dff_B_6JYjTF0m1_2),.dout(w_dff_B_GiFFH6du6_2),.clk(gclk));
	jdff dff_B_xaPCS9GA0_2(.din(w_dff_B_GiFFH6du6_2),.dout(w_dff_B_xaPCS9GA0_2),.clk(gclk));
	jdff dff_B_QupNyiK51_2(.din(w_dff_B_xaPCS9GA0_2),.dout(w_dff_B_QupNyiK51_2),.clk(gclk));
	jdff dff_B_zfECBIgh9_2(.din(w_dff_B_QupNyiK51_2),.dout(w_dff_B_zfECBIgh9_2),.clk(gclk));
	jdff dff_B_tZqpdtqD4_2(.din(w_dff_B_zfECBIgh9_2),.dout(w_dff_B_tZqpdtqD4_2),.clk(gclk));
	jdff dff_B_cb9E4iQu3_2(.din(w_dff_B_tZqpdtqD4_2),.dout(w_dff_B_cb9E4iQu3_2),.clk(gclk));
	jdff dff_B_lIxqaB019_2(.din(w_dff_B_cb9E4iQu3_2),.dout(w_dff_B_lIxqaB019_2),.clk(gclk));
	jdff dff_B_rebp5DpQ9_2(.din(w_dff_B_lIxqaB019_2),.dout(w_dff_B_rebp5DpQ9_2),.clk(gclk));
	jdff dff_B_qockIgX34_2(.din(w_dff_B_rebp5DpQ9_2),.dout(w_dff_B_qockIgX34_2),.clk(gclk));
	jdff dff_B_H1ZRfpr80_2(.din(w_dff_B_qockIgX34_2),.dout(w_dff_B_H1ZRfpr80_2),.clk(gclk));
	jdff dff_B_L9MWqCdD2_2(.din(w_dff_B_H1ZRfpr80_2),.dout(w_dff_B_L9MWqCdD2_2),.clk(gclk));
	jdff dff_B_MwCkCbO47_2(.din(w_dff_B_L9MWqCdD2_2),.dout(w_dff_B_MwCkCbO47_2),.clk(gclk));
	jdff dff_B_Tnvf8DVQ3_2(.din(w_dff_B_MwCkCbO47_2),.dout(w_dff_B_Tnvf8DVQ3_2),.clk(gclk));
	jdff dff_B_RDWDIazy7_2(.din(w_dff_B_Tnvf8DVQ3_2),.dout(w_dff_B_RDWDIazy7_2),.clk(gclk));
	jdff dff_B_ulTm7mSm4_2(.din(w_dff_B_RDWDIazy7_2),.dout(w_dff_B_ulTm7mSm4_2),.clk(gclk));
	jdff dff_B_7oVIdcJM4_2(.din(w_dff_B_ulTm7mSm4_2),.dout(w_dff_B_7oVIdcJM4_2),.clk(gclk));
	jdff dff_B_3dgdwS6e4_2(.din(w_dff_B_7oVIdcJM4_2),.dout(w_dff_B_3dgdwS6e4_2),.clk(gclk));
	jdff dff_B_McpLEPzu8_2(.din(w_dff_B_3dgdwS6e4_2),.dout(w_dff_B_McpLEPzu8_2),.clk(gclk));
	jdff dff_B_IcRXRP7O7_2(.din(w_dff_B_McpLEPzu8_2),.dout(w_dff_B_IcRXRP7O7_2),.clk(gclk));
	jdff dff_B_K7d4hIjO0_2(.din(w_dff_B_IcRXRP7O7_2),.dout(w_dff_B_K7d4hIjO0_2),.clk(gclk));
	jdff dff_B_GK5aTa5s1_2(.din(w_dff_B_K7d4hIjO0_2),.dout(w_dff_B_GK5aTa5s1_2),.clk(gclk));
	jdff dff_B_OfZUHjtI3_2(.din(w_dff_B_GK5aTa5s1_2),.dout(w_dff_B_OfZUHjtI3_2),.clk(gclk));
	jdff dff_B_MJKSD1ir7_2(.din(w_dff_B_OfZUHjtI3_2),.dout(w_dff_B_MJKSD1ir7_2),.clk(gclk));
	jdff dff_B_omBAHzXb1_2(.din(w_dff_B_MJKSD1ir7_2),.dout(w_dff_B_omBAHzXb1_2),.clk(gclk));
	jdff dff_B_cvsacRiZ6_2(.din(w_dff_B_omBAHzXb1_2),.dout(w_dff_B_cvsacRiZ6_2),.clk(gclk));
	jdff dff_B_5NNsqtcs0_2(.din(w_dff_B_cvsacRiZ6_2),.dout(w_dff_B_5NNsqtcs0_2),.clk(gclk));
	jdff dff_A_jtq9VIji0_0(.dout(w_n1022_0[0]),.din(w_dff_A_jtq9VIji0_0),.clk(gclk));
	jdff dff_B_L4bM11W03_1(.din(n1020),.dout(w_dff_B_L4bM11W03_1),.clk(gclk));
	jdff dff_B_NXpybWVb0_2(.din(n916),.dout(w_dff_B_NXpybWVb0_2),.clk(gclk));
	jdff dff_B_SNfaZxqY4_2(.din(w_dff_B_NXpybWVb0_2),.dout(w_dff_B_SNfaZxqY4_2),.clk(gclk));
	jdff dff_B_unmECFzh3_2(.din(w_dff_B_SNfaZxqY4_2),.dout(w_dff_B_unmECFzh3_2),.clk(gclk));
	jdff dff_B_lzeeD1D73_2(.din(w_dff_B_unmECFzh3_2),.dout(w_dff_B_lzeeD1D73_2),.clk(gclk));
	jdff dff_B_pV981ygm7_2(.din(w_dff_B_lzeeD1D73_2),.dout(w_dff_B_pV981ygm7_2),.clk(gclk));
	jdff dff_B_US0csvFV5_2(.din(w_dff_B_pV981ygm7_2),.dout(w_dff_B_US0csvFV5_2),.clk(gclk));
	jdff dff_B_gjQBVSZT0_2(.din(w_dff_B_US0csvFV5_2),.dout(w_dff_B_gjQBVSZT0_2),.clk(gclk));
	jdff dff_B_7XS5vAmo3_2(.din(w_dff_B_gjQBVSZT0_2),.dout(w_dff_B_7XS5vAmo3_2),.clk(gclk));
	jdff dff_B_y7jSaYIm2_2(.din(w_dff_B_7XS5vAmo3_2),.dout(w_dff_B_y7jSaYIm2_2),.clk(gclk));
	jdff dff_B_7X16aKI65_2(.din(w_dff_B_y7jSaYIm2_2),.dout(w_dff_B_7X16aKI65_2),.clk(gclk));
	jdff dff_B_dYzLpyIv9_2(.din(w_dff_B_7X16aKI65_2),.dout(w_dff_B_dYzLpyIv9_2),.clk(gclk));
	jdff dff_B_DEqnNIst6_2(.din(w_dff_B_dYzLpyIv9_2),.dout(w_dff_B_DEqnNIst6_2),.clk(gclk));
	jdff dff_B_ttTgWAgs7_2(.din(w_dff_B_DEqnNIst6_2),.dout(w_dff_B_ttTgWAgs7_2),.clk(gclk));
	jdff dff_B_aQr5yUPV7_2(.din(w_dff_B_ttTgWAgs7_2),.dout(w_dff_B_aQr5yUPV7_2),.clk(gclk));
	jdff dff_B_tkqZrdFq3_2(.din(w_dff_B_aQr5yUPV7_2),.dout(w_dff_B_tkqZrdFq3_2),.clk(gclk));
	jdff dff_B_UtvbkyQV0_2(.din(w_dff_B_tkqZrdFq3_2),.dout(w_dff_B_UtvbkyQV0_2),.clk(gclk));
	jdff dff_B_YYmzVbct7_2(.din(w_dff_B_UtvbkyQV0_2),.dout(w_dff_B_YYmzVbct7_2),.clk(gclk));
	jdff dff_B_yg1oDqeG3_2(.din(w_dff_B_YYmzVbct7_2),.dout(w_dff_B_yg1oDqeG3_2),.clk(gclk));
	jdff dff_B_QN6STyxv3_2(.din(w_dff_B_yg1oDqeG3_2),.dout(w_dff_B_QN6STyxv3_2),.clk(gclk));
	jdff dff_B_saMXTMqk2_2(.din(w_dff_B_QN6STyxv3_2),.dout(w_dff_B_saMXTMqk2_2),.clk(gclk));
	jdff dff_B_qO0D7mff5_2(.din(w_dff_B_saMXTMqk2_2),.dout(w_dff_B_qO0D7mff5_2),.clk(gclk));
	jdff dff_B_aNSdxiyd0_2(.din(w_dff_B_qO0D7mff5_2),.dout(w_dff_B_aNSdxiyd0_2),.clk(gclk));
	jdff dff_B_uM4KoRwI5_2(.din(w_dff_B_aNSdxiyd0_2),.dout(w_dff_B_uM4KoRwI5_2),.clk(gclk));
	jdff dff_B_eutStpg04_2(.din(w_dff_B_uM4KoRwI5_2),.dout(w_dff_B_eutStpg04_2),.clk(gclk));
	jdff dff_B_Fpge5zU09_2(.din(w_dff_B_eutStpg04_2),.dout(w_dff_B_Fpge5zU09_2),.clk(gclk));
	jdff dff_B_UDRrIOuF2_2(.din(w_dff_B_Fpge5zU09_2),.dout(w_dff_B_UDRrIOuF2_2),.clk(gclk));
	jdff dff_B_2M7o3Xm55_2(.din(w_dff_B_UDRrIOuF2_2),.dout(w_dff_B_2M7o3Xm55_2),.clk(gclk));
	jdff dff_B_NMt9eYEZ2_2(.din(w_dff_B_2M7o3Xm55_2),.dout(w_dff_B_NMt9eYEZ2_2),.clk(gclk));
	jdff dff_B_M8PEl6yE4_2(.din(w_dff_B_NMt9eYEZ2_2),.dout(w_dff_B_M8PEl6yE4_2),.clk(gclk));
	jdff dff_B_F8UOjfwp2_2(.din(w_dff_B_M8PEl6yE4_2),.dout(w_dff_B_F8UOjfwp2_2),.clk(gclk));
	jdff dff_B_BF8davyZ9_2(.din(w_dff_B_F8UOjfwp2_2),.dout(w_dff_B_BF8davyZ9_2),.clk(gclk));
	jdff dff_B_nH9dYGtR9_2(.din(w_dff_B_BF8davyZ9_2),.dout(w_dff_B_nH9dYGtR9_2),.clk(gclk));
	jdff dff_B_sVIqy5wP8_2(.din(w_dff_B_nH9dYGtR9_2),.dout(w_dff_B_sVIqy5wP8_2),.clk(gclk));
	jdff dff_B_Magq2tLW1_2(.din(w_dff_B_sVIqy5wP8_2),.dout(w_dff_B_Magq2tLW1_2),.clk(gclk));
	jdff dff_B_42odInzz4_2(.din(w_dff_B_Magq2tLW1_2),.dout(w_dff_B_42odInzz4_2),.clk(gclk));
	jdff dff_B_5JqZnrUw2_2(.din(w_dff_B_42odInzz4_2),.dout(w_dff_B_5JqZnrUw2_2),.clk(gclk));
	jdff dff_B_ySZqLxuy4_2(.din(w_dff_B_5JqZnrUw2_2),.dout(w_dff_B_ySZqLxuy4_2),.clk(gclk));
	jdff dff_B_E5urkzbu4_2(.din(w_dff_B_ySZqLxuy4_2),.dout(w_dff_B_E5urkzbu4_2),.clk(gclk));
	jdff dff_B_Gp3sfWDO7_2(.din(w_dff_B_E5urkzbu4_2),.dout(w_dff_B_Gp3sfWDO7_2),.clk(gclk));
	jdff dff_B_GiPGGvU81_2(.din(w_dff_B_Gp3sfWDO7_2),.dout(w_dff_B_GiPGGvU81_2),.clk(gclk));
	jdff dff_A_hYbFF23a1_1(.dout(w_n1006_0[1]),.din(w_dff_A_hYbFF23a1_1),.clk(gclk));
	jdff dff_A_UvLQDDSv5_0(.dout(w_n816_0[0]),.din(w_dff_A_UvLQDDSv5_0),.clk(gclk));
	jdff dff_A_kstmPLp70_0(.dout(w_dff_A_UvLQDDSv5_0),.din(w_dff_A_kstmPLp70_0),.clk(gclk));
	jdff dff_A_wFyE6uTZ6_0(.dout(w_dff_A_kstmPLp70_0),.din(w_dff_A_wFyE6uTZ6_0),.clk(gclk));
	jdff dff_A_nSRMrK0O5_0(.dout(w_dff_A_wFyE6uTZ6_0),.din(w_dff_A_nSRMrK0O5_0),.clk(gclk));
	jdff dff_A_MC0Qs3eK4_0(.dout(w_dff_A_nSRMrK0O5_0),.din(w_dff_A_MC0Qs3eK4_0),.clk(gclk));
	jdff dff_A_Bnu8nZuB0_0(.dout(w_dff_A_MC0Qs3eK4_0),.din(w_dff_A_Bnu8nZuB0_0),.clk(gclk));
	jdff dff_A_ljA7cAPy1_0(.dout(w_dff_A_Bnu8nZuB0_0),.din(w_dff_A_ljA7cAPy1_0),.clk(gclk));
	jdff dff_A_vFuPo2Il1_0(.dout(w_dff_A_ljA7cAPy1_0),.din(w_dff_A_vFuPo2Il1_0),.clk(gclk));
	jdff dff_A_RlpAuLPe3_0(.dout(w_dff_A_vFuPo2Il1_0),.din(w_dff_A_RlpAuLPe3_0),.clk(gclk));
	jdff dff_A_nXICAeIO3_0(.dout(w_dff_A_RlpAuLPe3_0),.din(w_dff_A_nXICAeIO3_0),.clk(gclk));
	jdff dff_A_BdIuxJW48_0(.dout(w_dff_A_nXICAeIO3_0),.din(w_dff_A_BdIuxJW48_0),.clk(gclk));
	jdff dff_A_iIRk5VLh5_0(.dout(w_dff_A_BdIuxJW48_0),.din(w_dff_A_iIRk5VLh5_0),.clk(gclk));
	jdff dff_A_ezUAFxHZ1_0(.dout(w_dff_A_iIRk5VLh5_0),.din(w_dff_A_ezUAFxHZ1_0),.clk(gclk));
	jdff dff_A_PeIArAzX7_0(.dout(w_dff_A_ezUAFxHZ1_0),.din(w_dff_A_PeIArAzX7_0),.clk(gclk));
	jdff dff_A_1zWLdJ3N7_0(.dout(w_dff_A_PeIArAzX7_0),.din(w_dff_A_1zWLdJ3N7_0),.clk(gclk));
	jdff dff_A_kB0tQKH79_0(.dout(w_dff_A_1zWLdJ3N7_0),.din(w_dff_A_kB0tQKH79_0),.clk(gclk));
	jdff dff_A_73wH3RgH5_0(.dout(w_dff_A_kB0tQKH79_0),.din(w_dff_A_73wH3RgH5_0),.clk(gclk));
	jdff dff_A_twPON9eS6_0(.dout(w_dff_A_73wH3RgH5_0),.din(w_dff_A_twPON9eS6_0),.clk(gclk));
	jdff dff_A_9O3gJxRv3_0(.dout(w_dff_A_twPON9eS6_0),.din(w_dff_A_9O3gJxRv3_0),.clk(gclk));
	jdff dff_A_7lk4NUJ14_0(.dout(w_dff_A_9O3gJxRv3_0),.din(w_dff_A_7lk4NUJ14_0),.clk(gclk));
	jdff dff_A_HKw6jIgO9_0(.dout(w_dff_A_7lk4NUJ14_0),.din(w_dff_A_HKw6jIgO9_0),.clk(gclk));
	jdff dff_A_U2qgJ6413_0(.dout(w_dff_A_HKw6jIgO9_0),.din(w_dff_A_U2qgJ6413_0),.clk(gclk));
	jdff dff_A_VQsAhFVy1_0(.dout(w_dff_A_U2qgJ6413_0),.din(w_dff_A_VQsAhFVy1_0),.clk(gclk));
	jdff dff_A_XdrIhCRw8_0(.dout(w_dff_A_VQsAhFVy1_0),.din(w_dff_A_XdrIhCRw8_0),.clk(gclk));
	jdff dff_A_HEXadBW79_0(.dout(w_dff_A_XdrIhCRw8_0),.din(w_dff_A_HEXadBW79_0),.clk(gclk));
	jdff dff_A_3PsCWxAH3_0(.dout(w_dff_A_HEXadBW79_0),.din(w_dff_A_3PsCWxAH3_0),.clk(gclk));
	jdff dff_A_KEHKnKex5_0(.dout(w_dff_A_3PsCWxAH3_0),.din(w_dff_A_KEHKnKex5_0),.clk(gclk));
	jdff dff_A_iodJtMTu7_0(.dout(w_dff_A_KEHKnKex5_0),.din(w_dff_A_iodJtMTu7_0),.clk(gclk));
	jdff dff_A_FWLtlRdZ9_0(.dout(w_dff_A_iodJtMTu7_0),.din(w_dff_A_FWLtlRdZ9_0),.clk(gclk));
	jdff dff_A_oQaM2Mvm7_0(.dout(w_dff_A_FWLtlRdZ9_0),.din(w_dff_A_oQaM2Mvm7_0),.clk(gclk));
	jdff dff_A_v3G458jc4_0(.dout(w_dff_A_oQaM2Mvm7_0),.din(w_dff_A_v3G458jc4_0),.clk(gclk));
	jdff dff_A_mFXfWBcB2_0(.dout(w_dff_A_v3G458jc4_0),.din(w_dff_A_mFXfWBcB2_0),.clk(gclk));
	jdff dff_A_ZB7ACmPt8_0(.dout(w_dff_A_mFXfWBcB2_0),.din(w_dff_A_ZB7ACmPt8_0),.clk(gclk));
	jdff dff_A_LcHzCn9O8_0(.dout(w_dff_A_ZB7ACmPt8_0),.din(w_dff_A_LcHzCn9O8_0),.clk(gclk));
	jdff dff_A_kOMYAdAY8_0(.dout(w_dff_A_LcHzCn9O8_0),.din(w_dff_A_kOMYAdAY8_0),.clk(gclk));
	jdff dff_A_H8PJtw943_0(.dout(w_dff_A_kOMYAdAY8_0),.din(w_dff_A_H8PJtw943_0),.clk(gclk));
	jdff dff_A_B8itLeCq2_0(.dout(w_dff_A_H8PJtw943_0),.din(w_dff_A_B8itLeCq2_0),.clk(gclk));
	jdff dff_A_Pt0afR317_1(.dout(w_n900_0[1]),.din(w_dff_A_Pt0afR317_1),.clk(gclk));
	jdff dff_A_0aocDaWj8_2(.dout(w_n900_0[2]),.din(w_dff_A_0aocDaWj8_2),.clk(gclk));
	jdff dff_B_dNQi9PLH0_1(.din(n818),.dout(w_dff_B_dNQi9PLH0_1),.clk(gclk));
	jdff dff_B_P5kqbM7h2_2(.din(n719),.dout(w_dff_B_P5kqbM7h2_2),.clk(gclk));
	jdff dff_B_PPyj4RN67_2(.din(w_dff_B_P5kqbM7h2_2),.dout(w_dff_B_PPyj4RN67_2),.clk(gclk));
	jdff dff_B_FTZvdhQU1_2(.din(w_dff_B_PPyj4RN67_2),.dout(w_dff_B_FTZvdhQU1_2),.clk(gclk));
	jdff dff_B_I5b0sp8H6_2(.din(w_dff_B_FTZvdhQU1_2),.dout(w_dff_B_I5b0sp8H6_2),.clk(gclk));
	jdff dff_B_ihd7apOB8_2(.din(w_dff_B_I5b0sp8H6_2),.dout(w_dff_B_ihd7apOB8_2),.clk(gclk));
	jdff dff_B_iNmPesNL5_2(.din(w_dff_B_ihd7apOB8_2),.dout(w_dff_B_iNmPesNL5_2),.clk(gclk));
	jdff dff_B_idfNLey56_2(.din(w_dff_B_iNmPesNL5_2),.dout(w_dff_B_idfNLey56_2),.clk(gclk));
	jdff dff_B_Eyv94Qvs4_2(.din(w_dff_B_idfNLey56_2),.dout(w_dff_B_Eyv94Qvs4_2),.clk(gclk));
	jdff dff_B_OMl5hO618_2(.din(w_dff_B_Eyv94Qvs4_2),.dout(w_dff_B_OMl5hO618_2),.clk(gclk));
	jdff dff_B_QO7kxPFe6_2(.din(w_dff_B_OMl5hO618_2),.dout(w_dff_B_QO7kxPFe6_2),.clk(gclk));
	jdff dff_B_vT1oA9iS5_2(.din(w_dff_B_QO7kxPFe6_2),.dout(w_dff_B_vT1oA9iS5_2),.clk(gclk));
	jdff dff_B_raYfew9D8_2(.din(w_dff_B_vT1oA9iS5_2),.dout(w_dff_B_raYfew9D8_2),.clk(gclk));
	jdff dff_B_tOGUTWXH3_2(.din(w_dff_B_raYfew9D8_2),.dout(w_dff_B_tOGUTWXH3_2),.clk(gclk));
	jdff dff_B_p2kaPQWR6_2(.din(w_dff_B_tOGUTWXH3_2),.dout(w_dff_B_p2kaPQWR6_2),.clk(gclk));
	jdff dff_B_UoFZvXiB8_2(.din(w_dff_B_p2kaPQWR6_2),.dout(w_dff_B_UoFZvXiB8_2),.clk(gclk));
	jdff dff_B_zT0Yk9Hi4_2(.din(w_dff_B_UoFZvXiB8_2),.dout(w_dff_B_zT0Yk9Hi4_2),.clk(gclk));
	jdff dff_B_rNqmNcCx6_2(.din(w_dff_B_zT0Yk9Hi4_2),.dout(w_dff_B_rNqmNcCx6_2),.clk(gclk));
	jdff dff_B_lv1SRQXi1_2(.din(w_dff_B_rNqmNcCx6_2),.dout(w_dff_B_lv1SRQXi1_2),.clk(gclk));
	jdff dff_B_MdZkpYz10_2(.din(w_dff_B_lv1SRQXi1_2),.dout(w_dff_B_MdZkpYz10_2),.clk(gclk));
	jdff dff_B_bZRHx9if7_2(.din(w_dff_B_MdZkpYz10_2),.dout(w_dff_B_bZRHx9if7_2),.clk(gclk));
	jdff dff_B_PY2wD7eq7_2(.din(w_dff_B_bZRHx9if7_2),.dout(w_dff_B_PY2wD7eq7_2),.clk(gclk));
	jdff dff_B_b8D34B625_2(.din(w_dff_B_PY2wD7eq7_2),.dout(w_dff_B_b8D34B625_2),.clk(gclk));
	jdff dff_B_fAxKGH039_2(.din(w_dff_B_b8D34B625_2),.dout(w_dff_B_fAxKGH039_2),.clk(gclk));
	jdff dff_B_3n01StlD6_2(.din(w_dff_B_fAxKGH039_2),.dout(w_dff_B_3n01StlD6_2),.clk(gclk));
	jdff dff_B_8AXscg2M5_2(.din(w_dff_B_3n01StlD6_2),.dout(w_dff_B_8AXscg2M5_2),.clk(gclk));
	jdff dff_B_stLbKPUz1_2(.din(w_dff_B_8AXscg2M5_2),.dout(w_dff_B_stLbKPUz1_2),.clk(gclk));
	jdff dff_B_4JcNNLnI1_2(.din(w_dff_B_stLbKPUz1_2),.dout(w_dff_B_4JcNNLnI1_2),.clk(gclk));
	jdff dff_B_KcbvCYKb7_2(.din(w_dff_B_4JcNNLnI1_2),.dout(w_dff_B_KcbvCYKb7_2),.clk(gclk));
	jdff dff_B_A5OQRGhH1_2(.din(w_dff_B_KcbvCYKb7_2),.dout(w_dff_B_A5OQRGhH1_2),.clk(gclk));
	jdff dff_B_E1rZKPON0_2(.din(w_dff_B_A5OQRGhH1_2),.dout(w_dff_B_E1rZKPON0_2),.clk(gclk));
	jdff dff_B_ErlpDTqi1_2(.din(w_dff_B_E1rZKPON0_2),.dout(w_dff_B_ErlpDTqi1_2),.clk(gclk));
	jdff dff_B_NJuq3n8J9_2(.din(w_dff_B_ErlpDTqi1_2),.dout(w_dff_B_NJuq3n8J9_2),.clk(gclk));
	jdff dff_B_LMMTeiyX9_2(.din(w_dff_B_NJuq3n8J9_2),.dout(w_dff_B_LMMTeiyX9_2),.clk(gclk));
	jdff dff_B_ah10LIvS1_2(.din(n797),.dout(w_dff_B_ah10LIvS1_2),.clk(gclk));
	jdff dff_B_Dlogfoix6_1(.din(n720),.dout(w_dff_B_Dlogfoix6_1),.clk(gclk));
	jdff dff_B_I5qByQ2b0_2(.din(n627),.dout(w_dff_B_I5qByQ2b0_2),.clk(gclk));
	jdff dff_B_AM9CuuDy7_2(.din(w_dff_B_I5qByQ2b0_2),.dout(w_dff_B_AM9CuuDy7_2),.clk(gclk));
	jdff dff_B_Ltm5NdKr8_2(.din(w_dff_B_AM9CuuDy7_2),.dout(w_dff_B_Ltm5NdKr8_2),.clk(gclk));
	jdff dff_B_F5yvn08P8_2(.din(w_dff_B_Ltm5NdKr8_2),.dout(w_dff_B_F5yvn08P8_2),.clk(gclk));
	jdff dff_B_2v9bMgNf8_2(.din(w_dff_B_F5yvn08P8_2),.dout(w_dff_B_2v9bMgNf8_2),.clk(gclk));
	jdff dff_B_7wzU8vK20_2(.din(w_dff_B_2v9bMgNf8_2),.dout(w_dff_B_7wzU8vK20_2),.clk(gclk));
	jdff dff_B_tb8bruCo5_2(.din(w_dff_B_7wzU8vK20_2),.dout(w_dff_B_tb8bruCo5_2),.clk(gclk));
	jdff dff_B_VS5c4Ex44_2(.din(w_dff_B_tb8bruCo5_2),.dout(w_dff_B_VS5c4Ex44_2),.clk(gclk));
	jdff dff_B_gPlquzEW3_2(.din(w_dff_B_VS5c4Ex44_2),.dout(w_dff_B_gPlquzEW3_2),.clk(gclk));
	jdff dff_B_kBc74Hlf1_2(.din(w_dff_B_gPlquzEW3_2),.dout(w_dff_B_kBc74Hlf1_2),.clk(gclk));
	jdff dff_B_9hlGbQcB1_2(.din(w_dff_B_kBc74Hlf1_2),.dout(w_dff_B_9hlGbQcB1_2),.clk(gclk));
	jdff dff_B_JKc2WJVm2_2(.din(w_dff_B_9hlGbQcB1_2),.dout(w_dff_B_JKc2WJVm2_2),.clk(gclk));
	jdff dff_B_DMgHGdz74_2(.din(w_dff_B_JKc2WJVm2_2),.dout(w_dff_B_DMgHGdz74_2),.clk(gclk));
	jdff dff_B_GjsClQzy5_2(.din(w_dff_B_DMgHGdz74_2),.dout(w_dff_B_GjsClQzy5_2),.clk(gclk));
	jdff dff_B_Y6EvD0z66_2(.din(w_dff_B_GjsClQzy5_2),.dout(w_dff_B_Y6EvD0z66_2),.clk(gclk));
	jdff dff_B_MOibOGLg5_2(.din(w_dff_B_Y6EvD0z66_2),.dout(w_dff_B_MOibOGLg5_2),.clk(gclk));
	jdff dff_B_Tp1Yx1iJ6_2(.din(w_dff_B_MOibOGLg5_2),.dout(w_dff_B_Tp1Yx1iJ6_2),.clk(gclk));
	jdff dff_B_5susflEF9_2(.din(w_dff_B_Tp1Yx1iJ6_2),.dout(w_dff_B_5susflEF9_2),.clk(gclk));
	jdff dff_B_p2w1ZfdA3_2(.din(w_dff_B_5susflEF9_2),.dout(w_dff_B_p2w1ZfdA3_2),.clk(gclk));
	jdff dff_B_hycbdnRu4_2(.din(w_dff_B_p2w1ZfdA3_2),.dout(w_dff_B_hycbdnRu4_2),.clk(gclk));
	jdff dff_B_0qEocB764_2(.din(w_dff_B_hycbdnRu4_2),.dout(w_dff_B_0qEocB764_2),.clk(gclk));
	jdff dff_B_E1EsZ7Zp7_2(.din(w_dff_B_0qEocB764_2),.dout(w_dff_B_E1EsZ7Zp7_2),.clk(gclk));
	jdff dff_B_fTpHpzeg2_2(.din(w_dff_B_E1EsZ7Zp7_2),.dout(w_dff_B_fTpHpzeg2_2),.clk(gclk));
	jdff dff_B_S4CnyiCq6_2(.din(w_dff_B_fTpHpzeg2_2),.dout(w_dff_B_S4CnyiCq6_2),.clk(gclk));
	jdff dff_B_vZTI7Q4v9_2(.din(w_dff_B_S4CnyiCq6_2),.dout(w_dff_B_vZTI7Q4v9_2),.clk(gclk));
	jdff dff_B_PYZxaz5r4_2(.din(w_dff_B_vZTI7Q4v9_2),.dout(w_dff_B_PYZxaz5r4_2),.clk(gclk));
	jdff dff_B_Oazy7wZj8_2(.din(w_dff_B_PYZxaz5r4_2),.dout(w_dff_B_Oazy7wZj8_2),.clk(gclk));
	jdff dff_B_Xg8h8zKW0_2(.din(w_dff_B_Oazy7wZj8_2),.dout(w_dff_B_Xg8h8zKW0_2),.clk(gclk));
	jdff dff_B_KwQq9Pvw0_2(.din(w_dff_B_Xg8h8zKW0_2),.dout(w_dff_B_KwQq9Pvw0_2),.clk(gclk));
	jdff dff_B_uCo2WFDQ7_2(.din(w_dff_B_KwQq9Pvw0_2),.dout(w_dff_B_uCo2WFDQ7_2),.clk(gclk));
	jdff dff_B_BpsdmnhP5_2(.din(n698),.dout(w_dff_B_BpsdmnhP5_2),.clk(gclk));
	jdff dff_B_VlAwclpH3_1(.din(n628),.dout(w_dff_B_VlAwclpH3_1),.clk(gclk));
	jdff dff_B_frsO1YE89_2(.din(n542),.dout(w_dff_B_frsO1YE89_2),.clk(gclk));
	jdff dff_B_q2OIXh6o9_2(.din(w_dff_B_frsO1YE89_2),.dout(w_dff_B_q2OIXh6o9_2),.clk(gclk));
	jdff dff_B_AOPQ8Cgv5_2(.din(w_dff_B_q2OIXh6o9_2),.dout(w_dff_B_AOPQ8Cgv5_2),.clk(gclk));
	jdff dff_B_3tgNZQ2M5_2(.din(w_dff_B_AOPQ8Cgv5_2),.dout(w_dff_B_3tgNZQ2M5_2),.clk(gclk));
	jdff dff_B_3tOvUodx0_2(.din(w_dff_B_3tgNZQ2M5_2),.dout(w_dff_B_3tOvUodx0_2),.clk(gclk));
	jdff dff_B_Qf7Ol6hQ5_2(.din(w_dff_B_3tOvUodx0_2),.dout(w_dff_B_Qf7Ol6hQ5_2),.clk(gclk));
	jdff dff_B_gvOhazXT0_2(.din(w_dff_B_Qf7Ol6hQ5_2),.dout(w_dff_B_gvOhazXT0_2),.clk(gclk));
	jdff dff_B_VHcLtPYa1_2(.din(w_dff_B_gvOhazXT0_2),.dout(w_dff_B_VHcLtPYa1_2),.clk(gclk));
	jdff dff_B_KjcNmx9n4_2(.din(w_dff_B_VHcLtPYa1_2),.dout(w_dff_B_KjcNmx9n4_2),.clk(gclk));
	jdff dff_B_OdAHMk085_2(.din(w_dff_B_KjcNmx9n4_2),.dout(w_dff_B_OdAHMk085_2),.clk(gclk));
	jdff dff_B_M08TkCT50_2(.din(w_dff_B_OdAHMk085_2),.dout(w_dff_B_M08TkCT50_2),.clk(gclk));
	jdff dff_B_KudcsrTK9_2(.din(w_dff_B_M08TkCT50_2),.dout(w_dff_B_KudcsrTK9_2),.clk(gclk));
	jdff dff_B_oYaIClRT9_2(.din(w_dff_B_KudcsrTK9_2),.dout(w_dff_B_oYaIClRT9_2),.clk(gclk));
	jdff dff_B_0yQqW5rK6_2(.din(w_dff_B_oYaIClRT9_2),.dout(w_dff_B_0yQqW5rK6_2),.clk(gclk));
	jdff dff_B_4NfDJ9Do6_2(.din(w_dff_B_0yQqW5rK6_2),.dout(w_dff_B_4NfDJ9Do6_2),.clk(gclk));
	jdff dff_B_21AlTdPx9_2(.din(w_dff_B_4NfDJ9Do6_2),.dout(w_dff_B_21AlTdPx9_2),.clk(gclk));
	jdff dff_B_9R50SdT34_2(.din(w_dff_B_21AlTdPx9_2),.dout(w_dff_B_9R50SdT34_2),.clk(gclk));
	jdff dff_B_fNBn6mQi5_2(.din(w_dff_B_9R50SdT34_2),.dout(w_dff_B_fNBn6mQi5_2),.clk(gclk));
	jdff dff_B_eyd7J8PN4_2(.din(w_dff_B_fNBn6mQi5_2),.dout(w_dff_B_eyd7J8PN4_2),.clk(gclk));
	jdff dff_B_mQ9i8Y283_2(.din(w_dff_B_eyd7J8PN4_2),.dout(w_dff_B_mQ9i8Y283_2),.clk(gclk));
	jdff dff_B_Pe5S1Bua7_2(.din(w_dff_B_mQ9i8Y283_2),.dout(w_dff_B_Pe5S1Bua7_2),.clk(gclk));
	jdff dff_B_8GmyEVhh7_2(.din(w_dff_B_Pe5S1Bua7_2),.dout(w_dff_B_8GmyEVhh7_2),.clk(gclk));
	jdff dff_B_KzNRgZlN9_2(.din(w_dff_B_8GmyEVhh7_2),.dout(w_dff_B_KzNRgZlN9_2),.clk(gclk));
	jdff dff_B_debyNz7m6_2(.din(w_dff_B_KzNRgZlN9_2),.dout(w_dff_B_debyNz7m6_2),.clk(gclk));
	jdff dff_B_71sD4LkC3_2(.din(w_dff_B_debyNz7m6_2),.dout(w_dff_B_71sD4LkC3_2),.clk(gclk));
	jdff dff_B_OKLa9Y4w5_2(.din(w_dff_B_71sD4LkC3_2),.dout(w_dff_B_OKLa9Y4w5_2),.clk(gclk));
	jdff dff_B_vAR6gnbU2_2(.din(w_dff_B_OKLa9Y4w5_2),.dout(w_dff_B_vAR6gnbU2_2),.clk(gclk));
	jdff dff_B_SQ2UFCHO7_2(.din(n606),.dout(w_dff_B_SQ2UFCHO7_2),.clk(gclk));
	jdff dff_B_L2nPKQmm2_1(.din(n543),.dout(w_dff_B_L2nPKQmm2_1),.clk(gclk));
	jdff dff_B_c4sq8zqR5_2(.din(n464),.dout(w_dff_B_c4sq8zqR5_2),.clk(gclk));
	jdff dff_B_mOoYf1Jb9_2(.din(w_dff_B_c4sq8zqR5_2),.dout(w_dff_B_mOoYf1Jb9_2),.clk(gclk));
	jdff dff_B_yCZhBPxp8_2(.din(w_dff_B_mOoYf1Jb9_2),.dout(w_dff_B_yCZhBPxp8_2),.clk(gclk));
	jdff dff_B_Mul37upJ9_2(.din(w_dff_B_yCZhBPxp8_2),.dout(w_dff_B_Mul37upJ9_2),.clk(gclk));
	jdff dff_B_Vr2Pzmrc5_2(.din(w_dff_B_Mul37upJ9_2),.dout(w_dff_B_Vr2Pzmrc5_2),.clk(gclk));
	jdff dff_B_qo8HQgrj5_2(.din(w_dff_B_Vr2Pzmrc5_2),.dout(w_dff_B_qo8HQgrj5_2),.clk(gclk));
	jdff dff_B_K3DD2AXb5_2(.din(w_dff_B_qo8HQgrj5_2),.dout(w_dff_B_K3DD2AXb5_2),.clk(gclk));
	jdff dff_B_HZkZjAfV5_2(.din(w_dff_B_K3DD2AXb5_2),.dout(w_dff_B_HZkZjAfV5_2),.clk(gclk));
	jdff dff_B_FH92ztJZ4_2(.din(w_dff_B_HZkZjAfV5_2),.dout(w_dff_B_FH92ztJZ4_2),.clk(gclk));
	jdff dff_B_w8i5aEmS3_2(.din(w_dff_B_FH92ztJZ4_2),.dout(w_dff_B_w8i5aEmS3_2),.clk(gclk));
	jdff dff_B_cjp2gP3k2_2(.din(w_dff_B_w8i5aEmS3_2),.dout(w_dff_B_cjp2gP3k2_2),.clk(gclk));
	jdff dff_B_Z5u0LZ2M7_2(.din(w_dff_B_cjp2gP3k2_2),.dout(w_dff_B_Z5u0LZ2M7_2),.clk(gclk));
	jdff dff_B_XiHaLHLS6_2(.din(w_dff_B_Z5u0LZ2M7_2),.dout(w_dff_B_XiHaLHLS6_2),.clk(gclk));
	jdff dff_B_IXsfg1ad6_2(.din(w_dff_B_XiHaLHLS6_2),.dout(w_dff_B_IXsfg1ad6_2),.clk(gclk));
	jdff dff_B_WaX5XqFb4_2(.din(w_dff_B_IXsfg1ad6_2),.dout(w_dff_B_WaX5XqFb4_2),.clk(gclk));
	jdff dff_B_7Ze0OYxt3_2(.din(w_dff_B_WaX5XqFb4_2),.dout(w_dff_B_7Ze0OYxt3_2),.clk(gclk));
	jdff dff_B_WTlshVem5_2(.din(w_dff_B_7Ze0OYxt3_2),.dout(w_dff_B_WTlshVem5_2),.clk(gclk));
	jdff dff_B_d9wXloB33_2(.din(w_dff_B_WTlshVem5_2),.dout(w_dff_B_d9wXloB33_2),.clk(gclk));
	jdff dff_B_RSoPvPgy5_2(.din(w_dff_B_d9wXloB33_2),.dout(w_dff_B_RSoPvPgy5_2),.clk(gclk));
	jdff dff_B_Xya5hZUY2_2(.din(w_dff_B_RSoPvPgy5_2),.dout(w_dff_B_Xya5hZUY2_2),.clk(gclk));
	jdff dff_B_zqATVwVs3_2(.din(w_dff_B_Xya5hZUY2_2),.dout(w_dff_B_zqATVwVs3_2),.clk(gclk));
	jdff dff_B_Xi5AxfYo5_2(.din(w_dff_B_zqATVwVs3_2),.dout(w_dff_B_Xi5AxfYo5_2),.clk(gclk));
	jdff dff_B_8Nz5cBEq1_2(.din(w_dff_B_Xi5AxfYo5_2),.dout(w_dff_B_8Nz5cBEq1_2),.clk(gclk));
	jdff dff_B_qarWrr7Y9_2(.din(w_dff_B_8Nz5cBEq1_2),.dout(w_dff_B_qarWrr7Y9_2),.clk(gclk));
	jdff dff_B_4CbSZ5vX4_2(.din(n521),.dout(w_dff_B_4CbSZ5vX4_2),.clk(gclk));
	jdff dff_B_X5omvm2U0_1(.din(n465),.dout(w_dff_B_X5omvm2U0_1),.clk(gclk));
	jdff dff_B_FL4oPBb72_2(.din(n393),.dout(w_dff_B_FL4oPBb72_2),.clk(gclk));
	jdff dff_B_LvPyXXkq7_2(.din(w_dff_B_FL4oPBb72_2),.dout(w_dff_B_LvPyXXkq7_2),.clk(gclk));
	jdff dff_B_2bilZ0N25_2(.din(w_dff_B_LvPyXXkq7_2),.dout(w_dff_B_2bilZ0N25_2),.clk(gclk));
	jdff dff_B_ENdoiEJq4_2(.din(w_dff_B_2bilZ0N25_2),.dout(w_dff_B_ENdoiEJq4_2),.clk(gclk));
	jdff dff_B_vese2wvk4_2(.din(w_dff_B_ENdoiEJq4_2),.dout(w_dff_B_vese2wvk4_2),.clk(gclk));
	jdff dff_B_WM4BWJ4s8_2(.din(w_dff_B_vese2wvk4_2),.dout(w_dff_B_WM4BWJ4s8_2),.clk(gclk));
	jdff dff_B_jNlVsGzh4_2(.din(w_dff_B_WM4BWJ4s8_2),.dout(w_dff_B_jNlVsGzh4_2),.clk(gclk));
	jdff dff_B_q0eth2wE1_2(.din(w_dff_B_jNlVsGzh4_2),.dout(w_dff_B_q0eth2wE1_2),.clk(gclk));
	jdff dff_B_WG9DLVO93_2(.din(w_dff_B_q0eth2wE1_2),.dout(w_dff_B_WG9DLVO93_2),.clk(gclk));
	jdff dff_B_FP48xxx35_2(.din(w_dff_B_WG9DLVO93_2),.dout(w_dff_B_FP48xxx35_2),.clk(gclk));
	jdff dff_B_WcOaV3KZ7_2(.din(w_dff_B_FP48xxx35_2),.dout(w_dff_B_WcOaV3KZ7_2),.clk(gclk));
	jdff dff_B_u5k8TSn71_2(.din(w_dff_B_WcOaV3KZ7_2),.dout(w_dff_B_u5k8TSn71_2),.clk(gclk));
	jdff dff_B_c4e9w2VA4_2(.din(w_dff_B_u5k8TSn71_2),.dout(w_dff_B_c4e9w2VA4_2),.clk(gclk));
	jdff dff_B_jXUeBYB18_2(.din(w_dff_B_c4e9w2VA4_2),.dout(w_dff_B_jXUeBYB18_2),.clk(gclk));
	jdff dff_B_hjc6npKu3_2(.din(w_dff_B_jXUeBYB18_2),.dout(w_dff_B_hjc6npKu3_2),.clk(gclk));
	jdff dff_B_TfLbHHsW6_2(.din(w_dff_B_hjc6npKu3_2),.dout(w_dff_B_TfLbHHsW6_2),.clk(gclk));
	jdff dff_B_r5XncUOe1_2(.din(w_dff_B_TfLbHHsW6_2),.dout(w_dff_B_r5XncUOe1_2),.clk(gclk));
	jdff dff_B_byJXfhuc8_2(.din(w_dff_B_r5XncUOe1_2),.dout(w_dff_B_byJXfhuc8_2),.clk(gclk));
	jdff dff_B_j3iwvC752_2(.din(w_dff_B_byJXfhuc8_2),.dout(w_dff_B_j3iwvC752_2),.clk(gclk));
	jdff dff_B_JfxA9DbI9_2(.din(w_dff_B_j3iwvC752_2),.dout(w_dff_B_JfxA9DbI9_2),.clk(gclk));
	jdff dff_B_ym3Zhri70_2(.din(w_dff_B_JfxA9DbI9_2),.dout(w_dff_B_ym3Zhri70_2),.clk(gclk));
	jdff dff_B_zx4XBNOA8_2(.din(n443),.dout(w_dff_B_zx4XBNOA8_2),.clk(gclk));
	jdff dff_B_Bs4DgqRc7_1(.din(n394),.dout(w_dff_B_Bs4DgqRc7_1),.clk(gclk));
	jdff dff_B_eVoHHgMh1_2(.din(n330),.dout(w_dff_B_eVoHHgMh1_2),.clk(gclk));
	jdff dff_B_ifv1llP13_2(.din(w_dff_B_eVoHHgMh1_2),.dout(w_dff_B_ifv1llP13_2),.clk(gclk));
	jdff dff_B_pncGDIyb2_2(.din(w_dff_B_ifv1llP13_2),.dout(w_dff_B_pncGDIyb2_2),.clk(gclk));
	jdff dff_B_dpQYugbH5_2(.din(w_dff_B_pncGDIyb2_2),.dout(w_dff_B_dpQYugbH5_2),.clk(gclk));
	jdff dff_B_sv95vB819_2(.din(w_dff_B_dpQYugbH5_2),.dout(w_dff_B_sv95vB819_2),.clk(gclk));
	jdff dff_B_u2QHBXNp3_2(.din(w_dff_B_sv95vB819_2),.dout(w_dff_B_u2QHBXNp3_2),.clk(gclk));
	jdff dff_B_6xU8DAjM9_2(.din(w_dff_B_u2QHBXNp3_2),.dout(w_dff_B_6xU8DAjM9_2),.clk(gclk));
	jdff dff_B_rVOc4Pvu7_2(.din(w_dff_B_6xU8DAjM9_2),.dout(w_dff_B_rVOc4Pvu7_2),.clk(gclk));
	jdff dff_B_Y867QQsv3_2(.din(w_dff_B_rVOc4Pvu7_2),.dout(w_dff_B_Y867QQsv3_2),.clk(gclk));
	jdff dff_B_IABYL4ue1_2(.din(w_dff_B_Y867QQsv3_2),.dout(w_dff_B_IABYL4ue1_2),.clk(gclk));
	jdff dff_B_aKZmd10S1_2(.din(w_dff_B_IABYL4ue1_2),.dout(w_dff_B_aKZmd10S1_2),.clk(gclk));
	jdff dff_B_P3GWNgdy4_2(.din(w_dff_B_aKZmd10S1_2),.dout(w_dff_B_P3GWNgdy4_2),.clk(gclk));
	jdff dff_B_ptWp9URN8_2(.din(w_dff_B_P3GWNgdy4_2),.dout(w_dff_B_ptWp9URN8_2),.clk(gclk));
	jdff dff_B_Pw44QFse8_2(.din(w_dff_B_ptWp9URN8_2),.dout(w_dff_B_Pw44QFse8_2),.clk(gclk));
	jdff dff_B_nJAi9NUS2_2(.din(w_dff_B_Pw44QFse8_2),.dout(w_dff_B_nJAi9NUS2_2),.clk(gclk));
	jdff dff_B_xgBntN4U4_2(.din(w_dff_B_nJAi9NUS2_2),.dout(w_dff_B_xgBntN4U4_2),.clk(gclk));
	jdff dff_B_UBMDuBur1_2(.din(w_dff_B_xgBntN4U4_2),.dout(w_dff_B_UBMDuBur1_2),.clk(gclk));
	jdff dff_B_GcmFsTjW1_2(.din(w_dff_B_UBMDuBur1_2),.dout(w_dff_B_GcmFsTjW1_2),.clk(gclk));
	jdff dff_B_hTY2G8Qz6_2(.din(n372),.dout(w_dff_B_hTY2G8Qz6_2),.clk(gclk));
	jdff dff_B_XaXDB1un7_1(.din(n331),.dout(w_dff_B_XaXDB1un7_1),.clk(gclk));
	jdff dff_B_3AYx6PUb7_2(.din(n274),.dout(w_dff_B_3AYx6PUb7_2),.clk(gclk));
	jdff dff_B_LQ3iHkdQ4_2(.din(w_dff_B_3AYx6PUb7_2),.dout(w_dff_B_LQ3iHkdQ4_2),.clk(gclk));
	jdff dff_B_H27fDRbF5_2(.din(w_dff_B_LQ3iHkdQ4_2),.dout(w_dff_B_H27fDRbF5_2),.clk(gclk));
	jdff dff_B_nKPtcQ663_2(.din(w_dff_B_H27fDRbF5_2),.dout(w_dff_B_nKPtcQ663_2),.clk(gclk));
	jdff dff_B_TEIh8Wse9_2(.din(w_dff_B_nKPtcQ663_2),.dout(w_dff_B_TEIh8Wse9_2),.clk(gclk));
	jdff dff_B_ktNZMjEI5_2(.din(w_dff_B_TEIh8Wse9_2),.dout(w_dff_B_ktNZMjEI5_2),.clk(gclk));
	jdff dff_B_BeC7EHWL6_2(.din(w_dff_B_ktNZMjEI5_2),.dout(w_dff_B_BeC7EHWL6_2),.clk(gclk));
	jdff dff_B_qJimZa2S7_2(.din(w_dff_B_BeC7EHWL6_2),.dout(w_dff_B_qJimZa2S7_2),.clk(gclk));
	jdff dff_B_Qu8p78dQ7_2(.din(w_dff_B_qJimZa2S7_2),.dout(w_dff_B_Qu8p78dQ7_2),.clk(gclk));
	jdff dff_B_p96mk8IX7_2(.din(w_dff_B_Qu8p78dQ7_2),.dout(w_dff_B_p96mk8IX7_2),.clk(gclk));
	jdff dff_B_VZOo691w6_2(.din(w_dff_B_p96mk8IX7_2),.dout(w_dff_B_VZOo691w6_2),.clk(gclk));
	jdff dff_B_D0bKMrlm2_2(.din(w_dff_B_VZOo691w6_2),.dout(w_dff_B_D0bKMrlm2_2),.clk(gclk));
	jdff dff_B_YHb5QV8n9_2(.din(w_dff_B_D0bKMrlm2_2),.dout(w_dff_B_YHb5QV8n9_2),.clk(gclk));
	jdff dff_B_2eL7hIAR7_2(.din(w_dff_B_YHb5QV8n9_2),.dout(w_dff_B_2eL7hIAR7_2),.clk(gclk));
	jdff dff_B_n0acGMyX6_2(.din(w_dff_B_2eL7hIAR7_2),.dout(w_dff_B_n0acGMyX6_2),.clk(gclk));
	jdff dff_B_MdHYQ9QH5_2(.din(n309),.dout(w_dff_B_MdHYQ9QH5_2),.clk(gclk));
	jdff dff_B_2zdPCp3j5_1(.din(n275),.dout(w_dff_B_2zdPCp3j5_1),.clk(gclk));
	jdff dff_B_fBUYFPWv9_2(.din(n225),.dout(w_dff_B_fBUYFPWv9_2),.clk(gclk));
	jdff dff_B_nLXPnEUn5_2(.din(w_dff_B_fBUYFPWv9_2),.dout(w_dff_B_nLXPnEUn5_2),.clk(gclk));
	jdff dff_B_Lb1EoDNV4_2(.din(w_dff_B_nLXPnEUn5_2),.dout(w_dff_B_Lb1EoDNV4_2),.clk(gclk));
	jdff dff_B_e5TTvIDn2_2(.din(w_dff_B_Lb1EoDNV4_2),.dout(w_dff_B_e5TTvIDn2_2),.clk(gclk));
	jdff dff_B_8xb3SKbj7_2(.din(w_dff_B_e5TTvIDn2_2),.dout(w_dff_B_8xb3SKbj7_2),.clk(gclk));
	jdff dff_B_8pmgmrqv9_2(.din(w_dff_B_8xb3SKbj7_2),.dout(w_dff_B_8pmgmrqv9_2),.clk(gclk));
	jdff dff_B_UUxAbdPb9_2(.din(w_dff_B_8pmgmrqv9_2),.dout(w_dff_B_UUxAbdPb9_2),.clk(gclk));
	jdff dff_B_tH1kPjGu9_2(.din(w_dff_B_UUxAbdPb9_2),.dout(w_dff_B_tH1kPjGu9_2),.clk(gclk));
	jdff dff_B_xiCsUoNt2_2(.din(w_dff_B_tH1kPjGu9_2),.dout(w_dff_B_xiCsUoNt2_2),.clk(gclk));
	jdff dff_B_CzKDmZqK4_2(.din(w_dff_B_xiCsUoNt2_2),.dout(w_dff_B_CzKDmZqK4_2),.clk(gclk));
	jdff dff_B_o71D0EqK8_2(.din(w_dff_B_CzKDmZqK4_2),.dout(w_dff_B_o71D0EqK8_2),.clk(gclk));
	jdff dff_B_lpY4cnop9_2(.din(w_dff_B_o71D0EqK8_2),.dout(w_dff_B_lpY4cnop9_2),.clk(gclk));
	jdff dff_B_u8z9iEiN3_2(.din(n253),.dout(w_dff_B_u8z9iEiN3_2),.clk(gclk));
	jdff dff_B_y8neqvKc3_1(.din(n226),.dout(w_dff_B_y8neqvKc3_1),.clk(gclk));
	jdff dff_B_kyr9crAz3_2(.din(n183),.dout(w_dff_B_kyr9crAz3_2),.clk(gclk));
	jdff dff_B_a1diWAbW8_2(.din(w_dff_B_kyr9crAz3_2),.dout(w_dff_B_a1diWAbW8_2),.clk(gclk));
	jdff dff_B_vWOEN5Am9_2(.din(w_dff_B_a1diWAbW8_2),.dout(w_dff_B_vWOEN5Am9_2),.clk(gclk));
	jdff dff_B_qTCT4rn00_2(.din(w_dff_B_vWOEN5Am9_2),.dout(w_dff_B_qTCT4rn00_2),.clk(gclk));
	jdff dff_B_OV1Rcg7f1_2(.din(w_dff_B_qTCT4rn00_2),.dout(w_dff_B_OV1Rcg7f1_2),.clk(gclk));
	jdff dff_B_jYusxhKz8_2(.din(w_dff_B_OV1Rcg7f1_2),.dout(w_dff_B_jYusxhKz8_2),.clk(gclk));
	jdff dff_B_OOlb4gtb7_2(.din(w_dff_B_jYusxhKz8_2),.dout(w_dff_B_OOlb4gtb7_2),.clk(gclk));
	jdff dff_B_p6zTNLbH6_2(.din(w_dff_B_OOlb4gtb7_2),.dout(w_dff_B_p6zTNLbH6_2),.clk(gclk));
	jdff dff_B_RQbxMgue5_2(.din(w_dff_B_p6zTNLbH6_2),.dout(w_dff_B_RQbxMgue5_2),.clk(gclk));
	jdff dff_B_YSaWgmih5_2(.din(n204),.dout(w_dff_B_YSaWgmih5_2),.clk(gclk));
	jdff dff_B_Ahgr0w2R0_1(.din(n184),.dout(w_dff_B_Ahgr0w2R0_1),.clk(gclk));
	jdff dff_B_f3hDQk3h4_2(.din(n148),.dout(w_dff_B_f3hDQk3h4_2),.clk(gclk));
	jdff dff_B_zeCKEgXy2_2(.din(w_dff_B_f3hDQk3h4_2),.dout(w_dff_B_zeCKEgXy2_2),.clk(gclk));
	jdff dff_B_ds9YZXoq9_2(.din(w_dff_B_zeCKEgXy2_2),.dout(w_dff_B_ds9YZXoq9_2),.clk(gclk));
	jdff dff_B_aeIqsUPX2_2(.din(w_dff_B_ds9YZXoq9_2),.dout(w_dff_B_aeIqsUPX2_2),.clk(gclk));
	jdff dff_B_b74r9Gi62_2(.din(w_dff_B_aeIqsUPX2_2),.dout(w_dff_B_b74r9Gi62_2),.clk(gclk));
	jdff dff_B_GKEotS8a1_2(.din(w_dff_B_b74r9Gi62_2),.dout(w_dff_B_GKEotS8a1_2),.clk(gclk));
	jdff dff_B_3qcV8KCs4_2(.din(n162),.dout(w_dff_B_3qcV8KCs4_2),.clk(gclk));
	jdff dff_B_aPUqMr1Q7_2(.din(n119),.dout(w_dff_B_aPUqMr1Q7_2),.clk(gclk));
	jdff dff_B_RrCKCGtT2_2(.din(w_dff_B_aPUqMr1Q7_2),.dout(w_dff_B_RrCKCGtT2_2),.clk(gclk));
	jdff dff_B_SKjCMl7v6_2(.din(w_dff_B_RrCKCGtT2_2),.dout(w_dff_B_SKjCMl7v6_2),.clk(gclk));
	jdff dff_B_Vp1e94050_0(.din(n126),.dout(w_dff_B_Vp1e94050_0),.clk(gclk));
	jdff dff_B_eXsPARqE7_0(.din(n1298),.dout(w_dff_B_eXsPARqE7_0),.clk(gclk));
	jdff dff_A_DlOdnnnI0_1(.dout(w_n1294_0[1]),.din(w_dff_A_DlOdnnnI0_1),.clk(gclk));
	jdff dff_A_SO1P2mKd0_1(.dout(w_dff_A_DlOdnnnI0_1),.din(w_dff_A_SO1P2mKd0_1),.clk(gclk));
	jdff dff_B_P9F6kZrV9_1(.din(n1214),.dout(w_dff_B_P9F6kZrV9_1),.clk(gclk));
	jdff dff_B_oqfRcZfn8_1(.din(w_dff_B_P9F6kZrV9_1),.dout(w_dff_B_oqfRcZfn8_1),.clk(gclk));
	jdff dff_B_EVVFRqZg9_2(.din(n1120),.dout(w_dff_B_EVVFRqZg9_2),.clk(gclk));
	jdff dff_B_awF2P6AN6_2(.din(w_dff_B_EVVFRqZg9_2),.dout(w_dff_B_awF2P6AN6_2),.clk(gclk));
	jdff dff_B_8EQXT19O0_2(.din(w_dff_B_awF2P6AN6_2),.dout(w_dff_B_8EQXT19O0_2),.clk(gclk));
	jdff dff_B_DfazqAdr5_2(.din(w_dff_B_8EQXT19O0_2),.dout(w_dff_B_DfazqAdr5_2),.clk(gclk));
	jdff dff_B_e4opkjwI4_2(.din(w_dff_B_DfazqAdr5_2),.dout(w_dff_B_e4opkjwI4_2),.clk(gclk));
	jdff dff_B_2am6qQWW5_2(.din(w_dff_B_e4opkjwI4_2),.dout(w_dff_B_2am6qQWW5_2),.clk(gclk));
	jdff dff_B_ADZmoE0x3_2(.din(w_dff_B_2am6qQWW5_2),.dout(w_dff_B_ADZmoE0x3_2),.clk(gclk));
	jdff dff_B_rRFl05J20_2(.din(w_dff_B_ADZmoE0x3_2),.dout(w_dff_B_rRFl05J20_2),.clk(gclk));
	jdff dff_B_Etxsq8lX1_2(.din(w_dff_B_rRFl05J20_2),.dout(w_dff_B_Etxsq8lX1_2),.clk(gclk));
	jdff dff_B_bdHEFPg50_2(.din(w_dff_B_Etxsq8lX1_2),.dout(w_dff_B_bdHEFPg50_2),.clk(gclk));
	jdff dff_B_WkyDX7Ym8_2(.din(w_dff_B_bdHEFPg50_2),.dout(w_dff_B_WkyDX7Ym8_2),.clk(gclk));
	jdff dff_B_VxLzf2U09_2(.din(w_dff_B_WkyDX7Ym8_2),.dout(w_dff_B_VxLzf2U09_2),.clk(gclk));
	jdff dff_B_0Op7r6oD3_2(.din(w_dff_B_VxLzf2U09_2),.dout(w_dff_B_0Op7r6oD3_2),.clk(gclk));
	jdff dff_B_aOsRYIrX9_2(.din(w_dff_B_0Op7r6oD3_2),.dout(w_dff_B_aOsRYIrX9_2),.clk(gclk));
	jdff dff_B_QkMcCj3B1_2(.din(w_dff_B_aOsRYIrX9_2),.dout(w_dff_B_QkMcCj3B1_2),.clk(gclk));
	jdff dff_B_43t4PVte6_2(.din(w_dff_B_QkMcCj3B1_2),.dout(w_dff_B_43t4PVte6_2),.clk(gclk));
	jdff dff_B_OT7JCWRn5_2(.din(w_dff_B_43t4PVte6_2),.dout(w_dff_B_OT7JCWRn5_2),.clk(gclk));
	jdff dff_B_YDaXchOg2_2(.din(w_dff_B_OT7JCWRn5_2),.dout(w_dff_B_YDaXchOg2_2),.clk(gclk));
	jdff dff_B_wgCOrgMY7_2(.din(w_dff_B_YDaXchOg2_2),.dout(w_dff_B_wgCOrgMY7_2),.clk(gclk));
	jdff dff_B_RhUz6OvF2_2(.din(w_dff_B_wgCOrgMY7_2),.dout(w_dff_B_RhUz6OvF2_2),.clk(gclk));
	jdff dff_B_2MlIBitM5_2(.din(w_dff_B_RhUz6OvF2_2),.dout(w_dff_B_2MlIBitM5_2),.clk(gclk));
	jdff dff_B_2VF38Yei9_2(.din(w_dff_B_2MlIBitM5_2),.dout(w_dff_B_2VF38Yei9_2),.clk(gclk));
	jdff dff_B_RgLwhXgw5_2(.din(w_dff_B_2VF38Yei9_2),.dout(w_dff_B_RgLwhXgw5_2),.clk(gclk));
	jdff dff_B_WjSiQqSf8_2(.din(w_dff_B_RgLwhXgw5_2),.dout(w_dff_B_WjSiQqSf8_2),.clk(gclk));
	jdff dff_B_2TAtEa473_2(.din(w_dff_B_WjSiQqSf8_2),.dout(w_dff_B_2TAtEa473_2),.clk(gclk));
	jdff dff_B_TsjUJFQZ1_2(.din(w_dff_B_2TAtEa473_2),.dout(w_dff_B_TsjUJFQZ1_2),.clk(gclk));
	jdff dff_B_D0KO3jPT7_2(.din(w_dff_B_TsjUJFQZ1_2),.dout(w_dff_B_D0KO3jPT7_2),.clk(gclk));
	jdff dff_B_Gm9f3XRR9_2(.din(w_dff_B_D0KO3jPT7_2),.dout(w_dff_B_Gm9f3XRR9_2),.clk(gclk));
	jdff dff_B_293qiK9z6_2(.din(w_dff_B_Gm9f3XRR9_2),.dout(w_dff_B_293qiK9z6_2),.clk(gclk));
	jdff dff_B_mvUxN0mq1_2(.din(w_dff_B_293qiK9z6_2),.dout(w_dff_B_mvUxN0mq1_2),.clk(gclk));
	jdff dff_B_SOCLBoWa4_2(.din(w_dff_B_mvUxN0mq1_2),.dout(w_dff_B_SOCLBoWa4_2),.clk(gclk));
	jdff dff_B_oKEjuQty0_2(.din(w_dff_B_SOCLBoWa4_2),.dout(w_dff_B_oKEjuQty0_2),.clk(gclk));
	jdff dff_B_ayF3F6j89_2(.din(w_dff_B_oKEjuQty0_2),.dout(w_dff_B_ayF3F6j89_2),.clk(gclk));
	jdff dff_B_fpGvMBxt1_2(.din(w_dff_B_ayF3F6j89_2),.dout(w_dff_B_fpGvMBxt1_2),.clk(gclk));
	jdff dff_B_NX1yYp398_2(.din(w_dff_B_fpGvMBxt1_2),.dout(w_dff_B_NX1yYp398_2),.clk(gclk));
	jdff dff_B_u3FVPYPI5_2(.din(w_dff_B_NX1yYp398_2),.dout(w_dff_B_u3FVPYPI5_2),.clk(gclk));
	jdff dff_B_Y5CJJox81_2(.din(w_dff_B_u3FVPYPI5_2),.dout(w_dff_B_Y5CJJox81_2),.clk(gclk));
	jdff dff_B_8eo7xoXf6_2(.din(w_dff_B_Y5CJJox81_2),.dout(w_dff_B_8eo7xoXf6_2),.clk(gclk));
	jdff dff_B_qISSE5J91_2(.din(w_dff_B_8eo7xoXf6_2),.dout(w_dff_B_qISSE5J91_2),.clk(gclk));
	jdff dff_B_LEndyedm0_2(.din(w_dff_B_qISSE5J91_2),.dout(w_dff_B_LEndyedm0_2),.clk(gclk));
	jdff dff_B_oyWtLiPE7_2(.din(w_dff_B_LEndyedm0_2),.dout(w_dff_B_oyWtLiPE7_2),.clk(gclk));
	jdff dff_B_fiNWfDKF5_2(.din(w_dff_B_oyWtLiPE7_2),.dout(w_dff_B_fiNWfDKF5_2),.clk(gclk));
	jdff dff_B_6HkBwK4T1_2(.din(w_dff_B_fiNWfDKF5_2),.dout(w_dff_B_6HkBwK4T1_2),.clk(gclk));
	jdff dff_B_nzO81hGf5_2(.din(w_dff_B_6HkBwK4T1_2),.dout(w_dff_B_nzO81hGf5_2),.clk(gclk));
	jdff dff_B_k6qpMpUd0_2(.din(w_dff_B_nzO81hGf5_2),.dout(w_dff_B_k6qpMpUd0_2),.clk(gclk));
	jdff dff_B_5rgbaAfY4_2(.din(n1203),.dout(w_dff_B_5rgbaAfY4_2),.clk(gclk));
	jdff dff_B_2agerOhh0_1(.din(n1122),.dout(w_dff_B_2agerOhh0_1),.clk(gclk));
	jdff dff_B_plRlcrQy1_2(.din(n1023),.dout(w_dff_B_plRlcrQy1_2),.clk(gclk));
	jdff dff_B_XHyuMrUU8_2(.din(w_dff_B_plRlcrQy1_2),.dout(w_dff_B_XHyuMrUU8_2),.clk(gclk));
	jdff dff_B_xRCoA3tL9_2(.din(w_dff_B_XHyuMrUU8_2),.dout(w_dff_B_xRCoA3tL9_2),.clk(gclk));
	jdff dff_B_bgdDR2Tq7_2(.din(w_dff_B_xRCoA3tL9_2),.dout(w_dff_B_bgdDR2Tq7_2),.clk(gclk));
	jdff dff_B_o8xBbSY07_2(.din(w_dff_B_bgdDR2Tq7_2),.dout(w_dff_B_o8xBbSY07_2),.clk(gclk));
	jdff dff_B_BppLBu097_2(.din(w_dff_B_o8xBbSY07_2),.dout(w_dff_B_BppLBu097_2),.clk(gclk));
	jdff dff_B_w7DjH2Zj6_2(.din(w_dff_B_BppLBu097_2),.dout(w_dff_B_w7DjH2Zj6_2),.clk(gclk));
	jdff dff_B_GwUYymFD8_2(.din(w_dff_B_w7DjH2Zj6_2),.dout(w_dff_B_GwUYymFD8_2),.clk(gclk));
	jdff dff_B_NLaVXcXC1_2(.din(w_dff_B_GwUYymFD8_2),.dout(w_dff_B_NLaVXcXC1_2),.clk(gclk));
	jdff dff_B_CvXsLa9q4_2(.din(w_dff_B_NLaVXcXC1_2),.dout(w_dff_B_CvXsLa9q4_2),.clk(gclk));
	jdff dff_B_aWKAKEWC6_2(.din(w_dff_B_CvXsLa9q4_2),.dout(w_dff_B_aWKAKEWC6_2),.clk(gclk));
	jdff dff_B_PCkpH6ki9_2(.din(w_dff_B_aWKAKEWC6_2),.dout(w_dff_B_PCkpH6ki9_2),.clk(gclk));
	jdff dff_B_IjzZGE777_2(.din(w_dff_B_PCkpH6ki9_2),.dout(w_dff_B_IjzZGE777_2),.clk(gclk));
	jdff dff_B_vwlhKaln2_2(.din(w_dff_B_IjzZGE777_2),.dout(w_dff_B_vwlhKaln2_2),.clk(gclk));
	jdff dff_B_4r9cV33p6_2(.din(w_dff_B_vwlhKaln2_2),.dout(w_dff_B_4r9cV33p6_2),.clk(gclk));
	jdff dff_B_bcFjwpJ61_2(.din(w_dff_B_4r9cV33p6_2),.dout(w_dff_B_bcFjwpJ61_2),.clk(gclk));
	jdff dff_B_g1QVrJ7F6_2(.din(w_dff_B_bcFjwpJ61_2),.dout(w_dff_B_g1QVrJ7F6_2),.clk(gclk));
	jdff dff_B_UqJogqPs6_2(.din(w_dff_B_g1QVrJ7F6_2),.dout(w_dff_B_UqJogqPs6_2),.clk(gclk));
	jdff dff_B_mqTMNk6f9_2(.din(w_dff_B_UqJogqPs6_2),.dout(w_dff_B_mqTMNk6f9_2),.clk(gclk));
	jdff dff_B_WRGjUugp9_2(.din(w_dff_B_mqTMNk6f9_2),.dout(w_dff_B_WRGjUugp9_2),.clk(gclk));
	jdff dff_B_R0w3avMd0_2(.din(w_dff_B_WRGjUugp9_2),.dout(w_dff_B_R0w3avMd0_2),.clk(gclk));
	jdff dff_B_NpBR11xX4_2(.din(w_dff_B_R0w3avMd0_2),.dout(w_dff_B_NpBR11xX4_2),.clk(gclk));
	jdff dff_B_VUN5HsKF1_2(.din(w_dff_B_NpBR11xX4_2),.dout(w_dff_B_VUN5HsKF1_2),.clk(gclk));
	jdff dff_B_HFrn3sbE3_2(.din(w_dff_B_VUN5HsKF1_2),.dout(w_dff_B_HFrn3sbE3_2),.clk(gclk));
	jdff dff_B_xXFSDG067_2(.din(w_dff_B_HFrn3sbE3_2),.dout(w_dff_B_xXFSDG067_2),.clk(gclk));
	jdff dff_B_sypxpxNa8_2(.din(w_dff_B_xXFSDG067_2),.dout(w_dff_B_sypxpxNa8_2),.clk(gclk));
	jdff dff_B_SVqo9Ppz3_2(.din(w_dff_B_sypxpxNa8_2),.dout(w_dff_B_SVqo9Ppz3_2),.clk(gclk));
	jdff dff_B_YnURCieT3_2(.din(w_dff_B_SVqo9Ppz3_2),.dout(w_dff_B_YnURCieT3_2),.clk(gclk));
	jdff dff_B_CZqbhFpD0_2(.din(w_dff_B_YnURCieT3_2),.dout(w_dff_B_CZqbhFpD0_2),.clk(gclk));
	jdff dff_B_3qa0X0CI2_2(.din(w_dff_B_CZqbhFpD0_2),.dout(w_dff_B_3qa0X0CI2_2),.clk(gclk));
	jdff dff_B_xjHt7fKf4_2(.din(w_dff_B_3qa0X0CI2_2),.dout(w_dff_B_xjHt7fKf4_2),.clk(gclk));
	jdff dff_B_BQP1rre78_2(.din(w_dff_B_xjHt7fKf4_2),.dout(w_dff_B_BQP1rre78_2),.clk(gclk));
	jdff dff_B_l59G6I9D3_2(.din(w_dff_B_BQP1rre78_2),.dout(w_dff_B_l59G6I9D3_2),.clk(gclk));
	jdff dff_B_bKRVCC3o7_2(.din(w_dff_B_l59G6I9D3_2),.dout(w_dff_B_bKRVCC3o7_2),.clk(gclk));
	jdff dff_B_pey6Gaoz4_2(.din(w_dff_B_bKRVCC3o7_2),.dout(w_dff_B_pey6Gaoz4_2),.clk(gclk));
	jdff dff_B_XvTtMi7d7_2(.din(w_dff_B_pey6Gaoz4_2),.dout(w_dff_B_XvTtMi7d7_2),.clk(gclk));
	jdff dff_B_R1QsuEeq6_2(.din(w_dff_B_XvTtMi7d7_2),.dout(w_dff_B_R1QsuEeq6_2),.clk(gclk));
	jdff dff_B_9Mpx2Jkw4_2(.din(w_dff_B_R1QsuEeq6_2),.dout(w_dff_B_9Mpx2Jkw4_2),.clk(gclk));
	jdff dff_B_X7HNuwVK1_2(.din(w_dff_B_9Mpx2Jkw4_2),.dout(w_dff_B_X7HNuwVK1_2),.clk(gclk));
	jdff dff_B_osmQoWUC6_2(.din(w_dff_B_X7HNuwVK1_2),.dout(w_dff_B_osmQoWUC6_2),.clk(gclk));
	jdff dff_B_zeGKJ73x9_2(.din(w_dff_B_osmQoWUC6_2),.dout(w_dff_B_zeGKJ73x9_2),.clk(gclk));
	jdff dff_B_SP7NRKBw2_2(.din(n1103),.dout(w_dff_B_SP7NRKBw2_2),.clk(gclk));
	jdff dff_B_JZOAAh0m7_1(.din(n1024),.dout(w_dff_B_JZOAAh0m7_1),.clk(gclk));
	jdff dff_B_SfGCj1NX8_2(.din(n924),.dout(w_dff_B_SfGCj1NX8_2),.clk(gclk));
	jdff dff_B_BKn5tQhV2_2(.din(w_dff_B_SfGCj1NX8_2),.dout(w_dff_B_BKn5tQhV2_2),.clk(gclk));
	jdff dff_B_z8sYq6UD6_2(.din(w_dff_B_BKn5tQhV2_2),.dout(w_dff_B_z8sYq6UD6_2),.clk(gclk));
	jdff dff_B_K5y0Uywy1_2(.din(w_dff_B_z8sYq6UD6_2),.dout(w_dff_B_K5y0Uywy1_2),.clk(gclk));
	jdff dff_B_yEYlMSue0_2(.din(w_dff_B_K5y0Uywy1_2),.dout(w_dff_B_yEYlMSue0_2),.clk(gclk));
	jdff dff_B_Y37g2gjH6_2(.din(w_dff_B_yEYlMSue0_2),.dout(w_dff_B_Y37g2gjH6_2),.clk(gclk));
	jdff dff_B_kbGAFFd82_2(.din(w_dff_B_Y37g2gjH6_2),.dout(w_dff_B_kbGAFFd82_2),.clk(gclk));
	jdff dff_B_jV8hqtSE5_2(.din(w_dff_B_kbGAFFd82_2),.dout(w_dff_B_jV8hqtSE5_2),.clk(gclk));
	jdff dff_B_qmC5z9LQ6_2(.din(w_dff_B_jV8hqtSE5_2),.dout(w_dff_B_qmC5z9LQ6_2),.clk(gclk));
	jdff dff_B_VXvuDzya9_2(.din(w_dff_B_qmC5z9LQ6_2),.dout(w_dff_B_VXvuDzya9_2),.clk(gclk));
	jdff dff_B_aYTOhepd7_2(.din(w_dff_B_VXvuDzya9_2),.dout(w_dff_B_aYTOhepd7_2),.clk(gclk));
	jdff dff_B_eFbGPJ9D4_2(.din(w_dff_B_aYTOhepd7_2),.dout(w_dff_B_eFbGPJ9D4_2),.clk(gclk));
	jdff dff_B_xJpviDem3_2(.din(w_dff_B_eFbGPJ9D4_2),.dout(w_dff_B_xJpviDem3_2),.clk(gclk));
	jdff dff_B_FsBFaBbz5_2(.din(w_dff_B_xJpviDem3_2),.dout(w_dff_B_FsBFaBbz5_2),.clk(gclk));
	jdff dff_B_3emKv7rM0_2(.din(w_dff_B_FsBFaBbz5_2),.dout(w_dff_B_3emKv7rM0_2),.clk(gclk));
	jdff dff_B_XC3gfv0r1_2(.din(w_dff_B_3emKv7rM0_2),.dout(w_dff_B_XC3gfv0r1_2),.clk(gclk));
	jdff dff_B_rMrBkCUc2_2(.din(w_dff_B_XC3gfv0r1_2),.dout(w_dff_B_rMrBkCUc2_2),.clk(gclk));
	jdff dff_B_BtrmtMzp4_2(.din(w_dff_B_rMrBkCUc2_2),.dout(w_dff_B_BtrmtMzp4_2),.clk(gclk));
	jdff dff_B_B1JvIKgZ8_2(.din(w_dff_B_BtrmtMzp4_2),.dout(w_dff_B_B1JvIKgZ8_2),.clk(gclk));
	jdff dff_B_UxY7OPnX1_2(.din(w_dff_B_B1JvIKgZ8_2),.dout(w_dff_B_UxY7OPnX1_2),.clk(gclk));
	jdff dff_B_pPFbDXp40_2(.din(w_dff_B_UxY7OPnX1_2),.dout(w_dff_B_pPFbDXp40_2),.clk(gclk));
	jdff dff_B_3UVQFIHO7_2(.din(w_dff_B_pPFbDXp40_2),.dout(w_dff_B_3UVQFIHO7_2),.clk(gclk));
	jdff dff_B_4Zi5bA0R3_2(.din(w_dff_B_3UVQFIHO7_2),.dout(w_dff_B_4Zi5bA0R3_2),.clk(gclk));
	jdff dff_B_xJY3JMIk0_2(.din(w_dff_B_4Zi5bA0R3_2),.dout(w_dff_B_xJY3JMIk0_2),.clk(gclk));
	jdff dff_B_o4TAkCq11_2(.din(w_dff_B_xJY3JMIk0_2),.dout(w_dff_B_o4TAkCq11_2),.clk(gclk));
	jdff dff_B_nBtW83Wj8_2(.din(w_dff_B_o4TAkCq11_2),.dout(w_dff_B_nBtW83Wj8_2),.clk(gclk));
	jdff dff_B_yrFlx6x65_2(.din(w_dff_B_nBtW83Wj8_2),.dout(w_dff_B_yrFlx6x65_2),.clk(gclk));
	jdff dff_B_odXFmtme4_2(.din(w_dff_B_yrFlx6x65_2),.dout(w_dff_B_odXFmtme4_2),.clk(gclk));
	jdff dff_B_xkzBdazl2_2(.din(w_dff_B_odXFmtme4_2),.dout(w_dff_B_xkzBdazl2_2),.clk(gclk));
	jdff dff_B_Uv6GYbcM8_2(.din(w_dff_B_xkzBdazl2_2),.dout(w_dff_B_Uv6GYbcM8_2),.clk(gclk));
	jdff dff_B_CHfjPQzu2_2(.din(w_dff_B_Uv6GYbcM8_2),.dout(w_dff_B_CHfjPQzu2_2),.clk(gclk));
	jdff dff_B_abwMh0ZC7_2(.din(w_dff_B_CHfjPQzu2_2),.dout(w_dff_B_abwMh0ZC7_2),.clk(gclk));
	jdff dff_B_2NZmxyyc6_2(.din(w_dff_B_abwMh0ZC7_2),.dout(w_dff_B_2NZmxyyc6_2),.clk(gclk));
	jdff dff_B_tnnsRXoL7_2(.din(w_dff_B_2NZmxyyc6_2),.dout(w_dff_B_tnnsRXoL7_2),.clk(gclk));
	jdff dff_B_NeNp9QR70_2(.din(w_dff_B_tnnsRXoL7_2),.dout(w_dff_B_NeNp9QR70_2),.clk(gclk));
	jdff dff_B_tA00dRxH2_2(.din(w_dff_B_NeNp9QR70_2),.dout(w_dff_B_tA00dRxH2_2),.clk(gclk));
	jdff dff_B_zPu8CIsz0_2(.din(n1004),.dout(w_dff_B_zPu8CIsz0_2),.clk(gclk));
	jdff dff_B_tWfpopR90_1(.din(n925),.dout(w_dff_B_tWfpopR90_1),.clk(gclk));
	jdff dff_B_5xmqKnFL5_2(.din(n822),.dout(w_dff_B_5xmqKnFL5_2),.clk(gclk));
	jdff dff_B_ZZbxtirt1_2(.din(w_dff_B_5xmqKnFL5_2),.dout(w_dff_B_ZZbxtirt1_2),.clk(gclk));
	jdff dff_B_9R46VbSd3_2(.din(w_dff_B_ZZbxtirt1_2),.dout(w_dff_B_9R46VbSd3_2),.clk(gclk));
	jdff dff_B_4qQeQjl38_2(.din(w_dff_B_9R46VbSd3_2),.dout(w_dff_B_4qQeQjl38_2),.clk(gclk));
	jdff dff_B_idy0wPN87_2(.din(w_dff_B_4qQeQjl38_2),.dout(w_dff_B_idy0wPN87_2),.clk(gclk));
	jdff dff_B_1m2z7O3Y4_2(.din(w_dff_B_idy0wPN87_2),.dout(w_dff_B_1m2z7O3Y4_2),.clk(gclk));
	jdff dff_B_OUWuT4dg8_2(.din(w_dff_B_1m2z7O3Y4_2),.dout(w_dff_B_OUWuT4dg8_2),.clk(gclk));
	jdff dff_B_Tmf8wHcL6_2(.din(w_dff_B_OUWuT4dg8_2),.dout(w_dff_B_Tmf8wHcL6_2),.clk(gclk));
	jdff dff_B_fOpeZru06_2(.din(w_dff_B_Tmf8wHcL6_2),.dout(w_dff_B_fOpeZru06_2),.clk(gclk));
	jdff dff_B_95d57tZi2_2(.din(w_dff_B_fOpeZru06_2),.dout(w_dff_B_95d57tZi2_2),.clk(gclk));
	jdff dff_B_CdyXRYiv6_2(.din(w_dff_B_95d57tZi2_2),.dout(w_dff_B_CdyXRYiv6_2),.clk(gclk));
	jdff dff_B_2a3lZlvX8_2(.din(w_dff_B_CdyXRYiv6_2),.dout(w_dff_B_2a3lZlvX8_2),.clk(gclk));
	jdff dff_B_UCKJ8daa0_2(.din(w_dff_B_2a3lZlvX8_2),.dout(w_dff_B_UCKJ8daa0_2),.clk(gclk));
	jdff dff_B_k40dRXGm8_2(.din(w_dff_B_UCKJ8daa0_2),.dout(w_dff_B_k40dRXGm8_2),.clk(gclk));
	jdff dff_B_5G0zsCcN3_2(.din(w_dff_B_k40dRXGm8_2),.dout(w_dff_B_5G0zsCcN3_2),.clk(gclk));
	jdff dff_B_o4Hb9KNs8_2(.din(w_dff_B_5G0zsCcN3_2),.dout(w_dff_B_o4Hb9KNs8_2),.clk(gclk));
	jdff dff_B_m9ajCnLM7_2(.din(w_dff_B_o4Hb9KNs8_2),.dout(w_dff_B_m9ajCnLM7_2),.clk(gclk));
	jdff dff_B_o2RQk1c75_2(.din(w_dff_B_m9ajCnLM7_2),.dout(w_dff_B_o2RQk1c75_2),.clk(gclk));
	jdff dff_B_jWFOf66m4_2(.din(w_dff_B_o2RQk1c75_2),.dout(w_dff_B_jWFOf66m4_2),.clk(gclk));
	jdff dff_B_CZszh0S51_2(.din(w_dff_B_jWFOf66m4_2),.dout(w_dff_B_CZszh0S51_2),.clk(gclk));
	jdff dff_B_RgbMZKsJ8_2(.din(w_dff_B_CZszh0S51_2),.dout(w_dff_B_RgbMZKsJ8_2),.clk(gclk));
	jdff dff_B_sOV6mkJm6_2(.din(w_dff_B_RgbMZKsJ8_2),.dout(w_dff_B_sOV6mkJm6_2),.clk(gclk));
	jdff dff_B_ZxU2XHPK0_2(.din(w_dff_B_sOV6mkJm6_2),.dout(w_dff_B_ZxU2XHPK0_2),.clk(gclk));
	jdff dff_B_izXJIk7T0_2(.din(w_dff_B_ZxU2XHPK0_2),.dout(w_dff_B_izXJIk7T0_2),.clk(gclk));
	jdff dff_B_YAhRNZkW1_2(.din(w_dff_B_izXJIk7T0_2),.dout(w_dff_B_YAhRNZkW1_2),.clk(gclk));
	jdff dff_B_Ct9c1h916_2(.din(w_dff_B_YAhRNZkW1_2),.dout(w_dff_B_Ct9c1h916_2),.clk(gclk));
	jdff dff_B_JxsqKyAW5_2(.din(w_dff_B_Ct9c1h916_2),.dout(w_dff_B_JxsqKyAW5_2),.clk(gclk));
	jdff dff_B_t1XGfg2G0_2(.din(w_dff_B_JxsqKyAW5_2),.dout(w_dff_B_t1XGfg2G0_2),.clk(gclk));
	jdff dff_B_FDFs0Ajd6_2(.din(w_dff_B_t1XGfg2G0_2),.dout(w_dff_B_FDFs0Ajd6_2),.clk(gclk));
	jdff dff_B_diqJhKW81_2(.din(w_dff_B_FDFs0Ajd6_2),.dout(w_dff_B_diqJhKW81_2),.clk(gclk));
	jdff dff_B_bb24lChW1_2(.din(w_dff_B_diqJhKW81_2),.dout(w_dff_B_bb24lChW1_2),.clk(gclk));
	jdff dff_B_nbpakffp1_2(.din(w_dff_B_bb24lChW1_2),.dout(w_dff_B_nbpakffp1_2),.clk(gclk));
	jdff dff_B_3JPXeLls3_2(.din(w_dff_B_nbpakffp1_2),.dout(w_dff_B_3JPXeLls3_2),.clk(gclk));
	jdff dff_B_8iCog5Rp9_2(.din(n898),.dout(w_dff_B_8iCog5Rp9_2),.clk(gclk));
	jdff dff_B_BysUlr9y6_1(.din(n823),.dout(w_dff_B_BysUlr9y6_1),.clk(gclk));
	jdff dff_B_qz2j93Cu9_2(.din(n724),.dout(w_dff_B_qz2j93Cu9_2),.clk(gclk));
	jdff dff_B_pzVR9Z3b0_2(.din(w_dff_B_qz2j93Cu9_2),.dout(w_dff_B_pzVR9Z3b0_2),.clk(gclk));
	jdff dff_B_RFuSuZLs4_2(.din(w_dff_B_pzVR9Z3b0_2),.dout(w_dff_B_RFuSuZLs4_2),.clk(gclk));
	jdff dff_B_VPhVP4Xt9_2(.din(w_dff_B_RFuSuZLs4_2),.dout(w_dff_B_VPhVP4Xt9_2),.clk(gclk));
	jdff dff_B_MxhLVDQj8_2(.din(w_dff_B_VPhVP4Xt9_2),.dout(w_dff_B_MxhLVDQj8_2),.clk(gclk));
	jdff dff_B_2LXPNHTf1_2(.din(w_dff_B_MxhLVDQj8_2),.dout(w_dff_B_2LXPNHTf1_2),.clk(gclk));
	jdff dff_B_yXpl13D91_2(.din(w_dff_B_2LXPNHTf1_2),.dout(w_dff_B_yXpl13D91_2),.clk(gclk));
	jdff dff_B_cX3mh0TA6_2(.din(w_dff_B_yXpl13D91_2),.dout(w_dff_B_cX3mh0TA6_2),.clk(gclk));
	jdff dff_B_HcaSunOj6_2(.din(w_dff_B_cX3mh0TA6_2),.dout(w_dff_B_HcaSunOj6_2),.clk(gclk));
	jdff dff_B_iS1G2Wt26_2(.din(w_dff_B_HcaSunOj6_2),.dout(w_dff_B_iS1G2Wt26_2),.clk(gclk));
	jdff dff_B_OuvjgAH26_2(.din(w_dff_B_iS1G2Wt26_2),.dout(w_dff_B_OuvjgAH26_2),.clk(gclk));
	jdff dff_B_gJfVkYUi5_2(.din(w_dff_B_OuvjgAH26_2),.dout(w_dff_B_gJfVkYUi5_2),.clk(gclk));
	jdff dff_B_w3JLBf8L0_2(.din(w_dff_B_gJfVkYUi5_2),.dout(w_dff_B_w3JLBf8L0_2),.clk(gclk));
	jdff dff_B_uvdapXKf3_2(.din(w_dff_B_w3JLBf8L0_2),.dout(w_dff_B_uvdapXKf3_2),.clk(gclk));
	jdff dff_B_mB0mnk9N8_2(.din(w_dff_B_uvdapXKf3_2),.dout(w_dff_B_mB0mnk9N8_2),.clk(gclk));
	jdff dff_B_XObe7jZ28_2(.din(w_dff_B_mB0mnk9N8_2),.dout(w_dff_B_XObe7jZ28_2),.clk(gclk));
	jdff dff_B_VzGhWh159_2(.din(w_dff_B_XObe7jZ28_2),.dout(w_dff_B_VzGhWh159_2),.clk(gclk));
	jdff dff_B_dSok3YC12_2(.din(w_dff_B_VzGhWh159_2),.dout(w_dff_B_dSok3YC12_2),.clk(gclk));
	jdff dff_B_ZOD1UMvF8_2(.din(w_dff_B_dSok3YC12_2),.dout(w_dff_B_ZOD1UMvF8_2),.clk(gclk));
	jdff dff_B_uIlMGlyK7_2(.din(w_dff_B_ZOD1UMvF8_2),.dout(w_dff_B_uIlMGlyK7_2),.clk(gclk));
	jdff dff_B_q5hiiK7n0_2(.din(w_dff_B_uIlMGlyK7_2),.dout(w_dff_B_q5hiiK7n0_2),.clk(gclk));
	jdff dff_B_1rXs8uF41_2(.din(w_dff_B_q5hiiK7n0_2),.dout(w_dff_B_1rXs8uF41_2),.clk(gclk));
	jdff dff_B_QItZIc6D2_2(.din(w_dff_B_1rXs8uF41_2),.dout(w_dff_B_QItZIc6D2_2),.clk(gclk));
	jdff dff_B_DrbFUlg39_2(.din(w_dff_B_QItZIc6D2_2),.dout(w_dff_B_DrbFUlg39_2),.clk(gclk));
	jdff dff_B_ScDjIgIN3_2(.din(w_dff_B_DrbFUlg39_2),.dout(w_dff_B_ScDjIgIN3_2),.clk(gclk));
	jdff dff_B_SDXyv6ay4_2(.din(w_dff_B_ScDjIgIN3_2),.dout(w_dff_B_SDXyv6ay4_2),.clk(gclk));
	jdff dff_B_BEQgbryD0_2(.din(w_dff_B_SDXyv6ay4_2),.dout(w_dff_B_BEQgbryD0_2),.clk(gclk));
	jdff dff_B_UImHBzLF6_2(.din(w_dff_B_BEQgbryD0_2),.dout(w_dff_B_UImHBzLF6_2),.clk(gclk));
	jdff dff_B_KwO1WfyY5_2(.din(w_dff_B_UImHBzLF6_2),.dout(w_dff_B_KwO1WfyY5_2),.clk(gclk));
	jdff dff_B_2FHoCyLs4_2(.din(w_dff_B_KwO1WfyY5_2),.dout(w_dff_B_2FHoCyLs4_2),.clk(gclk));
	jdff dff_B_9RmJStxt8_2(.din(n795),.dout(w_dff_B_9RmJStxt8_2),.clk(gclk));
	jdff dff_B_bl7gv11g3_1(.din(n725),.dout(w_dff_B_bl7gv11g3_1),.clk(gclk));
	jdff dff_B_sgctC2ms6_2(.din(n632),.dout(w_dff_B_sgctC2ms6_2),.clk(gclk));
	jdff dff_B_QDlLT5Dg2_2(.din(w_dff_B_sgctC2ms6_2),.dout(w_dff_B_QDlLT5Dg2_2),.clk(gclk));
	jdff dff_B_5PJko8JB2_2(.din(w_dff_B_QDlLT5Dg2_2),.dout(w_dff_B_5PJko8JB2_2),.clk(gclk));
	jdff dff_B_xg0tMxRL1_2(.din(w_dff_B_5PJko8JB2_2),.dout(w_dff_B_xg0tMxRL1_2),.clk(gclk));
	jdff dff_B_I9VxXEZz3_2(.din(w_dff_B_xg0tMxRL1_2),.dout(w_dff_B_I9VxXEZz3_2),.clk(gclk));
	jdff dff_B_tL0DKbUx6_2(.din(w_dff_B_I9VxXEZz3_2),.dout(w_dff_B_tL0DKbUx6_2),.clk(gclk));
	jdff dff_B_QuV1SDT26_2(.din(w_dff_B_tL0DKbUx6_2),.dout(w_dff_B_QuV1SDT26_2),.clk(gclk));
	jdff dff_B_BV28o4XO2_2(.din(w_dff_B_QuV1SDT26_2),.dout(w_dff_B_BV28o4XO2_2),.clk(gclk));
	jdff dff_B_70khY1v44_2(.din(w_dff_B_BV28o4XO2_2),.dout(w_dff_B_70khY1v44_2),.clk(gclk));
	jdff dff_B_6F2iZ29O1_2(.din(w_dff_B_70khY1v44_2),.dout(w_dff_B_6F2iZ29O1_2),.clk(gclk));
	jdff dff_B_jgAw1G9q7_2(.din(w_dff_B_6F2iZ29O1_2),.dout(w_dff_B_jgAw1G9q7_2),.clk(gclk));
	jdff dff_B_sOofq8fZ9_2(.din(w_dff_B_jgAw1G9q7_2),.dout(w_dff_B_sOofq8fZ9_2),.clk(gclk));
	jdff dff_B_mDwnVTuZ6_2(.din(w_dff_B_sOofq8fZ9_2),.dout(w_dff_B_mDwnVTuZ6_2),.clk(gclk));
	jdff dff_B_h4Szrg7x8_2(.din(w_dff_B_mDwnVTuZ6_2),.dout(w_dff_B_h4Szrg7x8_2),.clk(gclk));
	jdff dff_B_gEc78X3u3_2(.din(w_dff_B_h4Szrg7x8_2),.dout(w_dff_B_gEc78X3u3_2),.clk(gclk));
	jdff dff_B_FOoxqQW81_2(.din(w_dff_B_gEc78X3u3_2),.dout(w_dff_B_FOoxqQW81_2),.clk(gclk));
	jdff dff_B_zFZf0V4C5_2(.din(w_dff_B_FOoxqQW81_2),.dout(w_dff_B_zFZf0V4C5_2),.clk(gclk));
	jdff dff_B_ccihcXOc7_2(.din(w_dff_B_zFZf0V4C5_2),.dout(w_dff_B_ccihcXOc7_2),.clk(gclk));
	jdff dff_B_BYTy5ETk6_2(.din(w_dff_B_ccihcXOc7_2),.dout(w_dff_B_BYTy5ETk6_2),.clk(gclk));
	jdff dff_B_dgjtkW2T1_2(.din(w_dff_B_BYTy5ETk6_2),.dout(w_dff_B_dgjtkW2T1_2),.clk(gclk));
	jdff dff_B_h6GEwEum3_2(.din(w_dff_B_dgjtkW2T1_2),.dout(w_dff_B_h6GEwEum3_2),.clk(gclk));
	jdff dff_B_x0NX5xOp9_2(.din(w_dff_B_h6GEwEum3_2),.dout(w_dff_B_x0NX5xOp9_2),.clk(gclk));
	jdff dff_B_KKb1EUnh2_2(.din(w_dff_B_x0NX5xOp9_2),.dout(w_dff_B_KKb1EUnh2_2),.clk(gclk));
	jdff dff_B_lAiRSUL17_2(.din(w_dff_B_KKb1EUnh2_2),.dout(w_dff_B_lAiRSUL17_2),.clk(gclk));
	jdff dff_B_ZtL614pE9_2(.din(w_dff_B_lAiRSUL17_2),.dout(w_dff_B_ZtL614pE9_2),.clk(gclk));
	jdff dff_B_nJVDWohz7_2(.din(w_dff_B_ZtL614pE9_2),.dout(w_dff_B_nJVDWohz7_2),.clk(gclk));
	jdff dff_B_VjjXjdD76_2(.din(w_dff_B_nJVDWohz7_2),.dout(w_dff_B_VjjXjdD76_2),.clk(gclk));
	jdff dff_B_aBR7h1Hy2_2(.din(n696),.dout(w_dff_B_aBR7h1Hy2_2),.clk(gclk));
	jdff dff_B_aD7x3mA87_1(.din(n633),.dout(w_dff_B_aD7x3mA87_1),.clk(gclk));
	jdff dff_B_THAfjzzN6_2(.din(n547),.dout(w_dff_B_THAfjzzN6_2),.clk(gclk));
	jdff dff_B_fpMykrte6_2(.din(w_dff_B_THAfjzzN6_2),.dout(w_dff_B_fpMykrte6_2),.clk(gclk));
	jdff dff_B_i5MGwZqR6_2(.din(w_dff_B_fpMykrte6_2),.dout(w_dff_B_i5MGwZqR6_2),.clk(gclk));
	jdff dff_B_wrL4KYTs4_2(.din(w_dff_B_i5MGwZqR6_2),.dout(w_dff_B_wrL4KYTs4_2),.clk(gclk));
	jdff dff_B_up88BSOY2_2(.din(w_dff_B_wrL4KYTs4_2),.dout(w_dff_B_up88BSOY2_2),.clk(gclk));
	jdff dff_B_JXgeXzgy7_2(.din(w_dff_B_up88BSOY2_2),.dout(w_dff_B_JXgeXzgy7_2),.clk(gclk));
	jdff dff_B_S2FjTR3z9_2(.din(w_dff_B_JXgeXzgy7_2),.dout(w_dff_B_S2FjTR3z9_2),.clk(gclk));
	jdff dff_B_NE2Htc2V6_2(.din(w_dff_B_S2FjTR3z9_2),.dout(w_dff_B_NE2Htc2V6_2),.clk(gclk));
	jdff dff_B_ZDuH2iOY1_2(.din(w_dff_B_NE2Htc2V6_2),.dout(w_dff_B_ZDuH2iOY1_2),.clk(gclk));
	jdff dff_B_a2saWzPG6_2(.din(w_dff_B_ZDuH2iOY1_2),.dout(w_dff_B_a2saWzPG6_2),.clk(gclk));
	jdff dff_B_Ru4ExJ7l9_2(.din(w_dff_B_a2saWzPG6_2),.dout(w_dff_B_Ru4ExJ7l9_2),.clk(gclk));
	jdff dff_B_p4PIKxPn9_2(.din(w_dff_B_Ru4ExJ7l9_2),.dout(w_dff_B_p4PIKxPn9_2),.clk(gclk));
	jdff dff_B_IYBh4PKs9_2(.din(w_dff_B_p4PIKxPn9_2),.dout(w_dff_B_IYBh4PKs9_2),.clk(gclk));
	jdff dff_B_gn1RbeKP9_2(.din(w_dff_B_IYBh4PKs9_2),.dout(w_dff_B_gn1RbeKP9_2),.clk(gclk));
	jdff dff_B_JobxkEj82_2(.din(w_dff_B_gn1RbeKP9_2),.dout(w_dff_B_JobxkEj82_2),.clk(gclk));
	jdff dff_B_eyyG0nGG4_2(.din(w_dff_B_JobxkEj82_2),.dout(w_dff_B_eyyG0nGG4_2),.clk(gclk));
	jdff dff_B_SMrOrYep3_2(.din(w_dff_B_eyyG0nGG4_2),.dout(w_dff_B_SMrOrYep3_2),.clk(gclk));
	jdff dff_B_wQB0DR4o7_2(.din(w_dff_B_SMrOrYep3_2),.dout(w_dff_B_wQB0DR4o7_2),.clk(gclk));
	jdff dff_B_SnnuDMwd1_2(.din(w_dff_B_wQB0DR4o7_2),.dout(w_dff_B_SnnuDMwd1_2),.clk(gclk));
	jdff dff_B_yA9eEGGP0_2(.din(w_dff_B_SnnuDMwd1_2),.dout(w_dff_B_yA9eEGGP0_2),.clk(gclk));
	jdff dff_B_2AykSPL21_2(.din(w_dff_B_yA9eEGGP0_2),.dout(w_dff_B_2AykSPL21_2),.clk(gclk));
	jdff dff_B_F7yXKers5_2(.din(w_dff_B_2AykSPL21_2),.dout(w_dff_B_F7yXKers5_2),.clk(gclk));
	jdff dff_B_li0uOzq46_2(.din(w_dff_B_F7yXKers5_2),.dout(w_dff_B_li0uOzq46_2),.clk(gclk));
	jdff dff_B_0cTUdrvL2_2(.din(w_dff_B_li0uOzq46_2),.dout(w_dff_B_0cTUdrvL2_2),.clk(gclk));
	jdff dff_B_zTSUf4yg2_2(.din(n604),.dout(w_dff_B_zTSUf4yg2_2),.clk(gclk));
	jdff dff_B_JMosQLe99_1(.din(n548),.dout(w_dff_B_JMosQLe99_1),.clk(gclk));
	jdff dff_B_evkuoxgF7_2(.din(n469),.dout(w_dff_B_evkuoxgF7_2),.clk(gclk));
	jdff dff_B_vmepfc7l6_2(.din(w_dff_B_evkuoxgF7_2),.dout(w_dff_B_vmepfc7l6_2),.clk(gclk));
	jdff dff_B_Uv072pIe8_2(.din(w_dff_B_vmepfc7l6_2),.dout(w_dff_B_Uv072pIe8_2),.clk(gclk));
	jdff dff_B_WiOPty1Y5_2(.din(w_dff_B_Uv072pIe8_2),.dout(w_dff_B_WiOPty1Y5_2),.clk(gclk));
	jdff dff_B_COZ8HxcW5_2(.din(w_dff_B_WiOPty1Y5_2),.dout(w_dff_B_COZ8HxcW5_2),.clk(gclk));
	jdff dff_B_pkToUIgK6_2(.din(w_dff_B_COZ8HxcW5_2),.dout(w_dff_B_pkToUIgK6_2),.clk(gclk));
	jdff dff_B_SHoS1vMN9_2(.din(w_dff_B_pkToUIgK6_2),.dout(w_dff_B_SHoS1vMN9_2),.clk(gclk));
	jdff dff_B_tuZ4q8mk1_2(.din(w_dff_B_SHoS1vMN9_2),.dout(w_dff_B_tuZ4q8mk1_2),.clk(gclk));
	jdff dff_B_adbh6YNe3_2(.din(w_dff_B_tuZ4q8mk1_2),.dout(w_dff_B_adbh6YNe3_2),.clk(gclk));
	jdff dff_B_PicBMPJH2_2(.din(w_dff_B_adbh6YNe3_2),.dout(w_dff_B_PicBMPJH2_2),.clk(gclk));
	jdff dff_B_5lGIudHz2_2(.din(w_dff_B_PicBMPJH2_2),.dout(w_dff_B_5lGIudHz2_2),.clk(gclk));
	jdff dff_B_kVmSAe5U9_2(.din(w_dff_B_5lGIudHz2_2),.dout(w_dff_B_kVmSAe5U9_2),.clk(gclk));
	jdff dff_B_0EcuB2rK7_2(.din(w_dff_B_kVmSAe5U9_2),.dout(w_dff_B_0EcuB2rK7_2),.clk(gclk));
	jdff dff_B_xUEFUTM94_2(.din(w_dff_B_0EcuB2rK7_2),.dout(w_dff_B_xUEFUTM94_2),.clk(gclk));
	jdff dff_B_Yb3MFoWe3_2(.din(w_dff_B_xUEFUTM94_2),.dout(w_dff_B_Yb3MFoWe3_2),.clk(gclk));
	jdff dff_B_V3ysKATD7_2(.din(w_dff_B_Yb3MFoWe3_2),.dout(w_dff_B_V3ysKATD7_2),.clk(gclk));
	jdff dff_B_lki6xDrr8_2(.din(w_dff_B_V3ysKATD7_2),.dout(w_dff_B_lki6xDrr8_2),.clk(gclk));
	jdff dff_B_DgVIYWTG7_2(.din(w_dff_B_lki6xDrr8_2),.dout(w_dff_B_DgVIYWTG7_2),.clk(gclk));
	jdff dff_B_zB03IuIx7_2(.din(w_dff_B_DgVIYWTG7_2),.dout(w_dff_B_zB03IuIx7_2),.clk(gclk));
	jdff dff_B_xAiTgPQE0_2(.din(w_dff_B_zB03IuIx7_2),.dout(w_dff_B_xAiTgPQE0_2),.clk(gclk));
	jdff dff_B_VqpNoIgB5_2(.din(w_dff_B_xAiTgPQE0_2),.dout(w_dff_B_VqpNoIgB5_2),.clk(gclk));
	jdff dff_B_zFtsBFuG7_2(.din(n519),.dout(w_dff_B_zFtsBFuG7_2),.clk(gclk));
	jdff dff_B_U0htOr0J6_1(.din(n470),.dout(w_dff_B_U0htOr0J6_1),.clk(gclk));
	jdff dff_B_KUgqZjEE7_2(.din(n398),.dout(w_dff_B_KUgqZjEE7_2),.clk(gclk));
	jdff dff_B_wxUNL26q6_2(.din(w_dff_B_KUgqZjEE7_2),.dout(w_dff_B_wxUNL26q6_2),.clk(gclk));
	jdff dff_B_xiJ0v6c28_2(.din(w_dff_B_wxUNL26q6_2),.dout(w_dff_B_xiJ0v6c28_2),.clk(gclk));
	jdff dff_B_vQplVdSV2_2(.din(w_dff_B_xiJ0v6c28_2),.dout(w_dff_B_vQplVdSV2_2),.clk(gclk));
	jdff dff_B_Cl9pVdzs3_2(.din(w_dff_B_vQplVdSV2_2),.dout(w_dff_B_Cl9pVdzs3_2),.clk(gclk));
	jdff dff_B_KlkEIGIx6_2(.din(w_dff_B_Cl9pVdzs3_2),.dout(w_dff_B_KlkEIGIx6_2),.clk(gclk));
	jdff dff_B_FBu0J2Su7_2(.din(w_dff_B_KlkEIGIx6_2),.dout(w_dff_B_FBu0J2Su7_2),.clk(gclk));
	jdff dff_B_w6KgQCQM0_2(.din(w_dff_B_FBu0J2Su7_2),.dout(w_dff_B_w6KgQCQM0_2),.clk(gclk));
	jdff dff_B_i4Dilrae4_2(.din(w_dff_B_w6KgQCQM0_2),.dout(w_dff_B_i4Dilrae4_2),.clk(gclk));
	jdff dff_B_3KyqIZti9_2(.din(w_dff_B_i4Dilrae4_2),.dout(w_dff_B_3KyqIZti9_2),.clk(gclk));
	jdff dff_B_LwtuXjcv0_2(.din(w_dff_B_3KyqIZti9_2),.dout(w_dff_B_LwtuXjcv0_2),.clk(gclk));
	jdff dff_B_8fQ49QiS7_2(.din(w_dff_B_LwtuXjcv0_2),.dout(w_dff_B_8fQ49QiS7_2),.clk(gclk));
	jdff dff_B_fEVbJMi30_2(.din(w_dff_B_8fQ49QiS7_2),.dout(w_dff_B_fEVbJMi30_2),.clk(gclk));
	jdff dff_B_juLqisgc0_2(.din(w_dff_B_fEVbJMi30_2),.dout(w_dff_B_juLqisgc0_2),.clk(gclk));
	jdff dff_B_wfezRKVB2_2(.din(w_dff_B_juLqisgc0_2),.dout(w_dff_B_wfezRKVB2_2),.clk(gclk));
	jdff dff_B_GbsgmZ433_2(.din(w_dff_B_wfezRKVB2_2),.dout(w_dff_B_GbsgmZ433_2),.clk(gclk));
	jdff dff_B_iPrzVBwB6_2(.din(w_dff_B_GbsgmZ433_2),.dout(w_dff_B_iPrzVBwB6_2),.clk(gclk));
	jdff dff_B_mLPwvyRw6_2(.din(w_dff_B_iPrzVBwB6_2),.dout(w_dff_B_mLPwvyRw6_2),.clk(gclk));
	jdff dff_B_XQlWpnvd2_2(.din(n441),.dout(w_dff_B_XQlWpnvd2_2),.clk(gclk));
	jdff dff_B_Iyryb7Ag3_1(.din(n399),.dout(w_dff_B_Iyryb7Ag3_1),.clk(gclk));
	jdff dff_B_L0df6ITD8_2(.din(n335),.dout(w_dff_B_L0df6ITD8_2),.clk(gclk));
	jdff dff_B_aOQyFdbY0_2(.din(w_dff_B_L0df6ITD8_2),.dout(w_dff_B_aOQyFdbY0_2),.clk(gclk));
	jdff dff_B_znBRIrXq5_2(.din(w_dff_B_aOQyFdbY0_2),.dout(w_dff_B_znBRIrXq5_2),.clk(gclk));
	jdff dff_B_gN9lqP0x1_2(.din(w_dff_B_znBRIrXq5_2),.dout(w_dff_B_gN9lqP0x1_2),.clk(gclk));
	jdff dff_B_ktn6rVR98_2(.din(w_dff_B_gN9lqP0x1_2),.dout(w_dff_B_ktn6rVR98_2),.clk(gclk));
	jdff dff_B_a7BAjz0B0_2(.din(w_dff_B_ktn6rVR98_2),.dout(w_dff_B_a7BAjz0B0_2),.clk(gclk));
	jdff dff_B_WXQdLsEp9_2(.din(w_dff_B_a7BAjz0B0_2),.dout(w_dff_B_WXQdLsEp9_2),.clk(gclk));
	jdff dff_B_IZ0zSYvF3_2(.din(w_dff_B_WXQdLsEp9_2),.dout(w_dff_B_IZ0zSYvF3_2),.clk(gclk));
	jdff dff_B_ttIhVM3d9_2(.din(w_dff_B_IZ0zSYvF3_2),.dout(w_dff_B_ttIhVM3d9_2),.clk(gclk));
	jdff dff_B_ye0jgQYT3_2(.din(w_dff_B_ttIhVM3d9_2),.dout(w_dff_B_ye0jgQYT3_2),.clk(gclk));
	jdff dff_B_BW6TAmCM6_2(.din(w_dff_B_ye0jgQYT3_2),.dout(w_dff_B_BW6TAmCM6_2),.clk(gclk));
	jdff dff_B_0g5TJARm0_2(.din(w_dff_B_BW6TAmCM6_2),.dout(w_dff_B_0g5TJARm0_2),.clk(gclk));
	jdff dff_B_y88AwWPC6_2(.din(w_dff_B_0g5TJARm0_2),.dout(w_dff_B_y88AwWPC6_2),.clk(gclk));
	jdff dff_B_NSpNPeqM5_2(.din(w_dff_B_y88AwWPC6_2),.dout(w_dff_B_NSpNPeqM5_2),.clk(gclk));
	jdff dff_B_ZMuS2v2G9_2(.din(w_dff_B_NSpNPeqM5_2),.dout(w_dff_B_ZMuS2v2G9_2),.clk(gclk));
	jdff dff_B_6WoNTM9e2_2(.din(n370),.dout(w_dff_B_6WoNTM9e2_2),.clk(gclk));
	jdff dff_B_3fp6Nyge0_1(.din(n336),.dout(w_dff_B_3fp6Nyge0_1),.clk(gclk));
	jdff dff_B_HOEKbKf41_2(.din(n279),.dout(w_dff_B_HOEKbKf41_2),.clk(gclk));
	jdff dff_B_vuuZnh450_2(.din(w_dff_B_HOEKbKf41_2),.dout(w_dff_B_vuuZnh450_2),.clk(gclk));
	jdff dff_B_Zjcsl5wP6_2(.din(w_dff_B_vuuZnh450_2),.dout(w_dff_B_Zjcsl5wP6_2),.clk(gclk));
	jdff dff_B_nUi9cYoc0_2(.din(w_dff_B_Zjcsl5wP6_2),.dout(w_dff_B_nUi9cYoc0_2),.clk(gclk));
	jdff dff_B_NYBsgyeo4_2(.din(w_dff_B_nUi9cYoc0_2),.dout(w_dff_B_NYBsgyeo4_2),.clk(gclk));
	jdff dff_B_ZaJKuGs42_2(.din(w_dff_B_NYBsgyeo4_2),.dout(w_dff_B_ZaJKuGs42_2),.clk(gclk));
	jdff dff_B_5cZYg6TB4_2(.din(w_dff_B_ZaJKuGs42_2),.dout(w_dff_B_5cZYg6TB4_2),.clk(gclk));
	jdff dff_B_r93McewT1_2(.din(w_dff_B_5cZYg6TB4_2),.dout(w_dff_B_r93McewT1_2),.clk(gclk));
	jdff dff_B_P3Fm3UB04_2(.din(w_dff_B_r93McewT1_2),.dout(w_dff_B_P3Fm3UB04_2),.clk(gclk));
	jdff dff_B_2p6Rr5Ra2_2(.din(w_dff_B_P3Fm3UB04_2),.dout(w_dff_B_2p6Rr5Ra2_2),.clk(gclk));
	jdff dff_B_X7aUmSwt2_2(.din(w_dff_B_2p6Rr5Ra2_2),.dout(w_dff_B_X7aUmSwt2_2),.clk(gclk));
	jdff dff_B_lBNBFkrK6_2(.din(w_dff_B_X7aUmSwt2_2),.dout(w_dff_B_lBNBFkrK6_2),.clk(gclk));
	jdff dff_B_LAmdmyhz3_2(.din(n307),.dout(w_dff_B_LAmdmyhz3_2),.clk(gclk));
	jdff dff_B_yNEAHrJk0_1(.din(n280),.dout(w_dff_B_yNEAHrJk0_1),.clk(gclk));
	jdff dff_B_n9ZaYF507_2(.din(n230),.dout(w_dff_B_n9ZaYF507_2),.clk(gclk));
	jdff dff_B_02VdiIyv7_2(.din(w_dff_B_n9ZaYF507_2),.dout(w_dff_B_02VdiIyv7_2),.clk(gclk));
	jdff dff_B_gcgRUa4g5_2(.din(w_dff_B_02VdiIyv7_2),.dout(w_dff_B_gcgRUa4g5_2),.clk(gclk));
	jdff dff_B_pUFMYXEQ9_2(.din(w_dff_B_gcgRUa4g5_2),.dout(w_dff_B_pUFMYXEQ9_2),.clk(gclk));
	jdff dff_B_7KSL262Q3_2(.din(w_dff_B_pUFMYXEQ9_2),.dout(w_dff_B_7KSL262Q3_2),.clk(gclk));
	jdff dff_B_XhUVsXSg9_2(.din(w_dff_B_7KSL262Q3_2),.dout(w_dff_B_XhUVsXSg9_2),.clk(gclk));
	jdff dff_B_XXTPQTv89_2(.din(w_dff_B_XhUVsXSg9_2),.dout(w_dff_B_XXTPQTv89_2),.clk(gclk));
	jdff dff_B_5DEFtKar6_2(.din(w_dff_B_XXTPQTv89_2),.dout(w_dff_B_5DEFtKar6_2),.clk(gclk));
	jdff dff_B_B1atzNu17_2(.din(w_dff_B_5DEFtKar6_2),.dout(w_dff_B_B1atzNu17_2),.clk(gclk));
	jdff dff_B_nxiq51Ud2_2(.din(n251),.dout(w_dff_B_nxiq51Ud2_2),.clk(gclk));
	jdff dff_B_bmAOyLyk1_1(.din(n231),.dout(w_dff_B_bmAOyLyk1_1),.clk(gclk));
	jdff dff_B_0iZdEHEx9_2(.din(n188),.dout(w_dff_B_0iZdEHEx9_2),.clk(gclk));
	jdff dff_B_o53S9IqX2_2(.din(w_dff_B_0iZdEHEx9_2),.dout(w_dff_B_o53S9IqX2_2),.clk(gclk));
	jdff dff_B_lcyoUKLj0_2(.din(w_dff_B_o53S9IqX2_2),.dout(w_dff_B_lcyoUKLj0_2),.clk(gclk));
	jdff dff_B_SOX6ZN0Z6_2(.din(w_dff_B_lcyoUKLj0_2),.dout(w_dff_B_SOX6ZN0Z6_2),.clk(gclk));
	jdff dff_B_cxulTZoH0_2(.din(w_dff_B_SOX6ZN0Z6_2),.dout(w_dff_B_cxulTZoH0_2),.clk(gclk));
	jdff dff_B_8W3jZQuq6_2(.din(w_dff_B_cxulTZoH0_2),.dout(w_dff_B_8W3jZQuq6_2),.clk(gclk));
	jdff dff_B_iUG0sUcw6_2(.din(n202),.dout(w_dff_B_iUG0sUcw6_2),.clk(gclk));
	jdff dff_B_JuzekZtg4_2(.din(n154),.dout(w_dff_B_JuzekZtg4_2),.clk(gclk));
	jdff dff_B_xb9va1oA8_2(.din(w_dff_B_JuzekZtg4_2),.dout(w_dff_B_xb9va1oA8_2),.clk(gclk));
	jdff dff_B_xEacR6If5_2(.din(w_dff_B_xb9va1oA8_2),.dout(w_dff_B_xEacR6If5_2),.clk(gclk));
	jdff dff_B_r3s5Qos04_0(.din(n159),.dout(w_dff_B_r3s5Qos04_0),.clk(gclk));
	jdff dff_A_3QQsrz8h0_0(.dout(w_n123_0[0]),.din(w_dff_A_3QQsrz8h0_0),.clk(gclk));
	jdff dff_A_tqDlP7NW9_0(.dout(w_dff_A_3QQsrz8h0_0),.din(w_dff_A_tqDlP7NW9_0),.clk(gclk));
	jdff dff_A_qChiSjTT1_0(.dout(w_n122_0[0]),.din(w_dff_A_qChiSjTT1_0),.clk(gclk));
	jdff dff_A_9ki8toQ61_0(.dout(w_dff_A_qChiSjTT1_0),.din(w_dff_A_9ki8toQ61_0),.clk(gclk));
	jdff dff_B_0Tq9flrP8_1(.din(n1304),.dout(w_dff_B_0Tq9flrP8_1),.clk(gclk));
	jdff dff_B_RC3DzLJi9_2(.din(n1217),.dout(w_dff_B_RC3DzLJi9_2),.clk(gclk));
	jdff dff_B_41vVKmW97_2(.din(w_dff_B_RC3DzLJi9_2),.dout(w_dff_B_41vVKmW97_2),.clk(gclk));
	jdff dff_B_Vy2zL9cD0_2(.din(w_dff_B_41vVKmW97_2),.dout(w_dff_B_Vy2zL9cD0_2),.clk(gclk));
	jdff dff_B_xvNydhBx9_2(.din(w_dff_B_Vy2zL9cD0_2),.dout(w_dff_B_xvNydhBx9_2),.clk(gclk));
	jdff dff_B_yYeXScd81_2(.din(w_dff_B_xvNydhBx9_2),.dout(w_dff_B_yYeXScd81_2),.clk(gclk));
	jdff dff_B_xe1jJSAf0_2(.din(w_dff_B_yYeXScd81_2),.dout(w_dff_B_xe1jJSAf0_2),.clk(gclk));
	jdff dff_B_FMKqSaua2_2(.din(w_dff_B_xe1jJSAf0_2),.dout(w_dff_B_FMKqSaua2_2),.clk(gclk));
	jdff dff_B_H9R5l9Ci5_2(.din(w_dff_B_FMKqSaua2_2),.dout(w_dff_B_H9R5l9Ci5_2),.clk(gclk));
	jdff dff_B_RJ6utOV02_2(.din(w_dff_B_H9R5l9Ci5_2),.dout(w_dff_B_RJ6utOV02_2),.clk(gclk));
	jdff dff_B_CqkL9ZQR2_2(.din(w_dff_B_RJ6utOV02_2),.dout(w_dff_B_CqkL9ZQR2_2),.clk(gclk));
	jdff dff_B_8xhQzuQ41_2(.din(w_dff_B_CqkL9ZQR2_2),.dout(w_dff_B_8xhQzuQ41_2),.clk(gclk));
	jdff dff_B_qXaQoU6P6_2(.din(w_dff_B_8xhQzuQ41_2),.dout(w_dff_B_qXaQoU6P6_2),.clk(gclk));
	jdff dff_B_vOouALVs6_2(.din(w_dff_B_qXaQoU6P6_2),.dout(w_dff_B_vOouALVs6_2),.clk(gclk));
	jdff dff_B_4TpawNZv0_2(.din(w_dff_B_vOouALVs6_2),.dout(w_dff_B_4TpawNZv0_2),.clk(gclk));
	jdff dff_B_HkU3zgBf5_2(.din(w_dff_B_4TpawNZv0_2),.dout(w_dff_B_HkU3zgBf5_2),.clk(gclk));
	jdff dff_B_506aG5TU7_2(.din(w_dff_B_HkU3zgBf5_2),.dout(w_dff_B_506aG5TU7_2),.clk(gclk));
	jdff dff_B_iMfTyXVX4_2(.din(w_dff_B_506aG5TU7_2),.dout(w_dff_B_iMfTyXVX4_2),.clk(gclk));
	jdff dff_B_Psn9Xlde3_2(.din(w_dff_B_iMfTyXVX4_2),.dout(w_dff_B_Psn9Xlde3_2),.clk(gclk));
	jdff dff_B_MdIewARP2_2(.din(w_dff_B_Psn9Xlde3_2),.dout(w_dff_B_MdIewARP2_2),.clk(gclk));
	jdff dff_B_PyGevuDR5_2(.din(w_dff_B_MdIewARP2_2),.dout(w_dff_B_PyGevuDR5_2),.clk(gclk));
	jdff dff_B_vjyZ07B55_2(.din(w_dff_B_PyGevuDR5_2),.dout(w_dff_B_vjyZ07B55_2),.clk(gclk));
	jdff dff_B_yMMg5mFA0_2(.din(w_dff_B_vjyZ07B55_2),.dout(w_dff_B_yMMg5mFA0_2),.clk(gclk));
	jdff dff_B_p3mljQqH1_2(.din(w_dff_B_yMMg5mFA0_2),.dout(w_dff_B_p3mljQqH1_2),.clk(gclk));
	jdff dff_B_ga7XhXMp3_2(.din(w_dff_B_p3mljQqH1_2),.dout(w_dff_B_ga7XhXMp3_2),.clk(gclk));
	jdff dff_B_50FIKzDS2_2(.din(w_dff_B_ga7XhXMp3_2),.dout(w_dff_B_50FIKzDS2_2),.clk(gclk));
	jdff dff_B_gp9e7UAL7_2(.din(w_dff_B_50FIKzDS2_2),.dout(w_dff_B_gp9e7UAL7_2),.clk(gclk));
	jdff dff_B_8ZNOG0zT5_2(.din(w_dff_B_gp9e7UAL7_2),.dout(w_dff_B_8ZNOG0zT5_2),.clk(gclk));
	jdff dff_B_bTM5Vijz5_2(.din(w_dff_B_8ZNOG0zT5_2),.dout(w_dff_B_bTM5Vijz5_2),.clk(gclk));
	jdff dff_B_ghHWn50z7_2(.din(w_dff_B_bTM5Vijz5_2),.dout(w_dff_B_ghHWn50z7_2),.clk(gclk));
	jdff dff_B_MKu59GoH2_2(.din(w_dff_B_ghHWn50z7_2),.dout(w_dff_B_MKu59GoH2_2),.clk(gclk));
	jdff dff_B_UP3upJe72_2(.din(w_dff_B_MKu59GoH2_2),.dout(w_dff_B_UP3upJe72_2),.clk(gclk));
	jdff dff_B_Gt73K3dY1_2(.din(w_dff_B_UP3upJe72_2),.dout(w_dff_B_Gt73K3dY1_2),.clk(gclk));
	jdff dff_B_nmZshGw77_2(.din(w_dff_B_Gt73K3dY1_2),.dout(w_dff_B_nmZshGw77_2),.clk(gclk));
	jdff dff_B_TdlP5mEs6_2(.din(w_dff_B_nmZshGw77_2),.dout(w_dff_B_TdlP5mEs6_2),.clk(gclk));
	jdff dff_B_RCtarpdH5_2(.din(w_dff_B_TdlP5mEs6_2),.dout(w_dff_B_RCtarpdH5_2),.clk(gclk));
	jdff dff_B_TBChotMj6_2(.din(w_dff_B_RCtarpdH5_2),.dout(w_dff_B_TBChotMj6_2),.clk(gclk));
	jdff dff_B_admalDvB7_2(.din(w_dff_B_TBChotMj6_2),.dout(w_dff_B_admalDvB7_2),.clk(gclk));
	jdff dff_B_dVmmNH8Q3_2(.din(w_dff_B_admalDvB7_2),.dout(w_dff_B_dVmmNH8Q3_2),.clk(gclk));
	jdff dff_B_LgFQUSNZ4_2(.din(w_dff_B_dVmmNH8Q3_2),.dout(w_dff_B_LgFQUSNZ4_2),.clk(gclk));
	jdff dff_B_yPxKtyo95_2(.din(w_dff_B_LgFQUSNZ4_2),.dout(w_dff_B_yPxKtyo95_2),.clk(gclk));
	jdff dff_B_1UWqrAzI4_2(.din(w_dff_B_yPxKtyo95_2),.dout(w_dff_B_1UWqrAzI4_2),.clk(gclk));
	jdff dff_B_ViywdTj95_2(.din(w_dff_B_1UWqrAzI4_2),.dout(w_dff_B_ViywdTj95_2),.clk(gclk));
	jdff dff_B_RnfD60v84_2(.din(w_dff_B_ViywdTj95_2),.dout(w_dff_B_RnfD60v84_2),.clk(gclk));
	jdff dff_B_8NRw3rHp5_2(.din(w_dff_B_RnfD60v84_2),.dout(w_dff_B_8NRw3rHp5_2),.clk(gclk));
	jdff dff_B_DIbn7qAF3_0(.din(n1303),.dout(w_dff_B_DIbn7qAF3_0),.clk(gclk));
	jdff dff_A_lYf27aFO6_1(.dout(w_n1291_0[1]),.din(w_dff_A_lYf27aFO6_1),.clk(gclk));
	jdff dff_B_5b7MHFLe9_1(.din(n1218),.dout(w_dff_B_5b7MHFLe9_1),.clk(gclk));
	jdff dff_B_vbDbSqNB6_2(.din(n1126),.dout(w_dff_B_vbDbSqNB6_2),.clk(gclk));
	jdff dff_B_OSMIUIRZ4_2(.din(w_dff_B_vbDbSqNB6_2),.dout(w_dff_B_OSMIUIRZ4_2),.clk(gclk));
	jdff dff_B_LwqzFRSM7_2(.din(w_dff_B_OSMIUIRZ4_2),.dout(w_dff_B_LwqzFRSM7_2),.clk(gclk));
	jdff dff_B_UWrPxdzc7_2(.din(w_dff_B_LwqzFRSM7_2),.dout(w_dff_B_UWrPxdzc7_2),.clk(gclk));
	jdff dff_B_KnFwu6QV4_2(.din(w_dff_B_UWrPxdzc7_2),.dout(w_dff_B_KnFwu6QV4_2),.clk(gclk));
	jdff dff_B_qRFYBKY82_2(.din(w_dff_B_KnFwu6QV4_2),.dout(w_dff_B_qRFYBKY82_2),.clk(gclk));
	jdff dff_B_cZtzH5tg7_2(.din(w_dff_B_qRFYBKY82_2),.dout(w_dff_B_cZtzH5tg7_2),.clk(gclk));
	jdff dff_B_KRrw8Jvd2_2(.din(w_dff_B_cZtzH5tg7_2),.dout(w_dff_B_KRrw8Jvd2_2),.clk(gclk));
	jdff dff_B_ex9EOPU21_2(.din(w_dff_B_KRrw8Jvd2_2),.dout(w_dff_B_ex9EOPU21_2),.clk(gclk));
	jdff dff_B_O0tfZ5s76_2(.din(w_dff_B_ex9EOPU21_2),.dout(w_dff_B_O0tfZ5s76_2),.clk(gclk));
	jdff dff_B_4ilJbEqV7_2(.din(w_dff_B_O0tfZ5s76_2),.dout(w_dff_B_4ilJbEqV7_2),.clk(gclk));
	jdff dff_B_Z7PfLtWP3_2(.din(w_dff_B_4ilJbEqV7_2),.dout(w_dff_B_Z7PfLtWP3_2),.clk(gclk));
	jdff dff_B_ejOFnKkv3_2(.din(w_dff_B_Z7PfLtWP3_2),.dout(w_dff_B_ejOFnKkv3_2),.clk(gclk));
	jdff dff_B_CDZaLuLw8_2(.din(w_dff_B_ejOFnKkv3_2),.dout(w_dff_B_CDZaLuLw8_2),.clk(gclk));
	jdff dff_B_YKGkE7RC2_2(.din(w_dff_B_CDZaLuLw8_2),.dout(w_dff_B_YKGkE7RC2_2),.clk(gclk));
	jdff dff_B_VdZKIYkh7_2(.din(w_dff_B_YKGkE7RC2_2),.dout(w_dff_B_VdZKIYkh7_2),.clk(gclk));
	jdff dff_B_roL2bsNd8_2(.din(w_dff_B_VdZKIYkh7_2),.dout(w_dff_B_roL2bsNd8_2),.clk(gclk));
	jdff dff_B_B5cJly2x4_2(.din(w_dff_B_roL2bsNd8_2),.dout(w_dff_B_B5cJly2x4_2),.clk(gclk));
	jdff dff_B_WJc95NuN1_2(.din(w_dff_B_B5cJly2x4_2),.dout(w_dff_B_WJc95NuN1_2),.clk(gclk));
	jdff dff_B_9WeYMuTj5_2(.din(w_dff_B_WJc95NuN1_2),.dout(w_dff_B_9WeYMuTj5_2),.clk(gclk));
	jdff dff_B_lyxoAaqq6_2(.din(w_dff_B_9WeYMuTj5_2),.dout(w_dff_B_lyxoAaqq6_2),.clk(gclk));
	jdff dff_B_xaBHL6Jf8_2(.din(w_dff_B_lyxoAaqq6_2),.dout(w_dff_B_xaBHL6Jf8_2),.clk(gclk));
	jdff dff_B_237AxNRa0_2(.din(w_dff_B_xaBHL6Jf8_2),.dout(w_dff_B_237AxNRa0_2),.clk(gclk));
	jdff dff_B_zjWZUXKu3_2(.din(w_dff_B_237AxNRa0_2),.dout(w_dff_B_zjWZUXKu3_2),.clk(gclk));
	jdff dff_B_Totrr1c28_2(.din(w_dff_B_zjWZUXKu3_2),.dout(w_dff_B_Totrr1c28_2),.clk(gclk));
	jdff dff_B_yHnZ6pZd3_2(.din(w_dff_B_Totrr1c28_2),.dout(w_dff_B_yHnZ6pZd3_2),.clk(gclk));
	jdff dff_B_CaqJxvK11_2(.din(w_dff_B_yHnZ6pZd3_2),.dout(w_dff_B_CaqJxvK11_2),.clk(gclk));
	jdff dff_B_buvGEhHE4_2(.din(w_dff_B_CaqJxvK11_2),.dout(w_dff_B_buvGEhHE4_2),.clk(gclk));
	jdff dff_B_21VvH6B65_2(.din(w_dff_B_buvGEhHE4_2),.dout(w_dff_B_21VvH6B65_2),.clk(gclk));
	jdff dff_B_C1ONkMfs3_2(.din(w_dff_B_21VvH6B65_2),.dout(w_dff_B_C1ONkMfs3_2),.clk(gclk));
	jdff dff_B_MMXkNZlI3_2(.din(w_dff_B_C1ONkMfs3_2),.dout(w_dff_B_MMXkNZlI3_2),.clk(gclk));
	jdff dff_B_g2Wjjm5N4_2(.din(w_dff_B_MMXkNZlI3_2),.dout(w_dff_B_g2Wjjm5N4_2),.clk(gclk));
	jdff dff_B_v3Ri2d5g7_2(.din(w_dff_B_g2Wjjm5N4_2),.dout(w_dff_B_v3Ri2d5g7_2),.clk(gclk));
	jdff dff_B_mTtG2pcZ8_2(.din(w_dff_B_v3Ri2d5g7_2),.dout(w_dff_B_mTtG2pcZ8_2),.clk(gclk));
	jdff dff_B_sLrCaugh6_2(.din(w_dff_B_mTtG2pcZ8_2),.dout(w_dff_B_sLrCaugh6_2),.clk(gclk));
	jdff dff_B_WTcQIfv96_2(.din(w_dff_B_sLrCaugh6_2),.dout(w_dff_B_WTcQIfv96_2),.clk(gclk));
	jdff dff_B_qjvsO5PI5_2(.din(w_dff_B_WTcQIfv96_2),.dout(w_dff_B_qjvsO5PI5_2),.clk(gclk));
	jdff dff_B_2Z3H3mR92_2(.din(w_dff_B_qjvsO5PI5_2),.dout(w_dff_B_2Z3H3mR92_2),.clk(gclk));
	jdff dff_B_e1hx0Z8G3_2(.din(w_dff_B_2Z3H3mR92_2),.dout(w_dff_B_e1hx0Z8G3_2),.clk(gclk));
	jdff dff_B_xyI3tAO59_2(.din(n1200),.dout(w_dff_B_xyI3tAO59_2),.clk(gclk));
	jdff dff_B_ALbNq03a9_1(.din(n1127),.dout(w_dff_B_ALbNq03a9_1),.clk(gclk));
	jdff dff_B_v2dMiSA64_2(.din(n1028),.dout(w_dff_B_v2dMiSA64_2),.clk(gclk));
	jdff dff_B_bUR6Jbse2_2(.din(w_dff_B_v2dMiSA64_2),.dout(w_dff_B_bUR6Jbse2_2),.clk(gclk));
	jdff dff_B_LQiljXHt6_2(.din(w_dff_B_bUR6Jbse2_2),.dout(w_dff_B_LQiljXHt6_2),.clk(gclk));
	jdff dff_B_G0NB0KcF0_2(.din(w_dff_B_LQiljXHt6_2),.dout(w_dff_B_G0NB0KcF0_2),.clk(gclk));
	jdff dff_B_sXUbyWm39_2(.din(w_dff_B_G0NB0KcF0_2),.dout(w_dff_B_sXUbyWm39_2),.clk(gclk));
	jdff dff_B_PF3v1WVF3_2(.din(w_dff_B_sXUbyWm39_2),.dout(w_dff_B_PF3v1WVF3_2),.clk(gclk));
	jdff dff_B_vEeFK2NN9_2(.din(w_dff_B_PF3v1WVF3_2),.dout(w_dff_B_vEeFK2NN9_2),.clk(gclk));
	jdff dff_B_CTHnz4QK6_2(.din(w_dff_B_vEeFK2NN9_2),.dout(w_dff_B_CTHnz4QK6_2),.clk(gclk));
	jdff dff_B_KzRjYztY3_2(.din(w_dff_B_CTHnz4QK6_2),.dout(w_dff_B_KzRjYztY3_2),.clk(gclk));
	jdff dff_B_6YWGK0mB3_2(.din(w_dff_B_KzRjYztY3_2),.dout(w_dff_B_6YWGK0mB3_2),.clk(gclk));
	jdff dff_B_Ne9oEF0r1_2(.din(w_dff_B_6YWGK0mB3_2),.dout(w_dff_B_Ne9oEF0r1_2),.clk(gclk));
	jdff dff_B_kPvIBqUA6_2(.din(w_dff_B_Ne9oEF0r1_2),.dout(w_dff_B_kPvIBqUA6_2),.clk(gclk));
	jdff dff_B_DNHDwCFR7_2(.din(w_dff_B_kPvIBqUA6_2),.dout(w_dff_B_DNHDwCFR7_2),.clk(gclk));
	jdff dff_B_7h5yKv5G1_2(.din(w_dff_B_DNHDwCFR7_2),.dout(w_dff_B_7h5yKv5G1_2),.clk(gclk));
	jdff dff_B_vGzsnYHc3_2(.din(w_dff_B_7h5yKv5G1_2),.dout(w_dff_B_vGzsnYHc3_2),.clk(gclk));
	jdff dff_B_dSx3LZEv9_2(.din(w_dff_B_vGzsnYHc3_2),.dout(w_dff_B_dSx3LZEv9_2),.clk(gclk));
	jdff dff_B_D0yM60QO6_2(.din(w_dff_B_dSx3LZEv9_2),.dout(w_dff_B_D0yM60QO6_2),.clk(gclk));
	jdff dff_B_LlfVOZ4Y4_2(.din(w_dff_B_D0yM60QO6_2),.dout(w_dff_B_LlfVOZ4Y4_2),.clk(gclk));
	jdff dff_B_1ia5lneo8_2(.din(w_dff_B_LlfVOZ4Y4_2),.dout(w_dff_B_1ia5lneo8_2),.clk(gclk));
	jdff dff_B_fNdXa7x81_2(.din(w_dff_B_1ia5lneo8_2),.dout(w_dff_B_fNdXa7x81_2),.clk(gclk));
	jdff dff_B_mnScxryE3_2(.din(w_dff_B_fNdXa7x81_2),.dout(w_dff_B_mnScxryE3_2),.clk(gclk));
	jdff dff_B_mJ0XS2XH3_2(.din(w_dff_B_mnScxryE3_2),.dout(w_dff_B_mJ0XS2XH3_2),.clk(gclk));
	jdff dff_B_0LJkCJNO9_2(.din(w_dff_B_mJ0XS2XH3_2),.dout(w_dff_B_0LJkCJNO9_2),.clk(gclk));
	jdff dff_B_TYxXuLLp1_2(.din(w_dff_B_0LJkCJNO9_2),.dout(w_dff_B_TYxXuLLp1_2),.clk(gclk));
	jdff dff_B_NzfBssT10_2(.din(w_dff_B_TYxXuLLp1_2),.dout(w_dff_B_NzfBssT10_2),.clk(gclk));
	jdff dff_B_xqc7mgcY6_2(.din(w_dff_B_NzfBssT10_2),.dout(w_dff_B_xqc7mgcY6_2),.clk(gclk));
	jdff dff_B_NkXm7E5v4_2(.din(w_dff_B_xqc7mgcY6_2),.dout(w_dff_B_NkXm7E5v4_2),.clk(gclk));
	jdff dff_B_ki8dsgDd2_2(.din(w_dff_B_NkXm7E5v4_2),.dout(w_dff_B_ki8dsgDd2_2),.clk(gclk));
	jdff dff_B_KXl0rC2Y9_2(.din(w_dff_B_ki8dsgDd2_2),.dout(w_dff_B_KXl0rC2Y9_2),.clk(gclk));
	jdff dff_B_Olt5ViON0_2(.din(w_dff_B_KXl0rC2Y9_2),.dout(w_dff_B_Olt5ViON0_2),.clk(gclk));
	jdff dff_B_YPMijV1J2_2(.din(w_dff_B_Olt5ViON0_2),.dout(w_dff_B_YPMijV1J2_2),.clk(gclk));
	jdff dff_B_FWhOfQcU2_2(.din(w_dff_B_YPMijV1J2_2),.dout(w_dff_B_FWhOfQcU2_2),.clk(gclk));
	jdff dff_B_8DdjDPLX7_2(.din(w_dff_B_FWhOfQcU2_2),.dout(w_dff_B_8DdjDPLX7_2),.clk(gclk));
	jdff dff_B_daAklES03_2(.din(w_dff_B_8DdjDPLX7_2),.dout(w_dff_B_daAklES03_2),.clk(gclk));
	jdff dff_B_dTa0L80u3_2(.din(w_dff_B_daAklES03_2),.dout(w_dff_B_dTa0L80u3_2),.clk(gclk));
	jdff dff_B_DZtWG4YR4_2(.din(w_dff_B_dTa0L80u3_2),.dout(w_dff_B_DZtWG4YR4_2),.clk(gclk));
	jdff dff_B_b33kYsUA6_2(.din(n1101),.dout(w_dff_B_b33kYsUA6_2),.clk(gclk));
	jdff dff_B_tM9aG5Ne4_1(.din(n1029),.dout(w_dff_B_tM9aG5Ne4_1),.clk(gclk));
	jdff dff_B_X33akk7n2_2(.din(n929),.dout(w_dff_B_X33akk7n2_2),.clk(gclk));
	jdff dff_B_DtUVPjlF1_2(.din(w_dff_B_X33akk7n2_2),.dout(w_dff_B_DtUVPjlF1_2),.clk(gclk));
	jdff dff_B_rd3KiYXc9_2(.din(w_dff_B_DtUVPjlF1_2),.dout(w_dff_B_rd3KiYXc9_2),.clk(gclk));
	jdff dff_B_uCXfeUfO7_2(.din(w_dff_B_rd3KiYXc9_2),.dout(w_dff_B_uCXfeUfO7_2),.clk(gclk));
	jdff dff_B_1qA0kXFD1_2(.din(w_dff_B_uCXfeUfO7_2),.dout(w_dff_B_1qA0kXFD1_2),.clk(gclk));
	jdff dff_B_CALulnsx6_2(.din(w_dff_B_1qA0kXFD1_2),.dout(w_dff_B_CALulnsx6_2),.clk(gclk));
	jdff dff_B_KXVeKuOc5_2(.din(w_dff_B_CALulnsx6_2),.dout(w_dff_B_KXVeKuOc5_2),.clk(gclk));
	jdff dff_B_ZDdd0oX22_2(.din(w_dff_B_KXVeKuOc5_2),.dout(w_dff_B_ZDdd0oX22_2),.clk(gclk));
	jdff dff_B_qpVt4v6H0_2(.din(w_dff_B_ZDdd0oX22_2),.dout(w_dff_B_qpVt4v6H0_2),.clk(gclk));
	jdff dff_B_hhudREVW2_2(.din(w_dff_B_qpVt4v6H0_2),.dout(w_dff_B_hhudREVW2_2),.clk(gclk));
	jdff dff_B_cEVre46x1_2(.din(w_dff_B_hhudREVW2_2),.dout(w_dff_B_cEVre46x1_2),.clk(gclk));
	jdff dff_B_lBT0qaRG0_2(.din(w_dff_B_cEVre46x1_2),.dout(w_dff_B_lBT0qaRG0_2),.clk(gclk));
	jdff dff_B_uoSgA8na3_2(.din(w_dff_B_lBT0qaRG0_2),.dout(w_dff_B_uoSgA8na3_2),.clk(gclk));
	jdff dff_B_6ioeJRdx1_2(.din(w_dff_B_uoSgA8na3_2),.dout(w_dff_B_6ioeJRdx1_2),.clk(gclk));
	jdff dff_B_ohYpvn1y2_2(.din(w_dff_B_6ioeJRdx1_2),.dout(w_dff_B_ohYpvn1y2_2),.clk(gclk));
	jdff dff_B_mh1Qfucu0_2(.din(w_dff_B_ohYpvn1y2_2),.dout(w_dff_B_mh1Qfucu0_2),.clk(gclk));
	jdff dff_B_Km0WM7KA6_2(.din(w_dff_B_mh1Qfucu0_2),.dout(w_dff_B_Km0WM7KA6_2),.clk(gclk));
	jdff dff_B_yNq2aYil7_2(.din(w_dff_B_Km0WM7KA6_2),.dout(w_dff_B_yNq2aYil7_2),.clk(gclk));
	jdff dff_B_AsRD1YKj7_2(.din(w_dff_B_yNq2aYil7_2),.dout(w_dff_B_AsRD1YKj7_2),.clk(gclk));
	jdff dff_B_qH8dJJgq0_2(.din(w_dff_B_AsRD1YKj7_2),.dout(w_dff_B_qH8dJJgq0_2),.clk(gclk));
	jdff dff_B_oaSuyjv46_2(.din(w_dff_B_qH8dJJgq0_2),.dout(w_dff_B_oaSuyjv46_2),.clk(gclk));
	jdff dff_B_bl5Iuqq96_2(.din(w_dff_B_oaSuyjv46_2),.dout(w_dff_B_bl5Iuqq96_2),.clk(gclk));
	jdff dff_B_kxAFGSW07_2(.din(w_dff_B_bl5Iuqq96_2),.dout(w_dff_B_kxAFGSW07_2),.clk(gclk));
	jdff dff_B_FYRkc7Ru9_2(.din(w_dff_B_kxAFGSW07_2),.dout(w_dff_B_FYRkc7Ru9_2),.clk(gclk));
	jdff dff_B_yg0LnYqi5_2(.din(w_dff_B_FYRkc7Ru9_2),.dout(w_dff_B_yg0LnYqi5_2),.clk(gclk));
	jdff dff_B_I9GAGc4b3_2(.din(w_dff_B_yg0LnYqi5_2),.dout(w_dff_B_I9GAGc4b3_2),.clk(gclk));
	jdff dff_B_12DvJwqp2_2(.din(w_dff_B_I9GAGc4b3_2),.dout(w_dff_B_12DvJwqp2_2),.clk(gclk));
	jdff dff_B_3eo30jx80_2(.din(w_dff_B_12DvJwqp2_2),.dout(w_dff_B_3eo30jx80_2),.clk(gclk));
	jdff dff_B_uscUeEHA5_2(.din(w_dff_B_3eo30jx80_2),.dout(w_dff_B_uscUeEHA5_2),.clk(gclk));
	jdff dff_B_ULinil997_2(.din(w_dff_B_uscUeEHA5_2),.dout(w_dff_B_ULinil997_2),.clk(gclk));
	jdff dff_B_T2cedTRv7_2(.din(w_dff_B_ULinil997_2),.dout(w_dff_B_T2cedTRv7_2),.clk(gclk));
	jdff dff_B_GomBGRAp5_2(.din(w_dff_B_T2cedTRv7_2),.dout(w_dff_B_GomBGRAp5_2),.clk(gclk));
	jdff dff_B_UrvDxQ9U4_2(.din(w_dff_B_GomBGRAp5_2),.dout(w_dff_B_UrvDxQ9U4_2),.clk(gclk));
	jdff dff_B_WAhhwlNj0_2(.din(n1002),.dout(w_dff_B_WAhhwlNj0_2),.clk(gclk));
	jdff dff_B_ES8A9qFY2_1(.din(n930),.dout(w_dff_B_ES8A9qFY2_1),.clk(gclk));
	jdff dff_B_4OKM4cKp7_2(.din(n827),.dout(w_dff_B_4OKM4cKp7_2),.clk(gclk));
	jdff dff_B_GdG1bUWr0_2(.din(w_dff_B_4OKM4cKp7_2),.dout(w_dff_B_GdG1bUWr0_2),.clk(gclk));
	jdff dff_B_McEmyvUX2_2(.din(w_dff_B_GdG1bUWr0_2),.dout(w_dff_B_McEmyvUX2_2),.clk(gclk));
	jdff dff_B_a60qLhFd6_2(.din(w_dff_B_McEmyvUX2_2),.dout(w_dff_B_a60qLhFd6_2),.clk(gclk));
	jdff dff_B_YzeipnX85_2(.din(w_dff_B_a60qLhFd6_2),.dout(w_dff_B_YzeipnX85_2),.clk(gclk));
	jdff dff_B_lR4kSvH20_2(.din(w_dff_B_YzeipnX85_2),.dout(w_dff_B_lR4kSvH20_2),.clk(gclk));
	jdff dff_B_ndTj5aDB8_2(.din(w_dff_B_lR4kSvH20_2),.dout(w_dff_B_ndTj5aDB8_2),.clk(gclk));
	jdff dff_B_PAyzfLUT1_2(.din(w_dff_B_ndTj5aDB8_2),.dout(w_dff_B_PAyzfLUT1_2),.clk(gclk));
	jdff dff_B_g7jmvIFk6_2(.din(w_dff_B_PAyzfLUT1_2),.dout(w_dff_B_g7jmvIFk6_2),.clk(gclk));
	jdff dff_B_zoISVPjS2_2(.din(w_dff_B_g7jmvIFk6_2),.dout(w_dff_B_zoISVPjS2_2),.clk(gclk));
	jdff dff_B_PTJKGiy70_2(.din(w_dff_B_zoISVPjS2_2),.dout(w_dff_B_PTJKGiy70_2),.clk(gclk));
	jdff dff_B_Dp89tbBr2_2(.din(w_dff_B_PTJKGiy70_2),.dout(w_dff_B_Dp89tbBr2_2),.clk(gclk));
	jdff dff_B_u3fV66GJ7_2(.din(w_dff_B_Dp89tbBr2_2),.dout(w_dff_B_u3fV66GJ7_2),.clk(gclk));
	jdff dff_B_9H44FkjQ5_2(.din(w_dff_B_u3fV66GJ7_2),.dout(w_dff_B_9H44FkjQ5_2),.clk(gclk));
	jdff dff_B_b8HlkuWd3_2(.din(w_dff_B_9H44FkjQ5_2),.dout(w_dff_B_b8HlkuWd3_2),.clk(gclk));
	jdff dff_B_7sLHKdh51_2(.din(w_dff_B_b8HlkuWd3_2),.dout(w_dff_B_7sLHKdh51_2),.clk(gclk));
	jdff dff_B_XBBSYOyr6_2(.din(w_dff_B_7sLHKdh51_2),.dout(w_dff_B_XBBSYOyr6_2),.clk(gclk));
	jdff dff_B_AUNKYcOn9_2(.din(w_dff_B_XBBSYOyr6_2),.dout(w_dff_B_AUNKYcOn9_2),.clk(gclk));
	jdff dff_B_wAtPlfI39_2(.din(w_dff_B_AUNKYcOn9_2),.dout(w_dff_B_wAtPlfI39_2),.clk(gclk));
	jdff dff_B_25t42bdX4_2(.din(w_dff_B_wAtPlfI39_2),.dout(w_dff_B_25t42bdX4_2),.clk(gclk));
	jdff dff_B_gKD0Gxe66_2(.din(w_dff_B_25t42bdX4_2),.dout(w_dff_B_gKD0Gxe66_2),.clk(gclk));
	jdff dff_B_jFZoaqyw7_2(.din(w_dff_B_gKD0Gxe66_2),.dout(w_dff_B_jFZoaqyw7_2),.clk(gclk));
	jdff dff_B_HWCxjJ2i0_2(.din(w_dff_B_jFZoaqyw7_2),.dout(w_dff_B_HWCxjJ2i0_2),.clk(gclk));
	jdff dff_B_HvlRzSII5_2(.din(w_dff_B_HWCxjJ2i0_2),.dout(w_dff_B_HvlRzSII5_2),.clk(gclk));
	jdff dff_B_Eq8k8tt39_2(.din(w_dff_B_HvlRzSII5_2),.dout(w_dff_B_Eq8k8tt39_2),.clk(gclk));
	jdff dff_B_25aefGon7_2(.din(w_dff_B_Eq8k8tt39_2),.dout(w_dff_B_25aefGon7_2),.clk(gclk));
	jdff dff_B_UqxYYvQe9_2(.din(w_dff_B_25aefGon7_2),.dout(w_dff_B_UqxYYvQe9_2),.clk(gclk));
	jdff dff_B_psQDKeQz4_2(.din(w_dff_B_UqxYYvQe9_2),.dout(w_dff_B_psQDKeQz4_2),.clk(gclk));
	jdff dff_B_zpf0RMsl6_2(.din(w_dff_B_psQDKeQz4_2),.dout(w_dff_B_zpf0RMsl6_2),.clk(gclk));
	jdff dff_B_QxodiXm21_2(.din(w_dff_B_zpf0RMsl6_2),.dout(w_dff_B_QxodiXm21_2),.clk(gclk));
	jdff dff_B_J1SboDT76_2(.din(n896),.dout(w_dff_B_J1SboDT76_2),.clk(gclk));
	jdff dff_B_BEvijuvY2_1(.din(n828),.dout(w_dff_B_BEvijuvY2_1),.clk(gclk));
	jdff dff_B_GQ3QdFvL0_2(.din(n729),.dout(w_dff_B_GQ3QdFvL0_2),.clk(gclk));
	jdff dff_B_HFHh5zsi0_2(.din(w_dff_B_GQ3QdFvL0_2),.dout(w_dff_B_HFHh5zsi0_2),.clk(gclk));
	jdff dff_B_aF7loKUi6_2(.din(w_dff_B_HFHh5zsi0_2),.dout(w_dff_B_aF7loKUi6_2),.clk(gclk));
	jdff dff_B_yefhpsUQ8_2(.din(w_dff_B_aF7loKUi6_2),.dout(w_dff_B_yefhpsUQ8_2),.clk(gclk));
	jdff dff_B_AetPeZ4R5_2(.din(w_dff_B_yefhpsUQ8_2),.dout(w_dff_B_AetPeZ4R5_2),.clk(gclk));
	jdff dff_B_XXOV84DU6_2(.din(w_dff_B_AetPeZ4R5_2),.dout(w_dff_B_XXOV84DU6_2),.clk(gclk));
	jdff dff_B_B9Vgeurz8_2(.din(w_dff_B_XXOV84DU6_2),.dout(w_dff_B_B9Vgeurz8_2),.clk(gclk));
	jdff dff_B_cFhCzb1c5_2(.din(w_dff_B_B9Vgeurz8_2),.dout(w_dff_B_cFhCzb1c5_2),.clk(gclk));
	jdff dff_B_bHTPZ83v2_2(.din(w_dff_B_cFhCzb1c5_2),.dout(w_dff_B_bHTPZ83v2_2),.clk(gclk));
	jdff dff_B_7V3YVRwD4_2(.din(w_dff_B_bHTPZ83v2_2),.dout(w_dff_B_7V3YVRwD4_2),.clk(gclk));
	jdff dff_B_jrhUNSGX5_2(.din(w_dff_B_7V3YVRwD4_2),.dout(w_dff_B_jrhUNSGX5_2),.clk(gclk));
	jdff dff_B_HhUXOQlg9_2(.din(w_dff_B_jrhUNSGX5_2),.dout(w_dff_B_HhUXOQlg9_2),.clk(gclk));
	jdff dff_B_BcdhCkD81_2(.din(w_dff_B_HhUXOQlg9_2),.dout(w_dff_B_BcdhCkD81_2),.clk(gclk));
	jdff dff_B_NzrZNvWT0_2(.din(w_dff_B_BcdhCkD81_2),.dout(w_dff_B_NzrZNvWT0_2),.clk(gclk));
	jdff dff_B_V5hvzjcu8_2(.din(w_dff_B_NzrZNvWT0_2),.dout(w_dff_B_V5hvzjcu8_2),.clk(gclk));
	jdff dff_B_U0ueuIPn1_2(.din(w_dff_B_V5hvzjcu8_2),.dout(w_dff_B_U0ueuIPn1_2),.clk(gclk));
	jdff dff_B_kW9adihj2_2(.din(w_dff_B_U0ueuIPn1_2),.dout(w_dff_B_kW9adihj2_2),.clk(gclk));
	jdff dff_B_obvdkl5p8_2(.din(w_dff_B_kW9adihj2_2),.dout(w_dff_B_obvdkl5p8_2),.clk(gclk));
	jdff dff_B_a42tlBsV7_2(.din(w_dff_B_obvdkl5p8_2),.dout(w_dff_B_a42tlBsV7_2),.clk(gclk));
	jdff dff_B_nJmuKdlf0_2(.din(w_dff_B_a42tlBsV7_2),.dout(w_dff_B_nJmuKdlf0_2),.clk(gclk));
	jdff dff_B_IRynea0h1_2(.din(w_dff_B_nJmuKdlf0_2),.dout(w_dff_B_IRynea0h1_2),.clk(gclk));
	jdff dff_B_KwqeBfpv8_2(.din(w_dff_B_IRynea0h1_2),.dout(w_dff_B_KwqeBfpv8_2),.clk(gclk));
	jdff dff_B_8FlsdvU64_2(.din(w_dff_B_KwqeBfpv8_2),.dout(w_dff_B_8FlsdvU64_2),.clk(gclk));
	jdff dff_B_rfX2w4o63_2(.din(w_dff_B_8FlsdvU64_2),.dout(w_dff_B_rfX2w4o63_2),.clk(gclk));
	jdff dff_B_7jqHOznN0_2(.din(w_dff_B_rfX2w4o63_2),.dout(w_dff_B_7jqHOznN0_2),.clk(gclk));
	jdff dff_B_UtuN7ZTW3_2(.din(w_dff_B_7jqHOznN0_2),.dout(w_dff_B_UtuN7ZTW3_2),.clk(gclk));
	jdff dff_B_hrcXJnDK9_2(.din(w_dff_B_UtuN7ZTW3_2),.dout(w_dff_B_hrcXJnDK9_2),.clk(gclk));
	jdff dff_B_svrYkw6u9_2(.din(n793),.dout(w_dff_B_svrYkw6u9_2),.clk(gclk));
	jdff dff_B_FXe6CwUR4_1(.din(n730),.dout(w_dff_B_FXe6CwUR4_1),.clk(gclk));
	jdff dff_B_t1XBVJht3_2(.din(n637),.dout(w_dff_B_t1XBVJht3_2),.clk(gclk));
	jdff dff_B_rSySyf5D7_2(.din(w_dff_B_t1XBVJht3_2),.dout(w_dff_B_rSySyf5D7_2),.clk(gclk));
	jdff dff_B_iks8NdLb4_2(.din(w_dff_B_rSySyf5D7_2),.dout(w_dff_B_iks8NdLb4_2),.clk(gclk));
	jdff dff_B_ViliiN2U3_2(.din(w_dff_B_iks8NdLb4_2),.dout(w_dff_B_ViliiN2U3_2),.clk(gclk));
	jdff dff_B_gEyCpVS98_2(.din(w_dff_B_ViliiN2U3_2),.dout(w_dff_B_gEyCpVS98_2),.clk(gclk));
	jdff dff_B_qozLjBPJ2_2(.din(w_dff_B_gEyCpVS98_2),.dout(w_dff_B_qozLjBPJ2_2),.clk(gclk));
	jdff dff_B_61jcc8J72_2(.din(w_dff_B_qozLjBPJ2_2),.dout(w_dff_B_61jcc8J72_2),.clk(gclk));
	jdff dff_B_wcCzGFN59_2(.din(w_dff_B_61jcc8J72_2),.dout(w_dff_B_wcCzGFN59_2),.clk(gclk));
	jdff dff_B_RUamuXrZ0_2(.din(w_dff_B_wcCzGFN59_2),.dout(w_dff_B_RUamuXrZ0_2),.clk(gclk));
	jdff dff_B_X7mtnsEN2_2(.din(w_dff_B_RUamuXrZ0_2),.dout(w_dff_B_X7mtnsEN2_2),.clk(gclk));
	jdff dff_B_sEaYM43W3_2(.din(w_dff_B_X7mtnsEN2_2),.dout(w_dff_B_sEaYM43W3_2),.clk(gclk));
	jdff dff_B_JpJF7PRE8_2(.din(w_dff_B_sEaYM43W3_2),.dout(w_dff_B_JpJF7PRE8_2),.clk(gclk));
	jdff dff_B_xdYxnhQO8_2(.din(w_dff_B_JpJF7PRE8_2),.dout(w_dff_B_xdYxnhQO8_2),.clk(gclk));
	jdff dff_B_nRnL4E6W4_2(.din(w_dff_B_xdYxnhQO8_2),.dout(w_dff_B_nRnL4E6W4_2),.clk(gclk));
	jdff dff_B_lSIZ6eIi9_2(.din(w_dff_B_nRnL4E6W4_2),.dout(w_dff_B_lSIZ6eIi9_2),.clk(gclk));
	jdff dff_B_zlKdYJbH3_2(.din(w_dff_B_lSIZ6eIi9_2),.dout(w_dff_B_zlKdYJbH3_2),.clk(gclk));
	jdff dff_B_m1YmdJ9t1_2(.din(w_dff_B_zlKdYJbH3_2),.dout(w_dff_B_m1YmdJ9t1_2),.clk(gclk));
	jdff dff_B_0MKCJrkr1_2(.din(w_dff_B_m1YmdJ9t1_2),.dout(w_dff_B_0MKCJrkr1_2),.clk(gclk));
	jdff dff_B_jLR83C9x0_2(.din(w_dff_B_0MKCJrkr1_2),.dout(w_dff_B_jLR83C9x0_2),.clk(gclk));
	jdff dff_B_Qn3XVrj43_2(.din(w_dff_B_jLR83C9x0_2),.dout(w_dff_B_Qn3XVrj43_2),.clk(gclk));
	jdff dff_B_5EVpO9IP8_2(.din(w_dff_B_Qn3XVrj43_2),.dout(w_dff_B_5EVpO9IP8_2),.clk(gclk));
	jdff dff_B_6p0ufAyi4_2(.din(w_dff_B_5EVpO9IP8_2),.dout(w_dff_B_6p0ufAyi4_2),.clk(gclk));
	jdff dff_B_c3qKAM3p1_2(.din(w_dff_B_6p0ufAyi4_2),.dout(w_dff_B_c3qKAM3p1_2),.clk(gclk));
	jdff dff_B_96dG2lku2_2(.din(w_dff_B_c3qKAM3p1_2),.dout(w_dff_B_96dG2lku2_2),.clk(gclk));
	jdff dff_B_uPSobetU8_2(.din(n694),.dout(w_dff_B_uPSobetU8_2),.clk(gclk));
	jdff dff_B_1euSCDwy0_1(.din(n638),.dout(w_dff_B_1euSCDwy0_1),.clk(gclk));
	jdff dff_B_jdaWrV129_2(.din(n552),.dout(w_dff_B_jdaWrV129_2),.clk(gclk));
	jdff dff_B_Ws6j2AqG6_2(.din(w_dff_B_jdaWrV129_2),.dout(w_dff_B_Ws6j2AqG6_2),.clk(gclk));
	jdff dff_B_JEHKea2e6_2(.din(w_dff_B_Ws6j2AqG6_2),.dout(w_dff_B_JEHKea2e6_2),.clk(gclk));
	jdff dff_B_46kIN4dJ8_2(.din(w_dff_B_JEHKea2e6_2),.dout(w_dff_B_46kIN4dJ8_2),.clk(gclk));
	jdff dff_B_tEth13KY7_2(.din(w_dff_B_46kIN4dJ8_2),.dout(w_dff_B_tEth13KY7_2),.clk(gclk));
	jdff dff_B_BlB4pSDy7_2(.din(w_dff_B_tEth13KY7_2),.dout(w_dff_B_BlB4pSDy7_2),.clk(gclk));
	jdff dff_B_aomaS7Ha4_2(.din(w_dff_B_BlB4pSDy7_2),.dout(w_dff_B_aomaS7Ha4_2),.clk(gclk));
	jdff dff_B_opUpP3oK8_2(.din(w_dff_B_aomaS7Ha4_2),.dout(w_dff_B_opUpP3oK8_2),.clk(gclk));
	jdff dff_B_r8wvA1h25_2(.din(w_dff_B_opUpP3oK8_2),.dout(w_dff_B_r8wvA1h25_2),.clk(gclk));
	jdff dff_B_P0oLKxNr5_2(.din(w_dff_B_r8wvA1h25_2),.dout(w_dff_B_P0oLKxNr5_2),.clk(gclk));
	jdff dff_B_yTXSK4yW0_2(.din(w_dff_B_P0oLKxNr5_2),.dout(w_dff_B_yTXSK4yW0_2),.clk(gclk));
	jdff dff_B_2UHkJSm74_2(.din(w_dff_B_yTXSK4yW0_2),.dout(w_dff_B_2UHkJSm74_2),.clk(gclk));
	jdff dff_B_nzMkGFDw9_2(.din(w_dff_B_2UHkJSm74_2),.dout(w_dff_B_nzMkGFDw9_2),.clk(gclk));
	jdff dff_B_QyOBWDvR4_2(.din(w_dff_B_nzMkGFDw9_2),.dout(w_dff_B_QyOBWDvR4_2),.clk(gclk));
	jdff dff_B_PvIhAwNA1_2(.din(w_dff_B_QyOBWDvR4_2),.dout(w_dff_B_PvIhAwNA1_2),.clk(gclk));
	jdff dff_B_6f40NG5z5_2(.din(w_dff_B_PvIhAwNA1_2),.dout(w_dff_B_6f40NG5z5_2),.clk(gclk));
	jdff dff_B_b5xwAwts8_2(.din(w_dff_B_6f40NG5z5_2),.dout(w_dff_B_b5xwAwts8_2),.clk(gclk));
	jdff dff_B_mu7wUGIp4_2(.din(w_dff_B_b5xwAwts8_2),.dout(w_dff_B_mu7wUGIp4_2),.clk(gclk));
	jdff dff_B_OmTfFvBC3_2(.din(w_dff_B_mu7wUGIp4_2),.dout(w_dff_B_OmTfFvBC3_2),.clk(gclk));
	jdff dff_B_se3F7SJA5_2(.din(w_dff_B_OmTfFvBC3_2),.dout(w_dff_B_se3F7SJA5_2),.clk(gclk));
	jdff dff_B_QQcdNQza5_2(.din(w_dff_B_se3F7SJA5_2),.dout(w_dff_B_QQcdNQza5_2),.clk(gclk));
	jdff dff_B_lgr9fuJH8_2(.din(n602),.dout(w_dff_B_lgr9fuJH8_2),.clk(gclk));
	jdff dff_B_uy2SawVe8_1(.din(n553),.dout(w_dff_B_uy2SawVe8_1),.clk(gclk));
	jdff dff_B_vzemtAjL1_2(.din(n474),.dout(w_dff_B_vzemtAjL1_2),.clk(gclk));
	jdff dff_B_yFFYn2TD0_2(.din(w_dff_B_vzemtAjL1_2),.dout(w_dff_B_yFFYn2TD0_2),.clk(gclk));
	jdff dff_B_snmph6z98_2(.din(w_dff_B_yFFYn2TD0_2),.dout(w_dff_B_snmph6z98_2),.clk(gclk));
	jdff dff_B_sy3F2kV40_2(.din(w_dff_B_snmph6z98_2),.dout(w_dff_B_sy3F2kV40_2),.clk(gclk));
	jdff dff_B_qUdlNRve4_2(.din(w_dff_B_sy3F2kV40_2),.dout(w_dff_B_qUdlNRve4_2),.clk(gclk));
	jdff dff_B_hSyDXdHs6_2(.din(w_dff_B_qUdlNRve4_2),.dout(w_dff_B_hSyDXdHs6_2),.clk(gclk));
	jdff dff_B_zCYVFSva2_2(.din(w_dff_B_hSyDXdHs6_2),.dout(w_dff_B_zCYVFSva2_2),.clk(gclk));
	jdff dff_B_ovYZAF3U1_2(.din(w_dff_B_zCYVFSva2_2),.dout(w_dff_B_ovYZAF3U1_2),.clk(gclk));
	jdff dff_B_k47Nm3CI9_2(.din(w_dff_B_ovYZAF3U1_2),.dout(w_dff_B_k47Nm3CI9_2),.clk(gclk));
	jdff dff_B_iVMjVeeL9_2(.din(w_dff_B_k47Nm3CI9_2),.dout(w_dff_B_iVMjVeeL9_2),.clk(gclk));
	jdff dff_B_CfPIXJVu3_2(.din(w_dff_B_iVMjVeeL9_2),.dout(w_dff_B_CfPIXJVu3_2),.clk(gclk));
	jdff dff_B_77beoL2m7_2(.din(w_dff_B_CfPIXJVu3_2),.dout(w_dff_B_77beoL2m7_2),.clk(gclk));
	jdff dff_B_DSJn62HN1_2(.din(w_dff_B_77beoL2m7_2),.dout(w_dff_B_DSJn62HN1_2),.clk(gclk));
	jdff dff_B_laxTxQlK7_2(.din(w_dff_B_DSJn62HN1_2),.dout(w_dff_B_laxTxQlK7_2),.clk(gclk));
	jdff dff_B_V24fdcLu1_2(.din(w_dff_B_laxTxQlK7_2),.dout(w_dff_B_V24fdcLu1_2),.clk(gclk));
	jdff dff_B_5HOpSRCc4_2(.din(w_dff_B_V24fdcLu1_2),.dout(w_dff_B_5HOpSRCc4_2),.clk(gclk));
	jdff dff_B_k32OGgPv5_2(.din(w_dff_B_5HOpSRCc4_2),.dout(w_dff_B_k32OGgPv5_2),.clk(gclk));
	jdff dff_B_oIoefvFy9_2(.din(w_dff_B_k32OGgPv5_2),.dout(w_dff_B_oIoefvFy9_2),.clk(gclk));
	jdff dff_B_nZJmTAnu1_2(.din(n517),.dout(w_dff_B_nZJmTAnu1_2),.clk(gclk));
	jdff dff_B_GXqD2o435_1(.din(n475),.dout(w_dff_B_GXqD2o435_1),.clk(gclk));
	jdff dff_B_yQWoVcq78_2(.din(n403),.dout(w_dff_B_yQWoVcq78_2),.clk(gclk));
	jdff dff_B_OzxQIpyc3_2(.din(w_dff_B_yQWoVcq78_2),.dout(w_dff_B_OzxQIpyc3_2),.clk(gclk));
	jdff dff_B_bwWGxP5g0_2(.din(w_dff_B_OzxQIpyc3_2),.dout(w_dff_B_bwWGxP5g0_2),.clk(gclk));
	jdff dff_B_b5ciOZUC7_2(.din(w_dff_B_bwWGxP5g0_2),.dout(w_dff_B_b5ciOZUC7_2),.clk(gclk));
	jdff dff_B_jFdfFPbR8_2(.din(w_dff_B_b5ciOZUC7_2),.dout(w_dff_B_jFdfFPbR8_2),.clk(gclk));
	jdff dff_B_yj84MG5C4_2(.din(w_dff_B_jFdfFPbR8_2),.dout(w_dff_B_yj84MG5C4_2),.clk(gclk));
	jdff dff_B_ZnmMV5Gk3_2(.din(w_dff_B_yj84MG5C4_2),.dout(w_dff_B_ZnmMV5Gk3_2),.clk(gclk));
	jdff dff_B_BVD23hxG1_2(.din(w_dff_B_ZnmMV5Gk3_2),.dout(w_dff_B_BVD23hxG1_2),.clk(gclk));
	jdff dff_B_9ZRrLiv72_2(.din(w_dff_B_BVD23hxG1_2),.dout(w_dff_B_9ZRrLiv72_2),.clk(gclk));
	jdff dff_B_MtSGdIjF2_2(.din(w_dff_B_9ZRrLiv72_2),.dout(w_dff_B_MtSGdIjF2_2),.clk(gclk));
	jdff dff_B_IKjg6YUZ9_2(.din(w_dff_B_MtSGdIjF2_2),.dout(w_dff_B_IKjg6YUZ9_2),.clk(gclk));
	jdff dff_B_HRceJayX3_2(.din(w_dff_B_IKjg6YUZ9_2),.dout(w_dff_B_HRceJayX3_2),.clk(gclk));
	jdff dff_B_IVbcteM63_2(.din(w_dff_B_HRceJayX3_2),.dout(w_dff_B_IVbcteM63_2),.clk(gclk));
	jdff dff_B_SsTK8xTm0_2(.din(w_dff_B_IVbcteM63_2),.dout(w_dff_B_SsTK8xTm0_2),.clk(gclk));
	jdff dff_B_xobzKttg0_2(.din(w_dff_B_SsTK8xTm0_2),.dout(w_dff_B_xobzKttg0_2),.clk(gclk));
	jdff dff_B_Ef1UaLVG5_2(.din(n439),.dout(w_dff_B_Ef1UaLVG5_2),.clk(gclk));
	jdff dff_B_hSfTyuhW6_1(.din(n404),.dout(w_dff_B_hSfTyuhW6_1),.clk(gclk));
	jdff dff_B_PWQJ2Vnu3_2(.din(n340),.dout(w_dff_B_PWQJ2Vnu3_2),.clk(gclk));
	jdff dff_B_6B2YF9Ay1_2(.din(w_dff_B_PWQJ2Vnu3_2),.dout(w_dff_B_6B2YF9Ay1_2),.clk(gclk));
	jdff dff_B_y9ktx8Jb5_2(.din(w_dff_B_6B2YF9Ay1_2),.dout(w_dff_B_y9ktx8Jb5_2),.clk(gclk));
	jdff dff_B_rjQWH52K2_2(.din(w_dff_B_y9ktx8Jb5_2),.dout(w_dff_B_rjQWH52K2_2),.clk(gclk));
	jdff dff_B_KQm4MA0M9_2(.din(w_dff_B_rjQWH52K2_2),.dout(w_dff_B_KQm4MA0M9_2),.clk(gclk));
	jdff dff_B_gxsauXrw9_2(.din(w_dff_B_KQm4MA0M9_2),.dout(w_dff_B_gxsauXrw9_2),.clk(gclk));
	jdff dff_B_AjTY6Lo33_2(.din(w_dff_B_gxsauXrw9_2),.dout(w_dff_B_AjTY6Lo33_2),.clk(gclk));
	jdff dff_B_r84F0BXi2_2(.din(w_dff_B_AjTY6Lo33_2),.dout(w_dff_B_r84F0BXi2_2),.clk(gclk));
	jdff dff_B_BVhpNlmg8_2(.din(w_dff_B_r84F0BXi2_2),.dout(w_dff_B_BVhpNlmg8_2),.clk(gclk));
	jdff dff_B_1ZNcWDTJ4_2(.din(w_dff_B_BVhpNlmg8_2),.dout(w_dff_B_1ZNcWDTJ4_2),.clk(gclk));
	jdff dff_B_U1GybGGG9_2(.din(w_dff_B_1ZNcWDTJ4_2),.dout(w_dff_B_U1GybGGG9_2),.clk(gclk));
	jdff dff_B_b8fAa6Jb0_2(.din(w_dff_B_U1GybGGG9_2),.dout(w_dff_B_b8fAa6Jb0_2),.clk(gclk));
	jdff dff_B_IE4fTbbZ3_2(.din(n368),.dout(w_dff_B_IE4fTbbZ3_2),.clk(gclk));
	jdff dff_B_TBd7wztu5_1(.din(n341),.dout(w_dff_B_TBd7wztu5_1),.clk(gclk));
	jdff dff_B_nNKdS2049_2(.din(n284),.dout(w_dff_B_nNKdS2049_2),.clk(gclk));
	jdff dff_B_NURwZw7z5_2(.din(w_dff_B_nNKdS2049_2),.dout(w_dff_B_NURwZw7z5_2),.clk(gclk));
	jdff dff_B_zQUzFn1p0_2(.din(w_dff_B_NURwZw7z5_2),.dout(w_dff_B_zQUzFn1p0_2),.clk(gclk));
	jdff dff_B_7SibxeSs7_2(.din(w_dff_B_zQUzFn1p0_2),.dout(w_dff_B_7SibxeSs7_2),.clk(gclk));
	jdff dff_B_m9aJIOKE2_2(.din(w_dff_B_7SibxeSs7_2),.dout(w_dff_B_m9aJIOKE2_2),.clk(gclk));
	jdff dff_B_a0Se4UDH4_2(.din(w_dff_B_m9aJIOKE2_2),.dout(w_dff_B_a0Se4UDH4_2),.clk(gclk));
	jdff dff_B_V96D4y7W9_2(.din(w_dff_B_a0Se4UDH4_2),.dout(w_dff_B_V96D4y7W9_2),.clk(gclk));
	jdff dff_B_Y6VQH7IZ4_2(.din(w_dff_B_V96D4y7W9_2),.dout(w_dff_B_Y6VQH7IZ4_2),.clk(gclk));
	jdff dff_B_CbvTIG0O8_2(.din(w_dff_B_Y6VQH7IZ4_2),.dout(w_dff_B_CbvTIG0O8_2),.clk(gclk));
	jdff dff_B_n3Z6e0v41_2(.din(n305),.dout(w_dff_B_n3Z6e0v41_2),.clk(gclk));
	jdff dff_B_YoDQV3J86_1(.din(n285),.dout(w_dff_B_YoDQV3J86_1),.clk(gclk));
	jdff dff_B_GbOS7NLd1_2(.din(n235),.dout(w_dff_B_GbOS7NLd1_2),.clk(gclk));
	jdff dff_B_WQnTFrOB2_2(.din(w_dff_B_GbOS7NLd1_2),.dout(w_dff_B_WQnTFrOB2_2),.clk(gclk));
	jdff dff_B_Wors72lZ0_2(.din(w_dff_B_WQnTFrOB2_2),.dout(w_dff_B_Wors72lZ0_2),.clk(gclk));
	jdff dff_B_X0ggv1W10_2(.din(w_dff_B_Wors72lZ0_2),.dout(w_dff_B_X0ggv1W10_2),.clk(gclk));
	jdff dff_B_GkuqroHq8_2(.din(w_dff_B_X0ggv1W10_2),.dout(w_dff_B_GkuqroHq8_2),.clk(gclk));
	jdff dff_B_7mP3ZrFy4_2(.din(w_dff_B_GkuqroHq8_2),.dout(w_dff_B_7mP3ZrFy4_2),.clk(gclk));
	jdff dff_B_6moYWDCl8_2(.din(n249),.dout(w_dff_B_6moYWDCl8_2),.clk(gclk));
	jdff dff_B_tLxctWia2_2(.din(n194),.dout(w_dff_B_tLxctWia2_2),.clk(gclk));
	jdff dff_B_epZiYMrb5_2(.din(w_dff_B_tLxctWia2_2),.dout(w_dff_B_epZiYMrb5_2),.clk(gclk));
	jdff dff_B_5j9PqDcD1_2(.din(w_dff_B_epZiYMrb5_2),.dout(w_dff_B_5j9PqDcD1_2),.clk(gclk));
	jdff dff_B_vi41Mh5Q9_0(.din(n199),.dout(w_dff_B_vi41Mh5Q9_0),.clk(gclk));
	jdff dff_A_T32BztU16_0(.dout(w_n157_0[0]),.din(w_dff_A_T32BztU16_0),.clk(gclk));
	jdff dff_A_Rg6AGHtF7_0(.dout(w_dff_A_T32BztU16_0),.din(w_dff_A_Rg6AGHtF7_0),.clk(gclk));
	jdff dff_A_5EX1W2hZ4_0(.dout(w_n156_0[0]),.din(w_dff_A_5EX1W2hZ4_0),.clk(gclk));
	jdff dff_A_nGqydeaL0_0(.dout(w_dff_A_5EX1W2hZ4_0),.din(w_dff_A_nGqydeaL0_0),.clk(gclk));
	jdff dff_B_HsitQwma1_2(.din(n1389),.dout(w_dff_B_HsitQwma1_2),.clk(gclk));
	jdff dff_B_3Elpi5LQ4_1(.din(n1387),.dout(w_dff_B_3Elpi5LQ4_1),.clk(gclk));
	jdff dff_B_DRYQFlrp3_2(.din(n1307),.dout(w_dff_B_DRYQFlrp3_2),.clk(gclk));
	jdff dff_B_Gl0SiJCf0_2(.din(w_dff_B_DRYQFlrp3_2),.dout(w_dff_B_Gl0SiJCf0_2),.clk(gclk));
	jdff dff_B_SVeeDJSP8_2(.din(w_dff_B_Gl0SiJCf0_2),.dout(w_dff_B_SVeeDJSP8_2),.clk(gclk));
	jdff dff_B_C6iZAuX13_2(.din(w_dff_B_SVeeDJSP8_2),.dout(w_dff_B_C6iZAuX13_2),.clk(gclk));
	jdff dff_B_3IYusue31_2(.din(w_dff_B_C6iZAuX13_2),.dout(w_dff_B_3IYusue31_2),.clk(gclk));
	jdff dff_B_dEEzoEfp9_2(.din(w_dff_B_3IYusue31_2),.dout(w_dff_B_dEEzoEfp9_2),.clk(gclk));
	jdff dff_B_jrBR3hNx5_2(.din(w_dff_B_dEEzoEfp9_2),.dout(w_dff_B_jrBR3hNx5_2),.clk(gclk));
	jdff dff_B_TD39RoJ25_2(.din(w_dff_B_jrBR3hNx5_2),.dout(w_dff_B_TD39RoJ25_2),.clk(gclk));
	jdff dff_B_xE9dR0lx5_2(.din(w_dff_B_TD39RoJ25_2),.dout(w_dff_B_xE9dR0lx5_2),.clk(gclk));
	jdff dff_B_EgN0PYJT6_2(.din(w_dff_B_xE9dR0lx5_2),.dout(w_dff_B_EgN0PYJT6_2),.clk(gclk));
	jdff dff_B_zAIScBcD5_2(.din(w_dff_B_EgN0PYJT6_2),.dout(w_dff_B_zAIScBcD5_2),.clk(gclk));
	jdff dff_B_KgskRtnN4_2(.din(w_dff_B_zAIScBcD5_2),.dout(w_dff_B_KgskRtnN4_2),.clk(gclk));
	jdff dff_B_fsM45eLY9_2(.din(w_dff_B_KgskRtnN4_2),.dout(w_dff_B_fsM45eLY9_2),.clk(gclk));
	jdff dff_B_fbwW3KCr9_2(.din(w_dff_B_fsM45eLY9_2),.dout(w_dff_B_fbwW3KCr9_2),.clk(gclk));
	jdff dff_B_GiWfCGXA7_2(.din(w_dff_B_fbwW3KCr9_2),.dout(w_dff_B_GiWfCGXA7_2),.clk(gclk));
	jdff dff_B_hHjCLsR01_2(.din(w_dff_B_GiWfCGXA7_2),.dout(w_dff_B_hHjCLsR01_2),.clk(gclk));
	jdff dff_B_cJtUaC1u5_2(.din(w_dff_B_hHjCLsR01_2),.dout(w_dff_B_cJtUaC1u5_2),.clk(gclk));
	jdff dff_B_dgkr1E9x4_2(.din(w_dff_B_cJtUaC1u5_2),.dout(w_dff_B_dgkr1E9x4_2),.clk(gclk));
	jdff dff_B_VBvgpe0w2_2(.din(w_dff_B_dgkr1E9x4_2),.dout(w_dff_B_VBvgpe0w2_2),.clk(gclk));
	jdff dff_B_K0Mn1GUF2_2(.din(w_dff_B_VBvgpe0w2_2),.dout(w_dff_B_K0Mn1GUF2_2),.clk(gclk));
	jdff dff_B_TgK9lkI00_2(.din(w_dff_B_K0Mn1GUF2_2),.dout(w_dff_B_TgK9lkI00_2),.clk(gclk));
	jdff dff_B_D3UkFlhV2_2(.din(w_dff_B_TgK9lkI00_2),.dout(w_dff_B_D3UkFlhV2_2),.clk(gclk));
	jdff dff_B_X8FVcDj51_2(.din(w_dff_B_D3UkFlhV2_2),.dout(w_dff_B_X8FVcDj51_2),.clk(gclk));
	jdff dff_B_elgSfL0S3_2(.din(w_dff_B_X8FVcDj51_2),.dout(w_dff_B_elgSfL0S3_2),.clk(gclk));
	jdff dff_B_IR3vG3Zu1_2(.din(w_dff_B_elgSfL0S3_2),.dout(w_dff_B_IR3vG3Zu1_2),.clk(gclk));
	jdff dff_B_aWCy2cF89_2(.din(w_dff_B_IR3vG3Zu1_2),.dout(w_dff_B_aWCy2cF89_2),.clk(gclk));
	jdff dff_B_SoLQ3Xav9_2(.din(w_dff_B_aWCy2cF89_2),.dout(w_dff_B_SoLQ3Xav9_2),.clk(gclk));
	jdff dff_B_ezl1TwEr2_2(.din(w_dff_B_SoLQ3Xav9_2),.dout(w_dff_B_ezl1TwEr2_2),.clk(gclk));
	jdff dff_B_You15Nnr4_2(.din(w_dff_B_ezl1TwEr2_2),.dout(w_dff_B_You15Nnr4_2),.clk(gclk));
	jdff dff_B_Vl6gXDkl3_2(.din(w_dff_B_You15Nnr4_2),.dout(w_dff_B_Vl6gXDkl3_2),.clk(gclk));
	jdff dff_B_w4nqc8XN4_2(.din(w_dff_B_Vl6gXDkl3_2),.dout(w_dff_B_w4nqc8XN4_2),.clk(gclk));
	jdff dff_B_rIxlfcrw2_2(.din(w_dff_B_w4nqc8XN4_2),.dout(w_dff_B_rIxlfcrw2_2),.clk(gclk));
	jdff dff_B_YEzMr56n5_2(.din(w_dff_B_rIxlfcrw2_2),.dout(w_dff_B_YEzMr56n5_2),.clk(gclk));
	jdff dff_B_Kwqoe2np4_2(.din(w_dff_B_YEzMr56n5_2),.dout(w_dff_B_Kwqoe2np4_2),.clk(gclk));
	jdff dff_B_XzqoWY2q4_2(.din(w_dff_B_Kwqoe2np4_2),.dout(w_dff_B_XzqoWY2q4_2),.clk(gclk));
	jdff dff_B_N2nn0n0g0_2(.din(w_dff_B_XzqoWY2q4_2),.dout(w_dff_B_N2nn0n0g0_2),.clk(gclk));
	jdff dff_B_oybLVK4D8_2(.din(w_dff_B_N2nn0n0g0_2),.dout(w_dff_B_oybLVK4D8_2),.clk(gclk));
	jdff dff_B_izwdhGDY8_2(.din(w_dff_B_oybLVK4D8_2),.dout(w_dff_B_izwdhGDY8_2),.clk(gclk));
	jdff dff_B_LFpGHjxF6_2(.din(w_dff_B_izwdhGDY8_2),.dout(w_dff_B_LFpGHjxF6_2),.clk(gclk));
	jdff dff_B_MxUou9Hc5_2(.din(w_dff_B_LFpGHjxF6_2),.dout(w_dff_B_MxUou9Hc5_2),.clk(gclk));
	jdff dff_B_xvJ6aTvz4_2(.din(w_dff_B_MxUou9Hc5_2),.dout(w_dff_B_xvJ6aTvz4_2),.clk(gclk));
	jdff dff_B_JRknODPh7_2(.din(w_dff_B_xvJ6aTvz4_2),.dout(w_dff_B_JRknODPh7_2),.clk(gclk));
	jdff dff_B_t7ZsAJgh2_2(.din(w_dff_B_JRknODPh7_2),.dout(w_dff_B_t7ZsAJgh2_2),.clk(gclk));
	jdff dff_B_Lo8FIWC53_2(.din(w_dff_B_t7ZsAJgh2_2),.dout(w_dff_B_Lo8FIWC53_2),.clk(gclk));
	jdff dff_B_k8XlVUA97_1(.din(n1308),.dout(w_dff_B_k8XlVUA97_1),.clk(gclk));
	jdff dff_B_fAgyJvSN6_2(.din(n1222),.dout(w_dff_B_fAgyJvSN6_2),.clk(gclk));
	jdff dff_B_mwyaLb3v2_2(.din(w_dff_B_fAgyJvSN6_2),.dout(w_dff_B_mwyaLb3v2_2),.clk(gclk));
	jdff dff_B_tJPE0WFp3_2(.din(w_dff_B_mwyaLb3v2_2),.dout(w_dff_B_tJPE0WFp3_2),.clk(gclk));
	jdff dff_B_68CUfuxP7_2(.din(w_dff_B_tJPE0WFp3_2),.dout(w_dff_B_68CUfuxP7_2),.clk(gclk));
	jdff dff_B_zlNpVvvW0_2(.din(w_dff_B_68CUfuxP7_2),.dout(w_dff_B_zlNpVvvW0_2),.clk(gclk));
	jdff dff_B_OPM4i01Q4_2(.din(w_dff_B_zlNpVvvW0_2),.dout(w_dff_B_OPM4i01Q4_2),.clk(gclk));
	jdff dff_B_fpKwXHvc4_2(.din(w_dff_B_OPM4i01Q4_2),.dout(w_dff_B_fpKwXHvc4_2),.clk(gclk));
	jdff dff_B_poSb7Tcn7_2(.din(w_dff_B_fpKwXHvc4_2),.dout(w_dff_B_poSb7Tcn7_2),.clk(gclk));
	jdff dff_B_aoMWe0xT4_2(.din(w_dff_B_poSb7Tcn7_2),.dout(w_dff_B_aoMWe0xT4_2),.clk(gclk));
	jdff dff_B_rDrlEccx5_2(.din(w_dff_B_aoMWe0xT4_2),.dout(w_dff_B_rDrlEccx5_2),.clk(gclk));
	jdff dff_B_3FbUVB1E7_2(.din(w_dff_B_rDrlEccx5_2),.dout(w_dff_B_3FbUVB1E7_2),.clk(gclk));
	jdff dff_B_nnpi5Kj04_2(.din(w_dff_B_3FbUVB1E7_2),.dout(w_dff_B_nnpi5Kj04_2),.clk(gclk));
	jdff dff_B_wray5jyJ6_2(.din(w_dff_B_nnpi5Kj04_2),.dout(w_dff_B_wray5jyJ6_2),.clk(gclk));
	jdff dff_B_yJ6ZsH4o8_2(.din(w_dff_B_wray5jyJ6_2),.dout(w_dff_B_yJ6ZsH4o8_2),.clk(gclk));
	jdff dff_B_jXAZaE1N3_2(.din(w_dff_B_yJ6ZsH4o8_2),.dout(w_dff_B_jXAZaE1N3_2),.clk(gclk));
	jdff dff_B_iYXLo5l90_2(.din(w_dff_B_jXAZaE1N3_2),.dout(w_dff_B_iYXLo5l90_2),.clk(gclk));
	jdff dff_B_5FOah2fI3_2(.din(w_dff_B_iYXLo5l90_2),.dout(w_dff_B_5FOah2fI3_2),.clk(gclk));
	jdff dff_B_mnKdMAz65_2(.din(w_dff_B_5FOah2fI3_2),.dout(w_dff_B_mnKdMAz65_2),.clk(gclk));
	jdff dff_B_vo7eoJt71_2(.din(w_dff_B_mnKdMAz65_2),.dout(w_dff_B_vo7eoJt71_2),.clk(gclk));
	jdff dff_B_nEYU0SN60_2(.din(w_dff_B_vo7eoJt71_2),.dout(w_dff_B_nEYU0SN60_2),.clk(gclk));
	jdff dff_B_uSNmt1l58_2(.din(w_dff_B_nEYU0SN60_2),.dout(w_dff_B_uSNmt1l58_2),.clk(gclk));
	jdff dff_B_d5vHjC0C0_2(.din(w_dff_B_uSNmt1l58_2),.dout(w_dff_B_d5vHjC0C0_2),.clk(gclk));
	jdff dff_B_y0Oo2BPK8_2(.din(w_dff_B_d5vHjC0C0_2),.dout(w_dff_B_y0Oo2BPK8_2),.clk(gclk));
	jdff dff_B_yNKXbDM99_2(.din(w_dff_B_y0Oo2BPK8_2),.dout(w_dff_B_yNKXbDM99_2),.clk(gclk));
	jdff dff_B_m6cRa4Jl3_2(.din(w_dff_B_yNKXbDM99_2),.dout(w_dff_B_m6cRa4Jl3_2),.clk(gclk));
	jdff dff_B_DwibTo361_2(.din(w_dff_B_m6cRa4Jl3_2),.dout(w_dff_B_DwibTo361_2),.clk(gclk));
	jdff dff_B_hg03bV8v8_2(.din(w_dff_B_DwibTo361_2),.dout(w_dff_B_hg03bV8v8_2),.clk(gclk));
	jdff dff_B_RnFolPgg2_2(.din(w_dff_B_hg03bV8v8_2),.dout(w_dff_B_RnFolPgg2_2),.clk(gclk));
	jdff dff_B_CdCj96At8_2(.din(w_dff_B_RnFolPgg2_2),.dout(w_dff_B_CdCj96At8_2),.clk(gclk));
	jdff dff_B_arwfT5Ft4_2(.din(w_dff_B_CdCj96At8_2),.dout(w_dff_B_arwfT5Ft4_2),.clk(gclk));
	jdff dff_B_tYntJP816_2(.din(w_dff_B_arwfT5Ft4_2),.dout(w_dff_B_tYntJP816_2),.clk(gclk));
	jdff dff_B_jg6mtGK87_2(.din(w_dff_B_tYntJP816_2),.dout(w_dff_B_jg6mtGK87_2),.clk(gclk));
	jdff dff_B_O9ILECp82_2(.din(w_dff_B_jg6mtGK87_2),.dout(w_dff_B_O9ILECp82_2),.clk(gclk));
	jdff dff_B_swlrL67e4_2(.din(w_dff_B_O9ILECp82_2),.dout(w_dff_B_swlrL67e4_2),.clk(gclk));
	jdff dff_B_A66EmYzY5_2(.din(w_dff_B_swlrL67e4_2),.dout(w_dff_B_A66EmYzY5_2),.clk(gclk));
	jdff dff_B_VhcX5Szs4_2(.din(w_dff_B_A66EmYzY5_2),.dout(w_dff_B_VhcX5Szs4_2),.clk(gclk));
	jdff dff_B_D7wBaV4Z1_2(.din(w_dff_B_VhcX5Szs4_2),.dout(w_dff_B_D7wBaV4Z1_2),.clk(gclk));
	jdff dff_B_N1AHSpAn2_2(.din(w_dff_B_D7wBaV4Z1_2),.dout(w_dff_B_N1AHSpAn2_2),.clk(gclk));
	jdff dff_B_39RFgBUm3_2(.din(w_dff_B_N1AHSpAn2_2),.dout(w_dff_B_39RFgBUm3_2),.clk(gclk));
	jdff dff_B_fiwM2wYC8_1(.din(n1223),.dout(w_dff_B_fiwM2wYC8_1),.clk(gclk));
	jdff dff_B_tKDdBQqd8_2(.din(n1131),.dout(w_dff_B_tKDdBQqd8_2),.clk(gclk));
	jdff dff_B_qNEzsbKg7_2(.din(w_dff_B_tKDdBQqd8_2),.dout(w_dff_B_qNEzsbKg7_2),.clk(gclk));
	jdff dff_B_vUOUi9cH3_2(.din(w_dff_B_qNEzsbKg7_2),.dout(w_dff_B_vUOUi9cH3_2),.clk(gclk));
	jdff dff_B_lP8AAloD7_2(.din(w_dff_B_vUOUi9cH3_2),.dout(w_dff_B_lP8AAloD7_2),.clk(gclk));
	jdff dff_B_W0DFx3Zh8_2(.din(w_dff_B_lP8AAloD7_2),.dout(w_dff_B_W0DFx3Zh8_2),.clk(gclk));
	jdff dff_B_ONs93hSM2_2(.din(w_dff_B_W0DFx3Zh8_2),.dout(w_dff_B_ONs93hSM2_2),.clk(gclk));
	jdff dff_B_ShxoNOvX9_2(.din(w_dff_B_ONs93hSM2_2),.dout(w_dff_B_ShxoNOvX9_2),.clk(gclk));
	jdff dff_B_01LndCTO5_2(.din(w_dff_B_ShxoNOvX9_2),.dout(w_dff_B_01LndCTO5_2),.clk(gclk));
	jdff dff_B_aUKBCvj80_2(.din(w_dff_B_01LndCTO5_2),.dout(w_dff_B_aUKBCvj80_2),.clk(gclk));
	jdff dff_B_eCkCW5nx3_2(.din(w_dff_B_aUKBCvj80_2),.dout(w_dff_B_eCkCW5nx3_2),.clk(gclk));
	jdff dff_B_lqT8ZVYz1_2(.din(w_dff_B_eCkCW5nx3_2),.dout(w_dff_B_lqT8ZVYz1_2),.clk(gclk));
	jdff dff_B_o8jYEeQb0_2(.din(w_dff_B_lqT8ZVYz1_2),.dout(w_dff_B_o8jYEeQb0_2),.clk(gclk));
	jdff dff_B_mnKFgr1B9_2(.din(w_dff_B_o8jYEeQb0_2),.dout(w_dff_B_mnKFgr1B9_2),.clk(gclk));
	jdff dff_B_p60nv3tk8_2(.din(w_dff_B_mnKFgr1B9_2),.dout(w_dff_B_p60nv3tk8_2),.clk(gclk));
	jdff dff_B_0BZbX3UZ5_2(.din(w_dff_B_p60nv3tk8_2),.dout(w_dff_B_0BZbX3UZ5_2),.clk(gclk));
	jdff dff_B_I14t2u4i9_2(.din(w_dff_B_0BZbX3UZ5_2),.dout(w_dff_B_I14t2u4i9_2),.clk(gclk));
	jdff dff_B_x4KC1XaE7_2(.din(w_dff_B_I14t2u4i9_2),.dout(w_dff_B_x4KC1XaE7_2),.clk(gclk));
	jdff dff_B_t5gKtYkM3_2(.din(w_dff_B_x4KC1XaE7_2),.dout(w_dff_B_t5gKtYkM3_2),.clk(gclk));
	jdff dff_B_7k9cYEWR5_2(.din(w_dff_B_t5gKtYkM3_2),.dout(w_dff_B_7k9cYEWR5_2),.clk(gclk));
	jdff dff_B_35gFl6HC6_2(.din(w_dff_B_7k9cYEWR5_2),.dout(w_dff_B_35gFl6HC6_2),.clk(gclk));
	jdff dff_B_DvyTw6HX9_2(.din(w_dff_B_35gFl6HC6_2),.dout(w_dff_B_DvyTw6HX9_2),.clk(gclk));
	jdff dff_B_aRmcyMxX6_2(.din(w_dff_B_DvyTw6HX9_2),.dout(w_dff_B_aRmcyMxX6_2),.clk(gclk));
	jdff dff_B_qVlpD0Ka4_2(.din(w_dff_B_aRmcyMxX6_2),.dout(w_dff_B_qVlpD0Ka4_2),.clk(gclk));
	jdff dff_B_OsW73hAU7_2(.din(w_dff_B_qVlpD0Ka4_2),.dout(w_dff_B_OsW73hAU7_2),.clk(gclk));
	jdff dff_B_gxQu3uKK3_2(.din(w_dff_B_OsW73hAU7_2),.dout(w_dff_B_gxQu3uKK3_2),.clk(gclk));
	jdff dff_B_Ckf0V3sk5_2(.din(w_dff_B_gxQu3uKK3_2),.dout(w_dff_B_Ckf0V3sk5_2),.clk(gclk));
	jdff dff_B_TFONE8Ha0_2(.din(w_dff_B_Ckf0V3sk5_2),.dout(w_dff_B_TFONE8Ha0_2),.clk(gclk));
	jdff dff_B_WDDXFCA29_2(.din(w_dff_B_TFONE8Ha0_2),.dout(w_dff_B_WDDXFCA29_2),.clk(gclk));
	jdff dff_B_kUMuguP50_2(.din(w_dff_B_WDDXFCA29_2),.dout(w_dff_B_kUMuguP50_2),.clk(gclk));
	jdff dff_B_NakSXBwn8_2(.din(w_dff_B_kUMuguP50_2),.dout(w_dff_B_NakSXBwn8_2),.clk(gclk));
	jdff dff_B_qRjbkKcV6_2(.din(w_dff_B_NakSXBwn8_2),.dout(w_dff_B_qRjbkKcV6_2),.clk(gclk));
	jdff dff_B_n9cBxznM3_2(.din(w_dff_B_qRjbkKcV6_2),.dout(w_dff_B_n9cBxznM3_2),.clk(gclk));
	jdff dff_B_ijHw9koU1_2(.din(w_dff_B_n9cBxznM3_2),.dout(w_dff_B_ijHw9koU1_2),.clk(gclk));
	jdff dff_B_TUI4EmhO3_2(.din(w_dff_B_ijHw9koU1_2),.dout(w_dff_B_TUI4EmhO3_2),.clk(gclk));
	jdff dff_B_1vHsV6SF0_2(.din(w_dff_B_TUI4EmhO3_2),.dout(w_dff_B_1vHsV6SF0_2),.clk(gclk));
	jdff dff_B_J3NOWJQd2_2(.din(w_dff_B_1vHsV6SF0_2),.dout(w_dff_B_J3NOWJQd2_2),.clk(gclk));
	jdff dff_B_HfWrQ1Ho7_1(.din(n1132),.dout(w_dff_B_HfWrQ1Ho7_1),.clk(gclk));
	jdff dff_B_KODIlDmX1_2(.din(n1033),.dout(w_dff_B_KODIlDmX1_2),.clk(gclk));
	jdff dff_B_csCOtoNU4_2(.din(w_dff_B_KODIlDmX1_2),.dout(w_dff_B_csCOtoNU4_2),.clk(gclk));
	jdff dff_B_9wGhnw8x6_2(.din(w_dff_B_csCOtoNU4_2),.dout(w_dff_B_9wGhnw8x6_2),.clk(gclk));
	jdff dff_B_CMWpwJBe2_2(.din(w_dff_B_9wGhnw8x6_2),.dout(w_dff_B_CMWpwJBe2_2),.clk(gclk));
	jdff dff_B_5y4qAQ0k8_2(.din(w_dff_B_CMWpwJBe2_2),.dout(w_dff_B_5y4qAQ0k8_2),.clk(gclk));
	jdff dff_B_O1yL9swT8_2(.din(w_dff_B_5y4qAQ0k8_2),.dout(w_dff_B_O1yL9swT8_2),.clk(gclk));
	jdff dff_B_K2dzaRKH4_2(.din(w_dff_B_O1yL9swT8_2),.dout(w_dff_B_K2dzaRKH4_2),.clk(gclk));
	jdff dff_B_92z9Qms06_2(.din(w_dff_B_K2dzaRKH4_2),.dout(w_dff_B_92z9Qms06_2),.clk(gclk));
	jdff dff_B_cWxRY6Ya0_2(.din(w_dff_B_92z9Qms06_2),.dout(w_dff_B_cWxRY6Ya0_2),.clk(gclk));
	jdff dff_B_pPMpScHQ3_2(.din(w_dff_B_cWxRY6Ya0_2),.dout(w_dff_B_pPMpScHQ3_2),.clk(gclk));
	jdff dff_B_TYUblta39_2(.din(w_dff_B_pPMpScHQ3_2),.dout(w_dff_B_TYUblta39_2),.clk(gclk));
	jdff dff_B_XIiO30kZ4_2(.din(w_dff_B_TYUblta39_2),.dout(w_dff_B_XIiO30kZ4_2),.clk(gclk));
	jdff dff_B_dfNUeEuS9_2(.din(w_dff_B_XIiO30kZ4_2),.dout(w_dff_B_dfNUeEuS9_2),.clk(gclk));
	jdff dff_B_7uOR295C2_2(.din(w_dff_B_dfNUeEuS9_2),.dout(w_dff_B_7uOR295C2_2),.clk(gclk));
	jdff dff_B_hXbwctaK6_2(.din(w_dff_B_7uOR295C2_2),.dout(w_dff_B_hXbwctaK6_2),.clk(gclk));
	jdff dff_B_gtQMHRbk1_2(.din(w_dff_B_hXbwctaK6_2),.dout(w_dff_B_gtQMHRbk1_2),.clk(gclk));
	jdff dff_B_uzVLRekc5_2(.din(w_dff_B_gtQMHRbk1_2),.dout(w_dff_B_uzVLRekc5_2),.clk(gclk));
	jdff dff_B_CARo65hi7_2(.din(w_dff_B_uzVLRekc5_2),.dout(w_dff_B_CARo65hi7_2),.clk(gclk));
	jdff dff_B_FDTDgNN44_2(.din(w_dff_B_CARo65hi7_2),.dout(w_dff_B_FDTDgNN44_2),.clk(gclk));
	jdff dff_B_YZ4VpJSX8_2(.din(w_dff_B_FDTDgNN44_2),.dout(w_dff_B_YZ4VpJSX8_2),.clk(gclk));
	jdff dff_B_OK4Ukae05_2(.din(w_dff_B_YZ4VpJSX8_2),.dout(w_dff_B_OK4Ukae05_2),.clk(gclk));
	jdff dff_B_AMWiKE6O4_2(.din(w_dff_B_OK4Ukae05_2),.dout(w_dff_B_AMWiKE6O4_2),.clk(gclk));
	jdff dff_B_TigrChrE8_2(.din(w_dff_B_AMWiKE6O4_2),.dout(w_dff_B_TigrChrE8_2),.clk(gclk));
	jdff dff_B_lJhJMmwD4_2(.din(w_dff_B_TigrChrE8_2),.dout(w_dff_B_lJhJMmwD4_2),.clk(gclk));
	jdff dff_B_TZa3XLot5_2(.din(w_dff_B_lJhJMmwD4_2),.dout(w_dff_B_TZa3XLot5_2),.clk(gclk));
	jdff dff_B_Ac4cxLrh2_2(.din(w_dff_B_TZa3XLot5_2),.dout(w_dff_B_Ac4cxLrh2_2),.clk(gclk));
	jdff dff_B_zROXxUve7_2(.din(w_dff_B_Ac4cxLrh2_2),.dout(w_dff_B_zROXxUve7_2),.clk(gclk));
	jdff dff_B_UsFytzGm9_2(.din(w_dff_B_zROXxUve7_2),.dout(w_dff_B_UsFytzGm9_2),.clk(gclk));
	jdff dff_B_S6HvVgXo8_2(.din(w_dff_B_UsFytzGm9_2),.dout(w_dff_B_S6HvVgXo8_2),.clk(gclk));
	jdff dff_B_DshDVSHv6_2(.din(w_dff_B_S6HvVgXo8_2),.dout(w_dff_B_DshDVSHv6_2),.clk(gclk));
	jdff dff_B_N5EhLutR4_2(.din(w_dff_B_DshDVSHv6_2),.dout(w_dff_B_N5EhLutR4_2),.clk(gclk));
	jdff dff_B_rxpvaiXx5_2(.din(w_dff_B_N5EhLutR4_2),.dout(w_dff_B_rxpvaiXx5_2),.clk(gclk));
	jdff dff_B_lQyCJl4Y6_2(.din(w_dff_B_rxpvaiXx5_2),.dout(w_dff_B_lQyCJl4Y6_2),.clk(gclk));
	jdff dff_B_RhSaeNsr6_1(.din(n1034),.dout(w_dff_B_RhSaeNsr6_1),.clk(gclk));
	jdff dff_B_W1mFT3IN0_2(.din(n934),.dout(w_dff_B_W1mFT3IN0_2),.clk(gclk));
	jdff dff_B_uTZGI3sU8_2(.din(w_dff_B_W1mFT3IN0_2),.dout(w_dff_B_uTZGI3sU8_2),.clk(gclk));
	jdff dff_B_6hRcDbyc0_2(.din(w_dff_B_uTZGI3sU8_2),.dout(w_dff_B_6hRcDbyc0_2),.clk(gclk));
	jdff dff_B_fAL3bVqH2_2(.din(w_dff_B_6hRcDbyc0_2),.dout(w_dff_B_fAL3bVqH2_2),.clk(gclk));
	jdff dff_B_reVJgRRt1_2(.din(w_dff_B_fAL3bVqH2_2),.dout(w_dff_B_reVJgRRt1_2),.clk(gclk));
	jdff dff_B_iwxoP96i4_2(.din(w_dff_B_reVJgRRt1_2),.dout(w_dff_B_iwxoP96i4_2),.clk(gclk));
	jdff dff_B_92Jd6xJe0_2(.din(w_dff_B_iwxoP96i4_2),.dout(w_dff_B_92Jd6xJe0_2),.clk(gclk));
	jdff dff_B_1lN2lGqZ9_2(.din(w_dff_B_92Jd6xJe0_2),.dout(w_dff_B_1lN2lGqZ9_2),.clk(gclk));
	jdff dff_B_bk9xbFrT0_2(.din(w_dff_B_1lN2lGqZ9_2),.dout(w_dff_B_bk9xbFrT0_2),.clk(gclk));
	jdff dff_B_omEZxyTQ5_2(.din(w_dff_B_bk9xbFrT0_2),.dout(w_dff_B_omEZxyTQ5_2),.clk(gclk));
	jdff dff_B_BPrLBHMV3_2(.din(w_dff_B_omEZxyTQ5_2),.dout(w_dff_B_BPrLBHMV3_2),.clk(gclk));
	jdff dff_B_ZUwYEeX83_2(.din(w_dff_B_BPrLBHMV3_2),.dout(w_dff_B_ZUwYEeX83_2),.clk(gclk));
	jdff dff_B_K4w2dVa61_2(.din(w_dff_B_ZUwYEeX83_2),.dout(w_dff_B_K4w2dVa61_2),.clk(gclk));
	jdff dff_B_tIM5N5Zq1_2(.din(w_dff_B_K4w2dVa61_2),.dout(w_dff_B_tIM5N5Zq1_2),.clk(gclk));
	jdff dff_B_hGxe35nt6_2(.din(w_dff_B_tIM5N5Zq1_2),.dout(w_dff_B_hGxe35nt6_2),.clk(gclk));
	jdff dff_B_TIjSAsJ70_2(.din(w_dff_B_hGxe35nt6_2),.dout(w_dff_B_TIjSAsJ70_2),.clk(gclk));
	jdff dff_B_nGrFAuFj2_2(.din(w_dff_B_TIjSAsJ70_2),.dout(w_dff_B_nGrFAuFj2_2),.clk(gclk));
	jdff dff_B_CwTMXs6S7_2(.din(w_dff_B_nGrFAuFj2_2),.dout(w_dff_B_CwTMXs6S7_2),.clk(gclk));
	jdff dff_B_nlxyfOhE6_2(.din(w_dff_B_CwTMXs6S7_2),.dout(w_dff_B_nlxyfOhE6_2),.clk(gclk));
	jdff dff_B_ponracsk3_2(.din(w_dff_B_nlxyfOhE6_2),.dout(w_dff_B_ponracsk3_2),.clk(gclk));
	jdff dff_B_A3eNbX6Y6_2(.din(w_dff_B_ponracsk3_2),.dout(w_dff_B_A3eNbX6Y6_2),.clk(gclk));
	jdff dff_B_8iMnrbZi7_2(.din(w_dff_B_A3eNbX6Y6_2),.dout(w_dff_B_8iMnrbZi7_2),.clk(gclk));
	jdff dff_B_G91A9Xx24_2(.din(w_dff_B_8iMnrbZi7_2),.dout(w_dff_B_G91A9Xx24_2),.clk(gclk));
	jdff dff_B_vlQPEQfi2_2(.din(w_dff_B_G91A9Xx24_2),.dout(w_dff_B_vlQPEQfi2_2),.clk(gclk));
	jdff dff_B_dQVHuCkX2_2(.din(w_dff_B_vlQPEQfi2_2),.dout(w_dff_B_dQVHuCkX2_2),.clk(gclk));
	jdff dff_B_WQd0TssQ8_2(.din(w_dff_B_dQVHuCkX2_2),.dout(w_dff_B_WQd0TssQ8_2),.clk(gclk));
	jdff dff_B_Di5fBYKC8_2(.din(w_dff_B_WQd0TssQ8_2),.dout(w_dff_B_Di5fBYKC8_2),.clk(gclk));
	jdff dff_B_TpaGXncm5_2(.din(w_dff_B_Di5fBYKC8_2),.dout(w_dff_B_TpaGXncm5_2),.clk(gclk));
	jdff dff_B_rRbimV570_2(.din(w_dff_B_TpaGXncm5_2),.dout(w_dff_B_rRbimV570_2),.clk(gclk));
	jdff dff_B_8BHbKbWp9_2(.din(w_dff_B_rRbimV570_2),.dout(w_dff_B_8BHbKbWp9_2),.clk(gclk));
	jdff dff_B_QJ7JBseb2_1(.din(n935),.dout(w_dff_B_QJ7JBseb2_1),.clk(gclk));
	jdff dff_B_OHTtpgJ00_2(.din(n832),.dout(w_dff_B_OHTtpgJ00_2),.clk(gclk));
	jdff dff_B_AnhGii639_2(.din(w_dff_B_OHTtpgJ00_2),.dout(w_dff_B_AnhGii639_2),.clk(gclk));
	jdff dff_B_rrnvr8jj2_2(.din(w_dff_B_AnhGii639_2),.dout(w_dff_B_rrnvr8jj2_2),.clk(gclk));
	jdff dff_B_NnPK0t1N6_2(.din(w_dff_B_rrnvr8jj2_2),.dout(w_dff_B_NnPK0t1N6_2),.clk(gclk));
	jdff dff_B_hNpaOvIQ3_2(.din(w_dff_B_NnPK0t1N6_2),.dout(w_dff_B_hNpaOvIQ3_2),.clk(gclk));
	jdff dff_B_FTw4nQhW1_2(.din(w_dff_B_hNpaOvIQ3_2),.dout(w_dff_B_FTw4nQhW1_2),.clk(gclk));
	jdff dff_B_cXiKRgxT2_2(.din(w_dff_B_FTw4nQhW1_2),.dout(w_dff_B_cXiKRgxT2_2),.clk(gclk));
	jdff dff_B_VbYUTTOn2_2(.din(w_dff_B_cXiKRgxT2_2),.dout(w_dff_B_VbYUTTOn2_2),.clk(gclk));
	jdff dff_B_IKda24pJ4_2(.din(w_dff_B_VbYUTTOn2_2),.dout(w_dff_B_IKda24pJ4_2),.clk(gclk));
	jdff dff_B_QpfYUdSV3_2(.din(w_dff_B_IKda24pJ4_2),.dout(w_dff_B_QpfYUdSV3_2),.clk(gclk));
	jdff dff_B_4GN8XVSh0_2(.din(w_dff_B_QpfYUdSV3_2),.dout(w_dff_B_4GN8XVSh0_2),.clk(gclk));
	jdff dff_B_BPYizo1R5_2(.din(w_dff_B_4GN8XVSh0_2),.dout(w_dff_B_BPYizo1R5_2),.clk(gclk));
	jdff dff_B_Zi2Esws10_2(.din(w_dff_B_BPYizo1R5_2),.dout(w_dff_B_Zi2Esws10_2),.clk(gclk));
	jdff dff_B_DzL6x2KE2_2(.din(w_dff_B_Zi2Esws10_2),.dout(w_dff_B_DzL6x2KE2_2),.clk(gclk));
	jdff dff_B_W828Mu7m0_2(.din(w_dff_B_DzL6x2KE2_2),.dout(w_dff_B_W828Mu7m0_2),.clk(gclk));
	jdff dff_B_faAN3UCE9_2(.din(w_dff_B_W828Mu7m0_2),.dout(w_dff_B_faAN3UCE9_2),.clk(gclk));
	jdff dff_B_Y2TeiGFM2_2(.din(w_dff_B_faAN3UCE9_2),.dout(w_dff_B_Y2TeiGFM2_2),.clk(gclk));
	jdff dff_B_D1Mgrz1W5_2(.din(w_dff_B_Y2TeiGFM2_2),.dout(w_dff_B_D1Mgrz1W5_2),.clk(gclk));
	jdff dff_B_cWLBa6684_2(.din(w_dff_B_D1Mgrz1W5_2),.dout(w_dff_B_cWLBa6684_2),.clk(gclk));
	jdff dff_B_LA41AzYl7_2(.din(w_dff_B_cWLBa6684_2),.dout(w_dff_B_LA41AzYl7_2),.clk(gclk));
	jdff dff_B_hnH68s2H6_2(.din(w_dff_B_LA41AzYl7_2),.dout(w_dff_B_hnH68s2H6_2),.clk(gclk));
	jdff dff_B_kAYKam8T5_2(.din(w_dff_B_hnH68s2H6_2),.dout(w_dff_B_kAYKam8T5_2),.clk(gclk));
	jdff dff_B_ZxOyhqWS8_2(.din(w_dff_B_kAYKam8T5_2),.dout(w_dff_B_ZxOyhqWS8_2),.clk(gclk));
	jdff dff_B_XcjG0ExS7_2(.din(w_dff_B_ZxOyhqWS8_2),.dout(w_dff_B_XcjG0ExS7_2),.clk(gclk));
	jdff dff_B_1kkDEOlE6_2(.din(w_dff_B_XcjG0ExS7_2),.dout(w_dff_B_1kkDEOlE6_2),.clk(gclk));
	jdff dff_B_Hiw2Z4ik1_2(.din(w_dff_B_1kkDEOlE6_2),.dout(w_dff_B_Hiw2Z4ik1_2),.clk(gclk));
	jdff dff_B_0jYhmeDR2_2(.din(w_dff_B_Hiw2Z4ik1_2),.dout(w_dff_B_0jYhmeDR2_2),.clk(gclk));
	jdff dff_B_aKoY2FFS5_1(.din(n833),.dout(w_dff_B_aKoY2FFS5_1),.clk(gclk));
	jdff dff_B_7MdYhEU40_2(.din(n734),.dout(w_dff_B_7MdYhEU40_2),.clk(gclk));
	jdff dff_B_bYsAvfoF0_2(.din(w_dff_B_7MdYhEU40_2),.dout(w_dff_B_bYsAvfoF0_2),.clk(gclk));
	jdff dff_B_8SEpU9cv1_2(.din(w_dff_B_bYsAvfoF0_2),.dout(w_dff_B_8SEpU9cv1_2),.clk(gclk));
	jdff dff_B_IxA3BBVu1_2(.din(w_dff_B_8SEpU9cv1_2),.dout(w_dff_B_IxA3BBVu1_2),.clk(gclk));
	jdff dff_B_4VHLFzQw3_2(.din(w_dff_B_IxA3BBVu1_2),.dout(w_dff_B_4VHLFzQw3_2),.clk(gclk));
	jdff dff_B_jBQ4GdPP9_2(.din(w_dff_B_4VHLFzQw3_2),.dout(w_dff_B_jBQ4GdPP9_2),.clk(gclk));
	jdff dff_B_LPjKVJF13_2(.din(w_dff_B_jBQ4GdPP9_2),.dout(w_dff_B_LPjKVJF13_2),.clk(gclk));
	jdff dff_B_MOmlbwMm4_2(.din(w_dff_B_LPjKVJF13_2),.dout(w_dff_B_MOmlbwMm4_2),.clk(gclk));
	jdff dff_B_cr8VTA2l6_2(.din(w_dff_B_MOmlbwMm4_2),.dout(w_dff_B_cr8VTA2l6_2),.clk(gclk));
	jdff dff_B_qlilAu5e1_2(.din(w_dff_B_cr8VTA2l6_2),.dout(w_dff_B_qlilAu5e1_2),.clk(gclk));
	jdff dff_B_nqOWRDfA9_2(.din(w_dff_B_qlilAu5e1_2),.dout(w_dff_B_nqOWRDfA9_2),.clk(gclk));
	jdff dff_B_c95FA0pp0_2(.din(w_dff_B_nqOWRDfA9_2),.dout(w_dff_B_c95FA0pp0_2),.clk(gclk));
	jdff dff_B_7wpSharB5_2(.din(w_dff_B_c95FA0pp0_2),.dout(w_dff_B_7wpSharB5_2),.clk(gclk));
	jdff dff_B_iAoUph6s3_2(.din(w_dff_B_7wpSharB5_2),.dout(w_dff_B_iAoUph6s3_2),.clk(gclk));
	jdff dff_B_10zKxQgf3_2(.din(w_dff_B_iAoUph6s3_2),.dout(w_dff_B_10zKxQgf3_2),.clk(gclk));
	jdff dff_B_ebOEtC5u9_2(.din(w_dff_B_10zKxQgf3_2),.dout(w_dff_B_ebOEtC5u9_2),.clk(gclk));
	jdff dff_B_33YMv3sj6_2(.din(w_dff_B_ebOEtC5u9_2),.dout(w_dff_B_33YMv3sj6_2),.clk(gclk));
	jdff dff_B_oOUXpSxl3_2(.din(w_dff_B_33YMv3sj6_2),.dout(w_dff_B_oOUXpSxl3_2),.clk(gclk));
	jdff dff_B_nwcT9UN73_2(.din(w_dff_B_oOUXpSxl3_2),.dout(w_dff_B_nwcT9UN73_2),.clk(gclk));
	jdff dff_B_3u7FlmR44_2(.din(w_dff_B_nwcT9UN73_2),.dout(w_dff_B_3u7FlmR44_2),.clk(gclk));
	jdff dff_B_Db3Odp5g5_2(.din(w_dff_B_3u7FlmR44_2),.dout(w_dff_B_Db3Odp5g5_2),.clk(gclk));
	jdff dff_B_QywCoaMc4_2(.din(w_dff_B_Db3Odp5g5_2),.dout(w_dff_B_QywCoaMc4_2),.clk(gclk));
	jdff dff_B_aWxI0aVn1_2(.din(w_dff_B_QywCoaMc4_2),.dout(w_dff_B_aWxI0aVn1_2),.clk(gclk));
	jdff dff_B_oRp3NQyX5_2(.din(w_dff_B_aWxI0aVn1_2),.dout(w_dff_B_oRp3NQyX5_2),.clk(gclk));
	jdff dff_B_dKuj7UIM9_1(.din(n735),.dout(w_dff_B_dKuj7UIM9_1),.clk(gclk));
	jdff dff_B_q3QMKSYf2_2(.din(n642),.dout(w_dff_B_q3QMKSYf2_2),.clk(gclk));
	jdff dff_B_Aph4nQxB0_2(.din(w_dff_B_q3QMKSYf2_2),.dout(w_dff_B_Aph4nQxB0_2),.clk(gclk));
	jdff dff_B_cgHpw67p6_2(.din(w_dff_B_Aph4nQxB0_2),.dout(w_dff_B_cgHpw67p6_2),.clk(gclk));
	jdff dff_B_sl3PHFQe5_2(.din(w_dff_B_cgHpw67p6_2),.dout(w_dff_B_sl3PHFQe5_2),.clk(gclk));
	jdff dff_B_75yho7qO7_2(.din(w_dff_B_sl3PHFQe5_2),.dout(w_dff_B_75yho7qO7_2),.clk(gclk));
	jdff dff_B_oOhw1uEk5_2(.din(w_dff_B_75yho7qO7_2),.dout(w_dff_B_oOhw1uEk5_2),.clk(gclk));
	jdff dff_B_8eyCW8ID0_2(.din(w_dff_B_oOhw1uEk5_2),.dout(w_dff_B_8eyCW8ID0_2),.clk(gclk));
	jdff dff_B_0z2WCI0I5_2(.din(w_dff_B_8eyCW8ID0_2),.dout(w_dff_B_0z2WCI0I5_2),.clk(gclk));
	jdff dff_B_0iTd3ZHM4_2(.din(w_dff_B_0z2WCI0I5_2),.dout(w_dff_B_0iTd3ZHM4_2),.clk(gclk));
	jdff dff_B_ckLG8WYz6_2(.din(w_dff_B_0iTd3ZHM4_2),.dout(w_dff_B_ckLG8WYz6_2),.clk(gclk));
	jdff dff_B_FlSiSvfJ8_2(.din(w_dff_B_ckLG8WYz6_2),.dout(w_dff_B_FlSiSvfJ8_2),.clk(gclk));
	jdff dff_B_KSHntsTn6_2(.din(w_dff_B_FlSiSvfJ8_2),.dout(w_dff_B_KSHntsTn6_2),.clk(gclk));
	jdff dff_B_XbMv8Vz49_2(.din(w_dff_B_KSHntsTn6_2),.dout(w_dff_B_XbMv8Vz49_2),.clk(gclk));
	jdff dff_B_4CPKUTPl6_2(.din(w_dff_B_XbMv8Vz49_2),.dout(w_dff_B_4CPKUTPl6_2),.clk(gclk));
	jdff dff_B_RXc1X9gg8_2(.din(w_dff_B_4CPKUTPl6_2),.dout(w_dff_B_RXc1X9gg8_2),.clk(gclk));
	jdff dff_B_SrOlL3PA3_2(.din(w_dff_B_RXc1X9gg8_2),.dout(w_dff_B_SrOlL3PA3_2),.clk(gclk));
	jdff dff_B_boADKgOE7_2(.din(w_dff_B_SrOlL3PA3_2),.dout(w_dff_B_boADKgOE7_2),.clk(gclk));
	jdff dff_B_hG7l2ONS5_2(.din(w_dff_B_boADKgOE7_2),.dout(w_dff_B_hG7l2ONS5_2),.clk(gclk));
	jdff dff_B_V92Sy3Sx9_2(.din(w_dff_B_hG7l2ONS5_2),.dout(w_dff_B_V92Sy3Sx9_2),.clk(gclk));
	jdff dff_B_TuM6Ewv20_2(.din(w_dff_B_V92Sy3Sx9_2),.dout(w_dff_B_TuM6Ewv20_2),.clk(gclk));
	jdff dff_B_5qY27qCF0_2(.din(w_dff_B_TuM6Ewv20_2),.dout(w_dff_B_5qY27qCF0_2),.clk(gclk));
	jdff dff_B_aQcRGXAd3_1(.din(n643),.dout(w_dff_B_aQcRGXAd3_1),.clk(gclk));
	jdff dff_B_zf7qMEU36_2(.din(n557),.dout(w_dff_B_zf7qMEU36_2),.clk(gclk));
	jdff dff_B_H0CaMaGA1_2(.din(w_dff_B_zf7qMEU36_2),.dout(w_dff_B_H0CaMaGA1_2),.clk(gclk));
	jdff dff_B_oot3Kj9n4_2(.din(w_dff_B_H0CaMaGA1_2),.dout(w_dff_B_oot3Kj9n4_2),.clk(gclk));
	jdff dff_B_r4T12Dzd2_2(.din(w_dff_B_oot3Kj9n4_2),.dout(w_dff_B_r4T12Dzd2_2),.clk(gclk));
	jdff dff_B_0ge5Pz5b8_2(.din(w_dff_B_r4T12Dzd2_2),.dout(w_dff_B_0ge5Pz5b8_2),.clk(gclk));
	jdff dff_B_G5cskc422_2(.din(w_dff_B_0ge5Pz5b8_2),.dout(w_dff_B_G5cskc422_2),.clk(gclk));
	jdff dff_B_JxoS9pvz3_2(.din(w_dff_B_G5cskc422_2),.dout(w_dff_B_JxoS9pvz3_2),.clk(gclk));
	jdff dff_B_heZSkhma0_2(.din(w_dff_B_JxoS9pvz3_2),.dout(w_dff_B_heZSkhma0_2),.clk(gclk));
	jdff dff_B_wfBTfFld2_2(.din(w_dff_B_heZSkhma0_2),.dout(w_dff_B_wfBTfFld2_2),.clk(gclk));
	jdff dff_B_FXD2ZjPd2_2(.din(w_dff_B_wfBTfFld2_2),.dout(w_dff_B_FXD2ZjPd2_2),.clk(gclk));
	jdff dff_B_XJ9TIffT4_2(.din(w_dff_B_FXD2ZjPd2_2),.dout(w_dff_B_XJ9TIffT4_2),.clk(gclk));
	jdff dff_B_mQTIjlwR0_2(.din(w_dff_B_XJ9TIffT4_2),.dout(w_dff_B_mQTIjlwR0_2),.clk(gclk));
	jdff dff_B_E0WKH84L1_2(.din(w_dff_B_mQTIjlwR0_2),.dout(w_dff_B_E0WKH84L1_2),.clk(gclk));
	jdff dff_B_C7I1qSDs0_2(.din(w_dff_B_E0WKH84L1_2),.dout(w_dff_B_C7I1qSDs0_2),.clk(gclk));
	jdff dff_B_fssYfKpV7_2(.din(w_dff_B_C7I1qSDs0_2),.dout(w_dff_B_fssYfKpV7_2),.clk(gclk));
	jdff dff_B_Sdh0qhQX6_2(.din(w_dff_B_fssYfKpV7_2),.dout(w_dff_B_Sdh0qhQX6_2),.clk(gclk));
	jdff dff_B_fPtc7Jlv2_2(.din(w_dff_B_Sdh0qhQX6_2),.dout(w_dff_B_fPtc7Jlv2_2),.clk(gclk));
	jdff dff_B_5g0nQWiE2_2(.din(w_dff_B_fPtc7Jlv2_2),.dout(w_dff_B_5g0nQWiE2_2),.clk(gclk));
	jdff dff_B_P1aw5ykX6_1(.din(n558),.dout(w_dff_B_P1aw5ykX6_1),.clk(gclk));
	jdff dff_B_NXFFFSE95_2(.din(n479),.dout(w_dff_B_NXFFFSE95_2),.clk(gclk));
	jdff dff_B_qUFF4Dlu1_2(.din(w_dff_B_NXFFFSE95_2),.dout(w_dff_B_qUFF4Dlu1_2),.clk(gclk));
	jdff dff_B_PmlSuEvl6_2(.din(w_dff_B_qUFF4Dlu1_2),.dout(w_dff_B_PmlSuEvl6_2),.clk(gclk));
	jdff dff_B_9BnGul3M6_2(.din(w_dff_B_PmlSuEvl6_2),.dout(w_dff_B_9BnGul3M6_2),.clk(gclk));
	jdff dff_B_sIjyY2IA6_2(.din(w_dff_B_9BnGul3M6_2),.dout(w_dff_B_sIjyY2IA6_2),.clk(gclk));
	jdff dff_B_wNgmwsv64_2(.din(w_dff_B_sIjyY2IA6_2),.dout(w_dff_B_wNgmwsv64_2),.clk(gclk));
	jdff dff_B_8kIr1eeO8_2(.din(w_dff_B_wNgmwsv64_2),.dout(w_dff_B_8kIr1eeO8_2),.clk(gclk));
	jdff dff_B_JY2n58mY7_2(.din(w_dff_B_8kIr1eeO8_2),.dout(w_dff_B_JY2n58mY7_2),.clk(gclk));
	jdff dff_B_x1U1S38Z9_2(.din(w_dff_B_JY2n58mY7_2),.dout(w_dff_B_x1U1S38Z9_2),.clk(gclk));
	jdff dff_B_ZXqKzxfj4_2(.din(w_dff_B_x1U1S38Z9_2),.dout(w_dff_B_ZXqKzxfj4_2),.clk(gclk));
	jdff dff_B_hpZCRbIk6_2(.din(w_dff_B_ZXqKzxfj4_2),.dout(w_dff_B_hpZCRbIk6_2),.clk(gclk));
	jdff dff_B_3GJtlzYM1_2(.din(w_dff_B_hpZCRbIk6_2),.dout(w_dff_B_3GJtlzYM1_2),.clk(gclk));
	jdff dff_B_zgg8Tj2w8_2(.din(w_dff_B_3GJtlzYM1_2),.dout(w_dff_B_zgg8Tj2w8_2),.clk(gclk));
	jdff dff_B_4w8tkCCg1_2(.din(w_dff_B_zgg8Tj2w8_2),.dout(w_dff_B_4w8tkCCg1_2),.clk(gclk));
	jdff dff_B_L4ZbzIDi7_2(.din(w_dff_B_4w8tkCCg1_2),.dout(w_dff_B_L4ZbzIDi7_2),.clk(gclk));
	jdff dff_B_6HH7rVy35_1(.din(n480),.dout(w_dff_B_6HH7rVy35_1),.clk(gclk));
	jdff dff_B_gVsqYsu18_2(.din(n408),.dout(w_dff_B_gVsqYsu18_2),.clk(gclk));
	jdff dff_B_ytMNg9Lb1_2(.din(w_dff_B_gVsqYsu18_2),.dout(w_dff_B_ytMNg9Lb1_2),.clk(gclk));
	jdff dff_B_6WZRlhWR4_2(.din(w_dff_B_ytMNg9Lb1_2),.dout(w_dff_B_6WZRlhWR4_2),.clk(gclk));
	jdff dff_B_h0LQLSH50_2(.din(w_dff_B_6WZRlhWR4_2),.dout(w_dff_B_h0LQLSH50_2),.clk(gclk));
	jdff dff_B_I3EjWxr31_2(.din(w_dff_B_h0LQLSH50_2),.dout(w_dff_B_I3EjWxr31_2),.clk(gclk));
	jdff dff_B_SlXB7Bt70_2(.din(w_dff_B_I3EjWxr31_2),.dout(w_dff_B_SlXB7Bt70_2),.clk(gclk));
	jdff dff_B_HPsLlWeB0_2(.din(w_dff_B_SlXB7Bt70_2),.dout(w_dff_B_HPsLlWeB0_2),.clk(gclk));
	jdff dff_B_ulNJqK5x1_2(.din(w_dff_B_HPsLlWeB0_2),.dout(w_dff_B_ulNJqK5x1_2),.clk(gclk));
	jdff dff_B_vy5M9ujs3_2(.din(w_dff_B_ulNJqK5x1_2),.dout(w_dff_B_vy5M9ujs3_2),.clk(gclk));
	jdff dff_B_3FelmzPf6_2(.din(w_dff_B_vy5M9ujs3_2),.dout(w_dff_B_3FelmzPf6_2),.clk(gclk));
	jdff dff_B_I2vQsKeF9_2(.din(w_dff_B_3FelmzPf6_2),.dout(w_dff_B_I2vQsKeF9_2),.clk(gclk));
	jdff dff_B_hhHb4CZS5_2(.din(w_dff_B_I2vQsKeF9_2),.dout(w_dff_B_hhHb4CZS5_2),.clk(gclk));
	jdff dff_B_YL95S5n31_1(.din(n409),.dout(w_dff_B_YL95S5n31_1),.clk(gclk));
	jdff dff_B_87uMtoxF9_2(.din(n345),.dout(w_dff_B_87uMtoxF9_2),.clk(gclk));
	jdff dff_B_HJqRWbSf9_2(.din(w_dff_B_87uMtoxF9_2),.dout(w_dff_B_HJqRWbSf9_2),.clk(gclk));
	jdff dff_B_8yUtVIQm2_2(.din(w_dff_B_HJqRWbSf9_2),.dout(w_dff_B_8yUtVIQm2_2),.clk(gclk));
	jdff dff_B_L2En0x2s0_2(.din(w_dff_B_8yUtVIQm2_2),.dout(w_dff_B_L2En0x2s0_2),.clk(gclk));
	jdff dff_B_G4hiu4kD4_2(.din(w_dff_B_L2En0x2s0_2),.dout(w_dff_B_G4hiu4kD4_2),.clk(gclk));
	jdff dff_B_sceqQ9rB1_2(.din(w_dff_B_G4hiu4kD4_2),.dout(w_dff_B_sceqQ9rB1_2),.clk(gclk));
	jdff dff_B_Qh4mReII3_2(.din(w_dff_B_sceqQ9rB1_2),.dout(w_dff_B_Qh4mReII3_2),.clk(gclk));
	jdff dff_B_IZ53g2WM5_2(.din(w_dff_B_Qh4mReII3_2),.dout(w_dff_B_IZ53g2WM5_2),.clk(gclk));
	jdff dff_B_9RkqwVp20_2(.din(w_dff_B_IZ53g2WM5_2),.dout(w_dff_B_9RkqwVp20_2),.clk(gclk));
	jdff dff_B_D35Bkf912_2(.din(n366),.dout(w_dff_B_D35Bkf912_2),.clk(gclk));
	jdff dff_B_ir1ZwmwY5_1(.din(n346),.dout(w_dff_B_ir1ZwmwY5_1),.clk(gclk));
	jdff dff_B_EfvDEuPI7_2(.din(n289),.dout(w_dff_B_EfvDEuPI7_2),.clk(gclk));
	jdff dff_B_SFqcnKhA5_2(.din(w_dff_B_EfvDEuPI7_2),.dout(w_dff_B_SFqcnKhA5_2),.clk(gclk));
	jdff dff_B_OVN1Mg9T4_2(.din(w_dff_B_SFqcnKhA5_2),.dout(w_dff_B_OVN1Mg9T4_2),.clk(gclk));
	jdff dff_B_6kAhJTRB4_2(.din(w_dff_B_OVN1Mg9T4_2),.dout(w_dff_B_6kAhJTRB4_2),.clk(gclk));
	jdff dff_B_MKnRdFyu1_2(.din(w_dff_B_6kAhJTRB4_2),.dout(w_dff_B_MKnRdFyu1_2),.clk(gclk));
	jdff dff_B_EZJuavUv4_2(.din(w_dff_B_MKnRdFyu1_2),.dout(w_dff_B_EZJuavUv4_2),.clk(gclk));
	jdff dff_B_KrkZHRZ11_2(.din(n303),.dout(w_dff_B_KrkZHRZ11_2),.clk(gclk));
	jdff dff_B_HOBApmeT6_2(.din(n241),.dout(w_dff_B_HOBApmeT6_2),.clk(gclk));
	jdff dff_B_yNro1q3L6_2(.din(w_dff_B_HOBApmeT6_2),.dout(w_dff_B_yNro1q3L6_2),.clk(gclk));
	jdff dff_B_DPQAd0JT2_2(.din(w_dff_B_yNro1q3L6_2),.dout(w_dff_B_DPQAd0JT2_2),.clk(gclk));
	jdff dff_B_dFtM3qTM2_0(.din(n246),.dout(w_dff_B_dFtM3qTM2_0),.clk(gclk));
	jdff dff_A_ltPdOqju8_0(.dout(w_n196_0[0]),.din(w_dff_A_ltPdOqju8_0),.clk(gclk));
	jdff dff_A_JUhNNVgm0_0(.dout(w_dff_A_ltPdOqju8_0),.din(w_dff_A_JUhNNVgm0_0),.clk(gclk));
	jdff dff_A_Kt85JJ044_1(.dout(w_n196_0[1]),.din(w_dff_A_Kt85JJ044_1),.clk(gclk));
	jdff dff_A_ZLkAxtuN9_1(.dout(w_dff_A_Kt85JJ044_1),.din(w_dff_A_ZLkAxtuN9_1),.clk(gclk));
	jdff dff_B_8w74N4ai7_2(.din(n1465),.dout(w_dff_B_8w74N4ai7_2),.clk(gclk));
	jdff dff_B_tyeEbBLJ7_1(.din(n1463),.dout(w_dff_B_tyeEbBLJ7_1),.clk(gclk));
	jdff dff_B_fVuhJmVK5_2(.din(n1390),.dout(w_dff_B_fVuhJmVK5_2),.clk(gclk));
	jdff dff_B_ZJenFmRo7_2(.din(w_dff_B_fVuhJmVK5_2),.dout(w_dff_B_ZJenFmRo7_2),.clk(gclk));
	jdff dff_B_HPTKlO0P7_2(.din(w_dff_B_ZJenFmRo7_2),.dout(w_dff_B_HPTKlO0P7_2),.clk(gclk));
	jdff dff_B_QutrbreA6_2(.din(w_dff_B_HPTKlO0P7_2),.dout(w_dff_B_QutrbreA6_2),.clk(gclk));
	jdff dff_B_nk9i37RL3_2(.din(w_dff_B_QutrbreA6_2),.dout(w_dff_B_nk9i37RL3_2),.clk(gclk));
	jdff dff_B_Y8DcatZY5_2(.din(w_dff_B_nk9i37RL3_2),.dout(w_dff_B_Y8DcatZY5_2),.clk(gclk));
	jdff dff_B_daMRik372_2(.din(w_dff_B_Y8DcatZY5_2),.dout(w_dff_B_daMRik372_2),.clk(gclk));
	jdff dff_B_TuZLNalW6_2(.din(w_dff_B_daMRik372_2),.dout(w_dff_B_TuZLNalW6_2),.clk(gclk));
	jdff dff_B_cJyEoYtY8_2(.din(w_dff_B_TuZLNalW6_2),.dout(w_dff_B_cJyEoYtY8_2),.clk(gclk));
	jdff dff_B_uPwcfmdA8_2(.din(w_dff_B_cJyEoYtY8_2),.dout(w_dff_B_uPwcfmdA8_2),.clk(gclk));
	jdff dff_B_FdUkVYnb0_2(.din(w_dff_B_uPwcfmdA8_2),.dout(w_dff_B_FdUkVYnb0_2),.clk(gclk));
	jdff dff_B_M7U83DY40_2(.din(w_dff_B_FdUkVYnb0_2),.dout(w_dff_B_M7U83DY40_2),.clk(gclk));
	jdff dff_B_qhWFS2cL0_2(.din(w_dff_B_M7U83DY40_2),.dout(w_dff_B_qhWFS2cL0_2),.clk(gclk));
	jdff dff_B_jcnHWUJX7_2(.din(w_dff_B_qhWFS2cL0_2),.dout(w_dff_B_jcnHWUJX7_2),.clk(gclk));
	jdff dff_B_v5yd2RQ81_2(.din(w_dff_B_jcnHWUJX7_2),.dout(w_dff_B_v5yd2RQ81_2),.clk(gclk));
	jdff dff_B_IICoYyHR3_2(.din(w_dff_B_v5yd2RQ81_2),.dout(w_dff_B_IICoYyHR3_2),.clk(gclk));
	jdff dff_B_pmRUkfVb4_2(.din(w_dff_B_IICoYyHR3_2),.dout(w_dff_B_pmRUkfVb4_2),.clk(gclk));
	jdff dff_B_mh4S1d5X4_2(.din(w_dff_B_pmRUkfVb4_2),.dout(w_dff_B_mh4S1d5X4_2),.clk(gclk));
	jdff dff_B_S5gXFcqx8_2(.din(w_dff_B_mh4S1d5X4_2),.dout(w_dff_B_S5gXFcqx8_2),.clk(gclk));
	jdff dff_B_UdVJUrad3_2(.din(w_dff_B_S5gXFcqx8_2),.dout(w_dff_B_UdVJUrad3_2),.clk(gclk));
	jdff dff_B_CuWwkZcY5_2(.din(w_dff_B_UdVJUrad3_2),.dout(w_dff_B_CuWwkZcY5_2),.clk(gclk));
	jdff dff_B_w0cZCKHO9_2(.din(w_dff_B_CuWwkZcY5_2),.dout(w_dff_B_w0cZCKHO9_2),.clk(gclk));
	jdff dff_B_6Z3bVJ5f8_2(.din(w_dff_B_w0cZCKHO9_2),.dout(w_dff_B_6Z3bVJ5f8_2),.clk(gclk));
	jdff dff_B_yzFAqiAR7_2(.din(w_dff_B_6Z3bVJ5f8_2),.dout(w_dff_B_yzFAqiAR7_2),.clk(gclk));
	jdff dff_B_7iYX3Mei0_2(.din(w_dff_B_yzFAqiAR7_2),.dout(w_dff_B_7iYX3Mei0_2),.clk(gclk));
	jdff dff_B_6pPTLiTa6_2(.din(w_dff_B_7iYX3Mei0_2),.dout(w_dff_B_6pPTLiTa6_2),.clk(gclk));
	jdff dff_B_IoZO6PAx8_2(.din(w_dff_B_6pPTLiTa6_2),.dout(w_dff_B_IoZO6PAx8_2),.clk(gclk));
	jdff dff_B_yAXuRTv26_2(.din(w_dff_B_IoZO6PAx8_2),.dout(w_dff_B_yAXuRTv26_2),.clk(gclk));
	jdff dff_B_VNPO8uiN9_2(.din(w_dff_B_yAXuRTv26_2),.dout(w_dff_B_VNPO8uiN9_2),.clk(gclk));
	jdff dff_B_B79uhzjP3_2(.din(w_dff_B_VNPO8uiN9_2),.dout(w_dff_B_B79uhzjP3_2),.clk(gclk));
	jdff dff_B_BlxmijrU6_2(.din(w_dff_B_B79uhzjP3_2),.dout(w_dff_B_BlxmijrU6_2),.clk(gclk));
	jdff dff_B_58QYTuvJ5_2(.din(w_dff_B_BlxmijrU6_2),.dout(w_dff_B_58QYTuvJ5_2),.clk(gclk));
	jdff dff_B_QTjHgQ1H1_2(.din(w_dff_B_58QYTuvJ5_2),.dout(w_dff_B_QTjHgQ1H1_2),.clk(gclk));
	jdff dff_B_pbLRlp6D9_2(.din(w_dff_B_QTjHgQ1H1_2),.dout(w_dff_B_pbLRlp6D9_2),.clk(gclk));
	jdff dff_B_fGObqosS0_2(.din(w_dff_B_pbLRlp6D9_2),.dout(w_dff_B_fGObqosS0_2),.clk(gclk));
	jdff dff_B_ebXtDkaj5_2(.din(w_dff_B_fGObqosS0_2),.dout(w_dff_B_ebXtDkaj5_2),.clk(gclk));
	jdff dff_B_2y2RXh0P5_2(.din(w_dff_B_ebXtDkaj5_2),.dout(w_dff_B_2y2RXh0P5_2),.clk(gclk));
	jdff dff_B_frlZztg88_2(.din(w_dff_B_2y2RXh0P5_2),.dout(w_dff_B_frlZztg88_2),.clk(gclk));
	jdff dff_B_AzscMRNQ4_2(.din(w_dff_B_frlZztg88_2),.dout(w_dff_B_AzscMRNQ4_2),.clk(gclk));
	jdff dff_B_bWQfYQug0_2(.din(w_dff_B_AzscMRNQ4_2),.dout(w_dff_B_bWQfYQug0_2),.clk(gclk));
	jdff dff_B_IMR3K2bM4_2(.din(w_dff_B_bWQfYQug0_2),.dout(w_dff_B_IMR3K2bM4_2),.clk(gclk));
	jdff dff_B_wosXpw0K0_2(.din(w_dff_B_IMR3K2bM4_2),.dout(w_dff_B_wosXpw0K0_2),.clk(gclk));
	jdff dff_B_hpoS111w6_2(.din(w_dff_B_wosXpw0K0_2),.dout(w_dff_B_hpoS111w6_2),.clk(gclk));
	jdff dff_B_Sr0ExSmE5_2(.din(w_dff_B_hpoS111w6_2),.dout(w_dff_B_Sr0ExSmE5_2),.clk(gclk));
	jdff dff_B_RlCGGr5Y0_2(.din(w_dff_B_Sr0ExSmE5_2),.dout(w_dff_B_RlCGGr5Y0_2),.clk(gclk));
	jdff dff_B_NdHYw2Ji4_1(.din(n1391),.dout(w_dff_B_NdHYw2Ji4_1),.clk(gclk));
	jdff dff_B_U6Ubw3pp7_2(.din(n1312),.dout(w_dff_B_U6Ubw3pp7_2),.clk(gclk));
	jdff dff_B_8y31KhAG1_2(.din(w_dff_B_U6Ubw3pp7_2),.dout(w_dff_B_8y31KhAG1_2),.clk(gclk));
	jdff dff_B_WDuo4Wx99_2(.din(w_dff_B_8y31KhAG1_2),.dout(w_dff_B_WDuo4Wx99_2),.clk(gclk));
	jdff dff_B_wbsBZ0wh1_2(.din(w_dff_B_WDuo4Wx99_2),.dout(w_dff_B_wbsBZ0wh1_2),.clk(gclk));
	jdff dff_B_XQBzbO711_2(.din(w_dff_B_wbsBZ0wh1_2),.dout(w_dff_B_XQBzbO711_2),.clk(gclk));
	jdff dff_B_POkTLrYn1_2(.din(w_dff_B_XQBzbO711_2),.dout(w_dff_B_POkTLrYn1_2),.clk(gclk));
	jdff dff_B_3Z2dZ2y55_2(.din(w_dff_B_POkTLrYn1_2),.dout(w_dff_B_3Z2dZ2y55_2),.clk(gclk));
	jdff dff_B_5C0cvymz5_2(.din(w_dff_B_3Z2dZ2y55_2),.dout(w_dff_B_5C0cvymz5_2),.clk(gclk));
	jdff dff_B_KISb0sGm6_2(.din(w_dff_B_5C0cvymz5_2),.dout(w_dff_B_KISb0sGm6_2),.clk(gclk));
	jdff dff_B_fFfPC3k22_2(.din(w_dff_B_KISb0sGm6_2),.dout(w_dff_B_fFfPC3k22_2),.clk(gclk));
	jdff dff_B_UG0yZ99Q3_2(.din(w_dff_B_fFfPC3k22_2),.dout(w_dff_B_UG0yZ99Q3_2),.clk(gclk));
	jdff dff_B_SLXdx0D89_2(.din(w_dff_B_UG0yZ99Q3_2),.dout(w_dff_B_SLXdx0D89_2),.clk(gclk));
	jdff dff_B_oX0d8D2Y1_2(.din(w_dff_B_SLXdx0D89_2),.dout(w_dff_B_oX0d8D2Y1_2),.clk(gclk));
	jdff dff_B_Mxmc4wt85_2(.din(w_dff_B_oX0d8D2Y1_2),.dout(w_dff_B_Mxmc4wt85_2),.clk(gclk));
	jdff dff_B_mrGCGhk83_2(.din(w_dff_B_Mxmc4wt85_2),.dout(w_dff_B_mrGCGhk83_2),.clk(gclk));
	jdff dff_B_LAW0QPg33_2(.din(w_dff_B_mrGCGhk83_2),.dout(w_dff_B_LAW0QPg33_2),.clk(gclk));
	jdff dff_B_OQrWFPAw2_2(.din(w_dff_B_LAW0QPg33_2),.dout(w_dff_B_OQrWFPAw2_2),.clk(gclk));
	jdff dff_B_gzs3GLYf8_2(.din(w_dff_B_OQrWFPAw2_2),.dout(w_dff_B_gzs3GLYf8_2),.clk(gclk));
	jdff dff_B_D9EZcvwU9_2(.din(w_dff_B_gzs3GLYf8_2),.dout(w_dff_B_D9EZcvwU9_2),.clk(gclk));
	jdff dff_B_kn0MMw319_2(.din(w_dff_B_D9EZcvwU9_2),.dout(w_dff_B_kn0MMw319_2),.clk(gclk));
	jdff dff_B_xyfehsFM1_2(.din(w_dff_B_kn0MMw319_2),.dout(w_dff_B_xyfehsFM1_2),.clk(gclk));
	jdff dff_B_4OmD33P44_2(.din(w_dff_B_xyfehsFM1_2),.dout(w_dff_B_4OmD33P44_2),.clk(gclk));
	jdff dff_B_ONgPNZhT5_2(.din(w_dff_B_4OmD33P44_2),.dout(w_dff_B_ONgPNZhT5_2),.clk(gclk));
	jdff dff_B_hAyWX5ki0_2(.din(w_dff_B_ONgPNZhT5_2),.dout(w_dff_B_hAyWX5ki0_2),.clk(gclk));
	jdff dff_B_29g9LcSI1_2(.din(w_dff_B_hAyWX5ki0_2),.dout(w_dff_B_29g9LcSI1_2),.clk(gclk));
	jdff dff_B_yi1YVyiv9_2(.din(w_dff_B_29g9LcSI1_2),.dout(w_dff_B_yi1YVyiv9_2),.clk(gclk));
	jdff dff_B_MqMIe5CU8_2(.din(w_dff_B_yi1YVyiv9_2),.dout(w_dff_B_MqMIe5CU8_2),.clk(gclk));
	jdff dff_B_MJpMMPUn9_2(.din(w_dff_B_MqMIe5CU8_2),.dout(w_dff_B_MJpMMPUn9_2),.clk(gclk));
	jdff dff_B_WQ9ZA4Bg5_2(.din(w_dff_B_MJpMMPUn9_2),.dout(w_dff_B_WQ9ZA4Bg5_2),.clk(gclk));
	jdff dff_B_T6gQ6IyL3_2(.din(w_dff_B_WQ9ZA4Bg5_2),.dout(w_dff_B_T6gQ6IyL3_2),.clk(gclk));
	jdff dff_B_z4YkEEGY1_2(.din(w_dff_B_T6gQ6IyL3_2),.dout(w_dff_B_z4YkEEGY1_2),.clk(gclk));
	jdff dff_B_YDMz8jpm1_2(.din(w_dff_B_z4YkEEGY1_2),.dout(w_dff_B_YDMz8jpm1_2),.clk(gclk));
	jdff dff_B_S8lu1yTv5_2(.din(w_dff_B_YDMz8jpm1_2),.dout(w_dff_B_S8lu1yTv5_2),.clk(gclk));
	jdff dff_B_EOfLXsNi3_2(.din(w_dff_B_S8lu1yTv5_2),.dout(w_dff_B_EOfLXsNi3_2),.clk(gclk));
	jdff dff_B_DVaSfitn6_2(.din(w_dff_B_EOfLXsNi3_2),.dout(w_dff_B_DVaSfitn6_2),.clk(gclk));
	jdff dff_B_oc45YKuR1_2(.din(w_dff_B_DVaSfitn6_2),.dout(w_dff_B_oc45YKuR1_2),.clk(gclk));
	jdff dff_B_TpuK3uk54_2(.din(w_dff_B_oc45YKuR1_2),.dout(w_dff_B_TpuK3uk54_2),.clk(gclk));
	jdff dff_B_47ENbsaX8_2(.din(w_dff_B_TpuK3uk54_2),.dout(w_dff_B_47ENbsaX8_2),.clk(gclk));
	jdff dff_B_kyZA73wn3_2(.din(w_dff_B_47ENbsaX8_2),.dout(w_dff_B_kyZA73wn3_2),.clk(gclk));
	jdff dff_B_GTCAo03K0_2(.din(w_dff_B_kyZA73wn3_2),.dout(w_dff_B_GTCAo03K0_2),.clk(gclk));
	jdff dff_B_0H3Hy2HC2_1(.din(n1313),.dout(w_dff_B_0H3Hy2HC2_1),.clk(gclk));
	jdff dff_B_WaCNSFAD9_2(.din(n1227),.dout(w_dff_B_WaCNSFAD9_2),.clk(gclk));
	jdff dff_B_MmTj9uej6_2(.din(w_dff_B_WaCNSFAD9_2),.dout(w_dff_B_MmTj9uej6_2),.clk(gclk));
	jdff dff_B_iSPwaqOV4_2(.din(w_dff_B_MmTj9uej6_2),.dout(w_dff_B_iSPwaqOV4_2),.clk(gclk));
	jdff dff_B_IqpecuSu4_2(.din(w_dff_B_iSPwaqOV4_2),.dout(w_dff_B_IqpecuSu4_2),.clk(gclk));
	jdff dff_B_kboR52OL5_2(.din(w_dff_B_IqpecuSu4_2),.dout(w_dff_B_kboR52OL5_2),.clk(gclk));
	jdff dff_B_K1SfeoQm6_2(.din(w_dff_B_kboR52OL5_2),.dout(w_dff_B_K1SfeoQm6_2),.clk(gclk));
	jdff dff_B_UZ6rPx319_2(.din(w_dff_B_K1SfeoQm6_2),.dout(w_dff_B_UZ6rPx319_2),.clk(gclk));
	jdff dff_B_jldKp3rJ3_2(.din(w_dff_B_UZ6rPx319_2),.dout(w_dff_B_jldKp3rJ3_2),.clk(gclk));
	jdff dff_B_VMT8lu7f3_2(.din(w_dff_B_jldKp3rJ3_2),.dout(w_dff_B_VMT8lu7f3_2),.clk(gclk));
	jdff dff_B_koqA6MUA1_2(.din(w_dff_B_VMT8lu7f3_2),.dout(w_dff_B_koqA6MUA1_2),.clk(gclk));
	jdff dff_B_EKJKSklJ0_2(.din(w_dff_B_koqA6MUA1_2),.dout(w_dff_B_EKJKSklJ0_2),.clk(gclk));
	jdff dff_B_Tadc9CTp4_2(.din(w_dff_B_EKJKSklJ0_2),.dout(w_dff_B_Tadc9CTp4_2),.clk(gclk));
	jdff dff_B_9U5ceWEf9_2(.din(w_dff_B_Tadc9CTp4_2),.dout(w_dff_B_9U5ceWEf9_2),.clk(gclk));
	jdff dff_B_bdaHPO2g3_2(.din(w_dff_B_9U5ceWEf9_2),.dout(w_dff_B_bdaHPO2g3_2),.clk(gclk));
	jdff dff_B_5SFXbCKm4_2(.din(w_dff_B_bdaHPO2g3_2),.dout(w_dff_B_5SFXbCKm4_2),.clk(gclk));
	jdff dff_B_vjaOVjhX4_2(.din(w_dff_B_5SFXbCKm4_2),.dout(w_dff_B_vjaOVjhX4_2),.clk(gclk));
	jdff dff_B_tndIYSkn6_2(.din(w_dff_B_vjaOVjhX4_2),.dout(w_dff_B_tndIYSkn6_2),.clk(gclk));
	jdff dff_B_eYQBbDY71_2(.din(w_dff_B_tndIYSkn6_2),.dout(w_dff_B_eYQBbDY71_2),.clk(gclk));
	jdff dff_B_KfRiBqqk7_2(.din(w_dff_B_eYQBbDY71_2),.dout(w_dff_B_KfRiBqqk7_2),.clk(gclk));
	jdff dff_B_sVUntn618_2(.din(w_dff_B_KfRiBqqk7_2),.dout(w_dff_B_sVUntn618_2),.clk(gclk));
	jdff dff_B_5E0S7Mk61_2(.din(w_dff_B_sVUntn618_2),.dout(w_dff_B_5E0S7Mk61_2),.clk(gclk));
	jdff dff_B_AkPqbWMS6_2(.din(w_dff_B_5E0S7Mk61_2),.dout(w_dff_B_AkPqbWMS6_2),.clk(gclk));
	jdff dff_B_T29OzGGi0_2(.din(w_dff_B_AkPqbWMS6_2),.dout(w_dff_B_T29OzGGi0_2),.clk(gclk));
	jdff dff_B_dbHMGxAf7_2(.din(w_dff_B_T29OzGGi0_2),.dout(w_dff_B_dbHMGxAf7_2),.clk(gclk));
	jdff dff_B_VYi3cu8q2_2(.din(w_dff_B_dbHMGxAf7_2),.dout(w_dff_B_VYi3cu8q2_2),.clk(gclk));
	jdff dff_B_og7Gg05P5_2(.din(w_dff_B_VYi3cu8q2_2),.dout(w_dff_B_og7Gg05P5_2),.clk(gclk));
	jdff dff_B_nxteRPeU9_2(.din(w_dff_B_og7Gg05P5_2),.dout(w_dff_B_nxteRPeU9_2),.clk(gclk));
	jdff dff_B_2Q601fps1_2(.din(w_dff_B_nxteRPeU9_2),.dout(w_dff_B_2Q601fps1_2),.clk(gclk));
	jdff dff_B_LKcnht060_2(.din(w_dff_B_2Q601fps1_2),.dout(w_dff_B_LKcnht060_2),.clk(gclk));
	jdff dff_B_mp4znJFi8_2(.din(w_dff_B_LKcnht060_2),.dout(w_dff_B_mp4znJFi8_2),.clk(gclk));
	jdff dff_B_2TX2MUxa8_2(.din(w_dff_B_mp4znJFi8_2),.dout(w_dff_B_2TX2MUxa8_2),.clk(gclk));
	jdff dff_B_ybZWlAH97_2(.din(w_dff_B_2TX2MUxa8_2),.dout(w_dff_B_ybZWlAH97_2),.clk(gclk));
	jdff dff_B_mHMSWxFA9_2(.din(w_dff_B_ybZWlAH97_2),.dout(w_dff_B_mHMSWxFA9_2),.clk(gclk));
	jdff dff_B_o7MXoDFr3_2(.din(w_dff_B_mHMSWxFA9_2),.dout(w_dff_B_o7MXoDFr3_2),.clk(gclk));
	jdff dff_B_khC0GNDL1_2(.din(w_dff_B_o7MXoDFr3_2),.dout(w_dff_B_khC0GNDL1_2),.clk(gclk));
	jdff dff_B_fQN4zX1Q9_2(.din(w_dff_B_khC0GNDL1_2),.dout(w_dff_B_fQN4zX1Q9_2),.clk(gclk));
	jdff dff_B_d8wm2tPJ1_2(.din(w_dff_B_fQN4zX1Q9_2),.dout(w_dff_B_d8wm2tPJ1_2),.clk(gclk));
	jdff dff_B_mv68vdNy4_1(.din(n1228),.dout(w_dff_B_mv68vdNy4_1),.clk(gclk));
	jdff dff_B_N19jddEL1_2(.din(n1136),.dout(w_dff_B_N19jddEL1_2),.clk(gclk));
	jdff dff_B_zCSAdxRo9_2(.din(w_dff_B_N19jddEL1_2),.dout(w_dff_B_zCSAdxRo9_2),.clk(gclk));
	jdff dff_B_k7UHKrmN5_2(.din(w_dff_B_zCSAdxRo9_2),.dout(w_dff_B_k7UHKrmN5_2),.clk(gclk));
	jdff dff_B_QO4Wi0rH7_2(.din(w_dff_B_k7UHKrmN5_2),.dout(w_dff_B_QO4Wi0rH7_2),.clk(gclk));
	jdff dff_B_dlYknYU47_2(.din(w_dff_B_QO4Wi0rH7_2),.dout(w_dff_B_dlYknYU47_2),.clk(gclk));
	jdff dff_B_lf8cTiQT3_2(.din(w_dff_B_dlYknYU47_2),.dout(w_dff_B_lf8cTiQT3_2),.clk(gclk));
	jdff dff_B_jQKFDVaN3_2(.din(w_dff_B_lf8cTiQT3_2),.dout(w_dff_B_jQKFDVaN3_2),.clk(gclk));
	jdff dff_B_819MoxBQ6_2(.din(w_dff_B_jQKFDVaN3_2),.dout(w_dff_B_819MoxBQ6_2),.clk(gclk));
	jdff dff_B_ITXowIf06_2(.din(w_dff_B_819MoxBQ6_2),.dout(w_dff_B_ITXowIf06_2),.clk(gclk));
	jdff dff_B_9KJNCrAw7_2(.din(w_dff_B_ITXowIf06_2),.dout(w_dff_B_9KJNCrAw7_2),.clk(gclk));
	jdff dff_B_ghQBMAJ50_2(.din(w_dff_B_9KJNCrAw7_2),.dout(w_dff_B_ghQBMAJ50_2),.clk(gclk));
	jdff dff_B_crOhpl8S4_2(.din(w_dff_B_ghQBMAJ50_2),.dout(w_dff_B_crOhpl8S4_2),.clk(gclk));
	jdff dff_B_DBwlyrH25_2(.din(w_dff_B_crOhpl8S4_2),.dout(w_dff_B_DBwlyrH25_2),.clk(gclk));
	jdff dff_B_na5gIAp41_2(.din(w_dff_B_DBwlyrH25_2),.dout(w_dff_B_na5gIAp41_2),.clk(gclk));
	jdff dff_B_kvE4x7du9_2(.din(w_dff_B_na5gIAp41_2),.dout(w_dff_B_kvE4x7du9_2),.clk(gclk));
	jdff dff_B_RrvAzQYm0_2(.din(w_dff_B_kvE4x7du9_2),.dout(w_dff_B_RrvAzQYm0_2),.clk(gclk));
	jdff dff_B_1zxwHV1P6_2(.din(w_dff_B_RrvAzQYm0_2),.dout(w_dff_B_1zxwHV1P6_2),.clk(gclk));
	jdff dff_B_C2CwjGL09_2(.din(w_dff_B_1zxwHV1P6_2),.dout(w_dff_B_C2CwjGL09_2),.clk(gclk));
	jdff dff_B_omL9CEEb8_2(.din(w_dff_B_C2CwjGL09_2),.dout(w_dff_B_omL9CEEb8_2),.clk(gclk));
	jdff dff_B_Wv9QBvxG9_2(.din(w_dff_B_omL9CEEb8_2),.dout(w_dff_B_Wv9QBvxG9_2),.clk(gclk));
	jdff dff_B_86qSjaqv5_2(.din(w_dff_B_Wv9QBvxG9_2),.dout(w_dff_B_86qSjaqv5_2),.clk(gclk));
	jdff dff_B_a2EivDk55_2(.din(w_dff_B_86qSjaqv5_2),.dout(w_dff_B_a2EivDk55_2),.clk(gclk));
	jdff dff_B_2wwv2AWA8_2(.din(w_dff_B_a2EivDk55_2),.dout(w_dff_B_2wwv2AWA8_2),.clk(gclk));
	jdff dff_B_zgBzSHyD9_2(.din(w_dff_B_2wwv2AWA8_2),.dout(w_dff_B_zgBzSHyD9_2),.clk(gclk));
	jdff dff_B_OmoqOIOh3_2(.din(w_dff_B_zgBzSHyD9_2),.dout(w_dff_B_OmoqOIOh3_2),.clk(gclk));
	jdff dff_B_aVGXOIuJ0_2(.din(w_dff_B_OmoqOIOh3_2),.dout(w_dff_B_aVGXOIuJ0_2),.clk(gclk));
	jdff dff_B_mn1lX62U7_2(.din(w_dff_B_aVGXOIuJ0_2),.dout(w_dff_B_mn1lX62U7_2),.clk(gclk));
	jdff dff_B_3Yt60LoN1_2(.din(w_dff_B_mn1lX62U7_2),.dout(w_dff_B_3Yt60LoN1_2),.clk(gclk));
	jdff dff_B_zSuTzn4U3_2(.din(w_dff_B_3Yt60LoN1_2),.dout(w_dff_B_zSuTzn4U3_2),.clk(gclk));
	jdff dff_B_7qrznLfw0_2(.din(w_dff_B_zSuTzn4U3_2),.dout(w_dff_B_7qrznLfw0_2),.clk(gclk));
	jdff dff_B_803htx507_2(.din(w_dff_B_7qrznLfw0_2),.dout(w_dff_B_803htx507_2),.clk(gclk));
	jdff dff_B_rVW0ikC74_2(.din(w_dff_B_803htx507_2),.dout(w_dff_B_rVW0ikC74_2),.clk(gclk));
	jdff dff_B_Yl3UZDtS0_2(.din(w_dff_B_rVW0ikC74_2),.dout(w_dff_B_Yl3UZDtS0_2),.clk(gclk));
	jdff dff_B_mhXbmUcO0_2(.din(w_dff_B_Yl3UZDtS0_2),.dout(w_dff_B_mhXbmUcO0_2),.clk(gclk));
	jdff dff_B_RZrP3vIZ0_1(.din(n1137),.dout(w_dff_B_RZrP3vIZ0_1),.clk(gclk));
	jdff dff_B_emabwrZH3_2(.din(n1038),.dout(w_dff_B_emabwrZH3_2),.clk(gclk));
	jdff dff_B_ih9tL02v4_2(.din(w_dff_B_emabwrZH3_2),.dout(w_dff_B_ih9tL02v4_2),.clk(gclk));
	jdff dff_B_8LfxJpnY3_2(.din(w_dff_B_ih9tL02v4_2),.dout(w_dff_B_8LfxJpnY3_2),.clk(gclk));
	jdff dff_B_UnvWLgoe4_2(.din(w_dff_B_8LfxJpnY3_2),.dout(w_dff_B_UnvWLgoe4_2),.clk(gclk));
	jdff dff_B_sXLHwsOj3_2(.din(w_dff_B_UnvWLgoe4_2),.dout(w_dff_B_sXLHwsOj3_2),.clk(gclk));
	jdff dff_B_fJ4Ys15I5_2(.din(w_dff_B_sXLHwsOj3_2),.dout(w_dff_B_fJ4Ys15I5_2),.clk(gclk));
	jdff dff_B_4E0A09X87_2(.din(w_dff_B_fJ4Ys15I5_2),.dout(w_dff_B_4E0A09X87_2),.clk(gclk));
	jdff dff_B_mEMRNyYs0_2(.din(w_dff_B_4E0A09X87_2),.dout(w_dff_B_mEMRNyYs0_2),.clk(gclk));
	jdff dff_B_nX6BpL9K7_2(.din(w_dff_B_mEMRNyYs0_2),.dout(w_dff_B_nX6BpL9K7_2),.clk(gclk));
	jdff dff_B_kU34mXxB5_2(.din(w_dff_B_nX6BpL9K7_2),.dout(w_dff_B_kU34mXxB5_2),.clk(gclk));
	jdff dff_B_CHH1R1PH1_2(.din(w_dff_B_kU34mXxB5_2),.dout(w_dff_B_CHH1R1PH1_2),.clk(gclk));
	jdff dff_B_Z9Krbvwn0_2(.din(w_dff_B_CHH1R1PH1_2),.dout(w_dff_B_Z9Krbvwn0_2),.clk(gclk));
	jdff dff_B_6D06yrvc2_2(.din(w_dff_B_Z9Krbvwn0_2),.dout(w_dff_B_6D06yrvc2_2),.clk(gclk));
	jdff dff_B_evHTy8lh5_2(.din(w_dff_B_6D06yrvc2_2),.dout(w_dff_B_evHTy8lh5_2),.clk(gclk));
	jdff dff_B_tzBsdoiJ9_2(.din(w_dff_B_evHTy8lh5_2),.dout(w_dff_B_tzBsdoiJ9_2),.clk(gclk));
	jdff dff_B_8R8pBGxB7_2(.din(w_dff_B_tzBsdoiJ9_2),.dout(w_dff_B_8R8pBGxB7_2),.clk(gclk));
	jdff dff_B_PJHzxGPt8_2(.din(w_dff_B_8R8pBGxB7_2),.dout(w_dff_B_PJHzxGPt8_2),.clk(gclk));
	jdff dff_B_nkJlaTvE7_2(.din(w_dff_B_PJHzxGPt8_2),.dout(w_dff_B_nkJlaTvE7_2),.clk(gclk));
	jdff dff_B_Dqj2ac0W8_2(.din(w_dff_B_nkJlaTvE7_2),.dout(w_dff_B_Dqj2ac0W8_2),.clk(gclk));
	jdff dff_B_beOFBzPl8_2(.din(w_dff_B_Dqj2ac0W8_2),.dout(w_dff_B_beOFBzPl8_2),.clk(gclk));
	jdff dff_B_PfCkoZLF5_2(.din(w_dff_B_beOFBzPl8_2),.dout(w_dff_B_PfCkoZLF5_2),.clk(gclk));
	jdff dff_B_0vEl2Oyo4_2(.din(w_dff_B_PfCkoZLF5_2),.dout(w_dff_B_0vEl2Oyo4_2),.clk(gclk));
	jdff dff_B_CXTPmEgr7_2(.din(w_dff_B_0vEl2Oyo4_2),.dout(w_dff_B_CXTPmEgr7_2),.clk(gclk));
	jdff dff_B_5xyxvJKs0_2(.din(w_dff_B_CXTPmEgr7_2),.dout(w_dff_B_5xyxvJKs0_2),.clk(gclk));
	jdff dff_B_rvrh4gJu6_2(.din(w_dff_B_5xyxvJKs0_2),.dout(w_dff_B_rvrh4gJu6_2),.clk(gclk));
	jdff dff_B_jIP2ZTtx8_2(.din(w_dff_B_rvrh4gJu6_2),.dout(w_dff_B_jIP2ZTtx8_2),.clk(gclk));
	jdff dff_B_0MXe75ZF6_2(.din(w_dff_B_jIP2ZTtx8_2),.dout(w_dff_B_0MXe75ZF6_2),.clk(gclk));
	jdff dff_B_konae6BJ4_2(.din(w_dff_B_0MXe75ZF6_2),.dout(w_dff_B_konae6BJ4_2),.clk(gclk));
	jdff dff_B_byl4MSlQ5_2(.din(w_dff_B_konae6BJ4_2),.dout(w_dff_B_byl4MSlQ5_2),.clk(gclk));
	jdff dff_B_0BUPneNN4_2(.din(w_dff_B_byl4MSlQ5_2),.dout(w_dff_B_0BUPneNN4_2),.clk(gclk));
	jdff dff_B_rid0auL54_2(.din(w_dff_B_0BUPneNN4_2),.dout(w_dff_B_rid0auL54_2),.clk(gclk));
	jdff dff_B_CB0sktN81_1(.din(n1039),.dout(w_dff_B_CB0sktN81_1),.clk(gclk));
	jdff dff_B_ZuPv0UCP1_2(.din(n939),.dout(w_dff_B_ZuPv0UCP1_2),.clk(gclk));
	jdff dff_B_2PhOPdVE6_2(.din(w_dff_B_ZuPv0UCP1_2),.dout(w_dff_B_2PhOPdVE6_2),.clk(gclk));
	jdff dff_B_eF68Gr4u9_2(.din(w_dff_B_2PhOPdVE6_2),.dout(w_dff_B_eF68Gr4u9_2),.clk(gclk));
	jdff dff_B_OgHyAR9h0_2(.din(w_dff_B_eF68Gr4u9_2),.dout(w_dff_B_OgHyAR9h0_2),.clk(gclk));
	jdff dff_B_ntxEm7ok8_2(.din(w_dff_B_OgHyAR9h0_2),.dout(w_dff_B_ntxEm7ok8_2),.clk(gclk));
	jdff dff_B_Y1pRCgYT7_2(.din(w_dff_B_ntxEm7ok8_2),.dout(w_dff_B_Y1pRCgYT7_2),.clk(gclk));
	jdff dff_B_RQtvvaoB6_2(.din(w_dff_B_Y1pRCgYT7_2),.dout(w_dff_B_RQtvvaoB6_2),.clk(gclk));
	jdff dff_B_FWC5jXQF2_2(.din(w_dff_B_RQtvvaoB6_2),.dout(w_dff_B_FWC5jXQF2_2),.clk(gclk));
	jdff dff_B_CURFQNWl5_2(.din(w_dff_B_FWC5jXQF2_2),.dout(w_dff_B_CURFQNWl5_2),.clk(gclk));
	jdff dff_B_Zfz6R5ip9_2(.din(w_dff_B_CURFQNWl5_2),.dout(w_dff_B_Zfz6R5ip9_2),.clk(gclk));
	jdff dff_B_cI1z6C6B9_2(.din(w_dff_B_Zfz6R5ip9_2),.dout(w_dff_B_cI1z6C6B9_2),.clk(gclk));
	jdff dff_B_WdR5ugpk1_2(.din(w_dff_B_cI1z6C6B9_2),.dout(w_dff_B_WdR5ugpk1_2),.clk(gclk));
	jdff dff_B_5GxzGWHf3_2(.din(w_dff_B_WdR5ugpk1_2),.dout(w_dff_B_5GxzGWHf3_2),.clk(gclk));
	jdff dff_B_ioAtN6GD9_2(.din(w_dff_B_5GxzGWHf3_2),.dout(w_dff_B_ioAtN6GD9_2),.clk(gclk));
	jdff dff_B_NYbpLxkt9_2(.din(w_dff_B_ioAtN6GD9_2),.dout(w_dff_B_NYbpLxkt9_2),.clk(gclk));
	jdff dff_B_vYX7WNda7_2(.din(w_dff_B_NYbpLxkt9_2),.dout(w_dff_B_vYX7WNda7_2),.clk(gclk));
	jdff dff_B_yy1t4VSv5_2(.din(w_dff_B_vYX7WNda7_2),.dout(w_dff_B_yy1t4VSv5_2),.clk(gclk));
	jdff dff_B_BejsI9Wk5_2(.din(w_dff_B_yy1t4VSv5_2),.dout(w_dff_B_BejsI9Wk5_2),.clk(gclk));
	jdff dff_B_7JrZ1iPz7_2(.din(w_dff_B_BejsI9Wk5_2),.dout(w_dff_B_7JrZ1iPz7_2),.clk(gclk));
	jdff dff_B_O86Yp4628_2(.din(w_dff_B_7JrZ1iPz7_2),.dout(w_dff_B_O86Yp4628_2),.clk(gclk));
	jdff dff_B_FBoc3Kks4_2(.din(w_dff_B_O86Yp4628_2),.dout(w_dff_B_FBoc3Kks4_2),.clk(gclk));
	jdff dff_B_UzydEc451_2(.din(w_dff_B_FBoc3Kks4_2),.dout(w_dff_B_UzydEc451_2),.clk(gclk));
	jdff dff_B_790z7C9M9_2(.din(w_dff_B_UzydEc451_2),.dout(w_dff_B_790z7C9M9_2),.clk(gclk));
	jdff dff_B_4prvWc2y5_2(.din(w_dff_B_790z7C9M9_2),.dout(w_dff_B_4prvWc2y5_2),.clk(gclk));
	jdff dff_B_Mgx47BCv9_2(.din(w_dff_B_4prvWc2y5_2),.dout(w_dff_B_Mgx47BCv9_2),.clk(gclk));
	jdff dff_B_otfWY0iH9_2(.din(w_dff_B_Mgx47BCv9_2),.dout(w_dff_B_otfWY0iH9_2),.clk(gclk));
	jdff dff_B_PgAFMw7M5_2(.din(w_dff_B_otfWY0iH9_2),.dout(w_dff_B_PgAFMw7M5_2),.clk(gclk));
	jdff dff_B_guKhFquV9_2(.din(w_dff_B_PgAFMw7M5_2),.dout(w_dff_B_guKhFquV9_2),.clk(gclk));
	jdff dff_B_euu1EETl5_1(.din(n940),.dout(w_dff_B_euu1EETl5_1),.clk(gclk));
	jdff dff_B_140oDg3y9_2(.din(n837),.dout(w_dff_B_140oDg3y9_2),.clk(gclk));
	jdff dff_B_IYsYkObq8_2(.din(w_dff_B_140oDg3y9_2),.dout(w_dff_B_IYsYkObq8_2),.clk(gclk));
	jdff dff_B_foP3H1gP0_2(.din(w_dff_B_IYsYkObq8_2),.dout(w_dff_B_foP3H1gP0_2),.clk(gclk));
	jdff dff_B_u7Z2H9ci5_2(.din(w_dff_B_foP3H1gP0_2),.dout(w_dff_B_u7Z2H9ci5_2),.clk(gclk));
	jdff dff_B_RznP0vOC0_2(.din(w_dff_B_u7Z2H9ci5_2),.dout(w_dff_B_RznP0vOC0_2),.clk(gclk));
	jdff dff_B_IBCdzPW32_2(.din(w_dff_B_RznP0vOC0_2),.dout(w_dff_B_IBCdzPW32_2),.clk(gclk));
	jdff dff_B_KB20gC9q5_2(.din(w_dff_B_IBCdzPW32_2),.dout(w_dff_B_KB20gC9q5_2),.clk(gclk));
	jdff dff_B_S5VAJ7gx7_2(.din(w_dff_B_KB20gC9q5_2),.dout(w_dff_B_S5VAJ7gx7_2),.clk(gclk));
	jdff dff_B_6ftHPquV8_2(.din(w_dff_B_S5VAJ7gx7_2),.dout(w_dff_B_6ftHPquV8_2),.clk(gclk));
	jdff dff_B_Uhkxv0Ek3_2(.din(w_dff_B_6ftHPquV8_2),.dout(w_dff_B_Uhkxv0Ek3_2),.clk(gclk));
	jdff dff_B_GI15IjLD1_2(.din(w_dff_B_Uhkxv0Ek3_2),.dout(w_dff_B_GI15IjLD1_2),.clk(gclk));
	jdff dff_B_lIWNvGbD4_2(.din(w_dff_B_GI15IjLD1_2),.dout(w_dff_B_lIWNvGbD4_2),.clk(gclk));
	jdff dff_B_NWq41bgg1_2(.din(w_dff_B_lIWNvGbD4_2),.dout(w_dff_B_NWq41bgg1_2),.clk(gclk));
	jdff dff_B_8yRuhjn20_2(.din(w_dff_B_NWq41bgg1_2),.dout(w_dff_B_8yRuhjn20_2),.clk(gclk));
	jdff dff_B_Gh9Yabwx6_2(.din(w_dff_B_8yRuhjn20_2),.dout(w_dff_B_Gh9Yabwx6_2),.clk(gclk));
	jdff dff_B_PcXjcuxO7_2(.din(w_dff_B_Gh9Yabwx6_2),.dout(w_dff_B_PcXjcuxO7_2),.clk(gclk));
	jdff dff_B_zjBU6wvI0_2(.din(w_dff_B_PcXjcuxO7_2),.dout(w_dff_B_zjBU6wvI0_2),.clk(gclk));
	jdff dff_B_4wCIEq9L2_2(.din(w_dff_B_zjBU6wvI0_2),.dout(w_dff_B_4wCIEq9L2_2),.clk(gclk));
	jdff dff_B_OeccjMiK7_2(.din(w_dff_B_4wCIEq9L2_2),.dout(w_dff_B_OeccjMiK7_2),.clk(gclk));
	jdff dff_B_BpxqhOfG3_2(.din(w_dff_B_OeccjMiK7_2),.dout(w_dff_B_BpxqhOfG3_2),.clk(gclk));
	jdff dff_B_UVP3n2FV6_2(.din(w_dff_B_BpxqhOfG3_2),.dout(w_dff_B_UVP3n2FV6_2),.clk(gclk));
	jdff dff_B_MHLEkW565_2(.din(w_dff_B_UVP3n2FV6_2),.dout(w_dff_B_MHLEkW565_2),.clk(gclk));
	jdff dff_B_nxEQdo8F8_2(.din(w_dff_B_MHLEkW565_2),.dout(w_dff_B_nxEQdo8F8_2),.clk(gclk));
	jdff dff_B_Xeegg63e1_2(.din(w_dff_B_nxEQdo8F8_2),.dout(w_dff_B_Xeegg63e1_2),.clk(gclk));
	jdff dff_B_M7snh6mM0_2(.din(w_dff_B_Xeegg63e1_2),.dout(w_dff_B_M7snh6mM0_2),.clk(gclk));
	jdff dff_B_80NBw8E22_1(.din(n838),.dout(w_dff_B_80NBw8E22_1),.clk(gclk));
	jdff dff_B_gaHa6Ttn8_2(.din(n739),.dout(w_dff_B_gaHa6Ttn8_2),.clk(gclk));
	jdff dff_B_2qIe3AW63_2(.din(w_dff_B_gaHa6Ttn8_2),.dout(w_dff_B_2qIe3AW63_2),.clk(gclk));
	jdff dff_B_7fImEcFy5_2(.din(w_dff_B_2qIe3AW63_2),.dout(w_dff_B_7fImEcFy5_2),.clk(gclk));
	jdff dff_B_fUmlFteO5_2(.din(w_dff_B_7fImEcFy5_2),.dout(w_dff_B_fUmlFteO5_2),.clk(gclk));
	jdff dff_B_Vi6yQiHF6_2(.din(w_dff_B_fUmlFteO5_2),.dout(w_dff_B_Vi6yQiHF6_2),.clk(gclk));
	jdff dff_B_2rJ3BzyP8_2(.din(w_dff_B_Vi6yQiHF6_2),.dout(w_dff_B_2rJ3BzyP8_2),.clk(gclk));
	jdff dff_B_QfAQvCrZ5_2(.din(w_dff_B_2rJ3BzyP8_2),.dout(w_dff_B_QfAQvCrZ5_2),.clk(gclk));
	jdff dff_B_HbDuMGaU3_2(.din(w_dff_B_QfAQvCrZ5_2),.dout(w_dff_B_HbDuMGaU3_2),.clk(gclk));
	jdff dff_B_b6UI1FgC3_2(.din(w_dff_B_HbDuMGaU3_2),.dout(w_dff_B_b6UI1FgC3_2),.clk(gclk));
	jdff dff_B_2d1ULuW58_2(.din(w_dff_B_b6UI1FgC3_2),.dout(w_dff_B_2d1ULuW58_2),.clk(gclk));
	jdff dff_B_AAan1nW28_2(.din(w_dff_B_2d1ULuW58_2),.dout(w_dff_B_AAan1nW28_2),.clk(gclk));
	jdff dff_B_nEnGV00g8_2(.din(w_dff_B_AAan1nW28_2),.dout(w_dff_B_nEnGV00g8_2),.clk(gclk));
	jdff dff_B_XTBEhzw57_2(.din(w_dff_B_nEnGV00g8_2),.dout(w_dff_B_XTBEhzw57_2),.clk(gclk));
	jdff dff_B_jQLgfyHJ8_2(.din(w_dff_B_XTBEhzw57_2),.dout(w_dff_B_jQLgfyHJ8_2),.clk(gclk));
	jdff dff_B_4PbDtGpy8_2(.din(w_dff_B_jQLgfyHJ8_2),.dout(w_dff_B_4PbDtGpy8_2),.clk(gclk));
	jdff dff_B_61uNtf058_2(.din(w_dff_B_4PbDtGpy8_2),.dout(w_dff_B_61uNtf058_2),.clk(gclk));
	jdff dff_B_mV8Jujk52_2(.din(w_dff_B_61uNtf058_2),.dout(w_dff_B_mV8Jujk52_2),.clk(gclk));
	jdff dff_B_VYrb5c288_2(.din(w_dff_B_mV8Jujk52_2),.dout(w_dff_B_VYrb5c288_2),.clk(gclk));
	jdff dff_B_dwunB3z69_2(.din(w_dff_B_VYrb5c288_2),.dout(w_dff_B_dwunB3z69_2),.clk(gclk));
	jdff dff_B_WfLAAADk9_2(.din(w_dff_B_dwunB3z69_2),.dout(w_dff_B_WfLAAADk9_2),.clk(gclk));
	jdff dff_B_a8fZlPKO3_2(.din(w_dff_B_WfLAAADk9_2),.dout(w_dff_B_a8fZlPKO3_2),.clk(gclk));
	jdff dff_B_cBGvdRqR1_2(.din(w_dff_B_a8fZlPKO3_2),.dout(w_dff_B_cBGvdRqR1_2),.clk(gclk));
	jdff dff_B_hEuuqHdi4_1(.din(n740),.dout(w_dff_B_hEuuqHdi4_1),.clk(gclk));
	jdff dff_B_fbvPWilt2_2(.din(n647),.dout(w_dff_B_fbvPWilt2_2),.clk(gclk));
	jdff dff_B_I5wSJXMr1_2(.din(w_dff_B_fbvPWilt2_2),.dout(w_dff_B_I5wSJXMr1_2),.clk(gclk));
	jdff dff_B_FvnetU492_2(.din(w_dff_B_I5wSJXMr1_2),.dout(w_dff_B_FvnetU492_2),.clk(gclk));
	jdff dff_B_vyl0QTHK9_2(.din(w_dff_B_FvnetU492_2),.dout(w_dff_B_vyl0QTHK9_2),.clk(gclk));
	jdff dff_B_LfhKWCDh7_2(.din(w_dff_B_vyl0QTHK9_2),.dout(w_dff_B_LfhKWCDh7_2),.clk(gclk));
	jdff dff_B_ROchpxLD1_2(.din(w_dff_B_LfhKWCDh7_2),.dout(w_dff_B_ROchpxLD1_2),.clk(gclk));
	jdff dff_B_LJiSSg278_2(.din(w_dff_B_ROchpxLD1_2),.dout(w_dff_B_LJiSSg278_2),.clk(gclk));
	jdff dff_B_ZIoIHeRj5_2(.din(w_dff_B_LJiSSg278_2),.dout(w_dff_B_ZIoIHeRj5_2),.clk(gclk));
	jdff dff_B_8uFlPPON6_2(.din(w_dff_B_ZIoIHeRj5_2),.dout(w_dff_B_8uFlPPON6_2),.clk(gclk));
	jdff dff_B_OJGwLr494_2(.din(w_dff_B_8uFlPPON6_2),.dout(w_dff_B_OJGwLr494_2),.clk(gclk));
	jdff dff_B_ZDhRUGph2_2(.din(w_dff_B_OJGwLr494_2),.dout(w_dff_B_ZDhRUGph2_2),.clk(gclk));
	jdff dff_B_gN3O8cuC7_2(.din(w_dff_B_ZDhRUGph2_2),.dout(w_dff_B_gN3O8cuC7_2),.clk(gclk));
	jdff dff_B_1jTV0hhF5_2(.din(w_dff_B_gN3O8cuC7_2),.dout(w_dff_B_1jTV0hhF5_2),.clk(gclk));
	jdff dff_B_8zK6q8DU3_2(.din(w_dff_B_1jTV0hhF5_2),.dout(w_dff_B_8zK6q8DU3_2),.clk(gclk));
	jdff dff_B_s2CgjbII3_2(.din(w_dff_B_8zK6q8DU3_2),.dout(w_dff_B_s2CgjbII3_2),.clk(gclk));
	jdff dff_B_9yvpeUFL7_2(.din(w_dff_B_s2CgjbII3_2),.dout(w_dff_B_9yvpeUFL7_2),.clk(gclk));
	jdff dff_B_0OlITHCw5_2(.din(w_dff_B_9yvpeUFL7_2),.dout(w_dff_B_0OlITHCw5_2),.clk(gclk));
	jdff dff_B_DetLcREn6_2(.din(w_dff_B_0OlITHCw5_2),.dout(w_dff_B_DetLcREn6_2),.clk(gclk));
	jdff dff_B_i37JVgK58_2(.din(w_dff_B_DetLcREn6_2),.dout(w_dff_B_i37JVgK58_2),.clk(gclk));
	jdff dff_B_X2riWvgE7_1(.din(n648),.dout(w_dff_B_X2riWvgE7_1),.clk(gclk));
	jdff dff_B_RY9wnxnK4_2(.din(n562),.dout(w_dff_B_RY9wnxnK4_2),.clk(gclk));
	jdff dff_B_Pfpbnudr5_2(.din(w_dff_B_RY9wnxnK4_2),.dout(w_dff_B_Pfpbnudr5_2),.clk(gclk));
	jdff dff_B_jQwzLbSu8_2(.din(w_dff_B_Pfpbnudr5_2),.dout(w_dff_B_jQwzLbSu8_2),.clk(gclk));
	jdff dff_B_EN54tcqP5_2(.din(w_dff_B_jQwzLbSu8_2),.dout(w_dff_B_EN54tcqP5_2),.clk(gclk));
	jdff dff_B_JLwThOEh0_2(.din(w_dff_B_EN54tcqP5_2),.dout(w_dff_B_JLwThOEh0_2),.clk(gclk));
	jdff dff_B_OG9oEXUv6_2(.din(w_dff_B_JLwThOEh0_2),.dout(w_dff_B_OG9oEXUv6_2),.clk(gclk));
	jdff dff_B_URsgLQtx1_2(.din(w_dff_B_OG9oEXUv6_2),.dout(w_dff_B_URsgLQtx1_2),.clk(gclk));
	jdff dff_B_nyXakjjf5_2(.din(w_dff_B_URsgLQtx1_2),.dout(w_dff_B_nyXakjjf5_2),.clk(gclk));
	jdff dff_B_yNLoLpNb1_2(.din(w_dff_B_nyXakjjf5_2),.dout(w_dff_B_yNLoLpNb1_2),.clk(gclk));
	jdff dff_B_BzRJ3EN29_2(.din(w_dff_B_yNLoLpNb1_2),.dout(w_dff_B_BzRJ3EN29_2),.clk(gclk));
	jdff dff_B_a9tNjHic7_2(.din(w_dff_B_BzRJ3EN29_2),.dout(w_dff_B_a9tNjHic7_2),.clk(gclk));
	jdff dff_B_bb5Pwi2E8_2(.din(w_dff_B_a9tNjHic7_2),.dout(w_dff_B_bb5Pwi2E8_2),.clk(gclk));
	jdff dff_B_eVeuy8Od2_2(.din(w_dff_B_bb5Pwi2E8_2),.dout(w_dff_B_eVeuy8Od2_2),.clk(gclk));
	jdff dff_B_ZofbYMf14_2(.din(w_dff_B_eVeuy8Od2_2),.dout(w_dff_B_ZofbYMf14_2),.clk(gclk));
	jdff dff_B_ouWBy32k7_2(.din(w_dff_B_ZofbYMf14_2),.dout(w_dff_B_ouWBy32k7_2),.clk(gclk));
	jdff dff_B_HmOy9gdZ6_2(.din(w_dff_B_ouWBy32k7_2),.dout(w_dff_B_HmOy9gdZ6_2),.clk(gclk));
	jdff dff_B_npGZULCR8_1(.din(n563),.dout(w_dff_B_npGZULCR8_1),.clk(gclk));
	jdff dff_B_tP8yLYmi3_2(.din(n484),.dout(w_dff_B_tP8yLYmi3_2),.clk(gclk));
	jdff dff_B_KlMpgy0L5_2(.din(w_dff_B_tP8yLYmi3_2),.dout(w_dff_B_KlMpgy0L5_2),.clk(gclk));
	jdff dff_B_J4eLG92o3_2(.din(w_dff_B_KlMpgy0L5_2),.dout(w_dff_B_J4eLG92o3_2),.clk(gclk));
	jdff dff_B_eNBPa2Nn4_2(.din(w_dff_B_J4eLG92o3_2),.dout(w_dff_B_eNBPa2Nn4_2),.clk(gclk));
	jdff dff_B_CT5KwJnv4_2(.din(w_dff_B_eNBPa2Nn4_2),.dout(w_dff_B_CT5KwJnv4_2),.clk(gclk));
	jdff dff_B_sXqHW34T9_2(.din(w_dff_B_CT5KwJnv4_2),.dout(w_dff_B_sXqHW34T9_2),.clk(gclk));
	jdff dff_B_cWlML1WQ6_2(.din(w_dff_B_sXqHW34T9_2),.dout(w_dff_B_cWlML1WQ6_2),.clk(gclk));
	jdff dff_B_HcahgT2a9_2(.din(w_dff_B_cWlML1WQ6_2),.dout(w_dff_B_HcahgT2a9_2),.clk(gclk));
	jdff dff_B_u1HP4UEW7_2(.din(w_dff_B_HcahgT2a9_2),.dout(w_dff_B_u1HP4UEW7_2),.clk(gclk));
	jdff dff_B_IKWzQX9x2_2(.din(w_dff_B_u1HP4UEW7_2),.dout(w_dff_B_IKWzQX9x2_2),.clk(gclk));
	jdff dff_B_5SQtOB3W8_2(.din(w_dff_B_IKWzQX9x2_2),.dout(w_dff_B_5SQtOB3W8_2),.clk(gclk));
	jdff dff_B_eQOmFkzZ5_2(.din(w_dff_B_5SQtOB3W8_2),.dout(w_dff_B_eQOmFkzZ5_2),.clk(gclk));
	jdff dff_B_fkV0tacZ9_2(.din(w_dff_B_eQOmFkzZ5_2),.dout(w_dff_B_fkV0tacZ9_2),.clk(gclk));
	jdff dff_B_MhBtpbU40_1(.din(n485),.dout(w_dff_B_MhBtpbU40_1),.clk(gclk));
	jdff dff_B_AlzyFC0d4_2(.din(n413),.dout(w_dff_B_AlzyFC0d4_2),.clk(gclk));
	jdff dff_B_cAUyq2nS0_2(.din(w_dff_B_AlzyFC0d4_2),.dout(w_dff_B_cAUyq2nS0_2),.clk(gclk));
	jdff dff_B_nT4RwkNr1_2(.din(w_dff_B_cAUyq2nS0_2),.dout(w_dff_B_nT4RwkNr1_2),.clk(gclk));
	jdff dff_B_4aIHD7BG6_2(.din(w_dff_B_nT4RwkNr1_2),.dout(w_dff_B_4aIHD7BG6_2),.clk(gclk));
	jdff dff_B_kkV6g1UX2_2(.din(w_dff_B_4aIHD7BG6_2),.dout(w_dff_B_kkV6g1UX2_2),.clk(gclk));
	jdff dff_B_0VdfSvSY1_2(.din(w_dff_B_kkV6g1UX2_2),.dout(w_dff_B_0VdfSvSY1_2),.clk(gclk));
	jdff dff_B_D34umgtn8_2(.din(w_dff_B_0VdfSvSY1_2),.dout(w_dff_B_D34umgtn8_2),.clk(gclk));
	jdff dff_B_CDsU8MiW5_2(.din(w_dff_B_D34umgtn8_2),.dout(w_dff_B_CDsU8MiW5_2),.clk(gclk));
	jdff dff_B_3jElJUyu7_2(.din(w_dff_B_CDsU8MiW5_2),.dout(w_dff_B_3jElJUyu7_2),.clk(gclk));
	jdff dff_B_s9XxNWqf5_2(.din(w_dff_B_3jElJUyu7_2),.dout(w_dff_B_s9XxNWqf5_2),.clk(gclk));
	jdff dff_B_L38jzCHb3_2(.din(n416),.dout(w_dff_B_L38jzCHb3_2),.clk(gclk));
	jdff dff_B_hvejbr7D5_1(.din(n414),.dout(w_dff_B_hvejbr7D5_1),.clk(gclk));
	jdff dff_B_sKjMvSKJ5_2(.din(n350),.dout(w_dff_B_sKjMvSKJ5_2),.clk(gclk));
	jdff dff_B_F3xIrhsK2_2(.din(w_dff_B_sKjMvSKJ5_2),.dout(w_dff_B_F3xIrhsK2_2),.clk(gclk));
	jdff dff_B_JQ8vV1Ct7_2(.din(w_dff_B_F3xIrhsK2_2),.dout(w_dff_B_JQ8vV1Ct7_2),.clk(gclk));
	jdff dff_B_mV2s5AHh3_2(.din(w_dff_B_JQ8vV1Ct7_2),.dout(w_dff_B_mV2s5AHh3_2),.clk(gclk));
	jdff dff_B_JJN7KISF6_2(.din(w_dff_B_mV2s5AHh3_2),.dout(w_dff_B_JJN7KISF6_2),.clk(gclk));
	jdff dff_B_lM87nnUQ3_2(.din(w_dff_B_JJN7KISF6_2),.dout(w_dff_B_lM87nnUQ3_2),.clk(gclk));
	jdff dff_B_yrwF1j462_2(.din(n364),.dout(w_dff_B_yrwF1j462_2),.clk(gclk));
	jdff dff_B_8DhbLyL88_2(.din(n295),.dout(w_dff_B_8DhbLyL88_2),.clk(gclk));
	jdff dff_B_h6T7WqZy2_2(.din(w_dff_B_8DhbLyL88_2),.dout(w_dff_B_h6T7WqZy2_2),.clk(gclk));
	jdff dff_B_muOGxhGJ0_2(.din(w_dff_B_h6T7WqZy2_2),.dout(w_dff_B_muOGxhGJ0_2),.clk(gclk));
	jdff dff_B_KO48WI7V7_0(.din(n300),.dout(w_dff_B_KO48WI7V7_0),.clk(gclk));
	jdff dff_A_xjlCJ5fH0_0(.dout(w_n243_0[0]),.din(w_dff_A_xjlCJ5fH0_0),.clk(gclk));
	jdff dff_A_HYTriE2r8_0(.dout(w_dff_A_xjlCJ5fH0_0),.din(w_dff_A_HYTriE2r8_0),.clk(gclk));
	jdff dff_A_X4THlejH0_1(.dout(w_n243_0[1]),.din(w_dff_A_X4THlejH0_1),.clk(gclk));
	jdff dff_A_y8ecDZvJ4_1(.dout(w_dff_A_X4THlejH0_1),.din(w_dff_A_y8ecDZvJ4_1),.clk(gclk));
	jdff dff_B_ro5cP48Y3_1(.din(n1532),.dout(w_dff_B_ro5cP48Y3_1),.clk(gclk));
	jdff dff_B_e9hx0nUu3_2(.din(n1466),.dout(w_dff_B_e9hx0nUu3_2),.clk(gclk));
	jdff dff_B_rxRlKeHn5_2(.din(w_dff_B_e9hx0nUu3_2),.dout(w_dff_B_rxRlKeHn5_2),.clk(gclk));
	jdff dff_B_m3tKkT4H1_2(.din(w_dff_B_rxRlKeHn5_2),.dout(w_dff_B_m3tKkT4H1_2),.clk(gclk));
	jdff dff_B_eojPBsxJ9_2(.din(w_dff_B_m3tKkT4H1_2),.dout(w_dff_B_eojPBsxJ9_2),.clk(gclk));
	jdff dff_B_Aw5oXyTs3_2(.din(w_dff_B_eojPBsxJ9_2),.dout(w_dff_B_Aw5oXyTs3_2),.clk(gclk));
	jdff dff_B_XKXNnmcC7_2(.din(w_dff_B_Aw5oXyTs3_2),.dout(w_dff_B_XKXNnmcC7_2),.clk(gclk));
	jdff dff_B_Qnxulk1J9_2(.din(w_dff_B_XKXNnmcC7_2),.dout(w_dff_B_Qnxulk1J9_2),.clk(gclk));
	jdff dff_B_azXO8WOf0_2(.din(w_dff_B_Qnxulk1J9_2),.dout(w_dff_B_azXO8WOf0_2),.clk(gclk));
	jdff dff_B_x3FjfZDu1_2(.din(w_dff_B_azXO8WOf0_2),.dout(w_dff_B_x3FjfZDu1_2),.clk(gclk));
	jdff dff_B_cHwPmx7o9_2(.din(w_dff_B_x3FjfZDu1_2),.dout(w_dff_B_cHwPmx7o9_2),.clk(gclk));
	jdff dff_B_AunaTG8D8_2(.din(w_dff_B_cHwPmx7o9_2),.dout(w_dff_B_AunaTG8D8_2),.clk(gclk));
	jdff dff_B_IqUEvn7s6_2(.din(w_dff_B_AunaTG8D8_2),.dout(w_dff_B_IqUEvn7s6_2),.clk(gclk));
	jdff dff_B_E2NKaZ5a1_2(.din(w_dff_B_IqUEvn7s6_2),.dout(w_dff_B_E2NKaZ5a1_2),.clk(gclk));
	jdff dff_B_8fH1qxUN0_2(.din(w_dff_B_E2NKaZ5a1_2),.dout(w_dff_B_8fH1qxUN0_2),.clk(gclk));
	jdff dff_B_AXLrF5O73_2(.din(w_dff_B_8fH1qxUN0_2),.dout(w_dff_B_AXLrF5O73_2),.clk(gclk));
	jdff dff_B_Oi2AIzEE4_2(.din(w_dff_B_AXLrF5O73_2),.dout(w_dff_B_Oi2AIzEE4_2),.clk(gclk));
	jdff dff_B_iIs3XRv60_2(.din(w_dff_B_Oi2AIzEE4_2),.dout(w_dff_B_iIs3XRv60_2),.clk(gclk));
	jdff dff_B_Tu1j5mQB1_2(.din(w_dff_B_iIs3XRv60_2),.dout(w_dff_B_Tu1j5mQB1_2),.clk(gclk));
	jdff dff_B_tnlgnleI5_2(.din(w_dff_B_Tu1j5mQB1_2),.dout(w_dff_B_tnlgnleI5_2),.clk(gclk));
	jdff dff_B_XQHYbaeu4_2(.din(w_dff_B_tnlgnleI5_2),.dout(w_dff_B_XQHYbaeu4_2),.clk(gclk));
	jdff dff_B_BLFWJ7ha6_2(.din(w_dff_B_XQHYbaeu4_2),.dout(w_dff_B_BLFWJ7ha6_2),.clk(gclk));
	jdff dff_B_64pBxwNZ7_2(.din(w_dff_B_BLFWJ7ha6_2),.dout(w_dff_B_64pBxwNZ7_2),.clk(gclk));
	jdff dff_B_myrIGuL12_2(.din(w_dff_B_64pBxwNZ7_2),.dout(w_dff_B_myrIGuL12_2),.clk(gclk));
	jdff dff_B_nGXbkOdq6_2(.din(w_dff_B_myrIGuL12_2),.dout(w_dff_B_nGXbkOdq6_2),.clk(gclk));
	jdff dff_B_oe1UKJlG4_2(.din(w_dff_B_nGXbkOdq6_2),.dout(w_dff_B_oe1UKJlG4_2),.clk(gclk));
	jdff dff_B_EF9vJNIh7_2(.din(w_dff_B_oe1UKJlG4_2),.dout(w_dff_B_EF9vJNIh7_2),.clk(gclk));
	jdff dff_B_LPAoNBBK6_2(.din(w_dff_B_EF9vJNIh7_2),.dout(w_dff_B_LPAoNBBK6_2),.clk(gclk));
	jdff dff_B_HTfnSY413_2(.din(w_dff_B_LPAoNBBK6_2),.dout(w_dff_B_HTfnSY413_2),.clk(gclk));
	jdff dff_B_xlbU1lKx0_2(.din(w_dff_B_HTfnSY413_2),.dout(w_dff_B_xlbU1lKx0_2),.clk(gclk));
	jdff dff_B_dGee7S2H7_2(.din(w_dff_B_xlbU1lKx0_2),.dout(w_dff_B_dGee7S2H7_2),.clk(gclk));
	jdff dff_B_hekHXXVp8_2(.din(w_dff_B_dGee7S2H7_2),.dout(w_dff_B_hekHXXVp8_2),.clk(gclk));
	jdff dff_B_rLR9XlKF9_2(.din(w_dff_B_hekHXXVp8_2),.dout(w_dff_B_rLR9XlKF9_2),.clk(gclk));
	jdff dff_B_vBX8i7zp2_2(.din(w_dff_B_rLR9XlKF9_2),.dout(w_dff_B_vBX8i7zp2_2),.clk(gclk));
	jdff dff_B_tf1dHzvh9_2(.din(w_dff_B_vBX8i7zp2_2),.dout(w_dff_B_tf1dHzvh9_2),.clk(gclk));
	jdff dff_B_9LZ5ya752_2(.din(w_dff_B_tf1dHzvh9_2),.dout(w_dff_B_9LZ5ya752_2),.clk(gclk));
	jdff dff_B_062t9TBY1_2(.din(w_dff_B_9LZ5ya752_2),.dout(w_dff_B_062t9TBY1_2),.clk(gclk));
	jdff dff_B_vdsF2kNk9_2(.din(w_dff_B_062t9TBY1_2),.dout(w_dff_B_vdsF2kNk9_2),.clk(gclk));
	jdff dff_B_Xc4cmSKZ7_2(.din(w_dff_B_vdsF2kNk9_2),.dout(w_dff_B_Xc4cmSKZ7_2),.clk(gclk));
	jdff dff_B_TUAjzaQc5_2(.din(w_dff_B_Xc4cmSKZ7_2),.dout(w_dff_B_TUAjzaQc5_2),.clk(gclk));
	jdff dff_B_M1cXpTH12_2(.din(w_dff_B_TUAjzaQc5_2),.dout(w_dff_B_M1cXpTH12_2),.clk(gclk));
	jdff dff_B_9ZJrYBGp7_2(.din(w_dff_B_M1cXpTH12_2),.dout(w_dff_B_9ZJrYBGp7_2),.clk(gclk));
	jdff dff_B_eP63CA6Z8_2(.din(w_dff_B_9ZJrYBGp7_2),.dout(w_dff_B_eP63CA6Z8_2),.clk(gclk));
	jdff dff_B_XbFSq7fE1_2(.din(w_dff_B_eP63CA6Z8_2),.dout(w_dff_B_XbFSq7fE1_2),.clk(gclk));
	jdff dff_B_IESZAlaq7_2(.din(w_dff_B_XbFSq7fE1_2),.dout(w_dff_B_IESZAlaq7_2),.clk(gclk));
	jdff dff_B_lfyc2Dh14_2(.din(w_dff_B_IESZAlaq7_2),.dout(w_dff_B_lfyc2Dh14_2),.clk(gclk));
	jdff dff_B_KmYUFH5k9_2(.din(w_dff_B_lfyc2Dh14_2),.dout(w_dff_B_KmYUFH5k9_2),.clk(gclk));
	jdff dff_B_Ed9BH3408_0(.din(n1531),.dout(w_dff_B_Ed9BH3408_0),.clk(gclk));
	jdff dff_A_zDIQNUSH4_1(.dout(w_n1519_0[1]),.din(w_dff_A_zDIQNUSH4_1),.clk(gclk));
	jdff dff_B_SwruDX775_1(.din(n1467),.dout(w_dff_B_SwruDX775_1),.clk(gclk));
	jdff dff_B_ZFLKPJdI7_2(.din(n1395),.dout(w_dff_B_ZFLKPJdI7_2),.clk(gclk));
	jdff dff_B_5YUTvlny2_2(.din(w_dff_B_ZFLKPJdI7_2),.dout(w_dff_B_5YUTvlny2_2),.clk(gclk));
	jdff dff_B_fVq5IO5Z8_2(.din(w_dff_B_5YUTvlny2_2),.dout(w_dff_B_fVq5IO5Z8_2),.clk(gclk));
	jdff dff_B_UFTdSGGb8_2(.din(w_dff_B_fVq5IO5Z8_2),.dout(w_dff_B_UFTdSGGb8_2),.clk(gclk));
	jdff dff_B_F961kvvd6_2(.din(w_dff_B_UFTdSGGb8_2),.dout(w_dff_B_F961kvvd6_2),.clk(gclk));
	jdff dff_B_2tsZpQrR7_2(.din(w_dff_B_F961kvvd6_2),.dout(w_dff_B_2tsZpQrR7_2),.clk(gclk));
	jdff dff_B_3FqGXqHb6_2(.din(w_dff_B_2tsZpQrR7_2),.dout(w_dff_B_3FqGXqHb6_2),.clk(gclk));
	jdff dff_B_ukePDoKZ0_2(.din(w_dff_B_3FqGXqHb6_2),.dout(w_dff_B_ukePDoKZ0_2),.clk(gclk));
	jdff dff_B_43K46HWJ1_2(.din(w_dff_B_ukePDoKZ0_2),.dout(w_dff_B_43K46HWJ1_2),.clk(gclk));
	jdff dff_B_choCfG798_2(.din(w_dff_B_43K46HWJ1_2),.dout(w_dff_B_choCfG798_2),.clk(gclk));
	jdff dff_B_HB2ovhRj3_2(.din(w_dff_B_choCfG798_2),.dout(w_dff_B_HB2ovhRj3_2),.clk(gclk));
	jdff dff_B_v5Wb0iHJ4_2(.din(w_dff_B_HB2ovhRj3_2),.dout(w_dff_B_v5Wb0iHJ4_2),.clk(gclk));
	jdff dff_B_tV1mwPZ21_2(.din(w_dff_B_v5Wb0iHJ4_2),.dout(w_dff_B_tV1mwPZ21_2),.clk(gclk));
	jdff dff_B_OqHRrrz13_2(.din(w_dff_B_tV1mwPZ21_2),.dout(w_dff_B_OqHRrrz13_2),.clk(gclk));
	jdff dff_B_9znQpidB3_2(.din(w_dff_B_OqHRrrz13_2),.dout(w_dff_B_9znQpidB3_2),.clk(gclk));
	jdff dff_B_8ohYwqSV2_2(.din(w_dff_B_9znQpidB3_2),.dout(w_dff_B_8ohYwqSV2_2),.clk(gclk));
	jdff dff_B_Bf3ow6S36_2(.din(w_dff_B_8ohYwqSV2_2),.dout(w_dff_B_Bf3ow6S36_2),.clk(gclk));
	jdff dff_B_oF1ZgOQ17_2(.din(w_dff_B_Bf3ow6S36_2),.dout(w_dff_B_oF1ZgOQ17_2),.clk(gclk));
	jdff dff_B_UDrsoCEv9_2(.din(w_dff_B_oF1ZgOQ17_2),.dout(w_dff_B_UDrsoCEv9_2),.clk(gclk));
	jdff dff_B_7uFdHyHj5_2(.din(w_dff_B_UDrsoCEv9_2),.dout(w_dff_B_7uFdHyHj5_2),.clk(gclk));
	jdff dff_B_sSDQfO7u7_2(.din(w_dff_B_7uFdHyHj5_2),.dout(w_dff_B_sSDQfO7u7_2),.clk(gclk));
	jdff dff_B_rpZfSjZL3_2(.din(w_dff_B_sSDQfO7u7_2),.dout(w_dff_B_rpZfSjZL3_2),.clk(gclk));
	jdff dff_B_BYMxRWhV9_2(.din(w_dff_B_rpZfSjZL3_2),.dout(w_dff_B_BYMxRWhV9_2),.clk(gclk));
	jdff dff_B_hQpLa3C88_2(.din(w_dff_B_BYMxRWhV9_2),.dout(w_dff_B_hQpLa3C88_2),.clk(gclk));
	jdff dff_B_eOTUKhrR2_2(.din(w_dff_B_hQpLa3C88_2),.dout(w_dff_B_eOTUKhrR2_2),.clk(gclk));
	jdff dff_B_blWOgusu2_2(.din(w_dff_B_eOTUKhrR2_2),.dout(w_dff_B_blWOgusu2_2),.clk(gclk));
	jdff dff_B_aTiybGHH9_2(.din(w_dff_B_blWOgusu2_2),.dout(w_dff_B_aTiybGHH9_2),.clk(gclk));
	jdff dff_B_FZ0vuZHe8_2(.din(w_dff_B_aTiybGHH9_2),.dout(w_dff_B_FZ0vuZHe8_2),.clk(gclk));
	jdff dff_B_igVgbz570_2(.din(w_dff_B_FZ0vuZHe8_2),.dout(w_dff_B_igVgbz570_2),.clk(gclk));
	jdff dff_B_6tRHFwrC0_2(.din(w_dff_B_igVgbz570_2),.dout(w_dff_B_6tRHFwrC0_2),.clk(gclk));
	jdff dff_B_2QzioibU2_2(.din(w_dff_B_6tRHFwrC0_2),.dout(w_dff_B_2QzioibU2_2),.clk(gclk));
	jdff dff_B_7Lal1JNS0_2(.din(w_dff_B_2QzioibU2_2),.dout(w_dff_B_7Lal1JNS0_2),.clk(gclk));
	jdff dff_B_cxwcPxIW9_2(.din(w_dff_B_7Lal1JNS0_2),.dout(w_dff_B_cxwcPxIW9_2),.clk(gclk));
	jdff dff_B_UQiUkEWc3_2(.din(w_dff_B_cxwcPxIW9_2),.dout(w_dff_B_UQiUkEWc3_2),.clk(gclk));
	jdff dff_B_jKip5CG98_2(.din(w_dff_B_UQiUkEWc3_2),.dout(w_dff_B_jKip5CG98_2),.clk(gclk));
	jdff dff_B_LYtwX1wa1_2(.din(w_dff_B_jKip5CG98_2),.dout(w_dff_B_LYtwX1wa1_2),.clk(gclk));
	jdff dff_B_EjwOCjkJ8_2(.din(w_dff_B_LYtwX1wa1_2),.dout(w_dff_B_EjwOCjkJ8_2),.clk(gclk));
	jdff dff_B_P0Z487Ck5_2(.din(w_dff_B_EjwOCjkJ8_2),.dout(w_dff_B_P0Z487Ck5_2),.clk(gclk));
	jdff dff_B_lCGCcQDY8_2(.din(w_dff_B_P0Z487Ck5_2),.dout(w_dff_B_lCGCcQDY8_2),.clk(gclk));
	jdff dff_B_Nzm1NpCa4_2(.din(w_dff_B_lCGCcQDY8_2),.dout(w_dff_B_Nzm1NpCa4_2),.clk(gclk));
	jdff dff_B_jTp396Bm6_2(.din(w_dff_B_Nzm1NpCa4_2),.dout(w_dff_B_jTp396Bm6_2),.clk(gclk));
	jdff dff_B_jfnSrci08_2(.din(n1448),.dout(w_dff_B_jfnSrci08_2),.clk(gclk));
	jdff dff_B_72didT1E7_1(.din(n1396),.dout(w_dff_B_72didT1E7_1),.clk(gclk));
	jdff dff_B_koLmQBVx9_2(.din(n1317),.dout(w_dff_B_koLmQBVx9_2),.clk(gclk));
	jdff dff_B_2NeL1kKh4_2(.din(w_dff_B_koLmQBVx9_2),.dout(w_dff_B_2NeL1kKh4_2),.clk(gclk));
	jdff dff_B_RJ8OZ77n7_2(.din(w_dff_B_2NeL1kKh4_2),.dout(w_dff_B_RJ8OZ77n7_2),.clk(gclk));
	jdff dff_B_f3WxRuip5_2(.din(w_dff_B_RJ8OZ77n7_2),.dout(w_dff_B_f3WxRuip5_2),.clk(gclk));
	jdff dff_B_zUN74IGU2_2(.din(w_dff_B_f3WxRuip5_2),.dout(w_dff_B_zUN74IGU2_2),.clk(gclk));
	jdff dff_B_Ysqbm8bS8_2(.din(w_dff_B_zUN74IGU2_2),.dout(w_dff_B_Ysqbm8bS8_2),.clk(gclk));
	jdff dff_B_91ITMEux7_2(.din(w_dff_B_Ysqbm8bS8_2),.dout(w_dff_B_91ITMEux7_2),.clk(gclk));
	jdff dff_B_sjKZHQDI0_2(.din(w_dff_B_91ITMEux7_2),.dout(w_dff_B_sjKZHQDI0_2),.clk(gclk));
	jdff dff_B_MxphXzJP0_2(.din(w_dff_B_sjKZHQDI0_2),.dout(w_dff_B_MxphXzJP0_2),.clk(gclk));
	jdff dff_B_AarvnL5V8_2(.din(w_dff_B_MxphXzJP0_2),.dout(w_dff_B_AarvnL5V8_2),.clk(gclk));
	jdff dff_B_ICokY8lt5_2(.din(w_dff_B_AarvnL5V8_2),.dout(w_dff_B_ICokY8lt5_2),.clk(gclk));
	jdff dff_B_6Q24a3Lb8_2(.din(w_dff_B_ICokY8lt5_2),.dout(w_dff_B_6Q24a3Lb8_2),.clk(gclk));
	jdff dff_B_HZYMmhHe6_2(.din(w_dff_B_6Q24a3Lb8_2),.dout(w_dff_B_HZYMmhHe6_2),.clk(gclk));
	jdff dff_B_pkwZdyEq5_2(.din(w_dff_B_HZYMmhHe6_2),.dout(w_dff_B_pkwZdyEq5_2),.clk(gclk));
	jdff dff_B_xIGQhoHB5_2(.din(w_dff_B_pkwZdyEq5_2),.dout(w_dff_B_xIGQhoHB5_2),.clk(gclk));
	jdff dff_B_DZdqauXq5_2(.din(w_dff_B_xIGQhoHB5_2),.dout(w_dff_B_DZdqauXq5_2),.clk(gclk));
	jdff dff_B_CaLWwJJC1_2(.din(w_dff_B_DZdqauXq5_2),.dout(w_dff_B_CaLWwJJC1_2),.clk(gclk));
	jdff dff_B_Wbxpflml8_2(.din(w_dff_B_CaLWwJJC1_2),.dout(w_dff_B_Wbxpflml8_2),.clk(gclk));
	jdff dff_B_WltMCCl04_2(.din(w_dff_B_Wbxpflml8_2),.dout(w_dff_B_WltMCCl04_2),.clk(gclk));
	jdff dff_B_YADgxmS45_2(.din(w_dff_B_WltMCCl04_2),.dout(w_dff_B_YADgxmS45_2),.clk(gclk));
	jdff dff_B_AjzUHZIG9_2(.din(w_dff_B_YADgxmS45_2),.dout(w_dff_B_AjzUHZIG9_2),.clk(gclk));
	jdff dff_B_MD0dnGNm8_2(.din(w_dff_B_AjzUHZIG9_2),.dout(w_dff_B_MD0dnGNm8_2),.clk(gclk));
	jdff dff_B_3dZI2tTN6_2(.din(w_dff_B_MD0dnGNm8_2),.dout(w_dff_B_3dZI2tTN6_2),.clk(gclk));
	jdff dff_B_ftYZnWzI9_2(.din(w_dff_B_3dZI2tTN6_2),.dout(w_dff_B_ftYZnWzI9_2),.clk(gclk));
	jdff dff_B_xd2ONGLZ8_2(.din(w_dff_B_ftYZnWzI9_2),.dout(w_dff_B_xd2ONGLZ8_2),.clk(gclk));
	jdff dff_B_iZCDyWct0_2(.din(w_dff_B_xd2ONGLZ8_2),.dout(w_dff_B_iZCDyWct0_2),.clk(gclk));
	jdff dff_B_1K44OmuI2_2(.din(w_dff_B_iZCDyWct0_2),.dout(w_dff_B_1K44OmuI2_2),.clk(gclk));
	jdff dff_B_gc9JE6wK9_2(.din(w_dff_B_1K44OmuI2_2),.dout(w_dff_B_gc9JE6wK9_2),.clk(gclk));
	jdff dff_B_XNKZBaDe0_2(.din(w_dff_B_gc9JE6wK9_2),.dout(w_dff_B_XNKZBaDe0_2),.clk(gclk));
	jdff dff_B_mJ7nhXEv2_2(.din(w_dff_B_XNKZBaDe0_2),.dout(w_dff_B_mJ7nhXEv2_2),.clk(gclk));
	jdff dff_B_Avu5dUl02_2(.din(w_dff_B_mJ7nhXEv2_2),.dout(w_dff_B_Avu5dUl02_2),.clk(gclk));
	jdff dff_B_eZ9ABUN80_2(.din(w_dff_B_Avu5dUl02_2),.dout(w_dff_B_eZ9ABUN80_2),.clk(gclk));
	jdff dff_B_OlrDENrr0_2(.din(w_dff_B_eZ9ABUN80_2),.dout(w_dff_B_OlrDENrr0_2),.clk(gclk));
	jdff dff_B_PJyKYYJK4_2(.din(w_dff_B_OlrDENrr0_2),.dout(w_dff_B_PJyKYYJK4_2),.clk(gclk));
	jdff dff_B_7vwcqmpR6_2(.din(w_dff_B_PJyKYYJK4_2),.dout(w_dff_B_7vwcqmpR6_2),.clk(gclk));
	jdff dff_B_AY4AJOQO3_2(.din(w_dff_B_7vwcqmpR6_2),.dout(w_dff_B_AY4AJOQO3_2),.clk(gclk));
	jdff dff_B_b5ywJgcS4_2(.din(w_dff_B_AY4AJOQO3_2),.dout(w_dff_B_b5ywJgcS4_2),.clk(gclk));
	jdff dff_B_2Kdu6SYs4_2(.din(w_dff_B_b5ywJgcS4_2),.dout(w_dff_B_2Kdu6SYs4_2),.clk(gclk));
	jdff dff_B_SkmqDCMx4_2(.din(n1370),.dout(w_dff_B_SkmqDCMx4_2),.clk(gclk));
	jdff dff_B_m5BQ8Cor6_1(.din(n1318),.dout(w_dff_B_m5BQ8Cor6_1),.clk(gclk));
	jdff dff_B_ZFv2DbFa6_2(.din(n1232),.dout(w_dff_B_ZFv2DbFa6_2),.clk(gclk));
	jdff dff_B_Rgsdhu8z9_2(.din(w_dff_B_ZFv2DbFa6_2),.dout(w_dff_B_Rgsdhu8z9_2),.clk(gclk));
	jdff dff_B_4loedHyv2_2(.din(w_dff_B_Rgsdhu8z9_2),.dout(w_dff_B_4loedHyv2_2),.clk(gclk));
	jdff dff_B_1irYhlm43_2(.din(w_dff_B_4loedHyv2_2),.dout(w_dff_B_1irYhlm43_2),.clk(gclk));
	jdff dff_B_pKp2z2pW6_2(.din(w_dff_B_1irYhlm43_2),.dout(w_dff_B_pKp2z2pW6_2),.clk(gclk));
	jdff dff_B_4vPUwsJy7_2(.din(w_dff_B_pKp2z2pW6_2),.dout(w_dff_B_4vPUwsJy7_2),.clk(gclk));
	jdff dff_B_yW9mvhdH5_2(.din(w_dff_B_4vPUwsJy7_2),.dout(w_dff_B_yW9mvhdH5_2),.clk(gclk));
	jdff dff_B_qppZnRYI5_2(.din(w_dff_B_yW9mvhdH5_2),.dout(w_dff_B_qppZnRYI5_2),.clk(gclk));
	jdff dff_B_eFho2Ocr0_2(.din(w_dff_B_qppZnRYI5_2),.dout(w_dff_B_eFho2Ocr0_2),.clk(gclk));
	jdff dff_B_w6IdzP6c3_2(.din(w_dff_B_eFho2Ocr0_2),.dout(w_dff_B_w6IdzP6c3_2),.clk(gclk));
	jdff dff_B_eDyzI75j0_2(.din(w_dff_B_w6IdzP6c3_2),.dout(w_dff_B_eDyzI75j0_2),.clk(gclk));
	jdff dff_B_7x8o2d7b2_2(.din(w_dff_B_eDyzI75j0_2),.dout(w_dff_B_7x8o2d7b2_2),.clk(gclk));
	jdff dff_B_FsVR2xqC3_2(.din(w_dff_B_7x8o2d7b2_2),.dout(w_dff_B_FsVR2xqC3_2),.clk(gclk));
	jdff dff_B_zdSw8gB36_2(.din(w_dff_B_FsVR2xqC3_2),.dout(w_dff_B_zdSw8gB36_2),.clk(gclk));
	jdff dff_B_x75q6FaY7_2(.din(w_dff_B_zdSw8gB36_2),.dout(w_dff_B_x75q6FaY7_2),.clk(gclk));
	jdff dff_B_WmuiCPUb9_2(.din(w_dff_B_x75q6FaY7_2),.dout(w_dff_B_WmuiCPUb9_2),.clk(gclk));
	jdff dff_B_dMHStHUJ0_2(.din(w_dff_B_WmuiCPUb9_2),.dout(w_dff_B_dMHStHUJ0_2),.clk(gclk));
	jdff dff_B_RF6Zny4U8_2(.din(w_dff_B_dMHStHUJ0_2),.dout(w_dff_B_RF6Zny4U8_2),.clk(gclk));
	jdff dff_B_OWYIk00z9_2(.din(w_dff_B_RF6Zny4U8_2),.dout(w_dff_B_OWYIk00z9_2),.clk(gclk));
	jdff dff_B_DKJTnKOe5_2(.din(w_dff_B_OWYIk00z9_2),.dout(w_dff_B_DKJTnKOe5_2),.clk(gclk));
	jdff dff_B_CJJwGijn9_2(.din(w_dff_B_DKJTnKOe5_2),.dout(w_dff_B_CJJwGijn9_2),.clk(gclk));
	jdff dff_B_rkI5szww7_2(.din(w_dff_B_CJJwGijn9_2),.dout(w_dff_B_rkI5szww7_2),.clk(gclk));
	jdff dff_B_y0d4yNIv7_2(.din(w_dff_B_rkI5szww7_2),.dout(w_dff_B_y0d4yNIv7_2),.clk(gclk));
	jdff dff_B_s6rwE94m2_2(.din(w_dff_B_y0d4yNIv7_2),.dout(w_dff_B_s6rwE94m2_2),.clk(gclk));
	jdff dff_B_mSthmGMl1_2(.din(w_dff_B_s6rwE94m2_2),.dout(w_dff_B_mSthmGMl1_2),.clk(gclk));
	jdff dff_B_dp4bfbII8_2(.din(w_dff_B_mSthmGMl1_2),.dout(w_dff_B_dp4bfbII8_2),.clk(gclk));
	jdff dff_B_BaRpYuK41_2(.din(w_dff_B_dp4bfbII8_2),.dout(w_dff_B_BaRpYuK41_2),.clk(gclk));
	jdff dff_B_b6dAJ7fh2_2(.din(w_dff_B_BaRpYuK41_2),.dout(w_dff_B_b6dAJ7fh2_2),.clk(gclk));
	jdff dff_B_ppyBh3EC0_2(.din(w_dff_B_b6dAJ7fh2_2),.dout(w_dff_B_ppyBh3EC0_2),.clk(gclk));
	jdff dff_B_ZUFVAfxQ6_2(.din(w_dff_B_ppyBh3EC0_2),.dout(w_dff_B_ZUFVAfxQ6_2),.clk(gclk));
	jdff dff_B_pHgVYMsK1_2(.din(w_dff_B_ZUFVAfxQ6_2),.dout(w_dff_B_pHgVYMsK1_2),.clk(gclk));
	jdff dff_B_eDzazIj67_2(.din(w_dff_B_pHgVYMsK1_2),.dout(w_dff_B_eDzazIj67_2),.clk(gclk));
	jdff dff_B_fEp8Xi859_2(.din(w_dff_B_eDzazIj67_2),.dout(w_dff_B_fEp8Xi859_2),.clk(gclk));
	jdff dff_B_bhke1jhb5_2(.din(w_dff_B_fEp8Xi859_2),.dout(w_dff_B_bhke1jhb5_2),.clk(gclk));
	jdff dff_B_Gs5q38Ow6_2(.din(w_dff_B_bhke1jhb5_2),.dout(w_dff_B_Gs5q38Ow6_2),.clk(gclk));
	jdff dff_B_Fhg9wTZk4_2(.din(n1285),.dout(w_dff_B_Fhg9wTZk4_2),.clk(gclk));
	jdff dff_B_uK9k6vOp8_1(.din(n1233),.dout(w_dff_B_uK9k6vOp8_1),.clk(gclk));
	jdff dff_B_YT3Oav0l2_2(.din(n1141),.dout(w_dff_B_YT3Oav0l2_2),.clk(gclk));
	jdff dff_B_n7VUH4rp0_2(.din(w_dff_B_YT3Oav0l2_2),.dout(w_dff_B_n7VUH4rp0_2),.clk(gclk));
	jdff dff_B_tR6z7l7b3_2(.din(w_dff_B_n7VUH4rp0_2),.dout(w_dff_B_tR6z7l7b3_2),.clk(gclk));
	jdff dff_B_gRCHUCka2_2(.din(w_dff_B_tR6z7l7b3_2),.dout(w_dff_B_gRCHUCka2_2),.clk(gclk));
	jdff dff_B_kLCdBYPu0_2(.din(w_dff_B_gRCHUCka2_2),.dout(w_dff_B_kLCdBYPu0_2),.clk(gclk));
	jdff dff_B_LLvt2ApK3_2(.din(w_dff_B_kLCdBYPu0_2),.dout(w_dff_B_LLvt2ApK3_2),.clk(gclk));
	jdff dff_B_1QCdPEgW0_2(.din(w_dff_B_LLvt2ApK3_2),.dout(w_dff_B_1QCdPEgW0_2),.clk(gclk));
	jdff dff_B_EYsZsjDO7_2(.din(w_dff_B_1QCdPEgW0_2),.dout(w_dff_B_EYsZsjDO7_2),.clk(gclk));
	jdff dff_B_YuQ7oVd31_2(.din(w_dff_B_EYsZsjDO7_2),.dout(w_dff_B_YuQ7oVd31_2),.clk(gclk));
	jdff dff_B_m9rjNFu97_2(.din(w_dff_B_YuQ7oVd31_2),.dout(w_dff_B_m9rjNFu97_2),.clk(gclk));
	jdff dff_B_cUt6OpAC0_2(.din(w_dff_B_m9rjNFu97_2),.dout(w_dff_B_cUt6OpAC0_2),.clk(gclk));
	jdff dff_B_h8geLlOu5_2(.din(w_dff_B_cUt6OpAC0_2),.dout(w_dff_B_h8geLlOu5_2),.clk(gclk));
	jdff dff_B_PHxDSOKU6_2(.din(w_dff_B_h8geLlOu5_2),.dout(w_dff_B_PHxDSOKU6_2),.clk(gclk));
	jdff dff_B_7I1OUmOt6_2(.din(w_dff_B_PHxDSOKU6_2),.dout(w_dff_B_7I1OUmOt6_2),.clk(gclk));
	jdff dff_B_LHxuTWIV8_2(.din(w_dff_B_7I1OUmOt6_2),.dout(w_dff_B_LHxuTWIV8_2),.clk(gclk));
	jdff dff_B_iyQbVhyw3_2(.din(w_dff_B_LHxuTWIV8_2),.dout(w_dff_B_iyQbVhyw3_2),.clk(gclk));
	jdff dff_B_cQcIEMFr0_2(.din(w_dff_B_iyQbVhyw3_2),.dout(w_dff_B_cQcIEMFr0_2),.clk(gclk));
	jdff dff_B_hxj5GZfK8_2(.din(w_dff_B_cQcIEMFr0_2),.dout(w_dff_B_hxj5GZfK8_2),.clk(gclk));
	jdff dff_B_RuBPVcm53_2(.din(w_dff_B_hxj5GZfK8_2),.dout(w_dff_B_RuBPVcm53_2),.clk(gclk));
	jdff dff_B_n5h6j43O1_2(.din(w_dff_B_RuBPVcm53_2),.dout(w_dff_B_n5h6j43O1_2),.clk(gclk));
	jdff dff_B_7uNnuhgy3_2(.din(w_dff_B_n5h6j43O1_2),.dout(w_dff_B_7uNnuhgy3_2),.clk(gclk));
	jdff dff_B_vT9CQ6Jv2_2(.din(w_dff_B_7uNnuhgy3_2),.dout(w_dff_B_vT9CQ6Jv2_2),.clk(gclk));
	jdff dff_B_dW60OF9P0_2(.din(w_dff_B_vT9CQ6Jv2_2),.dout(w_dff_B_dW60OF9P0_2),.clk(gclk));
	jdff dff_B_W35zB9hd0_2(.din(w_dff_B_dW60OF9P0_2),.dout(w_dff_B_W35zB9hd0_2),.clk(gclk));
	jdff dff_B_QnuR2BcK0_2(.din(w_dff_B_W35zB9hd0_2),.dout(w_dff_B_QnuR2BcK0_2),.clk(gclk));
	jdff dff_B_W7CSpw3n6_2(.din(w_dff_B_QnuR2BcK0_2),.dout(w_dff_B_W7CSpw3n6_2),.clk(gclk));
	jdff dff_B_yzpa4i1u6_2(.din(w_dff_B_W7CSpw3n6_2),.dout(w_dff_B_yzpa4i1u6_2),.clk(gclk));
	jdff dff_B_mHYYZmXZ5_2(.din(w_dff_B_yzpa4i1u6_2),.dout(w_dff_B_mHYYZmXZ5_2),.clk(gclk));
	jdff dff_B_w1W6beGH7_2(.din(w_dff_B_mHYYZmXZ5_2),.dout(w_dff_B_w1W6beGH7_2),.clk(gclk));
	jdff dff_B_QxvQZhVJ9_2(.din(w_dff_B_w1W6beGH7_2),.dout(w_dff_B_QxvQZhVJ9_2),.clk(gclk));
	jdff dff_B_K6alEr3G9_2(.din(w_dff_B_QxvQZhVJ9_2),.dout(w_dff_B_K6alEr3G9_2),.clk(gclk));
	jdff dff_B_YzDpsTeH8_2(.din(w_dff_B_K6alEr3G9_2),.dout(w_dff_B_YzDpsTeH8_2),.clk(gclk));
	jdff dff_B_mToJob0I8_2(.din(n1194),.dout(w_dff_B_mToJob0I8_2),.clk(gclk));
	jdff dff_B_1LktRM5K5_1(.din(n1142),.dout(w_dff_B_1LktRM5K5_1),.clk(gclk));
	jdff dff_B_J6WTWbRu9_2(.din(n1043),.dout(w_dff_B_J6WTWbRu9_2),.clk(gclk));
	jdff dff_B_6ZHoQYwV3_2(.din(w_dff_B_J6WTWbRu9_2),.dout(w_dff_B_6ZHoQYwV3_2),.clk(gclk));
	jdff dff_B_W1xHsh0Y7_2(.din(w_dff_B_6ZHoQYwV3_2),.dout(w_dff_B_W1xHsh0Y7_2),.clk(gclk));
	jdff dff_B_N8Nrvvdr8_2(.din(w_dff_B_W1xHsh0Y7_2),.dout(w_dff_B_N8Nrvvdr8_2),.clk(gclk));
	jdff dff_B_ZgW69Ha32_2(.din(w_dff_B_N8Nrvvdr8_2),.dout(w_dff_B_ZgW69Ha32_2),.clk(gclk));
	jdff dff_B_966qRKTz0_2(.din(w_dff_B_ZgW69Ha32_2),.dout(w_dff_B_966qRKTz0_2),.clk(gclk));
	jdff dff_B_yxCLSotg3_2(.din(w_dff_B_966qRKTz0_2),.dout(w_dff_B_yxCLSotg3_2),.clk(gclk));
	jdff dff_B_eBvW2OIU5_2(.din(w_dff_B_yxCLSotg3_2),.dout(w_dff_B_eBvW2OIU5_2),.clk(gclk));
	jdff dff_B_fIOEa8zb1_2(.din(w_dff_B_eBvW2OIU5_2),.dout(w_dff_B_fIOEa8zb1_2),.clk(gclk));
	jdff dff_B_bWQjhRvE6_2(.din(w_dff_B_fIOEa8zb1_2),.dout(w_dff_B_bWQjhRvE6_2),.clk(gclk));
	jdff dff_B_Q2f95jkD5_2(.din(w_dff_B_bWQjhRvE6_2),.dout(w_dff_B_Q2f95jkD5_2),.clk(gclk));
	jdff dff_B_AYwitsEW3_2(.din(w_dff_B_Q2f95jkD5_2),.dout(w_dff_B_AYwitsEW3_2),.clk(gclk));
	jdff dff_B_jEKa6cXH1_2(.din(w_dff_B_AYwitsEW3_2),.dout(w_dff_B_jEKa6cXH1_2),.clk(gclk));
	jdff dff_B_TRTSBtWP8_2(.din(w_dff_B_jEKa6cXH1_2),.dout(w_dff_B_TRTSBtWP8_2),.clk(gclk));
	jdff dff_B_GXwVtD863_2(.din(w_dff_B_TRTSBtWP8_2),.dout(w_dff_B_GXwVtD863_2),.clk(gclk));
	jdff dff_B_7606xbX21_2(.din(w_dff_B_GXwVtD863_2),.dout(w_dff_B_7606xbX21_2),.clk(gclk));
	jdff dff_B_9jlg54Nl8_2(.din(w_dff_B_7606xbX21_2),.dout(w_dff_B_9jlg54Nl8_2),.clk(gclk));
	jdff dff_B_7ejpO0pr5_2(.din(w_dff_B_9jlg54Nl8_2),.dout(w_dff_B_7ejpO0pr5_2),.clk(gclk));
	jdff dff_B_izIltxwd8_2(.din(w_dff_B_7ejpO0pr5_2),.dout(w_dff_B_izIltxwd8_2),.clk(gclk));
	jdff dff_B_A6yHRtyG0_2(.din(w_dff_B_izIltxwd8_2),.dout(w_dff_B_A6yHRtyG0_2),.clk(gclk));
	jdff dff_B_D0Mjjkng0_2(.din(w_dff_B_A6yHRtyG0_2),.dout(w_dff_B_D0Mjjkng0_2),.clk(gclk));
	jdff dff_B_IN1IzNOB8_2(.din(w_dff_B_D0Mjjkng0_2),.dout(w_dff_B_IN1IzNOB8_2),.clk(gclk));
	jdff dff_B_qhIPU2ky0_2(.din(w_dff_B_IN1IzNOB8_2),.dout(w_dff_B_qhIPU2ky0_2),.clk(gclk));
	jdff dff_B_3oXBbsWI7_2(.din(w_dff_B_qhIPU2ky0_2),.dout(w_dff_B_3oXBbsWI7_2),.clk(gclk));
	jdff dff_B_YiHYoCaW1_2(.din(w_dff_B_3oXBbsWI7_2),.dout(w_dff_B_YiHYoCaW1_2),.clk(gclk));
	jdff dff_B_GsTU2seh5_2(.din(w_dff_B_YiHYoCaW1_2),.dout(w_dff_B_GsTU2seh5_2),.clk(gclk));
	jdff dff_B_UyWPELAZ8_2(.din(w_dff_B_GsTU2seh5_2),.dout(w_dff_B_UyWPELAZ8_2),.clk(gclk));
	jdff dff_B_miABNWeP6_2(.din(w_dff_B_UyWPELAZ8_2),.dout(w_dff_B_miABNWeP6_2),.clk(gclk));
	jdff dff_B_Y4ySdTZE1_2(.din(w_dff_B_miABNWeP6_2),.dout(w_dff_B_Y4ySdTZE1_2),.clk(gclk));
	jdff dff_B_Y6GAW0cI0_2(.din(n1095),.dout(w_dff_B_Y6GAW0cI0_2),.clk(gclk));
	jdff dff_B_sCOjvpwk7_1(.din(n1044),.dout(w_dff_B_sCOjvpwk7_1),.clk(gclk));
	jdff dff_B_s8t8Y6jC0_2(.din(n944),.dout(w_dff_B_s8t8Y6jC0_2),.clk(gclk));
	jdff dff_B_Fjg59sQk4_2(.din(w_dff_B_s8t8Y6jC0_2),.dout(w_dff_B_Fjg59sQk4_2),.clk(gclk));
	jdff dff_B_NIVnNRD34_2(.din(w_dff_B_Fjg59sQk4_2),.dout(w_dff_B_NIVnNRD34_2),.clk(gclk));
	jdff dff_B_cPctDPIu9_2(.din(w_dff_B_NIVnNRD34_2),.dout(w_dff_B_cPctDPIu9_2),.clk(gclk));
	jdff dff_B_ZDsRNgsI3_2(.din(w_dff_B_cPctDPIu9_2),.dout(w_dff_B_ZDsRNgsI3_2),.clk(gclk));
	jdff dff_B_2kZISSSF4_2(.din(w_dff_B_ZDsRNgsI3_2),.dout(w_dff_B_2kZISSSF4_2),.clk(gclk));
	jdff dff_B_GT4L85wp8_2(.din(w_dff_B_2kZISSSF4_2),.dout(w_dff_B_GT4L85wp8_2),.clk(gclk));
	jdff dff_B_fXI8qcWG4_2(.din(w_dff_B_GT4L85wp8_2),.dout(w_dff_B_fXI8qcWG4_2),.clk(gclk));
	jdff dff_B_3WbCNHrf9_2(.din(w_dff_B_fXI8qcWG4_2),.dout(w_dff_B_3WbCNHrf9_2),.clk(gclk));
	jdff dff_B_3a4zULMd1_2(.din(w_dff_B_3WbCNHrf9_2),.dout(w_dff_B_3a4zULMd1_2),.clk(gclk));
	jdff dff_B_SOBtObaT2_2(.din(w_dff_B_3a4zULMd1_2),.dout(w_dff_B_SOBtObaT2_2),.clk(gclk));
	jdff dff_B_cb9BPlpi5_2(.din(w_dff_B_SOBtObaT2_2),.dout(w_dff_B_cb9BPlpi5_2),.clk(gclk));
	jdff dff_B_mUR7WmDM7_2(.din(w_dff_B_cb9BPlpi5_2),.dout(w_dff_B_mUR7WmDM7_2),.clk(gclk));
	jdff dff_B_85fNOHrM6_2(.din(w_dff_B_mUR7WmDM7_2),.dout(w_dff_B_85fNOHrM6_2),.clk(gclk));
	jdff dff_B_d2lSzW5Z7_2(.din(w_dff_B_85fNOHrM6_2),.dout(w_dff_B_d2lSzW5Z7_2),.clk(gclk));
	jdff dff_B_XyPOo3FA9_2(.din(w_dff_B_d2lSzW5Z7_2),.dout(w_dff_B_XyPOo3FA9_2),.clk(gclk));
	jdff dff_B_iW40ZDY95_2(.din(w_dff_B_XyPOo3FA9_2),.dout(w_dff_B_iW40ZDY95_2),.clk(gclk));
	jdff dff_B_OaECFVQW8_2(.din(w_dff_B_iW40ZDY95_2),.dout(w_dff_B_OaECFVQW8_2),.clk(gclk));
	jdff dff_B_xAsIWQLc4_2(.din(w_dff_B_OaECFVQW8_2),.dout(w_dff_B_xAsIWQLc4_2),.clk(gclk));
	jdff dff_B_68NWWaE34_2(.din(w_dff_B_xAsIWQLc4_2),.dout(w_dff_B_68NWWaE34_2),.clk(gclk));
	jdff dff_B_c5F9Q2IR2_2(.din(w_dff_B_68NWWaE34_2),.dout(w_dff_B_c5F9Q2IR2_2),.clk(gclk));
	jdff dff_B_9TfUHFVB1_2(.din(w_dff_B_c5F9Q2IR2_2),.dout(w_dff_B_9TfUHFVB1_2),.clk(gclk));
	jdff dff_B_qaIPyx9p7_2(.din(w_dff_B_9TfUHFVB1_2),.dout(w_dff_B_qaIPyx9p7_2),.clk(gclk));
	jdff dff_B_3KuNxgML2_2(.din(w_dff_B_qaIPyx9p7_2),.dout(w_dff_B_3KuNxgML2_2),.clk(gclk));
	jdff dff_B_LBV9gPn63_2(.din(w_dff_B_3KuNxgML2_2),.dout(w_dff_B_LBV9gPn63_2),.clk(gclk));
	jdff dff_B_YADlhlg21_2(.din(w_dff_B_LBV9gPn63_2),.dout(w_dff_B_YADlhlg21_2),.clk(gclk));
	jdff dff_B_hc93bl1r7_2(.din(n996),.dout(w_dff_B_hc93bl1r7_2),.clk(gclk));
	jdff dff_B_6kM8FJQY9_1(.din(n945),.dout(w_dff_B_6kM8FJQY9_1),.clk(gclk));
	jdff dff_B_ZyzgSRoN8_2(.din(n842),.dout(w_dff_B_ZyzgSRoN8_2),.clk(gclk));
	jdff dff_B_OUeqsrJM9_2(.din(w_dff_B_ZyzgSRoN8_2),.dout(w_dff_B_OUeqsrJM9_2),.clk(gclk));
	jdff dff_B_jkVpC7Dy5_2(.din(w_dff_B_OUeqsrJM9_2),.dout(w_dff_B_jkVpC7Dy5_2),.clk(gclk));
	jdff dff_B_gkCR23mv0_2(.din(w_dff_B_jkVpC7Dy5_2),.dout(w_dff_B_gkCR23mv0_2),.clk(gclk));
	jdff dff_B_WrIzNfP32_2(.din(w_dff_B_gkCR23mv0_2),.dout(w_dff_B_WrIzNfP32_2),.clk(gclk));
	jdff dff_B_nkJYK7ve5_2(.din(w_dff_B_WrIzNfP32_2),.dout(w_dff_B_nkJYK7ve5_2),.clk(gclk));
	jdff dff_B_hThd8Uot6_2(.din(w_dff_B_nkJYK7ve5_2),.dout(w_dff_B_hThd8Uot6_2),.clk(gclk));
	jdff dff_B_vfo2Y41P6_2(.din(w_dff_B_hThd8Uot6_2),.dout(w_dff_B_vfo2Y41P6_2),.clk(gclk));
	jdff dff_B_qmqbmAq66_2(.din(w_dff_B_vfo2Y41P6_2),.dout(w_dff_B_qmqbmAq66_2),.clk(gclk));
	jdff dff_B_FynjsJbm4_2(.din(w_dff_B_qmqbmAq66_2),.dout(w_dff_B_FynjsJbm4_2),.clk(gclk));
	jdff dff_B_bsGDJrYI3_2(.din(w_dff_B_FynjsJbm4_2),.dout(w_dff_B_bsGDJrYI3_2),.clk(gclk));
	jdff dff_B_zBBQ3SDi4_2(.din(w_dff_B_bsGDJrYI3_2),.dout(w_dff_B_zBBQ3SDi4_2),.clk(gclk));
	jdff dff_B_FyKHuwoQ6_2(.din(w_dff_B_zBBQ3SDi4_2),.dout(w_dff_B_FyKHuwoQ6_2),.clk(gclk));
	jdff dff_B_l2R6oesL6_2(.din(w_dff_B_FyKHuwoQ6_2),.dout(w_dff_B_l2R6oesL6_2),.clk(gclk));
	jdff dff_B_GoeeFxNv9_2(.din(w_dff_B_l2R6oesL6_2),.dout(w_dff_B_GoeeFxNv9_2),.clk(gclk));
	jdff dff_B_zYinyuAT5_2(.din(w_dff_B_GoeeFxNv9_2),.dout(w_dff_B_zYinyuAT5_2),.clk(gclk));
	jdff dff_B_ZZD9bShk4_2(.din(w_dff_B_zYinyuAT5_2),.dout(w_dff_B_ZZD9bShk4_2),.clk(gclk));
	jdff dff_B_tUCneVk78_2(.din(w_dff_B_ZZD9bShk4_2),.dout(w_dff_B_tUCneVk78_2),.clk(gclk));
	jdff dff_B_4x9OCzuh4_2(.din(w_dff_B_tUCneVk78_2),.dout(w_dff_B_4x9OCzuh4_2),.clk(gclk));
	jdff dff_B_wXYqPP6c4_2(.din(w_dff_B_4x9OCzuh4_2),.dout(w_dff_B_wXYqPP6c4_2),.clk(gclk));
	jdff dff_B_LCmPTTOE9_2(.din(w_dff_B_wXYqPP6c4_2),.dout(w_dff_B_LCmPTTOE9_2),.clk(gclk));
	jdff dff_B_VgGuNdZS4_2(.din(w_dff_B_LCmPTTOE9_2),.dout(w_dff_B_VgGuNdZS4_2),.clk(gclk));
	jdff dff_B_WtYEZnw26_2(.din(w_dff_B_VgGuNdZS4_2),.dout(w_dff_B_WtYEZnw26_2),.clk(gclk));
	jdff dff_B_DI2KDhzz3_2(.din(n890),.dout(w_dff_B_DI2KDhzz3_2),.clk(gclk));
	jdff dff_B_i5rvOa3p3_1(.din(n843),.dout(w_dff_B_i5rvOa3p3_1),.clk(gclk));
	jdff dff_B_FGOo59EC6_2(.din(n744),.dout(w_dff_B_FGOo59EC6_2),.clk(gclk));
	jdff dff_B_0BzU38913_2(.din(w_dff_B_FGOo59EC6_2),.dout(w_dff_B_0BzU38913_2),.clk(gclk));
	jdff dff_B_A9EtvMiB6_2(.din(w_dff_B_0BzU38913_2),.dout(w_dff_B_A9EtvMiB6_2),.clk(gclk));
	jdff dff_B_NB5SXZe11_2(.din(w_dff_B_A9EtvMiB6_2),.dout(w_dff_B_NB5SXZe11_2),.clk(gclk));
	jdff dff_B_PxuWLaUL7_2(.din(w_dff_B_NB5SXZe11_2),.dout(w_dff_B_PxuWLaUL7_2),.clk(gclk));
	jdff dff_B_eAv1dQOL5_2(.din(w_dff_B_PxuWLaUL7_2),.dout(w_dff_B_eAv1dQOL5_2),.clk(gclk));
	jdff dff_B_R8wxR1fV5_2(.din(w_dff_B_eAv1dQOL5_2),.dout(w_dff_B_R8wxR1fV5_2),.clk(gclk));
	jdff dff_B_wlcobMyC5_2(.din(w_dff_B_R8wxR1fV5_2),.dout(w_dff_B_wlcobMyC5_2),.clk(gclk));
	jdff dff_B_DjF9SevS9_2(.din(w_dff_B_wlcobMyC5_2),.dout(w_dff_B_DjF9SevS9_2),.clk(gclk));
	jdff dff_B_gH3e6Los9_2(.din(w_dff_B_DjF9SevS9_2),.dout(w_dff_B_gH3e6Los9_2),.clk(gclk));
	jdff dff_B_3MImr5rk7_2(.din(w_dff_B_gH3e6Los9_2),.dout(w_dff_B_3MImr5rk7_2),.clk(gclk));
	jdff dff_B_niBvErOj2_2(.din(w_dff_B_3MImr5rk7_2),.dout(w_dff_B_niBvErOj2_2),.clk(gclk));
	jdff dff_B_uOWDBK3b1_2(.din(w_dff_B_niBvErOj2_2),.dout(w_dff_B_uOWDBK3b1_2),.clk(gclk));
	jdff dff_B_tEm9qimH6_2(.din(w_dff_B_uOWDBK3b1_2),.dout(w_dff_B_tEm9qimH6_2),.clk(gclk));
	jdff dff_B_0lvyRvPs7_2(.din(w_dff_B_tEm9qimH6_2),.dout(w_dff_B_0lvyRvPs7_2),.clk(gclk));
	jdff dff_B_4nU3qPdF6_2(.din(w_dff_B_0lvyRvPs7_2),.dout(w_dff_B_4nU3qPdF6_2),.clk(gclk));
	jdff dff_B_pV06f9Cc4_2(.din(w_dff_B_4nU3qPdF6_2),.dout(w_dff_B_pV06f9Cc4_2),.clk(gclk));
	jdff dff_B_YysPbcvA7_2(.din(w_dff_B_pV06f9Cc4_2),.dout(w_dff_B_YysPbcvA7_2),.clk(gclk));
	jdff dff_B_FuojEz9c7_2(.din(w_dff_B_YysPbcvA7_2),.dout(w_dff_B_FuojEz9c7_2),.clk(gclk));
	jdff dff_B_YF5CjkL67_2(.din(w_dff_B_FuojEz9c7_2),.dout(w_dff_B_YF5CjkL67_2),.clk(gclk));
	jdff dff_B_XofydX4J3_2(.din(n787),.dout(w_dff_B_XofydX4J3_2),.clk(gclk));
	jdff dff_B_cxqTMeGw6_1(.din(n745),.dout(w_dff_B_cxqTMeGw6_1),.clk(gclk));
	jdff dff_B_OYpVKsSp0_2(.din(n652),.dout(w_dff_B_OYpVKsSp0_2),.clk(gclk));
	jdff dff_B_oicXX7277_2(.din(w_dff_B_OYpVKsSp0_2),.dout(w_dff_B_oicXX7277_2),.clk(gclk));
	jdff dff_B_r1U5wM4T0_2(.din(w_dff_B_oicXX7277_2),.dout(w_dff_B_r1U5wM4T0_2),.clk(gclk));
	jdff dff_B_1dXnuMea1_2(.din(w_dff_B_r1U5wM4T0_2),.dout(w_dff_B_1dXnuMea1_2),.clk(gclk));
	jdff dff_B_CW7tpbTA8_2(.din(w_dff_B_1dXnuMea1_2),.dout(w_dff_B_CW7tpbTA8_2),.clk(gclk));
	jdff dff_B_qay6GDby2_2(.din(w_dff_B_CW7tpbTA8_2),.dout(w_dff_B_qay6GDby2_2),.clk(gclk));
	jdff dff_B_S5AWkLQn4_2(.din(w_dff_B_qay6GDby2_2),.dout(w_dff_B_S5AWkLQn4_2),.clk(gclk));
	jdff dff_B_4KoGR2c12_2(.din(w_dff_B_S5AWkLQn4_2),.dout(w_dff_B_4KoGR2c12_2),.clk(gclk));
	jdff dff_B_KtLuIGYF7_2(.din(w_dff_B_4KoGR2c12_2),.dout(w_dff_B_KtLuIGYF7_2),.clk(gclk));
	jdff dff_B_SVOeVH5J3_2(.din(w_dff_B_KtLuIGYF7_2),.dout(w_dff_B_SVOeVH5J3_2),.clk(gclk));
	jdff dff_B_RoFIz7MI8_2(.din(w_dff_B_SVOeVH5J3_2),.dout(w_dff_B_RoFIz7MI8_2),.clk(gclk));
	jdff dff_B_TvaTr2md3_2(.din(w_dff_B_RoFIz7MI8_2),.dout(w_dff_B_TvaTr2md3_2),.clk(gclk));
	jdff dff_B_lsZc9F6t0_2(.din(w_dff_B_TvaTr2md3_2),.dout(w_dff_B_lsZc9F6t0_2),.clk(gclk));
	jdff dff_B_IxLePcrZ7_2(.din(w_dff_B_lsZc9F6t0_2),.dout(w_dff_B_IxLePcrZ7_2),.clk(gclk));
	jdff dff_B_CxQRB3R63_2(.din(w_dff_B_IxLePcrZ7_2),.dout(w_dff_B_CxQRB3R63_2),.clk(gclk));
	jdff dff_B_I7nGwSX22_2(.din(w_dff_B_CxQRB3R63_2),.dout(w_dff_B_I7nGwSX22_2),.clk(gclk));
	jdff dff_B_1HcQjVsl8_2(.din(w_dff_B_I7nGwSX22_2),.dout(w_dff_B_1HcQjVsl8_2),.clk(gclk));
	jdff dff_B_aKw7mzUM2_2(.din(n688),.dout(w_dff_B_aKw7mzUM2_2),.clk(gclk));
	jdff dff_B_iYHSkoAI3_1(.din(n653),.dout(w_dff_B_iYHSkoAI3_1),.clk(gclk));
	jdff dff_B_Mgft5F382_2(.din(n567),.dout(w_dff_B_Mgft5F382_2),.clk(gclk));
	jdff dff_B_G47GsENl3_2(.din(w_dff_B_Mgft5F382_2),.dout(w_dff_B_G47GsENl3_2),.clk(gclk));
	jdff dff_B_VRctDRZy4_2(.din(w_dff_B_G47GsENl3_2),.dout(w_dff_B_VRctDRZy4_2),.clk(gclk));
	jdff dff_B_VdiWadEt1_2(.din(w_dff_B_VRctDRZy4_2),.dout(w_dff_B_VdiWadEt1_2),.clk(gclk));
	jdff dff_B_j5PSWXcg0_2(.din(w_dff_B_VdiWadEt1_2),.dout(w_dff_B_j5PSWXcg0_2),.clk(gclk));
	jdff dff_B_Czwk7QF38_2(.din(w_dff_B_j5PSWXcg0_2),.dout(w_dff_B_Czwk7QF38_2),.clk(gclk));
	jdff dff_B_5hQbSskh1_2(.din(w_dff_B_Czwk7QF38_2),.dout(w_dff_B_5hQbSskh1_2),.clk(gclk));
	jdff dff_B_f8ff7PKS8_2(.din(w_dff_B_5hQbSskh1_2),.dout(w_dff_B_f8ff7PKS8_2),.clk(gclk));
	jdff dff_B_NvncKvTK9_2(.din(w_dff_B_f8ff7PKS8_2),.dout(w_dff_B_NvncKvTK9_2),.clk(gclk));
	jdff dff_B_OLSWtFCH0_2(.din(w_dff_B_NvncKvTK9_2),.dout(w_dff_B_OLSWtFCH0_2),.clk(gclk));
	jdff dff_B_ECyh6JfX5_2(.din(w_dff_B_OLSWtFCH0_2),.dout(w_dff_B_ECyh6JfX5_2),.clk(gclk));
	jdff dff_B_0gSdxCt41_2(.din(w_dff_B_ECyh6JfX5_2),.dout(w_dff_B_0gSdxCt41_2),.clk(gclk));
	jdff dff_B_7UplmbCD0_2(.din(w_dff_B_0gSdxCt41_2),.dout(w_dff_B_7UplmbCD0_2),.clk(gclk));
	jdff dff_B_MuPLUmnB9_2(.din(w_dff_B_7UplmbCD0_2),.dout(w_dff_B_MuPLUmnB9_2),.clk(gclk));
	jdff dff_B_8FZDh62H1_2(.din(n596),.dout(w_dff_B_8FZDh62H1_2),.clk(gclk));
	jdff dff_B_LYvvcZlp2_1(.din(n568),.dout(w_dff_B_LYvvcZlp2_1),.clk(gclk));
	jdff dff_B_NHzErvfo8_2(.din(n489),.dout(w_dff_B_NHzErvfo8_2),.clk(gclk));
	jdff dff_B_Wh6ejkyV2_2(.din(w_dff_B_NHzErvfo8_2),.dout(w_dff_B_Wh6ejkyV2_2),.clk(gclk));
	jdff dff_B_e3MUNzrD9_2(.din(w_dff_B_Wh6ejkyV2_2),.dout(w_dff_B_e3MUNzrD9_2),.clk(gclk));
	jdff dff_B_zEGRgbGm4_2(.din(w_dff_B_e3MUNzrD9_2),.dout(w_dff_B_zEGRgbGm4_2),.clk(gclk));
	jdff dff_B_INOngRA77_2(.din(w_dff_B_zEGRgbGm4_2),.dout(w_dff_B_INOngRA77_2),.clk(gclk));
	jdff dff_B_KBYuhoZD1_2(.din(w_dff_B_INOngRA77_2),.dout(w_dff_B_KBYuhoZD1_2),.clk(gclk));
	jdff dff_B_hPmpx0wQ8_2(.din(w_dff_B_KBYuhoZD1_2),.dout(w_dff_B_hPmpx0wQ8_2),.clk(gclk));
	jdff dff_B_qT4cfSNC8_2(.din(w_dff_B_hPmpx0wQ8_2),.dout(w_dff_B_qT4cfSNC8_2),.clk(gclk));
	jdff dff_B_Be6lNEUY1_2(.din(w_dff_B_qT4cfSNC8_2),.dout(w_dff_B_Be6lNEUY1_2),.clk(gclk));
	jdff dff_B_G90Oi5jn9_2(.din(w_dff_B_Be6lNEUY1_2),.dout(w_dff_B_G90Oi5jn9_2),.clk(gclk));
	jdff dff_B_T7hkcrGP2_2(.din(w_dff_B_G90Oi5jn9_2),.dout(w_dff_B_T7hkcrGP2_2),.clk(gclk));
	jdff dff_B_KbVs6OG40_2(.din(n511),.dout(w_dff_B_KbVs6OG40_2),.clk(gclk));
	jdff dff_B_1Eksn2Zn3_1(.din(n490),.dout(w_dff_B_1Eksn2Zn3_1),.clk(gclk));
	jdff dff_B_O5gyWS1I6_2(.din(n418),.dout(w_dff_B_O5gyWS1I6_2),.clk(gclk));
	jdff dff_B_GvOStkZh7_2(.din(w_dff_B_O5gyWS1I6_2),.dout(w_dff_B_GvOStkZh7_2),.clk(gclk));
	jdff dff_B_QsIJ3ucJ6_2(.din(w_dff_B_GvOStkZh7_2),.dout(w_dff_B_QsIJ3ucJ6_2),.clk(gclk));
	jdff dff_B_4xyshxkA5_2(.din(w_dff_B_QsIJ3ucJ6_2),.dout(w_dff_B_4xyshxkA5_2),.clk(gclk));
	jdff dff_B_KmlJ57ou0_2(.din(w_dff_B_4xyshxkA5_2),.dout(w_dff_B_KmlJ57ou0_2),.clk(gclk));
	jdff dff_B_n4fHl4XQ7_2(.din(w_dff_B_KmlJ57ou0_2),.dout(w_dff_B_n4fHl4XQ7_2),.clk(gclk));
	jdff dff_B_V9mFu0RL1_2(.din(w_dff_B_n4fHl4XQ7_2),.dout(w_dff_B_V9mFu0RL1_2),.clk(gclk));
	jdff dff_B_3M5uY5Tr9_2(.din(w_dff_B_V9mFu0RL1_2),.dout(w_dff_B_3M5uY5Tr9_2),.clk(gclk));
	jdff dff_B_ZaWpwy740_2(.din(n433),.dout(w_dff_B_ZaWpwy740_2),.clk(gclk));
	jdff dff_B_RFwDKia83_2(.din(w_dff_B_ZaWpwy740_2),.dout(w_dff_B_RFwDKia83_2),.clk(gclk));
	jdff dff_B_mS9zbmyi8_2(.din(w_dff_B_RFwDKia83_2),.dout(w_dff_B_mS9zbmyi8_2),.clk(gclk));
	jdff dff_B_VbOJDbnY3_1(.din(n419),.dout(w_dff_B_VbOJDbnY3_1),.clk(gclk));
	jdff dff_B_9n09owlS0_1(.din(w_dff_B_VbOJDbnY3_1),.dout(w_dff_B_9n09owlS0_1),.clk(gclk));
	jdff dff_B_zQnT7X9Y1_2(.din(n356),.dout(w_dff_B_zQnT7X9Y1_2),.clk(gclk));
	jdff dff_B_DGmkYPqP0_2(.din(w_dff_B_zQnT7X9Y1_2),.dout(w_dff_B_DGmkYPqP0_2),.clk(gclk));
	jdff dff_B_E4u52Zoz7_2(.din(w_dff_B_DGmkYPqP0_2),.dout(w_dff_B_E4u52Zoz7_2),.clk(gclk));
	jdff dff_B_x2mpqGpk1_0(.din(n361),.dout(w_dff_B_x2mpqGpk1_0),.clk(gclk));
	jdff dff_A_hG4Qr7px8_0(.dout(w_n297_0[0]),.din(w_dff_A_hG4Qr7px8_0),.clk(gclk));
	jdff dff_A_nqIjHJqT2_0(.dout(w_dff_A_hG4Qr7px8_0),.din(w_dff_A_nqIjHJqT2_0),.clk(gclk));
	jdff dff_A_nHEdJLsC4_1(.dout(w_n297_0[1]),.din(w_dff_A_nHEdJLsC4_1),.clk(gclk));
	jdff dff_A_g1Mpap7a6_1(.dout(w_dff_A_nHEdJLsC4_1),.din(w_dff_A_g1Mpap7a6_1),.clk(gclk));
	jdff dff_B_9t040d6f3_1(.din(n1594),.dout(w_dff_B_9t040d6f3_1),.clk(gclk));
	jdff dff_B_Mev7A2tR5_2(.din(n1535),.dout(w_dff_B_Mev7A2tR5_2),.clk(gclk));
	jdff dff_B_EeKtMkSW3_2(.din(w_dff_B_Mev7A2tR5_2),.dout(w_dff_B_EeKtMkSW3_2),.clk(gclk));
	jdff dff_B_4jql7c3u4_2(.din(w_dff_B_EeKtMkSW3_2),.dout(w_dff_B_4jql7c3u4_2),.clk(gclk));
	jdff dff_B_hntGXt5R9_2(.din(w_dff_B_4jql7c3u4_2),.dout(w_dff_B_hntGXt5R9_2),.clk(gclk));
	jdff dff_B_CfNg9dQo8_2(.din(w_dff_B_hntGXt5R9_2),.dout(w_dff_B_CfNg9dQo8_2),.clk(gclk));
	jdff dff_B_6jojmauz7_2(.din(w_dff_B_CfNg9dQo8_2),.dout(w_dff_B_6jojmauz7_2),.clk(gclk));
	jdff dff_B_yxoYTJqx3_2(.din(w_dff_B_6jojmauz7_2),.dout(w_dff_B_yxoYTJqx3_2),.clk(gclk));
	jdff dff_B_p2NofYur5_2(.din(w_dff_B_yxoYTJqx3_2),.dout(w_dff_B_p2NofYur5_2),.clk(gclk));
	jdff dff_B_bAzpiuRG6_2(.din(w_dff_B_p2NofYur5_2),.dout(w_dff_B_bAzpiuRG6_2),.clk(gclk));
	jdff dff_B_5BKnZWRv1_2(.din(w_dff_B_bAzpiuRG6_2),.dout(w_dff_B_5BKnZWRv1_2),.clk(gclk));
	jdff dff_B_r05j243Y0_2(.din(w_dff_B_5BKnZWRv1_2),.dout(w_dff_B_r05j243Y0_2),.clk(gclk));
	jdff dff_B_kobXswfi0_2(.din(w_dff_B_r05j243Y0_2),.dout(w_dff_B_kobXswfi0_2),.clk(gclk));
	jdff dff_B_RSMXxXds7_2(.din(w_dff_B_kobXswfi0_2),.dout(w_dff_B_RSMXxXds7_2),.clk(gclk));
	jdff dff_B_YGSifZPw2_2(.din(w_dff_B_RSMXxXds7_2),.dout(w_dff_B_YGSifZPw2_2),.clk(gclk));
	jdff dff_B_YNwOSMAk9_2(.din(w_dff_B_YGSifZPw2_2),.dout(w_dff_B_YNwOSMAk9_2),.clk(gclk));
	jdff dff_B_NMYcZaMZ6_2(.din(w_dff_B_YNwOSMAk9_2),.dout(w_dff_B_NMYcZaMZ6_2),.clk(gclk));
	jdff dff_B_l5mBzfNd7_2(.din(w_dff_B_NMYcZaMZ6_2),.dout(w_dff_B_l5mBzfNd7_2),.clk(gclk));
	jdff dff_B_fu7N1rfx6_2(.din(w_dff_B_l5mBzfNd7_2),.dout(w_dff_B_fu7N1rfx6_2),.clk(gclk));
	jdff dff_B_mBDhIcze4_2(.din(w_dff_B_fu7N1rfx6_2),.dout(w_dff_B_mBDhIcze4_2),.clk(gclk));
	jdff dff_B_ISmq8vt38_2(.din(w_dff_B_mBDhIcze4_2),.dout(w_dff_B_ISmq8vt38_2),.clk(gclk));
	jdff dff_B_uMziZcN20_2(.din(w_dff_B_ISmq8vt38_2),.dout(w_dff_B_uMziZcN20_2),.clk(gclk));
	jdff dff_B_HWjKfqSf5_2(.din(w_dff_B_uMziZcN20_2),.dout(w_dff_B_HWjKfqSf5_2),.clk(gclk));
	jdff dff_B_63Qul5YC3_2(.din(w_dff_B_HWjKfqSf5_2),.dout(w_dff_B_63Qul5YC3_2),.clk(gclk));
	jdff dff_B_vCqWrtgW6_2(.din(w_dff_B_63Qul5YC3_2),.dout(w_dff_B_vCqWrtgW6_2),.clk(gclk));
	jdff dff_B_E1YEEBaE3_2(.din(w_dff_B_vCqWrtgW6_2),.dout(w_dff_B_E1YEEBaE3_2),.clk(gclk));
	jdff dff_B_jx82Vfhe2_2(.din(w_dff_B_E1YEEBaE3_2),.dout(w_dff_B_jx82Vfhe2_2),.clk(gclk));
	jdff dff_B_2pLYcsUD1_2(.din(w_dff_B_jx82Vfhe2_2),.dout(w_dff_B_2pLYcsUD1_2),.clk(gclk));
	jdff dff_B_x2wMZitc2_2(.din(w_dff_B_2pLYcsUD1_2),.dout(w_dff_B_x2wMZitc2_2),.clk(gclk));
	jdff dff_B_X6Ml1W8V8_2(.din(w_dff_B_x2wMZitc2_2),.dout(w_dff_B_X6Ml1W8V8_2),.clk(gclk));
	jdff dff_B_MxeULBOb2_2(.din(w_dff_B_X6Ml1W8V8_2),.dout(w_dff_B_MxeULBOb2_2),.clk(gclk));
	jdff dff_B_vzCeqZdo9_2(.din(w_dff_B_MxeULBOb2_2),.dout(w_dff_B_vzCeqZdo9_2),.clk(gclk));
	jdff dff_B_j8gJeYrE7_2(.din(w_dff_B_vzCeqZdo9_2),.dout(w_dff_B_j8gJeYrE7_2),.clk(gclk));
	jdff dff_B_uNiqXae08_2(.din(w_dff_B_j8gJeYrE7_2),.dout(w_dff_B_uNiqXae08_2),.clk(gclk));
	jdff dff_B_lgATJXxJ1_2(.din(w_dff_B_uNiqXae08_2),.dout(w_dff_B_lgATJXxJ1_2),.clk(gclk));
	jdff dff_B_EAoBZrwA9_2(.din(w_dff_B_lgATJXxJ1_2),.dout(w_dff_B_EAoBZrwA9_2),.clk(gclk));
	jdff dff_B_TMgvlIA79_2(.din(w_dff_B_EAoBZrwA9_2),.dout(w_dff_B_TMgvlIA79_2),.clk(gclk));
	jdff dff_B_RrR9zis70_2(.din(w_dff_B_TMgvlIA79_2),.dout(w_dff_B_RrR9zis70_2),.clk(gclk));
	jdff dff_B_GmA4Vr5K0_2(.din(w_dff_B_RrR9zis70_2),.dout(w_dff_B_GmA4Vr5K0_2),.clk(gclk));
	jdff dff_B_jz4ORJk21_2(.din(w_dff_B_GmA4Vr5K0_2),.dout(w_dff_B_jz4ORJk21_2),.clk(gclk));
	jdff dff_B_MO59b8JA7_2(.din(w_dff_B_jz4ORJk21_2),.dout(w_dff_B_MO59b8JA7_2),.clk(gclk));
	jdff dff_B_skBfKhuI0_2(.din(w_dff_B_MO59b8JA7_2),.dout(w_dff_B_skBfKhuI0_2),.clk(gclk));
	jdff dff_B_lTImN72h1_2(.din(w_dff_B_skBfKhuI0_2),.dout(w_dff_B_lTImN72h1_2),.clk(gclk));
	jdff dff_B_PND3Uvmr6_2(.din(w_dff_B_lTImN72h1_2),.dout(w_dff_B_PND3Uvmr6_2),.clk(gclk));
	jdff dff_B_KUj90Kln8_2(.din(w_dff_B_PND3Uvmr6_2),.dout(w_dff_B_KUj90Kln8_2),.clk(gclk));
	jdff dff_B_TiBUXKJU4_2(.din(w_dff_B_KUj90Kln8_2),.dout(w_dff_B_TiBUXKJU4_2),.clk(gclk));
	jdff dff_B_JtkMUbzs3_2(.din(w_dff_B_TiBUXKJU4_2),.dout(w_dff_B_JtkMUbzs3_2),.clk(gclk));
	jdff dff_B_wztV4xSX0_0(.din(n1593),.dout(w_dff_B_wztV4xSX0_0),.clk(gclk));
	jdff dff_A_s2XrVx6R2_1(.dout(w_n1581_0[1]),.din(w_dff_A_s2XrVx6R2_1),.clk(gclk));
	jdff dff_B_mwxOl5mb9_1(.din(n1536),.dout(w_dff_B_mwxOl5mb9_1),.clk(gclk));
	jdff dff_B_wXRiHMXH9_2(.din(n1471),.dout(w_dff_B_wXRiHMXH9_2),.clk(gclk));
	jdff dff_B_a0W6LTZY3_2(.din(w_dff_B_wXRiHMXH9_2),.dout(w_dff_B_a0W6LTZY3_2),.clk(gclk));
	jdff dff_B_gnTokJbh4_2(.din(w_dff_B_a0W6LTZY3_2),.dout(w_dff_B_gnTokJbh4_2),.clk(gclk));
	jdff dff_B_buhPrzya7_2(.din(w_dff_B_gnTokJbh4_2),.dout(w_dff_B_buhPrzya7_2),.clk(gclk));
	jdff dff_B_qmGOzqXB2_2(.din(w_dff_B_buhPrzya7_2),.dout(w_dff_B_qmGOzqXB2_2),.clk(gclk));
	jdff dff_B_2Rwtgp866_2(.din(w_dff_B_qmGOzqXB2_2),.dout(w_dff_B_2Rwtgp866_2),.clk(gclk));
	jdff dff_B_oB3l6RXp6_2(.din(w_dff_B_2Rwtgp866_2),.dout(w_dff_B_oB3l6RXp6_2),.clk(gclk));
	jdff dff_B_6TPLTBmE4_2(.din(w_dff_B_oB3l6RXp6_2),.dout(w_dff_B_6TPLTBmE4_2),.clk(gclk));
	jdff dff_B_iijzvRKa6_2(.din(w_dff_B_6TPLTBmE4_2),.dout(w_dff_B_iijzvRKa6_2),.clk(gclk));
	jdff dff_B_CDmkz72u0_2(.din(w_dff_B_iijzvRKa6_2),.dout(w_dff_B_CDmkz72u0_2),.clk(gclk));
	jdff dff_B_L1abFwff6_2(.din(w_dff_B_CDmkz72u0_2),.dout(w_dff_B_L1abFwff6_2),.clk(gclk));
	jdff dff_B_jpUODlBj1_2(.din(w_dff_B_L1abFwff6_2),.dout(w_dff_B_jpUODlBj1_2),.clk(gclk));
	jdff dff_B_MlXYdS4E5_2(.din(w_dff_B_jpUODlBj1_2),.dout(w_dff_B_MlXYdS4E5_2),.clk(gclk));
	jdff dff_B_zVo3CANZ2_2(.din(w_dff_B_MlXYdS4E5_2),.dout(w_dff_B_zVo3CANZ2_2),.clk(gclk));
	jdff dff_B_Y86smOFu3_2(.din(w_dff_B_zVo3CANZ2_2),.dout(w_dff_B_Y86smOFu3_2),.clk(gclk));
	jdff dff_B_1nIuf5JA9_2(.din(w_dff_B_Y86smOFu3_2),.dout(w_dff_B_1nIuf5JA9_2),.clk(gclk));
	jdff dff_B_F8T7Bx9u6_2(.din(w_dff_B_1nIuf5JA9_2),.dout(w_dff_B_F8T7Bx9u6_2),.clk(gclk));
	jdff dff_B_PBxRXUcp8_2(.din(w_dff_B_F8T7Bx9u6_2),.dout(w_dff_B_PBxRXUcp8_2),.clk(gclk));
	jdff dff_B_HEp7zFMA7_2(.din(w_dff_B_PBxRXUcp8_2),.dout(w_dff_B_HEp7zFMA7_2),.clk(gclk));
	jdff dff_B_dHRQ70XL4_2(.din(w_dff_B_HEp7zFMA7_2),.dout(w_dff_B_dHRQ70XL4_2),.clk(gclk));
	jdff dff_B_sxbtVEAB0_2(.din(w_dff_B_dHRQ70XL4_2),.dout(w_dff_B_sxbtVEAB0_2),.clk(gclk));
	jdff dff_B_lkfgfxll7_2(.din(w_dff_B_sxbtVEAB0_2),.dout(w_dff_B_lkfgfxll7_2),.clk(gclk));
	jdff dff_B_jEj45JqO5_2(.din(w_dff_B_lkfgfxll7_2),.dout(w_dff_B_jEj45JqO5_2),.clk(gclk));
	jdff dff_B_twt6vKDL5_2(.din(w_dff_B_jEj45JqO5_2),.dout(w_dff_B_twt6vKDL5_2),.clk(gclk));
	jdff dff_B_r17X3Flb5_2(.din(w_dff_B_twt6vKDL5_2),.dout(w_dff_B_r17X3Flb5_2),.clk(gclk));
	jdff dff_B_qpDD8kv18_2(.din(w_dff_B_r17X3Flb5_2),.dout(w_dff_B_qpDD8kv18_2),.clk(gclk));
	jdff dff_B_5kpM8K1R9_2(.din(w_dff_B_qpDD8kv18_2),.dout(w_dff_B_5kpM8K1R9_2),.clk(gclk));
	jdff dff_B_J7dseuea3_2(.din(w_dff_B_5kpM8K1R9_2),.dout(w_dff_B_J7dseuea3_2),.clk(gclk));
	jdff dff_B_6DoHxmma1_2(.din(w_dff_B_J7dseuea3_2),.dout(w_dff_B_6DoHxmma1_2),.clk(gclk));
	jdff dff_B_1RVTBdNJ0_2(.din(w_dff_B_6DoHxmma1_2),.dout(w_dff_B_1RVTBdNJ0_2),.clk(gclk));
	jdff dff_B_JE9RxYM24_2(.din(w_dff_B_1RVTBdNJ0_2),.dout(w_dff_B_JE9RxYM24_2),.clk(gclk));
	jdff dff_B_dmxwLxfi2_2(.din(w_dff_B_JE9RxYM24_2),.dout(w_dff_B_dmxwLxfi2_2),.clk(gclk));
	jdff dff_B_V5VCLTH43_2(.din(w_dff_B_dmxwLxfi2_2),.dout(w_dff_B_V5VCLTH43_2),.clk(gclk));
	jdff dff_B_a4osvAmc2_2(.din(w_dff_B_V5VCLTH43_2),.dout(w_dff_B_a4osvAmc2_2),.clk(gclk));
	jdff dff_B_N6AHXkbF5_2(.din(w_dff_B_a4osvAmc2_2),.dout(w_dff_B_N6AHXkbF5_2),.clk(gclk));
	jdff dff_B_O0JhIPw07_2(.din(w_dff_B_N6AHXkbF5_2),.dout(w_dff_B_O0JhIPw07_2),.clk(gclk));
	jdff dff_B_DQHEeKIw4_2(.din(w_dff_B_O0JhIPw07_2),.dout(w_dff_B_DQHEeKIw4_2),.clk(gclk));
	jdff dff_B_kcsrwiPU6_2(.din(w_dff_B_DQHEeKIw4_2),.dout(w_dff_B_kcsrwiPU6_2),.clk(gclk));
	jdff dff_B_L6Rp2KA26_2(.din(w_dff_B_kcsrwiPU6_2),.dout(w_dff_B_L6Rp2KA26_2),.clk(gclk));
	jdff dff_B_npZRYyU75_2(.din(w_dff_B_L6Rp2KA26_2),.dout(w_dff_B_npZRYyU75_2),.clk(gclk));
	jdff dff_B_tdWHgp7n9_2(.din(w_dff_B_npZRYyU75_2),.dout(w_dff_B_tdWHgp7n9_2),.clk(gclk));
	jdff dff_B_wuiWfaLW9_2(.din(n1517),.dout(w_dff_B_wuiWfaLW9_2),.clk(gclk));
	jdff dff_B_zcHUBgZ90_1(.din(n1472),.dout(w_dff_B_zcHUBgZ90_1),.clk(gclk));
	jdff dff_B_8LFVjVyH9_2(.din(n1400),.dout(w_dff_B_8LFVjVyH9_2),.clk(gclk));
	jdff dff_B_DpDWqd1R9_2(.din(w_dff_B_8LFVjVyH9_2),.dout(w_dff_B_DpDWqd1R9_2),.clk(gclk));
	jdff dff_B_FUWQD5aA9_2(.din(w_dff_B_DpDWqd1R9_2),.dout(w_dff_B_FUWQD5aA9_2),.clk(gclk));
	jdff dff_B_CMDEz6jy6_2(.din(w_dff_B_FUWQD5aA9_2),.dout(w_dff_B_CMDEz6jy6_2),.clk(gclk));
	jdff dff_B_o4Qq07tr2_2(.din(w_dff_B_CMDEz6jy6_2),.dout(w_dff_B_o4Qq07tr2_2),.clk(gclk));
	jdff dff_B_pXFwTl3J0_2(.din(w_dff_B_o4Qq07tr2_2),.dout(w_dff_B_pXFwTl3J0_2),.clk(gclk));
	jdff dff_B_SMUDMK8o4_2(.din(w_dff_B_pXFwTl3J0_2),.dout(w_dff_B_SMUDMK8o4_2),.clk(gclk));
	jdff dff_B_tYZcWdYQ0_2(.din(w_dff_B_SMUDMK8o4_2),.dout(w_dff_B_tYZcWdYQ0_2),.clk(gclk));
	jdff dff_B_gcYlqGOP8_2(.din(w_dff_B_tYZcWdYQ0_2),.dout(w_dff_B_gcYlqGOP8_2),.clk(gclk));
	jdff dff_B_rZoHJuAq7_2(.din(w_dff_B_gcYlqGOP8_2),.dout(w_dff_B_rZoHJuAq7_2),.clk(gclk));
	jdff dff_B_GdxRIVTI6_2(.din(w_dff_B_rZoHJuAq7_2),.dout(w_dff_B_GdxRIVTI6_2),.clk(gclk));
	jdff dff_B_wXGjJxQu8_2(.din(w_dff_B_GdxRIVTI6_2),.dout(w_dff_B_wXGjJxQu8_2),.clk(gclk));
	jdff dff_B_Z2TGY7Zb5_2(.din(w_dff_B_wXGjJxQu8_2),.dout(w_dff_B_Z2TGY7Zb5_2),.clk(gclk));
	jdff dff_B_dQJOBsL50_2(.din(w_dff_B_Z2TGY7Zb5_2),.dout(w_dff_B_dQJOBsL50_2),.clk(gclk));
	jdff dff_B_Hwl65rLE5_2(.din(w_dff_B_dQJOBsL50_2),.dout(w_dff_B_Hwl65rLE5_2),.clk(gclk));
	jdff dff_B_iDhMGPT26_2(.din(w_dff_B_Hwl65rLE5_2),.dout(w_dff_B_iDhMGPT26_2),.clk(gclk));
	jdff dff_B_TH1ZTvff4_2(.din(w_dff_B_iDhMGPT26_2),.dout(w_dff_B_TH1ZTvff4_2),.clk(gclk));
	jdff dff_B_MIcxA2Vq0_2(.din(w_dff_B_TH1ZTvff4_2),.dout(w_dff_B_MIcxA2Vq0_2),.clk(gclk));
	jdff dff_B_1gE1HjZl2_2(.din(w_dff_B_MIcxA2Vq0_2),.dout(w_dff_B_1gE1HjZl2_2),.clk(gclk));
	jdff dff_B_Cynb3zst0_2(.din(w_dff_B_1gE1HjZl2_2),.dout(w_dff_B_Cynb3zst0_2),.clk(gclk));
	jdff dff_B_YIwcJRkS7_2(.din(w_dff_B_Cynb3zst0_2),.dout(w_dff_B_YIwcJRkS7_2),.clk(gclk));
	jdff dff_B_gzp6AcP23_2(.din(w_dff_B_YIwcJRkS7_2),.dout(w_dff_B_gzp6AcP23_2),.clk(gclk));
	jdff dff_B_GyGQnDmy6_2(.din(w_dff_B_gzp6AcP23_2),.dout(w_dff_B_GyGQnDmy6_2),.clk(gclk));
	jdff dff_B_Cpaa194s9_2(.din(w_dff_B_GyGQnDmy6_2),.dout(w_dff_B_Cpaa194s9_2),.clk(gclk));
	jdff dff_B_Vscg8Jay6_2(.din(w_dff_B_Cpaa194s9_2),.dout(w_dff_B_Vscg8Jay6_2),.clk(gclk));
	jdff dff_B_vZUcsHqd7_2(.din(w_dff_B_Vscg8Jay6_2),.dout(w_dff_B_vZUcsHqd7_2),.clk(gclk));
	jdff dff_B_4PeIBbgi5_2(.din(w_dff_B_vZUcsHqd7_2),.dout(w_dff_B_4PeIBbgi5_2),.clk(gclk));
	jdff dff_B_a4f51BJZ3_2(.din(w_dff_B_4PeIBbgi5_2),.dout(w_dff_B_a4f51BJZ3_2),.clk(gclk));
	jdff dff_B_EJUCWQe28_2(.din(w_dff_B_a4f51BJZ3_2),.dout(w_dff_B_EJUCWQe28_2),.clk(gclk));
	jdff dff_B_0e1C559U2_2(.din(w_dff_B_EJUCWQe28_2),.dout(w_dff_B_0e1C559U2_2),.clk(gclk));
	jdff dff_B_AdZfayq25_2(.din(w_dff_B_0e1C559U2_2),.dout(w_dff_B_AdZfayq25_2),.clk(gclk));
	jdff dff_B_tfuUpwKE0_2(.din(w_dff_B_AdZfayq25_2),.dout(w_dff_B_tfuUpwKE0_2),.clk(gclk));
	jdff dff_B_2vbQGTsJ6_2(.din(w_dff_B_tfuUpwKE0_2),.dout(w_dff_B_2vbQGTsJ6_2),.clk(gclk));
	jdff dff_B_VZssfK2X6_2(.din(w_dff_B_2vbQGTsJ6_2),.dout(w_dff_B_VZssfK2X6_2),.clk(gclk));
	jdff dff_B_R6LeE3Ft7_2(.din(w_dff_B_VZssfK2X6_2),.dout(w_dff_B_R6LeE3Ft7_2),.clk(gclk));
	jdff dff_B_bljc86PX1_2(.din(w_dff_B_R6LeE3Ft7_2),.dout(w_dff_B_bljc86PX1_2),.clk(gclk));
	jdff dff_B_K8JRXiRX2_2(.din(w_dff_B_bljc86PX1_2),.dout(w_dff_B_K8JRXiRX2_2),.clk(gclk));
	jdff dff_B_lW0kk8354_2(.din(w_dff_B_K8JRXiRX2_2),.dout(w_dff_B_lW0kk8354_2),.clk(gclk));
	jdff dff_B_mbhr9m1M1_2(.din(n1446),.dout(w_dff_B_mbhr9m1M1_2),.clk(gclk));
	jdff dff_B_lqFfUgs60_1(.din(n1401),.dout(w_dff_B_lqFfUgs60_1),.clk(gclk));
	jdff dff_B_KBeKWEJB4_2(.din(n1322),.dout(w_dff_B_KBeKWEJB4_2),.clk(gclk));
	jdff dff_B_JyfXNeKL5_2(.din(w_dff_B_KBeKWEJB4_2),.dout(w_dff_B_JyfXNeKL5_2),.clk(gclk));
	jdff dff_B_qEnCukdO6_2(.din(w_dff_B_JyfXNeKL5_2),.dout(w_dff_B_qEnCukdO6_2),.clk(gclk));
	jdff dff_B_W2Rurbls0_2(.din(w_dff_B_qEnCukdO6_2),.dout(w_dff_B_W2Rurbls0_2),.clk(gclk));
	jdff dff_B_cjfsOv1y8_2(.din(w_dff_B_W2Rurbls0_2),.dout(w_dff_B_cjfsOv1y8_2),.clk(gclk));
	jdff dff_B_qV1g9Prs5_2(.din(w_dff_B_cjfsOv1y8_2),.dout(w_dff_B_qV1g9Prs5_2),.clk(gclk));
	jdff dff_B_ONi6J01R7_2(.din(w_dff_B_qV1g9Prs5_2),.dout(w_dff_B_ONi6J01R7_2),.clk(gclk));
	jdff dff_B_HniIYiJL6_2(.din(w_dff_B_ONi6J01R7_2),.dout(w_dff_B_HniIYiJL6_2),.clk(gclk));
	jdff dff_B_Jmj5DSi88_2(.din(w_dff_B_HniIYiJL6_2),.dout(w_dff_B_Jmj5DSi88_2),.clk(gclk));
	jdff dff_B_dHbY1vWt0_2(.din(w_dff_B_Jmj5DSi88_2),.dout(w_dff_B_dHbY1vWt0_2),.clk(gclk));
	jdff dff_B_wl19Ld9m2_2(.din(w_dff_B_dHbY1vWt0_2),.dout(w_dff_B_wl19Ld9m2_2),.clk(gclk));
	jdff dff_B_85UvMXL87_2(.din(w_dff_B_wl19Ld9m2_2),.dout(w_dff_B_85UvMXL87_2),.clk(gclk));
	jdff dff_B_k3iX4E0i5_2(.din(w_dff_B_85UvMXL87_2),.dout(w_dff_B_k3iX4E0i5_2),.clk(gclk));
	jdff dff_B_Caezq4bY2_2(.din(w_dff_B_k3iX4E0i5_2),.dout(w_dff_B_Caezq4bY2_2),.clk(gclk));
	jdff dff_B_YQrebjQp4_2(.din(w_dff_B_Caezq4bY2_2),.dout(w_dff_B_YQrebjQp4_2),.clk(gclk));
	jdff dff_B_QuE9XNyK1_2(.din(w_dff_B_YQrebjQp4_2),.dout(w_dff_B_QuE9XNyK1_2),.clk(gclk));
	jdff dff_B_I6lkS5e53_2(.din(w_dff_B_QuE9XNyK1_2),.dout(w_dff_B_I6lkS5e53_2),.clk(gclk));
	jdff dff_B_AWynAbvu6_2(.din(w_dff_B_I6lkS5e53_2),.dout(w_dff_B_AWynAbvu6_2),.clk(gclk));
	jdff dff_B_hgs86rlD8_2(.din(w_dff_B_AWynAbvu6_2),.dout(w_dff_B_hgs86rlD8_2),.clk(gclk));
	jdff dff_B_vgPhUIB04_2(.din(w_dff_B_hgs86rlD8_2),.dout(w_dff_B_vgPhUIB04_2),.clk(gclk));
	jdff dff_B_riKux56G7_2(.din(w_dff_B_vgPhUIB04_2),.dout(w_dff_B_riKux56G7_2),.clk(gclk));
	jdff dff_B_bUr5vGjO8_2(.din(w_dff_B_riKux56G7_2),.dout(w_dff_B_bUr5vGjO8_2),.clk(gclk));
	jdff dff_B_M86Ho1Bm1_2(.din(w_dff_B_bUr5vGjO8_2),.dout(w_dff_B_M86Ho1Bm1_2),.clk(gclk));
	jdff dff_B_m5GmsNR90_2(.din(w_dff_B_M86Ho1Bm1_2),.dout(w_dff_B_m5GmsNR90_2),.clk(gclk));
	jdff dff_B_bL3vy8Vl6_2(.din(w_dff_B_m5GmsNR90_2),.dout(w_dff_B_bL3vy8Vl6_2),.clk(gclk));
	jdff dff_B_m2sC1NEV4_2(.din(w_dff_B_bL3vy8Vl6_2),.dout(w_dff_B_m2sC1NEV4_2),.clk(gclk));
	jdff dff_B_1jNKTHhZ1_2(.din(w_dff_B_m2sC1NEV4_2),.dout(w_dff_B_1jNKTHhZ1_2),.clk(gclk));
	jdff dff_B_llysxnyL1_2(.din(w_dff_B_1jNKTHhZ1_2),.dout(w_dff_B_llysxnyL1_2),.clk(gclk));
	jdff dff_B_Lq9rmOH56_2(.din(w_dff_B_llysxnyL1_2),.dout(w_dff_B_Lq9rmOH56_2),.clk(gclk));
	jdff dff_B_W4zzFZB87_2(.din(w_dff_B_Lq9rmOH56_2),.dout(w_dff_B_W4zzFZB87_2),.clk(gclk));
	jdff dff_B_AFp6Rvfp9_2(.din(w_dff_B_W4zzFZB87_2),.dout(w_dff_B_AFp6Rvfp9_2),.clk(gclk));
	jdff dff_B_sJztinWD0_2(.din(w_dff_B_AFp6Rvfp9_2),.dout(w_dff_B_sJztinWD0_2),.clk(gclk));
	jdff dff_B_HKctigfB6_2(.din(w_dff_B_sJztinWD0_2),.dout(w_dff_B_HKctigfB6_2),.clk(gclk));
	jdff dff_B_GTtQcLjM1_2(.din(w_dff_B_HKctigfB6_2),.dout(w_dff_B_GTtQcLjM1_2),.clk(gclk));
	jdff dff_B_1yz24uV28_2(.din(w_dff_B_GTtQcLjM1_2),.dout(w_dff_B_1yz24uV28_2),.clk(gclk));
	jdff dff_B_FRdNxege6_2(.din(n1368),.dout(w_dff_B_FRdNxege6_2),.clk(gclk));
	jdff dff_B_1MmuV6Vb7_1(.din(n1323),.dout(w_dff_B_1MmuV6Vb7_1),.clk(gclk));
	jdff dff_B_2qajahL00_2(.din(n1237),.dout(w_dff_B_2qajahL00_2),.clk(gclk));
	jdff dff_B_zx5zGZ3z5_2(.din(w_dff_B_2qajahL00_2),.dout(w_dff_B_zx5zGZ3z5_2),.clk(gclk));
	jdff dff_B_qkXnfkjC3_2(.din(w_dff_B_zx5zGZ3z5_2),.dout(w_dff_B_qkXnfkjC3_2),.clk(gclk));
	jdff dff_B_QW1dHc2r4_2(.din(w_dff_B_qkXnfkjC3_2),.dout(w_dff_B_QW1dHc2r4_2),.clk(gclk));
	jdff dff_B_qXvLha4E2_2(.din(w_dff_B_QW1dHc2r4_2),.dout(w_dff_B_qXvLha4E2_2),.clk(gclk));
	jdff dff_B_VeBiJPly0_2(.din(w_dff_B_qXvLha4E2_2),.dout(w_dff_B_VeBiJPly0_2),.clk(gclk));
	jdff dff_B_QhKmzk4d2_2(.din(w_dff_B_VeBiJPly0_2),.dout(w_dff_B_QhKmzk4d2_2),.clk(gclk));
	jdff dff_B_xf8nfrmz8_2(.din(w_dff_B_QhKmzk4d2_2),.dout(w_dff_B_xf8nfrmz8_2),.clk(gclk));
	jdff dff_B_Amj9SR2e0_2(.din(w_dff_B_xf8nfrmz8_2),.dout(w_dff_B_Amj9SR2e0_2),.clk(gclk));
	jdff dff_B_yQXeHfFn3_2(.din(w_dff_B_Amj9SR2e0_2),.dout(w_dff_B_yQXeHfFn3_2),.clk(gclk));
	jdff dff_B_3YCtFFb71_2(.din(w_dff_B_yQXeHfFn3_2),.dout(w_dff_B_3YCtFFb71_2),.clk(gclk));
	jdff dff_B_4i5y2rlA0_2(.din(w_dff_B_3YCtFFb71_2),.dout(w_dff_B_4i5y2rlA0_2),.clk(gclk));
	jdff dff_B_FzeFKLdv1_2(.din(w_dff_B_4i5y2rlA0_2),.dout(w_dff_B_FzeFKLdv1_2),.clk(gclk));
	jdff dff_B_9fHz8tE97_2(.din(w_dff_B_FzeFKLdv1_2),.dout(w_dff_B_9fHz8tE97_2),.clk(gclk));
	jdff dff_B_kmk8lekL2_2(.din(w_dff_B_9fHz8tE97_2),.dout(w_dff_B_kmk8lekL2_2),.clk(gclk));
	jdff dff_B_3SClmbQ98_2(.din(w_dff_B_kmk8lekL2_2),.dout(w_dff_B_3SClmbQ98_2),.clk(gclk));
	jdff dff_B_xAnIGToR2_2(.din(w_dff_B_3SClmbQ98_2),.dout(w_dff_B_xAnIGToR2_2),.clk(gclk));
	jdff dff_B_Qlcq6qvH2_2(.din(w_dff_B_xAnIGToR2_2),.dout(w_dff_B_Qlcq6qvH2_2),.clk(gclk));
	jdff dff_B_s477KKrP8_2(.din(w_dff_B_Qlcq6qvH2_2),.dout(w_dff_B_s477KKrP8_2),.clk(gclk));
	jdff dff_B_qKTptbSZ1_2(.din(w_dff_B_s477KKrP8_2),.dout(w_dff_B_qKTptbSZ1_2),.clk(gclk));
	jdff dff_B_WlarPdLD0_2(.din(w_dff_B_qKTptbSZ1_2),.dout(w_dff_B_WlarPdLD0_2),.clk(gclk));
	jdff dff_B_45KLFwQS7_2(.din(w_dff_B_WlarPdLD0_2),.dout(w_dff_B_45KLFwQS7_2),.clk(gclk));
	jdff dff_B_TUyAwlTn3_2(.din(w_dff_B_45KLFwQS7_2),.dout(w_dff_B_TUyAwlTn3_2),.clk(gclk));
	jdff dff_B_b5ylFTOj4_2(.din(w_dff_B_TUyAwlTn3_2),.dout(w_dff_B_b5ylFTOj4_2),.clk(gclk));
	jdff dff_B_l91dVKwJ7_2(.din(w_dff_B_b5ylFTOj4_2),.dout(w_dff_B_l91dVKwJ7_2),.clk(gclk));
	jdff dff_B_96RTggfs1_2(.din(w_dff_B_l91dVKwJ7_2),.dout(w_dff_B_96RTggfs1_2),.clk(gclk));
	jdff dff_B_0qOC2W1v2_2(.din(w_dff_B_96RTggfs1_2),.dout(w_dff_B_0qOC2W1v2_2),.clk(gclk));
	jdff dff_B_NuO0l4nZ5_2(.din(w_dff_B_0qOC2W1v2_2),.dout(w_dff_B_NuO0l4nZ5_2),.clk(gclk));
	jdff dff_B_TBfQyYoT1_2(.din(w_dff_B_NuO0l4nZ5_2),.dout(w_dff_B_TBfQyYoT1_2),.clk(gclk));
	jdff dff_B_39pfXZz19_2(.din(w_dff_B_TBfQyYoT1_2),.dout(w_dff_B_39pfXZz19_2),.clk(gclk));
	jdff dff_B_8bu60b5c9_2(.din(w_dff_B_39pfXZz19_2),.dout(w_dff_B_8bu60b5c9_2),.clk(gclk));
	jdff dff_B_61PhXr827_2(.din(w_dff_B_8bu60b5c9_2),.dout(w_dff_B_61PhXr827_2),.clk(gclk));
	jdff dff_B_gQfjdZlo5_2(.din(n1283),.dout(w_dff_B_gQfjdZlo5_2),.clk(gclk));
	jdff dff_B_Gsa8nd0s8_1(.din(n1238),.dout(w_dff_B_Gsa8nd0s8_1),.clk(gclk));
	jdff dff_B_afuhBzha9_2(.din(n1146),.dout(w_dff_B_afuhBzha9_2),.clk(gclk));
	jdff dff_B_WtZzsr5W8_2(.din(w_dff_B_afuhBzha9_2),.dout(w_dff_B_WtZzsr5W8_2),.clk(gclk));
	jdff dff_B_Wwc8q2Rw4_2(.din(w_dff_B_WtZzsr5W8_2),.dout(w_dff_B_Wwc8q2Rw4_2),.clk(gclk));
	jdff dff_B_q5QB4lUo2_2(.din(w_dff_B_Wwc8q2Rw4_2),.dout(w_dff_B_q5QB4lUo2_2),.clk(gclk));
	jdff dff_B_swaUDdSF0_2(.din(w_dff_B_q5QB4lUo2_2),.dout(w_dff_B_swaUDdSF0_2),.clk(gclk));
	jdff dff_B_qDYt7nbd2_2(.din(w_dff_B_swaUDdSF0_2),.dout(w_dff_B_qDYt7nbd2_2),.clk(gclk));
	jdff dff_B_2qTqRvlW3_2(.din(w_dff_B_qDYt7nbd2_2),.dout(w_dff_B_2qTqRvlW3_2),.clk(gclk));
	jdff dff_B_vRuBQgIE4_2(.din(w_dff_B_2qTqRvlW3_2),.dout(w_dff_B_vRuBQgIE4_2),.clk(gclk));
	jdff dff_B_C6nCEh9i5_2(.din(w_dff_B_vRuBQgIE4_2),.dout(w_dff_B_C6nCEh9i5_2),.clk(gclk));
	jdff dff_B_pMm4pkmh7_2(.din(w_dff_B_C6nCEh9i5_2),.dout(w_dff_B_pMm4pkmh7_2),.clk(gclk));
	jdff dff_B_5I2ou4L92_2(.din(w_dff_B_pMm4pkmh7_2),.dout(w_dff_B_5I2ou4L92_2),.clk(gclk));
	jdff dff_B_dUH4GDyX4_2(.din(w_dff_B_5I2ou4L92_2),.dout(w_dff_B_dUH4GDyX4_2),.clk(gclk));
	jdff dff_B_kTw7f4GD7_2(.din(w_dff_B_dUH4GDyX4_2),.dout(w_dff_B_kTw7f4GD7_2),.clk(gclk));
	jdff dff_B_mdN2fhrM6_2(.din(w_dff_B_kTw7f4GD7_2),.dout(w_dff_B_mdN2fhrM6_2),.clk(gclk));
	jdff dff_B_mYzYfili8_2(.din(w_dff_B_mdN2fhrM6_2),.dout(w_dff_B_mYzYfili8_2),.clk(gclk));
	jdff dff_B_CfP76dGT1_2(.din(w_dff_B_mYzYfili8_2),.dout(w_dff_B_CfP76dGT1_2),.clk(gclk));
	jdff dff_B_EYDedzUd4_2(.din(w_dff_B_CfP76dGT1_2),.dout(w_dff_B_EYDedzUd4_2),.clk(gclk));
	jdff dff_B_PSKzpbiE1_2(.din(w_dff_B_EYDedzUd4_2),.dout(w_dff_B_PSKzpbiE1_2),.clk(gclk));
	jdff dff_B_z7sC5bZP5_2(.din(w_dff_B_PSKzpbiE1_2),.dout(w_dff_B_z7sC5bZP5_2),.clk(gclk));
	jdff dff_B_UEuPTdyw1_2(.din(w_dff_B_z7sC5bZP5_2),.dout(w_dff_B_UEuPTdyw1_2),.clk(gclk));
	jdff dff_B_fwIPDdqK3_2(.din(w_dff_B_UEuPTdyw1_2),.dout(w_dff_B_fwIPDdqK3_2),.clk(gclk));
	jdff dff_B_UnrrENxU3_2(.din(w_dff_B_fwIPDdqK3_2),.dout(w_dff_B_UnrrENxU3_2),.clk(gclk));
	jdff dff_B_wzpjEvUe5_2(.din(w_dff_B_UnrrENxU3_2),.dout(w_dff_B_wzpjEvUe5_2),.clk(gclk));
	jdff dff_B_SqVhbY4B1_2(.din(w_dff_B_wzpjEvUe5_2),.dout(w_dff_B_SqVhbY4B1_2),.clk(gclk));
	jdff dff_B_KhvejIkn0_2(.din(w_dff_B_SqVhbY4B1_2),.dout(w_dff_B_KhvejIkn0_2),.clk(gclk));
	jdff dff_B_rWSS7VCu7_2(.din(w_dff_B_KhvejIkn0_2),.dout(w_dff_B_rWSS7VCu7_2),.clk(gclk));
	jdff dff_B_RNsonPTE1_2(.din(w_dff_B_rWSS7VCu7_2),.dout(w_dff_B_RNsonPTE1_2),.clk(gclk));
	jdff dff_B_hs2zLa393_2(.din(w_dff_B_RNsonPTE1_2),.dout(w_dff_B_hs2zLa393_2),.clk(gclk));
	jdff dff_B_kzrcoXMJ4_2(.din(w_dff_B_hs2zLa393_2),.dout(w_dff_B_kzrcoXMJ4_2),.clk(gclk));
	jdff dff_B_agDZGcgb0_2(.din(n1192),.dout(w_dff_B_agDZGcgb0_2),.clk(gclk));
	jdff dff_B_KmONAJPs5_1(.din(n1147),.dout(w_dff_B_KmONAJPs5_1),.clk(gclk));
	jdff dff_B_9C3wDcnH7_2(.din(n1048),.dout(w_dff_B_9C3wDcnH7_2),.clk(gclk));
	jdff dff_B_aYjU6GZ77_2(.din(w_dff_B_9C3wDcnH7_2),.dout(w_dff_B_aYjU6GZ77_2),.clk(gclk));
	jdff dff_B_dAQ4DXwb0_2(.din(w_dff_B_aYjU6GZ77_2),.dout(w_dff_B_dAQ4DXwb0_2),.clk(gclk));
	jdff dff_B_GXnwgz5D6_2(.din(w_dff_B_dAQ4DXwb0_2),.dout(w_dff_B_GXnwgz5D6_2),.clk(gclk));
	jdff dff_B_wSezUTmB8_2(.din(w_dff_B_GXnwgz5D6_2),.dout(w_dff_B_wSezUTmB8_2),.clk(gclk));
	jdff dff_B_A9Q1NYPP4_2(.din(w_dff_B_wSezUTmB8_2),.dout(w_dff_B_A9Q1NYPP4_2),.clk(gclk));
	jdff dff_B_xn9GcnWh8_2(.din(w_dff_B_A9Q1NYPP4_2),.dout(w_dff_B_xn9GcnWh8_2),.clk(gclk));
	jdff dff_B_9j13FQdz2_2(.din(w_dff_B_xn9GcnWh8_2),.dout(w_dff_B_9j13FQdz2_2),.clk(gclk));
	jdff dff_B_7t34lPtK3_2(.din(w_dff_B_9j13FQdz2_2),.dout(w_dff_B_7t34lPtK3_2),.clk(gclk));
	jdff dff_B_Kagtc9w50_2(.din(w_dff_B_7t34lPtK3_2),.dout(w_dff_B_Kagtc9w50_2),.clk(gclk));
	jdff dff_B_H29SMceJ4_2(.din(w_dff_B_Kagtc9w50_2),.dout(w_dff_B_H29SMceJ4_2),.clk(gclk));
	jdff dff_B_QuDqRJX72_2(.din(w_dff_B_H29SMceJ4_2),.dout(w_dff_B_QuDqRJX72_2),.clk(gclk));
	jdff dff_B_FKa6rfTr3_2(.din(w_dff_B_QuDqRJX72_2),.dout(w_dff_B_FKa6rfTr3_2),.clk(gclk));
	jdff dff_B_gM8mhMaM2_2(.din(w_dff_B_FKa6rfTr3_2),.dout(w_dff_B_gM8mhMaM2_2),.clk(gclk));
	jdff dff_B_D6if3GDK8_2(.din(w_dff_B_gM8mhMaM2_2),.dout(w_dff_B_D6if3GDK8_2),.clk(gclk));
	jdff dff_B_k2LfXZY65_2(.din(w_dff_B_D6if3GDK8_2),.dout(w_dff_B_k2LfXZY65_2),.clk(gclk));
	jdff dff_B_ff1Wecaz5_2(.din(w_dff_B_k2LfXZY65_2),.dout(w_dff_B_ff1Wecaz5_2),.clk(gclk));
	jdff dff_B_BHTOasWb7_2(.din(w_dff_B_ff1Wecaz5_2),.dout(w_dff_B_BHTOasWb7_2),.clk(gclk));
	jdff dff_B_wdD4OTvt7_2(.din(w_dff_B_BHTOasWb7_2),.dout(w_dff_B_wdD4OTvt7_2),.clk(gclk));
	jdff dff_B_3AAbsJM04_2(.din(w_dff_B_wdD4OTvt7_2),.dout(w_dff_B_3AAbsJM04_2),.clk(gclk));
	jdff dff_B_IklaTZij1_2(.din(w_dff_B_3AAbsJM04_2),.dout(w_dff_B_IklaTZij1_2),.clk(gclk));
	jdff dff_B_wtlmhCxI6_2(.din(w_dff_B_IklaTZij1_2),.dout(w_dff_B_wtlmhCxI6_2),.clk(gclk));
	jdff dff_B_mwhgo5Sm6_2(.din(w_dff_B_wtlmhCxI6_2),.dout(w_dff_B_mwhgo5Sm6_2),.clk(gclk));
	jdff dff_B_0BakiQWU6_2(.din(w_dff_B_mwhgo5Sm6_2),.dout(w_dff_B_0BakiQWU6_2),.clk(gclk));
	jdff dff_B_QJHueJYm9_2(.din(w_dff_B_0BakiQWU6_2),.dout(w_dff_B_QJHueJYm9_2),.clk(gclk));
	jdff dff_B_bqaJiNvs7_2(.din(w_dff_B_QJHueJYm9_2),.dout(w_dff_B_bqaJiNvs7_2),.clk(gclk));
	jdff dff_B_X5KODBcQ8_2(.din(n1093),.dout(w_dff_B_X5KODBcQ8_2),.clk(gclk));
	jdff dff_B_Fm64XX5H4_1(.din(n1049),.dout(w_dff_B_Fm64XX5H4_1),.clk(gclk));
	jdff dff_B_oOHcAjoA9_2(.din(n949),.dout(w_dff_B_oOHcAjoA9_2),.clk(gclk));
	jdff dff_B_esaunbSb6_2(.din(w_dff_B_oOHcAjoA9_2),.dout(w_dff_B_esaunbSb6_2),.clk(gclk));
	jdff dff_B_UC16XmCD7_2(.din(w_dff_B_esaunbSb6_2),.dout(w_dff_B_UC16XmCD7_2),.clk(gclk));
	jdff dff_B_GPgHBzW92_2(.din(w_dff_B_UC16XmCD7_2),.dout(w_dff_B_GPgHBzW92_2),.clk(gclk));
	jdff dff_B_QC8QxRYn7_2(.din(w_dff_B_GPgHBzW92_2),.dout(w_dff_B_QC8QxRYn7_2),.clk(gclk));
	jdff dff_B_7PczbEzD1_2(.din(w_dff_B_QC8QxRYn7_2),.dout(w_dff_B_7PczbEzD1_2),.clk(gclk));
	jdff dff_B_KjjvChe66_2(.din(w_dff_B_7PczbEzD1_2),.dout(w_dff_B_KjjvChe66_2),.clk(gclk));
	jdff dff_B_qy9ut7mM2_2(.din(w_dff_B_KjjvChe66_2),.dout(w_dff_B_qy9ut7mM2_2),.clk(gclk));
	jdff dff_B_pVfqf9br4_2(.din(w_dff_B_qy9ut7mM2_2),.dout(w_dff_B_pVfqf9br4_2),.clk(gclk));
	jdff dff_B_Olcqf9OU1_2(.din(w_dff_B_pVfqf9br4_2),.dout(w_dff_B_Olcqf9OU1_2),.clk(gclk));
	jdff dff_B_wxZsCW0Z7_2(.din(w_dff_B_Olcqf9OU1_2),.dout(w_dff_B_wxZsCW0Z7_2),.clk(gclk));
	jdff dff_B_Tem6Ds3i6_2(.din(w_dff_B_wxZsCW0Z7_2),.dout(w_dff_B_Tem6Ds3i6_2),.clk(gclk));
	jdff dff_B_JpKp5glT1_2(.din(w_dff_B_Tem6Ds3i6_2),.dout(w_dff_B_JpKp5glT1_2),.clk(gclk));
	jdff dff_B_CXmYz1ss1_2(.din(w_dff_B_JpKp5glT1_2),.dout(w_dff_B_CXmYz1ss1_2),.clk(gclk));
	jdff dff_B_yOXM7FSi1_2(.din(w_dff_B_CXmYz1ss1_2),.dout(w_dff_B_yOXM7FSi1_2),.clk(gclk));
	jdff dff_B_fyk4inXr3_2(.din(w_dff_B_yOXM7FSi1_2),.dout(w_dff_B_fyk4inXr3_2),.clk(gclk));
	jdff dff_B_uUhqt12A2_2(.din(w_dff_B_fyk4inXr3_2),.dout(w_dff_B_uUhqt12A2_2),.clk(gclk));
	jdff dff_B_l6TdmEOG4_2(.din(w_dff_B_uUhqt12A2_2),.dout(w_dff_B_l6TdmEOG4_2),.clk(gclk));
	jdff dff_B_ipyvXdGK8_2(.din(w_dff_B_l6TdmEOG4_2),.dout(w_dff_B_ipyvXdGK8_2),.clk(gclk));
	jdff dff_B_FtuwAEjf2_2(.din(w_dff_B_ipyvXdGK8_2),.dout(w_dff_B_FtuwAEjf2_2),.clk(gclk));
	jdff dff_B_a9QQZFrk2_2(.din(w_dff_B_FtuwAEjf2_2),.dout(w_dff_B_a9QQZFrk2_2),.clk(gclk));
	jdff dff_B_3dB2SyH27_2(.din(w_dff_B_a9QQZFrk2_2),.dout(w_dff_B_3dB2SyH27_2),.clk(gclk));
	jdff dff_B_ezzIuTk95_2(.din(w_dff_B_3dB2SyH27_2),.dout(w_dff_B_ezzIuTk95_2),.clk(gclk));
	jdff dff_B_5zjqFYag2_2(.din(n994),.dout(w_dff_B_5zjqFYag2_2),.clk(gclk));
	jdff dff_B_8U4bRvfp3_1(.din(n950),.dout(w_dff_B_8U4bRvfp3_1),.clk(gclk));
	jdff dff_B_2KzRaxmx7_2(.din(n847),.dout(w_dff_B_2KzRaxmx7_2),.clk(gclk));
	jdff dff_B_9DUP62Jz3_2(.din(w_dff_B_2KzRaxmx7_2),.dout(w_dff_B_9DUP62Jz3_2),.clk(gclk));
	jdff dff_B_D9gNovTs7_2(.din(w_dff_B_9DUP62Jz3_2),.dout(w_dff_B_D9gNovTs7_2),.clk(gclk));
	jdff dff_B_OdEG0UGN2_2(.din(w_dff_B_D9gNovTs7_2),.dout(w_dff_B_OdEG0UGN2_2),.clk(gclk));
	jdff dff_B_XXCYUZkq1_2(.din(w_dff_B_OdEG0UGN2_2),.dout(w_dff_B_XXCYUZkq1_2),.clk(gclk));
	jdff dff_B_AiygU9vh8_2(.din(w_dff_B_XXCYUZkq1_2),.dout(w_dff_B_AiygU9vh8_2),.clk(gclk));
	jdff dff_B_dxEzX2fk8_2(.din(w_dff_B_AiygU9vh8_2),.dout(w_dff_B_dxEzX2fk8_2),.clk(gclk));
	jdff dff_B_fpa3Njoi2_2(.din(w_dff_B_dxEzX2fk8_2),.dout(w_dff_B_fpa3Njoi2_2),.clk(gclk));
	jdff dff_B_A3IYaeHX9_2(.din(w_dff_B_fpa3Njoi2_2),.dout(w_dff_B_A3IYaeHX9_2),.clk(gclk));
	jdff dff_B_AY4zyO7d9_2(.din(w_dff_B_A3IYaeHX9_2),.dout(w_dff_B_AY4zyO7d9_2),.clk(gclk));
	jdff dff_B_EjldRlN04_2(.din(w_dff_B_AY4zyO7d9_2),.dout(w_dff_B_EjldRlN04_2),.clk(gclk));
	jdff dff_B_O1AGV8Mj5_2(.din(w_dff_B_EjldRlN04_2),.dout(w_dff_B_O1AGV8Mj5_2),.clk(gclk));
	jdff dff_B_01r305D21_2(.din(w_dff_B_O1AGV8Mj5_2),.dout(w_dff_B_01r305D21_2),.clk(gclk));
	jdff dff_B_z4b6ezLd9_2(.din(w_dff_B_01r305D21_2),.dout(w_dff_B_z4b6ezLd9_2),.clk(gclk));
	jdff dff_B_O6uKpGyC9_2(.din(w_dff_B_z4b6ezLd9_2),.dout(w_dff_B_O6uKpGyC9_2),.clk(gclk));
	jdff dff_B_lJItwmgE8_2(.din(w_dff_B_O6uKpGyC9_2),.dout(w_dff_B_lJItwmgE8_2),.clk(gclk));
	jdff dff_B_mQKObdEv8_2(.din(w_dff_B_lJItwmgE8_2),.dout(w_dff_B_mQKObdEv8_2),.clk(gclk));
	jdff dff_B_s691kwsS4_2(.din(w_dff_B_mQKObdEv8_2),.dout(w_dff_B_s691kwsS4_2),.clk(gclk));
	jdff dff_B_ZaMaxq0z2_2(.din(w_dff_B_s691kwsS4_2),.dout(w_dff_B_ZaMaxq0z2_2),.clk(gclk));
	jdff dff_B_Az5yo4cW8_2(.din(w_dff_B_ZaMaxq0z2_2),.dout(w_dff_B_Az5yo4cW8_2),.clk(gclk));
	jdff dff_B_kPyJZvli6_2(.din(n888),.dout(w_dff_B_kPyJZvli6_2),.clk(gclk));
	jdff dff_B_GuYSHLCf0_1(.din(n848),.dout(w_dff_B_GuYSHLCf0_1),.clk(gclk));
	jdff dff_B_mUclxpru7_2(.din(n749),.dout(w_dff_B_mUclxpru7_2),.clk(gclk));
	jdff dff_B_UqD2P0ku7_2(.din(w_dff_B_mUclxpru7_2),.dout(w_dff_B_UqD2P0ku7_2),.clk(gclk));
	jdff dff_B_jYBafdmq0_2(.din(w_dff_B_UqD2P0ku7_2),.dout(w_dff_B_jYBafdmq0_2),.clk(gclk));
	jdff dff_B_Bqc89Xmn6_2(.din(w_dff_B_jYBafdmq0_2),.dout(w_dff_B_Bqc89Xmn6_2),.clk(gclk));
	jdff dff_B_velkgLsM1_2(.din(w_dff_B_Bqc89Xmn6_2),.dout(w_dff_B_velkgLsM1_2),.clk(gclk));
	jdff dff_B_RKygZ9z57_2(.din(w_dff_B_velkgLsM1_2),.dout(w_dff_B_RKygZ9z57_2),.clk(gclk));
	jdff dff_B_jRMC4n5K0_2(.din(w_dff_B_RKygZ9z57_2),.dout(w_dff_B_jRMC4n5K0_2),.clk(gclk));
	jdff dff_B_j4n2Vfjf3_2(.din(w_dff_B_jRMC4n5K0_2),.dout(w_dff_B_j4n2Vfjf3_2),.clk(gclk));
	jdff dff_B_KEqbxZAs4_2(.din(w_dff_B_j4n2Vfjf3_2),.dout(w_dff_B_KEqbxZAs4_2),.clk(gclk));
	jdff dff_B_ThCaaDeO8_2(.din(w_dff_B_KEqbxZAs4_2),.dout(w_dff_B_ThCaaDeO8_2),.clk(gclk));
	jdff dff_B_2mKLQ3yo5_2(.din(w_dff_B_ThCaaDeO8_2),.dout(w_dff_B_2mKLQ3yo5_2),.clk(gclk));
	jdff dff_B_vFPDQEYe6_2(.din(w_dff_B_2mKLQ3yo5_2),.dout(w_dff_B_vFPDQEYe6_2),.clk(gclk));
	jdff dff_B_wHyZ3VmD0_2(.din(w_dff_B_vFPDQEYe6_2),.dout(w_dff_B_wHyZ3VmD0_2),.clk(gclk));
	jdff dff_B_59OiT60s9_2(.din(w_dff_B_wHyZ3VmD0_2),.dout(w_dff_B_59OiT60s9_2),.clk(gclk));
	jdff dff_B_o5MepG8Q6_2(.din(w_dff_B_59OiT60s9_2),.dout(w_dff_B_o5MepG8Q6_2),.clk(gclk));
	jdff dff_B_fiHQYdtG8_2(.din(w_dff_B_o5MepG8Q6_2),.dout(w_dff_B_fiHQYdtG8_2),.clk(gclk));
	jdff dff_B_e8OA1mjm3_2(.din(w_dff_B_fiHQYdtG8_2),.dout(w_dff_B_e8OA1mjm3_2),.clk(gclk));
	jdff dff_B_1fONnGMT0_2(.din(n785),.dout(w_dff_B_1fONnGMT0_2),.clk(gclk));
	jdff dff_B_TyaiXiWX8_1(.din(n750),.dout(w_dff_B_TyaiXiWX8_1),.clk(gclk));
	jdff dff_B_kSAGYTcu8_2(.din(n657),.dout(w_dff_B_kSAGYTcu8_2),.clk(gclk));
	jdff dff_B_l915hsfN1_2(.din(w_dff_B_kSAGYTcu8_2),.dout(w_dff_B_l915hsfN1_2),.clk(gclk));
	jdff dff_B_7iAyFHPN8_2(.din(w_dff_B_l915hsfN1_2),.dout(w_dff_B_7iAyFHPN8_2),.clk(gclk));
	jdff dff_B_jVYgW8v39_2(.din(w_dff_B_7iAyFHPN8_2),.dout(w_dff_B_jVYgW8v39_2),.clk(gclk));
	jdff dff_B_PkLk4g3a4_2(.din(w_dff_B_jVYgW8v39_2),.dout(w_dff_B_PkLk4g3a4_2),.clk(gclk));
	jdff dff_B_r7RM0ham1_2(.din(w_dff_B_PkLk4g3a4_2),.dout(w_dff_B_r7RM0ham1_2),.clk(gclk));
	jdff dff_B_hW1pG5ih6_2(.din(w_dff_B_r7RM0ham1_2),.dout(w_dff_B_hW1pG5ih6_2),.clk(gclk));
	jdff dff_B_lK6Ho6Lu3_2(.din(w_dff_B_hW1pG5ih6_2),.dout(w_dff_B_lK6Ho6Lu3_2),.clk(gclk));
	jdff dff_B_69YT2YFB1_2(.din(w_dff_B_lK6Ho6Lu3_2),.dout(w_dff_B_69YT2YFB1_2),.clk(gclk));
	jdff dff_B_uJdAzTQq5_2(.din(w_dff_B_69YT2YFB1_2),.dout(w_dff_B_uJdAzTQq5_2),.clk(gclk));
	jdff dff_B_dwCyvl3u9_2(.din(w_dff_B_uJdAzTQq5_2),.dout(w_dff_B_dwCyvl3u9_2),.clk(gclk));
	jdff dff_B_puXUq43Z6_2(.din(w_dff_B_dwCyvl3u9_2),.dout(w_dff_B_puXUq43Z6_2),.clk(gclk));
	jdff dff_B_VdZ7G18k2_2(.din(w_dff_B_puXUq43Z6_2),.dout(w_dff_B_VdZ7G18k2_2),.clk(gclk));
	jdff dff_B_cutxkZDZ0_2(.din(w_dff_B_VdZ7G18k2_2),.dout(w_dff_B_cutxkZDZ0_2),.clk(gclk));
	jdff dff_B_1OLi2jHj4_2(.din(n686),.dout(w_dff_B_1OLi2jHj4_2),.clk(gclk));
	jdff dff_B_HLJpNWGj5_1(.din(n658),.dout(w_dff_B_HLJpNWGj5_1),.clk(gclk));
	jdff dff_B_mHi4H4Ha4_2(.din(n572),.dout(w_dff_B_mHi4H4Ha4_2),.clk(gclk));
	jdff dff_B_oaIatHEk3_2(.din(w_dff_B_mHi4H4Ha4_2),.dout(w_dff_B_oaIatHEk3_2),.clk(gclk));
	jdff dff_B_A3pP1mEA4_2(.din(w_dff_B_oaIatHEk3_2),.dout(w_dff_B_A3pP1mEA4_2),.clk(gclk));
	jdff dff_B_wb9IMQ4a4_2(.din(w_dff_B_A3pP1mEA4_2),.dout(w_dff_B_wb9IMQ4a4_2),.clk(gclk));
	jdff dff_B_7wzD5FRp2_2(.din(w_dff_B_wb9IMQ4a4_2),.dout(w_dff_B_7wzD5FRp2_2),.clk(gclk));
	jdff dff_B_e1HZEEES3_2(.din(w_dff_B_7wzD5FRp2_2),.dout(w_dff_B_e1HZEEES3_2),.clk(gclk));
	jdff dff_B_GK9OsL6K1_2(.din(w_dff_B_e1HZEEES3_2),.dout(w_dff_B_GK9OsL6K1_2),.clk(gclk));
	jdff dff_B_9NE4ZEbF7_2(.din(w_dff_B_GK9OsL6K1_2),.dout(w_dff_B_9NE4ZEbF7_2),.clk(gclk));
	jdff dff_B_RYKPiDi66_2(.din(w_dff_B_9NE4ZEbF7_2),.dout(w_dff_B_RYKPiDi66_2),.clk(gclk));
	jdff dff_B_NtiND1tn5_2(.din(w_dff_B_RYKPiDi66_2),.dout(w_dff_B_NtiND1tn5_2),.clk(gclk));
	jdff dff_B_CtZDk9d71_2(.din(w_dff_B_NtiND1tn5_2),.dout(w_dff_B_CtZDk9d71_2),.clk(gclk));
	jdff dff_B_uXYkKBb94_2(.din(n594),.dout(w_dff_B_uXYkKBb94_2),.clk(gclk));
	jdff dff_B_sfcCpwer7_1(.din(n573),.dout(w_dff_B_sfcCpwer7_1),.clk(gclk));
	jdff dff_B_cwChgFb36_2(.din(n494),.dout(w_dff_B_cwChgFb36_2),.clk(gclk));
	jdff dff_B_2jW0S4wf9_2(.din(w_dff_B_cwChgFb36_2),.dout(w_dff_B_2jW0S4wf9_2),.clk(gclk));
	jdff dff_B_4KFNpsED5_2(.din(w_dff_B_2jW0S4wf9_2),.dout(w_dff_B_4KFNpsED5_2),.clk(gclk));
	jdff dff_B_2THOlbMO2_2(.din(w_dff_B_4KFNpsED5_2),.dout(w_dff_B_2THOlbMO2_2),.clk(gclk));
	jdff dff_B_C8F8gtl95_2(.din(w_dff_B_2THOlbMO2_2),.dout(w_dff_B_C8F8gtl95_2),.clk(gclk));
	jdff dff_B_LMTNzjtw9_2(.din(w_dff_B_C8F8gtl95_2),.dout(w_dff_B_LMTNzjtw9_2),.clk(gclk));
	jdff dff_B_XpVCeBoh5_2(.din(w_dff_B_LMTNzjtw9_2),.dout(w_dff_B_XpVCeBoh5_2),.clk(gclk));
	jdff dff_B_JDMQXHZZ1_2(.din(w_dff_B_XpVCeBoh5_2),.dout(w_dff_B_JDMQXHZZ1_2),.clk(gclk));
	jdff dff_B_Q5RmVBP66_2(.din(n509),.dout(w_dff_B_Q5RmVBP66_2),.clk(gclk));
	jdff dff_B_jSyAlbkI4_2(.din(w_dff_B_Q5RmVBP66_2),.dout(w_dff_B_jSyAlbkI4_2),.clk(gclk));
	jdff dff_B_CHBlmuDm5_2(.din(w_dff_B_jSyAlbkI4_2),.dout(w_dff_B_CHBlmuDm5_2),.clk(gclk));
	jdff dff_B_3wmnwqtf4_1(.din(n495),.dout(w_dff_B_3wmnwqtf4_1),.clk(gclk));
	jdff dff_B_jCZ6uKDN9_1(.din(w_dff_B_3wmnwqtf4_1),.dout(w_dff_B_jCZ6uKDN9_1),.clk(gclk));
	jdff dff_B_vIMy7gBQ4_2(.din(n425),.dout(w_dff_B_vIMy7gBQ4_2),.clk(gclk));
	jdff dff_B_kJvLCQcI9_2(.din(w_dff_B_vIMy7gBQ4_2),.dout(w_dff_B_kJvLCQcI9_2),.clk(gclk));
	jdff dff_B_zDriRcux5_2(.din(w_dff_B_kJvLCQcI9_2),.dout(w_dff_B_zDriRcux5_2),.clk(gclk));
	jdff dff_B_pnrgftmm8_0(.din(n430),.dout(w_dff_B_pnrgftmm8_0),.clk(gclk));
	jdff dff_A_YpcDgDI45_0(.dout(w_n358_0[0]),.din(w_dff_A_YpcDgDI45_0),.clk(gclk));
	jdff dff_A_DeY9akHJ1_0(.dout(w_dff_A_YpcDgDI45_0),.din(w_dff_A_DeY9akHJ1_0),.clk(gclk));
	jdff dff_A_6dRNXfir4_1(.dout(w_n358_0[1]),.din(w_dff_A_6dRNXfir4_1),.clk(gclk));
	jdff dff_A_ae8Leg8q5_1(.dout(w_dff_A_6dRNXfir4_1),.din(w_dff_A_ae8Leg8q5_1),.clk(gclk));
	jdff dff_B_5UjToAl94_2(.din(n1651),.dout(w_dff_B_5UjToAl94_2),.clk(gclk));
	jdff dff_B_SP1HpvoC3_1(.din(n1649),.dout(w_dff_B_SP1HpvoC3_1),.clk(gclk));
	jdff dff_B_71cK37nZ6_2(.din(n1597),.dout(w_dff_B_71cK37nZ6_2),.clk(gclk));
	jdff dff_B_YK0SbFRt6_2(.din(w_dff_B_71cK37nZ6_2),.dout(w_dff_B_YK0SbFRt6_2),.clk(gclk));
	jdff dff_B_l9SbmwhF0_2(.din(w_dff_B_YK0SbFRt6_2),.dout(w_dff_B_l9SbmwhF0_2),.clk(gclk));
	jdff dff_B_jRxX2vNX1_2(.din(w_dff_B_l9SbmwhF0_2),.dout(w_dff_B_jRxX2vNX1_2),.clk(gclk));
	jdff dff_B_TXHHwfc74_2(.din(w_dff_B_jRxX2vNX1_2),.dout(w_dff_B_TXHHwfc74_2),.clk(gclk));
	jdff dff_B_VPUXu7tS8_2(.din(w_dff_B_TXHHwfc74_2),.dout(w_dff_B_VPUXu7tS8_2),.clk(gclk));
	jdff dff_B_P3CeeXQm7_2(.din(w_dff_B_VPUXu7tS8_2),.dout(w_dff_B_P3CeeXQm7_2),.clk(gclk));
	jdff dff_B_o9V35KRA9_2(.din(w_dff_B_P3CeeXQm7_2),.dout(w_dff_B_o9V35KRA9_2),.clk(gclk));
	jdff dff_B_nh9s3tTn1_2(.din(w_dff_B_o9V35KRA9_2),.dout(w_dff_B_nh9s3tTn1_2),.clk(gclk));
	jdff dff_B_vSbYCo453_2(.din(w_dff_B_nh9s3tTn1_2),.dout(w_dff_B_vSbYCo453_2),.clk(gclk));
	jdff dff_B_e9QocAal7_2(.din(w_dff_B_vSbYCo453_2),.dout(w_dff_B_e9QocAal7_2),.clk(gclk));
	jdff dff_B_wgWsdMIV8_2(.din(w_dff_B_e9QocAal7_2),.dout(w_dff_B_wgWsdMIV8_2),.clk(gclk));
	jdff dff_B_DAbkcINL6_2(.din(w_dff_B_wgWsdMIV8_2),.dout(w_dff_B_DAbkcINL6_2),.clk(gclk));
	jdff dff_B_8x9jV9B98_2(.din(w_dff_B_DAbkcINL6_2),.dout(w_dff_B_8x9jV9B98_2),.clk(gclk));
	jdff dff_B_G5xoHGjX5_2(.din(w_dff_B_8x9jV9B98_2),.dout(w_dff_B_G5xoHGjX5_2),.clk(gclk));
	jdff dff_B_mjikOwLC7_2(.din(w_dff_B_G5xoHGjX5_2),.dout(w_dff_B_mjikOwLC7_2),.clk(gclk));
	jdff dff_B_u8zQrG3z9_2(.din(w_dff_B_mjikOwLC7_2),.dout(w_dff_B_u8zQrG3z9_2),.clk(gclk));
	jdff dff_B_ZggIJJAC3_2(.din(w_dff_B_u8zQrG3z9_2),.dout(w_dff_B_ZggIJJAC3_2),.clk(gclk));
	jdff dff_B_WvfaBn5O1_2(.din(w_dff_B_ZggIJJAC3_2),.dout(w_dff_B_WvfaBn5O1_2),.clk(gclk));
	jdff dff_B_zqQtchwe3_2(.din(w_dff_B_WvfaBn5O1_2),.dout(w_dff_B_zqQtchwe3_2),.clk(gclk));
	jdff dff_B_IXOXLDQa0_2(.din(w_dff_B_zqQtchwe3_2),.dout(w_dff_B_IXOXLDQa0_2),.clk(gclk));
	jdff dff_B_R41Ituzw7_2(.din(w_dff_B_IXOXLDQa0_2),.dout(w_dff_B_R41Ituzw7_2),.clk(gclk));
	jdff dff_B_e92hMknu6_2(.din(w_dff_B_R41Ituzw7_2),.dout(w_dff_B_e92hMknu6_2),.clk(gclk));
	jdff dff_B_0ZkeI9lZ3_2(.din(w_dff_B_e92hMknu6_2),.dout(w_dff_B_0ZkeI9lZ3_2),.clk(gclk));
	jdff dff_B_tuLgRq3u5_2(.din(w_dff_B_0ZkeI9lZ3_2),.dout(w_dff_B_tuLgRq3u5_2),.clk(gclk));
	jdff dff_B_EM5gG7WT6_2(.din(w_dff_B_tuLgRq3u5_2),.dout(w_dff_B_EM5gG7WT6_2),.clk(gclk));
	jdff dff_B_2bCPBpfY4_2(.din(w_dff_B_EM5gG7WT6_2),.dout(w_dff_B_2bCPBpfY4_2),.clk(gclk));
	jdff dff_B_rFemxtgI9_2(.din(w_dff_B_2bCPBpfY4_2),.dout(w_dff_B_rFemxtgI9_2),.clk(gclk));
	jdff dff_B_TE82Mu566_2(.din(w_dff_B_rFemxtgI9_2),.dout(w_dff_B_TE82Mu566_2),.clk(gclk));
	jdff dff_B_YNoogsYC9_2(.din(w_dff_B_TE82Mu566_2),.dout(w_dff_B_YNoogsYC9_2),.clk(gclk));
	jdff dff_B_DEJEUtwu3_2(.din(w_dff_B_YNoogsYC9_2),.dout(w_dff_B_DEJEUtwu3_2),.clk(gclk));
	jdff dff_B_Qnw7XuIt0_2(.din(w_dff_B_DEJEUtwu3_2),.dout(w_dff_B_Qnw7XuIt0_2),.clk(gclk));
	jdff dff_B_Djj2TcPL3_2(.din(w_dff_B_Qnw7XuIt0_2),.dout(w_dff_B_Djj2TcPL3_2),.clk(gclk));
	jdff dff_B_bKHsVbBg8_2(.din(w_dff_B_Djj2TcPL3_2),.dout(w_dff_B_bKHsVbBg8_2),.clk(gclk));
	jdff dff_B_NV0MGv9q6_2(.din(w_dff_B_bKHsVbBg8_2),.dout(w_dff_B_NV0MGv9q6_2),.clk(gclk));
	jdff dff_B_kDOhS67u4_2(.din(w_dff_B_NV0MGv9q6_2),.dout(w_dff_B_kDOhS67u4_2),.clk(gclk));
	jdff dff_B_TLj0vM5f8_2(.din(w_dff_B_kDOhS67u4_2),.dout(w_dff_B_TLj0vM5f8_2),.clk(gclk));
	jdff dff_B_dWYwdqNx2_2(.din(w_dff_B_TLj0vM5f8_2),.dout(w_dff_B_dWYwdqNx2_2),.clk(gclk));
	jdff dff_B_lljg9htH9_2(.din(w_dff_B_dWYwdqNx2_2),.dout(w_dff_B_lljg9htH9_2),.clk(gclk));
	jdff dff_B_few84Wq91_2(.din(w_dff_B_lljg9htH9_2),.dout(w_dff_B_few84Wq91_2),.clk(gclk));
	jdff dff_B_0eo0p8Kg9_2(.din(w_dff_B_few84Wq91_2),.dout(w_dff_B_0eo0p8Kg9_2),.clk(gclk));
	jdff dff_B_MI4lqtHn0_2(.din(w_dff_B_0eo0p8Kg9_2),.dout(w_dff_B_MI4lqtHn0_2),.clk(gclk));
	jdff dff_B_ykau3p4K6_2(.din(w_dff_B_MI4lqtHn0_2),.dout(w_dff_B_ykau3p4K6_2),.clk(gclk));
	jdff dff_B_Mk0TUSzN9_2(.din(w_dff_B_ykau3p4K6_2),.dout(w_dff_B_Mk0TUSzN9_2),.clk(gclk));
	jdff dff_B_zOpO2JFm7_2(.din(w_dff_B_Mk0TUSzN9_2),.dout(w_dff_B_zOpO2JFm7_2),.clk(gclk));
	jdff dff_B_sg5RzDjZ8_2(.din(w_dff_B_zOpO2JFm7_2),.dout(w_dff_B_sg5RzDjZ8_2),.clk(gclk));
	jdff dff_B_ZnchbZUI3_1(.din(n1598),.dout(w_dff_B_ZnchbZUI3_1),.clk(gclk));
	jdff dff_B_wdAMPoaF0_2(.din(n1540),.dout(w_dff_B_wdAMPoaF0_2),.clk(gclk));
	jdff dff_B_5URAdbae0_2(.din(w_dff_B_wdAMPoaF0_2),.dout(w_dff_B_5URAdbae0_2),.clk(gclk));
	jdff dff_B_2wvz0KpW4_2(.din(w_dff_B_5URAdbae0_2),.dout(w_dff_B_2wvz0KpW4_2),.clk(gclk));
	jdff dff_B_BClbjmIh3_2(.din(w_dff_B_2wvz0KpW4_2),.dout(w_dff_B_BClbjmIh3_2),.clk(gclk));
	jdff dff_B_3RZ21tG67_2(.din(w_dff_B_BClbjmIh3_2),.dout(w_dff_B_3RZ21tG67_2),.clk(gclk));
	jdff dff_B_wRwX9GTn0_2(.din(w_dff_B_3RZ21tG67_2),.dout(w_dff_B_wRwX9GTn0_2),.clk(gclk));
	jdff dff_B_CeA2Fwuc8_2(.din(w_dff_B_wRwX9GTn0_2),.dout(w_dff_B_CeA2Fwuc8_2),.clk(gclk));
	jdff dff_B_wQ4XOuxH8_2(.din(w_dff_B_CeA2Fwuc8_2),.dout(w_dff_B_wQ4XOuxH8_2),.clk(gclk));
	jdff dff_B_MgCTk6jI1_2(.din(w_dff_B_wQ4XOuxH8_2),.dout(w_dff_B_MgCTk6jI1_2),.clk(gclk));
	jdff dff_B_w5cP2fYv4_2(.din(w_dff_B_MgCTk6jI1_2),.dout(w_dff_B_w5cP2fYv4_2),.clk(gclk));
	jdff dff_B_UDIBngJ91_2(.din(w_dff_B_w5cP2fYv4_2),.dout(w_dff_B_UDIBngJ91_2),.clk(gclk));
	jdff dff_B_bqyMLTma7_2(.din(w_dff_B_UDIBngJ91_2),.dout(w_dff_B_bqyMLTma7_2),.clk(gclk));
	jdff dff_B_AdknMspm5_2(.din(w_dff_B_bqyMLTma7_2),.dout(w_dff_B_AdknMspm5_2),.clk(gclk));
	jdff dff_B_1tY35QHh3_2(.din(w_dff_B_AdknMspm5_2),.dout(w_dff_B_1tY35QHh3_2),.clk(gclk));
	jdff dff_B_oxchOEEt4_2(.din(w_dff_B_1tY35QHh3_2),.dout(w_dff_B_oxchOEEt4_2),.clk(gclk));
	jdff dff_B_64Cmum3t4_2(.din(w_dff_B_oxchOEEt4_2),.dout(w_dff_B_64Cmum3t4_2),.clk(gclk));
	jdff dff_B_fzBkggOH7_2(.din(w_dff_B_64Cmum3t4_2),.dout(w_dff_B_fzBkggOH7_2),.clk(gclk));
	jdff dff_B_aHIko8rw1_2(.din(w_dff_B_fzBkggOH7_2),.dout(w_dff_B_aHIko8rw1_2),.clk(gclk));
	jdff dff_B_cSpqfCL07_2(.din(w_dff_B_aHIko8rw1_2),.dout(w_dff_B_cSpqfCL07_2),.clk(gclk));
	jdff dff_B_Kd4jgXSm8_2(.din(w_dff_B_cSpqfCL07_2),.dout(w_dff_B_Kd4jgXSm8_2),.clk(gclk));
	jdff dff_B_moHWxap25_2(.din(w_dff_B_Kd4jgXSm8_2),.dout(w_dff_B_moHWxap25_2),.clk(gclk));
	jdff dff_B_RRltPjFi3_2(.din(w_dff_B_moHWxap25_2),.dout(w_dff_B_RRltPjFi3_2),.clk(gclk));
	jdff dff_B_5wKUrzf65_2(.din(w_dff_B_RRltPjFi3_2),.dout(w_dff_B_5wKUrzf65_2),.clk(gclk));
	jdff dff_B_dGSAcWoX4_2(.din(w_dff_B_5wKUrzf65_2),.dout(w_dff_B_dGSAcWoX4_2),.clk(gclk));
	jdff dff_B_jsmUPEP30_2(.din(w_dff_B_dGSAcWoX4_2),.dout(w_dff_B_jsmUPEP30_2),.clk(gclk));
	jdff dff_B_fv9hfoGt9_2(.din(w_dff_B_jsmUPEP30_2),.dout(w_dff_B_fv9hfoGt9_2),.clk(gclk));
	jdff dff_B_5FZSmRek4_2(.din(w_dff_B_fv9hfoGt9_2),.dout(w_dff_B_5FZSmRek4_2),.clk(gclk));
	jdff dff_B_mjx9Eo4e7_2(.din(w_dff_B_5FZSmRek4_2),.dout(w_dff_B_mjx9Eo4e7_2),.clk(gclk));
	jdff dff_B_rUwZoaS78_2(.din(w_dff_B_mjx9Eo4e7_2),.dout(w_dff_B_rUwZoaS78_2),.clk(gclk));
	jdff dff_B_D0lFcWPB5_2(.din(w_dff_B_rUwZoaS78_2),.dout(w_dff_B_D0lFcWPB5_2),.clk(gclk));
	jdff dff_B_NjQMJKnR7_2(.din(w_dff_B_D0lFcWPB5_2),.dout(w_dff_B_NjQMJKnR7_2),.clk(gclk));
	jdff dff_B_X9DVy4Qx8_2(.din(w_dff_B_NjQMJKnR7_2),.dout(w_dff_B_X9DVy4Qx8_2),.clk(gclk));
	jdff dff_B_0XLoYU5T4_2(.din(w_dff_B_X9DVy4Qx8_2),.dout(w_dff_B_0XLoYU5T4_2),.clk(gclk));
	jdff dff_B_Vp3ifSjy0_2(.din(w_dff_B_0XLoYU5T4_2),.dout(w_dff_B_Vp3ifSjy0_2),.clk(gclk));
	jdff dff_B_okLpPXzQ2_2(.din(w_dff_B_Vp3ifSjy0_2),.dout(w_dff_B_okLpPXzQ2_2),.clk(gclk));
	jdff dff_B_xCEpiB3p3_2(.din(w_dff_B_okLpPXzQ2_2),.dout(w_dff_B_xCEpiB3p3_2),.clk(gclk));
	jdff dff_B_hH3DvJTQ0_2(.din(w_dff_B_xCEpiB3p3_2),.dout(w_dff_B_hH3DvJTQ0_2),.clk(gclk));
	jdff dff_B_umnE4FMY2_2(.din(w_dff_B_hH3DvJTQ0_2),.dout(w_dff_B_umnE4FMY2_2),.clk(gclk));
	jdff dff_B_dmCv4WHx8_2(.din(w_dff_B_umnE4FMY2_2),.dout(w_dff_B_dmCv4WHx8_2),.clk(gclk));
	jdff dff_B_45YYGLI79_2(.din(w_dff_B_dmCv4WHx8_2),.dout(w_dff_B_45YYGLI79_2),.clk(gclk));
	jdff dff_B_qf6KaGu87_2(.din(w_dff_B_45YYGLI79_2),.dout(w_dff_B_qf6KaGu87_2),.clk(gclk));
	jdff dff_B_f5jzpFwY9_2(.din(n1579),.dout(w_dff_B_f5jzpFwY9_2),.clk(gclk));
	jdff dff_B_CrfapjXi1_1(.din(n1541),.dout(w_dff_B_CrfapjXi1_1),.clk(gclk));
	jdff dff_B_V69YQsqG4_2(.din(n1476),.dout(w_dff_B_V69YQsqG4_2),.clk(gclk));
	jdff dff_B_6UawjIrV5_2(.din(w_dff_B_V69YQsqG4_2),.dout(w_dff_B_6UawjIrV5_2),.clk(gclk));
	jdff dff_B_EDDUXb4S1_2(.din(w_dff_B_6UawjIrV5_2),.dout(w_dff_B_EDDUXb4S1_2),.clk(gclk));
	jdff dff_B_ud80M0vy1_2(.din(w_dff_B_EDDUXb4S1_2),.dout(w_dff_B_ud80M0vy1_2),.clk(gclk));
	jdff dff_B_mXgA2FpI4_2(.din(w_dff_B_ud80M0vy1_2),.dout(w_dff_B_mXgA2FpI4_2),.clk(gclk));
	jdff dff_B_09ygmIav2_2(.din(w_dff_B_mXgA2FpI4_2),.dout(w_dff_B_09ygmIav2_2),.clk(gclk));
	jdff dff_B_Auv3TVh96_2(.din(w_dff_B_09ygmIav2_2),.dout(w_dff_B_Auv3TVh96_2),.clk(gclk));
	jdff dff_B_Xi8lea3v9_2(.din(w_dff_B_Auv3TVh96_2),.dout(w_dff_B_Xi8lea3v9_2),.clk(gclk));
	jdff dff_B_BGrSYvj22_2(.din(w_dff_B_Xi8lea3v9_2),.dout(w_dff_B_BGrSYvj22_2),.clk(gclk));
	jdff dff_B_F8gJViX73_2(.din(w_dff_B_BGrSYvj22_2),.dout(w_dff_B_F8gJViX73_2),.clk(gclk));
	jdff dff_B_dMF2Ni9S0_2(.din(w_dff_B_F8gJViX73_2),.dout(w_dff_B_dMF2Ni9S0_2),.clk(gclk));
	jdff dff_B_2HGrpTvm3_2(.din(w_dff_B_dMF2Ni9S0_2),.dout(w_dff_B_2HGrpTvm3_2),.clk(gclk));
	jdff dff_B_Z94lnMzP8_2(.din(w_dff_B_2HGrpTvm3_2),.dout(w_dff_B_Z94lnMzP8_2),.clk(gclk));
	jdff dff_B_CGHP00si3_2(.din(w_dff_B_Z94lnMzP8_2),.dout(w_dff_B_CGHP00si3_2),.clk(gclk));
	jdff dff_B_4raPXYEk1_2(.din(w_dff_B_CGHP00si3_2),.dout(w_dff_B_4raPXYEk1_2),.clk(gclk));
	jdff dff_B_RJ5hshh29_2(.din(w_dff_B_4raPXYEk1_2),.dout(w_dff_B_RJ5hshh29_2),.clk(gclk));
	jdff dff_B_vtNaouEg7_2(.din(w_dff_B_RJ5hshh29_2),.dout(w_dff_B_vtNaouEg7_2),.clk(gclk));
	jdff dff_B_28g9tOFh2_2(.din(w_dff_B_vtNaouEg7_2),.dout(w_dff_B_28g9tOFh2_2),.clk(gclk));
	jdff dff_B_FKJ3wFMO7_2(.din(w_dff_B_28g9tOFh2_2),.dout(w_dff_B_FKJ3wFMO7_2),.clk(gclk));
	jdff dff_B_prSK7DWw7_2(.din(w_dff_B_FKJ3wFMO7_2),.dout(w_dff_B_prSK7DWw7_2),.clk(gclk));
	jdff dff_B_BCAdCdye2_2(.din(w_dff_B_prSK7DWw7_2),.dout(w_dff_B_BCAdCdye2_2),.clk(gclk));
	jdff dff_B_Q8ulPfxt9_2(.din(w_dff_B_BCAdCdye2_2),.dout(w_dff_B_Q8ulPfxt9_2),.clk(gclk));
	jdff dff_B_bHpKbI9B6_2(.din(w_dff_B_Q8ulPfxt9_2),.dout(w_dff_B_bHpKbI9B6_2),.clk(gclk));
	jdff dff_B_K5ju37lr5_2(.din(w_dff_B_bHpKbI9B6_2),.dout(w_dff_B_K5ju37lr5_2),.clk(gclk));
	jdff dff_B_229QCfxt9_2(.din(w_dff_B_K5ju37lr5_2),.dout(w_dff_B_229QCfxt9_2),.clk(gclk));
	jdff dff_B_7v78ovQT2_2(.din(w_dff_B_229QCfxt9_2),.dout(w_dff_B_7v78ovQT2_2),.clk(gclk));
	jdff dff_B_JsVFV5wz2_2(.din(w_dff_B_7v78ovQT2_2),.dout(w_dff_B_JsVFV5wz2_2),.clk(gclk));
	jdff dff_B_SdNBurqI6_2(.din(w_dff_B_JsVFV5wz2_2),.dout(w_dff_B_SdNBurqI6_2),.clk(gclk));
	jdff dff_B_pODrh9r59_2(.din(w_dff_B_SdNBurqI6_2),.dout(w_dff_B_pODrh9r59_2),.clk(gclk));
	jdff dff_B_7zxmP5Zr7_2(.din(w_dff_B_pODrh9r59_2),.dout(w_dff_B_7zxmP5Zr7_2),.clk(gclk));
	jdff dff_B_x2Z4l0kg9_2(.din(w_dff_B_7zxmP5Zr7_2),.dout(w_dff_B_x2Z4l0kg9_2),.clk(gclk));
	jdff dff_B_jLFTsBHk6_2(.din(w_dff_B_x2Z4l0kg9_2),.dout(w_dff_B_jLFTsBHk6_2),.clk(gclk));
	jdff dff_B_9D1WOhjy7_2(.din(w_dff_B_jLFTsBHk6_2),.dout(w_dff_B_9D1WOhjy7_2),.clk(gclk));
	jdff dff_B_WFLJ8JVs3_2(.din(w_dff_B_9D1WOhjy7_2),.dout(w_dff_B_WFLJ8JVs3_2),.clk(gclk));
	jdff dff_B_z7olk5Sa9_2(.din(w_dff_B_WFLJ8JVs3_2),.dout(w_dff_B_z7olk5Sa9_2),.clk(gclk));
	jdff dff_B_pGQqjV7U0_2(.din(w_dff_B_z7olk5Sa9_2),.dout(w_dff_B_pGQqjV7U0_2),.clk(gclk));
	jdff dff_B_0hNEUiv10_2(.din(w_dff_B_pGQqjV7U0_2),.dout(w_dff_B_0hNEUiv10_2),.clk(gclk));
	jdff dff_B_ooaUOpmP9_2(.din(w_dff_B_0hNEUiv10_2),.dout(w_dff_B_ooaUOpmP9_2),.clk(gclk));
	jdff dff_B_y0v4w9nr6_2(.din(n1515),.dout(w_dff_B_y0v4w9nr6_2),.clk(gclk));
	jdff dff_B_m02Mw1jm9_1(.din(n1477),.dout(w_dff_B_m02Mw1jm9_1),.clk(gclk));
	jdff dff_B_cxFXrJTS5_2(.din(n1405),.dout(w_dff_B_cxFXrJTS5_2),.clk(gclk));
	jdff dff_B_kqS5ULAi3_2(.din(w_dff_B_cxFXrJTS5_2),.dout(w_dff_B_kqS5ULAi3_2),.clk(gclk));
	jdff dff_B_2yRIJCt79_2(.din(w_dff_B_kqS5ULAi3_2),.dout(w_dff_B_2yRIJCt79_2),.clk(gclk));
	jdff dff_B_2zxAJRTr3_2(.din(w_dff_B_2yRIJCt79_2),.dout(w_dff_B_2zxAJRTr3_2),.clk(gclk));
	jdff dff_B_WwHnwgwd0_2(.din(w_dff_B_2zxAJRTr3_2),.dout(w_dff_B_WwHnwgwd0_2),.clk(gclk));
	jdff dff_B_SuE322iB6_2(.din(w_dff_B_WwHnwgwd0_2),.dout(w_dff_B_SuE322iB6_2),.clk(gclk));
	jdff dff_B_9dmu7QGB2_2(.din(w_dff_B_SuE322iB6_2),.dout(w_dff_B_9dmu7QGB2_2),.clk(gclk));
	jdff dff_B_mLpTjJZh3_2(.din(w_dff_B_9dmu7QGB2_2),.dout(w_dff_B_mLpTjJZh3_2),.clk(gclk));
	jdff dff_B_w0Tf9ODh6_2(.din(w_dff_B_mLpTjJZh3_2),.dout(w_dff_B_w0Tf9ODh6_2),.clk(gclk));
	jdff dff_B_UFDaTRqW1_2(.din(w_dff_B_w0Tf9ODh6_2),.dout(w_dff_B_UFDaTRqW1_2),.clk(gclk));
	jdff dff_B_UYGEtdvl5_2(.din(w_dff_B_UFDaTRqW1_2),.dout(w_dff_B_UYGEtdvl5_2),.clk(gclk));
	jdff dff_B_x2XSTL6S0_2(.din(w_dff_B_UYGEtdvl5_2),.dout(w_dff_B_x2XSTL6S0_2),.clk(gclk));
	jdff dff_B_QiZuaDGp4_2(.din(w_dff_B_x2XSTL6S0_2),.dout(w_dff_B_QiZuaDGp4_2),.clk(gclk));
	jdff dff_B_3UsTOzIP5_2(.din(w_dff_B_QiZuaDGp4_2),.dout(w_dff_B_3UsTOzIP5_2),.clk(gclk));
	jdff dff_B_5P9KJta54_2(.din(w_dff_B_3UsTOzIP5_2),.dout(w_dff_B_5P9KJta54_2),.clk(gclk));
	jdff dff_B_v9sYggrd1_2(.din(w_dff_B_5P9KJta54_2),.dout(w_dff_B_v9sYggrd1_2),.clk(gclk));
	jdff dff_B_Ssl33oJn0_2(.din(w_dff_B_v9sYggrd1_2),.dout(w_dff_B_Ssl33oJn0_2),.clk(gclk));
	jdff dff_B_U1WXKmK53_2(.din(w_dff_B_Ssl33oJn0_2),.dout(w_dff_B_U1WXKmK53_2),.clk(gclk));
	jdff dff_B_wuZPX3pd1_2(.din(w_dff_B_U1WXKmK53_2),.dout(w_dff_B_wuZPX3pd1_2),.clk(gclk));
	jdff dff_B_HGWXxLhB5_2(.din(w_dff_B_wuZPX3pd1_2),.dout(w_dff_B_HGWXxLhB5_2),.clk(gclk));
	jdff dff_B_paDfDDmw0_2(.din(w_dff_B_HGWXxLhB5_2),.dout(w_dff_B_paDfDDmw0_2),.clk(gclk));
	jdff dff_B_6GFn8D1V1_2(.din(w_dff_B_paDfDDmw0_2),.dout(w_dff_B_6GFn8D1V1_2),.clk(gclk));
	jdff dff_B_tL76Uq5V2_2(.din(w_dff_B_6GFn8D1V1_2),.dout(w_dff_B_tL76Uq5V2_2),.clk(gclk));
	jdff dff_B_cGjkux6G4_2(.din(w_dff_B_tL76Uq5V2_2),.dout(w_dff_B_cGjkux6G4_2),.clk(gclk));
	jdff dff_B_mi4VUHIQ2_2(.din(w_dff_B_cGjkux6G4_2),.dout(w_dff_B_mi4VUHIQ2_2),.clk(gclk));
	jdff dff_B_ZMfxlqyd3_2(.din(w_dff_B_mi4VUHIQ2_2),.dout(w_dff_B_ZMfxlqyd3_2),.clk(gclk));
	jdff dff_B_iYhExfym0_2(.din(w_dff_B_ZMfxlqyd3_2),.dout(w_dff_B_iYhExfym0_2),.clk(gclk));
	jdff dff_B_wiwxmdGk2_2(.din(w_dff_B_iYhExfym0_2),.dout(w_dff_B_wiwxmdGk2_2),.clk(gclk));
	jdff dff_B_2WCuw5mT3_2(.din(w_dff_B_wiwxmdGk2_2),.dout(w_dff_B_2WCuw5mT3_2),.clk(gclk));
	jdff dff_B_Tb1vvtYi2_2(.din(w_dff_B_2WCuw5mT3_2),.dout(w_dff_B_Tb1vvtYi2_2),.clk(gclk));
	jdff dff_B_Ixm0xFCO7_2(.din(w_dff_B_Tb1vvtYi2_2),.dout(w_dff_B_Ixm0xFCO7_2),.clk(gclk));
	jdff dff_B_GR8kSYNR7_2(.din(w_dff_B_Ixm0xFCO7_2),.dout(w_dff_B_GR8kSYNR7_2),.clk(gclk));
	jdff dff_B_5Vy1W1Gf9_2(.din(w_dff_B_GR8kSYNR7_2),.dout(w_dff_B_5Vy1W1Gf9_2),.clk(gclk));
	jdff dff_B_6uS1MzVD9_2(.din(w_dff_B_5Vy1W1Gf9_2),.dout(w_dff_B_6uS1MzVD9_2),.clk(gclk));
	jdff dff_B_FlcmKFLv6_2(.din(w_dff_B_6uS1MzVD9_2),.dout(w_dff_B_FlcmKFLv6_2),.clk(gclk));
	jdff dff_B_9zXT8tMX6_2(.din(n1444),.dout(w_dff_B_9zXT8tMX6_2),.clk(gclk));
	jdff dff_B_g8XKJVFw3_1(.din(n1406),.dout(w_dff_B_g8XKJVFw3_1),.clk(gclk));
	jdff dff_B_79xcPeQN5_2(.din(n1327),.dout(w_dff_B_79xcPeQN5_2),.clk(gclk));
	jdff dff_B_NVgzO3NF1_2(.din(w_dff_B_79xcPeQN5_2),.dout(w_dff_B_NVgzO3NF1_2),.clk(gclk));
	jdff dff_B_XFdAogwm4_2(.din(w_dff_B_NVgzO3NF1_2),.dout(w_dff_B_XFdAogwm4_2),.clk(gclk));
	jdff dff_B_FtAlXc7k3_2(.din(w_dff_B_XFdAogwm4_2),.dout(w_dff_B_FtAlXc7k3_2),.clk(gclk));
	jdff dff_B_3wdPJEmg0_2(.din(w_dff_B_FtAlXc7k3_2),.dout(w_dff_B_3wdPJEmg0_2),.clk(gclk));
	jdff dff_B_dcIfVtK90_2(.din(w_dff_B_3wdPJEmg0_2),.dout(w_dff_B_dcIfVtK90_2),.clk(gclk));
	jdff dff_B_Zuw9jU3M8_2(.din(w_dff_B_dcIfVtK90_2),.dout(w_dff_B_Zuw9jU3M8_2),.clk(gclk));
	jdff dff_B_AmqrlRJz0_2(.din(w_dff_B_Zuw9jU3M8_2),.dout(w_dff_B_AmqrlRJz0_2),.clk(gclk));
	jdff dff_B_3ZkWtzQX2_2(.din(w_dff_B_AmqrlRJz0_2),.dout(w_dff_B_3ZkWtzQX2_2),.clk(gclk));
	jdff dff_B_Kx9IwpM71_2(.din(w_dff_B_3ZkWtzQX2_2),.dout(w_dff_B_Kx9IwpM71_2),.clk(gclk));
	jdff dff_B_HUmgC5bV4_2(.din(w_dff_B_Kx9IwpM71_2),.dout(w_dff_B_HUmgC5bV4_2),.clk(gclk));
	jdff dff_B_8zupik028_2(.din(w_dff_B_HUmgC5bV4_2),.dout(w_dff_B_8zupik028_2),.clk(gclk));
	jdff dff_B_lKR91fiW8_2(.din(w_dff_B_8zupik028_2),.dout(w_dff_B_lKR91fiW8_2),.clk(gclk));
	jdff dff_B_gmCZ4vL74_2(.din(w_dff_B_lKR91fiW8_2),.dout(w_dff_B_gmCZ4vL74_2),.clk(gclk));
	jdff dff_B_jd2WnOjq9_2(.din(w_dff_B_gmCZ4vL74_2),.dout(w_dff_B_jd2WnOjq9_2),.clk(gclk));
	jdff dff_B_ZiTPcUyT7_2(.din(w_dff_B_jd2WnOjq9_2),.dout(w_dff_B_ZiTPcUyT7_2),.clk(gclk));
	jdff dff_B_UsvavLb55_2(.din(w_dff_B_ZiTPcUyT7_2),.dout(w_dff_B_UsvavLb55_2),.clk(gclk));
	jdff dff_B_63O8CR9r1_2(.din(w_dff_B_UsvavLb55_2),.dout(w_dff_B_63O8CR9r1_2),.clk(gclk));
	jdff dff_B_iNrKj0ju9_2(.din(w_dff_B_63O8CR9r1_2),.dout(w_dff_B_iNrKj0ju9_2),.clk(gclk));
	jdff dff_B_rwpmIUYj5_2(.din(w_dff_B_iNrKj0ju9_2),.dout(w_dff_B_rwpmIUYj5_2),.clk(gclk));
	jdff dff_B_ak1xBx2U8_2(.din(w_dff_B_rwpmIUYj5_2),.dout(w_dff_B_ak1xBx2U8_2),.clk(gclk));
	jdff dff_B_xA4YWT8C0_2(.din(w_dff_B_ak1xBx2U8_2),.dout(w_dff_B_xA4YWT8C0_2),.clk(gclk));
	jdff dff_B_K77LXZyO8_2(.din(w_dff_B_xA4YWT8C0_2),.dout(w_dff_B_K77LXZyO8_2),.clk(gclk));
	jdff dff_B_o72rBbEI4_2(.din(w_dff_B_K77LXZyO8_2),.dout(w_dff_B_o72rBbEI4_2),.clk(gclk));
	jdff dff_B_Mymlih731_2(.din(w_dff_B_o72rBbEI4_2),.dout(w_dff_B_Mymlih731_2),.clk(gclk));
	jdff dff_B_t1oPpmXf2_2(.din(w_dff_B_Mymlih731_2),.dout(w_dff_B_t1oPpmXf2_2),.clk(gclk));
	jdff dff_B_vSj4aknc2_2(.din(w_dff_B_t1oPpmXf2_2),.dout(w_dff_B_vSj4aknc2_2),.clk(gclk));
	jdff dff_B_lluLUQWV3_2(.din(w_dff_B_vSj4aknc2_2),.dout(w_dff_B_lluLUQWV3_2),.clk(gclk));
	jdff dff_B_AKMhD39Q0_2(.din(w_dff_B_lluLUQWV3_2),.dout(w_dff_B_AKMhD39Q0_2),.clk(gclk));
	jdff dff_B_Yp1yWMb26_2(.din(w_dff_B_AKMhD39Q0_2),.dout(w_dff_B_Yp1yWMb26_2),.clk(gclk));
	jdff dff_B_5Zfa1MZy7_2(.din(w_dff_B_Yp1yWMb26_2),.dout(w_dff_B_5Zfa1MZy7_2),.clk(gclk));
	jdff dff_B_DoOjH9fV8_2(.din(w_dff_B_5Zfa1MZy7_2),.dout(w_dff_B_DoOjH9fV8_2),.clk(gclk));
	jdff dff_B_krZPfOzy8_2(.din(n1366),.dout(w_dff_B_krZPfOzy8_2),.clk(gclk));
	jdff dff_B_DgelcY9s0_1(.din(n1328),.dout(w_dff_B_DgelcY9s0_1),.clk(gclk));
	jdff dff_B_n2wlbCTp3_2(.din(n1242),.dout(w_dff_B_n2wlbCTp3_2),.clk(gclk));
	jdff dff_B_iV9qx05D7_2(.din(w_dff_B_n2wlbCTp3_2),.dout(w_dff_B_iV9qx05D7_2),.clk(gclk));
	jdff dff_B_va4LksZJ6_2(.din(w_dff_B_iV9qx05D7_2),.dout(w_dff_B_va4LksZJ6_2),.clk(gclk));
	jdff dff_B_wLd8OlM61_2(.din(w_dff_B_va4LksZJ6_2),.dout(w_dff_B_wLd8OlM61_2),.clk(gclk));
	jdff dff_B_8Tk36hCG3_2(.din(w_dff_B_wLd8OlM61_2),.dout(w_dff_B_8Tk36hCG3_2),.clk(gclk));
	jdff dff_B_WSdfvYBY5_2(.din(w_dff_B_8Tk36hCG3_2),.dout(w_dff_B_WSdfvYBY5_2),.clk(gclk));
	jdff dff_B_m0ZDxtK81_2(.din(w_dff_B_WSdfvYBY5_2),.dout(w_dff_B_m0ZDxtK81_2),.clk(gclk));
	jdff dff_B_lkPEqwj77_2(.din(w_dff_B_m0ZDxtK81_2),.dout(w_dff_B_lkPEqwj77_2),.clk(gclk));
	jdff dff_B_KC6Jr47j8_2(.din(w_dff_B_lkPEqwj77_2),.dout(w_dff_B_KC6Jr47j8_2),.clk(gclk));
	jdff dff_B_lwgW2GI17_2(.din(w_dff_B_KC6Jr47j8_2),.dout(w_dff_B_lwgW2GI17_2),.clk(gclk));
	jdff dff_B_I0V4xDrm2_2(.din(w_dff_B_lwgW2GI17_2),.dout(w_dff_B_I0V4xDrm2_2),.clk(gclk));
	jdff dff_B_IetvA6Mi8_2(.din(w_dff_B_I0V4xDrm2_2),.dout(w_dff_B_IetvA6Mi8_2),.clk(gclk));
	jdff dff_B_Iwr3XN9U5_2(.din(w_dff_B_IetvA6Mi8_2),.dout(w_dff_B_Iwr3XN9U5_2),.clk(gclk));
	jdff dff_B_6RMFK7qw7_2(.din(w_dff_B_Iwr3XN9U5_2),.dout(w_dff_B_6RMFK7qw7_2),.clk(gclk));
	jdff dff_B_iVQFYlep3_2(.din(w_dff_B_6RMFK7qw7_2),.dout(w_dff_B_iVQFYlep3_2),.clk(gclk));
	jdff dff_B_vmfQfqnN2_2(.din(w_dff_B_iVQFYlep3_2),.dout(w_dff_B_vmfQfqnN2_2),.clk(gclk));
	jdff dff_B_Icnrj4Bo2_2(.din(w_dff_B_vmfQfqnN2_2),.dout(w_dff_B_Icnrj4Bo2_2),.clk(gclk));
	jdff dff_B_johYvclZ3_2(.din(w_dff_B_Icnrj4Bo2_2),.dout(w_dff_B_johYvclZ3_2),.clk(gclk));
	jdff dff_B_s4nzUCk26_2(.din(w_dff_B_johYvclZ3_2),.dout(w_dff_B_s4nzUCk26_2),.clk(gclk));
	jdff dff_B_od5SsdDx4_2(.din(w_dff_B_s4nzUCk26_2),.dout(w_dff_B_od5SsdDx4_2),.clk(gclk));
	jdff dff_B_ok7elgaY6_2(.din(w_dff_B_od5SsdDx4_2),.dout(w_dff_B_ok7elgaY6_2),.clk(gclk));
	jdff dff_B_fB6TQAIy2_2(.din(w_dff_B_ok7elgaY6_2),.dout(w_dff_B_fB6TQAIy2_2),.clk(gclk));
	jdff dff_B_IVfJyvYH3_2(.din(w_dff_B_fB6TQAIy2_2),.dout(w_dff_B_IVfJyvYH3_2),.clk(gclk));
	jdff dff_B_KFP4rjqn8_2(.din(w_dff_B_IVfJyvYH3_2),.dout(w_dff_B_KFP4rjqn8_2),.clk(gclk));
	jdff dff_B_VvkALyYG6_2(.din(w_dff_B_KFP4rjqn8_2),.dout(w_dff_B_VvkALyYG6_2),.clk(gclk));
	jdff dff_B_4nNpd3uk5_2(.din(w_dff_B_VvkALyYG6_2),.dout(w_dff_B_4nNpd3uk5_2),.clk(gclk));
	jdff dff_B_3p8Vyoyk6_2(.din(w_dff_B_4nNpd3uk5_2),.dout(w_dff_B_3p8Vyoyk6_2),.clk(gclk));
	jdff dff_B_ixf2x6Qq0_2(.din(w_dff_B_3p8Vyoyk6_2),.dout(w_dff_B_ixf2x6Qq0_2),.clk(gclk));
	jdff dff_B_udHESU6A9_2(.din(w_dff_B_ixf2x6Qq0_2),.dout(w_dff_B_udHESU6A9_2),.clk(gclk));
	jdff dff_B_wqiKM8GG9_2(.din(n1281),.dout(w_dff_B_wqiKM8GG9_2),.clk(gclk));
	jdff dff_B_gdrGJvfb5_1(.din(n1243),.dout(w_dff_B_gdrGJvfb5_1),.clk(gclk));
	jdff dff_B_6LAxITUM1_2(.din(n1151),.dout(w_dff_B_6LAxITUM1_2),.clk(gclk));
	jdff dff_B_wqR3q3tK0_2(.din(w_dff_B_6LAxITUM1_2),.dout(w_dff_B_wqR3q3tK0_2),.clk(gclk));
	jdff dff_B_x46Z4r6u8_2(.din(w_dff_B_wqR3q3tK0_2),.dout(w_dff_B_x46Z4r6u8_2),.clk(gclk));
	jdff dff_B_bZT47peb1_2(.din(w_dff_B_x46Z4r6u8_2),.dout(w_dff_B_bZT47peb1_2),.clk(gclk));
	jdff dff_B_bRNfpkxY2_2(.din(w_dff_B_bZT47peb1_2),.dout(w_dff_B_bRNfpkxY2_2),.clk(gclk));
	jdff dff_B_2IO2lG6n8_2(.din(w_dff_B_bRNfpkxY2_2),.dout(w_dff_B_2IO2lG6n8_2),.clk(gclk));
	jdff dff_B_holTAT613_2(.din(w_dff_B_2IO2lG6n8_2),.dout(w_dff_B_holTAT613_2),.clk(gclk));
	jdff dff_B_mhZVSbhS8_2(.din(w_dff_B_holTAT613_2),.dout(w_dff_B_mhZVSbhS8_2),.clk(gclk));
	jdff dff_B_EL0OK4th6_2(.din(w_dff_B_mhZVSbhS8_2),.dout(w_dff_B_EL0OK4th6_2),.clk(gclk));
	jdff dff_B_wZD3fL640_2(.din(w_dff_B_EL0OK4th6_2),.dout(w_dff_B_wZD3fL640_2),.clk(gclk));
	jdff dff_B_OA5ufeU86_2(.din(w_dff_B_wZD3fL640_2),.dout(w_dff_B_OA5ufeU86_2),.clk(gclk));
	jdff dff_B_6XBoNMvw5_2(.din(w_dff_B_OA5ufeU86_2),.dout(w_dff_B_6XBoNMvw5_2),.clk(gclk));
	jdff dff_B_GNbxkuDy3_2(.din(w_dff_B_6XBoNMvw5_2),.dout(w_dff_B_GNbxkuDy3_2),.clk(gclk));
	jdff dff_B_aHllh0UQ8_2(.din(w_dff_B_GNbxkuDy3_2),.dout(w_dff_B_aHllh0UQ8_2),.clk(gclk));
	jdff dff_B_ORPEDbGn2_2(.din(w_dff_B_aHllh0UQ8_2),.dout(w_dff_B_ORPEDbGn2_2),.clk(gclk));
	jdff dff_B_0LQUf4Ah5_2(.din(w_dff_B_ORPEDbGn2_2),.dout(w_dff_B_0LQUf4Ah5_2),.clk(gclk));
	jdff dff_B_6JmgZ9PH7_2(.din(w_dff_B_0LQUf4Ah5_2),.dout(w_dff_B_6JmgZ9PH7_2),.clk(gclk));
	jdff dff_B_He58tmNP8_2(.din(w_dff_B_6JmgZ9PH7_2),.dout(w_dff_B_He58tmNP8_2),.clk(gclk));
	jdff dff_B_PrL1D6tf4_2(.din(w_dff_B_He58tmNP8_2),.dout(w_dff_B_PrL1D6tf4_2),.clk(gclk));
	jdff dff_B_aZCe5bF60_2(.din(w_dff_B_PrL1D6tf4_2),.dout(w_dff_B_aZCe5bF60_2),.clk(gclk));
	jdff dff_B_Ueu599mm7_2(.din(w_dff_B_aZCe5bF60_2),.dout(w_dff_B_Ueu599mm7_2),.clk(gclk));
	jdff dff_B_RHUtLhne3_2(.din(w_dff_B_Ueu599mm7_2),.dout(w_dff_B_RHUtLhne3_2),.clk(gclk));
	jdff dff_B_M4GdUuWq6_2(.din(w_dff_B_RHUtLhne3_2),.dout(w_dff_B_M4GdUuWq6_2),.clk(gclk));
	jdff dff_B_VZqh0cDT6_2(.din(w_dff_B_M4GdUuWq6_2),.dout(w_dff_B_VZqh0cDT6_2),.clk(gclk));
	jdff dff_B_IhLGXj228_2(.din(w_dff_B_VZqh0cDT6_2),.dout(w_dff_B_IhLGXj228_2),.clk(gclk));
	jdff dff_B_lGtpcAJp7_2(.din(w_dff_B_IhLGXj228_2),.dout(w_dff_B_lGtpcAJp7_2),.clk(gclk));
	jdff dff_B_03qnLCe22_2(.din(n1190),.dout(w_dff_B_03qnLCe22_2),.clk(gclk));
	jdff dff_B_hbAs9MRE7_1(.din(n1152),.dout(w_dff_B_hbAs9MRE7_1),.clk(gclk));
	jdff dff_B_7YSbfqLc6_2(.din(n1053),.dout(w_dff_B_7YSbfqLc6_2),.clk(gclk));
	jdff dff_B_br1dIeQV4_2(.din(w_dff_B_7YSbfqLc6_2),.dout(w_dff_B_br1dIeQV4_2),.clk(gclk));
	jdff dff_B_KpEuoHQc7_2(.din(w_dff_B_br1dIeQV4_2),.dout(w_dff_B_KpEuoHQc7_2),.clk(gclk));
	jdff dff_B_nH6yqGFt7_2(.din(w_dff_B_KpEuoHQc7_2),.dout(w_dff_B_nH6yqGFt7_2),.clk(gclk));
	jdff dff_B_k7FErPul7_2(.din(w_dff_B_nH6yqGFt7_2),.dout(w_dff_B_k7FErPul7_2),.clk(gclk));
	jdff dff_B_n9aGapcV5_2(.din(w_dff_B_k7FErPul7_2),.dout(w_dff_B_n9aGapcV5_2),.clk(gclk));
	jdff dff_B_NVE8bpjW7_2(.din(w_dff_B_n9aGapcV5_2),.dout(w_dff_B_NVE8bpjW7_2),.clk(gclk));
	jdff dff_B_bK2InPNT6_2(.din(w_dff_B_NVE8bpjW7_2),.dout(w_dff_B_bK2InPNT6_2),.clk(gclk));
	jdff dff_B_oWdkY0Gi6_2(.din(w_dff_B_bK2InPNT6_2),.dout(w_dff_B_oWdkY0Gi6_2),.clk(gclk));
	jdff dff_B_rfjTdLWg6_2(.din(w_dff_B_oWdkY0Gi6_2),.dout(w_dff_B_rfjTdLWg6_2),.clk(gclk));
	jdff dff_B_6OlVESxY9_2(.din(w_dff_B_rfjTdLWg6_2),.dout(w_dff_B_6OlVESxY9_2),.clk(gclk));
	jdff dff_B_uqLgkRFO9_2(.din(w_dff_B_6OlVESxY9_2),.dout(w_dff_B_uqLgkRFO9_2),.clk(gclk));
	jdff dff_B_Lnio3Zql7_2(.din(w_dff_B_uqLgkRFO9_2),.dout(w_dff_B_Lnio3Zql7_2),.clk(gclk));
	jdff dff_B_z4nlAwtf6_2(.din(w_dff_B_Lnio3Zql7_2),.dout(w_dff_B_z4nlAwtf6_2),.clk(gclk));
	jdff dff_B_DvKdE5fy1_2(.din(w_dff_B_z4nlAwtf6_2),.dout(w_dff_B_DvKdE5fy1_2),.clk(gclk));
	jdff dff_B_ZFyPLXeB2_2(.din(w_dff_B_DvKdE5fy1_2),.dout(w_dff_B_ZFyPLXeB2_2),.clk(gclk));
	jdff dff_B_PXKTojbK7_2(.din(w_dff_B_ZFyPLXeB2_2),.dout(w_dff_B_PXKTojbK7_2),.clk(gclk));
	jdff dff_B_qxRhpnAz0_2(.din(w_dff_B_PXKTojbK7_2),.dout(w_dff_B_qxRhpnAz0_2),.clk(gclk));
	jdff dff_B_OsCNhheQ6_2(.din(w_dff_B_qxRhpnAz0_2),.dout(w_dff_B_OsCNhheQ6_2),.clk(gclk));
	jdff dff_B_Z02BIdNg0_2(.din(w_dff_B_OsCNhheQ6_2),.dout(w_dff_B_Z02BIdNg0_2),.clk(gclk));
	jdff dff_B_Ebr1VH9l9_2(.din(w_dff_B_Z02BIdNg0_2),.dout(w_dff_B_Ebr1VH9l9_2),.clk(gclk));
	jdff dff_B_pVJGLeRL7_2(.din(w_dff_B_Ebr1VH9l9_2),.dout(w_dff_B_pVJGLeRL7_2),.clk(gclk));
	jdff dff_B_ao91obDv1_2(.din(w_dff_B_pVJGLeRL7_2),.dout(w_dff_B_ao91obDv1_2),.clk(gclk));
	jdff dff_B_4xpjW6mv9_2(.din(n1091),.dout(w_dff_B_4xpjW6mv9_2),.clk(gclk));
	jdff dff_B_LAVnKpcM7_1(.din(n1054),.dout(w_dff_B_LAVnKpcM7_1),.clk(gclk));
	jdff dff_B_3BT3or5H8_2(.din(n954),.dout(w_dff_B_3BT3or5H8_2),.clk(gclk));
	jdff dff_B_Z4EtcHTU7_2(.din(w_dff_B_3BT3or5H8_2),.dout(w_dff_B_Z4EtcHTU7_2),.clk(gclk));
	jdff dff_B_HU98oJWt6_2(.din(w_dff_B_Z4EtcHTU7_2),.dout(w_dff_B_HU98oJWt6_2),.clk(gclk));
	jdff dff_B_Z1xelDDy1_2(.din(w_dff_B_HU98oJWt6_2),.dout(w_dff_B_Z1xelDDy1_2),.clk(gclk));
	jdff dff_B_trYHmvBe8_2(.din(w_dff_B_Z1xelDDy1_2),.dout(w_dff_B_trYHmvBe8_2),.clk(gclk));
	jdff dff_B_4gKp8EFT8_2(.din(w_dff_B_trYHmvBe8_2),.dout(w_dff_B_4gKp8EFT8_2),.clk(gclk));
	jdff dff_B_AF0608h03_2(.din(w_dff_B_4gKp8EFT8_2),.dout(w_dff_B_AF0608h03_2),.clk(gclk));
	jdff dff_B_YtbohqzK5_2(.din(w_dff_B_AF0608h03_2),.dout(w_dff_B_YtbohqzK5_2),.clk(gclk));
	jdff dff_B_OkgsXH552_2(.din(w_dff_B_YtbohqzK5_2),.dout(w_dff_B_OkgsXH552_2),.clk(gclk));
	jdff dff_B_H5s0HGV35_2(.din(w_dff_B_OkgsXH552_2),.dout(w_dff_B_H5s0HGV35_2),.clk(gclk));
	jdff dff_B_frD7O9NK8_2(.din(w_dff_B_H5s0HGV35_2),.dout(w_dff_B_frD7O9NK8_2),.clk(gclk));
	jdff dff_B_1m8GGWQI6_2(.din(w_dff_B_frD7O9NK8_2),.dout(w_dff_B_1m8GGWQI6_2),.clk(gclk));
	jdff dff_B_CR7uknkT1_2(.din(w_dff_B_1m8GGWQI6_2),.dout(w_dff_B_CR7uknkT1_2),.clk(gclk));
	jdff dff_B_rq8TM1ly0_2(.din(w_dff_B_CR7uknkT1_2),.dout(w_dff_B_rq8TM1ly0_2),.clk(gclk));
	jdff dff_B_yZ2DPA2L6_2(.din(w_dff_B_rq8TM1ly0_2),.dout(w_dff_B_yZ2DPA2L6_2),.clk(gclk));
	jdff dff_B_qPRdAYD37_2(.din(w_dff_B_yZ2DPA2L6_2),.dout(w_dff_B_qPRdAYD37_2),.clk(gclk));
	jdff dff_B_kYnLVwGx9_2(.din(w_dff_B_qPRdAYD37_2),.dout(w_dff_B_kYnLVwGx9_2),.clk(gclk));
	jdff dff_B_ADDWrBKg7_2(.din(w_dff_B_kYnLVwGx9_2),.dout(w_dff_B_ADDWrBKg7_2),.clk(gclk));
	jdff dff_B_zNLnX71z2_2(.din(w_dff_B_ADDWrBKg7_2),.dout(w_dff_B_zNLnX71z2_2),.clk(gclk));
	jdff dff_B_d4nEiHRz9_2(.din(w_dff_B_zNLnX71z2_2),.dout(w_dff_B_d4nEiHRz9_2),.clk(gclk));
	jdff dff_B_aoIjgNAi7_2(.din(n992),.dout(w_dff_B_aoIjgNAi7_2),.clk(gclk));
	jdff dff_B_RYkSGtmM3_1(.din(n955),.dout(w_dff_B_RYkSGtmM3_1),.clk(gclk));
	jdff dff_B_YUD9nspG2_2(.din(n852),.dout(w_dff_B_YUD9nspG2_2),.clk(gclk));
	jdff dff_B_UUqmA8X71_2(.din(w_dff_B_YUD9nspG2_2),.dout(w_dff_B_UUqmA8X71_2),.clk(gclk));
	jdff dff_B_aubJzKXX8_2(.din(w_dff_B_UUqmA8X71_2),.dout(w_dff_B_aubJzKXX8_2),.clk(gclk));
	jdff dff_B_qhmQ3wqw2_2(.din(w_dff_B_aubJzKXX8_2),.dout(w_dff_B_qhmQ3wqw2_2),.clk(gclk));
	jdff dff_B_JRoSQOaS8_2(.din(w_dff_B_qhmQ3wqw2_2),.dout(w_dff_B_JRoSQOaS8_2),.clk(gclk));
	jdff dff_B_48cd8Bc66_2(.din(w_dff_B_JRoSQOaS8_2),.dout(w_dff_B_48cd8Bc66_2),.clk(gclk));
	jdff dff_B_EG6g5fEI9_2(.din(w_dff_B_48cd8Bc66_2),.dout(w_dff_B_EG6g5fEI9_2),.clk(gclk));
	jdff dff_B_n5FdlT3x7_2(.din(w_dff_B_EG6g5fEI9_2),.dout(w_dff_B_n5FdlT3x7_2),.clk(gclk));
	jdff dff_B_1ZaeDNct5_2(.din(w_dff_B_n5FdlT3x7_2),.dout(w_dff_B_1ZaeDNct5_2),.clk(gclk));
	jdff dff_B_bgmMBiAu4_2(.din(w_dff_B_1ZaeDNct5_2),.dout(w_dff_B_bgmMBiAu4_2),.clk(gclk));
	jdff dff_B_oJ3U0Udn5_2(.din(w_dff_B_bgmMBiAu4_2),.dout(w_dff_B_oJ3U0Udn5_2),.clk(gclk));
	jdff dff_B_6WqpbwZZ0_2(.din(w_dff_B_oJ3U0Udn5_2),.dout(w_dff_B_6WqpbwZZ0_2),.clk(gclk));
	jdff dff_B_EFo5p8J57_2(.din(w_dff_B_6WqpbwZZ0_2),.dout(w_dff_B_EFo5p8J57_2),.clk(gclk));
	jdff dff_B_J8iXcCjd8_2(.din(w_dff_B_EFo5p8J57_2),.dout(w_dff_B_J8iXcCjd8_2),.clk(gclk));
	jdff dff_B_AqMfvCMo8_2(.din(w_dff_B_J8iXcCjd8_2),.dout(w_dff_B_AqMfvCMo8_2),.clk(gclk));
	jdff dff_B_8C8LvwYj9_2(.din(w_dff_B_AqMfvCMo8_2),.dout(w_dff_B_8C8LvwYj9_2),.clk(gclk));
	jdff dff_B_atvicVez0_2(.din(w_dff_B_8C8LvwYj9_2),.dout(w_dff_B_atvicVez0_2),.clk(gclk));
	jdff dff_B_q9E9E1EZ5_2(.din(n886),.dout(w_dff_B_q9E9E1EZ5_2),.clk(gclk));
	jdff dff_B_pky1lf7R0_1(.din(n853),.dout(w_dff_B_pky1lf7R0_1),.clk(gclk));
	jdff dff_B_cop3KlzS0_2(.din(n754),.dout(w_dff_B_cop3KlzS0_2),.clk(gclk));
	jdff dff_B_7Pfajhzu8_2(.din(w_dff_B_cop3KlzS0_2),.dout(w_dff_B_7Pfajhzu8_2),.clk(gclk));
	jdff dff_B_Qa3fqE9G6_2(.din(w_dff_B_7Pfajhzu8_2),.dout(w_dff_B_Qa3fqE9G6_2),.clk(gclk));
	jdff dff_B_WL7rJb5t8_2(.din(w_dff_B_Qa3fqE9G6_2),.dout(w_dff_B_WL7rJb5t8_2),.clk(gclk));
	jdff dff_B_81MAUXDq3_2(.din(w_dff_B_WL7rJb5t8_2),.dout(w_dff_B_81MAUXDq3_2),.clk(gclk));
	jdff dff_B_bI8U3JD88_2(.din(w_dff_B_81MAUXDq3_2),.dout(w_dff_B_bI8U3JD88_2),.clk(gclk));
	jdff dff_B_SOrQUK9g3_2(.din(w_dff_B_bI8U3JD88_2),.dout(w_dff_B_SOrQUK9g3_2),.clk(gclk));
	jdff dff_B_bn8T6aC32_2(.din(w_dff_B_SOrQUK9g3_2),.dout(w_dff_B_bn8T6aC32_2),.clk(gclk));
	jdff dff_B_MxMY04SY1_2(.din(w_dff_B_bn8T6aC32_2),.dout(w_dff_B_MxMY04SY1_2),.clk(gclk));
	jdff dff_B_hoD6JlkO7_2(.din(w_dff_B_MxMY04SY1_2),.dout(w_dff_B_hoD6JlkO7_2),.clk(gclk));
	jdff dff_B_QCN9vbEl6_2(.din(w_dff_B_hoD6JlkO7_2),.dout(w_dff_B_QCN9vbEl6_2),.clk(gclk));
	jdff dff_B_XkTyAUcG1_2(.din(w_dff_B_QCN9vbEl6_2),.dout(w_dff_B_XkTyAUcG1_2),.clk(gclk));
	jdff dff_B_CkImynzt0_2(.din(w_dff_B_XkTyAUcG1_2),.dout(w_dff_B_CkImynzt0_2),.clk(gclk));
	jdff dff_B_vtGoz9zg2_2(.din(w_dff_B_CkImynzt0_2),.dout(w_dff_B_vtGoz9zg2_2),.clk(gclk));
	jdff dff_B_GvEQLVg08_2(.din(n783),.dout(w_dff_B_GvEQLVg08_2),.clk(gclk));
	jdff dff_B_QHE2z7Ie5_1(.din(n755),.dout(w_dff_B_QHE2z7Ie5_1),.clk(gclk));
	jdff dff_B_bLxyMb3P9_2(.din(n662),.dout(w_dff_B_bLxyMb3P9_2),.clk(gclk));
	jdff dff_B_cvBs6jAA5_2(.din(w_dff_B_bLxyMb3P9_2),.dout(w_dff_B_cvBs6jAA5_2),.clk(gclk));
	jdff dff_B_Kg8QyU639_2(.din(w_dff_B_cvBs6jAA5_2),.dout(w_dff_B_Kg8QyU639_2),.clk(gclk));
	jdff dff_B_WKoQoKNC6_2(.din(w_dff_B_Kg8QyU639_2),.dout(w_dff_B_WKoQoKNC6_2),.clk(gclk));
	jdff dff_B_IBDF3cDn0_2(.din(w_dff_B_WKoQoKNC6_2),.dout(w_dff_B_IBDF3cDn0_2),.clk(gclk));
	jdff dff_B_tzQdXW0o1_2(.din(w_dff_B_IBDF3cDn0_2),.dout(w_dff_B_tzQdXW0o1_2),.clk(gclk));
	jdff dff_B_9JWlaWHN3_2(.din(w_dff_B_tzQdXW0o1_2),.dout(w_dff_B_9JWlaWHN3_2),.clk(gclk));
	jdff dff_B_kYa6cxna7_2(.din(w_dff_B_9JWlaWHN3_2),.dout(w_dff_B_kYa6cxna7_2),.clk(gclk));
	jdff dff_B_PhvJ10wD4_2(.din(w_dff_B_kYa6cxna7_2),.dout(w_dff_B_PhvJ10wD4_2),.clk(gclk));
	jdff dff_B_z02FG4Ot5_2(.din(w_dff_B_PhvJ10wD4_2),.dout(w_dff_B_z02FG4Ot5_2),.clk(gclk));
	jdff dff_B_kjssqN031_2(.din(w_dff_B_z02FG4Ot5_2),.dout(w_dff_B_kjssqN031_2),.clk(gclk));
	jdff dff_B_R87REC4W0_2(.din(n684),.dout(w_dff_B_R87REC4W0_2),.clk(gclk));
	jdff dff_B_YlGTExVH1_1(.din(n663),.dout(w_dff_B_YlGTExVH1_1),.clk(gclk));
	jdff dff_B_ePkst0b07_2(.din(n577),.dout(w_dff_B_ePkst0b07_2),.clk(gclk));
	jdff dff_B_087CWndQ4_2(.din(w_dff_B_ePkst0b07_2),.dout(w_dff_B_087CWndQ4_2),.clk(gclk));
	jdff dff_B_UsXfUvZq6_2(.din(w_dff_B_087CWndQ4_2),.dout(w_dff_B_UsXfUvZq6_2),.clk(gclk));
	jdff dff_B_87JjQ5LB2_2(.din(w_dff_B_UsXfUvZq6_2),.dout(w_dff_B_87JjQ5LB2_2),.clk(gclk));
	jdff dff_B_hfEbtF9y3_2(.din(w_dff_B_87JjQ5LB2_2),.dout(w_dff_B_hfEbtF9y3_2),.clk(gclk));
	jdff dff_B_wIRjB66Y0_2(.din(w_dff_B_hfEbtF9y3_2),.dout(w_dff_B_wIRjB66Y0_2),.clk(gclk));
	jdff dff_B_va1fvv802_2(.din(w_dff_B_wIRjB66Y0_2),.dout(w_dff_B_va1fvv802_2),.clk(gclk));
	jdff dff_B_fFbYDQIW4_2(.din(w_dff_B_va1fvv802_2),.dout(w_dff_B_fFbYDQIW4_2),.clk(gclk));
	jdff dff_B_S4QVlaXz1_2(.din(n592),.dout(w_dff_B_S4QVlaXz1_2),.clk(gclk));
	jdff dff_B_VvMOypjG3_2(.din(w_dff_B_S4QVlaXz1_2),.dout(w_dff_B_VvMOypjG3_2),.clk(gclk));
	jdff dff_B_nCxF0Fs43_2(.din(w_dff_B_VvMOypjG3_2),.dout(w_dff_B_nCxF0Fs43_2),.clk(gclk));
	jdff dff_B_HWfi7Esq8_1(.din(n578),.dout(w_dff_B_HWfi7Esq8_1),.clk(gclk));
	jdff dff_B_6q58Zi7A0_1(.din(w_dff_B_HWfi7Esq8_1),.dout(w_dff_B_6q58Zi7A0_1),.clk(gclk));
	jdff dff_B_ATyUjume4_2(.din(n501),.dout(w_dff_B_ATyUjume4_2),.clk(gclk));
	jdff dff_B_HjpMqqJB6_2(.din(w_dff_B_ATyUjume4_2),.dout(w_dff_B_HjpMqqJB6_2),.clk(gclk));
	jdff dff_B_wPhdDcjg4_2(.din(w_dff_B_HjpMqqJB6_2),.dout(w_dff_B_wPhdDcjg4_2),.clk(gclk));
	jdff dff_B_JIdhCC2w7_0(.din(n506),.dout(w_dff_B_JIdhCC2w7_0),.clk(gclk));
	jdff dff_A_kmoZ7gjB8_0(.dout(w_n427_0[0]),.din(w_dff_A_kmoZ7gjB8_0),.clk(gclk));
	jdff dff_A_qgqYeQLl3_0(.dout(w_dff_A_kmoZ7gjB8_0),.din(w_dff_A_qgqYeQLl3_0),.clk(gclk));
	jdff dff_A_hGhDz4u86_1(.dout(w_n427_0[1]),.din(w_dff_A_hGhDz4u86_1),.clk(gclk));
	jdff dff_A_qSqHHLZm1_1(.dout(w_dff_A_hGhDz4u86_1),.din(w_dff_A_qSqHHLZm1_1),.clk(gclk));
	jdff dff_B_RNmKnxNj1_1(.din(n1729),.dout(w_dff_B_RNmKnxNj1_1),.clk(gclk));
	jdff dff_A_kB4EvvLH8_1(.dout(w_n1697_0[1]),.din(w_dff_A_kB4EvvLH8_1),.clk(gclk));
	jdff dff_B_EjhvP3lH5_1(.din(n1695),.dout(w_dff_B_EjhvP3lH5_1),.clk(gclk));
	jdff dff_B_86NpWNeW8_2(.din(n1653),.dout(w_dff_B_86NpWNeW8_2),.clk(gclk));
	jdff dff_B_MHrQKCMV5_2(.din(w_dff_B_86NpWNeW8_2),.dout(w_dff_B_MHrQKCMV5_2),.clk(gclk));
	jdff dff_B_2YxjOSjQ7_2(.din(w_dff_B_MHrQKCMV5_2),.dout(w_dff_B_2YxjOSjQ7_2),.clk(gclk));
	jdff dff_B_DxQyfBfM7_2(.din(w_dff_B_2YxjOSjQ7_2),.dout(w_dff_B_DxQyfBfM7_2),.clk(gclk));
	jdff dff_B_1ZJYhFPx1_2(.din(w_dff_B_DxQyfBfM7_2),.dout(w_dff_B_1ZJYhFPx1_2),.clk(gclk));
	jdff dff_B_ZGAvkeWZ3_2(.din(w_dff_B_1ZJYhFPx1_2),.dout(w_dff_B_ZGAvkeWZ3_2),.clk(gclk));
	jdff dff_B_wY2YYS6D7_2(.din(w_dff_B_ZGAvkeWZ3_2),.dout(w_dff_B_wY2YYS6D7_2),.clk(gclk));
	jdff dff_B_nwQcUs8N8_2(.din(w_dff_B_wY2YYS6D7_2),.dout(w_dff_B_nwQcUs8N8_2),.clk(gclk));
	jdff dff_B_rRVXfMNa0_2(.din(w_dff_B_nwQcUs8N8_2),.dout(w_dff_B_rRVXfMNa0_2),.clk(gclk));
	jdff dff_B_oYbLJG688_2(.din(w_dff_B_rRVXfMNa0_2),.dout(w_dff_B_oYbLJG688_2),.clk(gclk));
	jdff dff_B_I4PYwhX82_2(.din(w_dff_B_oYbLJG688_2),.dout(w_dff_B_I4PYwhX82_2),.clk(gclk));
	jdff dff_B_e4Ss7TB39_2(.din(w_dff_B_I4PYwhX82_2),.dout(w_dff_B_e4Ss7TB39_2),.clk(gclk));
	jdff dff_B_9US6O8uT3_2(.din(w_dff_B_e4Ss7TB39_2),.dout(w_dff_B_9US6O8uT3_2),.clk(gclk));
	jdff dff_B_swadolk93_2(.din(w_dff_B_9US6O8uT3_2),.dout(w_dff_B_swadolk93_2),.clk(gclk));
	jdff dff_B_HS4oMSVO2_2(.din(w_dff_B_swadolk93_2),.dout(w_dff_B_HS4oMSVO2_2),.clk(gclk));
	jdff dff_B_4TPCzsBT0_2(.din(w_dff_B_HS4oMSVO2_2),.dout(w_dff_B_4TPCzsBT0_2),.clk(gclk));
	jdff dff_B_PUCIrwSb8_2(.din(w_dff_B_4TPCzsBT0_2),.dout(w_dff_B_PUCIrwSb8_2),.clk(gclk));
	jdff dff_B_iS7dKMz94_2(.din(w_dff_B_PUCIrwSb8_2),.dout(w_dff_B_iS7dKMz94_2),.clk(gclk));
	jdff dff_B_ud2SorNx9_2(.din(w_dff_B_iS7dKMz94_2),.dout(w_dff_B_ud2SorNx9_2),.clk(gclk));
	jdff dff_B_44ClnKSg6_2(.din(w_dff_B_ud2SorNx9_2),.dout(w_dff_B_44ClnKSg6_2),.clk(gclk));
	jdff dff_B_AmEBpAcH4_2(.din(w_dff_B_44ClnKSg6_2),.dout(w_dff_B_AmEBpAcH4_2),.clk(gclk));
	jdff dff_B_D1n7xwRJ6_2(.din(w_dff_B_AmEBpAcH4_2),.dout(w_dff_B_D1n7xwRJ6_2),.clk(gclk));
	jdff dff_B_uga1Kz5B5_2(.din(w_dff_B_D1n7xwRJ6_2),.dout(w_dff_B_uga1Kz5B5_2),.clk(gclk));
	jdff dff_B_VFfhgVS75_2(.din(w_dff_B_uga1Kz5B5_2),.dout(w_dff_B_VFfhgVS75_2),.clk(gclk));
	jdff dff_B_HmIja5Vp0_2(.din(w_dff_B_VFfhgVS75_2),.dout(w_dff_B_HmIja5Vp0_2),.clk(gclk));
	jdff dff_B_C9x4hNgZ1_2(.din(w_dff_B_HmIja5Vp0_2),.dout(w_dff_B_C9x4hNgZ1_2),.clk(gclk));
	jdff dff_B_tkL76kbB1_2(.din(w_dff_B_C9x4hNgZ1_2),.dout(w_dff_B_tkL76kbB1_2),.clk(gclk));
	jdff dff_B_oG3I6i9v9_2(.din(w_dff_B_tkL76kbB1_2),.dout(w_dff_B_oG3I6i9v9_2),.clk(gclk));
	jdff dff_B_ab25Dm6h1_2(.din(w_dff_B_oG3I6i9v9_2),.dout(w_dff_B_ab25Dm6h1_2),.clk(gclk));
	jdff dff_B_bhFxR8fG6_2(.din(w_dff_B_ab25Dm6h1_2),.dout(w_dff_B_bhFxR8fG6_2),.clk(gclk));
	jdff dff_B_0ecvAmry6_2(.din(w_dff_B_bhFxR8fG6_2),.dout(w_dff_B_0ecvAmry6_2),.clk(gclk));
	jdff dff_B_A0HQTnRS5_2(.din(w_dff_B_0ecvAmry6_2),.dout(w_dff_B_A0HQTnRS5_2),.clk(gclk));
	jdff dff_B_1Ji9BOsi7_2(.din(w_dff_B_A0HQTnRS5_2),.dout(w_dff_B_1Ji9BOsi7_2),.clk(gclk));
	jdff dff_B_LaJRO3fp4_2(.din(w_dff_B_1Ji9BOsi7_2),.dout(w_dff_B_LaJRO3fp4_2),.clk(gclk));
	jdff dff_B_FV0XBqGk8_2(.din(w_dff_B_LaJRO3fp4_2),.dout(w_dff_B_FV0XBqGk8_2),.clk(gclk));
	jdff dff_B_NjCPu9Mz0_2(.din(w_dff_B_FV0XBqGk8_2),.dout(w_dff_B_NjCPu9Mz0_2),.clk(gclk));
	jdff dff_B_I0iEEkOt3_2(.din(w_dff_B_NjCPu9Mz0_2),.dout(w_dff_B_I0iEEkOt3_2),.clk(gclk));
	jdff dff_B_Lt0jMCye4_2(.din(w_dff_B_I0iEEkOt3_2),.dout(w_dff_B_Lt0jMCye4_2),.clk(gclk));
	jdff dff_B_GGFHYT3U8_2(.din(w_dff_B_Lt0jMCye4_2),.dout(w_dff_B_GGFHYT3U8_2),.clk(gclk));
	jdff dff_B_tkUk5iCJ8_2(.din(w_dff_B_GGFHYT3U8_2),.dout(w_dff_B_tkUk5iCJ8_2),.clk(gclk));
	jdff dff_B_kpk8K8ZK8_2(.din(w_dff_B_tkUk5iCJ8_2),.dout(w_dff_B_kpk8K8ZK8_2),.clk(gclk));
	jdff dff_B_VzYXxpMT1_2(.din(w_dff_B_kpk8K8ZK8_2),.dout(w_dff_B_VzYXxpMT1_2),.clk(gclk));
	jdff dff_B_jRGarOmj8_2(.din(w_dff_B_VzYXxpMT1_2),.dout(w_dff_B_jRGarOmj8_2),.clk(gclk));
	jdff dff_B_vwd53Nsd6_2(.din(w_dff_B_jRGarOmj8_2),.dout(w_dff_B_vwd53Nsd6_2),.clk(gclk));
	jdff dff_B_ogga8Sqf7_2(.din(w_dff_B_vwd53Nsd6_2),.dout(w_dff_B_ogga8Sqf7_2),.clk(gclk));
	jdff dff_B_pE3RY6EJ3_2(.din(w_dff_B_ogga8Sqf7_2),.dout(w_dff_B_pE3RY6EJ3_2),.clk(gclk));
	jdff dff_B_sNHG63tc4_2(.din(n1656),.dout(w_dff_B_sNHG63tc4_2),.clk(gclk));
	jdff dff_B_Hda611ca5_1(.din(n1654),.dout(w_dff_B_Hda611ca5_1),.clk(gclk));
	jdff dff_B_zXXELH222_2(.din(n1602),.dout(w_dff_B_zXXELH222_2),.clk(gclk));
	jdff dff_B_Q5Wo0zzI6_2(.din(w_dff_B_zXXELH222_2),.dout(w_dff_B_Q5Wo0zzI6_2),.clk(gclk));
	jdff dff_B_hFCgGp9V9_2(.din(w_dff_B_Q5Wo0zzI6_2),.dout(w_dff_B_hFCgGp9V9_2),.clk(gclk));
	jdff dff_B_ZIWHJBJw3_2(.din(w_dff_B_hFCgGp9V9_2),.dout(w_dff_B_ZIWHJBJw3_2),.clk(gclk));
	jdff dff_B_aIgN8ii19_2(.din(w_dff_B_ZIWHJBJw3_2),.dout(w_dff_B_aIgN8ii19_2),.clk(gclk));
	jdff dff_B_YZOVsGuE4_2(.din(w_dff_B_aIgN8ii19_2),.dout(w_dff_B_YZOVsGuE4_2),.clk(gclk));
	jdff dff_B_MGVTiXsw6_2(.din(w_dff_B_YZOVsGuE4_2),.dout(w_dff_B_MGVTiXsw6_2),.clk(gclk));
	jdff dff_B_78Qz7F2r8_2(.din(w_dff_B_MGVTiXsw6_2),.dout(w_dff_B_78Qz7F2r8_2),.clk(gclk));
	jdff dff_B_sfvx99TZ5_2(.din(w_dff_B_78Qz7F2r8_2),.dout(w_dff_B_sfvx99TZ5_2),.clk(gclk));
	jdff dff_B_0PMYyms69_2(.din(w_dff_B_sfvx99TZ5_2),.dout(w_dff_B_0PMYyms69_2),.clk(gclk));
	jdff dff_B_sOnGZSRu0_2(.din(w_dff_B_0PMYyms69_2),.dout(w_dff_B_sOnGZSRu0_2),.clk(gclk));
	jdff dff_B_jZsMk6Zv9_2(.din(w_dff_B_sOnGZSRu0_2),.dout(w_dff_B_jZsMk6Zv9_2),.clk(gclk));
	jdff dff_B_JmUourcI3_2(.din(w_dff_B_jZsMk6Zv9_2),.dout(w_dff_B_JmUourcI3_2),.clk(gclk));
	jdff dff_B_27738wuW2_2(.din(w_dff_B_JmUourcI3_2),.dout(w_dff_B_27738wuW2_2),.clk(gclk));
	jdff dff_B_C1SmVTst8_2(.din(w_dff_B_27738wuW2_2),.dout(w_dff_B_C1SmVTst8_2),.clk(gclk));
	jdff dff_B_QNWiyBi36_2(.din(w_dff_B_C1SmVTst8_2),.dout(w_dff_B_QNWiyBi36_2),.clk(gclk));
	jdff dff_B_xdFx4idk7_2(.din(w_dff_B_QNWiyBi36_2),.dout(w_dff_B_xdFx4idk7_2),.clk(gclk));
	jdff dff_B_cHjPVH1P8_2(.din(w_dff_B_xdFx4idk7_2),.dout(w_dff_B_cHjPVH1P8_2),.clk(gclk));
	jdff dff_B_J99FYGp43_2(.din(w_dff_B_cHjPVH1P8_2),.dout(w_dff_B_J99FYGp43_2),.clk(gclk));
	jdff dff_B_JP3qFZba7_2(.din(w_dff_B_J99FYGp43_2),.dout(w_dff_B_JP3qFZba7_2),.clk(gclk));
	jdff dff_B_3oMdCaRj7_2(.din(w_dff_B_JP3qFZba7_2),.dout(w_dff_B_3oMdCaRj7_2),.clk(gclk));
	jdff dff_B_QFVFKalo4_2(.din(w_dff_B_3oMdCaRj7_2),.dout(w_dff_B_QFVFKalo4_2),.clk(gclk));
	jdff dff_B_8T1GbwaS4_2(.din(w_dff_B_QFVFKalo4_2),.dout(w_dff_B_8T1GbwaS4_2),.clk(gclk));
	jdff dff_B_KPiNWqn23_2(.din(w_dff_B_8T1GbwaS4_2),.dout(w_dff_B_KPiNWqn23_2),.clk(gclk));
	jdff dff_B_lmoQQE0S4_2(.din(w_dff_B_KPiNWqn23_2),.dout(w_dff_B_lmoQQE0S4_2),.clk(gclk));
	jdff dff_B_gXzfq2pK9_2(.din(w_dff_B_lmoQQE0S4_2),.dout(w_dff_B_gXzfq2pK9_2),.clk(gclk));
	jdff dff_B_yVuYxYSV7_2(.din(w_dff_B_gXzfq2pK9_2),.dout(w_dff_B_yVuYxYSV7_2),.clk(gclk));
	jdff dff_B_5fYUDq1q6_2(.din(w_dff_B_yVuYxYSV7_2),.dout(w_dff_B_5fYUDq1q6_2),.clk(gclk));
	jdff dff_B_2WKPpk5e7_2(.din(w_dff_B_5fYUDq1q6_2),.dout(w_dff_B_2WKPpk5e7_2),.clk(gclk));
	jdff dff_B_zPGj7Znh0_2(.din(w_dff_B_2WKPpk5e7_2),.dout(w_dff_B_zPGj7Znh0_2),.clk(gclk));
	jdff dff_B_GML0Fae86_2(.din(w_dff_B_zPGj7Znh0_2),.dout(w_dff_B_GML0Fae86_2),.clk(gclk));
	jdff dff_B_pJOJ8wix4_2(.din(w_dff_B_GML0Fae86_2),.dout(w_dff_B_pJOJ8wix4_2),.clk(gclk));
	jdff dff_B_xemwHUVc7_2(.din(w_dff_B_pJOJ8wix4_2),.dout(w_dff_B_xemwHUVc7_2),.clk(gclk));
	jdff dff_B_ttnCY9od6_2(.din(w_dff_B_xemwHUVc7_2),.dout(w_dff_B_ttnCY9od6_2),.clk(gclk));
	jdff dff_B_E8XeTHSK4_2(.din(w_dff_B_ttnCY9od6_2),.dout(w_dff_B_E8XeTHSK4_2),.clk(gclk));
	jdff dff_B_SfNyBD0v8_2(.din(w_dff_B_E8XeTHSK4_2),.dout(w_dff_B_SfNyBD0v8_2),.clk(gclk));
	jdff dff_B_vZKQ6Mfu5_2(.din(w_dff_B_SfNyBD0v8_2),.dout(w_dff_B_vZKQ6Mfu5_2),.clk(gclk));
	jdff dff_B_w5g9bPqK3_2(.din(w_dff_B_vZKQ6Mfu5_2),.dout(w_dff_B_w5g9bPqK3_2),.clk(gclk));
	jdff dff_B_QoEsyjak3_2(.din(w_dff_B_w5g9bPqK3_2),.dout(w_dff_B_QoEsyjak3_2),.clk(gclk));
	jdff dff_B_CYpQHWUI5_2(.din(w_dff_B_QoEsyjak3_2),.dout(w_dff_B_CYpQHWUI5_2),.clk(gclk));
	jdff dff_B_7qTU7lys5_2(.din(w_dff_B_CYpQHWUI5_2),.dout(w_dff_B_7qTU7lys5_2),.clk(gclk));
	jdff dff_B_RQf5jV8H4_2(.din(w_dff_B_7qTU7lys5_2),.dout(w_dff_B_RQf5jV8H4_2),.clk(gclk));
	jdff dff_B_8O6FL66n5_2(.din(n1605),.dout(w_dff_B_8O6FL66n5_2),.clk(gclk));
	jdff dff_B_PWGUw7d86_1(.din(n1603),.dout(w_dff_B_PWGUw7d86_1),.clk(gclk));
	jdff dff_B_UjtCsIq95_2(.din(n1545),.dout(w_dff_B_UjtCsIq95_2),.clk(gclk));
	jdff dff_B_2FBFf7nb9_2(.din(w_dff_B_UjtCsIq95_2),.dout(w_dff_B_2FBFf7nb9_2),.clk(gclk));
	jdff dff_B_A3hZxBXW2_2(.din(w_dff_B_2FBFf7nb9_2),.dout(w_dff_B_A3hZxBXW2_2),.clk(gclk));
	jdff dff_B_IxevdxLc8_2(.din(w_dff_B_A3hZxBXW2_2),.dout(w_dff_B_IxevdxLc8_2),.clk(gclk));
	jdff dff_B_xQ3h8aY55_2(.din(w_dff_B_IxevdxLc8_2),.dout(w_dff_B_xQ3h8aY55_2),.clk(gclk));
	jdff dff_B_DkOgFsMV8_2(.din(w_dff_B_xQ3h8aY55_2),.dout(w_dff_B_DkOgFsMV8_2),.clk(gclk));
	jdff dff_B_fJBcM0qM6_2(.din(w_dff_B_DkOgFsMV8_2),.dout(w_dff_B_fJBcM0qM6_2),.clk(gclk));
	jdff dff_B_L7sjh2oX9_2(.din(w_dff_B_fJBcM0qM6_2),.dout(w_dff_B_L7sjh2oX9_2),.clk(gclk));
	jdff dff_B_IyDywO801_2(.din(w_dff_B_L7sjh2oX9_2),.dout(w_dff_B_IyDywO801_2),.clk(gclk));
	jdff dff_B_gE8xoJnz6_2(.din(w_dff_B_IyDywO801_2),.dout(w_dff_B_gE8xoJnz6_2),.clk(gclk));
	jdff dff_B_0TEbxsic0_2(.din(w_dff_B_gE8xoJnz6_2),.dout(w_dff_B_0TEbxsic0_2),.clk(gclk));
	jdff dff_B_o6TRXdeQ0_2(.din(w_dff_B_0TEbxsic0_2),.dout(w_dff_B_o6TRXdeQ0_2),.clk(gclk));
	jdff dff_B_p7CqJLlQ0_2(.din(w_dff_B_o6TRXdeQ0_2),.dout(w_dff_B_p7CqJLlQ0_2),.clk(gclk));
	jdff dff_B_ZneqRuYq6_2(.din(w_dff_B_p7CqJLlQ0_2),.dout(w_dff_B_ZneqRuYq6_2),.clk(gclk));
	jdff dff_B_45jqCXTn0_2(.din(w_dff_B_ZneqRuYq6_2),.dout(w_dff_B_45jqCXTn0_2),.clk(gclk));
	jdff dff_B_Qq7vmDBE6_2(.din(w_dff_B_45jqCXTn0_2),.dout(w_dff_B_Qq7vmDBE6_2),.clk(gclk));
	jdff dff_B_eA3vTREJ7_2(.din(w_dff_B_Qq7vmDBE6_2),.dout(w_dff_B_eA3vTREJ7_2),.clk(gclk));
	jdff dff_B_KcisPGXK9_2(.din(w_dff_B_eA3vTREJ7_2),.dout(w_dff_B_KcisPGXK9_2),.clk(gclk));
	jdff dff_B_WEDuEVWN1_2(.din(w_dff_B_KcisPGXK9_2),.dout(w_dff_B_WEDuEVWN1_2),.clk(gclk));
	jdff dff_B_plOaHfpE7_2(.din(w_dff_B_WEDuEVWN1_2),.dout(w_dff_B_plOaHfpE7_2),.clk(gclk));
	jdff dff_B_emkmWjAt8_2(.din(w_dff_B_plOaHfpE7_2),.dout(w_dff_B_emkmWjAt8_2),.clk(gclk));
	jdff dff_B_qvuQ9Hzb7_2(.din(w_dff_B_emkmWjAt8_2),.dout(w_dff_B_qvuQ9Hzb7_2),.clk(gclk));
	jdff dff_B_5Fzxgran2_2(.din(w_dff_B_qvuQ9Hzb7_2),.dout(w_dff_B_5Fzxgran2_2),.clk(gclk));
	jdff dff_B_dP9OO4NJ2_2(.din(w_dff_B_5Fzxgran2_2),.dout(w_dff_B_dP9OO4NJ2_2),.clk(gclk));
	jdff dff_B_1CLlZGws5_2(.din(w_dff_B_dP9OO4NJ2_2),.dout(w_dff_B_1CLlZGws5_2),.clk(gclk));
	jdff dff_B_bq2q6p1G5_2(.din(w_dff_B_1CLlZGws5_2),.dout(w_dff_B_bq2q6p1G5_2),.clk(gclk));
	jdff dff_B_pr619eye4_2(.din(w_dff_B_bq2q6p1G5_2),.dout(w_dff_B_pr619eye4_2),.clk(gclk));
	jdff dff_B_Hpxyhvh51_2(.din(w_dff_B_pr619eye4_2),.dout(w_dff_B_Hpxyhvh51_2),.clk(gclk));
	jdff dff_B_gbTO50EO7_2(.din(w_dff_B_Hpxyhvh51_2),.dout(w_dff_B_gbTO50EO7_2),.clk(gclk));
	jdff dff_B_jIfg9ag48_2(.din(w_dff_B_gbTO50EO7_2),.dout(w_dff_B_jIfg9ag48_2),.clk(gclk));
	jdff dff_B_NCdnn3Yy6_2(.din(w_dff_B_jIfg9ag48_2),.dout(w_dff_B_NCdnn3Yy6_2),.clk(gclk));
	jdff dff_B_yQ8ZbIFE5_2(.din(w_dff_B_NCdnn3Yy6_2),.dout(w_dff_B_yQ8ZbIFE5_2),.clk(gclk));
	jdff dff_B_KQnXlsq47_2(.din(w_dff_B_yQ8ZbIFE5_2),.dout(w_dff_B_KQnXlsq47_2),.clk(gclk));
	jdff dff_B_VYo8NXq32_2(.din(w_dff_B_KQnXlsq47_2),.dout(w_dff_B_VYo8NXq32_2),.clk(gclk));
	jdff dff_B_jetdDKut5_2(.din(w_dff_B_VYo8NXq32_2),.dout(w_dff_B_jetdDKut5_2),.clk(gclk));
	jdff dff_B_hodL1qM27_2(.din(w_dff_B_jetdDKut5_2),.dout(w_dff_B_hodL1qM27_2),.clk(gclk));
	jdff dff_B_weh610iE4_2(.din(w_dff_B_hodL1qM27_2),.dout(w_dff_B_weh610iE4_2),.clk(gclk));
	jdff dff_B_ryjsFclc7_2(.din(w_dff_B_weh610iE4_2),.dout(w_dff_B_ryjsFclc7_2),.clk(gclk));
	jdff dff_B_TkxqROVW5_1(.din(n1546),.dout(w_dff_B_TkxqROVW5_1),.clk(gclk));
	jdff dff_B_ILYBq7oC4_2(.din(n1481),.dout(w_dff_B_ILYBq7oC4_2),.clk(gclk));
	jdff dff_B_FhiqZvdu7_2(.din(w_dff_B_ILYBq7oC4_2),.dout(w_dff_B_FhiqZvdu7_2),.clk(gclk));
	jdff dff_B_jRvyvnNH2_2(.din(w_dff_B_FhiqZvdu7_2),.dout(w_dff_B_jRvyvnNH2_2),.clk(gclk));
	jdff dff_B_8SniH8HP9_2(.din(w_dff_B_jRvyvnNH2_2),.dout(w_dff_B_8SniH8HP9_2),.clk(gclk));
	jdff dff_B_7a3dHNp73_2(.din(w_dff_B_8SniH8HP9_2),.dout(w_dff_B_7a3dHNp73_2),.clk(gclk));
	jdff dff_B_qOPBmmdJ9_2(.din(w_dff_B_7a3dHNp73_2),.dout(w_dff_B_qOPBmmdJ9_2),.clk(gclk));
	jdff dff_B_hqkURLnP4_2(.din(w_dff_B_qOPBmmdJ9_2),.dout(w_dff_B_hqkURLnP4_2),.clk(gclk));
	jdff dff_B_dYMx2zw50_2(.din(w_dff_B_hqkURLnP4_2),.dout(w_dff_B_dYMx2zw50_2),.clk(gclk));
	jdff dff_B_e8kVhg791_2(.din(w_dff_B_dYMx2zw50_2),.dout(w_dff_B_e8kVhg791_2),.clk(gclk));
	jdff dff_B_F7tCiPu11_2(.din(w_dff_B_e8kVhg791_2),.dout(w_dff_B_F7tCiPu11_2),.clk(gclk));
	jdff dff_B_SjbfP5Z02_2(.din(w_dff_B_F7tCiPu11_2),.dout(w_dff_B_SjbfP5Z02_2),.clk(gclk));
	jdff dff_B_xX9DT0jS3_2(.din(w_dff_B_SjbfP5Z02_2),.dout(w_dff_B_xX9DT0jS3_2),.clk(gclk));
	jdff dff_B_pU3K24Qg8_2(.din(w_dff_B_xX9DT0jS3_2),.dout(w_dff_B_pU3K24Qg8_2),.clk(gclk));
	jdff dff_B_97WXnysl8_2(.din(w_dff_B_pU3K24Qg8_2),.dout(w_dff_B_97WXnysl8_2),.clk(gclk));
	jdff dff_B_wsh8o2237_2(.din(w_dff_B_97WXnysl8_2),.dout(w_dff_B_wsh8o2237_2),.clk(gclk));
	jdff dff_B_E3vO13B00_2(.din(w_dff_B_wsh8o2237_2),.dout(w_dff_B_E3vO13B00_2),.clk(gclk));
	jdff dff_B_BwToRSrO5_2(.din(w_dff_B_E3vO13B00_2),.dout(w_dff_B_BwToRSrO5_2),.clk(gclk));
	jdff dff_B_ta7y8tgH6_2(.din(w_dff_B_BwToRSrO5_2),.dout(w_dff_B_ta7y8tgH6_2),.clk(gclk));
	jdff dff_B_4dE50Gwp8_2(.din(w_dff_B_ta7y8tgH6_2),.dout(w_dff_B_4dE50Gwp8_2),.clk(gclk));
	jdff dff_B_4466LlwD0_2(.din(w_dff_B_4dE50Gwp8_2),.dout(w_dff_B_4466LlwD0_2),.clk(gclk));
	jdff dff_B_MXoQ7O9y8_2(.din(w_dff_B_4466LlwD0_2),.dout(w_dff_B_MXoQ7O9y8_2),.clk(gclk));
	jdff dff_B_D2wU16SM2_2(.din(w_dff_B_MXoQ7O9y8_2),.dout(w_dff_B_D2wU16SM2_2),.clk(gclk));
	jdff dff_B_TRmMkrUB4_2(.din(w_dff_B_D2wU16SM2_2),.dout(w_dff_B_TRmMkrUB4_2),.clk(gclk));
	jdff dff_B_wJ2AoZmT2_2(.din(w_dff_B_TRmMkrUB4_2),.dout(w_dff_B_wJ2AoZmT2_2),.clk(gclk));
	jdff dff_B_rJkbEKeZ2_2(.din(w_dff_B_wJ2AoZmT2_2),.dout(w_dff_B_rJkbEKeZ2_2),.clk(gclk));
	jdff dff_B_QiWiEkcq3_2(.din(w_dff_B_rJkbEKeZ2_2),.dout(w_dff_B_QiWiEkcq3_2),.clk(gclk));
	jdff dff_B_nz7xI0Ml6_2(.din(w_dff_B_QiWiEkcq3_2),.dout(w_dff_B_nz7xI0Ml6_2),.clk(gclk));
	jdff dff_B_PO2f7dKZ3_2(.din(w_dff_B_nz7xI0Ml6_2),.dout(w_dff_B_PO2f7dKZ3_2),.clk(gclk));
	jdff dff_B_cg2pk6Qf3_2(.din(w_dff_B_PO2f7dKZ3_2),.dout(w_dff_B_cg2pk6Qf3_2),.clk(gclk));
	jdff dff_B_7VfQK97E2_2(.din(w_dff_B_cg2pk6Qf3_2),.dout(w_dff_B_7VfQK97E2_2),.clk(gclk));
	jdff dff_B_0x1OAe0j3_2(.din(w_dff_B_7VfQK97E2_2),.dout(w_dff_B_0x1OAe0j3_2),.clk(gclk));
	jdff dff_B_77bUs3HG7_2(.din(w_dff_B_0x1OAe0j3_2),.dout(w_dff_B_77bUs3HG7_2),.clk(gclk));
	jdff dff_B_BikqO5xy9_2(.din(w_dff_B_77bUs3HG7_2),.dout(w_dff_B_BikqO5xy9_2),.clk(gclk));
	jdff dff_B_FUvRPWGM6_2(.din(w_dff_B_BikqO5xy9_2),.dout(w_dff_B_FUvRPWGM6_2),.clk(gclk));
	jdff dff_B_7kyonYWH5_2(.din(w_dff_B_FUvRPWGM6_2),.dout(w_dff_B_7kyonYWH5_2),.clk(gclk));
	jdff dff_B_Lxj1A7jA7_2(.din(n1513),.dout(w_dff_B_Lxj1A7jA7_2),.clk(gclk));
	jdff dff_B_hpSnetn01_1(.din(n1482),.dout(w_dff_B_hpSnetn01_1),.clk(gclk));
	jdff dff_B_WHa8wRvB1_2(.din(n1410),.dout(w_dff_B_WHa8wRvB1_2),.clk(gclk));
	jdff dff_B_49e0OhMy7_2(.din(w_dff_B_WHa8wRvB1_2),.dout(w_dff_B_49e0OhMy7_2),.clk(gclk));
	jdff dff_B_OhDGhI9z1_2(.din(w_dff_B_49e0OhMy7_2),.dout(w_dff_B_OhDGhI9z1_2),.clk(gclk));
	jdff dff_B_HnJpM4PZ3_2(.din(w_dff_B_OhDGhI9z1_2),.dout(w_dff_B_HnJpM4PZ3_2),.clk(gclk));
	jdff dff_B_y9xdCoen3_2(.din(w_dff_B_HnJpM4PZ3_2),.dout(w_dff_B_y9xdCoen3_2),.clk(gclk));
	jdff dff_B_TxxhFT373_2(.din(w_dff_B_y9xdCoen3_2),.dout(w_dff_B_TxxhFT373_2),.clk(gclk));
	jdff dff_B_FqhYvdZG8_2(.din(w_dff_B_TxxhFT373_2),.dout(w_dff_B_FqhYvdZG8_2),.clk(gclk));
	jdff dff_B_fRqZcGXX4_2(.din(w_dff_B_FqhYvdZG8_2),.dout(w_dff_B_fRqZcGXX4_2),.clk(gclk));
	jdff dff_B_iNo8s8U23_2(.din(w_dff_B_fRqZcGXX4_2),.dout(w_dff_B_iNo8s8U23_2),.clk(gclk));
	jdff dff_B_tikmd1Ny1_2(.din(w_dff_B_iNo8s8U23_2),.dout(w_dff_B_tikmd1Ny1_2),.clk(gclk));
	jdff dff_B_ikuEt39o1_2(.din(w_dff_B_tikmd1Ny1_2),.dout(w_dff_B_ikuEt39o1_2),.clk(gclk));
	jdff dff_B_O9CkpP3U1_2(.din(w_dff_B_ikuEt39o1_2),.dout(w_dff_B_O9CkpP3U1_2),.clk(gclk));
	jdff dff_B_r82IGXdZ6_2(.din(w_dff_B_O9CkpP3U1_2),.dout(w_dff_B_r82IGXdZ6_2),.clk(gclk));
	jdff dff_B_3grm17AD7_2(.din(w_dff_B_r82IGXdZ6_2),.dout(w_dff_B_3grm17AD7_2),.clk(gclk));
	jdff dff_B_xyafewkp7_2(.din(w_dff_B_3grm17AD7_2),.dout(w_dff_B_xyafewkp7_2),.clk(gclk));
	jdff dff_B_e4RXbdMU0_2(.din(w_dff_B_xyafewkp7_2),.dout(w_dff_B_e4RXbdMU0_2),.clk(gclk));
	jdff dff_B_I5hyxxs73_2(.din(w_dff_B_e4RXbdMU0_2),.dout(w_dff_B_I5hyxxs73_2),.clk(gclk));
	jdff dff_B_wqi8rNtI1_2(.din(w_dff_B_I5hyxxs73_2),.dout(w_dff_B_wqi8rNtI1_2),.clk(gclk));
	jdff dff_B_G2C80Fdd2_2(.din(w_dff_B_wqi8rNtI1_2),.dout(w_dff_B_G2C80Fdd2_2),.clk(gclk));
	jdff dff_B_oD2Hcv5r4_2(.din(w_dff_B_G2C80Fdd2_2),.dout(w_dff_B_oD2Hcv5r4_2),.clk(gclk));
	jdff dff_B_fog9XP5O2_2(.din(w_dff_B_oD2Hcv5r4_2),.dout(w_dff_B_fog9XP5O2_2),.clk(gclk));
	jdff dff_B_5HXJhtaF3_2(.din(w_dff_B_fog9XP5O2_2),.dout(w_dff_B_5HXJhtaF3_2),.clk(gclk));
	jdff dff_B_0NoRYcOp6_2(.din(w_dff_B_5HXJhtaF3_2),.dout(w_dff_B_0NoRYcOp6_2),.clk(gclk));
	jdff dff_B_btDNh6wR3_2(.din(w_dff_B_0NoRYcOp6_2),.dout(w_dff_B_btDNh6wR3_2),.clk(gclk));
	jdff dff_B_d87YSAsi0_2(.din(w_dff_B_btDNh6wR3_2),.dout(w_dff_B_d87YSAsi0_2),.clk(gclk));
	jdff dff_B_DGq3LQSS9_2(.din(w_dff_B_d87YSAsi0_2),.dout(w_dff_B_DGq3LQSS9_2),.clk(gclk));
	jdff dff_B_8mcX23te9_2(.din(w_dff_B_DGq3LQSS9_2),.dout(w_dff_B_8mcX23te9_2),.clk(gclk));
	jdff dff_B_FrAHjZAT7_2(.din(w_dff_B_8mcX23te9_2),.dout(w_dff_B_FrAHjZAT7_2),.clk(gclk));
	jdff dff_B_f3ceJS240_2(.din(w_dff_B_FrAHjZAT7_2),.dout(w_dff_B_f3ceJS240_2),.clk(gclk));
	jdff dff_B_nPrlUkPQ9_2(.din(w_dff_B_f3ceJS240_2),.dout(w_dff_B_nPrlUkPQ9_2),.clk(gclk));
	jdff dff_B_YkPAgCZk6_2(.din(w_dff_B_nPrlUkPQ9_2),.dout(w_dff_B_YkPAgCZk6_2),.clk(gclk));
	jdff dff_B_Hlxo0DKL6_2(.din(w_dff_B_YkPAgCZk6_2),.dout(w_dff_B_Hlxo0DKL6_2),.clk(gclk));
	jdff dff_B_tqh4Egzt0_2(.din(n1442),.dout(w_dff_B_tqh4Egzt0_2),.clk(gclk));
	jdff dff_B_AGOGhga26_1(.din(n1411),.dout(w_dff_B_AGOGhga26_1),.clk(gclk));
	jdff dff_B_iKkpZuvh2_2(.din(n1332),.dout(w_dff_B_iKkpZuvh2_2),.clk(gclk));
	jdff dff_B_d2JHRYAE6_2(.din(w_dff_B_iKkpZuvh2_2),.dout(w_dff_B_d2JHRYAE6_2),.clk(gclk));
	jdff dff_B_dQVzrfqs2_2(.din(w_dff_B_d2JHRYAE6_2),.dout(w_dff_B_dQVzrfqs2_2),.clk(gclk));
	jdff dff_B_Y2i3sSXZ1_2(.din(w_dff_B_dQVzrfqs2_2),.dout(w_dff_B_Y2i3sSXZ1_2),.clk(gclk));
	jdff dff_B_hoj4EpN59_2(.din(w_dff_B_Y2i3sSXZ1_2),.dout(w_dff_B_hoj4EpN59_2),.clk(gclk));
	jdff dff_B_itmNrREO9_2(.din(w_dff_B_hoj4EpN59_2),.dout(w_dff_B_itmNrREO9_2),.clk(gclk));
	jdff dff_B_f8KWNAef2_2(.din(w_dff_B_itmNrREO9_2),.dout(w_dff_B_f8KWNAef2_2),.clk(gclk));
	jdff dff_B_JUkqhfsD7_2(.din(w_dff_B_f8KWNAef2_2),.dout(w_dff_B_JUkqhfsD7_2),.clk(gclk));
	jdff dff_B_W1exKHoF5_2(.din(w_dff_B_JUkqhfsD7_2),.dout(w_dff_B_W1exKHoF5_2),.clk(gclk));
	jdff dff_B_dnQuA9eV7_2(.din(w_dff_B_W1exKHoF5_2),.dout(w_dff_B_dnQuA9eV7_2),.clk(gclk));
	jdff dff_B_OYrOFMKU8_2(.din(w_dff_B_dnQuA9eV7_2),.dout(w_dff_B_OYrOFMKU8_2),.clk(gclk));
	jdff dff_B_ru2tzxYP9_2(.din(w_dff_B_OYrOFMKU8_2),.dout(w_dff_B_ru2tzxYP9_2),.clk(gclk));
	jdff dff_B_q2WK9FCg1_2(.din(w_dff_B_ru2tzxYP9_2),.dout(w_dff_B_q2WK9FCg1_2),.clk(gclk));
	jdff dff_B_TRrY3cb73_2(.din(w_dff_B_q2WK9FCg1_2),.dout(w_dff_B_TRrY3cb73_2),.clk(gclk));
	jdff dff_B_L2hbt7Qv3_2(.din(w_dff_B_TRrY3cb73_2),.dout(w_dff_B_L2hbt7Qv3_2),.clk(gclk));
	jdff dff_B_bomolWtn5_2(.din(w_dff_B_L2hbt7Qv3_2),.dout(w_dff_B_bomolWtn5_2),.clk(gclk));
	jdff dff_B_ExVtAqnd6_2(.din(w_dff_B_bomolWtn5_2),.dout(w_dff_B_ExVtAqnd6_2),.clk(gclk));
	jdff dff_B_K8NCccEu6_2(.din(w_dff_B_ExVtAqnd6_2),.dout(w_dff_B_K8NCccEu6_2),.clk(gclk));
	jdff dff_B_eZaVu03u2_2(.din(w_dff_B_K8NCccEu6_2),.dout(w_dff_B_eZaVu03u2_2),.clk(gclk));
	jdff dff_B_WWe23Agw5_2(.din(w_dff_B_eZaVu03u2_2),.dout(w_dff_B_WWe23Agw5_2),.clk(gclk));
	jdff dff_B_6UxDvB6k9_2(.din(w_dff_B_WWe23Agw5_2),.dout(w_dff_B_6UxDvB6k9_2),.clk(gclk));
	jdff dff_B_9Cqae6962_2(.din(w_dff_B_6UxDvB6k9_2),.dout(w_dff_B_9Cqae6962_2),.clk(gclk));
	jdff dff_B_atxFZfKO9_2(.din(w_dff_B_9Cqae6962_2),.dout(w_dff_B_atxFZfKO9_2),.clk(gclk));
	jdff dff_B_BTNP1cHa8_2(.din(w_dff_B_atxFZfKO9_2),.dout(w_dff_B_BTNP1cHa8_2),.clk(gclk));
	jdff dff_B_JuGvrBSW0_2(.din(w_dff_B_BTNP1cHa8_2),.dout(w_dff_B_JuGvrBSW0_2),.clk(gclk));
	jdff dff_B_rj9OZnPs9_2(.din(w_dff_B_JuGvrBSW0_2),.dout(w_dff_B_rj9OZnPs9_2),.clk(gclk));
	jdff dff_B_Rwy09Gx62_2(.din(w_dff_B_rj9OZnPs9_2),.dout(w_dff_B_Rwy09Gx62_2),.clk(gclk));
	jdff dff_B_35y5uoGK4_2(.din(w_dff_B_Rwy09Gx62_2),.dout(w_dff_B_35y5uoGK4_2),.clk(gclk));
	jdff dff_B_efYzMPz54_2(.din(w_dff_B_35y5uoGK4_2),.dout(w_dff_B_efYzMPz54_2),.clk(gclk));
	jdff dff_B_SkDVNICh2_2(.din(n1364),.dout(w_dff_B_SkDVNICh2_2),.clk(gclk));
	jdff dff_B_aLxXaBkb0_1(.din(n1333),.dout(w_dff_B_aLxXaBkb0_1),.clk(gclk));
	jdff dff_B_9vvyijU41_2(.din(n1247),.dout(w_dff_B_9vvyijU41_2),.clk(gclk));
	jdff dff_B_Jc3wGxe92_2(.din(w_dff_B_9vvyijU41_2),.dout(w_dff_B_Jc3wGxe92_2),.clk(gclk));
	jdff dff_B_uQ6ZivpW7_2(.din(w_dff_B_Jc3wGxe92_2),.dout(w_dff_B_uQ6ZivpW7_2),.clk(gclk));
	jdff dff_B_PDOuhlgu0_2(.din(w_dff_B_uQ6ZivpW7_2),.dout(w_dff_B_PDOuhlgu0_2),.clk(gclk));
	jdff dff_B_NZfyBnrl7_2(.din(w_dff_B_PDOuhlgu0_2),.dout(w_dff_B_NZfyBnrl7_2),.clk(gclk));
	jdff dff_B_58NyR2xG8_2(.din(w_dff_B_NZfyBnrl7_2),.dout(w_dff_B_58NyR2xG8_2),.clk(gclk));
	jdff dff_B_QEhTsO0T2_2(.din(w_dff_B_58NyR2xG8_2),.dout(w_dff_B_QEhTsO0T2_2),.clk(gclk));
	jdff dff_B_iLLBdhIE1_2(.din(w_dff_B_QEhTsO0T2_2),.dout(w_dff_B_iLLBdhIE1_2),.clk(gclk));
	jdff dff_B_2ziVN1Cx5_2(.din(w_dff_B_iLLBdhIE1_2),.dout(w_dff_B_2ziVN1Cx5_2),.clk(gclk));
	jdff dff_B_XGkMAYdB5_2(.din(w_dff_B_2ziVN1Cx5_2),.dout(w_dff_B_XGkMAYdB5_2),.clk(gclk));
	jdff dff_B_AORQPlV59_2(.din(w_dff_B_XGkMAYdB5_2),.dout(w_dff_B_AORQPlV59_2),.clk(gclk));
	jdff dff_B_dzu6utUz2_2(.din(w_dff_B_AORQPlV59_2),.dout(w_dff_B_dzu6utUz2_2),.clk(gclk));
	jdff dff_B_9ObBPCfB6_2(.din(w_dff_B_dzu6utUz2_2),.dout(w_dff_B_9ObBPCfB6_2),.clk(gclk));
	jdff dff_B_kVeQ6qku3_2(.din(w_dff_B_9ObBPCfB6_2),.dout(w_dff_B_kVeQ6qku3_2),.clk(gclk));
	jdff dff_B_6coCRPyg8_2(.din(w_dff_B_kVeQ6qku3_2),.dout(w_dff_B_6coCRPyg8_2),.clk(gclk));
	jdff dff_B_dAI4pKjT4_2(.din(w_dff_B_6coCRPyg8_2),.dout(w_dff_B_dAI4pKjT4_2),.clk(gclk));
	jdff dff_B_J4mpgpSg0_2(.din(w_dff_B_dAI4pKjT4_2),.dout(w_dff_B_J4mpgpSg0_2),.clk(gclk));
	jdff dff_B_PDNZTc5s5_2(.din(w_dff_B_J4mpgpSg0_2),.dout(w_dff_B_PDNZTc5s5_2),.clk(gclk));
	jdff dff_B_zAeVcSGl7_2(.din(w_dff_B_PDNZTc5s5_2),.dout(w_dff_B_zAeVcSGl7_2),.clk(gclk));
	jdff dff_B_3hbZyOdU6_2(.din(w_dff_B_zAeVcSGl7_2),.dout(w_dff_B_3hbZyOdU6_2),.clk(gclk));
	jdff dff_B_CUOsoGQR6_2(.din(w_dff_B_3hbZyOdU6_2),.dout(w_dff_B_CUOsoGQR6_2),.clk(gclk));
	jdff dff_B_RPwjE7CU8_2(.din(w_dff_B_CUOsoGQR6_2),.dout(w_dff_B_RPwjE7CU8_2),.clk(gclk));
	jdff dff_B_aNEZFJig2_2(.din(w_dff_B_RPwjE7CU8_2),.dout(w_dff_B_aNEZFJig2_2),.clk(gclk));
	jdff dff_B_nnEA6jhf4_2(.din(w_dff_B_aNEZFJig2_2),.dout(w_dff_B_nnEA6jhf4_2),.clk(gclk));
	jdff dff_B_2FugCIN58_2(.din(w_dff_B_nnEA6jhf4_2),.dout(w_dff_B_2FugCIN58_2),.clk(gclk));
	jdff dff_B_Z2H3KzTz3_2(.din(w_dff_B_2FugCIN58_2),.dout(w_dff_B_Z2H3KzTz3_2),.clk(gclk));
	jdff dff_B_c3ouuaHN5_2(.din(n1279),.dout(w_dff_B_c3ouuaHN5_2),.clk(gclk));
	jdff dff_B_C3FFnonp9_1(.din(n1248),.dout(w_dff_B_C3FFnonp9_1),.clk(gclk));
	jdff dff_B_NMSto3Mm2_2(.din(n1156),.dout(w_dff_B_NMSto3Mm2_2),.clk(gclk));
	jdff dff_B_I1LkqqKz2_2(.din(w_dff_B_NMSto3Mm2_2),.dout(w_dff_B_I1LkqqKz2_2),.clk(gclk));
	jdff dff_B_GxBhb5m90_2(.din(w_dff_B_I1LkqqKz2_2),.dout(w_dff_B_GxBhb5m90_2),.clk(gclk));
	jdff dff_B_LkBNXGK29_2(.din(w_dff_B_GxBhb5m90_2),.dout(w_dff_B_LkBNXGK29_2),.clk(gclk));
	jdff dff_B_sLmW6l7F5_2(.din(w_dff_B_LkBNXGK29_2),.dout(w_dff_B_sLmW6l7F5_2),.clk(gclk));
	jdff dff_B_CF4SF6d23_2(.din(w_dff_B_sLmW6l7F5_2),.dout(w_dff_B_CF4SF6d23_2),.clk(gclk));
	jdff dff_B_RRYrR1jQ7_2(.din(w_dff_B_CF4SF6d23_2),.dout(w_dff_B_RRYrR1jQ7_2),.clk(gclk));
	jdff dff_B_DHizh3n91_2(.din(w_dff_B_RRYrR1jQ7_2),.dout(w_dff_B_DHizh3n91_2),.clk(gclk));
	jdff dff_B_9q7jPIU23_2(.din(w_dff_B_DHizh3n91_2),.dout(w_dff_B_9q7jPIU23_2),.clk(gclk));
	jdff dff_B_smlRYZrp1_2(.din(w_dff_B_9q7jPIU23_2),.dout(w_dff_B_smlRYZrp1_2),.clk(gclk));
	jdff dff_B_jKewHi7F5_2(.din(w_dff_B_smlRYZrp1_2),.dout(w_dff_B_jKewHi7F5_2),.clk(gclk));
	jdff dff_B_Zx0BdT2J9_2(.din(w_dff_B_jKewHi7F5_2),.dout(w_dff_B_Zx0BdT2J9_2),.clk(gclk));
	jdff dff_B_GwqkwY8C5_2(.din(w_dff_B_Zx0BdT2J9_2),.dout(w_dff_B_GwqkwY8C5_2),.clk(gclk));
	jdff dff_B_qMg2IR714_2(.din(w_dff_B_GwqkwY8C5_2),.dout(w_dff_B_qMg2IR714_2),.clk(gclk));
	jdff dff_B_8gFIau1v5_2(.din(w_dff_B_qMg2IR714_2),.dout(w_dff_B_8gFIau1v5_2),.clk(gclk));
	jdff dff_B_0RWu5RWr2_2(.din(w_dff_B_8gFIau1v5_2),.dout(w_dff_B_0RWu5RWr2_2),.clk(gclk));
	jdff dff_B_6YTeBN2C2_2(.din(w_dff_B_0RWu5RWr2_2),.dout(w_dff_B_6YTeBN2C2_2),.clk(gclk));
	jdff dff_B_VDewpwzq9_2(.din(w_dff_B_6YTeBN2C2_2),.dout(w_dff_B_VDewpwzq9_2),.clk(gclk));
	jdff dff_B_qqZ9UZjH3_2(.din(w_dff_B_VDewpwzq9_2),.dout(w_dff_B_qqZ9UZjH3_2),.clk(gclk));
	jdff dff_B_1bpYPDPy7_2(.din(w_dff_B_qqZ9UZjH3_2),.dout(w_dff_B_1bpYPDPy7_2),.clk(gclk));
	jdff dff_B_mbKxSyET4_2(.din(w_dff_B_1bpYPDPy7_2),.dout(w_dff_B_mbKxSyET4_2),.clk(gclk));
	jdff dff_B_zPTss1mL8_2(.din(w_dff_B_mbKxSyET4_2),.dout(w_dff_B_zPTss1mL8_2),.clk(gclk));
	jdff dff_B_fFzEiE7X7_2(.din(w_dff_B_zPTss1mL8_2),.dout(w_dff_B_fFzEiE7X7_2),.clk(gclk));
	jdff dff_B_gVfB6OuJ0_2(.din(n1188),.dout(w_dff_B_gVfB6OuJ0_2),.clk(gclk));
	jdff dff_B_6uAOIO527_1(.din(n1157),.dout(w_dff_B_6uAOIO527_1),.clk(gclk));
	jdff dff_B_Og1E3fEo7_2(.din(n1058),.dout(w_dff_B_Og1E3fEo7_2),.clk(gclk));
	jdff dff_B_p1K4nSmB2_2(.din(w_dff_B_Og1E3fEo7_2),.dout(w_dff_B_p1K4nSmB2_2),.clk(gclk));
	jdff dff_B_VtvaCsJW8_2(.din(w_dff_B_p1K4nSmB2_2),.dout(w_dff_B_VtvaCsJW8_2),.clk(gclk));
	jdff dff_B_GdcaahH54_2(.din(w_dff_B_VtvaCsJW8_2),.dout(w_dff_B_GdcaahH54_2),.clk(gclk));
	jdff dff_B_cNYtdx9M4_2(.din(w_dff_B_GdcaahH54_2),.dout(w_dff_B_cNYtdx9M4_2),.clk(gclk));
	jdff dff_B_lTAmXAox1_2(.din(w_dff_B_cNYtdx9M4_2),.dout(w_dff_B_lTAmXAox1_2),.clk(gclk));
	jdff dff_B_MrIi5FUd4_2(.din(w_dff_B_lTAmXAox1_2),.dout(w_dff_B_MrIi5FUd4_2),.clk(gclk));
	jdff dff_B_shbaHQVl7_2(.din(w_dff_B_MrIi5FUd4_2),.dout(w_dff_B_shbaHQVl7_2),.clk(gclk));
	jdff dff_B_kbqHaiSe3_2(.din(w_dff_B_shbaHQVl7_2),.dout(w_dff_B_kbqHaiSe3_2),.clk(gclk));
	jdff dff_B_UAKDsih58_2(.din(w_dff_B_kbqHaiSe3_2),.dout(w_dff_B_UAKDsih58_2),.clk(gclk));
	jdff dff_B_XPrKZe582_2(.din(w_dff_B_UAKDsih58_2),.dout(w_dff_B_XPrKZe582_2),.clk(gclk));
	jdff dff_B_XTgMDWXg5_2(.din(w_dff_B_XPrKZe582_2),.dout(w_dff_B_XTgMDWXg5_2),.clk(gclk));
	jdff dff_B_EBQ3XWoe6_2(.din(w_dff_B_XTgMDWXg5_2),.dout(w_dff_B_EBQ3XWoe6_2),.clk(gclk));
	jdff dff_B_ufxvtP217_2(.din(w_dff_B_EBQ3XWoe6_2),.dout(w_dff_B_ufxvtP217_2),.clk(gclk));
	jdff dff_B_zMjPcx6u5_2(.din(w_dff_B_ufxvtP217_2),.dout(w_dff_B_zMjPcx6u5_2),.clk(gclk));
	jdff dff_B_kFRRaUWn9_2(.din(w_dff_B_zMjPcx6u5_2),.dout(w_dff_B_kFRRaUWn9_2),.clk(gclk));
	jdff dff_B_QCFiVIu31_2(.din(w_dff_B_kFRRaUWn9_2),.dout(w_dff_B_QCFiVIu31_2),.clk(gclk));
	jdff dff_B_UkwlhGwZ4_2(.din(w_dff_B_QCFiVIu31_2),.dout(w_dff_B_UkwlhGwZ4_2),.clk(gclk));
	jdff dff_B_4ijmjSmD2_2(.din(w_dff_B_UkwlhGwZ4_2),.dout(w_dff_B_4ijmjSmD2_2),.clk(gclk));
	jdff dff_B_aeK2CoD29_2(.din(w_dff_B_4ijmjSmD2_2),.dout(w_dff_B_aeK2CoD29_2),.clk(gclk));
	jdff dff_B_642m3ZPH9_2(.din(n1089),.dout(w_dff_B_642m3ZPH9_2),.clk(gclk));
	jdff dff_B_V7jV1Ext4_1(.din(n1059),.dout(w_dff_B_V7jV1Ext4_1),.clk(gclk));
	jdff dff_B_H0eY1vCP7_2(.din(n959),.dout(w_dff_B_H0eY1vCP7_2),.clk(gclk));
	jdff dff_B_kGDEyA688_2(.din(w_dff_B_H0eY1vCP7_2),.dout(w_dff_B_kGDEyA688_2),.clk(gclk));
	jdff dff_B_7midFWKD9_2(.din(w_dff_B_kGDEyA688_2),.dout(w_dff_B_7midFWKD9_2),.clk(gclk));
	jdff dff_B_7RTBT8P87_2(.din(w_dff_B_7midFWKD9_2),.dout(w_dff_B_7RTBT8P87_2),.clk(gclk));
	jdff dff_B_O192w7cy9_2(.din(w_dff_B_7RTBT8P87_2),.dout(w_dff_B_O192w7cy9_2),.clk(gclk));
	jdff dff_B_MfCgHR8F5_2(.din(w_dff_B_O192w7cy9_2),.dout(w_dff_B_MfCgHR8F5_2),.clk(gclk));
	jdff dff_B_5xHweeaR5_2(.din(w_dff_B_MfCgHR8F5_2),.dout(w_dff_B_5xHweeaR5_2),.clk(gclk));
	jdff dff_B_UWykl13E0_2(.din(w_dff_B_5xHweeaR5_2),.dout(w_dff_B_UWykl13E0_2),.clk(gclk));
	jdff dff_B_S25beSWm8_2(.din(w_dff_B_UWykl13E0_2),.dout(w_dff_B_S25beSWm8_2),.clk(gclk));
	jdff dff_B_2ATTapyC3_2(.din(w_dff_B_S25beSWm8_2),.dout(w_dff_B_2ATTapyC3_2),.clk(gclk));
	jdff dff_B_vwNcG6CI9_2(.din(w_dff_B_2ATTapyC3_2),.dout(w_dff_B_vwNcG6CI9_2),.clk(gclk));
	jdff dff_B_fBp0edJv9_2(.din(w_dff_B_vwNcG6CI9_2),.dout(w_dff_B_fBp0edJv9_2),.clk(gclk));
	jdff dff_B_Zp6cFr067_2(.din(w_dff_B_fBp0edJv9_2),.dout(w_dff_B_Zp6cFr067_2),.clk(gclk));
	jdff dff_B_jIB7rih82_2(.din(w_dff_B_Zp6cFr067_2),.dout(w_dff_B_jIB7rih82_2),.clk(gclk));
	jdff dff_B_JEI8yRGU7_2(.din(w_dff_B_jIB7rih82_2),.dout(w_dff_B_JEI8yRGU7_2),.clk(gclk));
	jdff dff_B_Z4HN1GRr4_2(.din(w_dff_B_JEI8yRGU7_2),.dout(w_dff_B_Z4HN1GRr4_2),.clk(gclk));
	jdff dff_B_d7RAo6mC7_2(.din(w_dff_B_Z4HN1GRr4_2),.dout(w_dff_B_d7RAo6mC7_2),.clk(gclk));
	jdff dff_B_6ZVNhIwl0_2(.din(n990),.dout(w_dff_B_6ZVNhIwl0_2),.clk(gclk));
	jdff dff_B_hXdk3x3M0_1(.din(n960),.dout(w_dff_B_hXdk3x3M0_1),.clk(gclk));
	jdff dff_B_XJQ9mYHf9_2(.din(n857),.dout(w_dff_B_XJQ9mYHf9_2),.clk(gclk));
	jdff dff_B_nnmoNH6T1_2(.din(w_dff_B_XJQ9mYHf9_2),.dout(w_dff_B_nnmoNH6T1_2),.clk(gclk));
	jdff dff_B_qwE0HqvV7_2(.din(w_dff_B_nnmoNH6T1_2),.dout(w_dff_B_qwE0HqvV7_2),.clk(gclk));
	jdff dff_B_Vzqqvx1Y6_2(.din(w_dff_B_qwE0HqvV7_2),.dout(w_dff_B_Vzqqvx1Y6_2),.clk(gclk));
	jdff dff_B_ny6Xgr5Z5_2(.din(w_dff_B_Vzqqvx1Y6_2),.dout(w_dff_B_ny6Xgr5Z5_2),.clk(gclk));
	jdff dff_B_nKpA752d8_2(.din(w_dff_B_ny6Xgr5Z5_2),.dout(w_dff_B_nKpA752d8_2),.clk(gclk));
	jdff dff_B_Pq9P0IlF6_2(.din(w_dff_B_nKpA752d8_2),.dout(w_dff_B_Pq9P0IlF6_2),.clk(gclk));
	jdff dff_B_CijSerZ83_2(.din(w_dff_B_Pq9P0IlF6_2),.dout(w_dff_B_CijSerZ83_2),.clk(gclk));
	jdff dff_B_BY284Atr3_2(.din(w_dff_B_CijSerZ83_2),.dout(w_dff_B_BY284Atr3_2),.clk(gclk));
	jdff dff_B_MfOHYXdU4_2(.din(w_dff_B_BY284Atr3_2),.dout(w_dff_B_MfOHYXdU4_2),.clk(gclk));
	jdff dff_B_akuff64K9_2(.din(w_dff_B_MfOHYXdU4_2),.dout(w_dff_B_akuff64K9_2),.clk(gclk));
	jdff dff_B_0LkS7Hcw8_2(.din(w_dff_B_akuff64K9_2),.dout(w_dff_B_0LkS7Hcw8_2),.clk(gclk));
	jdff dff_B_cCZloNXb6_2(.din(w_dff_B_0LkS7Hcw8_2),.dout(w_dff_B_cCZloNXb6_2),.clk(gclk));
	jdff dff_B_FZkZf7sr3_2(.din(w_dff_B_cCZloNXb6_2),.dout(w_dff_B_FZkZf7sr3_2),.clk(gclk));
	jdff dff_B_KTLbZe9Y4_2(.din(n884),.dout(w_dff_B_KTLbZe9Y4_2),.clk(gclk));
	jdff dff_B_rEp1xRQD0_1(.din(n858),.dout(w_dff_B_rEp1xRQD0_1),.clk(gclk));
	jdff dff_B_P969pCJR7_2(.din(n759),.dout(w_dff_B_P969pCJR7_2),.clk(gclk));
	jdff dff_B_xE7UWh4n0_2(.din(w_dff_B_P969pCJR7_2),.dout(w_dff_B_xE7UWh4n0_2),.clk(gclk));
	jdff dff_B_nAKMsubZ1_2(.din(w_dff_B_xE7UWh4n0_2),.dout(w_dff_B_nAKMsubZ1_2),.clk(gclk));
	jdff dff_B_QdT3Hk797_2(.din(w_dff_B_nAKMsubZ1_2),.dout(w_dff_B_QdT3Hk797_2),.clk(gclk));
	jdff dff_B_NWTacWc16_2(.din(w_dff_B_QdT3Hk797_2),.dout(w_dff_B_NWTacWc16_2),.clk(gclk));
	jdff dff_B_0pBkhihE4_2(.din(w_dff_B_NWTacWc16_2),.dout(w_dff_B_0pBkhihE4_2),.clk(gclk));
	jdff dff_B_045Z5u9l8_2(.din(w_dff_B_0pBkhihE4_2),.dout(w_dff_B_045Z5u9l8_2),.clk(gclk));
	jdff dff_B_JI6TOvjV8_2(.din(w_dff_B_045Z5u9l8_2),.dout(w_dff_B_JI6TOvjV8_2),.clk(gclk));
	jdff dff_B_j6TlcuSh7_2(.din(w_dff_B_JI6TOvjV8_2),.dout(w_dff_B_j6TlcuSh7_2),.clk(gclk));
	jdff dff_B_1qYIf7LQ4_2(.din(w_dff_B_j6TlcuSh7_2),.dout(w_dff_B_1qYIf7LQ4_2),.clk(gclk));
	jdff dff_B_kkq1ZYEO4_2(.din(w_dff_B_1qYIf7LQ4_2),.dout(w_dff_B_kkq1ZYEO4_2),.clk(gclk));
	jdff dff_B_lqGQoYfm1_2(.din(n781),.dout(w_dff_B_lqGQoYfm1_2),.clk(gclk));
	jdff dff_B_vcmnjSc07_1(.din(n760),.dout(w_dff_B_vcmnjSc07_1),.clk(gclk));
	jdff dff_B_OQTaVFbh9_2(.din(n667),.dout(w_dff_B_OQTaVFbh9_2),.clk(gclk));
	jdff dff_B_WiQUQgJW6_2(.din(w_dff_B_OQTaVFbh9_2),.dout(w_dff_B_WiQUQgJW6_2),.clk(gclk));
	jdff dff_B_5Xp2TDOR3_2(.din(w_dff_B_WiQUQgJW6_2),.dout(w_dff_B_5Xp2TDOR3_2),.clk(gclk));
	jdff dff_B_GD8msEAh0_2(.din(w_dff_B_5Xp2TDOR3_2),.dout(w_dff_B_GD8msEAh0_2),.clk(gclk));
	jdff dff_B_vL374RAq1_2(.din(w_dff_B_GD8msEAh0_2),.dout(w_dff_B_vL374RAq1_2),.clk(gclk));
	jdff dff_B_jfRUn2a51_2(.din(w_dff_B_vL374RAq1_2),.dout(w_dff_B_jfRUn2a51_2),.clk(gclk));
	jdff dff_B_hW8sr8e47_2(.din(w_dff_B_jfRUn2a51_2),.dout(w_dff_B_hW8sr8e47_2),.clk(gclk));
	jdff dff_B_an79LytC2_2(.din(w_dff_B_hW8sr8e47_2),.dout(w_dff_B_an79LytC2_2),.clk(gclk));
	jdff dff_B_Tu7fwmsW0_2(.din(n682),.dout(w_dff_B_Tu7fwmsW0_2),.clk(gclk));
	jdff dff_B_C45puVrB0_2(.din(w_dff_B_Tu7fwmsW0_2),.dout(w_dff_B_C45puVrB0_2),.clk(gclk));
	jdff dff_B_TtyaOiSh6_2(.din(w_dff_B_C45puVrB0_2),.dout(w_dff_B_TtyaOiSh6_2),.clk(gclk));
	jdff dff_B_FFb2oKXS3_1(.din(n668),.dout(w_dff_B_FFb2oKXS3_1),.clk(gclk));
	jdff dff_B_bX1BMdYa4_1(.din(w_dff_B_FFb2oKXS3_1),.dout(w_dff_B_bX1BMdYa4_1),.clk(gclk));
	jdff dff_B_HaImst948_2(.din(n584),.dout(w_dff_B_HaImst948_2),.clk(gclk));
	jdff dff_B_viGk7c4i9_2(.din(w_dff_B_HaImst948_2),.dout(w_dff_B_viGk7c4i9_2),.clk(gclk));
	jdff dff_B_neDSvnNh6_2(.din(w_dff_B_viGk7c4i9_2),.dout(w_dff_B_neDSvnNh6_2),.clk(gclk));
	jdff dff_B_SDciChy19_0(.din(n589),.dout(w_dff_B_SDciChy19_0),.clk(gclk));
	jdff dff_A_CknfTZA03_0(.dout(w_n503_0[0]),.din(w_dff_A_CknfTZA03_0),.clk(gclk));
	jdff dff_A_W0GH72gf8_0(.dout(w_dff_A_CknfTZA03_0),.din(w_dff_A_W0GH72gf8_0),.clk(gclk));
	jdff dff_A_FaAUVDb87_1(.dout(w_n503_0[1]),.din(w_dff_A_FaAUVDb87_1),.clk(gclk));
	jdff dff_A_7j3bc8678_1(.dout(w_dff_A_FaAUVDb87_1),.din(w_dff_A_7j3bc8678_1),.clk(gclk));
	jdff dff_B_v8v4A7LS1_1(.din(n1762),.dout(w_dff_B_v8v4A7LS1_1),.clk(gclk));
	jdff dff_A_NtY58GGi5_1(.dout(w_n1737_0[1]),.din(w_dff_A_NtY58GGi5_1),.clk(gclk));
	jdff dff_B_xxwiKctb7_1(.din(n1735),.dout(w_dff_B_xxwiKctb7_1),.clk(gclk));
	jdff dff_B_LcJA5Bqi7_2(.din(n1699),.dout(w_dff_B_LcJA5Bqi7_2),.clk(gclk));
	jdff dff_B_UfNDRm7f6_2(.din(w_dff_B_LcJA5Bqi7_2),.dout(w_dff_B_UfNDRm7f6_2),.clk(gclk));
	jdff dff_B_GY7K8U8i0_2(.din(w_dff_B_UfNDRm7f6_2),.dout(w_dff_B_GY7K8U8i0_2),.clk(gclk));
	jdff dff_B_RrKfvWFU5_2(.din(w_dff_B_GY7K8U8i0_2),.dout(w_dff_B_RrKfvWFU5_2),.clk(gclk));
	jdff dff_B_OEJT5zoy2_2(.din(w_dff_B_RrKfvWFU5_2),.dout(w_dff_B_OEJT5zoy2_2),.clk(gclk));
	jdff dff_B_rLCi2IIq2_2(.din(w_dff_B_OEJT5zoy2_2),.dout(w_dff_B_rLCi2IIq2_2),.clk(gclk));
	jdff dff_B_Yu4juAjS4_2(.din(w_dff_B_rLCi2IIq2_2),.dout(w_dff_B_Yu4juAjS4_2),.clk(gclk));
	jdff dff_B_8btXofuv6_2(.din(w_dff_B_Yu4juAjS4_2),.dout(w_dff_B_8btXofuv6_2),.clk(gclk));
	jdff dff_B_y0ga9Pip0_2(.din(w_dff_B_8btXofuv6_2),.dout(w_dff_B_y0ga9Pip0_2),.clk(gclk));
	jdff dff_B_tMhWONbk2_2(.din(w_dff_B_y0ga9Pip0_2),.dout(w_dff_B_tMhWONbk2_2),.clk(gclk));
	jdff dff_B_fksUxnGO4_2(.din(w_dff_B_tMhWONbk2_2),.dout(w_dff_B_fksUxnGO4_2),.clk(gclk));
	jdff dff_B_cfaU7hET9_2(.din(w_dff_B_fksUxnGO4_2),.dout(w_dff_B_cfaU7hET9_2),.clk(gclk));
	jdff dff_B_Mc80C5zE7_2(.din(w_dff_B_cfaU7hET9_2),.dout(w_dff_B_Mc80C5zE7_2),.clk(gclk));
	jdff dff_B_d9Gem43W8_2(.din(w_dff_B_Mc80C5zE7_2),.dout(w_dff_B_d9Gem43W8_2),.clk(gclk));
	jdff dff_B_8SSLVOf56_2(.din(w_dff_B_d9Gem43W8_2),.dout(w_dff_B_8SSLVOf56_2),.clk(gclk));
	jdff dff_B_XAQOilhm9_2(.din(w_dff_B_8SSLVOf56_2),.dout(w_dff_B_XAQOilhm9_2),.clk(gclk));
	jdff dff_B_t5VqixS82_2(.din(w_dff_B_XAQOilhm9_2),.dout(w_dff_B_t5VqixS82_2),.clk(gclk));
	jdff dff_B_UWdIDvmW0_2(.din(w_dff_B_t5VqixS82_2),.dout(w_dff_B_UWdIDvmW0_2),.clk(gclk));
	jdff dff_B_GzsXwmeC3_2(.din(w_dff_B_UWdIDvmW0_2),.dout(w_dff_B_GzsXwmeC3_2),.clk(gclk));
	jdff dff_B_exzaH3Wo0_2(.din(w_dff_B_GzsXwmeC3_2),.dout(w_dff_B_exzaH3Wo0_2),.clk(gclk));
	jdff dff_B_9DKXb4LL4_2(.din(w_dff_B_exzaH3Wo0_2),.dout(w_dff_B_9DKXb4LL4_2),.clk(gclk));
	jdff dff_B_dBANWLne5_2(.din(w_dff_B_9DKXb4LL4_2),.dout(w_dff_B_dBANWLne5_2),.clk(gclk));
	jdff dff_B_mDhSZInk3_2(.din(w_dff_B_dBANWLne5_2),.dout(w_dff_B_mDhSZInk3_2),.clk(gclk));
	jdff dff_B_ftViZq3V6_2(.din(w_dff_B_mDhSZInk3_2),.dout(w_dff_B_ftViZq3V6_2),.clk(gclk));
	jdff dff_B_q92XC5u46_2(.din(w_dff_B_ftViZq3V6_2),.dout(w_dff_B_q92XC5u46_2),.clk(gclk));
	jdff dff_B_07zvVMdD3_2(.din(w_dff_B_q92XC5u46_2),.dout(w_dff_B_07zvVMdD3_2),.clk(gclk));
	jdff dff_B_eGdnURNa3_2(.din(w_dff_B_07zvVMdD3_2),.dout(w_dff_B_eGdnURNa3_2),.clk(gclk));
	jdff dff_B_fg9cwdkh9_2(.din(w_dff_B_eGdnURNa3_2),.dout(w_dff_B_fg9cwdkh9_2),.clk(gclk));
	jdff dff_B_jhWfGbIB8_2(.din(w_dff_B_fg9cwdkh9_2),.dout(w_dff_B_jhWfGbIB8_2),.clk(gclk));
	jdff dff_B_EcHovQZ33_2(.din(w_dff_B_jhWfGbIB8_2),.dout(w_dff_B_EcHovQZ33_2),.clk(gclk));
	jdff dff_B_wROgSLxf1_2(.din(w_dff_B_EcHovQZ33_2),.dout(w_dff_B_wROgSLxf1_2),.clk(gclk));
	jdff dff_B_A1qacFVr2_2(.din(w_dff_B_wROgSLxf1_2),.dout(w_dff_B_A1qacFVr2_2),.clk(gclk));
	jdff dff_B_Oyk20svl8_2(.din(w_dff_B_A1qacFVr2_2),.dout(w_dff_B_Oyk20svl8_2),.clk(gclk));
	jdff dff_B_UqmthsR98_2(.din(w_dff_B_Oyk20svl8_2),.dout(w_dff_B_UqmthsR98_2),.clk(gclk));
	jdff dff_B_YTU2SVhg0_2(.din(w_dff_B_UqmthsR98_2),.dout(w_dff_B_YTU2SVhg0_2),.clk(gclk));
	jdff dff_B_2KmRIrEo7_2(.din(w_dff_B_YTU2SVhg0_2),.dout(w_dff_B_2KmRIrEo7_2),.clk(gclk));
	jdff dff_B_MVrdaGf84_2(.din(w_dff_B_2KmRIrEo7_2),.dout(w_dff_B_MVrdaGf84_2),.clk(gclk));
	jdff dff_B_fxFJaqLv6_2(.din(w_dff_B_MVrdaGf84_2),.dout(w_dff_B_fxFJaqLv6_2),.clk(gclk));
	jdff dff_B_cLlliuTa4_2(.din(w_dff_B_fxFJaqLv6_2),.dout(w_dff_B_cLlliuTa4_2),.clk(gclk));
	jdff dff_B_S9w9TuCP7_2(.din(w_dff_B_cLlliuTa4_2),.dout(w_dff_B_S9w9TuCP7_2),.clk(gclk));
	jdff dff_B_hBCZ7gpB9_2(.din(w_dff_B_S9w9TuCP7_2),.dout(w_dff_B_hBCZ7gpB9_2),.clk(gclk));
	jdff dff_B_qoc6ogO33_2(.din(w_dff_B_hBCZ7gpB9_2),.dout(w_dff_B_qoc6ogO33_2),.clk(gclk));
	jdff dff_B_Xhm2qsxB3_2(.din(w_dff_B_qoc6ogO33_2),.dout(w_dff_B_Xhm2qsxB3_2),.clk(gclk));
	jdff dff_B_VJj0m1Do2_2(.din(w_dff_B_Xhm2qsxB3_2),.dout(w_dff_B_VJj0m1Do2_2),.clk(gclk));
	jdff dff_B_70PEJUXi4_2(.din(w_dff_B_VJj0m1Do2_2),.dout(w_dff_B_70PEJUXi4_2),.clk(gclk));
	jdff dff_B_13gBd8gh5_2(.din(w_dff_B_70PEJUXi4_2),.dout(w_dff_B_13gBd8gh5_2),.clk(gclk));
	jdff dff_B_i4eIiAC04_2(.din(w_dff_B_13gBd8gh5_2),.dout(w_dff_B_i4eIiAC04_2),.clk(gclk));
	jdff dff_B_6OjCEdhs7_2(.din(w_dff_B_i4eIiAC04_2),.dout(w_dff_B_6OjCEdhs7_2),.clk(gclk));
	jdff dff_B_JpN0rZj48_2(.din(n1702),.dout(w_dff_B_JpN0rZj48_2),.clk(gclk));
	jdff dff_B_nqvQXrCN6_1(.din(n1700),.dout(w_dff_B_nqvQXrCN6_1),.clk(gclk));
	jdff dff_B_xVGKKs8u1_2(.din(n1658),.dout(w_dff_B_xVGKKs8u1_2),.clk(gclk));
	jdff dff_B_71oxvSmr9_2(.din(w_dff_B_xVGKKs8u1_2),.dout(w_dff_B_71oxvSmr9_2),.clk(gclk));
	jdff dff_B_VDWJjfHx8_2(.din(w_dff_B_71oxvSmr9_2),.dout(w_dff_B_VDWJjfHx8_2),.clk(gclk));
	jdff dff_B_Xf5vl8hx4_2(.din(w_dff_B_VDWJjfHx8_2),.dout(w_dff_B_Xf5vl8hx4_2),.clk(gclk));
	jdff dff_B_irXO5eZF6_2(.din(w_dff_B_Xf5vl8hx4_2),.dout(w_dff_B_irXO5eZF6_2),.clk(gclk));
	jdff dff_B_PdQXvMXa8_2(.din(w_dff_B_irXO5eZF6_2),.dout(w_dff_B_PdQXvMXa8_2),.clk(gclk));
	jdff dff_B_sv9CjH9b1_2(.din(w_dff_B_PdQXvMXa8_2),.dout(w_dff_B_sv9CjH9b1_2),.clk(gclk));
	jdff dff_B_DU2dZiy92_2(.din(w_dff_B_sv9CjH9b1_2),.dout(w_dff_B_DU2dZiy92_2),.clk(gclk));
	jdff dff_B_AWhWqrac2_2(.din(w_dff_B_DU2dZiy92_2),.dout(w_dff_B_AWhWqrac2_2),.clk(gclk));
	jdff dff_B_3O9FsM545_2(.din(w_dff_B_AWhWqrac2_2),.dout(w_dff_B_3O9FsM545_2),.clk(gclk));
	jdff dff_B_RklGZo928_2(.din(w_dff_B_3O9FsM545_2),.dout(w_dff_B_RklGZo928_2),.clk(gclk));
	jdff dff_B_2RJ4PmOO0_2(.din(w_dff_B_RklGZo928_2),.dout(w_dff_B_2RJ4PmOO0_2),.clk(gclk));
	jdff dff_B_EsLEBkm56_2(.din(w_dff_B_2RJ4PmOO0_2),.dout(w_dff_B_EsLEBkm56_2),.clk(gclk));
	jdff dff_B_4dIAflDz6_2(.din(w_dff_B_EsLEBkm56_2),.dout(w_dff_B_4dIAflDz6_2),.clk(gclk));
	jdff dff_B_HGAKkdYK3_2(.din(w_dff_B_4dIAflDz6_2),.dout(w_dff_B_HGAKkdYK3_2),.clk(gclk));
	jdff dff_B_HNQ9b8yK1_2(.din(w_dff_B_HGAKkdYK3_2),.dout(w_dff_B_HNQ9b8yK1_2),.clk(gclk));
	jdff dff_B_R1W7SSfX6_2(.din(w_dff_B_HNQ9b8yK1_2),.dout(w_dff_B_R1W7SSfX6_2),.clk(gclk));
	jdff dff_B_rmX5oKrJ3_2(.din(w_dff_B_R1W7SSfX6_2),.dout(w_dff_B_rmX5oKrJ3_2),.clk(gclk));
	jdff dff_B_ua7b4t665_2(.din(w_dff_B_rmX5oKrJ3_2),.dout(w_dff_B_ua7b4t665_2),.clk(gclk));
	jdff dff_B_14X4e4YK8_2(.din(w_dff_B_ua7b4t665_2),.dout(w_dff_B_14X4e4YK8_2),.clk(gclk));
	jdff dff_B_rjQagSH03_2(.din(w_dff_B_14X4e4YK8_2),.dout(w_dff_B_rjQagSH03_2),.clk(gclk));
	jdff dff_B_tEFkfzHf9_2(.din(w_dff_B_rjQagSH03_2),.dout(w_dff_B_tEFkfzHf9_2),.clk(gclk));
	jdff dff_B_TKVOVmoL9_2(.din(w_dff_B_tEFkfzHf9_2),.dout(w_dff_B_TKVOVmoL9_2),.clk(gclk));
	jdff dff_B_wttPaOG69_2(.din(w_dff_B_TKVOVmoL9_2),.dout(w_dff_B_wttPaOG69_2),.clk(gclk));
	jdff dff_B_lqo5lrpD9_2(.din(w_dff_B_wttPaOG69_2),.dout(w_dff_B_lqo5lrpD9_2),.clk(gclk));
	jdff dff_B_fPe0kNB17_2(.din(w_dff_B_lqo5lrpD9_2),.dout(w_dff_B_fPe0kNB17_2),.clk(gclk));
	jdff dff_B_93UqPvIe5_2(.din(w_dff_B_fPe0kNB17_2),.dout(w_dff_B_93UqPvIe5_2),.clk(gclk));
	jdff dff_B_TyfrnoXd9_2(.din(w_dff_B_93UqPvIe5_2),.dout(w_dff_B_TyfrnoXd9_2),.clk(gclk));
	jdff dff_B_paY5ipUC3_2(.din(w_dff_B_TyfrnoXd9_2),.dout(w_dff_B_paY5ipUC3_2),.clk(gclk));
	jdff dff_B_GvR4kVTr4_2(.din(w_dff_B_paY5ipUC3_2),.dout(w_dff_B_GvR4kVTr4_2),.clk(gclk));
	jdff dff_B_qG3iUPF92_2(.din(w_dff_B_GvR4kVTr4_2),.dout(w_dff_B_qG3iUPF92_2),.clk(gclk));
	jdff dff_B_nZJLRNkM6_2(.din(w_dff_B_qG3iUPF92_2),.dout(w_dff_B_nZJLRNkM6_2),.clk(gclk));
	jdff dff_B_O8zeAHm31_2(.din(w_dff_B_nZJLRNkM6_2),.dout(w_dff_B_O8zeAHm31_2),.clk(gclk));
	jdff dff_B_s43PEsiD1_2(.din(w_dff_B_O8zeAHm31_2),.dout(w_dff_B_s43PEsiD1_2),.clk(gclk));
	jdff dff_B_k418u75v3_2(.din(w_dff_B_s43PEsiD1_2),.dout(w_dff_B_k418u75v3_2),.clk(gclk));
	jdff dff_B_gvo1yXTy3_2(.din(w_dff_B_k418u75v3_2),.dout(w_dff_B_gvo1yXTy3_2),.clk(gclk));
	jdff dff_B_tfm2uLff8_2(.din(w_dff_B_gvo1yXTy3_2),.dout(w_dff_B_tfm2uLff8_2),.clk(gclk));
	jdff dff_B_WnD1Q5Is7_2(.din(w_dff_B_tfm2uLff8_2),.dout(w_dff_B_WnD1Q5Is7_2),.clk(gclk));
	jdff dff_B_uoSSnGrC7_2(.din(w_dff_B_WnD1Q5Is7_2),.dout(w_dff_B_uoSSnGrC7_2),.clk(gclk));
	jdff dff_B_D2DtCYLZ9_2(.din(w_dff_B_uoSSnGrC7_2),.dout(w_dff_B_D2DtCYLZ9_2),.clk(gclk));
	jdff dff_B_PNkfvJ2l3_2(.din(w_dff_B_D2DtCYLZ9_2),.dout(w_dff_B_PNkfvJ2l3_2),.clk(gclk));
	jdff dff_B_DU0dxzrJ1_2(.din(w_dff_B_PNkfvJ2l3_2),.dout(w_dff_B_DU0dxzrJ1_2),.clk(gclk));
	jdff dff_B_gXL6O2rA7_2(.din(w_dff_B_DU0dxzrJ1_2),.dout(w_dff_B_gXL6O2rA7_2),.clk(gclk));
	jdff dff_B_XKc9uIkO5_2(.din(w_dff_B_gXL6O2rA7_2),.dout(w_dff_B_XKc9uIkO5_2),.clk(gclk));
	jdff dff_B_5O1Mhl5G7_2(.din(n1661),.dout(w_dff_B_5O1Mhl5G7_2),.clk(gclk));
	jdff dff_B_tJimsX8j4_1(.din(n1659),.dout(w_dff_B_tJimsX8j4_1),.clk(gclk));
	jdff dff_B_frIaj2RI6_2(.din(n1607),.dout(w_dff_B_frIaj2RI6_2),.clk(gclk));
	jdff dff_B_9GUPOc4G3_2(.din(w_dff_B_frIaj2RI6_2),.dout(w_dff_B_9GUPOc4G3_2),.clk(gclk));
	jdff dff_B_GyDejqQZ6_2(.din(w_dff_B_9GUPOc4G3_2),.dout(w_dff_B_GyDejqQZ6_2),.clk(gclk));
	jdff dff_B_iE8ZleQ34_2(.din(w_dff_B_GyDejqQZ6_2),.dout(w_dff_B_iE8ZleQ34_2),.clk(gclk));
	jdff dff_B_eDtJpeUn1_2(.din(w_dff_B_iE8ZleQ34_2),.dout(w_dff_B_eDtJpeUn1_2),.clk(gclk));
	jdff dff_B_HFfVIqOH7_2(.din(w_dff_B_eDtJpeUn1_2),.dout(w_dff_B_HFfVIqOH7_2),.clk(gclk));
	jdff dff_B_4dmr9fh66_2(.din(w_dff_B_HFfVIqOH7_2),.dout(w_dff_B_4dmr9fh66_2),.clk(gclk));
	jdff dff_B_cf7s3GCB7_2(.din(w_dff_B_4dmr9fh66_2),.dout(w_dff_B_cf7s3GCB7_2),.clk(gclk));
	jdff dff_B_BCl9MYeo6_2(.din(w_dff_B_cf7s3GCB7_2),.dout(w_dff_B_BCl9MYeo6_2),.clk(gclk));
	jdff dff_B_MSz9wcsF6_2(.din(w_dff_B_BCl9MYeo6_2),.dout(w_dff_B_MSz9wcsF6_2),.clk(gclk));
	jdff dff_B_El6EXcGj8_2(.din(w_dff_B_MSz9wcsF6_2),.dout(w_dff_B_El6EXcGj8_2),.clk(gclk));
	jdff dff_B_Z7TBncL22_2(.din(w_dff_B_El6EXcGj8_2),.dout(w_dff_B_Z7TBncL22_2),.clk(gclk));
	jdff dff_B_UQOTd3cL0_2(.din(w_dff_B_Z7TBncL22_2),.dout(w_dff_B_UQOTd3cL0_2),.clk(gclk));
	jdff dff_B_98lTtZWW4_2(.din(w_dff_B_UQOTd3cL0_2),.dout(w_dff_B_98lTtZWW4_2),.clk(gclk));
	jdff dff_B_BCGqecOT6_2(.din(w_dff_B_98lTtZWW4_2),.dout(w_dff_B_BCGqecOT6_2),.clk(gclk));
	jdff dff_B_VRL736xT1_2(.din(w_dff_B_BCGqecOT6_2),.dout(w_dff_B_VRL736xT1_2),.clk(gclk));
	jdff dff_B_xxQ2KoaD6_2(.din(w_dff_B_VRL736xT1_2),.dout(w_dff_B_xxQ2KoaD6_2),.clk(gclk));
	jdff dff_B_pNqlZkVh7_2(.din(w_dff_B_xxQ2KoaD6_2),.dout(w_dff_B_pNqlZkVh7_2),.clk(gclk));
	jdff dff_B_iNPiKcZZ0_2(.din(w_dff_B_pNqlZkVh7_2),.dout(w_dff_B_iNPiKcZZ0_2),.clk(gclk));
	jdff dff_B_71H4NSuf0_2(.din(w_dff_B_iNPiKcZZ0_2),.dout(w_dff_B_71H4NSuf0_2),.clk(gclk));
	jdff dff_B_Ne9kFWUv8_2(.din(w_dff_B_71H4NSuf0_2),.dout(w_dff_B_Ne9kFWUv8_2),.clk(gclk));
	jdff dff_B_CVGfMbPx2_2(.din(w_dff_B_Ne9kFWUv8_2),.dout(w_dff_B_CVGfMbPx2_2),.clk(gclk));
	jdff dff_B_uOr5SNYT5_2(.din(w_dff_B_CVGfMbPx2_2),.dout(w_dff_B_uOr5SNYT5_2),.clk(gclk));
	jdff dff_B_VFBjNAp29_2(.din(w_dff_B_uOr5SNYT5_2),.dout(w_dff_B_VFBjNAp29_2),.clk(gclk));
	jdff dff_B_79WfRfcl2_2(.din(w_dff_B_VFBjNAp29_2),.dout(w_dff_B_79WfRfcl2_2),.clk(gclk));
	jdff dff_B_9MKOUFEs4_2(.din(w_dff_B_79WfRfcl2_2),.dout(w_dff_B_9MKOUFEs4_2),.clk(gclk));
	jdff dff_B_gpppMwAA8_2(.din(w_dff_B_9MKOUFEs4_2),.dout(w_dff_B_gpppMwAA8_2),.clk(gclk));
	jdff dff_B_yGXQaSIF9_2(.din(w_dff_B_gpppMwAA8_2),.dout(w_dff_B_yGXQaSIF9_2),.clk(gclk));
	jdff dff_B_dIFafHB12_2(.din(w_dff_B_yGXQaSIF9_2),.dout(w_dff_B_dIFafHB12_2),.clk(gclk));
	jdff dff_B_NAyzPjTs6_2(.din(w_dff_B_dIFafHB12_2),.dout(w_dff_B_NAyzPjTs6_2),.clk(gclk));
	jdff dff_B_vdgNYJ4J5_2(.din(w_dff_B_NAyzPjTs6_2),.dout(w_dff_B_vdgNYJ4J5_2),.clk(gclk));
	jdff dff_B_i2HGev2t7_2(.din(w_dff_B_vdgNYJ4J5_2),.dout(w_dff_B_i2HGev2t7_2),.clk(gclk));
	jdff dff_B_P98oAzxN1_2(.din(w_dff_B_i2HGev2t7_2),.dout(w_dff_B_P98oAzxN1_2),.clk(gclk));
	jdff dff_B_acRU4ZJT8_2(.din(w_dff_B_P98oAzxN1_2),.dout(w_dff_B_acRU4ZJT8_2),.clk(gclk));
	jdff dff_B_Gaj7Yz0v5_2(.din(w_dff_B_acRU4ZJT8_2),.dout(w_dff_B_Gaj7Yz0v5_2),.clk(gclk));
	jdff dff_B_ygTh3g6T2_2(.din(w_dff_B_Gaj7Yz0v5_2),.dout(w_dff_B_ygTh3g6T2_2),.clk(gclk));
	jdff dff_B_1UjozB693_2(.din(w_dff_B_ygTh3g6T2_2),.dout(w_dff_B_1UjozB693_2),.clk(gclk));
	jdff dff_B_OhDQm7O98_2(.din(w_dff_B_1UjozB693_2),.dout(w_dff_B_OhDQm7O98_2),.clk(gclk));
	jdff dff_B_FcU1j5sf0_2(.din(w_dff_B_OhDQm7O98_2),.dout(w_dff_B_FcU1j5sf0_2),.clk(gclk));
	jdff dff_B_ak5udAVA0_2(.din(w_dff_B_FcU1j5sf0_2),.dout(w_dff_B_ak5udAVA0_2),.clk(gclk));
	jdff dff_B_Ft9mJuO39_2(.din(n1610),.dout(w_dff_B_Ft9mJuO39_2),.clk(gclk));
	jdff dff_B_Jm8IZ2yX3_1(.din(n1608),.dout(w_dff_B_Jm8IZ2yX3_1),.clk(gclk));
	jdff dff_B_TLMwKooz6_2(.din(n1550),.dout(w_dff_B_TLMwKooz6_2),.clk(gclk));
	jdff dff_B_NMoIyqNe9_2(.din(w_dff_B_TLMwKooz6_2),.dout(w_dff_B_NMoIyqNe9_2),.clk(gclk));
	jdff dff_B_3LDtzcG92_2(.din(w_dff_B_NMoIyqNe9_2),.dout(w_dff_B_3LDtzcG92_2),.clk(gclk));
	jdff dff_B_hsZxwD3n0_2(.din(w_dff_B_3LDtzcG92_2),.dout(w_dff_B_hsZxwD3n0_2),.clk(gclk));
	jdff dff_B_ho1mJ0n92_2(.din(w_dff_B_hsZxwD3n0_2),.dout(w_dff_B_ho1mJ0n92_2),.clk(gclk));
	jdff dff_B_tPMLtXZC4_2(.din(w_dff_B_ho1mJ0n92_2),.dout(w_dff_B_tPMLtXZC4_2),.clk(gclk));
	jdff dff_B_jxTAML3I4_2(.din(w_dff_B_tPMLtXZC4_2),.dout(w_dff_B_jxTAML3I4_2),.clk(gclk));
	jdff dff_B_TbalT7X48_2(.din(w_dff_B_jxTAML3I4_2),.dout(w_dff_B_TbalT7X48_2),.clk(gclk));
	jdff dff_B_wi6yv5YD4_2(.din(w_dff_B_TbalT7X48_2),.dout(w_dff_B_wi6yv5YD4_2),.clk(gclk));
	jdff dff_B_9ZMoTj7O2_2(.din(w_dff_B_wi6yv5YD4_2),.dout(w_dff_B_9ZMoTj7O2_2),.clk(gclk));
	jdff dff_B_XhlUlpmN9_2(.din(w_dff_B_9ZMoTj7O2_2),.dout(w_dff_B_XhlUlpmN9_2),.clk(gclk));
	jdff dff_B_0Cy7ds3L9_2(.din(w_dff_B_XhlUlpmN9_2),.dout(w_dff_B_0Cy7ds3L9_2),.clk(gclk));
	jdff dff_B_JEGO43Gh0_2(.din(w_dff_B_0Cy7ds3L9_2),.dout(w_dff_B_JEGO43Gh0_2),.clk(gclk));
	jdff dff_B_tlA6hnOO0_2(.din(w_dff_B_JEGO43Gh0_2),.dout(w_dff_B_tlA6hnOO0_2),.clk(gclk));
	jdff dff_B_zK57mf7V5_2(.din(w_dff_B_tlA6hnOO0_2),.dout(w_dff_B_zK57mf7V5_2),.clk(gclk));
	jdff dff_B_FVjx6qJ20_2(.din(w_dff_B_zK57mf7V5_2),.dout(w_dff_B_FVjx6qJ20_2),.clk(gclk));
	jdff dff_B_FvOmMJRH7_2(.din(w_dff_B_FVjx6qJ20_2),.dout(w_dff_B_FvOmMJRH7_2),.clk(gclk));
	jdff dff_B_ZGkvIe3P5_2(.din(w_dff_B_FvOmMJRH7_2),.dout(w_dff_B_ZGkvIe3P5_2),.clk(gclk));
	jdff dff_B_Ga7PixhE1_2(.din(w_dff_B_ZGkvIe3P5_2),.dout(w_dff_B_Ga7PixhE1_2),.clk(gclk));
	jdff dff_B_rQxouyCF0_2(.din(w_dff_B_Ga7PixhE1_2),.dout(w_dff_B_rQxouyCF0_2),.clk(gclk));
	jdff dff_B_DDpThMtg6_2(.din(w_dff_B_rQxouyCF0_2),.dout(w_dff_B_DDpThMtg6_2),.clk(gclk));
	jdff dff_B_XT9cGpH54_2(.din(w_dff_B_DDpThMtg6_2),.dout(w_dff_B_XT9cGpH54_2),.clk(gclk));
	jdff dff_B_G4qlP3tX2_2(.din(w_dff_B_XT9cGpH54_2),.dout(w_dff_B_G4qlP3tX2_2),.clk(gclk));
	jdff dff_B_o9Ov8vg08_2(.din(w_dff_B_G4qlP3tX2_2),.dout(w_dff_B_o9Ov8vg08_2),.clk(gclk));
	jdff dff_B_Gssfd7i91_2(.din(w_dff_B_o9Ov8vg08_2),.dout(w_dff_B_Gssfd7i91_2),.clk(gclk));
	jdff dff_B_gJP2y6Lp0_2(.din(w_dff_B_Gssfd7i91_2),.dout(w_dff_B_gJP2y6Lp0_2),.clk(gclk));
	jdff dff_B_LjADZ1Q38_2(.din(w_dff_B_gJP2y6Lp0_2),.dout(w_dff_B_LjADZ1Q38_2),.clk(gclk));
	jdff dff_B_KqkiHu1Y1_2(.din(w_dff_B_LjADZ1Q38_2),.dout(w_dff_B_KqkiHu1Y1_2),.clk(gclk));
	jdff dff_B_glA7izOQ6_2(.din(w_dff_B_KqkiHu1Y1_2),.dout(w_dff_B_glA7izOQ6_2),.clk(gclk));
	jdff dff_B_fdEBLbDe0_2(.din(w_dff_B_glA7izOQ6_2),.dout(w_dff_B_fdEBLbDe0_2),.clk(gclk));
	jdff dff_B_PiUtUxb49_2(.din(w_dff_B_fdEBLbDe0_2),.dout(w_dff_B_PiUtUxb49_2),.clk(gclk));
	jdff dff_B_2LgUiKan6_2(.din(w_dff_B_PiUtUxb49_2),.dout(w_dff_B_2LgUiKan6_2),.clk(gclk));
	jdff dff_B_GTlewXVx6_2(.din(w_dff_B_2LgUiKan6_2),.dout(w_dff_B_GTlewXVx6_2),.clk(gclk));
	jdff dff_B_fAhIAaFB0_2(.din(w_dff_B_GTlewXVx6_2),.dout(w_dff_B_fAhIAaFB0_2),.clk(gclk));
	jdff dff_B_dJfnV5gX4_2(.din(w_dff_B_fAhIAaFB0_2),.dout(w_dff_B_dJfnV5gX4_2),.clk(gclk));
	jdff dff_B_74fhHmmo4_2(.din(w_dff_B_dJfnV5gX4_2),.dout(w_dff_B_74fhHmmo4_2),.clk(gclk));
	jdff dff_B_zJmFRF1S3_2(.din(n1553),.dout(w_dff_B_zJmFRF1S3_2),.clk(gclk));
	jdff dff_B_Va8VTkjZ2_1(.din(n1551),.dout(w_dff_B_Va8VTkjZ2_1),.clk(gclk));
	jdff dff_B_evoA3u0e5_2(.din(n1486),.dout(w_dff_B_evoA3u0e5_2),.clk(gclk));
	jdff dff_B_9fjy1hcf7_2(.din(w_dff_B_evoA3u0e5_2),.dout(w_dff_B_9fjy1hcf7_2),.clk(gclk));
	jdff dff_B_jBbS5RuG5_2(.din(w_dff_B_9fjy1hcf7_2),.dout(w_dff_B_jBbS5RuG5_2),.clk(gclk));
	jdff dff_B_FMWHfMZr3_2(.din(w_dff_B_jBbS5RuG5_2),.dout(w_dff_B_FMWHfMZr3_2),.clk(gclk));
	jdff dff_B_DXSiYJu52_2(.din(w_dff_B_FMWHfMZr3_2),.dout(w_dff_B_DXSiYJu52_2),.clk(gclk));
	jdff dff_B_JpNzzsqb0_2(.din(w_dff_B_DXSiYJu52_2),.dout(w_dff_B_JpNzzsqb0_2),.clk(gclk));
	jdff dff_B_18VsRlV54_2(.din(w_dff_B_JpNzzsqb0_2),.dout(w_dff_B_18VsRlV54_2),.clk(gclk));
	jdff dff_B_s0Lwa2JG5_2(.din(w_dff_B_18VsRlV54_2),.dout(w_dff_B_s0Lwa2JG5_2),.clk(gclk));
	jdff dff_B_0ohXihXH0_2(.din(w_dff_B_s0Lwa2JG5_2),.dout(w_dff_B_0ohXihXH0_2),.clk(gclk));
	jdff dff_B_xE5GTrDl4_2(.din(w_dff_B_0ohXihXH0_2),.dout(w_dff_B_xE5GTrDl4_2),.clk(gclk));
	jdff dff_B_AJjxi0RM7_2(.din(w_dff_B_xE5GTrDl4_2),.dout(w_dff_B_AJjxi0RM7_2),.clk(gclk));
	jdff dff_B_kujdne955_2(.din(w_dff_B_AJjxi0RM7_2),.dout(w_dff_B_kujdne955_2),.clk(gclk));
	jdff dff_B_Z4LdgwLL5_2(.din(w_dff_B_kujdne955_2),.dout(w_dff_B_Z4LdgwLL5_2),.clk(gclk));
	jdff dff_B_bng3TENJ8_2(.din(w_dff_B_Z4LdgwLL5_2),.dout(w_dff_B_bng3TENJ8_2),.clk(gclk));
	jdff dff_B_Wt50lZFc8_2(.din(w_dff_B_bng3TENJ8_2),.dout(w_dff_B_Wt50lZFc8_2),.clk(gclk));
	jdff dff_B_BP5LinwD5_2(.din(w_dff_B_Wt50lZFc8_2),.dout(w_dff_B_BP5LinwD5_2),.clk(gclk));
	jdff dff_B_df3C4cg64_2(.din(w_dff_B_BP5LinwD5_2),.dout(w_dff_B_df3C4cg64_2),.clk(gclk));
	jdff dff_B_o6Oc50zP4_2(.din(w_dff_B_df3C4cg64_2),.dout(w_dff_B_o6Oc50zP4_2),.clk(gclk));
	jdff dff_B_sYraskPq2_2(.din(w_dff_B_o6Oc50zP4_2),.dout(w_dff_B_sYraskPq2_2),.clk(gclk));
	jdff dff_B_zdGGUdN12_2(.din(w_dff_B_sYraskPq2_2),.dout(w_dff_B_zdGGUdN12_2),.clk(gclk));
	jdff dff_B_Cy6oI1Cd3_2(.din(w_dff_B_zdGGUdN12_2),.dout(w_dff_B_Cy6oI1Cd3_2),.clk(gclk));
	jdff dff_B_eFwuzjGV8_2(.din(w_dff_B_Cy6oI1Cd3_2),.dout(w_dff_B_eFwuzjGV8_2),.clk(gclk));
	jdff dff_B_25Q8x9Lc6_2(.din(w_dff_B_eFwuzjGV8_2),.dout(w_dff_B_25Q8x9Lc6_2),.clk(gclk));
	jdff dff_B_B7XcN1c74_2(.din(w_dff_B_25Q8x9Lc6_2),.dout(w_dff_B_B7XcN1c74_2),.clk(gclk));
	jdff dff_B_kPP1PRpe4_2(.din(w_dff_B_B7XcN1c74_2),.dout(w_dff_B_kPP1PRpe4_2),.clk(gclk));
	jdff dff_B_LvV2Wnea5_2(.din(w_dff_B_kPP1PRpe4_2),.dout(w_dff_B_LvV2Wnea5_2),.clk(gclk));
	jdff dff_B_LDa4iBRi6_2(.din(w_dff_B_LvV2Wnea5_2),.dout(w_dff_B_LDa4iBRi6_2),.clk(gclk));
	jdff dff_B_9Sb2e7uA3_2(.din(w_dff_B_LDa4iBRi6_2),.dout(w_dff_B_9Sb2e7uA3_2),.clk(gclk));
	jdff dff_B_iaf79csc3_2(.din(w_dff_B_9Sb2e7uA3_2),.dout(w_dff_B_iaf79csc3_2),.clk(gclk));
	jdff dff_B_Jmpy6PLJ5_2(.din(w_dff_B_iaf79csc3_2),.dout(w_dff_B_Jmpy6PLJ5_2),.clk(gclk));
	jdff dff_B_2cvUCt7I8_2(.din(w_dff_B_Jmpy6PLJ5_2),.dout(w_dff_B_2cvUCt7I8_2),.clk(gclk));
	jdff dff_B_vgDz7HGl0_2(.din(w_dff_B_2cvUCt7I8_2),.dout(w_dff_B_vgDz7HGl0_2),.clk(gclk));
	jdff dff_B_NOMqsQbb7_1(.din(n1487),.dout(w_dff_B_NOMqsQbb7_1),.clk(gclk));
	jdff dff_B_rzAh5RcK6_2(.din(n1415),.dout(w_dff_B_rzAh5RcK6_2),.clk(gclk));
	jdff dff_B_TL3k3i9w3_2(.din(w_dff_B_rzAh5RcK6_2),.dout(w_dff_B_TL3k3i9w3_2),.clk(gclk));
	jdff dff_B_BdC1pYdW0_2(.din(w_dff_B_TL3k3i9w3_2),.dout(w_dff_B_BdC1pYdW0_2),.clk(gclk));
	jdff dff_B_vHZ2E8h42_2(.din(w_dff_B_BdC1pYdW0_2),.dout(w_dff_B_vHZ2E8h42_2),.clk(gclk));
	jdff dff_B_KDPvP8p84_2(.din(w_dff_B_vHZ2E8h42_2),.dout(w_dff_B_KDPvP8p84_2),.clk(gclk));
	jdff dff_B_EJm5QPb62_2(.din(w_dff_B_KDPvP8p84_2),.dout(w_dff_B_EJm5QPb62_2),.clk(gclk));
	jdff dff_B_js9r2Jih3_2(.din(w_dff_B_EJm5QPb62_2),.dout(w_dff_B_js9r2Jih3_2),.clk(gclk));
	jdff dff_B_lZryZs087_2(.din(w_dff_B_js9r2Jih3_2),.dout(w_dff_B_lZryZs087_2),.clk(gclk));
	jdff dff_B_KVTqR6m77_2(.din(w_dff_B_lZryZs087_2),.dout(w_dff_B_KVTqR6m77_2),.clk(gclk));
	jdff dff_B_ZrHoH6s26_2(.din(w_dff_B_KVTqR6m77_2),.dout(w_dff_B_ZrHoH6s26_2),.clk(gclk));
	jdff dff_B_iEursiol9_2(.din(w_dff_B_ZrHoH6s26_2),.dout(w_dff_B_iEursiol9_2),.clk(gclk));
	jdff dff_B_E0Pr9wZX7_2(.din(w_dff_B_iEursiol9_2),.dout(w_dff_B_E0Pr9wZX7_2),.clk(gclk));
	jdff dff_B_hwMIAubV0_2(.din(w_dff_B_E0Pr9wZX7_2),.dout(w_dff_B_hwMIAubV0_2),.clk(gclk));
	jdff dff_B_A8KORzvp6_2(.din(w_dff_B_hwMIAubV0_2),.dout(w_dff_B_A8KORzvp6_2),.clk(gclk));
	jdff dff_B_B1JptVA97_2(.din(w_dff_B_A8KORzvp6_2),.dout(w_dff_B_B1JptVA97_2),.clk(gclk));
	jdff dff_B_DruRNvMn3_2(.din(w_dff_B_B1JptVA97_2),.dout(w_dff_B_DruRNvMn3_2),.clk(gclk));
	jdff dff_B_wrziWZtS7_2(.din(w_dff_B_DruRNvMn3_2),.dout(w_dff_B_wrziWZtS7_2),.clk(gclk));
	jdff dff_B_qATlgHj86_2(.din(w_dff_B_wrziWZtS7_2),.dout(w_dff_B_qATlgHj86_2),.clk(gclk));
	jdff dff_B_oB2yIpW74_2(.din(w_dff_B_qATlgHj86_2),.dout(w_dff_B_oB2yIpW74_2),.clk(gclk));
	jdff dff_B_XqrWpKwt9_2(.din(w_dff_B_oB2yIpW74_2),.dout(w_dff_B_XqrWpKwt9_2),.clk(gclk));
	jdff dff_B_UuOQwWzo9_2(.din(w_dff_B_XqrWpKwt9_2),.dout(w_dff_B_UuOQwWzo9_2),.clk(gclk));
	jdff dff_B_df8D3KrU1_2(.din(w_dff_B_UuOQwWzo9_2),.dout(w_dff_B_df8D3KrU1_2),.clk(gclk));
	jdff dff_B_b4AD2SLo8_2(.din(w_dff_B_df8D3KrU1_2),.dout(w_dff_B_b4AD2SLo8_2),.clk(gclk));
	jdff dff_B_DNJKM7Bh8_2(.din(w_dff_B_b4AD2SLo8_2),.dout(w_dff_B_DNJKM7Bh8_2),.clk(gclk));
	jdff dff_B_mhtO42R30_2(.din(w_dff_B_DNJKM7Bh8_2),.dout(w_dff_B_mhtO42R30_2),.clk(gclk));
	jdff dff_B_ljmbFGL86_2(.din(w_dff_B_mhtO42R30_2),.dout(w_dff_B_ljmbFGL86_2),.clk(gclk));
	jdff dff_B_5KP6FtA28_2(.din(w_dff_B_ljmbFGL86_2),.dout(w_dff_B_5KP6FtA28_2),.clk(gclk));
	jdff dff_B_ztnEy9jo6_2(.din(w_dff_B_5KP6FtA28_2),.dout(w_dff_B_ztnEy9jo6_2),.clk(gclk));
	jdff dff_B_XmFqVPUy1_2(.din(w_dff_B_ztnEy9jo6_2),.dout(w_dff_B_XmFqVPUy1_2),.clk(gclk));
	jdff dff_B_uFhzbbnU0_2(.din(n1440),.dout(w_dff_B_uFhzbbnU0_2),.clk(gclk));
	jdff dff_B_JDhLY78t9_1(.din(n1416),.dout(w_dff_B_JDhLY78t9_1),.clk(gclk));
	jdff dff_B_5M1pZYK88_2(.din(n1337),.dout(w_dff_B_5M1pZYK88_2),.clk(gclk));
	jdff dff_B_riturfmM2_2(.din(w_dff_B_5M1pZYK88_2),.dout(w_dff_B_riturfmM2_2),.clk(gclk));
	jdff dff_B_7TW9ku0j0_2(.din(w_dff_B_riturfmM2_2),.dout(w_dff_B_7TW9ku0j0_2),.clk(gclk));
	jdff dff_B_c9TestuX8_2(.din(w_dff_B_7TW9ku0j0_2),.dout(w_dff_B_c9TestuX8_2),.clk(gclk));
	jdff dff_B_cahsJowi9_2(.din(w_dff_B_c9TestuX8_2),.dout(w_dff_B_cahsJowi9_2),.clk(gclk));
	jdff dff_B_nmQWsTmW6_2(.din(w_dff_B_cahsJowi9_2),.dout(w_dff_B_nmQWsTmW6_2),.clk(gclk));
	jdff dff_B_PXQIHeDt4_2(.din(w_dff_B_nmQWsTmW6_2),.dout(w_dff_B_PXQIHeDt4_2),.clk(gclk));
	jdff dff_B_I7y39cJ69_2(.din(w_dff_B_PXQIHeDt4_2),.dout(w_dff_B_I7y39cJ69_2),.clk(gclk));
	jdff dff_B_7f4shHJb2_2(.din(w_dff_B_I7y39cJ69_2),.dout(w_dff_B_7f4shHJb2_2),.clk(gclk));
	jdff dff_B_9p19iKxK6_2(.din(w_dff_B_7f4shHJb2_2),.dout(w_dff_B_9p19iKxK6_2),.clk(gclk));
	jdff dff_B_mv4b9fhm6_2(.din(w_dff_B_9p19iKxK6_2),.dout(w_dff_B_mv4b9fhm6_2),.clk(gclk));
	jdff dff_B_LRfPGIup0_2(.din(w_dff_B_mv4b9fhm6_2),.dout(w_dff_B_LRfPGIup0_2),.clk(gclk));
	jdff dff_B_PJk8RI6r2_2(.din(w_dff_B_LRfPGIup0_2),.dout(w_dff_B_PJk8RI6r2_2),.clk(gclk));
	jdff dff_B_O5bwz0rN8_2(.din(w_dff_B_PJk8RI6r2_2),.dout(w_dff_B_O5bwz0rN8_2),.clk(gclk));
	jdff dff_B_tFx8tzA56_2(.din(w_dff_B_O5bwz0rN8_2),.dout(w_dff_B_tFx8tzA56_2),.clk(gclk));
	jdff dff_B_sYCDs1rW4_2(.din(w_dff_B_tFx8tzA56_2),.dout(w_dff_B_sYCDs1rW4_2),.clk(gclk));
	jdff dff_B_2sZRzt4m7_2(.din(w_dff_B_sYCDs1rW4_2),.dout(w_dff_B_2sZRzt4m7_2),.clk(gclk));
	jdff dff_B_UYh72TEh3_2(.din(w_dff_B_2sZRzt4m7_2),.dout(w_dff_B_UYh72TEh3_2),.clk(gclk));
	jdff dff_B_Q97c5wcB6_2(.din(w_dff_B_UYh72TEh3_2),.dout(w_dff_B_Q97c5wcB6_2),.clk(gclk));
	jdff dff_B_VnPZuiPs2_2(.din(w_dff_B_Q97c5wcB6_2),.dout(w_dff_B_VnPZuiPs2_2),.clk(gclk));
	jdff dff_B_wXh85ooP8_2(.din(w_dff_B_VnPZuiPs2_2),.dout(w_dff_B_wXh85ooP8_2),.clk(gclk));
	jdff dff_B_WKA8rCtM8_2(.din(w_dff_B_wXh85ooP8_2),.dout(w_dff_B_WKA8rCtM8_2),.clk(gclk));
	jdff dff_B_60Sy6Wjk2_2(.din(w_dff_B_WKA8rCtM8_2),.dout(w_dff_B_60Sy6Wjk2_2),.clk(gclk));
	jdff dff_B_2x0X6PHW1_2(.din(w_dff_B_60Sy6Wjk2_2),.dout(w_dff_B_2x0X6PHW1_2),.clk(gclk));
	jdff dff_B_LCZc02rR6_2(.din(w_dff_B_2x0X6PHW1_2),.dout(w_dff_B_LCZc02rR6_2),.clk(gclk));
	jdff dff_B_YqVPXIAC4_2(.din(w_dff_B_LCZc02rR6_2),.dout(w_dff_B_YqVPXIAC4_2),.clk(gclk));
	jdff dff_B_R2EcHsrg1_2(.din(n1362),.dout(w_dff_B_R2EcHsrg1_2),.clk(gclk));
	jdff dff_B_c1etSVAc6_1(.din(n1338),.dout(w_dff_B_c1etSVAc6_1),.clk(gclk));
	jdff dff_B_M8gCdQYB7_2(.din(n1252),.dout(w_dff_B_M8gCdQYB7_2),.clk(gclk));
	jdff dff_B_MA7wPNC92_2(.din(w_dff_B_M8gCdQYB7_2),.dout(w_dff_B_MA7wPNC92_2),.clk(gclk));
	jdff dff_B_eMDarAP04_2(.din(w_dff_B_MA7wPNC92_2),.dout(w_dff_B_eMDarAP04_2),.clk(gclk));
	jdff dff_B_9RpXHOHZ2_2(.din(w_dff_B_eMDarAP04_2),.dout(w_dff_B_9RpXHOHZ2_2),.clk(gclk));
	jdff dff_B_8JK15M254_2(.din(w_dff_B_9RpXHOHZ2_2),.dout(w_dff_B_8JK15M254_2),.clk(gclk));
	jdff dff_B_JLmJrbDQ5_2(.din(w_dff_B_8JK15M254_2),.dout(w_dff_B_JLmJrbDQ5_2),.clk(gclk));
	jdff dff_B_EIoeWHHn1_2(.din(w_dff_B_JLmJrbDQ5_2),.dout(w_dff_B_EIoeWHHn1_2),.clk(gclk));
	jdff dff_B_49I5weLS8_2(.din(w_dff_B_EIoeWHHn1_2),.dout(w_dff_B_49I5weLS8_2),.clk(gclk));
	jdff dff_B_Z5jZu9IV5_2(.din(w_dff_B_49I5weLS8_2),.dout(w_dff_B_Z5jZu9IV5_2),.clk(gclk));
	jdff dff_B_8mrcuC5s8_2(.din(w_dff_B_Z5jZu9IV5_2),.dout(w_dff_B_8mrcuC5s8_2),.clk(gclk));
	jdff dff_B_AGxnscc05_2(.din(w_dff_B_8mrcuC5s8_2),.dout(w_dff_B_AGxnscc05_2),.clk(gclk));
	jdff dff_B_pN9nYxDw0_2(.din(w_dff_B_AGxnscc05_2),.dout(w_dff_B_pN9nYxDw0_2),.clk(gclk));
	jdff dff_B_tTQiORyZ9_2(.din(w_dff_B_pN9nYxDw0_2),.dout(w_dff_B_tTQiORyZ9_2),.clk(gclk));
	jdff dff_B_C7gKbrz84_2(.din(w_dff_B_tTQiORyZ9_2),.dout(w_dff_B_C7gKbrz84_2),.clk(gclk));
	jdff dff_B_fCFaMa1U8_2(.din(w_dff_B_C7gKbrz84_2),.dout(w_dff_B_fCFaMa1U8_2),.clk(gclk));
	jdff dff_B_nu8UxruK7_2(.din(w_dff_B_fCFaMa1U8_2),.dout(w_dff_B_nu8UxruK7_2),.clk(gclk));
	jdff dff_B_N1dwY88e5_2(.din(w_dff_B_nu8UxruK7_2),.dout(w_dff_B_N1dwY88e5_2),.clk(gclk));
	jdff dff_B_ntFrNRJQ9_2(.din(w_dff_B_N1dwY88e5_2),.dout(w_dff_B_ntFrNRJQ9_2),.clk(gclk));
	jdff dff_B_ZYJtKi7w4_2(.din(w_dff_B_ntFrNRJQ9_2),.dout(w_dff_B_ZYJtKi7w4_2),.clk(gclk));
	jdff dff_B_3COP6sPn6_2(.din(w_dff_B_ZYJtKi7w4_2),.dout(w_dff_B_3COP6sPn6_2),.clk(gclk));
	jdff dff_B_jZOdiYwE2_2(.din(w_dff_B_3COP6sPn6_2),.dout(w_dff_B_jZOdiYwE2_2),.clk(gclk));
	jdff dff_B_Fnt90ml08_2(.din(w_dff_B_jZOdiYwE2_2),.dout(w_dff_B_Fnt90ml08_2),.clk(gclk));
	jdff dff_B_im5OGiDU0_2(.din(w_dff_B_Fnt90ml08_2),.dout(w_dff_B_im5OGiDU0_2),.clk(gclk));
	jdff dff_B_N8V3kiDx4_2(.din(n1277),.dout(w_dff_B_N8V3kiDx4_2),.clk(gclk));
	jdff dff_B_QSeZHBz11_1(.din(n1253),.dout(w_dff_B_QSeZHBz11_1),.clk(gclk));
	jdff dff_B_P98EKWL35_2(.din(n1161),.dout(w_dff_B_P98EKWL35_2),.clk(gclk));
	jdff dff_B_EGITGzLL9_2(.din(w_dff_B_P98EKWL35_2),.dout(w_dff_B_EGITGzLL9_2),.clk(gclk));
	jdff dff_B_mZgwUsGu9_2(.din(w_dff_B_EGITGzLL9_2),.dout(w_dff_B_mZgwUsGu9_2),.clk(gclk));
	jdff dff_B_cA0kpSps9_2(.din(w_dff_B_mZgwUsGu9_2),.dout(w_dff_B_cA0kpSps9_2),.clk(gclk));
	jdff dff_B_goHPfu9Y0_2(.din(w_dff_B_cA0kpSps9_2),.dout(w_dff_B_goHPfu9Y0_2),.clk(gclk));
	jdff dff_B_Mb85K9bQ3_2(.din(w_dff_B_goHPfu9Y0_2),.dout(w_dff_B_Mb85K9bQ3_2),.clk(gclk));
	jdff dff_B_IXgUMDHr0_2(.din(w_dff_B_Mb85K9bQ3_2),.dout(w_dff_B_IXgUMDHr0_2),.clk(gclk));
	jdff dff_B_Cp5W3Rwi1_2(.din(w_dff_B_IXgUMDHr0_2),.dout(w_dff_B_Cp5W3Rwi1_2),.clk(gclk));
	jdff dff_B_IgGP0blm0_2(.din(w_dff_B_Cp5W3Rwi1_2),.dout(w_dff_B_IgGP0blm0_2),.clk(gclk));
	jdff dff_B_cGgvSC5R9_2(.din(w_dff_B_IgGP0blm0_2),.dout(w_dff_B_cGgvSC5R9_2),.clk(gclk));
	jdff dff_B_iWfOXjoi9_2(.din(w_dff_B_cGgvSC5R9_2),.dout(w_dff_B_iWfOXjoi9_2),.clk(gclk));
	jdff dff_B_N0bKsjRq7_2(.din(w_dff_B_iWfOXjoi9_2),.dout(w_dff_B_N0bKsjRq7_2),.clk(gclk));
	jdff dff_B_QI8I4yxY7_2(.din(w_dff_B_N0bKsjRq7_2),.dout(w_dff_B_QI8I4yxY7_2),.clk(gclk));
	jdff dff_B_4valJuJS9_2(.din(w_dff_B_QI8I4yxY7_2),.dout(w_dff_B_4valJuJS9_2),.clk(gclk));
	jdff dff_B_LeXv3NRD9_2(.din(w_dff_B_4valJuJS9_2),.dout(w_dff_B_LeXv3NRD9_2),.clk(gclk));
	jdff dff_B_7suEemPV6_2(.din(w_dff_B_LeXv3NRD9_2),.dout(w_dff_B_7suEemPV6_2),.clk(gclk));
	jdff dff_B_A2H9Q2iP2_2(.din(w_dff_B_7suEemPV6_2),.dout(w_dff_B_A2H9Q2iP2_2),.clk(gclk));
	jdff dff_B_vAKrdrEp2_2(.din(w_dff_B_A2H9Q2iP2_2),.dout(w_dff_B_vAKrdrEp2_2),.clk(gclk));
	jdff dff_B_YVbkSeii8_2(.din(w_dff_B_vAKrdrEp2_2),.dout(w_dff_B_YVbkSeii8_2),.clk(gclk));
	jdff dff_B_KiwMMxOK1_2(.din(w_dff_B_YVbkSeii8_2),.dout(w_dff_B_KiwMMxOK1_2),.clk(gclk));
	jdff dff_B_0SMno3DD3_2(.din(n1186),.dout(w_dff_B_0SMno3DD3_2),.clk(gclk));
	jdff dff_B_BuVg0Fal8_1(.din(n1162),.dout(w_dff_B_BuVg0Fal8_1),.clk(gclk));
	jdff dff_B_uRZnHjlG6_2(.din(n1063),.dout(w_dff_B_uRZnHjlG6_2),.clk(gclk));
	jdff dff_B_8JTEWFuK7_2(.din(w_dff_B_uRZnHjlG6_2),.dout(w_dff_B_8JTEWFuK7_2),.clk(gclk));
	jdff dff_B_puOSgXYT4_2(.din(w_dff_B_8JTEWFuK7_2),.dout(w_dff_B_puOSgXYT4_2),.clk(gclk));
	jdff dff_B_VJZf9ttj0_2(.din(w_dff_B_puOSgXYT4_2),.dout(w_dff_B_VJZf9ttj0_2),.clk(gclk));
	jdff dff_B_7XAjTZvt0_2(.din(w_dff_B_VJZf9ttj0_2),.dout(w_dff_B_7XAjTZvt0_2),.clk(gclk));
	jdff dff_B_4ySnrHkG9_2(.din(w_dff_B_7XAjTZvt0_2),.dout(w_dff_B_4ySnrHkG9_2),.clk(gclk));
	jdff dff_B_gutEjDEN5_2(.din(w_dff_B_4ySnrHkG9_2),.dout(w_dff_B_gutEjDEN5_2),.clk(gclk));
	jdff dff_B_jOfjCySS2_2(.din(w_dff_B_gutEjDEN5_2),.dout(w_dff_B_jOfjCySS2_2),.clk(gclk));
	jdff dff_B_4mPQlNFP8_2(.din(w_dff_B_jOfjCySS2_2),.dout(w_dff_B_4mPQlNFP8_2),.clk(gclk));
	jdff dff_B_uubFtQX79_2(.din(w_dff_B_4mPQlNFP8_2),.dout(w_dff_B_uubFtQX79_2),.clk(gclk));
	jdff dff_B_yOc8uIUD3_2(.din(w_dff_B_uubFtQX79_2),.dout(w_dff_B_yOc8uIUD3_2),.clk(gclk));
	jdff dff_B_YMadiFVo3_2(.din(w_dff_B_yOc8uIUD3_2),.dout(w_dff_B_YMadiFVo3_2),.clk(gclk));
	jdff dff_B_KaYKnkPc7_2(.din(w_dff_B_YMadiFVo3_2),.dout(w_dff_B_KaYKnkPc7_2),.clk(gclk));
	jdff dff_B_mmk0al6M9_2(.din(w_dff_B_KaYKnkPc7_2),.dout(w_dff_B_mmk0al6M9_2),.clk(gclk));
	jdff dff_B_ZDLXlVxL8_2(.din(w_dff_B_mmk0al6M9_2),.dout(w_dff_B_ZDLXlVxL8_2),.clk(gclk));
	jdff dff_B_b6mkOZUi2_2(.din(w_dff_B_ZDLXlVxL8_2),.dout(w_dff_B_b6mkOZUi2_2),.clk(gclk));
	jdff dff_B_lyy5Ss3G8_2(.din(w_dff_B_b6mkOZUi2_2),.dout(w_dff_B_lyy5Ss3G8_2),.clk(gclk));
	jdff dff_B_werfbEQm9_2(.din(n1087),.dout(w_dff_B_werfbEQm9_2),.clk(gclk));
	jdff dff_B_KfPZcrTp9_1(.din(n1064),.dout(w_dff_B_KfPZcrTp9_1),.clk(gclk));
	jdff dff_B_F9p8MiAC1_2(.din(n964),.dout(w_dff_B_F9p8MiAC1_2),.clk(gclk));
	jdff dff_B_RecbO2QY7_2(.din(w_dff_B_F9p8MiAC1_2),.dout(w_dff_B_RecbO2QY7_2),.clk(gclk));
	jdff dff_B_vAQcqUzf8_2(.din(w_dff_B_RecbO2QY7_2),.dout(w_dff_B_vAQcqUzf8_2),.clk(gclk));
	jdff dff_B_Jx2yanIf7_2(.din(w_dff_B_vAQcqUzf8_2),.dout(w_dff_B_Jx2yanIf7_2),.clk(gclk));
	jdff dff_B_PcsyNyJa7_2(.din(w_dff_B_Jx2yanIf7_2),.dout(w_dff_B_PcsyNyJa7_2),.clk(gclk));
	jdff dff_B_824f8WqV7_2(.din(w_dff_B_PcsyNyJa7_2),.dout(w_dff_B_824f8WqV7_2),.clk(gclk));
	jdff dff_B_7PsSyqiD1_2(.din(w_dff_B_824f8WqV7_2),.dout(w_dff_B_7PsSyqiD1_2),.clk(gclk));
	jdff dff_B_xsfhwwj28_2(.din(w_dff_B_7PsSyqiD1_2),.dout(w_dff_B_xsfhwwj28_2),.clk(gclk));
	jdff dff_B_ixAxE6Rj1_2(.din(w_dff_B_xsfhwwj28_2),.dout(w_dff_B_ixAxE6Rj1_2),.clk(gclk));
	jdff dff_B_ke8KQ10q4_2(.din(w_dff_B_ixAxE6Rj1_2),.dout(w_dff_B_ke8KQ10q4_2),.clk(gclk));
	jdff dff_B_aAbtQ7CG6_2(.din(w_dff_B_ke8KQ10q4_2),.dout(w_dff_B_aAbtQ7CG6_2),.clk(gclk));
	jdff dff_B_xwT7C5Bk9_2(.din(w_dff_B_aAbtQ7CG6_2),.dout(w_dff_B_xwT7C5Bk9_2),.clk(gclk));
	jdff dff_B_h4GS01EF2_2(.din(w_dff_B_xwT7C5Bk9_2),.dout(w_dff_B_h4GS01EF2_2),.clk(gclk));
	jdff dff_B_UUS9ub6Q8_2(.din(w_dff_B_h4GS01EF2_2),.dout(w_dff_B_UUS9ub6Q8_2),.clk(gclk));
	jdff dff_B_HTmzlJ4h1_2(.din(n988),.dout(w_dff_B_HTmzlJ4h1_2),.clk(gclk));
	jdff dff_B_9T1eoiix9_1(.din(n965),.dout(w_dff_B_9T1eoiix9_1),.clk(gclk));
	jdff dff_B_25xqsulN2_2(.din(n862),.dout(w_dff_B_25xqsulN2_2),.clk(gclk));
	jdff dff_B_uZE0YxWa2_2(.din(w_dff_B_25xqsulN2_2),.dout(w_dff_B_uZE0YxWa2_2),.clk(gclk));
	jdff dff_B_p22cGFRo2_2(.din(w_dff_B_uZE0YxWa2_2),.dout(w_dff_B_p22cGFRo2_2),.clk(gclk));
	jdff dff_B_gIUcLDhp8_2(.din(w_dff_B_p22cGFRo2_2),.dout(w_dff_B_gIUcLDhp8_2),.clk(gclk));
	jdff dff_B_APbCrZMR1_2(.din(w_dff_B_gIUcLDhp8_2),.dout(w_dff_B_APbCrZMR1_2),.clk(gclk));
	jdff dff_B_0Z5tLtuI7_2(.din(w_dff_B_APbCrZMR1_2),.dout(w_dff_B_0Z5tLtuI7_2),.clk(gclk));
	jdff dff_B_N2Yi987I9_2(.din(w_dff_B_0Z5tLtuI7_2),.dout(w_dff_B_N2Yi987I9_2),.clk(gclk));
	jdff dff_B_NijsNKhx4_2(.din(w_dff_B_N2Yi987I9_2),.dout(w_dff_B_NijsNKhx4_2),.clk(gclk));
	jdff dff_B_4SJ33FUb7_2(.din(w_dff_B_NijsNKhx4_2),.dout(w_dff_B_4SJ33FUb7_2),.clk(gclk));
	jdff dff_B_8Ky5uIpk2_2(.din(w_dff_B_4SJ33FUb7_2),.dout(w_dff_B_8Ky5uIpk2_2),.clk(gclk));
	jdff dff_B_5scgfOcd7_2(.din(w_dff_B_8Ky5uIpk2_2),.dout(w_dff_B_5scgfOcd7_2),.clk(gclk));
	jdff dff_B_uELAWVEd5_2(.din(n882),.dout(w_dff_B_uELAWVEd5_2),.clk(gclk));
	jdff dff_B_DhUnkwK37_1(.din(n863),.dout(w_dff_B_DhUnkwK37_1),.clk(gclk));
	jdff dff_B_ozPk56Ju1_2(.din(n764),.dout(w_dff_B_ozPk56Ju1_2),.clk(gclk));
	jdff dff_B_P8dCb00Q8_2(.din(w_dff_B_ozPk56Ju1_2),.dout(w_dff_B_P8dCb00Q8_2),.clk(gclk));
	jdff dff_B_VeOTDZB43_2(.din(w_dff_B_P8dCb00Q8_2),.dout(w_dff_B_VeOTDZB43_2),.clk(gclk));
	jdff dff_B_fqXulsCF2_2(.din(w_dff_B_VeOTDZB43_2),.dout(w_dff_B_fqXulsCF2_2),.clk(gclk));
	jdff dff_B_UT9xhlH88_2(.din(w_dff_B_fqXulsCF2_2),.dout(w_dff_B_UT9xhlH88_2),.clk(gclk));
	jdff dff_B_ZXbv9itt5_2(.din(w_dff_B_UT9xhlH88_2),.dout(w_dff_B_ZXbv9itt5_2),.clk(gclk));
	jdff dff_B_NfygFl5U8_2(.din(w_dff_B_ZXbv9itt5_2),.dout(w_dff_B_NfygFl5U8_2),.clk(gclk));
	jdff dff_B_mnqJR6yD3_2(.din(w_dff_B_NfygFl5U8_2),.dout(w_dff_B_mnqJR6yD3_2),.clk(gclk));
	jdff dff_B_SMblcq3r0_2(.din(n779),.dout(w_dff_B_SMblcq3r0_2),.clk(gclk));
	jdff dff_B_bkF6reiD2_2(.din(w_dff_B_SMblcq3r0_2),.dout(w_dff_B_bkF6reiD2_2),.clk(gclk));
	jdff dff_B_Ol1vyf5o2_2(.din(w_dff_B_bkF6reiD2_2),.dout(w_dff_B_Ol1vyf5o2_2),.clk(gclk));
	jdff dff_B_fnPsljRX7_1(.din(n765),.dout(w_dff_B_fnPsljRX7_1),.clk(gclk));
	jdff dff_B_728XF6378_1(.din(w_dff_B_fnPsljRX7_1),.dout(w_dff_B_728XF6378_1),.clk(gclk));
	jdff dff_B_ti08sdLI4_2(.din(n674),.dout(w_dff_B_ti08sdLI4_2),.clk(gclk));
	jdff dff_B_c9BN89Rz8_2(.din(w_dff_B_ti08sdLI4_2),.dout(w_dff_B_c9BN89Rz8_2),.clk(gclk));
	jdff dff_B_nKqnNbB13_2(.din(w_dff_B_c9BN89Rz8_2),.dout(w_dff_B_nKqnNbB13_2),.clk(gclk));
	jdff dff_B_HZOk2ILt2_0(.din(n679),.dout(w_dff_B_HZOk2ILt2_0),.clk(gclk));
	jdff dff_A_j9vhROl75_0(.dout(w_n586_0[0]),.din(w_dff_A_j9vhROl75_0),.clk(gclk));
	jdff dff_A_jYzDXLF64_0(.dout(w_dff_A_j9vhROl75_0),.din(w_dff_A_jYzDXLF64_0),.clk(gclk));
	jdff dff_A_Inffjh1N0_1(.dout(w_n586_0[1]),.din(w_dff_A_Inffjh1N0_1),.clk(gclk));
	jdff dff_A_Px009JHl6_1(.dout(w_dff_A_Inffjh1N0_1),.din(w_dff_A_Px009JHl6_1),.clk(gclk));
	jdff dff_B_ETaZKDi58_1(.din(n1788),.dout(w_dff_B_ETaZKDi58_1),.clk(gclk));
	jdff dff_A_bbY4ozxq3_1(.dout(w_n1770_0[1]),.din(w_dff_A_bbY4ozxq3_1),.clk(gclk));
	jdff dff_B_FpK85Rv57_1(.din(n1768),.dout(w_dff_B_FpK85Rv57_1),.clk(gclk));
	jdff dff_B_0J7Gc0SF7_2(.din(n1739),.dout(w_dff_B_0J7Gc0SF7_2),.clk(gclk));
	jdff dff_B_RItlMF0x6_2(.din(w_dff_B_0J7Gc0SF7_2),.dout(w_dff_B_RItlMF0x6_2),.clk(gclk));
	jdff dff_B_4MaYUbDN9_2(.din(w_dff_B_RItlMF0x6_2),.dout(w_dff_B_4MaYUbDN9_2),.clk(gclk));
	jdff dff_B_jlak0FYh3_2(.din(w_dff_B_4MaYUbDN9_2),.dout(w_dff_B_jlak0FYh3_2),.clk(gclk));
	jdff dff_B_aHf5LmA61_2(.din(w_dff_B_jlak0FYh3_2),.dout(w_dff_B_aHf5LmA61_2),.clk(gclk));
	jdff dff_B_akiJMh763_2(.din(w_dff_B_aHf5LmA61_2),.dout(w_dff_B_akiJMh763_2),.clk(gclk));
	jdff dff_B_ZOVKDJZA3_2(.din(w_dff_B_akiJMh763_2),.dout(w_dff_B_ZOVKDJZA3_2),.clk(gclk));
	jdff dff_B_IZZAaECC8_2(.din(w_dff_B_ZOVKDJZA3_2),.dout(w_dff_B_IZZAaECC8_2),.clk(gclk));
	jdff dff_B_Jxu8CMxU9_2(.din(w_dff_B_IZZAaECC8_2),.dout(w_dff_B_Jxu8CMxU9_2),.clk(gclk));
	jdff dff_B_5001brXV3_2(.din(w_dff_B_Jxu8CMxU9_2),.dout(w_dff_B_5001brXV3_2),.clk(gclk));
	jdff dff_B_dXcM6R285_2(.din(w_dff_B_5001brXV3_2),.dout(w_dff_B_dXcM6R285_2),.clk(gclk));
	jdff dff_B_Zaz86RKs9_2(.din(w_dff_B_dXcM6R285_2),.dout(w_dff_B_Zaz86RKs9_2),.clk(gclk));
	jdff dff_B_vkoTzYjQ7_2(.din(w_dff_B_Zaz86RKs9_2),.dout(w_dff_B_vkoTzYjQ7_2),.clk(gclk));
	jdff dff_B_UtflPp6t4_2(.din(w_dff_B_vkoTzYjQ7_2),.dout(w_dff_B_UtflPp6t4_2),.clk(gclk));
	jdff dff_B_aXq7BneS8_2(.din(w_dff_B_UtflPp6t4_2),.dout(w_dff_B_aXq7BneS8_2),.clk(gclk));
	jdff dff_B_lucdm2r45_2(.din(w_dff_B_aXq7BneS8_2),.dout(w_dff_B_lucdm2r45_2),.clk(gclk));
	jdff dff_B_cA9cdT9m0_2(.din(w_dff_B_lucdm2r45_2),.dout(w_dff_B_cA9cdT9m0_2),.clk(gclk));
	jdff dff_B_FTlwbQ8F2_2(.din(w_dff_B_cA9cdT9m0_2),.dout(w_dff_B_FTlwbQ8F2_2),.clk(gclk));
	jdff dff_B_IcLyjPpy4_2(.din(w_dff_B_FTlwbQ8F2_2),.dout(w_dff_B_IcLyjPpy4_2),.clk(gclk));
	jdff dff_B_vqs514OL9_2(.din(w_dff_B_IcLyjPpy4_2),.dout(w_dff_B_vqs514OL9_2),.clk(gclk));
	jdff dff_B_o7AcsVXJ5_2(.din(w_dff_B_vqs514OL9_2),.dout(w_dff_B_o7AcsVXJ5_2),.clk(gclk));
	jdff dff_B_SHJbi5ee7_2(.din(w_dff_B_o7AcsVXJ5_2),.dout(w_dff_B_SHJbi5ee7_2),.clk(gclk));
	jdff dff_B_ninwYxOX8_2(.din(w_dff_B_SHJbi5ee7_2),.dout(w_dff_B_ninwYxOX8_2),.clk(gclk));
	jdff dff_B_kYsFLzp61_2(.din(w_dff_B_ninwYxOX8_2),.dout(w_dff_B_kYsFLzp61_2),.clk(gclk));
	jdff dff_B_VxEM1pZE0_2(.din(w_dff_B_kYsFLzp61_2),.dout(w_dff_B_VxEM1pZE0_2),.clk(gclk));
	jdff dff_B_h1enl7NK4_2(.din(w_dff_B_VxEM1pZE0_2),.dout(w_dff_B_h1enl7NK4_2),.clk(gclk));
	jdff dff_B_B2evrgU36_2(.din(w_dff_B_h1enl7NK4_2),.dout(w_dff_B_B2evrgU36_2),.clk(gclk));
	jdff dff_B_AB64OUGE6_2(.din(w_dff_B_B2evrgU36_2),.dout(w_dff_B_AB64OUGE6_2),.clk(gclk));
	jdff dff_B_m2iV2cTa9_2(.din(w_dff_B_AB64OUGE6_2),.dout(w_dff_B_m2iV2cTa9_2),.clk(gclk));
	jdff dff_B_eiv1bLO56_2(.din(w_dff_B_m2iV2cTa9_2),.dout(w_dff_B_eiv1bLO56_2),.clk(gclk));
	jdff dff_B_ERwakILn1_2(.din(w_dff_B_eiv1bLO56_2),.dout(w_dff_B_ERwakILn1_2),.clk(gclk));
	jdff dff_B_3tSAaoF18_2(.din(w_dff_B_ERwakILn1_2),.dout(w_dff_B_3tSAaoF18_2),.clk(gclk));
	jdff dff_B_XNXOuQKM1_2(.din(w_dff_B_3tSAaoF18_2),.dout(w_dff_B_XNXOuQKM1_2),.clk(gclk));
	jdff dff_B_tEtmH9Uw5_2(.din(w_dff_B_XNXOuQKM1_2),.dout(w_dff_B_tEtmH9Uw5_2),.clk(gclk));
	jdff dff_B_ySQWxMvM9_2(.din(w_dff_B_tEtmH9Uw5_2),.dout(w_dff_B_ySQWxMvM9_2),.clk(gclk));
	jdff dff_B_2MHDgYqP0_2(.din(w_dff_B_ySQWxMvM9_2),.dout(w_dff_B_2MHDgYqP0_2),.clk(gclk));
	jdff dff_B_EibVGkX51_2(.din(w_dff_B_2MHDgYqP0_2),.dout(w_dff_B_EibVGkX51_2),.clk(gclk));
	jdff dff_B_hYSdxW9Z8_2(.din(w_dff_B_EibVGkX51_2),.dout(w_dff_B_hYSdxW9Z8_2),.clk(gclk));
	jdff dff_B_XTovOF3k0_2(.din(w_dff_B_hYSdxW9Z8_2),.dout(w_dff_B_XTovOF3k0_2),.clk(gclk));
	jdff dff_B_bLrhwQwU1_2(.din(w_dff_B_XTovOF3k0_2),.dout(w_dff_B_bLrhwQwU1_2),.clk(gclk));
	jdff dff_B_FB5yVCJj2_2(.din(w_dff_B_bLrhwQwU1_2),.dout(w_dff_B_FB5yVCJj2_2),.clk(gclk));
	jdff dff_B_ynNgCZhF8_2(.din(w_dff_B_FB5yVCJj2_2),.dout(w_dff_B_ynNgCZhF8_2),.clk(gclk));
	jdff dff_B_wfrMVCi33_2(.din(w_dff_B_ynNgCZhF8_2),.dout(w_dff_B_wfrMVCi33_2),.clk(gclk));
	jdff dff_B_9YhcK1cV7_2(.din(w_dff_B_wfrMVCi33_2),.dout(w_dff_B_9YhcK1cV7_2),.clk(gclk));
	jdff dff_B_3KexhzEF3_2(.din(w_dff_B_9YhcK1cV7_2),.dout(w_dff_B_3KexhzEF3_2),.clk(gclk));
	jdff dff_B_OOwgU4En3_2(.din(w_dff_B_3KexhzEF3_2),.dout(w_dff_B_OOwgU4En3_2),.clk(gclk));
	jdff dff_B_FkR01uEE7_2(.din(w_dff_B_OOwgU4En3_2),.dout(w_dff_B_FkR01uEE7_2),.clk(gclk));
	jdff dff_B_IXyeuhBa9_2(.din(w_dff_B_FkR01uEE7_2),.dout(w_dff_B_IXyeuhBa9_2),.clk(gclk));
	jdff dff_B_2ARDXNAx6_2(.din(w_dff_B_IXyeuhBa9_2),.dout(w_dff_B_2ARDXNAx6_2),.clk(gclk));
	jdff dff_B_LKZsNJGw4_2(.din(w_dff_B_2ARDXNAx6_2),.dout(w_dff_B_LKZsNJGw4_2),.clk(gclk));
	jdff dff_B_fNHkhFqF1_2(.din(n1742),.dout(w_dff_B_fNHkhFqF1_2),.clk(gclk));
	jdff dff_B_Fwtz0GBI3_1(.din(n1740),.dout(w_dff_B_Fwtz0GBI3_1),.clk(gclk));
	jdff dff_B_c3RRbHhk2_2(.din(n1704),.dout(w_dff_B_c3RRbHhk2_2),.clk(gclk));
	jdff dff_B_Lk9HF94M1_2(.din(w_dff_B_c3RRbHhk2_2),.dout(w_dff_B_Lk9HF94M1_2),.clk(gclk));
	jdff dff_B_rxSKNL5Y5_2(.din(w_dff_B_Lk9HF94M1_2),.dout(w_dff_B_rxSKNL5Y5_2),.clk(gclk));
	jdff dff_B_Y7U2s3x88_2(.din(w_dff_B_rxSKNL5Y5_2),.dout(w_dff_B_Y7U2s3x88_2),.clk(gclk));
	jdff dff_B_V6mELiII3_2(.din(w_dff_B_Y7U2s3x88_2),.dout(w_dff_B_V6mELiII3_2),.clk(gclk));
	jdff dff_B_ekMijgTn3_2(.din(w_dff_B_V6mELiII3_2),.dout(w_dff_B_ekMijgTn3_2),.clk(gclk));
	jdff dff_B_1ior7ngO6_2(.din(w_dff_B_ekMijgTn3_2),.dout(w_dff_B_1ior7ngO6_2),.clk(gclk));
	jdff dff_B_QLK2MV150_2(.din(w_dff_B_1ior7ngO6_2),.dout(w_dff_B_QLK2MV150_2),.clk(gclk));
	jdff dff_B_hHqeOXhU4_2(.din(w_dff_B_QLK2MV150_2),.dout(w_dff_B_hHqeOXhU4_2),.clk(gclk));
	jdff dff_B_gJrM9ugt1_2(.din(w_dff_B_hHqeOXhU4_2),.dout(w_dff_B_gJrM9ugt1_2),.clk(gclk));
	jdff dff_B_3Cucg19M1_2(.din(w_dff_B_gJrM9ugt1_2),.dout(w_dff_B_3Cucg19M1_2),.clk(gclk));
	jdff dff_B_ygluhhKe9_2(.din(w_dff_B_3Cucg19M1_2),.dout(w_dff_B_ygluhhKe9_2),.clk(gclk));
	jdff dff_B_pde6lBDY9_2(.din(w_dff_B_ygluhhKe9_2),.dout(w_dff_B_pde6lBDY9_2),.clk(gclk));
	jdff dff_B_JoOifMwG6_2(.din(w_dff_B_pde6lBDY9_2),.dout(w_dff_B_JoOifMwG6_2),.clk(gclk));
	jdff dff_B_mRU9JJE20_2(.din(w_dff_B_JoOifMwG6_2),.dout(w_dff_B_mRU9JJE20_2),.clk(gclk));
	jdff dff_B_pyQmTLtt9_2(.din(w_dff_B_mRU9JJE20_2),.dout(w_dff_B_pyQmTLtt9_2),.clk(gclk));
	jdff dff_B_56Cfhd2K9_2(.din(w_dff_B_pyQmTLtt9_2),.dout(w_dff_B_56Cfhd2K9_2),.clk(gclk));
	jdff dff_B_Mr5GeYhh2_2(.din(w_dff_B_56Cfhd2K9_2),.dout(w_dff_B_Mr5GeYhh2_2),.clk(gclk));
	jdff dff_B_WZBDpkOC1_2(.din(w_dff_B_Mr5GeYhh2_2),.dout(w_dff_B_WZBDpkOC1_2),.clk(gclk));
	jdff dff_B_m5k2qyLm4_2(.din(w_dff_B_WZBDpkOC1_2),.dout(w_dff_B_m5k2qyLm4_2),.clk(gclk));
	jdff dff_B_weMayPOr5_2(.din(w_dff_B_m5k2qyLm4_2),.dout(w_dff_B_weMayPOr5_2),.clk(gclk));
	jdff dff_B_vOTxNLKD4_2(.din(w_dff_B_weMayPOr5_2),.dout(w_dff_B_vOTxNLKD4_2),.clk(gclk));
	jdff dff_B_QKR0Eo2v2_2(.din(w_dff_B_vOTxNLKD4_2),.dout(w_dff_B_QKR0Eo2v2_2),.clk(gclk));
	jdff dff_B_X0qbQzhS3_2(.din(w_dff_B_QKR0Eo2v2_2),.dout(w_dff_B_X0qbQzhS3_2),.clk(gclk));
	jdff dff_B_RBpoRr485_2(.din(w_dff_B_X0qbQzhS3_2),.dout(w_dff_B_RBpoRr485_2),.clk(gclk));
	jdff dff_B_nOXV2j3n2_2(.din(w_dff_B_RBpoRr485_2),.dout(w_dff_B_nOXV2j3n2_2),.clk(gclk));
	jdff dff_B_695sRdqD8_2(.din(w_dff_B_nOXV2j3n2_2),.dout(w_dff_B_695sRdqD8_2),.clk(gclk));
	jdff dff_B_VcDi0xUx4_2(.din(w_dff_B_695sRdqD8_2),.dout(w_dff_B_VcDi0xUx4_2),.clk(gclk));
	jdff dff_B_FcldosAC6_2(.din(w_dff_B_VcDi0xUx4_2),.dout(w_dff_B_FcldosAC6_2),.clk(gclk));
	jdff dff_B_4a77vzdv1_2(.din(w_dff_B_FcldosAC6_2),.dout(w_dff_B_4a77vzdv1_2),.clk(gclk));
	jdff dff_B_8aF2ljsM5_2(.din(w_dff_B_4a77vzdv1_2),.dout(w_dff_B_8aF2ljsM5_2),.clk(gclk));
	jdff dff_B_lMk6uqgL8_2(.din(w_dff_B_8aF2ljsM5_2),.dout(w_dff_B_lMk6uqgL8_2),.clk(gclk));
	jdff dff_B_e2CVeWme4_2(.din(w_dff_B_lMk6uqgL8_2),.dout(w_dff_B_e2CVeWme4_2),.clk(gclk));
	jdff dff_B_w9DTsEyy9_2(.din(w_dff_B_e2CVeWme4_2),.dout(w_dff_B_w9DTsEyy9_2),.clk(gclk));
	jdff dff_B_kQjwzu7a3_2(.din(w_dff_B_w9DTsEyy9_2),.dout(w_dff_B_kQjwzu7a3_2),.clk(gclk));
	jdff dff_B_T1G30gkP9_2(.din(w_dff_B_kQjwzu7a3_2),.dout(w_dff_B_T1G30gkP9_2),.clk(gclk));
	jdff dff_B_1ORF6B2k3_2(.din(w_dff_B_T1G30gkP9_2),.dout(w_dff_B_1ORF6B2k3_2),.clk(gclk));
	jdff dff_B_ycRTIGjs3_2(.din(w_dff_B_1ORF6B2k3_2),.dout(w_dff_B_ycRTIGjs3_2),.clk(gclk));
	jdff dff_B_aAyhudJG6_2(.din(w_dff_B_ycRTIGjs3_2),.dout(w_dff_B_aAyhudJG6_2),.clk(gclk));
	jdff dff_B_oAdVFYEh6_2(.din(w_dff_B_aAyhudJG6_2),.dout(w_dff_B_oAdVFYEh6_2),.clk(gclk));
	jdff dff_B_J0HjeCu54_2(.din(w_dff_B_oAdVFYEh6_2),.dout(w_dff_B_J0HjeCu54_2),.clk(gclk));
	jdff dff_B_WgN7AWFO4_2(.din(w_dff_B_J0HjeCu54_2),.dout(w_dff_B_WgN7AWFO4_2),.clk(gclk));
	jdff dff_B_gzyMYr3q3_2(.din(w_dff_B_WgN7AWFO4_2),.dout(w_dff_B_gzyMYr3q3_2),.clk(gclk));
	jdff dff_B_tUHatfsD4_2(.din(w_dff_B_gzyMYr3q3_2),.dout(w_dff_B_tUHatfsD4_2),.clk(gclk));
	jdff dff_B_50REtMdL3_2(.din(w_dff_B_tUHatfsD4_2),.dout(w_dff_B_50REtMdL3_2),.clk(gclk));
	jdff dff_B_99nspnyh2_2(.din(w_dff_B_50REtMdL3_2),.dout(w_dff_B_99nspnyh2_2),.clk(gclk));
	jdff dff_B_9eIiVIDf5_2(.din(n1707),.dout(w_dff_B_9eIiVIDf5_2),.clk(gclk));
	jdff dff_B_bKvMIyeU2_1(.din(n1705),.dout(w_dff_B_bKvMIyeU2_1),.clk(gclk));
	jdff dff_B_yyktrpNm2_2(.din(n1663),.dout(w_dff_B_yyktrpNm2_2),.clk(gclk));
	jdff dff_B_bu44eu1B6_2(.din(w_dff_B_yyktrpNm2_2),.dout(w_dff_B_bu44eu1B6_2),.clk(gclk));
	jdff dff_B_Csz3AXj83_2(.din(w_dff_B_bu44eu1B6_2),.dout(w_dff_B_Csz3AXj83_2),.clk(gclk));
	jdff dff_B_5CIQqlsm6_2(.din(w_dff_B_Csz3AXj83_2),.dout(w_dff_B_5CIQqlsm6_2),.clk(gclk));
	jdff dff_B_ZDKXoh2w4_2(.din(w_dff_B_5CIQqlsm6_2),.dout(w_dff_B_ZDKXoh2w4_2),.clk(gclk));
	jdff dff_B_jsKNAhOB9_2(.din(w_dff_B_ZDKXoh2w4_2),.dout(w_dff_B_jsKNAhOB9_2),.clk(gclk));
	jdff dff_B_JAVoLa977_2(.din(w_dff_B_jsKNAhOB9_2),.dout(w_dff_B_JAVoLa977_2),.clk(gclk));
	jdff dff_B_HEN85mpg4_2(.din(w_dff_B_JAVoLa977_2),.dout(w_dff_B_HEN85mpg4_2),.clk(gclk));
	jdff dff_B_nbzo6lFV1_2(.din(w_dff_B_HEN85mpg4_2),.dout(w_dff_B_nbzo6lFV1_2),.clk(gclk));
	jdff dff_B_m8i7scyu2_2(.din(w_dff_B_nbzo6lFV1_2),.dout(w_dff_B_m8i7scyu2_2),.clk(gclk));
	jdff dff_B_jYT64vM47_2(.din(w_dff_B_m8i7scyu2_2),.dout(w_dff_B_jYT64vM47_2),.clk(gclk));
	jdff dff_B_4CLFUP2v3_2(.din(w_dff_B_jYT64vM47_2),.dout(w_dff_B_4CLFUP2v3_2),.clk(gclk));
	jdff dff_B_mATS5brh5_2(.din(w_dff_B_4CLFUP2v3_2),.dout(w_dff_B_mATS5brh5_2),.clk(gclk));
	jdff dff_B_YbI7v3Ie3_2(.din(w_dff_B_mATS5brh5_2),.dout(w_dff_B_YbI7v3Ie3_2),.clk(gclk));
	jdff dff_B_DlVDXHU01_2(.din(w_dff_B_YbI7v3Ie3_2),.dout(w_dff_B_DlVDXHU01_2),.clk(gclk));
	jdff dff_B_x8TSpmYQ5_2(.din(w_dff_B_DlVDXHU01_2),.dout(w_dff_B_x8TSpmYQ5_2),.clk(gclk));
	jdff dff_B_0jjHzCaj3_2(.din(w_dff_B_x8TSpmYQ5_2),.dout(w_dff_B_0jjHzCaj3_2),.clk(gclk));
	jdff dff_B_BzmtM4pE5_2(.din(w_dff_B_0jjHzCaj3_2),.dout(w_dff_B_BzmtM4pE5_2),.clk(gclk));
	jdff dff_B_8EGmo8Zb9_2(.din(w_dff_B_BzmtM4pE5_2),.dout(w_dff_B_8EGmo8Zb9_2),.clk(gclk));
	jdff dff_B_NBkEa6QD6_2(.din(w_dff_B_8EGmo8Zb9_2),.dout(w_dff_B_NBkEa6QD6_2),.clk(gclk));
	jdff dff_B_pBSoxbIG2_2(.din(w_dff_B_NBkEa6QD6_2),.dout(w_dff_B_pBSoxbIG2_2),.clk(gclk));
	jdff dff_B_6Pc5XPYD7_2(.din(w_dff_B_pBSoxbIG2_2),.dout(w_dff_B_6Pc5XPYD7_2),.clk(gclk));
	jdff dff_B_POEtoDlq7_2(.din(w_dff_B_6Pc5XPYD7_2),.dout(w_dff_B_POEtoDlq7_2),.clk(gclk));
	jdff dff_B_PPwdF0Rf0_2(.din(w_dff_B_POEtoDlq7_2),.dout(w_dff_B_PPwdF0Rf0_2),.clk(gclk));
	jdff dff_B_b4gHzTWo4_2(.din(w_dff_B_PPwdF0Rf0_2),.dout(w_dff_B_b4gHzTWo4_2),.clk(gclk));
	jdff dff_B_VXDnRktu9_2(.din(w_dff_B_b4gHzTWo4_2),.dout(w_dff_B_VXDnRktu9_2),.clk(gclk));
	jdff dff_B_I0Jg6Rsa1_2(.din(w_dff_B_VXDnRktu9_2),.dout(w_dff_B_I0Jg6Rsa1_2),.clk(gclk));
	jdff dff_B_JSnNrEa39_2(.din(w_dff_B_I0Jg6Rsa1_2),.dout(w_dff_B_JSnNrEa39_2),.clk(gclk));
	jdff dff_B_f3wVelXf8_2(.din(w_dff_B_JSnNrEa39_2),.dout(w_dff_B_f3wVelXf8_2),.clk(gclk));
	jdff dff_B_b6Qfe2ap6_2(.din(w_dff_B_f3wVelXf8_2),.dout(w_dff_B_b6Qfe2ap6_2),.clk(gclk));
	jdff dff_B_MmGvxAvq5_2(.din(w_dff_B_b6Qfe2ap6_2),.dout(w_dff_B_MmGvxAvq5_2),.clk(gclk));
	jdff dff_B_6IKtcY6Q6_2(.din(w_dff_B_MmGvxAvq5_2),.dout(w_dff_B_6IKtcY6Q6_2),.clk(gclk));
	jdff dff_B_eCb2YjhA9_2(.din(w_dff_B_6IKtcY6Q6_2),.dout(w_dff_B_eCb2YjhA9_2),.clk(gclk));
	jdff dff_B_JodLjeCh7_2(.din(w_dff_B_eCb2YjhA9_2),.dout(w_dff_B_JodLjeCh7_2),.clk(gclk));
	jdff dff_B_cbvCIZhe2_2(.din(w_dff_B_JodLjeCh7_2),.dout(w_dff_B_cbvCIZhe2_2),.clk(gclk));
	jdff dff_B_KCwQgi8Y7_2(.din(w_dff_B_cbvCIZhe2_2),.dout(w_dff_B_KCwQgi8Y7_2),.clk(gclk));
	jdff dff_B_vmF7H9uT4_2(.din(w_dff_B_KCwQgi8Y7_2),.dout(w_dff_B_vmF7H9uT4_2),.clk(gclk));
	jdff dff_B_tNCXlTSp5_2(.din(w_dff_B_vmF7H9uT4_2),.dout(w_dff_B_tNCXlTSp5_2),.clk(gclk));
	jdff dff_B_vik4YCF04_2(.din(w_dff_B_tNCXlTSp5_2),.dout(w_dff_B_vik4YCF04_2),.clk(gclk));
	jdff dff_B_hX7Hdih84_2(.din(w_dff_B_vik4YCF04_2),.dout(w_dff_B_hX7Hdih84_2),.clk(gclk));
	jdff dff_B_6lFIrJ2u2_2(.din(w_dff_B_hX7Hdih84_2),.dout(w_dff_B_6lFIrJ2u2_2),.clk(gclk));
	jdff dff_B_YReXbETt0_2(.din(w_dff_B_6lFIrJ2u2_2),.dout(w_dff_B_YReXbETt0_2),.clk(gclk));
	jdff dff_B_AIRwaqk58_2(.din(n1666),.dout(w_dff_B_AIRwaqk58_2),.clk(gclk));
	jdff dff_B_uWD0VSwd7_1(.din(n1664),.dout(w_dff_B_uWD0VSwd7_1),.clk(gclk));
	jdff dff_B_9EP9codA9_2(.din(n1612),.dout(w_dff_B_9EP9codA9_2),.clk(gclk));
	jdff dff_B_FUCf8NxE5_2(.din(w_dff_B_9EP9codA9_2),.dout(w_dff_B_FUCf8NxE5_2),.clk(gclk));
	jdff dff_B_NtOVCewy8_2(.din(w_dff_B_FUCf8NxE5_2),.dout(w_dff_B_NtOVCewy8_2),.clk(gclk));
	jdff dff_B_AAmU4A087_2(.din(w_dff_B_NtOVCewy8_2),.dout(w_dff_B_AAmU4A087_2),.clk(gclk));
	jdff dff_B_SbpVYm8w6_2(.din(w_dff_B_AAmU4A087_2),.dout(w_dff_B_SbpVYm8w6_2),.clk(gclk));
	jdff dff_B_ARybbmoo7_2(.din(w_dff_B_SbpVYm8w6_2),.dout(w_dff_B_ARybbmoo7_2),.clk(gclk));
	jdff dff_B_E7QsuqFe9_2(.din(w_dff_B_ARybbmoo7_2),.dout(w_dff_B_E7QsuqFe9_2),.clk(gclk));
	jdff dff_B_UY1f4PDI3_2(.din(w_dff_B_E7QsuqFe9_2),.dout(w_dff_B_UY1f4PDI3_2),.clk(gclk));
	jdff dff_B_Fva5N2Ee8_2(.din(w_dff_B_UY1f4PDI3_2),.dout(w_dff_B_Fva5N2Ee8_2),.clk(gclk));
	jdff dff_B_eO7YgJXN7_2(.din(w_dff_B_Fva5N2Ee8_2),.dout(w_dff_B_eO7YgJXN7_2),.clk(gclk));
	jdff dff_B_JswO11cn4_2(.din(w_dff_B_eO7YgJXN7_2),.dout(w_dff_B_JswO11cn4_2),.clk(gclk));
	jdff dff_B_fQ3JW1hU4_2(.din(w_dff_B_JswO11cn4_2),.dout(w_dff_B_fQ3JW1hU4_2),.clk(gclk));
	jdff dff_B_CdvN1CaH5_2(.din(w_dff_B_fQ3JW1hU4_2),.dout(w_dff_B_CdvN1CaH5_2),.clk(gclk));
	jdff dff_B_mIEG6yNy3_2(.din(w_dff_B_CdvN1CaH5_2),.dout(w_dff_B_mIEG6yNy3_2),.clk(gclk));
	jdff dff_B_51WJwNha8_2(.din(w_dff_B_mIEG6yNy3_2),.dout(w_dff_B_51WJwNha8_2),.clk(gclk));
	jdff dff_B_to2EVpos1_2(.din(w_dff_B_51WJwNha8_2),.dout(w_dff_B_to2EVpos1_2),.clk(gclk));
	jdff dff_B_pC4Hs9Zd0_2(.din(w_dff_B_to2EVpos1_2),.dout(w_dff_B_pC4Hs9Zd0_2),.clk(gclk));
	jdff dff_B_o3dLxQRK3_2(.din(w_dff_B_pC4Hs9Zd0_2),.dout(w_dff_B_o3dLxQRK3_2),.clk(gclk));
	jdff dff_B_t0hWqOuN2_2(.din(w_dff_B_o3dLxQRK3_2),.dout(w_dff_B_t0hWqOuN2_2),.clk(gclk));
	jdff dff_B_G3E3fsmW4_2(.din(w_dff_B_t0hWqOuN2_2),.dout(w_dff_B_G3E3fsmW4_2),.clk(gclk));
	jdff dff_B_g4wAVB2x1_2(.din(w_dff_B_G3E3fsmW4_2),.dout(w_dff_B_g4wAVB2x1_2),.clk(gclk));
	jdff dff_B_7k9fO9Rr3_2(.din(w_dff_B_g4wAVB2x1_2),.dout(w_dff_B_7k9fO9Rr3_2),.clk(gclk));
	jdff dff_B_OJA1FgMG0_2(.din(w_dff_B_7k9fO9Rr3_2),.dout(w_dff_B_OJA1FgMG0_2),.clk(gclk));
	jdff dff_B_sdiTLzAQ9_2(.din(w_dff_B_OJA1FgMG0_2),.dout(w_dff_B_sdiTLzAQ9_2),.clk(gclk));
	jdff dff_B_D6jVjiLH7_2(.din(w_dff_B_sdiTLzAQ9_2),.dout(w_dff_B_D6jVjiLH7_2),.clk(gclk));
	jdff dff_B_MNHBAXIj2_2(.din(w_dff_B_D6jVjiLH7_2),.dout(w_dff_B_MNHBAXIj2_2),.clk(gclk));
	jdff dff_B_FmG2Xsxj6_2(.din(w_dff_B_MNHBAXIj2_2),.dout(w_dff_B_FmG2Xsxj6_2),.clk(gclk));
	jdff dff_B_k7thOBWJ9_2(.din(w_dff_B_FmG2Xsxj6_2),.dout(w_dff_B_k7thOBWJ9_2),.clk(gclk));
	jdff dff_B_tOKQBhwO5_2(.din(w_dff_B_k7thOBWJ9_2),.dout(w_dff_B_tOKQBhwO5_2),.clk(gclk));
	jdff dff_B_gXboCuKn2_2(.din(w_dff_B_tOKQBhwO5_2),.dout(w_dff_B_gXboCuKn2_2),.clk(gclk));
	jdff dff_B_LY9pV0b29_2(.din(w_dff_B_gXboCuKn2_2),.dout(w_dff_B_LY9pV0b29_2),.clk(gclk));
	jdff dff_B_M1NuotcH0_2(.din(w_dff_B_LY9pV0b29_2),.dout(w_dff_B_M1NuotcH0_2),.clk(gclk));
	jdff dff_B_bPbudhif3_2(.din(w_dff_B_M1NuotcH0_2),.dout(w_dff_B_bPbudhif3_2),.clk(gclk));
	jdff dff_B_fXlLPqGG9_2(.din(w_dff_B_bPbudhif3_2),.dout(w_dff_B_fXlLPqGG9_2),.clk(gclk));
	jdff dff_B_Tz7bpof40_2(.din(w_dff_B_fXlLPqGG9_2),.dout(w_dff_B_Tz7bpof40_2),.clk(gclk));
	jdff dff_B_5pdr62VP2_2(.din(w_dff_B_Tz7bpof40_2),.dout(w_dff_B_5pdr62VP2_2),.clk(gclk));
	jdff dff_B_pD8rLnxO2_2(.din(w_dff_B_5pdr62VP2_2),.dout(w_dff_B_pD8rLnxO2_2),.clk(gclk));
	jdff dff_B_NU2VaBpl9_2(.din(w_dff_B_pD8rLnxO2_2),.dout(w_dff_B_NU2VaBpl9_2),.clk(gclk));
	jdff dff_B_eSWBskYx7_2(.din(n1615),.dout(w_dff_B_eSWBskYx7_2),.clk(gclk));
	jdff dff_B_td0WxbKe1_1(.din(n1613),.dout(w_dff_B_td0WxbKe1_1),.clk(gclk));
	jdff dff_B_lR1OHnT79_2(.din(n1555),.dout(w_dff_B_lR1OHnT79_2),.clk(gclk));
	jdff dff_B_xExEMAf12_2(.din(w_dff_B_lR1OHnT79_2),.dout(w_dff_B_xExEMAf12_2),.clk(gclk));
	jdff dff_B_VeUPoq5F9_2(.din(w_dff_B_xExEMAf12_2),.dout(w_dff_B_VeUPoq5F9_2),.clk(gclk));
	jdff dff_B_KrF5GXoG2_2(.din(w_dff_B_VeUPoq5F9_2),.dout(w_dff_B_KrF5GXoG2_2),.clk(gclk));
	jdff dff_B_aLsi9sQW2_2(.din(w_dff_B_KrF5GXoG2_2),.dout(w_dff_B_aLsi9sQW2_2),.clk(gclk));
	jdff dff_B_OGRPt5W52_2(.din(w_dff_B_aLsi9sQW2_2),.dout(w_dff_B_OGRPt5W52_2),.clk(gclk));
	jdff dff_B_QeMouNEn3_2(.din(w_dff_B_OGRPt5W52_2),.dout(w_dff_B_QeMouNEn3_2),.clk(gclk));
	jdff dff_B_oWAms1w90_2(.din(w_dff_B_QeMouNEn3_2),.dout(w_dff_B_oWAms1w90_2),.clk(gclk));
	jdff dff_B_1DjPtBAV0_2(.din(w_dff_B_oWAms1w90_2),.dout(w_dff_B_1DjPtBAV0_2),.clk(gclk));
	jdff dff_B_DVvfyar48_2(.din(w_dff_B_1DjPtBAV0_2),.dout(w_dff_B_DVvfyar48_2),.clk(gclk));
	jdff dff_B_SwY7dVbT8_2(.din(w_dff_B_DVvfyar48_2),.dout(w_dff_B_SwY7dVbT8_2),.clk(gclk));
	jdff dff_B_80SXZOAi3_2(.din(w_dff_B_SwY7dVbT8_2),.dout(w_dff_B_80SXZOAi3_2),.clk(gclk));
	jdff dff_B_cZWOhMBL1_2(.din(w_dff_B_80SXZOAi3_2),.dout(w_dff_B_cZWOhMBL1_2),.clk(gclk));
	jdff dff_B_QmLWvtGn2_2(.din(w_dff_B_cZWOhMBL1_2),.dout(w_dff_B_QmLWvtGn2_2),.clk(gclk));
	jdff dff_B_wvOn5yyw2_2(.din(w_dff_B_QmLWvtGn2_2),.dout(w_dff_B_wvOn5yyw2_2),.clk(gclk));
	jdff dff_B_d7pYEh2H7_2(.din(w_dff_B_wvOn5yyw2_2),.dout(w_dff_B_d7pYEh2H7_2),.clk(gclk));
	jdff dff_B_tUBTESTP5_2(.din(w_dff_B_d7pYEh2H7_2),.dout(w_dff_B_tUBTESTP5_2),.clk(gclk));
	jdff dff_B_u2ewzUzZ6_2(.din(w_dff_B_tUBTESTP5_2),.dout(w_dff_B_u2ewzUzZ6_2),.clk(gclk));
	jdff dff_B_fp0m2A314_2(.din(w_dff_B_u2ewzUzZ6_2),.dout(w_dff_B_fp0m2A314_2),.clk(gclk));
	jdff dff_B_Ob11gPZD2_2(.din(w_dff_B_fp0m2A314_2),.dout(w_dff_B_Ob11gPZD2_2),.clk(gclk));
	jdff dff_B_oB4Rfb6C3_2(.din(w_dff_B_Ob11gPZD2_2),.dout(w_dff_B_oB4Rfb6C3_2),.clk(gclk));
	jdff dff_B_kMjtllTd1_2(.din(w_dff_B_oB4Rfb6C3_2),.dout(w_dff_B_kMjtllTd1_2),.clk(gclk));
	jdff dff_B_ws5sLlAW8_2(.din(w_dff_B_kMjtllTd1_2),.dout(w_dff_B_ws5sLlAW8_2),.clk(gclk));
	jdff dff_B_L3Alvh2Z4_2(.din(w_dff_B_ws5sLlAW8_2),.dout(w_dff_B_L3Alvh2Z4_2),.clk(gclk));
	jdff dff_B_n0fR6AjL1_2(.din(w_dff_B_L3Alvh2Z4_2),.dout(w_dff_B_n0fR6AjL1_2),.clk(gclk));
	jdff dff_B_R92hkvZX9_2(.din(w_dff_B_n0fR6AjL1_2),.dout(w_dff_B_R92hkvZX9_2),.clk(gclk));
	jdff dff_B_woDCuFZ14_2(.din(w_dff_B_R92hkvZX9_2),.dout(w_dff_B_woDCuFZ14_2),.clk(gclk));
	jdff dff_B_sDLU0lsD2_2(.din(w_dff_B_woDCuFZ14_2),.dout(w_dff_B_sDLU0lsD2_2),.clk(gclk));
	jdff dff_B_BCpNfPXZ6_2(.din(w_dff_B_sDLU0lsD2_2),.dout(w_dff_B_BCpNfPXZ6_2),.clk(gclk));
	jdff dff_B_2HS8vD7d7_2(.din(w_dff_B_BCpNfPXZ6_2),.dout(w_dff_B_2HS8vD7d7_2),.clk(gclk));
	jdff dff_B_8ujHI00n8_2(.din(w_dff_B_2HS8vD7d7_2),.dout(w_dff_B_8ujHI00n8_2),.clk(gclk));
	jdff dff_B_NzcSzjJV8_2(.din(w_dff_B_8ujHI00n8_2),.dout(w_dff_B_NzcSzjJV8_2),.clk(gclk));
	jdff dff_B_4owFNBrb9_2(.din(w_dff_B_NzcSzjJV8_2),.dout(w_dff_B_4owFNBrb9_2),.clk(gclk));
	jdff dff_B_hVjhuHCc7_2(.din(w_dff_B_4owFNBrb9_2),.dout(w_dff_B_hVjhuHCc7_2),.clk(gclk));
	jdff dff_B_wI1VmqpV6_2(.din(n1558),.dout(w_dff_B_wI1VmqpV6_2),.clk(gclk));
	jdff dff_B_XibNqeFm6_1(.din(n1556),.dout(w_dff_B_XibNqeFm6_1),.clk(gclk));
	jdff dff_B_5pNB9v7M9_2(.din(n1491),.dout(w_dff_B_5pNB9v7M9_2),.clk(gclk));
	jdff dff_B_UcyDdDiE6_2(.din(w_dff_B_5pNB9v7M9_2),.dout(w_dff_B_UcyDdDiE6_2),.clk(gclk));
	jdff dff_B_NUu40z0f2_2(.din(w_dff_B_UcyDdDiE6_2),.dout(w_dff_B_NUu40z0f2_2),.clk(gclk));
	jdff dff_B_WepBRDtN2_2(.din(w_dff_B_NUu40z0f2_2),.dout(w_dff_B_WepBRDtN2_2),.clk(gclk));
	jdff dff_B_AZ0movJs3_2(.din(w_dff_B_WepBRDtN2_2),.dout(w_dff_B_AZ0movJs3_2),.clk(gclk));
	jdff dff_B_cYCPIotE5_2(.din(w_dff_B_AZ0movJs3_2),.dout(w_dff_B_cYCPIotE5_2),.clk(gclk));
	jdff dff_B_GbiYccTs0_2(.din(w_dff_B_cYCPIotE5_2),.dout(w_dff_B_GbiYccTs0_2),.clk(gclk));
	jdff dff_B_xJjZIcJk9_2(.din(w_dff_B_GbiYccTs0_2),.dout(w_dff_B_xJjZIcJk9_2),.clk(gclk));
	jdff dff_B_jZwxBOn14_2(.din(w_dff_B_xJjZIcJk9_2),.dout(w_dff_B_jZwxBOn14_2),.clk(gclk));
	jdff dff_B_qVWqC9VF1_2(.din(w_dff_B_jZwxBOn14_2),.dout(w_dff_B_qVWqC9VF1_2),.clk(gclk));
	jdff dff_B_KMZ0YBCs6_2(.din(w_dff_B_qVWqC9VF1_2),.dout(w_dff_B_KMZ0YBCs6_2),.clk(gclk));
	jdff dff_B_s8RtqUdJ7_2(.din(w_dff_B_KMZ0YBCs6_2),.dout(w_dff_B_s8RtqUdJ7_2),.clk(gclk));
	jdff dff_B_nIWwlrBD2_2(.din(w_dff_B_s8RtqUdJ7_2),.dout(w_dff_B_nIWwlrBD2_2),.clk(gclk));
	jdff dff_B_GMfgLclG6_2(.din(w_dff_B_nIWwlrBD2_2),.dout(w_dff_B_GMfgLclG6_2),.clk(gclk));
	jdff dff_B_0ZKYV8au2_2(.din(w_dff_B_GMfgLclG6_2),.dout(w_dff_B_0ZKYV8au2_2),.clk(gclk));
	jdff dff_B_BlNw9jrD4_2(.din(w_dff_B_0ZKYV8au2_2),.dout(w_dff_B_BlNw9jrD4_2),.clk(gclk));
	jdff dff_B_ouJldoFm3_2(.din(w_dff_B_BlNw9jrD4_2),.dout(w_dff_B_ouJldoFm3_2),.clk(gclk));
	jdff dff_B_NCxsBkjw6_2(.din(w_dff_B_ouJldoFm3_2),.dout(w_dff_B_NCxsBkjw6_2),.clk(gclk));
	jdff dff_B_6pBiAHQg1_2(.din(w_dff_B_NCxsBkjw6_2),.dout(w_dff_B_6pBiAHQg1_2),.clk(gclk));
	jdff dff_B_JepAfnws1_2(.din(w_dff_B_6pBiAHQg1_2),.dout(w_dff_B_JepAfnws1_2),.clk(gclk));
	jdff dff_B_A0zD2iT57_2(.din(w_dff_B_JepAfnws1_2),.dout(w_dff_B_A0zD2iT57_2),.clk(gclk));
	jdff dff_B_panCBQgy1_2(.din(w_dff_B_A0zD2iT57_2),.dout(w_dff_B_panCBQgy1_2),.clk(gclk));
	jdff dff_B_Tg96JtO59_2(.din(w_dff_B_panCBQgy1_2),.dout(w_dff_B_Tg96JtO59_2),.clk(gclk));
	jdff dff_B_JLp5wwiB9_2(.din(w_dff_B_Tg96JtO59_2),.dout(w_dff_B_JLp5wwiB9_2),.clk(gclk));
	jdff dff_B_VJ36D2oQ1_2(.din(w_dff_B_JLp5wwiB9_2),.dout(w_dff_B_VJ36D2oQ1_2),.clk(gclk));
	jdff dff_B_jpKFKqBO4_2(.din(w_dff_B_VJ36D2oQ1_2),.dout(w_dff_B_jpKFKqBO4_2),.clk(gclk));
	jdff dff_B_Z354jVBY8_2(.din(w_dff_B_jpKFKqBO4_2),.dout(w_dff_B_Z354jVBY8_2),.clk(gclk));
	jdff dff_B_3JIOsrOB6_2(.din(w_dff_B_Z354jVBY8_2),.dout(w_dff_B_3JIOsrOB6_2),.clk(gclk));
	jdff dff_B_6o2KRl8z8_2(.din(w_dff_B_3JIOsrOB6_2),.dout(w_dff_B_6o2KRl8z8_2),.clk(gclk));
	jdff dff_B_9zzKoBVo7_2(.din(w_dff_B_6o2KRl8z8_2),.dout(w_dff_B_9zzKoBVo7_2),.clk(gclk));
	jdff dff_B_Z5aK2Mqf8_2(.din(n1494),.dout(w_dff_B_Z5aK2Mqf8_2),.clk(gclk));
	jdff dff_B_1lgDSPcO0_1(.din(n1492),.dout(w_dff_B_1lgDSPcO0_1),.clk(gclk));
	jdff dff_B_lsal0nxM1_2(.din(n1420),.dout(w_dff_B_lsal0nxM1_2),.clk(gclk));
	jdff dff_B_4cOYH2Bv9_2(.din(w_dff_B_lsal0nxM1_2),.dout(w_dff_B_4cOYH2Bv9_2),.clk(gclk));
	jdff dff_B_tfd2igIn3_2(.din(w_dff_B_4cOYH2Bv9_2),.dout(w_dff_B_tfd2igIn3_2),.clk(gclk));
	jdff dff_B_6gupaslH9_2(.din(w_dff_B_tfd2igIn3_2),.dout(w_dff_B_6gupaslH9_2),.clk(gclk));
	jdff dff_B_sU53PKXp3_2(.din(w_dff_B_6gupaslH9_2),.dout(w_dff_B_sU53PKXp3_2),.clk(gclk));
	jdff dff_B_e6AALpjn5_2(.din(w_dff_B_sU53PKXp3_2),.dout(w_dff_B_e6AALpjn5_2),.clk(gclk));
	jdff dff_B_IR7MDgCE1_2(.din(w_dff_B_e6AALpjn5_2),.dout(w_dff_B_IR7MDgCE1_2),.clk(gclk));
	jdff dff_B_b3GhAzpq8_2(.din(w_dff_B_IR7MDgCE1_2),.dout(w_dff_B_b3GhAzpq8_2),.clk(gclk));
	jdff dff_B_PCdLxVcJ4_2(.din(w_dff_B_b3GhAzpq8_2),.dout(w_dff_B_PCdLxVcJ4_2),.clk(gclk));
	jdff dff_B_O2Kwrf1q8_2(.din(w_dff_B_PCdLxVcJ4_2),.dout(w_dff_B_O2Kwrf1q8_2),.clk(gclk));
	jdff dff_B_CRz5nzIH8_2(.din(w_dff_B_O2Kwrf1q8_2),.dout(w_dff_B_CRz5nzIH8_2),.clk(gclk));
	jdff dff_B_N0dTfSQ35_2(.din(w_dff_B_CRz5nzIH8_2),.dout(w_dff_B_N0dTfSQ35_2),.clk(gclk));
	jdff dff_B_lBy6FCxs8_2(.din(w_dff_B_N0dTfSQ35_2),.dout(w_dff_B_lBy6FCxs8_2),.clk(gclk));
	jdff dff_B_mpU0aF9C6_2(.din(w_dff_B_lBy6FCxs8_2),.dout(w_dff_B_mpU0aF9C6_2),.clk(gclk));
	jdff dff_B_s1C4YxQa4_2(.din(w_dff_B_mpU0aF9C6_2),.dout(w_dff_B_s1C4YxQa4_2),.clk(gclk));
	jdff dff_B_pz1SME7d8_2(.din(w_dff_B_s1C4YxQa4_2),.dout(w_dff_B_pz1SME7d8_2),.clk(gclk));
	jdff dff_B_SGkNHoRI2_2(.din(w_dff_B_pz1SME7d8_2),.dout(w_dff_B_SGkNHoRI2_2),.clk(gclk));
	jdff dff_B_oZc2EKs89_2(.din(w_dff_B_SGkNHoRI2_2),.dout(w_dff_B_oZc2EKs89_2),.clk(gclk));
	jdff dff_B_L5MuNCV12_2(.din(w_dff_B_oZc2EKs89_2),.dout(w_dff_B_L5MuNCV12_2),.clk(gclk));
	jdff dff_B_7ljeYh7z9_2(.din(w_dff_B_L5MuNCV12_2),.dout(w_dff_B_7ljeYh7z9_2),.clk(gclk));
	jdff dff_B_KrP08cMV3_2(.din(w_dff_B_7ljeYh7z9_2),.dout(w_dff_B_KrP08cMV3_2),.clk(gclk));
	jdff dff_B_be7HGxfU7_2(.din(w_dff_B_KrP08cMV3_2),.dout(w_dff_B_be7HGxfU7_2),.clk(gclk));
	jdff dff_B_XSatfJ2t5_2(.din(w_dff_B_be7HGxfU7_2),.dout(w_dff_B_XSatfJ2t5_2),.clk(gclk));
	jdff dff_B_Kha9fibu0_2(.din(w_dff_B_XSatfJ2t5_2),.dout(w_dff_B_Kha9fibu0_2),.clk(gclk));
	jdff dff_B_Do3CHlZJ4_2(.din(w_dff_B_Kha9fibu0_2),.dout(w_dff_B_Do3CHlZJ4_2),.clk(gclk));
	jdff dff_B_e40zLt7F6_2(.din(w_dff_B_Do3CHlZJ4_2),.dout(w_dff_B_e40zLt7F6_2),.clk(gclk));
	jdff dff_B_n19aq9WK1_1(.din(n1421),.dout(w_dff_B_n19aq9WK1_1),.clk(gclk));
	jdff dff_B_ocY5mxKI8_2(.din(n1342),.dout(w_dff_B_ocY5mxKI8_2),.clk(gclk));
	jdff dff_B_cxtn1Egs2_2(.din(w_dff_B_ocY5mxKI8_2),.dout(w_dff_B_cxtn1Egs2_2),.clk(gclk));
	jdff dff_B_1W71HvGN9_2(.din(w_dff_B_cxtn1Egs2_2),.dout(w_dff_B_1W71HvGN9_2),.clk(gclk));
	jdff dff_B_BD4TXV0W6_2(.din(w_dff_B_1W71HvGN9_2),.dout(w_dff_B_BD4TXV0W6_2),.clk(gclk));
	jdff dff_B_dGnguKrX3_2(.din(w_dff_B_BD4TXV0W6_2),.dout(w_dff_B_dGnguKrX3_2),.clk(gclk));
	jdff dff_B_9hSTjei00_2(.din(w_dff_B_dGnguKrX3_2),.dout(w_dff_B_9hSTjei00_2),.clk(gclk));
	jdff dff_B_tiimYwi14_2(.din(w_dff_B_9hSTjei00_2),.dout(w_dff_B_tiimYwi14_2),.clk(gclk));
	jdff dff_B_Hxj5JbAl9_2(.din(w_dff_B_tiimYwi14_2),.dout(w_dff_B_Hxj5JbAl9_2),.clk(gclk));
	jdff dff_B_jGtmp9vK8_2(.din(w_dff_B_Hxj5JbAl9_2),.dout(w_dff_B_jGtmp9vK8_2),.clk(gclk));
	jdff dff_B_JaunJOqk6_2(.din(w_dff_B_jGtmp9vK8_2),.dout(w_dff_B_JaunJOqk6_2),.clk(gclk));
	jdff dff_B_mKJ5yvwJ9_2(.din(w_dff_B_JaunJOqk6_2),.dout(w_dff_B_mKJ5yvwJ9_2),.clk(gclk));
	jdff dff_B_KHG8SNb73_2(.din(w_dff_B_mKJ5yvwJ9_2),.dout(w_dff_B_KHG8SNb73_2),.clk(gclk));
	jdff dff_B_5FD3ET3e4_2(.din(w_dff_B_KHG8SNb73_2),.dout(w_dff_B_5FD3ET3e4_2),.clk(gclk));
	jdff dff_B_7tHAWO2m6_2(.din(w_dff_B_5FD3ET3e4_2),.dout(w_dff_B_7tHAWO2m6_2),.clk(gclk));
	jdff dff_B_Rv9qCRPw6_2(.din(w_dff_B_7tHAWO2m6_2),.dout(w_dff_B_Rv9qCRPw6_2),.clk(gclk));
	jdff dff_B_ZJ6g7wCM7_2(.din(w_dff_B_Rv9qCRPw6_2),.dout(w_dff_B_ZJ6g7wCM7_2),.clk(gclk));
	jdff dff_B_YKz3RTM64_2(.din(w_dff_B_ZJ6g7wCM7_2),.dout(w_dff_B_YKz3RTM64_2),.clk(gclk));
	jdff dff_B_qrh9tmJJ1_2(.din(w_dff_B_YKz3RTM64_2),.dout(w_dff_B_qrh9tmJJ1_2),.clk(gclk));
	jdff dff_B_aafwFHd19_2(.din(w_dff_B_qrh9tmJJ1_2),.dout(w_dff_B_aafwFHd19_2),.clk(gclk));
	jdff dff_B_DZkDxv8R1_2(.din(w_dff_B_aafwFHd19_2),.dout(w_dff_B_DZkDxv8R1_2),.clk(gclk));
	jdff dff_B_ffShLiOs1_2(.din(w_dff_B_DZkDxv8R1_2),.dout(w_dff_B_ffShLiOs1_2),.clk(gclk));
	jdff dff_B_lHCWwTcy0_2(.din(w_dff_B_ffShLiOs1_2),.dout(w_dff_B_lHCWwTcy0_2),.clk(gclk));
	jdff dff_B_MxE3o1cU9_2(.din(w_dff_B_lHCWwTcy0_2),.dout(w_dff_B_MxE3o1cU9_2),.clk(gclk));
	jdff dff_B_9iqGyKXP9_2(.din(n1360),.dout(w_dff_B_9iqGyKXP9_2),.clk(gclk));
	jdff dff_B_hdB6e6E61_1(.din(n1343),.dout(w_dff_B_hdB6e6E61_1),.clk(gclk));
	jdff dff_B_M8Ag9vRB1_2(.din(n1257),.dout(w_dff_B_M8Ag9vRB1_2),.clk(gclk));
	jdff dff_B_Fcx6PIzr0_2(.din(w_dff_B_M8Ag9vRB1_2),.dout(w_dff_B_Fcx6PIzr0_2),.clk(gclk));
	jdff dff_B_CJ1gukER8_2(.din(w_dff_B_Fcx6PIzr0_2),.dout(w_dff_B_CJ1gukER8_2),.clk(gclk));
	jdff dff_B_6XjSYidV3_2(.din(w_dff_B_CJ1gukER8_2),.dout(w_dff_B_6XjSYidV3_2),.clk(gclk));
	jdff dff_B_UsYIXMgo5_2(.din(w_dff_B_6XjSYidV3_2),.dout(w_dff_B_UsYIXMgo5_2),.clk(gclk));
	jdff dff_B_UYI1MK2r4_2(.din(w_dff_B_UsYIXMgo5_2),.dout(w_dff_B_UYI1MK2r4_2),.clk(gclk));
	jdff dff_B_1cF1h3Hw3_2(.din(w_dff_B_UYI1MK2r4_2),.dout(w_dff_B_1cF1h3Hw3_2),.clk(gclk));
	jdff dff_B_bC9exOXa0_2(.din(w_dff_B_1cF1h3Hw3_2),.dout(w_dff_B_bC9exOXa0_2),.clk(gclk));
	jdff dff_B_1otDCR9r1_2(.din(w_dff_B_bC9exOXa0_2),.dout(w_dff_B_1otDCR9r1_2),.clk(gclk));
	jdff dff_B_FmaWGmFY1_2(.din(w_dff_B_1otDCR9r1_2),.dout(w_dff_B_FmaWGmFY1_2),.clk(gclk));
	jdff dff_B_6waAWmvV4_2(.din(w_dff_B_FmaWGmFY1_2),.dout(w_dff_B_6waAWmvV4_2),.clk(gclk));
	jdff dff_B_3EcrslVx7_2(.din(w_dff_B_6waAWmvV4_2),.dout(w_dff_B_3EcrslVx7_2),.clk(gclk));
	jdff dff_B_pEUeYrei9_2(.din(w_dff_B_3EcrslVx7_2),.dout(w_dff_B_pEUeYrei9_2),.clk(gclk));
	jdff dff_B_t3pldeuE7_2(.din(w_dff_B_pEUeYrei9_2),.dout(w_dff_B_t3pldeuE7_2),.clk(gclk));
	jdff dff_B_WppsMTJk8_2(.din(w_dff_B_t3pldeuE7_2),.dout(w_dff_B_WppsMTJk8_2),.clk(gclk));
	jdff dff_B_9DC59lOa2_2(.din(w_dff_B_WppsMTJk8_2),.dout(w_dff_B_9DC59lOa2_2),.clk(gclk));
	jdff dff_B_qh3rdMGx4_2(.din(w_dff_B_9DC59lOa2_2),.dout(w_dff_B_qh3rdMGx4_2),.clk(gclk));
	jdff dff_B_9aVeab610_2(.din(w_dff_B_qh3rdMGx4_2),.dout(w_dff_B_9aVeab610_2),.clk(gclk));
	jdff dff_B_hZIvGtRx0_2(.din(w_dff_B_9aVeab610_2),.dout(w_dff_B_hZIvGtRx0_2),.clk(gclk));
	jdff dff_B_bV6shDjr6_2(.din(w_dff_B_hZIvGtRx0_2),.dout(w_dff_B_bV6shDjr6_2),.clk(gclk));
	jdff dff_B_xxLYShRk6_2(.din(n1275),.dout(w_dff_B_xxLYShRk6_2),.clk(gclk));
	jdff dff_B_mjBQCs7h3_1(.din(n1258),.dout(w_dff_B_mjBQCs7h3_1),.clk(gclk));
	jdff dff_B_fRNpdsny8_2(.din(n1166),.dout(w_dff_B_fRNpdsny8_2),.clk(gclk));
	jdff dff_B_afn9dtFl0_2(.din(w_dff_B_fRNpdsny8_2),.dout(w_dff_B_afn9dtFl0_2),.clk(gclk));
	jdff dff_B_wtD52uC91_2(.din(w_dff_B_afn9dtFl0_2),.dout(w_dff_B_wtD52uC91_2),.clk(gclk));
	jdff dff_B_r4uCN1Ci0_2(.din(w_dff_B_wtD52uC91_2),.dout(w_dff_B_r4uCN1Ci0_2),.clk(gclk));
	jdff dff_B_j4ddA7yP4_2(.din(w_dff_B_r4uCN1Ci0_2),.dout(w_dff_B_j4ddA7yP4_2),.clk(gclk));
	jdff dff_B_yrUthAg95_2(.din(w_dff_B_j4ddA7yP4_2),.dout(w_dff_B_yrUthAg95_2),.clk(gclk));
	jdff dff_B_CMldEojj1_2(.din(w_dff_B_yrUthAg95_2),.dout(w_dff_B_CMldEojj1_2),.clk(gclk));
	jdff dff_B_xllfnvYM3_2(.din(w_dff_B_CMldEojj1_2),.dout(w_dff_B_xllfnvYM3_2),.clk(gclk));
	jdff dff_B_7s3mM2d98_2(.din(w_dff_B_xllfnvYM3_2),.dout(w_dff_B_7s3mM2d98_2),.clk(gclk));
	jdff dff_B_QyqQjF4b8_2(.din(w_dff_B_7s3mM2d98_2),.dout(w_dff_B_QyqQjF4b8_2),.clk(gclk));
	jdff dff_B_2RLERi4D3_2(.din(w_dff_B_QyqQjF4b8_2),.dout(w_dff_B_2RLERi4D3_2),.clk(gclk));
	jdff dff_B_hsEK8ghl4_2(.din(w_dff_B_2RLERi4D3_2),.dout(w_dff_B_hsEK8ghl4_2),.clk(gclk));
	jdff dff_B_VbBFQejO1_2(.din(w_dff_B_hsEK8ghl4_2),.dout(w_dff_B_VbBFQejO1_2),.clk(gclk));
	jdff dff_B_NeAIDJ7I6_2(.din(w_dff_B_VbBFQejO1_2),.dout(w_dff_B_NeAIDJ7I6_2),.clk(gclk));
	jdff dff_B_AXWu38c30_2(.din(w_dff_B_NeAIDJ7I6_2),.dout(w_dff_B_AXWu38c30_2),.clk(gclk));
	jdff dff_B_mSEpAkhb3_2(.din(w_dff_B_AXWu38c30_2),.dout(w_dff_B_mSEpAkhb3_2),.clk(gclk));
	jdff dff_B_AdX8cphv6_2(.din(w_dff_B_mSEpAkhb3_2),.dout(w_dff_B_AdX8cphv6_2),.clk(gclk));
	jdff dff_B_pDsZakwK6_2(.din(n1184),.dout(w_dff_B_pDsZakwK6_2),.clk(gclk));
	jdff dff_B_s9KZOleJ3_1(.din(n1167),.dout(w_dff_B_s9KZOleJ3_1),.clk(gclk));
	jdff dff_B_lnZdkdhu8_2(.din(n1068),.dout(w_dff_B_lnZdkdhu8_2),.clk(gclk));
	jdff dff_B_3uOXyjC45_2(.din(w_dff_B_lnZdkdhu8_2),.dout(w_dff_B_3uOXyjC45_2),.clk(gclk));
	jdff dff_B_XSQuYT9H0_2(.din(w_dff_B_3uOXyjC45_2),.dout(w_dff_B_XSQuYT9H0_2),.clk(gclk));
	jdff dff_B_1IHjAhvv0_2(.din(w_dff_B_XSQuYT9H0_2),.dout(w_dff_B_1IHjAhvv0_2),.clk(gclk));
	jdff dff_B_rJYqr7oy9_2(.din(w_dff_B_1IHjAhvv0_2),.dout(w_dff_B_rJYqr7oy9_2),.clk(gclk));
	jdff dff_B_YUxIifb32_2(.din(w_dff_B_rJYqr7oy9_2),.dout(w_dff_B_YUxIifb32_2),.clk(gclk));
	jdff dff_B_NcDSgTR24_2(.din(w_dff_B_YUxIifb32_2),.dout(w_dff_B_NcDSgTR24_2),.clk(gclk));
	jdff dff_B_21N4drx09_2(.din(w_dff_B_NcDSgTR24_2),.dout(w_dff_B_21N4drx09_2),.clk(gclk));
	jdff dff_B_kFATyO175_2(.din(w_dff_B_21N4drx09_2),.dout(w_dff_B_kFATyO175_2),.clk(gclk));
	jdff dff_B_zUtO91ct9_2(.din(w_dff_B_kFATyO175_2),.dout(w_dff_B_zUtO91ct9_2),.clk(gclk));
	jdff dff_B_BcBRBhx66_2(.din(w_dff_B_zUtO91ct9_2),.dout(w_dff_B_BcBRBhx66_2),.clk(gclk));
	jdff dff_B_96nKsbR15_2(.din(w_dff_B_BcBRBhx66_2),.dout(w_dff_B_96nKsbR15_2),.clk(gclk));
	jdff dff_B_axJgrRFr3_2(.din(w_dff_B_96nKsbR15_2),.dout(w_dff_B_axJgrRFr3_2),.clk(gclk));
	jdff dff_B_PrtgEQao9_2(.din(w_dff_B_axJgrRFr3_2),.dout(w_dff_B_PrtgEQao9_2),.clk(gclk));
	jdff dff_B_4OQ3Tr7o3_2(.din(n1085),.dout(w_dff_B_4OQ3Tr7o3_2),.clk(gclk));
	jdff dff_B_JEKq79lb7_1(.din(n1069),.dout(w_dff_B_JEKq79lb7_1),.clk(gclk));
	jdff dff_B_7qVTZSt23_2(.din(n969),.dout(w_dff_B_7qVTZSt23_2),.clk(gclk));
	jdff dff_B_x4LXLFhz1_2(.din(w_dff_B_7qVTZSt23_2),.dout(w_dff_B_x4LXLFhz1_2),.clk(gclk));
	jdff dff_B_vkMs8pXZ9_2(.din(w_dff_B_x4LXLFhz1_2),.dout(w_dff_B_vkMs8pXZ9_2),.clk(gclk));
	jdff dff_B_YP3WyDY45_2(.din(w_dff_B_vkMs8pXZ9_2),.dout(w_dff_B_YP3WyDY45_2),.clk(gclk));
	jdff dff_B_5dYUpLsq5_2(.din(w_dff_B_YP3WyDY45_2),.dout(w_dff_B_5dYUpLsq5_2),.clk(gclk));
	jdff dff_B_1Kun2Lk55_2(.din(w_dff_B_5dYUpLsq5_2),.dout(w_dff_B_1Kun2Lk55_2),.clk(gclk));
	jdff dff_B_FOpswNle6_2(.din(w_dff_B_1Kun2Lk55_2),.dout(w_dff_B_FOpswNle6_2),.clk(gclk));
	jdff dff_B_19sugaSe5_2(.din(w_dff_B_FOpswNle6_2),.dout(w_dff_B_19sugaSe5_2),.clk(gclk));
	jdff dff_B_YZjIsvaf6_2(.din(w_dff_B_19sugaSe5_2),.dout(w_dff_B_YZjIsvaf6_2),.clk(gclk));
	jdff dff_B_1zRM0Uim6_2(.din(w_dff_B_YZjIsvaf6_2),.dout(w_dff_B_1zRM0Uim6_2),.clk(gclk));
	jdff dff_B_jri7Ub2C6_2(.din(w_dff_B_1zRM0Uim6_2),.dout(w_dff_B_jri7Ub2C6_2),.clk(gclk));
	jdff dff_B_KpAjid0A5_2(.din(n986),.dout(w_dff_B_KpAjid0A5_2),.clk(gclk));
	jdff dff_B_XDYSzb834_1(.din(n970),.dout(w_dff_B_XDYSzb834_1),.clk(gclk));
	jdff dff_B_zpKd6K8c6_2(.din(n867),.dout(w_dff_B_zpKd6K8c6_2),.clk(gclk));
	jdff dff_B_pHrcQcCv0_2(.din(w_dff_B_zpKd6K8c6_2),.dout(w_dff_B_pHrcQcCv0_2),.clk(gclk));
	jdff dff_B_lUwl4kVV6_2(.din(w_dff_B_pHrcQcCv0_2),.dout(w_dff_B_lUwl4kVV6_2),.clk(gclk));
	jdff dff_B_MvZZh7PX7_2(.din(w_dff_B_lUwl4kVV6_2),.dout(w_dff_B_MvZZh7PX7_2),.clk(gclk));
	jdff dff_B_DbUaWsD48_2(.din(w_dff_B_MvZZh7PX7_2),.dout(w_dff_B_DbUaWsD48_2),.clk(gclk));
	jdff dff_B_qniCvI2i3_2(.din(w_dff_B_DbUaWsD48_2),.dout(w_dff_B_qniCvI2i3_2),.clk(gclk));
	jdff dff_B_Acp5b3Kh4_2(.din(w_dff_B_qniCvI2i3_2),.dout(w_dff_B_Acp5b3Kh4_2),.clk(gclk));
	jdff dff_B_EXMcD6pc9_2(.din(w_dff_B_Acp5b3Kh4_2),.dout(w_dff_B_EXMcD6pc9_2),.clk(gclk));
	jdff dff_B_xP5YrImD0_2(.din(n880),.dout(w_dff_B_xP5YrImD0_2),.clk(gclk));
	jdff dff_B_XTmIjNuN8_2(.din(w_dff_B_xP5YrImD0_2),.dout(w_dff_B_XTmIjNuN8_2),.clk(gclk));
	jdff dff_B_5wJlXDlD9_2(.din(w_dff_B_XTmIjNuN8_2),.dout(w_dff_B_5wJlXDlD9_2),.clk(gclk));
	jdff dff_B_et0YoBfi1_1(.din(n868),.dout(w_dff_B_et0YoBfi1_1),.clk(gclk));
	jdff dff_B_Rx5fQxCb1_1(.din(w_dff_B_et0YoBfi1_1),.dout(w_dff_B_Rx5fQxCb1_1),.clk(gclk));
	jdff dff_B_3tgqI8hW8_2(.din(n771),.dout(w_dff_B_3tgqI8hW8_2),.clk(gclk));
	jdff dff_B_7TqT456q7_2(.din(w_dff_B_3tgqI8hW8_2),.dout(w_dff_B_7TqT456q7_2),.clk(gclk));
	jdff dff_B_wYrutqXZ8_2(.din(w_dff_B_7TqT456q7_2),.dout(w_dff_B_wYrutqXZ8_2),.clk(gclk));
	jdff dff_B_scAyxHrg4_0(.din(n776),.dout(w_dff_B_scAyxHrg4_0),.clk(gclk));
	jdff dff_A_Ehqss91C2_0(.dout(w_n676_0[0]),.din(w_dff_A_Ehqss91C2_0),.clk(gclk));
	jdff dff_A_96WjFtJZ9_0(.dout(w_dff_A_Ehqss91C2_0),.din(w_dff_A_96WjFtJZ9_0),.clk(gclk));
	jdff dff_A_vxfMr52P9_1(.dout(w_n676_0[1]),.din(w_dff_A_vxfMr52P9_1),.clk(gclk));
	jdff dff_A_z1Kp4bwm6_1(.dout(w_dff_A_vxfMr52P9_1),.din(w_dff_A_z1Kp4bwm6_1),.clk(gclk));
	jdff dff_B_jsicA2br8_1(.din(n1812),.dout(w_dff_B_jsicA2br8_1),.clk(gclk));
	jdff dff_B_EqsQe0zZ2_1(.din(n1799),.dout(w_dff_B_EqsQe0zZ2_1),.clk(gclk));
	jdff dff_B_SQb1nkqy3_1(.din(w_dff_B_EqsQe0zZ2_1),.dout(w_dff_B_SQb1nkqy3_1),.clk(gclk));
	jdff dff_B_0ZC1Rhkb4_2(.din(n1798),.dout(w_dff_B_0ZC1Rhkb4_2),.clk(gclk));
	jdff dff_B_b9bKABFx3_2(.din(w_dff_B_0ZC1Rhkb4_2),.dout(w_dff_B_b9bKABFx3_2),.clk(gclk));
	jdff dff_B_v16KuXGp9_2(.din(w_dff_B_b9bKABFx3_2),.dout(w_dff_B_v16KuXGp9_2),.clk(gclk));
	jdff dff_B_wAqBbolL7_2(.din(w_dff_B_v16KuXGp9_2),.dout(w_dff_B_wAqBbolL7_2),.clk(gclk));
	jdff dff_B_Mq6sI9D28_2(.din(w_dff_B_wAqBbolL7_2),.dout(w_dff_B_Mq6sI9D28_2),.clk(gclk));
	jdff dff_B_HfCZ0BMs4_2(.din(w_dff_B_Mq6sI9D28_2),.dout(w_dff_B_HfCZ0BMs4_2),.clk(gclk));
	jdff dff_B_T9QlhBoH0_2(.din(w_dff_B_HfCZ0BMs4_2),.dout(w_dff_B_T9QlhBoH0_2),.clk(gclk));
	jdff dff_B_5bFb3YYt0_2(.din(w_dff_B_T9QlhBoH0_2),.dout(w_dff_B_5bFb3YYt0_2),.clk(gclk));
	jdff dff_B_CHTigQ4K6_2(.din(w_dff_B_5bFb3YYt0_2),.dout(w_dff_B_CHTigQ4K6_2),.clk(gclk));
	jdff dff_B_E1mwLwzD3_2(.din(w_dff_B_CHTigQ4K6_2),.dout(w_dff_B_E1mwLwzD3_2),.clk(gclk));
	jdff dff_B_KBkld3fv6_2(.din(w_dff_B_E1mwLwzD3_2),.dout(w_dff_B_KBkld3fv6_2),.clk(gclk));
	jdff dff_B_eyyxhrH93_2(.din(w_dff_B_KBkld3fv6_2),.dout(w_dff_B_eyyxhrH93_2),.clk(gclk));
	jdff dff_B_ViIgY6qx5_2(.din(w_dff_B_eyyxhrH93_2),.dout(w_dff_B_ViIgY6qx5_2),.clk(gclk));
	jdff dff_B_PSjB8nIS1_2(.din(w_dff_B_ViIgY6qx5_2),.dout(w_dff_B_PSjB8nIS1_2),.clk(gclk));
	jdff dff_B_BRTnTT3k5_2(.din(w_dff_B_PSjB8nIS1_2),.dout(w_dff_B_BRTnTT3k5_2),.clk(gclk));
	jdff dff_B_orq0XXey8_2(.din(w_dff_B_BRTnTT3k5_2),.dout(w_dff_B_orq0XXey8_2),.clk(gclk));
	jdff dff_B_w5otUtWB7_2(.din(w_dff_B_orq0XXey8_2),.dout(w_dff_B_w5otUtWB7_2),.clk(gclk));
	jdff dff_B_WvWMk6WC9_2(.din(w_dff_B_w5otUtWB7_2),.dout(w_dff_B_WvWMk6WC9_2),.clk(gclk));
	jdff dff_B_dKREafO36_2(.din(w_dff_B_WvWMk6WC9_2),.dout(w_dff_B_dKREafO36_2),.clk(gclk));
	jdff dff_B_1gzraluq6_2(.din(w_dff_B_dKREafO36_2),.dout(w_dff_B_1gzraluq6_2),.clk(gclk));
	jdff dff_B_AJVUYrpd2_2(.din(w_dff_B_1gzraluq6_2),.dout(w_dff_B_AJVUYrpd2_2),.clk(gclk));
	jdff dff_B_U6GHPRTR5_2(.din(w_dff_B_AJVUYrpd2_2),.dout(w_dff_B_U6GHPRTR5_2),.clk(gclk));
	jdff dff_B_ljxAg85k1_2(.din(w_dff_B_U6GHPRTR5_2),.dout(w_dff_B_ljxAg85k1_2),.clk(gclk));
	jdff dff_B_vELiSrbG3_2(.din(w_dff_B_ljxAg85k1_2),.dout(w_dff_B_vELiSrbG3_2),.clk(gclk));
	jdff dff_B_N6RIcCje6_2(.din(w_dff_B_vELiSrbG3_2),.dout(w_dff_B_N6RIcCje6_2),.clk(gclk));
	jdff dff_B_0AYq1ozq9_2(.din(w_dff_B_N6RIcCje6_2),.dout(w_dff_B_0AYq1ozq9_2),.clk(gclk));
	jdff dff_B_DhlcXIkj0_2(.din(w_dff_B_0AYq1ozq9_2),.dout(w_dff_B_DhlcXIkj0_2),.clk(gclk));
	jdff dff_B_rK11GMSa2_2(.din(w_dff_B_DhlcXIkj0_2),.dout(w_dff_B_rK11GMSa2_2),.clk(gclk));
	jdff dff_B_PZ38W6Yx2_2(.din(w_dff_B_rK11GMSa2_2),.dout(w_dff_B_PZ38W6Yx2_2),.clk(gclk));
	jdff dff_B_yjgVH1fF0_2(.din(w_dff_B_PZ38W6Yx2_2),.dout(w_dff_B_yjgVH1fF0_2),.clk(gclk));
	jdff dff_B_Au7sQFSe9_2(.din(w_dff_B_yjgVH1fF0_2),.dout(w_dff_B_Au7sQFSe9_2),.clk(gclk));
	jdff dff_B_IQtbwsbQ9_2(.din(w_dff_B_Au7sQFSe9_2),.dout(w_dff_B_IQtbwsbQ9_2),.clk(gclk));
	jdff dff_B_ZnVnleM24_2(.din(w_dff_B_IQtbwsbQ9_2),.dout(w_dff_B_ZnVnleM24_2),.clk(gclk));
	jdff dff_B_FhLgab0R5_2(.din(w_dff_B_ZnVnleM24_2),.dout(w_dff_B_FhLgab0R5_2),.clk(gclk));
	jdff dff_B_RmOZQAAW1_2(.din(w_dff_B_FhLgab0R5_2),.dout(w_dff_B_RmOZQAAW1_2),.clk(gclk));
	jdff dff_B_mcoHI9228_2(.din(w_dff_B_RmOZQAAW1_2),.dout(w_dff_B_mcoHI9228_2),.clk(gclk));
	jdff dff_B_nu9yuFi28_2(.din(w_dff_B_mcoHI9228_2),.dout(w_dff_B_nu9yuFi28_2),.clk(gclk));
	jdff dff_B_57nUGVQH7_2(.din(w_dff_B_nu9yuFi28_2),.dout(w_dff_B_57nUGVQH7_2),.clk(gclk));
	jdff dff_B_WZVjoAz74_2(.din(w_dff_B_57nUGVQH7_2),.dout(w_dff_B_WZVjoAz74_2),.clk(gclk));
	jdff dff_B_Dj8wHJUw3_2(.din(w_dff_B_WZVjoAz74_2),.dout(w_dff_B_Dj8wHJUw3_2),.clk(gclk));
	jdff dff_B_CxuOwJ9T4_2(.din(w_dff_B_Dj8wHJUw3_2),.dout(w_dff_B_CxuOwJ9T4_2),.clk(gclk));
	jdff dff_B_YE5usB9l5_2(.din(w_dff_B_CxuOwJ9T4_2),.dout(w_dff_B_YE5usB9l5_2),.clk(gclk));
	jdff dff_B_MaLZ22Bi4_2(.din(w_dff_B_YE5usB9l5_2),.dout(w_dff_B_MaLZ22Bi4_2),.clk(gclk));
	jdff dff_B_0vlqLkWt1_2(.din(w_dff_B_MaLZ22Bi4_2),.dout(w_dff_B_0vlqLkWt1_2),.clk(gclk));
	jdff dff_B_yF9Xkmon8_2(.din(w_dff_B_0vlqLkWt1_2),.dout(w_dff_B_yF9Xkmon8_2),.clk(gclk));
	jdff dff_B_oQREDpah4_2(.din(w_dff_B_yF9Xkmon8_2),.dout(w_dff_B_oQREDpah4_2),.clk(gclk));
	jdff dff_B_3bykjGzj4_2(.din(w_dff_B_oQREDpah4_2),.dout(w_dff_B_3bykjGzj4_2),.clk(gclk));
	jdff dff_B_olshoiTp9_2(.din(w_dff_B_3bykjGzj4_2),.dout(w_dff_B_olshoiTp9_2),.clk(gclk));
	jdff dff_B_HKO57Efn9_2(.din(w_dff_B_olshoiTp9_2),.dout(w_dff_B_HKO57Efn9_2),.clk(gclk));
	jdff dff_B_ngOwxPRj8_2(.din(w_dff_B_HKO57Efn9_2),.dout(w_dff_B_ngOwxPRj8_2),.clk(gclk));
	jdff dff_B_ez7O8DKz6_2(.din(w_dff_B_ngOwxPRj8_2),.dout(w_dff_B_ez7O8DKz6_2),.clk(gclk));
	jdff dff_B_CJrNqhDw9_2(.din(w_dff_B_ez7O8DKz6_2),.dout(w_dff_B_CJrNqhDw9_2),.clk(gclk));
	jdff dff_B_Yqe5obyU9_2(.din(w_dff_B_CJrNqhDw9_2),.dout(w_dff_B_Yqe5obyU9_2),.clk(gclk));
	jdff dff_B_MUkFS5jG6_2(.din(n1797),.dout(w_dff_B_MUkFS5jG6_2),.clk(gclk));
	jdff dff_B_OGwC6Rvn1_2(.din(w_dff_B_MUkFS5jG6_2),.dout(w_dff_B_OGwC6Rvn1_2),.clk(gclk));
	jdff dff_B_gUFxVDau1_2(.din(w_dff_B_OGwC6Rvn1_2),.dout(w_dff_B_gUFxVDau1_2),.clk(gclk));
	jdff dff_B_YCYUCBC63_2(.din(w_dff_B_gUFxVDau1_2),.dout(w_dff_B_YCYUCBC63_2),.clk(gclk));
	jdff dff_B_MDn3ANsS2_2(.din(w_dff_B_YCYUCBC63_2),.dout(w_dff_B_MDn3ANsS2_2),.clk(gclk));
	jdff dff_B_KJ8cCYY08_2(.din(w_dff_B_MDn3ANsS2_2),.dout(w_dff_B_KJ8cCYY08_2),.clk(gclk));
	jdff dff_B_TKVh6Ytz4_2(.din(w_dff_B_KJ8cCYY08_2),.dout(w_dff_B_TKVh6Ytz4_2),.clk(gclk));
	jdff dff_B_4liTS6k20_2(.din(w_dff_B_TKVh6Ytz4_2),.dout(w_dff_B_4liTS6k20_2),.clk(gclk));
	jdff dff_B_eOR086B22_2(.din(w_dff_B_4liTS6k20_2),.dout(w_dff_B_eOR086B22_2),.clk(gclk));
	jdff dff_B_Hvgmn9CN1_2(.din(w_dff_B_eOR086B22_2),.dout(w_dff_B_Hvgmn9CN1_2),.clk(gclk));
	jdff dff_B_gQPX1R127_2(.din(w_dff_B_Hvgmn9CN1_2),.dout(w_dff_B_gQPX1R127_2),.clk(gclk));
	jdff dff_B_bAiX3mxd1_2(.din(w_dff_B_gQPX1R127_2),.dout(w_dff_B_bAiX3mxd1_2),.clk(gclk));
	jdff dff_B_9QjRRC6G0_2(.din(w_dff_B_bAiX3mxd1_2),.dout(w_dff_B_9QjRRC6G0_2),.clk(gclk));
	jdff dff_B_iYUtJfo63_2(.din(w_dff_B_9QjRRC6G0_2),.dout(w_dff_B_iYUtJfo63_2),.clk(gclk));
	jdff dff_B_BEjzN3Tk8_2(.din(w_dff_B_iYUtJfo63_2),.dout(w_dff_B_BEjzN3Tk8_2),.clk(gclk));
	jdff dff_B_oPkqVb122_2(.din(w_dff_B_BEjzN3Tk8_2),.dout(w_dff_B_oPkqVb122_2),.clk(gclk));
	jdff dff_B_ybM8yBJc6_2(.din(w_dff_B_oPkqVb122_2),.dout(w_dff_B_ybM8yBJc6_2),.clk(gclk));
	jdff dff_B_AwW3Li6B4_2(.din(w_dff_B_ybM8yBJc6_2),.dout(w_dff_B_AwW3Li6B4_2),.clk(gclk));
	jdff dff_B_wDiSjjVo0_2(.din(w_dff_B_AwW3Li6B4_2),.dout(w_dff_B_wDiSjjVo0_2),.clk(gclk));
	jdff dff_B_IDfo7be52_2(.din(w_dff_B_wDiSjjVo0_2),.dout(w_dff_B_IDfo7be52_2),.clk(gclk));
	jdff dff_B_v6NPQO604_2(.din(w_dff_B_IDfo7be52_2),.dout(w_dff_B_v6NPQO604_2),.clk(gclk));
	jdff dff_B_oM8ZydWC4_2(.din(w_dff_B_v6NPQO604_2),.dout(w_dff_B_oM8ZydWC4_2),.clk(gclk));
	jdff dff_B_7gmdIUcN3_2(.din(w_dff_B_oM8ZydWC4_2),.dout(w_dff_B_7gmdIUcN3_2),.clk(gclk));
	jdff dff_B_VJn4hN5I0_2(.din(w_dff_B_7gmdIUcN3_2),.dout(w_dff_B_VJn4hN5I0_2),.clk(gclk));
	jdff dff_B_ywgb2ue65_2(.din(w_dff_B_VJn4hN5I0_2),.dout(w_dff_B_ywgb2ue65_2),.clk(gclk));
	jdff dff_B_AhWO7RTD7_2(.din(w_dff_B_ywgb2ue65_2),.dout(w_dff_B_AhWO7RTD7_2),.clk(gclk));
	jdff dff_B_dee6IbdF6_2(.din(w_dff_B_AhWO7RTD7_2),.dout(w_dff_B_dee6IbdF6_2),.clk(gclk));
	jdff dff_B_0sTGuZlx4_2(.din(w_dff_B_dee6IbdF6_2),.dout(w_dff_B_0sTGuZlx4_2),.clk(gclk));
	jdff dff_B_U15bZJxy9_2(.din(w_dff_B_0sTGuZlx4_2),.dout(w_dff_B_U15bZJxy9_2),.clk(gclk));
	jdff dff_B_CBzR9XnT5_2(.din(w_dff_B_U15bZJxy9_2),.dout(w_dff_B_CBzR9XnT5_2),.clk(gclk));
	jdff dff_B_hjGEk3FN1_2(.din(w_dff_B_CBzR9XnT5_2),.dout(w_dff_B_hjGEk3FN1_2),.clk(gclk));
	jdff dff_B_UwDtDREG3_2(.din(w_dff_B_hjGEk3FN1_2),.dout(w_dff_B_UwDtDREG3_2),.clk(gclk));
	jdff dff_B_eo8weaP44_2(.din(w_dff_B_UwDtDREG3_2),.dout(w_dff_B_eo8weaP44_2),.clk(gclk));
	jdff dff_B_kugiXiML7_2(.din(w_dff_B_eo8weaP44_2),.dout(w_dff_B_kugiXiML7_2),.clk(gclk));
	jdff dff_B_XGFTtA0G2_2(.din(w_dff_B_kugiXiML7_2),.dout(w_dff_B_XGFTtA0G2_2),.clk(gclk));
	jdff dff_B_KI8OEpS27_2(.din(w_dff_B_XGFTtA0G2_2),.dout(w_dff_B_KI8OEpS27_2),.clk(gclk));
	jdff dff_B_YM4G7ZiF1_2(.din(w_dff_B_KI8OEpS27_2),.dout(w_dff_B_YM4G7ZiF1_2),.clk(gclk));
	jdff dff_B_zwpbgDYE5_2(.din(w_dff_B_YM4G7ZiF1_2),.dout(w_dff_B_zwpbgDYE5_2),.clk(gclk));
	jdff dff_B_XtfTWcjP3_2(.din(w_dff_B_zwpbgDYE5_2),.dout(w_dff_B_XtfTWcjP3_2),.clk(gclk));
	jdff dff_B_czZGDbNt3_2(.din(w_dff_B_XtfTWcjP3_2),.dout(w_dff_B_czZGDbNt3_2),.clk(gclk));
	jdff dff_B_UsjuP7vh9_2(.din(w_dff_B_czZGDbNt3_2),.dout(w_dff_B_UsjuP7vh9_2),.clk(gclk));
	jdff dff_B_dVmPfubU1_2(.din(w_dff_B_UsjuP7vh9_2),.dout(w_dff_B_dVmPfubU1_2),.clk(gclk));
	jdff dff_B_4QP4v6QC2_2(.din(w_dff_B_dVmPfubU1_2),.dout(w_dff_B_4QP4v6QC2_2),.clk(gclk));
	jdff dff_B_u7vexqQJ7_2(.din(w_dff_B_4QP4v6QC2_2),.dout(w_dff_B_u7vexqQJ7_2),.clk(gclk));
	jdff dff_B_vwqbKnIa1_2(.din(w_dff_B_u7vexqQJ7_2),.dout(w_dff_B_vwqbKnIa1_2),.clk(gclk));
	jdff dff_B_hbIAKUDn3_2(.din(w_dff_B_vwqbKnIa1_2),.dout(w_dff_B_hbIAKUDn3_2),.clk(gclk));
	jdff dff_B_9xf7aOe23_2(.din(w_dff_B_hbIAKUDn3_2),.dout(w_dff_B_9xf7aOe23_2),.clk(gclk));
	jdff dff_B_Lh8zPf0H3_2(.din(w_dff_B_9xf7aOe23_2),.dout(w_dff_B_Lh8zPf0H3_2),.clk(gclk));
	jdff dff_B_z7Oi3qKz3_2(.din(w_dff_B_Lh8zPf0H3_2),.dout(w_dff_B_z7Oi3qKz3_2),.clk(gclk));
	jdff dff_B_mJTxB75M7_2(.din(w_dff_B_z7Oi3qKz3_2),.dout(w_dff_B_mJTxB75M7_2),.clk(gclk));
	jdff dff_B_GiZa1NzW1_2(.din(w_dff_B_mJTxB75M7_2),.dout(w_dff_B_GiZa1NzW1_2),.clk(gclk));
	jdff dff_B_dTjgFn7P7_2(.din(w_dff_B_GiZa1NzW1_2),.dout(w_dff_B_dTjgFn7P7_2),.clk(gclk));
	jdff dff_B_lMh2uqU83_2(.din(w_dff_B_dTjgFn7P7_2),.dout(w_dff_B_lMh2uqU83_2),.clk(gclk));
	jdff dff_B_bQhuycTN1_2(.din(w_dff_B_lMh2uqU83_2),.dout(w_dff_B_bQhuycTN1_2),.clk(gclk));
	jdff dff_B_hAmTZHFN2_2(.din(w_dff_B_bQhuycTN1_2),.dout(w_dff_B_hAmTZHFN2_2),.clk(gclk));
	jdff dff_A_WUTJTKWd2_1(.dout(w_n1796_0[1]),.din(w_dff_A_WUTJTKWd2_1),.clk(gclk));
	jdff dff_B_wGgdgUrc1_1(.din(n1794),.dout(w_dff_B_wGgdgUrc1_1),.clk(gclk));
	jdff dff_B_sCeb9wVt9_2(.din(n1772),.dout(w_dff_B_sCeb9wVt9_2),.clk(gclk));
	jdff dff_B_ylhITx530_2(.din(w_dff_B_sCeb9wVt9_2),.dout(w_dff_B_ylhITx530_2),.clk(gclk));
	jdff dff_B_WjBnJe5F8_2(.din(w_dff_B_ylhITx530_2),.dout(w_dff_B_WjBnJe5F8_2),.clk(gclk));
	jdff dff_B_Gg7w9Nh92_2(.din(w_dff_B_WjBnJe5F8_2),.dout(w_dff_B_Gg7w9Nh92_2),.clk(gclk));
	jdff dff_B_Tvph5wDM4_2(.din(w_dff_B_Gg7w9Nh92_2),.dout(w_dff_B_Tvph5wDM4_2),.clk(gclk));
	jdff dff_B_dPZPOFDB6_2(.din(w_dff_B_Tvph5wDM4_2),.dout(w_dff_B_dPZPOFDB6_2),.clk(gclk));
	jdff dff_B_vnzkRU5m8_2(.din(w_dff_B_dPZPOFDB6_2),.dout(w_dff_B_vnzkRU5m8_2),.clk(gclk));
	jdff dff_B_9c3FrUCK4_2(.din(w_dff_B_vnzkRU5m8_2),.dout(w_dff_B_9c3FrUCK4_2),.clk(gclk));
	jdff dff_B_C2GU6Yls0_2(.din(w_dff_B_9c3FrUCK4_2),.dout(w_dff_B_C2GU6Yls0_2),.clk(gclk));
	jdff dff_B_Lu3HTxUo6_2(.din(w_dff_B_C2GU6Yls0_2),.dout(w_dff_B_Lu3HTxUo6_2),.clk(gclk));
	jdff dff_B_j23Qzexu3_2(.din(w_dff_B_Lu3HTxUo6_2),.dout(w_dff_B_j23Qzexu3_2),.clk(gclk));
	jdff dff_B_1wzHLvu67_2(.din(w_dff_B_j23Qzexu3_2),.dout(w_dff_B_1wzHLvu67_2),.clk(gclk));
	jdff dff_B_kyItvtrt4_2(.din(w_dff_B_1wzHLvu67_2),.dout(w_dff_B_kyItvtrt4_2),.clk(gclk));
	jdff dff_B_SvUP6WzU9_2(.din(w_dff_B_kyItvtrt4_2),.dout(w_dff_B_SvUP6WzU9_2),.clk(gclk));
	jdff dff_B_nEcOhYSY9_2(.din(w_dff_B_SvUP6WzU9_2),.dout(w_dff_B_nEcOhYSY9_2),.clk(gclk));
	jdff dff_B_VGjiVPLY7_2(.din(w_dff_B_nEcOhYSY9_2),.dout(w_dff_B_VGjiVPLY7_2),.clk(gclk));
	jdff dff_B_KQWCpyzV0_2(.din(w_dff_B_VGjiVPLY7_2),.dout(w_dff_B_KQWCpyzV0_2),.clk(gclk));
	jdff dff_B_LB2brG6O6_2(.din(w_dff_B_KQWCpyzV0_2),.dout(w_dff_B_LB2brG6O6_2),.clk(gclk));
	jdff dff_B_mI1Zg0cW1_2(.din(w_dff_B_LB2brG6O6_2),.dout(w_dff_B_mI1Zg0cW1_2),.clk(gclk));
	jdff dff_B_OXIrjBbR2_2(.din(w_dff_B_mI1Zg0cW1_2),.dout(w_dff_B_OXIrjBbR2_2),.clk(gclk));
	jdff dff_B_g7im5osU3_2(.din(w_dff_B_OXIrjBbR2_2),.dout(w_dff_B_g7im5osU3_2),.clk(gclk));
	jdff dff_B_BHDgTPr90_2(.din(w_dff_B_g7im5osU3_2),.dout(w_dff_B_BHDgTPr90_2),.clk(gclk));
	jdff dff_B_J8HDxvDj5_2(.din(w_dff_B_BHDgTPr90_2),.dout(w_dff_B_J8HDxvDj5_2),.clk(gclk));
	jdff dff_B_DRquSYQP2_2(.din(w_dff_B_J8HDxvDj5_2),.dout(w_dff_B_DRquSYQP2_2),.clk(gclk));
	jdff dff_B_UFQstv0P5_2(.din(w_dff_B_DRquSYQP2_2),.dout(w_dff_B_UFQstv0P5_2),.clk(gclk));
	jdff dff_B_NiRYfbKi4_2(.din(w_dff_B_UFQstv0P5_2),.dout(w_dff_B_NiRYfbKi4_2),.clk(gclk));
	jdff dff_B_071mX1x89_2(.din(w_dff_B_NiRYfbKi4_2),.dout(w_dff_B_071mX1x89_2),.clk(gclk));
	jdff dff_B_7yCmUlGK8_2(.din(w_dff_B_071mX1x89_2),.dout(w_dff_B_7yCmUlGK8_2),.clk(gclk));
	jdff dff_B_3ZGp1siw2_2(.din(w_dff_B_7yCmUlGK8_2),.dout(w_dff_B_3ZGp1siw2_2),.clk(gclk));
	jdff dff_B_cuQKHB7k7_2(.din(w_dff_B_3ZGp1siw2_2),.dout(w_dff_B_cuQKHB7k7_2),.clk(gclk));
	jdff dff_B_FZ78vUyu4_2(.din(w_dff_B_cuQKHB7k7_2),.dout(w_dff_B_FZ78vUyu4_2),.clk(gclk));
	jdff dff_B_70P1lBrn5_2(.din(w_dff_B_FZ78vUyu4_2),.dout(w_dff_B_70P1lBrn5_2),.clk(gclk));
	jdff dff_B_wlbwh8KZ7_2(.din(w_dff_B_70P1lBrn5_2),.dout(w_dff_B_wlbwh8KZ7_2),.clk(gclk));
	jdff dff_B_iBMZxMjk1_2(.din(w_dff_B_wlbwh8KZ7_2),.dout(w_dff_B_iBMZxMjk1_2),.clk(gclk));
	jdff dff_B_mr4jFSFb6_2(.din(w_dff_B_iBMZxMjk1_2),.dout(w_dff_B_mr4jFSFb6_2),.clk(gclk));
	jdff dff_B_ui9HzCMJ7_2(.din(w_dff_B_mr4jFSFb6_2),.dout(w_dff_B_ui9HzCMJ7_2),.clk(gclk));
	jdff dff_B_t5Kw2i9u2_2(.din(w_dff_B_ui9HzCMJ7_2),.dout(w_dff_B_t5Kw2i9u2_2),.clk(gclk));
	jdff dff_B_NSouHv6q5_2(.din(w_dff_B_t5Kw2i9u2_2),.dout(w_dff_B_NSouHv6q5_2),.clk(gclk));
	jdff dff_B_gXo3zGkQ7_2(.din(w_dff_B_NSouHv6q5_2),.dout(w_dff_B_gXo3zGkQ7_2),.clk(gclk));
	jdff dff_B_Ynzsrzsp4_2(.din(w_dff_B_gXo3zGkQ7_2),.dout(w_dff_B_Ynzsrzsp4_2),.clk(gclk));
	jdff dff_B_3cnBLrxN6_2(.din(w_dff_B_Ynzsrzsp4_2),.dout(w_dff_B_3cnBLrxN6_2),.clk(gclk));
	jdff dff_B_VLdoh07G5_2(.din(w_dff_B_3cnBLrxN6_2),.dout(w_dff_B_VLdoh07G5_2),.clk(gclk));
	jdff dff_B_ZHJi1bYo6_2(.din(w_dff_B_VLdoh07G5_2),.dout(w_dff_B_ZHJi1bYo6_2),.clk(gclk));
	jdff dff_B_SXcydJgu3_2(.din(w_dff_B_ZHJi1bYo6_2),.dout(w_dff_B_SXcydJgu3_2),.clk(gclk));
	jdff dff_B_tWmGSrej7_2(.din(w_dff_B_SXcydJgu3_2),.dout(w_dff_B_tWmGSrej7_2),.clk(gclk));
	jdff dff_B_2lda7fOH1_2(.din(w_dff_B_tWmGSrej7_2),.dout(w_dff_B_2lda7fOH1_2),.clk(gclk));
	jdff dff_B_e867UfEX2_2(.din(w_dff_B_2lda7fOH1_2),.dout(w_dff_B_e867UfEX2_2),.clk(gclk));
	jdff dff_B_0cqTYGmW5_2(.din(w_dff_B_e867UfEX2_2),.dout(w_dff_B_0cqTYGmW5_2),.clk(gclk));
	jdff dff_B_CLZacbvV3_2(.din(w_dff_B_0cqTYGmW5_2),.dout(w_dff_B_CLZacbvV3_2),.clk(gclk));
	jdff dff_B_ygypAn457_2(.din(w_dff_B_CLZacbvV3_2),.dout(w_dff_B_ygypAn457_2),.clk(gclk));
	jdff dff_B_hWcQC6fp4_2(.din(w_dff_B_ygypAn457_2),.dout(w_dff_B_hWcQC6fp4_2),.clk(gclk));
	jdff dff_B_85nnEfjK5_2(.din(w_dff_B_hWcQC6fp4_2),.dout(w_dff_B_85nnEfjK5_2),.clk(gclk));
	jdff dff_B_W6rnKeD31_1(.din(n1778),.dout(w_dff_B_W6rnKeD31_1),.clk(gclk));
	jdff dff_B_RZnj8RYO2_1(.din(w_dff_B_W6rnKeD31_1),.dout(w_dff_B_RZnj8RYO2_1),.clk(gclk));
	jdff dff_B_2J865Ohu3_2(.din(n1777),.dout(w_dff_B_2J865Ohu3_2),.clk(gclk));
	jdff dff_B_HVZ3fHA36_2(.din(w_dff_B_2J865Ohu3_2),.dout(w_dff_B_HVZ3fHA36_2),.clk(gclk));
	jdff dff_B_TqHM9f793_2(.din(w_dff_B_HVZ3fHA36_2),.dout(w_dff_B_TqHM9f793_2),.clk(gclk));
	jdff dff_B_K8tauUjq6_2(.din(w_dff_B_TqHM9f793_2),.dout(w_dff_B_K8tauUjq6_2),.clk(gclk));
	jdff dff_B_7O5ZcEF10_2(.din(w_dff_B_K8tauUjq6_2),.dout(w_dff_B_7O5ZcEF10_2),.clk(gclk));
	jdff dff_B_4O5C7DOo9_2(.din(w_dff_B_7O5ZcEF10_2),.dout(w_dff_B_4O5C7DOo9_2),.clk(gclk));
	jdff dff_B_MbmSYfdq3_2(.din(w_dff_B_4O5C7DOo9_2),.dout(w_dff_B_MbmSYfdq3_2),.clk(gclk));
	jdff dff_B_8ZHRrLpp7_2(.din(w_dff_B_MbmSYfdq3_2),.dout(w_dff_B_8ZHRrLpp7_2),.clk(gclk));
	jdff dff_B_nth6Zzm01_2(.din(w_dff_B_8ZHRrLpp7_2),.dout(w_dff_B_nth6Zzm01_2),.clk(gclk));
	jdff dff_B_ZBCUt1NI2_2(.din(w_dff_B_nth6Zzm01_2),.dout(w_dff_B_ZBCUt1NI2_2),.clk(gclk));
	jdff dff_B_8FaVY4zQ0_2(.din(w_dff_B_ZBCUt1NI2_2),.dout(w_dff_B_8FaVY4zQ0_2),.clk(gclk));
	jdff dff_B_KFce92R43_2(.din(w_dff_B_8FaVY4zQ0_2),.dout(w_dff_B_KFce92R43_2),.clk(gclk));
	jdff dff_B_qgVSkdWw7_2(.din(w_dff_B_KFce92R43_2),.dout(w_dff_B_qgVSkdWw7_2),.clk(gclk));
	jdff dff_B_MfUfDEm14_2(.din(w_dff_B_qgVSkdWw7_2),.dout(w_dff_B_MfUfDEm14_2),.clk(gclk));
	jdff dff_B_SWgQFbfC1_2(.din(w_dff_B_MfUfDEm14_2),.dout(w_dff_B_SWgQFbfC1_2),.clk(gclk));
	jdff dff_B_WY7lLxqQ4_2(.din(w_dff_B_SWgQFbfC1_2),.dout(w_dff_B_WY7lLxqQ4_2),.clk(gclk));
	jdff dff_B_OoDwh6u38_2(.din(w_dff_B_WY7lLxqQ4_2),.dout(w_dff_B_OoDwh6u38_2),.clk(gclk));
	jdff dff_B_XyZwpfnq1_2(.din(w_dff_B_OoDwh6u38_2),.dout(w_dff_B_XyZwpfnq1_2),.clk(gclk));
	jdff dff_B_GULrO4eb3_2(.din(w_dff_B_XyZwpfnq1_2),.dout(w_dff_B_GULrO4eb3_2),.clk(gclk));
	jdff dff_B_6rEcWJbo5_2(.din(w_dff_B_GULrO4eb3_2),.dout(w_dff_B_6rEcWJbo5_2),.clk(gclk));
	jdff dff_B_dh9tn2rf4_2(.din(w_dff_B_6rEcWJbo5_2),.dout(w_dff_B_dh9tn2rf4_2),.clk(gclk));
	jdff dff_B_WXktlnfk4_2(.din(w_dff_B_dh9tn2rf4_2),.dout(w_dff_B_WXktlnfk4_2),.clk(gclk));
	jdff dff_B_BScdIvYp7_2(.din(w_dff_B_WXktlnfk4_2),.dout(w_dff_B_BScdIvYp7_2),.clk(gclk));
	jdff dff_B_fCJsykjG5_2(.din(w_dff_B_BScdIvYp7_2),.dout(w_dff_B_fCJsykjG5_2),.clk(gclk));
	jdff dff_B_13rVuZoF7_2(.din(w_dff_B_fCJsykjG5_2),.dout(w_dff_B_13rVuZoF7_2),.clk(gclk));
	jdff dff_B_8q6t7x9G8_2(.din(w_dff_B_13rVuZoF7_2),.dout(w_dff_B_8q6t7x9G8_2),.clk(gclk));
	jdff dff_B_UVZGFrqb4_2(.din(w_dff_B_8q6t7x9G8_2),.dout(w_dff_B_UVZGFrqb4_2),.clk(gclk));
	jdff dff_B_Thh2GDD83_2(.din(w_dff_B_UVZGFrqb4_2),.dout(w_dff_B_Thh2GDD83_2),.clk(gclk));
	jdff dff_B_qSWBQnpy2_2(.din(w_dff_B_Thh2GDD83_2),.dout(w_dff_B_qSWBQnpy2_2),.clk(gclk));
	jdff dff_B_jYR6UxKH7_2(.din(w_dff_B_qSWBQnpy2_2),.dout(w_dff_B_jYR6UxKH7_2),.clk(gclk));
	jdff dff_B_DbNIh9ig4_2(.din(w_dff_B_jYR6UxKH7_2),.dout(w_dff_B_DbNIh9ig4_2),.clk(gclk));
	jdff dff_B_GsJrEfF28_2(.din(w_dff_B_DbNIh9ig4_2),.dout(w_dff_B_GsJrEfF28_2),.clk(gclk));
	jdff dff_B_lDy8tTWb4_2(.din(w_dff_B_GsJrEfF28_2),.dout(w_dff_B_lDy8tTWb4_2),.clk(gclk));
	jdff dff_B_84DxAPml2_2(.din(w_dff_B_lDy8tTWb4_2),.dout(w_dff_B_84DxAPml2_2),.clk(gclk));
	jdff dff_B_qwVJrxPE7_2(.din(w_dff_B_84DxAPml2_2),.dout(w_dff_B_qwVJrxPE7_2),.clk(gclk));
	jdff dff_B_7y3vtOru1_2(.din(w_dff_B_qwVJrxPE7_2),.dout(w_dff_B_7y3vtOru1_2),.clk(gclk));
	jdff dff_B_jz9gIu8r3_2(.din(w_dff_B_7y3vtOru1_2),.dout(w_dff_B_jz9gIu8r3_2),.clk(gclk));
	jdff dff_B_0MtxO2Sz1_2(.din(w_dff_B_jz9gIu8r3_2),.dout(w_dff_B_0MtxO2Sz1_2),.clk(gclk));
	jdff dff_B_XyLSfHrD3_2(.din(w_dff_B_0MtxO2Sz1_2),.dout(w_dff_B_XyLSfHrD3_2),.clk(gclk));
	jdff dff_B_57i03B9h9_2(.din(w_dff_B_XyLSfHrD3_2),.dout(w_dff_B_57i03B9h9_2),.clk(gclk));
	jdff dff_B_adTaDt612_2(.din(w_dff_B_57i03B9h9_2),.dout(w_dff_B_adTaDt612_2),.clk(gclk));
	jdff dff_B_DaLsLcXI6_2(.din(w_dff_B_adTaDt612_2),.dout(w_dff_B_DaLsLcXI6_2),.clk(gclk));
	jdff dff_B_3kIobVxA7_2(.din(w_dff_B_DaLsLcXI6_2),.dout(w_dff_B_3kIobVxA7_2),.clk(gclk));
	jdff dff_B_oBF2lXrS3_2(.din(w_dff_B_3kIobVxA7_2),.dout(w_dff_B_oBF2lXrS3_2),.clk(gclk));
	jdff dff_B_sBWxF3Ru3_2(.din(w_dff_B_oBF2lXrS3_2),.dout(w_dff_B_sBWxF3Ru3_2),.clk(gclk));
	jdff dff_B_5jJWr6HJ8_2(.din(w_dff_B_sBWxF3Ru3_2),.dout(w_dff_B_5jJWr6HJ8_2),.clk(gclk));
	jdff dff_B_BKRyAMPI2_2(.din(w_dff_B_5jJWr6HJ8_2),.dout(w_dff_B_BKRyAMPI2_2),.clk(gclk));
	jdff dff_B_z22qLd3X2_2(.din(w_dff_B_BKRyAMPI2_2),.dout(w_dff_B_z22qLd3X2_2),.clk(gclk));
	jdff dff_B_Z6YhwrNl1_2(.din(w_dff_B_z22qLd3X2_2),.dout(w_dff_B_Z6YhwrNl1_2),.clk(gclk));
	jdff dff_B_BVZmH9Fj5_2(.din(n1776),.dout(w_dff_B_BVZmH9Fj5_2),.clk(gclk));
	jdff dff_B_7JXgpsbT1_2(.din(w_dff_B_BVZmH9Fj5_2),.dout(w_dff_B_7JXgpsbT1_2),.clk(gclk));
	jdff dff_B_zL97k3z71_2(.din(w_dff_B_7JXgpsbT1_2),.dout(w_dff_B_zL97k3z71_2),.clk(gclk));
	jdff dff_B_pqGf6b2E9_2(.din(w_dff_B_zL97k3z71_2),.dout(w_dff_B_pqGf6b2E9_2),.clk(gclk));
	jdff dff_B_q7YYC9048_2(.din(w_dff_B_pqGf6b2E9_2),.dout(w_dff_B_q7YYC9048_2),.clk(gclk));
	jdff dff_B_fs7uiKUb7_2(.din(w_dff_B_q7YYC9048_2),.dout(w_dff_B_fs7uiKUb7_2),.clk(gclk));
	jdff dff_B_lfjrS0234_2(.din(w_dff_B_fs7uiKUb7_2),.dout(w_dff_B_lfjrS0234_2),.clk(gclk));
	jdff dff_B_WsdavIZf1_2(.din(w_dff_B_lfjrS0234_2),.dout(w_dff_B_WsdavIZf1_2),.clk(gclk));
	jdff dff_B_C6gMaQTZ2_2(.din(w_dff_B_WsdavIZf1_2),.dout(w_dff_B_C6gMaQTZ2_2),.clk(gclk));
	jdff dff_B_qwozOQVE0_2(.din(w_dff_B_C6gMaQTZ2_2),.dout(w_dff_B_qwozOQVE0_2),.clk(gclk));
	jdff dff_B_nhX3f3B65_2(.din(w_dff_B_qwozOQVE0_2),.dout(w_dff_B_nhX3f3B65_2),.clk(gclk));
	jdff dff_B_hKYoVlqY9_2(.din(w_dff_B_nhX3f3B65_2),.dout(w_dff_B_hKYoVlqY9_2),.clk(gclk));
	jdff dff_B_12yvBWWU6_2(.din(w_dff_B_hKYoVlqY9_2),.dout(w_dff_B_12yvBWWU6_2),.clk(gclk));
	jdff dff_B_XiavbY4o8_2(.din(w_dff_B_12yvBWWU6_2),.dout(w_dff_B_XiavbY4o8_2),.clk(gclk));
	jdff dff_B_Tc3xqEJy7_2(.din(w_dff_B_XiavbY4o8_2),.dout(w_dff_B_Tc3xqEJy7_2),.clk(gclk));
	jdff dff_B_93kJDd5I0_2(.din(w_dff_B_Tc3xqEJy7_2),.dout(w_dff_B_93kJDd5I0_2),.clk(gclk));
	jdff dff_B_UrLgxFgP5_2(.din(w_dff_B_93kJDd5I0_2),.dout(w_dff_B_UrLgxFgP5_2),.clk(gclk));
	jdff dff_B_Q8DmjmFR8_2(.din(w_dff_B_UrLgxFgP5_2),.dout(w_dff_B_Q8DmjmFR8_2),.clk(gclk));
	jdff dff_B_aSdGkBWq0_2(.din(w_dff_B_Q8DmjmFR8_2),.dout(w_dff_B_aSdGkBWq0_2),.clk(gclk));
	jdff dff_B_6VEaBnXq3_2(.din(w_dff_B_aSdGkBWq0_2),.dout(w_dff_B_6VEaBnXq3_2),.clk(gclk));
	jdff dff_B_23Xr9Jzk4_2(.din(w_dff_B_6VEaBnXq3_2),.dout(w_dff_B_23Xr9Jzk4_2),.clk(gclk));
	jdff dff_B_onEYiaQZ5_2(.din(w_dff_B_23Xr9Jzk4_2),.dout(w_dff_B_onEYiaQZ5_2),.clk(gclk));
	jdff dff_B_k0aWeSkx5_2(.din(w_dff_B_onEYiaQZ5_2),.dout(w_dff_B_k0aWeSkx5_2),.clk(gclk));
	jdff dff_B_Qjb1zy3w3_2(.din(w_dff_B_k0aWeSkx5_2),.dout(w_dff_B_Qjb1zy3w3_2),.clk(gclk));
	jdff dff_B_cZke7L2V5_2(.din(w_dff_B_Qjb1zy3w3_2),.dout(w_dff_B_cZke7L2V5_2),.clk(gclk));
	jdff dff_B_bOhgOz0n7_2(.din(w_dff_B_cZke7L2V5_2),.dout(w_dff_B_bOhgOz0n7_2),.clk(gclk));
	jdff dff_B_lKP4KhVR3_2(.din(w_dff_B_bOhgOz0n7_2),.dout(w_dff_B_lKP4KhVR3_2),.clk(gclk));
	jdff dff_B_4cmNqf2c6_2(.din(w_dff_B_lKP4KhVR3_2),.dout(w_dff_B_4cmNqf2c6_2),.clk(gclk));
	jdff dff_B_hRg4920O2_2(.din(w_dff_B_4cmNqf2c6_2),.dout(w_dff_B_hRg4920O2_2),.clk(gclk));
	jdff dff_B_0nGkvphh9_2(.din(w_dff_B_hRg4920O2_2),.dout(w_dff_B_0nGkvphh9_2),.clk(gclk));
	jdff dff_B_c0oPyYeU3_2(.din(w_dff_B_0nGkvphh9_2),.dout(w_dff_B_c0oPyYeU3_2),.clk(gclk));
	jdff dff_B_5nOaUjMi0_2(.din(w_dff_B_c0oPyYeU3_2),.dout(w_dff_B_5nOaUjMi0_2),.clk(gclk));
	jdff dff_B_zstZZFWV7_2(.din(w_dff_B_5nOaUjMi0_2),.dout(w_dff_B_zstZZFWV7_2),.clk(gclk));
	jdff dff_B_bruJMJFn8_2(.din(w_dff_B_zstZZFWV7_2),.dout(w_dff_B_bruJMJFn8_2),.clk(gclk));
	jdff dff_B_qM5vG8ip3_2(.din(w_dff_B_bruJMJFn8_2),.dout(w_dff_B_qM5vG8ip3_2),.clk(gclk));
	jdff dff_B_Z2E20n928_2(.din(w_dff_B_qM5vG8ip3_2),.dout(w_dff_B_Z2E20n928_2),.clk(gclk));
	jdff dff_B_vdWqJbFJ6_2(.din(w_dff_B_Z2E20n928_2),.dout(w_dff_B_vdWqJbFJ6_2),.clk(gclk));
	jdff dff_B_CmabRUo87_2(.din(w_dff_B_vdWqJbFJ6_2),.dout(w_dff_B_CmabRUo87_2),.clk(gclk));
	jdff dff_B_KsfOcV4e3_2(.din(w_dff_B_CmabRUo87_2),.dout(w_dff_B_KsfOcV4e3_2),.clk(gclk));
	jdff dff_B_n5E5HmvU4_2(.din(w_dff_B_KsfOcV4e3_2),.dout(w_dff_B_n5E5HmvU4_2),.clk(gclk));
	jdff dff_B_GzRa2q4H0_2(.din(w_dff_B_n5E5HmvU4_2),.dout(w_dff_B_GzRa2q4H0_2),.clk(gclk));
	jdff dff_B_staIUWfV4_2(.din(w_dff_B_GzRa2q4H0_2),.dout(w_dff_B_staIUWfV4_2),.clk(gclk));
	jdff dff_B_CG8DoOEK9_2(.din(w_dff_B_staIUWfV4_2),.dout(w_dff_B_CG8DoOEK9_2),.clk(gclk));
	jdff dff_B_o3yT1ZIc1_2(.din(w_dff_B_CG8DoOEK9_2),.dout(w_dff_B_o3yT1ZIc1_2),.clk(gclk));
	jdff dff_B_qHfqmhz79_2(.din(w_dff_B_o3yT1ZIc1_2),.dout(w_dff_B_qHfqmhz79_2),.clk(gclk));
	jdff dff_B_4g1I6MsN8_2(.din(w_dff_B_qHfqmhz79_2),.dout(w_dff_B_4g1I6MsN8_2),.clk(gclk));
	jdff dff_B_dmRd39eB5_2(.din(w_dff_B_4g1I6MsN8_2),.dout(w_dff_B_dmRd39eB5_2),.clk(gclk));
	jdff dff_B_gsq2MKZ29_2(.din(w_dff_B_dmRd39eB5_2),.dout(w_dff_B_gsq2MKZ29_2),.clk(gclk));
	jdff dff_B_8057qEsG4_2(.din(w_dff_B_gsq2MKZ29_2),.dout(w_dff_B_8057qEsG4_2),.clk(gclk));
	jdff dff_B_QULvV8V88_2(.din(w_dff_B_8057qEsG4_2),.dout(w_dff_B_QULvV8V88_2),.clk(gclk));
	jdff dff_B_BMwC0cpx0_2(.din(w_dff_B_QULvV8V88_2),.dout(w_dff_B_BMwC0cpx0_2),.clk(gclk));
	jdff dff_B_xwJvQPur6_2(.din(n1775),.dout(w_dff_B_xwJvQPur6_2),.clk(gclk));
	jdff dff_B_7dpaZHxq8_1(.din(n1773),.dout(w_dff_B_7dpaZHxq8_1),.clk(gclk));
	jdff dff_B_av0Z4jtR1_2(.din(n1744),.dout(w_dff_B_av0Z4jtR1_2),.clk(gclk));
	jdff dff_B_6qEj3pS98_2(.din(w_dff_B_av0Z4jtR1_2),.dout(w_dff_B_6qEj3pS98_2),.clk(gclk));
	jdff dff_B_i9tYDqdD2_2(.din(w_dff_B_6qEj3pS98_2),.dout(w_dff_B_i9tYDqdD2_2),.clk(gclk));
	jdff dff_B_4syNUP6B8_2(.din(w_dff_B_i9tYDqdD2_2),.dout(w_dff_B_4syNUP6B8_2),.clk(gclk));
	jdff dff_B_TyzTntKf3_2(.din(w_dff_B_4syNUP6B8_2),.dout(w_dff_B_TyzTntKf3_2),.clk(gclk));
	jdff dff_B_yy1RzfvQ4_2(.din(w_dff_B_TyzTntKf3_2),.dout(w_dff_B_yy1RzfvQ4_2),.clk(gclk));
	jdff dff_B_gCtZIFNU9_2(.din(w_dff_B_yy1RzfvQ4_2),.dout(w_dff_B_gCtZIFNU9_2),.clk(gclk));
	jdff dff_B_RGmZhSRa0_2(.din(w_dff_B_gCtZIFNU9_2),.dout(w_dff_B_RGmZhSRa0_2),.clk(gclk));
	jdff dff_B_Y2dCptr67_2(.din(w_dff_B_RGmZhSRa0_2),.dout(w_dff_B_Y2dCptr67_2),.clk(gclk));
	jdff dff_B_pnUedo9w9_2(.din(w_dff_B_Y2dCptr67_2),.dout(w_dff_B_pnUedo9w9_2),.clk(gclk));
	jdff dff_B_nxtiiZGi9_2(.din(w_dff_B_pnUedo9w9_2),.dout(w_dff_B_nxtiiZGi9_2),.clk(gclk));
	jdff dff_B_WsO6rbGz8_2(.din(w_dff_B_nxtiiZGi9_2),.dout(w_dff_B_WsO6rbGz8_2),.clk(gclk));
	jdff dff_B_t2pv4I0G9_2(.din(w_dff_B_WsO6rbGz8_2),.dout(w_dff_B_t2pv4I0G9_2),.clk(gclk));
	jdff dff_B_dM1QLNk81_2(.din(w_dff_B_t2pv4I0G9_2),.dout(w_dff_B_dM1QLNk81_2),.clk(gclk));
	jdff dff_B_cPgayzv85_2(.din(w_dff_B_dM1QLNk81_2),.dout(w_dff_B_cPgayzv85_2),.clk(gclk));
	jdff dff_B_eZhtcYPL1_2(.din(w_dff_B_cPgayzv85_2),.dout(w_dff_B_eZhtcYPL1_2),.clk(gclk));
	jdff dff_B_UVmh4zAv5_2(.din(w_dff_B_eZhtcYPL1_2),.dout(w_dff_B_UVmh4zAv5_2),.clk(gclk));
	jdff dff_B_KSttIiVW9_2(.din(w_dff_B_UVmh4zAv5_2),.dout(w_dff_B_KSttIiVW9_2),.clk(gclk));
	jdff dff_B_NuZYHMkO0_2(.din(w_dff_B_KSttIiVW9_2),.dout(w_dff_B_NuZYHMkO0_2),.clk(gclk));
	jdff dff_B_su2KVq545_2(.din(w_dff_B_NuZYHMkO0_2),.dout(w_dff_B_su2KVq545_2),.clk(gclk));
	jdff dff_B_2P1inuRz5_2(.din(w_dff_B_su2KVq545_2),.dout(w_dff_B_2P1inuRz5_2),.clk(gclk));
	jdff dff_B_yY6onhTI9_2(.din(w_dff_B_2P1inuRz5_2),.dout(w_dff_B_yY6onhTI9_2),.clk(gclk));
	jdff dff_B_xoGKECVJ9_2(.din(w_dff_B_yY6onhTI9_2),.dout(w_dff_B_xoGKECVJ9_2),.clk(gclk));
	jdff dff_B_UVaiboU92_2(.din(w_dff_B_xoGKECVJ9_2),.dout(w_dff_B_UVaiboU92_2),.clk(gclk));
	jdff dff_B_ICW8Ev2L5_2(.din(w_dff_B_UVaiboU92_2),.dout(w_dff_B_ICW8Ev2L5_2),.clk(gclk));
	jdff dff_B_Nf6GLSV29_2(.din(w_dff_B_ICW8Ev2L5_2),.dout(w_dff_B_Nf6GLSV29_2),.clk(gclk));
	jdff dff_B_VrN9zv2U0_2(.din(w_dff_B_Nf6GLSV29_2),.dout(w_dff_B_VrN9zv2U0_2),.clk(gclk));
	jdff dff_B_ddmjZsiA7_2(.din(w_dff_B_VrN9zv2U0_2),.dout(w_dff_B_ddmjZsiA7_2),.clk(gclk));
	jdff dff_B_I6WMBrAw8_2(.din(w_dff_B_ddmjZsiA7_2),.dout(w_dff_B_I6WMBrAw8_2),.clk(gclk));
	jdff dff_B_VSHuEfxU0_2(.din(w_dff_B_I6WMBrAw8_2),.dout(w_dff_B_VSHuEfxU0_2),.clk(gclk));
	jdff dff_B_uDkSno7C4_2(.din(w_dff_B_VSHuEfxU0_2),.dout(w_dff_B_uDkSno7C4_2),.clk(gclk));
	jdff dff_B_PnF0CkH76_2(.din(w_dff_B_uDkSno7C4_2),.dout(w_dff_B_PnF0CkH76_2),.clk(gclk));
	jdff dff_B_hnNILBVt1_2(.din(w_dff_B_PnF0CkH76_2),.dout(w_dff_B_hnNILBVt1_2),.clk(gclk));
	jdff dff_B_t62sOwyR2_2(.din(w_dff_B_hnNILBVt1_2),.dout(w_dff_B_t62sOwyR2_2),.clk(gclk));
	jdff dff_B_dlcYo8dZ8_2(.din(w_dff_B_t62sOwyR2_2),.dout(w_dff_B_dlcYo8dZ8_2),.clk(gclk));
	jdff dff_B_5ZtZWLSG3_2(.din(w_dff_B_dlcYo8dZ8_2),.dout(w_dff_B_5ZtZWLSG3_2),.clk(gclk));
	jdff dff_B_iSX1nsKp7_2(.din(w_dff_B_5ZtZWLSG3_2),.dout(w_dff_B_iSX1nsKp7_2),.clk(gclk));
	jdff dff_B_Dkg3i56c5_2(.din(w_dff_B_iSX1nsKp7_2),.dout(w_dff_B_Dkg3i56c5_2),.clk(gclk));
	jdff dff_B_uhQ1kuob9_2(.din(w_dff_B_Dkg3i56c5_2),.dout(w_dff_B_uhQ1kuob9_2),.clk(gclk));
	jdff dff_B_1ivoFxOM5_2(.din(w_dff_B_uhQ1kuob9_2),.dout(w_dff_B_1ivoFxOM5_2),.clk(gclk));
	jdff dff_B_v0im1tBe6_2(.din(w_dff_B_1ivoFxOM5_2),.dout(w_dff_B_v0im1tBe6_2),.clk(gclk));
	jdff dff_B_9IkQZ6dB1_2(.din(w_dff_B_v0im1tBe6_2),.dout(w_dff_B_9IkQZ6dB1_2),.clk(gclk));
	jdff dff_B_daRRA12K6_2(.din(w_dff_B_9IkQZ6dB1_2),.dout(w_dff_B_daRRA12K6_2),.clk(gclk));
	jdff dff_B_DDDeFEzQ2_2(.din(w_dff_B_daRRA12K6_2),.dout(w_dff_B_DDDeFEzQ2_2),.clk(gclk));
	jdff dff_B_WXeeu8oa4_2(.din(w_dff_B_DDDeFEzQ2_2),.dout(w_dff_B_WXeeu8oa4_2),.clk(gclk));
	jdff dff_B_9Wo1o3nk9_2(.din(w_dff_B_WXeeu8oa4_2),.dout(w_dff_B_9Wo1o3nk9_2),.clk(gclk));
	jdff dff_B_piTGDidU7_2(.din(w_dff_B_9Wo1o3nk9_2),.dout(w_dff_B_piTGDidU7_2),.clk(gclk));
	jdff dff_B_J8pEQWx43_2(.din(w_dff_B_piTGDidU7_2),.dout(w_dff_B_J8pEQWx43_2),.clk(gclk));
	jdff dff_B_xOGJrbx65_1(.din(n1750),.dout(w_dff_B_xOGJrbx65_1),.clk(gclk));
	jdff dff_B_Eb1e4zv05_1(.din(w_dff_B_xOGJrbx65_1),.dout(w_dff_B_Eb1e4zv05_1),.clk(gclk));
	jdff dff_B_QTUrXhTB7_2(.din(n1749),.dout(w_dff_B_QTUrXhTB7_2),.clk(gclk));
	jdff dff_B_bDexCrgx5_2(.din(w_dff_B_QTUrXhTB7_2),.dout(w_dff_B_bDexCrgx5_2),.clk(gclk));
	jdff dff_B_Avs9lNBp1_2(.din(w_dff_B_bDexCrgx5_2),.dout(w_dff_B_Avs9lNBp1_2),.clk(gclk));
	jdff dff_B_2SVGwvrh9_2(.din(w_dff_B_Avs9lNBp1_2),.dout(w_dff_B_2SVGwvrh9_2),.clk(gclk));
	jdff dff_B_tlsCTcUM0_2(.din(w_dff_B_2SVGwvrh9_2),.dout(w_dff_B_tlsCTcUM0_2),.clk(gclk));
	jdff dff_B_N0zI1NNW1_2(.din(w_dff_B_tlsCTcUM0_2),.dout(w_dff_B_N0zI1NNW1_2),.clk(gclk));
	jdff dff_B_E3L3xIaM1_2(.din(w_dff_B_N0zI1NNW1_2),.dout(w_dff_B_E3L3xIaM1_2),.clk(gclk));
	jdff dff_B_DTvsiQKD0_2(.din(w_dff_B_E3L3xIaM1_2),.dout(w_dff_B_DTvsiQKD0_2),.clk(gclk));
	jdff dff_B_QaZTbXsw8_2(.din(w_dff_B_DTvsiQKD0_2),.dout(w_dff_B_QaZTbXsw8_2),.clk(gclk));
	jdff dff_B_QzNICzxk3_2(.din(w_dff_B_QaZTbXsw8_2),.dout(w_dff_B_QzNICzxk3_2),.clk(gclk));
	jdff dff_B_mjeW80UN4_2(.din(w_dff_B_QzNICzxk3_2),.dout(w_dff_B_mjeW80UN4_2),.clk(gclk));
	jdff dff_B_7kYzLfl41_2(.din(w_dff_B_mjeW80UN4_2),.dout(w_dff_B_7kYzLfl41_2),.clk(gclk));
	jdff dff_B_dQqgCHMh2_2(.din(w_dff_B_7kYzLfl41_2),.dout(w_dff_B_dQqgCHMh2_2),.clk(gclk));
	jdff dff_B_RMPISNWG4_2(.din(w_dff_B_dQqgCHMh2_2),.dout(w_dff_B_RMPISNWG4_2),.clk(gclk));
	jdff dff_B_8T9FbkBe1_2(.din(w_dff_B_RMPISNWG4_2),.dout(w_dff_B_8T9FbkBe1_2),.clk(gclk));
	jdff dff_B_x1xgvqI17_2(.din(w_dff_B_8T9FbkBe1_2),.dout(w_dff_B_x1xgvqI17_2),.clk(gclk));
	jdff dff_B_3aj5npzq6_2(.din(w_dff_B_x1xgvqI17_2),.dout(w_dff_B_3aj5npzq6_2),.clk(gclk));
	jdff dff_B_ZKXZdRes4_2(.din(w_dff_B_3aj5npzq6_2),.dout(w_dff_B_ZKXZdRes4_2),.clk(gclk));
	jdff dff_B_OOne1VRC8_2(.din(w_dff_B_ZKXZdRes4_2),.dout(w_dff_B_OOne1VRC8_2),.clk(gclk));
	jdff dff_B_cq6H0Ksa1_2(.din(w_dff_B_OOne1VRC8_2),.dout(w_dff_B_cq6H0Ksa1_2),.clk(gclk));
	jdff dff_B_TbOS0GcV4_2(.din(w_dff_B_cq6H0Ksa1_2),.dout(w_dff_B_TbOS0GcV4_2),.clk(gclk));
	jdff dff_B_TE7dmQcq4_2(.din(w_dff_B_TbOS0GcV4_2),.dout(w_dff_B_TE7dmQcq4_2),.clk(gclk));
	jdff dff_B_zPEcD1dR1_2(.din(w_dff_B_TE7dmQcq4_2),.dout(w_dff_B_zPEcD1dR1_2),.clk(gclk));
	jdff dff_B_OTgWJMc69_2(.din(w_dff_B_zPEcD1dR1_2),.dout(w_dff_B_OTgWJMc69_2),.clk(gclk));
	jdff dff_B_S0dumocq8_2(.din(w_dff_B_OTgWJMc69_2),.dout(w_dff_B_S0dumocq8_2),.clk(gclk));
	jdff dff_B_jgvt7n2v2_2(.din(w_dff_B_S0dumocq8_2),.dout(w_dff_B_jgvt7n2v2_2),.clk(gclk));
	jdff dff_B_nRTinHS83_2(.din(w_dff_B_jgvt7n2v2_2),.dout(w_dff_B_nRTinHS83_2),.clk(gclk));
	jdff dff_B_AAvTchCT3_2(.din(w_dff_B_nRTinHS83_2),.dout(w_dff_B_AAvTchCT3_2),.clk(gclk));
	jdff dff_B_Y6jvpiLY7_2(.din(w_dff_B_AAvTchCT3_2),.dout(w_dff_B_Y6jvpiLY7_2),.clk(gclk));
	jdff dff_B_PYTlLPgU2_2(.din(w_dff_B_Y6jvpiLY7_2),.dout(w_dff_B_PYTlLPgU2_2),.clk(gclk));
	jdff dff_B_g4p8XUGx3_2(.din(w_dff_B_PYTlLPgU2_2),.dout(w_dff_B_g4p8XUGx3_2),.clk(gclk));
	jdff dff_B_4Vgkvirh1_2(.din(w_dff_B_g4p8XUGx3_2),.dout(w_dff_B_4Vgkvirh1_2),.clk(gclk));
	jdff dff_B_sGD4DW2H3_2(.din(w_dff_B_4Vgkvirh1_2),.dout(w_dff_B_sGD4DW2H3_2),.clk(gclk));
	jdff dff_B_sozmydQQ7_2(.din(w_dff_B_sGD4DW2H3_2),.dout(w_dff_B_sozmydQQ7_2),.clk(gclk));
	jdff dff_B_J3qRzl3k4_2(.din(w_dff_B_sozmydQQ7_2),.dout(w_dff_B_J3qRzl3k4_2),.clk(gclk));
	jdff dff_B_aIvhg7WE1_2(.din(w_dff_B_J3qRzl3k4_2),.dout(w_dff_B_aIvhg7WE1_2),.clk(gclk));
	jdff dff_B_VOQUcd8l4_2(.din(w_dff_B_aIvhg7WE1_2),.dout(w_dff_B_VOQUcd8l4_2),.clk(gclk));
	jdff dff_B_LTv6hB2J8_2(.din(w_dff_B_VOQUcd8l4_2),.dout(w_dff_B_LTv6hB2J8_2),.clk(gclk));
	jdff dff_B_0FfXaU3J1_2(.din(w_dff_B_LTv6hB2J8_2),.dout(w_dff_B_0FfXaU3J1_2),.clk(gclk));
	jdff dff_B_hfjAzmzM9_2(.din(w_dff_B_0FfXaU3J1_2),.dout(w_dff_B_hfjAzmzM9_2),.clk(gclk));
	jdff dff_B_rM7khkJN1_2(.din(w_dff_B_hfjAzmzM9_2),.dout(w_dff_B_rM7khkJN1_2),.clk(gclk));
	jdff dff_B_OrhBpZSr5_2(.din(w_dff_B_rM7khkJN1_2),.dout(w_dff_B_OrhBpZSr5_2),.clk(gclk));
	jdff dff_B_RTdvRxML0_2(.din(w_dff_B_OrhBpZSr5_2),.dout(w_dff_B_RTdvRxML0_2),.clk(gclk));
	jdff dff_B_LtRtLIKV1_2(.din(w_dff_B_RTdvRxML0_2),.dout(w_dff_B_LtRtLIKV1_2),.clk(gclk));
	jdff dff_B_GdviRPqa7_2(.din(w_dff_B_LtRtLIKV1_2),.dout(w_dff_B_GdviRPqa7_2),.clk(gclk));
	jdff dff_B_s0ChG4Md8_2(.din(n1748),.dout(w_dff_B_s0ChG4Md8_2),.clk(gclk));
	jdff dff_B_zp14U6pT5_2(.din(w_dff_B_s0ChG4Md8_2),.dout(w_dff_B_zp14U6pT5_2),.clk(gclk));
	jdff dff_B_USgDcLoi1_2(.din(w_dff_B_zp14U6pT5_2),.dout(w_dff_B_USgDcLoi1_2),.clk(gclk));
	jdff dff_B_A1zY5Kij0_2(.din(w_dff_B_USgDcLoi1_2),.dout(w_dff_B_A1zY5Kij0_2),.clk(gclk));
	jdff dff_B_rFOK6I2c3_2(.din(w_dff_B_A1zY5Kij0_2),.dout(w_dff_B_rFOK6I2c3_2),.clk(gclk));
	jdff dff_B_wHKvree92_2(.din(w_dff_B_rFOK6I2c3_2),.dout(w_dff_B_wHKvree92_2),.clk(gclk));
	jdff dff_B_ypwBiEOp5_2(.din(w_dff_B_wHKvree92_2),.dout(w_dff_B_ypwBiEOp5_2),.clk(gclk));
	jdff dff_B_aVDZ4jek4_2(.din(w_dff_B_ypwBiEOp5_2),.dout(w_dff_B_aVDZ4jek4_2),.clk(gclk));
	jdff dff_B_gGL9Nctf8_2(.din(w_dff_B_aVDZ4jek4_2),.dout(w_dff_B_gGL9Nctf8_2),.clk(gclk));
	jdff dff_B_2dwFD92M6_2(.din(w_dff_B_gGL9Nctf8_2),.dout(w_dff_B_2dwFD92M6_2),.clk(gclk));
	jdff dff_B_dTB2xocl2_2(.din(w_dff_B_2dwFD92M6_2),.dout(w_dff_B_dTB2xocl2_2),.clk(gclk));
	jdff dff_B_WTI3i5HF6_2(.din(w_dff_B_dTB2xocl2_2),.dout(w_dff_B_WTI3i5HF6_2),.clk(gclk));
	jdff dff_B_BIaSBGVc9_2(.din(w_dff_B_WTI3i5HF6_2),.dout(w_dff_B_BIaSBGVc9_2),.clk(gclk));
	jdff dff_B_bCYW4vfu7_2(.din(w_dff_B_BIaSBGVc9_2),.dout(w_dff_B_bCYW4vfu7_2),.clk(gclk));
	jdff dff_B_doOVltAs6_2(.din(w_dff_B_bCYW4vfu7_2),.dout(w_dff_B_doOVltAs6_2),.clk(gclk));
	jdff dff_B_SNRvUApd2_2(.din(w_dff_B_doOVltAs6_2),.dout(w_dff_B_SNRvUApd2_2),.clk(gclk));
	jdff dff_B_il0aZ23A7_2(.din(w_dff_B_SNRvUApd2_2),.dout(w_dff_B_il0aZ23A7_2),.clk(gclk));
	jdff dff_B_oOKMVDjz3_2(.din(w_dff_B_il0aZ23A7_2),.dout(w_dff_B_oOKMVDjz3_2),.clk(gclk));
	jdff dff_B_6nf6vUhG4_2(.din(w_dff_B_oOKMVDjz3_2),.dout(w_dff_B_6nf6vUhG4_2),.clk(gclk));
	jdff dff_B_KU0hY5iM2_2(.din(w_dff_B_6nf6vUhG4_2),.dout(w_dff_B_KU0hY5iM2_2),.clk(gclk));
	jdff dff_B_ku4WOzi16_2(.din(w_dff_B_KU0hY5iM2_2),.dout(w_dff_B_ku4WOzi16_2),.clk(gclk));
	jdff dff_B_Q90A9N5n7_2(.din(w_dff_B_ku4WOzi16_2),.dout(w_dff_B_Q90A9N5n7_2),.clk(gclk));
	jdff dff_B_qTNOXtMI8_2(.din(w_dff_B_Q90A9N5n7_2),.dout(w_dff_B_qTNOXtMI8_2),.clk(gclk));
	jdff dff_B_Af15cCWq9_2(.din(w_dff_B_qTNOXtMI8_2),.dout(w_dff_B_Af15cCWq9_2),.clk(gclk));
	jdff dff_B_ZaVDupB09_2(.din(w_dff_B_Af15cCWq9_2),.dout(w_dff_B_ZaVDupB09_2),.clk(gclk));
	jdff dff_B_a79sutxU0_2(.din(w_dff_B_ZaVDupB09_2),.dout(w_dff_B_a79sutxU0_2),.clk(gclk));
	jdff dff_B_wPlm9PoA1_2(.din(w_dff_B_a79sutxU0_2),.dout(w_dff_B_wPlm9PoA1_2),.clk(gclk));
	jdff dff_B_3RIUMySV6_2(.din(w_dff_B_wPlm9PoA1_2),.dout(w_dff_B_3RIUMySV6_2),.clk(gclk));
	jdff dff_B_5VXRJeTX5_2(.din(w_dff_B_3RIUMySV6_2),.dout(w_dff_B_5VXRJeTX5_2),.clk(gclk));
	jdff dff_B_10E7R6jW3_2(.din(w_dff_B_5VXRJeTX5_2),.dout(w_dff_B_10E7R6jW3_2),.clk(gclk));
	jdff dff_B_4wxEo3nc5_2(.din(w_dff_B_10E7R6jW3_2),.dout(w_dff_B_4wxEo3nc5_2),.clk(gclk));
	jdff dff_B_kz4ZAxxS3_2(.din(w_dff_B_4wxEo3nc5_2),.dout(w_dff_B_kz4ZAxxS3_2),.clk(gclk));
	jdff dff_B_PJxYP14y4_2(.din(w_dff_B_kz4ZAxxS3_2),.dout(w_dff_B_PJxYP14y4_2),.clk(gclk));
	jdff dff_B_U8dQpLzK1_2(.din(w_dff_B_PJxYP14y4_2),.dout(w_dff_B_U8dQpLzK1_2),.clk(gclk));
	jdff dff_B_OMk2KzHJ8_2(.din(w_dff_B_U8dQpLzK1_2),.dout(w_dff_B_OMk2KzHJ8_2),.clk(gclk));
	jdff dff_B_eKIOurO45_2(.din(w_dff_B_OMk2KzHJ8_2),.dout(w_dff_B_eKIOurO45_2),.clk(gclk));
	jdff dff_B_zRAUS7gg5_2(.din(w_dff_B_eKIOurO45_2),.dout(w_dff_B_zRAUS7gg5_2),.clk(gclk));
	jdff dff_B_OqyqSyrB2_2(.din(w_dff_B_zRAUS7gg5_2),.dout(w_dff_B_OqyqSyrB2_2),.clk(gclk));
	jdff dff_B_l0R9GduR1_2(.din(w_dff_B_OqyqSyrB2_2),.dout(w_dff_B_l0R9GduR1_2),.clk(gclk));
	jdff dff_B_srBtELsK7_2(.din(w_dff_B_l0R9GduR1_2),.dout(w_dff_B_srBtELsK7_2),.clk(gclk));
	jdff dff_B_U0i14xFa9_2(.din(w_dff_B_srBtELsK7_2),.dout(w_dff_B_U0i14xFa9_2),.clk(gclk));
	jdff dff_B_wDQ379xY9_2(.din(w_dff_B_U0i14xFa9_2),.dout(w_dff_B_wDQ379xY9_2),.clk(gclk));
	jdff dff_B_fmd4f86b2_2(.din(w_dff_B_wDQ379xY9_2),.dout(w_dff_B_fmd4f86b2_2),.clk(gclk));
	jdff dff_B_ERW3I19F4_2(.din(w_dff_B_fmd4f86b2_2),.dout(w_dff_B_ERW3I19F4_2),.clk(gclk));
	jdff dff_B_DqXazg6O0_2(.din(w_dff_B_ERW3I19F4_2),.dout(w_dff_B_DqXazg6O0_2),.clk(gclk));
	jdff dff_B_xvv2OEut9_2(.din(w_dff_B_DqXazg6O0_2),.dout(w_dff_B_xvv2OEut9_2),.clk(gclk));
	jdff dff_B_sbxCKHqq8_2(.din(w_dff_B_xvv2OEut9_2),.dout(w_dff_B_sbxCKHqq8_2),.clk(gclk));
	jdff dff_B_pFri1iHH0_2(.din(n1747),.dout(w_dff_B_pFri1iHH0_2),.clk(gclk));
	jdff dff_B_8w4XTPpi9_1(.din(n1745),.dout(w_dff_B_8w4XTPpi9_1),.clk(gclk));
	jdff dff_B_4ZmHRJrV1_2(.din(n1709),.dout(w_dff_B_4ZmHRJrV1_2),.clk(gclk));
	jdff dff_B_9DNKNgt53_2(.din(w_dff_B_4ZmHRJrV1_2),.dout(w_dff_B_9DNKNgt53_2),.clk(gclk));
	jdff dff_B_FdlhnPA41_2(.din(w_dff_B_9DNKNgt53_2),.dout(w_dff_B_FdlhnPA41_2),.clk(gclk));
	jdff dff_B_vZU7n0tT8_2(.din(w_dff_B_FdlhnPA41_2),.dout(w_dff_B_vZU7n0tT8_2),.clk(gclk));
	jdff dff_B_3S5Vq60G4_2(.din(w_dff_B_vZU7n0tT8_2),.dout(w_dff_B_3S5Vq60G4_2),.clk(gclk));
	jdff dff_B_L96CCz5K7_2(.din(w_dff_B_3S5Vq60G4_2),.dout(w_dff_B_L96CCz5K7_2),.clk(gclk));
	jdff dff_B_SaIBBEzU0_2(.din(w_dff_B_L96CCz5K7_2),.dout(w_dff_B_SaIBBEzU0_2),.clk(gclk));
	jdff dff_B_Ayo4m5VA7_2(.din(w_dff_B_SaIBBEzU0_2),.dout(w_dff_B_Ayo4m5VA7_2),.clk(gclk));
	jdff dff_B_pcvehPN78_2(.din(w_dff_B_Ayo4m5VA7_2),.dout(w_dff_B_pcvehPN78_2),.clk(gclk));
	jdff dff_B_YOG5Umbu8_2(.din(w_dff_B_pcvehPN78_2),.dout(w_dff_B_YOG5Umbu8_2),.clk(gclk));
	jdff dff_B_pgx7HPXs2_2(.din(w_dff_B_YOG5Umbu8_2),.dout(w_dff_B_pgx7HPXs2_2),.clk(gclk));
	jdff dff_B_h9LwHkWn0_2(.din(w_dff_B_pgx7HPXs2_2),.dout(w_dff_B_h9LwHkWn0_2),.clk(gclk));
	jdff dff_B_5XRL5acR6_2(.din(w_dff_B_h9LwHkWn0_2),.dout(w_dff_B_5XRL5acR6_2),.clk(gclk));
	jdff dff_B_fkDkQe9K9_2(.din(w_dff_B_5XRL5acR6_2),.dout(w_dff_B_fkDkQe9K9_2),.clk(gclk));
	jdff dff_B_d0mRO7T62_2(.din(w_dff_B_fkDkQe9K9_2),.dout(w_dff_B_d0mRO7T62_2),.clk(gclk));
	jdff dff_B_LhW3JaGi3_2(.din(w_dff_B_d0mRO7T62_2),.dout(w_dff_B_LhW3JaGi3_2),.clk(gclk));
	jdff dff_B_A4c859rS3_2(.din(w_dff_B_LhW3JaGi3_2),.dout(w_dff_B_A4c859rS3_2),.clk(gclk));
	jdff dff_B_4HXw9Oxz5_2(.din(w_dff_B_A4c859rS3_2),.dout(w_dff_B_4HXw9Oxz5_2),.clk(gclk));
	jdff dff_B_BAH15Enk3_2(.din(w_dff_B_4HXw9Oxz5_2),.dout(w_dff_B_BAH15Enk3_2),.clk(gclk));
	jdff dff_B_AxzJNU8C1_2(.din(w_dff_B_BAH15Enk3_2),.dout(w_dff_B_AxzJNU8C1_2),.clk(gclk));
	jdff dff_B_y7VGyiwD9_2(.din(w_dff_B_AxzJNU8C1_2),.dout(w_dff_B_y7VGyiwD9_2),.clk(gclk));
	jdff dff_B_zS9rBlHi4_2(.din(w_dff_B_y7VGyiwD9_2),.dout(w_dff_B_zS9rBlHi4_2),.clk(gclk));
	jdff dff_B_z3DVdtej0_2(.din(w_dff_B_zS9rBlHi4_2),.dout(w_dff_B_z3DVdtej0_2),.clk(gclk));
	jdff dff_B_G6J0wWIt7_2(.din(w_dff_B_z3DVdtej0_2),.dout(w_dff_B_G6J0wWIt7_2),.clk(gclk));
	jdff dff_B_2oLprXB86_2(.din(w_dff_B_G6J0wWIt7_2),.dout(w_dff_B_2oLprXB86_2),.clk(gclk));
	jdff dff_B_WmSjZBjW8_2(.din(w_dff_B_2oLprXB86_2),.dout(w_dff_B_WmSjZBjW8_2),.clk(gclk));
	jdff dff_B_jTcoAEOm8_2(.din(w_dff_B_WmSjZBjW8_2),.dout(w_dff_B_jTcoAEOm8_2),.clk(gclk));
	jdff dff_B_ZzX2JLmr1_2(.din(w_dff_B_jTcoAEOm8_2),.dout(w_dff_B_ZzX2JLmr1_2),.clk(gclk));
	jdff dff_B_6VDsy6lD4_2(.din(w_dff_B_ZzX2JLmr1_2),.dout(w_dff_B_6VDsy6lD4_2),.clk(gclk));
	jdff dff_B_2moIeQY85_2(.din(w_dff_B_6VDsy6lD4_2),.dout(w_dff_B_2moIeQY85_2),.clk(gclk));
	jdff dff_B_Dsjxsjoh1_2(.din(w_dff_B_2moIeQY85_2),.dout(w_dff_B_Dsjxsjoh1_2),.clk(gclk));
	jdff dff_B_0z0GZMjg5_2(.din(w_dff_B_Dsjxsjoh1_2),.dout(w_dff_B_0z0GZMjg5_2),.clk(gclk));
	jdff dff_B_AWfUhAC55_2(.din(w_dff_B_0z0GZMjg5_2),.dout(w_dff_B_AWfUhAC55_2),.clk(gclk));
	jdff dff_B_EM9w7JRr1_2(.din(w_dff_B_AWfUhAC55_2),.dout(w_dff_B_EM9w7JRr1_2),.clk(gclk));
	jdff dff_B_ARSC4Ftf7_2(.din(w_dff_B_EM9w7JRr1_2),.dout(w_dff_B_ARSC4Ftf7_2),.clk(gclk));
	jdff dff_B_7WG6CZLr4_2(.din(w_dff_B_ARSC4Ftf7_2),.dout(w_dff_B_7WG6CZLr4_2),.clk(gclk));
	jdff dff_B_rBbTmy2f3_2(.din(w_dff_B_7WG6CZLr4_2),.dout(w_dff_B_rBbTmy2f3_2),.clk(gclk));
	jdff dff_B_1pfvS0JA0_2(.din(w_dff_B_rBbTmy2f3_2),.dout(w_dff_B_1pfvS0JA0_2),.clk(gclk));
	jdff dff_B_cBzBdBST9_2(.din(w_dff_B_1pfvS0JA0_2),.dout(w_dff_B_cBzBdBST9_2),.clk(gclk));
	jdff dff_B_q7Gqt4ro1_2(.din(w_dff_B_cBzBdBST9_2),.dout(w_dff_B_q7Gqt4ro1_2),.clk(gclk));
	jdff dff_B_M4eqRp689_2(.din(w_dff_B_q7Gqt4ro1_2),.dout(w_dff_B_M4eqRp689_2),.clk(gclk));
	jdff dff_B_e1L6mD2V7_2(.din(w_dff_B_M4eqRp689_2),.dout(w_dff_B_e1L6mD2V7_2),.clk(gclk));
	jdff dff_B_VmSCkBYu1_2(.din(w_dff_B_e1L6mD2V7_2),.dout(w_dff_B_VmSCkBYu1_2),.clk(gclk));
	jdff dff_B_RXpiju8U5_2(.din(w_dff_B_VmSCkBYu1_2),.dout(w_dff_B_RXpiju8U5_2),.clk(gclk));
	jdff dff_B_CqtpbViC8_1(.din(n1715),.dout(w_dff_B_CqtpbViC8_1),.clk(gclk));
	jdff dff_B_ongJG3EE9_1(.din(w_dff_B_CqtpbViC8_1),.dout(w_dff_B_ongJG3EE9_1),.clk(gclk));
	jdff dff_B_2CyJdK8Z7_2(.din(n1714),.dout(w_dff_B_2CyJdK8Z7_2),.clk(gclk));
	jdff dff_B_ncZPwi679_2(.din(w_dff_B_2CyJdK8Z7_2),.dout(w_dff_B_ncZPwi679_2),.clk(gclk));
	jdff dff_B_xop6ylVZ1_2(.din(w_dff_B_ncZPwi679_2),.dout(w_dff_B_xop6ylVZ1_2),.clk(gclk));
	jdff dff_B_DazW0yQB0_2(.din(w_dff_B_xop6ylVZ1_2),.dout(w_dff_B_DazW0yQB0_2),.clk(gclk));
	jdff dff_B_t9qFKXAZ4_2(.din(w_dff_B_DazW0yQB0_2),.dout(w_dff_B_t9qFKXAZ4_2),.clk(gclk));
	jdff dff_B_RnAt7tCc0_2(.din(w_dff_B_t9qFKXAZ4_2),.dout(w_dff_B_RnAt7tCc0_2),.clk(gclk));
	jdff dff_B_c4jEV9eq6_2(.din(w_dff_B_RnAt7tCc0_2),.dout(w_dff_B_c4jEV9eq6_2),.clk(gclk));
	jdff dff_B_8YgfvItd4_2(.din(w_dff_B_c4jEV9eq6_2),.dout(w_dff_B_8YgfvItd4_2),.clk(gclk));
	jdff dff_B_N7oLL6FB0_2(.din(w_dff_B_8YgfvItd4_2),.dout(w_dff_B_N7oLL6FB0_2),.clk(gclk));
	jdff dff_B_7U0dit3X6_2(.din(w_dff_B_N7oLL6FB0_2),.dout(w_dff_B_7U0dit3X6_2),.clk(gclk));
	jdff dff_B_49HGPpv23_2(.din(w_dff_B_7U0dit3X6_2),.dout(w_dff_B_49HGPpv23_2),.clk(gclk));
	jdff dff_B_nWfFf0ch5_2(.din(w_dff_B_49HGPpv23_2),.dout(w_dff_B_nWfFf0ch5_2),.clk(gclk));
	jdff dff_B_wK5urF5u2_2(.din(w_dff_B_nWfFf0ch5_2),.dout(w_dff_B_wK5urF5u2_2),.clk(gclk));
	jdff dff_B_HDQRt5lp3_2(.din(w_dff_B_wK5urF5u2_2),.dout(w_dff_B_HDQRt5lp3_2),.clk(gclk));
	jdff dff_B_b37Hy5GF2_2(.din(w_dff_B_HDQRt5lp3_2),.dout(w_dff_B_b37Hy5GF2_2),.clk(gclk));
	jdff dff_B_YyrSW5Ct5_2(.din(w_dff_B_b37Hy5GF2_2),.dout(w_dff_B_YyrSW5Ct5_2),.clk(gclk));
	jdff dff_B_EsY9RjQV9_2(.din(w_dff_B_YyrSW5Ct5_2),.dout(w_dff_B_EsY9RjQV9_2),.clk(gclk));
	jdff dff_B_QwVvic7U2_2(.din(w_dff_B_EsY9RjQV9_2),.dout(w_dff_B_QwVvic7U2_2),.clk(gclk));
	jdff dff_B_m5itEPoM5_2(.din(w_dff_B_QwVvic7U2_2),.dout(w_dff_B_m5itEPoM5_2),.clk(gclk));
	jdff dff_B_u3HUYTPv7_2(.din(w_dff_B_m5itEPoM5_2),.dout(w_dff_B_u3HUYTPv7_2),.clk(gclk));
	jdff dff_B_ghN2Zun31_2(.din(w_dff_B_u3HUYTPv7_2),.dout(w_dff_B_ghN2Zun31_2),.clk(gclk));
	jdff dff_B_7Ru9YPn77_2(.din(w_dff_B_ghN2Zun31_2),.dout(w_dff_B_7Ru9YPn77_2),.clk(gclk));
	jdff dff_B_nqV95iwg0_2(.din(w_dff_B_7Ru9YPn77_2),.dout(w_dff_B_nqV95iwg0_2),.clk(gclk));
	jdff dff_B_s5Q5PXGk8_2(.din(w_dff_B_nqV95iwg0_2),.dout(w_dff_B_s5Q5PXGk8_2),.clk(gclk));
	jdff dff_B_0gbvO4OC2_2(.din(w_dff_B_s5Q5PXGk8_2),.dout(w_dff_B_0gbvO4OC2_2),.clk(gclk));
	jdff dff_B_MJTELs1G5_2(.din(w_dff_B_0gbvO4OC2_2),.dout(w_dff_B_MJTELs1G5_2),.clk(gclk));
	jdff dff_B_YqQifkcW1_2(.din(w_dff_B_MJTELs1G5_2),.dout(w_dff_B_YqQifkcW1_2),.clk(gclk));
	jdff dff_B_vfPaTgFh9_2(.din(w_dff_B_YqQifkcW1_2),.dout(w_dff_B_vfPaTgFh9_2),.clk(gclk));
	jdff dff_B_N86eqlBb5_2(.din(w_dff_B_vfPaTgFh9_2),.dout(w_dff_B_N86eqlBb5_2),.clk(gclk));
	jdff dff_B_7z0q1ZVd8_2(.din(w_dff_B_N86eqlBb5_2),.dout(w_dff_B_7z0q1ZVd8_2),.clk(gclk));
	jdff dff_B_j1TY1evc6_2(.din(w_dff_B_7z0q1ZVd8_2),.dout(w_dff_B_j1TY1evc6_2),.clk(gclk));
	jdff dff_B_OUtOs0oT9_2(.din(w_dff_B_j1TY1evc6_2),.dout(w_dff_B_OUtOs0oT9_2),.clk(gclk));
	jdff dff_B_XBVwhZ5j4_2(.din(w_dff_B_OUtOs0oT9_2),.dout(w_dff_B_XBVwhZ5j4_2),.clk(gclk));
	jdff dff_B_EZrCr98L4_2(.din(w_dff_B_XBVwhZ5j4_2),.dout(w_dff_B_EZrCr98L4_2),.clk(gclk));
	jdff dff_B_TMTsCZeM5_2(.din(w_dff_B_EZrCr98L4_2),.dout(w_dff_B_TMTsCZeM5_2),.clk(gclk));
	jdff dff_B_KBGpHGoT8_2(.din(w_dff_B_TMTsCZeM5_2),.dout(w_dff_B_KBGpHGoT8_2),.clk(gclk));
	jdff dff_B_VUniCjIM8_2(.din(w_dff_B_KBGpHGoT8_2),.dout(w_dff_B_VUniCjIM8_2),.clk(gclk));
	jdff dff_B_QQSf4ZWy6_2(.din(w_dff_B_VUniCjIM8_2),.dout(w_dff_B_QQSf4ZWy6_2),.clk(gclk));
	jdff dff_B_3AcoKcs97_2(.din(w_dff_B_QQSf4ZWy6_2),.dout(w_dff_B_3AcoKcs97_2),.clk(gclk));
	jdff dff_B_9hxYjqaB7_2(.din(w_dff_B_3AcoKcs97_2),.dout(w_dff_B_9hxYjqaB7_2),.clk(gclk));
	jdff dff_B_c3ReEHRB7_2(.din(w_dff_B_9hxYjqaB7_2),.dout(w_dff_B_c3ReEHRB7_2),.clk(gclk));
	jdff dff_B_R6dPuvtn1_2(.din(n1713),.dout(w_dff_B_R6dPuvtn1_2),.clk(gclk));
	jdff dff_B_4IjTNubv8_2(.din(w_dff_B_R6dPuvtn1_2),.dout(w_dff_B_4IjTNubv8_2),.clk(gclk));
	jdff dff_B_KDL99OvQ5_2(.din(w_dff_B_4IjTNubv8_2),.dout(w_dff_B_KDL99OvQ5_2),.clk(gclk));
	jdff dff_B_z4YZp4Du2_2(.din(w_dff_B_KDL99OvQ5_2),.dout(w_dff_B_z4YZp4Du2_2),.clk(gclk));
	jdff dff_B_3RgO0TWM3_2(.din(w_dff_B_z4YZp4Du2_2),.dout(w_dff_B_3RgO0TWM3_2),.clk(gclk));
	jdff dff_B_eZXbr0V54_2(.din(w_dff_B_3RgO0TWM3_2),.dout(w_dff_B_eZXbr0V54_2),.clk(gclk));
	jdff dff_B_hVJTkY7K6_2(.din(w_dff_B_eZXbr0V54_2),.dout(w_dff_B_hVJTkY7K6_2),.clk(gclk));
	jdff dff_B_bUAIVfIs6_2(.din(w_dff_B_hVJTkY7K6_2),.dout(w_dff_B_bUAIVfIs6_2),.clk(gclk));
	jdff dff_B_BILmwwex7_2(.din(w_dff_B_bUAIVfIs6_2),.dout(w_dff_B_BILmwwex7_2),.clk(gclk));
	jdff dff_B_G7rGZoZ10_2(.din(w_dff_B_BILmwwex7_2),.dout(w_dff_B_G7rGZoZ10_2),.clk(gclk));
	jdff dff_B_TeLTNiLL3_2(.din(w_dff_B_G7rGZoZ10_2),.dout(w_dff_B_TeLTNiLL3_2),.clk(gclk));
	jdff dff_B_rCG0LvIx7_2(.din(w_dff_B_TeLTNiLL3_2),.dout(w_dff_B_rCG0LvIx7_2),.clk(gclk));
	jdff dff_B_DBn2FbCR2_2(.din(w_dff_B_rCG0LvIx7_2),.dout(w_dff_B_DBn2FbCR2_2),.clk(gclk));
	jdff dff_B_b1lEewrK5_2(.din(w_dff_B_DBn2FbCR2_2),.dout(w_dff_B_b1lEewrK5_2),.clk(gclk));
	jdff dff_B_xK1ZFrHW9_2(.din(w_dff_B_b1lEewrK5_2),.dout(w_dff_B_xK1ZFrHW9_2),.clk(gclk));
	jdff dff_B_VcdB7Ems5_2(.din(w_dff_B_xK1ZFrHW9_2),.dout(w_dff_B_VcdB7Ems5_2),.clk(gclk));
	jdff dff_B_FXNntc2K9_2(.din(w_dff_B_VcdB7Ems5_2),.dout(w_dff_B_FXNntc2K9_2),.clk(gclk));
	jdff dff_B_mYwqHzcf8_2(.din(w_dff_B_FXNntc2K9_2),.dout(w_dff_B_mYwqHzcf8_2),.clk(gclk));
	jdff dff_B_atQJYgGv5_2(.din(w_dff_B_mYwqHzcf8_2),.dout(w_dff_B_atQJYgGv5_2),.clk(gclk));
	jdff dff_B_1NwKVTvC7_2(.din(w_dff_B_atQJYgGv5_2),.dout(w_dff_B_1NwKVTvC7_2),.clk(gclk));
	jdff dff_B_h0WYMxQh4_2(.din(w_dff_B_1NwKVTvC7_2),.dout(w_dff_B_h0WYMxQh4_2),.clk(gclk));
	jdff dff_B_xgZmrLAf0_2(.din(w_dff_B_h0WYMxQh4_2),.dout(w_dff_B_xgZmrLAf0_2),.clk(gclk));
	jdff dff_B_S2YyZGEL4_2(.din(w_dff_B_xgZmrLAf0_2),.dout(w_dff_B_S2YyZGEL4_2),.clk(gclk));
	jdff dff_B_E1c6ZsQY3_2(.din(w_dff_B_S2YyZGEL4_2),.dout(w_dff_B_E1c6ZsQY3_2),.clk(gclk));
	jdff dff_B_lYb19zPu5_2(.din(w_dff_B_E1c6ZsQY3_2),.dout(w_dff_B_lYb19zPu5_2),.clk(gclk));
	jdff dff_B_hCE862NY2_2(.din(w_dff_B_lYb19zPu5_2),.dout(w_dff_B_hCE862NY2_2),.clk(gclk));
	jdff dff_B_3uhZAm128_2(.din(w_dff_B_hCE862NY2_2),.dout(w_dff_B_3uhZAm128_2),.clk(gclk));
	jdff dff_B_ppVyT4Hw5_2(.din(w_dff_B_3uhZAm128_2),.dout(w_dff_B_ppVyT4Hw5_2),.clk(gclk));
	jdff dff_B_KZxWwOwg2_2(.din(w_dff_B_ppVyT4Hw5_2),.dout(w_dff_B_KZxWwOwg2_2),.clk(gclk));
	jdff dff_B_eEqE2GBI5_2(.din(w_dff_B_KZxWwOwg2_2),.dout(w_dff_B_eEqE2GBI5_2),.clk(gclk));
	jdff dff_B_f1YAp7Xu1_2(.din(w_dff_B_eEqE2GBI5_2),.dout(w_dff_B_f1YAp7Xu1_2),.clk(gclk));
	jdff dff_B_yudoXnwW9_2(.din(w_dff_B_f1YAp7Xu1_2),.dout(w_dff_B_yudoXnwW9_2),.clk(gclk));
	jdff dff_B_icYVq9Sk3_2(.din(w_dff_B_yudoXnwW9_2),.dout(w_dff_B_icYVq9Sk3_2),.clk(gclk));
	jdff dff_B_06cP4HMr5_2(.din(w_dff_B_icYVq9Sk3_2),.dout(w_dff_B_06cP4HMr5_2),.clk(gclk));
	jdff dff_B_eSa1ax943_2(.din(w_dff_B_06cP4HMr5_2),.dout(w_dff_B_eSa1ax943_2),.clk(gclk));
	jdff dff_B_NLyXDzBG8_2(.din(w_dff_B_eSa1ax943_2),.dout(w_dff_B_NLyXDzBG8_2),.clk(gclk));
	jdff dff_B_hXHlc8EP3_2(.din(w_dff_B_NLyXDzBG8_2),.dout(w_dff_B_hXHlc8EP3_2),.clk(gclk));
	jdff dff_B_Mc8N4V6c1_2(.din(w_dff_B_hXHlc8EP3_2),.dout(w_dff_B_Mc8N4V6c1_2),.clk(gclk));
	jdff dff_B_vcIT8ORZ9_2(.din(w_dff_B_Mc8N4V6c1_2),.dout(w_dff_B_vcIT8ORZ9_2),.clk(gclk));
	jdff dff_B_MmA9o2Px5_2(.din(w_dff_B_vcIT8ORZ9_2),.dout(w_dff_B_MmA9o2Px5_2),.clk(gclk));
	jdff dff_B_U9sq9dXx5_2(.din(w_dff_B_MmA9o2Px5_2),.dout(w_dff_B_U9sq9dXx5_2),.clk(gclk));
	jdff dff_B_fjff3wPx7_2(.din(w_dff_B_U9sq9dXx5_2),.dout(w_dff_B_fjff3wPx7_2),.clk(gclk));
	jdff dff_B_VE9RbqXC4_2(.din(w_dff_B_fjff3wPx7_2),.dout(w_dff_B_VE9RbqXC4_2),.clk(gclk));
	jdff dff_B_tXWfrrrp7_2(.din(n1712),.dout(w_dff_B_tXWfrrrp7_2),.clk(gclk));
	jdff dff_B_RYVMzpN97_1(.din(n1710),.dout(w_dff_B_RYVMzpN97_1),.clk(gclk));
	jdff dff_B_x9c3PDcI7_2(.din(n1668),.dout(w_dff_B_x9c3PDcI7_2),.clk(gclk));
	jdff dff_B_BnFDsRGs0_2(.din(w_dff_B_x9c3PDcI7_2),.dout(w_dff_B_BnFDsRGs0_2),.clk(gclk));
	jdff dff_B_K2L8qRO92_2(.din(w_dff_B_BnFDsRGs0_2),.dout(w_dff_B_K2L8qRO92_2),.clk(gclk));
	jdff dff_B_5xNigKaC1_2(.din(w_dff_B_K2L8qRO92_2),.dout(w_dff_B_5xNigKaC1_2),.clk(gclk));
	jdff dff_B_GqmQDBGx2_2(.din(w_dff_B_5xNigKaC1_2),.dout(w_dff_B_GqmQDBGx2_2),.clk(gclk));
	jdff dff_B_0QCbbunV0_2(.din(w_dff_B_GqmQDBGx2_2),.dout(w_dff_B_0QCbbunV0_2),.clk(gclk));
	jdff dff_B_qUWE1KkA6_2(.din(w_dff_B_0QCbbunV0_2),.dout(w_dff_B_qUWE1KkA6_2),.clk(gclk));
	jdff dff_B_sj9Xg9yW2_2(.din(w_dff_B_qUWE1KkA6_2),.dout(w_dff_B_sj9Xg9yW2_2),.clk(gclk));
	jdff dff_B_TRHFsr1R0_2(.din(w_dff_B_sj9Xg9yW2_2),.dout(w_dff_B_TRHFsr1R0_2),.clk(gclk));
	jdff dff_B_LXdu0AkO8_2(.din(w_dff_B_TRHFsr1R0_2),.dout(w_dff_B_LXdu0AkO8_2),.clk(gclk));
	jdff dff_B_AKixe2ru9_2(.din(w_dff_B_LXdu0AkO8_2),.dout(w_dff_B_AKixe2ru9_2),.clk(gclk));
	jdff dff_B_30HM3AC04_2(.din(w_dff_B_AKixe2ru9_2),.dout(w_dff_B_30HM3AC04_2),.clk(gclk));
	jdff dff_B_N6nEW1yV9_2(.din(w_dff_B_30HM3AC04_2),.dout(w_dff_B_N6nEW1yV9_2),.clk(gclk));
	jdff dff_B_KKSF2tfy0_2(.din(w_dff_B_N6nEW1yV9_2),.dout(w_dff_B_KKSF2tfy0_2),.clk(gclk));
	jdff dff_B_ZwrOPPdG9_2(.din(w_dff_B_KKSF2tfy0_2),.dout(w_dff_B_ZwrOPPdG9_2),.clk(gclk));
	jdff dff_B_R15dqJNn9_2(.din(w_dff_B_ZwrOPPdG9_2),.dout(w_dff_B_R15dqJNn9_2),.clk(gclk));
	jdff dff_B_xii39iJq9_2(.din(w_dff_B_R15dqJNn9_2),.dout(w_dff_B_xii39iJq9_2),.clk(gclk));
	jdff dff_B_YKI5l6Hs2_2(.din(w_dff_B_xii39iJq9_2),.dout(w_dff_B_YKI5l6Hs2_2),.clk(gclk));
	jdff dff_B_aIPBVgCe1_2(.din(w_dff_B_YKI5l6Hs2_2),.dout(w_dff_B_aIPBVgCe1_2),.clk(gclk));
	jdff dff_B_5O9epzDr1_2(.din(w_dff_B_aIPBVgCe1_2),.dout(w_dff_B_5O9epzDr1_2),.clk(gclk));
	jdff dff_B_tzDgVItv0_2(.din(w_dff_B_5O9epzDr1_2),.dout(w_dff_B_tzDgVItv0_2),.clk(gclk));
	jdff dff_B_iA10L69m2_2(.din(w_dff_B_tzDgVItv0_2),.dout(w_dff_B_iA10L69m2_2),.clk(gclk));
	jdff dff_B_2oWl4rML9_2(.din(w_dff_B_iA10L69m2_2),.dout(w_dff_B_2oWl4rML9_2),.clk(gclk));
	jdff dff_B_13pGjisS0_2(.din(w_dff_B_2oWl4rML9_2),.dout(w_dff_B_13pGjisS0_2),.clk(gclk));
	jdff dff_B_C2Wc6Wvw6_2(.din(w_dff_B_13pGjisS0_2),.dout(w_dff_B_C2Wc6Wvw6_2),.clk(gclk));
	jdff dff_B_s78V3ezX4_2(.din(w_dff_B_C2Wc6Wvw6_2),.dout(w_dff_B_s78V3ezX4_2),.clk(gclk));
	jdff dff_B_Tv2e50Nm6_2(.din(w_dff_B_s78V3ezX4_2),.dout(w_dff_B_Tv2e50Nm6_2),.clk(gclk));
	jdff dff_B_V729JHOL8_2(.din(w_dff_B_Tv2e50Nm6_2),.dout(w_dff_B_V729JHOL8_2),.clk(gclk));
	jdff dff_B_ECinXe1W0_2(.din(w_dff_B_V729JHOL8_2),.dout(w_dff_B_ECinXe1W0_2),.clk(gclk));
	jdff dff_B_T98C3kRf7_2(.din(w_dff_B_ECinXe1W0_2),.dout(w_dff_B_T98C3kRf7_2),.clk(gclk));
	jdff dff_B_Ve65sJdP7_2(.din(w_dff_B_T98C3kRf7_2),.dout(w_dff_B_Ve65sJdP7_2),.clk(gclk));
	jdff dff_B_2NtWCb7J9_2(.din(w_dff_B_Ve65sJdP7_2),.dout(w_dff_B_2NtWCb7J9_2),.clk(gclk));
	jdff dff_B_ESrSLO466_2(.din(w_dff_B_2NtWCb7J9_2),.dout(w_dff_B_ESrSLO466_2),.clk(gclk));
	jdff dff_B_ffJ3eKLO3_2(.din(w_dff_B_ESrSLO466_2),.dout(w_dff_B_ffJ3eKLO3_2),.clk(gclk));
	jdff dff_B_sYSEjoPj5_2(.din(w_dff_B_ffJ3eKLO3_2),.dout(w_dff_B_sYSEjoPj5_2),.clk(gclk));
	jdff dff_B_cvo0OhbJ5_2(.din(w_dff_B_sYSEjoPj5_2),.dout(w_dff_B_cvo0OhbJ5_2),.clk(gclk));
	jdff dff_B_NBaznYtg5_2(.din(w_dff_B_cvo0OhbJ5_2),.dout(w_dff_B_NBaznYtg5_2),.clk(gclk));
	jdff dff_B_D9nY5kld8_2(.din(w_dff_B_NBaznYtg5_2),.dout(w_dff_B_D9nY5kld8_2),.clk(gclk));
	jdff dff_B_nxNT8YVZ2_2(.din(w_dff_B_D9nY5kld8_2),.dout(w_dff_B_nxNT8YVZ2_2),.clk(gclk));
	jdff dff_B_d19QqC920_2(.din(w_dff_B_nxNT8YVZ2_2),.dout(w_dff_B_d19QqC920_2),.clk(gclk));
	jdff dff_B_qFz2i5bZ3_1(.din(n1674),.dout(w_dff_B_qFz2i5bZ3_1),.clk(gclk));
	jdff dff_B_BS5jlJis8_1(.din(w_dff_B_qFz2i5bZ3_1),.dout(w_dff_B_BS5jlJis8_1),.clk(gclk));
	jdff dff_B_BCHZwWHr9_2(.din(n1673),.dout(w_dff_B_BCHZwWHr9_2),.clk(gclk));
	jdff dff_B_3NkGgqFD3_2(.din(w_dff_B_BCHZwWHr9_2),.dout(w_dff_B_3NkGgqFD3_2),.clk(gclk));
	jdff dff_B_iOzz3uqc4_2(.din(w_dff_B_3NkGgqFD3_2),.dout(w_dff_B_iOzz3uqc4_2),.clk(gclk));
	jdff dff_B_PeJBjRHi5_2(.din(w_dff_B_iOzz3uqc4_2),.dout(w_dff_B_PeJBjRHi5_2),.clk(gclk));
	jdff dff_B_R2pf6reC5_2(.din(w_dff_B_PeJBjRHi5_2),.dout(w_dff_B_R2pf6reC5_2),.clk(gclk));
	jdff dff_B_xrSvcZms1_2(.din(w_dff_B_R2pf6reC5_2),.dout(w_dff_B_xrSvcZms1_2),.clk(gclk));
	jdff dff_B_A4JIWXhJ2_2(.din(w_dff_B_xrSvcZms1_2),.dout(w_dff_B_A4JIWXhJ2_2),.clk(gclk));
	jdff dff_B_iJLRGmSm9_2(.din(w_dff_B_A4JIWXhJ2_2),.dout(w_dff_B_iJLRGmSm9_2),.clk(gclk));
	jdff dff_B_9wXZ4drW7_2(.din(w_dff_B_iJLRGmSm9_2),.dout(w_dff_B_9wXZ4drW7_2),.clk(gclk));
	jdff dff_B_H6k7qUr83_2(.din(w_dff_B_9wXZ4drW7_2),.dout(w_dff_B_H6k7qUr83_2),.clk(gclk));
	jdff dff_B_rnR2EMVn3_2(.din(w_dff_B_H6k7qUr83_2),.dout(w_dff_B_rnR2EMVn3_2),.clk(gclk));
	jdff dff_B_cyYKyTcW9_2(.din(w_dff_B_rnR2EMVn3_2),.dout(w_dff_B_cyYKyTcW9_2),.clk(gclk));
	jdff dff_B_LG6HglGr7_2(.din(w_dff_B_cyYKyTcW9_2),.dout(w_dff_B_LG6HglGr7_2),.clk(gclk));
	jdff dff_B_4dF0UD2E1_2(.din(w_dff_B_LG6HglGr7_2),.dout(w_dff_B_4dF0UD2E1_2),.clk(gclk));
	jdff dff_B_7sVx1Bbz7_2(.din(w_dff_B_4dF0UD2E1_2),.dout(w_dff_B_7sVx1Bbz7_2),.clk(gclk));
	jdff dff_B_Yk6VcBVx3_2(.din(w_dff_B_7sVx1Bbz7_2),.dout(w_dff_B_Yk6VcBVx3_2),.clk(gclk));
	jdff dff_B_SvkAqVdf6_2(.din(w_dff_B_Yk6VcBVx3_2),.dout(w_dff_B_SvkAqVdf6_2),.clk(gclk));
	jdff dff_B_eTpezwir6_2(.din(w_dff_B_SvkAqVdf6_2),.dout(w_dff_B_eTpezwir6_2),.clk(gclk));
	jdff dff_B_Fv2vJcsU0_2(.din(w_dff_B_eTpezwir6_2),.dout(w_dff_B_Fv2vJcsU0_2),.clk(gclk));
	jdff dff_B_yw91nAdB1_2(.din(w_dff_B_Fv2vJcsU0_2),.dout(w_dff_B_yw91nAdB1_2),.clk(gclk));
	jdff dff_B_nt4QY3Pc6_2(.din(w_dff_B_yw91nAdB1_2),.dout(w_dff_B_nt4QY3Pc6_2),.clk(gclk));
	jdff dff_B_OCJ0P7RE3_2(.din(w_dff_B_nt4QY3Pc6_2),.dout(w_dff_B_OCJ0P7RE3_2),.clk(gclk));
	jdff dff_B_TPbdEi4f0_2(.din(w_dff_B_OCJ0P7RE3_2),.dout(w_dff_B_TPbdEi4f0_2),.clk(gclk));
	jdff dff_B_hmxQUuYV9_2(.din(w_dff_B_TPbdEi4f0_2),.dout(w_dff_B_hmxQUuYV9_2),.clk(gclk));
	jdff dff_B_OVrobNsX7_2(.din(w_dff_B_hmxQUuYV9_2),.dout(w_dff_B_OVrobNsX7_2),.clk(gclk));
	jdff dff_B_QtWt3vGn0_2(.din(w_dff_B_OVrobNsX7_2),.dout(w_dff_B_QtWt3vGn0_2),.clk(gclk));
	jdff dff_B_EizkcA7N0_2(.din(w_dff_B_QtWt3vGn0_2),.dout(w_dff_B_EizkcA7N0_2),.clk(gclk));
	jdff dff_B_7iGNFEju4_2(.din(w_dff_B_EizkcA7N0_2),.dout(w_dff_B_7iGNFEju4_2),.clk(gclk));
	jdff dff_B_qDCwc2Dl8_2(.din(w_dff_B_7iGNFEju4_2),.dout(w_dff_B_qDCwc2Dl8_2),.clk(gclk));
	jdff dff_B_UhItJk2c3_2(.din(w_dff_B_qDCwc2Dl8_2),.dout(w_dff_B_UhItJk2c3_2),.clk(gclk));
	jdff dff_B_YRbCoiYw2_2(.din(w_dff_B_UhItJk2c3_2),.dout(w_dff_B_YRbCoiYw2_2),.clk(gclk));
	jdff dff_B_cDJB2DsX7_2(.din(w_dff_B_YRbCoiYw2_2),.dout(w_dff_B_cDJB2DsX7_2),.clk(gclk));
	jdff dff_B_sWYheQJS9_2(.din(w_dff_B_cDJB2DsX7_2),.dout(w_dff_B_sWYheQJS9_2),.clk(gclk));
	jdff dff_B_pq2DPpZI7_2(.din(w_dff_B_sWYheQJS9_2),.dout(w_dff_B_pq2DPpZI7_2),.clk(gclk));
	jdff dff_B_1vPSXQt52_2(.din(w_dff_B_pq2DPpZI7_2),.dout(w_dff_B_1vPSXQt52_2),.clk(gclk));
	jdff dff_B_MWLO8jro5_2(.din(w_dff_B_1vPSXQt52_2),.dout(w_dff_B_MWLO8jro5_2),.clk(gclk));
	jdff dff_B_uCOPYHHr4_2(.din(w_dff_B_MWLO8jro5_2),.dout(w_dff_B_uCOPYHHr4_2),.clk(gclk));
	jdff dff_B_cMaruJZQ5_2(.din(n1672),.dout(w_dff_B_cMaruJZQ5_2),.clk(gclk));
	jdff dff_B_uYUlhEFw7_2(.din(w_dff_B_cMaruJZQ5_2),.dout(w_dff_B_uYUlhEFw7_2),.clk(gclk));
	jdff dff_B_8IVAGVyn6_2(.din(w_dff_B_uYUlhEFw7_2),.dout(w_dff_B_8IVAGVyn6_2),.clk(gclk));
	jdff dff_B_DQwNWSSj5_2(.din(w_dff_B_8IVAGVyn6_2),.dout(w_dff_B_DQwNWSSj5_2),.clk(gclk));
	jdff dff_B_yVi6PexV2_2(.din(w_dff_B_DQwNWSSj5_2),.dout(w_dff_B_yVi6PexV2_2),.clk(gclk));
	jdff dff_B_2smYxZgT2_2(.din(w_dff_B_yVi6PexV2_2),.dout(w_dff_B_2smYxZgT2_2),.clk(gclk));
	jdff dff_B_Pi5g5RIl7_2(.din(w_dff_B_2smYxZgT2_2),.dout(w_dff_B_Pi5g5RIl7_2),.clk(gclk));
	jdff dff_B_HClIwoj19_2(.din(w_dff_B_Pi5g5RIl7_2),.dout(w_dff_B_HClIwoj19_2),.clk(gclk));
	jdff dff_B_FnMWYGRF4_2(.din(w_dff_B_HClIwoj19_2),.dout(w_dff_B_FnMWYGRF4_2),.clk(gclk));
	jdff dff_B_W6lJyYdW8_2(.din(w_dff_B_FnMWYGRF4_2),.dout(w_dff_B_W6lJyYdW8_2),.clk(gclk));
	jdff dff_B_e8CvEH3I0_2(.din(w_dff_B_W6lJyYdW8_2),.dout(w_dff_B_e8CvEH3I0_2),.clk(gclk));
	jdff dff_B_NGhIjFql9_2(.din(w_dff_B_e8CvEH3I0_2),.dout(w_dff_B_NGhIjFql9_2),.clk(gclk));
	jdff dff_B_IF2z2di74_2(.din(w_dff_B_NGhIjFql9_2),.dout(w_dff_B_IF2z2di74_2),.clk(gclk));
	jdff dff_B_JPAaHdeJ3_2(.din(w_dff_B_IF2z2di74_2),.dout(w_dff_B_JPAaHdeJ3_2),.clk(gclk));
	jdff dff_B_1Nh4SGeK5_2(.din(w_dff_B_JPAaHdeJ3_2),.dout(w_dff_B_1Nh4SGeK5_2),.clk(gclk));
	jdff dff_B_q1FL87Rh1_2(.din(w_dff_B_1Nh4SGeK5_2),.dout(w_dff_B_q1FL87Rh1_2),.clk(gclk));
	jdff dff_B_HsRMh7uS3_2(.din(w_dff_B_q1FL87Rh1_2),.dout(w_dff_B_HsRMh7uS3_2),.clk(gclk));
	jdff dff_B_sf0OTIXx8_2(.din(w_dff_B_HsRMh7uS3_2),.dout(w_dff_B_sf0OTIXx8_2),.clk(gclk));
	jdff dff_B_SvxVQAP35_2(.din(w_dff_B_sf0OTIXx8_2),.dout(w_dff_B_SvxVQAP35_2),.clk(gclk));
	jdff dff_B_NKRMDZ1O4_2(.din(w_dff_B_SvxVQAP35_2),.dout(w_dff_B_NKRMDZ1O4_2),.clk(gclk));
	jdff dff_B_XgX7ehYZ6_2(.din(w_dff_B_NKRMDZ1O4_2),.dout(w_dff_B_XgX7ehYZ6_2),.clk(gclk));
	jdff dff_B_HkMirg7a2_2(.din(w_dff_B_XgX7ehYZ6_2),.dout(w_dff_B_HkMirg7a2_2),.clk(gclk));
	jdff dff_B_M7ywZa7k3_2(.din(w_dff_B_HkMirg7a2_2),.dout(w_dff_B_M7ywZa7k3_2),.clk(gclk));
	jdff dff_B_cP0VlKjz8_2(.din(w_dff_B_M7ywZa7k3_2),.dout(w_dff_B_cP0VlKjz8_2),.clk(gclk));
	jdff dff_B_eA3Yygsi4_2(.din(w_dff_B_cP0VlKjz8_2),.dout(w_dff_B_eA3Yygsi4_2),.clk(gclk));
	jdff dff_B_S3H5TUMo6_2(.din(w_dff_B_eA3Yygsi4_2),.dout(w_dff_B_S3H5TUMo6_2),.clk(gclk));
	jdff dff_B_gtNkzfLy2_2(.din(w_dff_B_S3H5TUMo6_2),.dout(w_dff_B_gtNkzfLy2_2),.clk(gclk));
	jdff dff_B_T2vebjFV1_2(.din(w_dff_B_gtNkzfLy2_2),.dout(w_dff_B_T2vebjFV1_2),.clk(gclk));
	jdff dff_B_HX5HcSot8_2(.din(w_dff_B_T2vebjFV1_2),.dout(w_dff_B_HX5HcSot8_2),.clk(gclk));
	jdff dff_B_WLbUSyTF1_2(.din(w_dff_B_HX5HcSot8_2),.dout(w_dff_B_WLbUSyTF1_2),.clk(gclk));
	jdff dff_B_RCKDo9C86_2(.din(w_dff_B_WLbUSyTF1_2),.dout(w_dff_B_RCKDo9C86_2),.clk(gclk));
	jdff dff_B_cSOKipbt9_2(.din(w_dff_B_RCKDo9C86_2),.dout(w_dff_B_cSOKipbt9_2),.clk(gclk));
	jdff dff_B_OqUJ9lt96_2(.din(w_dff_B_cSOKipbt9_2),.dout(w_dff_B_OqUJ9lt96_2),.clk(gclk));
	jdff dff_B_4knkifYT9_2(.din(w_dff_B_OqUJ9lt96_2),.dout(w_dff_B_4knkifYT9_2),.clk(gclk));
	jdff dff_B_Y81BF20X9_2(.din(w_dff_B_4knkifYT9_2),.dout(w_dff_B_Y81BF20X9_2),.clk(gclk));
	jdff dff_B_E0W5cjBN1_2(.din(w_dff_B_Y81BF20X9_2),.dout(w_dff_B_E0W5cjBN1_2),.clk(gclk));
	jdff dff_B_tJ9cO7eA7_2(.din(w_dff_B_E0W5cjBN1_2),.dout(w_dff_B_tJ9cO7eA7_2),.clk(gclk));
	jdff dff_B_jDunCeCm0_2(.din(w_dff_B_tJ9cO7eA7_2),.dout(w_dff_B_jDunCeCm0_2),.clk(gclk));
	jdff dff_B_qm4Xdjn60_2(.din(w_dff_B_jDunCeCm0_2),.dout(w_dff_B_qm4Xdjn60_2),.clk(gclk));
	jdff dff_B_KI6zkGY98_2(.din(n1671),.dout(w_dff_B_KI6zkGY98_2),.clk(gclk));
	jdff dff_B_ntwO1BtR6_1(.din(n1669),.dout(w_dff_B_ntwO1BtR6_1),.clk(gclk));
	jdff dff_B_YMrTLbXo8_2(.din(n1617),.dout(w_dff_B_YMrTLbXo8_2),.clk(gclk));
	jdff dff_B_Dj5C2tG87_2(.din(w_dff_B_YMrTLbXo8_2),.dout(w_dff_B_Dj5C2tG87_2),.clk(gclk));
	jdff dff_B_B9Q1NcNt9_2(.din(w_dff_B_Dj5C2tG87_2),.dout(w_dff_B_B9Q1NcNt9_2),.clk(gclk));
	jdff dff_B_LJcV8DAo4_2(.din(w_dff_B_B9Q1NcNt9_2),.dout(w_dff_B_LJcV8DAo4_2),.clk(gclk));
	jdff dff_B_yU9GDdmy5_2(.din(w_dff_B_LJcV8DAo4_2),.dout(w_dff_B_yU9GDdmy5_2),.clk(gclk));
	jdff dff_B_oj6I1fhT7_2(.din(w_dff_B_yU9GDdmy5_2),.dout(w_dff_B_oj6I1fhT7_2),.clk(gclk));
	jdff dff_B_p1friQVX9_2(.din(w_dff_B_oj6I1fhT7_2),.dout(w_dff_B_p1friQVX9_2),.clk(gclk));
	jdff dff_B_EPbDH7YQ4_2(.din(w_dff_B_p1friQVX9_2),.dout(w_dff_B_EPbDH7YQ4_2),.clk(gclk));
	jdff dff_B_MAqHVTY94_2(.din(w_dff_B_EPbDH7YQ4_2),.dout(w_dff_B_MAqHVTY94_2),.clk(gclk));
	jdff dff_B_P2H9yM5T1_2(.din(w_dff_B_MAqHVTY94_2),.dout(w_dff_B_P2H9yM5T1_2),.clk(gclk));
	jdff dff_B_DC05vVfq0_2(.din(w_dff_B_P2H9yM5T1_2),.dout(w_dff_B_DC05vVfq0_2),.clk(gclk));
	jdff dff_B_CA1fzLZ38_2(.din(w_dff_B_DC05vVfq0_2),.dout(w_dff_B_CA1fzLZ38_2),.clk(gclk));
	jdff dff_B_RHvCyUSp5_2(.din(w_dff_B_CA1fzLZ38_2),.dout(w_dff_B_RHvCyUSp5_2),.clk(gclk));
	jdff dff_B_jqEfmEm42_2(.din(w_dff_B_RHvCyUSp5_2),.dout(w_dff_B_jqEfmEm42_2),.clk(gclk));
	jdff dff_B_WrKoJqVN5_2(.din(w_dff_B_jqEfmEm42_2),.dout(w_dff_B_WrKoJqVN5_2),.clk(gclk));
	jdff dff_B_mtWdbZf87_2(.din(w_dff_B_WrKoJqVN5_2),.dout(w_dff_B_mtWdbZf87_2),.clk(gclk));
	jdff dff_B_Cl1VHnoQ1_2(.din(w_dff_B_mtWdbZf87_2),.dout(w_dff_B_Cl1VHnoQ1_2),.clk(gclk));
	jdff dff_B_8nwFrqKH8_2(.din(w_dff_B_Cl1VHnoQ1_2),.dout(w_dff_B_8nwFrqKH8_2),.clk(gclk));
	jdff dff_B_7xNJ6RWm7_2(.din(w_dff_B_8nwFrqKH8_2),.dout(w_dff_B_7xNJ6RWm7_2),.clk(gclk));
	jdff dff_B_DuCTP03u4_2(.din(w_dff_B_7xNJ6RWm7_2),.dout(w_dff_B_DuCTP03u4_2),.clk(gclk));
	jdff dff_B_irzoq4BI7_2(.din(w_dff_B_DuCTP03u4_2),.dout(w_dff_B_irzoq4BI7_2),.clk(gclk));
	jdff dff_B_GPPHDsy27_2(.din(w_dff_B_irzoq4BI7_2),.dout(w_dff_B_GPPHDsy27_2),.clk(gclk));
	jdff dff_B_wCPdB5n86_2(.din(w_dff_B_GPPHDsy27_2),.dout(w_dff_B_wCPdB5n86_2),.clk(gclk));
	jdff dff_B_H55aBVAt2_2(.din(w_dff_B_wCPdB5n86_2),.dout(w_dff_B_H55aBVAt2_2),.clk(gclk));
	jdff dff_B_3qhzTdwb9_2(.din(w_dff_B_H55aBVAt2_2),.dout(w_dff_B_3qhzTdwb9_2),.clk(gclk));
	jdff dff_B_DTuG6Slf4_2(.din(w_dff_B_3qhzTdwb9_2),.dout(w_dff_B_DTuG6Slf4_2),.clk(gclk));
	jdff dff_B_wwpDl90J9_2(.din(w_dff_B_DTuG6Slf4_2),.dout(w_dff_B_wwpDl90J9_2),.clk(gclk));
	jdff dff_B_fjSPGuSj6_2(.din(w_dff_B_wwpDl90J9_2),.dout(w_dff_B_fjSPGuSj6_2),.clk(gclk));
	jdff dff_B_KmBnLnlX7_2(.din(w_dff_B_fjSPGuSj6_2),.dout(w_dff_B_KmBnLnlX7_2),.clk(gclk));
	jdff dff_B_mmDMY6Gu5_2(.din(w_dff_B_KmBnLnlX7_2),.dout(w_dff_B_mmDMY6Gu5_2),.clk(gclk));
	jdff dff_B_au2uUdBm4_2(.din(w_dff_B_mmDMY6Gu5_2),.dout(w_dff_B_au2uUdBm4_2),.clk(gclk));
	jdff dff_B_wB5uG7jW4_2(.din(w_dff_B_au2uUdBm4_2),.dout(w_dff_B_wB5uG7jW4_2),.clk(gclk));
	jdff dff_B_SK2KFuYW8_2(.din(w_dff_B_wB5uG7jW4_2),.dout(w_dff_B_SK2KFuYW8_2),.clk(gclk));
	jdff dff_B_RLTDLljs4_2(.din(w_dff_B_SK2KFuYW8_2),.dout(w_dff_B_RLTDLljs4_2),.clk(gclk));
	jdff dff_B_a3whaK1s3_2(.din(w_dff_B_RLTDLljs4_2),.dout(w_dff_B_a3whaK1s3_2),.clk(gclk));
	jdff dff_B_tYEo24vg1_2(.din(w_dff_B_a3whaK1s3_2),.dout(w_dff_B_tYEo24vg1_2),.clk(gclk));
	jdff dff_B_jL5LBRT13_1(.din(n1623),.dout(w_dff_B_jL5LBRT13_1),.clk(gclk));
	jdff dff_B_CDUyJ6Ha0_1(.din(w_dff_B_jL5LBRT13_1),.dout(w_dff_B_CDUyJ6Ha0_1),.clk(gclk));
	jdff dff_B_lu2c9jbA0_2(.din(n1622),.dout(w_dff_B_lu2c9jbA0_2),.clk(gclk));
	jdff dff_B_MLfHG4xb3_2(.din(w_dff_B_lu2c9jbA0_2),.dout(w_dff_B_MLfHG4xb3_2),.clk(gclk));
	jdff dff_B_cQ1pxbYt1_2(.din(w_dff_B_MLfHG4xb3_2),.dout(w_dff_B_cQ1pxbYt1_2),.clk(gclk));
	jdff dff_B_2U6o0fJL7_2(.din(w_dff_B_cQ1pxbYt1_2),.dout(w_dff_B_2U6o0fJL7_2),.clk(gclk));
	jdff dff_B_3F2oAwlg3_2(.din(w_dff_B_2U6o0fJL7_2),.dout(w_dff_B_3F2oAwlg3_2),.clk(gclk));
	jdff dff_B_xJSs3pD08_2(.din(w_dff_B_3F2oAwlg3_2),.dout(w_dff_B_xJSs3pD08_2),.clk(gclk));
	jdff dff_B_b2iPkQUb6_2(.din(w_dff_B_xJSs3pD08_2),.dout(w_dff_B_b2iPkQUb6_2),.clk(gclk));
	jdff dff_B_wt3HlLd44_2(.din(w_dff_B_b2iPkQUb6_2),.dout(w_dff_B_wt3HlLd44_2),.clk(gclk));
	jdff dff_B_uGAakRTN8_2(.din(w_dff_B_wt3HlLd44_2),.dout(w_dff_B_uGAakRTN8_2),.clk(gclk));
	jdff dff_B_rdEeYATn5_2(.din(w_dff_B_uGAakRTN8_2),.dout(w_dff_B_rdEeYATn5_2),.clk(gclk));
	jdff dff_B_60CvUXGm4_2(.din(w_dff_B_rdEeYATn5_2),.dout(w_dff_B_60CvUXGm4_2),.clk(gclk));
	jdff dff_B_p2OyUcxS9_2(.din(w_dff_B_60CvUXGm4_2),.dout(w_dff_B_p2OyUcxS9_2),.clk(gclk));
	jdff dff_B_9CfXGiuI0_2(.din(w_dff_B_p2OyUcxS9_2),.dout(w_dff_B_9CfXGiuI0_2),.clk(gclk));
	jdff dff_B_OvTsoxPy4_2(.din(w_dff_B_9CfXGiuI0_2),.dout(w_dff_B_OvTsoxPy4_2),.clk(gclk));
	jdff dff_B_rTQelcBA9_2(.din(w_dff_B_OvTsoxPy4_2),.dout(w_dff_B_rTQelcBA9_2),.clk(gclk));
	jdff dff_B_8D96CdCl9_2(.din(w_dff_B_rTQelcBA9_2),.dout(w_dff_B_8D96CdCl9_2),.clk(gclk));
	jdff dff_B_OVG0goZC9_2(.din(w_dff_B_8D96CdCl9_2),.dout(w_dff_B_OVG0goZC9_2),.clk(gclk));
	jdff dff_B_acOnO6Zc4_2(.din(w_dff_B_OVG0goZC9_2),.dout(w_dff_B_acOnO6Zc4_2),.clk(gclk));
	jdff dff_B_9J3eSEQu2_2(.din(w_dff_B_acOnO6Zc4_2),.dout(w_dff_B_9J3eSEQu2_2),.clk(gclk));
	jdff dff_B_35gb3vVg5_2(.din(w_dff_B_9J3eSEQu2_2),.dout(w_dff_B_35gb3vVg5_2),.clk(gclk));
	jdff dff_B_2SA6zfzj1_2(.din(w_dff_B_35gb3vVg5_2),.dout(w_dff_B_2SA6zfzj1_2),.clk(gclk));
	jdff dff_B_jd3EjMk98_2(.din(w_dff_B_2SA6zfzj1_2),.dout(w_dff_B_jd3EjMk98_2),.clk(gclk));
	jdff dff_B_6OpeuCrB2_2(.din(w_dff_B_jd3EjMk98_2),.dout(w_dff_B_6OpeuCrB2_2),.clk(gclk));
	jdff dff_B_aGn6E8B36_2(.din(w_dff_B_6OpeuCrB2_2),.dout(w_dff_B_aGn6E8B36_2),.clk(gclk));
	jdff dff_B_v1pevEXP2_2(.din(w_dff_B_aGn6E8B36_2),.dout(w_dff_B_v1pevEXP2_2),.clk(gclk));
	jdff dff_B_D4ssf82m6_2(.din(w_dff_B_v1pevEXP2_2),.dout(w_dff_B_D4ssf82m6_2),.clk(gclk));
	jdff dff_B_y1v2CbCH9_2(.din(w_dff_B_D4ssf82m6_2),.dout(w_dff_B_y1v2CbCH9_2),.clk(gclk));
	jdff dff_B_sYk5t9Lx0_2(.din(w_dff_B_y1v2CbCH9_2),.dout(w_dff_B_sYk5t9Lx0_2),.clk(gclk));
	jdff dff_B_AKirHMAn0_2(.din(w_dff_B_sYk5t9Lx0_2),.dout(w_dff_B_AKirHMAn0_2),.clk(gclk));
	jdff dff_B_8N6yDly67_2(.din(w_dff_B_AKirHMAn0_2),.dout(w_dff_B_8N6yDly67_2),.clk(gclk));
	jdff dff_B_DvTfPtjn5_2(.din(w_dff_B_8N6yDly67_2),.dout(w_dff_B_DvTfPtjn5_2),.clk(gclk));
	jdff dff_B_sQNQuede2_2(.din(w_dff_B_DvTfPtjn5_2),.dout(w_dff_B_sQNQuede2_2),.clk(gclk));
	jdff dff_B_Xpc4Xt2r4_2(.din(w_dff_B_sQNQuede2_2),.dout(w_dff_B_Xpc4Xt2r4_2),.clk(gclk));
	jdff dff_B_9sAn7Fcb6_2(.din(n1621),.dout(w_dff_B_9sAn7Fcb6_2),.clk(gclk));
	jdff dff_B_hFlYIM527_2(.din(w_dff_B_9sAn7Fcb6_2),.dout(w_dff_B_hFlYIM527_2),.clk(gclk));
	jdff dff_B_lsNPF1TA8_2(.din(w_dff_B_hFlYIM527_2),.dout(w_dff_B_lsNPF1TA8_2),.clk(gclk));
	jdff dff_B_j0qBV0LY6_2(.din(w_dff_B_lsNPF1TA8_2),.dout(w_dff_B_j0qBV0LY6_2),.clk(gclk));
	jdff dff_B_gCtvqu4I2_2(.din(w_dff_B_j0qBV0LY6_2),.dout(w_dff_B_gCtvqu4I2_2),.clk(gclk));
	jdff dff_B_RidqMonS5_2(.din(w_dff_B_gCtvqu4I2_2),.dout(w_dff_B_RidqMonS5_2),.clk(gclk));
	jdff dff_B_nYS2B4yV8_2(.din(w_dff_B_RidqMonS5_2),.dout(w_dff_B_nYS2B4yV8_2),.clk(gclk));
	jdff dff_B_mchIiVzc1_2(.din(w_dff_B_nYS2B4yV8_2),.dout(w_dff_B_mchIiVzc1_2),.clk(gclk));
	jdff dff_B_sNEh0Q967_2(.din(w_dff_B_mchIiVzc1_2),.dout(w_dff_B_sNEh0Q967_2),.clk(gclk));
	jdff dff_B_VCfgkNlf1_2(.din(w_dff_B_sNEh0Q967_2),.dout(w_dff_B_VCfgkNlf1_2),.clk(gclk));
	jdff dff_B_k1xKFdHo2_2(.din(w_dff_B_VCfgkNlf1_2),.dout(w_dff_B_k1xKFdHo2_2),.clk(gclk));
	jdff dff_B_mQq6qvaZ3_2(.din(w_dff_B_k1xKFdHo2_2),.dout(w_dff_B_mQq6qvaZ3_2),.clk(gclk));
	jdff dff_B_KYdAZ0ES2_2(.din(w_dff_B_mQq6qvaZ3_2),.dout(w_dff_B_KYdAZ0ES2_2),.clk(gclk));
	jdff dff_B_C8c0Fvhr1_2(.din(w_dff_B_KYdAZ0ES2_2),.dout(w_dff_B_C8c0Fvhr1_2),.clk(gclk));
	jdff dff_B_SSKgi54W2_2(.din(w_dff_B_C8c0Fvhr1_2),.dout(w_dff_B_SSKgi54W2_2),.clk(gclk));
	jdff dff_B_j8oz2q7E1_2(.din(w_dff_B_SSKgi54W2_2),.dout(w_dff_B_j8oz2q7E1_2),.clk(gclk));
	jdff dff_B_7tgUzNhT3_2(.din(w_dff_B_j8oz2q7E1_2),.dout(w_dff_B_7tgUzNhT3_2),.clk(gclk));
	jdff dff_B_kTTGrVnz1_2(.din(w_dff_B_7tgUzNhT3_2),.dout(w_dff_B_kTTGrVnz1_2),.clk(gclk));
	jdff dff_B_frKsoiuy9_2(.din(w_dff_B_kTTGrVnz1_2),.dout(w_dff_B_frKsoiuy9_2),.clk(gclk));
	jdff dff_B_hfd3emXe7_2(.din(w_dff_B_frKsoiuy9_2),.dout(w_dff_B_hfd3emXe7_2),.clk(gclk));
	jdff dff_B_jccaAOYS8_2(.din(w_dff_B_hfd3emXe7_2),.dout(w_dff_B_jccaAOYS8_2),.clk(gclk));
	jdff dff_B_rkUXDS3V5_2(.din(w_dff_B_jccaAOYS8_2),.dout(w_dff_B_rkUXDS3V5_2),.clk(gclk));
	jdff dff_B_wSPNl7ez7_2(.din(w_dff_B_rkUXDS3V5_2),.dout(w_dff_B_wSPNl7ez7_2),.clk(gclk));
	jdff dff_B_P0WkqwtZ3_2(.din(w_dff_B_wSPNl7ez7_2),.dout(w_dff_B_P0WkqwtZ3_2),.clk(gclk));
	jdff dff_B_Zk9YvXF85_2(.din(w_dff_B_P0WkqwtZ3_2),.dout(w_dff_B_Zk9YvXF85_2),.clk(gclk));
	jdff dff_B_G1TmgyV26_2(.din(w_dff_B_Zk9YvXF85_2),.dout(w_dff_B_G1TmgyV26_2),.clk(gclk));
	jdff dff_B_IeFKOpvN1_2(.din(w_dff_B_G1TmgyV26_2),.dout(w_dff_B_IeFKOpvN1_2),.clk(gclk));
	jdff dff_B_IigCEz2c6_2(.din(w_dff_B_IeFKOpvN1_2),.dout(w_dff_B_IigCEz2c6_2),.clk(gclk));
	jdff dff_B_L8vOQTb50_2(.din(w_dff_B_IigCEz2c6_2),.dout(w_dff_B_L8vOQTb50_2),.clk(gclk));
	jdff dff_B_bd73EToM2_2(.din(w_dff_B_L8vOQTb50_2),.dout(w_dff_B_bd73EToM2_2),.clk(gclk));
	jdff dff_B_oWdZxOkF7_2(.din(w_dff_B_bd73EToM2_2),.dout(w_dff_B_oWdZxOkF7_2),.clk(gclk));
	jdff dff_B_wMxHba9J7_2(.din(w_dff_B_oWdZxOkF7_2),.dout(w_dff_B_wMxHba9J7_2),.clk(gclk));
	jdff dff_B_PCX08hoM6_2(.din(w_dff_B_wMxHba9J7_2),.dout(w_dff_B_PCX08hoM6_2),.clk(gclk));
	jdff dff_B_3Ec1X0q09_2(.din(w_dff_B_PCX08hoM6_2),.dout(w_dff_B_3Ec1X0q09_2),.clk(gclk));
	jdff dff_B_fUIKiS5m0_2(.din(w_dff_B_3Ec1X0q09_2),.dout(w_dff_B_fUIKiS5m0_2),.clk(gclk));
	jdff dff_B_RXKSSsqR2_2(.din(n1620),.dout(w_dff_B_RXKSSsqR2_2),.clk(gclk));
	jdff dff_B_lVfrHDpd8_1(.din(n1618),.dout(w_dff_B_lVfrHDpd8_1),.clk(gclk));
	jdff dff_B_Tbwpf6xt9_2(.din(n1560),.dout(w_dff_B_Tbwpf6xt9_2),.clk(gclk));
	jdff dff_B_4p6H30yu9_2(.din(w_dff_B_Tbwpf6xt9_2),.dout(w_dff_B_4p6H30yu9_2),.clk(gclk));
	jdff dff_B_NCV5bwJ41_2(.din(w_dff_B_4p6H30yu9_2),.dout(w_dff_B_NCV5bwJ41_2),.clk(gclk));
	jdff dff_B_K5lzGnLK5_2(.din(w_dff_B_NCV5bwJ41_2),.dout(w_dff_B_K5lzGnLK5_2),.clk(gclk));
	jdff dff_B_bx0cJ6n45_2(.din(w_dff_B_K5lzGnLK5_2),.dout(w_dff_B_bx0cJ6n45_2),.clk(gclk));
	jdff dff_B_YIAzdPWe5_2(.din(w_dff_B_bx0cJ6n45_2),.dout(w_dff_B_YIAzdPWe5_2),.clk(gclk));
	jdff dff_B_nfE1RCyW4_2(.din(w_dff_B_YIAzdPWe5_2),.dout(w_dff_B_nfE1RCyW4_2),.clk(gclk));
	jdff dff_B_mRxCSs2z4_2(.din(w_dff_B_nfE1RCyW4_2),.dout(w_dff_B_mRxCSs2z4_2),.clk(gclk));
	jdff dff_B_XE5Bi9jw8_2(.din(w_dff_B_mRxCSs2z4_2),.dout(w_dff_B_XE5Bi9jw8_2),.clk(gclk));
	jdff dff_B_jUhfG1Wo0_2(.din(w_dff_B_XE5Bi9jw8_2),.dout(w_dff_B_jUhfG1Wo0_2),.clk(gclk));
	jdff dff_B_a345NiQz9_2(.din(w_dff_B_jUhfG1Wo0_2),.dout(w_dff_B_a345NiQz9_2),.clk(gclk));
	jdff dff_B_axaNYMEY7_2(.din(w_dff_B_a345NiQz9_2),.dout(w_dff_B_axaNYMEY7_2),.clk(gclk));
	jdff dff_B_VGkCPCOe3_2(.din(w_dff_B_axaNYMEY7_2),.dout(w_dff_B_VGkCPCOe3_2),.clk(gclk));
	jdff dff_B_v6XLbMiq2_2(.din(w_dff_B_VGkCPCOe3_2),.dout(w_dff_B_v6XLbMiq2_2),.clk(gclk));
	jdff dff_B_oZ5UZ9j75_2(.din(w_dff_B_v6XLbMiq2_2),.dout(w_dff_B_oZ5UZ9j75_2),.clk(gclk));
	jdff dff_B_tvbVsxWb7_2(.din(w_dff_B_oZ5UZ9j75_2),.dout(w_dff_B_tvbVsxWb7_2),.clk(gclk));
	jdff dff_B_HYtGl2de5_2(.din(w_dff_B_tvbVsxWb7_2),.dout(w_dff_B_HYtGl2de5_2),.clk(gclk));
	jdff dff_B_oJ8eMsRB8_2(.din(w_dff_B_HYtGl2de5_2),.dout(w_dff_B_oJ8eMsRB8_2),.clk(gclk));
	jdff dff_B_xNXjctV55_2(.din(w_dff_B_oJ8eMsRB8_2),.dout(w_dff_B_xNXjctV55_2),.clk(gclk));
	jdff dff_B_yn6Jz8C52_2(.din(w_dff_B_xNXjctV55_2),.dout(w_dff_B_yn6Jz8C52_2),.clk(gclk));
	jdff dff_B_gjSxjEzl5_2(.din(w_dff_B_yn6Jz8C52_2),.dout(w_dff_B_gjSxjEzl5_2),.clk(gclk));
	jdff dff_B_tpO9zrKX3_2(.din(w_dff_B_gjSxjEzl5_2),.dout(w_dff_B_tpO9zrKX3_2),.clk(gclk));
	jdff dff_B_7o4EZgzI3_2(.din(w_dff_B_tpO9zrKX3_2),.dout(w_dff_B_7o4EZgzI3_2),.clk(gclk));
	jdff dff_B_pBitbiE92_2(.din(w_dff_B_7o4EZgzI3_2),.dout(w_dff_B_pBitbiE92_2),.clk(gclk));
	jdff dff_B_7th584bH8_2(.din(w_dff_B_pBitbiE92_2),.dout(w_dff_B_7th584bH8_2),.clk(gclk));
	jdff dff_B_IL1auyot5_2(.din(w_dff_B_7th584bH8_2),.dout(w_dff_B_IL1auyot5_2),.clk(gclk));
	jdff dff_B_Kvf7tkbt7_2(.din(w_dff_B_IL1auyot5_2),.dout(w_dff_B_Kvf7tkbt7_2),.clk(gclk));
	jdff dff_B_ul3IkykT6_2(.din(w_dff_B_Kvf7tkbt7_2),.dout(w_dff_B_ul3IkykT6_2),.clk(gclk));
	jdff dff_B_8jLUi6t41_2(.din(w_dff_B_ul3IkykT6_2),.dout(w_dff_B_8jLUi6t41_2),.clk(gclk));
	jdff dff_B_Q8QnPVam5_2(.din(w_dff_B_8jLUi6t41_2),.dout(w_dff_B_Q8QnPVam5_2),.clk(gclk));
	jdff dff_B_dGEwiIKs9_2(.din(w_dff_B_Q8QnPVam5_2),.dout(w_dff_B_dGEwiIKs9_2),.clk(gclk));
	jdff dff_B_NCLO9bGl6_2(.din(w_dff_B_dGEwiIKs9_2),.dout(w_dff_B_NCLO9bGl6_2),.clk(gclk));
	jdff dff_B_JqBDnx6C6_1(.din(n1566),.dout(w_dff_B_JqBDnx6C6_1),.clk(gclk));
	jdff dff_B_akoQDKb85_1(.din(w_dff_B_JqBDnx6C6_1),.dout(w_dff_B_akoQDKb85_1),.clk(gclk));
	jdff dff_B_80egostb8_2(.din(n1565),.dout(w_dff_B_80egostb8_2),.clk(gclk));
	jdff dff_B_gcHEIEyP4_2(.din(w_dff_B_80egostb8_2),.dout(w_dff_B_gcHEIEyP4_2),.clk(gclk));
	jdff dff_B_Knq085FN6_2(.din(w_dff_B_gcHEIEyP4_2),.dout(w_dff_B_Knq085FN6_2),.clk(gclk));
	jdff dff_B_xVBIBO344_2(.din(w_dff_B_Knq085FN6_2),.dout(w_dff_B_xVBIBO344_2),.clk(gclk));
	jdff dff_B_9fHuaslc8_2(.din(w_dff_B_xVBIBO344_2),.dout(w_dff_B_9fHuaslc8_2),.clk(gclk));
	jdff dff_B_mnsJi2EB1_2(.din(w_dff_B_9fHuaslc8_2),.dout(w_dff_B_mnsJi2EB1_2),.clk(gclk));
	jdff dff_B_SMHASyAu4_2(.din(w_dff_B_mnsJi2EB1_2),.dout(w_dff_B_SMHASyAu4_2),.clk(gclk));
	jdff dff_B_7IqK6qEg9_2(.din(w_dff_B_SMHASyAu4_2),.dout(w_dff_B_7IqK6qEg9_2),.clk(gclk));
	jdff dff_B_G8JdxIRP1_2(.din(w_dff_B_7IqK6qEg9_2),.dout(w_dff_B_G8JdxIRP1_2),.clk(gclk));
	jdff dff_B_R4DsbbLR1_2(.din(w_dff_B_G8JdxIRP1_2),.dout(w_dff_B_R4DsbbLR1_2),.clk(gclk));
	jdff dff_B_P472hPn29_2(.din(w_dff_B_R4DsbbLR1_2),.dout(w_dff_B_P472hPn29_2),.clk(gclk));
	jdff dff_B_lIDlEYAf0_2(.din(w_dff_B_P472hPn29_2),.dout(w_dff_B_lIDlEYAf0_2),.clk(gclk));
	jdff dff_B_dzRvG1Lu5_2(.din(w_dff_B_lIDlEYAf0_2),.dout(w_dff_B_dzRvG1Lu5_2),.clk(gclk));
	jdff dff_B_9EzyEBcd5_2(.din(w_dff_B_dzRvG1Lu5_2),.dout(w_dff_B_9EzyEBcd5_2),.clk(gclk));
	jdff dff_B_FD3a6GpS4_2(.din(w_dff_B_9EzyEBcd5_2),.dout(w_dff_B_FD3a6GpS4_2),.clk(gclk));
	jdff dff_B_CtD1V4Bz7_2(.din(w_dff_B_FD3a6GpS4_2),.dout(w_dff_B_CtD1V4Bz7_2),.clk(gclk));
	jdff dff_B_aIZ82vB52_2(.din(w_dff_B_CtD1V4Bz7_2),.dout(w_dff_B_aIZ82vB52_2),.clk(gclk));
	jdff dff_B_JQSAppdZ4_2(.din(w_dff_B_aIZ82vB52_2),.dout(w_dff_B_JQSAppdZ4_2),.clk(gclk));
	jdff dff_B_zKhtu69H4_2(.din(w_dff_B_JQSAppdZ4_2),.dout(w_dff_B_zKhtu69H4_2),.clk(gclk));
	jdff dff_B_buyjAk7I1_2(.din(w_dff_B_zKhtu69H4_2),.dout(w_dff_B_buyjAk7I1_2),.clk(gclk));
	jdff dff_B_Bb1KFwxw0_2(.din(w_dff_B_buyjAk7I1_2),.dout(w_dff_B_Bb1KFwxw0_2),.clk(gclk));
	jdff dff_B_geQLz2po7_2(.din(w_dff_B_Bb1KFwxw0_2),.dout(w_dff_B_geQLz2po7_2),.clk(gclk));
	jdff dff_B_hU03qZzE1_2(.din(w_dff_B_geQLz2po7_2),.dout(w_dff_B_hU03qZzE1_2),.clk(gclk));
	jdff dff_B_O0DEJEvc6_2(.din(w_dff_B_hU03qZzE1_2),.dout(w_dff_B_O0DEJEvc6_2),.clk(gclk));
	jdff dff_B_eQ3Uy3G08_2(.din(w_dff_B_O0DEJEvc6_2),.dout(w_dff_B_eQ3Uy3G08_2),.clk(gclk));
	jdff dff_B_yh7kAaU98_2(.din(w_dff_B_eQ3Uy3G08_2),.dout(w_dff_B_yh7kAaU98_2),.clk(gclk));
	jdff dff_B_h74D9eKU0_2(.din(w_dff_B_yh7kAaU98_2),.dout(w_dff_B_h74D9eKU0_2),.clk(gclk));
	jdff dff_B_f6waqcye3_2(.din(w_dff_B_h74D9eKU0_2),.dout(w_dff_B_f6waqcye3_2),.clk(gclk));
	jdff dff_B_q34FxeZk2_2(.din(w_dff_B_f6waqcye3_2),.dout(w_dff_B_q34FxeZk2_2),.clk(gclk));
	jdff dff_B_Bf9YOSqe2_2(.din(n1564),.dout(w_dff_B_Bf9YOSqe2_2),.clk(gclk));
	jdff dff_B_7nlPZ1h67_2(.din(w_dff_B_Bf9YOSqe2_2),.dout(w_dff_B_7nlPZ1h67_2),.clk(gclk));
	jdff dff_B_XTMmf55n7_2(.din(w_dff_B_7nlPZ1h67_2),.dout(w_dff_B_XTMmf55n7_2),.clk(gclk));
	jdff dff_B_0wG04RyC6_2(.din(w_dff_B_XTMmf55n7_2),.dout(w_dff_B_0wG04RyC6_2),.clk(gclk));
	jdff dff_B_lsRLi1j21_2(.din(w_dff_B_0wG04RyC6_2),.dout(w_dff_B_lsRLi1j21_2),.clk(gclk));
	jdff dff_B_6ZCo8SuC1_2(.din(w_dff_B_lsRLi1j21_2),.dout(w_dff_B_6ZCo8SuC1_2),.clk(gclk));
	jdff dff_B_g0yROJRG7_2(.din(w_dff_B_6ZCo8SuC1_2),.dout(w_dff_B_g0yROJRG7_2),.clk(gclk));
	jdff dff_B_KvTcEe1y7_2(.din(w_dff_B_g0yROJRG7_2),.dout(w_dff_B_KvTcEe1y7_2),.clk(gclk));
	jdff dff_B_V56bjvL51_2(.din(w_dff_B_KvTcEe1y7_2),.dout(w_dff_B_V56bjvL51_2),.clk(gclk));
	jdff dff_B_O3GCq6kZ7_2(.din(w_dff_B_V56bjvL51_2),.dout(w_dff_B_O3GCq6kZ7_2),.clk(gclk));
	jdff dff_B_ihzPeJjK7_2(.din(w_dff_B_O3GCq6kZ7_2),.dout(w_dff_B_ihzPeJjK7_2),.clk(gclk));
	jdff dff_B_mYM5gCoF7_2(.din(w_dff_B_ihzPeJjK7_2),.dout(w_dff_B_mYM5gCoF7_2),.clk(gclk));
	jdff dff_B_1yDYon1F2_2(.din(w_dff_B_mYM5gCoF7_2),.dout(w_dff_B_1yDYon1F2_2),.clk(gclk));
	jdff dff_B_k8xZ3v2D6_2(.din(w_dff_B_1yDYon1F2_2),.dout(w_dff_B_k8xZ3v2D6_2),.clk(gclk));
	jdff dff_B_UDeZe4N71_2(.din(w_dff_B_k8xZ3v2D6_2),.dout(w_dff_B_UDeZe4N71_2),.clk(gclk));
	jdff dff_B_wQN9B2v33_2(.din(w_dff_B_UDeZe4N71_2),.dout(w_dff_B_wQN9B2v33_2),.clk(gclk));
	jdff dff_B_IgagyY0E8_2(.din(w_dff_B_wQN9B2v33_2),.dout(w_dff_B_IgagyY0E8_2),.clk(gclk));
	jdff dff_B_HrTCHcvK7_2(.din(w_dff_B_IgagyY0E8_2),.dout(w_dff_B_HrTCHcvK7_2),.clk(gclk));
	jdff dff_B_JEOpD9dL1_2(.din(w_dff_B_HrTCHcvK7_2),.dout(w_dff_B_JEOpD9dL1_2),.clk(gclk));
	jdff dff_B_wXmlrgGV1_2(.din(w_dff_B_JEOpD9dL1_2),.dout(w_dff_B_wXmlrgGV1_2),.clk(gclk));
	jdff dff_B_WvqBDI8O0_2(.din(w_dff_B_wXmlrgGV1_2),.dout(w_dff_B_WvqBDI8O0_2),.clk(gclk));
	jdff dff_B_vzhlZg3w8_2(.din(w_dff_B_WvqBDI8O0_2),.dout(w_dff_B_vzhlZg3w8_2),.clk(gclk));
	jdff dff_B_NRMato3z0_2(.din(w_dff_B_vzhlZg3w8_2),.dout(w_dff_B_NRMato3z0_2),.clk(gclk));
	jdff dff_B_ns0dDKnN3_2(.din(w_dff_B_NRMato3z0_2),.dout(w_dff_B_ns0dDKnN3_2),.clk(gclk));
	jdff dff_B_eLhoSjZo1_2(.din(w_dff_B_ns0dDKnN3_2),.dout(w_dff_B_eLhoSjZo1_2),.clk(gclk));
	jdff dff_B_nnGcM5Q27_2(.din(w_dff_B_eLhoSjZo1_2),.dout(w_dff_B_nnGcM5Q27_2),.clk(gclk));
	jdff dff_B_bbUPCRWi9_2(.din(w_dff_B_nnGcM5Q27_2),.dout(w_dff_B_bbUPCRWi9_2),.clk(gclk));
	jdff dff_B_CbRoJI7X7_2(.din(w_dff_B_bbUPCRWi9_2),.dout(w_dff_B_CbRoJI7X7_2),.clk(gclk));
	jdff dff_B_5o1gj5FO1_2(.din(w_dff_B_CbRoJI7X7_2),.dout(w_dff_B_5o1gj5FO1_2),.clk(gclk));
	jdff dff_B_3xWtFiSr9_2(.din(w_dff_B_5o1gj5FO1_2),.dout(w_dff_B_3xWtFiSr9_2),.clk(gclk));
	jdff dff_B_AtA3bWf96_2(.din(w_dff_B_3xWtFiSr9_2),.dout(w_dff_B_AtA3bWf96_2),.clk(gclk));
	jdff dff_B_Lc401koj9_2(.din(n1563),.dout(w_dff_B_Lc401koj9_2),.clk(gclk));
	jdff dff_B_yLu2oWlL0_1(.din(n1561),.dout(w_dff_B_yLu2oWlL0_1),.clk(gclk));
	jdff dff_B_BKTdhDnF2_2(.din(n1496),.dout(w_dff_B_BKTdhDnF2_2),.clk(gclk));
	jdff dff_B_LzXR7G6t2_2(.din(w_dff_B_BKTdhDnF2_2),.dout(w_dff_B_LzXR7G6t2_2),.clk(gclk));
	jdff dff_B_0YeTcVzn2_2(.din(w_dff_B_LzXR7G6t2_2),.dout(w_dff_B_0YeTcVzn2_2),.clk(gclk));
	jdff dff_B_E5IgPBqR5_2(.din(w_dff_B_0YeTcVzn2_2),.dout(w_dff_B_E5IgPBqR5_2),.clk(gclk));
	jdff dff_B_Mn1sDoBt9_2(.din(w_dff_B_E5IgPBqR5_2),.dout(w_dff_B_Mn1sDoBt9_2),.clk(gclk));
	jdff dff_B_NiGSt4u23_2(.din(w_dff_B_Mn1sDoBt9_2),.dout(w_dff_B_NiGSt4u23_2),.clk(gclk));
	jdff dff_B_tLyMQgIP1_2(.din(w_dff_B_NiGSt4u23_2),.dout(w_dff_B_tLyMQgIP1_2),.clk(gclk));
	jdff dff_B_s48nmVZq0_2(.din(w_dff_B_tLyMQgIP1_2),.dout(w_dff_B_s48nmVZq0_2),.clk(gclk));
	jdff dff_B_eC59fv107_2(.din(w_dff_B_s48nmVZq0_2),.dout(w_dff_B_eC59fv107_2),.clk(gclk));
	jdff dff_B_zE3yWCua2_2(.din(w_dff_B_eC59fv107_2),.dout(w_dff_B_zE3yWCua2_2),.clk(gclk));
	jdff dff_B_dVd6AblZ6_2(.din(w_dff_B_zE3yWCua2_2),.dout(w_dff_B_dVd6AblZ6_2),.clk(gclk));
	jdff dff_B_B8bFEOKm6_2(.din(w_dff_B_dVd6AblZ6_2),.dout(w_dff_B_B8bFEOKm6_2),.clk(gclk));
	jdff dff_B_CGsZb66e7_2(.din(w_dff_B_B8bFEOKm6_2),.dout(w_dff_B_CGsZb66e7_2),.clk(gclk));
	jdff dff_B_WPMMIjTt1_2(.din(w_dff_B_CGsZb66e7_2),.dout(w_dff_B_WPMMIjTt1_2),.clk(gclk));
	jdff dff_B_FsH3WjZB3_2(.din(w_dff_B_WPMMIjTt1_2),.dout(w_dff_B_FsH3WjZB3_2),.clk(gclk));
	jdff dff_B_ibr7ghrX1_2(.din(w_dff_B_FsH3WjZB3_2),.dout(w_dff_B_ibr7ghrX1_2),.clk(gclk));
	jdff dff_B_PnAfyQpd1_2(.din(w_dff_B_ibr7ghrX1_2),.dout(w_dff_B_PnAfyQpd1_2),.clk(gclk));
	jdff dff_B_rUVhrAsh8_2(.din(w_dff_B_PnAfyQpd1_2),.dout(w_dff_B_rUVhrAsh8_2),.clk(gclk));
	jdff dff_B_zUVLmAQs5_2(.din(w_dff_B_rUVhrAsh8_2),.dout(w_dff_B_zUVLmAQs5_2),.clk(gclk));
	jdff dff_B_Ka83XLPu8_2(.din(w_dff_B_zUVLmAQs5_2),.dout(w_dff_B_Ka83XLPu8_2),.clk(gclk));
	jdff dff_B_nqQDGSgw0_2(.din(w_dff_B_Ka83XLPu8_2),.dout(w_dff_B_nqQDGSgw0_2),.clk(gclk));
	jdff dff_B_6Hq6EAjJ8_2(.din(w_dff_B_nqQDGSgw0_2),.dout(w_dff_B_6Hq6EAjJ8_2),.clk(gclk));
	jdff dff_B_fMHUahLR0_2(.din(w_dff_B_6Hq6EAjJ8_2),.dout(w_dff_B_fMHUahLR0_2),.clk(gclk));
	jdff dff_B_Gzq7vYFc0_2(.din(w_dff_B_fMHUahLR0_2),.dout(w_dff_B_Gzq7vYFc0_2),.clk(gclk));
	jdff dff_B_eLFM84gq6_2(.din(w_dff_B_Gzq7vYFc0_2),.dout(w_dff_B_eLFM84gq6_2),.clk(gclk));
	jdff dff_B_37kdYW5B6_2(.din(w_dff_B_eLFM84gq6_2),.dout(w_dff_B_37kdYW5B6_2),.clk(gclk));
	jdff dff_B_ivKCltzi8_2(.din(w_dff_B_37kdYW5B6_2),.dout(w_dff_B_ivKCltzi8_2),.clk(gclk));
	jdff dff_B_xOdbxLaE6_2(.din(w_dff_B_ivKCltzi8_2),.dout(w_dff_B_xOdbxLaE6_2),.clk(gclk));
	jdff dff_B_pHyen3Vw5_1(.din(n1502),.dout(w_dff_B_pHyen3Vw5_1),.clk(gclk));
	jdff dff_B_O4pQZRa68_1(.din(w_dff_B_pHyen3Vw5_1),.dout(w_dff_B_O4pQZRa68_1),.clk(gclk));
	jdff dff_B_VfOPYxpv2_2(.din(n1501),.dout(w_dff_B_VfOPYxpv2_2),.clk(gclk));
	jdff dff_B_sjij758H7_2(.din(w_dff_B_VfOPYxpv2_2),.dout(w_dff_B_sjij758H7_2),.clk(gclk));
	jdff dff_B_Yr8CD6EF9_2(.din(w_dff_B_sjij758H7_2),.dout(w_dff_B_Yr8CD6EF9_2),.clk(gclk));
	jdff dff_B_hdpzD2fa8_2(.din(w_dff_B_Yr8CD6EF9_2),.dout(w_dff_B_hdpzD2fa8_2),.clk(gclk));
	jdff dff_B_WJPSR8797_2(.din(w_dff_B_hdpzD2fa8_2),.dout(w_dff_B_WJPSR8797_2),.clk(gclk));
	jdff dff_B_Nbpw8GSc4_2(.din(w_dff_B_WJPSR8797_2),.dout(w_dff_B_Nbpw8GSc4_2),.clk(gclk));
	jdff dff_B_ddQWk0ub5_2(.din(w_dff_B_Nbpw8GSc4_2),.dout(w_dff_B_ddQWk0ub5_2),.clk(gclk));
	jdff dff_B_SGmKyeeq2_2(.din(w_dff_B_ddQWk0ub5_2),.dout(w_dff_B_SGmKyeeq2_2),.clk(gclk));
	jdff dff_B_eAeMZbFl5_2(.din(w_dff_B_SGmKyeeq2_2),.dout(w_dff_B_eAeMZbFl5_2),.clk(gclk));
	jdff dff_B_ClXnvXk25_2(.din(w_dff_B_eAeMZbFl5_2),.dout(w_dff_B_ClXnvXk25_2),.clk(gclk));
	jdff dff_B_CbyZSHUz2_2(.din(w_dff_B_ClXnvXk25_2),.dout(w_dff_B_CbyZSHUz2_2),.clk(gclk));
	jdff dff_B_tsmT14vq1_2(.din(w_dff_B_CbyZSHUz2_2),.dout(w_dff_B_tsmT14vq1_2),.clk(gclk));
	jdff dff_B_crN3jRC43_2(.din(w_dff_B_tsmT14vq1_2),.dout(w_dff_B_crN3jRC43_2),.clk(gclk));
	jdff dff_B_48Iods5x4_2(.din(w_dff_B_crN3jRC43_2),.dout(w_dff_B_48Iods5x4_2),.clk(gclk));
	jdff dff_B_VQxXYS8l8_2(.din(w_dff_B_48Iods5x4_2),.dout(w_dff_B_VQxXYS8l8_2),.clk(gclk));
	jdff dff_B_RSIiPJIW6_2(.din(w_dff_B_VQxXYS8l8_2),.dout(w_dff_B_RSIiPJIW6_2),.clk(gclk));
	jdff dff_B_ow2pnKit8_2(.din(w_dff_B_RSIiPJIW6_2),.dout(w_dff_B_ow2pnKit8_2),.clk(gclk));
	jdff dff_B_oyZ706BL6_2(.din(w_dff_B_ow2pnKit8_2),.dout(w_dff_B_oyZ706BL6_2),.clk(gclk));
	jdff dff_B_E5yecxaX6_2(.din(w_dff_B_oyZ706BL6_2),.dout(w_dff_B_E5yecxaX6_2),.clk(gclk));
	jdff dff_B_TpjybKn51_2(.din(w_dff_B_E5yecxaX6_2),.dout(w_dff_B_TpjybKn51_2),.clk(gclk));
	jdff dff_B_3zbxahj84_2(.din(w_dff_B_TpjybKn51_2),.dout(w_dff_B_3zbxahj84_2),.clk(gclk));
	jdff dff_B_1CDqRsBU4_2(.din(w_dff_B_3zbxahj84_2),.dout(w_dff_B_1CDqRsBU4_2),.clk(gclk));
	jdff dff_B_iz3mqyXT3_2(.din(w_dff_B_1CDqRsBU4_2),.dout(w_dff_B_iz3mqyXT3_2),.clk(gclk));
	jdff dff_B_Q3bdpMSd8_2(.din(w_dff_B_iz3mqyXT3_2),.dout(w_dff_B_Q3bdpMSd8_2),.clk(gclk));
	jdff dff_B_YQMQaZxU4_2(.din(w_dff_B_Q3bdpMSd8_2),.dout(w_dff_B_YQMQaZxU4_2),.clk(gclk));
	jdff dff_B_2Gvn7DMy9_2(.din(n1500),.dout(w_dff_B_2Gvn7DMy9_2),.clk(gclk));
	jdff dff_B_cbBRVvAf0_2(.din(w_dff_B_2Gvn7DMy9_2),.dout(w_dff_B_cbBRVvAf0_2),.clk(gclk));
	jdff dff_B_AS76nUfd4_2(.din(w_dff_B_cbBRVvAf0_2),.dout(w_dff_B_AS76nUfd4_2),.clk(gclk));
	jdff dff_B_DFaZJEyd8_2(.din(w_dff_B_AS76nUfd4_2),.dout(w_dff_B_DFaZJEyd8_2),.clk(gclk));
	jdff dff_B_J24kzodN2_2(.din(w_dff_B_DFaZJEyd8_2),.dout(w_dff_B_J24kzodN2_2),.clk(gclk));
	jdff dff_B_zwzp4V0h1_2(.din(w_dff_B_J24kzodN2_2),.dout(w_dff_B_zwzp4V0h1_2),.clk(gclk));
	jdff dff_B_5qoBdjaB4_2(.din(w_dff_B_zwzp4V0h1_2),.dout(w_dff_B_5qoBdjaB4_2),.clk(gclk));
	jdff dff_B_cKip2Vh62_2(.din(w_dff_B_5qoBdjaB4_2),.dout(w_dff_B_cKip2Vh62_2),.clk(gclk));
	jdff dff_B_PwhUEkCO8_2(.din(w_dff_B_cKip2Vh62_2),.dout(w_dff_B_PwhUEkCO8_2),.clk(gclk));
	jdff dff_B_8Os835gu0_2(.din(w_dff_B_PwhUEkCO8_2),.dout(w_dff_B_8Os835gu0_2),.clk(gclk));
	jdff dff_B_qtYUzJo82_2(.din(w_dff_B_8Os835gu0_2),.dout(w_dff_B_qtYUzJo82_2),.clk(gclk));
	jdff dff_B_MkqOsuV71_2(.din(w_dff_B_qtYUzJo82_2),.dout(w_dff_B_MkqOsuV71_2),.clk(gclk));
	jdff dff_B_4lpmtRRx0_2(.din(w_dff_B_MkqOsuV71_2),.dout(w_dff_B_4lpmtRRx0_2),.clk(gclk));
	jdff dff_B_0TZ1s0dd0_2(.din(w_dff_B_4lpmtRRx0_2),.dout(w_dff_B_0TZ1s0dd0_2),.clk(gclk));
	jdff dff_B_Mu6pU7tz2_2(.din(w_dff_B_0TZ1s0dd0_2),.dout(w_dff_B_Mu6pU7tz2_2),.clk(gclk));
	jdff dff_B_D8GY4yPm3_2(.din(w_dff_B_Mu6pU7tz2_2),.dout(w_dff_B_D8GY4yPm3_2),.clk(gclk));
	jdff dff_B_l4ulICik2_2(.din(w_dff_B_D8GY4yPm3_2),.dout(w_dff_B_l4ulICik2_2),.clk(gclk));
	jdff dff_B_yNtCmOZx2_2(.din(w_dff_B_l4ulICik2_2),.dout(w_dff_B_yNtCmOZx2_2),.clk(gclk));
	jdff dff_B_hHLtnYpG6_2(.din(w_dff_B_yNtCmOZx2_2),.dout(w_dff_B_hHLtnYpG6_2),.clk(gclk));
	jdff dff_B_CVVMM4nl2_2(.din(w_dff_B_hHLtnYpG6_2),.dout(w_dff_B_CVVMM4nl2_2),.clk(gclk));
	jdff dff_B_iN4KO8l51_2(.din(w_dff_B_CVVMM4nl2_2),.dout(w_dff_B_iN4KO8l51_2),.clk(gclk));
	jdff dff_B_nv21DhVX8_2(.din(w_dff_B_iN4KO8l51_2),.dout(w_dff_B_nv21DhVX8_2),.clk(gclk));
	jdff dff_B_hMGg3jI35_2(.din(w_dff_B_nv21DhVX8_2),.dout(w_dff_B_hMGg3jI35_2),.clk(gclk));
	jdff dff_B_Gvxw6GEQ6_2(.din(w_dff_B_hMGg3jI35_2),.dout(w_dff_B_Gvxw6GEQ6_2),.clk(gclk));
	jdff dff_B_ObiDmNgP1_2(.din(w_dff_B_Gvxw6GEQ6_2),.dout(w_dff_B_ObiDmNgP1_2),.clk(gclk));
	jdff dff_B_kiGupozr8_2(.din(w_dff_B_ObiDmNgP1_2),.dout(w_dff_B_kiGupozr8_2),.clk(gclk));
	jdff dff_B_sF8K7eJt7_2(.din(w_dff_B_kiGupozr8_2),.dout(w_dff_B_sF8K7eJt7_2),.clk(gclk));
	jdff dff_B_63ITM0IV8_2(.din(n1499),.dout(w_dff_B_63ITM0IV8_2),.clk(gclk));
	jdff dff_B_Nxts0IYw7_1(.din(n1497),.dout(w_dff_B_Nxts0IYw7_1),.clk(gclk));
	jdff dff_B_OqXGtk0r7_2(.din(n1425),.dout(w_dff_B_OqXGtk0r7_2),.clk(gclk));
	jdff dff_B_Cvja5RD80_2(.din(w_dff_B_OqXGtk0r7_2),.dout(w_dff_B_Cvja5RD80_2),.clk(gclk));
	jdff dff_B_NY42Quuc6_2(.din(w_dff_B_Cvja5RD80_2),.dout(w_dff_B_NY42Quuc6_2),.clk(gclk));
	jdff dff_B_M7SOeoaH5_2(.din(w_dff_B_NY42Quuc6_2),.dout(w_dff_B_M7SOeoaH5_2),.clk(gclk));
	jdff dff_B_jpgXIRCc1_2(.din(w_dff_B_M7SOeoaH5_2),.dout(w_dff_B_jpgXIRCc1_2),.clk(gclk));
	jdff dff_B_tNWJ3hDc2_2(.din(w_dff_B_jpgXIRCc1_2),.dout(w_dff_B_tNWJ3hDc2_2),.clk(gclk));
	jdff dff_B_eivDyMDw4_2(.din(w_dff_B_tNWJ3hDc2_2),.dout(w_dff_B_eivDyMDw4_2),.clk(gclk));
	jdff dff_B_jFIeS7iS5_2(.din(w_dff_B_eivDyMDw4_2),.dout(w_dff_B_jFIeS7iS5_2),.clk(gclk));
	jdff dff_B_tE7sWGt58_2(.din(w_dff_B_jFIeS7iS5_2),.dout(w_dff_B_tE7sWGt58_2),.clk(gclk));
	jdff dff_B_Blo8dg376_2(.din(w_dff_B_tE7sWGt58_2),.dout(w_dff_B_Blo8dg376_2),.clk(gclk));
	jdff dff_B_ZAa6HCIe9_2(.din(w_dff_B_Blo8dg376_2),.dout(w_dff_B_ZAa6HCIe9_2),.clk(gclk));
	jdff dff_B_eGeEOhDo8_2(.din(w_dff_B_ZAa6HCIe9_2),.dout(w_dff_B_eGeEOhDo8_2),.clk(gclk));
	jdff dff_B_c3LSE7Jp7_2(.din(w_dff_B_eGeEOhDo8_2),.dout(w_dff_B_c3LSE7Jp7_2),.clk(gclk));
	jdff dff_B_7y4iZ9Np2_2(.din(w_dff_B_c3LSE7Jp7_2),.dout(w_dff_B_7y4iZ9Np2_2),.clk(gclk));
	jdff dff_B_2F2XMy2d5_2(.din(w_dff_B_7y4iZ9Np2_2),.dout(w_dff_B_2F2XMy2d5_2),.clk(gclk));
	jdff dff_B_368IqZiA5_2(.din(w_dff_B_2F2XMy2d5_2),.dout(w_dff_B_368IqZiA5_2),.clk(gclk));
	jdff dff_B_SB2h7UB99_2(.din(w_dff_B_368IqZiA5_2),.dout(w_dff_B_SB2h7UB99_2),.clk(gclk));
	jdff dff_B_cWwLyUxA9_2(.din(w_dff_B_SB2h7UB99_2),.dout(w_dff_B_cWwLyUxA9_2),.clk(gclk));
	jdff dff_B_AvTLrOPv5_2(.din(w_dff_B_cWwLyUxA9_2),.dout(w_dff_B_AvTLrOPv5_2),.clk(gclk));
	jdff dff_B_ZUAe7bqy3_2(.din(w_dff_B_AvTLrOPv5_2),.dout(w_dff_B_ZUAe7bqy3_2),.clk(gclk));
	jdff dff_B_HOAfO1VV0_2(.din(w_dff_B_ZUAe7bqy3_2),.dout(w_dff_B_HOAfO1VV0_2),.clk(gclk));
	jdff dff_B_0hpV2Lgu2_2(.din(w_dff_B_HOAfO1VV0_2),.dout(w_dff_B_0hpV2Lgu2_2),.clk(gclk));
	jdff dff_B_iDM6MtEK6_2(.din(w_dff_B_0hpV2Lgu2_2),.dout(w_dff_B_iDM6MtEK6_2),.clk(gclk));
	jdff dff_B_cW7nfghM3_2(.din(w_dff_B_iDM6MtEK6_2),.dout(w_dff_B_cW7nfghM3_2),.clk(gclk));
	jdff dff_B_PSOlWlRS9_1(.din(n1431),.dout(w_dff_B_PSOlWlRS9_1),.clk(gclk));
	jdff dff_B_kUPrBYtM2_1(.din(w_dff_B_PSOlWlRS9_1),.dout(w_dff_B_kUPrBYtM2_1),.clk(gclk));
	jdff dff_B_nYbFUOK69_2(.din(n1430),.dout(w_dff_B_nYbFUOK69_2),.clk(gclk));
	jdff dff_B_ArXbxpJ25_2(.din(w_dff_B_nYbFUOK69_2),.dout(w_dff_B_ArXbxpJ25_2),.clk(gclk));
	jdff dff_B_KTvJJh0v9_2(.din(w_dff_B_ArXbxpJ25_2),.dout(w_dff_B_KTvJJh0v9_2),.clk(gclk));
	jdff dff_B_MarX1VX68_2(.din(w_dff_B_KTvJJh0v9_2),.dout(w_dff_B_MarX1VX68_2),.clk(gclk));
	jdff dff_B_8RpZfeWw6_2(.din(w_dff_B_MarX1VX68_2),.dout(w_dff_B_8RpZfeWw6_2),.clk(gclk));
	jdff dff_B_F31DFCFA2_2(.din(w_dff_B_8RpZfeWw6_2),.dout(w_dff_B_F31DFCFA2_2),.clk(gclk));
	jdff dff_B_w9m4zXIC9_2(.din(w_dff_B_F31DFCFA2_2),.dout(w_dff_B_w9m4zXIC9_2),.clk(gclk));
	jdff dff_B_wDvJF5NS0_2(.din(w_dff_B_w9m4zXIC9_2),.dout(w_dff_B_wDvJF5NS0_2),.clk(gclk));
	jdff dff_B_BBLwHwkQ8_2(.din(w_dff_B_wDvJF5NS0_2),.dout(w_dff_B_BBLwHwkQ8_2),.clk(gclk));
	jdff dff_B_UuwrVsM92_2(.din(w_dff_B_BBLwHwkQ8_2),.dout(w_dff_B_UuwrVsM92_2),.clk(gclk));
	jdff dff_B_EpoIowCu8_2(.din(w_dff_B_UuwrVsM92_2),.dout(w_dff_B_EpoIowCu8_2),.clk(gclk));
	jdff dff_B_ia5N8OXy8_2(.din(w_dff_B_EpoIowCu8_2),.dout(w_dff_B_ia5N8OXy8_2),.clk(gclk));
	jdff dff_B_Pn8Pv91D0_2(.din(w_dff_B_ia5N8OXy8_2),.dout(w_dff_B_Pn8Pv91D0_2),.clk(gclk));
	jdff dff_B_svcJVEXU4_2(.din(w_dff_B_Pn8Pv91D0_2),.dout(w_dff_B_svcJVEXU4_2),.clk(gclk));
	jdff dff_B_bdYi72WB1_2(.din(w_dff_B_svcJVEXU4_2),.dout(w_dff_B_bdYi72WB1_2),.clk(gclk));
	jdff dff_B_3TUxJHuE5_2(.din(w_dff_B_bdYi72WB1_2),.dout(w_dff_B_3TUxJHuE5_2),.clk(gclk));
	jdff dff_B_2eJcINEF6_2(.din(w_dff_B_3TUxJHuE5_2),.dout(w_dff_B_2eJcINEF6_2),.clk(gclk));
	jdff dff_B_uV5GGtDX8_2(.din(w_dff_B_2eJcINEF6_2),.dout(w_dff_B_uV5GGtDX8_2),.clk(gclk));
	jdff dff_B_vUkUamBW4_2(.din(w_dff_B_uV5GGtDX8_2),.dout(w_dff_B_vUkUamBW4_2),.clk(gclk));
	jdff dff_B_nDOtVjXs8_2(.din(w_dff_B_vUkUamBW4_2),.dout(w_dff_B_nDOtVjXs8_2),.clk(gclk));
	jdff dff_B_y2SyWNyp8_2(.din(w_dff_B_nDOtVjXs8_2),.dout(w_dff_B_y2SyWNyp8_2),.clk(gclk));
	jdff dff_B_OAWrp7nW6_2(.din(n1429),.dout(w_dff_B_OAWrp7nW6_2),.clk(gclk));
	jdff dff_B_cc8BGGwY9_2(.din(w_dff_B_OAWrp7nW6_2),.dout(w_dff_B_cc8BGGwY9_2),.clk(gclk));
	jdff dff_B_Gx5uZHb87_2(.din(w_dff_B_cc8BGGwY9_2),.dout(w_dff_B_Gx5uZHb87_2),.clk(gclk));
	jdff dff_B_XDhq4FBF6_2(.din(w_dff_B_Gx5uZHb87_2),.dout(w_dff_B_XDhq4FBF6_2),.clk(gclk));
	jdff dff_B_OfWoQqJH2_2(.din(w_dff_B_XDhq4FBF6_2),.dout(w_dff_B_OfWoQqJH2_2),.clk(gclk));
	jdff dff_B_BR4Tjjvr4_2(.din(w_dff_B_OfWoQqJH2_2),.dout(w_dff_B_BR4Tjjvr4_2),.clk(gclk));
	jdff dff_B_ZaHkSOZg9_2(.din(w_dff_B_BR4Tjjvr4_2),.dout(w_dff_B_ZaHkSOZg9_2),.clk(gclk));
	jdff dff_B_w5vKRf4Z8_2(.din(w_dff_B_ZaHkSOZg9_2),.dout(w_dff_B_w5vKRf4Z8_2),.clk(gclk));
	jdff dff_B_iKbfZKgF7_2(.din(w_dff_B_w5vKRf4Z8_2),.dout(w_dff_B_iKbfZKgF7_2),.clk(gclk));
	jdff dff_B_Q9IKnMa38_2(.din(w_dff_B_iKbfZKgF7_2),.dout(w_dff_B_Q9IKnMa38_2),.clk(gclk));
	jdff dff_B_CQX2jHmG3_2(.din(w_dff_B_Q9IKnMa38_2),.dout(w_dff_B_CQX2jHmG3_2),.clk(gclk));
	jdff dff_B_f63iPIcQ4_2(.din(w_dff_B_CQX2jHmG3_2),.dout(w_dff_B_f63iPIcQ4_2),.clk(gclk));
	jdff dff_B_38x8kn8X4_2(.din(w_dff_B_f63iPIcQ4_2),.dout(w_dff_B_38x8kn8X4_2),.clk(gclk));
	jdff dff_B_C0vKHX3G1_2(.din(w_dff_B_38x8kn8X4_2),.dout(w_dff_B_C0vKHX3G1_2),.clk(gclk));
	jdff dff_B_hIz0nFUS3_2(.din(w_dff_B_C0vKHX3G1_2),.dout(w_dff_B_hIz0nFUS3_2),.clk(gclk));
	jdff dff_B_geBw50nT9_2(.din(w_dff_B_hIz0nFUS3_2),.dout(w_dff_B_geBw50nT9_2),.clk(gclk));
	jdff dff_B_lKA6DX5k0_2(.din(w_dff_B_geBw50nT9_2),.dout(w_dff_B_lKA6DX5k0_2),.clk(gclk));
	jdff dff_B_YsxI9lXF3_2(.din(w_dff_B_lKA6DX5k0_2),.dout(w_dff_B_YsxI9lXF3_2),.clk(gclk));
	jdff dff_B_vNTh4RgE6_2(.din(w_dff_B_YsxI9lXF3_2),.dout(w_dff_B_vNTh4RgE6_2),.clk(gclk));
	jdff dff_B_kEIsEVAr4_2(.din(w_dff_B_vNTh4RgE6_2),.dout(w_dff_B_kEIsEVAr4_2),.clk(gclk));
	jdff dff_B_8wSfaBW14_2(.din(w_dff_B_kEIsEVAr4_2),.dout(w_dff_B_8wSfaBW14_2),.clk(gclk));
	jdff dff_B_fNZgH5Ia3_2(.din(w_dff_B_8wSfaBW14_2),.dout(w_dff_B_fNZgH5Ia3_2),.clk(gclk));
	jdff dff_B_gF9ti5EF3_2(.din(w_dff_B_fNZgH5Ia3_2),.dout(w_dff_B_gF9ti5EF3_2),.clk(gclk));
	jdff dff_B_1XAPDj0M1_2(.din(n1428),.dout(w_dff_B_1XAPDj0M1_2),.clk(gclk));
	jdff dff_B_0bFHJie74_1(.din(n1426),.dout(w_dff_B_0bFHJie74_1),.clk(gclk));
	jdff dff_B_4UY19m043_2(.din(n1347),.dout(w_dff_B_4UY19m043_2),.clk(gclk));
	jdff dff_B_d9XBYaqX8_2(.din(w_dff_B_4UY19m043_2),.dout(w_dff_B_d9XBYaqX8_2),.clk(gclk));
	jdff dff_B_YVabvJQa1_2(.din(w_dff_B_d9XBYaqX8_2),.dout(w_dff_B_YVabvJQa1_2),.clk(gclk));
	jdff dff_B_eC30aI6f6_2(.din(w_dff_B_YVabvJQa1_2),.dout(w_dff_B_eC30aI6f6_2),.clk(gclk));
	jdff dff_B_CPXcp7ny7_2(.din(w_dff_B_eC30aI6f6_2),.dout(w_dff_B_CPXcp7ny7_2),.clk(gclk));
	jdff dff_B_6dNqTBbT2_2(.din(w_dff_B_CPXcp7ny7_2),.dout(w_dff_B_6dNqTBbT2_2),.clk(gclk));
	jdff dff_B_Q5O0HqW16_2(.din(w_dff_B_6dNqTBbT2_2),.dout(w_dff_B_Q5O0HqW16_2),.clk(gclk));
	jdff dff_B_efNjonfQ7_2(.din(w_dff_B_Q5O0HqW16_2),.dout(w_dff_B_efNjonfQ7_2),.clk(gclk));
	jdff dff_B_iDnnnMfs1_2(.din(w_dff_B_efNjonfQ7_2),.dout(w_dff_B_iDnnnMfs1_2),.clk(gclk));
	jdff dff_B_fYOrmObb1_2(.din(w_dff_B_iDnnnMfs1_2),.dout(w_dff_B_fYOrmObb1_2),.clk(gclk));
	jdff dff_B_jYhlo0RK9_2(.din(w_dff_B_fYOrmObb1_2),.dout(w_dff_B_jYhlo0RK9_2),.clk(gclk));
	jdff dff_B_o96tmtMv2_2(.din(w_dff_B_jYhlo0RK9_2),.dout(w_dff_B_o96tmtMv2_2),.clk(gclk));
	jdff dff_B_tggmTTTF3_2(.din(w_dff_B_o96tmtMv2_2),.dout(w_dff_B_tggmTTTF3_2),.clk(gclk));
	jdff dff_B_IbjrAGqq9_2(.din(w_dff_B_tggmTTTF3_2),.dout(w_dff_B_IbjrAGqq9_2),.clk(gclk));
	jdff dff_B_u5zh3mSe2_2(.din(w_dff_B_IbjrAGqq9_2),.dout(w_dff_B_u5zh3mSe2_2),.clk(gclk));
	jdff dff_B_MjBcxu072_2(.din(w_dff_B_u5zh3mSe2_2),.dout(w_dff_B_MjBcxu072_2),.clk(gclk));
	jdff dff_B_eUTUXKbM1_2(.din(w_dff_B_MjBcxu072_2),.dout(w_dff_B_eUTUXKbM1_2),.clk(gclk));
	jdff dff_B_Ffqu1yuv3_2(.din(w_dff_B_eUTUXKbM1_2),.dout(w_dff_B_Ffqu1yuv3_2),.clk(gclk));
	jdff dff_B_3qWJqvg82_2(.din(w_dff_B_Ffqu1yuv3_2),.dout(w_dff_B_3qWJqvg82_2),.clk(gclk));
	jdff dff_B_jfnFqI8W0_2(.din(w_dff_B_3qWJqvg82_2),.dout(w_dff_B_jfnFqI8W0_2),.clk(gclk));
	jdff dff_B_IUJTneI48_1(.din(n1353),.dout(w_dff_B_IUJTneI48_1),.clk(gclk));
	jdff dff_B_O9rLtxNu0_1(.din(w_dff_B_IUJTneI48_1),.dout(w_dff_B_O9rLtxNu0_1),.clk(gclk));
	jdff dff_B_Yo4NJgHU9_2(.din(n1352),.dout(w_dff_B_Yo4NJgHU9_2),.clk(gclk));
	jdff dff_B_nAYduoFH1_2(.din(w_dff_B_Yo4NJgHU9_2),.dout(w_dff_B_nAYduoFH1_2),.clk(gclk));
	jdff dff_B_uASePRO83_2(.din(w_dff_B_nAYduoFH1_2),.dout(w_dff_B_uASePRO83_2),.clk(gclk));
	jdff dff_B_4faQDMdp3_2(.din(w_dff_B_uASePRO83_2),.dout(w_dff_B_4faQDMdp3_2),.clk(gclk));
	jdff dff_B_CPE5SUUB5_2(.din(w_dff_B_4faQDMdp3_2),.dout(w_dff_B_CPE5SUUB5_2),.clk(gclk));
	jdff dff_B_IM3GGFyb2_2(.din(w_dff_B_CPE5SUUB5_2),.dout(w_dff_B_IM3GGFyb2_2),.clk(gclk));
	jdff dff_B_BbHgMiGc9_2(.din(w_dff_B_IM3GGFyb2_2),.dout(w_dff_B_BbHgMiGc9_2),.clk(gclk));
	jdff dff_B_uY2zE2uQ1_2(.din(w_dff_B_BbHgMiGc9_2),.dout(w_dff_B_uY2zE2uQ1_2),.clk(gclk));
	jdff dff_B_bCKBVgiw5_2(.din(w_dff_B_uY2zE2uQ1_2),.dout(w_dff_B_bCKBVgiw5_2),.clk(gclk));
	jdff dff_B_OUade5p45_2(.din(w_dff_B_bCKBVgiw5_2),.dout(w_dff_B_OUade5p45_2),.clk(gclk));
	jdff dff_B_urKKBo6M9_2(.din(w_dff_B_OUade5p45_2),.dout(w_dff_B_urKKBo6M9_2),.clk(gclk));
	jdff dff_B_4o4OIB594_2(.din(w_dff_B_urKKBo6M9_2),.dout(w_dff_B_4o4OIB594_2),.clk(gclk));
	jdff dff_B_6WX05CD52_2(.din(w_dff_B_4o4OIB594_2),.dout(w_dff_B_6WX05CD52_2),.clk(gclk));
	jdff dff_B_xw50NHlM0_2(.din(w_dff_B_6WX05CD52_2),.dout(w_dff_B_xw50NHlM0_2),.clk(gclk));
	jdff dff_B_dmkToIFs6_2(.din(w_dff_B_xw50NHlM0_2),.dout(w_dff_B_dmkToIFs6_2),.clk(gclk));
	jdff dff_B_7eMuuLbb2_2(.din(w_dff_B_dmkToIFs6_2),.dout(w_dff_B_7eMuuLbb2_2),.clk(gclk));
	jdff dff_B_id4ZkbFR2_2(.din(w_dff_B_7eMuuLbb2_2),.dout(w_dff_B_id4ZkbFR2_2),.clk(gclk));
	jdff dff_B_vnMnEEWT2_2(.din(n1351),.dout(w_dff_B_vnMnEEWT2_2),.clk(gclk));
	jdff dff_B_sbjTJYux0_2(.din(w_dff_B_vnMnEEWT2_2),.dout(w_dff_B_sbjTJYux0_2),.clk(gclk));
	jdff dff_B_BVFSdiRn2_2(.din(w_dff_B_sbjTJYux0_2),.dout(w_dff_B_BVFSdiRn2_2),.clk(gclk));
	jdff dff_B_O2Pq2xS98_2(.din(w_dff_B_BVFSdiRn2_2),.dout(w_dff_B_O2Pq2xS98_2),.clk(gclk));
	jdff dff_B_yWAG5Exw1_2(.din(w_dff_B_O2Pq2xS98_2),.dout(w_dff_B_yWAG5Exw1_2),.clk(gclk));
	jdff dff_B_7ON9MR2A7_2(.din(w_dff_B_yWAG5Exw1_2),.dout(w_dff_B_7ON9MR2A7_2),.clk(gclk));
	jdff dff_B_hRAbzofl0_2(.din(w_dff_B_7ON9MR2A7_2),.dout(w_dff_B_hRAbzofl0_2),.clk(gclk));
	jdff dff_B_vAjlP61A0_2(.din(w_dff_B_hRAbzofl0_2),.dout(w_dff_B_vAjlP61A0_2),.clk(gclk));
	jdff dff_B_GUiXVbHH3_2(.din(w_dff_B_vAjlP61A0_2),.dout(w_dff_B_GUiXVbHH3_2),.clk(gclk));
	jdff dff_B_2pkieY3j1_2(.din(w_dff_B_GUiXVbHH3_2),.dout(w_dff_B_2pkieY3j1_2),.clk(gclk));
	jdff dff_B_6MkznyUo3_2(.din(w_dff_B_2pkieY3j1_2),.dout(w_dff_B_6MkznyUo3_2),.clk(gclk));
	jdff dff_B_TJrw2N5p9_2(.din(w_dff_B_6MkznyUo3_2),.dout(w_dff_B_TJrw2N5p9_2),.clk(gclk));
	jdff dff_B_2kvg4Fv99_2(.din(w_dff_B_TJrw2N5p9_2),.dout(w_dff_B_2kvg4Fv99_2),.clk(gclk));
	jdff dff_B_nVoxdnes2_2(.din(w_dff_B_2kvg4Fv99_2),.dout(w_dff_B_nVoxdnes2_2),.clk(gclk));
	jdff dff_B_D5utOWhA6_2(.din(w_dff_B_nVoxdnes2_2),.dout(w_dff_B_D5utOWhA6_2),.clk(gclk));
	jdff dff_B_jF5xRy7D9_2(.din(w_dff_B_D5utOWhA6_2),.dout(w_dff_B_jF5xRy7D9_2),.clk(gclk));
	jdff dff_B_Kmmi47nv6_2(.din(w_dff_B_jF5xRy7D9_2),.dout(w_dff_B_Kmmi47nv6_2),.clk(gclk));
	jdff dff_B_LC3BOYRO6_2(.din(w_dff_B_Kmmi47nv6_2),.dout(w_dff_B_LC3BOYRO6_2),.clk(gclk));
	jdff dff_B_R1ismnub3_2(.din(w_dff_B_LC3BOYRO6_2),.dout(w_dff_B_R1ismnub3_2),.clk(gclk));
	jdff dff_B_3mVv4DRR9_1(.din(n1348),.dout(w_dff_B_3mVv4DRR9_1),.clk(gclk));
	jdff dff_B_IWHhk4Ln3_2(.din(n1262),.dout(w_dff_B_IWHhk4Ln3_2),.clk(gclk));
	jdff dff_B_leddj2aF4_2(.din(w_dff_B_IWHhk4Ln3_2),.dout(w_dff_B_leddj2aF4_2),.clk(gclk));
	jdff dff_B_8rkaynPQ6_2(.din(w_dff_B_leddj2aF4_2),.dout(w_dff_B_8rkaynPQ6_2),.clk(gclk));
	jdff dff_B_sijKPjN28_2(.din(w_dff_B_8rkaynPQ6_2),.dout(w_dff_B_sijKPjN28_2),.clk(gclk));
	jdff dff_B_K5YNOlXo8_2(.din(w_dff_B_sijKPjN28_2),.dout(w_dff_B_K5YNOlXo8_2),.clk(gclk));
	jdff dff_B_M3BiYllW4_2(.din(w_dff_B_K5YNOlXo8_2),.dout(w_dff_B_M3BiYllW4_2),.clk(gclk));
	jdff dff_B_QSITtQkT5_2(.din(w_dff_B_M3BiYllW4_2),.dout(w_dff_B_QSITtQkT5_2),.clk(gclk));
	jdff dff_B_R0G6dGWk8_2(.din(w_dff_B_QSITtQkT5_2),.dout(w_dff_B_R0G6dGWk8_2),.clk(gclk));
	jdff dff_B_378IHsSa2_2(.din(w_dff_B_R0G6dGWk8_2),.dout(w_dff_B_378IHsSa2_2),.clk(gclk));
	jdff dff_B_ZG6YCjww7_2(.din(w_dff_B_378IHsSa2_2),.dout(w_dff_B_ZG6YCjww7_2),.clk(gclk));
	jdff dff_B_tOv6AX2j9_2(.din(w_dff_B_ZG6YCjww7_2),.dout(w_dff_B_tOv6AX2j9_2),.clk(gclk));
	jdff dff_B_K0hzm4e26_2(.din(w_dff_B_tOv6AX2j9_2),.dout(w_dff_B_K0hzm4e26_2),.clk(gclk));
	jdff dff_B_I5UfBLWq2_2(.din(w_dff_B_K0hzm4e26_2),.dout(w_dff_B_I5UfBLWq2_2),.clk(gclk));
	jdff dff_B_m2EJuf2V9_2(.din(w_dff_B_I5UfBLWq2_2),.dout(w_dff_B_m2EJuf2V9_2),.clk(gclk));
	jdff dff_B_2gu2iADJ0_2(.din(w_dff_B_m2EJuf2V9_2),.dout(w_dff_B_2gu2iADJ0_2),.clk(gclk));
	jdff dff_B_elEvupHo3_2(.din(w_dff_B_2gu2iADJ0_2),.dout(w_dff_B_elEvupHo3_2),.clk(gclk));
	jdff dff_B_AteBDex17_2(.din(w_dff_B_elEvupHo3_2),.dout(w_dff_B_AteBDex17_2),.clk(gclk));
	jdff dff_B_PKQSLXiP0_2(.din(n1273),.dout(w_dff_B_PKQSLXiP0_2),.clk(gclk));
	jdff dff_B_z3lkp7JR6_1(.din(n1268),.dout(w_dff_B_z3lkp7JR6_1),.clk(gclk));
	jdff dff_B_CSsJu4ca9_1(.din(w_dff_B_z3lkp7JR6_1),.dout(w_dff_B_CSsJu4ca9_1),.clk(gclk));
	jdff dff_B_Xo2BpnRW5_2(.din(n1267),.dout(w_dff_B_Xo2BpnRW5_2),.clk(gclk));
	jdff dff_B_5XQ0nrF35_2(.din(w_dff_B_Xo2BpnRW5_2),.dout(w_dff_B_5XQ0nrF35_2),.clk(gclk));
	jdff dff_B_qEXWvxh97_2(.din(w_dff_B_5XQ0nrF35_2),.dout(w_dff_B_qEXWvxh97_2),.clk(gclk));
	jdff dff_B_ZQJPXZFV5_2(.din(w_dff_B_qEXWvxh97_2),.dout(w_dff_B_ZQJPXZFV5_2),.clk(gclk));
	jdff dff_B_5IxobdZq5_2(.din(w_dff_B_ZQJPXZFV5_2),.dout(w_dff_B_5IxobdZq5_2),.clk(gclk));
	jdff dff_B_Jcy3oZuD4_2(.din(w_dff_B_5IxobdZq5_2),.dout(w_dff_B_Jcy3oZuD4_2),.clk(gclk));
	jdff dff_B_sYLgovAu7_2(.din(w_dff_B_Jcy3oZuD4_2),.dout(w_dff_B_sYLgovAu7_2),.clk(gclk));
	jdff dff_B_IZ6bZz6v2_2(.din(w_dff_B_sYLgovAu7_2),.dout(w_dff_B_IZ6bZz6v2_2),.clk(gclk));
	jdff dff_B_zrOP94kH2_2(.din(w_dff_B_IZ6bZz6v2_2),.dout(w_dff_B_zrOP94kH2_2),.clk(gclk));
	jdff dff_B_zompo2d58_2(.din(w_dff_B_zrOP94kH2_2),.dout(w_dff_B_zompo2d58_2),.clk(gclk));
	jdff dff_B_7lUNFWuT8_2(.din(w_dff_B_zompo2d58_2),.dout(w_dff_B_7lUNFWuT8_2),.clk(gclk));
	jdff dff_B_usv94h986_2(.din(w_dff_B_7lUNFWuT8_2),.dout(w_dff_B_usv94h986_2),.clk(gclk));
	jdff dff_B_W5C7l31p9_2(.din(w_dff_B_usv94h986_2),.dout(w_dff_B_W5C7l31p9_2),.clk(gclk));
	jdff dff_B_qEfu1ZfZ0_2(.din(n1266),.dout(w_dff_B_qEfu1ZfZ0_2),.clk(gclk));
	jdff dff_B_ZkRmFNuL2_2(.din(w_dff_B_qEfu1ZfZ0_2),.dout(w_dff_B_ZkRmFNuL2_2),.clk(gclk));
	jdff dff_B_VeaPsWuT4_2(.din(w_dff_B_ZkRmFNuL2_2),.dout(w_dff_B_VeaPsWuT4_2),.clk(gclk));
	jdff dff_B_3lEBNQst8_2(.din(w_dff_B_VeaPsWuT4_2),.dout(w_dff_B_3lEBNQst8_2),.clk(gclk));
	jdff dff_B_wcFO4hM45_2(.din(w_dff_B_3lEBNQst8_2),.dout(w_dff_B_wcFO4hM45_2),.clk(gclk));
	jdff dff_B_WJpZxDEC1_2(.din(w_dff_B_wcFO4hM45_2),.dout(w_dff_B_WJpZxDEC1_2),.clk(gclk));
	jdff dff_B_E037uTcI2_2(.din(w_dff_B_WJpZxDEC1_2),.dout(w_dff_B_E037uTcI2_2),.clk(gclk));
	jdff dff_B_Jhkh5mMR1_2(.din(w_dff_B_E037uTcI2_2),.dout(w_dff_B_Jhkh5mMR1_2),.clk(gclk));
	jdff dff_B_UK9mqZU10_2(.din(w_dff_B_Jhkh5mMR1_2),.dout(w_dff_B_UK9mqZU10_2),.clk(gclk));
	jdff dff_B_avWyTI751_2(.din(w_dff_B_UK9mqZU10_2),.dout(w_dff_B_avWyTI751_2),.clk(gclk));
	jdff dff_B_GC9wIpFz2_2(.din(w_dff_B_avWyTI751_2),.dout(w_dff_B_GC9wIpFz2_2),.clk(gclk));
	jdff dff_B_EIgSh8By8_2(.din(w_dff_B_GC9wIpFz2_2),.dout(w_dff_B_EIgSh8By8_2),.clk(gclk));
	jdff dff_B_tysjgboV3_2(.din(w_dff_B_EIgSh8By8_2),.dout(w_dff_B_tysjgboV3_2),.clk(gclk));
	jdff dff_B_0d5u6kvY2_2(.din(w_dff_B_tysjgboV3_2),.dout(w_dff_B_0d5u6kvY2_2),.clk(gclk));
	jdff dff_B_E3ivLrTe7_2(.din(w_dff_B_0d5u6kvY2_2),.dout(w_dff_B_E3ivLrTe7_2),.clk(gclk));
	jdff dff_B_zd2kEF9W7_1(.din(n1263),.dout(w_dff_B_zd2kEF9W7_1),.clk(gclk));
	jdff dff_B_uDJOOt0d7_2(.din(n1171),.dout(w_dff_B_uDJOOt0d7_2),.clk(gclk));
	jdff dff_B_0nOHOJjq5_2(.din(w_dff_B_uDJOOt0d7_2),.dout(w_dff_B_0nOHOJjq5_2),.clk(gclk));
	jdff dff_B_IDCpIKvz6_2(.din(w_dff_B_0nOHOJjq5_2),.dout(w_dff_B_IDCpIKvz6_2),.clk(gclk));
	jdff dff_B_74qhtc2l4_2(.din(w_dff_B_IDCpIKvz6_2),.dout(w_dff_B_74qhtc2l4_2),.clk(gclk));
	jdff dff_B_lyUkxFj24_2(.din(w_dff_B_74qhtc2l4_2),.dout(w_dff_B_lyUkxFj24_2),.clk(gclk));
	jdff dff_B_ezwYcDka4_2(.din(w_dff_B_lyUkxFj24_2),.dout(w_dff_B_ezwYcDka4_2),.clk(gclk));
	jdff dff_B_ikgVUA8i4_2(.din(w_dff_B_ezwYcDka4_2),.dout(w_dff_B_ikgVUA8i4_2),.clk(gclk));
	jdff dff_B_D1X70OjW9_2(.din(w_dff_B_ikgVUA8i4_2),.dout(w_dff_B_D1X70OjW9_2),.clk(gclk));
	jdff dff_B_tVvhSEI03_2(.din(w_dff_B_D1X70OjW9_2),.dout(w_dff_B_tVvhSEI03_2),.clk(gclk));
	jdff dff_B_FaPaHFCc3_2(.din(w_dff_B_tVvhSEI03_2),.dout(w_dff_B_FaPaHFCc3_2),.clk(gclk));
	jdff dff_B_q11e93fA8_2(.din(w_dff_B_FaPaHFCc3_2),.dout(w_dff_B_q11e93fA8_2),.clk(gclk));
	jdff dff_B_CHQM5nyO9_2(.din(w_dff_B_q11e93fA8_2),.dout(w_dff_B_CHQM5nyO9_2),.clk(gclk));
	jdff dff_B_yAJlfnKR7_2(.din(w_dff_B_CHQM5nyO9_2),.dout(w_dff_B_yAJlfnKR7_2),.clk(gclk));
	jdff dff_B_7AgCoNZE4_2(.din(w_dff_B_yAJlfnKR7_2),.dout(w_dff_B_7AgCoNZE4_2),.clk(gclk));
	jdff dff_B_XS4WX4E57_2(.din(n1182),.dout(w_dff_B_XS4WX4E57_2),.clk(gclk));
	jdff dff_B_RkzEbBhT9_2(.din(w_dff_B_XS4WX4E57_2),.dout(w_dff_B_RkzEbBhT9_2),.clk(gclk));
	jdff dff_B_bIQlvcg20_1(.din(n1177),.dout(w_dff_B_bIQlvcg20_1),.clk(gclk));
	jdff dff_B_Gjt8d74j1_1(.din(w_dff_B_bIQlvcg20_1),.dout(w_dff_B_Gjt8d74j1_1),.clk(gclk));
	jdff dff_B_LXYLAeB95_2(.din(n1176),.dout(w_dff_B_LXYLAeB95_2),.clk(gclk));
	jdff dff_B_0n2a2h1X1_2(.din(w_dff_B_LXYLAeB95_2),.dout(w_dff_B_0n2a2h1X1_2),.clk(gclk));
	jdff dff_B_wFXnMAqk6_2(.din(w_dff_B_0n2a2h1X1_2),.dout(w_dff_B_wFXnMAqk6_2),.clk(gclk));
	jdff dff_B_CXqwzez22_2(.din(w_dff_B_wFXnMAqk6_2),.dout(w_dff_B_CXqwzez22_2),.clk(gclk));
	jdff dff_B_f59dO4s58_2(.din(w_dff_B_CXqwzez22_2),.dout(w_dff_B_f59dO4s58_2),.clk(gclk));
	jdff dff_B_AVFPRMmi6_2(.din(w_dff_B_f59dO4s58_2),.dout(w_dff_B_AVFPRMmi6_2),.clk(gclk));
	jdff dff_B_w8A3RxER3_2(.din(w_dff_B_AVFPRMmi6_2),.dout(w_dff_B_w8A3RxER3_2),.clk(gclk));
	jdff dff_B_l1bbskJE9_2(.din(w_dff_B_w8A3RxER3_2),.dout(w_dff_B_l1bbskJE9_2),.clk(gclk));
	jdff dff_B_Wjv0KT8C0_2(.din(w_dff_B_l1bbskJE9_2),.dout(w_dff_B_Wjv0KT8C0_2),.clk(gclk));
	jdff dff_B_WhlOOeS69_2(.din(n1175),.dout(w_dff_B_WhlOOeS69_2),.clk(gclk));
	jdff dff_B_IVbFDPnX4_2(.din(w_dff_B_WhlOOeS69_2),.dout(w_dff_B_IVbFDPnX4_2),.clk(gclk));
	jdff dff_B_bXLmwg2S1_2(.din(w_dff_B_IVbFDPnX4_2),.dout(w_dff_B_bXLmwg2S1_2),.clk(gclk));
	jdff dff_B_ERRyIOcK5_2(.din(w_dff_B_bXLmwg2S1_2),.dout(w_dff_B_ERRyIOcK5_2),.clk(gclk));
	jdff dff_B_7GO5bWIN1_2(.din(w_dff_B_ERRyIOcK5_2),.dout(w_dff_B_7GO5bWIN1_2),.clk(gclk));
	jdff dff_B_Lz2fwbes8_2(.din(w_dff_B_7GO5bWIN1_2),.dout(w_dff_B_Lz2fwbes8_2),.clk(gclk));
	jdff dff_B_ZCvR93kx6_2(.din(w_dff_B_Lz2fwbes8_2),.dout(w_dff_B_ZCvR93kx6_2),.clk(gclk));
	jdff dff_B_xz6pQ6NE1_2(.din(w_dff_B_ZCvR93kx6_2),.dout(w_dff_B_xz6pQ6NE1_2),.clk(gclk));
	jdff dff_B_bUScqbrk2_2(.din(w_dff_B_xz6pQ6NE1_2),.dout(w_dff_B_bUScqbrk2_2),.clk(gclk));
	jdff dff_B_4HW70j5j1_2(.din(w_dff_B_bUScqbrk2_2),.dout(w_dff_B_4HW70j5j1_2),.clk(gclk));
	jdff dff_B_WfUqXEjd0_2(.din(w_dff_B_4HW70j5j1_2),.dout(w_dff_B_WfUqXEjd0_2),.clk(gclk));
	jdff dff_B_Ufyikq8N9_1(.din(n1172),.dout(w_dff_B_Ufyikq8N9_1),.clk(gclk));
	jdff dff_B_UveMoWF14_2(.din(n1073),.dout(w_dff_B_UveMoWF14_2),.clk(gclk));
	jdff dff_B_ulyTI7Oq7_2(.din(w_dff_B_UveMoWF14_2),.dout(w_dff_B_ulyTI7Oq7_2),.clk(gclk));
	jdff dff_B_OnKaUG1J7_2(.din(w_dff_B_ulyTI7Oq7_2),.dout(w_dff_B_OnKaUG1J7_2),.clk(gclk));
	jdff dff_B_hNzvNxiS0_2(.din(w_dff_B_OnKaUG1J7_2),.dout(w_dff_B_hNzvNxiS0_2),.clk(gclk));
	jdff dff_B_3vonbvKI4_2(.din(w_dff_B_hNzvNxiS0_2),.dout(w_dff_B_3vonbvKI4_2),.clk(gclk));
	jdff dff_B_2PgK952V4_2(.din(w_dff_B_3vonbvKI4_2),.dout(w_dff_B_2PgK952V4_2),.clk(gclk));
	jdff dff_B_bF404Jso3_2(.din(w_dff_B_2PgK952V4_2),.dout(w_dff_B_bF404Jso3_2),.clk(gclk));
	jdff dff_B_9Lzn0eOn5_2(.din(w_dff_B_bF404Jso3_2),.dout(w_dff_B_9Lzn0eOn5_2),.clk(gclk));
	jdff dff_B_SsUnkEGl2_2(.din(w_dff_B_9Lzn0eOn5_2),.dout(w_dff_B_SsUnkEGl2_2),.clk(gclk));
	jdff dff_B_ScpWsRMN6_2(.din(w_dff_B_SsUnkEGl2_2),.dout(w_dff_B_ScpWsRMN6_2),.clk(gclk));
	jdff dff_B_REPYmE8F0_2(.din(w_dff_B_ScpWsRMN6_2),.dout(w_dff_B_REPYmE8F0_2),.clk(gclk));
	jdff dff_B_SuelSZ3s7_2(.din(n1083),.dout(w_dff_B_SuelSZ3s7_2),.clk(gclk));
	jdff dff_B_4160zYfZ2_2(.din(w_dff_B_SuelSZ3s7_2),.dout(w_dff_B_4160zYfZ2_2),.clk(gclk));
	jdff dff_B_VcfgjPsI0_2(.din(w_dff_B_4160zYfZ2_2),.dout(w_dff_B_VcfgjPsI0_2),.clk(gclk));
	jdff dff_B_GlaY8Bbk6_2(.din(n1078),.dout(w_dff_B_GlaY8Bbk6_2),.clk(gclk));
	jdff dff_B_T3ULk5nn6_2(.din(w_dff_B_GlaY8Bbk6_2),.dout(w_dff_B_T3ULk5nn6_2),.clk(gclk));
	jdff dff_B_mcsrWnJK6_2(.din(w_dff_B_T3ULk5nn6_2),.dout(w_dff_B_mcsrWnJK6_2),.clk(gclk));
	jdff dff_B_NbWDpy8r7_2(.din(w_dff_B_mcsrWnJK6_2),.dout(w_dff_B_NbWDpy8r7_2),.clk(gclk));
	jdff dff_B_XKFgzDIA2_2(.din(w_dff_B_NbWDpy8r7_2),.dout(w_dff_B_XKFgzDIA2_2),.clk(gclk));
	jdff dff_B_eBmO4flu4_2(.din(n1077),.dout(w_dff_B_eBmO4flu4_2),.clk(gclk));
	jdff dff_B_6YAPjww34_2(.din(w_dff_B_eBmO4flu4_2),.dout(w_dff_B_6YAPjww34_2),.clk(gclk));
	jdff dff_B_eadTlS2A1_2(.din(w_dff_B_6YAPjww34_2),.dout(w_dff_B_eadTlS2A1_2),.clk(gclk));
	jdff dff_B_H8eNOtfX5_2(.din(w_dff_B_eadTlS2A1_2),.dout(w_dff_B_H8eNOtfX5_2),.clk(gclk));
	jdff dff_B_TZmvMU6P3_2(.din(w_dff_B_H8eNOtfX5_2),.dout(w_dff_B_TZmvMU6P3_2),.clk(gclk));
	jdff dff_B_91W0zb4V7_2(.din(w_dff_B_TZmvMU6P3_2),.dout(w_dff_B_91W0zb4V7_2),.clk(gclk));
	jdff dff_B_WKGtY2ml4_2(.din(w_dff_B_91W0zb4V7_2),.dout(w_dff_B_WKGtY2ml4_2),.clk(gclk));
	jdff dff_B_vjml4cqS8_1(.din(n1074),.dout(w_dff_B_vjml4cqS8_1),.clk(gclk));
	jdff dff_B_KpVUuAJN5_2(.din(n974),.dout(w_dff_B_KpVUuAJN5_2),.clk(gclk));
	jdff dff_B_w9jauQoR8_2(.din(w_dff_B_KpVUuAJN5_2),.dout(w_dff_B_w9jauQoR8_2),.clk(gclk));
	jdff dff_B_EaHDlXP45_2(.din(w_dff_B_w9jauQoR8_2),.dout(w_dff_B_EaHDlXP45_2),.clk(gclk));
	jdff dff_B_m8IARHne9_2(.din(w_dff_B_EaHDlXP45_2),.dout(w_dff_B_m8IARHne9_2),.clk(gclk));
	jdff dff_B_SJ9DI1s79_2(.din(w_dff_B_m8IARHne9_2),.dout(w_dff_B_SJ9DI1s79_2),.clk(gclk));
	jdff dff_B_8CrwbxYA8_2(.din(w_dff_B_SJ9DI1s79_2),.dout(w_dff_B_8CrwbxYA8_2),.clk(gclk));
	jdff dff_B_Ttx1IJNK3_2(.din(w_dff_B_8CrwbxYA8_2),.dout(w_dff_B_Ttx1IJNK3_2),.clk(gclk));
	jdff dff_B_mRin9tCy3_2(.din(w_dff_B_Ttx1IJNK3_2),.dout(w_dff_B_mRin9tCy3_2),.clk(gclk));
	jdff dff_B_tDITpW1u6_2(.din(n984),.dout(w_dff_B_tDITpW1u6_2),.clk(gclk));
	jdff dff_B_3e9rjiZe8_2(.din(w_dff_B_tDITpW1u6_2),.dout(w_dff_B_3e9rjiZe8_2),.clk(gclk));
	jdff dff_B_cLrWZABO6_2(.din(w_dff_B_3e9rjiZe8_2),.dout(w_dff_B_cLrWZABO6_2),.clk(gclk));
	jdff dff_B_GaJSvwO06_2(.din(w_dff_B_cLrWZABO6_2),.dout(w_dff_B_GaJSvwO06_2),.clk(gclk));
	jdff dff_B_gMd2PrvX8_2(.din(n983),.dout(w_dff_B_gMd2PrvX8_2),.clk(gclk));
	jdff dff_B_kc3LZIYa9_2(.din(w_dff_B_gMd2PrvX8_2),.dout(w_dff_B_kc3LZIYa9_2),.clk(gclk));
	jdff dff_B_gOT3hRON5_2(.din(w_dff_B_kc3LZIYa9_2),.dout(w_dff_B_gOT3hRON5_2),.clk(gclk));
	jdff dff_A_mBmYYDfz3_0(.dout(w_n980_0[0]),.din(w_dff_A_mBmYYDfz3_0),.clk(gclk));
	jdff dff_A_9NCxbHb42_0(.dout(w_dff_A_mBmYYDfz3_0),.din(w_dff_A_9NCxbHb42_0),.clk(gclk));
	jdff dff_A_UX8pD6aF4_0(.dout(w_dff_A_9NCxbHb42_0),.din(w_dff_A_UX8pD6aF4_0),.clk(gclk));
	jdff dff_B_mbQs6htz1_2(.din(n980),.dout(w_dff_B_mbQs6htz1_2),.clk(gclk));
	jdff dff_A_Y79VpmHU5_0(.dout(w_n877_0[0]),.din(w_dff_A_Y79VpmHU5_0),.clk(gclk));
	jdff dff_A_7r8RQZfT3_0(.dout(w_dff_A_Y79VpmHU5_0),.din(w_dff_A_7r8RQZfT3_0),.clk(gclk));
	jdff dff_A_cs9E2wFq9_0(.dout(w_dff_A_7r8RQZfT3_0),.din(w_dff_A_cs9E2wFq9_0),.clk(gclk));
	jdff dff_B_2jQ3RK4d0_2(.din(n877),.dout(w_dff_B_2jQ3RK4d0_2),.clk(gclk));
	jdff dff_A_XBZdRkvs1_0(.dout(w_n875_0[0]),.din(w_dff_A_XBZdRkvs1_0),.clk(gclk));
	jdff dff_A_BkdLtBcM6_0(.dout(w_dff_A_XBZdRkvs1_0),.din(w_dff_A_BkdLtBcM6_0),.clk(gclk));
	jdff dff_B_lXjMKyo05_2(.din(n874),.dout(w_dff_B_lXjMKyo05_2),.clk(gclk));
	jdff dff_B_JasEiltx4_2(.din(w_dff_B_lXjMKyo05_2),.dout(w_dff_B_JasEiltx4_2),.clk(gclk));
	jdff dff_B_Q2iIP7Qg7_2(.din(w_dff_B_JasEiltx4_2),.dout(w_dff_B_Q2iIP7Qg7_2),.clk(gclk));
	jdff dff_A_ooBIzX3Q9_1(.dout(w_dff_A_ooalAoq50_0),.din(w_dff_A_ooBIzX3Q9_1),.clk(gclk));
	jdff dff_A_ooalAoq50_0(.dout(w_dff_A_DSr6ENMU4_0),.din(w_dff_A_ooalAoq50_0),.clk(gclk));
	jdff dff_A_DSr6ENMU4_0(.dout(w_dff_A_wNznkkHX1_0),.din(w_dff_A_DSr6ENMU4_0),.clk(gclk));
	jdff dff_A_wNznkkHX1_0(.dout(w_dff_A_FrQBhmAr8_0),.din(w_dff_A_wNznkkHX1_0),.clk(gclk));
	jdff dff_A_FrQBhmAr8_0(.dout(w_dff_A_Hhbenz899_0),.din(w_dff_A_FrQBhmAr8_0),.clk(gclk));
	jdff dff_A_Hhbenz899_0(.dout(w_dff_A_NxH2jbQk7_0),.din(w_dff_A_Hhbenz899_0),.clk(gclk));
	jdff dff_A_NxH2jbQk7_0(.dout(w_dff_A_TLX1PWnh2_0),.din(w_dff_A_NxH2jbQk7_0),.clk(gclk));
	jdff dff_A_TLX1PWnh2_0(.dout(w_dff_A_sN2TyrCa8_0),.din(w_dff_A_TLX1PWnh2_0),.clk(gclk));
	jdff dff_A_sN2TyrCa8_0(.dout(w_dff_A_K0FvvkJp9_0),.din(w_dff_A_sN2TyrCa8_0),.clk(gclk));
	jdff dff_A_K0FvvkJp9_0(.dout(w_dff_A_LifDZLrE0_0),.din(w_dff_A_K0FvvkJp9_0),.clk(gclk));
	jdff dff_A_LifDZLrE0_0(.dout(w_dff_A_N06ojCkr9_0),.din(w_dff_A_LifDZLrE0_0),.clk(gclk));
	jdff dff_A_N06ojCkr9_0(.dout(w_dff_A_PY0KxP1a2_0),.din(w_dff_A_N06ojCkr9_0),.clk(gclk));
	jdff dff_A_PY0KxP1a2_0(.dout(w_dff_A_wJFNUXW48_0),.din(w_dff_A_PY0KxP1a2_0),.clk(gclk));
	jdff dff_A_wJFNUXW48_0(.dout(w_dff_A_5iBuQOlB0_0),.din(w_dff_A_wJFNUXW48_0),.clk(gclk));
	jdff dff_A_5iBuQOlB0_0(.dout(w_dff_A_BlHXVJON3_0),.din(w_dff_A_5iBuQOlB0_0),.clk(gclk));
	jdff dff_A_BlHXVJON3_0(.dout(w_dff_A_cnCqwNHi6_0),.din(w_dff_A_BlHXVJON3_0),.clk(gclk));
	jdff dff_A_cnCqwNHi6_0(.dout(w_dff_A_GzQiZkhL6_0),.din(w_dff_A_cnCqwNHi6_0),.clk(gclk));
	jdff dff_A_GzQiZkhL6_0(.dout(w_dff_A_Wwvneifu8_0),.din(w_dff_A_GzQiZkhL6_0),.clk(gclk));
	jdff dff_A_Wwvneifu8_0(.dout(w_dff_A_KkzAZReB7_0),.din(w_dff_A_Wwvneifu8_0),.clk(gclk));
	jdff dff_A_KkzAZReB7_0(.dout(w_dff_A_p1jrxzGC0_0),.din(w_dff_A_KkzAZReB7_0),.clk(gclk));
	jdff dff_A_p1jrxzGC0_0(.dout(w_dff_A_qwlMhPvA7_0),.din(w_dff_A_p1jrxzGC0_0),.clk(gclk));
	jdff dff_A_qwlMhPvA7_0(.dout(w_dff_A_zhrHWjME2_0),.din(w_dff_A_qwlMhPvA7_0),.clk(gclk));
	jdff dff_A_zhrHWjME2_0(.dout(w_dff_A_KNVu0Ji99_0),.din(w_dff_A_zhrHWjME2_0),.clk(gclk));
	jdff dff_A_KNVu0Ji99_0(.dout(w_dff_A_JmNUEczm9_0),.din(w_dff_A_KNVu0Ji99_0),.clk(gclk));
	jdff dff_A_JmNUEczm9_0(.dout(w_dff_A_m0nE4OuU7_0),.din(w_dff_A_JmNUEczm9_0),.clk(gclk));
	jdff dff_A_m0nE4OuU7_0(.dout(w_dff_A_BxmNwcYk5_0),.din(w_dff_A_m0nE4OuU7_0),.clk(gclk));
	jdff dff_A_BxmNwcYk5_0(.dout(w_dff_A_3k6zDv6d1_0),.din(w_dff_A_BxmNwcYk5_0),.clk(gclk));
	jdff dff_A_3k6zDv6d1_0(.dout(w_dff_A_URc29qnp7_0),.din(w_dff_A_3k6zDv6d1_0),.clk(gclk));
	jdff dff_A_URc29qnp7_0(.dout(w_dff_A_3hSDRLeS9_0),.din(w_dff_A_URc29qnp7_0),.clk(gclk));
	jdff dff_A_3hSDRLeS9_0(.dout(w_dff_A_fV559tTN4_0),.din(w_dff_A_3hSDRLeS9_0),.clk(gclk));
	jdff dff_A_fV559tTN4_0(.dout(w_dff_A_471LQcjL6_0),.din(w_dff_A_fV559tTN4_0),.clk(gclk));
	jdff dff_A_471LQcjL6_0(.dout(w_dff_A_j16ILcqv7_0),.din(w_dff_A_471LQcjL6_0),.clk(gclk));
	jdff dff_A_j16ILcqv7_0(.dout(w_dff_A_xQF2nmdq4_0),.din(w_dff_A_j16ILcqv7_0),.clk(gclk));
	jdff dff_A_xQF2nmdq4_0(.dout(w_dff_A_9JTXxx1I4_0),.din(w_dff_A_xQF2nmdq4_0),.clk(gclk));
	jdff dff_A_9JTXxx1I4_0(.dout(w_dff_A_ZxzDFWJl7_0),.din(w_dff_A_9JTXxx1I4_0),.clk(gclk));
	jdff dff_A_ZxzDFWJl7_0(.dout(w_dff_A_ChmJP1dU7_0),.din(w_dff_A_ZxzDFWJl7_0),.clk(gclk));
	jdff dff_A_ChmJP1dU7_0(.dout(w_dff_A_Xr4LdzK80_0),.din(w_dff_A_ChmJP1dU7_0),.clk(gclk));
	jdff dff_A_Xr4LdzK80_0(.dout(w_dff_A_JccgSi2u0_0),.din(w_dff_A_Xr4LdzK80_0),.clk(gclk));
	jdff dff_A_JccgSi2u0_0(.dout(w_dff_A_8OcIxksp1_0),.din(w_dff_A_JccgSi2u0_0),.clk(gclk));
	jdff dff_A_8OcIxksp1_0(.dout(w_dff_A_QuCUHEMZ8_0),.din(w_dff_A_8OcIxksp1_0),.clk(gclk));
	jdff dff_A_QuCUHEMZ8_0(.dout(w_dff_A_fdOsw1VI3_0),.din(w_dff_A_QuCUHEMZ8_0),.clk(gclk));
	jdff dff_A_fdOsw1VI3_0(.dout(w_dff_A_SdXJdlXV0_0),.din(w_dff_A_fdOsw1VI3_0),.clk(gclk));
	jdff dff_A_SdXJdlXV0_0(.dout(w_dff_A_cb5J6VfX0_0),.din(w_dff_A_SdXJdlXV0_0),.clk(gclk));
	jdff dff_A_cb5J6VfX0_0(.dout(w_dff_A_oDRamxAK6_0),.din(w_dff_A_cb5J6VfX0_0),.clk(gclk));
	jdff dff_A_oDRamxAK6_0(.dout(w_dff_A_HxYkZiuK6_0),.din(w_dff_A_oDRamxAK6_0),.clk(gclk));
	jdff dff_A_HxYkZiuK6_0(.dout(w_dff_A_eeamE3s85_0),.din(w_dff_A_HxYkZiuK6_0),.clk(gclk));
	jdff dff_A_eeamE3s85_0(.dout(w_dff_A_rVm0TM4c4_0),.din(w_dff_A_eeamE3s85_0),.clk(gclk));
	jdff dff_A_rVm0TM4c4_0(.dout(w_dff_A_XY5LdrhZ4_0),.din(w_dff_A_rVm0TM4c4_0),.clk(gclk));
	jdff dff_A_XY5LdrhZ4_0(.dout(w_dff_A_dTmWJk0V3_0),.din(w_dff_A_XY5LdrhZ4_0),.clk(gclk));
	jdff dff_A_dTmWJk0V3_0(.dout(w_dff_A_tbuDP5oc9_0),.din(w_dff_A_dTmWJk0V3_0),.clk(gclk));
	jdff dff_A_tbuDP5oc9_0(.dout(w_dff_A_pFkx1aAh1_0),.din(w_dff_A_tbuDP5oc9_0),.clk(gclk));
	jdff dff_A_pFkx1aAh1_0(.dout(w_dff_A_rYeUySUg9_0),.din(w_dff_A_pFkx1aAh1_0),.clk(gclk));
	jdff dff_A_rYeUySUg9_0(.dout(w_dff_A_YfJtFXKK6_0),.din(w_dff_A_rYeUySUg9_0),.clk(gclk));
	jdff dff_A_YfJtFXKK6_0(.dout(w_dff_A_7EWBmJsn3_0),.din(w_dff_A_YfJtFXKK6_0),.clk(gclk));
	jdff dff_A_7EWBmJsn3_0(.dout(w_dff_A_hRb4Uy4R2_0),.din(w_dff_A_7EWBmJsn3_0),.clk(gclk));
	jdff dff_A_hRb4Uy4R2_0(.dout(w_dff_A_1MBESbvS7_0),.din(w_dff_A_hRb4Uy4R2_0),.clk(gclk));
	jdff dff_A_1MBESbvS7_0(.dout(w_dff_A_4iKiaaya0_0),.din(w_dff_A_1MBESbvS7_0),.clk(gclk));
	jdff dff_A_4iKiaaya0_0(.dout(w_dff_A_tPAHFVZ62_0),.din(w_dff_A_4iKiaaya0_0),.clk(gclk));
	jdff dff_A_tPAHFVZ62_0(.dout(w_dff_A_fyTdke9w0_0),.din(w_dff_A_tPAHFVZ62_0),.clk(gclk));
	jdff dff_A_fyTdke9w0_0(.dout(w_dff_A_sPx8JKZc8_0),.din(w_dff_A_fyTdke9w0_0),.clk(gclk));
	jdff dff_A_sPx8JKZc8_0(.dout(w_dff_A_BefKe4R87_0),.din(w_dff_A_sPx8JKZc8_0),.clk(gclk));
	jdff dff_A_BefKe4R87_0(.dout(w_dff_A_F2E10s9i9_0),.din(w_dff_A_BefKe4R87_0),.clk(gclk));
	jdff dff_A_F2E10s9i9_0(.dout(w_dff_A_gXzTkQsB0_0),.din(w_dff_A_F2E10s9i9_0),.clk(gclk));
	jdff dff_A_gXzTkQsB0_0(.dout(w_dff_A_KV3yWYH62_0),.din(w_dff_A_gXzTkQsB0_0),.clk(gclk));
	jdff dff_A_KV3yWYH62_0(.dout(w_dff_A_b4sTED5r7_0),.din(w_dff_A_KV3yWYH62_0),.clk(gclk));
	jdff dff_A_b4sTED5r7_0(.dout(w_dff_A_kEVgXev02_0),.din(w_dff_A_b4sTED5r7_0),.clk(gclk));
	jdff dff_A_kEVgXev02_0(.dout(w_dff_A_wOJOhcwG3_0),.din(w_dff_A_kEVgXev02_0),.clk(gclk));
	jdff dff_A_wOJOhcwG3_0(.dout(w_dff_A_twS3z4Md7_0),.din(w_dff_A_wOJOhcwG3_0),.clk(gclk));
	jdff dff_A_twS3z4Md7_0(.dout(w_dff_A_c6JWTf9y6_0),.din(w_dff_A_twS3z4Md7_0),.clk(gclk));
	jdff dff_A_c6JWTf9y6_0(.dout(w_dff_A_BEn3V9Gl9_0),.din(w_dff_A_c6JWTf9y6_0),.clk(gclk));
	jdff dff_A_BEn3V9Gl9_0(.dout(w_dff_A_YYHzYWnv7_0),.din(w_dff_A_BEn3V9Gl9_0),.clk(gclk));
	jdff dff_A_YYHzYWnv7_0(.dout(w_dff_A_xsrUDg8Q4_0),.din(w_dff_A_YYHzYWnv7_0),.clk(gclk));
	jdff dff_A_xsrUDg8Q4_0(.dout(w_dff_A_d5AloKRx0_0),.din(w_dff_A_xsrUDg8Q4_0),.clk(gclk));
	jdff dff_A_d5AloKRx0_0(.dout(G545gat),.din(w_dff_A_d5AloKRx0_0),.clk(gclk));
	jdff dff_A_ERwqQcch6_2(.dout(w_dff_A_n9GB75JS3_0),.din(w_dff_A_ERwqQcch6_2),.clk(gclk));
	jdff dff_A_n9GB75JS3_0(.dout(w_dff_A_hHvtGTlQ8_0),.din(w_dff_A_n9GB75JS3_0),.clk(gclk));
	jdff dff_A_hHvtGTlQ8_0(.dout(w_dff_A_AnFkQSy58_0),.din(w_dff_A_hHvtGTlQ8_0),.clk(gclk));
	jdff dff_A_AnFkQSy58_0(.dout(w_dff_A_alQvqies3_0),.din(w_dff_A_AnFkQSy58_0),.clk(gclk));
	jdff dff_A_alQvqies3_0(.dout(w_dff_A_NTsj793Y3_0),.din(w_dff_A_alQvqies3_0),.clk(gclk));
	jdff dff_A_NTsj793Y3_0(.dout(w_dff_A_UdfStCmJ6_0),.din(w_dff_A_NTsj793Y3_0),.clk(gclk));
	jdff dff_A_UdfStCmJ6_0(.dout(w_dff_A_M5Gc7Mn44_0),.din(w_dff_A_UdfStCmJ6_0),.clk(gclk));
	jdff dff_A_M5Gc7Mn44_0(.dout(w_dff_A_ZoPEDEal0_0),.din(w_dff_A_M5Gc7Mn44_0),.clk(gclk));
	jdff dff_A_ZoPEDEal0_0(.dout(w_dff_A_MmoN4ZXN2_0),.din(w_dff_A_ZoPEDEal0_0),.clk(gclk));
	jdff dff_A_MmoN4ZXN2_0(.dout(w_dff_A_GvgcWzc66_0),.din(w_dff_A_MmoN4ZXN2_0),.clk(gclk));
	jdff dff_A_GvgcWzc66_0(.dout(w_dff_A_CopCHs636_0),.din(w_dff_A_GvgcWzc66_0),.clk(gclk));
	jdff dff_A_CopCHs636_0(.dout(w_dff_A_j2VkvqY69_0),.din(w_dff_A_CopCHs636_0),.clk(gclk));
	jdff dff_A_j2VkvqY69_0(.dout(w_dff_A_hSgVIXjW7_0),.din(w_dff_A_j2VkvqY69_0),.clk(gclk));
	jdff dff_A_hSgVIXjW7_0(.dout(w_dff_A_j2ztsuy43_0),.din(w_dff_A_hSgVIXjW7_0),.clk(gclk));
	jdff dff_A_j2ztsuy43_0(.dout(w_dff_A_v62F2IWC7_0),.din(w_dff_A_j2ztsuy43_0),.clk(gclk));
	jdff dff_A_v62F2IWC7_0(.dout(w_dff_A_6mpWp5Zf8_0),.din(w_dff_A_v62F2IWC7_0),.clk(gclk));
	jdff dff_A_6mpWp5Zf8_0(.dout(w_dff_A_tdtMLX1A3_0),.din(w_dff_A_6mpWp5Zf8_0),.clk(gclk));
	jdff dff_A_tdtMLX1A3_0(.dout(w_dff_A_2bhDzNnD9_0),.din(w_dff_A_tdtMLX1A3_0),.clk(gclk));
	jdff dff_A_2bhDzNnD9_0(.dout(w_dff_A_HBngTINL3_0),.din(w_dff_A_2bhDzNnD9_0),.clk(gclk));
	jdff dff_A_HBngTINL3_0(.dout(w_dff_A_44ZYftsj8_0),.din(w_dff_A_HBngTINL3_0),.clk(gclk));
	jdff dff_A_44ZYftsj8_0(.dout(w_dff_A_1T0wmQ9Q7_0),.din(w_dff_A_44ZYftsj8_0),.clk(gclk));
	jdff dff_A_1T0wmQ9Q7_0(.dout(w_dff_A_uwwWCaAN5_0),.din(w_dff_A_1T0wmQ9Q7_0),.clk(gclk));
	jdff dff_A_uwwWCaAN5_0(.dout(w_dff_A_OOVUengi4_0),.din(w_dff_A_uwwWCaAN5_0),.clk(gclk));
	jdff dff_A_OOVUengi4_0(.dout(w_dff_A_RiNYpsUZ4_0),.din(w_dff_A_OOVUengi4_0),.clk(gclk));
	jdff dff_A_RiNYpsUZ4_0(.dout(w_dff_A_pAz4n5Ij9_0),.din(w_dff_A_RiNYpsUZ4_0),.clk(gclk));
	jdff dff_A_pAz4n5Ij9_0(.dout(w_dff_A_2OUaKl2z8_0),.din(w_dff_A_pAz4n5Ij9_0),.clk(gclk));
	jdff dff_A_2OUaKl2z8_0(.dout(w_dff_A_ji4ZwdNe3_0),.din(w_dff_A_2OUaKl2z8_0),.clk(gclk));
	jdff dff_A_ji4ZwdNe3_0(.dout(w_dff_A_LEi7ziF49_0),.din(w_dff_A_ji4ZwdNe3_0),.clk(gclk));
	jdff dff_A_LEi7ziF49_0(.dout(w_dff_A_hHqfrAqe9_0),.din(w_dff_A_LEi7ziF49_0),.clk(gclk));
	jdff dff_A_hHqfrAqe9_0(.dout(w_dff_A_iafQQNhc1_0),.din(w_dff_A_hHqfrAqe9_0),.clk(gclk));
	jdff dff_A_iafQQNhc1_0(.dout(w_dff_A_qqEazY6k9_0),.din(w_dff_A_iafQQNhc1_0),.clk(gclk));
	jdff dff_A_qqEazY6k9_0(.dout(w_dff_A_Zjv5WxxK8_0),.din(w_dff_A_qqEazY6k9_0),.clk(gclk));
	jdff dff_A_Zjv5WxxK8_0(.dout(w_dff_A_QStrNx3z2_0),.din(w_dff_A_Zjv5WxxK8_0),.clk(gclk));
	jdff dff_A_QStrNx3z2_0(.dout(w_dff_A_iWUXfyjK0_0),.din(w_dff_A_QStrNx3z2_0),.clk(gclk));
	jdff dff_A_iWUXfyjK0_0(.dout(w_dff_A_QHqd1eQe9_0),.din(w_dff_A_iWUXfyjK0_0),.clk(gclk));
	jdff dff_A_QHqd1eQe9_0(.dout(w_dff_A_s5bR2fBA6_0),.din(w_dff_A_QHqd1eQe9_0),.clk(gclk));
	jdff dff_A_s5bR2fBA6_0(.dout(w_dff_A_7CjraK4O8_0),.din(w_dff_A_s5bR2fBA6_0),.clk(gclk));
	jdff dff_A_7CjraK4O8_0(.dout(w_dff_A_sra1MCyW3_0),.din(w_dff_A_7CjraK4O8_0),.clk(gclk));
	jdff dff_A_sra1MCyW3_0(.dout(w_dff_A_NqVRCeBe6_0),.din(w_dff_A_sra1MCyW3_0),.clk(gclk));
	jdff dff_A_NqVRCeBe6_0(.dout(w_dff_A_gewLgLH49_0),.din(w_dff_A_NqVRCeBe6_0),.clk(gclk));
	jdff dff_A_gewLgLH49_0(.dout(w_dff_A_yeUuBgYH3_0),.din(w_dff_A_gewLgLH49_0),.clk(gclk));
	jdff dff_A_yeUuBgYH3_0(.dout(w_dff_A_e5RL9Fr17_0),.din(w_dff_A_yeUuBgYH3_0),.clk(gclk));
	jdff dff_A_e5RL9Fr17_0(.dout(w_dff_A_vkcrJACS5_0),.din(w_dff_A_e5RL9Fr17_0),.clk(gclk));
	jdff dff_A_vkcrJACS5_0(.dout(w_dff_A_FvGyzLDv6_0),.din(w_dff_A_vkcrJACS5_0),.clk(gclk));
	jdff dff_A_FvGyzLDv6_0(.dout(w_dff_A_ynJToruf2_0),.din(w_dff_A_FvGyzLDv6_0),.clk(gclk));
	jdff dff_A_ynJToruf2_0(.dout(w_dff_A_ibkW8z117_0),.din(w_dff_A_ynJToruf2_0),.clk(gclk));
	jdff dff_A_ibkW8z117_0(.dout(w_dff_A_xQSrxj0P4_0),.din(w_dff_A_ibkW8z117_0),.clk(gclk));
	jdff dff_A_xQSrxj0P4_0(.dout(w_dff_A_us00chUJ7_0),.din(w_dff_A_xQSrxj0P4_0),.clk(gclk));
	jdff dff_A_us00chUJ7_0(.dout(w_dff_A_v1nt2IXZ5_0),.din(w_dff_A_us00chUJ7_0),.clk(gclk));
	jdff dff_A_v1nt2IXZ5_0(.dout(w_dff_A_B2YdVD7m5_0),.din(w_dff_A_v1nt2IXZ5_0),.clk(gclk));
	jdff dff_A_B2YdVD7m5_0(.dout(w_dff_A_fBkfM7Dk9_0),.din(w_dff_A_B2YdVD7m5_0),.clk(gclk));
	jdff dff_A_fBkfM7Dk9_0(.dout(w_dff_A_T9ce9Asc0_0),.din(w_dff_A_fBkfM7Dk9_0),.clk(gclk));
	jdff dff_A_T9ce9Asc0_0(.dout(w_dff_A_yLpw7GaN3_0),.din(w_dff_A_T9ce9Asc0_0),.clk(gclk));
	jdff dff_A_yLpw7GaN3_0(.dout(w_dff_A_Zr3ERBvI4_0),.din(w_dff_A_yLpw7GaN3_0),.clk(gclk));
	jdff dff_A_Zr3ERBvI4_0(.dout(w_dff_A_xcp2VARa5_0),.din(w_dff_A_Zr3ERBvI4_0),.clk(gclk));
	jdff dff_A_xcp2VARa5_0(.dout(w_dff_A_zVbkba7S3_0),.din(w_dff_A_xcp2VARa5_0),.clk(gclk));
	jdff dff_A_zVbkba7S3_0(.dout(w_dff_A_sepVj1Tp8_0),.din(w_dff_A_zVbkba7S3_0),.clk(gclk));
	jdff dff_A_sepVj1Tp8_0(.dout(w_dff_A_22FGuTkW5_0),.din(w_dff_A_sepVj1Tp8_0),.clk(gclk));
	jdff dff_A_22FGuTkW5_0(.dout(w_dff_A_sVhuT3xV8_0),.din(w_dff_A_22FGuTkW5_0),.clk(gclk));
	jdff dff_A_sVhuT3xV8_0(.dout(w_dff_A_e975MbsB1_0),.din(w_dff_A_sVhuT3xV8_0),.clk(gclk));
	jdff dff_A_e975MbsB1_0(.dout(w_dff_A_l2UfLZWH9_0),.din(w_dff_A_e975MbsB1_0),.clk(gclk));
	jdff dff_A_l2UfLZWH9_0(.dout(w_dff_A_KRDcwiQT3_0),.din(w_dff_A_l2UfLZWH9_0),.clk(gclk));
	jdff dff_A_KRDcwiQT3_0(.dout(w_dff_A_U8omtxaO8_0),.din(w_dff_A_KRDcwiQT3_0),.clk(gclk));
	jdff dff_A_U8omtxaO8_0(.dout(w_dff_A_5AqRMy096_0),.din(w_dff_A_U8omtxaO8_0),.clk(gclk));
	jdff dff_A_5AqRMy096_0(.dout(w_dff_A_cnOOCoKZ5_0),.din(w_dff_A_5AqRMy096_0),.clk(gclk));
	jdff dff_A_cnOOCoKZ5_0(.dout(w_dff_A_TBTHLLdM3_0),.din(w_dff_A_cnOOCoKZ5_0),.clk(gclk));
	jdff dff_A_TBTHLLdM3_0(.dout(w_dff_A_cZdjRu643_0),.din(w_dff_A_TBTHLLdM3_0),.clk(gclk));
	jdff dff_A_cZdjRu643_0(.dout(w_dff_A_8e6dsy809_0),.din(w_dff_A_cZdjRu643_0),.clk(gclk));
	jdff dff_A_8e6dsy809_0(.dout(w_dff_A_v9hUv4tu3_0),.din(w_dff_A_8e6dsy809_0),.clk(gclk));
	jdff dff_A_v9hUv4tu3_0(.dout(G1581gat),.din(w_dff_A_v9hUv4tu3_0),.clk(gclk));
	jdff dff_A_JVhOTcac7_2(.dout(w_dff_A_NT76UVWY5_0),.din(w_dff_A_JVhOTcac7_2),.clk(gclk));
	jdff dff_A_NT76UVWY5_0(.dout(w_dff_A_824KkLKS4_0),.din(w_dff_A_NT76UVWY5_0),.clk(gclk));
	jdff dff_A_824KkLKS4_0(.dout(w_dff_A_fMtPH8fD4_0),.din(w_dff_A_824KkLKS4_0),.clk(gclk));
	jdff dff_A_fMtPH8fD4_0(.dout(w_dff_A_VJyafekE9_0),.din(w_dff_A_fMtPH8fD4_0),.clk(gclk));
	jdff dff_A_VJyafekE9_0(.dout(w_dff_A_ID3HfpM18_0),.din(w_dff_A_VJyafekE9_0),.clk(gclk));
	jdff dff_A_ID3HfpM18_0(.dout(w_dff_A_Xa9r3keL2_0),.din(w_dff_A_ID3HfpM18_0),.clk(gclk));
	jdff dff_A_Xa9r3keL2_0(.dout(w_dff_A_fGqx4EVW3_0),.din(w_dff_A_Xa9r3keL2_0),.clk(gclk));
	jdff dff_A_fGqx4EVW3_0(.dout(w_dff_A_u5QbZPUF0_0),.din(w_dff_A_fGqx4EVW3_0),.clk(gclk));
	jdff dff_A_u5QbZPUF0_0(.dout(w_dff_A_e9Mq2UPP9_0),.din(w_dff_A_u5QbZPUF0_0),.clk(gclk));
	jdff dff_A_e9Mq2UPP9_0(.dout(w_dff_A_HhxrEXQQ2_0),.din(w_dff_A_e9Mq2UPP9_0),.clk(gclk));
	jdff dff_A_HhxrEXQQ2_0(.dout(w_dff_A_Gnnlkr3h1_0),.din(w_dff_A_HhxrEXQQ2_0),.clk(gclk));
	jdff dff_A_Gnnlkr3h1_0(.dout(w_dff_A_pUiflOiD1_0),.din(w_dff_A_Gnnlkr3h1_0),.clk(gclk));
	jdff dff_A_pUiflOiD1_0(.dout(w_dff_A_2lKeuyZs8_0),.din(w_dff_A_pUiflOiD1_0),.clk(gclk));
	jdff dff_A_2lKeuyZs8_0(.dout(w_dff_A_NFITlDAY8_0),.din(w_dff_A_2lKeuyZs8_0),.clk(gclk));
	jdff dff_A_NFITlDAY8_0(.dout(w_dff_A_hNdIgJyg0_0),.din(w_dff_A_NFITlDAY8_0),.clk(gclk));
	jdff dff_A_hNdIgJyg0_0(.dout(w_dff_A_7CtlbZyX5_0),.din(w_dff_A_hNdIgJyg0_0),.clk(gclk));
	jdff dff_A_7CtlbZyX5_0(.dout(w_dff_A_8hqeXyt36_0),.din(w_dff_A_7CtlbZyX5_0),.clk(gclk));
	jdff dff_A_8hqeXyt36_0(.dout(w_dff_A_133QnD3y4_0),.din(w_dff_A_8hqeXyt36_0),.clk(gclk));
	jdff dff_A_133QnD3y4_0(.dout(w_dff_A_tGlBxxaP5_0),.din(w_dff_A_133QnD3y4_0),.clk(gclk));
	jdff dff_A_tGlBxxaP5_0(.dout(w_dff_A_D0bWv7nh6_0),.din(w_dff_A_tGlBxxaP5_0),.clk(gclk));
	jdff dff_A_D0bWv7nh6_0(.dout(w_dff_A_KBQxncBm3_0),.din(w_dff_A_D0bWv7nh6_0),.clk(gclk));
	jdff dff_A_KBQxncBm3_0(.dout(w_dff_A_07Znfa8p1_0),.din(w_dff_A_KBQxncBm3_0),.clk(gclk));
	jdff dff_A_07Znfa8p1_0(.dout(w_dff_A_UhdnXtKU9_0),.din(w_dff_A_07Znfa8p1_0),.clk(gclk));
	jdff dff_A_UhdnXtKU9_0(.dout(w_dff_A_WmTEDsOs8_0),.din(w_dff_A_UhdnXtKU9_0),.clk(gclk));
	jdff dff_A_WmTEDsOs8_0(.dout(w_dff_A_1xzJKcZs7_0),.din(w_dff_A_WmTEDsOs8_0),.clk(gclk));
	jdff dff_A_1xzJKcZs7_0(.dout(w_dff_A_QTjy2HHt2_0),.din(w_dff_A_1xzJKcZs7_0),.clk(gclk));
	jdff dff_A_QTjy2HHt2_0(.dout(w_dff_A_ngxFGTSy8_0),.din(w_dff_A_QTjy2HHt2_0),.clk(gclk));
	jdff dff_A_ngxFGTSy8_0(.dout(w_dff_A_Kwl2yqEI4_0),.din(w_dff_A_ngxFGTSy8_0),.clk(gclk));
	jdff dff_A_Kwl2yqEI4_0(.dout(w_dff_A_fqgXS9d36_0),.din(w_dff_A_Kwl2yqEI4_0),.clk(gclk));
	jdff dff_A_fqgXS9d36_0(.dout(w_dff_A_97CxQrb70_0),.din(w_dff_A_fqgXS9d36_0),.clk(gclk));
	jdff dff_A_97CxQrb70_0(.dout(w_dff_A_tYGfJabt2_0),.din(w_dff_A_97CxQrb70_0),.clk(gclk));
	jdff dff_A_tYGfJabt2_0(.dout(w_dff_A_wkMNkgim6_0),.din(w_dff_A_tYGfJabt2_0),.clk(gclk));
	jdff dff_A_wkMNkgim6_0(.dout(w_dff_A_xNUMPrWg3_0),.din(w_dff_A_wkMNkgim6_0),.clk(gclk));
	jdff dff_A_xNUMPrWg3_0(.dout(w_dff_A_0RGdBZxN3_0),.din(w_dff_A_xNUMPrWg3_0),.clk(gclk));
	jdff dff_A_0RGdBZxN3_0(.dout(w_dff_A_kFROo3MS8_0),.din(w_dff_A_0RGdBZxN3_0),.clk(gclk));
	jdff dff_A_kFROo3MS8_0(.dout(w_dff_A_WdROrC0j6_0),.din(w_dff_A_kFROo3MS8_0),.clk(gclk));
	jdff dff_A_WdROrC0j6_0(.dout(w_dff_A_Ej6knU7C6_0),.din(w_dff_A_WdROrC0j6_0),.clk(gclk));
	jdff dff_A_Ej6knU7C6_0(.dout(w_dff_A_68COWNWm6_0),.din(w_dff_A_Ej6knU7C6_0),.clk(gclk));
	jdff dff_A_68COWNWm6_0(.dout(w_dff_A_Fs6yXC0n1_0),.din(w_dff_A_68COWNWm6_0),.clk(gclk));
	jdff dff_A_Fs6yXC0n1_0(.dout(w_dff_A_FcdE4FeK9_0),.din(w_dff_A_Fs6yXC0n1_0),.clk(gclk));
	jdff dff_A_FcdE4FeK9_0(.dout(w_dff_A_8UgCSxG51_0),.din(w_dff_A_FcdE4FeK9_0),.clk(gclk));
	jdff dff_A_8UgCSxG51_0(.dout(w_dff_A_sXMumqT44_0),.din(w_dff_A_8UgCSxG51_0),.clk(gclk));
	jdff dff_A_sXMumqT44_0(.dout(w_dff_A_0HM10aIA2_0),.din(w_dff_A_sXMumqT44_0),.clk(gclk));
	jdff dff_A_0HM10aIA2_0(.dout(w_dff_A_8FeN6LaS6_0),.din(w_dff_A_0HM10aIA2_0),.clk(gclk));
	jdff dff_A_8FeN6LaS6_0(.dout(w_dff_A_x1E0F7KP0_0),.din(w_dff_A_8FeN6LaS6_0),.clk(gclk));
	jdff dff_A_x1E0F7KP0_0(.dout(w_dff_A_YjWzstNl3_0),.din(w_dff_A_x1E0F7KP0_0),.clk(gclk));
	jdff dff_A_YjWzstNl3_0(.dout(w_dff_A_ZXNeWPsI9_0),.din(w_dff_A_YjWzstNl3_0),.clk(gclk));
	jdff dff_A_ZXNeWPsI9_0(.dout(w_dff_A_C4jqsiD09_0),.din(w_dff_A_ZXNeWPsI9_0),.clk(gclk));
	jdff dff_A_C4jqsiD09_0(.dout(w_dff_A_aiXV3y6k9_0),.din(w_dff_A_C4jqsiD09_0),.clk(gclk));
	jdff dff_A_aiXV3y6k9_0(.dout(w_dff_A_PiXCjjyt8_0),.din(w_dff_A_aiXV3y6k9_0),.clk(gclk));
	jdff dff_A_PiXCjjyt8_0(.dout(w_dff_A_FIhdjpn42_0),.din(w_dff_A_PiXCjjyt8_0),.clk(gclk));
	jdff dff_A_FIhdjpn42_0(.dout(w_dff_A_psrtXOYz5_0),.din(w_dff_A_FIhdjpn42_0),.clk(gclk));
	jdff dff_A_psrtXOYz5_0(.dout(w_dff_A_Inpql7wC1_0),.din(w_dff_A_psrtXOYz5_0),.clk(gclk));
	jdff dff_A_Inpql7wC1_0(.dout(w_dff_A_uqk1M2Gx6_0),.din(w_dff_A_Inpql7wC1_0),.clk(gclk));
	jdff dff_A_uqk1M2Gx6_0(.dout(w_dff_A_Q2CUbeza0_0),.din(w_dff_A_uqk1M2Gx6_0),.clk(gclk));
	jdff dff_A_Q2CUbeza0_0(.dout(w_dff_A_g0oU4rgc8_0),.din(w_dff_A_Q2CUbeza0_0),.clk(gclk));
	jdff dff_A_g0oU4rgc8_0(.dout(w_dff_A_gDlYcnpp3_0),.din(w_dff_A_g0oU4rgc8_0),.clk(gclk));
	jdff dff_A_gDlYcnpp3_0(.dout(w_dff_A_p0MP5Sde4_0),.din(w_dff_A_gDlYcnpp3_0),.clk(gclk));
	jdff dff_A_p0MP5Sde4_0(.dout(w_dff_A_Q8nhhH208_0),.din(w_dff_A_p0MP5Sde4_0),.clk(gclk));
	jdff dff_A_Q8nhhH208_0(.dout(w_dff_A_9LIkbH8r7_0),.din(w_dff_A_Q8nhhH208_0),.clk(gclk));
	jdff dff_A_9LIkbH8r7_0(.dout(w_dff_A_xOmjsfo56_0),.din(w_dff_A_9LIkbH8r7_0),.clk(gclk));
	jdff dff_A_xOmjsfo56_0(.dout(w_dff_A_fpXNrvut3_0),.din(w_dff_A_xOmjsfo56_0),.clk(gclk));
	jdff dff_A_fpXNrvut3_0(.dout(w_dff_A_yEu7myOq6_0),.din(w_dff_A_fpXNrvut3_0),.clk(gclk));
	jdff dff_A_yEu7myOq6_0(.dout(w_dff_A_I7iEgpZ91_0),.din(w_dff_A_yEu7myOq6_0),.clk(gclk));
	jdff dff_A_I7iEgpZ91_0(.dout(w_dff_A_TFyM6XWr9_0),.din(w_dff_A_I7iEgpZ91_0),.clk(gclk));
	jdff dff_A_TFyM6XWr9_0(.dout(w_dff_A_170TZJca6_0),.din(w_dff_A_TFyM6XWr9_0),.clk(gclk));
	jdff dff_A_170TZJca6_0(.dout(w_dff_A_omAAnoaQ4_0),.din(w_dff_A_170TZJca6_0),.clk(gclk));
	jdff dff_A_omAAnoaQ4_0(.dout(w_dff_A_Ipkfrq3U1_0),.din(w_dff_A_omAAnoaQ4_0),.clk(gclk));
	jdff dff_A_Ipkfrq3U1_0(.dout(G1901gat),.din(w_dff_A_Ipkfrq3U1_0),.clk(gclk));
	jdff dff_A_1yMaWZic3_2(.dout(w_dff_A_8X9du1RG9_0),.din(w_dff_A_1yMaWZic3_2),.clk(gclk));
	jdff dff_A_8X9du1RG9_0(.dout(w_dff_A_rFVpRbud2_0),.din(w_dff_A_8X9du1RG9_0),.clk(gclk));
	jdff dff_A_rFVpRbud2_0(.dout(w_dff_A_ErdpTLjR2_0),.din(w_dff_A_rFVpRbud2_0),.clk(gclk));
	jdff dff_A_ErdpTLjR2_0(.dout(w_dff_A_s05MepAb6_0),.din(w_dff_A_ErdpTLjR2_0),.clk(gclk));
	jdff dff_A_s05MepAb6_0(.dout(w_dff_A_TWufy2BV1_0),.din(w_dff_A_s05MepAb6_0),.clk(gclk));
	jdff dff_A_TWufy2BV1_0(.dout(w_dff_A_x4kecnmA0_0),.din(w_dff_A_TWufy2BV1_0),.clk(gclk));
	jdff dff_A_x4kecnmA0_0(.dout(w_dff_A_KyKEaOsH1_0),.din(w_dff_A_x4kecnmA0_0),.clk(gclk));
	jdff dff_A_KyKEaOsH1_0(.dout(w_dff_A_PrEVD5yV7_0),.din(w_dff_A_KyKEaOsH1_0),.clk(gclk));
	jdff dff_A_PrEVD5yV7_0(.dout(w_dff_A_b0TfVYAn0_0),.din(w_dff_A_PrEVD5yV7_0),.clk(gclk));
	jdff dff_A_b0TfVYAn0_0(.dout(w_dff_A_IbuQTzem8_0),.din(w_dff_A_b0TfVYAn0_0),.clk(gclk));
	jdff dff_A_IbuQTzem8_0(.dout(w_dff_A_R8NDF07a2_0),.din(w_dff_A_IbuQTzem8_0),.clk(gclk));
	jdff dff_A_R8NDF07a2_0(.dout(w_dff_A_JElYusPA3_0),.din(w_dff_A_R8NDF07a2_0),.clk(gclk));
	jdff dff_A_JElYusPA3_0(.dout(w_dff_A_CFpjbw0M6_0),.din(w_dff_A_JElYusPA3_0),.clk(gclk));
	jdff dff_A_CFpjbw0M6_0(.dout(w_dff_A_jENwXvRN6_0),.din(w_dff_A_CFpjbw0M6_0),.clk(gclk));
	jdff dff_A_jENwXvRN6_0(.dout(w_dff_A_Re96E3ou3_0),.din(w_dff_A_jENwXvRN6_0),.clk(gclk));
	jdff dff_A_Re96E3ou3_0(.dout(w_dff_A_Yvw7I55z3_0),.din(w_dff_A_Re96E3ou3_0),.clk(gclk));
	jdff dff_A_Yvw7I55z3_0(.dout(w_dff_A_SY9Td5QQ8_0),.din(w_dff_A_Yvw7I55z3_0),.clk(gclk));
	jdff dff_A_SY9Td5QQ8_0(.dout(w_dff_A_cjVJyWL80_0),.din(w_dff_A_SY9Td5QQ8_0),.clk(gclk));
	jdff dff_A_cjVJyWL80_0(.dout(w_dff_A_xY6YpDOM2_0),.din(w_dff_A_cjVJyWL80_0),.clk(gclk));
	jdff dff_A_xY6YpDOM2_0(.dout(w_dff_A_wzuAUU8H2_0),.din(w_dff_A_xY6YpDOM2_0),.clk(gclk));
	jdff dff_A_wzuAUU8H2_0(.dout(w_dff_A_8JLkeZUI0_0),.din(w_dff_A_wzuAUU8H2_0),.clk(gclk));
	jdff dff_A_8JLkeZUI0_0(.dout(w_dff_A_uheqYr9h6_0),.din(w_dff_A_8JLkeZUI0_0),.clk(gclk));
	jdff dff_A_uheqYr9h6_0(.dout(w_dff_A_iVzxobba6_0),.din(w_dff_A_uheqYr9h6_0),.clk(gclk));
	jdff dff_A_iVzxobba6_0(.dout(w_dff_A_GMDtooMm0_0),.din(w_dff_A_iVzxobba6_0),.clk(gclk));
	jdff dff_A_GMDtooMm0_0(.dout(w_dff_A_8gG22on23_0),.din(w_dff_A_GMDtooMm0_0),.clk(gclk));
	jdff dff_A_8gG22on23_0(.dout(w_dff_A_igzkPXVb7_0),.din(w_dff_A_8gG22on23_0),.clk(gclk));
	jdff dff_A_igzkPXVb7_0(.dout(w_dff_A_RMxLWcNl9_0),.din(w_dff_A_igzkPXVb7_0),.clk(gclk));
	jdff dff_A_RMxLWcNl9_0(.dout(w_dff_A_vIpiASBy9_0),.din(w_dff_A_RMxLWcNl9_0),.clk(gclk));
	jdff dff_A_vIpiASBy9_0(.dout(w_dff_A_WV4kVZTz5_0),.din(w_dff_A_vIpiASBy9_0),.clk(gclk));
	jdff dff_A_WV4kVZTz5_0(.dout(w_dff_A_oAmK9mjk3_0),.din(w_dff_A_WV4kVZTz5_0),.clk(gclk));
	jdff dff_A_oAmK9mjk3_0(.dout(w_dff_A_Ar1CFKkr3_0),.din(w_dff_A_oAmK9mjk3_0),.clk(gclk));
	jdff dff_A_Ar1CFKkr3_0(.dout(w_dff_A_gAgW4Gp38_0),.din(w_dff_A_Ar1CFKkr3_0),.clk(gclk));
	jdff dff_A_gAgW4Gp38_0(.dout(w_dff_A_L782zogU6_0),.din(w_dff_A_gAgW4Gp38_0),.clk(gclk));
	jdff dff_A_L782zogU6_0(.dout(w_dff_A_q47g306l8_0),.din(w_dff_A_L782zogU6_0),.clk(gclk));
	jdff dff_A_q47g306l8_0(.dout(w_dff_A_vcwRjrh79_0),.din(w_dff_A_q47g306l8_0),.clk(gclk));
	jdff dff_A_vcwRjrh79_0(.dout(w_dff_A_PHocqwJc6_0),.din(w_dff_A_vcwRjrh79_0),.clk(gclk));
	jdff dff_A_PHocqwJc6_0(.dout(w_dff_A_xBN6Utg09_0),.din(w_dff_A_PHocqwJc6_0),.clk(gclk));
	jdff dff_A_xBN6Utg09_0(.dout(w_dff_A_sggvOKUn2_0),.din(w_dff_A_xBN6Utg09_0),.clk(gclk));
	jdff dff_A_sggvOKUn2_0(.dout(w_dff_A_4AZEIa1j1_0),.din(w_dff_A_sggvOKUn2_0),.clk(gclk));
	jdff dff_A_4AZEIa1j1_0(.dout(w_dff_A_j2Rwxy2r9_0),.din(w_dff_A_4AZEIa1j1_0),.clk(gclk));
	jdff dff_A_j2Rwxy2r9_0(.dout(w_dff_A_TKYfrazv0_0),.din(w_dff_A_j2Rwxy2r9_0),.clk(gclk));
	jdff dff_A_TKYfrazv0_0(.dout(w_dff_A_77NnLVCI7_0),.din(w_dff_A_TKYfrazv0_0),.clk(gclk));
	jdff dff_A_77NnLVCI7_0(.dout(w_dff_A_BeqkVDrE2_0),.din(w_dff_A_77NnLVCI7_0),.clk(gclk));
	jdff dff_A_BeqkVDrE2_0(.dout(w_dff_A_ZPJpWdwx2_0),.din(w_dff_A_BeqkVDrE2_0),.clk(gclk));
	jdff dff_A_ZPJpWdwx2_0(.dout(w_dff_A_X2SBdZSj6_0),.din(w_dff_A_ZPJpWdwx2_0),.clk(gclk));
	jdff dff_A_X2SBdZSj6_0(.dout(w_dff_A_uUOBhka81_0),.din(w_dff_A_X2SBdZSj6_0),.clk(gclk));
	jdff dff_A_uUOBhka81_0(.dout(w_dff_A_iRgeIgQo3_0),.din(w_dff_A_uUOBhka81_0),.clk(gclk));
	jdff dff_A_iRgeIgQo3_0(.dout(w_dff_A_KcS4N9bR1_0),.din(w_dff_A_iRgeIgQo3_0),.clk(gclk));
	jdff dff_A_KcS4N9bR1_0(.dout(w_dff_A_VwK39ooS6_0),.din(w_dff_A_KcS4N9bR1_0),.clk(gclk));
	jdff dff_A_VwK39ooS6_0(.dout(w_dff_A_16XwVVWG5_0),.din(w_dff_A_VwK39ooS6_0),.clk(gclk));
	jdff dff_A_16XwVVWG5_0(.dout(w_dff_A_wbdI8snT1_0),.din(w_dff_A_16XwVVWG5_0),.clk(gclk));
	jdff dff_A_wbdI8snT1_0(.dout(w_dff_A_irtJAX4c7_0),.din(w_dff_A_wbdI8snT1_0),.clk(gclk));
	jdff dff_A_irtJAX4c7_0(.dout(w_dff_A_Yr0yTxxK8_0),.din(w_dff_A_irtJAX4c7_0),.clk(gclk));
	jdff dff_A_Yr0yTxxK8_0(.dout(w_dff_A_JkE0mIGb2_0),.din(w_dff_A_Yr0yTxxK8_0),.clk(gclk));
	jdff dff_A_JkE0mIGb2_0(.dout(w_dff_A_vtt15bAz7_0),.din(w_dff_A_JkE0mIGb2_0),.clk(gclk));
	jdff dff_A_vtt15bAz7_0(.dout(w_dff_A_Lusgj4m97_0),.din(w_dff_A_vtt15bAz7_0),.clk(gclk));
	jdff dff_A_Lusgj4m97_0(.dout(w_dff_A_PNV4wddq2_0),.din(w_dff_A_Lusgj4m97_0),.clk(gclk));
	jdff dff_A_PNV4wddq2_0(.dout(w_dff_A_ViDl5Bzk1_0),.din(w_dff_A_PNV4wddq2_0),.clk(gclk));
	jdff dff_A_ViDl5Bzk1_0(.dout(w_dff_A_IMNEaPK70_0),.din(w_dff_A_ViDl5Bzk1_0),.clk(gclk));
	jdff dff_A_IMNEaPK70_0(.dout(w_dff_A_udqJLdeb9_0),.din(w_dff_A_IMNEaPK70_0),.clk(gclk));
	jdff dff_A_udqJLdeb9_0(.dout(w_dff_A_ryLHRJvm6_0),.din(w_dff_A_udqJLdeb9_0),.clk(gclk));
	jdff dff_A_ryLHRJvm6_0(.dout(w_dff_A_lLEhQVjI2_0),.din(w_dff_A_ryLHRJvm6_0),.clk(gclk));
	jdff dff_A_lLEhQVjI2_0(.dout(w_dff_A_CxReM8mW6_0),.din(w_dff_A_lLEhQVjI2_0),.clk(gclk));
	jdff dff_A_CxReM8mW6_0(.dout(w_dff_A_0FjEIobv2_0),.din(w_dff_A_CxReM8mW6_0),.clk(gclk));
	jdff dff_A_0FjEIobv2_0(.dout(w_dff_A_lY17I36C2_0),.din(w_dff_A_0FjEIobv2_0),.clk(gclk));
	jdff dff_A_lY17I36C2_0(.dout(G2223gat),.din(w_dff_A_lY17I36C2_0),.clk(gclk));
	jdff dff_A_THDtcXMv5_2(.dout(w_dff_A_ODbkMDGw9_0),.din(w_dff_A_THDtcXMv5_2),.clk(gclk));
	jdff dff_A_ODbkMDGw9_0(.dout(w_dff_A_yzRjjQb78_0),.din(w_dff_A_ODbkMDGw9_0),.clk(gclk));
	jdff dff_A_yzRjjQb78_0(.dout(w_dff_A_nx7lV8ZY8_0),.din(w_dff_A_yzRjjQb78_0),.clk(gclk));
	jdff dff_A_nx7lV8ZY8_0(.dout(w_dff_A_6GBtMk3S7_0),.din(w_dff_A_nx7lV8ZY8_0),.clk(gclk));
	jdff dff_A_6GBtMk3S7_0(.dout(w_dff_A_t4n3Vxnp3_0),.din(w_dff_A_6GBtMk3S7_0),.clk(gclk));
	jdff dff_A_t4n3Vxnp3_0(.dout(w_dff_A_gnWkttWm2_0),.din(w_dff_A_t4n3Vxnp3_0),.clk(gclk));
	jdff dff_A_gnWkttWm2_0(.dout(w_dff_A_Ws57iV842_0),.din(w_dff_A_gnWkttWm2_0),.clk(gclk));
	jdff dff_A_Ws57iV842_0(.dout(w_dff_A_IyKUKQ4n2_0),.din(w_dff_A_Ws57iV842_0),.clk(gclk));
	jdff dff_A_IyKUKQ4n2_0(.dout(w_dff_A_mcq8eNv20_0),.din(w_dff_A_IyKUKQ4n2_0),.clk(gclk));
	jdff dff_A_mcq8eNv20_0(.dout(w_dff_A_XRGRVtm78_0),.din(w_dff_A_mcq8eNv20_0),.clk(gclk));
	jdff dff_A_XRGRVtm78_0(.dout(w_dff_A_qXiDv2w52_0),.din(w_dff_A_XRGRVtm78_0),.clk(gclk));
	jdff dff_A_qXiDv2w52_0(.dout(w_dff_A_MUAd3p4d7_0),.din(w_dff_A_qXiDv2w52_0),.clk(gclk));
	jdff dff_A_MUAd3p4d7_0(.dout(w_dff_A_EAaQ7z5e5_0),.din(w_dff_A_MUAd3p4d7_0),.clk(gclk));
	jdff dff_A_EAaQ7z5e5_0(.dout(w_dff_A_BpGXNOAY0_0),.din(w_dff_A_EAaQ7z5e5_0),.clk(gclk));
	jdff dff_A_BpGXNOAY0_0(.dout(w_dff_A_g7OYbm2x0_0),.din(w_dff_A_BpGXNOAY0_0),.clk(gclk));
	jdff dff_A_g7OYbm2x0_0(.dout(w_dff_A_xHo15xPE7_0),.din(w_dff_A_g7OYbm2x0_0),.clk(gclk));
	jdff dff_A_xHo15xPE7_0(.dout(w_dff_A_gpvHEGao3_0),.din(w_dff_A_xHo15xPE7_0),.clk(gclk));
	jdff dff_A_gpvHEGao3_0(.dout(w_dff_A_aUF0kOJh8_0),.din(w_dff_A_gpvHEGao3_0),.clk(gclk));
	jdff dff_A_aUF0kOJh8_0(.dout(w_dff_A_Kj8vqFVc2_0),.din(w_dff_A_aUF0kOJh8_0),.clk(gclk));
	jdff dff_A_Kj8vqFVc2_0(.dout(w_dff_A_BKloISGC6_0),.din(w_dff_A_Kj8vqFVc2_0),.clk(gclk));
	jdff dff_A_BKloISGC6_0(.dout(w_dff_A_Zvmu7Wwi2_0),.din(w_dff_A_BKloISGC6_0),.clk(gclk));
	jdff dff_A_Zvmu7Wwi2_0(.dout(w_dff_A_fyaRnmnx2_0),.din(w_dff_A_Zvmu7Wwi2_0),.clk(gclk));
	jdff dff_A_fyaRnmnx2_0(.dout(w_dff_A_Ay3fC7ts7_0),.din(w_dff_A_fyaRnmnx2_0),.clk(gclk));
	jdff dff_A_Ay3fC7ts7_0(.dout(w_dff_A_hCAdJnNv5_0),.din(w_dff_A_Ay3fC7ts7_0),.clk(gclk));
	jdff dff_A_hCAdJnNv5_0(.dout(w_dff_A_pPlhb8708_0),.din(w_dff_A_hCAdJnNv5_0),.clk(gclk));
	jdff dff_A_pPlhb8708_0(.dout(w_dff_A_WbSZbNhz6_0),.din(w_dff_A_pPlhb8708_0),.clk(gclk));
	jdff dff_A_WbSZbNhz6_0(.dout(w_dff_A_oWvcKqrA4_0),.din(w_dff_A_WbSZbNhz6_0),.clk(gclk));
	jdff dff_A_oWvcKqrA4_0(.dout(w_dff_A_WW2TlCyv3_0),.din(w_dff_A_oWvcKqrA4_0),.clk(gclk));
	jdff dff_A_WW2TlCyv3_0(.dout(w_dff_A_f8uAFxet7_0),.din(w_dff_A_WW2TlCyv3_0),.clk(gclk));
	jdff dff_A_f8uAFxet7_0(.dout(w_dff_A_1pdyoYeS8_0),.din(w_dff_A_f8uAFxet7_0),.clk(gclk));
	jdff dff_A_1pdyoYeS8_0(.dout(w_dff_A_QD0p07Am6_0),.din(w_dff_A_1pdyoYeS8_0),.clk(gclk));
	jdff dff_A_QD0p07Am6_0(.dout(w_dff_A_d8P6ylwF7_0),.din(w_dff_A_QD0p07Am6_0),.clk(gclk));
	jdff dff_A_d8P6ylwF7_0(.dout(w_dff_A_Lgm8zHoN0_0),.din(w_dff_A_d8P6ylwF7_0),.clk(gclk));
	jdff dff_A_Lgm8zHoN0_0(.dout(w_dff_A_6t3link02_0),.din(w_dff_A_Lgm8zHoN0_0),.clk(gclk));
	jdff dff_A_6t3link02_0(.dout(w_dff_A_8d8p2Gyi8_0),.din(w_dff_A_6t3link02_0),.clk(gclk));
	jdff dff_A_8d8p2Gyi8_0(.dout(w_dff_A_hoTGXh7o0_0),.din(w_dff_A_8d8p2Gyi8_0),.clk(gclk));
	jdff dff_A_hoTGXh7o0_0(.dout(w_dff_A_AB0CsfNW1_0),.din(w_dff_A_hoTGXh7o0_0),.clk(gclk));
	jdff dff_A_AB0CsfNW1_0(.dout(w_dff_A_seXohdPi0_0),.din(w_dff_A_AB0CsfNW1_0),.clk(gclk));
	jdff dff_A_seXohdPi0_0(.dout(w_dff_A_mTmIwOWB9_0),.din(w_dff_A_seXohdPi0_0),.clk(gclk));
	jdff dff_A_mTmIwOWB9_0(.dout(w_dff_A_Po82cIcz8_0),.din(w_dff_A_mTmIwOWB9_0),.clk(gclk));
	jdff dff_A_Po82cIcz8_0(.dout(w_dff_A_NFQrKPGr7_0),.din(w_dff_A_Po82cIcz8_0),.clk(gclk));
	jdff dff_A_NFQrKPGr7_0(.dout(w_dff_A_x1aK2mS70_0),.din(w_dff_A_NFQrKPGr7_0),.clk(gclk));
	jdff dff_A_x1aK2mS70_0(.dout(w_dff_A_2eaFZj3w8_0),.din(w_dff_A_x1aK2mS70_0),.clk(gclk));
	jdff dff_A_2eaFZj3w8_0(.dout(w_dff_A_zFNlT83p8_0),.din(w_dff_A_2eaFZj3w8_0),.clk(gclk));
	jdff dff_A_zFNlT83p8_0(.dout(w_dff_A_tqjlsVox0_0),.din(w_dff_A_zFNlT83p8_0),.clk(gclk));
	jdff dff_A_tqjlsVox0_0(.dout(w_dff_A_yIwuicAw7_0),.din(w_dff_A_tqjlsVox0_0),.clk(gclk));
	jdff dff_A_yIwuicAw7_0(.dout(w_dff_A_0x4CTKnf7_0),.din(w_dff_A_yIwuicAw7_0),.clk(gclk));
	jdff dff_A_0x4CTKnf7_0(.dout(w_dff_A_0rSnzzPj4_0),.din(w_dff_A_0x4CTKnf7_0),.clk(gclk));
	jdff dff_A_0rSnzzPj4_0(.dout(w_dff_A_a2LNhgPD4_0),.din(w_dff_A_0rSnzzPj4_0),.clk(gclk));
	jdff dff_A_a2LNhgPD4_0(.dout(w_dff_A_dqVEAAbu3_0),.din(w_dff_A_a2LNhgPD4_0),.clk(gclk));
	jdff dff_A_dqVEAAbu3_0(.dout(w_dff_A_DCuBdoDz4_0),.din(w_dff_A_dqVEAAbu3_0),.clk(gclk));
	jdff dff_A_DCuBdoDz4_0(.dout(w_dff_A_7Pu2h7lu1_0),.din(w_dff_A_DCuBdoDz4_0),.clk(gclk));
	jdff dff_A_7Pu2h7lu1_0(.dout(w_dff_A_qQnBUnhz3_0),.din(w_dff_A_7Pu2h7lu1_0),.clk(gclk));
	jdff dff_A_qQnBUnhz3_0(.dout(w_dff_A_4O8ace7l1_0),.din(w_dff_A_qQnBUnhz3_0),.clk(gclk));
	jdff dff_A_4O8ace7l1_0(.dout(w_dff_A_gyS4asOc8_0),.din(w_dff_A_4O8ace7l1_0),.clk(gclk));
	jdff dff_A_gyS4asOc8_0(.dout(w_dff_A_MJqVFwi67_0),.din(w_dff_A_gyS4asOc8_0),.clk(gclk));
	jdff dff_A_MJqVFwi67_0(.dout(w_dff_A_fFFvfhWN2_0),.din(w_dff_A_MJqVFwi67_0),.clk(gclk));
	jdff dff_A_fFFvfhWN2_0(.dout(w_dff_A_xie6wb2G0_0),.din(w_dff_A_fFFvfhWN2_0),.clk(gclk));
	jdff dff_A_xie6wb2G0_0(.dout(w_dff_A_TLjKRVch2_0),.din(w_dff_A_xie6wb2G0_0),.clk(gclk));
	jdff dff_A_TLjKRVch2_0(.dout(w_dff_A_pNp79i8V9_0),.din(w_dff_A_TLjKRVch2_0),.clk(gclk));
	jdff dff_A_pNp79i8V9_0(.dout(w_dff_A_wXRBSrFY6_0),.din(w_dff_A_pNp79i8V9_0),.clk(gclk));
	jdff dff_A_wXRBSrFY6_0(.dout(w_dff_A_3sQIG0Ov2_0),.din(w_dff_A_wXRBSrFY6_0),.clk(gclk));
	jdff dff_A_3sQIG0Ov2_0(.dout(G2548gat),.din(w_dff_A_3sQIG0Ov2_0),.clk(gclk));
	jdff dff_A_w3mHM9Py5_2(.dout(w_dff_A_JakqqeV08_0),.din(w_dff_A_w3mHM9Py5_2),.clk(gclk));
	jdff dff_A_JakqqeV08_0(.dout(w_dff_A_SesUIdQv5_0),.din(w_dff_A_JakqqeV08_0),.clk(gclk));
	jdff dff_A_SesUIdQv5_0(.dout(w_dff_A_4E6N3AQ14_0),.din(w_dff_A_SesUIdQv5_0),.clk(gclk));
	jdff dff_A_4E6N3AQ14_0(.dout(w_dff_A_zxi2NWyo2_0),.din(w_dff_A_4E6N3AQ14_0),.clk(gclk));
	jdff dff_A_zxi2NWyo2_0(.dout(w_dff_A_7xLM1DEP4_0),.din(w_dff_A_zxi2NWyo2_0),.clk(gclk));
	jdff dff_A_7xLM1DEP4_0(.dout(w_dff_A_5m0orVSO7_0),.din(w_dff_A_7xLM1DEP4_0),.clk(gclk));
	jdff dff_A_5m0orVSO7_0(.dout(w_dff_A_yIZrjeEn3_0),.din(w_dff_A_5m0orVSO7_0),.clk(gclk));
	jdff dff_A_yIZrjeEn3_0(.dout(w_dff_A_Vpdpc3n28_0),.din(w_dff_A_yIZrjeEn3_0),.clk(gclk));
	jdff dff_A_Vpdpc3n28_0(.dout(w_dff_A_42hxcsI41_0),.din(w_dff_A_Vpdpc3n28_0),.clk(gclk));
	jdff dff_A_42hxcsI41_0(.dout(w_dff_A_b867YtuE9_0),.din(w_dff_A_42hxcsI41_0),.clk(gclk));
	jdff dff_A_b867YtuE9_0(.dout(w_dff_A_S0yvhFAL4_0),.din(w_dff_A_b867YtuE9_0),.clk(gclk));
	jdff dff_A_S0yvhFAL4_0(.dout(w_dff_A_S5gYA1oS1_0),.din(w_dff_A_S0yvhFAL4_0),.clk(gclk));
	jdff dff_A_S5gYA1oS1_0(.dout(w_dff_A_IZl7vllN8_0),.din(w_dff_A_S5gYA1oS1_0),.clk(gclk));
	jdff dff_A_IZl7vllN8_0(.dout(w_dff_A_GnplEB9y1_0),.din(w_dff_A_IZl7vllN8_0),.clk(gclk));
	jdff dff_A_GnplEB9y1_0(.dout(w_dff_A_6t176Plu5_0),.din(w_dff_A_GnplEB9y1_0),.clk(gclk));
	jdff dff_A_6t176Plu5_0(.dout(w_dff_A_uPyWJ8VS5_0),.din(w_dff_A_6t176Plu5_0),.clk(gclk));
	jdff dff_A_uPyWJ8VS5_0(.dout(w_dff_A_gwWJWCzu0_0),.din(w_dff_A_uPyWJ8VS5_0),.clk(gclk));
	jdff dff_A_gwWJWCzu0_0(.dout(w_dff_A_pfsJhVjh9_0),.din(w_dff_A_gwWJWCzu0_0),.clk(gclk));
	jdff dff_A_pfsJhVjh9_0(.dout(w_dff_A_OEn9XMKV7_0),.din(w_dff_A_pfsJhVjh9_0),.clk(gclk));
	jdff dff_A_OEn9XMKV7_0(.dout(w_dff_A_hByr6STF4_0),.din(w_dff_A_OEn9XMKV7_0),.clk(gclk));
	jdff dff_A_hByr6STF4_0(.dout(w_dff_A_n4IIHgRg9_0),.din(w_dff_A_hByr6STF4_0),.clk(gclk));
	jdff dff_A_n4IIHgRg9_0(.dout(w_dff_A_XVww6zG93_0),.din(w_dff_A_n4IIHgRg9_0),.clk(gclk));
	jdff dff_A_XVww6zG93_0(.dout(w_dff_A_15Khhkqz1_0),.din(w_dff_A_XVww6zG93_0),.clk(gclk));
	jdff dff_A_15Khhkqz1_0(.dout(w_dff_A_pkr9Ey5o5_0),.din(w_dff_A_15Khhkqz1_0),.clk(gclk));
	jdff dff_A_pkr9Ey5o5_0(.dout(w_dff_A_8oemvZsB0_0),.din(w_dff_A_pkr9Ey5o5_0),.clk(gclk));
	jdff dff_A_8oemvZsB0_0(.dout(w_dff_A_tHo5P9X98_0),.din(w_dff_A_8oemvZsB0_0),.clk(gclk));
	jdff dff_A_tHo5P9X98_0(.dout(w_dff_A_1itXeHyd3_0),.din(w_dff_A_tHo5P9X98_0),.clk(gclk));
	jdff dff_A_1itXeHyd3_0(.dout(w_dff_A_B8cJIMHg6_0),.din(w_dff_A_1itXeHyd3_0),.clk(gclk));
	jdff dff_A_B8cJIMHg6_0(.dout(w_dff_A_c5FiU9ow1_0),.din(w_dff_A_B8cJIMHg6_0),.clk(gclk));
	jdff dff_A_c5FiU9ow1_0(.dout(w_dff_A_W3nfsRFu4_0),.din(w_dff_A_c5FiU9ow1_0),.clk(gclk));
	jdff dff_A_W3nfsRFu4_0(.dout(w_dff_A_EutsRKl33_0),.din(w_dff_A_W3nfsRFu4_0),.clk(gclk));
	jdff dff_A_EutsRKl33_0(.dout(w_dff_A_HqVcCpro5_0),.din(w_dff_A_EutsRKl33_0),.clk(gclk));
	jdff dff_A_HqVcCpro5_0(.dout(w_dff_A_p5cCwLaK2_0),.din(w_dff_A_HqVcCpro5_0),.clk(gclk));
	jdff dff_A_p5cCwLaK2_0(.dout(w_dff_A_TwB8fXxc6_0),.din(w_dff_A_p5cCwLaK2_0),.clk(gclk));
	jdff dff_A_TwB8fXxc6_0(.dout(w_dff_A_oe575g4w7_0),.din(w_dff_A_TwB8fXxc6_0),.clk(gclk));
	jdff dff_A_oe575g4w7_0(.dout(w_dff_A_B5eLN9NM1_0),.din(w_dff_A_oe575g4w7_0),.clk(gclk));
	jdff dff_A_B5eLN9NM1_0(.dout(w_dff_A_65Yafg4d4_0),.din(w_dff_A_B5eLN9NM1_0),.clk(gclk));
	jdff dff_A_65Yafg4d4_0(.dout(w_dff_A_DqSOxroJ5_0),.din(w_dff_A_65Yafg4d4_0),.clk(gclk));
	jdff dff_A_DqSOxroJ5_0(.dout(w_dff_A_iE3Vw3Mv5_0),.din(w_dff_A_DqSOxroJ5_0),.clk(gclk));
	jdff dff_A_iE3Vw3Mv5_0(.dout(w_dff_A_V0pYOB5p6_0),.din(w_dff_A_iE3Vw3Mv5_0),.clk(gclk));
	jdff dff_A_V0pYOB5p6_0(.dout(w_dff_A_ioLgQfr38_0),.din(w_dff_A_V0pYOB5p6_0),.clk(gclk));
	jdff dff_A_ioLgQfr38_0(.dout(w_dff_A_vE0OYVYI0_0),.din(w_dff_A_ioLgQfr38_0),.clk(gclk));
	jdff dff_A_vE0OYVYI0_0(.dout(w_dff_A_PTniF9K56_0),.din(w_dff_A_vE0OYVYI0_0),.clk(gclk));
	jdff dff_A_PTniF9K56_0(.dout(w_dff_A_Sw2QX1vV9_0),.din(w_dff_A_PTniF9K56_0),.clk(gclk));
	jdff dff_A_Sw2QX1vV9_0(.dout(w_dff_A_YMOXujyN8_0),.din(w_dff_A_Sw2QX1vV9_0),.clk(gclk));
	jdff dff_A_YMOXujyN8_0(.dout(w_dff_A_2xejjWoa4_0),.din(w_dff_A_YMOXujyN8_0),.clk(gclk));
	jdff dff_A_2xejjWoa4_0(.dout(w_dff_A_xISFREAK2_0),.din(w_dff_A_2xejjWoa4_0),.clk(gclk));
	jdff dff_A_xISFREAK2_0(.dout(w_dff_A_RiW9sP6b9_0),.din(w_dff_A_xISFREAK2_0),.clk(gclk));
	jdff dff_A_RiW9sP6b9_0(.dout(w_dff_A_Iz342MBE6_0),.din(w_dff_A_RiW9sP6b9_0),.clk(gclk));
	jdff dff_A_Iz342MBE6_0(.dout(w_dff_A_QaB235Zq1_0),.din(w_dff_A_Iz342MBE6_0),.clk(gclk));
	jdff dff_A_QaB235Zq1_0(.dout(w_dff_A_x2WhwkiH1_0),.din(w_dff_A_QaB235Zq1_0),.clk(gclk));
	jdff dff_A_x2WhwkiH1_0(.dout(w_dff_A_RAtZtlxT2_0),.din(w_dff_A_x2WhwkiH1_0),.clk(gclk));
	jdff dff_A_RAtZtlxT2_0(.dout(w_dff_A_16GcYN2g3_0),.din(w_dff_A_RAtZtlxT2_0),.clk(gclk));
	jdff dff_A_16GcYN2g3_0(.dout(w_dff_A_6FrJqOY24_0),.din(w_dff_A_16GcYN2g3_0),.clk(gclk));
	jdff dff_A_6FrJqOY24_0(.dout(w_dff_A_wNfL901z5_0),.din(w_dff_A_6FrJqOY24_0),.clk(gclk));
	jdff dff_A_wNfL901z5_0(.dout(w_dff_A_B1di4oAW9_0),.din(w_dff_A_wNfL901z5_0),.clk(gclk));
	jdff dff_A_B1di4oAW9_0(.dout(w_dff_A_tg7uLbtY4_0),.din(w_dff_A_B1di4oAW9_0),.clk(gclk));
	jdff dff_A_tg7uLbtY4_0(.dout(w_dff_A_f5r53jkt1_0),.din(w_dff_A_tg7uLbtY4_0),.clk(gclk));
	jdff dff_A_f5r53jkt1_0(.dout(w_dff_A_pDzvdEB44_0),.din(w_dff_A_f5r53jkt1_0),.clk(gclk));
	jdff dff_A_pDzvdEB44_0(.dout(G2877gat),.din(w_dff_A_pDzvdEB44_0),.clk(gclk));
	jdff dff_A_QxM6dCu23_2(.dout(w_dff_A_e01wDhmm2_0),.din(w_dff_A_QxM6dCu23_2),.clk(gclk));
	jdff dff_A_e01wDhmm2_0(.dout(w_dff_A_71V0GWoh3_0),.din(w_dff_A_e01wDhmm2_0),.clk(gclk));
	jdff dff_A_71V0GWoh3_0(.dout(w_dff_A_QP9mgEJw6_0),.din(w_dff_A_71V0GWoh3_0),.clk(gclk));
	jdff dff_A_QP9mgEJw6_0(.dout(w_dff_A_q9ky4FRJ8_0),.din(w_dff_A_QP9mgEJw6_0),.clk(gclk));
	jdff dff_A_q9ky4FRJ8_0(.dout(w_dff_A_34nH5grt4_0),.din(w_dff_A_q9ky4FRJ8_0),.clk(gclk));
	jdff dff_A_34nH5grt4_0(.dout(w_dff_A_3YMOdVJu1_0),.din(w_dff_A_34nH5grt4_0),.clk(gclk));
	jdff dff_A_3YMOdVJu1_0(.dout(w_dff_A_QsP3bsdy1_0),.din(w_dff_A_3YMOdVJu1_0),.clk(gclk));
	jdff dff_A_QsP3bsdy1_0(.dout(w_dff_A_imBaBLJ17_0),.din(w_dff_A_QsP3bsdy1_0),.clk(gclk));
	jdff dff_A_imBaBLJ17_0(.dout(w_dff_A_5mat9fLD2_0),.din(w_dff_A_imBaBLJ17_0),.clk(gclk));
	jdff dff_A_5mat9fLD2_0(.dout(w_dff_A_Txf3lufu9_0),.din(w_dff_A_5mat9fLD2_0),.clk(gclk));
	jdff dff_A_Txf3lufu9_0(.dout(w_dff_A_IFFby4vZ6_0),.din(w_dff_A_Txf3lufu9_0),.clk(gclk));
	jdff dff_A_IFFby4vZ6_0(.dout(w_dff_A_cxD9eBeh3_0),.din(w_dff_A_IFFby4vZ6_0),.clk(gclk));
	jdff dff_A_cxD9eBeh3_0(.dout(w_dff_A_6yLmLBFt0_0),.din(w_dff_A_cxD9eBeh3_0),.clk(gclk));
	jdff dff_A_6yLmLBFt0_0(.dout(w_dff_A_0Idnk2Po7_0),.din(w_dff_A_6yLmLBFt0_0),.clk(gclk));
	jdff dff_A_0Idnk2Po7_0(.dout(w_dff_A_qgxjHXtH5_0),.din(w_dff_A_0Idnk2Po7_0),.clk(gclk));
	jdff dff_A_qgxjHXtH5_0(.dout(w_dff_A_u9Cu1s053_0),.din(w_dff_A_qgxjHXtH5_0),.clk(gclk));
	jdff dff_A_u9Cu1s053_0(.dout(w_dff_A_2KA2uSxb2_0),.din(w_dff_A_u9Cu1s053_0),.clk(gclk));
	jdff dff_A_2KA2uSxb2_0(.dout(w_dff_A_eMHFlnZR8_0),.din(w_dff_A_2KA2uSxb2_0),.clk(gclk));
	jdff dff_A_eMHFlnZR8_0(.dout(w_dff_A_KwjGTL4p3_0),.din(w_dff_A_eMHFlnZR8_0),.clk(gclk));
	jdff dff_A_KwjGTL4p3_0(.dout(w_dff_A_LAPk2opK5_0),.din(w_dff_A_KwjGTL4p3_0),.clk(gclk));
	jdff dff_A_LAPk2opK5_0(.dout(w_dff_A_ihZeLB9x2_0),.din(w_dff_A_LAPk2opK5_0),.clk(gclk));
	jdff dff_A_ihZeLB9x2_0(.dout(w_dff_A_HjWGw5N04_0),.din(w_dff_A_ihZeLB9x2_0),.clk(gclk));
	jdff dff_A_HjWGw5N04_0(.dout(w_dff_A_ZOF2eZb34_0),.din(w_dff_A_HjWGw5N04_0),.clk(gclk));
	jdff dff_A_ZOF2eZb34_0(.dout(w_dff_A_NpPYNAmR8_0),.din(w_dff_A_ZOF2eZb34_0),.clk(gclk));
	jdff dff_A_NpPYNAmR8_0(.dout(w_dff_A_Jp2DZEsI4_0),.din(w_dff_A_NpPYNAmR8_0),.clk(gclk));
	jdff dff_A_Jp2DZEsI4_0(.dout(w_dff_A_ALE353iQ5_0),.din(w_dff_A_Jp2DZEsI4_0),.clk(gclk));
	jdff dff_A_ALE353iQ5_0(.dout(w_dff_A_W5LgvVxC7_0),.din(w_dff_A_ALE353iQ5_0),.clk(gclk));
	jdff dff_A_W5LgvVxC7_0(.dout(w_dff_A_KXqU0ZAF2_0),.din(w_dff_A_W5LgvVxC7_0),.clk(gclk));
	jdff dff_A_KXqU0ZAF2_0(.dout(w_dff_A_tK7Da9dN1_0),.din(w_dff_A_KXqU0ZAF2_0),.clk(gclk));
	jdff dff_A_tK7Da9dN1_0(.dout(w_dff_A_BKfJM7F47_0),.din(w_dff_A_tK7Da9dN1_0),.clk(gclk));
	jdff dff_A_BKfJM7F47_0(.dout(w_dff_A_Gt0mGzhN3_0),.din(w_dff_A_BKfJM7F47_0),.clk(gclk));
	jdff dff_A_Gt0mGzhN3_0(.dout(w_dff_A_JnAzQUn49_0),.din(w_dff_A_Gt0mGzhN3_0),.clk(gclk));
	jdff dff_A_JnAzQUn49_0(.dout(w_dff_A_i90H7wnC5_0),.din(w_dff_A_JnAzQUn49_0),.clk(gclk));
	jdff dff_A_i90H7wnC5_0(.dout(w_dff_A_txonvOJh0_0),.din(w_dff_A_i90H7wnC5_0),.clk(gclk));
	jdff dff_A_txonvOJh0_0(.dout(w_dff_A_h0Np84wX3_0),.din(w_dff_A_txonvOJh0_0),.clk(gclk));
	jdff dff_A_h0Np84wX3_0(.dout(w_dff_A_5b33Sm3G3_0),.din(w_dff_A_h0Np84wX3_0),.clk(gclk));
	jdff dff_A_5b33Sm3G3_0(.dout(w_dff_A_zsL0Qf338_0),.din(w_dff_A_5b33Sm3G3_0),.clk(gclk));
	jdff dff_A_zsL0Qf338_0(.dout(w_dff_A_ZLXs3Jm23_0),.din(w_dff_A_zsL0Qf338_0),.clk(gclk));
	jdff dff_A_ZLXs3Jm23_0(.dout(w_dff_A_b4ZMHgzr0_0),.din(w_dff_A_ZLXs3Jm23_0),.clk(gclk));
	jdff dff_A_b4ZMHgzr0_0(.dout(w_dff_A_6UvraaLu0_0),.din(w_dff_A_b4ZMHgzr0_0),.clk(gclk));
	jdff dff_A_6UvraaLu0_0(.dout(w_dff_A_x5mWSqiO5_0),.din(w_dff_A_6UvraaLu0_0),.clk(gclk));
	jdff dff_A_x5mWSqiO5_0(.dout(w_dff_A_YsUpNSSN9_0),.din(w_dff_A_x5mWSqiO5_0),.clk(gclk));
	jdff dff_A_YsUpNSSN9_0(.dout(w_dff_A_uempqmzs8_0),.din(w_dff_A_YsUpNSSN9_0),.clk(gclk));
	jdff dff_A_uempqmzs8_0(.dout(w_dff_A_S6X3TZmz0_0),.din(w_dff_A_uempqmzs8_0),.clk(gclk));
	jdff dff_A_S6X3TZmz0_0(.dout(w_dff_A_gYSrY5SC0_0),.din(w_dff_A_S6X3TZmz0_0),.clk(gclk));
	jdff dff_A_gYSrY5SC0_0(.dout(w_dff_A_zMZZJ41B4_0),.din(w_dff_A_gYSrY5SC0_0),.clk(gclk));
	jdff dff_A_zMZZJ41B4_0(.dout(w_dff_A_mYWVpp0j7_0),.din(w_dff_A_zMZZJ41B4_0),.clk(gclk));
	jdff dff_A_mYWVpp0j7_0(.dout(w_dff_A_XmsPwX095_0),.din(w_dff_A_mYWVpp0j7_0),.clk(gclk));
	jdff dff_A_XmsPwX095_0(.dout(w_dff_A_C4p2jBQJ3_0),.din(w_dff_A_XmsPwX095_0),.clk(gclk));
	jdff dff_A_C4p2jBQJ3_0(.dout(w_dff_A_eFZQk3Eh1_0),.din(w_dff_A_C4p2jBQJ3_0),.clk(gclk));
	jdff dff_A_eFZQk3Eh1_0(.dout(w_dff_A_zM5vnYCu7_0),.din(w_dff_A_eFZQk3Eh1_0),.clk(gclk));
	jdff dff_A_zM5vnYCu7_0(.dout(w_dff_A_9Nsn4WGU2_0),.din(w_dff_A_zM5vnYCu7_0),.clk(gclk));
	jdff dff_A_9Nsn4WGU2_0(.dout(w_dff_A_EeliMwh14_0),.din(w_dff_A_9Nsn4WGU2_0),.clk(gclk));
	jdff dff_A_EeliMwh14_0(.dout(w_dff_A_TGvP4lDF0_0),.din(w_dff_A_EeliMwh14_0),.clk(gclk));
	jdff dff_A_TGvP4lDF0_0(.dout(w_dff_A_ERuSPKMK5_0),.din(w_dff_A_TGvP4lDF0_0),.clk(gclk));
	jdff dff_A_ERuSPKMK5_0(.dout(w_dff_A_vYRT9OcE8_0),.din(w_dff_A_ERuSPKMK5_0),.clk(gclk));
	jdff dff_A_vYRT9OcE8_0(.dout(G3211gat),.din(w_dff_A_vYRT9OcE8_0),.clk(gclk));
	jdff dff_A_0JP3jwNj8_2(.dout(w_dff_A_9y7nuPwr7_0),.din(w_dff_A_0JP3jwNj8_2),.clk(gclk));
	jdff dff_A_9y7nuPwr7_0(.dout(w_dff_A_rwDIbwDH8_0),.din(w_dff_A_9y7nuPwr7_0),.clk(gclk));
	jdff dff_A_rwDIbwDH8_0(.dout(w_dff_A_EC2jM1kI2_0),.din(w_dff_A_rwDIbwDH8_0),.clk(gclk));
	jdff dff_A_EC2jM1kI2_0(.dout(w_dff_A_sFFvZO1G5_0),.din(w_dff_A_EC2jM1kI2_0),.clk(gclk));
	jdff dff_A_sFFvZO1G5_0(.dout(w_dff_A_o69ULqdI8_0),.din(w_dff_A_sFFvZO1G5_0),.clk(gclk));
	jdff dff_A_o69ULqdI8_0(.dout(w_dff_A_vnvzQmvE8_0),.din(w_dff_A_o69ULqdI8_0),.clk(gclk));
	jdff dff_A_vnvzQmvE8_0(.dout(w_dff_A_vPYQKSFe7_0),.din(w_dff_A_vnvzQmvE8_0),.clk(gclk));
	jdff dff_A_vPYQKSFe7_0(.dout(w_dff_A_Q3xFXEYr9_0),.din(w_dff_A_vPYQKSFe7_0),.clk(gclk));
	jdff dff_A_Q3xFXEYr9_0(.dout(w_dff_A_2p1SoVej6_0),.din(w_dff_A_Q3xFXEYr9_0),.clk(gclk));
	jdff dff_A_2p1SoVej6_0(.dout(w_dff_A_gICOUGPW3_0),.din(w_dff_A_2p1SoVej6_0),.clk(gclk));
	jdff dff_A_gICOUGPW3_0(.dout(w_dff_A_wrJOAbeg2_0),.din(w_dff_A_gICOUGPW3_0),.clk(gclk));
	jdff dff_A_wrJOAbeg2_0(.dout(w_dff_A_OZNbhE6V0_0),.din(w_dff_A_wrJOAbeg2_0),.clk(gclk));
	jdff dff_A_OZNbhE6V0_0(.dout(w_dff_A_dXbCAxYc2_0),.din(w_dff_A_OZNbhE6V0_0),.clk(gclk));
	jdff dff_A_dXbCAxYc2_0(.dout(w_dff_A_DWCE28Yg2_0),.din(w_dff_A_dXbCAxYc2_0),.clk(gclk));
	jdff dff_A_DWCE28Yg2_0(.dout(w_dff_A_ZW80NjQM6_0),.din(w_dff_A_DWCE28Yg2_0),.clk(gclk));
	jdff dff_A_ZW80NjQM6_0(.dout(w_dff_A_S5US0VGX6_0),.din(w_dff_A_ZW80NjQM6_0),.clk(gclk));
	jdff dff_A_S5US0VGX6_0(.dout(w_dff_A_dD5cbYH40_0),.din(w_dff_A_S5US0VGX6_0),.clk(gclk));
	jdff dff_A_dD5cbYH40_0(.dout(w_dff_A_8Tbz3cTc1_0),.din(w_dff_A_dD5cbYH40_0),.clk(gclk));
	jdff dff_A_8Tbz3cTc1_0(.dout(w_dff_A_gAAIlYDy1_0),.din(w_dff_A_8Tbz3cTc1_0),.clk(gclk));
	jdff dff_A_gAAIlYDy1_0(.dout(w_dff_A_aVN2lUok7_0),.din(w_dff_A_gAAIlYDy1_0),.clk(gclk));
	jdff dff_A_aVN2lUok7_0(.dout(w_dff_A_EZkZivps6_0),.din(w_dff_A_aVN2lUok7_0),.clk(gclk));
	jdff dff_A_EZkZivps6_0(.dout(w_dff_A_Z6qNvanW8_0),.din(w_dff_A_EZkZivps6_0),.clk(gclk));
	jdff dff_A_Z6qNvanW8_0(.dout(w_dff_A_YosXUhTH6_0),.din(w_dff_A_Z6qNvanW8_0),.clk(gclk));
	jdff dff_A_YosXUhTH6_0(.dout(w_dff_A_SCZnhn4U6_0),.din(w_dff_A_YosXUhTH6_0),.clk(gclk));
	jdff dff_A_SCZnhn4U6_0(.dout(w_dff_A_QCZh84Pu6_0),.din(w_dff_A_SCZnhn4U6_0),.clk(gclk));
	jdff dff_A_QCZh84Pu6_0(.dout(w_dff_A_tmlCZHY94_0),.din(w_dff_A_QCZh84Pu6_0),.clk(gclk));
	jdff dff_A_tmlCZHY94_0(.dout(w_dff_A_UIsUUhaR9_0),.din(w_dff_A_tmlCZHY94_0),.clk(gclk));
	jdff dff_A_UIsUUhaR9_0(.dout(w_dff_A_N9aQ43IP4_0),.din(w_dff_A_UIsUUhaR9_0),.clk(gclk));
	jdff dff_A_N9aQ43IP4_0(.dout(w_dff_A_wU9Lxyep3_0),.din(w_dff_A_N9aQ43IP4_0),.clk(gclk));
	jdff dff_A_wU9Lxyep3_0(.dout(w_dff_A_c0efwtBe5_0),.din(w_dff_A_wU9Lxyep3_0),.clk(gclk));
	jdff dff_A_c0efwtBe5_0(.dout(w_dff_A_8SbIfut79_0),.din(w_dff_A_c0efwtBe5_0),.clk(gclk));
	jdff dff_A_8SbIfut79_0(.dout(w_dff_A_tr4GEd7E8_0),.din(w_dff_A_8SbIfut79_0),.clk(gclk));
	jdff dff_A_tr4GEd7E8_0(.dout(w_dff_A_x9Ksuv9a4_0),.din(w_dff_A_tr4GEd7E8_0),.clk(gclk));
	jdff dff_A_x9Ksuv9a4_0(.dout(w_dff_A_fKGrflfG7_0),.din(w_dff_A_x9Ksuv9a4_0),.clk(gclk));
	jdff dff_A_fKGrflfG7_0(.dout(w_dff_A_2FXSAPhw0_0),.din(w_dff_A_fKGrflfG7_0),.clk(gclk));
	jdff dff_A_2FXSAPhw0_0(.dout(w_dff_A_8fEcePn13_0),.din(w_dff_A_2FXSAPhw0_0),.clk(gclk));
	jdff dff_A_8fEcePn13_0(.dout(w_dff_A_dZ2Or8Zg3_0),.din(w_dff_A_8fEcePn13_0),.clk(gclk));
	jdff dff_A_dZ2Or8Zg3_0(.dout(w_dff_A_PicvuRuG1_0),.din(w_dff_A_dZ2Or8Zg3_0),.clk(gclk));
	jdff dff_A_PicvuRuG1_0(.dout(w_dff_A_8kdxz9Ch5_0),.din(w_dff_A_PicvuRuG1_0),.clk(gclk));
	jdff dff_A_8kdxz9Ch5_0(.dout(w_dff_A_JTlG9CDe6_0),.din(w_dff_A_8kdxz9Ch5_0),.clk(gclk));
	jdff dff_A_JTlG9CDe6_0(.dout(w_dff_A_nuB0GE4r1_0),.din(w_dff_A_JTlG9CDe6_0),.clk(gclk));
	jdff dff_A_nuB0GE4r1_0(.dout(w_dff_A_MR2XgASb7_0),.din(w_dff_A_nuB0GE4r1_0),.clk(gclk));
	jdff dff_A_MR2XgASb7_0(.dout(w_dff_A_tFWlQKnh6_0),.din(w_dff_A_MR2XgASb7_0),.clk(gclk));
	jdff dff_A_tFWlQKnh6_0(.dout(w_dff_A_bhnfYepS4_0),.din(w_dff_A_tFWlQKnh6_0),.clk(gclk));
	jdff dff_A_bhnfYepS4_0(.dout(w_dff_A_S9bBKKld1_0),.din(w_dff_A_bhnfYepS4_0),.clk(gclk));
	jdff dff_A_S9bBKKld1_0(.dout(w_dff_A_cHdYMAfi8_0),.din(w_dff_A_S9bBKKld1_0),.clk(gclk));
	jdff dff_A_cHdYMAfi8_0(.dout(w_dff_A_r9Nlqm7i4_0),.din(w_dff_A_cHdYMAfi8_0),.clk(gclk));
	jdff dff_A_r9Nlqm7i4_0(.dout(w_dff_A_XkHpznFV3_0),.din(w_dff_A_r9Nlqm7i4_0),.clk(gclk));
	jdff dff_A_XkHpznFV3_0(.dout(w_dff_A_CyXriHxa6_0),.din(w_dff_A_XkHpznFV3_0),.clk(gclk));
	jdff dff_A_CyXriHxa6_0(.dout(w_dff_A_GmIQqCmU1_0),.din(w_dff_A_CyXriHxa6_0),.clk(gclk));
	jdff dff_A_GmIQqCmU1_0(.dout(w_dff_A_W06CTYbN9_0),.din(w_dff_A_GmIQqCmU1_0),.clk(gclk));
	jdff dff_A_W06CTYbN9_0(.dout(w_dff_A_S5MkaSO17_0),.din(w_dff_A_W06CTYbN9_0),.clk(gclk));
	jdff dff_A_S5MkaSO17_0(.dout(w_dff_A_l4fMSMGb2_0),.din(w_dff_A_S5MkaSO17_0),.clk(gclk));
	jdff dff_A_l4fMSMGb2_0(.dout(G3552gat),.din(w_dff_A_l4fMSMGb2_0),.clk(gclk));
	jdff dff_A_tDHTbtHD9_2(.dout(w_dff_A_q8aFmGwZ4_0),.din(w_dff_A_tDHTbtHD9_2),.clk(gclk));
	jdff dff_A_q8aFmGwZ4_0(.dout(w_dff_A_A0jCiuli4_0),.din(w_dff_A_q8aFmGwZ4_0),.clk(gclk));
	jdff dff_A_A0jCiuli4_0(.dout(w_dff_A_h6HUAdhD6_0),.din(w_dff_A_A0jCiuli4_0),.clk(gclk));
	jdff dff_A_h6HUAdhD6_0(.dout(w_dff_A_yNxj5BwM7_0),.din(w_dff_A_h6HUAdhD6_0),.clk(gclk));
	jdff dff_A_yNxj5BwM7_0(.dout(w_dff_A_p7RJdatl3_0),.din(w_dff_A_yNxj5BwM7_0),.clk(gclk));
	jdff dff_A_p7RJdatl3_0(.dout(w_dff_A_CiDFMdkw8_0),.din(w_dff_A_p7RJdatl3_0),.clk(gclk));
	jdff dff_A_CiDFMdkw8_0(.dout(w_dff_A_ofCcrgmp4_0),.din(w_dff_A_CiDFMdkw8_0),.clk(gclk));
	jdff dff_A_ofCcrgmp4_0(.dout(w_dff_A_Xo7ZIekS3_0),.din(w_dff_A_ofCcrgmp4_0),.clk(gclk));
	jdff dff_A_Xo7ZIekS3_0(.dout(w_dff_A_RpFuB8Qn1_0),.din(w_dff_A_Xo7ZIekS3_0),.clk(gclk));
	jdff dff_A_RpFuB8Qn1_0(.dout(w_dff_A_14TbbzkY5_0),.din(w_dff_A_RpFuB8Qn1_0),.clk(gclk));
	jdff dff_A_14TbbzkY5_0(.dout(w_dff_A_uXxcj9tz7_0),.din(w_dff_A_14TbbzkY5_0),.clk(gclk));
	jdff dff_A_uXxcj9tz7_0(.dout(w_dff_A_BHFk1Yzt1_0),.din(w_dff_A_uXxcj9tz7_0),.clk(gclk));
	jdff dff_A_BHFk1Yzt1_0(.dout(w_dff_A_50bpTB1X7_0),.din(w_dff_A_BHFk1Yzt1_0),.clk(gclk));
	jdff dff_A_50bpTB1X7_0(.dout(w_dff_A_dIi3DsUF7_0),.din(w_dff_A_50bpTB1X7_0),.clk(gclk));
	jdff dff_A_dIi3DsUF7_0(.dout(w_dff_A_upeYc7wD8_0),.din(w_dff_A_dIi3DsUF7_0),.clk(gclk));
	jdff dff_A_upeYc7wD8_0(.dout(w_dff_A_5Ld78PMj9_0),.din(w_dff_A_upeYc7wD8_0),.clk(gclk));
	jdff dff_A_5Ld78PMj9_0(.dout(w_dff_A_SSt2Kutn2_0),.din(w_dff_A_5Ld78PMj9_0),.clk(gclk));
	jdff dff_A_SSt2Kutn2_0(.dout(w_dff_A_gDbYxs4x9_0),.din(w_dff_A_SSt2Kutn2_0),.clk(gclk));
	jdff dff_A_gDbYxs4x9_0(.dout(w_dff_A_uYgVlVl84_0),.din(w_dff_A_gDbYxs4x9_0),.clk(gclk));
	jdff dff_A_uYgVlVl84_0(.dout(w_dff_A_j2ctZomr5_0),.din(w_dff_A_uYgVlVl84_0),.clk(gclk));
	jdff dff_A_j2ctZomr5_0(.dout(w_dff_A_ZxJillTQ5_0),.din(w_dff_A_j2ctZomr5_0),.clk(gclk));
	jdff dff_A_ZxJillTQ5_0(.dout(w_dff_A_QJVAZTCR0_0),.din(w_dff_A_ZxJillTQ5_0),.clk(gclk));
	jdff dff_A_QJVAZTCR0_0(.dout(w_dff_A_tvh4sAEC5_0),.din(w_dff_A_QJVAZTCR0_0),.clk(gclk));
	jdff dff_A_tvh4sAEC5_0(.dout(w_dff_A_bKZ7AmGt4_0),.din(w_dff_A_tvh4sAEC5_0),.clk(gclk));
	jdff dff_A_bKZ7AmGt4_0(.dout(w_dff_A_U9GbU6Fx4_0),.din(w_dff_A_bKZ7AmGt4_0),.clk(gclk));
	jdff dff_A_U9GbU6Fx4_0(.dout(w_dff_A_GbUPDE3q6_0),.din(w_dff_A_U9GbU6Fx4_0),.clk(gclk));
	jdff dff_A_GbUPDE3q6_0(.dout(w_dff_A_QiHzXXPs8_0),.din(w_dff_A_GbUPDE3q6_0),.clk(gclk));
	jdff dff_A_QiHzXXPs8_0(.dout(w_dff_A_noWrcSJX8_0),.din(w_dff_A_QiHzXXPs8_0),.clk(gclk));
	jdff dff_A_noWrcSJX8_0(.dout(w_dff_A_3XzaxxNv0_0),.din(w_dff_A_noWrcSJX8_0),.clk(gclk));
	jdff dff_A_3XzaxxNv0_0(.dout(w_dff_A_3uePTLzI7_0),.din(w_dff_A_3XzaxxNv0_0),.clk(gclk));
	jdff dff_A_3uePTLzI7_0(.dout(w_dff_A_rzlm0Y8B9_0),.din(w_dff_A_3uePTLzI7_0),.clk(gclk));
	jdff dff_A_rzlm0Y8B9_0(.dout(w_dff_A_SdU8bPRz6_0),.din(w_dff_A_rzlm0Y8B9_0),.clk(gclk));
	jdff dff_A_SdU8bPRz6_0(.dout(w_dff_A_9gdr0Xiz7_0),.din(w_dff_A_SdU8bPRz6_0),.clk(gclk));
	jdff dff_A_9gdr0Xiz7_0(.dout(w_dff_A_R08VmBP44_0),.din(w_dff_A_9gdr0Xiz7_0),.clk(gclk));
	jdff dff_A_R08VmBP44_0(.dout(w_dff_A_Ik9SmEod2_0),.din(w_dff_A_R08VmBP44_0),.clk(gclk));
	jdff dff_A_Ik9SmEod2_0(.dout(w_dff_A_rUGlc7xG3_0),.din(w_dff_A_Ik9SmEod2_0),.clk(gclk));
	jdff dff_A_rUGlc7xG3_0(.dout(w_dff_A_NE0Xxvtv7_0),.din(w_dff_A_rUGlc7xG3_0),.clk(gclk));
	jdff dff_A_NE0Xxvtv7_0(.dout(w_dff_A_agiBJQfc9_0),.din(w_dff_A_NE0Xxvtv7_0),.clk(gclk));
	jdff dff_A_agiBJQfc9_0(.dout(w_dff_A_5OTMzzmz6_0),.din(w_dff_A_agiBJQfc9_0),.clk(gclk));
	jdff dff_A_5OTMzzmz6_0(.dout(w_dff_A_Pj0pm2Lm9_0),.din(w_dff_A_5OTMzzmz6_0),.clk(gclk));
	jdff dff_A_Pj0pm2Lm9_0(.dout(w_dff_A_3VPgA6oT7_0),.din(w_dff_A_Pj0pm2Lm9_0),.clk(gclk));
	jdff dff_A_3VPgA6oT7_0(.dout(w_dff_A_UU2TEuBj0_0),.din(w_dff_A_3VPgA6oT7_0),.clk(gclk));
	jdff dff_A_UU2TEuBj0_0(.dout(w_dff_A_P125C3pf9_0),.din(w_dff_A_UU2TEuBj0_0),.clk(gclk));
	jdff dff_A_P125C3pf9_0(.dout(w_dff_A_XFrQZNcg6_0),.din(w_dff_A_P125C3pf9_0),.clk(gclk));
	jdff dff_A_XFrQZNcg6_0(.dout(w_dff_A_emcMfYOC1_0),.din(w_dff_A_XFrQZNcg6_0),.clk(gclk));
	jdff dff_A_emcMfYOC1_0(.dout(w_dff_A_eq14Vo006_0),.din(w_dff_A_emcMfYOC1_0),.clk(gclk));
	jdff dff_A_eq14Vo006_0(.dout(w_dff_A_nGM6iWhg4_0),.din(w_dff_A_eq14Vo006_0),.clk(gclk));
	jdff dff_A_nGM6iWhg4_0(.dout(w_dff_A_0Tuq0Iiq2_0),.din(w_dff_A_nGM6iWhg4_0),.clk(gclk));
	jdff dff_A_0Tuq0Iiq2_0(.dout(w_dff_A_FDDth7LC2_0),.din(w_dff_A_0Tuq0Iiq2_0),.clk(gclk));
	jdff dff_A_FDDth7LC2_0(.dout(w_dff_A_YVygEv5j9_0),.din(w_dff_A_FDDth7LC2_0),.clk(gclk));
	jdff dff_A_YVygEv5j9_0(.dout(G3895gat),.din(w_dff_A_YVygEv5j9_0),.clk(gclk));
	jdff dff_A_yY8yxN6c1_2(.dout(w_dff_A_0b1wWLal0_0),.din(w_dff_A_yY8yxN6c1_2),.clk(gclk));
	jdff dff_A_0b1wWLal0_0(.dout(w_dff_A_9v1dS7BS6_0),.din(w_dff_A_0b1wWLal0_0),.clk(gclk));
	jdff dff_A_9v1dS7BS6_0(.dout(w_dff_A_vM9hfPwR7_0),.din(w_dff_A_9v1dS7BS6_0),.clk(gclk));
	jdff dff_A_vM9hfPwR7_0(.dout(w_dff_A_vwnSNPbd6_0),.din(w_dff_A_vM9hfPwR7_0),.clk(gclk));
	jdff dff_A_vwnSNPbd6_0(.dout(w_dff_A_t7Nr2H954_0),.din(w_dff_A_vwnSNPbd6_0),.clk(gclk));
	jdff dff_A_t7Nr2H954_0(.dout(w_dff_A_PRPqvJq75_0),.din(w_dff_A_t7Nr2H954_0),.clk(gclk));
	jdff dff_A_PRPqvJq75_0(.dout(w_dff_A_P8lKd5Ei4_0),.din(w_dff_A_PRPqvJq75_0),.clk(gclk));
	jdff dff_A_P8lKd5Ei4_0(.dout(w_dff_A_nClFaeR25_0),.din(w_dff_A_P8lKd5Ei4_0),.clk(gclk));
	jdff dff_A_nClFaeR25_0(.dout(w_dff_A_7OdD3DtH2_0),.din(w_dff_A_nClFaeR25_0),.clk(gclk));
	jdff dff_A_7OdD3DtH2_0(.dout(w_dff_A_i96Tcl8H9_0),.din(w_dff_A_7OdD3DtH2_0),.clk(gclk));
	jdff dff_A_i96Tcl8H9_0(.dout(w_dff_A_z53VELXU9_0),.din(w_dff_A_i96Tcl8H9_0),.clk(gclk));
	jdff dff_A_z53VELXU9_0(.dout(w_dff_A_JG4tHwD50_0),.din(w_dff_A_z53VELXU9_0),.clk(gclk));
	jdff dff_A_JG4tHwD50_0(.dout(w_dff_A_TB75Yj5y7_0),.din(w_dff_A_JG4tHwD50_0),.clk(gclk));
	jdff dff_A_TB75Yj5y7_0(.dout(w_dff_A_fCfZubvv1_0),.din(w_dff_A_TB75Yj5y7_0),.clk(gclk));
	jdff dff_A_fCfZubvv1_0(.dout(w_dff_A_1Sdie3if2_0),.din(w_dff_A_fCfZubvv1_0),.clk(gclk));
	jdff dff_A_1Sdie3if2_0(.dout(w_dff_A_lkQwCQPJ1_0),.din(w_dff_A_1Sdie3if2_0),.clk(gclk));
	jdff dff_A_lkQwCQPJ1_0(.dout(w_dff_A_j3Ohi46O8_0),.din(w_dff_A_lkQwCQPJ1_0),.clk(gclk));
	jdff dff_A_j3Ohi46O8_0(.dout(w_dff_A_UIP0i0cf1_0),.din(w_dff_A_j3Ohi46O8_0),.clk(gclk));
	jdff dff_A_UIP0i0cf1_0(.dout(w_dff_A_fmR0BYtz3_0),.din(w_dff_A_UIP0i0cf1_0),.clk(gclk));
	jdff dff_A_fmR0BYtz3_0(.dout(w_dff_A_of14nbZc5_0),.din(w_dff_A_fmR0BYtz3_0),.clk(gclk));
	jdff dff_A_of14nbZc5_0(.dout(w_dff_A_gAnzB6kQ3_0),.din(w_dff_A_of14nbZc5_0),.clk(gclk));
	jdff dff_A_gAnzB6kQ3_0(.dout(w_dff_A_brmmQzJT5_0),.din(w_dff_A_gAnzB6kQ3_0),.clk(gclk));
	jdff dff_A_brmmQzJT5_0(.dout(w_dff_A_NkbS25FG6_0),.din(w_dff_A_brmmQzJT5_0),.clk(gclk));
	jdff dff_A_NkbS25FG6_0(.dout(w_dff_A_rw3kTQKb0_0),.din(w_dff_A_NkbS25FG6_0),.clk(gclk));
	jdff dff_A_rw3kTQKb0_0(.dout(w_dff_A_40WdcH1w2_0),.din(w_dff_A_rw3kTQKb0_0),.clk(gclk));
	jdff dff_A_40WdcH1w2_0(.dout(w_dff_A_7BYduC8C8_0),.din(w_dff_A_40WdcH1w2_0),.clk(gclk));
	jdff dff_A_7BYduC8C8_0(.dout(w_dff_A_NeIWGPHg2_0),.din(w_dff_A_7BYduC8C8_0),.clk(gclk));
	jdff dff_A_NeIWGPHg2_0(.dout(w_dff_A_u7aqd18z4_0),.din(w_dff_A_NeIWGPHg2_0),.clk(gclk));
	jdff dff_A_u7aqd18z4_0(.dout(w_dff_A_G4ZC9E6f8_0),.din(w_dff_A_u7aqd18z4_0),.clk(gclk));
	jdff dff_A_G4ZC9E6f8_0(.dout(w_dff_A_9k9HSoWQ7_0),.din(w_dff_A_G4ZC9E6f8_0),.clk(gclk));
	jdff dff_A_9k9HSoWQ7_0(.dout(w_dff_A_1XGm5JsJ0_0),.din(w_dff_A_9k9HSoWQ7_0),.clk(gclk));
	jdff dff_A_1XGm5JsJ0_0(.dout(w_dff_A_EJ1X0jFs0_0),.din(w_dff_A_1XGm5JsJ0_0),.clk(gclk));
	jdff dff_A_EJ1X0jFs0_0(.dout(w_dff_A_YJ7iCCNq3_0),.din(w_dff_A_EJ1X0jFs0_0),.clk(gclk));
	jdff dff_A_YJ7iCCNq3_0(.dout(w_dff_A_gLNRFF4J1_0),.din(w_dff_A_YJ7iCCNq3_0),.clk(gclk));
	jdff dff_A_gLNRFF4J1_0(.dout(w_dff_A_mPZgSX809_0),.din(w_dff_A_gLNRFF4J1_0),.clk(gclk));
	jdff dff_A_mPZgSX809_0(.dout(w_dff_A_NnglkXpB4_0),.din(w_dff_A_mPZgSX809_0),.clk(gclk));
	jdff dff_A_NnglkXpB4_0(.dout(w_dff_A_B8fArUQK7_0),.din(w_dff_A_NnglkXpB4_0),.clk(gclk));
	jdff dff_A_B8fArUQK7_0(.dout(w_dff_A_CVW4O55p7_0),.din(w_dff_A_B8fArUQK7_0),.clk(gclk));
	jdff dff_A_CVW4O55p7_0(.dout(w_dff_A_RCwCBnkA9_0),.din(w_dff_A_CVW4O55p7_0),.clk(gclk));
	jdff dff_A_RCwCBnkA9_0(.dout(w_dff_A_E33sluXJ1_0),.din(w_dff_A_RCwCBnkA9_0),.clk(gclk));
	jdff dff_A_E33sluXJ1_0(.dout(w_dff_A_FnVM3lPo6_0),.din(w_dff_A_E33sluXJ1_0),.clk(gclk));
	jdff dff_A_FnVM3lPo6_0(.dout(w_dff_A_1J2KOAl32_0),.din(w_dff_A_FnVM3lPo6_0),.clk(gclk));
	jdff dff_A_1J2KOAl32_0(.dout(w_dff_A_R6MIg0XX3_0),.din(w_dff_A_1J2KOAl32_0),.clk(gclk));
	jdff dff_A_R6MIg0XX3_0(.dout(w_dff_A_aL2jgIDE2_0),.din(w_dff_A_R6MIg0XX3_0),.clk(gclk));
	jdff dff_A_aL2jgIDE2_0(.dout(w_dff_A_i1Q5XMKk5_0),.din(w_dff_A_aL2jgIDE2_0),.clk(gclk));
	jdff dff_A_i1Q5XMKk5_0(.dout(w_dff_A_Q36wvf1V6_0),.din(w_dff_A_i1Q5XMKk5_0),.clk(gclk));
	jdff dff_A_Q36wvf1V6_0(.dout(w_dff_A_BsgY16DA7_0),.din(w_dff_A_Q36wvf1V6_0),.clk(gclk));
	jdff dff_A_BsgY16DA7_0(.dout(G4241gat),.din(w_dff_A_BsgY16DA7_0),.clk(gclk));
	jdff dff_A_fbgsIzQB8_2(.dout(w_dff_A_qNCNU8F57_0),.din(w_dff_A_fbgsIzQB8_2),.clk(gclk));
	jdff dff_A_qNCNU8F57_0(.dout(w_dff_A_rfKRqyHU1_0),.din(w_dff_A_qNCNU8F57_0),.clk(gclk));
	jdff dff_A_rfKRqyHU1_0(.dout(w_dff_A_ovHxfjTD4_0),.din(w_dff_A_rfKRqyHU1_0),.clk(gclk));
	jdff dff_A_ovHxfjTD4_0(.dout(w_dff_A_OX1r2rZU1_0),.din(w_dff_A_ovHxfjTD4_0),.clk(gclk));
	jdff dff_A_OX1r2rZU1_0(.dout(w_dff_A_L5drJ2ae2_0),.din(w_dff_A_OX1r2rZU1_0),.clk(gclk));
	jdff dff_A_L5drJ2ae2_0(.dout(w_dff_A_bARdbM5a4_0),.din(w_dff_A_L5drJ2ae2_0),.clk(gclk));
	jdff dff_A_bARdbM5a4_0(.dout(w_dff_A_AuZTwuwb0_0),.din(w_dff_A_bARdbM5a4_0),.clk(gclk));
	jdff dff_A_AuZTwuwb0_0(.dout(w_dff_A_VA6UYDbr0_0),.din(w_dff_A_AuZTwuwb0_0),.clk(gclk));
	jdff dff_A_VA6UYDbr0_0(.dout(w_dff_A_nb2VvcMG1_0),.din(w_dff_A_VA6UYDbr0_0),.clk(gclk));
	jdff dff_A_nb2VvcMG1_0(.dout(w_dff_A_MePFNjtP3_0),.din(w_dff_A_nb2VvcMG1_0),.clk(gclk));
	jdff dff_A_MePFNjtP3_0(.dout(w_dff_A_ZiV2sNfm9_0),.din(w_dff_A_MePFNjtP3_0),.clk(gclk));
	jdff dff_A_ZiV2sNfm9_0(.dout(w_dff_A_q45HJ2GB2_0),.din(w_dff_A_ZiV2sNfm9_0),.clk(gclk));
	jdff dff_A_q45HJ2GB2_0(.dout(w_dff_A_CZP3qcSt4_0),.din(w_dff_A_q45HJ2GB2_0),.clk(gclk));
	jdff dff_A_CZP3qcSt4_0(.dout(w_dff_A_DS6MY5VM5_0),.din(w_dff_A_CZP3qcSt4_0),.clk(gclk));
	jdff dff_A_DS6MY5VM5_0(.dout(w_dff_A_DdPtjZeI8_0),.din(w_dff_A_DS6MY5VM5_0),.clk(gclk));
	jdff dff_A_DdPtjZeI8_0(.dout(w_dff_A_pFyblxKc4_0),.din(w_dff_A_DdPtjZeI8_0),.clk(gclk));
	jdff dff_A_pFyblxKc4_0(.dout(w_dff_A_f9CFv9jU8_0),.din(w_dff_A_pFyblxKc4_0),.clk(gclk));
	jdff dff_A_f9CFv9jU8_0(.dout(w_dff_A_asFNwthJ7_0),.din(w_dff_A_f9CFv9jU8_0),.clk(gclk));
	jdff dff_A_asFNwthJ7_0(.dout(w_dff_A_W6Apw8iQ4_0),.din(w_dff_A_asFNwthJ7_0),.clk(gclk));
	jdff dff_A_W6Apw8iQ4_0(.dout(w_dff_A_oFLy3QE49_0),.din(w_dff_A_W6Apw8iQ4_0),.clk(gclk));
	jdff dff_A_oFLy3QE49_0(.dout(w_dff_A_9HvlsRXd7_0),.din(w_dff_A_oFLy3QE49_0),.clk(gclk));
	jdff dff_A_9HvlsRXd7_0(.dout(w_dff_A_fYfG2ma35_0),.din(w_dff_A_9HvlsRXd7_0),.clk(gclk));
	jdff dff_A_fYfG2ma35_0(.dout(w_dff_A_SelniTRZ8_0),.din(w_dff_A_fYfG2ma35_0),.clk(gclk));
	jdff dff_A_SelniTRZ8_0(.dout(w_dff_A_rV80BmMk3_0),.din(w_dff_A_SelniTRZ8_0),.clk(gclk));
	jdff dff_A_rV80BmMk3_0(.dout(w_dff_A_qLroIxiw2_0),.din(w_dff_A_rV80BmMk3_0),.clk(gclk));
	jdff dff_A_qLroIxiw2_0(.dout(w_dff_A_a85xfeTt2_0),.din(w_dff_A_qLroIxiw2_0),.clk(gclk));
	jdff dff_A_a85xfeTt2_0(.dout(w_dff_A_jGDSUmUd3_0),.din(w_dff_A_a85xfeTt2_0),.clk(gclk));
	jdff dff_A_jGDSUmUd3_0(.dout(w_dff_A_eOOedJWz2_0),.din(w_dff_A_jGDSUmUd3_0),.clk(gclk));
	jdff dff_A_eOOedJWz2_0(.dout(w_dff_A_uDRtnHPv0_0),.din(w_dff_A_eOOedJWz2_0),.clk(gclk));
	jdff dff_A_uDRtnHPv0_0(.dout(w_dff_A_oxMhZN4T2_0),.din(w_dff_A_uDRtnHPv0_0),.clk(gclk));
	jdff dff_A_oxMhZN4T2_0(.dout(w_dff_A_ESxJ4YV42_0),.din(w_dff_A_oxMhZN4T2_0),.clk(gclk));
	jdff dff_A_ESxJ4YV42_0(.dout(w_dff_A_paPIw30Y4_0),.din(w_dff_A_ESxJ4YV42_0),.clk(gclk));
	jdff dff_A_paPIw30Y4_0(.dout(w_dff_A_qLEpEyQN5_0),.din(w_dff_A_paPIw30Y4_0),.clk(gclk));
	jdff dff_A_qLEpEyQN5_0(.dout(w_dff_A_qVyleftZ2_0),.din(w_dff_A_qLEpEyQN5_0),.clk(gclk));
	jdff dff_A_qVyleftZ2_0(.dout(w_dff_A_4foWbfZS4_0),.din(w_dff_A_qVyleftZ2_0),.clk(gclk));
	jdff dff_A_4foWbfZS4_0(.dout(w_dff_A_xKh5cuOz4_0),.din(w_dff_A_4foWbfZS4_0),.clk(gclk));
	jdff dff_A_xKh5cuOz4_0(.dout(w_dff_A_RmSzaXQB6_0),.din(w_dff_A_xKh5cuOz4_0),.clk(gclk));
	jdff dff_A_RmSzaXQB6_0(.dout(w_dff_A_0MObwkrQ2_0),.din(w_dff_A_RmSzaXQB6_0),.clk(gclk));
	jdff dff_A_0MObwkrQ2_0(.dout(w_dff_A_fgKlhONG3_0),.din(w_dff_A_0MObwkrQ2_0),.clk(gclk));
	jdff dff_A_fgKlhONG3_0(.dout(w_dff_A_7V7YIKOI2_0),.din(w_dff_A_fgKlhONG3_0),.clk(gclk));
	jdff dff_A_7V7YIKOI2_0(.dout(w_dff_A_bswxh8ik4_0),.din(w_dff_A_7V7YIKOI2_0),.clk(gclk));
	jdff dff_A_bswxh8ik4_0(.dout(w_dff_A_6frSAAOX8_0),.din(w_dff_A_bswxh8ik4_0),.clk(gclk));
	jdff dff_A_6frSAAOX8_0(.dout(w_dff_A_T8XkDwd88_0),.din(w_dff_A_6frSAAOX8_0),.clk(gclk));
	jdff dff_A_T8XkDwd88_0(.dout(w_dff_A_8pOYho5g0_0),.din(w_dff_A_T8XkDwd88_0),.clk(gclk));
	jdff dff_A_8pOYho5g0_0(.dout(G4591gat),.din(w_dff_A_8pOYho5g0_0),.clk(gclk));
	jdff dff_A_DQUJXFRm8_2(.dout(w_dff_A_JFTtzcUb4_0),.din(w_dff_A_DQUJXFRm8_2),.clk(gclk));
	jdff dff_A_JFTtzcUb4_0(.dout(w_dff_A_HFjeRtC20_0),.din(w_dff_A_JFTtzcUb4_0),.clk(gclk));
	jdff dff_A_HFjeRtC20_0(.dout(w_dff_A_wD8F8hqE4_0),.din(w_dff_A_HFjeRtC20_0),.clk(gclk));
	jdff dff_A_wD8F8hqE4_0(.dout(w_dff_A_wVjVJ9ib8_0),.din(w_dff_A_wD8F8hqE4_0),.clk(gclk));
	jdff dff_A_wVjVJ9ib8_0(.dout(w_dff_A_7GWRsU4V5_0),.din(w_dff_A_wVjVJ9ib8_0),.clk(gclk));
	jdff dff_A_7GWRsU4V5_0(.dout(w_dff_A_beufR2cX8_0),.din(w_dff_A_7GWRsU4V5_0),.clk(gclk));
	jdff dff_A_beufR2cX8_0(.dout(w_dff_A_9gbRHc2e8_0),.din(w_dff_A_beufR2cX8_0),.clk(gclk));
	jdff dff_A_9gbRHc2e8_0(.dout(w_dff_A_M5tnwTok7_0),.din(w_dff_A_9gbRHc2e8_0),.clk(gclk));
	jdff dff_A_M5tnwTok7_0(.dout(w_dff_A_dysjJHkp7_0),.din(w_dff_A_M5tnwTok7_0),.clk(gclk));
	jdff dff_A_dysjJHkp7_0(.dout(w_dff_A_5lTRNEKv6_0),.din(w_dff_A_dysjJHkp7_0),.clk(gclk));
	jdff dff_A_5lTRNEKv6_0(.dout(w_dff_A_fkkSoLPu0_0),.din(w_dff_A_5lTRNEKv6_0),.clk(gclk));
	jdff dff_A_fkkSoLPu0_0(.dout(w_dff_A_VTBh2ZbQ4_0),.din(w_dff_A_fkkSoLPu0_0),.clk(gclk));
	jdff dff_A_VTBh2ZbQ4_0(.dout(w_dff_A_61uc9PD59_0),.din(w_dff_A_VTBh2ZbQ4_0),.clk(gclk));
	jdff dff_A_61uc9PD59_0(.dout(w_dff_A_bWdrDN9S0_0),.din(w_dff_A_61uc9PD59_0),.clk(gclk));
	jdff dff_A_bWdrDN9S0_0(.dout(w_dff_A_F3zsr08B1_0),.din(w_dff_A_bWdrDN9S0_0),.clk(gclk));
	jdff dff_A_F3zsr08B1_0(.dout(w_dff_A_UjKGELjN8_0),.din(w_dff_A_F3zsr08B1_0),.clk(gclk));
	jdff dff_A_UjKGELjN8_0(.dout(w_dff_A_M23keRjl5_0),.din(w_dff_A_UjKGELjN8_0),.clk(gclk));
	jdff dff_A_M23keRjl5_0(.dout(w_dff_A_H2Ro9ix14_0),.din(w_dff_A_M23keRjl5_0),.clk(gclk));
	jdff dff_A_H2Ro9ix14_0(.dout(w_dff_A_WAHmXhtO6_0),.din(w_dff_A_H2Ro9ix14_0),.clk(gclk));
	jdff dff_A_WAHmXhtO6_0(.dout(w_dff_A_QKKsJc3r3_0),.din(w_dff_A_WAHmXhtO6_0),.clk(gclk));
	jdff dff_A_QKKsJc3r3_0(.dout(w_dff_A_hF66G8km0_0),.din(w_dff_A_QKKsJc3r3_0),.clk(gclk));
	jdff dff_A_hF66G8km0_0(.dout(w_dff_A_Wlx5e4gI1_0),.din(w_dff_A_hF66G8km0_0),.clk(gclk));
	jdff dff_A_Wlx5e4gI1_0(.dout(w_dff_A_L8ZrONbv7_0),.din(w_dff_A_Wlx5e4gI1_0),.clk(gclk));
	jdff dff_A_L8ZrONbv7_0(.dout(w_dff_A_cBCe8gcX8_0),.din(w_dff_A_L8ZrONbv7_0),.clk(gclk));
	jdff dff_A_cBCe8gcX8_0(.dout(w_dff_A_dH9tmkyX1_0),.din(w_dff_A_cBCe8gcX8_0),.clk(gclk));
	jdff dff_A_dH9tmkyX1_0(.dout(w_dff_A_imBoMl9G9_0),.din(w_dff_A_dH9tmkyX1_0),.clk(gclk));
	jdff dff_A_imBoMl9G9_0(.dout(w_dff_A_W1mS41bH9_0),.din(w_dff_A_imBoMl9G9_0),.clk(gclk));
	jdff dff_A_W1mS41bH9_0(.dout(w_dff_A_ACIeM6bW5_0),.din(w_dff_A_W1mS41bH9_0),.clk(gclk));
	jdff dff_A_ACIeM6bW5_0(.dout(w_dff_A_644sRsx45_0),.din(w_dff_A_ACIeM6bW5_0),.clk(gclk));
	jdff dff_A_644sRsx45_0(.dout(w_dff_A_LJUwWryI9_0),.din(w_dff_A_644sRsx45_0),.clk(gclk));
	jdff dff_A_LJUwWryI9_0(.dout(w_dff_A_bX0adZO72_0),.din(w_dff_A_LJUwWryI9_0),.clk(gclk));
	jdff dff_A_bX0adZO72_0(.dout(w_dff_A_TtQPRtxi8_0),.din(w_dff_A_bX0adZO72_0),.clk(gclk));
	jdff dff_A_TtQPRtxi8_0(.dout(w_dff_A_ZvkeB0Gf4_0),.din(w_dff_A_TtQPRtxi8_0),.clk(gclk));
	jdff dff_A_ZvkeB0Gf4_0(.dout(w_dff_A_ZYE6agFO2_0),.din(w_dff_A_ZvkeB0Gf4_0),.clk(gclk));
	jdff dff_A_ZYE6agFO2_0(.dout(w_dff_A_JTmjFYKV3_0),.din(w_dff_A_ZYE6agFO2_0),.clk(gclk));
	jdff dff_A_JTmjFYKV3_0(.dout(w_dff_A_HzLv7mXe8_0),.din(w_dff_A_JTmjFYKV3_0),.clk(gclk));
	jdff dff_A_HzLv7mXe8_0(.dout(w_dff_A_4jUeqfUz6_0),.din(w_dff_A_HzLv7mXe8_0),.clk(gclk));
	jdff dff_A_4jUeqfUz6_0(.dout(w_dff_A_YM0Fr3Pz8_0),.din(w_dff_A_4jUeqfUz6_0),.clk(gclk));
	jdff dff_A_YM0Fr3Pz8_0(.dout(w_dff_A_IRmNQcGl4_0),.din(w_dff_A_YM0Fr3Pz8_0),.clk(gclk));
	jdff dff_A_IRmNQcGl4_0(.dout(w_dff_A_hpYCYBbp1_0),.din(w_dff_A_IRmNQcGl4_0),.clk(gclk));
	jdff dff_A_hpYCYBbp1_0(.dout(w_dff_A_xdIs2me35_0),.din(w_dff_A_hpYCYBbp1_0),.clk(gclk));
	jdff dff_A_xdIs2me35_0(.dout(G4946gat),.din(w_dff_A_xdIs2me35_0),.clk(gclk));
	jdff dff_A_8ScMJPuv8_2(.dout(w_dff_A_1sXjWFsi8_0),.din(w_dff_A_8ScMJPuv8_2),.clk(gclk));
	jdff dff_A_1sXjWFsi8_0(.dout(w_dff_A_vTjFl9Rn3_0),.din(w_dff_A_1sXjWFsi8_0),.clk(gclk));
	jdff dff_A_vTjFl9Rn3_0(.dout(w_dff_A_NMYpmCh04_0),.din(w_dff_A_vTjFl9Rn3_0),.clk(gclk));
	jdff dff_A_NMYpmCh04_0(.dout(w_dff_A_XyPynqNI2_0),.din(w_dff_A_NMYpmCh04_0),.clk(gclk));
	jdff dff_A_XyPynqNI2_0(.dout(w_dff_A_CmQ5euX20_0),.din(w_dff_A_XyPynqNI2_0),.clk(gclk));
	jdff dff_A_CmQ5euX20_0(.dout(w_dff_A_kWoSzfOi0_0),.din(w_dff_A_CmQ5euX20_0),.clk(gclk));
	jdff dff_A_kWoSzfOi0_0(.dout(w_dff_A_7c1wBPh17_0),.din(w_dff_A_kWoSzfOi0_0),.clk(gclk));
	jdff dff_A_7c1wBPh17_0(.dout(w_dff_A_pbz9b6dE0_0),.din(w_dff_A_7c1wBPh17_0),.clk(gclk));
	jdff dff_A_pbz9b6dE0_0(.dout(w_dff_A_g1d3kRWY8_0),.din(w_dff_A_pbz9b6dE0_0),.clk(gclk));
	jdff dff_A_g1d3kRWY8_0(.dout(w_dff_A_cU7By3wf1_0),.din(w_dff_A_g1d3kRWY8_0),.clk(gclk));
	jdff dff_A_cU7By3wf1_0(.dout(w_dff_A_GsWeOOmM5_0),.din(w_dff_A_cU7By3wf1_0),.clk(gclk));
	jdff dff_A_GsWeOOmM5_0(.dout(w_dff_A_5ApPesxj5_0),.din(w_dff_A_GsWeOOmM5_0),.clk(gclk));
	jdff dff_A_5ApPesxj5_0(.dout(w_dff_A_kDEVRP9n3_0),.din(w_dff_A_5ApPesxj5_0),.clk(gclk));
	jdff dff_A_kDEVRP9n3_0(.dout(w_dff_A_g3OrA6nu4_0),.din(w_dff_A_kDEVRP9n3_0),.clk(gclk));
	jdff dff_A_g3OrA6nu4_0(.dout(w_dff_A_icC5L8Iv9_0),.din(w_dff_A_g3OrA6nu4_0),.clk(gclk));
	jdff dff_A_icC5L8Iv9_0(.dout(w_dff_A_w2HZqHfQ1_0),.din(w_dff_A_icC5L8Iv9_0),.clk(gclk));
	jdff dff_A_w2HZqHfQ1_0(.dout(w_dff_A_x3qiTCHS1_0),.din(w_dff_A_w2HZqHfQ1_0),.clk(gclk));
	jdff dff_A_x3qiTCHS1_0(.dout(w_dff_A_7ZqXSU3f2_0),.din(w_dff_A_x3qiTCHS1_0),.clk(gclk));
	jdff dff_A_7ZqXSU3f2_0(.dout(w_dff_A_lTpGPtBB9_0),.din(w_dff_A_7ZqXSU3f2_0),.clk(gclk));
	jdff dff_A_lTpGPtBB9_0(.dout(w_dff_A_eMUjKrFr8_0),.din(w_dff_A_lTpGPtBB9_0),.clk(gclk));
	jdff dff_A_eMUjKrFr8_0(.dout(w_dff_A_EEYxIu5s7_0),.din(w_dff_A_eMUjKrFr8_0),.clk(gclk));
	jdff dff_A_EEYxIu5s7_0(.dout(w_dff_A_4ZKLbhg75_0),.din(w_dff_A_EEYxIu5s7_0),.clk(gclk));
	jdff dff_A_4ZKLbhg75_0(.dout(w_dff_A_CZdMZ5Cv1_0),.din(w_dff_A_4ZKLbhg75_0),.clk(gclk));
	jdff dff_A_CZdMZ5Cv1_0(.dout(w_dff_A_UunUEequ1_0),.din(w_dff_A_CZdMZ5Cv1_0),.clk(gclk));
	jdff dff_A_UunUEequ1_0(.dout(w_dff_A_HyF0T5Xn1_0),.din(w_dff_A_UunUEequ1_0),.clk(gclk));
	jdff dff_A_HyF0T5Xn1_0(.dout(w_dff_A_soyjrbM79_0),.din(w_dff_A_HyF0T5Xn1_0),.clk(gclk));
	jdff dff_A_soyjrbM79_0(.dout(w_dff_A_t6fhRwBl7_0),.din(w_dff_A_soyjrbM79_0),.clk(gclk));
	jdff dff_A_t6fhRwBl7_0(.dout(w_dff_A_ZCBCQ7Wy8_0),.din(w_dff_A_t6fhRwBl7_0),.clk(gclk));
	jdff dff_A_ZCBCQ7Wy8_0(.dout(w_dff_A_4bwfYfC41_0),.din(w_dff_A_ZCBCQ7Wy8_0),.clk(gclk));
	jdff dff_A_4bwfYfC41_0(.dout(w_dff_A_wPQlhMFN9_0),.din(w_dff_A_4bwfYfC41_0),.clk(gclk));
	jdff dff_A_wPQlhMFN9_0(.dout(w_dff_A_CvB16kXw1_0),.din(w_dff_A_wPQlhMFN9_0),.clk(gclk));
	jdff dff_A_CvB16kXw1_0(.dout(w_dff_A_EFMkvWW48_0),.din(w_dff_A_CvB16kXw1_0),.clk(gclk));
	jdff dff_A_EFMkvWW48_0(.dout(w_dff_A_B5lzMnH01_0),.din(w_dff_A_EFMkvWW48_0),.clk(gclk));
	jdff dff_A_B5lzMnH01_0(.dout(w_dff_A_foGIT7xW2_0),.din(w_dff_A_B5lzMnH01_0),.clk(gclk));
	jdff dff_A_foGIT7xW2_0(.dout(w_dff_A_7aqBwVGZ2_0),.din(w_dff_A_foGIT7xW2_0),.clk(gclk));
	jdff dff_A_7aqBwVGZ2_0(.dout(w_dff_A_vP8nQb8o3_0),.din(w_dff_A_7aqBwVGZ2_0),.clk(gclk));
	jdff dff_A_vP8nQb8o3_0(.dout(w_dff_A_ogiUPDms9_0),.din(w_dff_A_vP8nQb8o3_0),.clk(gclk));
	jdff dff_A_ogiUPDms9_0(.dout(w_dff_A_mVvJiUQc0_0),.din(w_dff_A_ogiUPDms9_0),.clk(gclk));
	jdff dff_A_mVvJiUQc0_0(.dout(G5308gat),.din(w_dff_A_mVvJiUQc0_0),.clk(gclk));
	jdff dff_A_rUJAEsv64_2(.dout(w_dff_A_JYqPvBDT0_0),.din(w_dff_A_rUJAEsv64_2),.clk(gclk));
	jdff dff_A_JYqPvBDT0_0(.dout(w_dff_A_VYAN729f8_0),.din(w_dff_A_JYqPvBDT0_0),.clk(gclk));
	jdff dff_A_VYAN729f8_0(.dout(w_dff_A_qtCHvmpF5_0),.din(w_dff_A_VYAN729f8_0),.clk(gclk));
	jdff dff_A_qtCHvmpF5_0(.dout(w_dff_A_SrxwfNOz6_0),.din(w_dff_A_qtCHvmpF5_0),.clk(gclk));
	jdff dff_A_SrxwfNOz6_0(.dout(w_dff_A_BXNLoJpd5_0),.din(w_dff_A_SrxwfNOz6_0),.clk(gclk));
	jdff dff_A_BXNLoJpd5_0(.dout(w_dff_A_QhYkGcty4_0),.din(w_dff_A_BXNLoJpd5_0),.clk(gclk));
	jdff dff_A_QhYkGcty4_0(.dout(w_dff_A_t12lW47r2_0),.din(w_dff_A_QhYkGcty4_0),.clk(gclk));
	jdff dff_A_t12lW47r2_0(.dout(w_dff_A_hSiAqwwP3_0),.din(w_dff_A_t12lW47r2_0),.clk(gclk));
	jdff dff_A_hSiAqwwP3_0(.dout(w_dff_A_GwI3OZQm6_0),.din(w_dff_A_hSiAqwwP3_0),.clk(gclk));
	jdff dff_A_GwI3OZQm6_0(.dout(w_dff_A_r2Trua028_0),.din(w_dff_A_GwI3OZQm6_0),.clk(gclk));
	jdff dff_A_r2Trua028_0(.dout(w_dff_A_Fi9ds2FE8_0),.din(w_dff_A_r2Trua028_0),.clk(gclk));
	jdff dff_A_Fi9ds2FE8_0(.dout(w_dff_A_clqbhO766_0),.din(w_dff_A_Fi9ds2FE8_0),.clk(gclk));
	jdff dff_A_clqbhO766_0(.dout(w_dff_A_eCqlIYJn5_0),.din(w_dff_A_clqbhO766_0),.clk(gclk));
	jdff dff_A_eCqlIYJn5_0(.dout(w_dff_A_WJqIf4YB2_0),.din(w_dff_A_eCqlIYJn5_0),.clk(gclk));
	jdff dff_A_WJqIf4YB2_0(.dout(w_dff_A_fPTxrkDm3_0),.din(w_dff_A_WJqIf4YB2_0),.clk(gclk));
	jdff dff_A_fPTxrkDm3_0(.dout(w_dff_A_a2vJftVL1_0),.din(w_dff_A_fPTxrkDm3_0),.clk(gclk));
	jdff dff_A_a2vJftVL1_0(.dout(w_dff_A_x2fm1VxS0_0),.din(w_dff_A_a2vJftVL1_0),.clk(gclk));
	jdff dff_A_x2fm1VxS0_0(.dout(w_dff_A_OEf8OgmG6_0),.din(w_dff_A_x2fm1VxS0_0),.clk(gclk));
	jdff dff_A_OEf8OgmG6_0(.dout(w_dff_A_QCqVLBS73_0),.din(w_dff_A_OEf8OgmG6_0),.clk(gclk));
	jdff dff_A_QCqVLBS73_0(.dout(w_dff_A_nZiHrkMA3_0),.din(w_dff_A_QCqVLBS73_0),.clk(gclk));
	jdff dff_A_nZiHrkMA3_0(.dout(w_dff_A_vE1RCgDa7_0),.din(w_dff_A_nZiHrkMA3_0),.clk(gclk));
	jdff dff_A_vE1RCgDa7_0(.dout(w_dff_A_G56Oklg13_0),.din(w_dff_A_vE1RCgDa7_0),.clk(gclk));
	jdff dff_A_G56Oklg13_0(.dout(w_dff_A_CSodMM0w7_0),.din(w_dff_A_G56Oklg13_0),.clk(gclk));
	jdff dff_A_CSodMM0w7_0(.dout(w_dff_A_zcaXJL5A1_0),.din(w_dff_A_CSodMM0w7_0),.clk(gclk));
	jdff dff_A_zcaXJL5A1_0(.dout(w_dff_A_YWyc4epU3_0),.din(w_dff_A_zcaXJL5A1_0),.clk(gclk));
	jdff dff_A_YWyc4epU3_0(.dout(w_dff_A_Pjvj8V4g0_0),.din(w_dff_A_YWyc4epU3_0),.clk(gclk));
	jdff dff_A_Pjvj8V4g0_0(.dout(w_dff_A_Z0MHmglx6_0),.din(w_dff_A_Pjvj8V4g0_0),.clk(gclk));
	jdff dff_A_Z0MHmglx6_0(.dout(w_dff_A_ECyjikka2_0),.din(w_dff_A_Z0MHmglx6_0),.clk(gclk));
	jdff dff_A_ECyjikka2_0(.dout(w_dff_A_yYyqOtGw9_0),.din(w_dff_A_ECyjikka2_0),.clk(gclk));
	jdff dff_A_yYyqOtGw9_0(.dout(w_dff_A_tH8tLAvU3_0),.din(w_dff_A_yYyqOtGw9_0),.clk(gclk));
	jdff dff_A_tH8tLAvU3_0(.dout(w_dff_A_SSE78vj12_0),.din(w_dff_A_tH8tLAvU3_0),.clk(gclk));
	jdff dff_A_SSE78vj12_0(.dout(w_dff_A_TorGxQLr8_0),.din(w_dff_A_SSE78vj12_0),.clk(gclk));
	jdff dff_A_TorGxQLr8_0(.dout(w_dff_A_uww9Xvi05_0),.din(w_dff_A_TorGxQLr8_0),.clk(gclk));
	jdff dff_A_uww9Xvi05_0(.dout(w_dff_A_RyQFf0FN1_0),.din(w_dff_A_uww9Xvi05_0),.clk(gclk));
	jdff dff_A_RyQFf0FN1_0(.dout(w_dff_A_YBcaU1TX9_0),.din(w_dff_A_RyQFf0FN1_0),.clk(gclk));
	jdff dff_A_YBcaU1TX9_0(.dout(G5672gat),.din(w_dff_A_YBcaU1TX9_0),.clk(gclk));
	jdff dff_A_84xyMY4Y3_2(.dout(w_dff_A_XTJhTSGg9_0),.din(w_dff_A_84xyMY4Y3_2),.clk(gclk));
	jdff dff_A_XTJhTSGg9_0(.dout(w_dff_A_sXhMawUE8_0),.din(w_dff_A_XTJhTSGg9_0),.clk(gclk));
	jdff dff_A_sXhMawUE8_0(.dout(w_dff_A_sN2E6JPZ3_0),.din(w_dff_A_sXhMawUE8_0),.clk(gclk));
	jdff dff_A_sN2E6JPZ3_0(.dout(w_dff_A_b5ZxHcPc0_0),.din(w_dff_A_sN2E6JPZ3_0),.clk(gclk));
	jdff dff_A_b5ZxHcPc0_0(.dout(w_dff_A_FZyfrE312_0),.din(w_dff_A_b5ZxHcPc0_0),.clk(gclk));
	jdff dff_A_FZyfrE312_0(.dout(w_dff_A_QDPN4ozZ1_0),.din(w_dff_A_FZyfrE312_0),.clk(gclk));
	jdff dff_A_QDPN4ozZ1_0(.dout(w_dff_A_OY5geCES6_0),.din(w_dff_A_QDPN4ozZ1_0),.clk(gclk));
	jdff dff_A_OY5geCES6_0(.dout(w_dff_A_ZSWMtmIt5_0),.din(w_dff_A_OY5geCES6_0),.clk(gclk));
	jdff dff_A_ZSWMtmIt5_0(.dout(w_dff_A_MNDivmGy2_0),.din(w_dff_A_ZSWMtmIt5_0),.clk(gclk));
	jdff dff_A_MNDivmGy2_0(.dout(w_dff_A_lz1MYfga9_0),.din(w_dff_A_MNDivmGy2_0),.clk(gclk));
	jdff dff_A_lz1MYfga9_0(.dout(w_dff_A_s4EZuP6e6_0),.din(w_dff_A_lz1MYfga9_0),.clk(gclk));
	jdff dff_A_s4EZuP6e6_0(.dout(w_dff_A_afiW7GTk6_0),.din(w_dff_A_s4EZuP6e6_0),.clk(gclk));
	jdff dff_A_afiW7GTk6_0(.dout(w_dff_A_wQ7vsfjB9_0),.din(w_dff_A_afiW7GTk6_0),.clk(gclk));
	jdff dff_A_wQ7vsfjB9_0(.dout(w_dff_A_K8JOOwg21_0),.din(w_dff_A_wQ7vsfjB9_0),.clk(gclk));
	jdff dff_A_K8JOOwg21_0(.dout(w_dff_A_kr6VHYWe5_0),.din(w_dff_A_K8JOOwg21_0),.clk(gclk));
	jdff dff_A_kr6VHYWe5_0(.dout(w_dff_A_dEIxKwy43_0),.din(w_dff_A_kr6VHYWe5_0),.clk(gclk));
	jdff dff_A_dEIxKwy43_0(.dout(w_dff_A_nerKESo28_0),.din(w_dff_A_dEIxKwy43_0),.clk(gclk));
	jdff dff_A_nerKESo28_0(.dout(w_dff_A_wPxiTZLp4_0),.din(w_dff_A_nerKESo28_0),.clk(gclk));
	jdff dff_A_wPxiTZLp4_0(.dout(w_dff_A_YLDbwvF19_0),.din(w_dff_A_wPxiTZLp4_0),.clk(gclk));
	jdff dff_A_YLDbwvF19_0(.dout(w_dff_A_OdnUEPO55_0),.din(w_dff_A_YLDbwvF19_0),.clk(gclk));
	jdff dff_A_OdnUEPO55_0(.dout(w_dff_A_P9sAmqPJ3_0),.din(w_dff_A_OdnUEPO55_0),.clk(gclk));
	jdff dff_A_P9sAmqPJ3_0(.dout(w_dff_A_dFpb3NUm9_0),.din(w_dff_A_P9sAmqPJ3_0),.clk(gclk));
	jdff dff_A_dFpb3NUm9_0(.dout(w_dff_A_JLc2T2nW7_0),.din(w_dff_A_dFpb3NUm9_0),.clk(gclk));
	jdff dff_A_JLc2T2nW7_0(.dout(w_dff_A_fsLSZjJc9_0),.din(w_dff_A_JLc2T2nW7_0),.clk(gclk));
	jdff dff_A_fsLSZjJc9_0(.dout(w_dff_A_PO2quGnb2_0),.din(w_dff_A_fsLSZjJc9_0),.clk(gclk));
	jdff dff_A_PO2quGnb2_0(.dout(w_dff_A_d323YXze7_0),.din(w_dff_A_PO2quGnb2_0),.clk(gclk));
	jdff dff_A_d323YXze7_0(.dout(w_dff_A_gbjPXZff0_0),.din(w_dff_A_d323YXze7_0),.clk(gclk));
	jdff dff_A_gbjPXZff0_0(.dout(w_dff_A_gVATgN0m7_0),.din(w_dff_A_gbjPXZff0_0),.clk(gclk));
	jdff dff_A_gVATgN0m7_0(.dout(w_dff_A_L4cqZF7I6_0),.din(w_dff_A_gVATgN0m7_0),.clk(gclk));
	jdff dff_A_L4cqZF7I6_0(.dout(w_dff_A_bpGAAgeE1_0),.din(w_dff_A_L4cqZF7I6_0),.clk(gclk));
	jdff dff_A_bpGAAgeE1_0(.dout(w_dff_A_xB0BdyQL4_0),.din(w_dff_A_bpGAAgeE1_0),.clk(gclk));
	jdff dff_A_xB0BdyQL4_0(.dout(w_dff_A_hRShA0ed5_0),.din(w_dff_A_xB0BdyQL4_0),.clk(gclk));
	jdff dff_A_hRShA0ed5_0(.dout(G5971gat),.din(w_dff_A_hRShA0ed5_0),.clk(gclk));
	jdff dff_A_1raJBPiI7_2(.dout(w_dff_A_b0A700nA8_0),.din(w_dff_A_1raJBPiI7_2),.clk(gclk));
	jdff dff_A_b0A700nA8_0(.dout(w_dff_A_EtbUJt987_0),.din(w_dff_A_b0A700nA8_0),.clk(gclk));
	jdff dff_A_EtbUJt987_0(.dout(w_dff_A_0swVoc0V3_0),.din(w_dff_A_EtbUJt987_0),.clk(gclk));
	jdff dff_A_0swVoc0V3_0(.dout(w_dff_A_CHqs3Bxe6_0),.din(w_dff_A_0swVoc0V3_0),.clk(gclk));
	jdff dff_A_CHqs3Bxe6_0(.dout(w_dff_A_FyJscuXk5_0),.din(w_dff_A_CHqs3Bxe6_0),.clk(gclk));
	jdff dff_A_FyJscuXk5_0(.dout(w_dff_A_DgTOnl1P9_0),.din(w_dff_A_FyJscuXk5_0),.clk(gclk));
	jdff dff_A_DgTOnl1P9_0(.dout(w_dff_A_Ax5KdSXQ6_0),.din(w_dff_A_DgTOnl1P9_0),.clk(gclk));
	jdff dff_A_Ax5KdSXQ6_0(.dout(w_dff_A_mQf30PIE5_0),.din(w_dff_A_Ax5KdSXQ6_0),.clk(gclk));
	jdff dff_A_mQf30PIE5_0(.dout(w_dff_A_tbPuAVsh2_0),.din(w_dff_A_mQf30PIE5_0),.clk(gclk));
	jdff dff_A_tbPuAVsh2_0(.dout(w_dff_A_LP01NtDK9_0),.din(w_dff_A_tbPuAVsh2_0),.clk(gclk));
	jdff dff_A_LP01NtDK9_0(.dout(w_dff_A_21FkTXyp3_0),.din(w_dff_A_LP01NtDK9_0),.clk(gclk));
	jdff dff_A_21FkTXyp3_0(.dout(w_dff_A_qIWPi15m5_0),.din(w_dff_A_21FkTXyp3_0),.clk(gclk));
	jdff dff_A_qIWPi15m5_0(.dout(w_dff_A_lQbnPwvX5_0),.din(w_dff_A_qIWPi15m5_0),.clk(gclk));
	jdff dff_A_lQbnPwvX5_0(.dout(w_dff_A_NtDgGHN10_0),.din(w_dff_A_lQbnPwvX5_0),.clk(gclk));
	jdff dff_A_NtDgGHN10_0(.dout(w_dff_A_uYrhRVcn8_0),.din(w_dff_A_NtDgGHN10_0),.clk(gclk));
	jdff dff_A_uYrhRVcn8_0(.dout(w_dff_A_iF8emuVV5_0),.din(w_dff_A_uYrhRVcn8_0),.clk(gclk));
	jdff dff_A_iF8emuVV5_0(.dout(w_dff_A_S7Rt2u0W1_0),.din(w_dff_A_iF8emuVV5_0),.clk(gclk));
	jdff dff_A_S7Rt2u0W1_0(.dout(w_dff_A_T447om4z0_0),.din(w_dff_A_S7Rt2u0W1_0),.clk(gclk));
	jdff dff_A_T447om4z0_0(.dout(w_dff_A_VVqMdkWK7_0),.din(w_dff_A_T447om4z0_0),.clk(gclk));
	jdff dff_A_VVqMdkWK7_0(.dout(w_dff_A_AhsZsNcg0_0),.din(w_dff_A_VVqMdkWK7_0),.clk(gclk));
	jdff dff_A_AhsZsNcg0_0(.dout(w_dff_A_1B0OHMJC9_0),.din(w_dff_A_AhsZsNcg0_0),.clk(gclk));
	jdff dff_A_1B0OHMJC9_0(.dout(w_dff_A_XWSbTKbY2_0),.din(w_dff_A_1B0OHMJC9_0),.clk(gclk));
	jdff dff_A_XWSbTKbY2_0(.dout(w_dff_A_1lvipsKF1_0),.din(w_dff_A_XWSbTKbY2_0),.clk(gclk));
	jdff dff_A_1lvipsKF1_0(.dout(w_dff_A_2lzSU0s65_0),.din(w_dff_A_1lvipsKF1_0),.clk(gclk));
	jdff dff_A_2lzSU0s65_0(.dout(w_dff_A_KPlMCcWP0_0),.din(w_dff_A_2lzSU0s65_0),.clk(gclk));
	jdff dff_A_KPlMCcWP0_0(.dout(w_dff_A_YKhpwTBF5_0),.din(w_dff_A_KPlMCcWP0_0),.clk(gclk));
	jdff dff_A_YKhpwTBF5_0(.dout(w_dff_A_1lOkirMM1_0),.din(w_dff_A_YKhpwTBF5_0),.clk(gclk));
	jdff dff_A_1lOkirMM1_0(.dout(w_dff_A_NgKhnMyS0_0),.din(w_dff_A_1lOkirMM1_0),.clk(gclk));
	jdff dff_A_NgKhnMyS0_0(.dout(w_dff_A_4ZOHlOK03_0),.din(w_dff_A_NgKhnMyS0_0),.clk(gclk));
	jdff dff_A_4ZOHlOK03_0(.dout(G6123gat),.din(w_dff_A_4ZOHlOK03_0),.clk(gclk));
	jdff dff_A_y2Cx0Ugv4_2(.dout(w_dff_A_IM9zw3ip2_0),.din(w_dff_A_y2Cx0Ugv4_2),.clk(gclk));
	jdff dff_A_IM9zw3ip2_0(.dout(w_dff_A_GuG5kwK45_0),.din(w_dff_A_IM9zw3ip2_0),.clk(gclk));
	jdff dff_A_GuG5kwK45_0(.dout(w_dff_A_HQDaexNy9_0),.din(w_dff_A_GuG5kwK45_0),.clk(gclk));
	jdff dff_A_HQDaexNy9_0(.dout(w_dff_A_XFlsTBiF8_0),.din(w_dff_A_HQDaexNy9_0),.clk(gclk));
	jdff dff_A_XFlsTBiF8_0(.dout(w_dff_A_tLsJc26L9_0),.din(w_dff_A_XFlsTBiF8_0),.clk(gclk));
	jdff dff_A_tLsJc26L9_0(.dout(w_dff_A_YPpQaonI8_0),.din(w_dff_A_tLsJc26L9_0),.clk(gclk));
	jdff dff_A_YPpQaonI8_0(.dout(w_dff_A_JD7hAYLi4_0),.din(w_dff_A_YPpQaonI8_0),.clk(gclk));
	jdff dff_A_JD7hAYLi4_0(.dout(w_dff_A_iyCJsjJN7_0),.din(w_dff_A_JD7hAYLi4_0),.clk(gclk));
	jdff dff_A_iyCJsjJN7_0(.dout(w_dff_A_rR3kr6zM4_0),.din(w_dff_A_iyCJsjJN7_0),.clk(gclk));
	jdff dff_A_rR3kr6zM4_0(.dout(w_dff_A_sG66h2zR4_0),.din(w_dff_A_rR3kr6zM4_0),.clk(gclk));
	jdff dff_A_sG66h2zR4_0(.dout(w_dff_A_7VOJ2J6Z1_0),.din(w_dff_A_sG66h2zR4_0),.clk(gclk));
	jdff dff_A_7VOJ2J6Z1_0(.dout(w_dff_A_W3vTYauk0_0),.din(w_dff_A_7VOJ2J6Z1_0),.clk(gclk));
	jdff dff_A_W3vTYauk0_0(.dout(w_dff_A_NM2eYEB24_0),.din(w_dff_A_W3vTYauk0_0),.clk(gclk));
	jdff dff_A_NM2eYEB24_0(.dout(w_dff_A_8YuQDSsh2_0),.din(w_dff_A_NM2eYEB24_0),.clk(gclk));
	jdff dff_A_8YuQDSsh2_0(.dout(w_dff_A_T6skV5jX5_0),.din(w_dff_A_8YuQDSsh2_0),.clk(gclk));
	jdff dff_A_T6skV5jX5_0(.dout(w_dff_A_Vt2bouFW6_0),.din(w_dff_A_T6skV5jX5_0),.clk(gclk));
	jdff dff_A_Vt2bouFW6_0(.dout(w_dff_A_H0Wn6B0I3_0),.din(w_dff_A_Vt2bouFW6_0),.clk(gclk));
	jdff dff_A_H0Wn6B0I3_0(.dout(w_dff_A_1PG892WP2_0),.din(w_dff_A_H0Wn6B0I3_0),.clk(gclk));
	jdff dff_A_1PG892WP2_0(.dout(w_dff_A_agF66L0e9_0),.din(w_dff_A_1PG892WP2_0),.clk(gclk));
	jdff dff_A_agF66L0e9_0(.dout(w_dff_A_JACyKZqv6_0),.din(w_dff_A_agF66L0e9_0),.clk(gclk));
	jdff dff_A_JACyKZqv6_0(.dout(w_dff_A_YgNyNfM41_0),.din(w_dff_A_JACyKZqv6_0),.clk(gclk));
	jdff dff_A_YgNyNfM41_0(.dout(w_dff_A_hrW6acbg0_0),.din(w_dff_A_YgNyNfM41_0),.clk(gclk));
	jdff dff_A_hrW6acbg0_0(.dout(w_dff_A_WcMAmwaU7_0),.din(w_dff_A_hrW6acbg0_0),.clk(gclk));
	jdff dff_A_WcMAmwaU7_0(.dout(w_dff_A_6SV7dqQK4_0),.din(w_dff_A_WcMAmwaU7_0),.clk(gclk));
	jdff dff_A_6SV7dqQK4_0(.dout(w_dff_A_8apvyxvv6_0),.din(w_dff_A_6SV7dqQK4_0),.clk(gclk));
	jdff dff_A_8apvyxvv6_0(.dout(w_dff_A_gd8vqqrV6_0),.din(w_dff_A_8apvyxvv6_0),.clk(gclk));
	jdff dff_A_gd8vqqrV6_0(.dout(w_dff_A_SUNrvR1n8_0),.din(w_dff_A_gd8vqqrV6_0),.clk(gclk));
	jdff dff_A_SUNrvR1n8_0(.dout(G6150gat),.din(w_dff_A_SUNrvR1n8_0),.clk(gclk));
	jdff dff_A_SvwK5EUw5_2(.dout(w_dff_A_bjd83Vxj5_0),.din(w_dff_A_SvwK5EUw5_2),.clk(gclk));
	jdff dff_A_bjd83Vxj5_0(.dout(w_dff_A_x9BftWh56_0),.din(w_dff_A_bjd83Vxj5_0),.clk(gclk));
	jdff dff_A_x9BftWh56_0(.dout(w_dff_A_bwo486E10_0),.din(w_dff_A_x9BftWh56_0),.clk(gclk));
	jdff dff_A_bwo486E10_0(.dout(w_dff_A_xkMMLt5c7_0),.din(w_dff_A_bwo486E10_0),.clk(gclk));
	jdff dff_A_xkMMLt5c7_0(.dout(w_dff_A_ruSffF2E4_0),.din(w_dff_A_xkMMLt5c7_0),.clk(gclk));
	jdff dff_A_ruSffF2E4_0(.dout(w_dff_A_u83didJi9_0),.din(w_dff_A_ruSffF2E4_0),.clk(gclk));
	jdff dff_A_u83didJi9_0(.dout(w_dff_A_SX9Eezw61_0),.din(w_dff_A_u83didJi9_0),.clk(gclk));
	jdff dff_A_SX9Eezw61_0(.dout(w_dff_A_VywakCAI0_0),.din(w_dff_A_SX9Eezw61_0),.clk(gclk));
	jdff dff_A_VywakCAI0_0(.dout(w_dff_A_HHhOAcAy8_0),.din(w_dff_A_VywakCAI0_0),.clk(gclk));
	jdff dff_A_HHhOAcAy8_0(.dout(w_dff_A_RGovoSLq4_0),.din(w_dff_A_HHhOAcAy8_0),.clk(gclk));
	jdff dff_A_RGovoSLq4_0(.dout(w_dff_A_c6mK9v437_0),.din(w_dff_A_RGovoSLq4_0),.clk(gclk));
	jdff dff_A_c6mK9v437_0(.dout(w_dff_A_Mdxt7XPY9_0),.din(w_dff_A_c6mK9v437_0),.clk(gclk));
	jdff dff_A_Mdxt7XPY9_0(.dout(w_dff_A_5Jr7QOea1_0),.din(w_dff_A_Mdxt7XPY9_0),.clk(gclk));
	jdff dff_A_5Jr7QOea1_0(.dout(w_dff_A_hoZveZIZ4_0),.din(w_dff_A_5Jr7QOea1_0),.clk(gclk));
	jdff dff_A_hoZveZIZ4_0(.dout(w_dff_A_HVlW4p3D1_0),.din(w_dff_A_hoZveZIZ4_0),.clk(gclk));
	jdff dff_A_HVlW4p3D1_0(.dout(w_dff_A_nKuLprAn3_0),.din(w_dff_A_HVlW4p3D1_0),.clk(gclk));
	jdff dff_A_nKuLprAn3_0(.dout(w_dff_A_ofZYTtmx6_0),.din(w_dff_A_nKuLprAn3_0),.clk(gclk));
	jdff dff_A_ofZYTtmx6_0(.dout(w_dff_A_DiCHfkEQ6_0),.din(w_dff_A_ofZYTtmx6_0),.clk(gclk));
	jdff dff_A_DiCHfkEQ6_0(.dout(w_dff_A_x0CBrwWu5_0),.din(w_dff_A_DiCHfkEQ6_0),.clk(gclk));
	jdff dff_A_x0CBrwWu5_0(.dout(w_dff_A_u5hkAvVI5_0),.din(w_dff_A_x0CBrwWu5_0),.clk(gclk));
	jdff dff_A_u5hkAvVI5_0(.dout(w_dff_A_CiM46Hfy3_0),.din(w_dff_A_u5hkAvVI5_0),.clk(gclk));
	jdff dff_A_CiM46Hfy3_0(.dout(w_dff_A_H4TnNXJI2_0),.din(w_dff_A_CiM46Hfy3_0),.clk(gclk));
	jdff dff_A_H4TnNXJI2_0(.dout(w_dff_A_KLkNfKOu4_0),.din(w_dff_A_H4TnNXJI2_0),.clk(gclk));
	jdff dff_A_KLkNfKOu4_0(.dout(w_dff_A_4oFE5pXi0_0),.din(w_dff_A_KLkNfKOu4_0),.clk(gclk));
	jdff dff_A_4oFE5pXi0_0(.dout(w_dff_A_s39hK2rb3_0),.din(w_dff_A_4oFE5pXi0_0),.clk(gclk));
	jdff dff_A_s39hK2rb3_0(.dout(G6160gat),.din(w_dff_A_s39hK2rb3_0),.clk(gclk));
	jdff dff_A_EELcdX9T0_2(.dout(w_dff_A_gufvd4Sv1_0),.din(w_dff_A_EELcdX9T0_2),.clk(gclk));
	jdff dff_A_gufvd4Sv1_0(.dout(w_dff_A_EHNCK4Ft7_0),.din(w_dff_A_gufvd4Sv1_0),.clk(gclk));
	jdff dff_A_EHNCK4Ft7_0(.dout(w_dff_A_SZNA8S4J5_0),.din(w_dff_A_EHNCK4Ft7_0),.clk(gclk));
	jdff dff_A_SZNA8S4J5_0(.dout(w_dff_A_UP180uH48_0),.din(w_dff_A_SZNA8S4J5_0),.clk(gclk));
	jdff dff_A_UP180uH48_0(.dout(w_dff_A_7tOsaqMl7_0),.din(w_dff_A_UP180uH48_0),.clk(gclk));
	jdff dff_A_7tOsaqMl7_0(.dout(w_dff_A_EqdzPePq4_0),.din(w_dff_A_7tOsaqMl7_0),.clk(gclk));
	jdff dff_A_EqdzPePq4_0(.dout(w_dff_A_BFf5iGPR9_0),.din(w_dff_A_EqdzPePq4_0),.clk(gclk));
	jdff dff_A_BFf5iGPR9_0(.dout(w_dff_A_hSUBVtHL8_0),.din(w_dff_A_BFf5iGPR9_0),.clk(gclk));
	jdff dff_A_hSUBVtHL8_0(.dout(w_dff_A_gfs4PPv88_0),.din(w_dff_A_hSUBVtHL8_0),.clk(gclk));
	jdff dff_A_gfs4PPv88_0(.dout(w_dff_A_lEIKIGiG4_0),.din(w_dff_A_gfs4PPv88_0),.clk(gclk));
	jdff dff_A_lEIKIGiG4_0(.dout(w_dff_A_NJddlC4g2_0),.din(w_dff_A_lEIKIGiG4_0),.clk(gclk));
	jdff dff_A_NJddlC4g2_0(.dout(w_dff_A_omlpZSum4_0),.din(w_dff_A_NJddlC4g2_0),.clk(gclk));
	jdff dff_A_omlpZSum4_0(.dout(w_dff_A_qHPpO4G22_0),.din(w_dff_A_omlpZSum4_0),.clk(gclk));
	jdff dff_A_qHPpO4G22_0(.dout(w_dff_A_fYwezJSA2_0),.din(w_dff_A_qHPpO4G22_0),.clk(gclk));
	jdff dff_A_fYwezJSA2_0(.dout(w_dff_A_Xq5Ii9hC4_0),.din(w_dff_A_fYwezJSA2_0),.clk(gclk));
	jdff dff_A_Xq5Ii9hC4_0(.dout(w_dff_A_RkjQx0pg0_0),.din(w_dff_A_Xq5Ii9hC4_0),.clk(gclk));
	jdff dff_A_RkjQx0pg0_0(.dout(w_dff_A_posI18bm7_0),.din(w_dff_A_RkjQx0pg0_0),.clk(gclk));
	jdff dff_A_posI18bm7_0(.dout(w_dff_A_TsSkDL2w4_0),.din(w_dff_A_posI18bm7_0),.clk(gclk));
	jdff dff_A_TsSkDL2w4_0(.dout(w_dff_A_5DnQ9DTu6_0),.din(w_dff_A_TsSkDL2w4_0),.clk(gclk));
	jdff dff_A_5DnQ9DTu6_0(.dout(w_dff_A_jF8lu5fj3_0),.din(w_dff_A_5DnQ9DTu6_0),.clk(gclk));
	jdff dff_A_jF8lu5fj3_0(.dout(w_dff_A_Eb4STl0r7_0),.din(w_dff_A_jF8lu5fj3_0),.clk(gclk));
	jdff dff_A_Eb4STl0r7_0(.dout(w_dff_A_hW0BFO5Z8_0),.din(w_dff_A_Eb4STl0r7_0),.clk(gclk));
	jdff dff_A_hW0BFO5Z8_0(.dout(w_dff_A_L1grFQ8m3_0),.din(w_dff_A_hW0BFO5Z8_0),.clk(gclk));
	jdff dff_A_L1grFQ8m3_0(.dout(w_dff_A_nA71Rspl2_0),.din(w_dff_A_L1grFQ8m3_0),.clk(gclk));
	jdff dff_A_nA71Rspl2_0(.dout(G6170gat),.din(w_dff_A_nA71Rspl2_0),.clk(gclk));
	jdff dff_A_RRpqyqj39_2(.dout(w_dff_A_W05T6Vtq2_0),.din(w_dff_A_RRpqyqj39_2),.clk(gclk));
	jdff dff_A_W05T6Vtq2_0(.dout(w_dff_A_iB45JsjX3_0),.din(w_dff_A_W05T6Vtq2_0),.clk(gclk));
	jdff dff_A_iB45JsjX3_0(.dout(w_dff_A_WJcSqkwi3_0),.din(w_dff_A_iB45JsjX3_0),.clk(gclk));
	jdff dff_A_WJcSqkwi3_0(.dout(w_dff_A_23r1uK1y2_0),.din(w_dff_A_WJcSqkwi3_0),.clk(gclk));
	jdff dff_A_23r1uK1y2_0(.dout(w_dff_A_r2igO0z46_0),.din(w_dff_A_23r1uK1y2_0),.clk(gclk));
	jdff dff_A_r2igO0z46_0(.dout(w_dff_A_aJnIeCz43_0),.din(w_dff_A_r2igO0z46_0),.clk(gclk));
	jdff dff_A_aJnIeCz43_0(.dout(w_dff_A_oK8tOAyr2_0),.din(w_dff_A_aJnIeCz43_0),.clk(gclk));
	jdff dff_A_oK8tOAyr2_0(.dout(w_dff_A_OeqywrbW2_0),.din(w_dff_A_oK8tOAyr2_0),.clk(gclk));
	jdff dff_A_OeqywrbW2_0(.dout(w_dff_A_EROGwThe8_0),.din(w_dff_A_OeqywrbW2_0),.clk(gclk));
	jdff dff_A_EROGwThe8_0(.dout(w_dff_A_YvPWHAVr6_0),.din(w_dff_A_EROGwThe8_0),.clk(gclk));
	jdff dff_A_YvPWHAVr6_0(.dout(w_dff_A_AQ2TWwBn4_0),.din(w_dff_A_YvPWHAVr6_0),.clk(gclk));
	jdff dff_A_AQ2TWwBn4_0(.dout(w_dff_A_SjyFdkBI1_0),.din(w_dff_A_AQ2TWwBn4_0),.clk(gclk));
	jdff dff_A_SjyFdkBI1_0(.dout(w_dff_A_fYnjaFlm9_0),.din(w_dff_A_SjyFdkBI1_0),.clk(gclk));
	jdff dff_A_fYnjaFlm9_0(.dout(w_dff_A_R8zPP88j0_0),.din(w_dff_A_fYnjaFlm9_0),.clk(gclk));
	jdff dff_A_R8zPP88j0_0(.dout(w_dff_A_ZQQzkbON9_0),.din(w_dff_A_R8zPP88j0_0),.clk(gclk));
	jdff dff_A_ZQQzkbON9_0(.dout(w_dff_A_R9C4OhDh2_0),.din(w_dff_A_ZQQzkbON9_0),.clk(gclk));
	jdff dff_A_R9C4OhDh2_0(.dout(w_dff_A_ZruFFfjo8_0),.din(w_dff_A_R9C4OhDh2_0),.clk(gclk));
	jdff dff_A_ZruFFfjo8_0(.dout(w_dff_A_34NIgfUP0_0),.din(w_dff_A_ZruFFfjo8_0),.clk(gclk));
	jdff dff_A_34NIgfUP0_0(.dout(w_dff_A_hEit6H518_0),.din(w_dff_A_34NIgfUP0_0),.clk(gclk));
	jdff dff_A_hEit6H518_0(.dout(w_dff_A_iNBAwf6Y9_0),.din(w_dff_A_hEit6H518_0),.clk(gclk));
	jdff dff_A_iNBAwf6Y9_0(.dout(w_dff_A_eS1NZCvx0_0),.din(w_dff_A_iNBAwf6Y9_0),.clk(gclk));
	jdff dff_A_eS1NZCvx0_0(.dout(w_dff_A_D9cfx2J05_0),.din(w_dff_A_eS1NZCvx0_0),.clk(gclk));
	jdff dff_A_D9cfx2J05_0(.dout(G6180gat),.din(w_dff_A_D9cfx2J05_0),.clk(gclk));
	jdff dff_A_qnZGkGXX4_2(.dout(w_dff_A_MrUqgbmz4_0),.din(w_dff_A_qnZGkGXX4_2),.clk(gclk));
	jdff dff_A_MrUqgbmz4_0(.dout(w_dff_A_YzHzUYsy2_0),.din(w_dff_A_MrUqgbmz4_0),.clk(gclk));
	jdff dff_A_YzHzUYsy2_0(.dout(w_dff_A_BQpyPue48_0),.din(w_dff_A_YzHzUYsy2_0),.clk(gclk));
	jdff dff_A_BQpyPue48_0(.dout(w_dff_A_ToE0Uzaa1_0),.din(w_dff_A_BQpyPue48_0),.clk(gclk));
	jdff dff_A_ToE0Uzaa1_0(.dout(w_dff_A_GTcSazS79_0),.din(w_dff_A_ToE0Uzaa1_0),.clk(gclk));
	jdff dff_A_GTcSazS79_0(.dout(w_dff_A_e1O9BePz0_0),.din(w_dff_A_GTcSazS79_0),.clk(gclk));
	jdff dff_A_e1O9BePz0_0(.dout(w_dff_A_L34fsglg0_0),.din(w_dff_A_e1O9BePz0_0),.clk(gclk));
	jdff dff_A_L34fsglg0_0(.dout(w_dff_A_5SBShVGD5_0),.din(w_dff_A_L34fsglg0_0),.clk(gclk));
	jdff dff_A_5SBShVGD5_0(.dout(w_dff_A_Cac4DcrY6_0),.din(w_dff_A_5SBShVGD5_0),.clk(gclk));
	jdff dff_A_Cac4DcrY6_0(.dout(w_dff_A_dbFnQviG9_0),.din(w_dff_A_Cac4DcrY6_0),.clk(gclk));
	jdff dff_A_dbFnQviG9_0(.dout(w_dff_A_dxRFwI2D7_0),.din(w_dff_A_dbFnQviG9_0),.clk(gclk));
	jdff dff_A_dxRFwI2D7_0(.dout(w_dff_A_IKDAjMqW5_0),.din(w_dff_A_dxRFwI2D7_0),.clk(gclk));
	jdff dff_A_IKDAjMqW5_0(.dout(w_dff_A_3b0H7rvu6_0),.din(w_dff_A_IKDAjMqW5_0),.clk(gclk));
	jdff dff_A_3b0H7rvu6_0(.dout(w_dff_A_SdRXAC8i4_0),.din(w_dff_A_3b0H7rvu6_0),.clk(gclk));
	jdff dff_A_SdRXAC8i4_0(.dout(w_dff_A_CmQM7OPJ6_0),.din(w_dff_A_SdRXAC8i4_0),.clk(gclk));
	jdff dff_A_CmQM7OPJ6_0(.dout(w_dff_A_Xl1H6DCG8_0),.din(w_dff_A_CmQM7OPJ6_0),.clk(gclk));
	jdff dff_A_Xl1H6DCG8_0(.dout(w_dff_A_pXI6Kagq6_0),.din(w_dff_A_Xl1H6DCG8_0),.clk(gclk));
	jdff dff_A_pXI6Kagq6_0(.dout(w_dff_A_ijoNJwum0_0),.din(w_dff_A_pXI6Kagq6_0),.clk(gclk));
	jdff dff_A_ijoNJwum0_0(.dout(w_dff_A_WVQpKK2N9_0),.din(w_dff_A_ijoNJwum0_0),.clk(gclk));
	jdff dff_A_WVQpKK2N9_0(.dout(w_dff_A_Xo1pRnTM3_0),.din(w_dff_A_WVQpKK2N9_0),.clk(gclk));
	jdff dff_A_Xo1pRnTM3_0(.dout(G6190gat),.din(w_dff_A_Xo1pRnTM3_0),.clk(gclk));
	jdff dff_A_WXOrmoWW8_2(.dout(w_dff_A_YD9nUo5Y2_0),.din(w_dff_A_WXOrmoWW8_2),.clk(gclk));
	jdff dff_A_YD9nUo5Y2_0(.dout(w_dff_A_6222Yix48_0),.din(w_dff_A_YD9nUo5Y2_0),.clk(gclk));
	jdff dff_A_6222Yix48_0(.dout(w_dff_A_VLK1D3XO4_0),.din(w_dff_A_6222Yix48_0),.clk(gclk));
	jdff dff_A_VLK1D3XO4_0(.dout(w_dff_A_qqwnvcOY4_0),.din(w_dff_A_VLK1D3XO4_0),.clk(gclk));
	jdff dff_A_qqwnvcOY4_0(.dout(w_dff_A_HhTak8JX4_0),.din(w_dff_A_qqwnvcOY4_0),.clk(gclk));
	jdff dff_A_HhTak8JX4_0(.dout(w_dff_A_XeoNVGQX0_0),.din(w_dff_A_HhTak8JX4_0),.clk(gclk));
	jdff dff_A_XeoNVGQX0_0(.dout(w_dff_A_L9N8ivgX5_0),.din(w_dff_A_XeoNVGQX0_0),.clk(gclk));
	jdff dff_A_L9N8ivgX5_0(.dout(w_dff_A_UwsvkvX28_0),.din(w_dff_A_L9N8ivgX5_0),.clk(gclk));
	jdff dff_A_UwsvkvX28_0(.dout(w_dff_A_f94bDBZ40_0),.din(w_dff_A_UwsvkvX28_0),.clk(gclk));
	jdff dff_A_f94bDBZ40_0(.dout(w_dff_A_ugLDeNNj6_0),.din(w_dff_A_f94bDBZ40_0),.clk(gclk));
	jdff dff_A_ugLDeNNj6_0(.dout(w_dff_A_9EmocGAs7_0),.din(w_dff_A_ugLDeNNj6_0),.clk(gclk));
	jdff dff_A_9EmocGAs7_0(.dout(w_dff_A_XOfhhKrZ3_0),.din(w_dff_A_9EmocGAs7_0),.clk(gclk));
	jdff dff_A_XOfhhKrZ3_0(.dout(w_dff_A_EA5B83wV8_0),.din(w_dff_A_XOfhhKrZ3_0),.clk(gclk));
	jdff dff_A_EA5B83wV8_0(.dout(w_dff_A_292ORCPw0_0),.din(w_dff_A_EA5B83wV8_0),.clk(gclk));
	jdff dff_A_292ORCPw0_0(.dout(w_dff_A_scfpyQbO1_0),.din(w_dff_A_292ORCPw0_0),.clk(gclk));
	jdff dff_A_scfpyQbO1_0(.dout(w_dff_A_7aiN5HCM8_0),.din(w_dff_A_scfpyQbO1_0),.clk(gclk));
	jdff dff_A_7aiN5HCM8_0(.dout(w_dff_A_eLb1kdS36_0),.din(w_dff_A_7aiN5HCM8_0),.clk(gclk));
	jdff dff_A_eLb1kdS36_0(.dout(w_dff_A_0C9Oi0wz7_0),.din(w_dff_A_eLb1kdS36_0),.clk(gclk));
	jdff dff_A_0C9Oi0wz7_0(.dout(G6200gat),.din(w_dff_A_0C9Oi0wz7_0),.clk(gclk));
	jdff dff_A_zBf6HHia3_2(.dout(w_dff_A_Cu2Gj7gW1_0),.din(w_dff_A_zBf6HHia3_2),.clk(gclk));
	jdff dff_A_Cu2Gj7gW1_0(.dout(w_dff_A_mbzG29En6_0),.din(w_dff_A_Cu2Gj7gW1_0),.clk(gclk));
	jdff dff_A_mbzG29En6_0(.dout(w_dff_A_1lPBvm1B0_0),.din(w_dff_A_mbzG29En6_0),.clk(gclk));
	jdff dff_A_1lPBvm1B0_0(.dout(w_dff_A_0oyWFeur6_0),.din(w_dff_A_1lPBvm1B0_0),.clk(gclk));
	jdff dff_A_0oyWFeur6_0(.dout(w_dff_A_QbFecoML7_0),.din(w_dff_A_0oyWFeur6_0),.clk(gclk));
	jdff dff_A_QbFecoML7_0(.dout(w_dff_A_YuUqoDk83_0),.din(w_dff_A_QbFecoML7_0),.clk(gclk));
	jdff dff_A_YuUqoDk83_0(.dout(w_dff_A_6B1ZG7hd4_0),.din(w_dff_A_YuUqoDk83_0),.clk(gclk));
	jdff dff_A_6B1ZG7hd4_0(.dout(w_dff_A_RGKk3GKA7_0),.din(w_dff_A_6B1ZG7hd4_0),.clk(gclk));
	jdff dff_A_RGKk3GKA7_0(.dout(w_dff_A_Y2WspOBJ8_0),.din(w_dff_A_RGKk3GKA7_0),.clk(gclk));
	jdff dff_A_Y2WspOBJ8_0(.dout(w_dff_A_2FOAFc9a3_0),.din(w_dff_A_Y2WspOBJ8_0),.clk(gclk));
	jdff dff_A_2FOAFc9a3_0(.dout(w_dff_A_gbxlx1kB9_0),.din(w_dff_A_2FOAFc9a3_0),.clk(gclk));
	jdff dff_A_gbxlx1kB9_0(.dout(w_dff_A_ygU1NomP4_0),.din(w_dff_A_gbxlx1kB9_0),.clk(gclk));
	jdff dff_A_ygU1NomP4_0(.dout(w_dff_A_D51HS72s5_0),.din(w_dff_A_ygU1NomP4_0),.clk(gclk));
	jdff dff_A_D51HS72s5_0(.dout(w_dff_A_3SlxXx1b3_0),.din(w_dff_A_D51HS72s5_0),.clk(gclk));
	jdff dff_A_3SlxXx1b3_0(.dout(w_dff_A_PNUJ3g586_0),.din(w_dff_A_3SlxXx1b3_0),.clk(gclk));
	jdff dff_A_PNUJ3g586_0(.dout(w_dff_A_vkEGzOEX2_0),.din(w_dff_A_PNUJ3g586_0),.clk(gclk));
	jdff dff_A_vkEGzOEX2_0(.dout(G6210gat),.din(w_dff_A_vkEGzOEX2_0),.clk(gclk));
	jdff dff_A_VdYZ4TDy2_2(.dout(w_dff_A_QqM89tHL5_0),.din(w_dff_A_VdYZ4TDy2_2),.clk(gclk));
	jdff dff_A_QqM89tHL5_0(.dout(w_dff_A_bQEtXRSJ5_0),.din(w_dff_A_QqM89tHL5_0),.clk(gclk));
	jdff dff_A_bQEtXRSJ5_0(.dout(w_dff_A_Xqh191pB3_0),.din(w_dff_A_bQEtXRSJ5_0),.clk(gclk));
	jdff dff_A_Xqh191pB3_0(.dout(w_dff_A_MNYBlyGd7_0),.din(w_dff_A_Xqh191pB3_0),.clk(gclk));
	jdff dff_A_MNYBlyGd7_0(.dout(w_dff_A_QEuc27FI9_0),.din(w_dff_A_MNYBlyGd7_0),.clk(gclk));
	jdff dff_A_QEuc27FI9_0(.dout(w_dff_A_3Q6eYBmT0_0),.din(w_dff_A_QEuc27FI9_0),.clk(gclk));
	jdff dff_A_3Q6eYBmT0_0(.dout(w_dff_A_HwoLkaH27_0),.din(w_dff_A_3Q6eYBmT0_0),.clk(gclk));
	jdff dff_A_HwoLkaH27_0(.dout(w_dff_A_JWFBjUrt6_0),.din(w_dff_A_HwoLkaH27_0),.clk(gclk));
	jdff dff_A_JWFBjUrt6_0(.dout(w_dff_A_TnUyeyoj9_0),.din(w_dff_A_JWFBjUrt6_0),.clk(gclk));
	jdff dff_A_TnUyeyoj9_0(.dout(w_dff_A_mBhYgjfA1_0),.din(w_dff_A_TnUyeyoj9_0),.clk(gclk));
	jdff dff_A_mBhYgjfA1_0(.dout(w_dff_A_26BAZ0Yn0_0),.din(w_dff_A_mBhYgjfA1_0),.clk(gclk));
	jdff dff_A_26BAZ0Yn0_0(.dout(w_dff_A_jbabzuMu4_0),.din(w_dff_A_26BAZ0Yn0_0),.clk(gclk));
	jdff dff_A_jbabzuMu4_0(.dout(w_dff_A_vc4KjUy91_0),.din(w_dff_A_jbabzuMu4_0),.clk(gclk));
	jdff dff_A_vc4KjUy91_0(.dout(w_dff_A_rdeBYawA9_0),.din(w_dff_A_vc4KjUy91_0),.clk(gclk));
	jdff dff_A_rdeBYawA9_0(.dout(G6220gat),.din(w_dff_A_rdeBYawA9_0),.clk(gclk));
	jdff dff_A_AlZA3pCn3_2(.dout(w_dff_A_IjYaULZR8_0),.din(w_dff_A_AlZA3pCn3_2),.clk(gclk));
	jdff dff_A_IjYaULZR8_0(.dout(w_dff_A_TbbjLwsR9_0),.din(w_dff_A_IjYaULZR8_0),.clk(gclk));
	jdff dff_A_TbbjLwsR9_0(.dout(w_dff_A_CC1v8XDI2_0),.din(w_dff_A_TbbjLwsR9_0),.clk(gclk));
	jdff dff_A_CC1v8XDI2_0(.dout(w_dff_A_WuSmD3gK6_0),.din(w_dff_A_CC1v8XDI2_0),.clk(gclk));
	jdff dff_A_WuSmD3gK6_0(.dout(w_dff_A_HXNWaxWZ9_0),.din(w_dff_A_WuSmD3gK6_0),.clk(gclk));
	jdff dff_A_HXNWaxWZ9_0(.dout(w_dff_A_f5cnWkfv1_0),.din(w_dff_A_HXNWaxWZ9_0),.clk(gclk));
	jdff dff_A_f5cnWkfv1_0(.dout(w_dff_A_kuvEhMcr4_0),.din(w_dff_A_f5cnWkfv1_0),.clk(gclk));
	jdff dff_A_kuvEhMcr4_0(.dout(w_dff_A_hnGk9Q8V0_0),.din(w_dff_A_kuvEhMcr4_0),.clk(gclk));
	jdff dff_A_hnGk9Q8V0_0(.dout(w_dff_A_UeqvxuhD3_0),.din(w_dff_A_hnGk9Q8V0_0),.clk(gclk));
	jdff dff_A_UeqvxuhD3_0(.dout(w_dff_A_h6LR23uM8_0),.din(w_dff_A_UeqvxuhD3_0),.clk(gclk));
	jdff dff_A_h6LR23uM8_0(.dout(w_dff_A_4yqZ4Pre6_0),.din(w_dff_A_h6LR23uM8_0),.clk(gclk));
	jdff dff_A_4yqZ4Pre6_0(.dout(w_dff_A_VzHzPI6Y7_0),.din(w_dff_A_4yqZ4Pre6_0),.clk(gclk));
	jdff dff_A_VzHzPI6Y7_0(.dout(G6230gat),.din(w_dff_A_VzHzPI6Y7_0),.clk(gclk));
	jdff dff_A_x9YO84OD2_2(.dout(w_dff_A_q9IerLkm3_0),.din(w_dff_A_x9YO84OD2_2),.clk(gclk));
	jdff dff_A_q9IerLkm3_0(.dout(w_dff_A_EVgzEf1Q6_0),.din(w_dff_A_q9IerLkm3_0),.clk(gclk));
	jdff dff_A_EVgzEf1Q6_0(.dout(w_dff_A_sl9KLPig2_0),.din(w_dff_A_EVgzEf1Q6_0),.clk(gclk));
	jdff dff_A_sl9KLPig2_0(.dout(w_dff_A_yxgyofFe1_0),.din(w_dff_A_sl9KLPig2_0),.clk(gclk));
	jdff dff_A_yxgyofFe1_0(.dout(w_dff_A_5rflpenG1_0),.din(w_dff_A_yxgyofFe1_0),.clk(gclk));
	jdff dff_A_5rflpenG1_0(.dout(w_dff_A_WzzfEBtd4_0),.din(w_dff_A_5rflpenG1_0),.clk(gclk));
	jdff dff_A_WzzfEBtd4_0(.dout(w_dff_A_iKVcCPPa2_0),.din(w_dff_A_WzzfEBtd4_0),.clk(gclk));
	jdff dff_A_iKVcCPPa2_0(.dout(w_dff_A_MREacc6p1_0),.din(w_dff_A_iKVcCPPa2_0),.clk(gclk));
	jdff dff_A_MREacc6p1_0(.dout(w_dff_A_AcLskXXc1_0),.din(w_dff_A_MREacc6p1_0),.clk(gclk));
	jdff dff_A_AcLskXXc1_0(.dout(w_dff_A_1g6mJbci7_0),.din(w_dff_A_AcLskXXc1_0),.clk(gclk));
	jdff dff_A_1g6mJbci7_0(.dout(G6240gat),.din(w_dff_A_1g6mJbci7_0),.clk(gclk));
	jdff dff_A_YgTyAIea9_2(.dout(w_dff_A_FdapSK7r3_0),.din(w_dff_A_YgTyAIea9_2),.clk(gclk));
	jdff dff_A_FdapSK7r3_0(.dout(w_dff_A_OQPZteuG2_0),.din(w_dff_A_FdapSK7r3_0),.clk(gclk));
	jdff dff_A_OQPZteuG2_0(.dout(w_dff_A_iKWHgDRZ0_0),.din(w_dff_A_OQPZteuG2_0),.clk(gclk));
	jdff dff_A_iKWHgDRZ0_0(.dout(w_dff_A_TtcaAFp44_0),.din(w_dff_A_iKWHgDRZ0_0),.clk(gclk));
	jdff dff_A_TtcaAFp44_0(.dout(w_dff_A_pWpLbvuA9_0),.din(w_dff_A_TtcaAFp44_0),.clk(gclk));
	jdff dff_A_pWpLbvuA9_0(.dout(w_dff_A_N5GSayY97_0),.din(w_dff_A_pWpLbvuA9_0),.clk(gclk));
	jdff dff_A_N5GSayY97_0(.dout(w_dff_A_LIox8mrh5_0),.din(w_dff_A_N5GSayY97_0),.clk(gclk));
	jdff dff_A_LIox8mrh5_0(.dout(w_dff_A_CjxTm4vc0_0),.din(w_dff_A_LIox8mrh5_0),.clk(gclk));
	jdff dff_A_CjxTm4vc0_0(.dout(G6250gat),.din(w_dff_A_CjxTm4vc0_0),.clk(gclk));
	jdff dff_A_1aNiPV9I1_2(.dout(w_dff_A_yw6ZvmmJ6_0),.din(w_dff_A_1aNiPV9I1_2),.clk(gclk));
	jdff dff_A_yw6ZvmmJ6_0(.dout(w_dff_A_RUHFp4pu4_0),.din(w_dff_A_yw6ZvmmJ6_0),.clk(gclk));
	jdff dff_A_RUHFp4pu4_0(.dout(w_dff_A_QqBqEDwE9_0),.din(w_dff_A_RUHFp4pu4_0),.clk(gclk));
	jdff dff_A_QqBqEDwE9_0(.dout(w_dff_A_V0roDClD2_0),.din(w_dff_A_QqBqEDwE9_0),.clk(gclk));
	jdff dff_A_V0roDClD2_0(.dout(w_dff_A_4dMcpDyQ8_0),.din(w_dff_A_V0roDClD2_0),.clk(gclk));
	jdff dff_A_4dMcpDyQ8_0(.dout(w_dff_A_FBcr8KZO8_0),.din(w_dff_A_4dMcpDyQ8_0),.clk(gclk));
	jdff dff_A_FBcr8KZO8_0(.dout(G6260gat),.din(w_dff_A_FBcr8KZO8_0),.clk(gclk));
	jdff dff_A_xYpvdcGX7_2(.dout(w_dff_A_boGHSrLK5_0),.din(w_dff_A_xYpvdcGX7_2),.clk(gclk));
	jdff dff_A_boGHSrLK5_0(.dout(w_dff_A_setKgQZu2_0),.din(w_dff_A_boGHSrLK5_0),.clk(gclk));
	jdff dff_A_setKgQZu2_0(.dout(w_dff_A_pB90dIRx5_0),.din(w_dff_A_setKgQZu2_0),.clk(gclk));
	jdff dff_A_pB90dIRx5_0(.dout(w_dff_A_7SeyXxwC1_0),.din(w_dff_A_pB90dIRx5_0),.clk(gclk));
	jdff dff_A_7SeyXxwC1_0(.dout(G6270gat),.din(w_dff_A_7SeyXxwC1_0),.clk(gclk));
	jdff dff_A_oBPVQzMN0_2(.dout(w_dff_A_XdEtSXX40_0),.din(w_dff_A_oBPVQzMN0_2),.clk(gclk));
	jdff dff_A_XdEtSXX40_0(.dout(w_dff_A_JZUSrm1M4_0),.din(w_dff_A_XdEtSXX40_0),.clk(gclk));
	jdff dff_A_JZUSrm1M4_0(.dout(G6280gat),.din(w_dff_A_JZUSrm1M4_0),.clk(gclk));
	jdff dff_A_i6yb8BNW4_2(.dout(G6288gat),.din(w_dff_A_i6yb8BNW4_2),.clk(gclk));
endmodule

