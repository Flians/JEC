// Benchmark "top" written by ABC on Thu May 28 22:01:50 2020

module rf_log2 ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] ;
  wire n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
    n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
    n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
    n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
    n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
    n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
    n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
    n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
    n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
    n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
    n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
    n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
    n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
    n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
    n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
    n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
    n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
    n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
    n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
    n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
    n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
    n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
    n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
    n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
    n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
    n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
    n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
    n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
    n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
    n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
    n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
    n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
    n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
    n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
    n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
    n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
    n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
    n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
    n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
    n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
    n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
    n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
    n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
    n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
    n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
    n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
    n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
    n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
    n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
    n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
    n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
    n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
    n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
    n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
    n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
    n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
    n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
    n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
    n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
    n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
    n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
    n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
    n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
    n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
    n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
    n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
    n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
    n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
    n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
    n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
    n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
    n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
    n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
    n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
    n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
    n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
    n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
    n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
    n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
    n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
    n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
    n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
    n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
    n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
    n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
    n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
    n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
    n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
    n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
    n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
    n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
    n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
    n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
    n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
    n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
    n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
    n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
    n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
    n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
    n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
    n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
    n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
    n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
    n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
    n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
    n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
    n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
    n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
    n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
    n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
    n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
    n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
    n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
    n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
    n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
    n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
    n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
    n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
    n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
    n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
    n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
    n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
    n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
    n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
    n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
    n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
    n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
    n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
    n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
    n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
    n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
    n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
    n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
    n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
    n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
    n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
    n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
    n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
    n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
    n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
    n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
    n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
    n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
    n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
    n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
    n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
    n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
    n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
    n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
    n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
    n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
    n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
    n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
    n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
    n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
    n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
    n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
    n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
    n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
    n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
    n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
    n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
    n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
    n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
    n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
    n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
    n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
    n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
    n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
    n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
    n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
    n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
    n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
    n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
    n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
    n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
    n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
    n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
    n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
    n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
    n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
    n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
    n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
    n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
    n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
    n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
    n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
    n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
    n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
    n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
    n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
    n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
    n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
    n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
    n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
    n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
    n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
    n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
    n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
    n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
    n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
    n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
    n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
    n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
    n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
    n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
    n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
    n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
    n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
    n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
    n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
    n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
    n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
    n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
    n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
    n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
    n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
    n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
    n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
    n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
    n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
    n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
    n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
    n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
    n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
    n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
    n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
    n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
    n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
    n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
    n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
    n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
    n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
    n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
    n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
    n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
    n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
    n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
    n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
    n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
    n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
    n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
    n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
    n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
    n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
    n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
    n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
    n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
    n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
    n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
    n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
    n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
    n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
    n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
    n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
    n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
    n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
    n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
    n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
    n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
    n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
    n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
    n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
    n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
    n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
    n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
    n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
    n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
    n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
    n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
    n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
    n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
    n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
    n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
    n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
    n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
    n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
    n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
    n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
    n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
    n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
    n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
    n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
    n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
    n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
    n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
    n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
    n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
    n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
    n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
    n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
    n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
    n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
    n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
    n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
    n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
    n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
    n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
    n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
    n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
    n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
    n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
    n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
    n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
    n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
    n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
    n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
    n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
    n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
    n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
    n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
    n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
    n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
    n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
    n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
    n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
    n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
    n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
    n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
    n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
    n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
    n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
    n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
    n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
    n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
    n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
    n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
    n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
    n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
    n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
    n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
    n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
    n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
    n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
    n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
    n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
    n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
    n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
    n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
    n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
    n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
    n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
    n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
    n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
    n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
    n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
    n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
    n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
    n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
    n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
    n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
    n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
    n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
    n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
    n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
    n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
    n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
    n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
    n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
    n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
    n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
    n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
    n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
    n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
    n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
    n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
    n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
    n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
    n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
    n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
    n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
    n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
    n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
    n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
    n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
    n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
    n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
    n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
    n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
    n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
    n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
    n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
    n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
    n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
    n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
    n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
    n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
    n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
    n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
    n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
    n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
    n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
    n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
    n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
    n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
    n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
    n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
    n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
    n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
    n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
    n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
    n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
    n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
    n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
    n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
    n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
    n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
    n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
    n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
    n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
    n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
    n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
    n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
    n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
    n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
    n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
    n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
    n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
    n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
    n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
    n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
    n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
    n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
    n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
    n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
    n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
    n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
    n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
    n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
    n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
    n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
    n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
    n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
    n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
    n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
    n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
    n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
    n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
    n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
    n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
    n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
    n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
    n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
    n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
    n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
    n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
    n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
    n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
    n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
    n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
    n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
    n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
    n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
    n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
    n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
    n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
    n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
    n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
    n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
    n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
    n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
    n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
    n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
    n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
    n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
    n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
    n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
    n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
    n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
    n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
    n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
    n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
    n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
    n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
    n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
    n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
    n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
    n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
    n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
    n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
    n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
    n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
    n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
    n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
    n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
    n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
    n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
    n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
    n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
    n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
    n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
    n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
    n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
    n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
    n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
    n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
    n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
    n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
    n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
    n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
    n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
    n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
    n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
    n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
    n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
    n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
    n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
    n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
    n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
    n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
    n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
    n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
    n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
    n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
    n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
    n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
    n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
    n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
    n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
    n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
    n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
    n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
    n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
    n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
    n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
    n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
    n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
    n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
    n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
    n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
    n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
    n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
    n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
    n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
    n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
    n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
    n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
    n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
    n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
    n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
    n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
    n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
    n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
    n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
    n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
    n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
    n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
    n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
    n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
    n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
    n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
    n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
    n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
    n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
    n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
    n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
    n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
    n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
    n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
    n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
    n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
    n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
    n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
    n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
    n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
    n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
    n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
    n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
    n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
    n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
    n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
    n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
    n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
    n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
    n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
    n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
    n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
    n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
    n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
    n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
    n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
    n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
    n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
    n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
    n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
    n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
    n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
    n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
    n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
    n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
    n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
    n11479, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
    n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
    n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
    n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
    n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
    n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
    n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
    n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
    n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
    n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
    n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
    n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
    n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
    n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
    n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
    n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
    n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
    n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
    n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
    n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
    n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
    n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
    n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
    n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
    n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
    n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
    n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
    n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
    n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
    n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
    n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
    n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
    n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
    n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
    n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
    n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
    n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
    n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
    n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
    n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
    n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
    n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
    n12323, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
    n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
    n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
    n12352, n12353, n12354, n12355, n12357, n12359, n12360, n12361, n12362,
    n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
    n12372, n12373, n12374, n12375, n12378, n12379, n12380, n12381, n12382,
    n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
    n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
    n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
    n12437, n12438, n12439, n12455, n12456, n12457, n12458, n12459, n12460,
    n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
    n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
    n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
    n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
    n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
    n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
    n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
    n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
    n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
    n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
    n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
    n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
    n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
    n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
    n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
    n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
    n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
    n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
    n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
    n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
    n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
    n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
    n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
    n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
    n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
    n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
    n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
    n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
    n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
    n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
    n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
    n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
    n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
    n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
    n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
    n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
    n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
    n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
    n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
    n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
    n12822, n12823, n12824, n12825, n12829, n12834, n12835, n12836, n12837,
    n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
    n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
    n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
    n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
    n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
    n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
    n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
    n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
    n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
    n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
    n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
    n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
    n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
    n12955, n12956, n12957, n12958, n12959, n12961, n12962, n12963, n12964,
    n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
    n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
    n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
    n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
    n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
    n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
    n13021, n13022, n13023, n13025, n13026, n13027, n13028, n13029, n13030,
    n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
    n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
    n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
    n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
    n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
    n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
    n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
    n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
    n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
    n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
    n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
    n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
    n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
    n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
    n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
    n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
    n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
    n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
    n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
    n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
    n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
    n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
    n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
    n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
    n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
    n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
    n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
    n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
    n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
    n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
    n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
    n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
    n13346, n13347, n13348, n13349, n13350, n13352, n13353, n13354, n13356,
    n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
    n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
    n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
    n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
    n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
    n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
    n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
    n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
    n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
    n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
    n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
    n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
    n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
    n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
    n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
    n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
    n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
    n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
    n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
    n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
    n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
    n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13559,
    n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
    n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
    n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
    n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
    n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
    n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
    n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
    n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
    n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
    n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
    n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
    n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
    n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
    n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
    n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
    n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
    n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
    n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
    n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
    n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
    n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
    n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
    n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
    n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
    n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
    n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
    n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
    n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
    n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
    n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
    n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
    n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
    n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
    n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
    n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
    n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
    n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
    n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
    n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
    n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
    n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
    n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
    n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
    n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
    n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
    n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
    n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
    n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
    n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
    n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
    n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
    n14023, n14024, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
    n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
    n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
    n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
    n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
    n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
    n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
    n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
    n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
    n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
    n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
    n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
    n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
    n14141, n14142, n14143, n14144, n14147, n14152, n14153, n14154, n14155,
    n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
    n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
    n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
    n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
    n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
    n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
    n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
    n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
    n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
    n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
    n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
    n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
    n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
    n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
    n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
    n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
    n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
    n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
    n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
    n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
    n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
    n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
    n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
    n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
    n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
    n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
    n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
    n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
    n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
    n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
    n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
    n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
    n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
    n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
    n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
    n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
    n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
    n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
    n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
    n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
    n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
    n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
    n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
    n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
    n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
    n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14705,
    n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
    n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
    n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
    n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
    n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
    n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
    n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
    n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
    n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
    n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
    n14835, n14836, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
    n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
    n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
    n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
    n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
    n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
    n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
    n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
    n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
    n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
    n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
    n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
    n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
    n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
    n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
    n14971, n14972, n14975, n14980, n14981, n14982, n14983, n14984, n14985,
    n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
    n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
    n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
    n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
    n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
    n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
    n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
    n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
    n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
    n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
    n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
    n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
    n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
    n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
    n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
    n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
    n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
    n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
    n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
    n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
    n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
    n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
    n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
    n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
    n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
    n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
    n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
    n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
    n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
    n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
    n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
    n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
    n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15283,
    n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
    n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
    n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
    n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
    n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
    n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
    n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
    n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
    n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
    n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
    n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
    n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
    n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
    n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
    n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
    n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
    n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
    n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
    n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
    n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
    n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
    n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
    n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
    n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
    n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
    n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
    n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
    n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
    n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
    n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
    n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
    n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
    n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
    n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
    n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
    n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
    n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
    n15620, n15621, n15622, n15623, n15624, n15625, n15627, n15628, n15629,
    n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
    n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
    n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
    n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
    n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
    n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
    n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
    n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
    n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
    n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
    n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
    n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
    n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
    n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
    n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
    n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
    n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
    n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
    n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
    n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
    n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
    n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
    n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
    n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
    n15981, n15982, n15985, n15990, n15991, n15992, n15993, n15994, n15995,
    n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
    n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
    n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
    n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
    n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
    n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
    n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
    n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
    n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
    n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
    n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
    n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
    n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
    n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
    n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
    n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
    n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
    n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
    n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
    n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
    n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
    n16392, n16393, n16395, n16399, n16400, n16401, n16402, n16403, n16404,
    n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
    n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
    n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
    n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
    n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
    n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
    n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
    n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
    n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
    n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
    n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
    n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
    n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
    n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
    n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
    n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
    n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
    n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
    n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
    n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
    n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
    n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
    n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
    n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
    n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
    n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
    n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
    n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
    n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
    n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
    n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
    n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
    n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
    n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
    n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
    n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
    n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
    n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
    n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
    n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
    n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
    n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
    n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
    n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
    n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16809, n16810,
    n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
    n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
    n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
    n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
    n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
    n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
    n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
    n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
    n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
    n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
    n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
    n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
    n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
    n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
    n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
    n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
    n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
    n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
    n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
    n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
    n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
    n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
    n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
    n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
    n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
    n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
    n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
    n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
    n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
    n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
    n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
    n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
    n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
    n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
    n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
    n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
    n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
    n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
    n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
    n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
    n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
    n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
    n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
    n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
    n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
    n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
    n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
    n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
    n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
    n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
    n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
    n17270, n17273, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
    n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
    n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
    n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
    n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
    n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
    n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
    n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
    n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
    n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
    n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
    n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
    n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
    n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
    n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
    n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
    n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
    n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
    n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
    n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
    n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
    n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
    n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
    n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
    n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
    n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
    n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
    n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
    n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
    n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
    n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
    n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
    n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
    n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
    n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
    n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
    n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
    n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
    n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
    n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
    n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
    n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
    n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
    n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
    n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
    n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
    n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
    n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
    n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
    n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
    n17744, n17745, n17746, n17747, n17748, n17749, n17751, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
    n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
    n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
    n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
    n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
    n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
    n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
    n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
    n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
    n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
    n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
    n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
    n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
    n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
    n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
    n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
    n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
    n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
    n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
    n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
    n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
    n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
    n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
    n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
    n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
    n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
    n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
    n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
    n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
    n18270, n18271, n18272, n18273, n18274, n18275, n18277, n18278, n18279,
    n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
    n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
    n18298, n18299, n18300, n18301, n18309, n18310, n18311, n18312, n18313,
    n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
    n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
    n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
    n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
    n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
    n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
    n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
    n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
    n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
    n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
    n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
    n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
    n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
    n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439,
    n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
    n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
    n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
    n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
    n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
    n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
    n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
    n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511,
    n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
    n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
    n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
    n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
    n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
    n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
    n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
    n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583,
    n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
    n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
    n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
    n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
    n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
    n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
    n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
    n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
    n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
    n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
    n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
    n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
    n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
    n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
    n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
    n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727,
    n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
    n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
    n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
    n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
    n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
    n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
    n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
    n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799,
    n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
    n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
    n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
    n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
    n18836, n18837, n18838, n18839, n18840, n18841, n18843, n18847, n18848,
    n18849, n18850, n18851, n18852, n18853, n18855, n18856, n18857, n18858,
    n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
    n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
    n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
    n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
    n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903,
    n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
    n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
    n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
    n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
    n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
    n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
    n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
    n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975,
    n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
    n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
    n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
    n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
    n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
    n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
    n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
    n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047,
    n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
    n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
    n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
    n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
    n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
    n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
    n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
    n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
    n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
    n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
    n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
    n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
    n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
    n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
    n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
    n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191,
    n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
    n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
    n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
    n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
    n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
    n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
    n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
    n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263,
    n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
    n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
    n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
    n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
    n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
    n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
    n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
    n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335,
    n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
    n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
    n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
    n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
    n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
    n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
    n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
    n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407,
    n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
    n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
    n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
    n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
    n19444, n19445, n19446, n19447, n19448, n19449, n19452, n19454, n19455,
    n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
    n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
    n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
    n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
    n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
    n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
    n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
    n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
    n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
    n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
    n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
    n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
    n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
    n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
    n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
    n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599,
    n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
    n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
    n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
    n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
    n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
    n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
    n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
    n19663, n19664, n19665, n19666, n19674, n19675, n19676, n19677, n19678,
    n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
    n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
    n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
    n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
    n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
    n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
    n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
    n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
    n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
    n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
    n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
    n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
    n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
    n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
    n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
    n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
    n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
    n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
    n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
    n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
    n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
    n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
    n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
    n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
    n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
    n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
    n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
    n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
    n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
    n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
    n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
    n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
    n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
    n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
    n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
    n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
    n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
    n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
    n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
    n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
    n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
    n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
    n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
    n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
    n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
    n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
    n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
    n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
    n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
    n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
    n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
    n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
    n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
    n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
    n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
    n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
    n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335,
    n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344,
    n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
    n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
    n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
    n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
    n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
    n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407,
    n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416,
    n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
    n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
    n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
    n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488,
    n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
    n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
    n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
    n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560,
    n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
    n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
    n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
    n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632,
    n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
    n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
    n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
    n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
    n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
    n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
    n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695,
    n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704,
    n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
    n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
    n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
    n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
    n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
    n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
    n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
    n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776,
    n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
    n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
    n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
    n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
    n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
    n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
    n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
    n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848,
    n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
    n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
    n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
    n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
    n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
    n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
    n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
    n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920,
    n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
    n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
    n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
    n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
    n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
    n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992,
    n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
    n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
    n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
    n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
    n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
    n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
    n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
    n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064,
    n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
    n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
    n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
    n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
    n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
    n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
    n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127,
    n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136,
    n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
    n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
    n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
    n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
    n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
    n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
    n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199,
    n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208,
    n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
    n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
    n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
    n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244,
    n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
    n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
    n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271,
    n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280,
    n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
    n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
    n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
    n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316,
    n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
    n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
    n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343,
    n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352,
    n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
    n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
    n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
    n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388,
    n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
    n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
    n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
    n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424,
    n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
    n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
    n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
    n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460,
    n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
    n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
    n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
    n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496,
    n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
    n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
    n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
    n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532,
    n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
    n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
    n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
    n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568,
    n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
    n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
    n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
    n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604,
    n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
    n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
    n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
    n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640,
    n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
    n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
    n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
    n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676,
    n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
    n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
    n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
    n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712,
    n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
    n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
    n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
    n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748,
    n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
    n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
    n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
    n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784,
    n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
    n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
    n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
    n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820,
    n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
    n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
    n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
    n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856,
    n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
    n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
    n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
    n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892,
    n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
    n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
    n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
    n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928,
    n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
    n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
    n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964,
    n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
    n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
    n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
    n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000,
    n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
    n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
    n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
    n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036,
    n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
    n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054,
    n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
    n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072,
    n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
    n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
    n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
    n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108,
    n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
    n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
    n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
    n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144,
    n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
    n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
    n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
    n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180,
    n22181, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
    n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
    n22200, n22201, n22202, n22204, n22205, n22206, n22207, n22208, n22209,
    n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
    n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
    n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
    n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245,
    n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
    n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
    n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
    n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
    n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
    n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
    n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
    n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317,
    n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326,
    n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
    n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
    n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
    n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
    n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
    n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
    n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389,
    n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
    n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
    n22408, n22409, n22410, n22411, n22412, n22413, n22416, n22418, n22419,
    n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428,
    n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437,
    n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446,
    n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
    n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464,
    n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
    n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
    n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
    n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500,
    n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509,
    n22510, n22511, n22512, n22513, n22521, n22522, n22523, n22524, n22525,
    n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534,
    n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
    n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552,
    n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22562,
    n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
    n22572, n22573, n22574, n22575, n22577, n22578, n22579, n22580, n22581,
    n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590,
    n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
    n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608,
    n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
    n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
    n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
    n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644,
    n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653,
    n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662,
    n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
    n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680,
    n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
    n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698,
    n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
    n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716,
    n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
    n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734,
    n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
    n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752,
    n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
    n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
    n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
    n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788,
    n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797,
    n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806,
    n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
    n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824,
    n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
    n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
    n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
    n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860,
    n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869,
    n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878,
    n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887,
    n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896,
    n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
    n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914,
    n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
    n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932,
    n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941,
    n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950,
    n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959,
    n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968,
    n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
    n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986,
    n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
    n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004,
    n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013,
    n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022,
    n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031,
    n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040,
    n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
    n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058,
    n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
    n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076,
    n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085,
    n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094,
    n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103,
    n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112,
    n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
    n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130,
    n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
    n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148,
    n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157,
    n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166,
    n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175,
    n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184,
    n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
    n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202,
    n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
    n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220,
    n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229,
    n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238,
    n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248,
    n23249, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
    n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23275,
    n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284,
    n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293,
    n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302,
    n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311,
    n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320,
    n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
    n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
    n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
    n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356,
    n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365,
    n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374,
    n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383,
    n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392,
    n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
    n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
    n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
    n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428,
    n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
    n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446,
    n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455,
    n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464,
    n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
    n23481, n23482, n23484, n23485, n23486, n23487, n23488, n23489, n23490,
    n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
    n23500, n23501, n23502, n23503, n23504, n23505, n23507, n23508, n23509,
    n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518,
    n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527,
    n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536,
    n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
    n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
    n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
    n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572,
    n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
    n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590,
    n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599,
    n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608,
    n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
    n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626,
    n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
    n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644,
    n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
    n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662,
    n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671,
    n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680,
    n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
    n23690, n23691, n23693, n23694, n23695, n23696, n23697, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711,
    n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23721,
    n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730,
    n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
    n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748,
    n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757,
    n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766,
    n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775,
    n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784,
    n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
    n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
    n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
    n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820,
    n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829,
    n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838,
    n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847,
    n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856,
    n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
    n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874,
    n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
    n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892,
    n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23902, n23903,
    n23904, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916,
    n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925,
    n23926, n23927, n23928, n23929, n23930, n23932, n23933, n23934, n23935,
    n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944,
    n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
    n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
    n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
    n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980,
    n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
    n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998,
    n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007,
    n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016,
    n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
    n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034,
    n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
    n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052,
    n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
    n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070,
    n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079,
    n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088,
    n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
    n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
    n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
    n24116, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
    n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142,
    n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151,
    n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
    n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170,
    n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
    n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188,
    n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197,
    n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206,
    n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215,
    n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224,
    n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
    n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242,
    n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
    n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260,
    n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269,
    n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278,
    n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287,
    n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296,
    n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
    n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314,
    n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
    n24324, n24325, n24326, n24328, n24329, n24330, n24331, n24332, n24333,
    n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342,
    n24343, n24344, n24345, n24346, n24347, n24349, n24350, n24351, n24352,
    n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
    n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370,
    n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
    n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388,
    n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397,
    n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406,
    n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
    n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
    n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
    n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
    n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
    n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460,
    n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469,
    n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478,
    n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
    n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,
    n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
    n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
    n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
    n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532,
    n24533, n24534, n24535, n24537, n24538, n24539, n24540, n24541, n24542,
    n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551,
    n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560,
    n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
    n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
    n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
    n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596,
    n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605,
    n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614,
    n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623,
    n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632,
    n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
    n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
    n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
    n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668,
    n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677,
    n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686,
    n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695,
    n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704,
    n24705, n24706, n24707, n24708, n24710, n24711, n24712, n24713, n24714,
    n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
    n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732,
    n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741,
    n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750,
    n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759,
    n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768,
    n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
    n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
    n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
    n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804,
    n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813,
    n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
    n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831,
    n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840,
    n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
    n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
    n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
    n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
    n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885,
    n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894,
    n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
    n24904, n24905, n24906, n24908, n24909, n24910, n24911, n24912, n24913,
    n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
    n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
    n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940,
    n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949,
    n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958,
    n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967,
    n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976,
    n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
    n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
    n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
    n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012,
    n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021,
    n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030,
    n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039,
    n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048,
    n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
    n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
    n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
    n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084,
    n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
    n25094, n25095, n25096, n25097, n25099, n25100, n25101, n25102, n25103,
    n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112,
    n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
    n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
    n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
    n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148,
    n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157,
    n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166,
    n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175,
    n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184,
    n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
    n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
    n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
    n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220,
    n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229,
    n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238,
    n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247,
    n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256,
    n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
    n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
    n25275, n25276, n25277, n25278, n25280, n25281, n25282, n25283, n25284,
    n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293,
    n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302,
    n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311,
    n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320,
    n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
    n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
    n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
    n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356,
    n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365,
    n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374,
    n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383,
    n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392,
    n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
    n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
    n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
    n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428,
    n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437,
    n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446,
    n25447, n25448, n25449, n25450, n25452, n25453, n25454, n25455, n25456,
    n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
    n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
    n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
    n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492,
    n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501,
    n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510,
    n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528,
    n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
    n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
    n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564,
    n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573,
    n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582,
    n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591,
    n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600,
    n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
    n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
    n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
    n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636,
    n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25647, n25648, n25649, n25651, n25652, n25653, n25654, n25655,
    n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664,
    n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
    n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
    n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
    n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700,
    n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709,
    n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718,
    n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727,
    n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736,
    n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
    n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
    n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
    n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772,
    n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781,
    n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790,
    n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799,
    n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808,
    n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25817, n25818,
    n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
    n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836,
    n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845,
    n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854,
    n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863,
    n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872,
    n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
    n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
    n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
    n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908,
    n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917,
    n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926,
    n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935,
    n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944,
    n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25954,
    n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
    n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972,
    n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981,
    n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990,
    n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999,
    n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008,
    n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
    n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
    n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
    n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044,
    n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053,
    n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062,
    n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071,
    n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080,
    n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
    n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
    n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26108,
    n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
    n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126,
    n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
    n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
    n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
    n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
    n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
    n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180,
    n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189,
    n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
    n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207,
    n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
    n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
    n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
    n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
    n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252,
    n26253, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262,
    n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271,
    n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280,
    n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
    n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
    n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
    n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316,
    n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325,
    n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334,
    n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343,
    n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
    n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
    n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
    n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26380,
    n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398,
    n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
    n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
    n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
    n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452,
    n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461,
    n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470,
    n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479,
    n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488,
    n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
    n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
    n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26515, n26516,
    n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525,
    n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534,
    n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
    n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552,
    n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
    n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
    n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
    n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588,
    n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597,
    n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606,
    n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615,
    n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624,
    n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
    n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
    n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652,
    n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661,
    n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670,
    n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679,
    n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688,
    n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
    n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
    n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715,
    n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724,
    n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733,
    n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742,
    n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751,
    n26752, n26753, n26754, n26755, n26756, n26758, n26759, n26760, n26761,
    n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
    n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
    n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788,
    n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
    n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806,
    n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815,
    n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824,
    n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
    n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
    n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
    n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860,
    n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
    n26870, n26871, n26872, n26873, n26875, n26876, n26877, n26878, n26879,
    n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888,
    n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
    n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
    n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
    n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924,
    n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933,
    n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942,
    n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951,
    n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960,
    n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
    n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
    n26979, n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988,
    n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997,
    n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006,
    n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015,
    n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024,
    n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
    n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
    n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
    n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060,
    n27061, n27062, n27063, n27064, n27067, n27070, n27071, n27072, n27073,
    n27074, n27075, n27077, n27084, n27085, n27086, n27087, n27088, n27089,
    n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
    n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
    n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
    n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125,
    n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
    n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
    n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
    n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
    n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
    n27171, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180,
    n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189,
    n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198,
    n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207,
    n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216,
    n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
    n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
    n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
    n27245, n27246, n27247, n27249, n27250, n27251, n27252, n27253, n27254,
    n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263,
    n27264, n27265, n27266, n27268, n27269, n27270, n27271, n27272, n27273,
    n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
    n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
    n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300,
    n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309,
    n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318,
    n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327,
    n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336,
    n27337, n27340, n27343, n27344, n27345, n27346, n27347, n27348, n27350,
    n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365,
    n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374,
    n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
    n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
    n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
    n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
    n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
    n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
    n27429, n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438,
    n27439, n27441, n27442, n27443, n27445, n27446, n27447, n27448, n27449,
    n27450, n27451, n27452, n27453, n27456, n27457, n27458, n27459, n27460,
    n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
    n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478,
    n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487,
    n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496,
    n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
    n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
    n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524,
    n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533,
    n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542,
    n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551,
    n27552, n27553, n27554, n27555, n27556, n27557, n27560, n27563, n27564,
    n27565, n27566, n27567, n27568, n27570, n27571, n27572, n27573, n27574,
    n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583,
    n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592,
    n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
    n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616,
    n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27625, n27626,
    n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
    n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644,
    n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
    n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662,
    n27663, n27664, n27665, n27666, n27667, n27668;
  jnot g00000(.din(\a[5] ), .dout(n64));
  jxor g00001(.dina(\a[3] ), .dinb(\a[2] ), .dout(n65));
  jxor g00002(.dina(\a[5] ), .dinb(\a[4] ), .dout(n66));
  jand g00003(.dina(n66), .dinb(n65), .dout(n67));
  jnot g00004(.din(\a[26] ), .dout(n68));
  jnot g00005(.din(\a[25] ), .dout(n69));
  jxor g00006(.dina(\a[26] ), .dinb(n69), .dout(n70));
  jnot g00007(.din(n70), .dout(n71));
  jnot g00008(.din(\a[23] ), .dout(n72));
  jxor g00009(.dina(\a[24] ), .dinb(n72), .dout(n73));
  jnot g00010(.din(n73), .dout(n74));
  jand g00011(.dina(n74), .dinb(n71), .dout(n75));
  jor  g00012(.dina(\a[30] ), .dinb(\a[29] ), .dout(n76));
  jor  g00013(.dina(\a[28] ), .dinb(\a[27] ), .dout(n77));
  jor  g00014(.dina(n77), .dinb(n76), .dout(n78));
  jor  g00015(.dina(\a[25] ), .dinb(\a[24] ), .dout(n79));
  jor  g00016(.dina(n68), .dinb(\a[23] ), .dout(n80));
  jor  g00017(.dina(n80), .dinb(n79), .dout(n81));
  jor  g00018(.dina(n81), .dinb(n78), .dout(n82));
  jor  g00019(.dina(\a[26] ), .dinb(n72), .dout(n83));
  jor  g00020(.dina(n69), .dinb(\a[24] ), .dout(n84));
  jor  g00021(.dina(n84), .dinb(n83), .dout(n85));
  jnot g00022(.din(\a[28] ), .dout(n86));
  jor  g00023(.dina(n86), .dinb(\a[27] ), .dout(n87));
  jnot g00024(.din(\a[29] ), .dout(n88));
  jnot g00025(.din(\a[30] ), .dout(n89));
  jor  g00026(.dina(n89), .dinb(n88), .dout(n90));
  jor  g00027(.dina(n90), .dinb(n87), .dout(n91));
  jor  g00028(.dina(n91), .dinb(n85), .dout(n92));
  jand g00029(.dina(n92), .dinb(n82), .dout(n93));
  jnot g00030(.din(\a[24] ), .dout(n94));
  jand g00031(.dina(n69), .dinb(n94), .dout(n95));
  jand g00032(.dina(\a[26] ), .dinb(\a[23] ), .dout(n96));
  jand g00033(.dina(n96), .dinb(n95), .dout(n97));
  jnot g00034(.din(\a[27] ), .dout(n98));
  jand g00035(.dina(n86), .dinb(n98), .dout(n99));
  jand g00036(.dina(n89), .dinb(\a[29] ), .dout(n100));
  jand g00037(.dina(n100), .dinb(n99), .dout(n101));
  jand g00038(.dina(n101), .dinb(n97), .dout(n102));
  jnot g00039(.din(n102), .dout(n103));
  jand g00040(.dina(\a[30] ), .dinb(\a[29] ), .dout(n104));
  jand g00041(.dina(\a[28] ), .dinb(\a[27] ), .dout(n105));
  jand g00042(.dina(n105), .dinb(n104), .dout(n106));
  jand g00043(.dina(n106), .dinb(n97), .dout(n107));
  jnot g00044(.din(n107), .dout(n108));
  jand g00045(.dina(n108), .dinb(n103), .dout(n109));
  jor  g00046(.dina(\a[30] ), .dinb(n88), .dout(n110));
  jor  g00047(.dina(n86), .dinb(n98), .dout(n111));
  jor  g00048(.dina(n111), .dinb(n110), .dout(n112));
  jor  g00049(.dina(n112), .dinb(n81), .dout(n113));
  jand g00050(.dina(\a[25] ), .dinb(n94), .dout(n114));
  jand g00051(.dina(n68), .dinb(n72), .dout(n115));
  jand g00052(.dina(n115), .dinb(n114), .dout(n116));
  jand g00053(.dina(\a[30] ), .dinb(n88), .dout(n117));
  jand g00054(.dina(n117), .dinb(n105), .dout(n118));
  jand g00055(.dina(n118), .dinb(n116), .dout(n119));
  jnot g00056(.din(n119), .dout(n120));
  jand g00057(.dina(n120), .dinb(n113), .dout(n121));
  jand g00058(.dina(n121), .dinb(n109), .dout(n122));
  jand g00059(.dina(n122), .dinb(n93), .dout(n123));
  jand g00060(.dina(n69), .dinb(\a[24] ), .dout(n124));
  jand g00061(.dina(n124), .dinb(n96), .dout(n125));
  jand g00062(.dina(n89), .dinb(n88), .dout(n126));
  jand g00063(.dina(\a[28] ), .dinb(n98), .dout(n127));
  jand g00064(.dina(n127), .dinb(n126), .dout(n128));
  jand g00065(.dina(n128), .dinb(n125), .dout(n129));
  jnot g00066(.din(n129), .dout(n130));
  jand g00067(.dina(\a[26] ), .dinb(n72), .dout(n131));
  jand g00068(.dina(n131), .dinb(n95), .dout(n132));
  jand g00069(.dina(n128), .dinb(n132), .dout(n133));
  jnot g00070(.din(n133), .dout(n134));
  jand g00071(.dina(n125), .dinb(n106), .dout(n135));
  jnot g00072(.din(n135), .dout(n136));
  jand g00073(.dina(n136), .dinb(n134), .dout(n137));
  jand g00074(.dina(n137), .dinb(n130), .dout(n138));
  jor  g00075(.dina(\a[26] ), .dinb(\a[23] ), .dout(n139));
  jor  g00076(.dina(n69), .dinb(n94), .dout(n140));
  jor  g00077(.dina(n140), .dinb(n139), .dout(n141));
  jor  g00078(.dina(n110), .dinb(n87), .dout(n142));
  jor  g00079(.dina(n142), .dinb(n141), .dout(n143));
  jor  g00080(.dina(n68), .dinb(n72), .dout(n144));
  jor  g00081(.dina(n140), .dinb(n144), .dout(n145));
  jor  g00082(.dina(n145), .dinb(n78), .dout(n146));
  jand g00083(.dina(n105), .dinb(n100), .dout(n147));
  jand g00084(.dina(n125), .dinb(n147), .dout(n148));
  jnot g00085(.din(n148), .dout(n149));
  jand g00086(.dina(n149), .dinb(n146), .dout(n150));
  jand g00087(.dina(n150), .dinb(n143), .dout(n151));
  jor  g00088(.dina(n111), .dinb(n76), .dout(n152));
  jor  g00089(.dina(n144), .dinb(n84), .dout(n153));
  jor  g00090(.dina(n153), .dinb(n152), .dout(n154));
  jand g00091(.dina(n124), .dinb(n115), .dout(n155));
  jand g00092(.dina(n155), .dinb(n118), .dout(n156));
  jnot g00093(.din(n156), .dout(n157));
  jand g00094(.dina(n157), .dinb(n154), .dout(n158));
  jand g00095(.dina(n114), .dinb(n131), .dout(n159));
  jand g00096(.dina(n159), .dinb(n101), .dout(n160));
  jnot g00097(.din(n160), .dout(n161));
  jor  g00098(.dina(n140), .dinb(n80), .dout(n162));
  jor  g00099(.dina(\a[28] ), .dinb(n98), .dout(n163));
  jor  g00100(.dina(n163), .dinb(n90), .dout(n164));
  jor  g00101(.dina(n164), .dinb(n162), .dout(n165));
  jand g00102(.dina(n165), .dinb(n161), .dout(n166));
  jand g00103(.dina(n166), .dinb(n158), .dout(n167));
  jand g00104(.dina(n167), .dinb(n151), .dout(n168));
  jand g00105(.dina(n168), .dinb(n138), .dout(n169));
  jand g00106(.dina(n169), .dinb(n123), .dout(n170));
  jand g00107(.dina(n86), .dinb(\a[27] ), .dout(n171));
  jand g00108(.dina(n171), .dinb(n104), .dout(n172));
  jand g00109(.dina(n172), .dinb(n132), .dout(n173));
  jnot g00110(.din(n173), .dout(n174));
  jor  g00111(.dina(n89), .dinb(\a[29] ), .dout(n175));
  jor  g00112(.dina(n175), .dinb(n77), .dout(n176));
  jor  g00113(.dina(n176), .dinb(n141), .dout(n177));
  jand g00114(.dina(n177), .dinb(n174), .dout(n178));
  jand g00115(.dina(n155), .dinb(n147), .dout(n179));
  jnot g00116(.din(n179), .dout(n180));
  jand g00117(.dina(\a[25] ), .dinb(\a[24] ), .dout(n181));
  jand g00118(.dina(n181), .dinb(n96), .dout(n182));
  jand g00119(.dina(n182), .dinb(n106), .dout(n183));
  jnot g00120(.din(n183), .dout(n184));
  jand g00121(.dina(n184), .dinb(n180), .dout(n185));
  jand g00122(.dina(n185), .dinb(n178), .dout(n186));
  jor  g00123(.dina(\a[25] ), .dinb(n94), .dout(n187));
  jor  g00124(.dina(n187), .dinb(n80), .dout(n188));
  jor  g00125(.dina(n163), .dinb(n110), .dout(n189));
  jor  g00126(.dina(n189), .dinb(n188), .dout(n190));
  jand g00127(.dina(n68), .dinb(\a[23] ), .dout(n191));
  jand g00128(.dina(n124), .dinb(n191), .dout(n192));
  jand g00129(.dina(n192), .dinb(n101), .dout(n193));
  jnot g00130(.din(n193), .dout(n194));
  jand g00131(.dina(n115), .dinb(n95), .dout(n195));
  jand g00132(.dina(n195), .dinb(n118), .dout(n196));
  jnot g00133(.din(n196), .dout(n197));
  jand g00134(.dina(n197), .dinb(n194), .dout(n198));
  jand g00135(.dina(n198), .dinb(n190), .dout(n199));
  jand g00136(.dina(n100), .dinb(n127), .dout(n200));
  jand g00137(.dina(n182), .dinb(n200), .dout(n201));
  jnot g00138(.din(n201), .dout(n202));
  jand g00139(.dina(n104), .dinb(n127), .dout(n203));
  jand g00140(.dina(n116), .dinb(n203), .dout(n204));
  jnot g00141(.din(n204), .dout(n205));
  jor  g00142(.dina(n140), .dinb(n83), .dout(n206));
  jor  g00143(.dina(n163), .dinb(n76), .dout(n207));
  jor  g00144(.dina(n207), .dinb(n206), .dout(n208));
  jand g00145(.dina(n208), .dinb(n205), .dout(n209));
  jand g00146(.dina(n209), .dinb(n202), .dout(n210));
  jand g00147(.dina(n210), .dinb(n199), .dout(n211));
  jand g00148(.dina(n211), .dinb(n186), .dout(n212));
  jor  g00149(.dina(n84), .dinb(n80), .dout(n213));
  jor  g00150(.dina(n213), .dinb(n112), .dout(n214));
  jand g00151(.dina(n181), .dinb(n131), .dout(n215));
  jand g00152(.dina(n215), .dinb(n147), .dout(n216));
  jnot g00153(.din(n216), .dout(n217));
  jand g00154(.dina(n217), .dinb(n214), .dout(n218));
  jand g00155(.dina(n181), .dinb(n115), .dout(n219));
  jand g00156(.dina(n172), .dinb(n219), .dout(n220));
  jnot g00157(.din(n220), .dout(n221));
  jand g00158(.dina(n104), .dinb(n99), .dout(n222));
  jand g00159(.dina(n222), .dinb(n132), .dout(n223));
  jnot g00160(.din(n223), .dout(n224));
  jand g00161(.dina(n224), .dinb(n221), .dout(n225));
  jand g00162(.dina(n225), .dinb(n218), .dout(n226));
  jand g00163(.dina(n195), .dinb(n200), .dout(n227));
  jnot g00164(.din(n227), .dout(n228));
  jand g00165(.dina(n128), .dinb(n97), .dout(n229));
  jnot g00166(.din(n229), .dout(n230));
  jand g00167(.dina(n230), .dinb(n228), .dout(n231));
  jand g00168(.dina(n171), .dinb(n100), .dout(n232));
  jand g00169(.dina(n232), .dinb(n159), .dout(n233));
  jnot g00170(.din(n233), .dout(n234));
  jand g00171(.dina(n191), .dinb(n95), .dout(n235));
  jand g00172(.dina(n117), .dinb(n127), .dout(n236));
  jand g00173(.dina(n236), .dinb(n235), .dout(n237));
  jnot g00174(.din(n237), .dout(n238));
  jand g00175(.dina(n238), .dinb(n234), .dout(n239));
  jand g00176(.dina(n239), .dinb(n231), .dout(n240));
  jand g00177(.dina(n240), .dinb(n226), .dout(n241));
  jand g00178(.dina(n232), .dinb(n155), .dout(n242));
  jnot g00179(.din(n242), .dout(n243));
  jor  g00180(.dina(n187), .dinb(n139), .dout(n244));
  jor  g00181(.dina(n244), .dinb(n142), .dout(n245));
  jand g00182(.dina(n245), .dinb(n243), .dout(n246));
  jnot g00183(.din(n78), .dout(n247));
  jand g00184(.dina(n219), .dinb(n247), .dout(n248));
  jnot g00185(.din(n248), .dout(n249));
  jand g00186(.dina(n124), .dinb(n131), .dout(n250));
  jand g00187(.dina(n222), .dinb(n250), .dout(n251));
  jnot g00188(.din(n251), .dout(n252));
  jand g00189(.dina(n252), .dinb(n249), .dout(n253));
  jand g00190(.dina(n253), .dinb(n246), .dout(n254));
  jor  g00191(.dina(n162), .dinb(n142), .dout(n255));
  jor  g00192(.dina(n139), .dinb(n79), .dout(n256));
  jor  g00193(.dina(n207), .dinb(n256), .dout(n257));
  jand g00194(.dina(n257), .dinb(n255), .dout(n258));
  jor  g00195(.dina(n90), .dinb(n77), .dout(n259));
  jor  g00196(.dina(n259), .dinb(n145), .dout(n260));
  jand g00197(.dina(n182), .dinb(n147), .dout(n261));
  jnot g00198(.din(n261), .dout(n262));
  jand g00199(.dina(n262), .dinb(n260), .dout(n263));
  jand g00200(.dina(n263), .dinb(n258), .dout(n264));
  jand g00201(.dina(n264), .dinb(n254), .dout(n265));
  jand g00202(.dina(n265), .dinb(n241), .dout(n266));
  jand g00203(.dina(n219), .dinb(n147), .dout(n267));
  jnot g00204(.din(n267), .dout(n268));
  jor  g00205(.dina(n175), .dinb(n87), .dout(n269));
  jor  g00206(.dina(n269), .dinb(n85), .dout(n270));
  jand g00207(.dina(n270), .dinb(n268), .dout(n271));
  jand g00208(.dina(n181), .dinb(n191), .dout(n272));
  jand g00209(.dina(n272), .dinb(n101), .dout(n273));
  jnot g00210(.din(n273), .dout(n274));
  jor  g00211(.dina(n110), .dinb(n77), .dout(n275));
  jor  g00212(.dina(n145), .dinb(n275), .dout(n276));
  jand g00213(.dina(n276), .dinb(n274), .dout(n277));
  jand g00214(.dina(n171), .dinb(n126), .dout(n278));
  jand g00215(.dina(n278), .dinb(n192), .dout(n279));
  jnot g00216(.din(n279), .dout(n280));
  jand g00217(.dina(n280), .dinb(n277), .dout(n281));
  jand g00218(.dina(n281), .dinb(n271), .dout(n282));
  jand g00219(.dina(n128), .dinb(n116), .dout(n283));
  jnot g00220(.din(n283), .dout(n284));
  jor  g00221(.dina(n187), .dinb(n144), .dout(n285));
  jor  g00222(.dina(n164), .dinb(n285), .dout(n286));
  jand g00223(.dina(n286), .dinb(n284), .dout(n287));
  jor  g00224(.dina(n207), .dinb(n213), .dout(n288));
  jand g00225(.dina(n219), .dinb(n101), .dout(n289));
  jnot g00226(.din(n289), .dout(n290));
  jand g00227(.dina(n215), .dinb(n203), .dout(n291));
  jnot g00228(.din(n291), .dout(n292));
  jand g00229(.dina(n292), .dinb(n290), .dout(n293));
  jand g00230(.dina(n293), .dinb(n288), .dout(n294));
  jand g00231(.dina(n294), .dinb(n287), .dout(n295));
  jand g00232(.dina(n295), .dinb(n282), .dout(n296));
  jand g00233(.dina(n296), .dinb(n266), .dout(n297));
  jand g00234(.dina(n297), .dinb(n212), .dout(n298));
  jand g00235(.dina(n298), .dinb(n170), .dout(n299));
  jand g00236(.dina(n114), .dinb(n191), .dout(n300));
  jand g00237(.dina(n300), .dinb(n247), .dout(n301));
  jnot g00238(.din(n301), .dout(n302));
  jand g00239(.dina(n215), .dinb(n101), .dout(n303));
  jnot g00240(.din(n303), .dout(n304));
  jor  g00241(.dina(n188), .dinb(n275), .dout(n305));
  jand g00242(.dina(n305), .dinb(n304), .dout(n306));
  jand g00243(.dina(n306), .dinb(n302), .dout(n307));
  jand g00244(.dina(n106), .dinb(n300), .dout(n308));
  jnot g00245(.din(n308), .dout(n309));
  jor  g00246(.dina(n163), .dinb(n175), .dout(n310));
  jor  g00247(.dina(n310), .dinb(n285), .dout(n311));
  jand g00248(.dina(n311), .dinb(n309), .dout(n312));
  jand g00249(.dina(n219), .dinb(n118), .dout(n313));
  jnot g00250(.din(n313), .dout(n314));
  jand g00251(.dina(n96), .dinb(n114), .dout(n315));
  jand g00252(.dina(n222), .dinb(n315), .dout(n316));
  jnot g00253(.din(n316), .dout(n317));
  jand g00254(.dina(n317), .dinb(n314), .dout(n318));
  jand g00255(.dina(n318), .dinb(n312), .dout(n319));
  jand g00256(.dina(n319), .dinb(n307), .dout(n320));
  jand g00257(.dina(n125), .dinb(n101), .dout(n321));
  jnot g00258(.din(n321), .dout(n322));
  jand g00259(.dina(n278), .dinb(n250), .dout(n323));
  jnot g00260(.din(n323), .dout(n324));
  jor  g00261(.dina(n269), .dinb(n145), .dout(n325));
  jand g00262(.dina(n325), .dinb(n324), .dout(n326));
  jand g00263(.dina(n326), .dinb(n322), .dout(n327));
  jand g00264(.dina(n125), .dinb(n203), .dout(n328));
  jnot g00265(.din(n328), .dout(n329));
  jor  g00266(.dina(n310), .dinb(n256), .dout(n330));
  jor  g00267(.dina(n206), .dinb(n176), .dout(n331));
  jand g00268(.dina(n331), .dinb(n330), .dout(n332));
  jand g00269(.dina(n332), .dinb(n329), .dout(n333));
  jand g00270(.dina(n333), .dinb(n327), .dout(n334));
  jand g00271(.dina(n334), .dinb(n320), .dout(n335));
  jor  g00272(.dina(n310), .dinb(n145), .dout(n336));
  jor  g00273(.dina(n310), .dinb(n244), .dout(n337));
  jand g00274(.dina(n171), .dinb(n117), .dout(n338));
  jand g00275(.dina(n338), .dinb(n315), .dout(n339));
  jnot g00276(.din(n339), .dout(n340));
  jand g00277(.dina(n340), .dinb(n337), .dout(n341));
  jand g00278(.dina(n341), .dinb(n336), .dout(n342));
  jor  g00279(.dina(n142), .dinb(n285), .dout(n343));
  jand g00280(.dina(n105), .dinb(n126), .dout(n344));
  jand g00281(.dina(n155), .dinb(n344), .dout(n345));
  jnot g00282(.din(n345), .dout(n346));
  jor  g00283(.dina(n83), .dinb(n79), .dout(n347));
  jor  g00284(.dina(n347), .dinb(n176), .dout(n348));
  jand g00285(.dina(n348), .dinb(n346), .dout(n349));
  jand g00286(.dina(n349), .dinb(n343), .dout(n350));
  jand g00287(.dina(n272), .dinb(n247), .dout(n351));
  jnot g00288(.din(n351), .dout(n352));
  jand g00289(.dina(n101), .dinb(n300), .dout(n353));
  jnot g00290(.din(n353), .dout(n354));
  jand g00291(.dina(n354), .dinb(n352), .dout(n355));
  jor  g00292(.dina(n87), .dinb(n76), .dout(n356));
  jor  g00293(.dina(n141), .dinb(n356), .dout(n357));
  jand g00294(.dina(n222), .dinb(n195), .dout(n358));
  jnot g00295(.din(n358), .dout(n359));
  jand g00296(.dina(n359), .dinb(n357), .dout(n360));
  jand g00297(.dina(n360), .dinb(n355), .dout(n361));
  jand g00298(.dina(n361), .dinb(n350), .dout(n362));
  jand g00299(.dina(n362), .dinb(n342), .dout(n363));
  jor  g00300(.dina(n144), .dinb(n79), .dout(n364));
  jor  g00301(.dina(n189), .dinb(n364), .dout(n365));
  jor  g00302(.dina(n112), .dinb(n85), .dout(n366));
  jor  g00303(.dina(n256), .dinb(n356), .dout(n367));
  jand g00304(.dina(n367), .dinb(n366), .dout(n368));
  jand g00305(.dina(n368), .dinb(n365), .dout(n369));
  jor  g00306(.dina(n111), .dinb(n90), .dout(n370));
  jor  g00307(.dina(n244), .dinb(n370), .dout(n371));
  jor  g00308(.dina(n310), .dinb(n364), .dout(n372));
  jand g00309(.dina(n372), .dinb(n371), .dout(n373));
  jand g00310(.dina(n222), .dinb(n192), .dout(n374));
  jnot g00311(.din(n374), .dout(n375));
  jand g00312(.dina(n236), .dinb(n125), .dout(n376));
  jnot g00313(.din(n376), .dout(n377));
  jand g00314(.dina(n377), .dinb(n375), .dout(n378));
  jand g00315(.dina(n378), .dinb(n373), .dout(n379));
  jand g00316(.dina(n379), .dinb(n369), .dout(n380));
  jand g00317(.dina(n195), .dinb(n232), .dout(n381));
  jnot g00318(.din(n381), .dout(n382));
  jor  g00319(.dina(n164), .dinb(n85), .dout(n383));
  jand g00320(.dina(n383), .dinb(n382), .dout(n384));
  jor  g00321(.dina(n206), .dinb(n91), .dout(n385));
  jor  g00322(.dina(n164), .dinb(n244), .dout(n386));
  jand g00323(.dina(n386), .dinb(n385), .dout(n387));
  jand g00324(.dina(n387), .dinb(n384), .dout(n388));
  jand g00325(.dina(n117), .dinb(n99), .dout(n389));
  jand g00326(.dina(n389), .dinb(n215), .dout(n390));
  jnot g00327(.din(n390), .dout(n391));
  jor  g00328(.dina(n269), .dinb(n153), .dout(n392));
  jand g00329(.dina(n392), .dinb(n391), .dout(n393));
  jor  g00330(.dina(n139), .dinb(n84), .dout(n394));
  jor  g00331(.dina(n176), .dinb(n394), .dout(n395));
  jor  g00332(.dina(n269), .dinb(n364), .dout(n396));
  jand g00333(.dina(n396), .dinb(n395), .dout(n397));
  jand g00334(.dina(n397), .dinb(n393), .dout(n398));
  jand g00335(.dina(n398), .dinb(n388), .dout(n399));
  jand g00336(.dina(n399), .dinb(n380), .dout(n400));
  jand g00337(.dina(n400), .dinb(n363), .dout(n401));
  jand g00338(.dina(n401), .dinb(n335), .dout(n402));
  jand g00339(.dina(n159), .dinb(n128), .dout(n403));
  jnot g00340(.din(n403), .dout(n404));
  jor  g00341(.dina(n310), .dinb(n206), .dout(n405));
  jand g00342(.dina(n405), .dinb(n404), .dout(n406));
  jor  g00343(.dina(n142), .dinb(n85), .dout(n407));
  jand g00344(.dina(n236), .dinb(n192), .dout(n408));
  jnot g00345(.din(n408), .dout(n409));
  jand g00346(.dina(n409), .dinb(n407), .dout(n410));
  jand g00347(.dina(n410), .dinb(n406), .dout(n411));
  jand g00348(.dina(n192), .dinb(n232), .dout(n412));
  jnot g00349(.din(n412), .dout(n413));
  jor  g00350(.dina(n259), .dinb(n206), .dout(n414));
  jand g00351(.dina(n414), .dinb(n413), .dout(n415));
  jor  g00352(.dina(n175), .dinb(n111), .dout(n416));
  jor  g00353(.dina(n162), .dinb(n416), .dout(n417));
  jor  g00354(.dina(n188), .dinb(n91), .dout(n418));
  jand g00355(.dina(n418), .dinb(n417), .dout(n419));
  jand g00356(.dina(n419), .dinb(n415), .dout(n420));
  jand g00357(.dina(n420), .dinb(n411), .dout(n421));
  jand g00358(.dina(n182), .dinb(n128), .dout(n422));
  jnot g00359(.din(n422), .dout(n423));
  jor  g00360(.dina(n416), .dinb(n364), .dout(n424));
  jand g00361(.dina(n424), .dinb(n423), .dout(n425));
  jand g00362(.dina(n192), .dinb(n172), .dout(n426));
  jnot g00363(.din(n426), .dout(n427));
  jor  g00364(.dina(n310), .dinb(n85), .dout(n428));
  jand g00365(.dina(n428), .dinb(n427), .dout(n429));
  jand g00366(.dina(n429), .dinb(n425), .dout(n430));
  jor  g00367(.dina(n275), .dinb(n81), .dout(n431));
  jor  g00368(.dina(n394), .dinb(n275), .dout(n432));
  jand g00369(.dina(n432), .dinb(n431), .dout(n433));
  jor  g00370(.dina(n347), .dinb(n189), .dout(n434));
  jor  g00371(.dina(n244), .dinb(n356), .dout(n435));
  jand g00372(.dina(n435), .dinb(n434), .dout(n436));
  jand g00373(.dina(n436), .dinb(n433), .dout(n437));
  jand g00374(.dina(n437), .dinb(n430), .dout(n438));
  jor  g00375(.dina(n188), .dinb(n142), .dout(n439));
  jand g00376(.dina(n159), .dinb(n106), .dout(n440));
  jnot g00377(.din(n440), .dout(n441));
  jand g00378(.dina(n441), .dinb(n439), .dout(n442));
  jor  g00379(.dina(n347), .dinb(n370), .dout(n443));
  jand g00380(.dina(n125), .dinb(n118), .dout(n444));
  jnot g00381(.din(n444), .dout(n445));
  jand g00382(.dina(n445), .dinb(n443), .dout(n446));
  jand g00383(.dina(n446), .dinb(n442), .dout(n447));
  jand g00384(.dina(n315), .dinb(n101), .dout(n448));
  jnot g00385(.din(n448), .dout(n449));
  jor  g00386(.dina(n259), .dinb(n85), .dout(n450));
  jand g00387(.dina(n450), .dinb(n449), .dout(n451));
  jand g00388(.dina(n159), .dinb(n344), .dout(n452));
  jand g00389(.dina(n215), .dinb(n247), .dout(n453));
  jor  g00390(.dina(n453), .dinb(n452), .dout(n454));
  jnot g00391(.din(n454), .dout(n455));
  jand g00392(.dina(n455), .dinb(n451), .dout(n456));
  jand g00393(.dina(n456), .dinb(n447), .dout(n457));
  jand g00394(.dina(n457), .dinb(n438), .dout(n458));
  jand g00395(.dina(n458), .dinb(n421), .dout(n459));
  jand g00396(.dina(n344), .dinb(n125), .dout(n460));
  jnot g00397(.din(n460), .dout(n461));
  jor  g00398(.dina(n152), .dinb(n141), .dout(n462));
  jand g00399(.dina(n462), .dinb(n461), .dout(n463));
  jand g00400(.dina(n235), .dinb(n203), .dout(n464));
  jnot g00401(.din(n464), .dout(n465));
  jand g00402(.dina(n278), .dinb(n97), .dout(n466));
  jnot g00403(.din(n466), .dout(n467));
  jand g00404(.dina(n467), .dinb(n465), .dout(n468));
  jand g00405(.dina(n235), .dinb(n200), .dout(n469));
  jnot g00406(.din(n469), .dout(n470));
  jand g00407(.dina(n278), .dinb(n219), .dout(n471));
  jnot g00408(.din(n471), .dout(n472));
  jand g00409(.dina(n472), .dinb(n470), .dout(n473));
  jand g00410(.dina(n473), .dinb(n468), .dout(n474));
  jand g00411(.dina(n474), .dinb(n463), .dout(n475));
  jor  g00412(.dina(n153), .dinb(n416), .dout(n476));
  jand g00413(.dina(n222), .dinb(n155), .dout(n477));
  jnot g00414(.din(n477), .dout(n478));
  jand g00415(.dina(n478), .dinb(n476), .dout(n479));
  jand g00416(.dina(n195), .dinb(n172), .dout(n480));
  jnot g00417(.din(n480), .dout(n481));
  jand g00418(.dina(n278), .dinb(n116), .dout(n482));
  jnot g00419(.din(n482), .dout(n483));
  jand g00420(.dina(n483), .dinb(n481), .dout(n484));
  jand g00421(.dina(n484), .dinb(n479), .dout(n485));
  jor  g00422(.dina(n206), .dinb(n152), .dout(n486));
  jnot g00423(.din(n486), .dout(n487));
  jand g00424(.dina(n203), .dinb(n132), .dout(n488));
  jor  g00425(.dina(n488), .dinb(n487), .dout(n489));
  jnot g00426(.din(n489), .dout(n490));
  jand g00427(.dina(n106), .dinb(n132), .dout(n491));
  jnot g00428(.din(n491), .dout(n492));
  jand g00429(.dina(n278), .dinb(n215), .dout(n493));
  jnot g00430(.din(n493), .dout(n494));
  jand g00431(.dina(n494), .dinb(n492), .dout(n495));
  jand g00432(.dina(n495), .dinb(n490), .dout(n496));
  jand g00433(.dina(n496), .dinb(n485), .dout(n497));
  jand g00434(.dina(n497), .dinb(n475), .dout(n498));
  jor  g00435(.dina(n176), .dinb(n213), .dout(n499));
  jor  g00436(.dina(n176), .dinb(n364), .dout(n500));
  jand g00437(.dina(n500), .dinb(n499), .dout(n501));
  jand g00438(.dina(n236), .dinb(n272), .dout(n502));
  jnot g00439(.din(n502), .dout(n503));
  jand g00440(.dina(n338), .dinb(n192), .dout(n504));
  jnot g00441(.din(n504), .dout(n505));
  jand g00442(.dina(n505), .dinb(n503), .dout(n506));
  jand g00443(.dina(n506), .dinb(n501), .dout(n507));
  jor  g00444(.dina(n189), .dinb(n285), .dout(n508));
  jor  g00445(.dina(n162), .dinb(n356), .dout(n509));
  jand g00446(.dina(n389), .dinb(n125), .dout(n510));
  jnot g00447(.din(n510), .dout(n511));
  jand g00448(.dina(n511), .dinb(n509), .dout(n512));
  jand g00449(.dina(n512), .dinb(n508), .dout(n513));
  jand g00450(.dina(n147), .dinb(n97), .dout(n514));
  jnot g00451(.din(n514), .dout(n515));
  jor  g00452(.dina(n206), .dinb(n142), .dout(n516));
  jor  g00453(.dina(n394), .dinb(n370), .dout(n517));
  jand g00454(.dina(n517), .dinb(n516), .dout(n518));
  jand g00455(.dina(n518), .dinb(n515), .dout(n519));
  jand g00456(.dina(n519), .dinb(n513), .dout(n520));
  jand g00457(.dina(n520), .dinb(n507), .dout(n521));
  jand g00458(.dina(n521), .dinb(n498), .dout(n522));
  jand g00459(.dina(n522), .dinb(n459), .dout(n523));
  jand g00460(.dina(n523), .dinb(n402), .dout(n524));
  jand g00461(.dina(n524), .dinb(n299), .dout(n525));
  jnot g00462(.din(n525), .dout(n526));
  jor  g00463(.dina(n189), .dinb(n145), .dout(n527));
  jand g00464(.dina(n172), .dinb(n182), .dout(n528));
  jnot g00465(.din(n528), .dout(n529));
  jand g00466(.dina(n529), .dinb(n439), .dout(n530));
  jand g00467(.dina(n530), .dinb(n527), .dout(n531));
  jor  g00468(.dina(n162), .dinb(n152), .dout(n532));
  jor  g00469(.dina(n310), .dinb(n213), .dout(n533));
  jand g00470(.dina(n533), .dinb(n532), .dout(n534));
  jor  g00471(.dina(n187), .dinb(n83), .dout(n535));
  jor  g00472(.dina(n535), .dinb(n176), .dout(n536));
  jand g00473(.dina(n536), .dinb(n395), .dout(n537));
  jand g00474(.dina(n428), .dinb(n304), .dout(n538));
  jand g00475(.dina(n538), .dinb(n537), .dout(n539));
  jand g00476(.dina(n539), .dinb(n534), .dout(n540));
  jand g00477(.dina(n540), .dinb(n531), .dout(n541));
  jor  g00478(.dina(n259), .dinb(n394), .dout(n542));
  jor  g00479(.dina(n256), .dinb(n91), .dout(n543));
  jand g00480(.dina(n543), .dinb(n542), .dout(n544));
  jand g00481(.dina(n338), .dinb(n132), .dout(n545));
  jor  g00482(.dina(n545), .dinb(n471), .dout(n546));
  jnot g00483(.din(n546), .dout(n547));
  jand g00484(.dina(n208), .dinb(n136), .dout(n548));
  jand g00485(.dina(n548), .dinb(n547), .dout(n549));
  jand g00486(.dina(n549), .dinb(n544), .dout(n550));
  jor  g00487(.dina(n310), .dinb(n347), .dout(n551));
  jand g00488(.dina(n551), .dinb(n396), .dout(n552));
  jor  g00489(.dina(n213), .dinb(n91), .dout(n553));
  jand g00490(.dina(n553), .dinb(n348), .dout(n554));
  jand g00491(.dina(n554), .dinb(n552), .dout(n555));
  jand g00492(.dina(n315), .dinb(n203), .dout(n556));
  jnot g00493(.din(n556), .dout(n557));
  jand g00494(.dina(n557), .dinb(n202), .dout(n558));
  jand g00495(.dina(n517), .dinb(n314), .dout(n559));
  jand g00496(.dina(n559), .dinb(n558), .dout(n560));
  jand g00497(.dina(n560), .dinb(n555), .dout(n561));
  jor  g00498(.dina(n152), .dinb(n394), .dout(n562));
  jand g00499(.dina(n562), .dinb(n149), .dout(n563));
  jand g00500(.dina(n481), .dinb(n445), .dout(n564));
  jand g00501(.dina(n564), .dinb(n563), .dout(n565));
  jor  g00502(.dina(n347), .dinb(n416), .dout(n566));
  jand g00503(.dina(n566), .dinb(n252), .dout(n567));
  jand g00504(.dina(n567), .dinb(n260), .dout(n568));
  jand g00505(.dina(n568), .dinb(n565), .dout(n569));
  jand g00506(.dina(n569), .dinb(n561), .dout(n570));
  jand g00507(.dina(n570), .dinb(n550), .dout(n571));
  jand g00508(.dina(n571), .dinb(n541), .dout(n572));
  jand g00509(.dina(n232), .dinb(n132), .dout(n573));
  jnot g00510(.din(n573), .dout(n574));
  jand g00511(.dina(n574), .dinb(n130), .dout(n575));
  jand g00512(.dina(n367), .dinb(n238), .dout(n576));
  jand g00513(.dina(n576), .dinb(n575), .dout(n577));
  jor  g00514(.dina(n206), .dinb(n112), .dout(n578));
  jand g00515(.dina(n578), .dinb(n366), .dout(n579));
  jand g00516(.dina(n579), .dinb(n433), .dout(n580));
  jand g00517(.dina(n580), .dinb(n577), .dout(n581));
  jand g00518(.dina(n172), .dinb(n97), .dout(n582));
  jnot g00519(.din(n582), .dout(n583));
  jand g00520(.dina(n583), .dinb(n391), .dout(n584));
  jand g00521(.dina(n584), .dinb(n461), .dout(n585));
  jor  g00522(.dina(n153), .dinb(n112), .dout(n586));
  jand g00523(.dina(n586), .dinb(n221), .dout(n587));
  jand g00524(.dina(n587), .dinb(n382), .dout(n588));
  jand g00525(.dina(n588), .dinb(n585), .dout(n589));
  jand g00526(.dina(n589), .dinb(n581), .dout(n590));
  jand g00527(.dina(n590), .dinb(n572), .dout(n591));
  jand g00528(.dina(n200), .dinb(n97), .dout(n592));
  jor  g00529(.dina(n592), .dinb(n510), .dout(n593));
  jnot g00530(.din(n593), .dout(n594));
  jor  g00531(.dina(n207), .dinb(n153), .dout(n595));
  jand g00532(.dina(n595), .dinb(n509), .dout(n596));
  jand g00533(.dina(n236), .dinb(n300), .dout(n597));
  jor  g00534(.dina(n347), .dinb(n152), .dout(n598));
  jnot g00535(.din(n598), .dout(n599));
  jor  g00536(.dina(n599), .dinb(n597), .dout(n600));
  jnot g00537(.din(n600), .dout(n601));
  jand g00538(.dina(n601), .dinb(n596), .dout(n602));
  jand g00539(.dina(n602), .dinb(n594), .dout(n603));
  jand g00540(.dina(n116), .dinb(n147), .dout(n604));
  jnot g00541(.din(n604), .dout(n605));
  jand g00542(.dina(n605), .dinb(n113), .dout(n606));
  jor  g00543(.dina(n152), .dinb(n364), .dout(n607));
  jand g00544(.dina(n250), .dinb(n106), .dout(n608));
  jnot g00545(.din(n608), .dout(n609));
  jand g00546(.dina(n609), .dinb(n607), .dout(n610));
  jand g00547(.dina(n610), .dinb(n606), .dout(n611));
  jor  g00548(.dina(n189), .dinb(n394), .dout(n612));
  jand g00549(.dina(n612), .dinb(n243), .dout(n613));
  jor  g00550(.dina(n310), .dinb(n394), .dout(n614));
  jand g00551(.dina(n614), .dinb(n331), .dout(n615));
  jand g00552(.dina(n615), .dinb(n613), .dout(n616));
  jand g00553(.dina(n616), .dinb(n611), .dout(n617));
  jand g00554(.dina(n236), .dinb(n195), .dout(n618));
  jnot g00555(.din(n618), .dout(n619));
  jand g00556(.dina(n619), .dinb(n516), .dout(n620));
  jand g00557(.dina(n195), .dinb(n389), .dout(n621));
  jnot g00558(.din(n621), .dout(n622));
  jand g00559(.dina(n622), .dinb(n383), .dout(n623));
  jand g00560(.dina(n623), .dinb(n620), .dout(n624));
  jand g00561(.dina(n118), .dinb(n300), .dout(n625));
  jnot g00562(.din(n625), .dout(n626));
  jand g00563(.dina(n626), .dinb(n217), .dout(n627));
  jand g00564(.dina(n627), .dinb(n180), .dout(n628));
  jand g00565(.dina(n628), .dinb(n624), .dout(n629));
  jand g00566(.dina(n629), .dinb(n617), .dout(n630));
  jand g00567(.dina(n630), .dinb(n603), .dout(n631));
  jand g00568(.dina(n250), .dinb(n118), .dout(n632));
  jnot g00569(.din(n632), .dout(n633));
  jand g00570(.dina(n633), .dinb(n337), .dout(n634));
  jor  g00571(.dina(n145), .dinb(n416), .dout(n635));
  jand g00572(.dina(n635), .dinb(n365), .dout(n636));
  jand g00573(.dina(n465), .dinb(n161), .dout(n637));
  jand g00574(.dina(n637), .dinb(n636), .dout(n638));
  jand g00575(.dina(n638), .dinb(n634), .dout(n639));
  jand g00576(.dina(n222), .dinb(n215), .dout(n640));
  jnot g00577(.din(n640), .dout(n641));
  jand g00578(.dina(n250), .dinb(n147), .dout(n642));
  jnot g00579(.din(n642), .dout(n643));
  jand g00580(.dina(n643), .dinb(n641), .dout(n644));
  jand g00581(.dina(n232), .dinb(n219), .dout(n645));
  jnot g00582(.din(n645), .dout(n646));
  jand g00583(.dina(n646), .dinb(n508), .dout(n647));
  jand g00584(.dina(n462), .dinb(n441), .dout(n648));
  jand g00585(.dina(n648), .dinb(n647), .dout(n649));
  jand g00586(.dina(n649), .dinb(n644), .dout(n650));
  jand g00587(.dina(n650), .dinb(n639), .dout(n651));
  jand g00588(.dina(n651), .dinb(n295), .dout(n652));
  jand g00589(.dina(n372), .dinb(n134), .dout(n653));
  jand g00590(.dina(n653), .dinb(n228), .dout(n654));
  jnot g00591(.din(n488), .dout(n655));
  jand g00592(.dina(n655), .dinb(n407), .dout(n656));
  jand g00593(.dina(n656), .dinb(n340), .dout(n657));
  jor  g00594(.dina(n269), .dinb(n213), .dout(n658));
  jand g00595(.dina(n658), .dinb(n450), .dout(n659));
  jand g00596(.dina(n236), .dinb(n315), .dout(n660));
  jand g00597(.dina(n236), .dinb(n132), .dout(n661));
  jor  g00598(.dina(n661), .dinb(n660), .dout(n662));
  jnot g00599(.din(n662), .dout(n663));
  jand g00600(.dina(n663), .dinb(n659), .dout(n664));
  jand g00601(.dina(n664), .dinb(n657), .dout(n665));
  jand g00602(.dina(n665), .dinb(n654), .dout(n666));
  jor  g00603(.dina(n188), .dinb(n164), .dout(n667));
  jand g00604(.dina(n667), .dinb(n385), .dout(n668));
  jand g00605(.dina(n668), .dinb(n154), .dout(n669));
  jand g00606(.dina(n172), .dinb(n116), .dout(n670));
  jnot g00607(.din(n670), .dout(n671));
  jand g00608(.dina(n671), .dinb(n359), .dout(n672));
  jand g00609(.dina(n672), .dinb(n157), .dout(n673));
  jand g00610(.dina(n195), .dinb(n101), .dout(n674));
  jnot g00611(.din(n674), .dout(n675));
  jand g00612(.dina(n675), .dinb(n245), .dout(n676));
  jand g00613(.dina(n389), .dinb(n315), .dout(n677));
  jnot g00614(.din(n677), .dout(n678));
  jand g00615(.dina(n678), .dinb(n309), .dout(n679));
  jand g00616(.dina(n679), .dinb(n676), .dout(n680));
  jand g00617(.dina(n680), .dinb(n673), .dout(n681));
  jand g00618(.dina(n681), .dinb(n669), .dout(n682));
  jand g00619(.dina(n682), .dinb(n666), .dout(n683));
  jand g00620(.dina(n683), .dinb(n652), .dout(n684));
  jand g00621(.dina(n684), .dinb(n631), .dout(n685));
  jand g00622(.dina(n235), .dinb(n278), .dout(n686));
  jnot g00623(.din(n686), .dout(n687));
  jand g00624(.dina(n687), .dinb(n257), .dout(n688));
  jnot g00625(.din(n453), .dout(n689));
  jand g00626(.dina(n689), .dinb(n146), .dout(n690));
  jand g00627(.dina(n690), .dinb(n688), .dout(n691));
  jor  g00628(.dina(n356), .dinb(n85), .dout(n692));
  jand g00629(.dina(n692), .dinb(n305), .dout(n693));
  jor  g00630(.dina(n207), .dinb(n81), .dout(n694));
  jand g00631(.dina(n236), .dinb(n116), .dout(n695));
  jnot g00632(.din(n695), .dout(n696));
  jand g00633(.dina(n696), .dinb(n694), .dout(n697));
  jand g00634(.dina(n697), .dinb(n693), .dout(n698));
  jand g00635(.dina(n698), .dinb(n691), .dout(n699));
  jor  g00636(.dina(n189), .dinb(n153), .dout(n700));
  jor  g00637(.dina(n141), .dinb(n91), .dout(n701));
  jand g00638(.dina(n222), .dinb(n97), .dout(n702));
  jnot g00639(.din(n702), .dout(n703));
  jand g00640(.dina(n703), .dinb(n701), .dout(n704));
  jand g00641(.dina(n704), .dinb(n700), .dout(n705));
  jand g00642(.dina(n235), .dinb(n147), .dout(n706));
  jnot g00643(.din(n706), .dout(n707));
  jor  g00644(.dina(n347), .dinb(n356), .dout(n708));
  jand g00645(.dina(n708), .dinb(n707), .dout(n709));
  jand g00646(.dina(n200), .dinb(n116), .dout(n710));
  jnot g00647(.din(n710), .dout(n711));
  jor  g00648(.dina(n188), .dinb(n176), .dout(n712));
  jand g00649(.dina(n712), .dinb(n711), .dout(n713));
  jand g00650(.dina(n713), .dinb(n709), .dout(n714));
  jor  g00651(.dina(n244), .dinb(n275), .dout(n715));
  jor  g00652(.dina(n207), .dinb(n244), .dout(n716));
  jand g00653(.dina(n716), .dinb(n715), .dout(n717));
  jand g00654(.dina(n159), .dinb(n200), .dout(n718));
  jnot g00655(.din(n718), .dout(n719));
  jand g00656(.dina(n192), .dinb(n106), .dout(n720));
  jnot g00657(.din(n720), .dout(n721));
  jand g00658(.dina(n721), .dinb(n719), .dout(n722));
  jand g00659(.dina(n722), .dinb(n717), .dout(n723));
  jand g00660(.dina(n723), .dinb(n714), .dout(n724));
  jand g00661(.dina(n724), .dinb(n705), .dout(n725));
  jand g00662(.dina(n725), .dinb(n699), .dout(n726));
  jand g00663(.dina(n726), .dinb(n685), .dout(n727));
  jand g00664(.dina(n727), .dinb(n591), .dout(n728));
  jxor g00665(.dina(n728), .dinb(n526), .dout(n729));
  jxor g00666(.dina(\a[30] ), .dinb(n88), .dout(n730));
  jnot g00667(.din(n730), .dout(n731));
  jand g00668(.dina(n731), .dinb(\a[31] ), .dout(n732));
  jand g00669(.dina(n286), .dinb(n82), .dout(n733));
  jand g00670(.dina(n733), .dinb(n268), .dout(n734));
  jand g00671(.dina(n192), .dinb(n344), .dout(n735));
  jnot g00672(.din(n735), .dout(n736));
  jand g00673(.dina(n736), .dinb(n646), .dout(n737));
  jand g00674(.dina(n236), .dinb(n219), .dout(n738));
  jnot g00675(.din(n738), .dout(n739));
  jand g00676(.dina(n739), .dinb(n494), .dout(n740));
  jand g00677(.dina(n372), .dinb(n165), .dout(n741));
  jand g00678(.dina(n741), .dinb(n740), .dout(n742));
  jand g00679(.dina(n742), .dinb(n737), .dout(n743));
  jand g00680(.dina(n743), .dinb(n734), .dout(n744));
  jand g00681(.dina(n375), .dinb(n134), .dout(n745));
  jand g00682(.dina(n578), .dinb(n536), .dout(n746));
  jand g00683(.dina(n746), .dinb(n745), .dout(n747));
  jand g00684(.dina(n272), .dinb(n172), .dout(n748));
  jnot g00685(.din(n748), .dout(n749));
  jand g00686(.dina(n389), .dinb(n300), .dout(n750));
  jnot g00687(.din(n750), .dout(n751));
  jand g00688(.dina(n751), .dinb(n749), .dout(n752));
  jand g00689(.dina(n396), .dinb(n221), .dout(n753));
  jand g00690(.dina(n753), .dinb(n752), .dout(n754));
  jand g00691(.dina(n754), .dinb(n747), .dout(n755));
  jor  g00692(.dina(n256), .dinb(n78), .dout(n756));
  jnot g00693(.din(n592), .dout(n757));
  jand g00694(.dina(n236), .dinb(n250), .dout(n758));
  jnot g00695(.din(n758), .dout(n759));
  jand g00696(.dina(n759), .dinb(n757), .dout(n760));
  jand g00697(.dina(n760), .dinb(n756), .dout(n761));
  jand g00698(.dina(n172), .dinb(n315), .dout(n762));
  jnot g00699(.din(n762), .dout(n763));
  jand g00700(.dina(n763), .dinb(n431), .dout(n764));
  jand g00701(.dina(n605), .dinb(n365), .dout(n765));
  jand g00702(.dina(n765), .dinb(n764), .dout(n766));
  jand g00703(.dina(n766), .dinb(n761), .dout(n767));
  jand g00704(.dina(n767), .dinb(n755), .dout(n768));
  jand g00705(.dina(n395), .dinb(n208), .dout(n769));
  jnot g00706(.din(n545), .dout(n770));
  jand g00707(.dina(n449), .dinb(n257), .dout(n771));
  jand g00708(.dina(n771), .dinb(n770), .dout(n772));
  jand g00709(.dina(n772), .dinb(n769), .dout(n773));
  jand g00710(.dina(n315), .dinb(n118), .dout(n774));
  jand g00711(.dina(n344), .dinb(n182), .dout(n775));
  jor  g00712(.dina(n775), .dinb(n774), .dout(n776));
  jnot g00713(.din(n776), .dout(n777));
  jnot g00714(.din(n661), .dout(n778));
  jand g00715(.dina(n778), .dinb(n478), .dout(n779));
  jand g00716(.dina(n779), .dinb(n445), .dout(n780));
  jand g00717(.dina(n780), .dinb(n777), .dout(n781));
  jand g00718(.dina(n781), .dinb(n773), .dout(n782));
  jand g00719(.dina(n782), .dinb(n768), .dout(n783));
  jand g00720(.dina(n783), .dinb(n744), .dout(n784));
  jand g00721(.dina(n159), .dinb(n118), .dout(n785));
  jnot g00722(.din(n785), .dout(n786));
  jand g00723(.dina(n786), .dinb(n635), .dout(n787));
  jand g00724(.dina(n542), .dinb(n417), .dout(n788));
  jand g00725(.dina(n788), .dinb(n450), .dout(n789));
  jand g00726(.dina(n789), .dinb(n787), .dout(n790));
  jand g00727(.dina(n562), .dinb(n405), .dout(n791));
  jand g00728(.dina(n389), .dinb(n155), .dout(n792));
  jnot g00729(.din(n792), .dout(n793));
  jand g00730(.dina(n793), .dinb(n346), .dout(n794));
  jnot g00731(.din(n113), .dout(n795));
  jand g00732(.dina(n389), .dinb(n132), .dout(n796));
  jor  g00733(.dina(n796), .dinb(n795), .dout(n797));
  jnot g00734(.din(n797), .dout(n798));
  jand g00735(.dina(n798), .dinb(n794), .dout(n799));
  jand g00736(.dina(n799), .dinb(n791), .dout(n800));
  jor  g00737(.dina(n347), .dinb(n275), .dout(n801));
  jand g00738(.dina(n801), .dinb(n532), .dout(n802));
  jand g00739(.dina(n583), .dinb(n383), .dout(n803));
  jand g00740(.dina(n803), .dinb(n802), .dout(n804));
  jor  g00741(.dina(n207), .dinb(n145), .dout(n805));
  jand g00742(.dina(n805), .dinb(n367), .dout(n806));
  jand g00743(.dina(n609), .dinb(n359), .dout(n807));
  jand g00744(.dina(n807), .dinb(n806), .dout(n808));
  jand g00745(.dina(n808), .dinb(n804), .dout(n809));
  jand g00746(.dina(n809), .dinb(n800), .dout(n810));
  jand g00747(.dina(n810), .dinb(n790), .dout(n811));
  jand g00748(.dina(n392), .dinb(n302), .dout(n812));
  jand g00749(.dina(n658), .dinb(n574), .dout(n813));
  jand g00750(.dina(n813), .dinb(n812), .dout(n814));
  jor  g00751(.dina(n164), .dinb(n213), .dout(n815));
  jand g00752(.dina(n815), .dinb(n146), .dout(n816));
  jor  g00753(.dina(n310), .dinb(n141), .dout(n817));
  jand g00754(.dina(n817), .dinb(n428), .dout(n818));
  jor  g00755(.dina(n347), .dinb(n259), .dout(n819));
  jand g00756(.dina(n819), .dinb(n249), .dout(n820));
  jand g00757(.dina(n820), .dinb(n818), .dout(n821));
  jand g00758(.dina(n821), .dinb(n816), .dout(n822));
  jand g00759(.dina(n822), .dinb(n814), .dout(n823));
  jor  g00760(.dina(n189), .dinb(n85), .dout(n824));
  jand g00761(.dina(n272), .dinb(n232), .dout(n825));
  jnot g00762(.din(n825), .dout(n826));
  jand g00763(.dina(n826), .dinb(n824), .dout(n827));
  jand g00764(.dina(n675), .dinb(n366), .dout(n828));
  jand g00765(.dina(n828), .dinb(n827), .dout(n829));
  jand g00766(.dina(n667), .dinb(n472), .dout(n830));
  jand g00767(.dina(n830), .dinb(n178), .dout(n831));
  jand g00768(.dina(n831), .dinb(n829), .dout(n832));
  jand g00769(.dina(n230), .dinb(n108), .dout(n833));
  jand g00770(.dina(n833), .dinb(n506), .dout(n834));
  jand g00771(.dina(n615), .dinb(n377), .dout(n835));
  jand g00772(.dina(n835), .dinb(n834), .dout(n836));
  jand g00773(.dina(n836), .dinb(n832), .dout(n837));
  jand g00774(.dina(n837), .dinb(n823), .dout(n838));
  jand g00775(.dina(n838), .dinb(n811), .dout(n839));
  jand g00776(.dina(n839), .dinb(n784), .dout(n840));
  jand g00777(.dina(n155), .dinb(n247), .dout(n841));
  jnot g00778(.din(n841), .dout(n842));
  jor  g00779(.dina(n244), .dinb(n91), .dout(n843));
  jand g00780(.dina(n843), .dinb(n284), .dout(n844));
  jand g00781(.dina(n844), .dinb(n842), .dout(n845));
  jand g00782(.dina(n215), .dinb(n106), .dout(n846));
  jnot g00783(.din(n846), .dout(n847));
  jand g00784(.dina(n847), .dinb(n382), .dout(n848));
  jand g00785(.dina(n633), .dinb(n245), .dout(n849));
  jand g00786(.dina(n849), .dinb(n848), .dout(n850));
  jand g00787(.dina(n850), .dinb(n845), .dout(n851));
  jand g00788(.dina(n125), .dinb(n247), .dout(n852));
  jnot g00789(.din(n852), .dout(n853));
  jand g00790(.dina(n853), .dinb(n716), .dout(n854));
  jand g00791(.dina(n854), .dinb(n280), .dout(n855));
  jand g00792(.dina(n232), .dinb(n215), .dout(n856));
  jnot g00793(.din(n856), .dout(n857));
  jand g00794(.dina(n857), .dinb(n515), .dout(n858));
  jand g00795(.dina(n315), .dinb(n106), .dout(n859));
  jnot g00796(.din(n859), .dout(n860));
  jand g00797(.dina(n860), .dinb(n290), .dout(n861));
  jand g00798(.dina(n861), .dinb(n858), .dout(n862));
  jand g00799(.dina(n862), .dinb(n855), .dout(n863));
  jand g00800(.dina(n863), .dinb(n851), .dout(n864));
  jor  g00801(.dina(n535), .dinb(n91), .dout(n865));
  jnot g00802(.din(n865), .dout(n866));
  jor  g00803(.dina(n866), .dinb(n323), .dout(n867));
  jnot g00804(.din(n867), .dout(n868));
  jand g00805(.dina(n551), .dinb(n337), .dout(n869));
  jand g00806(.dina(n543), .dinb(n527), .dout(n870));
  jand g00807(.dina(n870), .dinb(n869), .dout(n871));
  jand g00808(.dina(n871), .dinb(n868), .dout(n872));
  jand g00809(.dina(n278), .dinb(n125), .dout(n873));
  jnot g00810(.din(n873), .dout(n874));
  jand g00811(.dina(n159), .dinb(n247), .dout(n875));
  jnot g00812(.din(n875), .dout(n876));
  jand g00813(.dina(n876), .dinb(n874), .dout(n877));
  jand g00814(.dina(n719), .dinb(n228), .dout(n878));
  jand g00815(.dina(n878), .dinb(n877), .dout(n879));
  jand g00816(.dina(n184), .dinb(n136), .dout(n880));
  jand g00817(.dina(n250), .dinb(n344), .dout(n881));
  jnot g00818(.din(n881), .dout(n882));
  jand g00819(.dina(n882), .dinb(n304), .dout(n883));
  jand g00820(.dina(n883), .dinb(n880), .dout(n884));
  jand g00821(.dina(n884), .dinb(n879), .dout(n885));
  jand g00822(.dina(n885), .dinb(n872), .dout(n886));
  jand g00823(.dina(n886), .dinb(n864), .dout(n887));
  jor  g00824(.dina(n364), .dinb(n78), .dout(n888));
  jand g00825(.dina(n888), .dinb(n509), .dout(n889));
  jand g00826(.dina(n889), .dinb(n442), .dout(n890));
  jand g00827(.dina(n696), .dinb(n409), .dout(n891));
  jand g00828(.dina(n344), .dinb(n132), .dout(n892));
  jnot g00829(.din(n892), .dout(n893));
  jand g00830(.dina(n893), .dinb(n205), .dout(n894));
  jand g00831(.dina(n894), .dinb(n891), .dout(n895));
  jand g00832(.dina(n895), .dinb(n890), .dout(n896));
  jor  g00833(.dina(n535), .dinb(n78), .dout(n897));
  jnot g00834(.din(n897), .dout(n898));
  jor  g00835(.dina(n528), .dinb(n464), .dout(n899));
  jor  g00836(.dina(n899), .dinb(n898), .dout(n900));
  jnot g00837(.din(n900), .dout(n901));
  jand g00838(.dina(n470), .dinb(n270), .dout(n902));
  jand g00839(.dina(n902), .dinb(n92), .dout(n903));
  jand g00840(.dina(n903), .dinb(n901), .dout(n904));
  jand g00841(.dina(n904), .dinb(n896), .dout(n905));
  jand g00842(.dina(n192), .dinb(n128), .dout(n906));
  jnot g00843(.din(n906), .dout(n907));
  jand g00844(.dina(n315), .dinb(n128), .dout(n908));
  jnot g00845(.din(n908), .dout(n909));
  jand g00846(.dina(n909), .dinb(n907), .dout(n910));
  jand g00847(.dina(n910), .dinb(n354), .dout(n911));
  jand g00848(.dina(n315), .dinb(n200), .dout(n912));
  jnot g00849(.din(n912), .dout(n913));
  jand g00850(.dina(n913), .dinb(n607), .dout(n914));
  jand g00851(.dina(n643), .dinb(n343), .dout(n915));
  jand g00852(.dina(n915), .dinb(n277), .dout(n916));
  jand g00853(.dina(n916), .dinb(n914), .dout(n917));
  jand g00854(.dina(n917), .dinb(n911), .dout(n918));
  jand g00855(.dina(n918), .dinb(n905), .dout(n919));
  jand g00856(.dina(n919), .dinb(n887), .dout(n920));
  jand g00857(.dina(n920), .dinb(n840), .dout(n921));
  jnot g00858(.din(n921), .dout(n922));
  jand g00859(.dina(n909), .dinb(n302), .dout(n923));
  jor  g00860(.dina(n535), .dinb(n142), .dout(n924));
  jand g00861(.dina(n192), .dinb(n118), .dout(n925));
  jnot g00862(.din(n925), .dout(n926));
  jand g00863(.dina(n926), .dinb(n924), .dout(n927));
  jor  g00864(.dina(n856), .dinb(n604), .dout(n928));
  jnot g00865(.din(n928), .dout(n929));
  jand g00866(.dina(n929), .dinb(n927), .dout(n930));
  jand g00867(.dina(n930), .dinb(n923), .dout(n931));
  jand g00868(.dina(n579), .dinb(n268), .dout(n932));
  jand g00869(.dina(n633), .dinb(n82), .dout(n933));
  jand g00870(.dina(n708), .dinb(n494), .dout(n934));
  jand g00871(.dina(n934), .dinb(n933), .dout(n935));
  jand g00872(.dina(n935), .dinb(n932), .dout(n936));
  jand g00873(.dina(n936), .dinb(n931), .dout(n937));
  jand g00874(.dina(n711), .dinb(n255), .dout(n938));
  jand g00875(.dina(n434), .dinb(n202), .dout(n939));
  jand g00876(.dina(n939), .dinb(n190), .dout(n940));
  jand g00877(.dina(n940), .dinb(n938), .dout(n941));
  jor  g00878(.dina(n846), .dinb(n291), .dout(n942));
  jnot g00879(.din(n942), .dout(n943));
  jand g00880(.dina(n553), .dinb(n108), .dout(n944));
  jand g00881(.dina(n944), .dinb(n860), .dout(n945));
  jand g00882(.dina(n945), .dinb(n943), .dout(n946));
  jand g00883(.dina(n946), .dinb(n941), .dout(n947));
  jand g00884(.dina(n947), .dinb(n937), .dout(n948));
  jand g00885(.dina(n250), .dinb(n247), .dout(n949));
  jnot g00886(.din(n949), .dout(n950));
  jand g00887(.dina(n950), .dinb(n324), .dout(n951));
  jand g00888(.dina(n778), .dinb(n385), .dout(n952));
  jand g00889(.dina(n952), .dinb(n951), .dout(n953));
  jand g00890(.dina(n716), .dinb(n184), .dout(n954));
  jand g00891(.dina(n954), .dinb(n506), .dout(n955));
  jand g00892(.dina(n955), .dinb(n953), .dout(n956));
  jand g00893(.dina(n354), .dinb(n103), .dout(n957));
  jand g00894(.dina(n957), .dinb(n566), .dout(n958));
  jor  g00895(.dina(n152), .dinb(n145), .dout(n959));
  jand g00896(.dina(n959), .dinb(n586), .dout(n960));
  jand g00897(.dina(n960), .dinb(n198), .dout(n961));
  jand g00898(.dina(n961), .dinb(n958), .dout(n962));
  jand g00899(.dina(n736), .dinb(n536), .dout(n963));
  jand g00900(.dina(n97), .dinb(n203), .dout(n964));
  jnot g00901(.din(n964), .dout(n965));
  jand g00902(.dina(n236), .dinb(n215), .dout(n966));
  jnot g00903(.din(n966), .dout(n967));
  jand g00904(.dina(n967), .dinb(n965), .dout(n968));
  jand g00905(.dina(n968), .dinb(n963), .dout(n969));
  jand g00906(.dina(n418), .dinb(n290), .dout(n970));
  jand g00907(.dina(n614), .dinb(n304), .dout(n971));
  jand g00908(.dina(n971), .dinb(n970), .dout(n972));
  jand g00909(.dina(n972), .dinb(n969), .dout(n973));
  jand g00910(.dina(n973), .dinb(n962), .dout(n974));
  jand g00911(.dina(n974), .dinb(n956), .dout(n975));
  jand g00912(.dina(n461), .dinb(n243), .dout(n976));
  jand g00913(.dina(n976), .dinb(n149), .dout(n977));
  jand g00914(.dina(n749), .dinb(n703), .dout(n978));
  jor  g00915(.dina(n259), .dinb(n285), .dout(n979));
  jand g00916(.dina(n979), .dinb(n325), .dout(n980));
  jand g00917(.dina(n980), .dinb(n978), .dout(n981));
  jand g00918(.dina(n739), .dinb(n441), .dout(n982));
  jand g00919(.dina(n815), .dinb(n667), .dout(n983));
  jand g00920(.dina(n983), .dinb(n982), .dout(n984));
  jand g00921(.dina(n984), .dinb(n981), .dout(n985));
  jand g00922(.dina(n985), .dinb(n977), .dout(n986));
  jand g00923(.dina(n338), .dinb(n215), .dout(n987));
  jnot g00924(.din(n987), .dout(n988));
  jand g00925(.dina(n988), .dinb(n511), .dout(n989));
  jand g00926(.dina(n786), .dinb(n607), .dout(n990));
  jand g00927(.dina(n990), .dinb(n989), .dout(n991));
  jand g00928(.dina(n338), .dinb(n250), .dout(n992));
  jnot g00929(.din(n992), .dout(n993));
  jand g00930(.dina(n993), .dinb(n500), .dout(n994));
  jand g00931(.dina(n824), .dinb(n174), .dout(n995));
  jand g00932(.dina(n995), .dinb(n994), .dout(n996));
  jor  g00933(.dina(n256), .dinb(n112), .dout(n997));
  jand g00934(.dina(n583), .dinb(n228), .dout(n998));
  jand g00935(.dina(n998), .dinb(n997), .dout(n999));
  jand g00936(.dina(n999), .dinb(n996), .dout(n1000));
  jand g00937(.dina(n1000), .dinb(n991), .dout(n1001));
  jand g00938(.dina(n1001), .dinb(n986), .dout(n1002));
  jand g00939(.dina(n1002), .dinb(n975), .dout(n1003));
  jand g00940(.dina(n1003), .dinb(n948), .dout(n1004));
  jand g00941(.dina(n449), .dinb(n270), .dout(n1005));
  jand g00942(.dina(n1005), .dinb(n136), .dout(n1006));
  jand g00943(.dina(n701), .dinb(n499), .dout(n1007));
  jand g00944(.dina(n1007), .dinb(n527), .dout(n1008));
  jand g00945(.dina(n712), .dinb(n439), .dout(n1009));
  jand g00946(.dina(n1009), .dinb(n697), .dout(n1010));
  jand g00947(.dina(n1010), .dinb(n1008), .dout(n1011));
  jand g00948(.dina(n1011), .dinb(n1006), .dout(n1012));
  jand g00949(.dina(n315), .dinb(n247), .dout(n1013));
  jnot g00950(.din(n1013), .dout(n1014));
  jand g00951(.dina(n1014), .dinb(n757), .dout(n1015));
  jand g00952(.dina(n793), .dinb(n715), .dout(n1016));
  jand g00953(.dina(n1016), .dinb(n134), .dout(n1017));
  jand g00954(.dina(n1017), .dinb(n1015), .dout(n1018));
  jand g00955(.dina(n842), .dinb(n472), .dout(n1019));
  jand g00956(.dina(n907), .dinb(n221), .dout(n1020));
  jand g00957(.dina(n1020), .dinb(n635), .dout(n1021));
  jand g00958(.dina(n1021), .dinb(n1019), .dout(n1022));
  jand g00959(.dina(n655), .dinb(n317), .dout(n1023));
  jand g00960(.dina(n476), .dinb(n414), .dout(n1024));
  jand g00961(.dina(n383), .dinb(n343), .dout(n1025));
  jand g00962(.dina(n1025), .dinb(n1024), .dout(n1026));
  jand g00963(.dina(n1026), .dinb(n1023), .dout(n1027));
  jand g00964(.dina(n1027), .dinb(n1022), .dout(n1028));
  jand g00965(.dina(n1028), .dinb(n1018), .dout(n1029));
  jand g00966(.dina(n1029), .dinb(n1012), .dout(n1030));
  jnot g00967(.din(n452), .dout(n1031));
  jand g00968(.dina(n1031), .dinb(n288), .dout(n1032));
  jand g00969(.dina(n250), .dinb(n128), .dout(n1033));
  jnot g00970(.din(n1033), .dout(n1034));
  jand g00971(.dina(n1034), .dinb(n551), .dout(n1035));
  jand g00972(.dina(n407), .dinb(n311), .dout(n1036));
  jand g00973(.dina(n1036), .dinb(n1035), .dout(n1037));
  jand g00974(.dina(n1037), .dinb(n1032), .dout(n1038));
  jor  g00975(.dina(n256), .dinb(n152), .dout(n1039));
  jor  g00976(.dina(n259), .dinb(n141), .dout(n1040));
  jand g00977(.dina(n1040), .dinb(n557), .dout(n1041));
  jand g00978(.dina(n1041), .dinb(n1039), .dout(n1042));
  jand g00979(.dina(n532), .dinb(n423), .dout(n1043));
  jand g00980(.dina(n1043), .dinb(n417), .dout(n1044));
  jand g00981(.dina(n1044), .dinb(n1042), .dout(n1045));
  jand g00982(.dina(n1045), .dinb(n1038), .dout(n1046));
  jor  g00983(.dina(n152), .dinb(n85), .dout(n1047));
  jand g00984(.dina(n1047), .dinb(n609), .dout(n1048));
  jand g00985(.dina(n1048), .dinb(n693), .dout(n1049));
  jand g00986(.dina(n647), .dinb(n329), .dout(n1050));
  jand g00987(.dina(n893), .dinb(n337), .dout(n1051));
  jand g00988(.dina(n1051), .dinb(n224), .dout(n1052));
  jand g00989(.dina(n1052), .dinb(n1050), .dout(n1053));
  jand g00990(.dina(n1053), .dinb(n1049), .dout(n1054));
  jand g00991(.dina(n182), .dinb(n247), .dout(n1055));
  jor  g00992(.dina(n482), .dinb(n1055), .dout(n1056));
  jnot g00993(.din(n1056), .dout(n1057));
  jand g00994(.dina(n409), .dinb(n214), .dout(n1058));
  jand g00995(.dina(n340), .dinb(n157), .dout(n1059));
  jand g00996(.dina(n1059), .dinb(n1058), .dout(n1060));
  jand g00997(.dina(n1060), .dinb(n1057), .dout(n1061));
  jand g00998(.dina(n853), .dinb(n533), .dout(n1062));
  jand g00999(.dina(n395), .dinb(n252), .dout(n1063));
  jand g01000(.dina(n1063), .dinb(n1062), .dout(n1064));
  jand g01001(.dina(n222), .dinb(n159), .dout(n1065));
  jnot g01002(.din(n1065), .dout(n1066));
  jand g01003(.dina(n1066), .dinb(n445), .dout(n1067));
  jand g01004(.dina(n346), .dinb(n286), .dout(n1068));
  jand g01005(.dina(n1068), .dinb(n1067), .dout(n1069));
  jand g01006(.dina(n1069), .dinb(n1064), .dout(n1070));
  jand g01007(.dina(n1070), .dinb(n1061), .dout(n1071));
  jand g01008(.dina(n1071), .dinb(n1054), .dout(n1072));
  jand g01009(.dina(n1072), .dinb(n1046), .dout(n1073));
  jand g01010(.dina(n1073), .dinb(n1030), .dout(n1074));
  jand g01011(.dina(n1074), .dinb(n1004), .dout(n1075));
  jnot g01012(.din(n1075), .dout(n1076));
  jand g01013(.dina(n1076), .dinb(n922), .dout(n1077));
  jand g01014(.dina(n707), .dinb(n352), .dout(n1078));
  jand g01015(.dina(n692), .dinb(n543), .dout(n1079));
  jand g01016(.dina(n1079), .dinb(n1078), .dout(n1080));
  jand g01017(.dina(n826), .dinb(n396), .dout(n1081));
  jand g01018(.dina(n759), .dinb(n180), .dout(n1082));
  jand g01019(.dina(n1082), .dinb(n1081), .dout(n1083));
  jand g01020(.dina(n1083), .dinb(n1080), .dout(n1084));
  jand g01021(.dina(n423), .dinb(n280), .dout(n1085));
  jand g01022(.dina(n414), .dinb(n391), .dout(n1086));
  jand g01023(.dina(n1086), .dinb(n1085), .dout(n1087));
  jand g01024(.dina(n385), .dinb(n130), .dout(n1088));
  jand g01025(.dina(n1088), .dinb(n752), .dout(n1089));
  jand g01026(.dina(n719), .dinb(n224), .dout(n1090));
  jand g01027(.dina(n1090), .dinb(n1019), .dout(n1091));
  jand g01028(.dina(n1091), .dinb(n1089), .dout(n1092));
  jand g01029(.dina(n1092), .dinb(n1087), .dout(n1093));
  jand g01030(.dina(n1093), .dinb(n1084), .dout(n1094));
  jand g01031(.dina(n847), .dinb(n609), .dout(n1095));
  jand g01032(.dina(n1095), .dinb(n190), .dout(n1096));
  jand g01033(.dina(n712), .dinb(n500), .dout(n1097));
  jand g01034(.dina(n1097), .dinb(n277), .dout(n1098));
  jand g01035(.dina(n481), .dinb(n428), .dout(n1099));
  jand g01036(.dina(n383), .dinb(n120), .dout(n1100));
  jand g01037(.dina(n1100), .dinb(n1099), .dout(n1101));
  jand g01038(.dina(n1101), .dinb(n1098), .dout(n1102));
  jand g01039(.dina(n1102), .dinb(n1096), .dout(n1103));
  jand g01040(.dina(n357), .dinb(n284), .dout(n1104));
  jand g01041(.dina(n763), .dinb(n509), .dout(n1105));
  jand g01042(.dina(n1105), .dinb(n1104), .dout(n1106));
  jand g01043(.dina(n1106), .dinb(n109), .dout(n1107));
  jand g01044(.dina(n462), .dinb(n434), .dout(n1108));
  jand g01045(.dina(n1108), .dinb(n924), .dout(n1109));
  jand g01046(.dina(n824), .dinb(n154), .dout(n1110));
  jand g01047(.dina(n819), .dinb(n336), .dout(n1111));
  jand g01048(.dina(n1111), .dinb(n1110), .dout(n1112));
  jand g01049(.dina(n1112), .dinb(n1109), .dout(n1113));
  jand g01050(.dina(n1113), .dinb(n1107), .dout(n1114));
  jand g01051(.dina(n1114), .dinb(n1103), .dout(n1115));
  jand g01052(.dina(n1115), .dinb(n1094), .dout(n1116));
  jand g01053(.dina(n876), .dinb(n197), .dout(n1117));
  jand g01054(.dina(n1117), .dinb(n302), .dout(n1118));
  jand g01055(.dina(n696), .dinb(n354), .dout(n1119));
  jand g01056(.dina(n1119), .dinb(n1035), .dout(n1120));
  jand g01057(.dina(n1120), .dinb(n1118), .dout(n1121));
  jand g01058(.dina(n606), .dinb(n468), .dout(n1122));
  jand g01059(.dina(n993), .dinb(n529), .dout(n1123));
  jand g01060(.dina(n1123), .dinb(n443), .dout(n1124));
  jand g01061(.dina(n1124), .dinb(n1122), .dout(n1125));
  jand g01062(.dina(n1125), .dinb(n1121), .dout(n1126));
  jand g01063(.dina(n1126), .dinb(n1116), .dout(n1127));
  jand g01064(.dina(n1040), .dinb(n967), .dout(n1128));
  jand g01065(.dina(n721), .dinb(n655), .dout(n1129));
  jand g01066(.dina(n371), .dinb(n234), .dout(n1130));
  jand g01067(.dina(n1130), .dinb(n1129), .dout(n1131));
  jand g01068(.dina(n1131), .dinb(n1128), .dout(n1132));
  jor  g01069(.dina(n640), .dinb(n148), .dout(n1133));
  jnot g01070(.din(n1133), .dout(n1134));
  jand g01071(.dina(n853), .dinb(n461), .dout(n1135));
  jand g01072(.dina(n1135), .dinb(n1134), .dout(n1136));
  jand g01073(.dina(n703), .dinb(n143), .dout(n1137));
  jand g01074(.dina(n1137), .dinb(n717), .dout(n1138));
  jand g01075(.dina(n1138), .dinb(n1136), .dout(n1139));
  jand g01076(.dina(n532), .dinb(n441), .dout(n1140));
  jand g01077(.dina(n1140), .dinb(n626), .dout(n1141));
  jand g01078(.dina(n874), .dinb(n288), .dout(n1142));
  jand g01079(.dina(n182), .dinb(n203), .dout(n1143));
  jnot g01080(.din(n1143), .dout(n1144));
  jand g01081(.dina(n1144), .dinb(n337), .dout(n1145));
  jand g01082(.dina(n1145), .dinb(n1142), .dout(n1146));
  jand g01083(.dina(n1146), .dinb(n1141), .dout(n1147));
  jand g01084(.dina(n1147), .dinb(n1139), .dout(n1148));
  jand g01085(.dina(n1148), .dinb(n1132), .dout(n1149));
  jand g01086(.dina(n619), .dinb(n366), .dout(n1150));
  jand g01087(.dina(n1150), .dinb(n1014), .dout(n1151));
  jand g01088(.dina(n278), .dinb(n300), .dout(n1152));
  jnot g01089(.din(n1152), .dout(n1153));
  jand g01090(.dina(n1153), .dinb(n595), .dout(n1154));
  jand g01091(.dina(n418), .dinb(n311), .dout(n1155));
  jand g01092(.dina(n527), .dinb(n202), .dout(n1156));
  jand g01093(.dina(n1156), .dinb(n1155), .dout(n1157));
  jand g01094(.dina(n1157), .dinb(n1154), .dout(n1158));
  jand g01095(.dina(n1158), .dinb(n1151), .dout(n1159));
  jand g01096(.dina(n478), .dinb(n325), .dout(n1160));
  jand g01097(.dina(n711), .dinb(n270), .dout(n1161));
  jand g01098(.dina(n1161), .dinb(n1160), .dout(n1162));
  jand g01099(.dina(n786), .dinb(n445), .dout(n1163));
  jand g01100(.dina(n1163), .dinb(n494), .dout(n1164));
  jand g01101(.dina(n965), .dinb(n793), .dout(n1165));
  jand g01102(.dina(n116), .dinb(n247), .dout(n1166));
  jnot g01103(.din(n1166), .dout(n1167));
  jand g01104(.dina(n1167), .dinb(n805), .dout(n1168));
  jand g01105(.dina(n1168), .dinb(n1165), .dout(n1169));
  jand g01106(.dina(n1169), .dinb(n1164), .dout(n1170));
  jand g01107(.dina(n1170), .dinb(n1162), .dout(n1171));
  jand g01108(.dina(n1171), .dinb(n1159), .dout(n1172));
  jand g01109(.dina(n1172), .dinb(n1149), .dout(n1173));
  jand g01110(.dina(n893), .dinb(n359), .dout(n1174));
  jand g01111(.dina(n1174), .dinb(n857), .dout(n1175));
  jand g01112(.dina(n633), .dinb(n221), .dout(n1176));
  jand g01113(.dina(n235), .dinb(n247), .dout(n1177));
  jnot g01114(.din(n1177), .dout(n1178));
  jand g01115(.dina(n1178), .dinb(n165), .dout(n1179));
  jand g01116(.dina(n1179), .dinb(n1176), .dout(n1180));
  jand g01117(.dina(n1180), .dinb(n1175), .dout(n1181));
  jand g01118(.dina(n346), .dinb(n324), .dout(n1182));
  jand g01119(.dina(n1182), .dinb(n405), .dout(n1183));
  jor  g01120(.dina(n256), .dinb(n370), .dout(n1184));
  jand g01121(.dina(n1184), .dinb(n208), .dout(n1185));
  jand g01122(.dina(n1047), .dinb(n217), .dout(n1186));
  jand g01123(.dina(n1186), .dinb(n1185), .dout(n1187));
  jand g01124(.dina(n1187), .dinb(n1183), .dout(n1188));
  jand g01125(.dina(n1188), .dinb(n1181), .dout(n1189));
  jand g01126(.dina(n694), .dinb(n82), .dout(n1190));
  jand g01127(.dina(n1190), .dinb(n817), .dout(n1191));
  jand g01128(.dina(n675), .dinb(n449), .dout(n1192));
  jand g01129(.dina(n574), .dinb(n470), .dout(n1193));
  jand g01130(.dina(n1193), .dinb(n1192), .dout(n1194));
  jand g01131(.dina(n1194), .dinb(n1191), .dout(n1195));
  jand g01132(.dina(n678), .dinb(n262), .dout(n1196));
  jand g01133(.dina(n413), .dinb(n136), .dout(n1197));
  jand g01134(.dina(n1197), .dinb(n1196), .dout(n1198));
  jand g01135(.dina(n687), .dinb(n757), .dout(n1199));
  jand g01136(.dina(n1199), .dinb(n178), .dout(n1200));
  jand g01137(.dina(n1200), .dinb(n1198), .dout(n1201));
  jand g01138(.dina(n701), .dinb(n255), .dout(n1202));
  jand g01139(.dina(n1202), .dinb(n483), .dout(n1203));
  jand g01140(.dina(n860), .dinb(n409), .dout(n1204));
  jand g01141(.dina(n322), .dinb(n260), .dout(n1205));
  jand g01142(.dina(n1205), .dinb(n1204), .dout(n1206));
  jand g01143(.dina(n1206), .dinb(n1203), .dout(n1207));
  jand g01144(.dina(n1207), .dinb(n1201), .dout(n1208));
  jand g01145(.dina(n1208), .dinb(n1195), .dout(n1209));
  jand g01146(.dina(n1209), .dinb(n1189), .dout(n1210));
  jand g01147(.dina(n1210), .dinb(n1173), .dout(n1211));
  jand g01148(.dina(n1211), .dinb(n1127), .dout(n1212));
  jnot g01149(.din(n1212), .dout(n1213));
  jand g01150(.dina(n1213), .dinb(n1076), .dout(n1214));
  jor  g01151(.dina(n852), .dinb(n545), .dout(n1215));
  jnot g01152(.din(n1215), .dout(n1216));
  jand g01153(.dina(n997), .dinb(n658), .dout(n1217));
  jand g01154(.dina(n913), .dinb(n605), .dout(n1218));
  jand g01155(.dina(n1218), .dinb(n1217), .dout(n1219));
  jand g01156(.dina(n1219), .dinb(n1216), .dout(n1220));
  jor  g01157(.dina(n535), .dinb(n112), .dout(n1221));
  jand g01158(.dina(n1221), .dinb(n609), .dout(n1222));
  jand g01159(.dina(n1144), .dinb(n909), .dout(n1223));
  jand g01160(.dina(n1223), .dinb(n1222), .dout(n1224));
  jand g01161(.dina(n622), .dinb(n230), .dout(n1225));
  jand g01162(.dina(n993), .dinb(n542), .dout(n1226));
  jand g01163(.dina(n1226), .dinb(n1225), .dout(n1227));
  jand g01164(.dina(n1227), .dinb(n1224), .dout(n1228));
  jand g01165(.dina(n1228), .dinb(n1220), .dout(n1229));
  jand g01166(.dina(n219), .dinb(n106), .dout(n1230));
  jnot g01167(.din(n1230), .dout(n1231));
  jand g01168(.dina(n1231), .dinb(n553), .dout(n1232));
  jand g01169(.dina(n1232), .dinb(n409), .dout(n1233));
  jand g01170(.dina(n598), .dinb(n500), .dout(n1234));
  jand g01171(.dina(n739), .dinb(n432), .dout(n1235));
  jand g01172(.dina(n1235), .dinb(n1234), .dout(n1236));
  jand g01173(.dina(n428), .dinb(n238), .dout(n1237));
  jand g01174(.dina(n516), .dinb(n461), .dout(n1238));
  jand g01175(.dina(n1238), .dinb(n1237), .dout(n1239));
  jand g01176(.dina(n1239), .dinb(n1236), .dout(n1240));
  jand g01177(.dina(n1240), .dinb(n1233), .dout(n1241));
  jand g01178(.dina(n352), .dinb(n252), .dout(n1242));
  jand g01179(.dina(n907), .dinb(n826), .dout(n1243));
  jand g01180(.dina(n1243), .dinb(n716), .dout(n1244));
  jand g01181(.dina(n1244), .dinb(n1242), .dout(n1245));
  jand g01182(.dina(n882), .dinb(n136), .dout(n1246));
  jand g01183(.dina(n763), .dinb(n443), .dout(n1247));
  jand g01184(.dina(n1247), .dinb(n1246), .dout(n1248));
  jand g01185(.dina(n536), .dinb(n413), .dout(n1249));
  jand g01186(.dina(n486), .dinb(n357), .dout(n1250));
  jand g01187(.dina(n1250), .dinb(n1249), .dout(n1251));
  jand g01188(.dina(n1251), .dinb(n1248), .dout(n1252));
  jand g01189(.dina(n1252), .dinb(n1245), .dout(n1253));
  jand g01190(.dina(n1253), .dinb(n1241), .dout(n1254));
  jand g01191(.dina(n1254), .dinb(n1229), .dout(n1255));
  jand g01192(.dina(n979), .dinb(n274), .dout(n1256));
  jand g01193(.dina(n824), .dinb(n707), .dout(n1257));
  jand g01194(.dina(n1257), .dinb(n1256), .dout(n1258));
  jand g01195(.dina(n1184), .dinb(n532), .dout(n1259));
  jand g01196(.dina(n290), .dinb(n234), .dout(n1260));
  jand g01197(.dina(n1260), .dinb(n1259), .dout(n1261));
  jand g01198(.dina(n1261), .dinb(n1258), .dout(n1262));
  jand g01199(.dina(n389), .dinb(n182), .dout(n1263));
  jnot g01200(.din(n1263), .dout(n1264));
  jand g01201(.dina(n1264), .dinb(n511), .dout(n1265));
  jand g01202(.dina(n793), .dinb(n331), .dout(n1266));
  jand g01203(.dina(n1266), .dinb(n1265), .dout(n1267));
  jor  g01204(.dina(n206), .dinb(n416), .dout(n1268));
  jand g01205(.dina(n1268), .dinb(n515), .dout(n1269));
  jand g01206(.dina(n1269), .dinb(n959), .dout(n1270));
  jand g01207(.dina(n1270), .dinb(n1267), .dout(n1271));
  jand g01208(.dina(n1271), .dinb(n1262), .dout(n1272));
  jand g01209(.dina(n888), .dinb(n143), .dout(n1273));
  jand g01210(.dina(n865), .dinb(n696), .dout(n1274));
  jand g01211(.dina(n633), .dinb(n595), .dout(n1275));
  jand g01212(.dina(n1275), .dinb(n1274), .dout(n1276));
  jand g01213(.dina(n1276), .dinb(n1273), .dout(n1277));
  jand g01214(.dina(n667), .dinb(n336), .dout(n1278));
  jor  g01215(.dina(n966), .dinb(n220), .dout(n1279));
  jnot g01216(.din(n1279), .dout(n1280));
  jand g01217(.dina(n678), .dinb(n396), .dout(n1281));
  jand g01218(.dina(n1281), .dinb(n1280), .dout(n1282));
  jand g01219(.dina(n1282), .dinb(n1278), .dout(n1283));
  jand g01220(.dina(n924), .dinb(n439), .dout(n1284));
  jand g01221(.dina(n687), .dinb(n309), .dout(n1285));
  jand g01222(.dina(n1285), .dinb(n1284), .dout(n1286));
  jand g01223(.dina(n641), .dinb(n386), .dout(n1287));
  jand g01224(.dina(n1287), .dinb(n1085), .dout(n1288));
  jand g01225(.dina(n1288), .dinb(n1286), .dout(n1289));
  jand g01226(.dina(n1289), .dinb(n1283), .dout(n1290));
  jand g01227(.dina(n1290), .dinb(n1277), .dout(n1291));
  jand g01228(.dina(n1291), .dinb(n1272), .dout(n1292));
  jand g01229(.dina(n354), .dinb(n243), .dout(n1293));
  jand g01230(.dina(n1293), .dinb(n494), .dout(n1294));
  jand g01231(.dina(n1167), .dinb(n689), .dout(n1295));
  jand g01232(.dina(n701), .dinb(n375), .dout(n1296));
  jand g01233(.dina(n1296), .dinb(n1295), .dout(n1297));
  jand g01234(.dina(n1297), .dinb(n1294), .dout(n1298));
  jand g01235(.dina(n700), .dinb(n533), .dout(n1299));
  jand g01236(.dina(n751), .dinb(n612), .dout(n1300));
  jand g01237(.dina(n1300), .dinb(n1299), .dout(n1301));
  jand g01238(.dina(n1301), .dinb(n563), .dout(n1302));
  jand g01239(.dina(n646), .dinb(n255), .dout(n1303));
  jand g01240(.dina(n1303), .dinb(n1100), .dout(n1304));
  jand g01241(.dina(n329), .dinb(n165), .dout(n1305));
  jand g01242(.dina(n462), .dinb(n314), .dout(n1306));
  jand g01243(.dina(n1306), .dinb(n1305), .dout(n1307));
  jand g01244(.dina(n1307), .dinb(n1304), .dout(n1308));
  jand g01245(.dina(n1308), .dinb(n1302), .dout(n1309));
  jand g01246(.dina(n1309), .dinb(n1298), .dout(n1310));
  jand g01247(.dina(n101), .dinb(n132), .dout(n1311));
  jor  g01248(.dina(n1311), .dinb(n267), .dout(n1312));
  jand g01249(.dina(n235), .dinb(n172), .dout(n1313));
  jnot g01250(.din(n1313), .dout(n1314));
  jand g01251(.dina(n1314), .dinb(n130), .dout(n1315));
  jnot g01252(.din(n1315), .dout(n1316));
  jor  g01253(.dina(n1316), .dinb(n1312), .dout(n1317));
  jnot g01254(.din(n1317), .dout(n1318));
  jand g01255(.dina(n805), .dinb(n551), .dout(n1319));
  jand g01256(.dina(n470), .dinb(n245), .dout(n1320));
  jand g01257(.dina(n1320), .dinb(n1319), .dout(n1321));
  jand g01258(.dina(n1178), .dinb(n756), .dout(n1322));
  jand g01259(.dina(n583), .dinb(n517), .dout(n1323));
  jand g01260(.dina(n1323), .dinb(n1322), .dout(n1324));
  jand g01261(.dina(n1324), .dinb(n1321), .dout(n1325));
  jand g01262(.dina(n1325), .dinb(n1318), .dout(n1326));
  jand g01263(.dina(n377), .dinb(n184), .dout(n1327));
  jand g01264(.dina(n1327), .dinb(n108), .dout(n1328));
  jand g01265(.dina(n435), .dinb(n385), .dout(n1329));
  jand g01266(.dina(n1329), .dinb(n218), .dout(n1330));
  jand g01267(.dina(n1330), .dinb(n1328), .dout(n1331));
  jand g01268(.dina(n857), .dinb(n843), .dout(n1332));
  jand g01269(.dina(n1332), .dinb(n1024), .dout(n1333));
  jand g01270(.dina(n1040), .dinb(n359), .dout(n1334));
  jand g01271(.dina(n566), .dinb(n505), .dout(n1335));
  jand g01272(.dina(n1335), .dinb(n1334), .dout(n1336));
  jand g01273(.dina(n1336), .dinb(n1333), .dout(n1337));
  jand g01274(.dina(n1337), .dinb(n1331), .dout(n1338));
  jand g01275(.dina(n1338), .dinb(n1326), .dout(n1339));
  jand g01276(.dina(n1339), .dinb(n1310), .dout(n1340));
  jand g01277(.dina(n1340), .dinb(n1292), .dout(n1341));
  jand g01278(.dina(n1341), .dinb(n1255), .dout(n1342));
  jnot g01279(.din(n1342), .dout(n1343));
  jand g01280(.dina(n1343), .dinb(n1213), .dout(n1344));
  jand g01281(.dina(n907), .dinb(n708), .dout(n1345));
  jor  g01282(.dina(n269), .dinb(n244), .dout(n1346));
  jand g01283(.dina(n1346), .dinb(n359), .dout(n1347));
  jand g01284(.dina(n1347), .dinb(n1345), .dout(n1348));
  jand g01285(.dina(n322), .dinb(n161), .dout(n1349));
  jand g01286(.dina(n536), .dinb(n377), .dout(n1350));
  jand g01287(.dina(n1350), .dinb(n1349), .dout(n1351));
  jand g01288(.dina(n1351), .dinb(n1348), .dout(n1352));
  jand g01289(.dina(n843), .dinb(n177), .dout(n1353));
  jand g01290(.dina(n1353), .dinb(n501), .dout(n1354));
  jand g01291(.dina(n1354), .dinb(n109), .dout(n1355));
  jand g01292(.dina(n1184), .dinb(n113), .dout(n1356));
  jand g01293(.dina(n272), .dinb(n106), .dout(n1357));
  jor  g01294(.dina(n1357), .dinb(n133), .dout(n1358));
  jnot g01295(.din(n1358), .dout(n1359));
  jand g01296(.dina(n1359), .dinb(n1356), .dout(n1360));
  jand g01297(.dina(n1360), .dinb(n451), .dout(n1361));
  jand g01298(.dina(n1361), .dinb(n1355), .dout(n1362));
  jand g01299(.dina(n1362), .dinb(n1352), .dout(n1363));
  jand g01300(.dina(n805), .dinb(n757), .dout(n1364));
  jnot g01301(.din(n1364), .dout(n1365));
  jor  g01302(.dina(n796), .dinb(n625), .dout(n1366));
  jand g01303(.dina(n116), .dinb(n101), .dout(n1367));
  jor  g01304(.dina(n1143), .dinb(n1367), .dout(n1368));
  jor  g01305(.dina(n1368), .dinb(n1366), .dout(n1369));
  jor  g01306(.dina(n1369), .dinb(n1365), .dout(n1370));
  jnot g01307(.din(n924), .dout(n1371));
  jor  g01308(.dina(n1371), .dinb(n204), .dout(n1372));
  jor  g01309(.dina(n1372), .dinb(n928), .dout(n1373));
  jand g01310(.dina(n338), .dinb(n300), .dout(n1374));
  jnot g01311(.din(n701), .dout(n1375));
  jor  g01312(.dina(n1375), .dinb(n1374), .dout(n1376));
  jand g01313(.dina(n338), .dinb(n195), .dout(n1377));
  jor  g01314(.dina(n1377), .dinb(n183), .dout(n1378));
  jor  g01315(.dina(n1378), .dinb(n1376), .dout(n1379));
  jor  g01316(.dina(n1379), .dinb(n1373), .dout(n1380));
  jor  g01317(.dina(n1380), .dinb(n1370), .dout(n1381));
  jnot g01318(.din(n1381), .dout(n1382));
  jand g01319(.dina(n763), .dinb(n517), .dout(n1383));
  jand g01320(.dina(n1383), .dinb(n355), .dout(n1384));
  jand g01321(.dina(n756), .dinb(n255), .dout(n1385));
  jand g01322(.dina(n1385), .dinb(n506), .dout(n1386));
  jand g01323(.dina(n1386), .dinb(n1384), .dout(n1387));
  jand g01324(.dina(n897), .dinb(n427), .dout(n1388));
  jand g01325(.dina(n1388), .dinb(n826), .dout(n1389));
  jand g01326(.dina(n366), .dinb(n325), .dout(n1390));
  jand g01327(.dina(n1390), .dinb(n304), .dout(n1391));
  jand g01328(.dina(n1391), .dinb(n1389), .dout(n1392));
  jand g01329(.dina(n1392), .dinb(n1387), .dout(n1393));
  jand g01330(.dina(n1393), .dinb(n1382), .dout(n1394));
  jand g01331(.dina(n1394), .dinb(n1363), .dout(n1395));
  jand g01332(.dina(n315), .dinb(n147), .dout(n1396));
  jor  g01333(.dina(n1396), .dinb(n510), .dout(n1397));
  jnot g01334(.din(n1397), .dout(n1398));
  jand g01335(.dina(n1398), .dinb(n655), .dout(n1399));
  jand g01336(.dina(n260), .dinb(n217), .dout(n1400));
  jand g01337(.dina(n1400), .dinb(n391), .dout(n1401));
  jand g01338(.dina(n801), .dinb(n700), .dout(n1402));
  jand g01339(.dina(n232), .dinb(n250), .dout(n1403));
  jor  g01340(.dina(n966), .dinb(n1403), .dout(n1404));
  jnot g01341(.din(n1404), .dout(n1405));
  jand g01342(.dina(n1405), .dinb(n1402), .dout(n1406));
  jand g01343(.dina(n1406), .dinb(n1401), .dout(n1407));
  jand g01344(.dina(n1407), .dinb(n1399), .dout(n1408));
  jor  g01345(.dina(n416), .dinb(n81), .dout(n1409));
  jand g01346(.dina(n1409), .dinb(n371), .dout(n1410));
  jand g01347(.dina(n707), .dinb(n529), .dout(n1411));
  jand g01348(.dina(n882), .dinb(n641), .dout(n1412));
  jand g01349(.dina(n1412), .dinb(n1411), .dout(n1413));
  jand g01350(.dina(n1413), .dinb(n1410), .dout(n1414));
  jand g01351(.dina(n877), .dinb(n384), .dout(n1415));
  jand g01352(.dina(n817), .dinb(n678), .dout(n1416));
  jand g01353(.dina(n1416), .dinb(n1306), .dout(n1417));
  jand g01354(.dina(n1417), .dinb(n1415), .dout(n1418));
  jand g01355(.dina(n1418), .dinb(n1414), .dout(n1419));
  jand g01356(.dina(n1419), .dinb(n1408), .dout(n1420));
  jand g01357(.dina(n675), .dinb(n238), .dout(n1421));
  jand g01358(.dina(n1153), .dinb(n719), .dout(n1422));
  jand g01359(.dina(n1422), .dinb(n1421), .dout(n1423));
  jand g01360(.dina(n1178), .dinb(n712), .dout(n1424));
  jand g01361(.dina(n1424), .dinb(n1285), .dout(n1425));
  jand g01362(.dina(n1425), .dinb(n1423), .dout(n1426));
  jand g01363(.dina(n583), .dinb(n231), .dout(n1427));
  jand g01364(.dina(n515), .dinb(n130), .dout(n1428));
  jand g01365(.dina(n1428), .dinb(n598), .dout(n1429));
  jand g01366(.dina(n1429), .dinb(n1427), .dout(n1430));
  jand g01367(.dina(n1430), .dinb(n1426), .dout(n1431));
  jand g01368(.dina(n1264), .dinb(n516), .dout(n1432));
  jand g01369(.dina(n1432), .dinb(n615), .dout(n1433));
  jand g01370(.dina(n1433), .dinb(n752), .dout(n1434));
  jand g01371(.dina(n1314), .dinb(n276), .dout(n1435));
  jand g01372(.dina(n1435), .dinb(n820), .dout(n1436));
  jand g01373(.dina(n434), .dinb(n375), .dout(n1437));
  jand g01374(.dina(n1437), .dinb(n982), .dout(n1438));
  jand g01375(.dina(n1438), .dinb(n1436), .dout(n1439));
  jand g01376(.dina(n1439), .dinb(n1434), .dout(n1440));
  jand g01377(.dina(n1440), .dinb(n1431), .dout(n1441));
  jand g01378(.dina(n1441), .dinb(n1420), .dout(n1442));
  jand g01379(.dina(n1442), .dinb(n1395), .dout(n1443));
  jand g01380(.dina(n1443), .dinb(n1073), .dout(n1444));
  jnot g01381(.din(n1444), .dout(n1445));
  jand g01382(.dina(n1445), .dinb(n1343), .dout(n1446));
  jand g01383(.dina(n508), .dinb(n268), .dout(n1447));
  jand g01384(.dina(n1447), .dinb(n643), .dout(n1448));
  jand g01385(.dina(n1448), .dinb(n1182), .dout(n1449));
  jand g01386(.dina(n993), .dinb(n467), .dout(n1450));
  jand g01387(.dina(n1450), .dinb(n427), .dout(n1451));
  jand g01388(.dina(n562), .dinb(n409), .dout(n1452));
  jand g01389(.dina(n1452), .dinb(n258), .dout(n1453));
  jand g01390(.dina(n759), .dinb(n614), .dout(n1454));
  jand g01391(.dina(n1454), .dinb(n1137), .dout(n1455));
  jand g01392(.dina(n1455), .dinb(n1453), .dout(n1456));
  jand g01393(.dina(n1456), .dinb(n1451), .dout(n1457));
  jand g01394(.dina(n1457), .dinb(n1449), .dout(n1458));
  jand g01395(.dina(n909), .dinb(n270), .dout(n1459));
  jand g01396(.dina(n1459), .dinb(n827), .dout(n1460));
  jand g01397(.dina(n817), .dinb(n605), .dout(n1461));
  jand g01398(.dina(n1461), .dinb(n492), .dout(n1462));
  jand g01399(.dina(n1462), .dinb(n1460), .dout(n1463));
  jand g01400(.dina(n1463), .dinb(n1180), .dout(n1464));
  jand g01401(.dina(n382), .dinb(n365), .dout(n1465));
  jand g01402(.dina(n1465), .dinb(n751), .dout(n1466));
  jand g01403(.dina(n1314), .dinb(n687), .dout(n1467));
  jand g01404(.dina(n1467), .dinb(n1295), .dout(n1468));
  jand g01405(.dina(n1468), .dinb(n1466), .dout(n1469));
  jand g01406(.dina(n711), .dinb(n214), .dout(n1470));
  jand g01407(.dina(n1470), .dinb(n1024), .dout(n1471));
  jand g01408(.dina(n1471), .dinb(n1160), .dout(n1472));
  jand g01409(.dina(n693), .dinb(n490), .dout(n1473));
  jand g01410(.dina(n950), .dinb(n286), .dout(n1474));
  jand g01411(.dina(n675), .dinb(n180), .dout(n1475));
  jand g01412(.dina(n1475), .dinb(n1474), .dout(n1476));
  jand g01413(.dina(n1476), .dinb(n1473), .dout(n1477));
  jand g01414(.dina(n1477), .dinb(n1472), .dout(n1478));
  jand g01415(.dina(n1478), .dinb(n1469), .dout(n1479));
  jand g01416(.dina(n1479), .dinb(n1464), .dout(n1480));
  jand g01417(.dina(n1480), .dinb(n1458), .dout(n1481));
  jnot g01418(.din(n439), .dout(n1482));
  jor  g01419(.dina(n856), .dinb(n1482), .dout(n1483));
  jnot g01420(.din(n1483), .dout(n1484));
  jand g01421(.dina(n1484), .dinb(n924), .dout(n1485));
  jand g01422(.dina(n1485), .dinb(n612), .dout(n1486));
  jand g01423(.dina(n897), .dinb(n842), .dout(n1487));
  jand g01424(.dina(n1487), .dinb(n82), .dout(n1488));
  jand g01425(.dina(n249), .dinb(n103), .dout(n1489));
  jand g01426(.dina(n1489), .dinb(n1488), .dout(n1490));
  jand g01427(.dina(n1383), .dinb(n1205), .dout(n1491));
  jand g01428(.dina(n385), .dinb(n113), .dout(n1492));
  jand g01429(.dina(n1492), .dinb(n939), .dout(n1493));
  jand g01430(.dina(n1493), .dinb(n1491), .dout(n1494));
  jand g01431(.dina(n1494), .dinb(n1490), .dout(n1495));
  jand g01432(.dina(n1495), .dinb(n1486), .dout(n1496));
  jand g01433(.dina(n965), .dinb(n598), .dout(n1497));
  jand g01434(.dina(n1497), .dinb(n815), .dout(n1498));
  jand g01435(.dina(n757), .dinb(n407), .dout(n1499));
  jand g01436(.dina(n1268), .dinb(n245), .dout(n1500));
  jand g01437(.dina(n1500), .dinb(n833), .dout(n1501));
  jand g01438(.dina(n1501), .dinb(n1499), .dout(n1502));
  jand g01439(.dina(n1502), .dinb(n1498), .dout(n1503));
  jand g01440(.dina(n876), .dinb(n224), .dout(n1504));
  jand g01441(.dina(n1504), .dinb(n1296), .dout(n1505));
  jand g01442(.dina(n536), .dinb(n120), .dout(n1506));
  jand g01443(.dina(n529), .dinb(n372), .dout(n1507));
  jand g01444(.dina(n1507), .dinb(n1506), .dout(n1508));
  jand g01445(.dina(n1508), .dinb(n1505), .dout(n1509));
  jand g01446(.dina(n583), .dinb(n505), .dout(n1510));
  jand g01447(.dina(n1510), .dinb(n386), .dout(n1511));
  jand g01448(.dina(n959), .dinb(n417), .dout(n1512));
  jand g01449(.dina(n1512), .dinb(n208), .dout(n1513));
  jand g01450(.dina(n1513), .dinb(n1511), .dout(n1514));
  jand g01451(.dina(n1514), .dinb(n1509), .dout(n1515));
  jand g01452(.dina(n1515), .dinb(n1503), .dout(n1516));
  jand g01453(.dina(n1516), .dinb(n1496), .dout(n1517));
  jand g01454(.dina(n1057), .dinb(n860), .dout(n1518));
  jor  g01455(.dina(n142), .dinb(n81), .dout(n1519));
  jand g01456(.dina(n494), .dinb(n262), .dout(n1520));
  jand g01457(.dina(n1520), .dinb(n1519), .dout(n1521));
  jand g01458(.dina(n1521), .dinb(n1518), .dout(n1522));
  jand g01459(.dina(n1522), .dinb(n624), .dout(n1523));
  jand g01460(.dina(n717), .dinb(n543), .dout(n1524));
  jand g01461(.dina(n1524), .dinb(n888), .dout(n1525));
  jand g01462(.dina(n509), .dinb(n290), .dout(n1526));
  jand g01463(.dina(n1526), .dinb(n395), .dout(n1527));
  jand g01464(.dina(n707), .dinb(n404), .dout(n1528));
  jand g01465(.dina(n1528), .dinb(n648), .dout(n1529));
  jand g01466(.dina(n1529), .dinb(n1527), .dout(n1530));
  jand g01467(.dina(n1530), .dinb(n1525), .dout(n1531));
  jand g01468(.dina(n1531), .dinb(n1523), .dout(n1532));
  jand g01469(.dina(n472), .dinb(n314), .dout(n1533));
  jand g01470(.dina(n1533), .dinb(n340), .dout(n1534));
  jand g01471(.dina(n749), .dinb(n586), .dout(n1535));
  jand g01472(.dina(n357), .dinb(n288), .dout(n1536));
  jand g01473(.dina(n694), .dinb(n292), .dout(n1537));
  jand g01474(.dina(n1537), .dinb(n1536), .dout(n1538));
  jand g01475(.dina(n1538), .dinb(n1535), .dout(n1539));
  jand g01476(.dina(n1539), .dinb(n1534), .dout(n1540));
  jand g01477(.dina(n1040), .dinb(n174), .dout(n1541));
  jand g01478(.dina(n819), .dinb(n392), .dout(n1542));
  jand g01479(.dina(n1542), .dinb(n1541), .dout(n1543));
  jnot g01480(.din(n566), .dout(n1544));
  jor  g01481(.dina(n1143), .dinb(n1544), .dout(n1545));
  jnot g01482(.din(n1545), .dout(n1546));
  jand g01483(.dina(n1546), .dinb(n1099), .dout(n1547));
  jand g01484(.dina(n1547), .dinb(n1543), .dout(n1548));
  jand g01485(.dina(n671), .dinb(n667), .dout(n1549));
  jand g01486(.dina(n1549), .dinb(n134), .dout(n1550));
  jand g01487(.dina(n721), .dinb(n503), .dout(n1551));
  jand g01488(.dina(n432), .dinb(n276), .dout(n1552));
  jand g01489(.dina(n1552), .dinb(n1551), .dout(n1553));
  jand g01490(.dina(n1553), .dinb(n1550), .dout(n1554));
  jand g01491(.dina(n1554), .dinb(n1548), .dout(n1555));
  jand g01492(.dina(n1555), .dinb(n1540), .dout(n1556));
  jand g01493(.dina(n1556), .dinb(n1532), .dout(n1557));
  jand g01494(.dina(n1557), .dinb(n1517), .dout(n1558));
  jand g01495(.dina(n1558), .dinb(n1481), .dout(n1559));
  jnot g01496(.din(n1559), .dout(n1560));
  jand g01497(.dina(n1560), .dinb(n1445), .dout(n1561));
  jand g01498(.dina(n950), .dinb(n165), .dout(n1562));
  jand g01499(.dina(n1562), .dinb(n386), .dout(n1563));
  jand g01500(.dina(n1034), .dinb(n414), .dout(n1564));
  jand g01501(.dina(n626), .dinb(n262), .dout(n1565));
  jand g01502(.dina(n1565), .dinb(n1564), .dout(n1566));
  jnot g01503(.din(n716), .dout(n1567));
  jor  g01504(.dina(n1567), .dinb(n345), .dout(n1568));
  jnot g01505(.din(n1568), .dout(n1569));
  jand g01506(.dina(n1569), .dinb(n914), .dout(n1570));
  jand g01507(.dina(n1570), .dinb(n1566), .dout(n1571));
  jand g01508(.dina(n1571), .dinb(n1563), .dout(n1572));
  jand g01509(.dina(n324), .dinb(n245), .dout(n1573));
  jand g01510(.dina(n635), .dinb(n274), .dout(n1574));
  jand g01511(.dina(n1574), .dinb(n331), .dout(n1575));
  jand g01512(.dina(n1575), .dinb(n1573), .dout(n1576));
  jand g01513(.dina(n1221), .dinb(n92), .dout(n1577));
  jand g01514(.dina(n1314), .dinb(n993), .dout(n1578));
  jand g01515(.dina(n1578), .dinb(n1577), .dout(n1579));
  jand g01516(.dina(n759), .dinb(n177), .dout(n1580));
  jand g01517(.dina(n689), .dinb(n413), .dout(n1581));
  jand g01518(.dina(n1581), .dinb(n1580), .dout(n1582));
  jand g01519(.dina(n1582), .dinb(n1579), .dout(n1583));
  jand g01520(.dina(n1178), .dinb(n888), .dout(n1584));
  jand g01521(.dina(n1346), .dinb(n161), .dout(n1585));
  jand g01522(.dina(n1585), .dinb(n1475), .dout(n1586));
  jand g01523(.dina(n1586), .dinb(n1584), .dout(n1587));
  jand g01524(.dina(n1587), .dinb(n1583), .dout(n1588));
  jand g01525(.dina(n1588), .dinb(n1576), .dout(n1589));
  jand g01526(.dina(n1589), .dinb(n1572), .dout(n1590));
  jand g01527(.dina(n1047), .dinb(n979), .dout(n1591));
  jand g01528(.dina(n449), .dinb(n404), .dout(n1592));
  jand g01529(.dina(n1592), .dinb(n1591), .dout(n1593));
  jand g01530(.dina(n1040), .dinb(n377), .dout(n1594));
  jand g01531(.dina(n1594), .dinb(n1130), .dout(n1595));
  jand g01532(.dina(n1595), .dinb(n1593), .dout(n1596));
  jnot g01533(.din(n796), .dout(n1597));
  jand g01534(.dina(n1597), .dinb(n205), .dout(n1598));
  jand g01535(.dina(n1598), .dinb(n218), .dout(n1599));
  jand g01536(.dina(n893), .dinb(n817), .dout(n1600));
  jand g01537(.dina(n1600), .dinb(n1145), .dout(n1601));
  jand g01538(.dina(n1601), .dinb(n1599), .dout(n1602));
  jand g01539(.dina(n736), .dinb(n157), .dout(n1603));
  jand g01540(.dina(n1603), .dinb(n647), .dout(n1604));
  jand g01541(.dina(n1364), .dinb(n1204), .dout(n1605));
  jand g01542(.dina(n1605), .dinb(n1604), .dout(n1606));
  jand g01543(.dina(n1606), .dinb(n1602), .dout(n1607));
  jand g01544(.dina(n1607), .dinb(n1596), .dout(n1608));
  jnot g01545(.din(n1409), .dout(n1609));
  jor  g01546(.dina(n1609), .dinb(n1358), .dout(n1610));
  jnot g01547(.din(n1610), .dout(n1611));
  jand g01548(.dina(n909), .dinb(n476), .dout(n1612));
  jand g01549(.dina(n1612), .dinb(n82), .dout(n1613));
  jand g01550(.dina(n272), .dinb(n128), .dout(n1614));
  jnot g01551(.din(n1614), .dout(n1615));
  jand g01552(.dina(n965), .dinb(n184), .dout(n1616));
  jand g01553(.dina(n1616), .dinb(n1615), .dout(n1617));
  jand g01554(.dina(n1617), .dinb(n1613), .dout(n1618));
  jand g01555(.dina(n1618), .dinb(n1611), .dout(n1619));
  jand g01556(.dina(n1619), .dinb(n1114), .dout(n1620));
  jand g01557(.dina(n1620), .dinb(n1608), .dout(n1621));
  jand g01558(.dina(n1621), .dinb(n572), .dout(n1622));
  jand g01559(.dina(n1622), .dinb(n1590), .dout(n1623));
  jnot g01560(.din(n1623), .dout(n1624));
  jand g01561(.dina(n1624), .dinb(n1560), .dout(n1625));
  jor  g01562(.dina(n608), .dinb(n440), .dout(n1626));
  jnot g01563(.din(n1626), .dout(n1627));
  jand g01564(.dina(n467), .dinb(n352), .dout(n1628));
  jand g01565(.dina(n696), .dinb(n234), .dout(n1629));
  jand g01566(.dina(n1629), .dinb(n1628), .dout(n1630));
  jand g01567(.dina(n1630), .dinb(n1627), .dout(n1631));
  jand g01568(.dina(n228), .dinb(n190), .dout(n1632));
  jand g01569(.dina(n1632), .dinb(n1518), .dout(n1633));
  jnot g01570(.din(n1350), .dout(n1634));
  jor  g01571(.dina(n632), .dinb(n279), .dout(n1635));
  jor  g01572(.dina(n1635), .dinb(n426), .dout(n1636));
  jor  g01573(.dina(n1636), .dinb(n1634), .dout(n1637));
  jnot g01574(.din(n1637), .dout(n1638));
  jand g01575(.dina(n1638), .dinb(n1633), .dout(n1639));
  jand g01576(.dina(n1639), .dinb(n1631), .dout(n1640));
  jnot g01577(.din(n1357), .dout(n1641));
  jand g01578(.dina(n1066), .dinb(n270), .dout(n1642));
  jand g01579(.dina(n1642), .dinb(n1641), .dout(n1643));
  jand g01580(.dina(n888), .dinb(n857), .dout(n1644));
  jand g01581(.dina(n509), .dinb(n500), .dout(n1645));
  jand g01582(.dina(n1645), .dinb(n1644), .dout(n1646));
  jand g01583(.dina(n687), .dinb(n286), .dout(n1647));
  jand g01584(.dina(n1647), .dinb(n225), .dout(n1648));
  jand g01585(.dina(n1648), .dinb(n1646), .dout(n1649));
  jand g01586(.dina(n1649), .dinb(n1643), .dout(n1650));
  jand g01587(.dina(n366), .dinb(n354), .dout(n1651));
  jand g01588(.dina(n1167), .dinb(n751), .dout(n1652));
  jand g01589(.dina(n1652), .dinb(n1651), .dout(n1653));
  jand g01590(.dina(n938), .dinb(n93), .dout(n1654));
  jand g01591(.dina(n1654), .dinb(n1653), .dout(n1655));
  jand g01592(.dina(n1039), .dinb(n305), .dout(n1656));
  jand g01593(.dina(n1656), .dinb(n245), .dout(n1657));
  jand g01594(.dina(n529), .dinb(n404), .dout(n1658));
  jand g01595(.dina(n583), .dinb(n314), .dout(n1659));
  jand g01596(.dina(n1659), .dinb(n1658), .dout(n1660));
  jand g01597(.dina(n1660), .dinb(n1657), .dout(n1661));
  jand g01598(.dina(n1661), .dinb(n1655), .dout(n1662));
  jand g01599(.dina(n893), .dinb(n543), .dout(n1663));
  jand g01600(.dina(n643), .dinb(n329), .dout(n1664));
  jand g01601(.dina(n1664), .dinb(n1663), .dout(n1665));
  jand g01602(.dina(n802), .dinb(n384), .dout(n1666));
  jand g01603(.dina(n1666), .dinb(n1665), .dout(n1667));
  jand g01604(.dina(n461), .dinb(n1031), .dout(n1668));
  jand g01605(.dina(n1668), .dinb(n443), .dout(n1669));
  jand g01606(.dina(n1669), .dinb(n1164), .dout(n1670));
  jand g01607(.dina(n1670), .dinb(n1667), .dout(n1671));
  jand g01608(.dina(n1671), .dinb(n1662), .dout(n1672));
  jand g01609(.dina(n1672), .dinb(n1650), .dout(n1673));
  jand g01610(.dina(n1673), .dinb(n1640), .dout(n1674));
  jand g01611(.dina(n478), .dinb(n252), .dout(n1675));
  jand g01612(.dina(n712), .dinb(n533), .dout(n1676));
  jand g01613(.dina(n1676), .dinb(n1675), .dout(n1677));
  jand g01614(.dina(n1677), .dinb(n868), .dout(n1678));
  jnot g01615(.din(n1678), .dout(n1679));
  jand g01616(.dina(n770), .dinb(n274), .dout(n1680));
  jand g01617(.dina(n1680), .dinb(n527), .dout(n1681));
  jnot g01618(.din(n1681), .dout(n1682));
  jnot g01619(.din(n417), .dout(n1683));
  jand g01620(.dina(n235), .dinb(n389), .dout(n1684));
  jor  g01621(.dina(n912), .dinb(n1684), .dout(n1685));
  jor  g01622(.dina(n1685), .dinb(n1683), .dout(n1686));
  jor  g01623(.dina(n825), .dinb(n261), .dout(n1687));
  jand g01624(.dina(n462), .dinb(n371), .dout(n1688));
  jnot g01625(.din(n1688), .dout(n1689));
  jor  g01626(.dina(n1689), .dinb(n1687), .dout(n1690));
  jor  g01627(.dina(n1690), .dinb(n1686), .dout(n1691));
  jor  g01628(.dina(n1691), .dinb(n1682), .dout(n1692));
  jor  g01629(.dina(n1692), .dinb(n1679), .dout(n1693));
  jnot g01630(.din(n1270), .dout(n1694));
  jor  g01631(.dina(n1152), .dinb(n949), .dout(n1695));
  jor  g01632(.dina(n471), .dinb(n133), .dout(n1696));
  jor  g01633(.dina(n1696), .dinb(n1695), .dout(n1697));
  jor  g01634(.dina(n621), .dinb(n119), .dout(n1698));
  jand g01635(.dina(n614), .dinb(n439), .dout(n1699));
  jnot g01636(.din(n1699), .dout(n1700));
  jor  g01637(.dina(n1700), .dinb(n1698), .dout(n1701));
  jor  g01638(.dina(n1701), .dinb(n1697), .dout(n1702));
  jor  g01639(.dina(n1702), .dinb(n1694), .dout(n1703));
  jand g01640(.dina(n1231), .dinb(n359), .dout(n1704));
  jnot g01641(.din(n1704), .dout(n1705));
  jand g01642(.dina(n200), .dinb(n132), .dout(n1706));
  jor  g01643(.dina(n1706), .dinb(n718), .dout(n1707));
  jor  g01644(.dina(n873), .dinb(n774), .dout(n1708));
  jor  g01645(.dina(n1708), .dinb(n1707), .dout(n1709));
  jor  g01646(.dina(n1709), .dinb(n1705), .dout(n1710));
  jand g01647(.dina(n372), .dinb(n184), .dout(n1711));
  jnot g01648(.din(n1711), .dout(n1712));
  jor  g01649(.dina(n1712), .dinb(n489), .dout(n1713));
  jor  g01650(.dina(n964), .dinb(n291), .dout(n1714));
  jand g01651(.dina(n338), .dinb(n272), .dout(n1715));
  jand g01652(.dina(n338), .dinb(n219), .dout(n1716));
  jor  g01653(.dina(n1716), .dinb(n1715), .dout(n1717));
  jor  g01654(.dina(n1717), .dinb(n1714), .dout(n1718));
  jor  g01655(.dina(n1718), .dinb(n1713), .dout(n1719));
  jor  g01656(.dina(n1719), .dinb(n1710), .dout(n1720));
  jor  g01657(.dina(n1720), .dinb(n1703), .dout(n1721));
  jor  g01658(.dina(n1721), .dinb(n1693), .dout(n1722));
  jnot g01659(.din(n1722), .dout(n1723));
  jand g01660(.dina(n793), .dinb(n214), .dout(n1724));
  jand g01661(.dina(n909), .dinb(n853), .dout(n1725));
  jand g01662(.dina(n1725), .dinb(n1724), .dout(n1726));
  jand g01663(.dina(n997), .dinb(n365), .dout(n1727));
  jand g01664(.dina(n574), .dinb(n136), .dout(n1728));
  jand g01665(.dina(n1728), .dinb(n1727), .dout(n1729));
  jand g01666(.dina(n694), .dinb(n337), .dout(n1730));
  jand g01667(.dina(n819), .dinb(n290), .dout(n1731));
  jand g01668(.dina(n1731), .dinb(n1730), .dout(n1732));
  jand g01669(.dina(n1732), .dinb(n1729), .dout(n1733));
  jand g01670(.dina(n1733), .dinb(n1726), .dout(n1734));
  jand g01671(.dina(n451), .dinb(n340), .dout(n1735));
  jand g01672(.dina(n1735), .dinb(n1585), .dout(n1736));
  jand g01673(.dina(n619), .dinb(n260), .dout(n1737));
  jand g01674(.dina(n1737), .dinb(n197), .dout(n1738));
  jand g01675(.dina(n396), .dinb(n177), .dout(n1739));
  jand g01676(.dina(n1739), .dinb(n1738), .dout(n1740));
  jand g01677(.dina(n1740), .dinb(n1736), .dout(n1741));
  jand g01678(.dina(n1741), .dinb(n1734), .dout(n1742));
  jor  g01679(.dina(n881), .dinb(n156), .dout(n1743));
  jor  g01680(.dina(n670), .dinb(n102), .dout(n1744));
  jor  g01681(.dina(n1744), .dinb(n1743), .dout(n1745));
  jand g01682(.dina(n236), .dinb(n182), .dout(n1746));
  jor  g01683(.dina(n758), .dinb(n1746), .dout(n1747));
  jor  g01684(.dina(n846), .dinb(n604), .dout(n1748));
  jor  g01685(.dina(n1748), .dinb(n1747), .dout(n1749));
  jor  g01686(.dina(n1749), .dinb(n1745), .dout(n1750));
  jor  g01687(.dina(n748), .dinb(n107), .dout(n1751));
  jor  g01688(.dina(n1751), .dinb(n674), .dout(n1752));
  jor  g01689(.dina(n1263), .dinb(n1377), .dout(n1753));
  jnot g01690(.din(n756), .dout(n1754));
  jor  g01691(.dina(n1754), .dinb(n491), .dout(n1755));
  jor  g01692(.dina(n1755), .dinb(n1753), .dout(n1756));
  jor  g01693(.dina(n1756), .dinb(n1752), .dout(n1757));
  jor  g01694(.dina(n1757), .dinb(n1750), .dout(n1758));
  jnot g01695(.din(n1758), .dout(n1759));
  jand g01696(.dina(n824), .dinb(n635), .dout(n1760));
  jand g01697(.dina(n876), .dinb(n407), .dout(n1761));
  jand g01698(.dina(n1761), .dinb(n1760), .dout(n1762));
  jand g01699(.dina(n1541), .dinb(n558), .dout(n1763));
  jand g01700(.dina(n1763), .dinb(n1762), .dout(n1764));
  jand g01701(.dina(n516), .dinb(n304), .dout(n1765));
  jand g01702(.dina(n357), .dinb(n180), .dout(n1766));
  jand g01703(.dina(n1766), .dinb(n1765), .dout(n1767));
  jand g01704(.dina(n1014), .dinb(n311), .dout(n1768));
  jand g01705(.dina(n1768), .dinb(n983), .dout(n1769));
  jand g01706(.dina(n1769), .dinb(n1767), .dout(n1770));
  jand g01707(.dina(n1770), .dinb(n1764), .dout(n1771));
  jand g01708(.dina(n1771), .dinb(n1759), .dout(n1772));
  jand g01709(.dina(n1772), .dinb(n1742), .dout(n1773));
  jand g01710(.dina(n1773), .dinb(n1723), .dout(n1774));
  jand g01711(.dina(n1774), .dinb(n1674), .dout(n1775));
  jnot g01712(.din(n1775), .dout(n1776));
  jand g01713(.dina(n1776), .dinb(n1624), .dout(n1777));
  jand g01714(.dina(n805), .dinb(n317), .dout(n1778));
  jand g01715(.dina(n1778), .dinb(n1232), .dout(n1779));
  jand g01716(.dina(n857), .dinb(n759), .dout(n1780));
  jnot g01717(.din(n1780), .dout(n1781));
  jor  g01718(.dina(n1781), .dinb(n1312), .dout(n1782));
  jnot g01719(.din(n1782), .dout(n1783));
  jand g01720(.dina(n1783), .dinb(n1779), .dout(n1784));
  jand g01721(.dina(n1153), .dinb(n304), .dout(n1785));
  jand g01722(.dina(n1785), .dinb(n1546), .dout(n1786));
  jand g01723(.dina(n467), .dinb(n290), .dout(n1787));
  jand g01724(.dina(n1787), .dinb(n1409), .dout(n1788));
  jand g01725(.dina(n1788), .dinb(n1786), .dout(n1789));
  jand g01726(.dina(n1789), .dinb(n1784), .dout(n1790));
  jand g01727(.dina(n1790), .dinb(n1740), .dout(n1791));
  jand g01728(.dina(n542), .dinb(n184), .dout(n1792));
  jand g01729(.dina(n1792), .dinb(n694), .dout(n1793));
  jand g01730(.dina(n414), .dinb(n194), .dout(n1794));
  jand g01731(.dina(n1794), .dinb(n979), .dout(n1795));
  jand g01732(.dina(n993), .dinb(n262), .dout(n1796));
  jand g01733(.dina(n643), .dinb(n478), .dout(n1797));
  jand g01734(.dina(n1797), .dinb(n1796), .dout(n1798));
  jand g01735(.dina(n1798), .dinb(n1795), .dout(n1799));
  jand g01736(.dina(n1799), .dinb(n1793), .dout(n1800));
  jand g01737(.dina(n509), .dinb(n499), .dout(n1801));
  jnot g01738(.din(n1801), .dout(n1802));
  jor  g01739(.dina(n1802), .dinb(n1637), .dout(n1803));
  jnot g01740(.din(n1803), .dout(n1804));
  jand g01741(.dina(n1492), .dinb(n1349), .dout(n1805));
  jand g01742(.dina(n1805), .dinb(n1524), .dout(n1806));
  jand g01743(.dina(n1806), .dinb(n1488), .dout(n1807));
  jand g01744(.dina(n1807), .dinb(n1804), .dout(n1808));
  jand g01745(.dina(n1808), .dinb(n1800), .dout(n1809));
  jand g01746(.dina(n1809), .dinb(n1791), .dout(n1810));
  jand g01747(.dina(n330), .dinb(n165), .dout(n1811));
  jand g01748(.dina(n893), .dinb(n721), .dout(n1812));
  jand g01749(.dina(n1812), .dinb(n1811), .dout(n1813));
  jand g01750(.dina(n865), .dinb(n801), .dout(n1814));
  jand g01751(.dina(n678), .dinb(n340), .dout(n1815));
  jand g01752(.dina(n1815), .dinb(n1814), .dout(n1816));
  jand g01753(.dina(n1816), .dinb(n1813), .dout(n1817));
  jand g01754(.dina(n1615), .dinb(n409), .dout(n1818));
  jand g01755(.dina(n907), .dinb(n149), .dout(n1819));
  jand g01756(.dina(n1819), .dinb(n1818), .dout(n1820));
  jand g01757(.dina(n997), .dinb(n428), .dout(n1821));
  jand g01758(.dina(n1821), .dinb(n314), .dout(n1822));
  jand g01759(.dina(n1822), .dinb(n1042), .dout(n1823));
  jand g01760(.dina(n1823), .dinb(n1820), .dout(n1824));
  jand g01761(.dina(n1824), .dinb(n1817), .dout(n1825));
  jand g01762(.dina(n432), .dinb(n336), .dout(n1826));
  jand g01763(.dina(n1047), .dinb(n578), .dout(n1827));
  jand g01764(.dina(n1827), .dinb(n1826), .dout(n1828));
  jand g01765(.dina(n626), .dinb(n443), .dout(n1829));
  jand g01766(.dina(n815), .dinb(n739), .dout(n1830));
  jand g01767(.dina(n1830), .dinb(n1829), .dout(n1831));
  jand g01768(.dina(n1831), .dinb(n1828), .dout(n1832));
  jand g01769(.dina(n843), .dinb(n331), .dout(n1833));
  jand g01770(.dina(n1833), .dinb(n527), .dout(n1834));
  jand g01771(.dina(n1834), .dinb(n771), .dout(n1835));
  jand g01772(.dina(n1090), .dinb(n794), .dout(n1836));
  jand g01773(.dina(n1836), .dinb(n1470), .dout(n1837));
  jand g01774(.dina(n1837), .dinb(n1835), .dout(n1838));
  jand g01775(.dina(n1838), .dinb(n1832), .dout(n1839));
  jand g01776(.dina(n367), .dinb(n143), .dout(n1840));
  jand g01777(.dina(n1295), .dinb(n853), .dout(n1841));
  jand g01778(.dina(n1841), .dinb(n1840), .dout(n1842));
  jand g01779(.dina(n1842), .dinb(n1399), .dout(n1843));
  jand g01780(.dina(n696), .dinb(n481), .dout(n1844));
  jand g01781(.dina(n1844), .dinb(n1474), .dout(n1845));
  jand g01782(.dina(n462), .dinb(n391), .dout(n1846));
  jand g01783(.dina(n967), .dinb(n434), .dout(n1847));
  jand g01784(.dina(n1847), .dinb(n1846), .dout(n1848));
  jand g01785(.dina(n1848), .dinb(n1845), .dout(n1849));
  jand g01786(.dina(n1066), .dinb(n847), .dout(n1850));
  jand g01787(.dina(n817), .dinb(n228), .dout(n1851));
  jand g01788(.dina(n1851), .dinb(n1850), .dout(n1852));
  jand g01789(.dina(n1641), .dinb(n305), .dout(n1853));
  jand g01790(.dina(n500), .dinb(n472), .dout(n1854));
  jand g01791(.dina(n1854), .dinb(n1853), .dout(n1855));
  jand g01792(.dina(n1855), .dinb(n1852), .dout(n1856));
  jand g01793(.dina(n1856), .dinb(n1849), .dout(n1857));
  jand g01794(.dina(n1857), .dinb(n1843), .dout(n1858));
  jand g01795(.dina(n1858), .dinb(n1839), .dout(n1859));
  jand g01796(.dina(n1859), .dinb(n1825), .dout(n1860));
  jand g01797(.dina(n1860), .dinb(n1810), .dout(n1861));
  jnot g01798(.din(n1861), .dout(n1862));
  jand g01799(.dina(n1862), .dinb(n1776), .dout(n1863));
  jand g01800(.dina(n687), .dinb(n329), .dout(n1864));
  jand g01801(.dina(n1864), .dinb(n826), .dout(n1865));
  jand g01802(.dina(n595), .dinb(n450), .dout(n1866));
  jand g01803(.dina(n1866), .dinb(n205), .dout(n1867));
  jand g01804(.dina(n1039), .dinb(n483), .dout(n1868));
  jand g01805(.dina(n1868), .dinb(n833), .dout(n1869));
  jand g01806(.dina(n1869), .dinb(n1867), .dout(n1870));
  jand g01807(.dina(n1870), .dinb(n1865), .dout(n1871));
  jand g01808(.dina(n396), .dinb(n252), .dout(n1872));
  jand g01809(.dina(n1872), .dinb(n1231), .dout(n1873));
  jand g01810(.dina(n696), .dinb(n325), .dout(n1874));
  jand g01811(.dina(n1874), .dinb(n1040), .dout(n1875));
  jand g01812(.dina(n1875), .dinb(n1873), .dout(n1876));
  jand g01813(.dina(n880), .dinb(n384), .dout(n1877));
  jand g01814(.dina(n1435), .dinb(n478), .dout(n1878));
  jand g01815(.dina(n1878), .dinb(n1877), .dout(n1879));
  jand g01816(.dina(n1879), .dinb(n1876), .dout(n1880));
  jand g01817(.dina(n348), .dinb(n177), .dout(n1881));
  jand g01818(.dina(n1881), .dinb(n1250), .dout(n1882));
  jand g01819(.dina(n1882), .dinb(n1405), .dout(n1883));
  jand g01820(.dina(n857), .dinb(n532), .dout(n1884));
  jand g01821(.dina(n736), .dinb(n161), .dout(n1885));
  jand g01822(.dina(n1885), .dinb(n1884), .dout(n1886));
  jand g01823(.dina(n200), .dinb(n219), .dout(n1887));
  jor  g01824(.dina(n1614), .dinb(n1887), .dout(n1888));
  jnot g01825(.din(n1888), .dout(n1889));
  jand g01826(.dina(n1889), .dinb(n1506), .dout(n1890));
  jand g01827(.dina(n1890), .dinb(n1886), .dout(n1891));
  jand g01828(.dina(n1891), .dinb(n1883), .dout(n1892));
  jand g01829(.dina(n1892), .dinb(n1880), .dout(n1893));
  jand g01830(.dina(n1893), .dinb(n1871), .dout(n1894));
  jand g01831(.dina(n926), .dinb(n527), .dout(n1895));
  jand g01832(.dina(n1519), .dinb(n367), .dout(n1896));
  jand g01833(.dina(n1896), .dinb(n1895), .dout(n1897));
  jand g01834(.dina(n907), .dinb(n470), .dout(n1898));
  jand g01835(.dina(n913), .dinb(n481), .dout(n1899));
  jand g01836(.dina(n759), .dinb(n703), .dout(n1900));
  jand g01837(.dina(n1900), .dinb(n1899), .dout(n1901));
  jand g01838(.dina(n1901), .dinb(n1898), .dout(n1902));
  jand g01839(.dina(n1902), .dinb(n1897), .dout(n1903));
  jand g01840(.dina(n1346), .dinb(n492), .dout(n1904));
  jand g01841(.dina(n993), .dinb(n801), .dout(n1905));
  jand g01842(.dina(n1905), .dinb(n1904), .dout(n1906));
  jand g01843(.dina(n950), .dinb(n853), .dout(n1907));
  jand g01844(.dina(n1907), .dinb(n1306), .dout(n1908));
  jand g01845(.dina(n1908), .dinb(n1906), .dout(n1909));
  jand g01846(.dina(n1550), .dinb(n1183), .dout(n1910));
  jand g01847(.dina(n1910), .dinb(n1909), .dout(n1911));
  jand g01848(.dina(n391), .dinb(n157), .dout(n1912));
  jand g01849(.dina(n860), .dinb(n655), .dout(n1913));
  jand g01850(.dina(n1913), .dinb(n707), .dout(n1914));
  jand g01851(.dina(n1914), .dinb(n1912), .dout(n1915));
  jand g01852(.dina(n445), .dinb(n130), .dout(n1916));
  jand g01853(.dina(n1916), .dinb(n1627), .dout(n1917));
  jand g01854(.dina(n1917), .dinb(n1299), .dout(n1918));
  jand g01855(.dina(n1918), .dinb(n1915), .dout(n1919));
  jand g01856(.dina(n1919), .dinb(n1911), .dout(n1920));
  jand g01857(.dina(n1920), .dinb(n1903), .dout(n1921));
  jand g01858(.dina(n551), .dinb(n395), .dout(n1922));
  jand g01859(.dina(n1922), .dinb(n197), .dout(n1923));
  jand g01860(.dina(n622), .dinb(n228), .dout(n1924));
  jand g01861(.dina(n1924), .dinb(n717), .dout(n1925));
  jand g01862(.dina(n1925), .dinb(n1923), .dout(n1926));
  jand g01863(.dina(n882), .dinb(n517), .dout(n1927));
  jand g01864(.dina(n843), .dinb(n317), .dout(n1928));
  jand g01865(.dina(n1928), .dinb(n1927), .dout(n1929));
  jand g01866(.dina(n817), .dinb(n503), .dout(n1930));
  jand g01867(.dina(n1930), .dinb(n812), .dout(n1931));
  jand g01868(.dina(n1931), .dinb(n1929), .dout(n1932));
  jor  g01869(.dina(n642), .dinb(n403), .dout(n1933));
  jnot g01870(.din(n1933), .dout(n1934));
  jand g01871(.dina(n1934), .dinb(n558), .dout(n1935));
  jand g01872(.dina(n1935), .dinb(n1785), .dout(n1936));
  jand g01873(.dina(n1936), .dinb(n1932), .dout(n1937));
  jand g01874(.dina(n1937), .dinb(n1926), .dout(n1938));
  jand g01875(.dina(n1014), .dinb(n612), .dout(n1939));
  jand g01876(.dina(n815), .dinb(n1031), .dout(n1940));
  jand g01877(.dina(n1940), .dinb(n1939), .dout(n1941));
  jand g01878(.dina(n431), .dinb(n238), .dout(n1942));
  jand g01879(.dina(n1731), .dinb(n606), .dout(n1943));
  jand g01880(.dina(n1943), .dinb(n1942), .dout(n1944));
  jand g01881(.dina(n1944), .dinb(n1941), .dout(n1945));
  jand g01882(.dina(n1142), .dinb(n423), .dout(n1946));
  jand g01883(.dina(n692), .dinb(n336), .dout(n1947));
  jand g01884(.dina(n467), .dinb(n385), .dout(n1948));
  jand g01885(.dina(n1948), .dinb(n1947), .dout(n1949));
  jand g01886(.dina(n1949), .dinb(n835), .dout(n1950));
  jand g01887(.dina(n1950), .dinb(n1946), .dout(n1951));
  jand g01888(.dina(n1951), .dinb(n1945), .dout(n1952));
  jand g01889(.dina(n1952), .dinb(n1938), .dout(n1953));
  jand g01890(.dina(n1953), .dinb(n1921), .dout(n1954));
  jand g01891(.dina(n1954), .dinb(n1894), .dout(n1955));
  jnot g01892(.din(n1955), .dout(n1956));
  jand g01893(.dina(n1956), .dinb(n1862), .dout(n1957));
  jand g01894(.dina(n392), .dinb(n377), .dout(n1958));
  jand g01895(.dina(n988), .dinb(n486), .dout(n1959));
  jand g01896(.dina(n703), .dinb(n322), .dout(n1960));
  jand g01897(.dina(n1960), .dinb(n1959), .dout(n1961));
  jand g01898(.dina(n1961), .dinb(n1958), .dout(n1962));
  jand g01899(.dina(n786), .dinb(n551), .dout(n1963));
  jand g01900(.dina(n1963), .dinb(n574), .dout(n1964));
  jand g01901(.dina(n997), .dinb(n284), .dout(n1965));
  jand g01902(.dina(n1965), .dinb(n246), .dout(n1966));
  jand g01903(.dina(n633), .dinb(n418), .dout(n1967));
  jand g01904(.dina(n721), .dinb(n197), .dout(n1968));
  jand g01905(.dina(n1968), .dinb(n1967), .dout(n1969));
  jand g01906(.dina(n1969), .dinb(n1966), .dout(n1970));
  jand g01907(.dina(n1970), .dinb(n1964), .dout(n1971));
  jand g01908(.dina(n1971), .dinb(n1962), .dout(n1972));
  jand g01909(.dina(n874), .dinb(n641), .dout(n1973));
  jand g01910(.dina(n1973), .dinb(n130), .dout(n1974));
  jand g01911(.dina(n508), .dinb(n280), .dout(n1975));
  jand g01912(.dina(n671), .dinb(n346), .dout(n1976));
  jand g01913(.dina(n1976), .dinb(n757), .dout(n1977));
  jand g01914(.dina(n1977), .dinb(n1975), .dout(n1978));
  jand g01915(.dina(n1978), .dinb(n1974), .dout(n1979));
  jand g01916(.dina(n292), .dinb(n262), .dout(n1980));
  jand g01917(.dina(n1980), .dinb(n753), .dout(n1981));
  jand g01918(.dina(n1787), .dinb(n771), .dout(n1982));
  jand g01919(.dina(n1982), .dinb(n1981), .dout(n1983));
  jand g01920(.dina(n583), .dinb(n276), .dout(n1984));
  jand g01921(.dina(n1984), .dinb(n352), .dout(n1985));
  jand g01922(.dina(n909), .dinb(n146), .dout(n1986));
  jand g01923(.dina(n461), .dinb(n331), .dout(n1987));
  jand g01924(.dina(n1987), .dinb(n1986), .dout(n1988));
  jand g01925(.dina(n1988), .dinb(n1985), .dout(n1989));
  jand g01926(.dina(n1989), .dinb(n1983), .dout(n1990));
  jnot g01927(.din(n1743), .dout(n1991));
  jand g01928(.dina(n1221), .dinb(n708), .dout(n1992));
  jand g01929(.dina(n1992), .dinb(n1881), .dout(n1993));
  jand g01930(.dina(n1993), .dinb(n1991), .dout(n1994));
  jnot g01931(.din(n1753), .dout(n1995));
  jor  g01932(.dina(n469), .dinb(n227), .dout(n1996));
  jnot g01933(.din(n1996), .dout(n1997));
  jand g01934(.dina(n1997), .dinb(n1995), .dout(n1998));
  jand g01935(.dina(n1998), .dinb(n1584), .dout(n1999));
  jand g01936(.dina(n1999), .dinb(n1994), .dout(n2000));
  jand g01937(.dina(n2000), .dinb(n1990), .dout(n2001));
  jand g01938(.dina(n2001), .dinb(n1979), .dout(n2002));
  jand g01939(.dina(n2002), .dinb(n1972), .dout(n2003));
  jnot g01940(.din(n1695), .dout(n2004));
  jand g01941(.dina(n365), .dinb(n340), .dout(n2005));
  jand g01942(.dina(n2005), .dinb(n842), .dout(n2006));
  jand g01943(.dina(n2006), .dinb(n2004), .dout(n2007));
  jand g01944(.dina(n605), .dinb(n414), .dout(n2008));
  jand g01945(.dina(n2008), .dinb(n926), .dout(n2009));
  jand g01946(.dina(n578), .dinb(n566), .dout(n2010));
  jand g01947(.dina(n481), .dinb(n288), .dout(n2011));
  jand g01948(.dina(n2011), .dinb(n2010), .dout(n2012));
  jand g01949(.dina(n2012), .dinb(n2009), .dout(n2013));
  jand g01950(.dina(n1040), .dinb(n492), .dout(n2014));
  jand g01951(.dina(n612), .dinb(n598), .dout(n2015));
  jand g01952(.dina(n2015), .dinb(n693), .dout(n2016));
  jand g01953(.dina(n2016), .dinb(n2014), .dout(n2017));
  jand g01954(.dina(n2017), .dinb(n2013), .dout(n2018));
  jand g01955(.dina(n2018), .dinb(n2007), .dout(n2019));
  jand g01956(.dina(n739), .dinb(n770), .dout(n2020));
  jand g01957(.dina(n2020), .dinb(n763), .dout(n2021));
  jand g01958(.dina(n700), .dinb(n120), .dout(n2022));
  jand g01959(.dina(n1039), .dinb(n252), .dout(n2023));
  jand g01960(.dina(n2023), .dinb(n2022), .dout(n2024));
  jand g01961(.dina(n1031), .dinb(n190), .dout(n2025));
  jand g01962(.dina(n1066), .dinb(n658), .dout(n2026));
  jand g01963(.dina(n2026), .dinb(n2025), .dout(n2027));
  jand g01964(.dina(n2027), .dinb(n2024), .dout(n2028));
  jand g01965(.dina(n2028), .dinb(n2021), .dout(n2029));
  jand g01966(.dina(n924), .dinb(n255), .dout(n2030));
  jand g01967(.dina(n675), .dinb(n505), .dout(n2031));
  jand g01968(.dina(n2031), .dinb(n2030), .dout(n2032));
  jand g01969(.dina(n1615), .dinb(n826), .dout(n2033));
  jand g01970(.dina(n465), .dinb(n249), .dout(n2034));
  jand g01971(.dina(n2034), .dinb(n2033), .dout(n2035));
  jand g01972(.dina(n1416), .dinb(n717), .dout(n2036));
  jand g01973(.dina(n2036), .dinb(n2035), .dout(n2037));
  jand g01974(.dina(n2037), .dinb(n2032), .dout(n2038));
  jand g01975(.dina(n2038), .dinb(n2029), .dout(n2039));
  jand g01976(.dina(n2039), .dinb(n2019), .dout(n2040));
  jand g01977(.dina(n1314), .dinb(n1047), .dout(n2041));
  jand g01978(.dina(n2041), .dinb(n1519), .dout(n2042));
  jand g01979(.dina(n423), .dinb(n375), .dout(n2043));
  jand g01980(.dina(n2043), .dinb(n858), .dout(n2044));
  jand g01981(.dina(n2044), .dinb(n2042), .dout(n2045));
  jand g01982(.dina(n359), .dinb(n274), .dout(n2046));
  jand g01983(.dina(n860), .dinb(n238), .dout(n2047));
  jand g01984(.dina(n2047), .dinb(n2046), .dout(n2048));
  jand g01985(.dina(n622), .dinb(n337), .dout(n2049));
  jand g01986(.dina(n2049), .dinb(n385), .dout(n2050));
  jand g01987(.dina(n2050), .dinb(n2048), .dout(n2051));
  jand g01988(.dina(n2051), .dinb(n2045), .dout(n2052));
  jand g01989(.dina(n431), .dinb(n343), .dout(n2053));
  jand g01990(.dina(n2053), .dinb(n1585), .dout(n2054));
  jand g01991(.dina(n2054), .dinb(n791), .dout(n2055));
  jand g01992(.dina(n993), .dinb(n607), .dout(n2056));
  jand g01993(.dina(n819), .dinb(n404), .dout(n2057));
  jand g01994(.dina(n2057), .dinb(n2056), .dout(n2058));
  jand g01995(.dina(n542), .dinb(n427), .dout(n2059));
  jand g01996(.dina(n2059), .dinb(n271), .dout(n2060));
  jand g01997(.dina(n2060), .dinb(n2058), .dout(n2061));
  jand g01998(.dina(n2061), .dinb(n2055), .dout(n2062));
  jand g01999(.dina(n2062), .dinb(n2052), .dout(n2063));
  jand g02000(.dina(n2063), .dinb(n1843), .dout(n2064));
  jand g02001(.dina(n2064), .dinb(n2040), .dout(n2065));
  jand g02002(.dina(n2065), .dinb(n2003), .dout(n2066));
  jnot g02003(.din(n2066), .dout(n2067));
  jand g02004(.dina(n2067), .dinb(n1956), .dout(n2068));
  jnot g02005(.din(n1631), .dout(n2069));
  jnot g02006(.din(n257), .dout(n2070));
  jor  g02007(.dina(n448), .dinb(n2070), .dout(n2071));
  jor  g02008(.dina(n1404), .dinb(n408), .dout(n2072));
  jor  g02009(.dina(n2072), .dinb(n2071), .dout(n2073));
  jnot g02010(.din(n414), .dout(n2074));
  jor  g02011(.dina(n702), .dinb(n2074), .dout(n2075));
  jor  g02012(.dina(n2075), .dinb(n797), .dout(n2076));
  jor  g02013(.dina(n502), .dinb(n283), .dout(n2077));
  jor  g02014(.dina(n2077), .dinb(n1996), .dout(n2078));
  jor  g02015(.dina(n2078), .dinb(n2076), .dout(n2079));
  jor  g02016(.dina(n2079), .dinb(n2073), .dout(n2080));
  jor  g02017(.dina(n2080), .dinb(n2069), .dout(n2081));
  jand g02018(.dina(n1221), .dinb(n1039), .dout(n2082));
  jand g02019(.dina(n2082), .dinb(n82), .dout(n2083));
  jnot g02020(.din(n2083), .dout(n2084));
  jor  g02021(.dina(n738), .dinb(n390), .dout(n2085));
  jor  g02022(.dina(n2085), .dinb(n1568), .dout(n2086));
  jand g02023(.dina(n532), .dinb(n499), .dout(n2087));
  jnot g02024(.din(n2087), .dout(n2088));
  jor  g02025(.dina(n376), .dinb(n316), .dout(n2089));
  jor  g02026(.dina(n2089), .dinb(n2088), .dout(n2090));
  jor  g02027(.dina(n2090), .dinb(n2086), .dout(n2091));
  jor  g02028(.dina(n2091), .dinb(n2084), .dout(n2092));
  jor  g02029(.dina(n2092), .dinb(n1758), .dout(n2093));
  jor  g02030(.dina(n2093), .dinb(n2081), .dout(n2094));
  jnot g02031(.din(n2094), .dout(n2095));
  jand g02032(.dina(n719), .dinb(n646), .dout(n2096));
  jand g02033(.dina(n2096), .dinb(n154), .dout(n2097));
  jand g02034(.dina(n2097), .dinb(n1865), .dout(n2098));
  jand g02035(.dina(n950), .dinb(n217), .dout(n2099));
  jand g02036(.dina(n2099), .dinb(n92), .dout(n2100));
  jand g02037(.dina(n801), .dinb(n494), .dout(n2101));
  jand g02038(.dina(n288), .dinb(n230), .dout(n2102));
  jand g02039(.dina(n2102), .dinb(n2101), .dout(n2103));
  jand g02040(.dina(n2103), .dinb(n2100), .dout(n2104));
  jand g02041(.dina(n2104), .dinb(n2098), .dout(n2105));
  jand g02042(.dina(n1615), .dinb(n445), .dout(n2106));
  jand g02043(.dina(n517), .dinb(n481), .dout(n2107));
  jand g02044(.dina(n817), .dinb(n805), .dout(n2108));
  jand g02045(.dina(n2108), .dinb(n2107), .dout(n2109));
  jand g02046(.dina(n2109), .dinb(n2106), .dout(n2110));
  jand g02047(.dina(n1641), .dinb(n1268), .dout(n2111));
  jand g02048(.dina(n2111), .dinb(n1249), .dout(n2112));
  jand g02049(.dina(n2112), .dinb(n769), .dout(n2113));
  jand g02050(.dina(n2113), .dinb(n2110), .dout(n2114));
  jand g02051(.dina(n2114), .dinb(n2105), .dout(n2115));
  jand g02052(.dina(n578), .dinb(n386), .dout(n2116));
  jand g02053(.dina(n2116), .dinb(n924), .dout(n2117));
  jand g02054(.dina(n715), .dinb(n595), .dout(n2118));
  jnot g02055(.din(n1368), .dout(n2119));
  jand g02056(.dina(n435), .dinb(n371), .dout(n2120));
  jand g02057(.dina(n2120), .dinb(n2119), .dout(n2121));
  jand g02058(.dina(n2121), .dinb(n2118), .dout(n2122));
  jand g02059(.dina(n2122), .dinb(n2117), .dout(n2123));
  jand g02060(.dina(n2123), .dinb(n1771), .dout(n2124));
  jand g02061(.dina(n2124), .dinb(n2115), .dout(n2125));
  jand g02062(.dina(n2125), .dinb(n2095), .dout(n2126));
  jand g02063(.dina(n2126), .dinb(n2064), .dout(n2127));
  jnot g02064(.din(n2127), .dout(n2128));
  jand g02065(.dina(n2128), .dinb(n2067), .dout(n2129));
  jand g02066(.dina(n959), .dinb(n255), .dout(n2130));
  jand g02067(.dina(n2130), .dinb(n1196), .dout(n2131));
  jand g02068(.dina(n1153), .dinb(n292), .dout(n2132));
  jand g02069(.dina(n2132), .dinb(n1078), .dout(n2133));
  jand g02070(.dina(n2133), .dinb(n2131), .dout(n2134));
  jand g02071(.dina(n997), .dinb(n897), .dout(n2135));
  jand g02072(.dina(n888), .dinb(n302), .dout(n2136));
  jand g02073(.dina(n2136), .dinb(n2135), .dout(n2137));
  jand g02074(.dina(n2137), .dinb(n1657), .dout(n2138));
  jand g02075(.dina(n2138), .dinb(n1681), .dout(n2139));
  jand g02076(.dina(n2139), .dinb(n2134), .dout(n2140));
  jand g02077(.dina(n367), .dinb(n309), .dout(n2141));
  jand g02078(.dina(n2141), .dinb(n715), .dout(n2142));
  jand g02079(.dina(n2142), .dinb(n1399), .dout(n2143));
  jand g02080(.dina(n1597), .dinb(n317), .dout(n2144));
  jand g02081(.dina(n2144), .dinb(n1082), .dout(n2145));
  jand g02082(.dina(n566), .dinb(n396), .dout(n2146));
  jand g02083(.dina(n2146), .dinb(n1284), .dout(n2147));
  jand g02084(.dina(n2147), .dinb(n2145), .dout(n2148));
  jand g02085(.dina(n2148), .dinb(n2143), .dout(n2149));
  jand g02086(.dina(n843), .dinb(n418), .dout(n2150));
  jand g02087(.dina(n965), .dinb(n445), .dout(n2151));
  jand g02088(.dina(n993), .dinb(n340), .dout(n2152));
  jand g02089(.dina(n2152), .dinb(n2151), .dout(n2153));
  jand g02090(.dina(n2153), .dinb(n2150), .dout(n2154));
  jand g02091(.dina(n424), .dinb(n221), .dout(n2155));
  jand g02092(.dina(n2155), .dinb(n1424), .dout(n2156));
  jand g02093(.dina(n1959), .dinb(n601), .dout(n2157));
  jand g02094(.dina(n2157), .dinb(n2156), .dout(n2158));
  jand g02095(.dina(n2158), .dinb(n2154), .dout(n2159));
  jand g02096(.dina(n1034), .dinb(n842), .dout(n2160));
  jand g02097(.dina(n595), .dinb(n304), .dout(n2161));
  jand g02098(.dina(n2161), .dinb(n2160), .dout(n2162));
  jand g02099(.dina(n2162), .dinb(n1306), .dout(n2163));
  jand g02100(.dina(n801), .dinb(n483), .dout(n2164));
  jand g02101(.dina(n2164), .dinb(n607), .dout(n2165));
  jand g02102(.dina(n2165), .dinb(n982), .dout(n2166));
  jand g02103(.dina(n2166), .dinb(n2163), .dout(n2167));
  jand g02104(.dina(n2167), .dinb(n2159), .dout(n2168));
  jand g02105(.dina(n2168), .dinb(n2149), .dout(n2169));
  jand g02106(.dina(n2169), .dinb(n2140), .dout(n2170));
  jand g02107(.dina(n646), .dinb(n407), .dout(n2171));
  jand g02108(.dina(n2171), .dinb(n819), .dout(n2172));
  jand g02109(.dina(n428), .dinb(n331), .dout(n2173));
  jand g02110(.dina(n641), .dinb(n383), .dout(n2174));
  jand g02111(.dina(n2174), .dinb(n2173), .dout(n2175));
  jand g02112(.dina(n2175), .dinb(n2172), .dout(n2176));
  jand g02113(.dina(n2176), .dinb(n199), .dout(n2177));
  jand g02114(.dina(n824), .dinb(n692), .dout(n2178));
  jand g02115(.dina(n1268), .dinb(n716), .dout(n2179));
  jand g02116(.dina(n413), .dinb(n268), .dout(n2180));
  jand g02117(.dina(n2180), .dinb(n2179), .dout(n2181));
  jand g02118(.dina(n2181), .dinb(n2178), .dout(n2182));
  jand g02119(.dina(n336), .dinb(n252), .dout(n2183));
  jand g02120(.dina(n696), .dinb(n505), .dout(n2184));
  jand g02121(.dina(n2184), .dinb(n1663), .dout(n2185));
  jand g02122(.dina(n2185), .dinb(n2183), .dout(n2186));
  jand g02123(.dina(n2186), .dinb(n2182), .dout(n2187));
  jand g02124(.dina(n2187), .dinb(n2177), .dout(n2188));
  jand g02125(.dina(n1167), .dinb(n721), .dout(n2189));
  jand g02126(.dina(n2189), .dinb(n736), .dout(n2190));
  jand g02127(.dina(n778), .dinb(n553), .dout(n2191));
  jand g02128(.dina(n805), .dinb(n749), .dout(n2192));
  jand g02129(.dina(n2192), .dinb(n515), .dout(n2193));
  jand g02130(.dina(n2193), .dinb(n2191), .dout(n2194));
  jand g02131(.dina(n2194), .dinb(n2190), .dout(n2195));
  jand g02132(.dina(n626), .dinb(n286), .dout(n2196));
  jand g02133(.dina(n472), .dinb(n461), .dout(n2197));
  jand g02134(.dina(n2197), .dinb(n2196), .dout(n2198));
  jand g02135(.dina(n2198), .dinb(n2041), .dout(n2199));
  jand g02136(.dina(n404), .dinb(n174), .dout(n2200));
  jand g02137(.dina(n2200), .dinb(n365), .dout(n2201));
  jand g02138(.dina(n228), .dinb(n205), .dout(n2202));
  jand g02139(.dina(n2202), .dinb(n605), .dout(n2203));
  jand g02140(.dina(n2203), .dinb(n2201), .dout(n2204));
  jand g02141(.dina(n2204), .dinb(n2199), .dout(n2205));
  jand g02142(.dina(n2205), .dinb(n2195), .dout(n2206));
  jand g02143(.dina(n2206), .dinb(n2188), .dout(n2207));
  jand g02144(.dina(n1641), .dinb(n533), .dout(n2208));
  jand g02145(.dina(n583), .dinb(n478), .dout(n2209));
  jand g02146(.dina(n2209), .dinb(n2208), .dout(n2210));
  jand g02147(.dina(n671), .dinb(n516), .dout(n2211));
  jand g02148(.dina(n694), .dinb(n562), .dout(n2212));
  jand g02149(.dina(n2212), .dinb(n2211), .dout(n2213));
  jand g02150(.dina(n2213), .dinb(n218), .dout(n2214));
  jand g02151(.dina(n2214), .dinb(n2210), .dout(n2215));
  jand g02152(.dina(n909), .dinb(n330), .dout(n2216));
  jand g02153(.dina(n612), .dinb(n557), .dout(n2217));
  jand g02154(.dina(n2217), .dinb(n2216), .dout(n2218));
  jand g02155(.dina(n826), .dinb(n409), .dout(n2219));
  jand g02156(.dina(n950), .dinb(n542), .dout(n2220));
  jand g02157(.dina(n2220), .dinb(n2219), .dout(n2221));
  jand g02158(.dina(n499), .dinb(n450), .dout(n2222));
  jand g02159(.dina(n2222), .dinb(n393), .dout(n2223));
  jand g02160(.dina(n2223), .dinb(n2221), .dout(n2224));
  jand g02161(.dina(n2224), .dinb(n2218), .dout(n2225));
  jnot g02162(.din(n1710), .dout(n2226));
  jand g02163(.dina(n481), .dinb(n427), .dout(n2227));
  jand g02164(.dina(n619), .dinb(n405), .dout(n2228));
  jand g02165(.dina(n2228), .dinb(n2227), .dout(n2229));
  jand g02166(.dina(n2229), .dinb(n771), .dout(n2230));
  jand g02167(.dina(n2230), .dinb(n2226), .dout(n2231));
  jand g02168(.dina(n2231), .dinb(n2225), .dout(n2232));
  jand g02169(.dina(n2232), .dinb(n2215), .dout(n2233));
  jand g02170(.dina(n2233), .dinb(n170), .dout(n2234));
  jand g02171(.dina(n2234), .dinb(n2207), .dout(n2235));
  jand g02172(.dina(n2235), .dinb(n2170), .dout(n2236));
  jnot g02173(.din(n2236), .dout(n2237));
  jand g02174(.dina(n2237), .dinb(n2128), .dout(n2238));
  jand g02175(.dina(n997), .dinb(n553), .dout(n2239));
  jand g02176(.dina(n1031), .dinb(n292), .dout(n2240));
  jand g02177(.dina(n2240), .dinb(n2239), .dout(n2241));
  jand g02178(.dina(n2241), .dinb(n2014), .dout(n2242));
  jand g02179(.dina(n736), .dinb(n643), .dout(n2243));
  jand g02180(.dina(n2243), .dinb(n239), .dout(n2244));
  jand g02181(.dina(n586), .dinb(n517), .dout(n2245));
  jand g02182(.dina(n2245), .dinb(n386), .dout(n2246));
  jand g02183(.dina(n2246), .dinb(n2103), .dout(n2247));
  jand g02184(.dina(n2247), .dinb(n2244), .dout(n2248));
  jand g02185(.dina(n2248), .dinb(n2242), .dout(n2249));
  jand g02186(.dina(n1231), .dinb(n543), .dout(n2250));
  jand g02187(.dina(n2250), .dinb(n721), .dout(n2251));
  jand g02188(.dina(n1039), .dinb(n371), .dout(n2252));
  jand g02189(.dina(n2252), .dinb(n354), .dout(n2253));
  jand g02190(.dina(n2253), .dinb(n2251), .dout(n2254));
  jand g02191(.dina(n533), .dinb(n336), .dout(n2255));
  jand g02192(.dina(n2255), .dinb(n770), .dout(n2256));
  jand g02193(.dina(n2256), .dinb(n2009), .dout(n2257));
  jand g02194(.dina(n2257), .dinb(n2254), .dout(n2258));
  jand g02195(.dina(n2041), .dinb(n1104), .dout(n2259));
  jand g02196(.dina(n2259), .dinb(n468), .dout(n2260));
  jnot g02197(.din(n1707), .dout(n2261));
  jand g02198(.dina(n478), .dinb(n197), .dout(n2262));
  jand g02199(.dina(n2262), .dinb(n2261), .dout(n2263));
  jand g02200(.dina(n751), .dinb(n290), .dout(n2264));
  jand g02201(.dina(n2264), .dinb(n393), .dout(n2265));
  jand g02202(.dina(n2265), .dinb(n2263), .dout(n2266));
  jand g02203(.dina(n2266), .dinb(n2260), .dout(n2267));
  jand g02204(.dina(n2267), .dinb(n2258), .dout(n2268));
  jand g02205(.dina(n2268), .dinb(n2249), .dout(n2269));
  jand g02206(.dina(n1295), .dinb(n136), .dout(n2270));
  jand g02207(.dina(n2270), .dinb(n2269), .dout(n2271));
  jor  g02208(.dina(n1013), .dinb(n1715), .dout(n2272));
  jor  g02209(.dina(n1754), .dinb(n625), .dout(n2273));
  jor  g02210(.dina(n2273), .dinb(n2272), .dout(n2274));
  jnot g02211(.din(n2274), .dout(n2275));
  jand g02212(.dina(n348), .dinb(n245), .dout(n2276));
  jand g02213(.dina(n2276), .dinb(n1305), .dout(n2277));
  jand g02214(.dina(n778), .dinb(n612), .dout(n2278));
  jand g02215(.dina(n2278), .dinb(n2053), .dout(n2279));
  jand g02216(.dina(n2279), .dinb(n2277), .dout(n2280));
  jand g02217(.dina(n2280), .dinb(n2275), .dout(n2281));
  jand g02218(.dina(n527), .dinb(n511), .dout(n2282));
  jand g02219(.dina(n2282), .dinb(n806), .dout(n2283));
  jand g02220(.dina(n2283), .dinb(n1249), .dout(n2284));
  jand g02221(.dina(n988), .dinb(n667), .dout(n2285));
  jand g02222(.dina(n2285), .dinb(n646), .dout(n2286));
  jand g02223(.dina(n633), .dinb(n260), .dout(n2287));
  jand g02224(.dina(n2287), .dinb(n745), .dout(n2288));
  jand g02225(.dina(n2288), .dinb(n2286), .dout(n2289));
  jand g02226(.dina(n2289), .dinb(n2284), .dout(n2290));
  jand g02227(.dina(n1153), .dinb(n499), .dout(n2291));
  jand g02228(.dina(n1597), .dinb(n711), .dout(n2292));
  jand g02229(.dina(n1615), .dinb(n1409), .dout(n2293));
  jand g02230(.dina(n2293), .dinb(n2292), .dout(n2294));
  jand g02231(.dina(n2294), .dinb(n2291), .dout(n2295));
  jand g02232(.dina(n2295), .dinb(n1736), .dout(n2296));
  jand g02233(.dina(n2296), .dinb(n2290), .dout(n2297));
  jand g02234(.dina(n2297), .dinb(n2281), .dout(n2298));
  jand g02235(.dina(n671), .dinb(n252), .dout(n2299));
  jand g02236(.dina(n2299), .dinb(n1259), .dout(n2300));
  jand g02237(.dina(n382), .dinb(n154), .dout(n2301));
  jand g02238(.dina(n2301), .dinb(n1082), .dout(n2302));
  jand g02239(.dina(n2302), .dinb(n2300), .dout(n2303));
  jand g02240(.dina(n694), .dinb(n304), .dout(n2304));
  jand g02241(.dina(n607), .dinb(n427), .dout(n2305));
  jand g02242(.dina(n2305), .dinb(n2304), .dout(n2306));
  jand g02243(.dina(n407), .dinb(n395), .dout(n2307));
  jand g02244(.dina(n2307), .dinb(n888), .dout(n2308));
  jand g02245(.dina(n619), .dinb(n120), .dout(n2309));
  jand g02246(.dina(n847), .dinb(n708), .dout(n2310));
  jand g02247(.dina(n2310), .dinb(n2309), .dout(n2311));
  jand g02248(.dina(n2311), .dinb(n2308), .dout(n2312));
  jand g02249(.dina(n2312), .dinb(n2306), .dout(n2313));
  jand g02250(.dina(n2313), .dinb(n2303), .dout(n2314));
  jand g02251(.dina(n1034), .dinb(n130), .dout(n2315));
  jand g02252(.dina(n441), .dinb(n224), .dout(n2316));
  jand g02253(.dina(n503), .dinb(n317), .dout(n2317));
  jand g02254(.dina(n2317), .dinb(n2316), .dout(n2318));
  jand g02255(.dina(n2318), .dinb(n2315), .dout(n2319));
  jand g02256(.dina(n434), .dinb(n146), .dout(n2320));
  jand g02257(.dina(n2320), .dinb(n843), .dout(n2321));
  jand g02258(.dina(n874), .dinb(n574), .dout(n2322));
  jand g02259(.dina(n583), .dinb(n385), .dout(n2323));
  jand g02260(.dina(n2323), .dinb(n2322), .dout(n2324));
  jand g02261(.dina(n2324), .dinb(n2321), .dout(n2325));
  jand g02262(.dina(n2325), .dinb(n2319), .dout(n2326));
  jand g02263(.dina(n302), .dinb(n149), .dout(n2327));
  jand g02264(.dina(n1760), .dinb(n1247), .dout(n2328));
  jand g02265(.dina(n2328), .dinb(n2327), .dout(n2329));
  jor  g02266(.dina(n1263), .dinb(n351), .dout(n2330));
  jor  g02267(.dina(n912), .dinb(n785), .dout(n2331));
  jor  g02268(.dina(n2331), .dinb(n2330), .dout(n2332));
  jor  g02269(.dina(n859), .dinb(n183), .dout(n2333));
  jor  g02270(.dina(n892), .dinb(n674), .dout(n2334));
  jor  g02271(.dina(n2334), .dinb(n2333), .dout(n2335));
  jor  g02272(.dina(n2335), .dinb(n2332), .dout(n2336));
  jnot g02273(.din(n2336), .dout(n2337));
  jand g02274(.dina(n2337), .dinb(n2329), .dout(n2338));
  jand g02275(.dina(n2338), .dinb(n2326), .dout(n2339));
  jand g02276(.dina(n2339), .dinb(n2314), .dout(n2340));
  jand g02277(.dina(n2340), .dinb(n2298), .dout(n2341));
  jand g02278(.dina(n2341), .dinb(n2271), .dout(n2342));
  jnot g02279(.din(n2342), .dout(n2343));
  jand g02280(.dina(n2343), .dinb(n2237), .dout(n2344));
  jand g02281(.dina(n443), .dinb(n404), .dout(n2345));
  jand g02282(.dina(n2345), .dinb(n708), .dout(n2346));
  jand g02283(.dina(n824), .dinb(n712), .dout(n2347));
  jand g02284(.dina(n470), .dinb(n305), .dout(n2348));
  jand g02285(.dina(n2348), .dinb(n2347), .dout(n2349));
  jand g02286(.dina(n2349), .dinb(n1402), .dout(n2350));
  jand g02287(.dina(n2350), .dinb(n2346), .dout(n2351));
  jand g02288(.dina(n2351), .dinb(n2295), .dout(n2352));
  jand g02289(.dina(n1034), .dinb(n763), .dout(n2353));
  jand g02290(.dina(n2353), .dinb(n926), .dout(n2354));
  jand g02291(.dina(n719), .dinb(n692), .dout(n2355));
  jand g02292(.dina(n2355), .dinb(n1778), .dout(n2356));
  jand g02293(.dina(n2356), .dinb(n1960), .dout(n2357));
  jand g02294(.dina(n2357), .dinb(n2354), .dout(n2358));
  jand g02295(.dina(n1066), .dinb(n865), .dout(n2359));
  jand g02296(.dina(n2359), .dinb(n697), .dout(n2360));
  jand g02297(.dina(n1039), .dinb(n515), .dout(n2361));
  jand g02298(.dina(n701), .dinb(n336), .dout(n2362));
  jand g02299(.dina(n2362), .dinb(n2361), .dout(n2363));
  jand g02300(.dina(n2363), .dinb(n2360), .dout(n2364));
  jand g02301(.dina(n1641), .dinb(n721), .dout(n2365));
  jand g02302(.dina(n2365), .dinb(n492), .dout(n2366));
  jand g02303(.dina(n786), .dinb(n467), .dout(n2367));
  jand g02304(.dina(n2367), .dinb(n815), .dout(n2368));
  jand g02305(.dina(n1221), .dinb(n707), .dout(n2369));
  jand g02306(.dina(n715), .dinb(n413), .dout(n2370));
  jand g02307(.dina(n2370), .dinb(n2369), .dout(n2371));
  jand g02308(.dina(n2371), .dinb(n2368), .dout(n2372));
  jand g02309(.dina(n2372), .dinb(n2366), .dout(n2373));
  jand g02310(.dina(n2373), .dinb(n2364), .dout(n2374));
  jand g02311(.dina(n2374), .dinb(n2358), .dout(n2375));
  jand g02312(.dina(n2375), .dinb(n2352), .dout(n2376));
  jand g02313(.dina(n1285), .dinb(n594), .dout(n2377));
  jand g02314(.dina(n675), .dinb(n633), .dout(n2378));
  jand g02315(.dina(n2378), .dinb(n2278), .dout(n2379));
  jand g02316(.dina(n2379), .dinb(n2377), .dout(n2380));
  jor  g02317(.dina(n1177), .dinb(n758), .dout(n2381));
  jnot g02318(.din(n2381), .dout(n2382));
  jand g02319(.dina(n2382), .dinb(n716), .dout(n2383));
  jand g02320(.dina(n643), .dinb(n562), .dout(n2384));
  jand g02321(.dina(n2384), .dinb(n842), .dout(n2385));
  jand g02322(.dina(n1047), .dinb(n407), .dout(n2386));
  jand g02323(.dina(n2386), .dinb(n1243), .dout(n2387));
  jand g02324(.dina(n2387), .dinb(n2385), .dout(n2388));
  jand g02325(.dina(n2388), .dinb(n2383), .dout(n2389));
  jand g02326(.dina(n2389), .dinb(n2380), .dout(n2390));
  jand g02327(.dina(n1040), .dinb(n325), .dout(n2391));
  jand g02328(.dina(n1346), .dinb(n997), .dout(n2392));
  jand g02329(.dina(n2392), .dinb(n2391), .dout(n2393));
  jand g02330(.dina(n1231), .dinb(n882), .dout(n2394));
  jand g02331(.dina(n1144), .dinb(n793), .dout(n2395));
  jand g02332(.dina(n2395), .dinb(n2394), .dout(n2396));
  jand g02333(.dina(n1930), .dinb(n1437), .dout(n2397));
  jand g02334(.dina(n2397), .dinb(n2396), .dout(n2398));
  jand g02335(.dina(n2398), .dinb(n2393), .dout(n2399));
  jand g02336(.dina(n1167), .dinb(n647), .dout(n2400));
  jand g02337(.dina(n619), .dinb(n598), .dout(n2401));
  jand g02338(.dina(n595), .dinb(n516), .dout(n2402));
  jand g02339(.dina(n2402), .dinb(n615), .dout(n2403));
  jand g02340(.dina(n2403), .dinb(n2401), .dout(n2404));
  jand g02341(.dina(n2404), .dinb(n2400), .dout(n2405));
  jand g02342(.dina(n2405), .dinb(n541), .dout(n2406));
  jand g02343(.dina(n2406), .dinb(n2399), .dout(n2407));
  jand g02344(.dina(n2407), .dinb(n2390), .dout(n2408));
  jand g02345(.dina(n2408), .dinb(n299), .dout(n2409));
  jand g02346(.dina(n2409), .dinb(n2376), .dout(n2410));
  jnot g02347(.din(n2410), .dout(n2411));
  jand g02348(.dina(n2411), .dinb(n2343), .dout(n2412));
  jand g02349(.dina(n926), .dinb(n284), .dout(n2413));
  jand g02350(.dina(n874), .dinb(n694), .dout(n2414));
  jand g02351(.dina(n2414), .dinb(n2413), .dout(n2415));
  jand g02352(.dina(n614), .dinb(n157), .dout(n2416));
  jand g02353(.dina(n2416), .dinb(n1435), .dout(n2417));
  jand g02354(.dina(n2417), .dinb(n2107), .dout(n2418));
  jand g02355(.dina(n2418), .dinb(n2415), .dout(n2419));
  jand g02356(.dina(n499), .dinb(n407), .dout(n2420));
  jand g02357(.dina(n527), .dinb(n165), .dout(n2421));
  jand g02358(.dina(n2421), .dinb(n2420), .dout(n2422));
  jand g02359(.dina(n492), .dinb(n290), .dout(n2423));
  jand g02360(.dina(n2423), .dinb(n620), .dout(n2424));
  jand g02361(.dina(n2424), .dinb(n2422), .dout(n2425));
  jand g02362(.dina(n913), .dinb(n503), .dout(n2426));
  jand g02363(.dina(n2426), .dinb(n154), .dout(n2427));
  jand g02364(.dina(n1184), .dinb(n739), .dout(n2428));
  jand g02365(.dina(n909), .dinb(n897), .dout(n2429));
  jand g02366(.dina(n2429), .dinb(n2428), .dout(n2430));
  jand g02367(.dina(n2430), .dinb(n2427), .dout(n2431));
  jand g02368(.dina(n2431), .dinb(n2425), .dout(n2432));
  jand g02369(.dina(n424), .dinb(n257), .dout(n2433));
  jand g02370(.dina(n1144), .dinb(n542), .dout(n2434));
  jand g02371(.dina(n2434), .dinb(n2433), .dout(n2435));
  jand g02372(.dina(n2435), .dinb(n473), .dout(n2436));
  jand g02373(.dina(n595), .dinb(n180), .dout(n2437));
  jand g02374(.dina(n1597), .dinb(n605), .dout(n2438));
  jand g02375(.dina(n2438), .dinb(n348), .dout(n2439));
  jand g02376(.dina(n2439), .dinb(n2437), .dout(n2440));
  jand g02377(.dina(n2440), .dinb(n2436), .dout(n2441));
  jand g02378(.dina(n2441), .dinb(n2432), .dout(n2442));
  jand g02379(.dina(n2442), .dinb(n2419), .dout(n2443));
  jand g02380(.dina(n794), .dinb(n436), .dout(n2444));
  jand g02381(.dina(n2444), .dinb(n769), .dout(n2445));
  jand g02382(.dina(n1727), .dinb(n689), .dout(n2446));
  jand g02383(.dina(n396), .dinb(n304), .dout(n2447));
  jand g02384(.dina(n2447), .dinb(n375), .dout(n2448));
  jand g02385(.dina(n2448), .dinb(n1399), .dout(n2449));
  jand g02386(.dina(n2449), .dinb(n2446), .dout(n2450));
  jand g02387(.dina(n2450), .dinb(n2445), .dout(n2451));
  jand g02388(.dina(n1135), .dinb(n1067), .dout(n2452));
  jand g02389(.dina(n1197), .dinb(n451), .dout(n2453));
  jand g02390(.dina(n2453), .dinb(n2452), .dout(n2454));
  jand g02391(.dina(n959), .dinb(n598), .dout(n2455));
  jand g02392(.dina(n2455), .dinb(n508), .dout(n2456));
  jand g02393(.dina(n817), .dinb(n770), .dout(n2457));
  jand g02394(.dina(n551), .dinb(n309), .dout(n2458));
  jand g02395(.dina(n2458), .dinb(n2457), .dout(n2459));
  jand g02396(.dina(n2459), .dinb(n2456), .dout(n2460));
  jand g02397(.dina(n2369), .dinb(n1663), .dout(n2461));
  jand g02398(.dina(n2461), .dinb(n2244), .dout(n2462));
  jand g02399(.dina(n2462), .dinb(n2460), .dout(n2463));
  jand g02400(.dina(n2463), .dinb(n2454), .dout(n2464));
  jand g02401(.dina(n2464), .dinb(n2451), .dout(n2465));
  jand g02402(.dina(n344), .dinb(n116), .dout(n2466));
  jor  g02403(.dina(n661), .dinb(n2466), .dout(n2467));
  jnot g02404(.din(n2467), .dout(n2468));
  jand g02405(.dina(n1641), .dinb(n1264), .dout(n2469));
  jand g02406(.dina(n801), .dinb(n553), .dout(n2470));
  jand g02407(.dina(n2470), .dinb(n2469), .dout(n2471));
  jand g02408(.dina(n2471), .dinb(n2468), .dout(n2472));
  jand g02409(.dina(n337), .dinb(n243), .dout(n2473));
  jand g02410(.dina(n2150), .dinb(n954), .dout(n2474));
  jand g02411(.dina(n2474), .dinb(n2473), .dout(n2475));
  jand g02412(.dina(n1128), .dinb(n1009), .dout(n2476));
  jand g02413(.dina(n1474), .dinb(n109), .dout(n2477));
  jand g02414(.dina(n2477), .dinb(n2476), .dout(n2478));
  jand g02415(.dina(n2478), .dinb(n2475), .dout(n2479));
  jand g02416(.dina(n2479), .dinb(n2472), .dout(n2480));
  jand g02417(.dina(n888), .dinb(n675), .dout(n2481));
  jand g02418(.dina(n2481), .dinb(n687), .dout(n2482));
  jand g02419(.dina(n1034), .dinb(n330), .dout(n2483));
  jand g02420(.dina(n847), .dinb(n371), .dout(n2484));
  jand g02421(.dina(n2484), .dinb(n2483), .dout(n2485));
  jand g02422(.dina(n2485), .dinb(n2482), .dout(n2486));
  jand g02423(.dina(n759), .dinb(n205), .dout(n2487));
  jand g02424(.dina(n2487), .dinb(n575), .dout(n2488));
  jand g02425(.dina(n805), .dinb(n260), .dout(n2489));
  jand g02426(.dina(n2489), .dinb(n1196), .dout(n2490));
  jand g02427(.dina(n2490), .dinb(n2488), .dout(n2491));
  jand g02428(.dina(n2491), .dinb(n2486), .dout(n2492));
  jand g02429(.dina(n2492), .dinb(n1662), .dout(n2493));
  jand g02430(.dina(n2493), .dinb(n2480), .dout(n2494));
  jand g02431(.dina(n2494), .dinb(n2465), .dout(n2495));
  jand g02432(.dina(n2495), .dinb(n2443), .dout(n2496));
  jnot g02433(.din(n2496), .dout(n2497));
  jand g02434(.dina(n2497), .dinb(n2411), .dout(n2498));
  jand g02435(.dina(n1184), .dinb(n633), .dout(n2499));
  jand g02436(.dina(n1615), .dinb(n586), .dout(n2500));
  jand g02437(.dina(n2500), .dinb(n2499), .dout(n2501));
  jand g02438(.dina(n2501), .dinb(n1840), .dout(n2502));
  jand g02439(.dina(n612), .dinb(n503), .dout(n2503));
  jand g02440(.dina(n467), .dinb(n280), .dout(n2504));
  jand g02441(.dina(n2504), .dinb(n2503), .dout(n2505));
  jand g02442(.dina(n2505), .dinb(n1738), .dout(n2506));
  jand g02443(.dina(n357), .dinb(n268), .dout(n2507));
  jand g02444(.dina(n2507), .dinb(n304), .dout(n2508));
  jand g02445(.dina(n2508), .dinb(n2383), .dout(n2509));
  jand g02446(.dina(n2509), .dinb(n2506), .dout(n2510));
  jand g02447(.dina(n2510), .dinb(n2502), .dout(n2511));
  jand g02448(.dina(n1066), .dinb(n897), .dout(n2512));
  jand g02449(.dina(n2512), .dinb(n366), .dout(n2513));
  jand g02450(.dina(n819), .dinb(n377), .dout(n2514));
  jand g02451(.dina(n711), .dinb(n529), .dout(n2515));
  jand g02452(.dina(n2515), .dinb(n2514), .dout(n2516));
  jand g02453(.dina(n924), .dinb(n756), .dout(n2517));
  jand g02454(.dina(n2517), .dinb(n312), .dout(n2518));
  jand g02455(.dina(n2518), .dinb(n2516), .dout(n2519));
  jand g02456(.dina(n2519), .dinb(n2513), .dout(n2520));
  jand g02457(.dina(n340), .dinb(n154), .dout(n2521));
  jand g02458(.dina(n721), .dinb(n417), .dout(n2522));
  jand g02459(.dina(n2522), .dinb(n509), .dout(n2523));
  jand g02460(.dina(n2523), .dinb(n2521), .dout(n2524));
  jnot g02461(.din(n1748), .dout(n2525));
  jand g02462(.dina(n1268), .dinb(n643), .dout(n2526));
  jand g02463(.dina(n2526), .dinb(n709), .dout(n2527));
  jand g02464(.dina(n2527), .dinb(n2525), .dout(n2528));
  jand g02465(.dina(n2528), .dinb(n2524), .dout(n2529));
  jand g02466(.dina(n2529), .dinb(n2520), .dout(n2530));
  jand g02467(.dina(n2530), .dinb(n986), .dout(n2531));
  jand g02468(.dina(n2531), .dinb(n2511), .dout(n2532));
  jand g02469(.dina(n876), .dinb(n751), .dout(n2533));
  jand g02470(.dina(n2533), .dinb(n1986), .dout(n2534));
  jand g02471(.dina(n2534), .dinb(n2183), .dout(n2535));
  jand g02472(.dina(n443), .dinb(n286), .dout(n2536));
  jand g02473(.dina(n2536), .dinb(n609), .dout(n2537));
  jand g02474(.dina(n486), .dinb(n82), .dout(n2538));
  jand g02475(.dina(n395), .dinb(n305), .dout(n2539));
  jand g02476(.dina(n2539), .dinb(n2538), .dout(n2540));
  jand g02477(.dina(n2540), .dinb(n2537), .dout(n2541));
  jand g02478(.dina(n2541), .dinb(n2535), .dout(n2542));
  jand g02479(.dina(n2542), .dinb(n2532), .dout(n2543));
  jand g02480(.dina(n1040), .dinb(n993), .dout(n2544));
  jand g02481(.dina(n626), .dinb(n418), .dout(n2545));
  jand g02482(.dina(n2545), .dinb(n2544), .dout(n2546));
  jand g02483(.dina(n449), .dinb(n292), .dout(n2547));
  jand g02484(.dina(n888), .dinb(n551), .dout(n2548));
  jand g02485(.dina(n2548), .dinb(n2547), .dout(n2549));
  jand g02486(.dina(n2549), .dinb(n2546), .dout(n2550));
  jand g02487(.dina(n860), .dinb(n801), .dout(n2551));
  jand g02488(.dina(n2551), .dinb(n2416), .dout(n2552));
  jand g02489(.dina(n2552), .dinb(n2324), .dout(n2553));
  jand g02490(.dina(n2553), .dinb(n2550), .dout(n2554));
  jand g02491(.dina(n598), .dinb(n290), .dout(n2555));
  jand g02492(.dina(n354), .dinb(n274), .dout(n2556));
  jand g02493(.dina(n409), .dinb(n324), .dout(n2557));
  jand g02494(.dina(n2557), .dinb(n2556), .dout(n2558));
  jand g02495(.dina(n2558), .dinb(n2555), .dout(n2559));
  jand g02496(.dina(n658), .dinb(n177), .dout(n2560));
  jand g02497(.dina(n392), .dinb(n180), .dout(n2561));
  jand g02498(.dina(n2561), .dinb(n423), .dout(n2562));
  jand g02499(.dina(n2562), .dinb(n2560), .dout(n2563));
  jand g02500(.dina(n557), .dinb(n371), .dout(n2564));
  jand g02501(.dina(n542), .dinb(n462), .dout(n2565));
  jand g02502(.dina(n2565), .dinb(n2564), .dout(n2566));
  jand g02503(.dina(n764), .dinb(n384), .dout(n2567));
  jand g02504(.dina(n2567), .dinb(n2566), .dout(n2568));
  jand g02505(.dina(n2568), .dinb(n2563), .dout(n2569));
  jand g02506(.dina(n2569), .dinb(n2559), .dout(n2570));
  jand g02507(.dina(n2570), .dinb(n2554), .dout(n2571));
  jand g02508(.dina(n646), .dinb(n689), .dout(n2572));
  jand g02509(.dina(n2572), .dinb(n245), .dout(n2573));
  jand g02510(.dina(n1346), .dinb(n424), .dout(n2574));
  jand g02511(.dina(n2574), .dinb(n500), .dout(n2575));
  jand g02512(.dina(n2575), .dinb(n2573), .dout(n2576));
  jand g02513(.dina(n2576), .dinb(n138), .dout(n2577));
  jand g02514(.dina(n959), .dinb(n494), .dout(n2578));
  jand g02515(.dina(n2578), .dinb(n1265), .dout(n2579));
  jnot g02516(.din(n1744), .dout(n2580));
  jand g02517(.dina(n2580), .dinb(n218), .dout(n2581));
  jand g02518(.dina(n2581), .dinb(n2579), .dout(n2582));
  jand g02519(.dina(n736), .dinb(n562), .dout(n2583));
  jand g02520(.dina(n391), .dinb(n270), .dout(n2584));
  jand g02521(.dina(n2584), .dinb(n2583), .dout(n2585));
  jand g02522(.dina(n532), .dinb(n481), .dout(n2586));
  jand g02523(.dina(n2586), .dinb(n432), .dout(n2587));
  jand g02524(.dina(n2587), .dinb(n2585), .dout(n2588));
  jand g02525(.dina(n2588), .dinb(n2582), .dout(n2589));
  jand g02526(.dina(n786), .dinb(n655), .dout(n2590));
  jand g02527(.dina(n913), .dinb(n346), .dout(n2591));
  jand g02528(.dina(n1221), .dinb(n1014), .dout(n2592));
  jand g02529(.dina(n2592), .dinb(n2591), .dout(n2593));
  jand g02530(.dina(n2593), .dinb(n2590), .dout(n2594));
  jand g02531(.dina(n1600), .dinb(n798), .dout(n2595));
  jand g02532(.dina(n2595), .dinb(n746), .dout(n2596));
  jand g02533(.dina(n2596), .dinb(n2594), .dout(n2597));
  jand g02534(.dina(n2597), .dinb(n2589), .dout(n2598));
  jand g02535(.dina(n2598), .dinb(n2577), .dout(n2599));
  jand g02536(.dina(n2599), .dinb(n2571), .dout(n2600));
  jand g02537(.dina(n2600), .dinb(n2543), .dout(n2601));
  jnot g02538(.din(n2601), .dout(n2602));
  jand g02539(.dina(n2602), .dinb(n2497), .dout(n2603));
  jand g02540(.dina(n418), .dinb(n383), .dout(n2604));
  jand g02541(.dina(n2604), .dinb(n1204), .dout(n2605));
  jand g02542(.dina(n847), .dinb(n486), .dout(n2606));
  jand g02543(.dina(n2606), .dinb(n709), .dout(n2607));
  jand g02544(.dina(n2607), .dinb(n2605), .dout(n2608));
  jand g02545(.dina(n465), .dinb(n208), .dout(n2609));
  jand g02546(.dina(n2609), .dinb(n749), .dout(n2610));
  jand g02547(.dina(n605), .dinb(n255), .dout(n2611));
  jand g02548(.dina(n715), .dinb(n612), .dout(n2612));
  jand g02549(.dina(n2612), .dinb(n2611), .dout(n2613));
  jand g02550(.dina(n2613), .dinb(n2610), .dout(n2614));
  jand g02551(.dina(n2614), .dinb(n2608), .dout(n2615));
  jand g02552(.dina(n646), .dinb(n292), .dout(n2616));
  jand g02553(.dina(n543), .dinb(n197), .dout(n2617));
  jand g02554(.dina(n2617), .dinb(n2616), .dout(n2618));
  jnot g02555(.din(n1708), .dout(n2619));
  jand g02556(.dina(n305), .dinb(n161), .dout(n2620));
  jand g02557(.dina(n2620), .dinb(n2619), .dout(n2621));
  jand g02558(.dina(n1597), .dinb(n405), .dout(n2622));
  jand g02559(.dina(n2622), .dinb(n1135), .dout(n2623));
  jand g02560(.dina(n2623), .dinb(n2621), .dout(n2624));
  jand g02561(.dina(n2624), .dinb(n2618), .dout(n2625));
  jand g02562(.dina(n414), .dinb(n284), .dout(n2626));
  jand g02563(.dina(n533), .dinb(n500), .dout(n2627));
  jand g02564(.dina(n2627), .dinb(n2626), .dout(n2628));
  jand g02565(.dina(n359), .dinb(n82), .dout(n2629));
  jand g02566(.dina(n2629), .dinb(n812), .dout(n2630));
  jand g02567(.dina(n2630), .dinb(n2628), .dout(n2631));
  jand g02568(.dina(n1278), .dinb(n960), .dout(n2632));
  jand g02569(.dina(n2632), .dinb(n1500), .dout(n2633));
  jand g02570(.dina(n2633), .dinb(n2631), .dout(n2634));
  jand g02571(.dina(n2634), .dinb(n2625), .dout(n2635));
  jand g02572(.dina(n2635), .dinb(n2615), .dout(n2636));
  jand g02573(.dina(n472), .dinb(n136), .dout(n2637));
  jand g02574(.dina(n2637), .dinb(n2636), .dout(n2638));
  jand g02575(.dina(n553), .dinb(n428), .dout(n2639));
  jand g02576(.dina(n2639), .dinb(n257), .dout(n2640));
  jand g02577(.dina(n598), .dinb(n551), .dout(n2641));
  jand g02578(.dina(n1153), .dinb(n377), .dout(n2642));
  jand g02579(.dina(n2642), .dinb(n2641), .dout(n2643));
  jand g02580(.dina(n478), .dinb(n214), .dout(n2644));
  jand g02581(.dina(n2644), .dinb(n1536), .dout(n2645));
  jand g02582(.dina(n2645), .dinb(n2643), .dout(n2646));
  jand g02583(.dina(n2646), .dinb(n2640), .dout(n2647));
  jand g02584(.dina(n965), .dinb(n843), .dout(n2648));
  jand g02585(.dina(n366), .dinb(n260), .dout(n2649));
  jand g02586(.dina(n2649), .dinb(n815), .dout(n2650));
  jand g02587(.dina(n2650), .dinb(n2648), .dout(n2651));
  jand g02588(.dina(n1247), .dinb(n833), .dout(n2652));
  jand g02589(.dina(n756), .dinb(n194), .dout(n2653));
  jand g02590(.dina(n2653), .dinb(n1057), .dout(n2654));
  jand g02591(.dina(n2654), .dinb(n2652), .dout(n2655));
  jand g02592(.dina(n2655), .dinb(n2651), .dout(n2656));
  jand g02593(.dina(n2656), .dinb(n2647), .dout(n2657));
  jand g02594(.dina(n2657), .dinb(n1903), .dout(n2658));
  jand g02595(.dina(n435), .dinb(n423), .dout(n2659));
  jand g02596(.dina(n340), .dinb(n234), .dout(n2660));
  jand g02597(.dina(n2660), .dinb(n2659), .dout(n2661));
  jand g02598(.dina(n2661), .dinb(n1787), .dout(n2662));
  jand g02599(.dina(n819), .dinb(n445), .dout(n2663));
  jand g02600(.dina(n2663), .dinb(n988), .dout(n2664));
  jand g02601(.dina(n805), .dinb(n221), .dout(n2665));
  jand g02602(.dina(n2665), .dinb(n736), .dout(n2666));
  jand g02603(.dina(n2590), .dinb(n387), .dout(n2667));
  jand g02604(.dina(n2667), .dinb(n2666), .dout(n2668));
  jand g02605(.dina(n2668), .dinb(n2664), .dout(n2669));
  jand g02606(.dina(n2669), .dinb(n2662), .dout(n2670));
  jand g02607(.dina(n1995), .dinb(n277), .dout(n2671));
  jand g02608(.dina(n1231), .dinb(n1221), .dout(n2672));
  jand g02609(.dina(n2672), .dinb(n1924), .dout(n2673));
  jand g02610(.dina(n2673), .dinb(n2671), .dout(n2674));
  jand g02611(.dina(n711), .dinb(n427), .dout(n2675));
  jand g02612(.dina(n2675), .dinb(n1409), .dout(n2676));
  jand g02613(.dina(n801), .dinb(n395), .dout(n2677));
  jand g02614(.dina(n641), .dinb(n309), .dout(n2678));
  jand g02615(.dina(n2678), .dinb(n2677), .dout(n2679));
  jand g02616(.dina(n2679), .dinb(n2676), .dout(n2680));
  jand g02617(.dina(n2680), .dinb(n2674), .dout(n2681));
  jand g02618(.dina(n770), .dinb(n329), .dout(n2682));
  jand g02619(.dina(n583), .dinb(n578), .dout(n2683));
  jand g02620(.dina(n675), .dinb(n270), .dout(n2684));
  jand g02621(.dina(n2684), .dinb(n2683), .dout(n2685));
  jand g02622(.dina(n2685), .dinb(n2682), .dout(n2686));
  jand g02623(.dina(n1546), .dinb(n1284), .dout(n2687));
  jand g02624(.dina(n2687), .dinb(n615), .dout(n2688));
  jand g02625(.dina(n2688), .dinb(n2686), .dout(n2689));
  jand g02626(.dina(n2689), .dinb(n1298), .dout(n2690));
  jand g02627(.dina(n2690), .dinb(n2681), .dout(n2691));
  jand g02628(.dina(n2691), .dinb(n2670), .dout(n2692));
  jand g02629(.dina(n2692), .dinb(n2658), .dout(n2693));
  jand g02630(.dina(n2693), .dinb(n2638), .dout(n2694));
  jnot g02631(.din(n2694), .dout(n2695));
  jand g02632(.dina(n2695), .dinb(n2602), .dout(n2696));
  jand g02633(.dina(n635), .dinb(n614), .dout(n2697));
  jand g02634(.dina(n552), .dinb(n224), .dout(n2698));
  jand g02635(.dina(n2698), .dinb(n2697), .dout(n2699));
  jand g02636(.dina(n1264), .dinb(n876), .dout(n2700));
  jand g02637(.dina(n865), .dinb(n317), .dout(n2701));
  jand g02638(.dina(n2701), .dinb(n2700), .dout(n2702));
  jand g02639(.dina(n1178), .dinb(n847), .dout(n2703));
  jand g02640(.dina(n2703), .dinb(n322), .dout(n2704));
  jand g02641(.dina(n2704), .dinb(n2702), .dout(n2705));
  jand g02642(.dina(n988), .dinb(n234), .dout(n2706));
  jand g02643(.dina(n2706), .dinb(n594), .dout(n2707));
  jand g02644(.dina(n2707), .dinb(n1128), .dout(n2708));
  jand g02645(.dina(n2708), .dinb(n2705), .dout(n2709));
  jand g02646(.dina(n2709), .dinb(n2699), .dout(n2710));
  jand g02647(.dina(n574), .dinb(n352), .dout(n2711));
  jand g02648(.dina(n2711), .dinb(n566), .dout(n2712));
  jand g02649(.dina(n751), .dinb(n465), .dout(n2713));
  jand g02650(.dina(n601), .dinb(n455), .dout(n2714));
  jand g02651(.dina(n2714), .dinb(n2713), .dout(n2715));
  jand g02652(.dina(n2715), .dinb(n2712), .dout(n2716));
  jand g02653(.dina(n372), .dinb(n276), .dout(n2717));
  jand g02654(.dina(n2717), .dinb(n305), .dout(n2718));
  jand g02655(.dina(n979), .dinb(n414), .dout(n2719));
  jand g02656(.dina(n2719), .dinb(n443), .dout(n2720));
  jand g02657(.dina(n2720), .dinb(n2718), .dout(n2721));
  jand g02658(.dina(n377), .dinb(n249), .dout(n2722));
  jand g02659(.dina(n508), .dinb(n309), .dout(n2723));
  jand g02660(.dina(n2723), .dinb(n2722), .dout(n2724));
  jand g02661(.dina(n2724), .dinb(n2513), .dout(n2725));
  jand g02662(.dina(n2725), .dinb(n2721), .dout(n2726));
  jand g02663(.dina(n2726), .dinb(n2123), .dout(n2727));
  jand g02664(.dina(n2727), .dinb(n2716), .dout(n2728));
  jand g02665(.dina(n2728), .dinb(n2710), .dout(n2729));
  jand g02666(.dina(n2207), .dinb(n1921), .dout(n2730));
  jand g02667(.dina(n2730), .dinb(n2729), .dout(n2731));
  jnot g02668(.din(n2731), .dout(n2732));
  jand g02669(.dina(n2732), .dinb(n2695), .dout(n2733));
  jnot g02670(.din(n2733), .dout(n2734));
  jand g02671(.dina(n1073), .dinb(n360), .dout(n2735));
  jand g02672(.dina(n993), .dinb(n756), .dout(n2736));
  jand g02673(.dina(n2736), .dinb(n165), .dout(n2737));
  jand g02674(.dina(n2737), .dinb(n1306), .dout(n2738));
  jand g02675(.dina(n770), .dinb(n205), .dout(n2739));
  jand g02676(.dina(n516), .dinb(n130), .dout(n2740));
  jand g02677(.dina(n2740), .dinb(n2739), .dout(n2741));
  jand g02678(.dina(n965), .dinb(n432), .dout(n2742));
  jand g02679(.dina(n2742), .dinb(n1847), .dout(n2743));
  jand g02680(.dina(n2378), .dinb(n239), .dout(n2744));
  jand g02681(.dina(n2744), .dinb(n2743), .dout(n2745));
  jand g02682(.dina(n2745), .dinb(n2741), .dout(n2746));
  jand g02683(.dina(n2746), .dinb(n2738), .dout(n2747));
  jand g02684(.dina(n907), .dinb(n819), .dout(n2748));
  jand g02685(.dina(n2748), .dinb(n243), .dout(n2749));
  jand g02686(.dina(n739), .dinb(n317), .dout(n2750));
  jand g02687(.dina(n2750), .dinb(n1641), .dout(n2751));
  jand g02688(.dina(n2751), .dinb(n991), .dout(n2752));
  jand g02689(.dina(n2752), .dinb(n2749), .dout(n2753));
  jand g02690(.dina(n1889), .dinb(n1487), .dout(n2754));
  jand g02691(.dina(n2754), .dinb(n1934), .dout(n2755));
  jand g02692(.dina(n1178), .dinb(n1014), .dout(n2756));
  jand g02693(.dina(n435), .dinb(n113), .dout(n2757));
  jand g02694(.dina(n2757), .dinb(n2756), .dout(n2758));
  jand g02695(.dina(n882), .dinb(n450), .dout(n2759));
  jand g02696(.dina(n470), .dinb(n217), .dout(n2760));
  jand g02697(.dina(n2760), .dinb(n2759), .dout(n2761));
  jand g02698(.dina(n2761), .dinb(n2758), .dout(n2762));
  jand g02699(.dina(n2762), .dinb(n2755), .dout(n2763));
  jand g02700(.dina(n2763), .dinb(n2753), .dout(n2764));
  jand g02701(.dina(n2764), .dinb(n2747), .dout(n2765));
  jand g02702(.dina(n427), .dinb(n202), .dout(n2766));
  jand g02703(.dina(n2766), .dinb(n1727), .dout(n2767));
  jand g02704(.dina(n2767), .dinb(n1787), .dout(n2768));
  jand g02705(.dina(n703), .dinb(n414), .dout(n2769));
  jand g02706(.dina(n2769), .dinb(n1507), .dout(n2770));
  jand g02707(.dina(n721), .dinb(n103), .dout(n2771));
  jand g02708(.dina(n2771), .dinb(n396), .dout(n2772));
  jand g02709(.dina(n2772), .dinb(n2770), .dout(n2773));
  jand g02710(.dina(n2773), .dinb(n1006), .dout(n2774));
  jand g02711(.dina(n2774), .dinb(n2768), .dout(n2775));
  jand g02712(.dina(n700), .dinb(n658), .dout(n2776));
  jand g02713(.dina(n2776), .dinb(n793), .dout(n2777));
  jand g02714(.dina(n1597), .dinb(n228), .dout(n2778));
  jand g02715(.dina(n865), .dinb(n280), .dout(n2779));
  jand g02716(.dina(n708), .dinb(n441), .dout(n2780));
  jand g02717(.dina(n2780), .dinb(n2779), .dout(n2781));
  jand g02718(.dina(n2781), .dinb(n2778), .dout(n2782));
  jand g02719(.dina(n2782), .dinb(n2777), .dout(n2783));
  jand g02720(.dina(n612), .dinb(n391), .dout(n2784));
  jand g02721(.dina(n2784), .dinb(n833), .dout(n2785));
  jand g02722(.dina(n1581), .dinb(n1287), .dout(n2786));
  jand g02723(.dina(n2786), .dinb(n2785), .dout(n2787));
  jand g02724(.dina(n562), .dinb(n208), .dout(n2788));
  jand g02725(.dina(n1153), .dinb(n276), .dout(n2789));
  jand g02726(.dina(n2789), .dinb(n2788), .dout(n2790));
  jand g02727(.dina(n338), .dinb(n116), .dout(n2791));
  jor  g02728(.dina(n2791), .dinb(n491), .dout(n2792));
  jnot g02729(.din(n2792), .dout(n2793));
  jand g02730(.dina(n619), .dinb(n515), .dout(n2794));
  jand g02731(.dina(n2794), .dinb(n2793), .dout(n2795));
  jand g02732(.dina(n2795), .dinb(n2790), .dout(n2796));
  jand g02733(.dina(n2796), .dinb(n2787), .dout(n2797));
  jand g02734(.dina(n1160), .dinb(n354), .dout(n2798));
  jand g02735(.dina(n2798), .dinb(n2150), .dout(n2799));
  jand g02736(.dina(n1009), .dinb(n870), .dout(n2800));
  jand g02737(.dina(n2800), .dinb(n1829), .dout(n2801));
  jand g02738(.dina(n2801), .dinb(n2799), .dout(n2802));
  jand g02739(.dina(n2802), .dinb(n2797), .dout(n2803));
  jand g02740(.dina(n2803), .dinb(n2783), .dout(n2804));
  jand g02741(.dina(n2804), .dinb(n2775), .dout(n2805));
  jand g02742(.dina(n2805), .dinb(n2765), .dout(n2806));
  jand g02743(.dina(n2806), .dinb(n2735), .dout(n2807));
  jnot g02744(.din(n2807), .dout(n2808));
  jand g02745(.dina(n2808), .dinb(n2732), .dout(n2809));
  jnot g02746(.din(n2809), .dout(n2810));
  jand g02747(.dina(n1761), .dinb(n970), .dout(n2811));
  jand g02748(.dina(n988), .dinb(n441), .dout(n2812));
  jand g02749(.dina(n2812), .dinb(n1422), .dout(n2813));
  jand g02750(.dina(n2813), .dinb(n2811), .dout(n2814));
  jand g02751(.dina(n1615), .dinb(n311), .dout(n2815));
  jand g02752(.dina(n2815), .dinb(n392), .dout(n2816));
  jand g02753(.dina(n578), .dinb(n343), .dout(n2817));
  jand g02754(.dina(n1047), .dinb(n146), .dout(n2818));
  jand g02755(.dina(n2818), .dinb(n2817), .dout(n2819));
  jand g02756(.dina(n2819), .dinb(n2816), .dout(n2820));
  jand g02757(.dina(n2820), .dinb(n2718), .dout(n2821));
  jand g02758(.dina(n2821), .dinb(n2814), .dout(n2822));
  jand g02759(.dina(n224), .dinb(n120), .dout(n2823));
  jand g02760(.dina(n500), .dinb(n255), .dout(n2824));
  jand g02761(.dina(n2824), .dinb(n2823), .dout(n2825));
  jand g02762(.dina(n749), .dinb(n619), .dout(n2826));
  jand g02763(.dina(n517), .dinb(n329), .dout(n2827));
  jand g02764(.dina(n2827), .dinb(n2826), .dout(n2828));
  jand g02765(.dina(n562), .dinb(n262), .dout(n2829));
  jand g02766(.dina(n2829), .dinb(n2648), .dout(n2830));
  jand g02767(.dina(n2830), .dinb(n2828), .dout(n2831));
  jand g02768(.dina(n2831), .dinb(n2825), .dout(n2832));
  jand g02769(.dina(n1167), .dinb(n927), .dout(n2833));
  jand g02770(.dina(n882), .dinb(n1031), .dout(n2834));
  jand g02771(.dina(n2834), .dinb(n246), .dout(n2835));
  jand g02772(.dina(n2835), .dinb(n2833), .dout(n2836));
  jand g02773(.dina(n2347), .dinb(n802), .dout(n2837));
  jand g02774(.dina(n2837), .dinb(n2769), .dout(n2838));
  jand g02775(.dina(n2838), .dinb(n2836), .dout(n2839));
  jnot g02776(.din(n1376), .dout(n2840));
  jand g02777(.dina(n2840), .dinb(n756), .dout(n2841));
  jand g02778(.dina(n2841), .dinb(n1881), .dout(n2842));
  jand g02779(.dina(n2842), .dinb(n1022), .dout(n2843));
  jand g02780(.dina(n2843), .dinb(n2839), .dout(n2844));
  jand g02781(.dina(n2844), .dinb(n2832), .dout(n2845));
  jand g02782(.dina(n2845), .dinb(n2822), .dout(n2846));
  jand g02783(.dina(n950), .dinb(n325), .dout(n2847));
  jand g02784(.dina(n826), .dinb(n609), .dout(n2848));
  jand g02785(.dina(n2848), .dinb(n2847), .dout(n2849));
  jand g02786(.dina(n483), .dinb(n143), .dout(n2850));
  jand g02787(.dina(n2850), .dinb(n909), .dout(n2851));
  jand g02788(.dina(n2851), .dinb(n1511), .dout(n2852));
  jand g02789(.dina(n2852), .dinb(n2849), .dout(n2853));
  jand g02790(.dina(n2183), .dinb(n1085), .dout(n2854));
  jand g02791(.dina(n1119), .dinb(n198), .dout(n2855));
  jand g02792(.dina(n2855), .dinb(n2854), .dout(n2856));
  jand g02793(.dina(n715), .dinb(n553), .dout(n2857));
  jand g02794(.dina(n2857), .dinb(n1299), .dout(n2858));
  jand g02795(.dina(n257), .dinb(n217), .dout(n2859));
  jand g02796(.dina(n2859), .dinb(n2499), .dout(n2860));
  jand g02797(.dina(n2860), .dinb(n2858), .dout(n2861));
  jand g02798(.dina(n2861), .dinb(n2856), .dout(n2862));
  jand g02799(.dina(n2862), .dinb(n2524), .dout(n2863));
  jand g02800(.dina(n2863), .dinb(n2853), .dout(n2864));
  jand g02801(.dina(n2864), .dinb(n2465), .dout(n2865));
  jand g02802(.dina(n2865), .dinb(n2846), .dout(n2866));
  jnot g02803(.din(n2866), .dout(n2867));
  jand g02804(.dina(n2867), .dinb(n2808), .dout(n2868));
  jnot g02805(.din(n2868), .dout(n2869));
  jand g02806(.dina(n352), .dinb(n260), .dout(n2870));
  jand g02807(.dina(n2870), .dinb(n534), .dout(n2871));
  jand g02808(.dina(n385), .dinb(n288), .dout(n2872));
  jand g02809(.dina(n2872), .dinb(n1216), .dout(n2873));
  jand g02810(.dina(n2873), .dinb(n2871), .dout(n2874));
  jand g02811(.dina(n325), .dinb(n271), .dout(n2875));
  jand g02812(.dina(n756), .dinb(n509), .dout(n2876));
  jand g02813(.dina(n2876), .dinb(n1597), .dout(n2877));
  jand g02814(.dina(n317), .dinb(n202), .dout(n2878));
  jand g02815(.dina(n2878), .dinb(n1150), .dout(n2879));
  jand g02816(.dina(n2879), .dinb(n2877), .dout(n2880));
  jand g02817(.dina(n2880), .dinb(n2875), .dout(n2881));
  jand g02818(.dina(n2881), .dinb(n2874), .dout(n2882));
  jand g02819(.dina(n907), .dinb(n703), .dout(n2883));
  jand g02820(.dina(n1221), .dinb(n715), .dout(n2884));
  jand g02821(.dina(n2884), .dinb(n2883), .dout(n2885));
  jand g02822(.dina(n1470), .dinb(n451), .dout(n2886));
  jand g02823(.dina(n1268), .dinb(n337), .dout(n2887));
  jand g02824(.dina(n184), .dinb(n165), .dout(n2888));
  jand g02825(.dina(n2888), .dinb(n2887), .dout(n2889));
  jand g02826(.dina(n2889), .dinb(n2886), .dout(n2890));
  jand g02827(.dina(n2890), .dinb(n2885), .dout(n2891));
  jand g02828(.dina(n876), .dinb(n527), .dout(n2892));
  jand g02829(.dina(n392), .dinb(n386), .dout(n2893));
  jand g02830(.dina(n2893), .dinb(n2892), .dout(n2894));
  jand g02831(.dina(n2894), .dinb(n1644), .dout(n2895));
  jand g02832(.dina(n2512), .dinb(n501), .dout(n2896));
  jand g02833(.dina(n815), .dinb(n465), .dout(n2897));
  jand g02834(.dina(n2897), .dinb(n927), .dout(n2898));
  jand g02835(.dina(n2898), .dinb(n2896), .dout(n2899));
  jand g02836(.dina(n2899), .dinb(n2166), .dout(n2900));
  jand g02837(.dina(n2900), .dinb(n2895), .dout(n2901));
  jand g02838(.dina(n2901), .dinb(n2891), .dout(n2902));
  jand g02839(.dina(n2902), .dinb(n2882), .dout(n2903));
  jand g02840(.dina(n658), .dinb(n286), .dout(n2904));
  jand g02841(.dina(n2904), .dinb(n2053), .dout(n2905));
  jand g02842(.dina(n1085), .dinb(n979), .dout(n2906));
  jand g02843(.dina(n2906), .dinb(n2488), .dout(n2907));
  jand g02844(.dina(n2907), .dinb(n2905), .dout(n2908));
  jand g02845(.dina(n1034), .dinb(n635), .dout(n2909));
  jand g02846(.dina(n1409), .dinb(n874), .dout(n2910));
  jand g02847(.dina(n2910), .dinb(n2909), .dout(n2911));
  jand g02848(.dina(n993), .dinb(n505), .dout(n2912));
  jand g02849(.dina(n2912), .dinb(n2362), .dout(n2913));
  jand g02850(.dina(n2913), .dinb(n2911), .dout(n2914));
  jand g02851(.dina(n329), .dinb(n309), .dout(n2915));
  jand g02852(.dina(n2915), .dinb(n1165), .dout(n2916));
  jand g02853(.dina(n2916), .dinb(n1899), .dout(n2917));
  jand g02854(.dina(n1383), .dinb(n455), .dout(n2918));
  jand g02855(.dina(n2014), .dinb(n1100), .dout(n2919));
  jand g02856(.dina(n2919), .dinb(n2918), .dout(n2920));
  jand g02857(.dina(n2920), .dinb(n2917), .dout(n2921));
  jand g02858(.dina(n2921), .dinb(n2914), .dout(n2922));
  jand g02859(.dina(n2922), .dinb(n2908), .dout(n2923));
  jand g02860(.dina(n2264), .dinb(n678), .dout(n2924));
  jand g02861(.dina(n2150), .dinb(n2130), .dout(n2925));
  jand g02862(.dina(n2925), .dinb(n2924), .dout(n2926));
  jand g02863(.dina(n2015), .dinb(n833), .dout(n2927));
  jand g02864(.dina(n1048), .dinb(n791), .dout(n2928));
  jand g02865(.dina(n2928), .dinb(n2927), .dout(n2929));
  jand g02866(.dina(n414), .dinb(n154), .dout(n2930));
  jand g02867(.dina(n2930), .dinb(n622), .dout(n2931));
  jand g02868(.dina(n2931), .dinb(n2664), .dout(n2932));
  jand g02869(.dina(n2932), .dinb(n2929), .dout(n2933));
  jand g02870(.dina(n2933), .dinb(n2926), .dout(n2934));
  jand g02871(.dina(n865), .dinb(n511), .dout(n2935));
  jand g02872(.dina(n2935), .dinb(n93), .dout(n2936));
  jand g02873(.dina(n2936), .dinb(n1204), .dout(n2937));
  jand g02874(.dina(n605), .dinb(n149), .dout(n2938));
  jand g02875(.dina(n2938), .dinb(n694), .dout(n2939));
  jand g02876(.dina(n395), .dinb(n157), .dout(n2940));
  jand g02877(.dina(n346), .dinb(n249), .dout(n2941));
  jand g02878(.dina(n2941), .dinb(n2940), .dout(n2942));
  jand g02879(.dina(n2942), .dinb(n2939), .dout(n2943));
  jand g02880(.dina(n2943), .dinb(n2937), .dout(n2944));
  jand g02881(.dina(n529), .dinb(n243), .dout(n2945));
  jand g02882(.dina(n2945), .dinb(n788), .dout(n2946));
  jand g02883(.dina(n1675), .dinb(n174), .dout(n2947));
  jand g02884(.dina(n2947), .dinb(n1822), .dout(n2948));
  jand g02885(.dina(n2948), .dinb(n2946), .dout(n2949));
  jand g02886(.dina(n2949), .dinb(n2944), .dout(n2950));
  jand g02887(.dina(n2950), .dinb(n2934), .dout(n2951));
  jand g02888(.dina(n2951), .dinb(n2923), .dout(n2952));
  jand g02889(.dina(n2952), .dinb(n2903), .dout(n2953));
  jnot g02890(.din(n2953), .dout(n2954));
  jand g02891(.dina(n2954), .dinb(n2867), .dout(n2955));
  jnot g02892(.din(n2955), .dout(n2956));
  jand g02893(.dina(n788), .dinb(n659), .dout(n2957));
  jand g02894(.dina(n853), .dinb(n409), .dout(n2958));
  jand g02895(.dina(n2958), .dinb(n108), .dout(n2959));
  jand g02896(.dina(n2959), .dinb(n2957), .dout(n2960));
  jand g02897(.dina(n2960), .dinb(n2279), .dout(n2961));
  jand g02898(.dina(n703), .dinb(n405), .dout(n2962));
  jnot g02899(.din(n1372), .dout(n2963));
  jand g02900(.dina(n675), .dinb(n424), .dout(n2964));
  jand g02901(.dina(n2964), .dinb(n2963), .dout(n2965));
  jand g02902(.dina(n2965), .dinb(n2962), .dout(n2966));
  jand g02903(.dina(n2966), .dinb(n2705), .dout(n2967));
  jand g02904(.dina(n2967), .dinb(n2182), .dout(n2968));
  jand g02905(.dina(n2968), .dinb(n2961), .dout(n2969));
  jand g02906(.dina(n501), .dinb(n221), .dout(n2970));
  jand g02907(.dina(n2970), .dinb(n596), .dout(n2971));
  jand g02908(.dina(n1633), .dinb(n1576), .dout(n2972));
  jand g02909(.dina(n2972), .dinb(n2971), .dout(n2973));
  jand g02910(.dina(n2499), .dinb(n1474), .dout(n2974));
  jand g02911(.dina(n2974), .dinb(n1296), .dout(n2975));
  jand g02912(.dina(n965), .dinb(n472), .dout(n2976));
  jand g02913(.dina(n2976), .dinb(n202), .dout(n2977));
  jand g02914(.dina(n793), .dinb(n462), .dout(n2978));
  jand g02915(.dina(n2978), .dinb(n601), .dout(n2979));
  jand g02916(.dina(n2979), .dinb(n2977), .dout(n2980));
  jand g02917(.dina(n2980), .dinb(n2975), .dout(n2981));
  jand g02918(.dina(n1991), .dinb(n858), .dout(n2982));
  jand g02919(.dina(n2982), .dinb(n1627), .dout(n2983));
  jand g02920(.dina(n1067), .dinb(n557), .dout(n2984));
  jand g02921(.dina(n2984), .dinb(n2724), .dout(n2985));
  jand g02922(.dina(n2985), .dinb(n2983), .dout(n2986));
  jand g02923(.dina(n2986), .dinb(n2981), .dout(n2987));
  jand g02924(.dina(n2987), .dinb(n2973), .dout(n2988));
  jand g02925(.dina(n2988), .dinb(n2969), .dout(n2989));
  jand g02926(.dina(n2989), .dinb(n2271), .dout(n2990));
  jnot g02927(.din(n2990), .dout(n2991));
  jand g02928(.dina(n2991), .dinb(n2954), .dout(n2992));
  jnot g02929(.din(n2992), .dout(n2993));
  jand g02930(.dina(n499), .dinb(n405), .dout(n2994));
  jand g02931(.dina(n2994), .dinb(n1647), .dout(n2995));
  jand g02932(.dina(n1591), .dinb(n1088), .dout(n2996));
  jand g02933(.dina(n876), .dinb(n427), .dout(n2997));
  jand g02934(.dina(n2997), .dinb(n2870), .dout(n2998));
  jand g02935(.dina(n2998), .dinb(n2996), .dout(n2999));
  jand g02936(.dina(n2999), .dinb(n2995), .dout(n3000));
  jand g02937(.dina(n3000), .dinb(n2013), .dout(n3001));
  jand g02938(.dina(n1167), .dinb(n786), .dout(n3002));
  jand g02939(.dina(n3002), .dinb(n1280), .dout(n3003));
  jand g02940(.dina(n3003), .dinb(n1345), .dout(n3004));
  jand g02941(.dina(n404), .dinb(n340), .dout(n3005));
  jand g02942(.dina(n3005), .dinb(n478), .dout(n3006));
  jand g02943(.dina(n3006), .dinb(n2751), .dout(n3007));
  jand g02944(.dina(n3007), .dinb(n3004), .dout(n3008));
  jand g02945(.dina(n763), .dinb(n494), .dout(n3009));
  jand g02946(.dina(n3009), .dinb(n1305), .dout(n3010));
  jand g02947(.dina(n3010), .dinb(n1233), .dout(n3011));
  jnot g02948(.din(n1697), .dout(n3012));
  jand g02949(.dina(n2585), .dinb(n3012), .dout(n3013));
  jand g02950(.dina(n3013), .dinb(n3011), .dout(n3014));
  jand g02951(.dina(n377), .dinb(n174), .dout(n3015));
  jand g02952(.dina(n1314), .dinb(n529), .dout(n3016));
  jand g02953(.dina(n3016), .dinb(n3015), .dout(n3017));
  jand g02954(.dina(n2812), .dinb(n506), .dout(n3018));
  jand g02955(.dina(n3018), .dinb(n3017), .dout(n3019));
  jand g02956(.dina(n843), .dinb(n476), .dout(n3020));
  jand g02957(.dina(n423), .dinb(n208), .dout(n3021));
  jand g02958(.dina(n3021), .dinb(n3020), .dout(n3022));
  jand g02959(.dina(n749), .dinb(n770), .dout(n3023));
  jand g02960(.dina(n888), .dinb(n793), .dout(n3024));
  jand g02961(.dina(n3024), .dinb(n3023), .dout(n3025));
  jand g02962(.dina(n3025), .dinb(n3022), .dout(n3026));
  jand g02963(.dina(n3026), .dinb(n3019), .dout(n3027));
  jand g02964(.dina(n3027), .dinb(n3014), .dout(n3028));
  jand g02965(.dina(n3028), .dinb(n3008), .dout(n3029));
  jand g02966(.dina(n3029), .dinb(n3001), .dout(n3030));
  jand g02967(.dina(n913), .dinb(n407), .dout(n3031));
  jand g02968(.dina(n3031), .dinb(n647), .dout(n3032));
  jand g02969(.dina(n527), .dinb(n143), .dout(n3033));
  jand g02970(.dina(n3033), .dinb(n574), .dout(n3034));
  jand g02971(.dina(n3034), .dinb(n1997), .dout(n3035));
  jand g02972(.dina(n3035), .dinb(n3032), .dout(n3036));
  jand g02973(.dina(n1486), .dinb(n941), .dout(n3037));
  jand g02974(.dina(n3037), .dinb(n3036), .dout(n3038));
  jand g02975(.dina(n382), .dinb(n305), .dout(n3039));
  jand g02976(.dina(n3039), .dinb(n3038), .dout(n3040));
  jand g02977(.dina(n418), .dinb(n346), .dout(n3041));
  jand g02978(.dina(n3041), .dinb(n2401), .dout(n3042));
  jand g02979(.dina(n3042), .dinb(n1278), .dout(n3043));
  jand g02980(.dina(n1264), .dinb(n157), .dout(n3044));
  jand g02981(.dina(n3044), .dinb(n1039), .dout(n3045));
  jand g02982(.dina(n692), .dinb(n238), .dout(n3046));
  jand g02983(.dina(n375), .dinb(n359), .dout(n3047));
  jand g02984(.dina(n3047), .dinb(n3046), .dout(n3048));
  jand g02985(.dina(n3048), .dinb(n3045), .dout(n3049));
  jand g02986(.dina(n3049), .dinb(n2957), .dout(n3050));
  jand g02987(.dina(n3050), .dinb(n3043), .dout(n3051));
  jand g02988(.dina(n1390), .dinb(n1274), .dout(n3052));
  jand g02989(.dina(n3052), .dinb(n1506), .dout(n3053));
  jand g02990(.dina(n694), .dinb(n154), .dout(n3054));
  jand g02991(.dina(n395), .dinb(n108), .dout(n3055));
  jand g02992(.dina(n3055), .dinb(n3054), .dout(n3056));
  jand g02993(.dina(n678), .dinb(n348), .dout(n3057));
  jand g02994(.dina(n3057), .dinb(n500), .dout(n3058));
  jand g02995(.dina(n3058), .dinb(n3056), .dout(n3059));
  jand g02996(.dina(n3059), .dinb(n3053), .dout(n3060));
  jand g02997(.dina(n2606), .dinb(n815), .dout(n3061));
  jand g02998(.dina(n644), .dinb(n552), .dout(n3062));
  jand g02999(.dina(n3062), .dinb(n3061), .dout(n3063));
  jand g03000(.dina(n3063), .dinb(n2163), .dout(n3064));
  jand g03001(.dina(n3064), .dinb(n3060), .dout(n3065));
  jand g03002(.dina(n959), .dinb(n675), .dout(n3066));
  jand g03003(.dina(n3066), .dinb(n354), .dout(n3067));
  jand g03004(.dina(n194), .dinb(n103), .dout(n3068));
  jand g03005(.dina(n802), .dinb(n277), .dout(n3069));
  jand g03006(.dina(n3069), .dinb(n3068), .dout(n3070));
  jand g03007(.dina(n3070), .dinb(n3067), .dout(n3071));
  jand g03008(.dina(n371), .dinb(n331), .dout(n3072));
  jand g03009(.dina(n3072), .dinb(n280), .dout(n3073));
  jand g03010(.dina(n483), .dinb(n224), .dout(n3074));
  jand g03011(.dina(n461), .dinb(n302), .dout(n3075));
  jand g03012(.dina(n3075), .dinb(n3074), .dout(n3076));
  jand g03013(.dina(n622), .dinb(n543), .dout(n3077));
  jand g03014(.dina(n3077), .dinb(n1796), .dout(n3078));
  jand g03015(.dina(n3078), .dinb(n3076), .dout(n3079));
  jand g03016(.dina(n3079), .dinb(n3073), .dout(n3080));
  jand g03017(.dina(n3080), .dinb(n3071), .dout(n3081));
  jand g03018(.dina(n3081), .dinb(n3065), .dout(n3082));
  jand g03019(.dina(n3082), .dinb(n3051), .dout(n3083));
  jand g03020(.dina(n3083), .dinb(n3040), .dout(n3084));
  jand g03021(.dina(n3084), .dinb(n3030), .dout(n3085));
  jnot g03022(.din(n3085), .dout(n3086));
  jand g03023(.dina(n3086), .dinb(n2991), .dout(n3087));
  jnot g03024(.din(n3087), .dout(n3088));
  jand g03025(.dina(n1412), .dinb(n923), .dout(n3089));
  jand g03026(.dina(n2468), .dinb(n764), .dout(n3090));
  jand g03027(.dina(n3090), .dinb(n3089), .dout(n3091));
  jand g03028(.dina(n607), .dinb(n494), .dout(n3092));
  jand g03029(.dina(n3092), .dinb(n557), .dout(n3093));
  jand g03030(.dina(n711), .dinb(n324), .dout(n3094));
  jand g03031(.dina(n988), .dinb(n435), .dout(n3095));
  jand g03032(.dina(n3095), .dinb(n3094), .dout(n3096));
  jand g03033(.dina(n1615), .dinb(n424), .dout(n3097));
  jand g03034(.dina(n1144), .dinb(n979), .dout(n3098));
  jand g03035(.dina(n3098), .dinb(n3097), .dout(n3099));
  jand g03036(.dina(n3099), .dinb(n3096), .dout(n3100));
  jand g03037(.dina(n3100), .dinb(n3093), .dout(n3101));
  jand g03038(.dina(n3101), .dinb(n3091), .dout(n3102));
  jand g03039(.dina(n1184), .dinb(n853), .dout(n3103));
  jand g03040(.dina(n3103), .dinb(n1268), .dout(n3104));
  jand g03041(.dina(n578), .dinb(n224), .dout(n3105));
  jand g03042(.dina(n357), .dinb(n103), .dout(n3106));
  jand g03043(.dina(n3106), .dinb(n3105), .dout(n3107));
  jand g03044(.dina(n1014), .dinb(n331), .dout(n3108));
  jand g03045(.dina(n3108), .dinb(n442), .dout(n3109));
  jand g03046(.dina(n3109), .dinb(n3107), .dout(n3110));
  jand g03047(.dina(n3110), .dinb(n3104), .dout(n3111));
  jand g03048(.dina(n1761), .dinb(n709), .dout(n3112));
  jand g03049(.dina(n2130), .dinb(n1912), .dout(n3113));
  jand g03050(.dina(n3113), .dinb(n3112), .dout(n3114));
  jand g03051(.dina(n443), .dinb(n432), .dout(n3115));
  jand g03052(.dina(n3115), .dinb(n2629), .dout(n3116));
  jand g03053(.dina(n715), .dinb(n330), .dout(n3117));
  jand g03054(.dina(n3117), .dinb(n771), .dout(n3118));
  jand g03055(.dina(n3118), .dinb(n3116), .dout(n3119));
  jand g03056(.dina(n586), .dinb(n194), .dout(n3120));
  jand g03057(.dina(n692), .dinb(n633), .dout(n3121));
  jand g03058(.dina(n3121), .dinb(n3120), .dout(n3122));
  jand g03059(.dina(n3122), .dinb(n1427), .dout(n3123));
  jand g03060(.dina(n3123), .dinb(n3119), .dout(n3124));
  jand g03061(.dina(n3124), .dinb(n3114), .dout(n3125));
  jand g03062(.dina(n3125), .dinb(n3111), .dout(n3126));
  jand g03063(.dina(n3126), .dinb(n3102), .dout(n3127));
  jand g03064(.dina(n2548), .dinb(n483), .dout(n3128));
  jand g03065(.dina(n1314), .dinb(n375), .dout(n3129));
  jand g03066(.dina(n2793), .dinb(n2087), .dout(n3130));
  jand g03067(.dina(n3130), .dinb(n3129), .dout(n3131));
  jand g03068(.dina(n3131), .dinb(n3128), .dout(n3132));
  jand g03069(.dina(n805), .dinb(n288), .dout(n3133));
  jand g03070(.dina(n3133), .dinb(n700), .dout(n3134));
  jand g03071(.dina(n635), .dinb(n605), .dout(n3135));
  jand g03072(.dina(n3135), .dinb(n154), .dout(n3136));
  jand g03073(.dina(n1066), .dinb(n177), .dout(n3137));
  jand g03074(.dina(n476), .dinb(n343), .dout(n3138));
  jand g03075(.dina(n3138), .dinb(n3137), .dout(n3139));
  jand g03076(.dina(n3139), .dinb(n3136), .dout(n3140));
  jand g03077(.dina(n3140), .dinb(n3134), .dout(n3141));
  jand g03078(.dina(n214), .dinb(n108), .dout(n3142));
  jand g03079(.dina(n3142), .dinb(n703), .dout(n3143));
  jand g03080(.dina(n739), .dinb(n143), .dout(n3144));
  jand g03081(.dina(n413), .dinb(n205), .dout(n3145));
  jand g03082(.dina(n3145), .dinb(n3144), .dout(n3146));
  jand g03083(.dina(n3146), .dinb(n3143), .dout(n3147));
  jand g03084(.dina(n1796), .dinb(n1787), .dout(n3148));
  jand g03085(.dina(n1405), .dinb(n559), .dout(n3149));
  jand g03086(.dina(n3149), .dinb(n3148), .dout(n3150));
  jand g03087(.dina(n3150), .dinb(n3147), .dout(n3151));
  jand g03088(.dina(n3151), .dinb(n3141), .dout(n3152));
  jand g03089(.dina(n3152), .dinb(n3132), .dout(n3153));
  jand g03090(.dina(n462), .dinb(n427), .dout(n3154));
  jand g03091(.dina(n824), .dinb(n371), .dout(n3155));
  jand g03092(.dina(n3155), .dinb(n842), .dout(n3156));
  jand g03093(.dina(n3156), .dinb(n3154), .dout(n3157));
  jand g03094(.dina(n749), .dinb(n197), .dout(n3158));
  jand g03095(.dina(n3158), .dinb(n533), .dout(n3159));
  jand g03096(.dina(n286), .dinb(n221), .dout(n3160));
  jand g03097(.dina(n3160), .dinb(n2261), .dout(n3161));
  jand g03098(.dina(n3161), .dinb(n3159), .dout(n3162));
  jand g03099(.dina(n3162), .dinb(n3157), .dout(n3163));
  jand g03100(.dina(n3163), .dinb(n282), .dout(n3164));
  jand g03101(.dina(n847), .dinb(n309), .dout(n3165));
  jand g03102(.dina(n3165), .dinb(n243), .dout(n3166));
  jand g03103(.dina(n1409), .dinb(n284), .dout(n3167));
  jand g03104(.dina(n3167), .dinb(n1278), .dout(n3168));
  jand g03105(.dina(n3168), .dinb(n3166), .dout(n3169));
  jnot g03106(.din(n1686), .dout(n3170));
  jand g03107(.dina(n2977), .dinb(n3170), .dout(n3171));
  jand g03108(.dina(n3171), .dinb(n3169), .dout(n3172));
  jor  g03109(.dina(n695), .dinb(n593), .dout(n3173));
  jnot g03110(.din(n3173), .dout(n3174));
  jand g03111(.dina(n3174), .dinb(n2050), .dout(n3175));
  jand g03112(.dina(n1916), .dinb(n1048), .dout(n3176));
  jand g03113(.dina(n3176), .dinb(n1150), .dout(n3177));
  jand g03114(.dina(n3177), .dinb(n3175), .dout(n3178));
  jand g03115(.dina(n3178), .dinb(n3172), .dout(n3179));
  jand g03116(.dina(n3179), .dinb(n3164), .dout(n3180));
  jand g03117(.dina(n3180), .dinb(n3153), .dout(n3181));
  jand g03118(.dina(n3181), .dinb(n3127), .dout(n3182));
  jnot g03119(.din(n3182), .dout(n3183));
  jand g03120(.dina(n3183), .dinb(n3086), .dout(n3184));
  jnot g03121(.din(n3184), .dout(n3185));
  jand g03122(.dina(n1231), .dinb(n756), .dout(n3186));
  jand g03123(.dina(n1615), .dinb(n893), .dout(n3187));
  jand g03124(.dina(n3187), .dinb(n3186), .dout(n3188));
  jand g03125(.dina(n675), .dinb(n224), .dout(n3189));
  jand g03126(.dina(n2179), .dinb(n1246), .dout(n3190));
  jand g03127(.dina(n3190), .dinb(n3189), .dout(n3191));
  jand g03128(.dina(n3191), .dinb(n3188), .dout(n3192));
  jnot g03129(.din(n3192), .dout(n3193));
  jand g03130(.dina(n1067), .dinb(n367), .dout(n3194));
  jnot g03131(.din(n3194), .dout(n3195));
  jand g03132(.dina(n250), .dinb(n389), .dout(n3196));
  jor  g03133(.dina(n906), .dinb(n179), .dout(n3197));
  jor  g03134(.dina(n3197), .dinb(n3196), .dout(n3198));
  jor  g03135(.dina(n3198), .dinb(n3195), .dout(n3199));
  jnot g03136(.din(n385), .dout(n3200));
  jnot g03137(.din(n337), .dout(n3201));
  jor  g03138(.dina(n621), .dinb(n3201), .dout(n3202));
  jor  g03139(.dina(n3202), .dinb(n3200), .dout(n3203));
  jor  g03140(.dina(n3203), .dinb(n900), .dout(n3204));
  jor  g03141(.dina(n3204), .dinb(n3199), .dout(n3205));
  jnot g03142(.din(n2706), .dout(n3206));
  jand g03143(.dina(n222), .dinb(n116), .dout(n3207));
  jand g03144(.dina(n344), .dinb(n300), .dout(n3208));
  jor  g03145(.dina(n3208), .dinb(n3207), .dout(n3209));
  jnot g03146(.din(n435), .dout(n3210));
  jnot g03147(.din(n824), .dout(n3211));
  jor  g03148(.dina(n3211), .dinb(n3210), .dout(n3212));
  jor  g03149(.dina(n3212), .dinb(n3209), .dout(n3213));
  jor  g03150(.dina(n3213), .dinb(n3206), .dout(n3214));
  jnot g03151(.din(n260), .dout(n3215));
  jor  g03152(.dina(n2074), .dinb(n3215), .dout(n3216));
  jor  g03153(.dina(n966), .dinb(n313), .dout(n3217));
  jor  g03154(.dina(n3217), .dinb(n3216), .dout(n3218));
  jor  g03155(.dina(n852), .dinb(n448), .dout(n3219));
  jor  g03156(.dina(n3219), .dinb(n600), .dout(n3220));
  jor  g03157(.dina(n3220), .dinb(n3218), .dout(n3221));
  jor  g03158(.dina(n3221), .dinb(n3214), .dout(n3222));
  jor  g03159(.dina(n3222), .dinb(n3205), .dout(n3223));
  jor  g03160(.dina(n3223), .dinb(n3193), .dout(n3224));
  jnot g03161(.din(n3224), .dout(n3225));
  jand g03162(.dina(n1285), .dinb(n643), .dout(n3226));
  jand g03163(.dina(n3226), .dinb(n3225), .dout(n3227));
  jnot g03164(.din(n3227), .dout(n3228));
  jnot g03165(.din(n2864), .dout(n3229));
  jand g03166(.dina(n450), .dinb(n343), .dout(n3230));
  jand g03167(.dina(n842), .dinb(n478), .dout(n3231));
  jand g03168(.dina(n3231), .dinb(n3230), .dout(n3232));
  jand g03169(.dina(n646), .dinb(n434), .dout(n3233));
  jand g03170(.dina(n1346), .dinb(n749), .dout(n3234));
  jand g03171(.dina(n3234), .dinb(n3233), .dout(n3235));
  jand g03172(.dina(n1519), .dinb(n1039), .dout(n3236));
  jand g03173(.dina(n847), .dinb(n372), .dout(n3237));
  jand g03174(.dina(n3237), .dinb(n3236), .dout(n3238));
  jand g03175(.dina(n3238), .dinb(n3235), .dout(n3239));
  jand g03176(.dina(n3239), .dinb(n3232), .dout(n3240));
  jand g03177(.dina(n2292), .dinb(n1963), .dout(n3241));
  jand g03178(.dina(n2583), .dinb(n455), .dout(n3242));
  jand g03179(.dina(n3242), .dinb(n3241), .dout(n3243));
  jand g03180(.dina(n3243), .dinb(n1355), .dout(n3244));
  jand g03181(.dina(n3244), .dinb(n3240), .dout(n3245));
  jnot g03182(.din(n3245), .dout(n3246));
  jnot g03183(.din(n2944), .dout(n3247));
  jnot g03184(.din(n2421), .dout(n3248));
  jor  g03185(.dina(n3248), .dinb(n1483), .dout(n3249));
  jand g03186(.dina(n365), .dinb(n352), .dout(n3250));
  jand g03187(.dina(n3250), .dinb(n1584), .dout(n3251));
  jnot g03188(.din(n3251), .dout(n3252));
  jor  g03189(.dina(n3252), .dinb(n3249), .dout(n3253));
  jand g03190(.dina(n793), .dinb(n274), .dout(n3254));
  jand g03191(.dina(n692), .dinb(n655), .dout(n3255));
  jand g03192(.dina(n3255), .dinb(n3254), .dout(n3256));
  jnot g03193(.din(n3256), .dout(n3257));
  jor  g03194(.dina(n3257), .dinb(n1317), .dout(n3258));
  jor  g03195(.dina(n3258), .dinb(n3253), .dout(n3259));
  jand g03196(.dina(n739), .dinb(n574), .dout(n3260));
  jand g03197(.dina(n3260), .dinb(n1014), .dout(n3261));
  jand g03198(.dina(n467), .dinb(n413), .dout(n3262));
  jand g03199(.dina(n3262), .dinb(n3261), .dout(n3263));
  jnot g03200(.din(n3263), .dout(n3264));
  jnot g03201(.din(n709), .dout(n3265));
  jor  g03202(.dina(n1545), .dinb(n3265), .dout(n3266));
  jand g03203(.dina(n1104), .dinb(n983), .dout(n3267));
  jnot g03204(.din(n3267), .dout(n3268));
  jor  g03205(.dina(n3268), .dinb(n3266), .dout(n3269));
  jor  g03206(.dina(n3269), .dinb(n3264), .dout(n3270));
  jor  g03207(.dina(n3270), .dinb(n3259), .dout(n3271));
  jor  g03208(.dina(n3271), .dinb(n3247), .dout(n3272));
  jor  g03209(.dina(n3272), .dinb(n3246), .dout(n3273));
  jor  g03210(.dina(n3273), .dinb(n3229), .dout(n3274));
  jor  g03211(.dina(n3274), .dinb(n3228), .dout(n3275));
  jand g03212(.dina(n3275), .dinb(n3183), .dout(n3276));
  jnot g03213(.din(n3276), .dout(n3277));
  jand g03214(.dina(n1390), .dinb(n820), .dout(n3278));
  jand g03215(.dina(n715), .dinb(n304), .dout(n3279));
  jand g03216(.dina(n3279), .dinb(n2784), .dout(n3280));
  jand g03217(.dina(n3280), .dinb(n3278), .dout(n3281));
  jand g03218(.dina(n503), .dinb(n470), .dout(n3282));
  jand g03219(.dina(n865), .dinb(n359), .dout(n3283));
  jand g03220(.dina(n3283), .dinb(n3282), .dout(n3284));
  jand g03221(.dina(n1217), .dinb(n1154), .dout(n3285));
  jand g03222(.dina(n3285), .dinb(n3284), .dout(n3286));
  jand g03223(.dina(n1641), .dinb(n860), .dout(n3287));
  jand g03224(.dina(n965), .dinb(n284), .dout(n3288));
  jand g03225(.dina(n3288), .dinb(n3287), .dout(n3289));
  jand g03226(.dina(n1787), .dinb(n554), .dout(n3290));
  jand g03227(.dina(n3290), .dinb(n3289), .dout(n3291));
  jand g03228(.dina(n3291), .dinb(n3286), .dout(n3292));
  jand g03229(.dina(n3292), .dinb(n3281), .dout(n3293));
  jnot g03230(.din(n3293), .dout(n3294));
  jand g03231(.dina(n979), .dinb(n413), .dout(n3295));
  jand g03232(.dina(n3295), .dinb(n462), .dout(n3296));
  jand g03233(.dina(n609), .dinb(n221), .dout(n3297));
  jand g03234(.dina(n3297), .dinb(n3031), .dout(n3298));
  jand g03235(.dina(n3298), .dinb(n3296), .dout(n3299));
  jnot g03236(.din(n3299), .dout(n3300));
  jnot g03237(.din(n245), .dout(n3301));
  jor  g03238(.dina(n1313), .dinb(n702), .dout(n3302));
  jor  g03239(.dina(n3302), .dinb(n3301), .dout(n3303));
  jor  g03240(.dina(n776), .dinb(n546), .dout(n3304));
  jor  g03241(.dina(n3304), .dinb(n3303), .dout(n3305));
  jand g03242(.dina(n272), .dinb(n389), .dout(n3306));
  jor  g03243(.dina(n2791), .dinb(n3306), .dout(n3307));
  jor  g03244(.dina(n1397), .dinb(n792), .dout(n3308));
  jor  g03245(.dina(n3308), .dinb(n3307), .dout(n3309));
  jor  g03246(.dina(n3309), .dinb(n3305), .dout(n3310));
  jor  g03247(.dina(n3310), .dinb(n3300), .dout(n3311));
  jand g03248(.dina(n215), .dinb(n344), .dout(n3312));
  jand g03249(.dina(n235), .dinb(n101), .dout(n3313));
  jor  g03250(.dina(n3313), .dinb(n3312), .dout(n3314));
  jand g03251(.dina(n172), .dinb(n300), .dout(n3315));
  jor  g03252(.dina(n718), .dinb(n3315), .dout(n3316));
  jor  g03253(.dina(n3316), .dinb(n3314), .dout(n3317));
  jnot g03254(.din(n424), .dout(n3318));
  jor  g03255(.dina(n3318), .dinb(n422), .dout(n3319));
  jnot g03256(.din(n288), .dout(n3320));
  jor  g03257(.dina(n323), .dinb(n3320), .dout(n3321));
  jor  g03258(.dina(n3321), .dinb(n3319), .dout(n3322));
  jor  g03259(.dina(n3322), .dinb(n3317), .dout(n3323));
  jor  g03260(.dina(n493), .dinb(n2070), .dout(n3324));
  jor  g03261(.dina(n3324), .dinb(n1013), .dout(n3325));
  jnot g03262(.din(n276), .dout(n3326));
  jor  g03263(.dina(n477), .dinb(n3326), .dout(n3327));
  jor  g03264(.dina(n640), .dinb(n339), .dout(n3328));
  jor  g03265(.dina(n3328), .dinb(n3327), .dout(n3329));
  jor  g03266(.dina(n3329), .dinb(n3325), .dout(n3330));
  jor  g03267(.dina(n3330), .dinb(n3323), .dout(n3331));
  jor  g03268(.dina(n3331), .dinb(n1381), .dout(n3332));
  jor  g03269(.dina(n3332), .dinb(n3311), .dout(n3333));
  jor  g03270(.dina(n3333), .dinb(n3294), .dout(n3334));
  jand g03271(.dina(n1250), .dinb(n923), .dout(n3335));
  jand g03272(.dina(n3335), .dinb(n1281), .dout(n3336));
  jnot g03273(.din(n3336), .dout(n3337));
  jand g03274(.dina(n232), .dinb(n97), .dout(n3338));
  jor  g03275(.dina(n582), .dinb(n3338), .dout(n3339));
  jand g03276(.dina(n250), .dinb(n101), .dout(n3340));
  jand g03277(.dina(n192), .dinb(n147), .dout(n3341));
  jor  g03278(.dina(n3341), .dinb(n3340), .dout(n3342));
  jor  g03279(.dina(n3342), .dinb(n3339), .dout(n3343));
  jor  g03280(.dina(n825), .dinb(n735), .dout(n3344));
  jor  g03281(.dina(n3344), .dinb(n1056), .dout(n3345));
  jor  g03282(.dina(n3345), .dinb(n3343), .dout(n3346));
  jnot g03283(.din(n647), .dout(n3347));
  jnot g03284(.din(n700), .dout(n3348));
  jor  g03285(.dina(n3348), .dinb(n291), .dout(n3349));
  jor  g03286(.dina(n3349), .dinb(n3347), .dout(n3350));
  jor  g03287(.dina(n748), .dinb(n173), .dout(n3351));
  jor  g03288(.dina(n1177), .dinb(n201), .dout(n3352));
  jor  g03289(.dina(n3352), .dinb(n3351), .dout(n3353));
  jor  g03290(.dina(n3353), .dinb(n3350), .dout(n3354));
  jor  g03291(.dina(n3354), .dinb(n3346), .dout(n3355));
  jor  g03292(.dina(n3355), .dinb(n3337), .dout(n3356));
  jor  g03293(.dina(n3356), .dinb(n1803), .dout(n3357));
  jor  g03294(.dina(n3357), .dinb(n3224), .dout(n3358));
  jor  g03295(.dina(n3358), .dinb(n3334), .dout(n3359));
  jand g03296(.dina(n3359), .dinb(n3275), .dout(n3360));
  jnot g03297(.din(n3360), .dout(n3361));
  jnot g03298(.din(n596), .dout(n3362));
  jand g03299(.dina(n979), .dinb(n566), .dout(n3363));
  jnot g03300(.din(n3363), .dout(n3364));
  jand g03301(.dina(n215), .dinb(n200), .dout(n3365));
  jor  g03302(.dina(n677), .dinb(n3365), .dout(n3366));
  jor  g03303(.dina(n3366), .dinb(n3364), .dout(n3367));
  jor  g03304(.dina(n3367), .dinb(n3362), .dout(n3368));
  jnot g03305(.din(n3368), .dout(n3369));
  jand g03306(.dina(n278), .dinb(n272), .dout(n3370));
  jand g03307(.dina(n128), .dinb(n300), .dout(n3371));
  jor  g03308(.dina(n3371), .dinb(n3370), .dout(n3372));
  jor  g03309(.dina(n3372), .dinb(n313), .dout(n3373));
  jnot g03310(.din(n3373), .dout(n3374));
  jand g03311(.dina(n586), .dinb(n553), .dout(n3375));
  jand g03312(.dina(n309), .dinb(n230), .dout(n3376));
  jand g03313(.dina(n3376), .dinb(n3375), .dout(n3377));
  jand g03314(.dina(n3377), .dinb(n3194), .dout(n3378));
  jand g03315(.dina(n3378), .dinb(n3374), .dout(n3379));
  jand g03316(.dina(n3379), .dinb(n3369), .dout(n3380));
  jnot g03317(.din(n3380), .dout(n3381));
  jand g03318(.dina(n195), .dinb(n106), .dout(n3382));
  jor  g03319(.dina(n3382), .dinb(n528), .dout(n3383));
  jor  g03320(.dina(n1143), .dinb(n129), .dout(n3384));
  jor  g03321(.dina(n3384), .dinb(n3383), .dout(n3385));
  jnot g03322(.din(n3385), .dout(n3386));
  jand g03323(.dina(n700), .dinb(n382), .dout(n3387));
  jand g03324(.dina(n3387), .dinb(n907), .dout(n3388));
  jand g03325(.dina(n354), .dinb(n302), .dout(n3389));
  jand g03326(.dina(n3389), .dinb(n537), .dout(n3390));
  jand g03327(.dina(n3390), .dinb(n3388), .dout(n3391));
  jand g03328(.dina(n3391), .dinb(n3386), .dout(n3392));
  jnot g03329(.din(n3392), .dout(n3393));
  jand g03330(.dina(n1305), .dinb(n544), .dout(n3394));
  jand g03331(.dina(n3394), .dinb(n455), .dout(n3395));
  jnot g03332(.din(n3395), .dout(n3396));
  jand g03333(.dina(n786), .dinb(n715), .dout(n3397));
  jand g03334(.dina(n763), .dinb(n280), .dout(n3398));
  jand g03335(.dina(n3398), .dinb(n3397), .dout(n3399));
  jnot g03336(.din(n3399), .dout(n3400));
  jand g03337(.dina(n701), .dinb(n612), .dout(n3401));
  jnot g03338(.din(n3401), .dout(n3402));
  jor  g03339(.dina(n3402), .dinb(n662), .dout(n3403));
  jor  g03340(.dina(n1888), .dinb(n1133), .dout(n3404));
  jor  g03341(.dina(n3404), .dinb(n3403), .dout(n3405));
  jor  g03342(.dina(n3405), .dinb(n3400), .dout(n3406));
  jor  g03343(.dina(n3406), .dinb(n3396), .dout(n3407));
  jor  g03344(.dina(n3407), .dinb(n3393), .dout(n3408));
  jor  g03345(.dina(n3408), .dinb(n3381), .dout(n3409));
  jor  g03346(.dina(n2094), .dinb(n1722), .dout(n3410));
  jor  g03347(.dina(n3410), .dinb(n3409), .dout(n3411));
  jand g03348(.dina(n3411), .dinb(n3359), .dout(n3412));
  jnot g03349(.din(n3412), .dout(n3413));
  jnot g03350(.din(n3411), .dout(n3414));
  jand g03351(.dina(n794), .dinb(n354), .dout(n3415));
  jand g03352(.dina(n3415), .dinb(n1249), .dout(n3416));
  jand g03353(.dina(n439), .dinb(n113), .dout(n3417));
  jand g03354(.dina(n3417), .dinb(n3097), .dout(n3418));
  jand g03355(.dina(n2629), .dinb(n1934), .dout(n3419));
  jand g03356(.dina(n3419), .dinb(n3418), .dout(n3420));
  jand g03357(.dina(n876), .dinb(n435), .dout(n3421));
  jand g03358(.dina(n3421), .dinb(n882), .dout(n3422));
  jor  g03359(.dina(n702), .dinb(n504), .dout(n3423));
  jor  g03360(.dina(n964), .dinb(n381), .dout(n3424));
  jor  g03361(.dina(n3424), .dinb(n3423), .dout(n3425));
  jnot g03362(.din(n3425), .dout(n3426));
  jand g03363(.dina(n3426), .dinb(n3422), .dout(n3427));
  jand g03364(.dina(n3427), .dinb(n3420), .dout(n3428));
  jand g03365(.dina(n3428), .dinb(n3416), .dout(n3429));
  jand g03366(.dina(n909), .dinb(n566), .dout(n3430));
  jand g03367(.dina(n3430), .dinb(n716), .dout(n3431));
  jand g03368(.dina(n343), .dinb(n260), .dout(n3432));
  jand g03369(.dina(n3432), .dinb(n557), .dout(n3433));
  jand g03370(.dina(n924), .dinb(n197), .dout(n3434));
  jand g03371(.dina(n3434), .dinb(n1216), .dout(n3435));
  jand g03372(.dina(n3435), .dinb(n3433), .dout(n3436));
  jand g03373(.dina(n3436), .dinb(n3431), .dout(n3437));
  jand g03374(.dina(n842), .dinb(n417), .dout(n3438));
  jand g03375(.dina(n3438), .dinb(n202), .dout(n3439));
  jand g03376(.dina(n325), .dinb(n311), .dout(n3440));
  jand g03377(.dina(n607), .dinb(n562), .dout(n3441));
  jand g03378(.dina(n3441), .dinb(n3440), .dout(n3442));
  jand g03379(.dina(n3442), .dinb(n2640), .dout(n3443));
  jand g03380(.dina(n3443), .dinb(n3439), .dout(n3444));
  jand g03381(.dina(n527), .dinb(n120), .dout(n3445));
  jand g03382(.dina(n2420), .dinb(n579), .dout(n3446));
  jand g03383(.dina(n3446), .dinb(n3445), .dout(n3447));
  jand g03384(.dina(n843), .dinb(n450), .dout(n3448));
  jand g03385(.dina(n3448), .dinb(n983), .dout(n3449));
  jand g03386(.dina(n959), .dinb(n165), .dout(n3450));
  jand g03387(.dina(n3450), .dinb(n1591), .dout(n3451));
  jand g03388(.dina(n3451), .dinb(n3449), .dout(n3452));
  jand g03389(.dina(n3452), .dinb(n3447), .dout(n3453));
  jand g03390(.dina(n3453), .dinb(n3444), .dout(n3454));
  jand g03391(.dina(n3454), .dinb(n3437), .dout(n3455));
  jand g03392(.dina(n3455), .dinb(n3429), .dout(n3456));
  jand g03393(.dina(n517), .dinb(n190), .dout(n3457));
  jand g03394(.dina(n1221), .dinb(n392), .dout(n3458));
  jand g03395(.dina(n3458), .dinb(n3457), .dout(n3459));
  jand g03396(.dina(n2565), .dinb(n1840), .dout(n3460));
  jand g03397(.dina(n3460), .dinb(n3459), .dout(n3461));
  jand g03398(.dina(n1346), .dinb(n509), .dout(n3462));
  jand g03399(.dina(n3462), .dinb(n262), .dout(n3463));
  jand g03400(.dina(n3463), .dinb(n2446), .dout(n3464));
  jand g03401(.dina(n3464), .dinb(n3461), .dout(n3465));
  jand g03402(.dina(n1040), .dinb(n508), .dout(n3466));
  jand g03403(.dina(n3466), .dinb(n700), .dout(n3467));
  jor  g03404(.dina(n608), .dinb(n102), .dout(n3468));
  jnot g03405(.din(n3468), .dout(n3469));
  jand g03406(.dina(n3469), .dinb(n3467), .dout(n3470));
  jand g03407(.dina(n324), .dinb(n288), .dout(n3471));
  jand g03408(.dina(n2604), .dinb(n1676), .dout(n3472));
  jand g03409(.dina(n3472), .dinb(n3471), .dout(n3473));
  jand g03410(.dina(n3473), .dinb(n3470), .dout(n3474));
  jand g03411(.dina(n3474), .dinb(n3465), .dout(n3475));
  jand g03412(.dina(n3475), .dinb(n2338), .dout(n3476));
  jand g03413(.dina(n907), .dinb(n372), .dout(n3477));
  jand g03414(.dina(n3477), .dinb(n1611), .dout(n3478));
  jor  g03415(.dina(n618), .dinb(n460), .dout(n3479));
  jor  g03416(.dina(n3479), .dinb(n408), .dout(n3480));
  jnot g03417(.din(n3480), .dout(n3481));
  jor  g03418(.dina(n313), .dinb(n107), .dout(n3482));
  jnot g03419(.din(n3482), .dout(n3483));
  jand g03420(.dina(n3117), .dinb(n574), .dout(n3484));
  jand g03421(.dina(n3484), .dinb(n3483), .dout(n3485));
  jand g03422(.dina(n3485), .dinb(n3481), .dout(n3486));
  jand g03423(.dina(n3486), .dinb(n3478), .dout(n3487));
  jor  g03424(.dina(n2381), .dinb(n289), .dout(n3488));
  jnot g03425(.din(n3488), .dout(n3489));
  jand g03426(.dina(n817), .dinb(n405), .dout(n3490));
  jand g03427(.dina(n371), .dinb(n146), .dout(n3491));
  jand g03428(.dina(n3491), .dinb(n3490), .dout(n3492));
  jand g03429(.dina(n3492), .dinb(n1081), .dout(n3493));
  jand g03430(.dina(n3493), .dinb(n3489), .dout(n3494));
  jand g03431(.dina(n658), .dinb(n586), .dout(n3495));
  jand g03432(.dina(n1519), .dinb(n1268), .dout(n3496));
  jand g03433(.dina(n3496), .dinb(n3495), .dout(n3497));
  jand g03434(.dina(n802), .dinb(n693), .dout(n3498));
  jand g03435(.dina(n3498), .dinb(n3497), .dout(n3499));
  jand g03436(.dina(n1039), .dinb(n357), .dout(n3500));
  jand g03437(.dina(n476), .dinb(n336), .dout(n3501));
  jand g03438(.dina(n3501), .dinb(n3500), .dout(n3502));
  jand g03439(.dina(n270), .dinb(n255), .dout(n3503));
  jand g03440(.dina(n3503), .dinb(n214), .dout(n3504));
  jand g03441(.dina(n3504), .dinb(n3502), .dout(n3505));
  jand g03442(.dina(n3505), .dinb(n3499), .dout(n3506));
  jand g03443(.dina(n1185), .dinb(n386), .dout(n3507));
  jand g03444(.dina(n3507), .dinb(n615), .dout(n3508));
  jand g03445(.dina(n2402), .dinb(n433), .dout(n3509));
  jand g03446(.dina(n3509), .dinb(n1881), .dout(n3510));
  jand g03447(.dina(n3510), .dinb(n3508), .dout(n3511));
  jand g03448(.dina(n3511), .dinb(n3506), .dout(n3512));
  jand g03449(.dina(n3512), .dinb(n3494), .dout(n3513));
  jand g03450(.dina(n3513), .dinb(n3487), .dout(n3514));
  jand g03451(.dina(n3514), .dinb(n3476), .dout(n3515));
  jand g03452(.dina(n3515), .dinb(n3456), .dout(n3516));
  jor  g03453(.dina(n3516), .dinb(n3414), .dout(n3517));
  jxor g03454(.dina(n3516), .dinb(n3411), .dout(n3518));
  jand g03455(.dina(n993), .dinb(n427), .dout(n3519));
  jand g03456(.dina(n3519), .dinb(n893), .dout(n3520));
  jand g03457(.dina(n3520), .dinb(n2556), .dout(n3521));
  jand g03458(.dina(n3521), .dinb(n1521), .dout(n3522));
  jand g03459(.dina(n509), .dinb(n461), .dout(n3523));
  jand g03460(.dina(n3523), .dinb(n393), .dout(n3524));
  jand g03461(.dina(n563), .dinb(n559), .dout(n3525));
  jand g03462(.dina(n3525), .dinb(n3524), .dout(n3526));
  jand g03463(.dina(n876), .dinb(n472), .dout(n3527));
  jand g03464(.dina(n3527), .dinb(n1160), .dout(n3528));
  jand g03465(.dina(n3528), .dinb(n1050), .dout(n3529));
  jand g03466(.dina(n3529), .dinb(n3526), .dout(n3530));
  jand g03467(.dina(n696), .dinb(n583), .dout(n3531));
  jand g03468(.dina(n3531), .dinb(n255), .dout(n3532));
  jand g03469(.dina(n1231), .dinb(n671), .dout(n3533));
  jand g03470(.dina(n926), .dinb(n913), .dout(n3534));
  jand g03471(.dina(n3534), .dinb(n3533), .dout(n3535));
  jand g03472(.dina(n3535), .dinb(n3532), .dout(n3536));
  jand g03473(.dina(n2812), .dinb(n2423), .dout(n3537));
  jand g03474(.dina(n3537), .dinb(n833), .dout(n3538));
  jand g03475(.dina(n3538), .dinb(n3536), .dout(n3539));
  jand g03476(.dina(n3539), .dinb(n3530), .dout(n3540));
  jand g03477(.dina(n3540), .dinb(n3522), .dout(n3541));
  jand g03478(.dina(n450), .dinb(n397), .dout(n3542));
  jand g03479(.dina(n3542), .dinb(n2200), .dout(n3543));
  jand g03480(.dina(n1409), .dinb(n424), .dout(n3544));
  jand g03481(.dina(n3544), .dinb(n1492), .dout(n3545));
  jand g03482(.dina(n3363), .dinb(n1185), .dout(n3546));
  jand g03483(.dina(n3546), .dinb(n3545), .dout(n3547));
  jand g03484(.dina(n3547), .dinb(n3543), .dout(n3548));
  jand g03485(.dina(n3548), .dinb(n3263), .dout(n3549));
  jand g03486(.dina(n701), .dinb(n92), .dout(n3550));
  jand g03487(.dina(n865), .dinb(n700), .dout(n3551));
  jand g03488(.dina(n3551), .dinb(n3550), .dout(n3552));
  jand g03489(.dina(n2053), .dinb(n869), .dout(n3553));
  jand g03490(.dina(n3553), .dinb(n3552), .dout(n3554));
  jand g03491(.dina(n578), .dinb(n500), .dout(n3555));
  jand g03492(.dina(n3555), .dinb(n1711), .dout(n3556));
  jand g03493(.dina(n536), .dinb(n260), .dout(n3557));
  jand g03494(.dina(n443), .dinb(n257), .dout(n3558));
  jand g03495(.dina(n3558), .dinb(n3557), .dout(n3559));
  jand g03496(.dina(n3559), .dinb(n3556), .dout(n3560));
  jand g03497(.dina(n3560), .dinb(n3554), .dout(n3561));
  jand g03498(.dina(n2135), .dinb(n1536), .dout(n3562));
  jand g03499(.dina(n817), .dinb(n462), .dout(n3563));
  jand g03500(.dina(n3563), .dinb(n1273), .dout(n3564));
  jand g03501(.dina(n3564), .dinb(n3562), .dout(n3565));
  jand g03502(.dina(n1500), .dinb(n481), .dout(n3566));
  jand g03503(.dina(n716), .dinb(n330), .dout(n3567));
  jand g03504(.dina(n819), .dinb(n612), .dout(n3568));
  jand g03505(.dina(n3568), .dinb(n3567), .dout(n3569));
  jand g03506(.dina(n3569), .dinb(n3566), .dout(n3570));
  jand g03507(.dina(n3570), .dinb(n3565), .dout(n3571));
  jand g03508(.dina(n3571), .dinb(n3561), .dout(n3572));
  jand g03509(.dina(n3572), .dinb(n3549), .dout(n3573));
  jand g03510(.dina(n2823), .dinb(n2420), .dout(n3574));
  jand g03511(.dina(n1916), .dinb(n1585), .dout(n3575));
  jand g03512(.dina(n3575), .dinb(n3574), .dout(n3576));
  jand g03513(.dina(n1221), .dinb(n907), .dout(n3577));
  jand g03514(.dina(n3577), .dinb(n322), .dout(n3578));
  jand g03515(.dina(n658), .dinb(n202), .dout(n3579));
  jand g03516(.dina(n3579), .dinb(n239), .dout(n3580));
  jand g03517(.dina(n3580), .dinb(n3578), .dout(n3581));
  jand g03518(.dina(n3581), .dinb(n3576), .dout(n3582));
  jand g03519(.dina(n805), .dinb(n286), .dout(n3583));
  jand g03520(.dina(n3583), .dinb(n1760), .dout(n3584));
  jand g03521(.dina(n712), .dinb(n598), .dout(n3585));
  jand g03522(.dina(n3585), .dinb(n1024), .dout(n3586));
  jand g03523(.dina(n3586), .dinb(n3584), .dout(n3587));
  jand g03524(.dina(n532), .dinb(n516), .dout(n3588));
  jand g03525(.dina(n3588), .dinb(n788), .dout(n3589));
  jand g03526(.dina(n756), .dinb(n276), .dout(n3590));
  jand g03527(.dina(n3590), .dinb(n3054), .dout(n3591));
  jand g03528(.dina(n3591), .dinb(n3589), .dout(n3592));
  jand g03529(.dina(n3592), .dinb(n3587), .dout(n3593));
  jand g03530(.dina(n409), .dinb(n194), .dout(n3594));
  jand g03531(.dina(n708), .dinb(n432), .dout(n3595));
  jand g03532(.dina(n3595), .dinb(n436), .dout(n3596));
  jand g03533(.dina(n3596), .dinb(n3594), .dout(n3597));
  jand g03534(.dina(n2604), .dinb(n2538), .dout(n3598));
  jand g03535(.dina(n1284), .dinb(n870), .dout(n3599));
  jand g03536(.dina(n3599), .dinb(n3598), .dout(n3600));
  jand g03537(.dina(n3600), .dinb(n3597), .dout(n3601));
  jand g03538(.dina(n3601), .dinb(n3593), .dout(n3602));
  jand g03539(.dina(n3602), .dinb(n3582), .dout(n3603));
  jand g03540(.dina(n3603), .dinb(n3573), .dout(n3604));
  jand g03541(.dina(n3604), .dinb(n3541), .dout(n3605));
  jand g03542(.dina(n3605), .dinb(n3516), .dout(n3606));
  jand g03543(.dina(n2897), .dinb(n798), .dout(n3607));
  jand g03544(.dina(n431), .dinb(n243), .dout(n3608));
  jand g03545(.dina(n3608), .dinb(n3236), .dout(n3609));
  jand g03546(.dina(n3609), .dinb(n3607), .dout(n3610));
  jor  g03547(.dina(n308), .dinb(n216), .dout(n3611));
  jor  g03548(.dina(n3611), .dinb(n504), .dout(n3612));
  jor  g03549(.dina(n353), .dinb(n173), .dout(n3613));
  jor  g03550(.dina(n3613), .dinb(n1683), .dout(n3614));
  jor  g03551(.dina(n3614), .dinb(n3612), .dout(n3615));
  jnot g03552(.din(n3615), .dout(n3616));
  jand g03553(.dina(n3445), .dinb(n1881), .dout(n3617));
  jand g03554(.dina(n3617), .dinb(n2275), .dout(n3618));
  jand g03555(.dina(n3618), .dinb(n3616), .dout(n3619));
  jand g03556(.dina(n3619), .dinb(n3610), .dout(n3620));
  jand g03557(.dina(n435), .dinb(n284), .dout(n3621));
  jand g03558(.dina(n3621), .dinb(n612), .dout(n3622));
  jand g03559(.dina(n3622), .dinb(n1349), .dout(n3623));
  jand g03560(.dina(n3623), .dinb(n1974), .dout(n3624));
  jand g03561(.dina(n3624), .dinb(n3132), .dout(n3625));
  jand g03562(.dina(n3625), .dinb(n3620), .dout(n3626));
  jand g03563(.dina(n959), .dinb(n500), .dout(n3627));
  jand g03564(.dina(n3627), .dinb(n228), .dout(n3628));
  jand g03565(.dina(n3628), .dinb(n882), .dout(n3629));
  jor  g03566(.dina(n1166), .dinb(n229), .dout(n3630));
  jor  g03567(.dina(n3630), .dinb(n706), .dout(n3631));
  jnot g03568(.din(n3631), .dout(n3632));
  jand g03569(.dina(n3632), .dinb(n2660), .dout(n3633));
  jand g03570(.dina(n3633), .dinb(n3629), .dout(n3634));
  jand g03571(.dina(n865), .dinb(n543), .dout(n3635));
  jnot g03572(.din(n3635), .dout(n3636));
  jor  g03573(.dina(n964), .dinb(n204), .dout(n3637));
  jor  g03574(.dina(n528), .dinb(n488), .dout(n3638));
  jor  g03575(.dina(n3638), .dinb(n3637), .dout(n3639));
  jor  g03576(.dina(n3639), .dinb(n3636), .dout(n3640));
  jnot g03577(.din(n3640), .dout(n3641));
  jand g03578(.dina(n3641), .dinb(n3175), .dout(n3642));
  jand g03579(.dina(n3642), .dinb(n3634), .dout(n3643));
  jand g03580(.dina(n578), .dinb(n154), .dout(n3644));
  jand g03581(.dina(n3644), .dinb(n2468), .dout(n3645));
  jor  g03582(.dina(n718), .dinb(n556), .dout(n3646));
  jor  g03583(.dina(n3646), .dinb(n942), .dout(n3647));
  jnot g03584(.din(n3647), .dout(n3648));
  jand g03585(.dina(n3648), .dinb(n3645), .dout(n3649));
  jor  g03586(.dina(n925), .dinb(n514), .dout(n3650));
  jand g03587(.dina(n222), .dinb(n300), .dout(n3651));
  jor  g03588(.dina(n3651), .dinb(n403), .dout(n3652));
  jor  g03589(.dina(n3652), .dinb(n3650), .dout(n3653));
  jnot g03590(.din(n3653), .dout(n3654));
  jor  g03591(.dina(n480), .dinb(n193), .dout(n3655));
  jnot g03592(.din(n3655), .dout(n3656));
  jand g03593(.dina(n3656), .dinb(n425), .dout(n3657));
  jand g03594(.dina(n3657), .dinb(n3654), .dout(n3658));
  jand g03595(.dina(n3658), .dinb(n3649), .dout(n3659));
  jand g03596(.dina(n2769), .dinb(n1280), .dout(n3660));
  jor  g03597(.dina(n949), .dinb(n201), .dout(n3661));
  jnot g03598(.din(n3661), .dout(n3662));
  jand g03599(.dina(n3662), .dinb(n771), .dout(n3663));
  jand g03600(.dina(n3663), .dinb(n3660), .dout(n3664));
  jor  g03601(.dina(n493), .dinb(n303), .dout(n3665));
  jor  g03602(.dina(n3665), .dinb(n677), .dout(n3666));
  jand g03603(.dina(n159), .dinb(n203), .dout(n3667));
  jor  g03604(.dina(n3667), .dinb(n469), .dout(n3668));
  jor  g03605(.dina(n645), .dinb(n135), .dout(n3669));
  jor  g03606(.dina(n3669), .dinb(n3668), .dout(n3670));
  jor  g03607(.dina(n3670), .dinb(n3666), .dout(n3671));
  jnot g03608(.din(n3671), .dout(n3672));
  jand g03609(.dina(n3672), .dinb(n3664), .dout(n3673));
  jand g03610(.dina(n3673), .dinb(n3659), .dout(n3674));
  jand g03611(.dina(n3674), .dinb(n3643), .dout(n3675));
  jand g03612(.dina(n3675), .dinb(n3626), .dout(n3676));
  jand g03613(.dina(n3676), .dinb(n3476), .dout(n3677));
  jor  g03614(.dina(n3677), .dinb(n3606), .dout(n3678));
  jor  g03615(.dina(n3678), .dinb(n3518), .dout(n3679));
  jand g03616(.dina(n3679), .dinb(n3517), .dout(n3680));
  jxor g03617(.dina(n3414), .dinb(n3359), .dout(n3681));
  jor  g03618(.dina(n3681), .dinb(n3680), .dout(n3682));
  jand g03619(.dina(n3682), .dinb(n3413), .dout(n3683));
  jnot g03620(.din(n3359), .dout(n3684));
  jxor g03621(.dina(n3684), .dinb(n3275), .dout(n3685));
  jor  g03622(.dina(n3685), .dinb(n3683), .dout(n3686));
  jand g03623(.dina(n3686), .dinb(n3361), .dout(n3687));
  jxor g03624(.dina(n3275), .dinb(n3183), .dout(n3688));
  jnot g03625(.din(n3688), .dout(n3689));
  jor  g03626(.dina(n3689), .dinb(n3687), .dout(n3690));
  jand g03627(.dina(n3690), .dinb(n3277), .dout(n3691));
  jxor g03628(.dina(n3182), .dinb(n3085), .dout(n3692));
  jnot g03629(.din(n3692), .dout(n3693));
  jor  g03630(.dina(n3693), .dinb(n3691), .dout(n3694));
  jand g03631(.dina(n3694), .dinb(n3185), .dout(n3695));
  jxor g03632(.dina(n3085), .dinb(n2990), .dout(n3696));
  jnot g03633(.din(n3696), .dout(n3697));
  jor  g03634(.dina(n3697), .dinb(n3695), .dout(n3698));
  jand g03635(.dina(n3698), .dinb(n3088), .dout(n3699));
  jxor g03636(.dina(n2990), .dinb(n2953), .dout(n3700));
  jnot g03637(.din(n3700), .dout(n3701));
  jor  g03638(.dina(n3701), .dinb(n3699), .dout(n3702));
  jand g03639(.dina(n3702), .dinb(n2993), .dout(n3703));
  jxor g03640(.dina(n2953), .dinb(n2866), .dout(n3704));
  jnot g03641(.din(n3704), .dout(n3705));
  jor  g03642(.dina(n3705), .dinb(n3703), .dout(n3706));
  jand g03643(.dina(n3706), .dinb(n2956), .dout(n3707));
  jxor g03644(.dina(n2866), .dinb(n2807), .dout(n3708));
  jnot g03645(.din(n3708), .dout(n3709));
  jor  g03646(.dina(n3709), .dinb(n3707), .dout(n3710));
  jand g03647(.dina(n3710), .dinb(n2869), .dout(n3711));
  jxor g03648(.dina(n2807), .dinb(n2731), .dout(n3712));
  jnot g03649(.din(n3712), .dout(n3713));
  jor  g03650(.dina(n3713), .dinb(n3711), .dout(n3714));
  jand g03651(.dina(n3714), .dinb(n2810), .dout(n3715));
  jxor g03652(.dina(n2731), .dinb(n2694), .dout(n3716));
  jnot g03653(.din(n3716), .dout(n3717));
  jor  g03654(.dina(n3717), .dinb(n3715), .dout(n3718));
  jand g03655(.dina(n3718), .dinb(n2734), .dout(n3719));
  jnot g03656(.din(n3719), .dout(n3720));
  jxor g03657(.dina(n2694), .dinb(n2601), .dout(n3721));
  jand g03658(.dina(n3721), .dinb(n3720), .dout(n3722));
  jor  g03659(.dina(n3722), .dinb(n2696), .dout(n3723));
  jxor g03660(.dina(n2601), .dinb(n2496), .dout(n3724));
  jand g03661(.dina(n3724), .dinb(n3723), .dout(n3725));
  jor  g03662(.dina(n3725), .dinb(n2603), .dout(n3726));
  jxor g03663(.dina(n2496), .dinb(n2410), .dout(n3727));
  jand g03664(.dina(n3727), .dinb(n3726), .dout(n3728));
  jor  g03665(.dina(n3728), .dinb(n2498), .dout(n3729));
  jxor g03666(.dina(n2410), .dinb(n2342), .dout(n3730));
  jand g03667(.dina(n3730), .dinb(n3729), .dout(n3731));
  jor  g03668(.dina(n3731), .dinb(n2412), .dout(n3732));
  jxor g03669(.dina(n2342), .dinb(n2236), .dout(n3733));
  jand g03670(.dina(n3733), .dinb(n3732), .dout(n3734));
  jor  g03671(.dina(n3734), .dinb(n2344), .dout(n3735));
  jxor g03672(.dina(n2236), .dinb(n2127), .dout(n3736));
  jand g03673(.dina(n3736), .dinb(n3735), .dout(n3737));
  jor  g03674(.dina(n3737), .dinb(n2238), .dout(n3738));
  jxor g03675(.dina(n2127), .dinb(n2066), .dout(n3739));
  jand g03676(.dina(n3739), .dinb(n3738), .dout(n3740));
  jor  g03677(.dina(n3740), .dinb(n2129), .dout(n3741));
  jxor g03678(.dina(n2066), .dinb(n1955), .dout(n3742));
  jand g03679(.dina(n3742), .dinb(n3741), .dout(n3743));
  jor  g03680(.dina(n3743), .dinb(n2068), .dout(n3744));
  jxor g03681(.dina(n1955), .dinb(n1861), .dout(n3745));
  jand g03682(.dina(n3745), .dinb(n3744), .dout(n3746));
  jor  g03683(.dina(n3746), .dinb(n1957), .dout(n3747));
  jxor g03684(.dina(n1861), .dinb(n1775), .dout(n3748));
  jand g03685(.dina(n3748), .dinb(n3747), .dout(n3749));
  jor  g03686(.dina(n3749), .dinb(n1863), .dout(n3750));
  jxor g03687(.dina(n1775), .dinb(n1623), .dout(n3751));
  jand g03688(.dina(n3751), .dinb(n3750), .dout(n3752));
  jor  g03689(.dina(n3752), .dinb(n1777), .dout(n3753));
  jxor g03690(.dina(n1623), .dinb(n1559), .dout(n3754));
  jand g03691(.dina(n3754), .dinb(n3753), .dout(n3755));
  jor  g03692(.dina(n3755), .dinb(n1625), .dout(n3756));
  jxor g03693(.dina(n1559), .dinb(n1444), .dout(n3757));
  jand g03694(.dina(n3757), .dinb(n3756), .dout(n3758));
  jor  g03695(.dina(n3758), .dinb(n1561), .dout(n3759));
  jxor g03696(.dina(n1444), .dinb(n1342), .dout(n3760));
  jand g03697(.dina(n3760), .dinb(n3759), .dout(n3761));
  jor  g03698(.dina(n3761), .dinb(n1446), .dout(n3762));
  jxor g03699(.dina(n1342), .dinb(n1212), .dout(n3763));
  jand g03700(.dina(n3763), .dinb(n3762), .dout(n3764));
  jor  g03701(.dina(n3764), .dinb(n1344), .dout(n3765));
  jxor g03702(.dina(n1212), .dinb(n1075), .dout(n3766));
  jand g03703(.dina(n3766), .dinb(n3765), .dout(n3767));
  jor  g03704(.dina(n3767), .dinb(n1214), .dout(n3768));
  jxor g03705(.dina(n1075), .dinb(n921), .dout(n3769));
  jand g03706(.dina(n3769), .dinb(n3768), .dout(n3770));
  jor  g03707(.dina(n3770), .dinb(n1077), .dout(n3771));
  jand g03708(.dina(n1346), .dinb(n586), .dout(n3772));
  jand g03709(.dina(n3772), .dinb(n533), .dout(n3773));
  jand g03710(.dina(n3773), .dinb(n548), .dout(n3774));
  jand g03711(.dina(n3774), .dinb(n1800), .dout(n3775));
  jand g03712(.dina(n1040), .dinb(n405), .dout(n3776));
  jand g03713(.dina(n3776), .dinb(n467), .dout(n3777));
  jand g03714(.dina(n1099), .dinb(n802), .dout(n3778));
  jand g03715(.dina(n833), .dinb(n579), .dout(n3779));
  jand g03716(.dina(n3779), .dinb(n3778), .dout(n3780));
  jand g03717(.dina(n3780), .dinb(n3777), .dout(n3781));
  jand g03718(.dina(n622), .dinb(n527), .dout(n3782));
  jand g03719(.dina(n3782), .dinb(n787), .dout(n3783));
  jand g03720(.dina(n2629), .dinb(n1737), .dout(n3784));
  jand g03721(.dina(n3784), .dinb(n3783), .dout(n3785));
  jand g03722(.dina(n614), .dinb(n505), .dout(n3786));
  jand g03723(.dina(n3786), .dinb(n340), .dout(n3787));
  jand g03724(.dina(n888), .dinb(n417), .dout(n3788));
  jand g03725(.dina(n860), .dinb(n252), .dout(n3789));
  jand g03726(.dina(n3789), .dinb(n3788), .dout(n3790));
  jand g03727(.dina(n3790), .dinb(n3787), .dout(n3791));
  jand g03728(.dina(n2315), .dinb(n858), .dout(n3792));
  jand g03729(.dina(n372), .dinb(n224), .dout(n3793));
  jand g03730(.dina(n3793), .dinb(n1134), .dout(n3794));
  jand g03731(.dina(n3794), .dinb(n3792), .dout(n3795));
  jand g03732(.dina(n3795), .dinb(n3791), .dout(n3796));
  jand g03733(.dina(n3796), .dinb(n3785), .dout(n3797));
  jand g03734(.dina(n3797), .dinb(n3781), .dout(n3798));
  jand g03735(.dina(n3798), .dinb(n3775), .dout(n3799));
  jand g03736(.dina(n606), .dinb(n311), .dout(n3800));
  jand g03737(.dina(n450), .dinb(n386), .dout(n3801));
  jand g03738(.dina(n3801), .dinb(n745), .dout(n3802));
  jand g03739(.dina(n3802), .dinb(n218), .dout(n3803));
  jand g03740(.dina(n3803), .dinb(n3800), .dout(n3804));
  jand g03741(.dina(n404), .dinb(n317), .dout(n3805));
  jand g03742(.dina(n3805), .dinb(n268), .dout(n3806));
  jand g03743(.dina(n1826), .dinb(n1421), .dout(n3807));
  jand g03744(.dina(n3807), .dinb(n3806), .dout(n3808));
  jand g03745(.dina(n2664), .dinb(n1852), .dout(n3809));
  jand g03746(.dina(n3809), .dinb(n3808), .dout(n3810));
  jand g03747(.dina(n950), .dinb(n715), .dout(n3811));
  jand g03748(.dina(n3811), .dinb(n470), .dout(n3812));
  jand g03749(.dina(n3812), .dinb(n1627), .dout(n3813));
  jnot g03750(.din(n3813), .dout(n3814));
  jor  g03751(.dina(n3814), .dinb(n3305), .dout(n3815));
  jnot g03752(.din(n3815), .dout(n3816));
  jand g03753(.dina(n3816), .dinb(n3810), .dout(n3817));
  jand g03754(.dina(n3817), .dinb(n3804), .dout(n3818));
  jand g03755(.dina(n1167), .dinb(n687), .dout(n3819));
  jand g03756(.dina(n3819), .dinb(n869), .dout(n3820));
  jand g03757(.dina(n3820), .dinb(n2211), .dout(n3821));
  jand g03758(.dina(n486), .dinb(n146), .dout(n3822));
  jand g03759(.dina(n3822), .dinb(n346), .dout(n3823));
  jand g03760(.dina(n633), .dinb(n276), .dout(n3824));
  jand g03761(.dina(n3824), .dinb(n771), .dout(n3825));
  jand g03762(.dina(n2583), .dinb(n1487), .dout(n3826));
  jand g03763(.dina(n3826), .dinb(n3825), .dout(n3827));
  jand g03764(.dina(n3827), .dinb(n3823), .dout(n3828));
  jand g03765(.dina(n3828), .dinb(n3821), .dout(n3829));
  jand g03766(.dina(n708), .dinb(n413), .dout(n3830));
  jand g03767(.dina(n3830), .dinb(n382), .dout(n3831));
  jnot g03768(.din(n3665), .dout(n3832));
  jand g03769(.dina(n3832), .dinb(n806), .dout(n3833));
  jand g03770(.dina(n613), .dinb(n436), .dout(n3834));
  jand g03771(.dina(n3834), .dinb(n3833), .dout(n3835));
  jand g03772(.dina(n3835), .dinb(n3831), .dout(n3836));
  jand g03773(.dina(n2386), .dinb(n1519), .dout(n3837));
  jand g03774(.dina(n711), .dinb(n348), .dout(n3838));
  jand g03775(.dina(n924), .dinb(n143), .dout(n3839));
  jand g03776(.dina(n3839), .dinb(n3154), .dout(n3840));
  jand g03777(.dina(n3840), .dinb(n3838), .dout(n3841));
  jand g03778(.dina(n3841), .dinb(n3837), .dout(n3842));
  jand g03779(.dina(n3842), .dinb(n3836), .dout(n3843));
  jand g03780(.dina(n3843), .dinb(n3829), .dout(n3844));
  jand g03781(.dina(n3844), .dinb(n3818), .dout(n3845));
  jand g03782(.dina(n3845), .dinb(n3799), .dout(n3846));
  jxor g03783(.dina(n3846), .dinb(n921), .dout(n3847));
  jxor g03784(.dina(n3847), .dinb(n3771), .dout(n3848));
  jand g03785(.dina(n3848), .dinb(n732), .dout(n3849));
  jand g03786(.dina(\a[31] ), .dinb(\a[30] ), .dout(n3850));
  jand g03787(.dina(n3850), .dinb(n730), .dout(n3851));
  jand g03788(.dina(n3851), .dinb(n1076), .dout(n3852));
  jnot g03789(.din(n3846), .dout(n3853));
  jor  g03790(.dina(n730), .dinb(\a[31] ), .dout(n3854));
  jnot g03791(.din(n3854), .dout(n3855));
  jand g03792(.dina(n3855), .dinb(n3853), .dout(n3856));
  jxor g03793(.dina(\a[31] ), .dinb(\a[30] ), .dout(n3857));
  jand g03794(.dina(n3857), .dinb(n730), .dout(n3858));
  jand g03795(.dina(n3858), .dinb(n922), .dout(n3859));
  jor  g03796(.dina(n3859), .dinb(n3856), .dout(n3860));
  jor  g03797(.dina(n3860), .dinb(n3852), .dout(n3861));
  jor  g03798(.dina(n3861), .dinb(n3849), .dout(n3862));
  jxor g03799(.dina(n3862), .dinb(n729), .dout(n3863));
  jnot g03800(.din(n3863), .dout(n3864));
  jand g03801(.dina(n1039), .dinb(n383), .dout(n3865));
  jand g03802(.dina(n819), .dinb(n511), .dout(n3866));
  jand g03803(.dina(n3866), .dinb(n3865), .dout(n3867));
  jand g03804(.dina(n3867), .dinb(n1247), .dout(n3868));
  jand g03805(.dina(n897), .dinb(n108), .dout(n3869));
  jand g03806(.dina(n3869), .dinb(n354), .dout(n3870));
  jand g03807(.dina(n1641), .dinb(n566), .dout(n3871));
  jand g03808(.dina(n551), .dinb(n149), .dout(n3872));
  jand g03809(.dina(n3872), .dinb(n3871), .dout(n3873));
  jand g03810(.dina(n3873), .dinb(n3870), .dout(n3874));
  jand g03811(.dina(n2308), .dinb(n1169), .dout(n3875));
  jand g03812(.dina(n3875), .dinb(n3874), .dout(n3876));
  jand g03813(.dina(n3876), .dinb(n3868), .dout(n3877));
  jand g03814(.dina(n598), .dinb(n486), .dout(n3878));
  jand g03815(.dina(n1221), .dinb(n467), .dout(n3879));
  jand g03816(.dina(n3879), .dinb(n1412), .dout(n3880));
  jand g03817(.dina(n3880), .dinb(n3878), .dout(n3881));
  jand g03818(.dina(n553), .dinb(n277), .dout(n3882));
  jand g03819(.dina(n950), .dinb(n857), .dout(n3883));
  jand g03820(.dina(n3883), .dinb(n377), .dout(n3884));
  jand g03821(.dina(n3884), .dinb(n3882), .dout(n3885));
  jand g03822(.dina(n3885), .dinb(n3881), .dout(n3886));
  jand g03823(.dina(n3886), .dinb(n3494), .dout(n3887));
  jand g03824(.dina(n465), .dinb(n252), .dout(n3888));
  jand g03825(.dina(n372), .dinb(n92), .dout(n3889));
  jand g03826(.dina(n3889), .dinb(n3888), .dout(n3890));
  jand g03827(.dina(n1129), .dinb(n121), .dout(n3891));
  jand g03828(.dina(n3891), .dinb(n2997), .dout(n3892));
  jand g03829(.dina(n3892), .dinb(n3890), .dout(n3893));
  jand g03830(.dina(n622), .dinb(n462), .dout(n3894));
  jand g03831(.dina(n3894), .dinb(n557), .dout(n3895));
  jand g03832(.dina(n708), .dinb(n423), .dout(n3896));
  jand g03833(.dina(n715), .dinb(n177), .dout(n3897));
  jand g03834(.dina(n3897), .dinb(n647), .dout(n3898));
  jand g03835(.dina(n3898), .dinb(n3896), .dout(n3899));
  jand g03836(.dina(n3899), .dinb(n3895), .dout(n3900));
  jand g03837(.dina(n3900), .dinb(n3893), .dout(n3901));
  jand g03838(.dina(n3901), .dinb(n3887), .dout(n3902));
  jand g03839(.dina(n3902), .dinb(n3877), .dout(n3903));
  jand g03840(.dina(n470), .dinb(n357), .dout(n3904));
  jand g03841(.dina(n3904), .dinb(n2292), .dout(n3905));
  jand g03842(.dina(n689), .dinb(n417), .dout(n3906));
  jand g03843(.dina(n609), .dinb(n450), .dout(n3907));
  jand g03844(.dina(n3907), .dinb(n3906), .dout(n3908));
  jand g03845(.dina(n3908), .dinb(n3194), .dout(n3909));
  jand g03846(.dina(n3909), .dinb(n3905), .dout(n3910));
  jand g03847(.dina(n434), .dinb(n230), .dout(n3911));
  jand g03848(.dina(n959), .dinb(n217), .dout(n3912));
  jand g03849(.dina(n3912), .dinb(n770), .dout(n3913));
  jand g03850(.dina(n3913), .dinb(n3911), .dout(n3914));
  jand g03851(.dina(n337), .dinb(n197), .dout(n3915));
  jand g03852(.dina(n3915), .dinb(n2784), .dout(n3916));
  jand g03853(.dina(n2301), .dinb(n225), .dout(n3917));
  jand g03854(.dina(n3917), .dinb(n3916), .dout(n3918));
  jand g03855(.dina(n3918), .dinb(n3914), .dout(n3919));
  jand g03856(.dina(n3919), .dinb(n3910), .dout(n3920));
  jand g03857(.dina(n492), .dinb(n375), .dout(n3921));
  jand g03858(.dina(n3921), .dinb(n165), .dout(n3922));
  jand g03859(.dina(n1409), .dinb(n435), .dout(n3923));
  jand g03860(.dina(n3923), .dinb(n2776), .dout(n3924));
  jand g03861(.dina(n3924), .dinb(n1142), .dout(n3925));
  jand g03862(.dina(n3925), .dinb(n3922), .dout(n3926));
  jand g03863(.dina(n3926), .dinb(n2205), .dout(n3927));
  jand g03864(.dina(n3927), .dinb(n3920), .dout(n3928));
  jand g03865(.dina(n3928), .dinb(n3903), .dout(n3929));
  jnot g03866(.din(n3929), .dout(n3930));
  jand g03867(.dina(n1167), .dinb(n557), .dout(n3931));
  jand g03868(.dina(n3931), .dinb(n180), .dout(n3932));
  jand g03869(.dina(n431), .dinb(n404), .dout(n3933));
  jand g03870(.dina(n3933), .dinb(n284), .dout(n3934));
  jand g03871(.dina(n3934), .dinb(n3932), .dout(n3935));
  jand g03872(.dina(n612), .dinb(n407), .dout(n3936));
  jand g03873(.dina(n228), .dinb(n217), .dout(n3937));
  jand g03874(.dina(n3937), .dinb(n3936), .dout(n3938));
  jand g03875(.dina(n3938), .dinb(n342), .dout(n3939));
  jand g03876(.dina(n3939), .dinb(n3935), .dout(n3940));
  jand g03877(.dina(n1995), .dinb(n788), .dout(n3941));
  jand g03878(.dina(n3941), .dinb(n2620), .dout(n3942));
  jand g03879(.dina(n950), .dinb(n280), .dout(n3943));
  jand g03880(.dina(n3943), .dinb(n794), .dout(n3944));
  jand g03881(.dina(n3544), .dinb(n490), .dout(n3945));
  jand g03882(.dina(n3945), .dinb(n3944), .dout(n3946));
  jand g03883(.dina(n3946), .dinb(n3942), .dout(n3947));
  jand g03884(.dina(n3947), .dinb(n1022), .dout(n3948));
  jand g03885(.dina(n3948), .dinb(n3940), .dout(n3949));
  jand g03886(.dina(n667), .dinb(n224), .dout(n3950));
  jand g03887(.dina(n409), .dinb(n329), .dout(n3951));
  jand g03888(.dina(n3951), .dinb(n3950), .dout(n3952));
  jand g03889(.dina(n2025), .dinb(n1284), .dout(n3953));
  jand g03890(.dina(n3953), .dinb(n3952), .dout(n3954));
  jand g03891(.dina(n2812), .dinb(n1676), .dout(n3955));
  jand g03892(.dina(n1785), .dinb(n2580), .dout(n3956));
  jand g03893(.dina(n3956), .dinb(n3955), .dout(n3957));
  jand g03894(.dina(n3957), .dinb(n3954), .dout(n3958));
  jand g03895(.dina(n749), .dinb(n689), .dout(n3959));
  jand g03896(.dina(n3959), .dinb(n230), .dout(n3960));
  jand g03897(.dina(n3960), .dinb(n3092), .dout(n3961));
  jand g03898(.dina(n3961), .dinb(n1277), .dout(n3962));
  jand g03899(.dina(n3962), .dinb(n3958), .dout(n3963));
  jand g03900(.dina(n500), .dinb(n238), .dout(n3964));
  jand g03901(.dina(n3964), .dinb(n562), .dout(n3965));
  jand g03902(.dina(n365), .dinb(n197), .dout(n3966));
  jand g03903(.dina(n3966), .dinb(n1356), .dout(n3967));
  jand g03904(.dina(n2484), .dinb(n2135), .dout(n3968));
  jand g03905(.dina(n3968), .dinb(n3967), .dout(n3969));
  jand g03906(.dina(n3969), .dinb(n3965), .dout(n3970));
  jand g03907(.dina(n3970), .dinb(n2358), .dout(n3971));
  jand g03908(.dina(n3971), .dinb(n3963), .dout(n3972));
  jand g03909(.dina(n3972), .dinb(n3949), .dout(n3973));
  jand g03910(.dina(n3054), .dinb(n1285), .dout(n3974));
  jand g03911(.dina(n3974), .dinb(n3772), .dout(n3975));
  jand g03912(.dina(n427), .dinb(n292), .dout(n3976));
  jand g03913(.dina(n3976), .dinb(n1047), .dout(n3977));
  jand g03914(.dina(n3977), .dinb(n1296), .dout(n3978));
  jand g03915(.dina(n551), .dinb(n359), .dout(n3979));
  jand g03916(.dina(n3979), .dinb(n423), .dout(n3980));
  jand g03917(.dina(n3430), .dinb(n579), .dout(n3981));
  jand g03918(.dina(n3981), .dinb(n3980), .dout(n3982));
  jand g03919(.dina(n3982), .dinb(n3978), .dout(n3983));
  jand g03920(.dina(n3983), .dinb(n3975), .dout(n3984));
  jand g03921(.dina(n503), .dinb(n367), .dout(n3985));
  jand g03922(.dina(n993), .dinb(n751), .dout(n3986));
  jand g03923(.dina(n3986), .dinb(n3985), .dout(n3987));
  jand g03924(.dina(n824), .dinb(n675), .dout(n3988));
  jand g03925(.dina(n481), .dinb(n435), .dout(n3989));
  jand g03926(.dina(n3989), .dinb(n2401), .dout(n3990));
  jand g03927(.dina(n3990), .dinb(n3988), .dout(n3991));
  jand g03928(.dina(n3991), .dinb(n3987), .dout(n3992));
  jand g03929(.dina(n543), .dinb(n511), .dout(n3993));
  jand g03930(.dina(n3993), .dinb(n255), .dout(n3994));
  jand g03931(.dina(n715), .dinb(n108), .dout(n3995));
  jand g03932(.dina(n778), .dinb(n92), .dout(n3996));
  jand g03933(.dina(n3996), .dinb(n3995), .dout(n3997));
  jand g03934(.dina(n3997), .dinb(n3994), .dout(n3998));
  jand g03935(.dina(n853), .dinb(n149), .dout(n3999));
  jand g03936(.dina(n1519), .dinb(n739), .dout(n4000));
  jand g03937(.dina(n4000), .dinb(n3999), .dout(n4001));
  jand g03938(.dina(n4001), .dinb(n1643), .dout(n4002));
  jand g03939(.dina(n4002), .dinb(n3998), .dout(n4003));
  jand g03940(.dina(n467), .dinb(n311), .dout(n4004));
  jand g03941(.dina(n643), .dinb(n449), .dout(n4005));
  jand g03942(.dina(n4005), .dinb(n4004), .dout(n4006));
  jand g03943(.dina(n4006), .dinb(n1402), .dout(n4007));
  jand g03944(.dina(n4007), .dinb(n1994), .dout(n4008));
  jand g03945(.dina(n4008), .dinb(n4003), .dout(n4009));
  jand g03946(.dina(n4009), .dinb(n3992), .dout(n4010));
  jand g03947(.dina(n4010), .dinb(n3984), .dout(n4011));
  jand g03948(.dina(n4011), .dinb(n3973), .dout(n4012));
  jnot g03949(.din(n4012), .dout(n4013));
  jand g03950(.dina(n4013), .dinb(n3930), .dout(n4014));
  jnot g03951(.din(n4014), .dout(n4015));
  jand g03952(.dina(n4012), .dinb(n3929), .dout(n4016));
  jnot g03953(.din(n4016), .dout(n4017));
  jand g03954(.dina(n4017), .dinb(n72), .dout(n4018));
  jand g03955(.dina(n4018), .dinb(n4015), .dout(n4019));
  jnot g03956(.din(n4019), .dout(n4020));
  jand g03957(.dina(n4020), .dinb(n4015), .dout(n4021));
  jnot g03958(.din(n4021), .dout(n4022));
  jand g03959(.dina(n4022), .dinb(n525), .dout(n4023));
  jnot g03960(.din(n4023), .dout(n4024));
  jand g03961(.dina(n4021), .dinb(n526), .dout(n4025));
  jxor g03962(.dina(n3769), .dinb(n3768), .dout(n4026));
  jand g03963(.dina(n4026), .dinb(n732), .dout(n4027));
  jand g03964(.dina(n3851), .dinb(n1213), .dout(n4028));
  jand g03965(.dina(n3855), .dinb(n922), .dout(n4029));
  jand g03966(.dina(n3858), .dinb(n1076), .dout(n4030));
  jor  g03967(.dina(n4030), .dinb(n4029), .dout(n4031));
  jor  g03968(.dina(n4031), .dinb(n4028), .dout(n4032));
  jor  g03969(.dina(n4032), .dinb(n4027), .dout(n4033));
  jnot g03970(.din(n4033), .dout(n4034));
  jor  g03971(.dina(n4034), .dinb(n4025), .dout(n4035));
  jand g03972(.dina(n4035), .dinb(n4024), .dout(n4036));
  jor  g03973(.dina(n4036), .dinb(n3864), .dout(n4037));
  jxor g03974(.dina(n4036), .dinb(n3864), .dout(n4038));
  jnot g03975(.din(n4038), .dout(n4039));
  jand g03976(.dina(n4020), .dinb(n72), .dout(n4040));
  jand g03977(.dina(n4021), .dinb(n4017), .dout(n4041));
  jor  g03978(.dina(n4041), .dinb(n4040), .dout(n4042));
  jxor g03979(.dina(n3766), .dinb(n3765), .dout(n4043));
  jand g03980(.dina(n4043), .dinb(n732), .dout(n4044));
  jand g03981(.dina(n3855), .dinb(n1076), .dout(n4045));
  jand g03982(.dina(n3851), .dinb(n1343), .dout(n4046));
  jand g03983(.dina(n3858), .dinb(n1213), .dout(n4047));
  jor  g03984(.dina(n4047), .dinb(n4046), .dout(n4048));
  jor  g03985(.dina(n4048), .dinb(n4045), .dout(n4049));
  jor  g03986(.dina(n4049), .dinb(n4044), .dout(n4050));
  jand g03987(.dina(n4050), .dinb(n4042), .dout(n4051));
  jand g03988(.dina(n786), .dinb(n770), .dout(n4052));
  jand g03989(.dina(n4052), .dinb(n542), .dout(n4053));
  jand g03990(.dina(n470), .dinb(n392), .dout(n4054));
  jand g03991(.dina(n4054), .dinb(n2171), .dout(n4055));
  jand g03992(.dina(n4055), .dinb(n2047), .dout(n4056));
  jand g03993(.dina(n4056), .dinb(n4053), .dout(n4057));
  jand g03994(.dina(n1711), .dinb(n1385), .dout(n4058));
  jand g03995(.dina(n1580), .dinb(n1185), .dout(n4059));
  jand g03996(.dina(n4059), .dinb(n4058), .dout(n4060));
  jand g03997(.dina(n882), .dinb(n329), .dout(n4061));
  jand g03998(.dina(n4061), .dinb(n988), .dout(n4062));
  jand g03999(.dina(n2713), .dinb(n1536), .dout(n4063));
  jand g04000(.dina(n4063), .dinb(n4062), .dout(n4064));
  jand g04001(.dina(n4064), .dinb(n4060), .dout(n4065));
  jand g04002(.dina(n536), .dinb(n424), .dout(n4066));
  jand g04003(.dina(n4066), .dinb(n3463), .dout(n4067));
  jand g04004(.dina(n4067), .dinb(n1525), .dout(n4068));
  jand g04005(.dina(n4068), .dinb(n4065), .dout(n4069));
  jand g04006(.dina(n4069), .dinb(n4057), .dout(n4070));
  jand g04007(.dina(n4070), .dinb(n1825), .dout(n4071));
  jand g04008(.dina(n2892), .dinb(n108), .dout(n4072));
  jand g04009(.dina(n3129), .dinb(n2555), .dout(n4073));
  jand g04010(.dina(n4073), .dinb(n4072), .dout(n4074));
  jand g04011(.dina(n4074), .dinb(n3543), .dout(n4075));
  jand g04012(.dina(n432), .dinb(n343), .dout(n4076));
  jand g04013(.dina(n4076), .dinb(n3819), .dout(n4077));
  jand g04014(.dina(n386), .dinb(n157), .dout(n4078));
  jand g04015(.dina(n4078), .dinb(n2672), .dout(n4079));
  jand g04016(.dina(n4079), .dinb(n4077), .dout(n4080));
  jand g04017(.dina(n635), .dinb(n515), .dout(n4081));
  jand g04018(.dina(n494), .dinb(n120), .dout(n4082));
  jand g04019(.dina(n4082), .dinb(n4081), .dout(n4083));
  jand g04020(.dina(n214), .dinb(n92), .dout(n4084));
  jand g04021(.dina(n4084), .dinb(n1424), .dout(n4085));
  jand g04022(.dina(n4085), .dinb(n4083), .dout(n4086));
  jand g04023(.dina(n793), .dinb(n481), .dout(n4087));
  jand g04024(.dina(n4087), .dinb(n146), .dout(n4088));
  jand g04025(.dina(n4088), .dinb(n1485), .dout(n4089));
  jand g04026(.dina(n4089), .dinb(n4086), .dout(n4090));
  jand g04027(.dina(n4090), .dinb(n4080), .dout(n4091));
  jand g04028(.dina(n4091), .dinb(n4075), .dout(n4092));
  jand g04029(.dina(n4092), .dinb(n3180), .dout(n4093));
  jand g04030(.dina(n4093), .dinb(n4071), .dout(n4094));
  jnot g04031(.din(n4094), .dout(n4095));
  jand g04032(.dina(n4095), .dinb(n3929), .dout(n4096));
  jnot g04033(.din(n4096), .dout(n4097));
  jxor g04034(.dina(n4094), .dinb(n3930), .dout(n4098));
  jnot g04035(.din(n4098), .dout(n4099));
  jand g04036(.dina(n1780), .dinb(n1507), .dout(n4100));
  jand g04037(.dina(n552), .dinb(n197), .dout(n4101));
  jand g04038(.dina(n675), .dinb(n165), .dout(n4102));
  jand g04039(.dina(n4102), .dinb(n1150), .dout(n4103));
  jand g04040(.dina(n4103), .dinb(n4101), .dout(n4104));
  jand g04041(.dina(n4104), .dinb(n4100), .dout(n4105));
  jand g04042(.dina(n2812), .dinb(n393), .dout(n4106));
  jand g04043(.dina(n4106), .dinb(n1603), .dout(n4107));
  jand g04044(.dina(n472), .dinb(n423), .dout(n4108));
  jand g04045(.dina(n667), .dinb(n778), .dout(n4109));
  jand g04046(.dina(n4109), .dinb(n4108), .dout(n4110));
  jand g04047(.dina(n2963), .dinb(n258), .dout(n4111));
  jand g04048(.dina(n4111), .dinb(n4110), .dout(n4112));
  jand g04049(.dina(n4112), .dinb(n4107), .dout(n4113));
  jand g04050(.dina(n4113), .dinb(n4105), .dout(n4114));
  jand g04051(.dina(n4114), .dinb(n1979), .dout(n4115));
  jand g04052(.dina(n4115), .dinb(n2352), .dout(n4116));
  jand g04053(.dina(n2606), .dinb(n1594), .dout(n4117));
  jand g04054(.dina(n3662), .dinb(n433), .dout(n4118));
  jand g04055(.dina(n4118), .dinb(n4117), .dout(n4119));
  jand g04056(.dina(n450), .dinb(n371), .dout(n4120));
  jand g04057(.dina(n309), .dinb(n208), .dout(n4121));
  jand g04058(.dina(n4121), .dinb(n4120), .dout(n4122));
  jand g04059(.dina(n1034), .dinb(n274), .dout(n4123));
  jand g04060(.dina(n4123), .dinb(n1537), .dout(n4124));
  jand g04061(.dina(n4124), .dinb(n4122), .dout(n4125));
  jand g04062(.dina(n4125), .dinb(n4053), .dout(n4126));
  jand g04063(.dina(n4126), .dinb(n4119), .dout(n4127));
  jand g04064(.dina(n853), .dinb(n302), .dout(n4128));
  jand g04065(.dina(n4128), .dinb(n4066), .dout(n4129));
  jand g04066(.dina(n1145), .dinb(n225), .dout(n4130));
  jand g04067(.dina(n4130), .dinb(n4129), .dout(n4131));
  jand g04068(.dina(n1014), .dinb(n439), .dout(n4132));
  jand g04069(.dina(n4132), .dinb(n329), .dout(n4133));
  jand g04070(.dina(n749), .dinb(n103), .dout(n4134));
  jand g04071(.dina(n4134), .dinb(n330), .dout(n4135));
  jand g04072(.dina(n4135), .dinb(n4133), .dout(n4136));
  jand g04073(.dina(n4136), .dinb(n4131), .dout(n4137));
  jand g04074(.dina(n4137), .dinb(n2716), .dout(n4138));
  jand g04075(.dina(n4138), .dinb(n4127), .dout(n4139));
  jand g04076(.dina(n314), .dinb(n146), .dout(n4140));
  jand g04077(.dina(n4140), .dinb(n322), .dout(n4141));
  jand g04078(.dina(n2672), .dinb(n791), .dout(n4142));
  jand g04079(.dina(n4142), .dinb(n4141), .dout(n4143));
  jand g04080(.dina(n3800), .dinb(n2172), .dout(n4144));
  jand g04081(.dina(n4144), .dinb(n4143), .dout(n4145));
  jand g04082(.dina(n2150), .dinb(n870), .dout(n4146));
  jand g04083(.dina(n4146), .dinb(n2301), .dout(n4147));
  jand g04084(.dina(n4147), .dinb(n3629), .dout(n4148));
  jand g04085(.dina(n3093), .dinb(n375), .dout(n4149));
  jand g04086(.dina(n1039), .dinb(n633), .dout(n4150));
  jand g04087(.dina(n4150), .dinb(n435), .dout(n4151));
  jand g04088(.dina(n3046), .dinb(n1266), .dout(n4152));
  jand g04089(.dina(n4152), .dinb(n4151), .dout(n4153));
  jand g04090(.dina(n4153), .dinb(n4149), .dout(n4154));
  jand g04091(.dina(n4154), .dinb(n4148), .dout(n4155));
  jand g04092(.dina(n4155), .dinb(n4145), .dout(n4156));
  jand g04093(.dina(n4156), .dinb(n4139), .dout(n4157));
  jand g04094(.dina(n4157), .dinb(n4116), .dout(n4158));
  jnot g04095(.din(n4158), .dout(n4159));
  jand g04096(.dina(n678), .dinb(n377), .dout(n4160));
  jand g04097(.dina(n478), .dinb(n92), .dout(n4161));
  jand g04098(.dina(n4161), .dinb(n4160), .dout(n4162));
  jand g04099(.dina(n432), .dinb(n405), .dout(n4163));
  jand g04100(.dina(n4163), .dinb(n2041), .dout(n4164));
  jand g04101(.dina(n4164), .dinb(n4162), .dout(n4165));
  jand g04102(.dina(n1627), .dinb(n1193), .dout(n4166));
  jand g04103(.dina(n711), .dinb(n217), .dout(n4167));
  jand g04104(.dina(n4167), .dinb(n4004), .dout(n4168));
  jand g04105(.dina(n4168), .dinb(n4166), .dout(n4169));
  jand g04106(.dina(n4169), .dinb(n4165), .dout(n4170));
  jand g04107(.dina(n671), .dinb(n249), .dout(n4171));
  jand g04108(.dina(n4171), .dinb(n221), .dout(n4172));
  jand g04109(.dina(n3594), .dinb(n1830), .dout(n4173));
  jand g04110(.dina(n4173), .dinb(n4172), .dout(n4174));
  jand g04111(.dina(n3462), .dinb(n2014), .dout(n4175));
  jand g04112(.dina(n4175), .dinb(n2963), .dout(n4176));
  jand g04113(.dina(n3097), .dinb(n1711), .dout(n4177));
  jand g04114(.dina(n1584), .dinb(n868), .dout(n4178));
  jand g04115(.dina(n4178), .dinb(n4177), .dout(n4179));
  jand g04116(.dina(n4179), .dinb(n4176), .dout(n4180));
  jand g04117(.dina(n4180), .dinb(n4174), .dout(n4181));
  jand g04118(.dina(n4181), .dinb(n4170), .dout(n4182));
  jand g04119(.dina(n2130), .dinb(n336), .dout(n4183));
  jand g04120(.dina(n4183), .dinb(n667), .dout(n4184));
  jand g04121(.dina(n1144), .dinb(n965), .dout(n4185));
  jand g04122(.dina(n853), .dinb(n352), .dout(n4186));
  jand g04123(.dina(n4186), .dinb(n4185), .dout(n4187));
  jand g04124(.dina(n1663), .dinb(n1259), .dout(n4188));
  jand g04125(.dina(n4188), .dinb(n4187), .dout(n4189));
  jand g04126(.dina(n1492), .dinb(n926), .dout(n4190));
  jand g04127(.dina(n626), .dinb(n395), .dout(n4191));
  jand g04128(.dina(n4191), .dinb(n238), .dout(n4192));
  jand g04129(.dina(n4192), .dinb(n4190), .dout(n4193));
  jand g04130(.dina(n4193), .dinb(n4189), .dout(n4194));
  jand g04131(.dina(n4194), .dinb(n4184), .dout(n4195));
  jand g04132(.dina(n1506), .dinb(n1428), .dout(n4196));
  jand g04133(.dina(n1099), .dinb(n1057), .dout(n4197));
  jand g04134(.dina(n4197), .dinb(n4196), .dout(n4198));
  jand g04135(.dina(n503), .dinb(n329), .dout(n4199));
  jand g04136(.dina(n4199), .dinb(n719), .dout(n4200));
  jand g04137(.dina(n423), .dinb(n190), .dout(n4201));
  jand g04138(.dina(n897), .dinb(n382), .dout(n4202));
  jand g04139(.dina(n4202), .dinb(n4201), .dout(n4203));
  jand g04140(.dina(n4203), .dinb(n4200), .dout(n4204));
  jand g04141(.dina(n4204), .dinb(n4198), .dout(n4205));
  jand g04142(.dina(n4205), .dinb(n2405), .dout(n4206));
  jand g04143(.dina(n4206), .dinb(n4195), .dout(n4207));
  jand g04144(.dina(n1231), .dinb(n234), .dout(n4208));
  jand g04145(.dina(n1014), .dinb(n214), .dout(n4209));
  jand g04146(.dina(n4209), .dinb(n4208), .dout(n4210));
  jand g04147(.dina(n1597), .dinb(n391), .dout(n4211));
  jand g04148(.dina(n786), .dinb(n418), .dout(n4212));
  jand g04149(.dina(n4212), .dinb(n4211), .dout(n4213));
  jand g04150(.dina(n4213), .dinb(n4210), .dout(n4214));
  jand g04151(.dina(n967), .dinb(n857), .dout(n4215));
  jand g04152(.dina(n4215), .dinb(n476), .dout(n4216));
  jand g04153(.dina(n396), .dinb(n288), .dout(n4217));
  jand g04154(.dina(n529), .dinb(n517), .dout(n4218));
  jand g04155(.dina(n4218), .dinb(n4217), .dout(n4219));
  jand g04156(.dina(n4219), .dinb(n4216), .dout(n4220));
  jand g04157(.dina(n4220), .dinb(n4214), .dout(n4221));
  jand g04158(.dina(n1129), .dinb(n554), .dout(n4222));
  jand g04159(.dina(n1009), .dinb(n451), .dout(n4223));
  jand g04160(.dina(n4223), .dinb(n4222), .dout(n4224));
  jand g04161(.dina(n793), .dinb(n103), .dout(n4225));
  jand g04162(.dina(n707), .dinb(n305), .dout(n4226));
  jand g04163(.dina(n4226), .dinb(n4225), .dout(n4227));
  jand g04164(.dina(n4227), .dinb(n3136), .dout(n4228));
  jand g04165(.dina(n4228), .dinb(n4224), .dout(n4229));
  jand g04166(.dina(n4229), .dinb(n4221), .dout(n4230));
  jnot g04167(.din(n3339), .dout(n4231));
  jand g04168(.dina(n486), .dinb(n208), .dout(n4232));
  jand g04169(.dina(n4232), .dinb(n1349), .dout(n4233));
  jand g04170(.dina(n4233), .dinb(n4231), .dout(n4234));
  jand g04171(.dina(n3401), .dinb(n633), .dout(n4235));
  jand g04172(.dina(n366), .dinb(n245), .dout(n4236));
  jand g04173(.dina(n4236), .dinb(n801), .dout(n4237));
  jand g04174(.dina(n4237), .dinb(n4235), .dout(n4238));
  jand g04175(.dina(n4238), .dinb(n4234), .dout(n4239));
  jand g04176(.dina(n4239), .dinb(n918), .dout(n4240));
  jand g04177(.dina(n4240), .dinb(n4230), .dout(n4241));
  jand g04178(.dina(n4241), .dinb(n4207), .dout(n4242));
  jand g04179(.dina(n4242), .dinb(n4182), .dout(n4243));
  jnot g04180(.din(n4243), .dout(n4244));
  jand g04181(.dina(n4244), .dinb(n4159), .dout(n4245));
  jnot g04182(.din(n4245), .dout(n4246));
  jnot g04183(.din(\a[20] ), .dout(n4247));
  jand g04184(.dina(n4243), .dinb(n4158), .dout(n4248));
  jnot g04185(.din(n4248), .dout(n4249));
  jand g04186(.dina(n4249), .dinb(n4247), .dout(n4250));
  jand g04187(.dina(n4250), .dinb(n4246), .dout(n4251));
  jnot g04188(.din(n4251), .dout(n4252));
  jand g04189(.dina(n4252), .dinb(n4246), .dout(n4253));
  jnot g04190(.din(n4253), .dout(n4254));
  jand g04191(.dina(n4254), .dinb(n4094), .dout(n4255));
  jnot g04192(.din(n4255), .dout(n4256));
  jand g04193(.dina(n4253), .dinb(n4095), .dout(n4257));
  jxor g04194(.dina(n3760), .dinb(n3759), .dout(n4258));
  jand g04195(.dina(n4258), .dinb(n732), .dout(n4259));
  jand g04196(.dina(n3855), .dinb(n1343), .dout(n4260));
  jand g04197(.dina(n3851), .dinb(n1560), .dout(n4261));
  jand g04198(.dina(n3858), .dinb(n1445), .dout(n4262));
  jor  g04199(.dina(n4262), .dinb(n4261), .dout(n4263));
  jor  g04200(.dina(n4263), .dinb(n4260), .dout(n4264));
  jor  g04201(.dina(n4264), .dinb(n4259), .dout(n4265));
  jnot g04202(.din(n4265), .dout(n4266));
  jor  g04203(.dina(n4266), .dinb(n4257), .dout(n4267));
  jand g04204(.dina(n4267), .dinb(n4256), .dout(n4268));
  jor  g04205(.dina(n4268), .dinb(n4099), .dout(n4269));
  jand g04206(.dina(n4269), .dinb(n4097), .dout(n4270));
  jnot g04207(.din(n4270), .dout(n4271));
  jxor g04208(.dina(n4050), .dinb(n4042), .dout(n4272));
  jand g04209(.dina(n4272), .dinb(n4271), .dout(n4273));
  jor  g04210(.dina(n4273), .dinb(n4051), .dout(n4274));
  jxor g04211(.dina(n4021), .dinb(n526), .dout(n4275));
  jxor g04212(.dina(n4275), .dinb(n4033), .dout(n4276));
  jand g04213(.dina(n4276), .dinb(n4274), .dout(n4277));
  jnot g04214(.din(n4277), .dout(n4278));
  jxor g04215(.dina(n4276), .dinb(n4274), .dout(n4279));
  jnot g04216(.din(n4279), .dout(n4280));
  jand g04217(.dina(n4108), .dinb(n3462), .dout(n4281));
  jand g04218(.dina(n4281), .dinb(n697), .dout(n4282));
  jand g04219(.dina(n1034), .dinb(n197), .dout(n4283));
  jand g04220(.dina(n4283), .dinb(n3236), .dout(n4284));
  jand g04221(.dina(n4076), .dinb(n3839), .dout(n4285));
  jand g04222(.dina(n4285), .dinb(n4284), .dout(n4286));
  jand g04223(.dina(n516), .dinb(n322), .dout(n4287));
  jand g04224(.dina(n4287), .dinb(n2620), .dout(n4288));
  jand g04225(.dina(n913), .dinb(n847), .dout(n4289));
  jand g04226(.dina(n157), .dinb(n103), .dout(n4290));
  jand g04227(.dina(n4290), .dinb(n4289), .dout(n4291));
  jand g04228(.dina(n4291), .dinb(n4288), .dout(n4292));
  jand g04229(.dina(n4292), .dinb(n4286), .dout(n4293));
  jand g04230(.dina(n4293), .dinb(n4282), .dout(n4294));
  jand g04231(.dina(n404), .dinb(n134), .dout(n4295));
  jand g04232(.dina(n503), .dinb(n431), .dout(n4296));
  jand g04233(.dina(n4296), .dinb(n208), .dout(n4297));
  jand g04234(.dina(n4297), .dinb(n4295), .dout(n4298));
  jand g04235(.dina(n194), .dinb(n130), .dout(n4299));
  jand g04236(.dina(n4299), .dinb(n938), .dout(n4300));
  jand g04237(.dina(n439), .dinb(n396), .dout(n4301));
  jand g04238(.dina(n4301), .dinb(n1499), .dout(n4302));
  jand g04239(.dina(n4302), .dinb(n4300), .dout(n4303));
  jand g04240(.dina(n4303), .dinb(n4298), .dout(n4304));
  jand g04241(.dina(n4304), .dinb(n2559), .dout(n4305));
  jand g04242(.dina(n778), .dinb(n566), .dout(n4306));
  jand g04243(.dina(n4306), .dinb(n270), .dout(n4307));
  jand g04244(.dina(n967), .dinb(n739), .dout(n4308));
  jand g04245(.dina(n4308), .dinb(n1958), .dout(n4309));
  jand g04246(.dina(n4309), .dinb(n4307), .dout(n4310));
  jnot g04247(.din(n1747), .dout(n4311));
  jand g04248(.dina(n4311), .dinb(n658), .dout(n4312));
  jand g04249(.dina(n4312), .dinb(n4310), .dout(n4313));
  jand g04250(.dina(n1627), .dinb(n880), .dout(n4314));
  jand g04251(.dina(n909), .dinb(n833), .dout(n4315));
  jand g04252(.dina(n719), .dinb(n467), .dout(n4316));
  jand g04253(.dina(n860), .dinb(n715), .dout(n4317));
  jand g04254(.dina(n4317), .dinb(n4316), .dout(n4318));
  jand g04255(.dina(n4318), .dinb(n4315), .dout(n4319));
  jand g04256(.dina(n4319), .dinb(n4314), .dout(n4320));
  jand g04257(.dina(n4320), .dinb(n4313), .dout(n4321));
  jand g04258(.dina(n4321), .dinb(n4305), .dout(n4322));
  jand g04259(.dina(n4322), .dinb(n4294), .dout(n4323));
  jand g04260(.dina(n988), .dinb(n372), .dout(n4324));
  jand g04261(.dina(n4324), .dinb(n818), .dout(n4325));
  jand g04262(.dina(n4325), .dinb(n2228), .dout(n4326));
  jand g04263(.dina(n993), .dinb(n311), .dout(n4327));
  jand g04264(.dina(n4327), .dinb(n238), .dout(n4328));
  jand g04265(.dina(n4328), .dinb(n2256), .dout(n4329));
  jand g04266(.dina(n4329), .dinb(n3787), .dout(n4330));
  jand g04267(.dina(n4330), .dinb(n4326), .dout(n4331));
  jand g04268(.dina(n3544), .dinb(n314), .dout(n4332));
  jand g04269(.dina(n4332), .dinb(n626), .dout(n4333));
  jand g04270(.dina(n1014), .dinb(n888), .dout(n4334));
  jand g04271(.dina(n4334), .dinb(n997), .dout(n4335));
  jand g04272(.dina(n876), .dinb(n853), .dout(n4336));
  jand g04273(.dina(n4336), .dinb(n3066), .dout(n4337));
  jand g04274(.dina(n4337), .dinb(n3662), .dout(n4338));
  jand g04275(.dina(n4338), .dinb(n4335), .dout(n4339));
  jand g04276(.dina(n4339), .dinb(n4333), .dout(n4340));
  jand g04277(.dina(n595), .dinb(n82), .dout(n4341));
  jand g04278(.dina(n926), .dinb(n857), .dout(n4342));
  jand g04279(.dina(n4342), .dinb(n4341), .dout(n4343));
  jand g04280(.dina(n1178), .dinb(n689), .dout(n4344));
  jand g04281(.dina(n4344), .dinb(n3445), .dout(n4345));
  jand g04282(.dina(n1500), .dinb(n1142), .dout(n4346));
  jand g04283(.dina(n4346), .dinb(n4345), .dout(n4347));
  jand g04284(.dina(n4347), .dinb(n4343), .dout(n4348));
  jand g04285(.dina(n2369), .dinb(n180), .dout(n4349));
  jand g04286(.dina(n4349), .dinb(n756), .dout(n4350));
  jand g04287(.dina(n1997), .dinb(n802), .dout(n4351));
  jand g04288(.dina(n4351), .dinb(n869), .dout(n4352));
  jand g04289(.dina(n4352), .dinb(n4350), .dout(n4353));
  jand g04290(.dina(n4353), .dinb(n4348), .dout(n4354));
  jand g04291(.dina(n4354), .dinb(n4340), .dout(n4355));
  jand g04292(.dina(n4355), .dinb(n4331), .dout(n4356));
  jand g04293(.dina(n4356), .dinb(n4323), .dout(n4357));
  jnot g04294(.din(n4357), .dout(n4358));
  jand g04295(.dina(n4358), .dinb(n3853), .dout(n4359));
  jand g04296(.dina(n3853), .dinb(n922), .dout(n4360));
  jand g04297(.dina(n3847), .dinb(n3771), .dout(n4361));
  jor  g04298(.dina(n4361), .dinb(n4360), .dout(n4362));
  jxor g04299(.dina(n4357), .dinb(n3846), .dout(n4363));
  jand g04300(.dina(n4363), .dinb(n4362), .dout(n4364));
  jor  g04301(.dina(n4364), .dinb(n4359), .dout(n4365));
  jand g04302(.dina(n926), .dinb(n120), .dout(n4366));
  jand g04303(.dina(n4366), .dinb(n2887), .dout(n4367));
  jand g04304(.dina(n4367), .dinb(n891), .dout(n4368));
  jand g04305(.dina(n503), .dinb(n157), .dout(n4369));
  jand g04306(.dina(n1346), .dinb(n633), .dout(n4370));
  jand g04307(.dina(n4370), .dinb(n4369), .dout(n4371));
  jand g04308(.dina(n4371), .dinb(n4101), .dout(n4372));
  jand g04309(.dina(n4372), .dinb(n4368), .dout(n4373));
  jand g04310(.dina(n4373), .dinb(n4333), .dout(n4374));
  jand g04311(.dina(n4374), .dinb(n4313), .dout(n4375));
  jand g04312(.dina(n4375), .dinb(n4331), .dout(n4376));
  jand g04313(.dina(n979), .dinb(n260), .dout(n4377));
  jand g04314(.dina(n4377), .dinb(n1287), .dout(n4378));
  jand g04315(.dina(n3160), .dinb(n803), .dout(n4379));
  jand g04316(.dina(n4379), .dinb(n2299), .dout(n4380));
  jand g04317(.dina(n4380), .dinb(n4378), .dout(n4381));
  jand g04318(.dina(n749), .dinb(n317), .dout(n4382));
  jand g04319(.dina(n4382), .dinb(n3950), .dout(n4383));
  jand g04320(.dina(n1066), .dinb(n174), .dout(n4384));
  jand g04321(.dina(n4384), .dinb(n2227), .dout(n4385));
  jand g04322(.dina(n4385), .dinb(n4383), .dout(n4386));
  jnot g04323(.din(n1487), .dout(n4387));
  jor  g04324(.dina(n3302), .dinb(n4387), .dout(n4388));
  jnot g04325(.din(n4388), .dout(n4389));
  jand g04326(.dina(n4389), .dinb(n1322), .dout(n4390));
  jand g04327(.dina(n4390), .dinb(n4386), .dout(n4391));
  jand g04328(.dina(n4391), .dinb(n4381), .dout(n4392));
  jand g04329(.dina(n763), .dinb(n385), .dout(n4393));
  jand g04330(.dina(n4393), .dinb(n1305), .dout(n4394));
  jand g04331(.dina(n3550), .dinb(n2897), .dout(n4395));
  jand g04332(.dina(n4395), .dinb(n2150), .dout(n4396));
  jand g04333(.dina(n4396), .dinb(n4394), .dout(n4397));
  jand g04334(.dina(n4397), .dinb(n3641), .dout(n4398));
  jand g04335(.dina(n478), .dinb(n375), .dout(n4399));
  jand g04336(.dina(n4399), .dinb(n1334), .dout(n4400));
  jand g04337(.dina(n2663), .dinb(n1167), .dout(n4401));
  jand g04338(.dina(n4401), .dinb(n1024), .dout(n4402));
  jand g04339(.dina(n4402), .dinb(n4400), .dout(n4403));
  jand g04340(.dina(n4403), .dinb(n790), .dout(n4404));
  jand g04341(.dina(n4404), .dinb(n4398), .dout(n4405));
  jand g04342(.dina(n4405), .dinb(n4392), .dout(n4406));
  jand g04343(.dina(n1144), .dinb(n443), .dout(n4407));
  jand g04344(.dina(n4407), .dinb(n309), .dout(n4408));
  jand g04345(.dina(n1184), .dinb(n517), .dout(n4409));
  jand g04346(.dina(n4409), .dinb(n2564), .dout(n4410));
  jand g04347(.dina(n4410), .dinb(n4408), .dout(n4411));
  jand g04348(.dina(n4411), .dinb(n2366), .dout(n4412));
  jand g04349(.dina(n4412), .dinb(n1231), .dout(n4413));
  jand g04350(.dina(n4413), .dinb(n352), .dout(n4414));
  jand g04351(.dina(n4414), .dinb(n4406), .dout(n4415));
  jand g04352(.dina(n4415), .dinb(n4376), .dout(n4416));
  jand g04353(.dina(n449), .dinb(n290), .dout(n4417));
  jand g04354(.dina(n4417), .dinb(n433), .dout(n4418));
  jand g04355(.dina(n4418), .dinb(n1349), .dout(n4419));
  jand g04356(.dina(n4419), .dinb(n3071), .dout(n4420));
  jand g04357(.dina(n2118), .dinb(n357), .dout(n4421));
  jand g04358(.dina(n907), .dinb(n284), .dout(n4422));
  jand g04359(.dina(n4422), .dinb(n1142), .dout(n4423));
  jand g04360(.dina(n4423), .dinb(n693), .dout(n4424));
  jand g04361(.dina(n4424), .dinb(n4421), .dout(n4425));
  jand g04362(.dina(n4425), .dinb(n3836), .dout(n4426));
  jand g04363(.dina(n4426), .dinb(n4420), .dout(n4427));
  jnot g04364(.din(n3350), .dout(n4428));
  jand g04365(.dina(n574), .dinb(n365), .dout(n4429));
  jand g04366(.dina(n4429), .dinb(n234), .dout(n4430));
  jand g04367(.dina(n302), .dinb(n249), .dout(n4431));
  jand g04368(.dina(n553), .dinb(n190), .dout(n4432));
  jand g04369(.dina(n4432), .dinb(n4431), .dout(n4433));
  jand g04370(.dina(n4433), .dinb(n4430), .dout(n4434));
  jand g04371(.dina(n4434), .dinb(n4428), .dout(n4435));
  jand g04372(.dina(n694), .dinb(n324), .dout(n4436));
  jand g04373(.dina(n472), .dinb(n208), .dout(n4437));
  jand g04374(.dina(n4437), .dinb(n467), .dout(n4438));
  jand g04375(.dina(n4438), .dinb(n4436), .dout(n4439));
  jand g04376(.dina(n2033), .dinb(n824), .dout(n4440));
  jand g04377(.dina(n4440), .dinb(n4439), .dout(n4441));
  jand g04378(.dina(n4441), .dinb(n4435), .dout(n4442));
  jand g04379(.dina(n4442), .dinb(n4427), .dout(n4443));
  jand g04380(.dina(n4443), .dinb(n4416), .dout(n4444));
  jxor g04381(.dina(n4444), .dinb(n4357), .dout(n4445));
  jxor g04382(.dina(n4445), .dinb(n4365), .dout(n4446));
  jxor g04383(.dina(\a[27] ), .dinb(\a[26] ), .dout(n4447));
  jxor g04384(.dina(\a[29] ), .dinb(\a[28] ), .dout(n4448));
  jand g04385(.dina(n4448), .dinb(n4447), .dout(n4449));
  jand g04386(.dina(n4449), .dinb(n4446), .dout(n4450));
  jnot g04387(.din(n4444), .dout(n4451));
  jnot g04388(.din(n4448), .dout(n4452));
  jand g04389(.dina(n4452), .dinb(n4447), .dout(n4453));
  jand g04390(.dina(n4453), .dinb(n4451), .dout(n4454));
  jnot g04391(.din(n4447), .dout(n4455));
  jxor g04392(.dina(\a[28] ), .dinb(\a[27] ), .dout(n4456));
  jand g04393(.dina(n4456), .dinb(n4455), .dout(n4457));
  jand g04394(.dina(n4457), .dinb(n4358), .dout(n4458));
  jor  g04395(.dina(n4456), .dinb(n4447), .dout(n4459));
  jnot g04396(.din(n4459), .dout(n4460));
  jand g04397(.dina(n4460), .dinb(n4448), .dout(n4461));
  jand g04398(.dina(n4461), .dinb(n3853), .dout(n4462));
  jor  g04399(.dina(n4462), .dinb(n4458), .dout(n4463));
  jor  g04400(.dina(n4463), .dinb(n4454), .dout(n4464));
  jor  g04401(.dina(n4464), .dinb(n4450), .dout(n4465));
  jxor g04402(.dina(n4465), .dinb(n88), .dout(n4466));
  jor  g04403(.dina(n4466), .dinb(n4280), .dout(n4467));
  jand g04404(.dina(n4467), .dinb(n4278), .dout(n4468));
  jor  g04405(.dina(n4468), .dinb(n4039), .dout(n4469));
  jand g04406(.dina(n4469), .dinb(n4037), .dout(n4470));
  jnot g04407(.din(n4470), .dout(n4471));
  jor  g04408(.dina(n728), .dinb(n526), .dout(n4472));
  jand g04409(.dina(n3862), .dinb(n729), .dout(n4473));
  jnot g04410(.din(n4473), .dout(n4474));
  jand g04411(.dina(n4474), .dinb(n4472), .dout(n4475));
  jand g04412(.dina(n583), .dinb(n157), .dout(n4476));
  jand g04413(.dina(n641), .dinb(n542), .dout(n4477));
  jand g04414(.dina(n4477), .dinb(n4476), .dout(n4478));
  jand g04415(.dina(n1898), .dinb(n239), .dout(n4479));
  jand g04416(.dina(n4479), .dinb(n2484), .dout(n4480));
  jand g04417(.dina(n4480), .dinb(n4478), .dout(n4481));
  jand g04418(.dina(n793), .dinb(n322), .dout(n4482));
  jand g04419(.dina(n4482), .dinb(n286), .dout(n4483));
  jand g04420(.dina(n778), .dinb(n483), .dout(n4484));
  jand g04421(.dina(n988), .dinb(n274), .dout(n4485));
  jand g04422(.dina(n4485), .dinb(n4484), .dout(n4486));
  jand g04423(.dina(n860), .dinb(n309), .dout(n4487));
  jand g04424(.dina(n4487), .dinb(n1424), .dout(n4488));
  jand g04425(.dina(n4488), .dinb(n4486), .dout(n4489));
  jand g04426(.dina(n4489), .dinb(n4483), .dout(n4490));
  jand g04427(.dina(n1278), .dinb(n1023), .dout(n4491));
  jand g04428(.dina(n4491), .dinb(n2228), .dout(n4492));
  jand g04429(.dina(n1598), .dinb(n722), .dout(n4493));
  jand g04430(.dina(n967), .dinb(n874), .dout(n4494));
  jand g04431(.dina(n4494), .dinb(n2301), .dout(n4495));
  jand g04432(.dina(n4495), .dinb(n4493), .dout(n4496));
  jand g04433(.dina(n4496), .dinb(n4492), .dout(n4497));
  jand g04434(.dina(n4497), .dinb(n4490), .dout(n4498));
  jand g04435(.dina(n4498), .dinb(n4481), .dout(n4499));
  jand g04436(.dina(n707), .dinb(n375), .dout(n4500));
  jand g04437(.dina(n1047), .dinb(n302), .dout(n4501));
  jand g04438(.dina(n4501), .dinb(n4500), .dout(n4502));
  jand g04439(.dina(n843), .dinb(n346), .dout(n4503));
  jand g04440(.dina(n432), .dinb(n180), .dout(n4504));
  jand g04441(.dina(n4504), .dinb(n4503), .dout(n4505));
  jand g04442(.dina(n1160), .dinb(n960), .dout(n4506));
  jand g04443(.dina(n4506), .dinb(n4505), .dout(n4507));
  jand g04444(.dina(n4507), .dinb(n4502), .dout(n4508));
  jand g04445(.dina(n4508), .dinb(n3961), .dout(n4509));
  jand g04446(.dina(n1216), .dinb(n1067), .dout(n4510));
  jand g04447(.dina(n1432), .dinb(n198), .dout(n4511));
  jand g04448(.dina(n4511), .dinb(n4510), .dout(n4512));
  jnot g04449(.din(n2077), .dout(n4513));
  jand g04450(.dina(n517), .dinb(n276), .dout(n4514));
  jand g04451(.dina(n4514), .dinb(n4513), .dout(n4515));
  jand g04452(.dina(n511), .dinb(n1031), .dout(n4516));
  jand g04453(.dina(n1144), .dinb(n893), .dout(n4517));
  jand g04454(.dina(n4517), .dinb(n4516), .dout(n4518));
  jand g04455(.dina(n4518), .dinb(n4515), .dout(n4519));
  jand g04456(.dina(n4519), .dinb(n4512), .dout(n4520));
  jand g04457(.dina(n268), .dinb(n161), .dout(n4521));
  jand g04458(.dina(n4521), .dinb(n826), .dout(n4522));
  jand g04459(.dina(n4522), .dinb(n218), .dout(n4523));
  jand g04460(.dina(n3896), .dinb(n3250), .dout(n4524));
  jand g04461(.dina(n4524), .dinb(n2378), .dout(n4525));
  jand g04462(.dina(n4525), .dinb(n4523), .dout(n4526));
  jand g04463(.dina(n4526), .dinb(n4520), .dout(n4527));
  jand g04464(.dina(n4527), .dinb(n4509), .dout(n4528));
  jand g04465(.dina(n4528), .dinb(n4499), .dout(n4529));
  jand g04466(.dina(n4529), .dinb(n3573), .dout(n4530));
  jnot g04467(.din(n4530), .dout(n4531));
  jand g04468(.dina(n4531), .dinb(n526), .dout(n4532));
  jnot g04469(.din(n4532), .dout(n4533));
  jand g04470(.dina(n4530), .dinb(n525), .dout(n4534));
  jnot g04471(.din(n4534), .dout(n4535));
  jand g04472(.dina(n4535), .dinb(n68), .dout(n4536));
  jand g04473(.dina(n4536), .dinb(n4533), .dout(n4537));
  jor  g04474(.dina(n4537), .dinb(\a[26] ), .dout(n4538));
  jor  g04475(.dina(n4536), .dinb(n4532), .dout(n4539));
  jnot g04476(.din(n4539), .dout(n4540));
  jand g04477(.dina(n4540), .dinb(n4535), .dout(n4541));
  jnot g04478(.din(n4541), .dout(n4542));
  jand g04479(.dina(n4542), .dinb(n4538), .dout(n4543));
  jxor g04480(.dina(n4543), .dinb(n4475), .dout(n4544));
  jxor g04481(.dina(n4363), .dinb(n4362), .dout(n4545));
  jand g04482(.dina(n4545), .dinb(n732), .dout(n4546));
  jand g04483(.dina(n3851), .dinb(n922), .dout(n4547));
  jand g04484(.dina(n4358), .dinb(n3855), .dout(n4548));
  jand g04485(.dina(n3858), .dinb(n3853), .dout(n4549));
  jor  g04486(.dina(n4549), .dinb(n4548), .dout(n4550));
  jor  g04487(.dina(n4550), .dinb(n4547), .dout(n4551));
  jor  g04488(.dina(n4551), .dinb(n4546), .dout(n4552));
  jxor g04489(.dina(n4552), .dinb(n4544), .dout(n4553));
  jand g04490(.dina(n4553), .dinb(n4471), .dout(n4554));
  jand g04491(.dina(n757), .dinb(n413), .dout(n4555));
  jand g04492(.dina(n4555), .dinb(n246), .dout(n4556));
  jand g04493(.dina(n4556), .dinb(n1727), .dout(n4557));
  jand g04494(.dina(n2261), .dinb(n827), .dout(n4558));
  jand g04495(.dina(n700), .dinb(n234), .dout(n4559));
  jand g04496(.dina(n516), .dinb(n343), .dout(n4560));
  jand g04497(.dina(n4560), .dinb(n4559), .dout(n4561));
  jand g04498(.dina(n4561), .dinb(n4558), .dout(n4562));
  jand g04499(.dina(n4562), .dinb(n4557), .dout(n4563));
  jand g04500(.dina(n4563), .dinb(n3279), .dout(n4564));
  jand g04501(.dina(n4564), .dinb(n4420), .dout(n4565));
  jand g04502(.dina(n4565), .dinb(n3040), .dout(n4566));
  jand g04503(.dina(n751), .dinb(n622), .dout(n4567));
  jand g04504(.dina(n537), .dinb(n501), .dout(n4568));
  jand g04505(.dina(n4568), .dinb(n4567), .dout(n4569));
  jand g04506(.dina(n4211), .dinb(n712), .dout(n4570));
  jand g04507(.dina(n1881), .dinb(n1196), .dout(n4571));
  jand g04508(.dina(n4571), .dinb(n4570), .dout(n4572));
  jand g04509(.dina(n4572), .dinb(n1267), .dout(n4573));
  jand g04510(.dina(n4573), .dinb(n4569), .dout(n4574));
  jand g04511(.dina(n643), .dinb(n586), .dout(n4575));
  jand g04512(.dina(n4575), .dinb(n218), .dout(n4576));
  jand g04513(.dina(n515), .dinb(n149), .dout(n4577));
  jand g04514(.dina(n4577), .dinb(n4576), .dout(n4578));
  jand g04515(.dina(n4578), .dinb(n4574), .dout(n4579));
  jand g04516(.dina(n932), .dinb(n606), .dout(n4580));
  jand g04517(.dina(n4580), .dinb(n4349), .dout(n4581));
  jand g04518(.dina(n4581), .dinb(n4579), .dout(n4582));
  jand g04519(.dina(n4582), .dinb(n4566), .dout(n4583));
  jand g04520(.dina(n950), .dinb(n876), .dout(n4584));
  jand g04521(.dina(n4584), .dinb(n1014), .dout(n4585));
  jand g04522(.dina(n4585), .dinb(n688), .dout(n4586));
  jand g04523(.dina(n4586), .dinb(n855), .dout(n4587));
  jand g04524(.dina(n1584), .dinb(n1295), .dout(n4588));
  jand g04525(.dina(n4588), .dinb(n1057), .dout(n4589));
  jand g04526(.dina(n756), .dinb(n352), .dout(n4590));
  jand g04527(.dina(n4590), .dinb(n4431), .dout(n4591));
  jand g04528(.dina(n4591), .dinb(n1488), .dout(n4592));
  jand g04529(.dina(n4592), .dinb(n4589), .dout(n4593));
  jand g04530(.dina(n4593), .dinb(n4587), .dout(n4594));
  jand g04531(.dina(n1153), .dinb(n330), .dout(n4595));
  jand g04532(.dina(n4595), .dinb(n4594), .dout(n4596));
  jand g04533(.dina(n4596), .dinb(n4583), .dout(n4597));
  jnot g04534(.din(n4597), .dout(n4598));
  jand g04535(.dina(n4598), .dinb(n4451), .dout(n4599));
  jand g04536(.dina(n4451), .dinb(n4358), .dout(n4600));
  jand g04537(.dina(n4445), .dinb(n4365), .dout(n4601));
  jor  g04538(.dina(n4601), .dinb(n4600), .dout(n4602));
  jxor g04539(.dina(n4597), .dinb(n4444), .dout(n4603));
  jand g04540(.dina(n4603), .dinb(n4602), .dout(n4604));
  jor  g04541(.dina(n4604), .dinb(n4599), .dout(n4605));
  jand g04542(.dina(n4439), .dinb(n1153), .dout(n4606));
  jand g04543(.dina(n806), .dinb(n596), .dout(n4607));
  jand g04544(.dina(n4607), .dinb(n1104), .dout(n4608));
  jand g04545(.dina(n1039), .dinb(n346), .dout(n4609));
  jand g04546(.dina(n4609), .dinb(n4295), .dout(n4610));
  jand g04547(.dina(n692), .dinb(n230), .dout(n4611));
  jand g04548(.dina(n4611), .dinb(n2659), .dout(n4612));
  jand g04549(.dina(n4612), .dinb(n4610), .dout(n4613));
  jand g04550(.dina(n4613), .dinb(n4608), .dout(n4614));
  jand g04551(.dina(n1047), .dinb(n893), .dout(n4615));
  jand g04552(.dina(n4615), .dinb(n486), .dout(n4616));
  jand g04553(.dina(n2834), .dinb(n463), .dout(n4617));
  jand g04554(.dina(n4617), .dinb(n4616), .dout(n4618));
  jand g04555(.dina(n1615), .dinb(n909), .dout(n4619));
  jand g04556(.dina(n4619), .dinb(n2315), .dout(n4620));
  jand g04557(.dina(n4620), .dinb(n2583), .dout(n4621));
  jand g04558(.dina(n3092), .dinb(n598), .dout(n4622));
  jand g04559(.dina(n1345), .dinb(n1142), .dout(n4623));
  jand g04560(.dina(n4623), .dinb(n4622), .dout(n4624));
  jand g04561(.dina(n4624), .dinb(n4621), .dout(n4625));
  jand g04562(.dina(n4625), .dinb(n4618), .dout(n4626));
  jand g04563(.dina(n4626), .dinb(n4614), .dout(n4627));
  jand g04564(.dina(n4627), .dinb(n154), .dout(n4628));
  jand g04565(.dina(n4628), .dinb(n4606), .dout(n4629));
  jand g04566(.dina(n4629), .dinb(n4594), .dout(n4630));
  jnot g04567(.din(n4630), .dout(n4631));
  jand g04568(.dina(n4631), .dinb(n4598), .dout(n4632));
  jand g04569(.dina(n4629), .dinb(n4597), .dout(n4633));
  jor  g04570(.dina(n4633), .dinb(n4632), .dout(n4634));
  jnot g04571(.din(n4634), .dout(n4635));
  jxor g04572(.dina(n4635), .dinb(n4605), .dout(n4636));
  jand g04573(.dina(n4636), .dinb(n4449), .dout(n4637));
  jand g04574(.dina(n4461), .dinb(n4451), .dout(n4638));
  jand g04575(.dina(n4598), .dinb(n4457), .dout(n4639));
  jand g04576(.dina(n4631), .dinb(n4453), .dout(n4640));
  jor  g04577(.dina(n4640), .dinb(n4639), .dout(n4641));
  jor  g04578(.dina(n4641), .dinb(n4638), .dout(n4642));
  jor  g04579(.dina(n4642), .dinb(n4637), .dout(n4643));
  jxor g04580(.dina(n4643), .dinb(n88), .dout(n4644));
  jnot g04581(.din(n4644), .dout(n4645));
  jxor g04582(.dina(n4553), .dinb(n4471), .dout(n4646));
  jand g04583(.dina(n4646), .dinb(n4645), .dout(n4647));
  jor  g04584(.dina(n4647), .dinb(n4554), .dout(n4648));
  jor  g04585(.dina(n4543), .dinb(n4475), .dout(n4649));
  jand g04586(.dina(n4552), .dinb(n4544), .dout(n4650));
  jnot g04587(.din(n4650), .dout(n4651));
  jand g04588(.dina(n4651), .dinb(n4649), .dout(n4652));
  jnot g04589(.din(n4652), .dout(n4653));
  jand g04590(.dina(n4446), .dinb(n732), .dout(n4654));
  jand g04591(.dina(n4451), .dinb(n3855), .dout(n4655));
  jand g04592(.dina(n4358), .dinb(n3858), .dout(n4656));
  jand g04593(.dina(n3851), .dinb(n3853), .dout(n4657));
  jor  g04594(.dina(n4657), .dinb(n4656), .dout(n4658));
  jor  g04595(.dina(n4658), .dinb(n4655), .dout(n4659));
  jor  g04596(.dina(n4659), .dinb(n4654), .dout(n4660));
  jand g04597(.dina(n988), .dinb(n377), .dout(n4661));
  jand g04598(.dina(n4661), .dinb(n340), .dout(n4662));
  jand g04599(.dina(n4662), .dinb(n1786), .dout(n4663));
  jand g04600(.dina(n2817), .dinb(n967), .dout(n4664));
  jand g04601(.dina(n4664), .dinb(n4133), .dout(n4665));
  jand g04602(.dina(n4665), .dinb(n4663), .dout(n4666));
  jnot g04603(.din(n1714), .dout(n4667));
  jand g04604(.dina(n635), .dinb(n574), .dout(n4668));
  jand g04605(.dina(n4668), .dinb(n4667), .dout(n4669));
  jand g04606(.dina(n324), .dinb(n174), .dout(n4670));
  jand g04607(.dina(n4670), .dinb(n384), .dout(n4671));
  jand g04608(.dina(n4671), .dinb(n4669), .dout(n4672));
  jand g04609(.dina(n4672), .dinb(n2895), .dout(n4673));
  jand g04610(.dina(n4673), .dinb(n3162), .dout(n4674));
  jand g04611(.dina(n4674), .dinb(n4666), .dout(n4675));
  jand g04612(.dina(n4675), .dinb(n3051), .dout(n4676));
  jand g04613(.dina(n721), .dinb(n689), .dout(n4677));
  jand g04614(.dina(n4677), .dinb(n290), .dout(n4678));
  jand g04615(.dina(n786), .dinb(n671), .dout(n4679));
  jand g04616(.dina(n757), .dinb(n499), .dout(n4680));
  jand g04617(.dina(n4680), .dinb(n4679), .dout(n4681));
  jand g04618(.dina(n4681), .dinb(n4678), .dout(n4682));
  jand g04619(.dina(n4682), .dinb(n2058), .dout(n4683));
  jand g04620(.dina(n3389), .dinb(n2564), .dout(n4684));
  jand g04621(.dina(n4684), .dinb(n827), .dout(n4685));
  jand g04622(.dina(n1924), .dinb(n1285), .dout(n4686));
  jand g04623(.dina(n4232), .dinb(n4311), .dout(n4687));
  jand g04624(.dina(n4687), .dinb(n4686), .dout(n4688));
  jand g04625(.dina(n4688), .dinb(n4685), .dout(n4689));
  jand g04626(.dina(n4689), .dinb(n4683), .dout(n4690));
  jand g04627(.dina(n893), .dinb(n532), .dout(n4691));
  jand g04628(.dina(n4691), .dinb(n82), .dout(n4692));
  jand g04629(.dina(n4692), .dinb(n369), .dout(n4693));
  jand g04630(.dina(n4693), .dinb(n3800), .dout(n4694));
  jand g04631(.dina(n1536), .dinb(n277), .dout(n4695));
  jand g04632(.dina(n1196), .dinb(n537), .dout(n4696));
  jand g04633(.dina(n4696), .dinb(n4695), .dout(n4697));
  jand g04634(.dina(n472), .dinb(n443), .dout(n4698));
  jand g04635(.dina(n4698), .dinb(n1034), .dout(n4699));
  jand g04636(.dina(n1167), .dinb(n716), .dout(n4700));
  jand g04637(.dina(n959), .dinb(n391), .dout(n4701));
  jand g04638(.dina(n4701), .dinb(n4700), .dout(n4702));
  jand g04639(.dina(n4702), .dinb(n4699), .dout(n4703));
  jand g04640(.dina(n4703), .dinb(n4697), .dout(n4704));
  jand g04641(.dina(n4704), .dinb(n4694), .dout(n4705));
  jand g04642(.dina(n1992), .dinb(n2619), .dout(n4706));
  jand g04643(.dina(n1192), .dinb(n554), .dout(n4707));
  jand g04644(.dina(n4707), .dinb(n4706), .dout(n4708));
  jand g04645(.dina(n793), .dinb(n330), .dout(n4709));
  jand g04646(.dina(n4709), .dinb(n646), .dout(n4710));
  jand g04647(.dina(n427), .dinb(n337), .dout(n4711));
  jand g04648(.dina(n1184), .dinb(n478), .dout(n4712));
  jand g04649(.dina(n4712), .dinb(n4711), .dout(n4713));
  jand g04650(.dina(n4713), .dinb(n4710), .dout(n4714));
  jand g04651(.dina(n4714), .dinb(n4708), .dout(n4715));
  jand g04652(.dina(n4715), .dinb(n1326), .dout(n4716));
  jand g04653(.dina(n4716), .dinb(n4705), .dout(n4717));
  jand g04654(.dina(n4717), .dinb(n4690), .dout(n4718));
  jand g04655(.dina(n4718), .dinb(n4676), .dout(n4719));
  jxor g04656(.dina(n4719), .dinb(n4539), .dout(n4720));
  jxor g04657(.dina(n4720), .dinb(n4660), .dout(n4721));
  jxor g04658(.dina(n4721), .dinb(n4653), .dout(n4722));
  jnot g04659(.din(n4722), .dout(n4723));
  jnot g04660(.din(n4449), .dout(n4724));
  jand g04661(.dina(n4635), .dinb(n4605), .dout(n4725));
  jnot g04662(.din(n4725), .dout(n4726));
  jand g04663(.dina(n4726), .dinb(n4630), .dout(n4727));
  jand g04664(.dina(n4726), .dinb(n4597), .dout(n4728));
  jnot g04665(.din(n4728), .dout(n4729));
  jand g04666(.dina(n4729), .dinb(n4631), .dout(n4730));
  jor  g04667(.dina(n4730), .dinb(n4727), .dout(n4731));
  jor  g04668(.dina(n4731), .dinb(n4724), .dout(n4732));
  jnot g04669(.din(n4461), .dout(n4733));
  jor  g04670(.dina(n4597), .dinb(n4733), .dout(n4734));
  jnot g04671(.din(n4457), .dout(n4735));
  jor  g04672(.dina(n4630), .dinb(n4735), .dout(n4736));
  jand g04673(.dina(n4736), .dinb(n4734), .dout(n4737));
  jand g04674(.dina(n4737), .dinb(n4732), .dout(n4738));
  jxor g04675(.dina(n4738), .dinb(\a[29] ), .dout(n4739));
  jxor g04676(.dina(n4739), .dinb(n4723), .dout(n4740));
  jxor g04677(.dina(n4740), .dinb(n4648), .dout(n4741));
  jxor g04678(.dina(\a[25] ), .dinb(\a[24] ), .dout(n4742));
  jnot g04679(.din(n4742), .dout(n4743));
  jand g04680(.dina(n4743), .dinb(n73), .dout(n4744));
  jand g04681(.dina(n4744), .dinb(n71), .dout(n4745));
  jnot g04682(.din(n4745), .dout(n4746));
  jnot g04683(.din(n75), .dout(n4747));
  jor  g04684(.dina(n4728), .dinb(n4747), .dout(n4748));
  jand g04685(.dina(n4748), .dinb(n4746), .dout(n4749));
  jor  g04686(.dina(n4749), .dinb(n4630), .dout(n4750));
  jxor g04687(.dina(n4750), .dinb(\a[26] ), .dout(n4751));
  jxor g04688(.dina(n4603), .dinb(n4602), .dout(n4752));
  jand g04689(.dina(n4752), .dinb(n4449), .dout(n4753));
  jand g04690(.dina(n4457), .dinb(n4451), .dout(n4754));
  jand g04691(.dina(n4461), .dinb(n4358), .dout(n4755));
  jand g04692(.dina(n4598), .dinb(n4453), .dout(n4756));
  jor  g04693(.dina(n4756), .dinb(n4755), .dout(n4757));
  jor  g04694(.dina(n4757), .dinb(n4754), .dout(n4758));
  jor  g04695(.dina(n4758), .dinb(n4753), .dout(n4759));
  jxor g04696(.dina(n4759), .dinb(n88), .dout(n4760));
  jor  g04697(.dina(n4760), .dinb(n4751), .dout(n4761));
  jxor g04698(.dina(n4468), .dinb(n4039), .dout(n4762));
  jxor g04699(.dina(n4760), .dinb(n4751), .dout(n4763));
  jand g04700(.dina(n4763), .dinb(n4762), .dout(n4764));
  jnot g04701(.din(n4764), .dout(n4765));
  jand g04702(.dina(n4765), .dinb(n4761), .dout(n4766));
  jnot g04703(.din(n4766), .dout(n4767));
  jxor g04704(.dina(n4646), .dinb(n4645), .dout(n4768));
  jand g04705(.dina(n4768), .dinb(n4767), .dout(n4769));
  jxor g04706(.dina(n4466), .dinb(n4280), .dout(n4770));
  jxor g04707(.dina(n4268), .dinb(n4099), .dout(n4771));
  jxor g04708(.dina(n3763), .dinb(n3762), .dout(n4772));
  jand g04709(.dina(n4772), .dinb(n732), .dout(n4773));
  jand g04710(.dina(n3855), .dinb(n1213), .dout(n4774));
  jand g04711(.dina(n3851), .dinb(n1445), .dout(n4775));
  jand g04712(.dina(n3858), .dinb(n1343), .dout(n4776));
  jor  g04713(.dina(n4776), .dinb(n4775), .dout(n4777));
  jor  g04714(.dina(n4777), .dinb(n4774), .dout(n4778));
  jor  g04715(.dina(n4778), .dinb(n4773), .dout(n4779));
  jand g04716(.dina(n4779), .dinb(n4771), .dout(n4780));
  jand g04717(.dina(n2014), .dinb(n382), .dout(n4781));
  jand g04718(.dina(n4781), .dinb(n2053), .dout(n4782));
  jand g04719(.dina(n1899), .dinb(n1353), .dout(n4783));
  jand g04720(.dina(n1991), .dinb(n752), .dout(n4784));
  jand g04721(.dina(n4784), .dinb(n4783), .dout(n4785));
  jand g04722(.dina(n4785), .dinb(n4782), .dout(n4786));
  jand g04723(.dina(n678), .dinb(n130), .dout(n4787));
  jand g04724(.dina(n4787), .dinb(n2286), .dout(n4788));
  jand g04725(.dina(n499), .dinb(n274), .dout(n4789));
  jand g04726(.dina(n4789), .dinb(n391), .dout(n4790));
  jand g04727(.dina(n4790), .dinb(n1488), .dout(n4791));
  jand g04728(.dina(n4791), .dinb(n4788), .dout(n4792));
  jand g04729(.dina(n4792), .dinb(n4786), .dout(n4793));
  jand g04730(.dina(n566), .dinb(n542), .dout(n4794));
  jand g04731(.dina(n4794), .dinb(n483), .dout(n4795));
  jnot g04732(.din(n3646), .dout(n4796));
  jand g04733(.dina(n445), .dinb(n92), .dout(n4797));
  jand g04734(.dina(n4797), .dinb(n4796), .dout(n4798));
  jand g04735(.dina(n4798), .dinb(n3108), .dout(n4799));
  jand g04736(.dina(n4799), .dinb(n4795), .dout(n4800));
  jand g04737(.dina(n770), .dinb(n214), .dout(n4801));
  jand g04738(.dina(n494), .dinb(n149), .dout(n4802));
  jand g04739(.dina(n4802), .dinb(n4801), .dout(n4803));
  jand g04740(.dina(n4803), .dinb(n829), .dout(n4804));
  jand g04741(.dina(n4804), .dinb(n1224), .dout(n4805));
  jand g04742(.dina(n4805), .dinb(n4800), .dout(n4806));
  jand g04743(.dina(n4806), .dinb(n4793), .dout(n4807));
  jand g04744(.dina(n405), .dinb(n202), .dout(n4808));
  jand g04745(.dina(n4808), .dinb(n424), .dout(n4809));
  jand g04746(.dina(n622), .dinb(n136), .dout(n4810));
  jand g04747(.dina(n701), .dinb(n386), .dout(n4811));
  jand g04748(.dina(n819), .dinb(n515), .dout(n4812));
  jand g04749(.dina(n4812), .dinb(n4811), .dout(n4813));
  jand g04750(.dina(n4813), .dinb(n4810), .dout(n4814));
  jand g04751(.dina(n4814), .dinb(n4809), .dout(n4815));
  jand g04752(.dina(n586), .dinb(n509), .dout(n4816));
  jand g04753(.dina(n4816), .dinb(n365), .dout(n4817));
  jand g04754(.dina(n4817), .dinb(n1805), .dout(n4818));
  jand g04755(.dina(n4678), .dinb(n1187), .dout(n4819));
  jand g04756(.dina(n4819), .dinb(n4818), .dout(n4820));
  jand g04757(.dina(n612), .dinb(n367), .dout(n4821));
  jand g04758(.dina(n614), .dinb(n443), .dout(n4822));
  jand g04759(.dina(n4822), .dinb(n4821), .dout(n4823));
  jand g04760(.dina(n4128), .dinb(n802), .dout(n4824));
  jand g04761(.dina(n4824), .dinb(n4823), .dout(n4825));
  jand g04762(.dina(n1663), .dinb(n697), .dout(n4826));
  jand g04763(.dina(n1474), .dinb(n253), .dout(n4827));
  jand g04764(.dina(n4827), .dinb(n4826), .dout(n4828));
  jand g04765(.dina(n4828), .dinb(n4825), .dout(n4829));
  jand g04766(.dina(n4829), .dinb(n4820), .dout(n4830));
  jand g04767(.dina(n4830), .dinb(n4815), .dout(n4831));
  jand g04768(.dina(n392), .dinb(n257), .dout(n4832));
  jand g04769(.dina(n4832), .dinb(n703), .dout(n4833));
  jand g04770(.dina(n655), .dinb(n305), .dout(n4834));
  jand g04771(.dina(n4834), .dinb(n979), .dout(n4835));
  jand g04772(.dina(n4835), .dinb(n4833), .dout(n4836));
  jand g04773(.dina(n4836), .dinb(n1852), .dout(n4837));
  jand g04774(.dina(n3865), .dinb(n717), .dout(n4838));
  jand g04775(.dina(n2025), .dinb(n1711), .dout(n4839));
  jand g04776(.dina(n4839), .dinb(n4838), .dout(n4840));
  jand g04777(.dina(n4840), .dinb(n2738), .dout(n4841));
  jand g04778(.dina(n4841), .dinb(n4837), .dout(n4842));
  jand g04779(.dina(n3008), .dinb(n1503), .dout(n4843));
  jand g04780(.dina(n4843), .dinb(n4842), .dout(n4844));
  jand g04781(.dina(n4844), .dinb(n4831), .dout(n4845));
  jand g04782(.dina(n4845), .dinb(n4807), .dout(n4846));
  jor  g04783(.dina(n4846), .dinb(n4159), .dout(n4847));
  jxor g04784(.dina(n4846), .dinb(n4159), .dout(n4848));
  jxor g04785(.dina(n3754), .dinb(n3753), .dout(n4849));
  jand g04786(.dina(n4849), .dinb(n732), .dout(n4850));
  jand g04787(.dina(n3855), .dinb(n1560), .dout(n4851));
  jand g04788(.dina(n3851), .dinb(n1776), .dout(n4852));
  jand g04789(.dina(n3858), .dinb(n1624), .dout(n4853));
  jor  g04790(.dina(n4853), .dinb(n4852), .dout(n4854));
  jor  g04791(.dina(n4854), .dinb(n4851), .dout(n4855));
  jor  g04792(.dina(n4855), .dinb(n4850), .dout(n4856));
  jand g04793(.dina(n4856), .dinb(n4848), .dout(n4857));
  jnot g04794(.din(n4857), .dout(n4858));
  jand g04795(.dina(n4858), .dinb(n4847), .dout(n4859));
  jnot g04796(.din(n4859), .dout(n4860));
  jand g04797(.dina(n4252), .dinb(n4247), .dout(n4861));
  jand g04798(.dina(n4253), .dinb(n4249), .dout(n4862));
  jor  g04799(.dina(n4862), .dinb(n4861), .dout(n4863));
  jand g04800(.dina(n4863), .dinb(n4860), .dout(n4864));
  jxor g04801(.dina(n4863), .dinb(n4860), .dout(n4865));
  jxor g04802(.dina(n3757), .dinb(n3756), .dout(n4866));
  jand g04803(.dina(n4866), .dinb(n732), .dout(n4867));
  jand g04804(.dina(n3855), .dinb(n1445), .dout(n4868));
  jand g04805(.dina(n3851), .dinb(n1624), .dout(n4869));
  jand g04806(.dina(n3858), .dinb(n1560), .dout(n4870));
  jor  g04807(.dina(n4870), .dinb(n4869), .dout(n4871));
  jor  g04808(.dina(n4871), .dinb(n4868), .dout(n4872));
  jor  g04809(.dina(n4872), .dinb(n4867), .dout(n4873));
  jand g04810(.dina(n4873), .dinb(n4865), .dout(n4874));
  jor  g04811(.dina(n4874), .dinb(n4864), .dout(n4875));
  jxor g04812(.dina(n4253), .dinb(n4095), .dout(n4876));
  jxor g04813(.dina(n4876), .dinb(n4265), .dout(n4877));
  jand g04814(.dina(n4877), .dinb(n4875), .dout(n4878));
  jnot g04815(.din(n4878), .dout(n4879));
  jxor g04816(.dina(n4877), .dinb(n4875), .dout(n4880));
  jnot g04817(.din(n4880), .dout(n4881));
  jand g04818(.dina(n4449), .dinb(n4026), .dout(n4882));
  jand g04819(.dina(n4461), .dinb(n1213), .dout(n4883));
  jand g04820(.dina(n4457), .dinb(n1076), .dout(n4884));
  jand g04821(.dina(n4453), .dinb(n922), .dout(n4885));
  jor  g04822(.dina(n4885), .dinb(n4884), .dout(n4886));
  jor  g04823(.dina(n4886), .dinb(n4883), .dout(n4887));
  jor  g04824(.dina(n4887), .dinb(n4882), .dout(n4888));
  jxor g04825(.dina(n4888), .dinb(n88), .dout(n4889));
  jor  g04826(.dina(n4889), .dinb(n4881), .dout(n4890));
  jand g04827(.dina(n4890), .dinb(n4879), .dout(n4891));
  jnot g04828(.din(n4891), .dout(n4892));
  jxor g04829(.dina(n4779), .dinb(n4771), .dout(n4893));
  jand g04830(.dina(n4893), .dinb(n4892), .dout(n4894));
  jor  g04831(.dina(n4894), .dinb(n4780), .dout(n4895));
  jnot g04832(.din(n4895), .dout(n4896));
  jxor g04833(.dina(n4272), .dinb(n4271), .dout(n4897));
  jnot g04834(.din(n4897), .dout(n4898));
  jand g04835(.dina(n4898), .dinb(n4896), .dout(n4899));
  jnot g04836(.din(n4899), .dout(n4900));
  jand g04837(.dina(n4897), .dinb(n4895), .dout(n4901));
  jnot g04838(.din(n4545), .dout(n4902));
  jor  g04839(.dina(n4902), .dinb(n4724), .dout(n4903));
  jor  g04840(.dina(n4735), .dinb(n3846), .dout(n4904));
  jnot g04841(.din(n4453), .dout(n4905));
  jor  g04842(.dina(n4905), .dinb(n4357), .dout(n4906));
  jor  g04843(.dina(n4733), .dinb(n921), .dout(n4907));
  jand g04844(.dina(n4907), .dinb(n4906), .dout(n4908));
  jand g04845(.dina(n4908), .dinb(n4904), .dout(n4909));
  jand g04846(.dina(n4909), .dinb(n4903), .dout(n4910));
  jxor g04847(.dina(n4910), .dinb(\a[29] ), .dout(n4911));
  jnot g04848(.din(n4911), .dout(n4912));
  jor  g04849(.dina(n4912), .dinb(n4901), .dout(n4913));
  jand g04850(.dina(n4913), .dinb(n4900), .dout(n4914));
  jand g04851(.dina(n4914), .dinb(n4770), .dout(n4915));
  jor  g04852(.dina(n4731), .dinb(n4747), .dout(n4916));
  jor  g04853(.dina(n4746), .dinb(n4597), .dout(n4917));
  jand g04854(.dina(n4742), .dinb(n73), .dout(n4918));
  jnot g04855(.din(n4918), .dout(n4919));
  jor  g04856(.dina(n4919), .dinb(n4630), .dout(n4920));
  jand g04857(.dina(n4920), .dinb(n4917), .dout(n4921));
  jand g04858(.dina(n4921), .dinb(n4916), .dout(n4922));
  jxor g04859(.dina(n4922), .dinb(\a[26] ), .dout(n4923));
  jnot g04860(.din(n4923), .dout(n4924));
  jxor g04861(.dina(n4914), .dinb(n4770), .dout(n4925));
  jand g04862(.dina(n4925), .dinb(n4924), .dout(n4926));
  jor  g04863(.dina(n4926), .dinb(n4915), .dout(n4927));
  jxor g04864(.dina(n4763), .dinb(n4762), .dout(n4928));
  jand g04865(.dina(n4928), .dinb(n4927), .dout(n4929));
  jand g04866(.dina(n4636), .dinb(n75), .dout(n4930));
  jand g04867(.dina(n4745), .dinb(n4451), .dout(n4931));
  jand g04868(.dina(n4918), .dinb(n4598), .dout(n4932));
  jand g04869(.dina(n74), .dinb(n70), .dout(n4933));
  jand g04870(.dina(n4933), .dinb(n4631), .dout(n4934));
  jor  g04871(.dina(n4934), .dinb(n4932), .dout(n4935));
  jor  g04872(.dina(n4935), .dinb(n4931), .dout(n4936));
  jor  g04873(.dina(n4936), .dinb(n4930), .dout(n4937));
  jxor g04874(.dina(n4937), .dinb(n68), .dout(n4938));
  jnot g04875(.din(n4938), .dout(n4939));
  jnot g04876(.din(n3848), .dout(n4940));
  jor  g04877(.dina(n4724), .dinb(n4940), .dout(n4941));
  jor  g04878(.dina(n4733), .dinb(n1075), .dout(n4942));
  jor  g04879(.dina(n4735), .dinb(n921), .dout(n4943));
  jor  g04880(.dina(n4905), .dinb(n3846), .dout(n4944));
  jand g04881(.dina(n4944), .dinb(n4943), .dout(n4945));
  jand g04882(.dina(n4945), .dinb(n4942), .dout(n4946));
  jand g04883(.dina(n4946), .dinb(n4941), .dout(n4947));
  jxor g04884(.dina(n4947), .dinb(\a[29] ), .dout(n4948));
  jxor g04885(.dina(n4893), .dinb(n4892), .dout(n4949));
  jnot g04886(.din(n4949), .dout(n4950));
  jand g04887(.dina(n4950), .dinb(n4948), .dout(n4951));
  jnot g04888(.din(n4951), .dout(n4952));
  jnot g04889(.din(n4948), .dout(n4953));
  jand g04890(.dina(n4949), .dinb(n4953), .dout(n4954));
  jnot g04891(.din(n4752), .dout(n4955));
  jor  g04892(.dina(n4955), .dinb(n4747), .dout(n4956));
  jor  g04893(.dina(n4919), .dinb(n4444), .dout(n4957));
  jor  g04894(.dina(n4746), .dinb(n4357), .dout(n4958));
  jnot g04895(.din(n4933), .dout(n4959));
  jor  g04896(.dina(n4959), .dinb(n4597), .dout(n4960));
  jand g04897(.dina(n4960), .dinb(n4958), .dout(n4961));
  jand g04898(.dina(n4961), .dinb(n4957), .dout(n4962));
  jand g04899(.dina(n4962), .dinb(n4956), .dout(n4963));
  jxor g04900(.dina(n4963), .dinb(\a[26] ), .dout(n4964));
  jnot g04901(.din(n4964), .dout(n4965));
  jor  g04902(.dina(n4965), .dinb(n4954), .dout(n4966));
  jand g04903(.dina(n4966), .dinb(n4952), .dout(n4967));
  jand g04904(.dina(n4967), .dinb(n4939), .dout(n4968));
  jnot g04905(.din(n4968), .dout(n4969));
  jxor g04906(.dina(n4967), .dinb(n4939), .dout(n4970));
  jnot g04907(.din(n4970), .dout(n4971));
  jxor g04908(.dina(n4897), .dinb(n4895), .dout(n4972));
  jxor g04909(.dina(n4972), .dinb(n4911), .dout(n4973));
  jor  g04910(.dina(n4973), .dinb(n4971), .dout(n4974));
  jand g04911(.dina(n4974), .dinb(n4969), .dout(n4975));
  jnot g04912(.din(n4975), .dout(n4976));
  jxor g04913(.dina(n4925), .dinb(n4924), .dout(n4977));
  jand g04914(.dina(n4977), .dinb(n4976), .dout(n4978));
  jxor g04915(.dina(n4973), .dinb(n4971), .dout(n4979));
  jand g04916(.dina(n4449), .dinb(n4043), .dout(n4980));
  jand g04917(.dina(n4453), .dinb(n1076), .dout(n4981));
  jand g04918(.dina(n4457), .dinb(n1213), .dout(n4982));
  jand g04919(.dina(n4461), .dinb(n1343), .dout(n4983));
  jor  g04920(.dina(n4983), .dinb(n4982), .dout(n4984));
  jor  g04921(.dina(n4984), .dinb(n4981), .dout(n4985));
  jor  g04922(.dina(n4985), .dinb(n4980), .dout(n4986));
  jxor g04923(.dina(n4986), .dinb(n88), .dout(n4987));
  jnot g04924(.din(n4987), .dout(n4988));
  jxor g04925(.dina(n4873), .dinb(n4865), .dout(n4989));
  jand g04926(.dina(n4989), .dinb(n4988), .dout(n4990));
  jxor g04927(.dina(n4856), .dinb(n4848), .dout(n4991));
  jnot g04928(.din(n4991), .dout(n4992));
  jand g04929(.dina(n3041), .dinb(n1768), .dout(n4993));
  jand g04930(.dina(n1829), .dinb(n1492), .dout(n4994));
  jand g04931(.dina(n4994), .dinb(n4993), .dout(n4995));
  jand g04932(.dina(n1040), .dinb(n499), .dout(n4996));
  jand g04933(.dina(n926), .dinb(n427), .dout(n4997));
  jand g04934(.dina(n4997), .dinb(n4996), .dout(n4998));
  jand g04935(.dina(n1144), .dinb(n243), .dout(n4999));
  jand g04936(.dina(n4999), .dinb(n1265), .dout(n5000));
  jand g04937(.dina(n5000), .dinb(n4998), .dout(n5001));
  jand g04938(.dina(n5001), .dinb(n4995), .dout(n5002));
  jand g04939(.dina(n979), .dinb(n721), .dout(n5003));
  jand g04940(.dina(n5003), .dinb(n2769), .dout(n5004));
  jand g04941(.dina(n1467), .dinb(n1411), .dout(n5005));
  jand g04942(.dina(n5005), .dinb(n5004), .dout(n5006));
  jand g04943(.dina(n5006), .dinb(n1245), .dout(n5007));
  jand g04944(.dina(n5007), .dinb(n5002), .dout(n5008));
  jand g04945(.dina(n5008), .dinb(n3080), .dout(n5009));
  jand g04946(.dina(n4294), .dinb(n3293), .dout(n5010));
  jand g04947(.dina(n5010), .dinb(n5009), .dout(n5011));
  jand g04948(.dina(n5011), .dinb(n784), .dout(n5012));
  jnot g04949(.din(n5012), .dout(n5013));
  jand g04950(.dina(n701), .dinb(n418), .dout(n5014));
  jand g04951(.dina(n1346), .dinb(n243), .dout(n5015));
  jand g04952(.dina(n5015), .dinb(n5014), .dout(n5016));
  jand g04953(.dina(n5016), .dinb(n835), .dout(n5017));
  jand g04954(.dina(n671), .dinb(n492), .dout(n5018));
  jand g04955(.dina(n5018), .dinb(n769), .dout(n5019));
  jand g04956(.dina(n5019), .dinb(n862), .dout(n5020));
  jand g04957(.dina(n5020), .dinb(n5017), .dout(n5021));
  jand g04958(.dina(n314), .dinb(n262), .dout(n5022));
  jand g04959(.dina(n5022), .dinb(n2672), .dout(n5023));
  jand g04960(.dina(n5023), .dinb(n2041), .dout(n5024));
  jand g04961(.dina(n1675), .dinb(n737), .dout(n5025));
  jand g04962(.dina(n979), .dinb(n386), .dout(n5026));
  jand g04963(.dina(n5026), .dinb(n2526), .dout(n5027));
  jand g04964(.dina(n5027), .dinb(n5025), .dout(n5028));
  jand g04965(.dina(n5028), .dinb(n5024), .dout(n5029));
  jand g04966(.dina(n1031), .dinb(n134), .dout(n5030));
  jand g04967(.dina(n595), .dinb(n367), .dout(n5031));
  jand g04968(.dina(n5031), .dinb(n5030), .dout(n5032));
  jand g04969(.dina(n721), .dinb(n304), .dout(n5033));
  jand g04970(.dina(n5033), .dinb(n2026), .dout(n5034));
  jand g04971(.dina(n5034), .dinb(n5032), .dout(n5035));
  jand g04972(.dina(n5035), .dinb(n2166), .dout(n5036));
  jand g04973(.dina(n5036), .dinb(n5029), .dout(n5037));
  jand g04974(.dina(n5037), .dinb(n5021), .dout(n5038));
  jand g04975(.dina(n311), .dinb(n214), .dout(n5039));
  jand g04976(.dina(n435), .dinb(n194), .dout(n5040));
  jand g04977(.dina(n5040), .dinb(n5039), .dout(n5041));
  jand g04978(.dina(n5041), .dinb(n1399), .dout(n5042));
  jand g04979(.dina(n1615), .dinb(n404), .dout(n5043));
  jand g04980(.dina(n5043), .dinb(n1432), .dout(n5044));
  jand g04981(.dina(n1991), .dinb(n286), .dout(n5045));
  jand g04982(.dina(n5045), .dinb(n5044), .dout(n5046));
  jand g04983(.dina(n5046), .dinb(n5042), .dout(n5047));
  jand g04984(.dina(n1924), .dinb(n1295), .dout(n5048));
  jand g04985(.dina(n4832), .dinb(n2285), .dout(n5049));
  jand g04986(.dina(n5049), .dinb(n5048), .dout(n5050));
  jand g04987(.dina(n1144), .dinb(n292), .dout(n5051));
  jand g04988(.dina(n5051), .dinb(n508), .dout(n5052));
  jand g04989(.dina(n499), .dinb(n184), .dout(n5053));
  jand g04990(.dina(n5053), .dinb(n3117), .dout(n5054));
  jand g04991(.dina(n5054), .dinb(n5052), .dout(n5055));
  jand g04992(.dina(n5055), .dinb(n5050), .dout(n5056));
  jand g04993(.dina(n5056), .dinb(n790), .dout(n5057));
  jand g04994(.dina(n5057), .dinb(n5047), .dout(n5058));
  jand g04995(.dina(n5058), .dinb(n5038), .dout(n5059));
  jand g04996(.dina(n5059), .dinb(n1127), .dout(n5060));
  jnot g04997(.din(n5060), .dout(n5061));
  jand g04998(.dina(n5061), .dinb(n5013), .dout(n5062));
  jnot g04999(.din(n5062), .dout(n5063));
  jnot g05000(.din(\a[17] ), .dout(n5064));
  jand g05001(.dina(n5060), .dinb(n5012), .dout(n5065));
  jnot g05002(.din(n5065), .dout(n5066));
  jand g05003(.dina(n5066), .dinb(n5064), .dout(n5067));
  jand g05004(.dina(n5067), .dinb(n5063), .dout(n5068));
  jnot g05005(.din(n5068), .dout(n5069));
  jand g05006(.dina(n5069), .dinb(n5063), .dout(n5070));
  jnot g05007(.din(n5070), .dout(n5071));
  jand g05008(.dina(n5071), .dinb(n4158), .dout(n5072));
  jnot g05009(.din(n5072), .dout(n5073));
  jand g05010(.dina(n5070), .dinb(n4159), .dout(n5074));
  jxor g05011(.dina(n3751), .dinb(n3750), .dout(n5075));
  jand g05012(.dina(n5075), .dinb(n732), .dout(n5076));
  jand g05013(.dina(n3855), .dinb(n1624), .dout(n5077));
  jand g05014(.dina(n3851), .dinb(n1862), .dout(n5078));
  jand g05015(.dina(n3858), .dinb(n1776), .dout(n5079));
  jor  g05016(.dina(n5079), .dinb(n5078), .dout(n5080));
  jor  g05017(.dina(n5080), .dinb(n5077), .dout(n5081));
  jor  g05018(.dina(n5081), .dinb(n5076), .dout(n5082));
  jnot g05019(.din(n5082), .dout(n5083));
  jor  g05020(.dina(n5083), .dinb(n5074), .dout(n5084));
  jand g05021(.dina(n5084), .dinb(n5073), .dout(n5085));
  jor  g05022(.dina(n5085), .dinb(n4992), .dout(n5086));
  jxor g05023(.dina(n5085), .dinb(n4992), .dout(n5087));
  jnot g05024(.din(n5087), .dout(n5088));
  jand g05025(.dina(n5069), .dinb(n5064), .dout(n5089));
  jand g05026(.dina(n5070), .dinb(n5066), .dout(n5090));
  jor  g05027(.dina(n5090), .dinb(n5089), .dout(n5091));
  jxor g05028(.dina(n3748), .dinb(n3747), .dout(n5092));
  jand g05029(.dina(n5092), .dinb(n732), .dout(n5093));
  jand g05030(.dina(n3855), .dinb(n1776), .dout(n5094));
  jand g05031(.dina(n3851), .dinb(n1956), .dout(n5095));
  jand g05032(.dina(n3858), .dinb(n1862), .dout(n5096));
  jor  g05033(.dina(n5096), .dinb(n5095), .dout(n5097));
  jor  g05034(.dina(n5097), .dinb(n5094), .dout(n5098));
  jor  g05035(.dina(n5098), .dinb(n5093), .dout(n5099));
  jand g05036(.dina(n5099), .dinb(n5091), .dout(n5100));
  jand g05037(.dina(n2888), .dinb(n2672), .dout(n5101));
  jand g05038(.dina(n3009), .dinb(n425), .dout(n5102));
  jand g05039(.dina(n5102), .dinb(n5101), .dout(n5103));
  jand g05040(.dina(n5103), .dinb(n1490), .dout(n5104));
  jand g05041(.dina(n5104), .dinb(n3147), .dout(n5105));
  jand g05042(.dina(n759), .dinb(n194), .dout(n5106));
  jand g05043(.dina(n997), .dinb(n461), .dout(n5107));
  jand g05044(.dina(n5107), .dinb(n5106), .dout(n5108));
  jand g05045(.dina(n371), .dinb(n228), .dout(n5109));
  jand g05046(.dina(n721), .dinb(n274), .dout(n5110));
  jand g05047(.dina(n5110), .dinb(n5109), .dout(n5111));
  jand g05048(.dina(n5111), .dinb(n5108), .dout(n5112));
  jand g05049(.dina(n5112), .dinb(n3467), .dout(n5113));
  jand g05050(.dina(n5113), .dinb(n3624), .dout(n5114));
  jand g05051(.dina(n5114), .dinb(n5105), .dout(n5115));
  jnot g05052(.din(n3309), .dout(n5116));
  jand g05053(.dina(n1216), .dinb(n180), .dout(n5117));
  jand g05054(.dina(n1934), .dinb(n1651), .dout(n5118));
  jand g05055(.dina(n5118), .dinb(n923), .dout(n5119));
  jand g05056(.dina(n5119), .dinb(n5117), .dout(n5120));
  jand g05057(.dina(n5120), .dinb(n5116), .dout(n5121));
  jnot g05058(.din(n3344), .dout(n5122));
  jand g05059(.dina(n694), .dinb(n431), .dout(n5123));
  jand g05060(.dina(n5123), .dinb(n5122), .dout(n5124));
  jand g05061(.dina(n505), .dinb(n136), .dout(n5125));
  jand g05062(.dina(n1346), .dinb(n655), .dout(n5126));
  jand g05063(.dina(n5126), .dinb(n5125), .dout(n5127));
  jand g05064(.dina(n230), .dinb(n177), .dout(n5128));
  jand g05065(.dina(n5128), .dinb(n1628), .dout(n5129));
  jand g05066(.dina(n5129), .dinb(n5127), .dout(n5130));
  jand g05067(.dina(n5130), .dinb(n5124), .dout(n5131));
  jand g05068(.dina(n2525), .dinb(n869), .dout(n5132));
  jand g05069(.dina(n1067), .dinb(n688), .dout(n5133));
  jand g05070(.dina(n5133), .dinb(n5132), .dout(n5134));
  jand g05071(.dina(n5134), .dinb(n2836), .dout(n5135));
  jand g05072(.dina(n5135), .dinb(n5131), .dout(n5136));
  jand g05073(.dina(n5136), .dinb(n5121), .dout(n5137));
  jand g05074(.dina(n5137), .dinb(n5115), .dout(n5138));
  jand g05075(.dina(n5138), .dinb(n4676), .dout(n5139));
  jnot g05076(.din(n5139), .dout(n5140));
  jand g05077(.dina(n5140), .dinb(n5012), .dout(n5141));
  jnot g05078(.din(n5141), .dout(n5142));
  jxor g05079(.dina(n5139), .dinb(n5013), .dout(n5143));
  jnot g05080(.din(n5143), .dout(n5144));
  jand g05081(.dina(n1323), .dinb(n870), .dout(n5145));
  jand g05082(.dina(n5145), .dinb(n2749), .dout(n5146));
  jnot g05083(.din(n3612), .dout(n5147));
  jand g05084(.dina(n5045), .dinb(n5147), .dout(n5148));
  jand g05085(.dina(n5148), .dinb(n5146), .dout(n5149));
  jand g05086(.dina(n667), .dinb(n562), .dout(n5150));
  jand g05087(.dina(n5150), .dinb(n1564), .dout(n5151));
  jand g05088(.dina(n5151), .dinb(n1942), .dout(n5152));
  jand g05089(.dina(n1066), .dinb(n533), .dout(n5153));
  jand g05090(.dina(n324), .dinb(n268), .dout(n5154));
  jand g05091(.dina(n5154), .dinb(n5153), .dout(n5155));
  jand g05092(.dina(n4679), .dinb(n1411), .dout(n5156));
  jand g05093(.dina(n5156), .dinb(n5155), .dout(n5157));
  jand g05094(.dina(n1264), .dinb(n367), .dout(n5158));
  jand g05095(.dina(n1303), .dinb(n393), .dout(n5159));
  jand g05096(.dina(n5159), .dinb(n5158), .dout(n5160));
  jand g05097(.dina(n5160), .dinb(n5157), .dout(n5161));
  jand g05098(.dina(n5161), .dinb(n5152), .dout(n5162));
  jand g05099(.dina(n5162), .dinb(n5149), .dout(n5163));
  jand g05100(.dina(n5163), .dinb(n5121), .dout(n5164));
  jand g05101(.dina(n1641), .dinb(n205), .dout(n5165));
  jand g05102(.dina(n5165), .dinb(n857), .dout(n5166));
  jand g05103(.dina(n626), .dinb(n352), .dout(n5167));
  jand g05104(.dina(n5167), .dinb(n2178), .dout(n5168));
  jand g05105(.dina(n5168), .dinb(n5166), .dout(n5169));
  jand g05106(.dina(n5169), .dinb(n4664), .dout(n5170));
  jand g05107(.dina(n619), .dinb(n130), .dout(n5171));
  jand g05108(.dina(n1519), .dinb(n252), .dout(n5172));
  jand g05109(.dina(n5172), .dinb(n5171), .dout(n5173));
  jand g05110(.dina(n5173), .dinb(n3544), .dout(n5174));
  jand g05111(.dina(n1346), .dinb(n386), .dout(n5175));
  jand g05112(.dina(n5175), .dinb(n959), .dout(n5176));
  jand g05113(.dina(n5176), .dinb(n1946), .dout(n5177));
  jand g05114(.dina(n5177), .dinb(n5174), .dout(n5178));
  jand g05115(.dina(n3470), .dinb(n1195), .dout(n5179));
  jand g05116(.dina(n5179), .dinb(n5178), .dout(n5180));
  jand g05117(.dina(n5180), .dinb(n5170), .dout(n5181));
  jand g05118(.dina(n1014), .dinb(n249), .dout(n5182));
  jand g05119(.dina(n5182), .dinb(n1090), .dout(n5183));
  jand g05120(.dina(n5183), .dinb(n2420), .dout(n5184));
  jand g05121(.dina(n4344), .dinb(n536), .dout(n5185));
  jand g05122(.dina(n553), .dinb(n445), .dout(n5186));
  jand g05123(.dina(n359), .dinb(n174), .dout(n5187));
  jand g05124(.dina(n5187), .dinb(n5186), .dout(n5188));
  jand g05125(.dina(n979), .dinb(n847), .dout(n5189));
  jand g05126(.dina(n467), .dinb(n184), .dout(n5190));
  jand g05127(.dina(n5190), .dinb(n5189), .dout(n5191));
  jand g05128(.dina(n5191), .dinb(n5188), .dout(n5192));
  jand g05129(.dina(n5192), .dinb(n5185), .dout(n5193));
  jand g05130(.dina(n5193), .dinb(n5184), .dout(n5194));
  jand g05131(.dina(n993), .dinb(n149), .dout(n5195));
  jand g05132(.dina(n5195), .dinb(n598), .dout(n5196));
  jand g05133(.dina(n3117), .dinb(n372), .dout(n5197));
  jand g05134(.dina(n413), .dinb(n92), .dout(n5198));
  jand g05135(.dina(n5198), .dinb(n788), .dout(n5199));
  jand g05136(.dina(n5199), .dinb(n5197), .dout(n5200));
  jand g05137(.dina(n5200), .dinb(n5196), .dout(n5201));
  jand g05138(.dina(n913), .dinb(n450), .dout(n5202));
  jand g05139(.dina(n304), .dinb(n214), .dout(n5203));
  jand g05140(.dina(n5203), .dinb(n5202), .dout(n5204));
  jand g05141(.dina(n869), .dinb(n861), .dout(n5205));
  jand g05142(.dina(n5205), .dinb(n5204), .dout(n5206));
  jand g05143(.dina(n483), .dinb(n120), .dout(n5207));
  jand g05144(.dina(n5207), .dinb(n924), .dout(n5208));
  jand g05145(.dina(n5208), .dinb(n2977), .dout(n5209));
  jand g05146(.dina(n5209), .dinb(n5206), .dout(n5210));
  jand g05147(.dina(n655), .dinb(n443), .dout(n5211));
  jand g05148(.dina(n736), .dinb(n516), .dout(n5212));
  jand g05149(.dina(n5212), .dinb(n5211), .dout(n5213));
  jand g05150(.dina(n5213), .dinb(n798), .dout(n5214));
  jand g05151(.dina(n5214), .dinb(n4149), .dout(n5215));
  jand g05152(.dina(n5215), .dinb(n5210), .dout(n5216));
  jand g05153(.dina(n5216), .dinb(n5201), .dout(n5217));
  jand g05154(.dina(n5217), .dinb(n5194), .dout(n5218));
  jand g05155(.dina(n5218), .dinb(n5181), .dout(n5219));
  jand g05156(.dina(n5219), .dinb(n5164), .dout(n5220));
  jnot g05157(.din(n5220), .dout(n5221));
  jand g05158(.dina(n4514), .dinb(n1830), .dout(n5222));
  jand g05159(.dina(n5222), .dinb(n3074), .dout(n5223));
  jand g05160(.dina(n703), .dinb(n157), .dout(n5224));
  jand g05161(.dina(n5224), .dinb(n417), .dout(n5225));
  jand g05162(.dina(n3595), .dinb(n927), .dout(n5226));
  jand g05163(.dina(n5226), .dinb(n5225), .dout(n5227));
  jand g05164(.dina(n5227), .dinb(n5044), .dout(n5228));
  jand g05165(.dina(n5228), .dinb(n5223), .dout(n5229));
  jand g05166(.dina(n759), .dinb(n508), .dout(n5230));
  jand g05167(.dina(n5230), .dinb(n2151), .dout(n5231));
  jand g05168(.dina(n5231), .dinb(n258), .dout(n5232));
  jand g05169(.dina(n675), .dinb(n286), .dout(n5233));
  jand g05170(.dina(n707), .dinb(n476), .dout(n5234));
  jand g05171(.dina(n5234), .dinb(n5233), .dout(n5235));
  jand g05172(.dina(n2401), .dinb(n1154), .dout(n5236));
  jand g05173(.dina(n5236), .dinb(n5235), .dout(n5237));
  jand g05174(.dina(n5237), .dinb(n5124), .dout(n5238));
  jand g05175(.dina(n5238), .dinb(n5232), .dout(n5239));
  jand g05176(.dina(n5239), .dinb(n905), .dout(n5240));
  jand g05177(.dina(n5240), .dinb(n5229), .dout(n5241));
  jand g05178(.dina(n395), .dinb(n372), .dout(n5242));
  jand g05179(.dina(n635), .dinb(n500), .dout(n5243));
  jand g05180(.dina(n5243), .dinb(n5242), .dout(n5244));
  jand g05181(.dina(n857), .dinb(n763), .dout(n5245));
  jand g05182(.dina(n5245), .dinb(n1761), .dout(n5246));
  jand g05183(.dina(n5246), .dinb(n5244), .dout(n5247));
  jand g05184(.dina(n2261), .dinb(n198), .dout(n5248));
  jand g05185(.dina(n979), .dinb(n284), .dout(n5249));
  jand g05186(.dina(n542), .dinb(n154), .dout(n5250));
  jand g05187(.dina(n5250), .dinb(n5249), .dout(n5251));
  jand g05188(.dina(n5251), .dinb(n5248), .dout(n5252));
  jand g05189(.dina(n5252), .dinb(n5247), .dout(n5253));
  jand g05190(.dina(n1145), .dinb(n880), .dout(n5254));
  jand g05191(.dina(n5254), .dinb(n218), .dout(n5255));
  jand g05192(.dina(n5255), .dinb(n4825), .dout(n5256));
  jand g05193(.dina(n5256), .dinb(n3157), .dout(n5257));
  jand g05194(.dina(n5257), .dinb(n5253), .dout(n5258));
  jand g05195(.dina(n778), .dinb(n607), .dout(n5259));
  jand g05196(.dina(n5259), .dinb(n1924), .dout(n5260));
  jand g05197(.dina(n5260), .dinb(n2935), .dout(n5261));
  jand g05198(.dina(n641), .dinb(n329), .dout(n5262));
  jand g05199(.dina(n756), .dinb(n678), .dout(n5263));
  jand g05200(.dina(n5263), .dinb(n5262), .dout(n5264));
  jand g05201(.dina(n5264), .dinb(n2048), .dout(n5265));
  jand g05202(.dina(n5265), .dinb(n3134), .dout(n5266));
  jand g05203(.dina(n5266), .dinb(n5261), .dout(n5267));
  jand g05204(.dina(n751), .dinb(n424), .dout(n5268));
  jand g05205(.dina(n366), .dinb(n165), .dout(n5269));
  jand g05206(.dina(n5269), .dinb(n262), .dout(n5270));
  jand g05207(.dina(n5270), .dinb(n5268), .dout(n5271));
  jand g05208(.dina(n5271), .dinb(n2508), .dout(n5272));
  jand g05209(.dina(n967), .dinb(n494), .dout(n5273));
  jand g05210(.dina(n5273), .dinb(n392), .dout(n5274));
  jand g05211(.dina(n5274), .dinb(n834), .dout(n5275));
  jand g05212(.dina(n5275), .dinb(n1873), .dout(n5276));
  jand g05213(.dina(n2580), .dinb(n1424), .dout(n5277));
  jand g05214(.dina(n5277), .dinb(n2834), .dout(n5278));
  jand g05215(.dina(n428), .dinb(n290), .dout(n5279));
  jand g05216(.dina(n5279), .dinb(n2659), .dout(n5280));
  jand g05217(.dina(n3662), .dinb(n2222), .dout(n5281));
  jand g05218(.dina(n5281), .dinb(n5280), .dout(n5282));
  jand g05219(.dina(n5282), .dinb(n5278), .dout(n5283));
  jand g05220(.dina(n5283), .dinb(n5276), .dout(n5284));
  jand g05221(.dina(n5284), .dinb(n5272), .dout(n5285));
  jand g05222(.dina(n5285), .dinb(n5267), .dout(n5286));
  jand g05223(.dina(n5286), .dinb(n5258), .dout(n5287));
  jand g05224(.dina(n5287), .dinb(n5241), .dout(n5288));
  jnot g05225(.din(n5288), .dout(n5289));
  jand g05226(.dina(n5289), .dinb(n5221), .dout(n5290));
  jnot g05227(.din(n5290), .dout(n5291));
  jnot g05228(.din(\a[14] ), .dout(n5292));
  jand g05229(.dina(n5288), .dinb(n5220), .dout(n5293));
  jnot g05230(.din(n5293), .dout(n5294));
  jand g05231(.dina(n5294), .dinb(n5292), .dout(n5295));
  jand g05232(.dina(n5295), .dinb(n5291), .dout(n5296));
  jnot g05233(.din(n5296), .dout(n5297));
  jand g05234(.dina(n5297), .dinb(n5291), .dout(n5298));
  jnot g05235(.din(n5298), .dout(n5299));
  jand g05236(.dina(n5299), .dinb(n5139), .dout(n5300));
  jnot g05237(.din(n5300), .dout(n5301));
  jand g05238(.dina(n5298), .dinb(n5140), .dout(n5302));
  jxor g05239(.dina(n3742), .dinb(n3741), .dout(n5303));
  jand g05240(.dina(n5303), .dinb(n732), .dout(n5304));
  jand g05241(.dina(n3851), .dinb(n2128), .dout(n5305));
  jand g05242(.dina(n3855), .dinb(n1956), .dout(n5306));
  jand g05243(.dina(n3858), .dinb(n2067), .dout(n5307));
  jor  g05244(.dina(n5307), .dinb(n5306), .dout(n5308));
  jor  g05245(.dina(n5308), .dinb(n5305), .dout(n5309));
  jor  g05246(.dina(n5309), .dinb(n5304), .dout(n5310));
  jnot g05247(.din(n5310), .dout(n5311));
  jor  g05248(.dina(n5311), .dinb(n5302), .dout(n5312));
  jand g05249(.dina(n5312), .dinb(n5301), .dout(n5313));
  jor  g05250(.dina(n5313), .dinb(n5144), .dout(n5314));
  jand g05251(.dina(n5314), .dinb(n5142), .dout(n5315));
  jnot g05252(.din(n5315), .dout(n5316));
  jxor g05253(.dina(n5099), .dinb(n5091), .dout(n5317));
  jand g05254(.dina(n5317), .dinb(n5316), .dout(n5318));
  jor  g05255(.dina(n5318), .dinb(n5100), .dout(n5319));
  jxor g05256(.dina(n5070), .dinb(n4159), .dout(n5320));
  jxor g05257(.dina(n5320), .dinb(n5082), .dout(n5321));
  jand g05258(.dina(n5321), .dinb(n5319), .dout(n5322));
  jnot g05259(.din(n5322), .dout(n5323));
  jxor g05260(.dina(n5321), .dinb(n5319), .dout(n5324));
  jnot g05261(.din(n5324), .dout(n5325));
  jand g05262(.dina(n4449), .dinb(n4258), .dout(n5326));
  jand g05263(.dina(n4457), .dinb(n1445), .dout(n5327));
  jand g05264(.dina(n4461), .dinb(n1560), .dout(n5328));
  jand g05265(.dina(n4453), .dinb(n1343), .dout(n5329));
  jor  g05266(.dina(n5329), .dinb(n5328), .dout(n5330));
  jor  g05267(.dina(n5330), .dinb(n5327), .dout(n5331));
  jor  g05268(.dina(n5331), .dinb(n5326), .dout(n5332));
  jxor g05269(.dina(n5332), .dinb(n88), .dout(n5333));
  jor  g05270(.dina(n5333), .dinb(n5325), .dout(n5334));
  jand g05271(.dina(n5334), .dinb(n5323), .dout(n5335));
  jor  g05272(.dina(n5335), .dinb(n5088), .dout(n5336));
  jand g05273(.dina(n5336), .dinb(n5086), .dout(n5337));
  jnot g05274(.din(n5337), .dout(n5338));
  jxor g05275(.dina(n4989), .dinb(n4988), .dout(n5339));
  jand g05276(.dina(n5339), .dinb(n5338), .dout(n5340));
  jor  g05277(.dina(n5340), .dinb(n4990), .dout(n5341));
  jxor g05278(.dina(n4889), .dinb(n4881), .dout(n5342));
  jand g05279(.dina(n5342), .dinb(n5341), .dout(n5343));
  jand g05280(.dina(n4446), .dinb(n75), .dout(n5344));
  jand g05281(.dina(n4933), .dinb(n4451), .dout(n5345));
  jand g05282(.dina(n4918), .dinb(n4358), .dout(n5346));
  jand g05283(.dina(n4745), .dinb(n3853), .dout(n5347));
  jor  g05284(.dina(n5347), .dinb(n5346), .dout(n5348));
  jor  g05285(.dina(n5348), .dinb(n5345), .dout(n5349));
  jor  g05286(.dina(n5349), .dinb(n5344), .dout(n5350));
  jxor g05287(.dina(n5350), .dinb(n68), .dout(n5351));
  jnot g05288(.din(n5351), .dout(n5352));
  jxor g05289(.dina(n5342), .dinb(n5341), .dout(n5353));
  jand g05290(.dina(n5353), .dinb(n5352), .dout(n5354));
  jor  g05291(.dina(n5354), .dinb(n5343), .dout(n5355));
  jnot g05292(.din(n5355), .dout(n5356));
  jxor g05293(.dina(\a[23] ), .dinb(\a[22] ), .dout(n5357));
  jxor g05294(.dina(\a[21] ), .dinb(\a[20] ), .dout(n5358));
  jnot g05295(.din(n5358), .dout(n5359));
  jxor g05296(.dina(\a[22] ), .dinb(\a[21] ), .dout(n5360));
  jnot g05297(.din(n5360), .dout(n5361));
  jand g05298(.dina(n5361), .dinb(n5359), .dout(n5362));
  jand g05299(.dina(n5362), .dinb(n5357), .dout(n5363));
  jnot g05300(.din(n5363), .dout(n5364));
  jand g05301(.dina(n5358), .dinb(n5357), .dout(n5365));
  jnot g05302(.din(n5365), .dout(n5366));
  jor  g05303(.dina(n5366), .dinb(n4728), .dout(n5367));
  jand g05304(.dina(n5367), .dinb(n5364), .dout(n5368));
  jor  g05305(.dina(n5368), .dinb(n4630), .dout(n5369));
  jxor g05306(.dina(n5369), .dinb(\a[23] ), .dout(n5370));
  jand g05307(.dina(n5370), .dinb(n5356), .dout(n5371));
  jor  g05308(.dina(n5370), .dinb(n5356), .dout(n5372));
  jxor g05309(.dina(n4949), .dinb(n4953), .dout(n5373));
  jxor g05310(.dina(n5373), .dinb(n4964), .dout(n5374));
  jand g05311(.dina(n5374), .dinb(n5372), .dout(n5375));
  jor  g05312(.dina(n5375), .dinb(n5371), .dout(n5376));
  jnot g05313(.din(n5376), .dout(n5377));
  jand g05314(.dina(n5377), .dinb(n4979), .dout(n5378));
  jxor g05315(.dina(n5339), .dinb(n5338), .dout(n5379));
  jnot g05316(.din(n5379), .dout(n5380));
  jand g05317(.dina(n4545), .dinb(n75), .dout(n5381));
  jand g05318(.dina(n4745), .dinb(n922), .dout(n5382));
  jand g05319(.dina(n4918), .dinb(n3853), .dout(n5383));
  jand g05320(.dina(n4933), .dinb(n4358), .dout(n5384));
  jor  g05321(.dina(n5384), .dinb(n5383), .dout(n5385));
  jor  g05322(.dina(n5385), .dinb(n5382), .dout(n5386));
  jor  g05323(.dina(n5386), .dinb(n5381), .dout(n5387));
  jxor g05324(.dina(n5387), .dinb(n68), .dout(n5388));
  jor  g05325(.dina(n5388), .dinb(n5380), .dout(n5389));
  jxor g05326(.dina(n5335), .dinb(n5088), .dout(n5390));
  jnot g05327(.din(n5390), .dout(n5391));
  jand g05328(.dina(n4772), .dinb(n4449), .dout(n5392));
  jand g05329(.dina(n4457), .dinb(n1343), .dout(n5393));
  jand g05330(.dina(n4461), .dinb(n1445), .dout(n5394));
  jand g05331(.dina(n4453), .dinb(n1213), .dout(n5395));
  jor  g05332(.dina(n5395), .dinb(n5394), .dout(n5396));
  jor  g05333(.dina(n5396), .dinb(n5393), .dout(n5397));
  jor  g05334(.dina(n5397), .dinb(n5392), .dout(n5398));
  jxor g05335(.dina(n5398), .dinb(n88), .dout(n5399));
  jor  g05336(.dina(n5399), .dinb(n5391), .dout(n5400));
  jand g05337(.dina(n3848), .dinb(n75), .dout(n5401));
  jand g05338(.dina(n4918), .dinb(n922), .dout(n5402));
  jand g05339(.dina(n4933), .dinb(n3853), .dout(n5403));
  jand g05340(.dina(n4745), .dinb(n1076), .dout(n5404));
  jor  g05341(.dina(n5404), .dinb(n5403), .dout(n5405));
  jor  g05342(.dina(n5405), .dinb(n5402), .dout(n5406));
  jor  g05343(.dina(n5406), .dinb(n5401), .dout(n5407));
  jxor g05344(.dina(n5407), .dinb(n68), .dout(n5408));
  jnot g05345(.din(n5408), .dout(n5409));
  jxor g05346(.dina(n5399), .dinb(n5391), .dout(n5410));
  jand g05347(.dina(n5410), .dinb(n5409), .dout(n5411));
  jnot g05348(.din(n5411), .dout(n5412));
  jand g05349(.dina(n5412), .dinb(n5400), .dout(n5413));
  jnot g05350(.din(n5413), .dout(n5414));
  jxor g05351(.dina(n5388), .dinb(n5380), .dout(n5415));
  jand g05352(.dina(n5415), .dinb(n5414), .dout(n5416));
  jnot g05353(.din(n5416), .dout(n5417));
  jand g05354(.dina(n5417), .dinb(n5389), .dout(n5418));
  jnot g05355(.din(n5418), .dout(n5419));
  jxor g05356(.dina(n5353), .dinb(n5352), .dout(n5420));
  jand g05357(.dina(n5420), .dinb(n5419), .dout(n5421));
  jor  g05358(.dina(n5366), .dinb(n4731), .dout(n5422));
  jor  g05359(.dina(n5364), .dinb(n4597), .dout(n5423));
  jand g05360(.dina(n5360), .dinb(n5359), .dout(n5424));
  jnot g05361(.din(n5424), .dout(n5425));
  jor  g05362(.dina(n5425), .dinb(n4630), .dout(n5426));
  jand g05363(.dina(n5426), .dinb(n5423), .dout(n5427));
  jand g05364(.dina(n5427), .dinb(n5422), .dout(n5428));
  jxor g05365(.dina(n5428), .dinb(\a[23] ), .dout(n5429));
  jnot g05366(.din(n5429), .dout(n5430));
  jxor g05367(.dina(n5420), .dinb(n5419), .dout(n5431));
  jand g05368(.dina(n5431), .dinb(n5430), .dout(n5432));
  jor  g05369(.dina(n5432), .dinb(n5421), .dout(n5433));
  jxor g05370(.dina(n5370), .dinb(n5356), .dout(n5434));
  jxor g05371(.dina(n5434), .dinb(n5374), .dout(n5435));
  jnot g05372(.din(n5435), .dout(n5436));
  jand g05373(.dina(n5436), .dinb(n5433), .dout(n5437));
  jxor g05374(.dina(n5436), .dinb(n5433), .dout(n5438));
  jxor g05375(.dina(n5313), .dinb(n5144), .dout(n5439));
  jxor g05376(.dina(n3745), .dinb(n3744), .dout(n5440));
  jand g05377(.dina(n5440), .dinb(n732), .dout(n5441));
  jand g05378(.dina(n3851), .dinb(n2067), .dout(n5442));
  jand g05379(.dina(n3855), .dinb(n1862), .dout(n5443));
  jand g05380(.dina(n3858), .dinb(n1956), .dout(n5444));
  jor  g05381(.dina(n5444), .dinb(n5443), .dout(n5445));
  jor  g05382(.dina(n5445), .dinb(n5442), .dout(n5446));
  jor  g05383(.dina(n5446), .dinb(n5441), .dout(n5447));
  jand g05384(.dina(n5447), .dinb(n5439), .dout(n5448));
  jand g05385(.dina(n4849), .dinb(n4449), .dout(n5449));
  jand g05386(.dina(n4453), .dinb(n1560), .dout(n5450));
  jand g05387(.dina(n4457), .dinb(n1624), .dout(n5451));
  jand g05388(.dina(n4461), .dinb(n1776), .dout(n5452));
  jor  g05389(.dina(n5452), .dinb(n5451), .dout(n5453));
  jor  g05390(.dina(n5453), .dinb(n5450), .dout(n5454));
  jor  g05391(.dina(n5454), .dinb(n5449), .dout(n5455));
  jxor g05392(.dina(n5455), .dinb(n88), .dout(n5456));
  jnot g05393(.din(n5456), .dout(n5457));
  jxor g05394(.dina(n5447), .dinb(n5439), .dout(n5458));
  jand g05395(.dina(n5458), .dinb(n5457), .dout(n5459));
  jor  g05396(.dina(n5459), .dinb(n5448), .dout(n5460));
  jxor g05397(.dina(n5317), .dinb(n5316), .dout(n5461));
  jand g05398(.dina(n5461), .dinb(n5460), .dout(n5462));
  jand g05399(.dina(n4866), .dinb(n4449), .dout(n5463));
  jand g05400(.dina(n4453), .dinb(n1445), .dout(n5464));
  jand g05401(.dina(n4457), .dinb(n1560), .dout(n5465));
  jand g05402(.dina(n4461), .dinb(n1624), .dout(n5466));
  jor  g05403(.dina(n5466), .dinb(n5465), .dout(n5467));
  jor  g05404(.dina(n5467), .dinb(n5464), .dout(n5468));
  jor  g05405(.dina(n5468), .dinb(n5463), .dout(n5469));
  jxor g05406(.dina(n5469), .dinb(n88), .dout(n5470));
  jnot g05407(.din(n5470), .dout(n5471));
  jxor g05408(.dina(n5461), .dinb(n5460), .dout(n5472));
  jand g05409(.dina(n5472), .dinb(n5471), .dout(n5473));
  jor  g05410(.dina(n5473), .dinb(n5462), .dout(n5474));
  jxor g05411(.dina(n5333), .dinb(n5325), .dout(n5475));
  jand g05412(.dina(n5475), .dinb(n5474), .dout(n5476));
  jnot g05413(.din(n5476), .dout(n5477));
  jxor g05414(.dina(n5475), .dinb(n5474), .dout(n5478));
  jnot g05415(.din(n5478), .dout(n5479));
  jand g05416(.dina(n4026), .dinb(n75), .dout(n5480));
  jand g05417(.dina(n4918), .dinb(n1076), .dout(n5481));
  jand g05418(.dina(n4933), .dinb(n922), .dout(n5482));
  jand g05419(.dina(n4745), .dinb(n1213), .dout(n5483));
  jor  g05420(.dina(n5483), .dinb(n5482), .dout(n5484));
  jor  g05421(.dina(n5484), .dinb(n5481), .dout(n5485));
  jor  g05422(.dina(n5485), .dinb(n5480), .dout(n5486));
  jxor g05423(.dina(n5486), .dinb(n68), .dout(n5487));
  jor  g05424(.dina(n5487), .dinb(n5479), .dout(n5488));
  jand g05425(.dina(n5488), .dinb(n5477), .dout(n5489));
  jnot g05426(.din(n5489), .dout(n5490));
  jxor g05427(.dina(n5410), .dinb(n5409), .dout(n5491));
  jand g05428(.dina(n5491), .dinb(n5490), .dout(n5492));
  jnot g05429(.din(n5492), .dout(n5493));
  jxor g05430(.dina(n5491), .dinb(n5490), .dout(n5494));
  jnot g05431(.din(n5494), .dout(n5495));
  jand g05432(.dina(n5365), .dinb(n4752), .dout(n5496));
  jand g05433(.dina(n5424), .dinb(n4451), .dout(n5497));
  jand g05434(.dina(n5363), .dinb(n4358), .dout(n5498));
  jor  g05435(.dina(n5359), .dinb(n5357), .dout(n5499));
  jnot g05436(.din(n5499), .dout(n5500));
  jand g05437(.dina(n5500), .dinb(n4598), .dout(n5501));
  jor  g05438(.dina(n5501), .dinb(n5498), .dout(n5502));
  jor  g05439(.dina(n5502), .dinb(n5497), .dout(n5503));
  jor  g05440(.dina(n5503), .dinb(n5496), .dout(n5504));
  jxor g05441(.dina(n5504), .dinb(n72), .dout(n5505));
  jor  g05442(.dina(n5505), .dinb(n5495), .dout(n5506));
  jand g05443(.dina(n5506), .dinb(n5493), .dout(n5507));
  jand g05444(.dina(n5365), .dinb(n4636), .dout(n5508));
  jand g05445(.dina(n5363), .dinb(n4451), .dout(n5509));
  jand g05446(.dina(n5424), .dinb(n4598), .dout(n5510));
  jand g05447(.dina(n5500), .dinb(n4631), .dout(n5511));
  jor  g05448(.dina(n5511), .dinb(n5510), .dout(n5512));
  jor  g05449(.dina(n5512), .dinb(n5509), .dout(n5513));
  jor  g05450(.dina(n5513), .dinb(n5508), .dout(n5514));
  jxor g05451(.dina(n5514), .dinb(n72), .dout(n5515));
  jor  g05452(.dina(n5515), .dinb(n5507), .dout(n5516));
  jxor g05453(.dina(n5515), .dinb(n5507), .dout(n5517));
  jxor g05454(.dina(n5415), .dinb(n5414), .dout(n5518));
  jand g05455(.dina(n5518), .dinb(n5517), .dout(n5519));
  jnot g05456(.din(n5519), .dout(n5520));
  jand g05457(.dina(n5520), .dinb(n5516), .dout(n5521));
  jnot g05458(.din(n5521), .dout(n5522));
  jxor g05459(.dina(n5431), .dinb(n5430), .dout(n5523));
  jand g05460(.dina(n5523), .dinb(n5522), .dout(n5524));
  jand g05461(.dina(n4043), .dinb(n75), .dout(n5525));
  jand g05462(.dina(n4918), .dinb(n1213), .dout(n5526));
  jand g05463(.dina(n4745), .dinb(n1343), .dout(n5527));
  jand g05464(.dina(n4933), .dinb(n1076), .dout(n5528));
  jor  g05465(.dina(n5528), .dinb(n5527), .dout(n5529));
  jor  g05466(.dina(n5529), .dinb(n5526), .dout(n5530));
  jor  g05467(.dina(n5530), .dinb(n5525), .dout(n5531));
  jxor g05468(.dina(n5531), .dinb(n68), .dout(n5532));
  jnot g05469(.din(n5532), .dout(n5533));
  jxor g05470(.dina(n5472), .dinb(n5471), .dout(n5534));
  jand g05471(.dina(n5534), .dinb(n5533), .dout(n5535));
  jand g05472(.dina(n913), .dinb(n842), .dout(n5536));
  jand g05473(.dina(n619), .dinb(n532), .dout(n5537));
  jand g05474(.dina(n5537), .dinb(n646), .dout(n5538));
  jand g05475(.dina(n5538), .dinb(n5536), .dout(n5539));
  jand g05476(.dina(n749), .dinb(n715), .dout(n5540));
  jand g05477(.dina(n5540), .dinb(n874), .dout(n5541));
  jand g05478(.dina(n926), .dinb(n509), .dout(n5542));
  jand g05479(.dina(n5542), .dinb(n2564), .dout(n5543));
  jand g05480(.dina(n5543), .dinb(n5541), .dout(n5544));
  jnot g05481(.din(n3666), .dout(n5545));
  jand g05482(.dina(n5545), .dinb(n3431), .dout(n5546));
  jand g05483(.dina(n5546), .dinb(n5544), .dout(n5547));
  jand g05484(.dina(n5547), .dinb(n5539), .dout(n5548));
  jand g05485(.dina(n694), .dinb(n317), .dout(n5549));
  jand g05486(.dina(n5549), .dinb(n1474), .dout(n5550));
  jand g05487(.dina(n1184), .dinb(n82), .dout(n5551));
  jand g05488(.dina(n5551), .dinb(n635), .dout(n5552));
  jand g05489(.dina(n5552), .dinb(n991), .dout(n5553));
  jand g05490(.dina(n5553), .dinb(n5550), .dout(n5554));
  jand g05491(.dina(n404), .dinb(n396), .dout(n5555));
  jand g05492(.dina(n445), .dinb(n330), .dout(n5556));
  jand g05493(.dina(n5556), .dinb(n5555), .dout(n5557));
  jand g05494(.dina(n4078), .dinb(n1680), .dout(n5558));
  jand g05495(.dina(n5558), .dinb(n5557), .dout(n5559));
  jand g05496(.dina(n675), .dinb(n190), .dout(n5560));
  jand g05497(.dina(n1178), .dinb(n462), .dout(n5561));
  jand g05498(.dina(n5561), .dinb(n5560), .dout(n5562));
  jand g05499(.dina(n4231), .dinb(n1135), .dout(n5563));
  jand g05500(.dina(n5563), .dinb(n5562), .dout(n5564));
  jand g05501(.dina(n5564), .dinb(n2799), .dout(n5565));
  jand g05502(.dina(n5565), .dinb(n5559), .dout(n5566));
  jand g05503(.dina(n5566), .dinb(n5554), .dout(n5567));
  jand g05504(.dina(n5567), .dinb(n5548), .dout(n5568));
  jand g05505(.dina(n4514), .dinb(n2583), .dout(n5569));
  jand g05506(.dina(n5569), .dinb(n443), .dout(n5570));
  jand g05507(.dina(n1840), .dinb(n1422), .dout(n5571));
  jand g05508(.dina(n5571), .dinb(n2255), .dout(n5572));
  jand g05509(.dina(n1014), .dinb(n622), .dout(n5573));
  jand g05510(.dina(n5573), .dinb(n429), .dout(n5574));
  jand g05511(.dina(n5574), .dinb(n4111), .dout(n5575));
  jand g05512(.dina(n5575), .dinb(n5572), .dout(n5576));
  jand g05513(.dina(n5576), .dinb(n5570), .dout(n5577));
  jand g05514(.dina(n270), .dinb(n238), .dout(n5578));
  jand g05515(.dina(n492), .dinb(n146), .dout(n5579));
  jand g05516(.dina(n5579), .dinb(n5578), .dout(n5580));
  jand g05517(.dina(n5580), .dinb(n1233), .dout(n5581));
  jand g05518(.dina(n5581), .dinb(n4502), .dout(n5582));
  jand g05519(.dina(n5582), .dinb(n666), .dout(n5583));
  jand g05520(.dina(n5583), .dinb(n5577), .dout(n5584));
  jand g05521(.dina(n5003), .dinb(n2606), .dout(n5585));
  jand g05522(.dina(n3865), .dinb(n442), .dout(n5586));
  jand g05523(.dina(n5586), .dinb(n5585), .dout(n5587));
  jand g05524(.dina(n1519), .dinb(n194), .dout(n5588));
  jand g05525(.dina(n5588), .dinb(n1079), .dout(n5589));
  jand g05526(.dina(n1615), .dinb(n687), .dout(n5590));
  jand g05527(.dina(n700), .dinb(n417), .dout(n5591));
  jand g05528(.dina(n5591), .dinb(n5590), .dout(n5592));
  jand g05529(.dina(n5592), .dinb(n5589), .dout(n5593));
  jand g05530(.dina(n5593), .dinb(n5587), .dout(n5594));
  jand g05531(.dina(n1364), .dinb(n180), .dout(n5595));
  jand g05532(.dina(n5595), .dinb(n1305), .dout(n5596));
  jand g05533(.dina(n1847), .dinb(n606), .dout(n5597));
  jand g05534(.dina(n3445), .dinb(n769), .dout(n5598));
  jand g05535(.dina(n5598), .dinb(n5597), .dout(n5599));
  jand g05536(.dina(n5599), .dinb(n1352), .dout(n5600));
  jand g05537(.dina(n5600), .dinb(n5596), .dout(n5601));
  jand g05538(.dina(n5601), .dinb(n5594), .dout(n5602));
  jand g05539(.dina(n5602), .dinb(n5584), .dout(n5603));
  jand g05540(.dina(n5603), .dinb(n5568), .dout(n5604));
  jor  g05541(.dina(n5604), .dinb(n5221), .dout(n5605));
  jxor g05542(.dina(n5604), .dinb(n5221), .dout(n5606));
  jxor g05543(.dina(n3736), .dinb(n3735), .dout(n5607));
  jand g05544(.dina(n5607), .dinb(n732), .dout(n5608));
  jand g05545(.dina(n3858), .dinb(n2237), .dout(n5609));
  jand g05546(.dina(n3851), .dinb(n2343), .dout(n5610));
  jand g05547(.dina(n3855), .dinb(n2128), .dout(n5611));
  jor  g05548(.dina(n5611), .dinb(n5610), .dout(n5612));
  jor  g05549(.dina(n5612), .dinb(n5609), .dout(n5613));
  jor  g05550(.dina(n5613), .dinb(n5608), .dout(n5614));
  jand g05551(.dina(n5614), .dinb(n5606), .dout(n5615));
  jnot g05552(.din(n5615), .dout(n5616));
  jand g05553(.dina(n5616), .dinb(n5605), .dout(n5617));
  jnot g05554(.din(n5617), .dout(n5618));
  jand g05555(.dina(n5297), .dinb(n5292), .dout(n5619));
  jand g05556(.dina(n5298), .dinb(n5294), .dout(n5620));
  jor  g05557(.dina(n5620), .dinb(n5619), .dout(n5621));
  jand g05558(.dina(n5621), .dinb(n5618), .dout(n5622));
  jxor g05559(.dina(n5621), .dinb(n5618), .dout(n5623));
  jxor g05560(.dina(n3739), .dinb(n3738), .dout(n5624));
  jand g05561(.dina(n5624), .dinb(n732), .dout(n5625));
  jand g05562(.dina(n3851), .dinb(n2237), .dout(n5626));
  jand g05563(.dina(n3858), .dinb(n2128), .dout(n5627));
  jand g05564(.dina(n3855), .dinb(n2067), .dout(n5628));
  jor  g05565(.dina(n5628), .dinb(n5627), .dout(n5629));
  jor  g05566(.dina(n5629), .dinb(n5626), .dout(n5630));
  jor  g05567(.dina(n5630), .dinb(n5625), .dout(n5631));
  jand g05568(.dina(n5631), .dinb(n5623), .dout(n5632));
  jor  g05569(.dina(n5632), .dinb(n5622), .dout(n5633));
  jxor g05570(.dina(n5298), .dinb(n5140), .dout(n5634));
  jxor g05571(.dina(n5634), .dinb(n5310), .dout(n5635));
  jand g05572(.dina(n5635), .dinb(n5633), .dout(n5636));
  jnot g05573(.din(n5636), .dout(n5637));
  jxor g05574(.dina(n5635), .dinb(n5633), .dout(n5638));
  jnot g05575(.din(n5638), .dout(n5639));
  jand g05576(.dina(n5075), .dinb(n4449), .dout(n5640));
  jand g05577(.dina(n4457), .dinb(n1776), .dout(n5641));
  jand g05578(.dina(n4461), .dinb(n1862), .dout(n5642));
  jand g05579(.dina(n4453), .dinb(n1624), .dout(n5643));
  jor  g05580(.dina(n5643), .dinb(n5642), .dout(n5644));
  jor  g05581(.dina(n5644), .dinb(n5641), .dout(n5645));
  jor  g05582(.dina(n5645), .dinb(n5640), .dout(n5646));
  jxor g05583(.dina(n5646), .dinb(n88), .dout(n5647));
  jor  g05584(.dina(n5647), .dinb(n5639), .dout(n5648));
  jand g05585(.dina(n5648), .dinb(n5637), .dout(n5649));
  jnot g05586(.din(n5649), .dout(n5650));
  jxor g05587(.dina(n5458), .dinb(n5457), .dout(n5651));
  jand g05588(.dina(n5651), .dinb(n5650), .dout(n5652));
  jnot g05589(.din(n5652), .dout(n5653));
  jxor g05590(.dina(n5651), .dinb(n5650), .dout(n5654));
  jnot g05591(.din(n5654), .dout(n5655));
  jand g05592(.dina(n4772), .dinb(n75), .dout(n5656));
  jand g05593(.dina(n4933), .dinb(n1213), .dout(n5657));
  jand g05594(.dina(n4918), .dinb(n1343), .dout(n5658));
  jand g05595(.dina(n4745), .dinb(n1445), .dout(n5659));
  jor  g05596(.dina(n5659), .dinb(n5658), .dout(n5660));
  jor  g05597(.dina(n5660), .dinb(n5657), .dout(n5661));
  jor  g05598(.dina(n5661), .dinb(n5656), .dout(n5662));
  jxor g05599(.dina(n5662), .dinb(n68), .dout(n5663));
  jor  g05600(.dina(n5663), .dinb(n5655), .dout(n5664));
  jand g05601(.dina(n5664), .dinb(n5653), .dout(n5665));
  jnot g05602(.din(n5665), .dout(n5666));
  jxor g05603(.dina(n5534), .dinb(n5533), .dout(n5667));
  jand g05604(.dina(n5667), .dinb(n5666), .dout(n5668));
  jor  g05605(.dina(n5668), .dinb(n5535), .dout(n5669));
  jxor g05606(.dina(n5487), .dinb(n5479), .dout(n5670));
  jand g05607(.dina(n5670), .dinb(n5669), .dout(n5671));
  jnot g05608(.din(n5671), .dout(n5672));
  jxor g05609(.dina(n5670), .dinb(n5669), .dout(n5673));
  jnot g05610(.din(n5673), .dout(n5674));
  jand g05611(.dina(n5365), .dinb(n4446), .dout(n5675));
  jand g05612(.dina(n5500), .dinb(n4451), .dout(n5676));
  jand g05613(.dina(n5424), .dinb(n4358), .dout(n5677));
  jand g05614(.dina(n5363), .dinb(n3853), .dout(n5678));
  jor  g05615(.dina(n5678), .dinb(n5677), .dout(n5679));
  jor  g05616(.dina(n5679), .dinb(n5676), .dout(n5680));
  jor  g05617(.dina(n5680), .dinb(n5675), .dout(n5681));
  jxor g05618(.dina(n5681), .dinb(n72), .dout(n5682));
  jor  g05619(.dina(n5682), .dinb(n5674), .dout(n5683));
  jand g05620(.dina(n5683), .dinb(n5672), .dout(n5684));
  jxor g05621(.dina(\a[19] ), .dinb(\a[18] ), .dout(n5685));
  jnot g05622(.din(n5685), .dout(n5686));
  jxor g05623(.dina(\a[18] ), .dinb(\a[17] ), .dout(n5687));
  jnot g05624(.din(n5687), .dout(n5688));
  jand g05625(.dina(n5688), .dinb(n5686), .dout(n5689));
  jxor g05626(.dina(\a[20] ), .dinb(\a[19] ), .dout(n5690));
  jand g05627(.dina(n5690), .dinb(n5689), .dout(n5691));
  jnot g05628(.din(n5691), .dout(n5692));
  jand g05629(.dina(n5690), .dinb(n5687), .dout(n5693));
  jnot g05630(.din(n5693), .dout(n5694));
  jor  g05631(.dina(n5694), .dinb(n4728), .dout(n5695));
  jand g05632(.dina(n5695), .dinb(n5692), .dout(n5696));
  jor  g05633(.dina(n5696), .dinb(n4630), .dout(n5697));
  jxor g05634(.dina(n5697), .dinb(\a[20] ), .dout(n5698));
  jor  g05635(.dina(n5698), .dinb(n5684), .dout(n5699));
  jxor g05636(.dina(n5698), .dinb(n5684), .dout(n5700));
  jxor g05637(.dina(n5505), .dinb(n5495), .dout(n5701));
  jand g05638(.dina(n5701), .dinb(n5700), .dout(n5702));
  jnot g05639(.din(n5702), .dout(n5703));
  jand g05640(.dina(n5703), .dinb(n5699), .dout(n5704));
  jnot g05641(.din(n5704), .dout(n5705));
  jxor g05642(.dina(n5518), .dinb(n5517), .dout(n5706));
  jand g05643(.dina(n5706), .dinb(n5705), .dout(n5707));
  jxor g05644(.dina(n5706), .dinb(n5705), .dout(n5708));
  jand g05645(.dina(n5365), .dinb(n4545), .dout(n5709));
  jand g05646(.dina(n5424), .dinb(n3853), .dout(n5710));
  jand g05647(.dina(n5500), .dinb(n4358), .dout(n5711));
  jand g05648(.dina(n5363), .dinb(n922), .dout(n5712));
  jor  g05649(.dina(n5712), .dinb(n5711), .dout(n5713));
  jor  g05650(.dina(n5713), .dinb(n5710), .dout(n5714));
  jor  g05651(.dina(n5714), .dinb(n5709), .dout(n5715));
  jxor g05652(.dina(n5715), .dinb(n72), .dout(n5716));
  jnot g05653(.din(n5716), .dout(n5717));
  jxor g05654(.dina(n5667), .dinb(n5666), .dout(n5718));
  jand g05655(.dina(n5718), .dinb(n5717), .dout(n5719));
  jand g05656(.dina(n5092), .dinb(n4449), .dout(n5720));
  jand g05657(.dina(n4453), .dinb(n1776), .dout(n5721));
  jand g05658(.dina(n4457), .dinb(n1862), .dout(n5722));
  jand g05659(.dina(n4461), .dinb(n1956), .dout(n5723));
  jor  g05660(.dina(n5723), .dinb(n5722), .dout(n5724));
  jor  g05661(.dina(n5724), .dinb(n5721), .dout(n5725));
  jor  g05662(.dina(n5725), .dinb(n5720), .dout(n5726));
  jxor g05663(.dina(n5726), .dinb(n88), .dout(n5727));
  jnot g05664(.din(n5727), .dout(n5728));
  jxor g05665(.dina(n5631), .dinb(n5623), .dout(n5729));
  jand g05666(.dina(n5729), .dinb(n5728), .dout(n5730));
  jxor g05667(.dina(n5614), .dinb(n5606), .dout(n5731));
  jnot g05668(.din(n5731), .dout(n5732));
  jand g05669(.dina(n815), .dinb(n801), .dout(n5733));
  jand g05670(.dina(n5733), .dinb(n228), .dout(n5734));
  jand g05671(.dina(n1178), .dinb(n566), .dout(n5735));
  jand g05672(.dina(n5735), .dinb(n205), .dout(n5736));
  jand g05673(.dina(n5736), .dinb(n5734), .dout(n5737));
  jand g05674(.dina(n5737), .dinb(n2947), .dout(n5738));
  jand g05675(.dina(n1881), .dinb(n658), .dout(n5739));
  jand g05676(.dina(n5739), .dinb(n3250), .dout(n5740));
  jand g05677(.dina(n508), .dinb(n324), .dout(n5741));
  jand g05678(.dina(n5741), .dinb(n262), .dout(n5742));
  jand g05679(.dina(n5742), .dinb(n4212), .dout(n5743));
  jand g05680(.dina(n5743), .dinb(n5740), .dout(n5744));
  jand g05681(.dina(n5744), .dinb(n5738), .dout(n5745));
  jand g05682(.dina(n5201), .dinb(n2419), .dout(n5746));
  jand g05683(.dina(n5746), .dinb(n5745), .dout(n5747));
  jand g05684(.dina(n1231), .dinb(n245), .dout(n5748));
  jand g05685(.dina(n5748), .dinb(n1034), .dout(n5749));
  jand g05686(.dina(n988), .dinb(n445), .dout(n5750));
  jand g05687(.dina(n5750), .dinb(n963), .dout(n5751));
  jand g05688(.dina(n5751), .dinb(n5749), .dout(n5752));
  jand g05689(.dina(n2676), .dinb(n199), .dout(n5753));
  jand g05690(.dina(n5753), .dinb(n5752), .dout(n5754));
  jand g05691(.dina(n432), .dinb(n305), .dout(n5755));
  jand g05692(.dina(n907), .dinb(n359), .dout(n5756));
  jand g05693(.dina(n5756), .dinb(n5755), .dout(n5757));
  jand g05694(.dina(n2847), .dinb(n2538), .dout(n5758));
  jand g05695(.dina(n5758), .dinb(n5757), .dout(n5759));
  jand g05696(.dina(n1641), .dinb(n671), .dout(n5760));
  jand g05697(.dina(n5760), .dinb(n1535), .dout(n5761));
  jand g05698(.dina(n4004), .dinb(n1676), .dout(n5762));
  jand g05699(.dina(n5762), .dinb(n5761), .dout(n5763));
  jand g05700(.dina(n5763), .dinb(n5759), .dout(n5764));
  jand g05701(.dina(n5764), .dinb(n5754), .dout(n5765));
  jand g05702(.dina(n4287), .dinb(n393), .dout(n5766));
  jand g05703(.dina(n5766), .dinb(n4619), .dout(n5767));
  jand g05704(.dina(n465), .dinb(n404), .dout(n5768));
  jand g05705(.dina(n5768), .dinb(n1024), .dout(n5769));
  jand g05706(.dina(n5259), .dinb(n883), .dout(n5770));
  jand g05707(.dina(n5770), .dinb(n5769), .dout(n5771));
  jand g05708(.dina(n441), .dinb(n431), .dout(n5772));
  jand g05709(.dina(n5772), .dinb(n583), .dout(n5773));
  jand g05710(.dina(n5773), .dinb(n3374), .dout(n5774));
  jand g05711(.dina(n5774), .dinb(n5771), .dout(n5775));
  jand g05712(.dina(n5775), .dinb(n5767), .dout(n5776));
  jand g05713(.dina(n5776), .dinb(n5765), .dout(n5777));
  jand g05714(.dina(n5777), .dinb(n5747), .dout(n5778));
  jand g05715(.dina(n5778), .dinb(n1292), .dout(n5779));
  jnot g05716(.din(n5779), .dout(n5780));
  jand g05717(.dina(n492), .dinb(n346), .dout(n5781));
  jand g05718(.dina(n5781), .dinb(n667), .dout(n5782));
  jand g05719(.dina(n4078), .dinb(n3450), .dout(n5783));
  jand g05720(.dina(n5783), .dinb(n5782), .dout(n5784));
  jand g05721(.dina(n1178), .dinb(n262), .dout(n5785));
  jand g05722(.dina(n696), .dinb(n372), .dout(n5786));
  jand g05723(.dina(n5786), .dinb(n5785), .dout(n5787));
  jand g05724(.dina(n5787), .dinb(n3290), .dout(n5788));
  jand g05725(.dina(n5788), .dinb(n5784), .dout(n5789));
  jand g05726(.dina(n382), .dinb(n280), .dout(n5790));
  jand g05727(.dina(n435), .dinb(n428), .dout(n5791));
  jand g05728(.dina(n5791), .dinb(n5790), .dout(n5792));
  jand g05729(.dina(n2622), .dinb(n709), .dout(n5793));
  jand g05730(.dina(n5793), .dinb(n5792), .dout(n5794));
  jand g05731(.dina(n614), .dinb(n197), .dout(n5795));
  jand g05732(.dina(n5795), .dinb(n671), .dout(n5796));
  jand g05733(.dina(n396), .dinb(n134), .dout(n5797));
  jand g05734(.dina(n417), .dinb(n305), .dout(n5798));
  jand g05735(.dina(n5798), .dinb(n5797), .dout(n5799));
  jand g05736(.dina(n5799), .dinb(n5796), .dout(n5800));
  jand g05737(.dina(n5800), .dinb(n5794), .dout(n5801));
  jand g05738(.dina(n1924), .dinb(n501), .dout(n5802));
  jand g05739(.dina(n2499), .dinb(n2164), .dout(n5803));
  jand g05740(.dina(n5803), .dinb(n5802), .dout(n5804));
  jand g05741(.dina(n5804), .dinb(n1583), .dout(n5805));
  jand g05742(.dina(n5805), .dinb(n5801), .dout(n5806));
  jand g05743(.dina(n5806), .dinb(n5789), .dout(n5807));
  jand g05744(.dina(n687), .dinb(n605), .dout(n5808));
  jand g05745(.dina(n5808), .dinb(n385), .dout(n5809));
  jand g05746(.dina(n979), .dinb(n924), .dout(n5810));
  jand g05747(.dina(n5810), .dinb(n1760), .dout(n5811));
  jand g05748(.dina(n5811), .dinb(n5809), .dout(n5812));
  jand g05749(.dina(n907), .dinb(n249), .dout(n5813));
  jand g05750(.dina(n1231), .dinb(n357), .dout(n5814));
  jand g05751(.dina(n5814), .dinb(n5813), .dout(n5815));
  jand g05752(.dina(n5815), .dinb(n1966), .dout(n5816));
  jand g05753(.dina(n5816), .dinb(n5812), .dout(n5817));
  jand g05754(.dina(n1899), .dinb(n1296), .dout(n5818));
  jand g05755(.dina(n1160), .dinb(n506), .dout(n5819));
  jand g05756(.dina(n5819), .dinb(n5818), .dout(n5820));
  jand g05757(.dina(n5158), .dinb(n596), .dout(n5821));
  jand g05758(.dina(n2384), .dinb(n1676), .dout(n5822));
  jand g05759(.dina(n5822), .dinb(n5821), .dout(n5823));
  jand g05760(.dina(n5823), .dinb(n5820), .dout(n5824));
  jand g05761(.dina(n5824), .dinb(n5817), .dout(n5825));
  jand g05762(.dina(n5825), .dinb(n4137), .dout(n5826));
  jand g05763(.dina(n5776), .dinb(n3877), .dout(n5827));
  jand g05764(.dina(n5827), .dinb(n5826), .dout(n5828));
  jand g05765(.dina(n5828), .dinb(n5807), .dout(n5829));
  jnot g05766(.din(n5829), .dout(n5830));
  jand g05767(.dina(n5830), .dinb(n5780), .dout(n5831));
  jnot g05768(.din(n5831), .dout(n5832));
  jnot g05769(.din(\a[11] ), .dout(n5833));
  jand g05770(.dina(n5829), .dinb(n5779), .dout(n5834));
  jnot g05771(.din(n5834), .dout(n5835));
  jand g05772(.dina(n5835), .dinb(n5833), .dout(n5836));
  jand g05773(.dina(n5836), .dinb(n5832), .dout(n5837));
  jnot g05774(.din(n5837), .dout(n5838));
  jand g05775(.dina(n5838), .dinb(n5832), .dout(n5839));
  jnot g05776(.din(n5839), .dout(n5840));
  jand g05777(.dina(n5840), .dinb(n5220), .dout(n5841));
  jnot g05778(.din(n5841), .dout(n5842));
  jand g05779(.dina(n5839), .dinb(n5221), .dout(n5843));
  jxor g05780(.dina(n3733), .dinb(n3732), .dout(n5844));
  jand g05781(.dina(n5844), .dinb(n732), .dout(n5845));
  jand g05782(.dina(n3851), .dinb(n2411), .dout(n5846));
  jand g05783(.dina(n3855), .dinb(n2237), .dout(n5847));
  jand g05784(.dina(n3858), .dinb(n2343), .dout(n5848));
  jor  g05785(.dina(n5848), .dinb(n5847), .dout(n5849));
  jor  g05786(.dina(n5849), .dinb(n5846), .dout(n5850));
  jor  g05787(.dina(n5850), .dinb(n5845), .dout(n5851));
  jnot g05788(.din(n5851), .dout(n5852));
  jor  g05789(.dina(n5852), .dinb(n5843), .dout(n5853));
  jand g05790(.dina(n5853), .dinb(n5842), .dout(n5854));
  jor  g05791(.dina(n5854), .dinb(n5732), .dout(n5855));
  jxor g05792(.dina(n5854), .dinb(n5732), .dout(n5856));
  jnot g05793(.din(n5856), .dout(n5857));
  jand g05794(.dina(n5838), .dinb(n5833), .dout(n5858));
  jand g05795(.dina(n5839), .dinb(n5835), .dout(n5859));
  jor  g05796(.dina(n5859), .dinb(n5858), .dout(n5860));
  jxor g05797(.dina(n3730), .dinb(n3729), .dout(n5861));
  jand g05798(.dina(n5861), .dinb(n732), .dout(n5862));
  jand g05799(.dina(n3858), .dinb(n2411), .dout(n5863));
  jand g05800(.dina(n3855), .dinb(n2343), .dout(n5864));
  jand g05801(.dina(n3851), .dinb(n2497), .dout(n5865));
  jor  g05802(.dina(n5865), .dinb(n5864), .dout(n5866));
  jor  g05803(.dina(n5866), .dinb(n5863), .dout(n5867));
  jor  g05804(.dina(n5867), .dinb(n5862), .dout(n5868));
  jand g05805(.dina(n5868), .dinb(n5860), .dout(n5869));
  jand g05806(.dina(n700), .dinb(n311), .dout(n5870));
  jand g05807(.dina(n5870), .dinb(n198), .dout(n5871));
  jand g05808(.dina(n842), .dinb(n749), .dout(n5872));
  jand g05809(.dina(n5872), .dinb(n607), .dout(n5873));
  jand g05810(.dina(n5873), .dinb(n5871), .dout(n5874));
  jand g05811(.dina(n515), .dinb(n268), .dout(n5875));
  jand g05812(.dina(n5875), .dinb(n253), .dout(n5876));
  jand g05813(.dina(n5876), .dinb(n1820), .dout(n5877));
  jand g05814(.dina(n5877), .dinb(n5874), .dout(n5878));
  jand g05815(.dina(n1519), .dinb(n763), .dout(n5879));
  jand g05816(.dina(n1047), .dinb(n505), .dout(n5880));
  jand g05817(.dina(n5880), .dinb(n5879), .dout(n5881));
  jand g05818(.dina(n5881), .dinb(n2769), .dout(n5882));
  jand g05819(.dina(n1231), .dinb(n658), .dout(n5883));
  jand g05820(.dina(n5883), .dinb(n3471), .dout(n5884));
  jand g05821(.dina(n2784), .dinb(n2742), .dout(n5885));
  jand g05822(.dina(n5885), .dinb(n5884), .dout(n5886));
  jand g05823(.dina(n5886), .dinb(n5882), .dout(n5887));
  jand g05824(.dina(n5887), .dinb(n5878), .dout(n5888));
  jand g05825(.dina(n5888), .dinb(n3900), .dout(n5889));
  jand g05826(.dina(n5889), .dinb(n2451), .dout(n5890));
  jand g05827(.dina(n5890), .dinb(n2443), .dout(n5891));
  jand g05828(.dina(n5891), .dinb(n1674), .dout(n5892));
  jor  g05829(.dina(n5892), .dinb(n5780), .dout(n5893));
  jxor g05830(.dina(n5892), .dinb(n5780), .dout(n5894));
  jnot g05831(.din(n5894), .dout(n5895));
  jand g05832(.dina(n687), .dinb(n417), .dout(n5896));
  jand g05833(.dina(n5896), .dinb(n633), .dout(n5897));
  jnot g05834(.din(n3219), .dout(n5898));
  jand g05835(.dina(n1144), .dinb(n926), .dout(n5899));
  jand g05836(.dina(n5899), .dinb(n5898), .dout(n5900));
  jand g05837(.dina(n5900), .dinb(n5897), .dout(n5901));
  jand g05838(.dina(n643), .dinb(n336), .dout(n5902));
  jand g05839(.dina(n793), .dinb(n418), .dout(n5903));
  jand g05840(.dina(n5903), .dinb(n894), .dout(n5904));
  jand g05841(.dina(n5904), .dinb(n5902), .dout(n5905));
  jand g05842(.dina(n5905), .dinb(n5901), .dout(n5906));
  jand g05843(.dina(n5906), .dinb(n2686), .dout(n5907));
  jand g05844(.dina(n678), .dinb(n386), .dout(n5908));
  jand g05845(.dina(n5908), .dinb(n305), .dout(n5909));
  jand g05846(.dina(n2897), .dinb(n2560), .dout(n5910));
  jand g05847(.dina(n5910), .dinb(n3866), .dout(n5911));
  jand g05848(.dina(n5911), .dinb(n5909), .dout(n5912));
  jand g05849(.dina(n2015), .dinb(n1273), .dout(n5913));
  jand g05850(.dina(n5913), .dinb(n1997), .dout(n5914));
  jand g05851(.dina(n626), .dinb(n574), .dout(n5915));
  jand g05852(.dina(n5915), .dinb(n5813), .dout(n5916));
  jand g05853(.dina(n3417), .dinb(n2315), .dout(n5917));
  jand g05854(.dina(n5917), .dinb(n5916), .dout(n5918));
  jand g05855(.dina(n5918), .dinb(n5914), .dout(n5919));
  jand g05856(.dina(n508), .dinb(n274), .dout(n5920));
  jand g05857(.dina(n5920), .dinb(n605), .dout(n5921));
  jand g05858(.dina(n5921), .dinb(n565), .dout(n5922));
  jand g05859(.dina(n5922), .dinb(n5796), .dout(n5923));
  jand g05860(.dina(n5923), .dinb(n5919), .dout(n5924));
  jand g05861(.dina(n5924), .dinb(n5912), .dout(n5925));
  jand g05862(.dina(n5925), .dinb(n5907), .dout(n5926));
  jand g05863(.dina(n1039), .dinb(n527), .dout(n5927));
  jand g05864(.dina(n5927), .dinb(n478), .dout(n5928));
  jand g05865(.dina(n715), .dinb(n243), .dout(n5929));
  jand g05866(.dina(n503), .dinb(n288), .dout(n5930));
  jand g05867(.dina(n5930), .dinb(n5929), .dout(n5931));
  jand g05868(.dina(n5931), .dinb(n5928), .dout(n5932));
  jand g05869(.dina(n5185), .dinb(n2050), .dout(n5933));
  jand g05870(.dina(n5933), .dinb(n5932), .dout(n5934));
  jand g05871(.dina(n3160), .dinb(n1130), .dout(n5935));
  jand g05872(.dina(n5935), .dinb(n3838), .dout(n5936));
  jand g05873(.dina(n5936), .dinb(n1915), .dout(n5937));
  jand g05874(.dina(n5937), .dinb(n5934), .dout(n5938));
  jand g05875(.dina(n284), .dinb(n194), .dout(n5939));
  jand g05876(.dina(n826), .dinb(n302), .dout(n5940));
  jand g05877(.dina(n607), .dinb(n184), .dout(n5941));
  jand g05878(.dina(n5941), .dinb(n5940), .dout(n5942));
  jand g05879(.dina(n5942), .dinb(n5939), .dout(n5943));
  jand g05880(.dina(n5943), .dinb(n3022), .dout(n5944));
  jand g05881(.dina(n462), .dinb(n257), .dout(n5945));
  jand g05882(.dina(n756), .dinb(n533), .dout(n5946));
  jand g05883(.dina(n5946), .dinb(n5945), .dout(n5947));
  jand g05884(.dina(n1221), .dinb(n696), .dout(n5948));
  jand g05885(.dina(n1409), .dinb(n967), .dout(n5949));
  jand g05886(.dina(n5949), .dinb(n5948), .dout(n5950));
  jand g05887(.dina(n5950), .dinb(n5947), .dout(n5951));
  jand g05888(.dina(n5951), .dinb(n3932), .dout(n5952));
  jand g05889(.dina(n5952), .dinb(n5944), .dout(n5953));
  jand g05890(.dina(n5953), .dinb(n5938), .dout(n5954));
  jand g05891(.dina(n330), .dinb(n309), .dout(n5955));
  jand g05892(.dina(n5955), .dinb(n2053), .dout(n5956));
  jand g05893(.dina(n5956), .dinb(n3056), .dout(n5957));
  jand g05894(.dina(n5957), .dinb(n4100), .dout(n5958));
  jand g05895(.dina(n3233), .dinb(n501), .dout(n5959));
  jand g05896(.dina(n5959), .dinb(n1585), .dout(n5960));
  jand g05897(.dina(n595), .dinb(n174), .dout(n5961));
  jand g05898(.dina(n543), .dinb(n136), .dout(n5962));
  jand g05899(.dina(n5962), .dinb(n5961), .dout(n5963));
  jnot g05900(.din(n4004), .dout(n5964));
  jor  g05901(.dina(n5964), .dinb(n3316), .dout(n5965));
  jnot g05902(.din(n5965), .dout(n5966));
  jand g05903(.dina(n5966), .dinb(n5963), .dout(n5967));
  jand g05904(.dina(n5967), .dinb(n5960), .dout(n5968));
  jand g05905(.dina(n5968), .dinb(n5958), .dout(n5969));
  jand g05906(.dina(n5969), .dinb(n5272), .dout(n5970));
  jand g05907(.dina(n5970), .dinb(n5954), .dout(n5971));
  jand g05908(.dina(n5971), .dinb(n5926), .dout(n5972));
  jnot g05909(.din(n5972), .dout(n5973));
  jand g05910(.dina(n882), .dinb(n214), .dout(n5974));
  jand g05911(.dina(n5974), .dinb(n4500), .dout(n5975));
  jand g05912(.dina(n771), .dinb(n563), .dout(n5976));
  jand g05913(.dina(n5976), .dinb(n5975), .dout(n5977));
  jand g05914(.dina(n1130), .dinb(n554), .dout(n5978));
  jand g05915(.dina(n3092), .dinb(n2483), .dout(n5979));
  jand g05916(.dina(n5979), .dinb(n5978), .dout(n5980));
  jand g05917(.dina(n5980), .dinb(n5977), .dout(n5981));
  jand g05918(.dina(n647), .dinb(n268), .dout(n5982));
  jand g05919(.dina(n5982), .dinb(n815), .dout(n5983));
  jand g05920(.dina(n5983), .dinb(n4782), .dout(n5984));
  jand g05921(.dina(n5984), .dinb(n5981), .dout(n5985));
  jand g05922(.dina(n317), .dinb(n180), .dout(n5986));
  jand g05923(.dina(n395), .dinb(n146), .dout(n5987));
  jand g05924(.dina(n5987), .dinb(n5986), .dout(n5988));
  jnot g05925(.din(n3216), .dout(n5989));
  jand g05926(.dina(n3819), .dinb(n5989), .dout(n5990));
  jand g05927(.dina(n5990), .dinb(n5988), .dout(n5991));
  jand g05928(.dina(n1085), .dinb(n243), .dout(n5992));
  jand g05929(.dina(n505), .dinb(n325), .dout(n5993));
  jand g05930(.dina(n5993), .dinb(n500), .dout(n5994));
  jand g05931(.dina(n5994), .dinb(n5992), .dout(n5995));
  jand g05932(.dina(n5995), .dinb(n5991), .dout(n5996));
  jand g05933(.dina(n712), .dinb(n245), .dout(n5997));
  jand g05934(.dina(n778), .dinb(n467), .dout(n5998));
  jand g05935(.dina(n5998), .dinb(n5997), .dout(n5999));
  jand g05936(.dina(n4611), .dinb(n794), .dout(n6000));
  jand g05937(.dina(n6000), .dinb(n5999), .dout(n6001));
  jand g05938(.dina(n6001), .dinb(n1852), .dout(n6002));
  jand g05939(.dina(n6002), .dinb(n5996), .dout(n6003));
  jand g05940(.dina(n6003), .dinb(n5985), .dout(n6004));
  jand g05941(.dina(n1231), .dinb(n483), .dout(n6005));
  jand g05942(.dina(n1153), .dinb(n643), .dout(n6006));
  jand g05943(.dina(n6006), .dinb(n6005), .dout(n6007));
  jand g05944(.dina(n671), .dinb(n428), .dout(n6008));
  jand g05945(.dina(n6008), .dinb(n355), .dout(n6009));
  jand g05946(.dina(n6009), .dinb(n6007), .dout(n6010));
  jand g05947(.dina(n6010), .dinb(n3481), .dout(n6011));
  jand g05948(.dina(n1145), .dinb(n877), .dout(n6012));
  jand g05949(.dina(n1196), .dinb(n436), .dout(n6013));
  jand g05950(.dina(n6013), .dinb(n6012), .dout(n6014));
  jand g05951(.dina(n6014), .dinb(n4791), .dout(n6015));
  jand g05952(.dina(n6015), .dinb(n6011), .dout(n6016));
  jand g05953(.dina(n4487), .dinb(n2413), .dout(n6017));
  jand g05954(.dina(n1584), .dinb(n777), .dout(n6018));
  jand g05955(.dina(n6018), .dinb(n6017), .dout(n6019));
  jand g05956(.dina(n1346), .dinb(n134), .dout(n6020));
  jand g05957(.dina(n6020), .dinb(n763), .dout(n6021));
  jand g05958(.dina(n583), .dinb(n516), .dout(n6022));
  jand g05959(.dina(n6022), .dinb(n1959), .dout(n6023));
  jand g05960(.dina(n6023), .dinb(n6021), .dout(n6024));
  jand g05961(.dina(n6024), .dinb(n6019), .dout(n6025));
  jand g05962(.dina(n857), .dinb(n103), .dout(n6026));
  jand g05963(.dina(n1519), .dinb(n1264), .dout(n6027));
  jand g05964(.dina(n6027), .dinb(n6026), .dout(n6028));
  jand g05965(.dina(n2150), .dinb(n2106), .dout(n6029));
  jand g05966(.dina(n6029), .dinb(n4668), .dout(n6030));
  jand g05967(.dina(n6030), .dinb(n6028), .dout(n6031));
  jand g05968(.dina(n6031), .dinb(n6025), .dout(n6032));
  jand g05969(.dina(n6032), .dinb(n6016), .dout(n6033));
  jand g05970(.dina(n6033), .dinb(n6004), .dout(n6034));
  jand g05971(.dina(n6034), .dinb(n4831), .dout(n6035));
  jnot g05972(.din(n6035), .dout(n6036));
  jand g05973(.dina(n6036), .dinb(n5973), .dout(n6037));
  jnot g05974(.din(n6037), .dout(n6038));
  jnot g05975(.din(\a[8] ), .dout(n6039));
  jand g05976(.dina(n6035), .dinb(n5972), .dout(n6040));
  jnot g05977(.din(n6040), .dout(n6041));
  jand g05978(.dina(n6041), .dinb(n6039), .dout(n6042));
  jand g05979(.dina(n6042), .dinb(n6038), .dout(n6043));
  jnot g05980(.din(n6043), .dout(n6044));
  jand g05981(.dina(n6044), .dinb(n6038), .dout(n6045));
  jnot g05982(.din(n6045), .dout(n6046));
  jand g05983(.dina(n6046), .dinb(n5779), .dout(n6047));
  jnot g05984(.din(n6047), .dout(n6048));
  jand g05985(.dina(n6045), .dinb(n5780), .dout(n6049));
  jxor g05986(.dina(n3724), .dinb(n3723), .dout(n6050));
  jand g05987(.dina(n6050), .dinb(n732), .dout(n6051));
  jand g05988(.dina(n3858), .dinb(n2602), .dout(n6052));
  jand g05989(.dina(n3851), .dinb(n2695), .dout(n6053));
  jand g05990(.dina(n3855), .dinb(n2497), .dout(n6054));
  jor  g05991(.dina(n6054), .dinb(n6053), .dout(n6055));
  jor  g05992(.dina(n6055), .dinb(n6052), .dout(n6056));
  jor  g05993(.dina(n6056), .dinb(n6051), .dout(n6057));
  jnot g05994(.din(n6057), .dout(n6058));
  jor  g05995(.dina(n6058), .dinb(n6049), .dout(n6059));
  jand g05996(.dina(n6059), .dinb(n6048), .dout(n6060));
  jor  g05997(.dina(n6060), .dinb(n5895), .dout(n6061));
  jand g05998(.dina(n6061), .dinb(n5893), .dout(n6062));
  jnot g05999(.din(n6062), .dout(n6063));
  jxor g06000(.dina(n5868), .dinb(n5860), .dout(n6064));
  jand g06001(.dina(n6064), .dinb(n6063), .dout(n6065));
  jor  g06002(.dina(n6065), .dinb(n5869), .dout(n6066));
  jxor g06003(.dina(n5839), .dinb(n5221), .dout(n6067));
  jxor g06004(.dina(n6067), .dinb(n5851), .dout(n6068));
  jand g06005(.dina(n6068), .dinb(n6066), .dout(n6069));
  jnot g06006(.din(n6069), .dout(n6070));
  jxor g06007(.dina(n6068), .dinb(n6066), .dout(n6071));
  jnot g06008(.din(n6071), .dout(n6072));
  jand g06009(.dina(n5303), .dinb(n4449), .dout(n6073));
  jand g06010(.dina(n4461), .dinb(n2128), .dout(n6074));
  jand g06011(.dina(n4457), .dinb(n2067), .dout(n6075));
  jand g06012(.dina(n4453), .dinb(n1956), .dout(n6076));
  jor  g06013(.dina(n6076), .dinb(n6075), .dout(n6077));
  jor  g06014(.dina(n6077), .dinb(n6074), .dout(n6078));
  jor  g06015(.dina(n6078), .dinb(n6073), .dout(n6079));
  jxor g06016(.dina(n6079), .dinb(n88), .dout(n6080));
  jor  g06017(.dina(n6080), .dinb(n6072), .dout(n6081));
  jand g06018(.dina(n6081), .dinb(n6070), .dout(n6082));
  jor  g06019(.dina(n6082), .dinb(n5857), .dout(n6083));
  jand g06020(.dina(n6083), .dinb(n5855), .dout(n6084));
  jnot g06021(.din(n6084), .dout(n6085));
  jxor g06022(.dina(n5729), .dinb(n5728), .dout(n6086));
  jand g06023(.dina(n6086), .dinb(n6085), .dout(n6087));
  jor  g06024(.dina(n6087), .dinb(n5730), .dout(n6088));
  jxor g06025(.dina(n5647), .dinb(n5639), .dout(n6089));
  jand g06026(.dina(n6089), .dinb(n6088), .dout(n6090));
  jnot g06027(.din(n6090), .dout(n6091));
  jxor g06028(.dina(n6089), .dinb(n6088), .dout(n6092));
  jnot g06029(.din(n6092), .dout(n6093));
  jand g06030(.dina(n4258), .dinb(n75), .dout(n6094));
  jand g06031(.dina(n4933), .dinb(n1343), .dout(n6095));
  jand g06032(.dina(n4918), .dinb(n1445), .dout(n6096));
  jand g06033(.dina(n4745), .dinb(n1560), .dout(n6097));
  jor  g06034(.dina(n6097), .dinb(n6096), .dout(n6098));
  jor  g06035(.dina(n6098), .dinb(n6095), .dout(n6099));
  jor  g06036(.dina(n6099), .dinb(n6094), .dout(n6100));
  jxor g06037(.dina(n6100), .dinb(n68), .dout(n6101));
  jor  g06038(.dina(n6101), .dinb(n6093), .dout(n6102));
  jand g06039(.dina(n6102), .dinb(n6091), .dout(n6103));
  jnot g06040(.din(n6103), .dout(n6104));
  jxor g06041(.dina(n5663), .dinb(n5655), .dout(n6105));
  jand g06042(.dina(n6105), .dinb(n6104), .dout(n6106));
  jnot g06043(.din(n6106), .dout(n6107));
  jxor g06044(.dina(n6105), .dinb(n6104), .dout(n6108));
  jnot g06045(.din(n6108), .dout(n6109));
  jand g06046(.dina(n5365), .dinb(n3848), .dout(n6110));
  jand g06047(.dina(n5424), .dinb(n922), .dout(n6111));
  jand g06048(.dina(n5500), .dinb(n3853), .dout(n6112));
  jand g06049(.dina(n5363), .dinb(n1076), .dout(n6113));
  jor  g06050(.dina(n6113), .dinb(n6112), .dout(n6114));
  jor  g06051(.dina(n6114), .dinb(n6111), .dout(n6115));
  jor  g06052(.dina(n6115), .dinb(n6110), .dout(n6116));
  jxor g06053(.dina(n6116), .dinb(n72), .dout(n6117));
  jor  g06054(.dina(n6117), .dinb(n6109), .dout(n6118));
  jand g06055(.dina(n6118), .dinb(n6107), .dout(n6119));
  jnot g06056(.din(n6119), .dout(n6120));
  jxor g06057(.dina(n5718), .dinb(n5717), .dout(n6121));
  jand g06058(.dina(n6121), .dinb(n6120), .dout(n6122));
  jor  g06059(.dina(n6122), .dinb(n5719), .dout(n6123));
  jxor g06060(.dina(n5682), .dinb(n5674), .dout(n6124));
  jand g06061(.dina(n6124), .dinb(n6123), .dout(n6125));
  jnot g06062(.din(n6125), .dout(n6126));
  jxor g06063(.dina(n6124), .dinb(n6123), .dout(n6127));
  jnot g06064(.din(n6127), .dout(n6128));
  jor  g06065(.dina(n5694), .dinb(n4731), .dout(n6129));
  jor  g06066(.dina(n5692), .dinb(n4597), .dout(n6130));
  jand g06067(.dina(n5688), .dinb(n5685), .dout(n6131));
  jnot g06068(.din(n6131), .dout(n6132));
  jor  g06069(.dina(n6132), .dinb(n4630), .dout(n6133));
  jand g06070(.dina(n6133), .dinb(n6130), .dout(n6134));
  jand g06071(.dina(n6134), .dinb(n6129), .dout(n6135));
  jxor g06072(.dina(n6135), .dinb(\a[20] ), .dout(n6136));
  jor  g06073(.dina(n6136), .dinb(n6128), .dout(n6137));
  jand g06074(.dina(n6137), .dinb(n6126), .dout(n6138));
  jnot g06075(.din(n6138), .dout(n6139));
  jxor g06076(.dina(n5701), .dinb(n5700), .dout(n6140));
  jand g06077(.dina(n6140), .dinb(n6139), .dout(n6141));
  jxor g06078(.dina(n6140), .dinb(n6139), .dout(n6142));
  jxor g06079(.dina(n6086), .dinb(n6085), .dout(n6143));
  jnot g06080(.din(n6143), .dout(n6144));
  jand g06081(.dina(n4866), .dinb(n75), .dout(n6145));
  jand g06082(.dina(n4918), .dinb(n1560), .dout(n6146));
  jand g06083(.dina(n4745), .dinb(n1624), .dout(n6147));
  jand g06084(.dina(n4933), .dinb(n1445), .dout(n6148));
  jor  g06085(.dina(n6148), .dinb(n6147), .dout(n6149));
  jor  g06086(.dina(n6149), .dinb(n6146), .dout(n6150));
  jor  g06087(.dina(n6150), .dinb(n6145), .dout(n6151));
  jxor g06088(.dina(n6151), .dinb(n68), .dout(n6152));
  jor  g06089(.dina(n6152), .dinb(n6144), .dout(n6153));
  jxor g06090(.dina(n6082), .dinb(n5857), .dout(n6154));
  jnot g06091(.din(n6154), .dout(n6155));
  jand g06092(.dina(n5440), .dinb(n4449), .dout(n6156));
  jand g06093(.dina(n4461), .dinb(n2067), .dout(n6157));
  jand g06094(.dina(n4457), .dinb(n1956), .dout(n6158));
  jand g06095(.dina(n4453), .dinb(n1862), .dout(n6159));
  jor  g06096(.dina(n6159), .dinb(n6158), .dout(n6160));
  jor  g06097(.dina(n6160), .dinb(n6157), .dout(n6161));
  jor  g06098(.dina(n6161), .dinb(n6156), .dout(n6162));
  jxor g06099(.dina(n6162), .dinb(n88), .dout(n6163));
  jor  g06100(.dina(n6163), .dinb(n6155), .dout(n6164));
  jand g06101(.dina(n4849), .dinb(n75), .dout(n6165));
  jand g06102(.dina(n4933), .dinb(n1560), .dout(n6166));
  jand g06103(.dina(n4918), .dinb(n1624), .dout(n6167));
  jand g06104(.dina(n4745), .dinb(n1776), .dout(n6168));
  jor  g06105(.dina(n6168), .dinb(n6167), .dout(n6169));
  jor  g06106(.dina(n6169), .dinb(n6166), .dout(n6170));
  jor  g06107(.dina(n6170), .dinb(n6165), .dout(n6171));
  jxor g06108(.dina(n6171), .dinb(n68), .dout(n6172));
  jnot g06109(.din(n6172), .dout(n6173));
  jxor g06110(.dina(n6163), .dinb(n6155), .dout(n6174));
  jand g06111(.dina(n6174), .dinb(n6173), .dout(n6175));
  jnot g06112(.din(n6175), .dout(n6176));
  jand g06113(.dina(n6176), .dinb(n6164), .dout(n6177));
  jnot g06114(.din(n6177), .dout(n6178));
  jxor g06115(.dina(n6152), .dinb(n6144), .dout(n6179));
  jand g06116(.dina(n6179), .dinb(n6178), .dout(n6180));
  jnot g06117(.din(n6180), .dout(n6181));
  jand g06118(.dina(n6181), .dinb(n6153), .dout(n6182));
  jnot g06119(.din(n6182), .dout(n6183));
  jxor g06120(.dina(n6101), .dinb(n6093), .dout(n6184));
  jand g06121(.dina(n6184), .dinb(n6183), .dout(n6185));
  jnot g06122(.din(n6185), .dout(n6186));
  jxor g06123(.dina(n6184), .dinb(n6183), .dout(n6187));
  jnot g06124(.din(n6187), .dout(n6188));
  jand g06125(.dina(n5365), .dinb(n4026), .dout(n6189));
  jand g06126(.dina(n5424), .dinb(n1076), .dout(n6190));
  jand g06127(.dina(n5500), .dinb(n922), .dout(n6191));
  jand g06128(.dina(n5363), .dinb(n1213), .dout(n6192));
  jor  g06129(.dina(n6192), .dinb(n6191), .dout(n6193));
  jor  g06130(.dina(n6193), .dinb(n6190), .dout(n6194));
  jor  g06131(.dina(n6194), .dinb(n6189), .dout(n6195));
  jxor g06132(.dina(n6195), .dinb(n72), .dout(n6196));
  jor  g06133(.dina(n6196), .dinb(n6188), .dout(n6197));
  jand g06134(.dina(n6197), .dinb(n6186), .dout(n6198));
  jnot g06135(.din(n6198), .dout(n6199));
  jxor g06136(.dina(n6117), .dinb(n6109), .dout(n6200));
  jand g06137(.dina(n6200), .dinb(n6199), .dout(n6201));
  jnot g06138(.din(n6201), .dout(n6202));
  jxor g06139(.dina(n6200), .dinb(n6199), .dout(n6203));
  jnot g06140(.din(n6203), .dout(n6204));
  jand g06141(.dina(n5693), .dinb(n4752), .dout(n6205));
  jand g06142(.dina(n6131), .dinb(n4451), .dout(n6206));
  jand g06143(.dina(n5691), .dinb(n4358), .dout(n6207));
  jor  g06144(.dina(n5690), .dinb(n5688), .dout(n6208));
  jnot g06145(.din(n6208), .dout(n6209));
  jand g06146(.dina(n6209), .dinb(n4598), .dout(n6210));
  jor  g06147(.dina(n6210), .dinb(n6207), .dout(n6211));
  jor  g06148(.dina(n6211), .dinb(n6206), .dout(n6212));
  jor  g06149(.dina(n6212), .dinb(n6205), .dout(n6213));
  jxor g06150(.dina(n6213), .dinb(n4247), .dout(n6214));
  jor  g06151(.dina(n6214), .dinb(n6204), .dout(n6215));
  jand g06152(.dina(n6215), .dinb(n6202), .dout(n6216));
  jand g06153(.dina(n5693), .dinb(n4636), .dout(n6217));
  jand g06154(.dina(n5691), .dinb(n4451), .dout(n6218));
  jand g06155(.dina(n6131), .dinb(n4598), .dout(n6219));
  jand g06156(.dina(n6209), .dinb(n4631), .dout(n6220));
  jor  g06157(.dina(n6220), .dinb(n6219), .dout(n6221));
  jor  g06158(.dina(n6221), .dinb(n6218), .dout(n6222));
  jor  g06159(.dina(n6222), .dinb(n6217), .dout(n6223));
  jxor g06160(.dina(n6223), .dinb(n4247), .dout(n6224));
  jor  g06161(.dina(n6224), .dinb(n6216), .dout(n6225));
  jxor g06162(.dina(n6121), .dinb(n6120), .dout(n6226));
  jxor g06163(.dina(n6224), .dinb(n6216), .dout(n6227));
  jand g06164(.dina(n6227), .dinb(n6226), .dout(n6228));
  jnot g06165(.din(n6228), .dout(n6229));
  jand g06166(.dina(n6229), .dinb(n6225), .dout(n6230));
  jnot g06167(.din(n6230), .dout(n6231));
  jxor g06168(.dina(n6136), .dinb(n6128), .dout(n6232));
  jand g06169(.dina(n6232), .dinb(n6231), .dout(n6233));
  jxor g06170(.dina(n6232), .dinb(n6231), .dout(n6234));
  jand g06171(.dina(n5365), .dinb(n4043), .dout(n6235));
  jand g06172(.dina(n5500), .dinb(n1076), .dout(n6236));
  jand g06173(.dina(n5424), .dinb(n1213), .dout(n6237));
  jand g06174(.dina(n5363), .dinb(n1343), .dout(n6238));
  jor  g06175(.dina(n6238), .dinb(n6237), .dout(n6239));
  jor  g06176(.dina(n6239), .dinb(n6236), .dout(n6240));
  jor  g06177(.dina(n6240), .dinb(n6235), .dout(n6241));
  jxor g06178(.dina(n6241), .dinb(n72), .dout(n6242));
  jnot g06179(.din(n6242), .dout(n6243));
  jxor g06180(.dina(n6179), .dinb(n6178), .dout(n6244));
  jand g06181(.dina(n6244), .dinb(n6243), .dout(n6245));
  jxor g06182(.dina(n6060), .dinb(n5895), .dout(n6246));
  jxor g06183(.dina(n3727), .dinb(n3726), .dout(n6247));
  jand g06184(.dina(n6247), .dinb(n732), .dout(n6248));
  jand g06185(.dina(n3855), .dinb(n2411), .dout(n6249));
  jand g06186(.dina(n3851), .dinb(n2602), .dout(n6250));
  jand g06187(.dina(n3858), .dinb(n2497), .dout(n6251));
  jor  g06188(.dina(n6251), .dinb(n6250), .dout(n6252));
  jor  g06189(.dina(n6252), .dinb(n6249), .dout(n6253));
  jor  g06190(.dina(n6253), .dinb(n6248), .dout(n6254));
  jand g06191(.dina(n6254), .dinb(n6246), .dout(n6255));
  jand g06192(.dina(n5607), .dinb(n4449), .dout(n6256));
  jand g06193(.dina(n4457), .dinb(n2237), .dout(n6257));
  jand g06194(.dina(n4461), .dinb(n2343), .dout(n6258));
  jand g06195(.dina(n4453), .dinb(n2128), .dout(n6259));
  jor  g06196(.dina(n6259), .dinb(n6258), .dout(n6260));
  jor  g06197(.dina(n6260), .dinb(n6257), .dout(n6261));
  jor  g06198(.dina(n6261), .dinb(n6256), .dout(n6262));
  jxor g06199(.dina(n6262), .dinb(n88), .dout(n6263));
  jnot g06200(.din(n6263), .dout(n6264));
  jxor g06201(.dina(n6254), .dinb(n6246), .dout(n6265));
  jand g06202(.dina(n6265), .dinb(n6264), .dout(n6266));
  jor  g06203(.dina(n6266), .dinb(n6255), .dout(n6267));
  jxor g06204(.dina(n6064), .dinb(n6063), .dout(n6268));
  jand g06205(.dina(n6268), .dinb(n6267), .dout(n6269));
  jand g06206(.dina(n5624), .dinb(n4449), .dout(n6270));
  jand g06207(.dina(n4461), .dinb(n2237), .dout(n6271));
  jand g06208(.dina(n4457), .dinb(n2128), .dout(n6272));
  jand g06209(.dina(n4453), .dinb(n2067), .dout(n6273));
  jor  g06210(.dina(n6273), .dinb(n6272), .dout(n6274));
  jor  g06211(.dina(n6274), .dinb(n6271), .dout(n6275));
  jor  g06212(.dina(n6275), .dinb(n6270), .dout(n6276));
  jxor g06213(.dina(n6276), .dinb(n88), .dout(n6277));
  jnot g06214(.din(n6277), .dout(n6278));
  jxor g06215(.dina(n6268), .dinb(n6267), .dout(n6279));
  jand g06216(.dina(n6279), .dinb(n6278), .dout(n6280));
  jor  g06217(.dina(n6280), .dinb(n6269), .dout(n6281));
  jxor g06218(.dina(n6080), .dinb(n6072), .dout(n6282));
  jand g06219(.dina(n6282), .dinb(n6281), .dout(n6283));
  jnot g06220(.din(n6283), .dout(n6284));
  jxor g06221(.dina(n6282), .dinb(n6281), .dout(n6285));
  jnot g06222(.din(n6285), .dout(n6286));
  jand g06223(.dina(n5075), .dinb(n75), .dout(n6287));
  jand g06224(.dina(n4933), .dinb(n1624), .dout(n6288));
  jand g06225(.dina(n4918), .dinb(n1776), .dout(n6289));
  jand g06226(.dina(n4745), .dinb(n1862), .dout(n6290));
  jor  g06227(.dina(n6290), .dinb(n6289), .dout(n6291));
  jor  g06228(.dina(n6291), .dinb(n6288), .dout(n6292));
  jor  g06229(.dina(n6292), .dinb(n6287), .dout(n6293));
  jxor g06230(.dina(n6293), .dinb(n68), .dout(n6294));
  jor  g06231(.dina(n6294), .dinb(n6286), .dout(n6295));
  jand g06232(.dina(n6295), .dinb(n6284), .dout(n6296));
  jnot g06233(.din(n6296), .dout(n6297));
  jxor g06234(.dina(n6174), .dinb(n6173), .dout(n6298));
  jand g06235(.dina(n6298), .dinb(n6297), .dout(n6299));
  jnot g06236(.din(n6299), .dout(n6300));
  jxor g06237(.dina(n6298), .dinb(n6297), .dout(n6301));
  jnot g06238(.din(n6301), .dout(n6302));
  jand g06239(.dina(n5365), .dinb(n4772), .dout(n6303));
  jand g06240(.dina(n5500), .dinb(n1213), .dout(n6304));
  jand g06241(.dina(n5424), .dinb(n1343), .dout(n6305));
  jand g06242(.dina(n5363), .dinb(n1445), .dout(n6306));
  jor  g06243(.dina(n6306), .dinb(n6305), .dout(n6307));
  jor  g06244(.dina(n6307), .dinb(n6304), .dout(n6308));
  jor  g06245(.dina(n6308), .dinb(n6303), .dout(n6309));
  jxor g06246(.dina(n6309), .dinb(n72), .dout(n6310));
  jor  g06247(.dina(n6310), .dinb(n6302), .dout(n6311));
  jand g06248(.dina(n6311), .dinb(n6300), .dout(n6312));
  jnot g06249(.din(n6312), .dout(n6313));
  jxor g06250(.dina(n6244), .dinb(n6243), .dout(n6314));
  jand g06251(.dina(n6314), .dinb(n6313), .dout(n6315));
  jor  g06252(.dina(n6315), .dinb(n6245), .dout(n6316));
  jxor g06253(.dina(n6196), .dinb(n6188), .dout(n6317));
  jand g06254(.dina(n6317), .dinb(n6316), .dout(n6318));
  jnot g06255(.din(n6318), .dout(n6319));
  jxor g06256(.dina(n6317), .dinb(n6316), .dout(n6320));
  jnot g06257(.din(n6320), .dout(n6321));
  jand g06258(.dina(n5693), .dinb(n4446), .dout(n6322));
  jand g06259(.dina(n6209), .dinb(n4451), .dout(n6323));
  jand g06260(.dina(n6131), .dinb(n4358), .dout(n6324));
  jand g06261(.dina(n5691), .dinb(n3853), .dout(n6325));
  jor  g06262(.dina(n6325), .dinb(n6324), .dout(n6326));
  jor  g06263(.dina(n6326), .dinb(n6323), .dout(n6327));
  jor  g06264(.dina(n6327), .dinb(n6322), .dout(n6328));
  jxor g06265(.dina(n6328), .dinb(n4247), .dout(n6329));
  jor  g06266(.dina(n6329), .dinb(n6321), .dout(n6330));
  jand g06267(.dina(n6330), .dinb(n6319), .dout(n6331));
  jxor g06268(.dina(\a[16] ), .dinb(\a[15] ), .dout(n6332));
  jnot g06269(.din(n6332), .dout(n6333));
  jxor g06270(.dina(\a[15] ), .dinb(\a[14] ), .dout(n6334));
  jnot g06271(.din(n6334), .dout(n6335));
  jand g06272(.dina(n6335), .dinb(n6333), .dout(n6336));
  jxor g06273(.dina(\a[17] ), .dinb(\a[16] ), .dout(n6337));
  jand g06274(.dina(n6337), .dinb(n6336), .dout(n6338));
  jnot g06275(.din(n6338), .dout(n6339));
  jand g06276(.dina(n6337), .dinb(n6334), .dout(n6340));
  jnot g06277(.din(n6340), .dout(n6341));
  jor  g06278(.dina(n6341), .dinb(n4728), .dout(n6342));
  jand g06279(.dina(n6342), .dinb(n6339), .dout(n6343));
  jor  g06280(.dina(n6343), .dinb(n4630), .dout(n6344));
  jxor g06281(.dina(n6344), .dinb(\a[17] ), .dout(n6345));
  jor  g06282(.dina(n6345), .dinb(n6331), .dout(n6346));
  jxor g06283(.dina(n6345), .dinb(n6331), .dout(n6347));
  jxor g06284(.dina(n6214), .dinb(n6204), .dout(n6348));
  jand g06285(.dina(n6348), .dinb(n6347), .dout(n6349));
  jnot g06286(.din(n6349), .dout(n6350));
  jand g06287(.dina(n6350), .dinb(n6346), .dout(n6351));
  jnot g06288(.din(n6351), .dout(n6352));
  jxor g06289(.dina(n6227), .dinb(n6226), .dout(n6353));
  jand g06290(.dina(n6353), .dinb(n6352), .dout(n6354));
  jxor g06291(.dina(n6314), .dinb(n6313), .dout(n6355));
  jnot g06292(.din(n6355), .dout(n6356));
  jand g06293(.dina(n5693), .dinb(n4545), .dout(n6357));
  jand g06294(.dina(n5691), .dinb(n922), .dout(n6358));
  jand g06295(.dina(n6131), .dinb(n3853), .dout(n6359));
  jand g06296(.dina(n6209), .dinb(n4358), .dout(n6360));
  jor  g06297(.dina(n6360), .dinb(n6359), .dout(n6361));
  jor  g06298(.dina(n6361), .dinb(n6358), .dout(n6362));
  jor  g06299(.dina(n6362), .dinb(n6357), .dout(n6363));
  jxor g06300(.dina(n6363), .dinb(n4247), .dout(n6364));
  jor  g06301(.dina(n6364), .dinb(n6356), .dout(n6365));
  jand g06302(.dina(n5092), .dinb(n75), .dout(n6366));
  jand g06303(.dina(n4918), .dinb(n1862), .dout(n6367));
  jand g06304(.dina(n4745), .dinb(n1956), .dout(n6368));
  jand g06305(.dina(n4933), .dinb(n1776), .dout(n6369));
  jor  g06306(.dina(n6369), .dinb(n6368), .dout(n6370));
  jor  g06307(.dina(n6370), .dinb(n6367), .dout(n6371));
  jor  g06308(.dina(n6371), .dinb(n6366), .dout(n6372));
  jxor g06309(.dina(n6372), .dinb(n68), .dout(n6373));
  jnot g06310(.din(n6373), .dout(n6374));
  jxor g06311(.dina(n6279), .dinb(n6278), .dout(n6375));
  jand g06312(.dina(n6375), .dinb(n6374), .dout(n6376));
  jand g06313(.dina(n751), .dinb(n325), .dout(n6377));
  jand g06314(.dina(n6377), .dinb(n309), .dout(n6378));
  jand g06315(.dina(n505), .dinb(n494), .dout(n6379));
  jand g06316(.dina(n1178), .dinb(n108), .dout(n6380));
  jand g06317(.dina(n6380), .dinb(n6379), .dout(n6381));
  jand g06318(.dina(n4996), .dinb(n1581), .dout(n6382));
  jand g06319(.dina(n6382), .dinb(n6381), .dout(n6383));
  jand g06320(.dina(n6383), .dinb(n6378), .dout(n6384));
  jand g06321(.dina(n1039), .dinb(n154), .dout(n6385));
  jand g06322(.dina(n6385), .dinb(n717), .dout(n6386));
  jand g06323(.dina(n3462), .dinb(n1383), .dout(n6387));
  jand g06324(.dina(n6387), .dinb(n6386), .dout(n6388));
  jand g06325(.dina(n6388), .dinb(n5977), .dout(n6389));
  jand g06326(.dina(n6389), .dinb(n6384), .dout(n6390));
  jand g06327(.dina(n6390), .dinb(n5912), .dout(n6391));
  jnot g06328(.din(n1693), .dout(n6392));
  jand g06329(.dina(n1221), .dinb(n435), .dout(n6393));
  jand g06330(.dina(n842), .dinb(n270), .dout(n6394));
  jand g06331(.dina(n6394), .dinb(n6393), .dout(n6395));
  jand g06332(.dina(n4163), .dinb(n2240), .dout(n6396));
  jand g06333(.dina(n6396), .dinb(n6395), .dout(n6397));
  jand g06334(.dina(n3905), .dinb(n996), .dout(n6398));
  jand g06335(.dina(n6398), .dinb(n6397), .dout(n6399));
  jand g06336(.dina(n1284), .dinb(n1153), .dout(n6400));
  jand g06337(.dina(n6400), .dinb(n1204), .dout(n6401));
  jand g06338(.dina(n5986), .dinb(n1934), .dout(n6402));
  jand g06339(.dina(n6402), .dinb(n2483), .dout(n6403));
  jand g06340(.dina(n6403), .dinb(n6401), .dout(n6404));
  jand g06341(.dina(n6404), .dinb(n6399), .dout(n6405));
  jand g06342(.dina(n6405), .dinb(n6392), .dout(n6406));
  jand g06343(.dina(n6406), .dinb(n6391), .dout(n6407));
  jand g06344(.dina(n6407), .dinb(n4207), .dout(n6408));
  jor  g06345(.dina(n6408), .dinb(n5973), .dout(n6409));
  jand g06346(.dina(n793), .dinb(n221), .dout(n6410));
  jand g06347(.dina(n6410), .dinb(n197), .dout(n6411));
  jand g06348(.dina(n874), .dinb(n527), .dout(n6412));
  jand g06349(.dina(n6412), .dinb(n1319), .dout(n6413));
  jand g06350(.dina(n6413), .dinb(n6411), .dout(n6414));
  jand g06351(.dina(n1611), .dinb(n628), .dout(n6415));
  jand g06352(.dina(n6415), .dinb(n6414), .dout(n6416));
  jand g06353(.dina(n586), .dinb(n113), .dout(n6417));
  jand g06354(.dina(n1500), .dinb(n1185), .dout(n6418));
  jand g06355(.dina(n6418), .dinb(n6417), .dout(n6419));
  jand g06356(.dina(n6419), .dinb(n1302), .dout(n6420));
  jand g06357(.dina(n6420), .dinb(n6416), .dout(n6421));
  jand g06358(.dina(n967), .dinb(n959), .dout(n6422));
  jand g06359(.dina(n6422), .dinb(n842), .dout(n6423));
  jand g06360(.dina(n1047), .dinb(n274), .dout(n6424));
  jand g06361(.dina(n6424), .dinb(n1199), .dout(n6425));
  jand g06362(.dina(n6425), .dinb(n2359), .dout(n6426));
  jand g06363(.dina(n6426), .dinb(n6423), .dout(n6427));
  jand g06364(.dina(n6427), .dinb(n1229), .dout(n6428));
  jand g06365(.dina(n6428), .dinb(n6421), .dout(n6429));
  jand g06366(.dina(n6429), .dinb(n402), .dout(n6430));
  jand g06367(.dina(n6430), .dinb(n5241), .dout(n6431));
  jor  g06368(.dina(n6431), .dinb(\a[2] ), .dout(n6432));
  jxor g06369(.dina(n6431), .dinb(\a[2] ), .dout(n6433));
  jand g06370(.dina(n6433), .dinb(n64), .dout(n6434));
  jnot g06371(.din(n6434), .dout(n6435));
  jand g06372(.dina(n6435), .dinb(n6432), .dout(n6436));
  jor  g06373(.dina(n6436), .dinb(n5973), .dout(n6437));
  jxor g06374(.dina(n6436), .dinb(n5973), .dout(n6438));
  jxor g06375(.dina(n3713), .dinb(n3711), .dout(n6439));
  jand g06376(.dina(n6439), .dinb(n732), .dout(n6440));
  jand g06377(.dina(n3858), .dinb(n2808), .dout(n6441));
  jand g06378(.dina(n3855), .dinb(n2732), .dout(n6442));
  jand g06379(.dina(n3851), .dinb(n2867), .dout(n6443));
  jor  g06380(.dina(n6443), .dinb(n6442), .dout(n6444));
  jor  g06381(.dina(n6444), .dinb(n6441), .dout(n6445));
  jor  g06382(.dina(n6445), .dinb(n6440), .dout(n6446));
  jand g06383(.dina(n6446), .dinb(n6438), .dout(n6447));
  jnot g06384(.din(n6447), .dout(n6448));
  jand g06385(.dina(n6448), .dinb(n6437), .dout(n6449));
  jnot g06386(.din(n6449), .dout(n6450));
  jxor g06387(.dina(n6408), .dinb(n5973), .dout(n6451));
  jand g06388(.dina(n6451), .dinb(n6450), .dout(n6452));
  jnot g06389(.din(n6452), .dout(n6453));
  jand g06390(.dina(n6453), .dinb(n6409), .dout(n6454));
  jnot g06391(.din(n6454), .dout(n6455));
  jand g06392(.dina(n6044), .dinb(n6039), .dout(n6456));
  jand g06393(.dina(n6045), .dinb(n6041), .dout(n6457));
  jor  g06394(.dina(n6457), .dinb(n6456), .dout(n6458));
  jand g06395(.dina(n6458), .dinb(n6455), .dout(n6459));
  jnot g06396(.din(n6459), .dout(n6460));
  jxor g06397(.dina(n6458), .dinb(n6455), .dout(n6461));
  jnot g06398(.din(n6461), .dout(n6462));
  jnot g06399(.din(n732), .dout(n6463));
  jxor g06400(.dina(n3721), .dinb(n3719), .dout(n6464));
  jor  g06401(.dina(n6464), .dinb(n6463), .dout(n6465));
  jand g06402(.dina(n3855), .dinb(n2602), .dout(n6466));
  jand g06403(.dina(n3858), .dinb(n2695), .dout(n6467));
  jand g06404(.dina(n3851), .dinb(n2732), .dout(n6468));
  jor  g06405(.dina(n6468), .dinb(n6467), .dout(n6469));
  jor  g06406(.dina(n6469), .dinb(n6466), .dout(n6470));
  jnot g06407(.din(n6470), .dout(n6471));
  jand g06408(.dina(n6471), .dinb(n6465), .dout(n6472));
  jor  g06409(.dina(n6472), .dinb(n6462), .dout(n6473));
  jand g06410(.dina(n6473), .dinb(n6460), .dout(n6474));
  jnot g06411(.din(n6474), .dout(n6475));
  jxor g06412(.dina(n6045), .dinb(n5780), .dout(n6476));
  jxor g06413(.dina(n6476), .dinb(n6057), .dout(n6477));
  jand g06414(.dina(n6477), .dinb(n6475), .dout(n6478));
  jnot g06415(.din(n6478), .dout(n6479));
  jxor g06416(.dina(n6477), .dinb(n6475), .dout(n6480));
  jnot g06417(.din(n6480), .dout(n6481));
  jand g06418(.dina(n5844), .dinb(n4449), .dout(n6482));
  jand g06419(.dina(n4461), .dinb(n2411), .dout(n6483));
  jand g06420(.dina(n4453), .dinb(n2237), .dout(n6484));
  jand g06421(.dina(n4457), .dinb(n2343), .dout(n6485));
  jor  g06422(.dina(n6485), .dinb(n6484), .dout(n6486));
  jor  g06423(.dina(n6486), .dinb(n6483), .dout(n6487));
  jor  g06424(.dina(n6487), .dinb(n6482), .dout(n6488));
  jxor g06425(.dina(n6488), .dinb(n88), .dout(n6489));
  jor  g06426(.dina(n6489), .dinb(n6481), .dout(n6490));
  jand g06427(.dina(n6490), .dinb(n6479), .dout(n6491));
  jnot g06428(.din(n6491), .dout(n6492));
  jxor g06429(.dina(n6265), .dinb(n6264), .dout(n6493));
  jand g06430(.dina(n6493), .dinb(n6492), .dout(n6494));
  jnot g06431(.din(n6494), .dout(n6495));
  jxor g06432(.dina(n6493), .dinb(n6492), .dout(n6496));
  jnot g06433(.din(n6496), .dout(n6497));
  jand g06434(.dina(n5440), .dinb(n75), .dout(n6498));
  jand g06435(.dina(n4918), .dinb(n1956), .dout(n6499));
  jand g06436(.dina(n4933), .dinb(n1862), .dout(n6500));
  jand g06437(.dina(n4745), .dinb(n2067), .dout(n6501));
  jor  g06438(.dina(n6501), .dinb(n6500), .dout(n6502));
  jor  g06439(.dina(n6502), .dinb(n6499), .dout(n6503));
  jor  g06440(.dina(n6503), .dinb(n6498), .dout(n6504));
  jxor g06441(.dina(n6504), .dinb(n68), .dout(n6505));
  jor  g06442(.dina(n6505), .dinb(n6497), .dout(n6506));
  jand g06443(.dina(n6506), .dinb(n6495), .dout(n6507));
  jnot g06444(.din(n6507), .dout(n6508));
  jxor g06445(.dina(n6375), .dinb(n6374), .dout(n6509));
  jand g06446(.dina(n6509), .dinb(n6508), .dout(n6510));
  jor  g06447(.dina(n6510), .dinb(n6376), .dout(n6511));
  jxor g06448(.dina(n6294), .dinb(n6286), .dout(n6512));
  jand g06449(.dina(n6512), .dinb(n6511), .dout(n6513));
  jnot g06450(.din(n6513), .dout(n6514));
  jxor g06451(.dina(n6512), .dinb(n6511), .dout(n6515));
  jnot g06452(.din(n6515), .dout(n6516));
  jand g06453(.dina(n5365), .dinb(n4258), .dout(n6517));
  jand g06454(.dina(n5500), .dinb(n1343), .dout(n6518));
  jand g06455(.dina(n5424), .dinb(n1445), .dout(n6519));
  jand g06456(.dina(n5363), .dinb(n1560), .dout(n6520));
  jor  g06457(.dina(n6520), .dinb(n6519), .dout(n6521));
  jor  g06458(.dina(n6521), .dinb(n6518), .dout(n6522));
  jor  g06459(.dina(n6522), .dinb(n6517), .dout(n6523));
  jxor g06460(.dina(n6523), .dinb(n72), .dout(n6524));
  jor  g06461(.dina(n6524), .dinb(n6516), .dout(n6525));
  jand g06462(.dina(n6525), .dinb(n6514), .dout(n6526));
  jnot g06463(.din(n6526), .dout(n6527));
  jxor g06464(.dina(n6310), .dinb(n6302), .dout(n6528));
  jand g06465(.dina(n6528), .dinb(n6527), .dout(n6529));
  jnot g06466(.din(n6529), .dout(n6530));
  jxor g06467(.dina(n6528), .dinb(n6527), .dout(n6531));
  jnot g06468(.din(n6531), .dout(n6532));
  jand g06469(.dina(n5693), .dinb(n3848), .dout(n6533));
  jand g06470(.dina(n6131), .dinb(n922), .dout(n6534));
  jand g06471(.dina(n6209), .dinb(n3853), .dout(n6535));
  jand g06472(.dina(n5691), .dinb(n1076), .dout(n6536));
  jor  g06473(.dina(n6536), .dinb(n6535), .dout(n6537));
  jor  g06474(.dina(n6537), .dinb(n6534), .dout(n6538));
  jor  g06475(.dina(n6538), .dinb(n6533), .dout(n6539));
  jxor g06476(.dina(n6539), .dinb(n4247), .dout(n6540));
  jor  g06477(.dina(n6540), .dinb(n6532), .dout(n6541));
  jand g06478(.dina(n6541), .dinb(n6530), .dout(n6542));
  jnot g06479(.din(n6542), .dout(n6543));
  jxor g06480(.dina(n6364), .dinb(n6356), .dout(n6544));
  jand g06481(.dina(n6544), .dinb(n6543), .dout(n6545));
  jnot g06482(.din(n6545), .dout(n6546));
  jand g06483(.dina(n6546), .dinb(n6365), .dout(n6547));
  jnot g06484(.din(n6547), .dout(n6548));
  jxor g06485(.dina(n6329), .dinb(n6321), .dout(n6549));
  jand g06486(.dina(n6549), .dinb(n6548), .dout(n6550));
  jnot g06487(.din(n6550), .dout(n6551));
  jxor g06488(.dina(n6549), .dinb(n6548), .dout(n6552));
  jnot g06489(.din(n6552), .dout(n6553));
  jor  g06490(.dina(n6341), .dinb(n4731), .dout(n6554));
  jor  g06491(.dina(n6339), .dinb(n4597), .dout(n6555));
  jand g06492(.dina(n6335), .dinb(n6332), .dout(n6556));
  jnot g06493(.din(n6556), .dout(n6557));
  jor  g06494(.dina(n6557), .dinb(n4630), .dout(n6558));
  jand g06495(.dina(n6558), .dinb(n6555), .dout(n6559));
  jand g06496(.dina(n6559), .dinb(n6554), .dout(n6560));
  jxor g06497(.dina(n6560), .dinb(\a[17] ), .dout(n6561));
  jor  g06498(.dina(n6561), .dinb(n6553), .dout(n6562));
  jand g06499(.dina(n6562), .dinb(n6551), .dout(n6563));
  jnot g06500(.din(n6563), .dout(n6564));
  jxor g06501(.dina(n6348), .dinb(n6347), .dout(n6565));
  jand g06502(.dina(n6565), .dinb(n6564), .dout(n6566));
  jxor g06503(.dina(n6565), .dinb(n6564), .dout(n6567));
  jand g06504(.dina(n5365), .dinb(n4866), .dout(n6568));
  jand g06505(.dina(n5500), .dinb(n1445), .dout(n6569));
  jand g06506(.dina(n5424), .dinb(n1560), .dout(n6570));
  jand g06507(.dina(n5363), .dinb(n1624), .dout(n6571));
  jor  g06508(.dina(n6571), .dinb(n6570), .dout(n6572));
  jor  g06509(.dina(n6572), .dinb(n6569), .dout(n6573));
  jor  g06510(.dina(n6573), .dinb(n6568), .dout(n6574));
  jxor g06511(.dina(n6574), .dinb(n72), .dout(n6575));
  jnot g06512(.din(n6575), .dout(n6576));
  jxor g06513(.dina(n6509), .dinb(n6508), .dout(n6577));
  jand g06514(.dina(n6577), .dinb(n6576), .dout(n6578));
  jand g06515(.dina(n5861), .dinb(n4449), .dout(n6579));
  jand g06516(.dina(n4457), .dinb(n2411), .dout(n6580));
  jand g06517(.dina(n4453), .dinb(n2343), .dout(n6581));
  jand g06518(.dina(n4461), .dinb(n2497), .dout(n6582));
  jor  g06519(.dina(n6582), .dinb(n6581), .dout(n6583));
  jor  g06520(.dina(n6583), .dinb(n6580), .dout(n6584));
  jor  g06521(.dina(n6584), .dinb(n6579), .dout(n6585));
  jxor g06522(.dina(n6585), .dinb(n88), .dout(n6586));
  jnot g06523(.din(n6586), .dout(n6587));
  jxor g06524(.dina(n6472), .dinb(n6462), .dout(n6588));
  jand g06525(.dina(n6588), .dinb(n6587), .dout(n6589));
  jxor g06526(.dina(n6451), .dinb(n6450), .dout(n6590));
  jxor g06527(.dina(n3717), .dinb(n3715), .dout(n6591));
  jand g06528(.dina(n6591), .dinb(n732), .dout(n6592));
  jand g06529(.dina(n3855), .dinb(n2695), .dout(n6593));
  jand g06530(.dina(n3851), .dinb(n2808), .dout(n6594));
  jand g06531(.dina(n3858), .dinb(n2732), .dout(n6595));
  jor  g06532(.dina(n6595), .dinb(n6594), .dout(n6596));
  jor  g06533(.dina(n6596), .dinb(n6593), .dout(n6597));
  jor  g06534(.dina(n6597), .dinb(n6592), .dout(n6598));
  jand g06535(.dina(n6598), .dinb(n6590), .dout(n6599));
  jnot g06536(.din(\a[2] ), .dout(n6600));
  jand g06537(.dina(n404), .dinb(n348), .dout(n6601));
  jand g06538(.dina(n6601), .dinb(n751), .dout(n6602));
  jand g06539(.dina(n2940), .dinb(n844), .dout(n6603));
  jand g06540(.dina(n6603), .dinb(n6602), .dout(n6604));
  jand g06541(.dina(n5211), .dinb(n552), .dout(n6605));
  jand g06542(.dina(n6605), .dinb(n429), .dout(n6606));
  jand g06543(.dina(n6606), .dinb(n2007), .dout(n6607));
  jand g06544(.dina(n6607), .dinb(n6604), .dout(n6608));
  jand g06545(.dina(n626), .dinb(n515), .dout(n6609));
  jand g06546(.dina(n6609), .dinb(n486), .dout(n6610));
  jand g06547(.dina(n4796), .dinb(n2556), .dout(n6611));
  jand g06548(.dina(n1134), .dinb(n976), .dout(n6612));
  jand g06549(.dina(n6612), .dinb(n6611), .dout(n6613));
  jand g06550(.dina(n6613), .dinb(n6610), .dout(n6614));
  jand g06551(.dina(n462), .dinb(n113), .dout(n6615));
  jand g06552(.dina(n322), .dinb(n245), .dout(n6616));
  jand g06553(.dina(n6616), .dinb(n6615), .dout(n6617));
  jand g06554(.dina(n6617), .dinb(n1183), .dout(n6618));
  jand g06555(.dina(n5871), .dinb(n5787), .dout(n6619));
  jand g06556(.dina(n6619), .dinb(n6618), .dout(n6620));
  jand g06557(.dina(n6620), .dinb(n6614), .dout(n6621));
  jand g06558(.dina(n6621), .dinb(n6608), .dout(n6622));
  jand g06559(.dina(n6622), .dinb(n948), .dout(n6623));
  jand g06560(.dina(n3225), .dinb(n2923), .dout(n6624));
  jand g06561(.dina(n6624), .dinb(n6623), .dout(n6625));
  jor  g06562(.dina(n6625), .dinb(n6600), .dout(n6626));
  jand g06563(.dina(n1014), .dinb(n194), .dout(n6627));
  jand g06564(.dina(n6627), .dinb(n1104), .dout(n6628));
  jand g06565(.dina(n6628), .dinb(n1295), .dout(n6629));
  jand g06566(.dina(n6629), .dinb(n1277), .dout(n6630));
  jand g06567(.dina(n3865), .dinb(n1603), .dout(n6631));
  jand g06568(.dina(n6631), .dinb(n552), .dout(n6632));
  jand g06569(.dina(n6632), .dinb(n5157), .dout(n6633));
  jand g06570(.dina(n6633), .dinb(n6630), .dout(n6634));
  jand g06571(.dina(n874), .dinb(n252), .dout(n6635));
  jand g06572(.dina(n234), .dinb(n180), .dout(n6636));
  jand g06573(.dina(n6636), .dinb(n6635), .dout(n6637));
  jand g06574(.dina(n2278), .dinb(n1663), .dout(n6638));
  jand g06575(.dina(n6638), .dinb(n6637), .dout(n6639));
  jand g06576(.dina(n5550), .dinb(n1050), .dout(n6640));
  jand g06577(.dina(n6640), .dinb(n6639), .dout(n6641));
  jand g06578(.dina(n6641), .dinb(n498), .dout(n6642));
  jand g06579(.dina(n6642), .dinb(n6634), .dout(n6643));
  jand g06580(.dina(n6643), .dinb(n1441), .dout(n6644));
  jand g06581(.dina(n6644), .dinb(n3456), .dout(n6645));
  jor  g06582(.dina(n6645), .dinb(n6600), .dout(n6646));
  jand g06583(.dina(n5876), .dinb(n3422), .dout(n6647));
  jand g06584(.dina(n6647), .dinb(n1183), .dout(n6648));
  jand g06585(.dina(n2713), .dinb(n722), .dout(n6649));
  jand g06586(.dina(n1295), .dinb(n1128), .dout(n6650));
  jand g06587(.dina(n6650), .dinb(n6649), .dout(n6651));
  jand g06588(.dina(n391), .dinb(n375), .dout(n6652));
  jand g06589(.dina(n6652), .dinb(n786), .dout(n6653));
  jand g06590(.dina(n383), .dinb(n365), .dout(n6654));
  jand g06591(.dina(n6654), .dinb(n1881), .dout(n6655));
  jand g06592(.dina(n6655), .dinb(n6653), .dout(n6656));
  jand g06593(.dina(n6656), .dinb(n6651), .dout(n6657));
  jand g06594(.dina(n6657), .dinb(n5901), .dout(n6658));
  jand g06595(.dina(n6658), .dinb(n6648), .dout(n6659));
  jand g06596(.dina(n508), .dinb(n290), .dout(n6660));
  jand g06597(.dina(n6660), .dinb(n429), .dout(n6661));
  jand g06598(.dina(n5588), .dinb(n1364), .dout(n6662));
  jand g06599(.dina(n6662), .dinb(n6661), .dout(n6663));
  jand g06600(.dina(n6663), .dinb(n4515), .dout(n6664));
  jand g06601(.dina(n658), .dinb(n461), .dout(n6665));
  jand g06602(.dina(n6665), .dinb(n609), .dout(n6666));
  jand g06603(.dina(n736), .dinb(n711), .dout(n6667));
  jand g06604(.dina(n6667), .dinb(n218), .dout(n6668));
  jand g06605(.dina(n6668), .dinb(n6666), .dout(n6669));
  jand g06606(.dina(n3595), .dinb(n3009), .dout(n6670));
  jand g06607(.dina(n6670), .dinb(n5153), .dout(n6671));
  jand g06608(.dina(n6671), .dinb(n6669), .dout(n6672));
  jand g06609(.dina(n6672), .dinb(n6664), .dout(n6673));
  jand g06610(.dina(n4481), .dinb(n3561), .dout(n6674));
  jand g06611(.dina(n6674), .dinb(n6673), .dout(n6675));
  jand g06612(.dina(n6675), .dinb(n6659), .dout(n6676));
  jand g06613(.dina(n6676), .dinb(n2170), .dout(n6677));
  jor  g06614(.dina(n6677), .dinb(n6600), .dout(n6678));
  jxor g06615(.dina(n6677), .dinb(n6600), .dout(n6679));
  jnot g06616(.din(n6679), .dout(n6680));
  jxor g06617(.dina(n3696), .dinb(n3695), .dout(n6681));
  jor  g06618(.dina(n6681), .dinb(n6463), .dout(n6682));
  jand g06619(.dina(n3858), .dinb(n3086), .dout(n6683));
  jand g06620(.dina(n3855), .dinb(n2991), .dout(n6684));
  jand g06621(.dina(n3851), .dinb(n3183), .dout(n6685));
  jor  g06622(.dina(n6685), .dinb(n6684), .dout(n6686));
  jor  g06623(.dina(n6686), .dinb(n6683), .dout(n6687));
  jnot g06624(.din(n6687), .dout(n6688));
  jand g06625(.dina(n6688), .dinb(n6682), .dout(n6689));
  jor  g06626(.dina(n6689), .dinb(n6680), .dout(n6690));
  jand g06627(.dina(n6690), .dinb(n6678), .dout(n6691));
  jnot g06628(.din(n6691), .dout(n6692));
  jxor g06629(.dina(n6645), .dinb(n6600), .dout(n6693));
  jand g06630(.dina(n6693), .dinb(n6692), .dout(n6694));
  jnot g06631(.din(n6694), .dout(n6695));
  jand g06632(.dina(n6695), .dinb(n6646), .dout(n6696));
  jnot g06633(.din(n6696), .dout(n6697));
  jxor g06634(.dina(n6625), .dinb(n6600), .dout(n6698));
  jand g06635(.dina(n6698), .dinb(n6697), .dout(n6699));
  jnot g06636(.din(n6699), .dout(n6700));
  jand g06637(.dina(n6700), .dinb(n6626), .dout(n6701));
  jnot g06638(.din(n6701), .dout(n6702));
  jxor g06639(.dina(n6433), .dinb(n64), .dout(n6703));
  jand g06640(.dina(n6703), .dinb(n6702), .dout(n6704));
  jxor g06641(.dina(n6703), .dinb(n6702), .dout(n6705));
  jxor g06642(.dina(n3709), .dinb(n3707), .dout(n6706));
  jand g06643(.dina(n6706), .dinb(n732), .dout(n6707));
  jand g06644(.dina(n3855), .dinb(n2808), .dout(n6708));
  jand g06645(.dina(n3851), .dinb(n2954), .dout(n6709));
  jand g06646(.dina(n3858), .dinb(n2867), .dout(n6710));
  jor  g06647(.dina(n6710), .dinb(n6709), .dout(n6711));
  jor  g06648(.dina(n6711), .dinb(n6708), .dout(n6712));
  jor  g06649(.dina(n6712), .dinb(n6707), .dout(n6713));
  jand g06650(.dina(n6713), .dinb(n6705), .dout(n6714));
  jor  g06651(.dina(n6714), .dinb(n6704), .dout(n6715));
  jxor g06652(.dina(n6446), .dinb(n6438), .dout(n6716));
  jand g06653(.dina(n6716), .dinb(n6715), .dout(n6717));
  jnot g06654(.din(n6717), .dout(n6718));
  jxor g06655(.dina(n6716), .dinb(n6715), .dout(n6719));
  jnot g06656(.din(n6719), .dout(n6720));
  jand g06657(.dina(n6050), .dinb(n4449), .dout(n6721));
  jand g06658(.dina(n4457), .dinb(n2602), .dout(n6722));
  jand g06659(.dina(n4461), .dinb(n2695), .dout(n6723));
  jand g06660(.dina(n4453), .dinb(n2497), .dout(n6724));
  jor  g06661(.dina(n6724), .dinb(n6723), .dout(n6725));
  jor  g06662(.dina(n6725), .dinb(n6722), .dout(n6726));
  jor  g06663(.dina(n6726), .dinb(n6721), .dout(n6727));
  jxor g06664(.dina(n6727), .dinb(n88), .dout(n6728));
  jor  g06665(.dina(n6728), .dinb(n6720), .dout(n6729));
  jand g06666(.dina(n6729), .dinb(n6718), .dout(n6730));
  jnot g06667(.din(n6730), .dout(n6731));
  jxor g06668(.dina(n6598), .dinb(n6590), .dout(n6732));
  jand g06669(.dina(n6732), .dinb(n6731), .dout(n6733));
  jor  g06670(.dina(n6733), .dinb(n6599), .dout(n6734));
  jxor g06671(.dina(n6588), .dinb(n6587), .dout(n6735));
  jand g06672(.dina(n6735), .dinb(n6734), .dout(n6736));
  jor  g06673(.dina(n6736), .dinb(n6589), .dout(n6737));
  jxor g06674(.dina(n6489), .dinb(n6481), .dout(n6738));
  jand g06675(.dina(n6738), .dinb(n6737), .dout(n6739));
  jnot g06676(.din(n6739), .dout(n6740));
  jxor g06677(.dina(n6738), .dinb(n6737), .dout(n6741));
  jnot g06678(.din(n6741), .dout(n6742));
  jand g06679(.dina(n5303), .dinb(n75), .dout(n6743));
  jand g06680(.dina(n4918), .dinb(n2067), .dout(n6744));
  jand g06681(.dina(n4933), .dinb(n1956), .dout(n6745));
  jand g06682(.dina(n4745), .dinb(n2128), .dout(n6746));
  jor  g06683(.dina(n6746), .dinb(n6745), .dout(n6747));
  jor  g06684(.dina(n6747), .dinb(n6744), .dout(n6748));
  jor  g06685(.dina(n6748), .dinb(n6743), .dout(n6749));
  jxor g06686(.dina(n6749), .dinb(n68), .dout(n6750));
  jor  g06687(.dina(n6750), .dinb(n6742), .dout(n6751));
  jand g06688(.dina(n6751), .dinb(n6740), .dout(n6752));
  jnot g06689(.din(n6752), .dout(n6753));
  jxor g06690(.dina(n6505), .dinb(n6497), .dout(n6754));
  jand g06691(.dina(n6754), .dinb(n6753), .dout(n6755));
  jnot g06692(.din(n6755), .dout(n6756));
  jxor g06693(.dina(n6754), .dinb(n6753), .dout(n6757));
  jnot g06694(.din(n6757), .dout(n6758));
  jand g06695(.dina(n5365), .dinb(n4849), .dout(n6759));
  jand g06696(.dina(n5500), .dinb(n1560), .dout(n6760));
  jand g06697(.dina(n5424), .dinb(n1624), .dout(n6761));
  jand g06698(.dina(n5363), .dinb(n1776), .dout(n6762));
  jor  g06699(.dina(n6762), .dinb(n6761), .dout(n6763));
  jor  g06700(.dina(n6763), .dinb(n6760), .dout(n6764));
  jor  g06701(.dina(n6764), .dinb(n6759), .dout(n6765));
  jxor g06702(.dina(n6765), .dinb(n72), .dout(n6766));
  jor  g06703(.dina(n6766), .dinb(n6758), .dout(n6767));
  jand g06704(.dina(n6767), .dinb(n6756), .dout(n6768));
  jnot g06705(.din(n6768), .dout(n6769));
  jxor g06706(.dina(n6577), .dinb(n6576), .dout(n6770));
  jand g06707(.dina(n6770), .dinb(n6769), .dout(n6771));
  jor  g06708(.dina(n6771), .dinb(n6578), .dout(n6772));
  jxor g06709(.dina(n6524), .dinb(n6516), .dout(n6773));
  jand g06710(.dina(n6773), .dinb(n6772), .dout(n6774));
  jnot g06711(.din(n6774), .dout(n6775));
  jxor g06712(.dina(n6773), .dinb(n6772), .dout(n6776));
  jnot g06713(.din(n6776), .dout(n6777));
  jand g06714(.dina(n5693), .dinb(n4026), .dout(n6778));
  jand g06715(.dina(n6131), .dinb(n1076), .dout(n6779));
  jand g06716(.dina(n6209), .dinb(n922), .dout(n6780));
  jand g06717(.dina(n5691), .dinb(n1213), .dout(n6781));
  jor  g06718(.dina(n6781), .dinb(n6780), .dout(n6782));
  jor  g06719(.dina(n6782), .dinb(n6779), .dout(n6783));
  jor  g06720(.dina(n6783), .dinb(n6778), .dout(n6784));
  jxor g06721(.dina(n6784), .dinb(n4247), .dout(n6785));
  jor  g06722(.dina(n6785), .dinb(n6777), .dout(n6786));
  jand g06723(.dina(n6786), .dinb(n6775), .dout(n6787));
  jnot g06724(.din(n6787), .dout(n6788));
  jxor g06725(.dina(n6540), .dinb(n6532), .dout(n6789));
  jand g06726(.dina(n6789), .dinb(n6788), .dout(n6790));
  jnot g06727(.din(n6790), .dout(n6791));
  jxor g06728(.dina(n6789), .dinb(n6788), .dout(n6792));
  jnot g06729(.din(n6792), .dout(n6793));
  jand g06730(.dina(n6340), .dinb(n4752), .dout(n6794));
  jand g06731(.dina(n6556), .dinb(n4451), .dout(n6795));
  jand g06732(.dina(n6338), .dinb(n4358), .dout(n6796));
  jor  g06733(.dina(n6337), .dinb(n6335), .dout(n6797));
  jnot g06734(.din(n6797), .dout(n6798));
  jand g06735(.dina(n6798), .dinb(n4598), .dout(n6799));
  jor  g06736(.dina(n6799), .dinb(n6796), .dout(n6800));
  jor  g06737(.dina(n6800), .dinb(n6795), .dout(n6801));
  jor  g06738(.dina(n6801), .dinb(n6794), .dout(n6802));
  jxor g06739(.dina(n6802), .dinb(n5064), .dout(n6803));
  jor  g06740(.dina(n6803), .dinb(n6793), .dout(n6804));
  jand g06741(.dina(n6804), .dinb(n6791), .dout(n6805));
  jand g06742(.dina(n6340), .dinb(n4636), .dout(n6806));
  jand g06743(.dina(n6338), .dinb(n4451), .dout(n6807));
  jand g06744(.dina(n6556), .dinb(n4598), .dout(n6808));
  jand g06745(.dina(n6798), .dinb(n4631), .dout(n6809));
  jor  g06746(.dina(n6809), .dinb(n6808), .dout(n6810));
  jor  g06747(.dina(n6810), .dinb(n6807), .dout(n6811));
  jor  g06748(.dina(n6811), .dinb(n6806), .dout(n6812));
  jxor g06749(.dina(n6812), .dinb(n5064), .dout(n6813));
  jor  g06750(.dina(n6813), .dinb(n6805), .dout(n6814));
  jxor g06751(.dina(n6813), .dinb(n6805), .dout(n6815));
  jxor g06752(.dina(n6544), .dinb(n6543), .dout(n6816));
  jand g06753(.dina(n6816), .dinb(n6815), .dout(n6817));
  jnot g06754(.din(n6817), .dout(n6818));
  jand g06755(.dina(n6818), .dinb(n6814), .dout(n6819));
  jnot g06756(.din(n6819), .dout(n6820));
  jxor g06757(.dina(n6561), .dinb(n6553), .dout(n6821));
  jand g06758(.dina(n6821), .dinb(n6820), .dout(n6822));
  jxor g06759(.dina(n6821), .dinb(n6820), .dout(n6823));
  jxor g06760(.dina(n6770), .dinb(n6769), .dout(n6824));
  jnot g06761(.din(n6824), .dout(n6825));
  jand g06762(.dina(n5693), .dinb(n4043), .dout(n6826));
  jand g06763(.dina(n6131), .dinb(n1213), .dout(n6827));
  jand g06764(.dina(n5691), .dinb(n1343), .dout(n6828));
  jand g06765(.dina(n6209), .dinb(n1076), .dout(n6829));
  jor  g06766(.dina(n6829), .dinb(n6828), .dout(n6830));
  jor  g06767(.dina(n6830), .dinb(n6827), .dout(n6831));
  jor  g06768(.dina(n6831), .dinb(n6826), .dout(n6832));
  jxor g06769(.dina(n6832), .dinb(n4247), .dout(n6833));
  jor  g06770(.dina(n6833), .dinb(n6825), .dout(n6834));
  jxor g06771(.dina(n6735), .dinb(n6734), .dout(n6835));
  jnot g06772(.din(n6835), .dout(n6836));
  jand g06773(.dina(n5624), .dinb(n75), .dout(n6837));
  jand g06774(.dina(n4745), .dinb(n2237), .dout(n6838));
  jand g06775(.dina(n4918), .dinb(n2128), .dout(n6839));
  jand g06776(.dina(n4933), .dinb(n2067), .dout(n6840));
  jor  g06777(.dina(n6840), .dinb(n6839), .dout(n6841));
  jor  g06778(.dina(n6841), .dinb(n6838), .dout(n6842));
  jor  g06779(.dina(n6842), .dinb(n6837), .dout(n6843));
  jxor g06780(.dina(n6843), .dinb(n68), .dout(n6844));
  jor  g06781(.dina(n6844), .dinb(n6836), .dout(n6845));
  jand g06782(.dina(n6247), .dinb(n4449), .dout(n6846));
  jand g06783(.dina(n4453), .dinb(n2411), .dout(n6847));
  jand g06784(.dina(n4461), .dinb(n2602), .dout(n6848));
  jand g06785(.dina(n4457), .dinb(n2497), .dout(n6849));
  jor  g06786(.dina(n6849), .dinb(n6848), .dout(n6850));
  jor  g06787(.dina(n6850), .dinb(n6847), .dout(n6851));
  jor  g06788(.dina(n6851), .dinb(n6846), .dout(n6852));
  jxor g06789(.dina(n6852), .dinb(n88), .dout(n6853));
  jnot g06790(.din(n6853), .dout(n6854));
  jxor g06791(.dina(n6732), .dinb(n6731), .dout(n6855));
  jand g06792(.dina(n6855), .dinb(n6854), .dout(n6856));
  jnot g06793(.din(n6856), .dout(n6857));
  jxor g06794(.dina(n6855), .dinb(n6854), .dout(n6858));
  jnot g06795(.din(n6858), .dout(n6859));
  jand g06796(.dina(n5607), .dinb(n75), .dout(n6860));
  jand g06797(.dina(n4918), .dinb(n2237), .dout(n6861));
  jand g06798(.dina(n4745), .dinb(n2343), .dout(n6862));
  jand g06799(.dina(n4933), .dinb(n2128), .dout(n6863));
  jor  g06800(.dina(n6863), .dinb(n6862), .dout(n6864));
  jor  g06801(.dina(n6864), .dinb(n6861), .dout(n6865));
  jor  g06802(.dina(n6865), .dinb(n6860), .dout(n6866));
  jxor g06803(.dina(n6866), .dinb(n68), .dout(n6867));
  jor  g06804(.dina(n6867), .dinb(n6859), .dout(n6868));
  jand g06805(.dina(n6868), .dinb(n6857), .dout(n6869));
  jnot g06806(.din(n6869), .dout(n6870));
  jxor g06807(.dina(n6844), .dinb(n6836), .dout(n6871));
  jand g06808(.dina(n6871), .dinb(n6870), .dout(n6872));
  jnot g06809(.din(n6872), .dout(n6873));
  jand g06810(.dina(n6873), .dinb(n6845), .dout(n6874));
  jnot g06811(.din(n6874), .dout(n6875));
  jxor g06812(.dina(n6750), .dinb(n6742), .dout(n6876));
  jand g06813(.dina(n6876), .dinb(n6875), .dout(n6877));
  jnot g06814(.din(n6877), .dout(n6878));
  jxor g06815(.dina(n6876), .dinb(n6875), .dout(n6879));
  jnot g06816(.din(n6879), .dout(n6880));
  jand g06817(.dina(n5365), .dinb(n5075), .dout(n6881));
  jand g06818(.dina(n5500), .dinb(n1624), .dout(n6882));
  jand g06819(.dina(n5424), .dinb(n1776), .dout(n6883));
  jand g06820(.dina(n5363), .dinb(n1862), .dout(n6884));
  jor  g06821(.dina(n6884), .dinb(n6883), .dout(n6885));
  jor  g06822(.dina(n6885), .dinb(n6882), .dout(n6886));
  jor  g06823(.dina(n6886), .dinb(n6881), .dout(n6887));
  jxor g06824(.dina(n6887), .dinb(n72), .dout(n6888));
  jor  g06825(.dina(n6888), .dinb(n6880), .dout(n6889));
  jand g06826(.dina(n6889), .dinb(n6878), .dout(n6890));
  jnot g06827(.din(n6890), .dout(n6891));
  jxor g06828(.dina(n6766), .dinb(n6758), .dout(n6892));
  jand g06829(.dina(n6892), .dinb(n6891), .dout(n6893));
  jnot g06830(.din(n6893), .dout(n6894));
  jxor g06831(.dina(n6892), .dinb(n6891), .dout(n6895));
  jnot g06832(.din(n6895), .dout(n6896));
  jand g06833(.dina(n5693), .dinb(n4772), .dout(n6897));
  jand g06834(.dina(n6209), .dinb(n1213), .dout(n6898));
  jand g06835(.dina(n6131), .dinb(n1343), .dout(n6899));
  jand g06836(.dina(n5691), .dinb(n1445), .dout(n6900));
  jor  g06837(.dina(n6900), .dinb(n6899), .dout(n6901));
  jor  g06838(.dina(n6901), .dinb(n6898), .dout(n6902));
  jor  g06839(.dina(n6902), .dinb(n6897), .dout(n6903));
  jxor g06840(.dina(n6903), .dinb(n4247), .dout(n6904));
  jor  g06841(.dina(n6904), .dinb(n6896), .dout(n6905));
  jand g06842(.dina(n6905), .dinb(n6894), .dout(n6906));
  jnot g06843(.din(n6906), .dout(n6907));
  jxor g06844(.dina(n6833), .dinb(n6825), .dout(n6908));
  jand g06845(.dina(n6908), .dinb(n6907), .dout(n6909));
  jnot g06846(.din(n6909), .dout(n6910));
  jand g06847(.dina(n6910), .dinb(n6834), .dout(n6911));
  jnot g06848(.din(n6911), .dout(n6912));
  jxor g06849(.dina(n6785), .dinb(n6777), .dout(n6913));
  jand g06850(.dina(n6913), .dinb(n6912), .dout(n6914));
  jnot g06851(.din(n6914), .dout(n6915));
  jxor g06852(.dina(n6913), .dinb(n6912), .dout(n6916));
  jnot g06853(.din(n6916), .dout(n6917));
  jand g06854(.dina(n6340), .dinb(n4446), .dout(n6918));
  jand g06855(.dina(n6798), .dinb(n4451), .dout(n6919));
  jand g06856(.dina(n6556), .dinb(n4358), .dout(n6920));
  jand g06857(.dina(n6338), .dinb(n3853), .dout(n6921));
  jor  g06858(.dina(n6921), .dinb(n6920), .dout(n6922));
  jor  g06859(.dina(n6922), .dinb(n6919), .dout(n6923));
  jor  g06860(.dina(n6923), .dinb(n6918), .dout(n6924));
  jxor g06861(.dina(n6924), .dinb(n5064), .dout(n6925));
  jor  g06862(.dina(n6925), .dinb(n6917), .dout(n6926));
  jand g06863(.dina(n6926), .dinb(n6915), .dout(n6927));
  jxor g06864(.dina(\a[12] ), .dinb(\a[11] ), .dout(n6928));
  jnot g06865(.din(n6928), .dout(n6929));
  jxor g06866(.dina(\a[13] ), .dinb(\a[12] ), .dout(n6930));
  jnot g06867(.din(n6930), .dout(n6931));
  jand g06868(.dina(n6931), .dinb(n6929), .dout(n6932));
  jxor g06869(.dina(\a[14] ), .dinb(\a[13] ), .dout(n6933));
  jand g06870(.dina(n6933), .dinb(n6932), .dout(n6934));
  jnot g06871(.din(n6934), .dout(n6935));
  jand g06872(.dina(n6933), .dinb(n6928), .dout(n6936));
  jnot g06873(.din(n6936), .dout(n6937));
  jor  g06874(.dina(n6937), .dinb(n4728), .dout(n6938));
  jand g06875(.dina(n6938), .dinb(n6935), .dout(n6939));
  jor  g06876(.dina(n6939), .dinb(n4630), .dout(n6940));
  jxor g06877(.dina(n6940), .dinb(\a[14] ), .dout(n6941));
  jor  g06878(.dina(n6941), .dinb(n6927), .dout(n6942));
  jxor g06879(.dina(n6941), .dinb(n6927), .dout(n6943));
  jxor g06880(.dina(n6803), .dinb(n6793), .dout(n6944));
  jand g06881(.dina(n6944), .dinb(n6943), .dout(n6945));
  jnot g06882(.din(n6945), .dout(n6946));
  jand g06883(.dina(n6946), .dinb(n6942), .dout(n6947));
  jnot g06884(.din(n6947), .dout(n6948));
  jxor g06885(.dina(n6816), .dinb(n6815), .dout(n6949));
  jand g06886(.dina(n6949), .dinb(n6948), .dout(n6950));
  jxor g06887(.dina(n6949), .dinb(n6948), .dout(n6951));
  jand g06888(.dina(n6340), .dinb(n4545), .dout(n6952));
  jand g06889(.dina(n6556), .dinb(n3853), .dout(n6953));
  jand g06890(.dina(n6798), .dinb(n4358), .dout(n6954));
  jand g06891(.dina(n6338), .dinb(n922), .dout(n6955));
  jor  g06892(.dina(n6955), .dinb(n6954), .dout(n6956));
  jor  g06893(.dina(n6956), .dinb(n6953), .dout(n6957));
  jor  g06894(.dina(n6957), .dinb(n6952), .dout(n6958));
  jxor g06895(.dina(n6958), .dinb(n5064), .dout(n6959));
  jnot g06896(.din(n6959), .dout(n6960));
  jxor g06897(.dina(n6908), .dinb(n6907), .dout(n6961));
  jand g06898(.dina(n6961), .dinb(n6960), .dout(n6962));
  jand g06899(.dina(n5365), .dinb(n5092), .dout(n6963));
  jand g06900(.dina(n5500), .dinb(n1776), .dout(n6964));
  jand g06901(.dina(n5424), .dinb(n1862), .dout(n6965));
  jand g06902(.dina(n5363), .dinb(n1956), .dout(n6966));
  jor  g06903(.dina(n6966), .dinb(n6965), .dout(n6967));
  jor  g06904(.dina(n6967), .dinb(n6964), .dout(n6968));
  jor  g06905(.dina(n6968), .dinb(n6963), .dout(n6969));
  jxor g06906(.dina(n6969), .dinb(n72), .dout(n6970));
  jnot g06907(.din(n6970), .dout(n6971));
  jxor g06908(.dina(n6871), .dinb(n6870), .dout(n6972));
  jand g06909(.dina(n6972), .dinb(n6971), .dout(n6973));
  jxor g06910(.dina(n6698), .dinb(n6697), .dout(n6974));
  jnot g06911(.din(n6974), .dout(n6975));
  jxor g06912(.dina(n3704), .dinb(n3703), .dout(n6976));
  jor  g06913(.dina(n6976), .dinb(n6463), .dout(n6977));
  jand g06914(.dina(n3855), .dinb(n2867), .dout(n6978));
  jand g06915(.dina(n3851), .dinb(n2991), .dout(n6979));
  jand g06916(.dina(n3858), .dinb(n2954), .dout(n6980));
  jor  g06917(.dina(n6980), .dinb(n6979), .dout(n6981));
  jor  g06918(.dina(n6981), .dinb(n6978), .dout(n6982));
  jnot g06919(.din(n6982), .dout(n6983));
  jand g06920(.dina(n6983), .dinb(n6977), .dout(n6984));
  jor  g06921(.dina(n6984), .dinb(n6975), .dout(n6985));
  jxor g06922(.dina(n6693), .dinb(n6692), .dout(n6986));
  jnot g06923(.din(n6986), .dout(n6987));
  jxor g06924(.dina(n3700), .dinb(n3699), .dout(n6988));
  jor  g06925(.dina(n6988), .dinb(n6463), .dout(n6989));
  jand g06926(.dina(n3851), .dinb(n3086), .dout(n6990));
  jand g06927(.dina(n3855), .dinb(n2954), .dout(n6991));
  jand g06928(.dina(n3858), .dinb(n2991), .dout(n6992));
  jor  g06929(.dina(n6992), .dinb(n6991), .dout(n6993));
  jor  g06930(.dina(n6993), .dinb(n6990), .dout(n6994));
  jnot g06931(.din(n6994), .dout(n6995));
  jand g06932(.dina(n6995), .dinb(n6989), .dout(n6996));
  jor  g06933(.dina(n6996), .dinb(n6987), .dout(n6997));
  jand g06934(.dina(n1346), .dinb(n692), .dout(n6998));
  jand g06935(.dina(n6998), .dinb(n1269), .dout(n6999));
  jand g06936(.dina(n6999), .dinb(n2366), .dout(n7000));
  jand g06937(.dina(n7000), .dinb(n327), .dout(n7001));
  jand g06938(.dina(n5903), .dinb(n557), .dout(n7002));
  jand g06939(.dina(n7002), .dinb(n1222), .dout(n7003));
  jand g06940(.dina(n529), .dinb(n143), .dout(n7004));
  jand g06941(.dina(n7004), .dinb(n1295), .dout(n7005));
  jand g06942(.dina(n2722), .dinb(n1199), .dout(n7006));
  jand g06943(.dina(n7006), .dinb(n7005), .dout(n7007));
  jand g06944(.dina(n2538), .dinb(n130), .dout(n7008));
  jand g06945(.dina(n1663), .dinb(n1598), .dout(n7009));
  jand g06946(.dina(n7009), .dinb(n7008), .dout(n7010));
  jand g06947(.dina(n7010), .dinb(n7007), .dout(n7011));
  jand g06948(.dina(n7011), .dinb(n7003), .dout(n7012));
  jand g06949(.dina(n7012), .dinb(n7001), .dout(n7013));
  jand g06950(.dina(n7013), .dinb(n5229), .dout(n7014));
  jand g06951(.dina(n3450), .dinb(n2228), .dout(n7015));
  jand g06952(.dina(n5259), .dinb(n2041), .dout(n7016));
  jand g06953(.dina(n7016), .dinb(n7015), .dout(n7017));
  jand g06954(.dina(n865), .dinb(n817), .dout(n7018));
  jand g06955(.dina(n7018), .dinb(n396), .dout(n7019));
  jand g06956(.dina(n1014), .dinb(n897), .dout(n7020));
  jand g06957(.dina(n7020), .dinb(n1847), .dout(n7021));
  jand g06958(.dina(n7021), .dinb(n7019), .dout(n7022));
  jand g06959(.dina(n7022), .dinb(n7017), .dout(n7023));
  jand g06960(.dina(n5549), .dinb(n1334), .dout(n7024));
  jand g06961(.dina(n7024), .dinb(n506), .dout(n7025));
  jand g06962(.dina(n7025), .dinb(n5152), .dout(n7026));
  jand g06963(.dina(n7026), .dinb(n7023), .dout(n7027));
  jand g06964(.dina(n7027), .dinb(n2670), .dout(n7028));
  jand g06965(.dina(n7028), .dinb(n5258), .dout(n7029));
  jand g06966(.dina(n7029), .dinb(n7014), .dout(n7030));
  jxor g06967(.dina(n3692), .dinb(n3691), .dout(n7031));
  jor  g06968(.dina(n7031), .dinb(n6463), .dout(n7032));
  jand g06969(.dina(n3855), .dinb(n3086), .dout(n7033));
  jand g06970(.dina(n3851), .dinb(n3275), .dout(n7034));
  jand g06971(.dina(n3858), .dinb(n3183), .dout(n7035));
  jor  g06972(.dina(n7035), .dinb(n7034), .dout(n7036));
  jor  g06973(.dina(n7036), .dinb(n7033), .dout(n7037));
  jnot g06974(.din(n7037), .dout(n7038));
  jand g06975(.dina(n7038), .dinb(n7032), .dout(n7039));
  jor  g06976(.dina(n7039), .dinb(n7030), .dout(n7040));
  jand g06977(.dina(n2878), .dinb(n2034), .dout(n7041));
  jand g06978(.dina(n7041), .dinb(n1474), .dout(n7042));
  jand g06979(.dina(n375), .dinb(n337), .dout(n7043));
  jand g06980(.dina(n7043), .dinb(n1475), .dout(n7044));
  jand g06981(.dina(n7044), .dinb(n2526), .dout(n7045));
  jand g06982(.dina(n3500), .dinb(n2538), .dout(n7046));
  jand g06983(.dina(n1829), .dinb(n1088), .dout(n7047));
  jand g06984(.dina(n7047), .dinb(n7046), .dout(n7048));
  jand g06985(.dina(n7048), .dinb(n7045), .dout(n7049));
  jand g06986(.dina(n7049), .dinb(n7042), .dout(n7050));
  jand g06987(.dina(n646), .dinb(n409), .dout(n7051));
  jand g06988(.dina(n7051), .dinb(n2547), .dout(n7052));
  jand g06989(.dina(n7052), .dinb(n834), .dout(n7053));
  jand g06990(.dina(n712), .dinb(n221), .dout(n7054));
  jand g06991(.dina(n7054), .dinb(n2053), .dout(n7055));
  jand g06992(.dina(n7055), .dinb(n5569), .dout(n7056));
  jand g06993(.dina(n7056), .dinb(n7053), .dout(n7057));
  jand g06994(.dina(n7057), .dinb(n5789), .dout(n7058));
  jand g06995(.dina(n7058), .dinb(n7050), .dout(n7059));
  jand g06996(.dina(n635), .dinb(n340), .dout(n7060));
  jand g06997(.dina(n7060), .dinb(n770), .dout(n7061));
  jand g06998(.dina(n5879), .dinb(n1197), .dout(n7062));
  jand g06999(.dina(n7062), .dinb(n7061), .dout(n7063));
  jand g07000(.dina(n1264), .dinb(n174), .dout(n7064));
  jand g07001(.dina(n7064), .dinb(n439), .dout(n7065));
  jand g07002(.dina(n7065), .dinb(n5749), .dout(n7066));
  jand g07003(.dina(n7066), .dinb(n7063), .dout(n7067));
  jand g07004(.dina(n2659), .dinb(n355), .dout(n7068));
  jand g07005(.dina(n847), .dinb(n113), .dout(n7069));
  jand g07006(.dina(n7069), .dinb(n3445), .dout(n7070));
  jand g07007(.dina(n7070), .dinb(n7068), .dout(n7071));
  jand g07008(.dina(n7071), .dinb(n5035), .dout(n7072));
  jand g07009(.dina(n7072), .dinb(n7067), .dout(n7073));
  jand g07010(.dina(n7073), .dinb(n1420), .dout(n7074));
  jand g07011(.dina(n7074), .dinb(n7059), .dout(n7075));
  jxor g07012(.dina(n3688), .dinb(n3687), .dout(n7076));
  jor  g07013(.dina(n7076), .dinb(n6463), .dout(n7077));
  jand g07014(.dina(n3858), .dinb(n3275), .dout(n7078));
  jand g07015(.dina(n3855), .dinb(n3183), .dout(n7079));
  jand g07016(.dina(n3851), .dinb(n3359), .dout(n7080));
  jor  g07017(.dina(n7080), .dinb(n7079), .dout(n7081));
  jor  g07018(.dina(n7081), .dinb(n7078), .dout(n7082));
  jnot g07019(.din(n7082), .dout(n7083));
  jand g07020(.dina(n7083), .dinb(n7077), .dout(n7084));
  jor  g07021(.dina(n7084), .dinb(n7075), .dout(n7085));
  jand g07022(.dina(n619), .dinb(n205), .dout(n7086));
  jand g07023(.dina(n7086), .dinb(n1144), .dout(n7087));
  jand g07024(.dina(n7087), .dinb(n2977), .dout(n7088));
  jand g07025(.dina(n177), .dinb(n143), .dout(n7089));
  jand g07026(.dina(n382), .dinb(n146), .dout(n7090));
  jand g07027(.dina(n7090), .dinb(n7089), .dout(n7091));
  jand g07028(.dina(n1231), .dinb(n427), .dout(n7092));
  jand g07029(.dina(n7092), .dinb(n1035), .dout(n7093));
  jand g07030(.dina(n7093), .dinb(n2359), .dout(n7094));
  jand g07031(.dina(n7094), .dinb(n7091), .dout(n7095));
  jand g07032(.dina(n7095), .dinb(n7088), .dout(n7096));
  jand g07033(.dina(n751), .dinb(n405), .dout(n7097));
  jand g07034(.dina(n7097), .dinb(n355), .dout(n7098));
  jand g07035(.dina(n3046), .dinb(n1432), .dout(n7099));
  jand g07036(.dina(n7099), .dinb(n7098), .dout(n7100));
  jand g07037(.dina(n913), .dinb(n874), .dout(n7101));
  jand g07038(.dina(n7101), .dinb(n486), .dout(n7102));
  jand g07039(.dina(n7102), .dinb(n1822), .dout(n7103));
  jand g07040(.dina(n7103), .dinb(n7100), .dout(n7104));
  jand g07041(.dina(n3804), .dinb(n3111), .dout(n7105));
  jand g07042(.dina(n7105), .dinb(n7104), .dout(n7106));
  jand g07043(.dina(n7106), .dinb(n7096), .dout(n7107));
  jand g07044(.dina(n897), .dinb(n499), .dout(n7108));
  jand g07045(.dina(n7108), .dinb(n367), .dout(n7109));
  jand g07046(.dina(n566), .dinb(n434), .dout(n7110));
  jand g07047(.dina(n847), .dinb(n574), .dout(n7111));
  jand g07048(.dina(n7111), .dinb(n7110), .dout(n7112));
  jand g07049(.dina(n7112), .dinb(n7109), .dout(n7113));
  jand g07050(.dina(n7113), .dinb(n2456), .dout(n7114));
  jand g07051(.dina(n786), .dinb(n280), .dout(n7115));
  jand g07052(.dina(n7115), .dinb(n290), .dout(n7116));
  jand g07053(.dina(n7116), .dinb(n2620), .dout(n7117));
  jand g07054(.dina(n492), .dinb(n395), .dout(n7118));
  jand g07055(.dina(n7118), .dinb(n563), .dout(n7119));
  jand g07056(.dina(n2240), .dinb(n802), .dout(n7120));
  jand g07057(.dina(n7120), .dinb(n7119), .dout(n7121));
  jand g07058(.dina(n7121), .dinb(n7117), .dout(n7122));
  jand g07059(.dina(n330), .dinb(n174), .dout(n7123));
  jand g07060(.dina(n7123), .dinb(n4315), .dout(n7124));
  jand g07061(.dina(n7124), .dinb(n5882), .dout(n7125));
  jand g07062(.dina(n7125), .dinb(n7122), .dout(n7126));
  jand g07063(.dina(n7126), .dinb(n7114), .dout(n7127));
  jand g07064(.dina(n7127), .dinb(n5954), .dout(n7128));
  jand g07065(.dina(n7128), .dinb(n7107), .dout(n7129));
  jnot g07066(.din(n3685), .dout(n7130));
  jxor g07067(.dina(n7130), .dinb(n3683), .dout(n7131));
  jor  g07068(.dina(n7131), .dinb(n6463), .dout(n7132));
  jand g07069(.dina(n3855), .dinb(n3275), .dout(n7133));
  jand g07070(.dina(n3858), .dinb(n3359), .dout(n7134));
  jand g07071(.dina(n3851), .dinb(n3411), .dout(n7135));
  jor  g07072(.dina(n7135), .dinb(n7134), .dout(n7136));
  jor  g07073(.dina(n7136), .dinb(n7133), .dout(n7137));
  jnot g07074(.din(n7137), .dout(n7138));
  jand g07075(.dina(n7138), .dinb(n7132), .dout(n7139));
  jor  g07076(.dina(n7139), .dinb(n7129), .dout(n7140));
  jand g07077(.dina(n1025), .dinb(n818), .dout(n7141));
  jand g07078(.dina(n7141), .dinb(n254), .dout(n7142));
  jand g07079(.dina(n330), .dinb(n324), .dout(n7143));
  jand g07080(.dina(n7143), .dinb(n671), .dout(n7144));
  jand g07081(.dina(n1346), .dinb(n1597), .dout(n7145));
  jand g07082(.dina(n924), .dinb(n759), .dout(n7146));
  jand g07083(.dina(n7146), .dinb(n7145), .dout(n7147));
  jand g07084(.dina(n7147), .dinb(n7144), .dout(n7148));
  jand g07085(.dina(n7148), .dinb(n4833), .dout(n7149));
  jand g07086(.dina(n7149), .dinb(n7142), .dout(n7150));
  jand g07087(.dina(n614), .dinb(n757), .dout(n7151));
  jand g07088(.dina(n7151), .dinb(n1104), .dout(n7152));
  jand g07089(.dina(n860), .dinb(n527), .dout(n7153));
  jand g07090(.dina(n819), .dinb(n716), .dout(n7154));
  jand g07091(.dina(n7154), .dinb(n7153), .dout(n7155));
  jand g07092(.dina(n7155), .dinb(n7152), .dout(n7156));
  jand g07093(.dina(n3938), .dinb(n2446), .dout(n7157));
  jand g07094(.dina(n7157), .dinb(n7156), .dout(n7158));
  jand g07095(.dina(n1268), .dinb(n103), .dout(n7159));
  jand g07096(.dina(n7159), .dinb(n268), .dout(n7160));
  jand g07097(.dina(n305), .dinb(n230), .dout(n7161));
  jand g07098(.dina(n7161), .dinb(n2261), .dout(n7162));
  jand g07099(.dina(n7162), .dinb(n7160), .dout(n7163));
  jand g07100(.dina(n433), .dinb(n277), .dout(n7164));
  jand g07101(.dina(n1986), .dinb(n880), .dout(n7165));
  jand g07102(.dina(n7165), .dinb(n7164), .dout(n7166));
  jand g07103(.dina(n532), .dinb(n177), .dout(n7167));
  jand g07104(.dina(n7167), .dinb(n5153), .dout(n7168));
  jand g07105(.dina(n4667), .dinb(n858), .dout(n7169));
  jand g07106(.dina(n7169), .dinb(n7168), .dout(n7170));
  jand g07107(.dina(n7170), .dinb(n7166), .dout(n7171));
  jand g07108(.dina(n7171), .dinb(n7163), .dout(n7172));
  jand g07109(.dina(n7172), .dinb(n7158), .dout(n7173));
  jand g07110(.dina(n7173), .dinb(n7150), .dout(n7174));
  jand g07111(.dina(n7174), .dinb(n3030), .dout(n7175));
  jnot g07112(.din(n3681), .dout(n7176));
  jxor g07113(.dina(n7176), .dinb(n3680), .dout(n7177));
  jor  g07114(.dina(n7177), .dinb(n6463), .dout(n7178));
  jnot g07115(.din(n3416), .dout(n7179));
  jor  g07116(.dina(n1614), .dinb(n3318), .dout(n7180));
  jnot g07117(.din(n3417), .dout(n7181));
  jor  g07118(.dina(n7181), .dinb(n7180), .dout(n7182));
  jnot g07119(.din(n82), .dout(n7183));
  jor  g07120(.dina(n358), .dinb(n7183), .dout(n7184));
  jor  g07121(.dina(n7184), .dinb(n1933), .dout(n7185));
  jor  g07122(.dina(n7185), .dinb(n7182), .dout(n7186));
  jor  g07123(.dina(n875), .dinb(n3210), .dout(n7187));
  jor  g07124(.dina(n7187), .dinb(n881), .dout(n7188));
  jor  g07125(.dina(n3425), .dinb(n7188), .dout(n7189));
  jor  g07126(.dina(n7189), .dinb(n7186), .dout(n7190));
  jor  g07127(.dina(n7190), .dinb(n7179), .dout(n7191));
  jnot g07128(.din(n3431), .dout(n7192));
  jnot g07129(.din(n3433), .dout(n7193));
  jor  g07130(.dina(n1371), .dinb(n196), .dout(n7194));
  jor  g07131(.dina(n7194), .dinb(n1215), .dout(n7195));
  jor  g07132(.dina(n7195), .dinb(n7193), .dout(n7196));
  jor  g07133(.dina(n7196), .dinb(n7192), .dout(n7197));
  jor  g07134(.dina(n841), .dinb(n1683), .dout(n7198));
  jor  g07135(.dina(n7198), .dinb(n201), .dout(n7199));
  jor  g07136(.dina(n3667), .dinb(n1374), .dout(n7200));
  jor  g07137(.dina(n7200), .dinb(n2070), .dout(n7201));
  jand g07138(.dina(n338), .dinb(n125), .dout(n7202));
  jor  g07139(.dina(n1746), .dinb(n7202), .dout(n7203));
  jand g07140(.dina(n344), .dinb(n97), .dout(n7204));
  jor  g07141(.dina(n7204), .dinb(n2466), .dout(n7205));
  jor  g07142(.dina(n7205), .dinb(n7203), .dout(n7206));
  jor  g07143(.dina(n7206), .dinb(n7201), .dout(n7207));
  jor  g07144(.dina(n7207), .dinb(n7199), .dout(n7208));
  jnot g07145(.din(n527), .dout(n7209));
  jor  g07146(.dina(n7209), .dinb(n119), .dout(n7210));
  jand g07147(.dina(n147), .dinb(n300), .dout(n7211));
  jand g07148(.dina(n272), .dinb(n147), .dout(n7212));
  jor  g07149(.dina(n7212), .dinb(n7211), .dout(n7213));
  jand g07150(.dina(n200), .dinb(n300), .dout(n7214));
  jand g07151(.dina(n389), .dinb(n159), .dout(n7215));
  jor  g07152(.dina(n7215), .dinb(n7214), .dout(n7216));
  jor  g07153(.dina(n7216), .dinb(n7213), .dout(n7217));
  jor  g07154(.dina(n7217), .dinb(n7210), .dout(n7218));
  jand g07155(.dina(n250), .dinb(n172), .dout(n7219));
  jand g07156(.dina(n172), .dinb(n159), .dout(n7220));
  jor  g07157(.dina(n7220), .dinb(n7219), .dout(n7221));
  jand g07158(.dina(n155), .dinb(n203), .dout(n7222));
  jor  g07159(.dina(n7222), .dinb(n3651), .dout(n7223));
  jor  g07160(.dina(n7223), .dinb(n7221), .dout(n7224));
  jand g07161(.dina(n222), .dinb(n125), .dout(n7225));
  jor  g07162(.dina(n3208), .dinb(n7225), .dout(n7226));
  jand g07163(.dina(n172), .dinb(n215), .dout(n7227));
  jor  g07164(.dina(n775), .dinb(n7227), .dout(n7228));
  jor  g07165(.dina(n7228), .dinb(n7226), .dout(n7229));
  jor  g07166(.dina(n7229), .dinb(n7224), .dout(n7230));
  jor  g07167(.dina(n7230), .dinb(n7218), .dout(n7231));
  jor  g07168(.dina(n7231), .dinb(n7208), .dout(n7232));
  jor  g07169(.dina(n7232), .dinb(n7197), .dout(n7233));
  jor  g07170(.dina(n7233), .dinb(n7191), .dout(n7234));
  jnot g07171(.din(n2327), .dout(n7235));
  jnot g07172(.din(n443), .dout(n7236));
  jor  g07173(.dina(n762), .dinb(n7236), .dout(n7237));
  jnot g07174(.din(n1760), .dout(n7238));
  jor  g07175(.dina(n7238), .dinb(n7237), .dout(n7239));
  jor  g07176(.dina(n7239), .dinb(n7235), .dout(n7240));
  jor  g07177(.dina(n2336), .dinb(n7240), .dout(n7241));
  jand g07178(.dina(n116), .dinb(n106), .dout(n7242));
  jor  g07179(.dina(n7242), .dinb(n1403), .dout(n7243));
  jor  g07180(.dina(n3341), .dinb(n660), .dout(n7244));
  jor  g07181(.dina(n7244), .dinb(n7243), .dout(n7245));
  jand g07182(.dina(n195), .dinb(n128), .dout(n7246));
  jor  g07183(.dina(n7246), .dinb(n1887), .dout(n7247));
  jand g07184(.dina(n344), .dinb(n219), .dout(n7248));
  jor  g07185(.dina(n3207), .dinb(n7248), .dout(n7249));
  jor  g07186(.dina(n7249), .dinb(n7247), .dout(n7250));
  jor  g07187(.dina(n7250), .dinb(n7245), .dout(n7251));
  jand g07188(.dina(n195), .dinb(n147), .dout(n7252));
  jor  g07189(.dina(n7252), .dinb(n3338), .dout(n7253));
  jor  g07190(.dina(n7253), .dinb(n453), .dout(n7254));
  jand g07191(.dina(n215), .dinb(n128), .dout(n7255));
  jand g07192(.dina(n236), .dinb(n155), .dout(n7256));
  jor  g07193(.dina(n7256), .dinb(n7255), .dout(n7257));
  jor  g07194(.dina(n7257), .dinb(n261), .dout(n7258));
  jor  g07195(.dina(n7258), .dinb(n7254), .dout(n7259));
  jor  g07196(.dina(n7259), .dinb(n7251), .dout(n7260));
  jand g07197(.dina(n232), .dinb(n125), .dout(n7261));
  jand g07198(.dina(n222), .dinb(n219), .dout(n7262));
  jor  g07199(.dina(n7262), .dinb(n7261), .dout(n7263));
  jor  g07200(.dina(n7263), .dinb(n3348), .dout(n7264));
  jor  g07201(.dina(n3468), .dinb(n7264), .dout(n7265));
  jand g07202(.dina(n338), .dinb(n159), .dout(n7266));
  jor  g07203(.dina(n3196), .dinb(n7266), .dout(n7267));
  jand g07204(.dina(n250), .dinb(n203), .dout(n7268));
  jor  g07205(.dina(n7268), .dinb(n3315), .dout(n7269));
  jor  g07206(.dina(n7269), .dinb(n7267), .dout(n7270));
  jor  g07207(.dina(n7270), .dinb(n3321), .dout(n7271));
  jor  g07208(.dina(n7271), .dinb(n7265), .dout(n7272));
  jor  g07209(.dina(n7272), .dinb(n7260), .dout(n7273));
  jor  g07210(.dina(n7273), .dinb(n7241), .dout(n7274));
  jnot g07211(.din(n3477), .dout(n7275));
  jor  g07212(.dina(n7275), .dinb(n1610), .dout(n7276));
  jand g07213(.dina(n155), .dinb(n101), .dout(n7277));
  jor  g07214(.dina(n7277), .dinb(n1377), .dout(n7278));
  jor  g07215(.dina(n7278), .dinb(n573), .dout(n7279));
  jor  g07216(.dina(n7279), .dinb(n3482), .dout(n7280));
  jor  g07217(.dina(n7280), .dinb(n3480), .dout(n7281));
  jor  g07218(.dina(n7281), .dinb(n7276), .dout(n7282));
  jnot g07219(.din(n396), .dout(n7283));
  jor  g07220(.dina(n825), .dinb(n7283), .dout(n7284));
  jand g07221(.dina(n155), .dinb(n106), .dout(n7285));
  jor  g07222(.dina(n7285), .dinb(n1055), .dout(n7286));
  jor  g07223(.dina(n7286), .dinb(n1717), .dout(n7287));
  jor  g07224(.dina(n7287), .dinb(n7284), .dout(n7288));
  jor  g07225(.dina(n7288), .dinb(n3488), .dout(n7289));
  jand g07226(.dina(n236), .dinb(n159), .dout(n7290));
  jor  g07227(.dina(n7290), .dinb(n1396), .dout(n7291));
  jand g07228(.dina(n272), .dinb(n118), .dout(n7292));
  jor  g07229(.dina(n1706), .dinb(n7292), .dout(n7293));
  jor  g07230(.dina(n7293), .dinb(n7291), .dout(n7294));
  jor  g07231(.dina(n3371), .dinb(n3340), .dout(n7295));
  jor  g07232(.dina(n3314), .dinb(n7295), .dout(n7296));
  jor  g07233(.dina(n7296), .dinb(n7294), .dout(n7297));
  jand g07234(.dina(n219), .dinb(n128), .dout(n7298));
  jand g07235(.dina(n195), .dinb(n344), .dout(n7299));
  jor  g07236(.dina(n7299), .dinb(n7298), .dout(n7300));
  jand g07237(.dina(n338), .dinb(n182), .dout(n7301));
  jor  g07238(.dina(n774), .dinb(n7301), .dout(n7302));
  jor  g07239(.dina(n7302), .dinb(n7300), .dout(n7303));
  jand g07240(.dina(n159), .dinb(n147), .dout(n7304));
  jor  g07241(.dina(n597), .dinb(n3365), .dout(n7305));
  jor  g07242(.dina(n7305), .dinb(n7304), .dout(n7306));
  jor  g07243(.dina(n7306), .dinb(n7303), .dout(n7307));
  jor  g07244(.dina(n7307), .dinb(n7297), .dout(n7308));
  jand g07245(.dina(n172), .dinb(n155), .dout(n7309));
  jor  g07246(.dina(n3382), .dinb(n3370), .dout(n7310));
  jor  g07247(.dina(n7310), .dinb(n7309), .dout(n7311));
  jor  g07248(.dina(n7311), .dinb(n3307), .dout(n7312));
  jand g07249(.dina(n389), .dinb(n219), .dout(n7313));
  jor  g07250(.dina(n1684), .dinb(n7313), .dout(n7314));
  jor  g07251(.dina(n1367), .dinb(n1311), .dout(n7315));
  jand g07252(.dina(n272), .dinb(n200), .dout(n7316));
  jand g07253(.dina(n278), .dinb(n315), .dout(n7317));
  jor  g07254(.dina(n7317), .dinb(n7316), .dout(n7318));
  jor  g07255(.dina(n7318), .dinb(n7315), .dout(n7319));
  jor  g07256(.dina(n7319), .dinb(n7314), .dout(n7320));
  jor  g07257(.dina(n7320), .dinb(n7312), .dout(n7321));
  jor  g07258(.dina(n7321), .dinb(n7308), .dout(n7322));
  jor  g07259(.dina(n7322), .dinb(n7289), .dout(n7323));
  jor  g07260(.dina(n7323), .dinb(n7282), .dout(n7324));
  jor  g07261(.dina(n7324), .dinb(n7274), .dout(n7325));
  jor  g07262(.dina(n7325), .dinb(n7234), .dout(n7326));
  jand g07263(.dina(n3851), .dinb(n7326), .dout(n7327));
  jand g07264(.dina(n3855), .dinb(n3359), .dout(n7328));
  jand g07265(.dina(n3858), .dinb(n3411), .dout(n7329));
  jor  g07266(.dina(n7329), .dinb(n7328), .dout(n7330));
  jor  g07267(.dina(n7330), .dinb(n7327), .dout(n7331));
  jnot g07268(.din(n7331), .dout(n7332));
  jand g07269(.dina(n7332), .dinb(n7178), .dout(n7333));
  jor  g07270(.dina(n7333), .dinb(n7175), .dout(n7334));
  jand g07271(.dina(n805), .dinb(n503), .dout(n7335));
  jand g07272(.dina(n1641), .dinb(n255), .dout(n7336));
  jand g07273(.dina(n7336), .dinb(n7335), .dout(n7337));
  jand g07274(.dina(n778), .dinb(n494), .dout(n7338));
  jand g07275(.dina(n7338), .dinb(n820), .dout(n7339));
  jand g07276(.dina(n7339), .dinb(n3644), .dout(n7340));
  jand g07277(.dina(n7340), .dinb(n7337), .dout(n7341));
  jand g07278(.dina(n1285), .dinb(n1197), .dout(n7342));
  jand g07279(.dina(n1846), .dinb(n1506), .dout(n7343));
  jand g07280(.dina(n7343), .dinb(n7342), .dout(n7344));
  jand g07281(.dina(n817), .dinb(n751), .dout(n7345));
  jand g07282(.dina(n427), .dinb(n329), .dout(n7346));
  jand g07283(.dina(n7346), .dinb(n7345), .dout(n7347));
  jand g07284(.dina(n4494), .dinb(n868), .dout(n7348));
  jand g07285(.dina(n7348), .dinb(n7347), .dout(n7349));
  jand g07286(.dina(n7349), .dinb(n7344), .dout(n7350));
  jand g07287(.dina(n343), .dinb(n149), .dout(n7351));
  jand g07288(.dina(n7351), .dinb(n3882), .dout(n7352));
  jand g07289(.dina(n3237), .dinb(n2499), .dout(n7353));
  jand g07290(.dina(n1281), .dinb(n93), .dout(n7354));
  jand g07291(.dina(n7354), .dinb(n7353), .dout(n7355));
  jand g07292(.dina(n7355), .dinb(n7352), .dout(n7356));
  jand g07293(.dina(n7356), .dinb(n7350), .dout(n7357));
  jand g07294(.dina(n7357), .dinb(n7341), .dout(n7358));
  jand g07295(.dina(n7358), .dinb(n2882), .dout(n7359));
  jand g07296(.dina(n5038), .dinb(n3949), .dout(n7360));
  jand g07297(.dina(n7360), .dinb(n7359), .dout(n7361));
  jnot g07298(.din(n7361), .dout(n7362));
  jnot g07299(.din(n2897), .dout(n7363));
  jor  g07300(.dina(n7363), .dinb(n797), .dout(n7364));
  jnot g07301(.din(n3609), .dout(n7365));
  jor  g07302(.dina(n7365), .dinb(n7364), .dout(n7366));
  jor  g07303(.dina(n7210), .dinb(n7314), .dout(n7367));
  jor  g07304(.dina(n7367), .dinb(n2274), .dout(n7368));
  jor  g07305(.dina(n7368), .dinb(n3615), .dout(n7369));
  jor  g07306(.dina(n7369), .dinb(n7366), .dout(n7370));
  jnot g07307(.din(n3128), .dout(n7371));
  jnot g07308(.din(n3129), .dout(n7372));
  jor  g07309(.dina(n2792), .dinb(n2088), .dout(n7373));
  jor  g07310(.dina(n7373), .dinb(n7372), .dout(n7374));
  jor  g07311(.dina(n7374), .dinb(n7371), .dout(n7375));
  jnot g07312(.din(n1974), .dout(n7376));
  jnot g07313(.din(n1349), .dout(n7377));
  jnot g07314(.din(n612), .dout(n7378));
  jor  g07315(.dina(n3210), .dinb(n283), .dout(n7379));
  jor  g07316(.dina(n7379), .dinb(n7378), .dout(n7380));
  jor  g07317(.dina(n7380), .dinb(n7377), .dout(n7381));
  jor  g07318(.dina(n7381), .dinb(n7376), .dout(n7382));
  jor  g07319(.dina(n7382), .dinb(n7375), .dout(n7383));
  jor  g07320(.dina(n7383), .dinb(n7370), .dout(n7384));
  jnot g07321(.din(n3629), .dout(n7385));
  jnot g07322(.din(n2660), .dout(n7386));
  jor  g07323(.dina(n3631), .dinb(n7386), .dout(n7387));
  jor  g07324(.dina(n7387), .dinb(n7385), .dout(n7388));
  jor  g07325(.dina(n3173), .dinb(n3203), .dout(n7389));
  jor  g07326(.dina(n3640), .dinb(n7389), .dout(n7390));
  jor  g07327(.dina(n7390), .dinb(n7388), .dout(n7391));
  jnot g07328(.din(n3644), .dout(n7392));
  jor  g07329(.dina(n7392), .dinb(n2467), .dout(n7393));
  jor  g07330(.dina(n3647), .dinb(n7393), .dout(n7394));
  jor  g07331(.dina(n3655), .dinb(n3319), .dout(n7395));
  jor  g07332(.dina(n7395), .dinb(n3653), .dout(n7396));
  jor  g07333(.dina(n7396), .dinb(n7394), .dout(n7397));
  jor  g07334(.dina(n2075), .dinb(n1279), .dout(n7398));
  jor  g07335(.dina(n3661), .dinb(n2071), .dout(n7399));
  jor  g07336(.dina(n7399), .dinb(n7398), .dout(n7400));
  jor  g07337(.dina(n3671), .dinb(n7400), .dout(n7401));
  jor  g07338(.dina(n7401), .dinb(n7397), .dout(n7402));
  jor  g07339(.dina(n7402), .dinb(n7391), .dout(n7403));
  jor  g07340(.dina(n7403), .dinb(n7384), .dout(n7404));
  jor  g07341(.dina(n7404), .dinb(n7274), .dout(n7405));
  jand g07342(.dina(n7405), .dinb(n3605), .dout(n7406));
  jxor g07343(.dina(n7406), .dinb(n7326), .dout(n7407));
  jand g07344(.dina(n7407), .dinb(n732), .dout(n7408));
  jand g07345(.dina(n3855), .dinb(n7326), .dout(n7409));
  jand g07346(.dina(n3858), .dinb(n7405), .dout(n7410));
  jnot g07347(.din(n3605), .dout(n7411));
  jand g07348(.dina(n3851), .dinb(n7411), .dout(n7412));
  jor  g07349(.dina(n7412), .dinb(n7410), .dout(n7413));
  jor  g07350(.dina(n7413), .dinb(n7409), .dout(n7414));
  jor  g07351(.dina(n7414), .dinb(n7408), .dout(n7415));
  jand g07352(.dina(n7415), .dinb(n7362), .dout(n7416));
  jnot g07353(.din(n7416), .dout(n7417));
  jand g07354(.dina(n5992), .dinb(n4692), .dout(n7418));
  jand g07355(.dina(n7418), .dinb(n2100), .dout(n7419));
  jand g07356(.dina(n805), .dinb(n365), .dout(n7420));
  jand g07357(.dina(n1221), .dinb(n434), .dout(n7421));
  jand g07358(.dina(n7421), .dinb(n262), .dout(n7422));
  jand g07359(.dina(n7422), .dinb(n7420), .dout(n7423));
  jand g07360(.dina(n7423), .dinb(n2436), .dout(n7424));
  jand g07361(.dina(n1785), .dinb(n346), .dout(n7425));
  jand g07362(.dina(n7425), .dinb(n655), .dout(n7426));
  jand g07363(.dina(n739), .dinb(n184), .dout(n7427));
  jand g07364(.dina(n7427), .dinb(n988), .dout(n7428));
  jand g07365(.dina(n2915), .dinb(n820), .dout(n7429));
  jand g07366(.dina(n7429), .dinb(n7428), .dout(n7430));
  jand g07367(.dina(n7430), .dinb(n7426), .dout(n7431));
  jand g07368(.dina(n7431), .dinb(n7424), .dout(n7432));
  jand g07369(.dina(n7432), .dinb(n7419), .dout(n7433));
  jand g07370(.dina(n7433), .dinb(n3487), .dout(n7434));
  jand g07371(.dina(n3462), .dinb(n178), .dout(n7435));
  jand g07372(.dina(n7435), .dinb(n4287), .dout(n7436));
  jand g07373(.dina(n826), .dinb(n443), .dout(n7437));
  jand g07374(.dina(n756), .dinb(n149), .dout(n7438));
  jand g07375(.dina(n7438), .dinb(n7437), .dout(n7439));
  jand g07376(.dina(n7439), .dinb(n2427), .dout(n7440));
  jand g07377(.dina(n7440), .dinb(n7436), .dout(n7441));
  jand g07378(.dina(n1268), .dinb(n367), .dout(n7442));
  jand g07379(.dina(n7442), .dinb(n1644), .dout(n7443));
  jand g07380(.dina(n5898), .dinb(n2619), .dout(n7444));
  jand g07381(.dina(n7444), .dinb(n7443), .dout(n7445));
  jand g07382(.dina(n708), .dinb(n508), .dout(n7446));
  jand g07383(.dina(n7446), .dinb(n994), .dout(n7447));
  jand g07384(.dina(n483), .dinb(n418), .dout(n7448));
  jand g07385(.dina(n711), .dinb(n439), .dout(n7449));
  jand g07386(.dina(n7449), .dinb(n7448), .dout(n7450));
  jand g07387(.dina(n7450), .dinb(n7447), .dout(n7451));
  jand g07388(.dina(n7451), .dinb(n7445), .dout(n7452));
  jand g07389(.dina(n2875), .dinb(n622), .dout(n7453));
  jand g07390(.dina(n594), .dinb(n384), .dout(n7454));
  jand g07391(.dina(n2382), .dinb(n277), .dout(n7455));
  jand g07392(.dina(n7455), .dinb(n7454), .dout(n7456));
  jand g07393(.dina(n7456), .dinb(n7453), .dout(n7457));
  jand g07394(.dina(n7457), .dinb(n7452), .dout(n7458));
  jand g07395(.dina(n7458), .dinb(n7441), .dout(n7459));
  jand g07396(.dina(n7459), .dinb(n2269), .dout(n7460));
  jand g07397(.dina(n7460), .dinb(n7434), .dout(n7461));
  jor  g07398(.dina(n7461), .dinb(n7417), .dout(n7462));
  jxor g07399(.dina(n7461), .dinb(n7417), .dout(n7463));
  jnot g07400(.din(n7463), .dout(n7464));
  jnot g07401(.din(n3518), .dout(n7465));
  jxor g07402(.dina(n3678), .dinb(n7465), .dout(n7466));
  jor  g07403(.dina(n7466), .dinb(n6463), .dout(n7467));
  jand g07404(.dina(n3858), .dinb(n7326), .dout(n7468));
  jand g07405(.dina(n3855), .dinb(n3411), .dout(n7469));
  jand g07406(.dina(n3851), .dinb(n7405), .dout(n7470));
  jor  g07407(.dina(n7470), .dinb(n7469), .dout(n7471));
  jor  g07408(.dina(n7471), .dinb(n7468), .dout(n7472));
  jnot g07409(.din(n7472), .dout(n7473));
  jand g07410(.dina(n7473), .dinb(n7467), .dout(n7474));
  jor  g07411(.dina(n7474), .dinb(n7464), .dout(n7475));
  jand g07412(.dina(n7475), .dinb(n7462), .dout(n7476));
  jnot g07413(.din(n7476), .dout(n7477));
  jxor g07414(.dina(n7333), .dinb(n7175), .dout(n7478));
  jand g07415(.dina(n7478), .dinb(n7477), .dout(n7479));
  jnot g07416(.din(n7479), .dout(n7480));
  jand g07417(.dina(n7480), .dinb(n7334), .dout(n7481));
  jnot g07418(.din(n7481), .dout(n7482));
  jxor g07419(.dina(n7139), .dinb(n7129), .dout(n7483));
  jand g07420(.dina(n7483), .dinb(n7482), .dout(n7484));
  jnot g07421(.din(n7484), .dout(n7485));
  jand g07422(.dina(n7485), .dinb(n7140), .dout(n7486));
  jnot g07423(.din(n7486), .dout(n7487));
  jxor g07424(.dina(n7084), .dinb(n7075), .dout(n7488));
  jand g07425(.dina(n7488), .dinb(n7487), .dout(n7489));
  jnot g07426(.din(n7489), .dout(n7490));
  jand g07427(.dina(n7490), .dinb(n7085), .dout(n7491));
  jnot g07428(.din(n7491), .dout(n7492));
  jxor g07429(.dina(n7039), .dinb(n7030), .dout(n7493));
  jand g07430(.dina(n7493), .dinb(n7492), .dout(n7494));
  jnot g07431(.din(n7494), .dout(n7495));
  jand g07432(.dina(n7495), .dinb(n7040), .dout(n7496));
  jnot g07433(.din(n7496), .dout(n7497));
  jxor g07434(.dina(n6689), .dinb(n6680), .dout(n7498));
  jand g07435(.dina(n7498), .dinb(n7497), .dout(n7499));
  jnot g07436(.din(n7499), .dout(n7500));
  jxor g07437(.dina(n7498), .dinb(n7497), .dout(n7501));
  jnot g07438(.din(n7501), .dout(n7502));
  jand g07439(.dina(n6706), .dinb(n4449), .dout(n7503));
  jand g07440(.dina(n4453), .dinb(n2808), .dout(n7504));
  jand g07441(.dina(n4461), .dinb(n2954), .dout(n7505));
  jand g07442(.dina(n4457), .dinb(n2867), .dout(n7506));
  jor  g07443(.dina(n7506), .dinb(n7505), .dout(n7507));
  jor  g07444(.dina(n7507), .dinb(n7504), .dout(n7508));
  jor  g07445(.dina(n7508), .dinb(n7503), .dout(n7509));
  jxor g07446(.dina(n7509), .dinb(n88), .dout(n7510));
  jor  g07447(.dina(n7510), .dinb(n7502), .dout(n7511));
  jand g07448(.dina(n7511), .dinb(n7500), .dout(n7512));
  jnot g07449(.din(n7512), .dout(n7513));
  jxor g07450(.dina(n6996), .dinb(n6987), .dout(n7514));
  jand g07451(.dina(n7514), .dinb(n7513), .dout(n7515));
  jnot g07452(.din(n7515), .dout(n7516));
  jand g07453(.dina(n7516), .dinb(n6997), .dout(n7517));
  jnot g07454(.din(n7517), .dout(n7518));
  jxor g07455(.dina(n6984), .dinb(n6975), .dout(n7519));
  jand g07456(.dina(n7519), .dinb(n7518), .dout(n7520));
  jnot g07457(.din(n7520), .dout(n7521));
  jand g07458(.dina(n7521), .dinb(n6985), .dout(n7522));
  jnot g07459(.din(n7522), .dout(n7523));
  jxor g07460(.dina(n6713), .dinb(n6705), .dout(n7524));
  jand g07461(.dina(n7524), .dinb(n7523), .dout(n7525));
  jnot g07462(.din(n7525), .dout(n7526));
  jxor g07463(.dina(n7524), .dinb(n7523), .dout(n7527));
  jnot g07464(.din(n7527), .dout(n7528));
  jor  g07465(.dina(n6464), .dinb(n4724), .dout(n7529));
  jor  g07466(.dina(n4905), .dinb(n2601), .dout(n7530));
  jor  g07467(.dina(n4735), .dinb(n2694), .dout(n7531));
  jor  g07468(.dina(n4733), .dinb(n2731), .dout(n7532));
  jand g07469(.dina(n7532), .dinb(n7531), .dout(n7533));
  jand g07470(.dina(n7533), .dinb(n7530), .dout(n7534));
  jand g07471(.dina(n7534), .dinb(n7529), .dout(n7535));
  jxor g07472(.dina(n7535), .dinb(\a[29] ), .dout(n7536));
  jor  g07473(.dina(n7536), .dinb(n7528), .dout(n7537));
  jand g07474(.dina(n7537), .dinb(n7526), .dout(n7538));
  jnot g07475(.din(n7538), .dout(n7539));
  jxor g07476(.dina(n6728), .dinb(n6720), .dout(n7540));
  jand g07477(.dina(n7540), .dinb(n7539), .dout(n7541));
  jnot g07478(.din(n7541), .dout(n7542));
  jxor g07479(.dina(n7540), .dinb(n7539), .dout(n7543));
  jnot g07480(.din(n7543), .dout(n7544));
  jand g07481(.dina(n5844), .dinb(n75), .dout(n7545));
  jand g07482(.dina(n4745), .dinb(n2411), .dout(n7546));
  jand g07483(.dina(n4933), .dinb(n2237), .dout(n7547));
  jand g07484(.dina(n4918), .dinb(n2343), .dout(n7548));
  jor  g07485(.dina(n7548), .dinb(n7547), .dout(n7549));
  jor  g07486(.dina(n7549), .dinb(n7546), .dout(n7550));
  jor  g07487(.dina(n7550), .dinb(n7545), .dout(n7551));
  jxor g07488(.dina(n7551), .dinb(n68), .dout(n7552));
  jor  g07489(.dina(n7552), .dinb(n7544), .dout(n7553));
  jand g07490(.dina(n7553), .dinb(n7542), .dout(n7554));
  jnot g07491(.din(n7554), .dout(n7555));
  jxor g07492(.dina(n6867), .dinb(n6859), .dout(n7556));
  jand g07493(.dina(n7556), .dinb(n7555), .dout(n7557));
  jnot g07494(.din(n7557), .dout(n7558));
  jxor g07495(.dina(n7556), .dinb(n7555), .dout(n7559));
  jnot g07496(.din(n7559), .dout(n7560));
  jand g07497(.dina(n5440), .dinb(n5365), .dout(n7561));
  jand g07498(.dina(n5424), .dinb(n1956), .dout(n7562));
  jand g07499(.dina(n5500), .dinb(n1862), .dout(n7563));
  jand g07500(.dina(n5363), .dinb(n2067), .dout(n7564));
  jor  g07501(.dina(n7564), .dinb(n7563), .dout(n7565));
  jor  g07502(.dina(n7565), .dinb(n7562), .dout(n7566));
  jor  g07503(.dina(n7566), .dinb(n7561), .dout(n7567));
  jxor g07504(.dina(n7567), .dinb(n72), .dout(n7568));
  jor  g07505(.dina(n7568), .dinb(n7560), .dout(n7569));
  jand g07506(.dina(n7569), .dinb(n7558), .dout(n7570));
  jnot g07507(.din(n7570), .dout(n7571));
  jxor g07508(.dina(n6972), .dinb(n6971), .dout(n7572));
  jand g07509(.dina(n7572), .dinb(n7571), .dout(n7573));
  jor  g07510(.dina(n7573), .dinb(n6973), .dout(n7574));
  jxor g07511(.dina(n6888), .dinb(n6880), .dout(n7575));
  jand g07512(.dina(n7575), .dinb(n7574), .dout(n7576));
  jnot g07513(.din(n7576), .dout(n7577));
  jxor g07514(.dina(n7575), .dinb(n7574), .dout(n7578));
  jnot g07515(.din(n7578), .dout(n7579));
  jand g07516(.dina(n5693), .dinb(n4258), .dout(n7580));
  jand g07517(.dina(n6209), .dinb(n1343), .dout(n7581));
  jand g07518(.dina(n6131), .dinb(n1445), .dout(n7582));
  jand g07519(.dina(n5691), .dinb(n1560), .dout(n7583));
  jor  g07520(.dina(n7583), .dinb(n7582), .dout(n7584));
  jor  g07521(.dina(n7584), .dinb(n7581), .dout(n7585));
  jor  g07522(.dina(n7585), .dinb(n7580), .dout(n7586));
  jxor g07523(.dina(n7586), .dinb(n4247), .dout(n7587));
  jor  g07524(.dina(n7587), .dinb(n7579), .dout(n7588));
  jand g07525(.dina(n7588), .dinb(n7577), .dout(n7589));
  jnot g07526(.din(n7589), .dout(n7590));
  jxor g07527(.dina(n6904), .dinb(n6896), .dout(n7591));
  jand g07528(.dina(n7591), .dinb(n7590), .dout(n7592));
  jnot g07529(.din(n7592), .dout(n7593));
  jxor g07530(.dina(n7591), .dinb(n7590), .dout(n7594));
  jnot g07531(.din(n7594), .dout(n7595));
  jand g07532(.dina(n6340), .dinb(n3848), .dout(n7596));
  jand g07533(.dina(n6556), .dinb(n922), .dout(n7597));
  jand g07534(.dina(n6798), .dinb(n3853), .dout(n7598));
  jand g07535(.dina(n6338), .dinb(n1076), .dout(n7599));
  jor  g07536(.dina(n7599), .dinb(n7598), .dout(n7600));
  jor  g07537(.dina(n7600), .dinb(n7597), .dout(n7601));
  jor  g07538(.dina(n7601), .dinb(n7596), .dout(n7602));
  jxor g07539(.dina(n7602), .dinb(n5064), .dout(n7603));
  jor  g07540(.dina(n7603), .dinb(n7595), .dout(n7604));
  jand g07541(.dina(n7604), .dinb(n7593), .dout(n7605));
  jnot g07542(.din(n7605), .dout(n7606));
  jxor g07543(.dina(n6961), .dinb(n6960), .dout(n7607));
  jand g07544(.dina(n7607), .dinb(n7606), .dout(n7608));
  jor  g07545(.dina(n7608), .dinb(n6962), .dout(n7609));
  jnot g07546(.din(n7609), .dout(n7610));
  jor  g07547(.dina(n6937), .dinb(n4731), .dout(n7611));
  jor  g07548(.dina(n6935), .dinb(n4597), .dout(n7612));
  jand g07549(.dina(n6930), .dinb(n6929), .dout(n7613));
  jnot g07550(.din(n7613), .dout(n7614));
  jor  g07551(.dina(n7614), .dinb(n4630), .dout(n7615));
  jand g07552(.dina(n7615), .dinb(n7612), .dout(n7616));
  jand g07553(.dina(n7616), .dinb(n7611), .dout(n7617));
  jxor g07554(.dina(n7617), .dinb(\a[14] ), .dout(n7618));
  jor  g07555(.dina(n7618), .dinb(n7610), .dout(n7619));
  jxor g07556(.dina(n7618), .dinb(n7610), .dout(n7620));
  jxor g07557(.dina(n6925), .dinb(n6917), .dout(n7621));
  jand g07558(.dina(n7621), .dinb(n7620), .dout(n7622));
  jnot g07559(.din(n7622), .dout(n7623));
  jand g07560(.dina(n7623), .dinb(n7619), .dout(n7624));
  jnot g07561(.din(n7624), .dout(n7625));
  jxor g07562(.dina(n6944), .dinb(n6943), .dout(n7626));
  jand g07563(.dina(n7626), .dinb(n7625), .dout(n7627));
  jxor g07564(.dina(n7626), .dinb(n7625), .dout(n7628));
  jxor g07565(.dina(n7572), .dinb(n7571), .dout(n7629));
  jnot g07566(.din(n7629), .dout(n7630));
  jand g07567(.dina(n5693), .dinb(n4866), .dout(n7631));
  jand g07568(.dina(n6131), .dinb(n1560), .dout(n7632));
  jand g07569(.dina(n5691), .dinb(n1624), .dout(n7633));
  jand g07570(.dina(n6209), .dinb(n1445), .dout(n7634));
  jor  g07571(.dina(n7634), .dinb(n7633), .dout(n7635));
  jor  g07572(.dina(n7635), .dinb(n7632), .dout(n7636));
  jor  g07573(.dina(n7636), .dinb(n7631), .dout(n7637));
  jxor g07574(.dina(n7637), .dinb(n4247), .dout(n7638));
  jor  g07575(.dina(n7638), .dinb(n7630), .dout(n7639));
  jand g07576(.dina(n5861), .dinb(n75), .dout(n7640));
  jand g07577(.dina(n4918), .dinb(n2411), .dout(n7641));
  jand g07578(.dina(n4933), .dinb(n2343), .dout(n7642));
  jand g07579(.dina(n4745), .dinb(n2497), .dout(n7643));
  jor  g07580(.dina(n7643), .dinb(n7642), .dout(n7644));
  jor  g07581(.dina(n7644), .dinb(n7641), .dout(n7645));
  jor  g07582(.dina(n7645), .dinb(n7640), .dout(n7646));
  jxor g07583(.dina(n7646), .dinb(n68), .dout(n7647));
  jnot g07584(.din(n7647), .dout(n7648));
  jxor g07585(.dina(n7536), .dinb(n7528), .dout(n7649));
  jand g07586(.dina(n7649), .dinb(n7648), .dout(n7650));
  jand g07587(.dina(n6591), .dinb(n4449), .dout(n7651));
  jand g07588(.dina(n4453), .dinb(n2695), .dout(n7652));
  jand g07589(.dina(n4461), .dinb(n2808), .dout(n7653));
  jand g07590(.dina(n4457), .dinb(n2732), .dout(n7654));
  jor  g07591(.dina(n7654), .dinb(n7653), .dout(n7655));
  jor  g07592(.dina(n7655), .dinb(n7652), .dout(n7656));
  jor  g07593(.dina(n7656), .dinb(n7651), .dout(n7657));
  jxor g07594(.dina(n7657), .dinb(n88), .dout(n7658));
  jnot g07595(.din(n7658), .dout(n7659));
  jxor g07596(.dina(n7519), .dinb(n7518), .dout(n7660));
  jand g07597(.dina(n7660), .dinb(n7659), .dout(n7661));
  jnot g07598(.din(n7661), .dout(n7662));
  jxor g07599(.dina(n7660), .dinb(n7659), .dout(n7663));
  jnot g07600(.din(n7663), .dout(n7664));
  jand g07601(.dina(n6247), .dinb(n75), .dout(n7665));
  jand g07602(.dina(n4933), .dinb(n2411), .dout(n7666));
  jand g07603(.dina(n4745), .dinb(n2602), .dout(n7667));
  jand g07604(.dina(n4918), .dinb(n2497), .dout(n7668));
  jor  g07605(.dina(n7668), .dinb(n7667), .dout(n7669));
  jor  g07606(.dina(n7669), .dinb(n7666), .dout(n7670));
  jor  g07607(.dina(n7670), .dinb(n7665), .dout(n7671));
  jxor g07608(.dina(n7671), .dinb(n68), .dout(n7672));
  jor  g07609(.dina(n7672), .dinb(n7664), .dout(n7673));
  jand g07610(.dina(n7673), .dinb(n7662), .dout(n7674));
  jnot g07611(.din(n7674), .dout(n7675));
  jxor g07612(.dina(n7649), .dinb(n7648), .dout(n7676));
  jand g07613(.dina(n7676), .dinb(n7675), .dout(n7677));
  jor  g07614(.dina(n7677), .dinb(n7650), .dout(n7678));
  jxor g07615(.dina(n7552), .dinb(n7544), .dout(n7679));
  jand g07616(.dina(n7679), .dinb(n7678), .dout(n7680));
  jnot g07617(.din(n7680), .dout(n7681));
  jxor g07618(.dina(n7679), .dinb(n7678), .dout(n7682));
  jnot g07619(.din(n7682), .dout(n7683));
  jand g07620(.dina(n5365), .dinb(n5303), .dout(n7684));
  jand g07621(.dina(n5424), .dinb(n2067), .dout(n7685));
  jand g07622(.dina(n5500), .dinb(n1956), .dout(n7686));
  jand g07623(.dina(n5363), .dinb(n2128), .dout(n7687));
  jor  g07624(.dina(n7687), .dinb(n7686), .dout(n7688));
  jor  g07625(.dina(n7688), .dinb(n7685), .dout(n7689));
  jor  g07626(.dina(n7689), .dinb(n7684), .dout(n7690));
  jxor g07627(.dina(n7690), .dinb(n72), .dout(n7691));
  jor  g07628(.dina(n7691), .dinb(n7683), .dout(n7692));
  jand g07629(.dina(n7692), .dinb(n7681), .dout(n7693));
  jnot g07630(.din(n7693), .dout(n7694));
  jxor g07631(.dina(n7568), .dinb(n7560), .dout(n7695));
  jand g07632(.dina(n7695), .dinb(n7694), .dout(n7696));
  jnot g07633(.din(n7696), .dout(n7697));
  jxor g07634(.dina(n7695), .dinb(n7694), .dout(n7698));
  jnot g07635(.din(n7698), .dout(n7699));
  jand g07636(.dina(n5693), .dinb(n4849), .dout(n7700));
  jand g07637(.dina(n6209), .dinb(n1560), .dout(n7701));
  jand g07638(.dina(n6131), .dinb(n1624), .dout(n7702));
  jand g07639(.dina(n5691), .dinb(n1776), .dout(n7703));
  jor  g07640(.dina(n7703), .dinb(n7702), .dout(n7704));
  jor  g07641(.dina(n7704), .dinb(n7701), .dout(n7705));
  jor  g07642(.dina(n7705), .dinb(n7700), .dout(n7706));
  jxor g07643(.dina(n7706), .dinb(n4247), .dout(n7707));
  jor  g07644(.dina(n7707), .dinb(n7699), .dout(n7708));
  jand g07645(.dina(n7708), .dinb(n7697), .dout(n7709));
  jnot g07646(.din(n7709), .dout(n7710));
  jxor g07647(.dina(n7638), .dinb(n7630), .dout(n7711));
  jand g07648(.dina(n7711), .dinb(n7710), .dout(n7712));
  jnot g07649(.din(n7712), .dout(n7713));
  jand g07650(.dina(n7713), .dinb(n7639), .dout(n7714));
  jnot g07651(.din(n7714), .dout(n7715));
  jxor g07652(.dina(n7587), .dinb(n7579), .dout(n7716));
  jand g07653(.dina(n7716), .dinb(n7715), .dout(n7717));
  jnot g07654(.din(n7717), .dout(n7718));
  jxor g07655(.dina(n7716), .dinb(n7715), .dout(n7719));
  jnot g07656(.din(n7719), .dout(n7720));
  jand g07657(.dina(n6340), .dinb(n4026), .dout(n7721));
  jand g07658(.dina(n6556), .dinb(n1076), .dout(n7722));
  jand g07659(.dina(n6798), .dinb(n922), .dout(n7723));
  jand g07660(.dina(n6338), .dinb(n1213), .dout(n7724));
  jor  g07661(.dina(n7724), .dinb(n7723), .dout(n7725));
  jor  g07662(.dina(n7725), .dinb(n7722), .dout(n7726));
  jor  g07663(.dina(n7726), .dinb(n7721), .dout(n7727));
  jxor g07664(.dina(n7727), .dinb(n5064), .dout(n7728));
  jor  g07665(.dina(n7728), .dinb(n7720), .dout(n7729));
  jand g07666(.dina(n7729), .dinb(n7718), .dout(n7730));
  jnot g07667(.din(n7730), .dout(n7731));
  jxor g07668(.dina(n7603), .dinb(n7595), .dout(n7732));
  jand g07669(.dina(n7732), .dinb(n7731), .dout(n7733));
  jnot g07670(.din(n7733), .dout(n7734));
  jxor g07671(.dina(n7732), .dinb(n7731), .dout(n7735));
  jnot g07672(.din(n7735), .dout(n7736));
  jand g07673(.dina(n6936), .dinb(n4752), .dout(n7737));
  jand g07674(.dina(n7613), .dinb(n4451), .dout(n7738));
  jand g07675(.dina(n6934), .dinb(n4358), .dout(n7739));
  jor  g07676(.dina(n6933), .dinb(n6929), .dout(n7740));
  jnot g07677(.din(n7740), .dout(n7741));
  jand g07678(.dina(n7741), .dinb(n4598), .dout(n7742));
  jor  g07679(.dina(n7742), .dinb(n7739), .dout(n7743));
  jor  g07680(.dina(n7743), .dinb(n7738), .dout(n7744));
  jor  g07681(.dina(n7744), .dinb(n7737), .dout(n7745));
  jxor g07682(.dina(n7745), .dinb(n5292), .dout(n7746));
  jor  g07683(.dina(n7746), .dinb(n7736), .dout(n7747));
  jand g07684(.dina(n7747), .dinb(n7734), .dout(n7748));
  jand g07685(.dina(n6936), .dinb(n4636), .dout(n7749));
  jand g07686(.dina(n6934), .dinb(n4451), .dout(n7750));
  jand g07687(.dina(n7613), .dinb(n4598), .dout(n7751));
  jand g07688(.dina(n7741), .dinb(n4631), .dout(n7752));
  jor  g07689(.dina(n7752), .dinb(n7751), .dout(n7753));
  jor  g07690(.dina(n7753), .dinb(n7750), .dout(n7754));
  jor  g07691(.dina(n7754), .dinb(n7749), .dout(n7755));
  jxor g07692(.dina(n7755), .dinb(n5292), .dout(n7756));
  jor  g07693(.dina(n7756), .dinb(n7748), .dout(n7757));
  jxor g07694(.dina(n7607), .dinb(n7606), .dout(n7758));
  jxor g07695(.dina(n7756), .dinb(n7748), .dout(n7759));
  jand g07696(.dina(n7759), .dinb(n7758), .dout(n7760));
  jnot g07697(.din(n7760), .dout(n7761));
  jand g07698(.dina(n7761), .dinb(n7757), .dout(n7762));
  jnot g07699(.din(n7762), .dout(n7763));
  jxor g07700(.dina(n7621), .dinb(n7620), .dout(n7764));
  jand g07701(.dina(n7764), .dinb(n7763), .dout(n7765));
  jand g07702(.dina(n6340), .dinb(n4043), .dout(n7766));
  jand g07703(.dina(n6798), .dinb(n1076), .dout(n7767));
  jand g07704(.dina(n6556), .dinb(n1213), .dout(n7768));
  jand g07705(.dina(n6338), .dinb(n1343), .dout(n7769));
  jor  g07706(.dina(n7769), .dinb(n7768), .dout(n7770));
  jor  g07707(.dina(n7770), .dinb(n7767), .dout(n7771));
  jor  g07708(.dina(n7771), .dinb(n7766), .dout(n7772));
  jxor g07709(.dina(n7772), .dinb(n5064), .dout(n7773));
  jnot g07710(.din(n7773), .dout(n7774));
  jxor g07711(.dina(n7711), .dinb(n7710), .dout(n7775));
  jand g07712(.dina(n7775), .dinb(n7774), .dout(n7776));
  jand g07713(.dina(n5624), .dinb(n5365), .dout(n7777));
  jand g07714(.dina(n5363), .dinb(n2237), .dout(n7778));
  jand g07715(.dina(n5424), .dinb(n2128), .dout(n7779));
  jand g07716(.dina(n5500), .dinb(n2067), .dout(n7780));
  jor  g07717(.dina(n7780), .dinb(n7779), .dout(n7781));
  jor  g07718(.dina(n7781), .dinb(n7778), .dout(n7782));
  jor  g07719(.dina(n7782), .dinb(n7777), .dout(n7783));
  jxor g07720(.dina(n7783), .dinb(n72), .dout(n7784));
  jnot g07721(.din(n7784), .dout(n7785));
  jxor g07722(.dina(n7676), .dinb(n7675), .dout(n7786));
  jand g07723(.dina(n7786), .dinb(n7785), .dout(n7787));
  jand g07724(.dina(n6439), .dinb(n4449), .dout(n7788));
  jand g07725(.dina(n4457), .dinb(n2808), .dout(n7789));
  jand g07726(.dina(n4453), .dinb(n2732), .dout(n7790));
  jand g07727(.dina(n4461), .dinb(n2867), .dout(n7791));
  jor  g07728(.dina(n7791), .dinb(n7790), .dout(n7792));
  jor  g07729(.dina(n7792), .dinb(n7789), .dout(n7793));
  jor  g07730(.dina(n7793), .dinb(n7788), .dout(n7794));
  jxor g07731(.dina(n7794), .dinb(n88), .dout(n7795));
  jnot g07732(.din(n7795), .dout(n7796));
  jxor g07733(.dina(n7514), .dinb(n7513), .dout(n7797));
  jand g07734(.dina(n7797), .dinb(n7796), .dout(n7798));
  jnot g07735(.din(n7798), .dout(n7799));
  jxor g07736(.dina(n7797), .dinb(n7796), .dout(n7800));
  jnot g07737(.din(n7800), .dout(n7801));
  jand g07738(.dina(n6050), .dinb(n75), .dout(n7802));
  jand g07739(.dina(n4745), .dinb(n2695), .dout(n7803));
  jand g07740(.dina(n4918), .dinb(n2602), .dout(n7804));
  jand g07741(.dina(n4933), .dinb(n2497), .dout(n7805));
  jor  g07742(.dina(n7805), .dinb(n7804), .dout(n7806));
  jor  g07743(.dina(n7806), .dinb(n7803), .dout(n7807));
  jor  g07744(.dina(n7807), .dinb(n7802), .dout(n7808));
  jxor g07745(.dina(n7808), .dinb(n68), .dout(n7809));
  jor  g07746(.dina(n7809), .dinb(n7801), .dout(n7810));
  jand g07747(.dina(n7810), .dinb(n7799), .dout(n7811));
  jnot g07748(.din(n7811), .dout(n7812));
  jxor g07749(.dina(n7672), .dinb(n7664), .dout(n7813));
  jand g07750(.dina(n7813), .dinb(n7812), .dout(n7814));
  jnot g07751(.din(n7814), .dout(n7815));
  jxor g07752(.dina(n7813), .dinb(n7812), .dout(n7816));
  jnot g07753(.din(n7816), .dout(n7817));
  jand g07754(.dina(n5607), .dinb(n5365), .dout(n7818));
  jand g07755(.dina(n5424), .dinb(n2237), .dout(n7819));
  jand g07756(.dina(n5363), .dinb(n2343), .dout(n7820));
  jand g07757(.dina(n5500), .dinb(n2128), .dout(n7821));
  jor  g07758(.dina(n7821), .dinb(n7820), .dout(n7822));
  jor  g07759(.dina(n7822), .dinb(n7819), .dout(n7823));
  jor  g07760(.dina(n7823), .dinb(n7818), .dout(n7824));
  jxor g07761(.dina(n7824), .dinb(n72), .dout(n7825));
  jor  g07762(.dina(n7825), .dinb(n7817), .dout(n7826));
  jand g07763(.dina(n7826), .dinb(n7815), .dout(n7827));
  jnot g07764(.din(n7827), .dout(n7828));
  jxor g07765(.dina(n7786), .dinb(n7785), .dout(n7829));
  jand g07766(.dina(n7829), .dinb(n7828), .dout(n7830));
  jor  g07767(.dina(n7830), .dinb(n7787), .dout(n7831));
  jxor g07768(.dina(n7691), .dinb(n7683), .dout(n7832));
  jand g07769(.dina(n7832), .dinb(n7831), .dout(n7833));
  jnot g07770(.din(n7833), .dout(n7834));
  jxor g07771(.dina(n7832), .dinb(n7831), .dout(n7835));
  jnot g07772(.din(n7835), .dout(n7836));
  jand g07773(.dina(n5693), .dinb(n5075), .dout(n7837));
  jand g07774(.dina(n6209), .dinb(n1624), .dout(n7838));
  jand g07775(.dina(n6131), .dinb(n1776), .dout(n7839));
  jand g07776(.dina(n5691), .dinb(n1862), .dout(n7840));
  jor  g07777(.dina(n7840), .dinb(n7839), .dout(n7841));
  jor  g07778(.dina(n7841), .dinb(n7838), .dout(n7842));
  jor  g07779(.dina(n7842), .dinb(n7837), .dout(n7843));
  jxor g07780(.dina(n7843), .dinb(n4247), .dout(n7844));
  jor  g07781(.dina(n7844), .dinb(n7836), .dout(n7845));
  jand g07782(.dina(n7845), .dinb(n7834), .dout(n7846));
  jnot g07783(.din(n7846), .dout(n7847));
  jxor g07784(.dina(n7707), .dinb(n7699), .dout(n7848));
  jand g07785(.dina(n7848), .dinb(n7847), .dout(n7849));
  jnot g07786(.din(n7849), .dout(n7850));
  jxor g07787(.dina(n7848), .dinb(n7847), .dout(n7851));
  jnot g07788(.din(n7851), .dout(n7852));
  jand g07789(.dina(n6340), .dinb(n4772), .dout(n7853));
  jand g07790(.dina(n6798), .dinb(n1213), .dout(n7854));
  jand g07791(.dina(n6556), .dinb(n1343), .dout(n7855));
  jand g07792(.dina(n6338), .dinb(n1445), .dout(n7856));
  jor  g07793(.dina(n7856), .dinb(n7855), .dout(n7857));
  jor  g07794(.dina(n7857), .dinb(n7854), .dout(n7858));
  jor  g07795(.dina(n7858), .dinb(n7853), .dout(n7859));
  jxor g07796(.dina(n7859), .dinb(n5064), .dout(n7860));
  jor  g07797(.dina(n7860), .dinb(n7852), .dout(n7861));
  jand g07798(.dina(n7861), .dinb(n7850), .dout(n7862));
  jnot g07799(.din(n7862), .dout(n7863));
  jxor g07800(.dina(n7775), .dinb(n7774), .dout(n7864));
  jand g07801(.dina(n7864), .dinb(n7863), .dout(n7865));
  jor  g07802(.dina(n7865), .dinb(n7776), .dout(n7866));
  jxor g07803(.dina(n7728), .dinb(n7720), .dout(n7867));
  jand g07804(.dina(n7867), .dinb(n7866), .dout(n7868));
  jnot g07805(.din(n7868), .dout(n7869));
  jxor g07806(.dina(n7867), .dinb(n7866), .dout(n7870));
  jnot g07807(.din(n7870), .dout(n7871));
  jand g07808(.dina(n6936), .dinb(n4446), .dout(n7872));
  jand g07809(.dina(n7741), .dinb(n4451), .dout(n7873));
  jand g07810(.dina(n7613), .dinb(n4358), .dout(n7874));
  jand g07811(.dina(n6934), .dinb(n3853), .dout(n7875));
  jor  g07812(.dina(n7875), .dinb(n7874), .dout(n7876));
  jor  g07813(.dina(n7876), .dinb(n7873), .dout(n7877));
  jor  g07814(.dina(n7877), .dinb(n7872), .dout(n7878));
  jxor g07815(.dina(n7878), .dinb(n5292), .dout(n7879));
  jor  g07816(.dina(n7879), .dinb(n7871), .dout(n7880));
  jand g07817(.dina(n7880), .dinb(n7869), .dout(n7881));
  jxor g07818(.dina(\a[10] ), .dinb(\a[9] ), .dout(n7882));
  jnot g07819(.din(n7882), .dout(n7883));
  jxor g07820(.dina(\a[9] ), .dinb(\a[8] ), .dout(n7884));
  jnot g07821(.din(n7884), .dout(n7885));
  jand g07822(.dina(n7885), .dinb(n7883), .dout(n7886));
  jxor g07823(.dina(\a[11] ), .dinb(\a[10] ), .dout(n7887));
  jand g07824(.dina(n7887), .dinb(n7886), .dout(n7888));
  jnot g07825(.din(n7888), .dout(n7889));
  jand g07826(.dina(n7887), .dinb(n7884), .dout(n7890));
  jnot g07827(.din(n7890), .dout(n7891));
  jor  g07828(.dina(n7891), .dinb(n4728), .dout(n7892));
  jand g07829(.dina(n7892), .dinb(n7889), .dout(n7893));
  jor  g07830(.dina(n7893), .dinb(n4630), .dout(n7894));
  jxor g07831(.dina(n7894), .dinb(\a[11] ), .dout(n7895));
  jor  g07832(.dina(n7895), .dinb(n7881), .dout(n7896));
  jxor g07833(.dina(n7895), .dinb(n7881), .dout(n7897));
  jxor g07834(.dina(n7746), .dinb(n7736), .dout(n7898));
  jand g07835(.dina(n7898), .dinb(n7897), .dout(n7899));
  jnot g07836(.din(n7899), .dout(n7900));
  jand g07837(.dina(n7900), .dinb(n7896), .dout(n7901));
  jnot g07838(.din(n7901), .dout(n7902));
  jxor g07839(.dina(n7759), .dinb(n7758), .dout(n7903));
  jand g07840(.dina(n7903), .dinb(n7902), .dout(n7904));
  jxor g07841(.dina(n7864), .dinb(n7863), .dout(n7905));
  jnot g07842(.din(n7905), .dout(n7906));
  jand g07843(.dina(n6936), .dinb(n4545), .dout(n7907));
  jand g07844(.dina(n6934), .dinb(n922), .dout(n7908));
  jand g07845(.dina(n7613), .dinb(n3853), .dout(n7909));
  jand g07846(.dina(n7741), .dinb(n4358), .dout(n7910));
  jor  g07847(.dina(n7910), .dinb(n7909), .dout(n7911));
  jor  g07848(.dina(n7911), .dinb(n7908), .dout(n7912));
  jor  g07849(.dina(n7912), .dinb(n7907), .dout(n7913));
  jxor g07850(.dina(n7913), .dinb(n5292), .dout(n7914));
  jor  g07851(.dina(n7914), .dinb(n7906), .dout(n7915));
  jxor g07852(.dina(n7829), .dinb(n7828), .dout(n7916));
  jnot g07853(.din(n7916), .dout(n7917));
  jand g07854(.dina(n5693), .dinb(n5092), .dout(n7918));
  jand g07855(.dina(n6131), .dinb(n1862), .dout(n7919));
  jand g07856(.dina(n5691), .dinb(n1956), .dout(n7920));
  jand g07857(.dina(n6209), .dinb(n1776), .dout(n7921));
  jor  g07858(.dina(n7921), .dinb(n7920), .dout(n7922));
  jor  g07859(.dina(n7922), .dinb(n7919), .dout(n7923));
  jor  g07860(.dina(n7923), .dinb(n7918), .dout(n7924));
  jxor g07861(.dina(n7924), .dinb(n4247), .dout(n7925));
  jor  g07862(.dina(n7925), .dinb(n7917), .dout(n7926));
  jor  g07863(.dina(n6976), .dinb(n4724), .dout(n7927));
  jor  g07864(.dina(n4735), .dinb(n2953), .dout(n7928));
  jor  g07865(.dina(n4733), .dinb(n2990), .dout(n7929));
  jor  g07866(.dina(n4905), .dinb(n2866), .dout(n7930));
  jand g07867(.dina(n7930), .dinb(n7929), .dout(n7931));
  jand g07868(.dina(n7931), .dinb(n7928), .dout(n7932));
  jand g07869(.dina(n7932), .dinb(n7927), .dout(n7933));
  jxor g07870(.dina(n7933), .dinb(\a[29] ), .dout(n7934));
  jnot g07871(.din(n7934), .dout(n7935));
  jxor g07872(.dina(n7493), .dinb(n7492), .dout(n7936));
  jand g07873(.dina(n7936), .dinb(n7935), .dout(n7937));
  jor  g07874(.dina(n6988), .dinb(n4724), .dout(n7938));
  jor  g07875(.dina(n4733), .dinb(n3085), .dout(n7939));
  jor  g07876(.dina(n4905), .dinb(n2953), .dout(n7940));
  jor  g07877(.dina(n4735), .dinb(n2990), .dout(n7941));
  jand g07878(.dina(n7941), .dinb(n7940), .dout(n7942));
  jand g07879(.dina(n7942), .dinb(n7939), .dout(n7943));
  jand g07880(.dina(n7943), .dinb(n7938), .dout(n7944));
  jxor g07881(.dina(n7944), .dinb(\a[29] ), .dout(n7945));
  jnot g07882(.din(n7945), .dout(n7946));
  jxor g07883(.dina(n7488), .dinb(n7487), .dout(n7947));
  jand g07884(.dina(n7947), .dinb(n7946), .dout(n7948));
  jor  g07885(.dina(n6681), .dinb(n4724), .dout(n7949));
  jor  g07886(.dina(n4735), .dinb(n3085), .dout(n7950));
  jor  g07887(.dina(n4905), .dinb(n2990), .dout(n7951));
  jor  g07888(.dina(n4733), .dinb(n3182), .dout(n7952));
  jand g07889(.dina(n7952), .dinb(n7951), .dout(n7953));
  jand g07890(.dina(n7953), .dinb(n7950), .dout(n7954));
  jand g07891(.dina(n7954), .dinb(n7949), .dout(n7955));
  jxor g07892(.dina(n7955), .dinb(\a[29] ), .dout(n7956));
  jnot g07893(.din(n7956), .dout(n7957));
  jxor g07894(.dina(n7483), .dinb(n7482), .dout(n7958));
  jand g07895(.dina(n7958), .dinb(n7957), .dout(n7959));
  jor  g07896(.dina(n7031), .dinb(n4724), .dout(n7960));
  jor  g07897(.dina(n4905), .dinb(n3085), .dout(n7961));
  jnot g07898(.din(n3275), .dout(n7962));
  jor  g07899(.dina(n4733), .dinb(n7962), .dout(n7963));
  jor  g07900(.dina(n4735), .dinb(n3182), .dout(n7964));
  jand g07901(.dina(n7964), .dinb(n7963), .dout(n7965));
  jand g07902(.dina(n7965), .dinb(n7961), .dout(n7966));
  jand g07903(.dina(n7966), .dinb(n7960), .dout(n7967));
  jxor g07904(.dina(n7967), .dinb(\a[29] ), .dout(n7968));
  jnot g07905(.din(n7968), .dout(n7969));
  jxor g07906(.dina(n7478), .dinb(n7477), .dout(n7970));
  jand g07907(.dina(n7970), .dinb(n7969), .dout(n7971));
  jor  g07908(.dina(n7076), .dinb(n4724), .dout(n7972));
  jor  g07909(.dina(n4735), .dinb(n7962), .dout(n7973));
  jor  g07910(.dina(n4905), .dinb(n3182), .dout(n7974));
  jor  g07911(.dina(n4733), .dinb(n3684), .dout(n7975));
  jand g07912(.dina(n7975), .dinb(n7974), .dout(n7976));
  jand g07913(.dina(n7976), .dinb(n7973), .dout(n7977));
  jand g07914(.dina(n7977), .dinb(n7972), .dout(n7978));
  jxor g07915(.dina(n7978), .dinb(\a[29] ), .dout(n7979));
  jnot g07916(.din(n7979), .dout(n7980));
  jxor g07917(.dina(n7474), .dinb(n7464), .dout(n7981));
  jand g07918(.dina(n7981), .dinb(n7980), .dout(n7982));
  jor  g07919(.dina(n7131), .dinb(n4724), .dout(n7983));
  jor  g07920(.dina(n4905), .dinb(n7962), .dout(n7984));
  jor  g07921(.dina(n4733), .dinb(n3414), .dout(n7985));
  jor  g07922(.dina(n4735), .dinb(n3684), .dout(n7986));
  jand g07923(.dina(n7986), .dinb(n7985), .dout(n7987));
  jand g07924(.dina(n7987), .dinb(n7984), .dout(n7988));
  jand g07925(.dina(n7988), .dinb(n7983), .dout(n7989));
  jxor g07926(.dina(n7989), .dinb(\a[29] ), .dout(n7990));
  jnot g07927(.din(n7990), .dout(n7991));
  jxor g07928(.dina(n7415), .dinb(n7362), .dout(n7992));
  jand g07929(.dina(n7992), .dinb(n7991), .dout(n7993));
  jor  g07930(.dina(n7177), .dinb(n4724), .dout(n7994));
  jor  g07931(.dina(n4733), .dinb(n3516), .dout(n7995));
  jor  g07932(.dina(n4905), .dinb(n3684), .dout(n7996));
  jor  g07933(.dina(n4735), .dinb(n3414), .dout(n7997));
  jand g07934(.dina(n7997), .dinb(n7996), .dout(n7998));
  jand g07935(.dina(n7998), .dinb(n7995), .dout(n7999));
  jand g07936(.dina(n7999), .dinb(n7994), .dout(n8000));
  jxor g07937(.dina(n8000), .dinb(\a[29] ), .dout(n8001));
  jnot g07938(.din(n8001), .dout(n8002));
  jxor g07939(.dina(n3677), .dinb(n7411), .dout(n8003));
  jnot g07940(.din(n8003), .dout(n8004));
  jand g07941(.dina(n8004), .dinb(n732), .dout(n8005));
  jand g07942(.dina(n3858), .dinb(n7411), .dout(n8006));
  jand g07943(.dina(n3855), .dinb(n7405), .dout(n8007));
  jor  g07944(.dina(n8007), .dinb(n8006), .dout(n8008));
  jor  g07945(.dina(n8008), .dinb(n8005), .dout(n8009));
  jand g07946(.dina(n8009), .dinb(n8002), .dout(n8010));
  jand g07947(.dina(n7411), .dinb(n731), .dout(n8011));
  jand g07948(.dina(n8004), .dinb(n4449), .dout(n8012));
  jand g07949(.dina(n4457), .dinb(n7411), .dout(n8013));
  jand g07950(.dina(n4453), .dinb(n7405), .dout(n8014));
  jor  g07951(.dina(n8014), .dinb(n8013), .dout(n8015));
  jor  g07952(.dina(n8015), .dinb(n8012), .dout(n8016));
  jnot g07953(.din(n8016), .dout(n8017));
  jand g07954(.dina(n4447), .dinb(n7411), .dout(n8018));
  jnot g07955(.din(n8018), .dout(n8019));
  jand g07956(.dina(n8019), .dinb(\a[29] ), .dout(n8020));
  jand g07957(.dina(n8020), .dinb(n8017), .dout(n8021));
  jand g07958(.dina(n7407), .dinb(n4449), .dout(n8022));
  jand g07959(.dina(n4453), .dinb(n7326), .dout(n8023));
  jand g07960(.dina(n4461), .dinb(n7411), .dout(n8024));
  jand g07961(.dina(n4457), .dinb(n7405), .dout(n8025));
  jor  g07962(.dina(n8025), .dinb(n8024), .dout(n8026));
  jor  g07963(.dina(n8026), .dinb(n8023), .dout(n8027));
  jor  g07964(.dina(n8027), .dinb(n8022), .dout(n8028));
  jnot g07965(.din(n8028), .dout(n8029));
  jand g07966(.dina(n8029), .dinb(n8021), .dout(n8030));
  jand g07967(.dina(n8030), .dinb(n8011), .dout(n8031));
  jor  g07968(.dina(n7466), .dinb(n4724), .dout(n8032));
  jor  g07969(.dina(n4735), .dinb(n3516), .dout(n8033));
  jor  g07970(.dina(n4905), .dinb(n3414), .dout(n8034));
  jor  g07971(.dina(n4733), .dinb(n3677), .dout(n8035));
  jand g07972(.dina(n8035), .dinb(n8034), .dout(n8036));
  jand g07973(.dina(n8036), .dinb(n8033), .dout(n8037));
  jand g07974(.dina(n8037), .dinb(n8032), .dout(n8038));
  jxor g07975(.dina(n8038), .dinb(\a[29] ), .dout(n8039));
  jnot g07976(.din(n8039), .dout(n8040));
  jxor g07977(.dina(n8030), .dinb(n8011), .dout(n8041));
  jand g07978(.dina(n8041), .dinb(n8040), .dout(n8042));
  jor  g07979(.dina(n8042), .dinb(n8031), .dout(n8043));
  jxor g07980(.dina(n8009), .dinb(n8002), .dout(n8044));
  jand g07981(.dina(n8044), .dinb(n8043), .dout(n8045));
  jor  g07982(.dina(n8045), .dinb(n8010), .dout(n8046));
  jxor g07983(.dina(n7992), .dinb(n7991), .dout(n8047));
  jand g07984(.dina(n8047), .dinb(n8046), .dout(n8048));
  jor  g07985(.dina(n8048), .dinb(n7993), .dout(n8049));
  jxor g07986(.dina(n7981), .dinb(n7980), .dout(n8050));
  jand g07987(.dina(n8050), .dinb(n8049), .dout(n8051));
  jor  g07988(.dina(n8051), .dinb(n7982), .dout(n8052));
  jxor g07989(.dina(n7970), .dinb(n7969), .dout(n8053));
  jand g07990(.dina(n8053), .dinb(n8052), .dout(n8054));
  jor  g07991(.dina(n8054), .dinb(n7971), .dout(n8055));
  jxor g07992(.dina(n7958), .dinb(n7957), .dout(n8056));
  jand g07993(.dina(n8056), .dinb(n8055), .dout(n8057));
  jor  g07994(.dina(n8057), .dinb(n7959), .dout(n8058));
  jxor g07995(.dina(n7947), .dinb(n7946), .dout(n8059));
  jand g07996(.dina(n8059), .dinb(n8058), .dout(n8060));
  jor  g07997(.dina(n8060), .dinb(n7948), .dout(n8061));
  jxor g07998(.dina(n7936), .dinb(n7935), .dout(n8062));
  jand g07999(.dina(n8062), .dinb(n8061), .dout(n8063));
  jor  g08000(.dina(n8063), .dinb(n7937), .dout(n8064));
  jxor g08001(.dina(n7510), .dinb(n7502), .dout(n8065));
  jand g08002(.dina(n8065), .dinb(n8064), .dout(n8066));
  jor  g08003(.dina(n6464), .dinb(n4747), .dout(n8067));
  jor  g08004(.dina(n4959), .dinb(n2601), .dout(n8068));
  jor  g08005(.dina(n4919), .dinb(n2694), .dout(n8069));
  jor  g08006(.dina(n4746), .dinb(n2731), .dout(n8070));
  jand g08007(.dina(n8070), .dinb(n8069), .dout(n8071));
  jand g08008(.dina(n8071), .dinb(n8068), .dout(n8072));
  jand g08009(.dina(n8072), .dinb(n8067), .dout(n8073));
  jxor g08010(.dina(n8073), .dinb(\a[26] ), .dout(n8074));
  jnot g08011(.din(n8074), .dout(n8075));
  jxor g08012(.dina(n8065), .dinb(n8064), .dout(n8076));
  jand g08013(.dina(n8076), .dinb(n8075), .dout(n8077));
  jor  g08014(.dina(n8077), .dinb(n8066), .dout(n8078));
  jxor g08015(.dina(n7809), .dinb(n7801), .dout(n8079));
  jand g08016(.dina(n8079), .dinb(n8078), .dout(n8080));
  jnot g08017(.din(n8080), .dout(n8081));
  jxor g08018(.dina(n8079), .dinb(n8078), .dout(n8082));
  jnot g08019(.din(n8082), .dout(n8083));
  jand g08020(.dina(n5844), .dinb(n5365), .dout(n8084));
  jand g08021(.dina(n5363), .dinb(n2411), .dout(n8085));
  jand g08022(.dina(n5500), .dinb(n2237), .dout(n8086));
  jand g08023(.dina(n5424), .dinb(n2343), .dout(n8087));
  jor  g08024(.dina(n8087), .dinb(n8086), .dout(n8088));
  jor  g08025(.dina(n8088), .dinb(n8085), .dout(n8089));
  jor  g08026(.dina(n8089), .dinb(n8084), .dout(n8090));
  jxor g08027(.dina(n8090), .dinb(n72), .dout(n8091));
  jor  g08028(.dina(n8091), .dinb(n8083), .dout(n8092));
  jand g08029(.dina(n8092), .dinb(n8081), .dout(n8093));
  jnot g08030(.din(n8093), .dout(n8094));
  jxor g08031(.dina(n7825), .dinb(n7817), .dout(n8095));
  jand g08032(.dina(n8095), .dinb(n8094), .dout(n8096));
  jnot g08033(.din(n8096), .dout(n8097));
  jxor g08034(.dina(n8095), .dinb(n8094), .dout(n8098));
  jnot g08035(.din(n8098), .dout(n8099));
  jand g08036(.dina(n5693), .dinb(n5440), .dout(n8100));
  jand g08037(.dina(n6131), .dinb(n1956), .dout(n8101));
  jand g08038(.dina(n6209), .dinb(n1862), .dout(n8102));
  jand g08039(.dina(n5691), .dinb(n2067), .dout(n8103));
  jor  g08040(.dina(n8103), .dinb(n8102), .dout(n8104));
  jor  g08041(.dina(n8104), .dinb(n8101), .dout(n8105));
  jor  g08042(.dina(n8105), .dinb(n8100), .dout(n8106));
  jxor g08043(.dina(n8106), .dinb(n4247), .dout(n8107));
  jor  g08044(.dina(n8107), .dinb(n8099), .dout(n8108));
  jand g08045(.dina(n8108), .dinb(n8097), .dout(n8109));
  jnot g08046(.din(n8109), .dout(n8110));
  jxor g08047(.dina(n7925), .dinb(n7917), .dout(n8111));
  jand g08048(.dina(n8111), .dinb(n8110), .dout(n8112));
  jnot g08049(.din(n8112), .dout(n8113));
  jand g08050(.dina(n8113), .dinb(n7926), .dout(n8114));
  jnot g08051(.din(n8114), .dout(n8115));
  jxor g08052(.dina(n7844), .dinb(n7836), .dout(n8116));
  jand g08053(.dina(n8116), .dinb(n8115), .dout(n8117));
  jnot g08054(.din(n8117), .dout(n8118));
  jxor g08055(.dina(n8116), .dinb(n8115), .dout(n8119));
  jnot g08056(.din(n8119), .dout(n8120));
  jand g08057(.dina(n6340), .dinb(n4258), .dout(n8121));
  jand g08058(.dina(n6798), .dinb(n1343), .dout(n8122));
  jand g08059(.dina(n6556), .dinb(n1445), .dout(n8123));
  jand g08060(.dina(n6338), .dinb(n1560), .dout(n8124));
  jor  g08061(.dina(n8124), .dinb(n8123), .dout(n8125));
  jor  g08062(.dina(n8125), .dinb(n8122), .dout(n8126));
  jor  g08063(.dina(n8126), .dinb(n8121), .dout(n8127));
  jxor g08064(.dina(n8127), .dinb(n5064), .dout(n8128));
  jor  g08065(.dina(n8128), .dinb(n8120), .dout(n8129));
  jand g08066(.dina(n8129), .dinb(n8118), .dout(n8130));
  jnot g08067(.din(n8130), .dout(n8131));
  jxor g08068(.dina(n7860), .dinb(n7852), .dout(n8132));
  jand g08069(.dina(n8132), .dinb(n8131), .dout(n8133));
  jnot g08070(.din(n8133), .dout(n8134));
  jxor g08071(.dina(n8132), .dinb(n8131), .dout(n8135));
  jnot g08072(.din(n8135), .dout(n8136));
  jand g08073(.dina(n6936), .dinb(n3848), .dout(n8137));
  jand g08074(.dina(n7613), .dinb(n922), .dout(n8138));
  jand g08075(.dina(n7741), .dinb(n3853), .dout(n8139));
  jand g08076(.dina(n6934), .dinb(n1076), .dout(n8140));
  jor  g08077(.dina(n8140), .dinb(n8139), .dout(n8141));
  jor  g08078(.dina(n8141), .dinb(n8138), .dout(n8142));
  jor  g08079(.dina(n8142), .dinb(n8137), .dout(n8143));
  jxor g08080(.dina(n8143), .dinb(n5292), .dout(n8144));
  jor  g08081(.dina(n8144), .dinb(n8136), .dout(n8145));
  jand g08082(.dina(n8145), .dinb(n8134), .dout(n8146));
  jnot g08083(.din(n8146), .dout(n8147));
  jxor g08084(.dina(n7914), .dinb(n7906), .dout(n8148));
  jand g08085(.dina(n8148), .dinb(n8147), .dout(n8149));
  jnot g08086(.din(n8149), .dout(n8150));
  jand g08087(.dina(n8150), .dinb(n7915), .dout(n8151));
  jor  g08088(.dina(n7891), .dinb(n4731), .dout(n8152));
  jor  g08089(.dina(n7889), .dinb(n4597), .dout(n8153));
  jand g08090(.dina(n7885), .dinb(n7882), .dout(n8154));
  jnot g08091(.din(n8154), .dout(n8155));
  jor  g08092(.dina(n8155), .dinb(n4630), .dout(n8156));
  jand g08093(.dina(n8156), .dinb(n8153), .dout(n8157));
  jand g08094(.dina(n8157), .dinb(n8152), .dout(n8158));
  jxor g08095(.dina(n8158), .dinb(\a[11] ), .dout(n8159));
  jor  g08096(.dina(n8159), .dinb(n8151), .dout(n8160));
  jxor g08097(.dina(n8159), .dinb(n8151), .dout(n8161));
  jxor g08098(.dina(n7879), .dinb(n7871), .dout(n8162));
  jand g08099(.dina(n8162), .dinb(n8161), .dout(n8163));
  jnot g08100(.din(n8163), .dout(n8164));
  jand g08101(.dina(n8164), .dinb(n8160), .dout(n8165));
  jnot g08102(.din(n8165), .dout(n8166));
  jxor g08103(.dina(n7898), .dinb(n7897), .dout(n8167));
  jand g08104(.dina(n8167), .dinb(n8166), .dout(n8168));
  jxor g08105(.dina(n8167), .dinb(n8166), .dout(n8169));
  jand g08106(.dina(n6340), .dinb(n4866), .dout(n8170));
  jand g08107(.dina(n6798), .dinb(n1445), .dout(n8171));
  jand g08108(.dina(n6556), .dinb(n1560), .dout(n8172));
  jand g08109(.dina(n6338), .dinb(n1624), .dout(n8173));
  jor  g08110(.dina(n8173), .dinb(n8172), .dout(n8174));
  jor  g08111(.dina(n8174), .dinb(n8171), .dout(n8175));
  jor  g08112(.dina(n8175), .dinb(n8170), .dout(n8176));
  jxor g08113(.dina(n8176), .dinb(n5064), .dout(n8177));
  jnot g08114(.din(n8177), .dout(n8178));
  jxor g08115(.dina(n8111), .dinb(n8110), .dout(n8179));
  jand g08116(.dina(n8179), .dinb(n8178), .dout(n8180));
  jxor g08117(.dina(n8062), .dinb(n8061), .dout(n8181));
  jnot g08118(.din(n8181), .dout(n8182));
  jand g08119(.dina(n6591), .dinb(n75), .dout(n8183));
  jand g08120(.dina(n4933), .dinb(n2695), .dout(n8184));
  jand g08121(.dina(n4745), .dinb(n2808), .dout(n8185));
  jand g08122(.dina(n4918), .dinb(n2732), .dout(n8186));
  jor  g08123(.dina(n8186), .dinb(n8185), .dout(n8187));
  jor  g08124(.dina(n8187), .dinb(n8184), .dout(n8188));
  jor  g08125(.dina(n8188), .dinb(n8183), .dout(n8189));
  jxor g08126(.dina(n8189), .dinb(n68), .dout(n8190));
  jor  g08127(.dina(n8190), .dinb(n8182), .dout(n8191));
  jxor g08128(.dina(n8059), .dinb(n8058), .dout(n8192));
  jnot g08129(.din(n8192), .dout(n8193));
  jand g08130(.dina(n6439), .dinb(n75), .dout(n8194));
  jand g08131(.dina(n4918), .dinb(n2808), .dout(n8195));
  jand g08132(.dina(n4933), .dinb(n2732), .dout(n8196));
  jand g08133(.dina(n4745), .dinb(n2867), .dout(n8197));
  jor  g08134(.dina(n8197), .dinb(n8196), .dout(n8198));
  jor  g08135(.dina(n8198), .dinb(n8195), .dout(n8199));
  jor  g08136(.dina(n8199), .dinb(n8194), .dout(n8200));
  jxor g08137(.dina(n8200), .dinb(n68), .dout(n8201));
  jor  g08138(.dina(n8201), .dinb(n8193), .dout(n8202));
  jxor g08139(.dina(n8056), .dinb(n8055), .dout(n8203));
  jnot g08140(.din(n8203), .dout(n8204));
  jand g08141(.dina(n6706), .dinb(n75), .dout(n8205));
  jand g08142(.dina(n4933), .dinb(n2808), .dout(n8206));
  jand g08143(.dina(n4745), .dinb(n2954), .dout(n8207));
  jand g08144(.dina(n4918), .dinb(n2867), .dout(n8208));
  jor  g08145(.dina(n8208), .dinb(n8207), .dout(n8209));
  jor  g08146(.dina(n8209), .dinb(n8206), .dout(n8210));
  jor  g08147(.dina(n8210), .dinb(n8205), .dout(n8211));
  jxor g08148(.dina(n8211), .dinb(n68), .dout(n8212));
  jor  g08149(.dina(n8212), .dinb(n8204), .dout(n8213));
  jxor g08150(.dina(n8053), .dinb(n8052), .dout(n8214));
  jnot g08151(.din(n8214), .dout(n8215));
  jor  g08152(.dina(n6976), .dinb(n4747), .dout(n8216));
  jor  g08153(.dina(n4919), .dinb(n2953), .dout(n8217));
  jor  g08154(.dina(n4746), .dinb(n2990), .dout(n8218));
  jor  g08155(.dina(n4959), .dinb(n2866), .dout(n8219));
  jand g08156(.dina(n8219), .dinb(n8218), .dout(n8220));
  jand g08157(.dina(n8220), .dinb(n8217), .dout(n8221));
  jand g08158(.dina(n8221), .dinb(n8216), .dout(n8222));
  jxor g08159(.dina(n8222), .dinb(\a[26] ), .dout(n8223));
  jor  g08160(.dina(n8223), .dinb(n8215), .dout(n8224));
  jxor g08161(.dina(n8050), .dinb(n8049), .dout(n8225));
  jnot g08162(.din(n8225), .dout(n8226));
  jor  g08163(.dina(n6988), .dinb(n4747), .dout(n8227));
  jor  g08164(.dina(n4746), .dinb(n3085), .dout(n8228));
  jor  g08165(.dina(n4959), .dinb(n2953), .dout(n8229));
  jor  g08166(.dina(n4919), .dinb(n2990), .dout(n8230));
  jand g08167(.dina(n8230), .dinb(n8229), .dout(n8231));
  jand g08168(.dina(n8231), .dinb(n8228), .dout(n8232));
  jand g08169(.dina(n8232), .dinb(n8227), .dout(n8233));
  jxor g08170(.dina(n8233), .dinb(\a[26] ), .dout(n8234));
  jor  g08171(.dina(n8234), .dinb(n8226), .dout(n8235));
  jxor g08172(.dina(n8047), .dinb(n8046), .dout(n8236));
  jnot g08173(.din(n8236), .dout(n8237));
  jor  g08174(.dina(n6681), .dinb(n4747), .dout(n8238));
  jor  g08175(.dina(n4919), .dinb(n3085), .dout(n8239));
  jor  g08176(.dina(n4959), .dinb(n2990), .dout(n8240));
  jor  g08177(.dina(n4746), .dinb(n3182), .dout(n8241));
  jand g08178(.dina(n8241), .dinb(n8240), .dout(n8242));
  jand g08179(.dina(n8242), .dinb(n8239), .dout(n8243));
  jand g08180(.dina(n8243), .dinb(n8238), .dout(n8244));
  jxor g08181(.dina(n8244), .dinb(\a[26] ), .dout(n8245));
  jor  g08182(.dina(n8245), .dinb(n8237), .dout(n8246));
  jor  g08183(.dina(n7031), .dinb(n4747), .dout(n8247));
  jor  g08184(.dina(n4959), .dinb(n3085), .dout(n8248));
  jor  g08185(.dina(n4746), .dinb(n7962), .dout(n8249));
  jor  g08186(.dina(n4919), .dinb(n3182), .dout(n8250));
  jand g08187(.dina(n8250), .dinb(n8249), .dout(n8251));
  jand g08188(.dina(n8251), .dinb(n8248), .dout(n8252));
  jand g08189(.dina(n8252), .dinb(n8247), .dout(n8253));
  jxor g08190(.dina(n8253), .dinb(\a[26] ), .dout(n8254));
  jnot g08191(.din(n8254), .dout(n8255));
  jxor g08192(.dina(n8044), .dinb(n8043), .dout(n8256));
  jand g08193(.dina(n8256), .dinb(n8255), .dout(n8257));
  jor  g08194(.dina(n7076), .dinb(n4747), .dout(n8258));
  jor  g08195(.dina(n4919), .dinb(n7962), .dout(n8259));
  jor  g08196(.dina(n4959), .dinb(n3182), .dout(n8260));
  jor  g08197(.dina(n4746), .dinb(n3684), .dout(n8261));
  jand g08198(.dina(n8261), .dinb(n8260), .dout(n8262));
  jand g08199(.dina(n8262), .dinb(n8259), .dout(n8263));
  jand g08200(.dina(n8263), .dinb(n8258), .dout(n8264));
  jxor g08201(.dina(n8264), .dinb(\a[26] ), .dout(n8265));
  jnot g08202(.din(n8265), .dout(n8266));
  jxor g08203(.dina(n8041), .dinb(n8040), .dout(n8267));
  jand g08204(.dina(n8267), .dinb(n8266), .dout(n8268));
  jor  g08205(.dina(n7131), .dinb(n4747), .dout(n8269));
  jor  g08206(.dina(n4959), .dinb(n7962), .dout(n8270));
  jor  g08207(.dina(n4746), .dinb(n3414), .dout(n8271));
  jor  g08208(.dina(n4919), .dinb(n3684), .dout(n8272));
  jand g08209(.dina(n8272), .dinb(n8271), .dout(n8273));
  jand g08210(.dina(n8273), .dinb(n8270), .dout(n8274));
  jand g08211(.dina(n8274), .dinb(n8269), .dout(n8275));
  jxor g08212(.dina(n8275), .dinb(\a[26] ), .dout(n8276));
  jnot g08213(.din(n8276), .dout(n8277));
  jor  g08214(.dina(n8021), .dinb(n88), .dout(n8278));
  jxor g08215(.dina(n8278), .dinb(n8029), .dout(n8279));
  jand g08216(.dina(n8279), .dinb(n8277), .dout(n8280));
  jor  g08217(.dina(n7177), .dinb(n4747), .dout(n8281));
  jor  g08218(.dina(n4746), .dinb(n3516), .dout(n8282));
  jor  g08219(.dina(n4959), .dinb(n3684), .dout(n8283));
  jor  g08220(.dina(n4919), .dinb(n3414), .dout(n8284));
  jand g08221(.dina(n8284), .dinb(n8283), .dout(n8285));
  jand g08222(.dina(n8285), .dinb(n8282), .dout(n8286));
  jand g08223(.dina(n8286), .dinb(n8281), .dout(n8287));
  jxor g08224(.dina(n8287), .dinb(\a[26] ), .dout(n8288));
  jnot g08225(.din(n8288), .dout(n8289));
  jand g08226(.dina(n8018), .dinb(\a[29] ), .dout(n8290));
  jxor g08227(.dina(n8290), .dinb(n8016), .dout(n8291));
  jand g08228(.dina(n8291), .dinb(n8289), .dout(n8292));
  jand g08229(.dina(n8004), .dinb(n75), .dout(n8293));
  jand g08230(.dina(n4918), .dinb(n7411), .dout(n8294));
  jand g08231(.dina(n4933), .dinb(n7405), .dout(n8295));
  jor  g08232(.dina(n8295), .dinb(n8294), .dout(n8296));
  jor  g08233(.dina(n8296), .dinb(n8293), .dout(n8297));
  jnot g08234(.din(n8297), .dout(n8298));
  jand g08235(.dina(n7411), .dinb(n74), .dout(n8299));
  jnot g08236(.din(n8299), .dout(n8300));
  jand g08237(.dina(n8300), .dinb(\a[26] ), .dout(n8301));
  jand g08238(.dina(n8301), .dinb(n8298), .dout(n8302));
  jand g08239(.dina(n7407), .dinb(n75), .dout(n8303));
  jand g08240(.dina(n4933), .dinb(n7326), .dout(n8304));
  jand g08241(.dina(n4745), .dinb(n7411), .dout(n8305));
  jand g08242(.dina(n4918), .dinb(n7405), .dout(n8306));
  jor  g08243(.dina(n8306), .dinb(n8305), .dout(n8307));
  jor  g08244(.dina(n8307), .dinb(n8304), .dout(n8308));
  jor  g08245(.dina(n8308), .dinb(n8303), .dout(n8309));
  jnot g08246(.din(n8309), .dout(n8310));
  jand g08247(.dina(n8310), .dinb(n8302), .dout(n8311));
  jand g08248(.dina(n8311), .dinb(n8018), .dout(n8312));
  jor  g08249(.dina(n7466), .dinb(n4747), .dout(n8313));
  jor  g08250(.dina(n4919), .dinb(n3516), .dout(n8314));
  jor  g08251(.dina(n4959), .dinb(n3414), .dout(n8315));
  jor  g08252(.dina(n4746), .dinb(n3677), .dout(n8316));
  jand g08253(.dina(n8316), .dinb(n8315), .dout(n8317));
  jand g08254(.dina(n8317), .dinb(n8314), .dout(n8318));
  jand g08255(.dina(n8318), .dinb(n8313), .dout(n8319));
  jxor g08256(.dina(n8319), .dinb(\a[26] ), .dout(n8320));
  jnot g08257(.din(n8320), .dout(n8321));
  jxor g08258(.dina(n8311), .dinb(n8018), .dout(n8322));
  jand g08259(.dina(n8322), .dinb(n8321), .dout(n8323));
  jor  g08260(.dina(n8323), .dinb(n8312), .dout(n8324));
  jxor g08261(.dina(n8291), .dinb(n8289), .dout(n8325));
  jand g08262(.dina(n8325), .dinb(n8324), .dout(n8326));
  jor  g08263(.dina(n8326), .dinb(n8292), .dout(n8327));
  jxor g08264(.dina(n8279), .dinb(n8277), .dout(n8328));
  jand g08265(.dina(n8328), .dinb(n8327), .dout(n8329));
  jor  g08266(.dina(n8329), .dinb(n8280), .dout(n8330));
  jxor g08267(.dina(n8267), .dinb(n8266), .dout(n8331));
  jand g08268(.dina(n8331), .dinb(n8330), .dout(n8332));
  jor  g08269(.dina(n8332), .dinb(n8268), .dout(n8333));
  jxor g08270(.dina(n8256), .dinb(n8255), .dout(n8334));
  jand g08271(.dina(n8334), .dinb(n8333), .dout(n8335));
  jor  g08272(.dina(n8335), .dinb(n8257), .dout(n8336));
  jxor g08273(.dina(n8245), .dinb(n8237), .dout(n8337));
  jand g08274(.dina(n8337), .dinb(n8336), .dout(n8338));
  jnot g08275(.din(n8338), .dout(n8339));
  jand g08276(.dina(n8339), .dinb(n8246), .dout(n8340));
  jnot g08277(.din(n8340), .dout(n8341));
  jxor g08278(.dina(n8234), .dinb(n8226), .dout(n8342));
  jand g08279(.dina(n8342), .dinb(n8341), .dout(n8343));
  jnot g08280(.din(n8343), .dout(n8344));
  jand g08281(.dina(n8344), .dinb(n8235), .dout(n8345));
  jnot g08282(.din(n8345), .dout(n8346));
  jxor g08283(.dina(n8223), .dinb(n8215), .dout(n8347));
  jand g08284(.dina(n8347), .dinb(n8346), .dout(n8348));
  jnot g08285(.din(n8348), .dout(n8349));
  jand g08286(.dina(n8349), .dinb(n8224), .dout(n8350));
  jnot g08287(.din(n8350), .dout(n8351));
  jxor g08288(.dina(n8212), .dinb(n8204), .dout(n8352));
  jand g08289(.dina(n8352), .dinb(n8351), .dout(n8353));
  jnot g08290(.din(n8353), .dout(n8354));
  jand g08291(.dina(n8354), .dinb(n8213), .dout(n8355));
  jnot g08292(.din(n8355), .dout(n8356));
  jxor g08293(.dina(n8201), .dinb(n8193), .dout(n8357));
  jand g08294(.dina(n8357), .dinb(n8356), .dout(n8358));
  jnot g08295(.din(n8358), .dout(n8359));
  jand g08296(.dina(n8359), .dinb(n8202), .dout(n8360));
  jnot g08297(.din(n8360), .dout(n8361));
  jxor g08298(.dina(n8190), .dinb(n8182), .dout(n8362));
  jand g08299(.dina(n8362), .dinb(n8361), .dout(n8363));
  jnot g08300(.din(n8363), .dout(n8364));
  jand g08301(.dina(n8364), .dinb(n8191), .dout(n8365));
  jnot g08302(.din(n8365), .dout(n8366));
  jxor g08303(.dina(n8076), .dinb(n8075), .dout(n8367));
  jand g08304(.dina(n8367), .dinb(n8366), .dout(n8368));
  jand g08305(.dina(n5861), .dinb(n5365), .dout(n8369));
  jand g08306(.dina(n5424), .dinb(n2411), .dout(n8370));
  jand g08307(.dina(n5500), .dinb(n2343), .dout(n8371));
  jand g08308(.dina(n5363), .dinb(n2497), .dout(n8372));
  jor  g08309(.dina(n8372), .dinb(n8371), .dout(n8373));
  jor  g08310(.dina(n8373), .dinb(n8370), .dout(n8374));
  jor  g08311(.dina(n8374), .dinb(n8369), .dout(n8375));
  jxor g08312(.dina(n8375), .dinb(n72), .dout(n8376));
  jnot g08313(.din(n8376), .dout(n8377));
  jxor g08314(.dina(n8367), .dinb(n8366), .dout(n8378));
  jand g08315(.dina(n8378), .dinb(n8377), .dout(n8379));
  jor  g08316(.dina(n8379), .dinb(n8368), .dout(n8380));
  jxor g08317(.dina(n8091), .dinb(n8083), .dout(n8381));
  jand g08318(.dina(n8381), .dinb(n8380), .dout(n8382));
  jnot g08319(.din(n8382), .dout(n8383));
  jxor g08320(.dina(n8381), .dinb(n8380), .dout(n8384));
  jnot g08321(.din(n8384), .dout(n8385));
  jand g08322(.dina(n5693), .dinb(n5303), .dout(n8386));
  jand g08323(.dina(n6131), .dinb(n2067), .dout(n8387));
  jand g08324(.dina(n6209), .dinb(n1956), .dout(n8388));
  jand g08325(.dina(n5691), .dinb(n2128), .dout(n8389));
  jor  g08326(.dina(n8389), .dinb(n8388), .dout(n8390));
  jor  g08327(.dina(n8390), .dinb(n8387), .dout(n8391));
  jor  g08328(.dina(n8391), .dinb(n8386), .dout(n8392));
  jxor g08329(.dina(n8392), .dinb(n4247), .dout(n8393));
  jor  g08330(.dina(n8393), .dinb(n8385), .dout(n8394));
  jand g08331(.dina(n8394), .dinb(n8383), .dout(n8395));
  jnot g08332(.din(n8395), .dout(n8396));
  jxor g08333(.dina(n8107), .dinb(n8099), .dout(n8397));
  jand g08334(.dina(n8397), .dinb(n8396), .dout(n8398));
  jnot g08335(.din(n8398), .dout(n8399));
  jxor g08336(.dina(n8397), .dinb(n8396), .dout(n8400));
  jnot g08337(.din(n8400), .dout(n8401));
  jand g08338(.dina(n6340), .dinb(n4849), .dout(n8402));
  jand g08339(.dina(n6798), .dinb(n1560), .dout(n8403));
  jand g08340(.dina(n6556), .dinb(n1624), .dout(n8404));
  jand g08341(.dina(n6338), .dinb(n1776), .dout(n8405));
  jor  g08342(.dina(n8405), .dinb(n8404), .dout(n8406));
  jor  g08343(.dina(n8406), .dinb(n8403), .dout(n8407));
  jor  g08344(.dina(n8407), .dinb(n8402), .dout(n8408));
  jxor g08345(.dina(n8408), .dinb(n5064), .dout(n8409));
  jor  g08346(.dina(n8409), .dinb(n8401), .dout(n8410));
  jand g08347(.dina(n8410), .dinb(n8399), .dout(n8411));
  jnot g08348(.din(n8411), .dout(n8412));
  jxor g08349(.dina(n8179), .dinb(n8178), .dout(n8413));
  jand g08350(.dina(n8413), .dinb(n8412), .dout(n8414));
  jor  g08351(.dina(n8414), .dinb(n8180), .dout(n8415));
  jxor g08352(.dina(n8128), .dinb(n8120), .dout(n8416));
  jand g08353(.dina(n8416), .dinb(n8415), .dout(n8417));
  jnot g08354(.din(n8417), .dout(n8418));
  jxor g08355(.dina(n8416), .dinb(n8415), .dout(n8419));
  jnot g08356(.din(n8419), .dout(n8420));
  jand g08357(.dina(n6936), .dinb(n4026), .dout(n8421));
  jand g08358(.dina(n7613), .dinb(n1076), .dout(n8422));
  jand g08359(.dina(n7741), .dinb(n922), .dout(n8423));
  jand g08360(.dina(n6934), .dinb(n1213), .dout(n8424));
  jor  g08361(.dina(n8424), .dinb(n8423), .dout(n8425));
  jor  g08362(.dina(n8425), .dinb(n8422), .dout(n8426));
  jor  g08363(.dina(n8426), .dinb(n8421), .dout(n8427));
  jxor g08364(.dina(n8427), .dinb(n5292), .dout(n8428));
  jor  g08365(.dina(n8428), .dinb(n8420), .dout(n8429));
  jand g08366(.dina(n8429), .dinb(n8418), .dout(n8430));
  jnot g08367(.din(n8430), .dout(n8431));
  jxor g08368(.dina(n8144), .dinb(n8136), .dout(n8432));
  jand g08369(.dina(n8432), .dinb(n8431), .dout(n8433));
  jnot g08370(.din(n8433), .dout(n8434));
  jxor g08371(.dina(n8432), .dinb(n8431), .dout(n8435));
  jnot g08372(.din(n8435), .dout(n8436));
  jand g08373(.dina(n7890), .dinb(n4752), .dout(n8437));
  jand g08374(.dina(n8154), .dinb(n4451), .dout(n8438));
  jand g08375(.dina(n7888), .dinb(n4358), .dout(n8439));
  jor  g08376(.dina(n7887), .dinb(n7885), .dout(n8440));
  jnot g08377(.din(n8440), .dout(n8441));
  jand g08378(.dina(n8441), .dinb(n4598), .dout(n8442));
  jor  g08379(.dina(n8442), .dinb(n8439), .dout(n8443));
  jor  g08380(.dina(n8443), .dinb(n8438), .dout(n8444));
  jor  g08381(.dina(n8444), .dinb(n8437), .dout(n8445));
  jxor g08382(.dina(n8445), .dinb(n5833), .dout(n8446));
  jor  g08383(.dina(n8446), .dinb(n8436), .dout(n8447));
  jand g08384(.dina(n8447), .dinb(n8434), .dout(n8448));
  jand g08385(.dina(n7890), .dinb(n4636), .dout(n8449));
  jand g08386(.dina(n7888), .dinb(n4451), .dout(n8450));
  jand g08387(.dina(n8154), .dinb(n4598), .dout(n8451));
  jand g08388(.dina(n8441), .dinb(n4631), .dout(n8452));
  jor  g08389(.dina(n8452), .dinb(n8451), .dout(n8453));
  jor  g08390(.dina(n8453), .dinb(n8450), .dout(n8454));
  jor  g08391(.dina(n8454), .dinb(n8449), .dout(n8455));
  jxor g08392(.dina(n8455), .dinb(n5833), .dout(n8456));
  jor  g08393(.dina(n8456), .dinb(n8448), .dout(n8457));
  jxor g08394(.dina(n8456), .dinb(n8448), .dout(n8458));
  jxor g08395(.dina(n8148), .dinb(n8147), .dout(n8459));
  jand g08396(.dina(n8459), .dinb(n8458), .dout(n8460));
  jnot g08397(.din(n8460), .dout(n8461));
  jand g08398(.dina(n8461), .dinb(n8457), .dout(n8462));
  jnot g08399(.din(n8462), .dout(n8463));
  jxor g08400(.dina(n8162), .dinb(n8161), .dout(n8464));
  jand g08401(.dina(n8464), .dinb(n8463), .dout(n8465));
  jxor g08402(.dina(n8413), .dinb(n8412), .dout(n8466));
  jnot g08403(.din(n8466), .dout(n8467));
  jand g08404(.dina(n6936), .dinb(n4043), .dout(n8468));
  jand g08405(.dina(n7613), .dinb(n1213), .dout(n8469));
  jand g08406(.dina(n6934), .dinb(n1343), .dout(n8470));
  jand g08407(.dina(n7741), .dinb(n1076), .dout(n8471));
  jor  g08408(.dina(n8471), .dinb(n8470), .dout(n8472));
  jor  g08409(.dina(n8472), .dinb(n8469), .dout(n8473));
  jor  g08410(.dina(n8473), .dinb(n8468), .dout(n8474));
  jxor g08411(.dina(n8474), .dinb(n5292), .dout(n8475));
  jor  g08412(.dina(n8475), .dinb(n8467), .dout(n8476));
  jand g08413(.dina(n6247), .dinb(n5365), .dout(n8477));
  jand g08414(.dina(n5500), .dinb(n2411), .dout(n8478));
  jand g08415(.dina(n5363), .dinb(n2602), .dout(n8479));
  jand g08416(.dina(n5424), .dinb(n2497), .dout(n8480));
  jor  g08417(.dina(n8480), .dinb(n8479), .dout(n8481));
  jor  g08418(.dina(n8481), .dinb(n8478), .dout(n8482));
  jor  g08419(.dina(n8482), .dinb(n8477), .dout(n8483));
  jxor g08420(.dina(n8483), .dinb(n72), .dout(n8484));
  jnot g08421(.din(n8484), .dout(n8485));
  jxor g08422(.dina(n8362), .dinb(n8361), .dout(n8486));
  jand g08423(.dina(n8486), .dinb(n8485), .dout(n8487));
  jand g08424(.dina(n6050), .dinb(n5365), .dout(n8488));
  jand g08425(.dina(n5363), .dinb(n2695), .dout(n8489));
  jand g08426(.dina(n5424), .dinb(n2602), .dout(n8490));
  jand g08427(.dina(n5500), .dinb(n2497), .dout(n8491));
  jor  g08428(.dina(n8491), .dinb(n8490), .dout(n8492));
  jor  g08429(.dina(n8492), .dinb(n8489), .dout(n8493));
  jor  g08430(.dina(n8493), .dinb(n8488), .dout(n8494));
  jxor g08431(.dina(n8494), .dinb(n72), .dout(n8495));
  jnot g08432(.din(n8495), .dout(n8496));
  jxor g08433(.dina(n8357), .dinb(n8356), .dout(n8497));
  jand g08434(.dina(n8497), .dinb(n8496), .dout(n8498));
  jor  g08435(.dina(n6464), .dinb(n5366), .dout(n8499));
  jor  g08436(.dina(n5499), .dinb(n2601), .dout(n8500));
  jor  g08437(.dina(n5425), .dinb(n2694), .dout(n8501));
  jor  g08438(.dina(n5364), .dinb(n2731), .dout(n8502));
  jand g08439(.dina(n8502), .dinb(n8501), .dout(n8503));
  jand g08440(.dina(n8503), .dinb(n8500), .dout(n8504));
  jand g08441(.dina(n8504), .dinb(n8499), .dout(n8505));
  jxor g08442(.dina(n8505), .dinb(\a[23] ), .dout(n8506));
  jnot g08443(.din(n8506), .dout(n8507));
  jxor g08444(.dina(n8352), .dinb(n8351), .dout(n8508));
  jand g08445(.dina(n8508), .dinb(n8507), .dout(n8509));
  jand g08446(.dina(n6591), .dinb(n5365), .dout(n8510));
  jand g08447(.dina(n5500), .dinb(n2695), .dout(n8511));
  jand g08448(.dina(n5363), .dinb(n2808), .dout(n8512));
  jand g08449(.dina(n5424), .dinb(n2732), .dout(n8513));
  jor  g08450(.dina(n8513), .dinb(n8512), .dout(n8514));
  jor  g08451(.dina(n8514), .dinb(n8511), .dout(n8515));
  jor  g08452(.dina(n8515), .dinb(n8510), .dout(n8516));
  jxor g08453(.dina(n8516), .dinb(n72), .dout(n8517));
  jnot g08454(.din(n8517), .dout(n8518));
  jxor g08455(.dina(n8347), .dinb(n8346), .dout(n8519));
  jand g08456(.dina(n8519), .dinb(n8518), .dout(n8520));
  jand g08457(.dina(n6439), .dinb(n5365), .dout(n8521));
  jand g08458(.dina(n5424), .dinb(n2808), .dout(n8522));
  jand g08459(.dina(n5500), .dinb(n2732), .dout(n8523));
  jand g08460(.dina(n5363), .dinb(n2867), .dout(n8524));
  jor  g08461(.dina(n8524), .dinb(n8523), .dout(n8525));
  jor  g08462(.dina(n8525), .dinb(n8522), .dout(n8526));
  jor  g08463(.dina(n8526), .dinb(n8521), .dout(n8527));
  jxor g08464(.dina(n8527), .dinb(n72), .dout(n8528));
  jnot g08465(.din(n8528), .dout(n8529));
  jxor g08466(.dina(n8342), .dinb(n8341), .dout(n8530));
  jand g08467(.dina(n8530), .dinb(n8529), .dout(n8531));
  jand g08468(.dina(n6706), .dinb(n5365), .dout(n8532));
  jand g08469(.dina(n5500), .dinb(n2808), .dout(n8533));
  jand g08470(.dina(n5363), .dinb(n2954), .dout(n8534));
  jand g08471(.dina(n5424), .dinb(n2867), .dout(n8535));
  jor  g08472(.dina(n8535), .dinb(n8534), .dout(n8536));
  jor  g08473(.dina(n8536), .dinb(n8533), .dout(n8537));
  jor  g08474(.dina(n8537), .dinb(n8532), .dout(n8538));
  jxor g08475(.dina(n8538), .dinb(n72), .dout(n8539));
  jnot g08476(.din(n8539), .dout(n8540));
  jxor g08477(.dina(n8337), .dinb(n8336), .dout(n8541));
  jand g08478(.dina(n8541), .dinb(n8540), .dout(n8542));
  jor  g08479(.dina(n6976), .dinb(n5366), .dout(n8543));
  jor  g08480(.dina(n5499), .dinb(n2866), .dout(n8544));
  jor  g08481(.dina(n5425), .dinb(n2953), .dout(n8545));
  jor  g08482(.dina(n5364), .dinb(n2990), .dout(n8546));
  jand g08483(.dina(n8546), .dinb(n8545), .dout(n8547));
  jand g08484(.dina(n8547), .dinb(n8544), .dout(n8548));
  jand g08485(.dina(n8548), .dinb(n8543), .dout(n8549));
  jxor g08486(.dina(n8549), .dinb(\a[23] ), .dout(n8550));
  jnot g08487(.din(n8550), .dout(n8551));
  jxor g08488(.dina(n8334), .dinb(n8333), .dout(n8552));
  jand g08489(.dina(n8552), .dinb(n8551), .dout(n8553));
  jxor g08490(.dina(n8331), .dinb(n8330), .dout(n8554));
  jnot g08491(.din(n8554), .dout(n8555));
  jor  g08492(.dina(n6988), .dinb(n5366), .dout(n8556));
  jor  g08493(.dina(n5364), .dinb(n3085), .dout(n8557));
  jor  g08494(.dina(n5499), .dinb(n2953), .dout(n8558));
  jor  g08495(.dina(n5425), .dinb(n2990), .dout(n8559));
  jand g08496(.dina(n8559), .dinb(n8558), .dout(n8560));
  jand g08497(.dina(n8560), .dinb(n8557), .dout(n8561));
  jand g08498(.dina(n8561), .dinb(n8556), .dout(n8562));
  jxor g08499(.dina(n8562), .dinb(\a[23] ), .dout(n8563));
  jor  g08500(.dina(n8563), .dinb(n8555), .dout(n8564));
  jxor g08501(.dina(n8328), .dinb(n8327), .dout(n8565));
  jnot g08502(.din(n8565), .dout(n8566));
  jor  g08503(.dina(n6681), .dinb(n5366), .dout(n8567));
  jor  g08504(.dina(n5425), .dinb(n3085), .dout(n8568));
  jor  g08505(.dina(n5499), .dinb(n2990), .dout(n8569));
  jor  g08506(.dina(n5364), .dinb(n3182), .dout(n8570));
  jand g08507(.dina(n8570), .dinb(n8569), .dout(n8571));
  jand g08508(.dina(n8571), .dinb(n8568), .dout(n8572));
  jand g08509(.dina(n8572), .dinb(n8567), .dout(n8573));
  jxor g08510(.dina(n8573), .dinb(\a[23] ), .dout(n8574));
  jor  g08511(.dina(n8574), .dinb(n8566), .dout(n8575));
  jor  g08512(.dina(n7031), .dinb(n5366), .dout(n8576));
  jor  g08513(.dina(n5499), .dinb(n3085), .dout(n8577));
  jor  g08514(.dina(n5364), .dinb(n7962), .dout(n8578));
  jor  g08515(.dina(n5425), .dinb(n3182), .dout(n8579));
  jand g08516(.dina(n8579), .dinb(n8578), .dout(n8580));
  jand g08517(.dina(n8580), .dinb(n8577), .dout(n8581));
  jand g08518(.dina(n8581), .dinb(n8576), .dout(n8582));
  jxor g08519(.dina(n8582), .dinb(\a[23] ), .dout(n8583));
  jnot g08520(.din(n8583), .dout(n8584));
  jxor g08521(.dina(n8325), .dinb(n8324), .dout(n8585));
  jand g08522(.dina(n8585), .dinb(n8584), .dout(n8586));
  jor  g08523(.dina(n7076), .dinb(n5366), .dout(n8587));
  jor  g08524(.dina(n5425), .dinb(n7962), .dout(n8588));
  jor  g08525(.dina(n5499), .dinb(n3182), .dout(n8589));
  jor  g08526(.dina(n5364), .dinb(n3684), .dout(n8590));
  jand g08527(.dina(n8590), .dinb(n8589), .dout(n8591));
  jand g08528(.dina(n8591), .dinb(n8588), .dout(n8592));
  jand g08529(.dina(n8592), .dinb(n8587), .dout(n8593));
  jxor g08530(.dina(n8593), .dinb(\a[23] ), .dout(n8594));
  jnot g08531(.din(n8594), .dout(n8595));
  jxor g08532(.dina(n8322), .dinb(n8321), .dout(n8596));
  jand g08533(.dina(n8596), .dinb(n8595), .dout(n8597));
  jor  g08534(.dina(n7131), .dinb(n5366), .dout(n8598));
  jor  g08535(.dina(n5499), .dinb(n7962), .dout(n8599));
  jor  g08536(.dina(n5364), .dinb(n3414), .dout(n8600));
  jor  g08537(.dina(n5425), .dinb(n3684), .dout(n8601));
  jand g08538(.dina(n8601), .dinb(n8600), .dout(n8602));
  jand g08539(.dina(n8602), .dinb(n8599), .dout(n8603));
  jand g08540(.dina(n8603), .dinb(n8598), .dout(n8604));
  jxor g08541(.dina(n8604), .dinb(\a[23] ), .dout(n8605));
  jnot g08542(.din(n8605), .dout(n8606));
  jor  g08543(.dina(n8302), .dinb(n68), .dout(n8607));
  jxor g08544(.dina(n8607), .dinb(n8310), .dout(n8608));
  jand g08545(.dina(n8608), .dinb(n8606), .dout(n8609));
  jor  g08546(.dina(n7177), .dinb(n5366), .dout(n8610));
  jor  g08547(.dina(n5364), .dinb(n3516), .dout(n8611));
  jor  g08548(.dina(n5499), .dinb(n3684), .dout(n8612));
  jor  g08549(.dina(n5425), .dinb(n3414), .dout(n8613));
  jand g08550(.dina(n8613), .dinb(n8612), .dout(n8614));
  jand g08551(.dina(n8614), .dinb(n8611), .dout(n8615));
  jand g08552(.dina(n8615), .dinb(n8610), .dout(n8616));
  jxor g08553(.dina(n8616), .dinb(\a[23] ), .dout(n8617));
  jnot g08554(.din(n8617), .dout(n8618));
  jand g08555(.dina(n8299), .dinb(\a[26] ), .dout(n8619));
  jxor g08556(.dina(n8619), .dinb(n8297), .dout(n8620));
  jand g08557(.dina(n8620), .dinb(n8618), .dout(n8621));
  jand g08558(.dina(n8004), .dinb(n5365), .dout(n8622));
  jand g08559(.dina(n5424), .dinb(n7411), .dout(n8623));
  jand g08560(.dina(n5500), .dinb(n7405), .dout(n8624));
  jor  g08561(.dina(n8624), .dinb(n8623), .dout(n8625));
  jor  g08562(.dina(n8625), .dinb(n8622), .dout(n8626));
  jnot g08563(.din(n8626), .dout(n8627));
  jand g08564(.dina(n5358), .dinb(n7411), .dout(n8628));
  jnot g08565(.din(n8628), .dout(n8629));
  jand g08566(.dina(n8629), .dinb(\a[23] ), .dout(n8630));
  jand g08567(.dina(n8630), .dinb(n8627), .dout(n8631));
  jand g08568(.dina(n7407), .dinb(n5365), .dout(n8632));
  jand g08569(.dina(n5500), .dinb(n7326), .dout(n8633));
  jand g08570(.dina(n5363), .dinb(n7411), .dout(n8634));
  jand g08571(.dina(n5424), .dinb(n7405), .dout(n8635));
  jor  g08572(.dina(n8635), .dinb(n8634), .dout(n8636));
  jor  g08573(.dina(n8636), .dinb(n8633), .dout(n8637));
  jor  g08574(.dina(n8637), .dinb(n8632), .dout(n8638));
  jnot g08575(.din(n8638), .dout(n8639));
  jand g08576(.dina(n8639), .dinb(n8631), .dout(n8640));
  jand g08577(.dina(n8640), .dinb(n8299), .dout(n8641));
  jor  g08578(.dina(n7466), .dinb(n5366), .dout(n8642));
  jor  g08579(.dina(n5425), .dinb(n3516), .dout(n8643));
  jor  g08580(.dina(n5499), .dinb(n3414), .dout(n8644));
  jor  g08581(.dina(n5364), .dinb(n3677), .dout(n8645));
  jand g08582(.dina(n8645), .dinb(n8644), .dout(n8646));
  jand g08583(.dina(n8646), .dinb(n8643), .dout(n8647));
  jand g08584(.dina(n8647), .dinb(n8642), .dout(n8648));
  jxor g08585(.dina(n8648), .dinb(\a[23] ), .dout(n8649));
  jnot g08586(.din(n8649), .dout(n8650));
  jxor g08587(.dina(n8640), .dinb(n8299), .dout(n8651));
  jand g08588(.dina(n8651), .dinb(n8650), .dout(n8652));
  jor  g08589(.dina(n8652), .dinb(n8641), .dout(n8653));
  jxor g08590(.dina(n8620), .dinb(n8618), .dout(n8654));
  jand g08591(.dina(n8654), .dinb(n8653), .dout(n8655));
  jor  g08592(.dina(n8655), .dinb(n8621), .dout(n8656));
  jxor g08593(.dina(n8608), .dinb(n8606), .dout(n8657));
  jand g08594(.dina(n8657), .dinb(n8656), .dout(n8658));
  jor  g08595(.dina(n8658), .dinb(n8609), .dout(n8659));
  jxor g08596(.dina(n8596), .dinb(n8595), .dout(n8660));
  jand g08597(.dina(n8660), .dinb(n8659), .dout(n8661));
  jor  g08598(.dina(n8661), .dinb(n8597), .dout(n8662));
  jxor g08599(.dina(n8585), .dinb(n8584), .dout(n8663));
  jand g08600(.dina(n8663), .dinb(n8662), .dout(n8664));
  jor  g08601(.dina(n8664), .dinb(n8586), .dout(n8665));
  jxor g08602(.dina(n8574), .dinb(n8566), .dout(n8666));
  jand g08603(.dina(n8666), .dinb(n8665), .dout(n8667));
  jnot g08604(.din(n8667), .dout(n8668));
  jand g08605(.dina(n8668), .dinb(n8575), .dout(n8669));
  jnot g08606(.din(n8669), .dout(n8670));
  jxor g08607(.dina(n8563), .dinb(n8555), .dout(n8671));
  jand g08608(.dina(n8671), .dinb(n8670), .dout(n8672));
  jnot g08609(.din(n8672), .dout(n8673));
  jand g08610(.dina(n8673), .dinb(n8564), .dout(n8674));
  jnot g08611(.din(n8674), .dout(n8675));
  jxor g08612(.dina(n8552), .dinb(n8551), .dout(n8676));
  jand g08613(.dina(n8676), .dinb(n8675), .dout(n8677));
  jor  g08614(.dina(n8677), .dinb(n8553), .dout(n8678));
  jxor g08615(.dina(n8541), .dinb(n8540), .dout(n8679));
  jand g08616(.dina(n8679), .dinb(n8678), .dout(n8680));
  jor  g08617(.dina(n8680), .dinb(n8542), .dout(n8681));
  jxor g08618(.dina(n8530), .dinb(n8529), .dout(n8682));
  jand g08619(.dina(n8682), .dinb(n8681), .dout(n8683));
  jor  g08620(.dina(n8683), .dinb(n8531), .dout(n8684));
  jxor g08621(.dina(n8519), .dinb(n8518), .dout(n8685));
  jand g08622(.dina(n8685), .dinb(n8684), .dout(n8686));
  jor  g08623(.dina(n8686), .dinb(n8520), .dout(n8687));
  jxor g08624(.dina(n8508), .dinb(n8507), .dout(n8688));
  jand g08625(.dina(n8688), .dinb(n8687), .dout(n8689));
  jor  g08626(.dina(n8689), .dinb(n8509), .dout(n8690));
  jxor g08627(.dina(n8497), .dinb(n8496), .dout(n8691));
  jand g08628(.dina(n8691), .dinb(n8690), .dout(n8692));
  jor  g08629(.dina(n8692), .dinb(n8498), .dout(n8693));
  jxor g08630(.dina(n8486), .dinb(n8485), .dout(n8694));
  jand g08631(.dina(n8694), .dinb(n8693), .dout(n8695));
  jor  g08632(.dina(n8695), .dinb(n8487), .dout(n8696));
  jxor g08633(.dina(n8378), .dinb(n8377), .dout(n8697));
  jand g08634(.dina(n8697), .dinb(n8696), .dout(n8698));
  jand g08635(.dina(n5693), .dinb(n5624), .dout(n8699));
  jand g08636(.dina(n5691), .dinb(n2237), .dout(n8700));
  jand g08637(.dina(n6131), .dinb(n2128), .dout(n8701));
  jand g08638(.dina(n6209), .dinb(n2067), .dout(n8702));
  jor  g08639(.dina(n8702), .dinb(n8701), .dout(n8703));
  jor  g08640(.dina(n8703), .dinb(n8700), .dout(n8704));
  jor  g08641(.dina(n8704), .dinb(n8699), .dout(n8705));
  jxor g08642(.dina(n8705), .dinb(n4247), .dout(n8706));
  jnot g08643(.din(n8706), .dout(n8707));
  jxor g08644(.dina(n8697), .dinb(n8696), .dout(n8708));
  jand g08645(.dina(n8708), .dinb(n8707), .dout(n8709));
  jor  g08646(.dina(n8709), .dinb(n8698), .dout(n8710));
  jxor g08647(.dina(n8393), .dinb(n8385), .dout(n8711));
  jand g08648(.dina(n8711), .dinb(n8710), .dout(n8712));
  jnot g08649(.din(n8712), .dout(n8713));
  jxor g08650(.dina(n8711), .dinb(n8710), .dout(n8714));
  jnot g08651(.din(n8714), .dout(n8715));
  jand g08652(.dina(n6340), .dinb(n5075), .dout(n8716));
  jand g08653(.dina(n6798), .dinb(n1624), .dout(n8717));
  jand g08654(.dina(n6556), .dinb(n1776), .dout(n8718));
  jand g08655(.dina(n6338), .dinb(n1862), .dout(n8719));
  jor  g08656(.dina(n8719), .dinb(n8718), .dout(n8720));
  jor  g08657(.dina(n8720), .dinb(n8717), .dout(n8721));
  jor  g08658(.dina(n8721), .dinb(n8716), .dout(n8722));
  jxor g08659(.dina(n8722), .dinb(n5064), .dout(n8723));
  jor  g08660(.dina(n8723), .dinb(n8715), .dout(n8724));
  jand g08661(.dina(n8724), .dinb(n8713), .dout(n8725));
  jnot g08662(.din(n8725), .dout(n8726));
  jxor g08663(.dina(n8409), .dinb(n8401), .dout(n8727));
  jand g08664(.dina(n8727), .dinb(n8726), .dout(n8728));
  jnot g08665(.din(n8728), .dout(n8729));
  jxor g08666(.dina(n8727), .dinb(n8726), .dout(n8730));
  jnot g08667(.din(n8730), .dout(n8731));
  jand g08668(.dina(n6936), .dinb(n4772), .dout(n8732));
  jand g08669(.dina(n7741), .dinb(n1213), .dout(n8733));
  jand g08670(.dina(n7613), .dinb(n1343), .dout(n8734));
  jand g08671(.dina(n6934), .dinb(n1445), .dout(n8735));
  jor  g08672(.dina(n8735), .dinb(n8734), .dout(n8736));
  jor  g08673(.dina(n8736), .dinb(n8733), .dout(n8737));
  jor  g08674(.dina(n8737), .dinb(n8732), .dout(n8738));
  jxor g08675(.dina(n8738), .dinb(n5292), .dout(n8739));
  jor  g08676(.dina(n8739), .dinb(n8731), .dout(n8740));
  jand g08677(.dina(n8740), .dinb(n8729), .dout(n8741));
  jnot g08678(.din(n8741), .dout(n8742));
  jxor g08679(.dina(n8475), .dinb(n8467), .dout(n8743));
  jand g08680(.dina(n8743), .dinb(n8742), .dout(n8744));
  jnot g08681(.din(n8744), .dout(n8745));
  jand g08682(.dina(n8745), .dinb(n8476), .dout(n8746));
  jnot g08683(.din(n8746), .dout(n8747));
  jxor g08684(.dina(n8428), .dinb(n8420), .dout(n8748));
  jand g08685(.dina(n8748), .dinb(n8747), .dout(n8749));
  jnot g08686(.din(n8749), .dout(n8750));
  jxor g08687(.dina(n8748), .dinb(n8747), .dout(n8751));
  jnot g08688(.din(n8751), .dout(n8752));
  jand g08689(.dina(n7890), .dinb(n4446), .dout(n8753));
  jand g08690(.dina(n8441), .dinb(n4451), .dout(n8754));
  jand g08691(.dina(n8154), .dinb(n4358), .dout(n8755));
  jand g08692(.dina(n7888), .dinb(n3853), .dout(n8756));
  jor  g08693(.dina(n8756), .dinb(n8755), .dout(n8757));
  jor  g08694(.dina(n8757), .dinb(n8754), .dout(n8758));
  jor  g08695(.dina(n8758), .dinb(n8753), .dout(n8759));
  jxor g08696(.dina(n8759), .dinb(n5833), .dout(n8760));
  jor  g08697(.dina(n8760), .dinb(n8752), .dout(n8761));
  jand g08698(.dina(n8761), .dinb(n8750), .dout(n8762));
  jxor g08699(.dina(\a[7] ), .dinb(\a[6] ), .dout(n8763));
  jnot g08700(.din(n8763), .dout(n8764));
  jxor g08701(.dina(\a[6] ), .dinb(\a[5] ), .dout(n8765));
  jnot g08702(.din(n8765), .dout(n8766));
  jand g08703(.dina(n8766), .dinb(n8764), .dout(n8767));
  jxor g08704(.dina(\a[8] ), .dinb(\a[7] ), .dout(n8768));
  jand g08705(.dina(n8768), .dinb(n8767), .dout(n8769));
  jnot g08706(.din(n8769), .dout(n8770));
  jand g08707(.dina(n8768), .dinb(n8765), .dout(n8771));
  jnot g08708(.din(n8771), .dout(n8772));
  jor  g08709(.dina(n8772), .dinb(n4728), .dout(n8773));
  jand g08710(.dina(n8773), .dinb(n8770), .dout(n8774));
  jor  g08711(.dina(n8774), .dinb(n4630), .dout(n8775));
  jxor g08712(.dina(n8775), .dinb(\a[8] ), .dout(n8776));
  jor  g08713(.dina(n8776), .dinb(n8762), .dout(n8777));
  jxor g08714(.dina(n8776), .dinb(n8762), .dout(n8778));
  jxor g08715(.dina(n8446), .dinb(n8436), .dout(n8779));
  jand g08716(.dina(n8779), .dinb(n8778), .dout(n8780));
  jnot g08717(.din(n8780), .dout(n8781));
  jand g08718(.dina(n8781), .dinb(n8777), .dout(n8782));
  jnot g08719(.din(n8782), .dout(n8783));
  jxor g08720(.dina(n8459), .dinb(n8458), .dout(n8784));
  jand g08721(.dina(n8784), .dinb(n8783), .dout(n8785));
  jxor g08722(.dina(n8784), .dinb(n8783), .dout(n8786));
  jxor g08723(.dina(n8694), .dinb(n8693), .dout(n8787));
  jnot g08724(.din(n8787), .dout(n8788));
  jand g08725(.dina(n5693), .dinb(n5607), .dout(n8789));
  jand g08726(.dina(n6131), .dinb(n2237), .dout(n8790));
  jand g08727(.dina(n5691), .dinb(n2343), .dout(n8791));
  jand g08728(.dina(n6209), .dinb(n2128), .dout(n8792));
  jor  g08729(.dina(n8792), .dinb(n8791), .dout(n8793));
  jor  g08730(.dina(n8793), .dinb(n8790), .dout(n8794));
  jor  g08731(.dina(n8794), .dinb(n8789), .dout(n8795));
  jxor g08732(.dina(n8795), .dinb(n4247), .dout(n8796));
  jor  g08733(.dina(n8796), .dinb(n8788), .dout(n8797));
  jxor g08734(.dina(n8691), .dinb(n8690), .dout(n8798));
  jnot g08735(.din(n8798), .dout(n8799));
  jand g08736(.dina(n5844), .dinb(n5693), .dout(n8800));
  jand g08737(.dina(n5691), .dinb(n2411), .dout(n8801));
  jand g08738(.dina(n6209), .dinb(n2237), .dout(n8802));
  jand g08739(.dina(n6131), .dinb(n2343), .dout(n8803));
  jor  g08740(.dina(n8803), .dinb(n8802), .dout(n8804));
  jor  g08741(.dina(n8804), .dinb(n8801), .dout(n8805));
  jor  g08742(.dina(n8805), .dinb(n8800), .dout(n8806));
  jxor g08743(.dina(n8806), .dinb(n4247), .dout(n8807));
  jor  g08744(.dina(n8807), .dinb(n8799), .dout(n8808));
  jxor g08745(.dina(n8688), .dinb(n8687), .dout(n8809));
  jnot g08746(.din(n8809), .dout(n8810));
  jand g08747(.dina(n5861), .dinb(n5693), .dout(n8811));
  jand g08748(.dina(n6131), .dinb(n2411), .dout(n8812));
  jand g08749(.dina(n6209), .dinb(n2343), .dout(n8813));
  jand g08750(.dina(n5691), .dinb(n2497), .dout(n8814));
  jor  g08751(.dina(n8814), .dinb(n8813), .dout(n8815));
  jor  g08752(.dina(n8815), .dinb(n8812), .dout(n8816));
  jor  g08753(.dina(n8816), .dinb(n8811), .dout(n8817));
  jxor g08754(.dina(n8817), .dinb(n4247), .dout(n8818));
  jor  g08755(.dina(n8818), .dinb(n8810), .dout(n8819));
  jxor g08756(.dina(n8685), .dinb(n8684), .dout(n8820));
  jnot g08757(.din(n8820), .dout(n8821));
  jand g08758(.dina(n6247), .dinb(n5693), .dout(n8822));
  jand g08759(.dina(n6209), .dinb(n2411), .dout(n8823));
  jand g08760(.dina(n5691), .dinb(n2602), .dout(n8824));
  jand g08761(.dina(n6131), .dinb(n2497), .dout(n8825));
  jor  g08762(.dina(n8825), .dinb(n8824), .dout(n8826));
  jor  g08763(.dina(n8826), .dinb(n8823), .dout(n8827));
  jor  g08764(.dina(n8827), .dinb(n8822), .dout(n8828));
  jxor g08765(.dina(n8828), .dinb(n4247), .dout(n8829));
  jor  g08766(.dina(n8829), .dinb(n8821), .dout(n8830));
  jxor g08767(.dina(n8682), .dinb(n8681), .dout(n8831));
  jnot g08768(.din(n8831), .dout(n8832));
  jand g08769(.dina(n6050), .dinb(n5693), .dout(n8833));
  jand g08770(.dina(n6131), .dinb(n2602), .dout(n8834));
  jand g08771(.dina(n5691), .dinb(n2695), .dout(n8835));
  jand g08772(.dina(n6209), .dinb(n2497), .dout(n8836));
  jor  g08773(.dina(n8836), .dinb(n8835), .dout(n8837));
  jor  g08774(.dina(n8837), .dinb(n8834), .dout(n8838));
  jor  g08775(.dina(n8838), .dinb(n8833), .dout(n8839));
  jxor g08776(.dina(n8839), .dinb(n4247), .dout(n8840));
  jor  g08777(.dina(n8840), .dinb(n8832), .dout(n8841));
  jxor g08778(.dina(n8679), .dinb(n8678), .dout(n8842));
  jnot g08779(.din(n8842), .dout(n8843));
  jor  g08780(.dina(n6464), .dinb(n5694), .dout(n8844));
  jor  g08781(.dina(n6208), .dinb(n2601), .dout(n8845));
  jor  g08782(.dina(n6132), .dinb(n2694), .dout(n8846));
  jor  g08783(.dina(n5692), .dinb(n2731), .dout(n8847));
  jand g08784(.dina(n8847), .dinb(n8846), .dout(n8848));
  jand g08785(.dina(n8848), .dinb(n8845), .dout(n8849));
  jand g08786(.dina(n8849), .dinb(n8844), .dout(n8850));
  jxor g08787(.dina(n8850), .dinb(\a[20] ), .dout(n8851));
  jor  g08788(.dina(n8851), .dinb(n8843), .dout(n8852));
  jxor g08789(.dina(n8676), .dinb(n8675), .dout(n8853));
  jnot g08790(.din(n8853), .dout(n8854));
  jand g08791(.dina(n6591), .dinb(n5693), .dout(n8855));
  jand g08792(.dina(n6209), .dinb(n2695), .dout(n8856));
  jand g08793(.dina(n5691), .dinb(n2808), .dout(n8857));
  jand g08794(.dina(n6131), .dinb(n2732), .dout(n8858));
  jor  g08795(.dina(n8858), .dinb(n8857), .dout(n8859));
  jor  g08796(.dina(n8859), .dinb(n8856), .dout(n8860));
  jor  g08797(.dina(n8860), .dinb(n8855), .dout(n8861));
  jxor g08798(.dina(n8861), .dinb(n4247), .dout(n8862));
  jor  g08799(.dina(n8862), .dinb(n8854), .dout(n8863));
  jand g08800(.dina(n6439), .dinb(n5693), .dout(n8864));
  jand g08801(.dina(n6131), .dinb(n2808), .dout(n8865));
  jand g08802(.dina(n6209), .dinb(n2732), .dout(n8866));
  jand g08803(.dina(n5691), .dinb(n2867), .dout(n8867));
  jor  g08804(.dina(n8867), .dinb(n8866), .dout(n8868));
  jor  g08805(.dina(n8868), .dinb(n8865), .dout(n8869));
  jor  g08806(.dina(n8869), .dinb(n8864), .dout(n8870));
  jxor g08807(.dina(n8870), .dinb(n4247), .dout(n8871));
  jnot g08808(.din(n8871), .dout(n8872));
  jxor g08809(.dina(n8671), .dinb(n8670), .dout(n8873));
  jand g08810(.dina(n8873), .dinb(n8872), .dout(n8874));
  jand g08811(.dina(n6706), .dinb(n5693), .dout(n8875));
  jand g08812(.dina(n6209), .dinb(n2808), .dout(n8876));
  jand g08813(.dina(n5691), .dinb(n2954), .dout(n8877));
  jand g08814(.dina(n6131), .dinb(n2867), .dout(n8878));
  jor  g08815(.dina(n8878), .dinb(n8877), .dout(n8879));
  jor  g08816(.dina(n8879), .dinb(n8876), .dout(n8880));
  jor  g08817(.dina(n8880), .dinb(n8875), .dout(n8881));
  jxor g08818(.dina(n8881), .dinb(n4247), .dout(n8882));
  jnot g08819(.din(n8882), .dout(n8883));
  jxor g08820(.dina(n8666), .dinb(n8665), .dout(n8884));
  jand g08821(.dina(n8884), .dinb(n8883), .dout(n8885));
  jxor g08822(.dina(n8663), .dinb(n8662), .dout(n8886));
  jnot g08823(.din(n8886), .dout(n8887));
  jor  g08824(.dina(n6976), .dinb(n5694), .dout(n8888));
  jor  g08825(.dina(n6132), .dinb(n2953), .dout(n8889));
  jor  g08826(.dina(n5692), .dinb(n2990), .dout(n8890));
  jor  g08827(.dina(n6208), .dinb(n2866), .dout(n8891));
  jand g08828(.dina(n8891), .dinb(n8890), .dout(n8892));
  jand g08829(.dina(n8892), .dinb(n8889), .dout(n8893));
  jand g08830(.dina(n8893), .dinb(n8888), .dout(n8894));
  jxor g08831(.dina(n8894), .dinb(\a[20] ), .dout(n8895));
  jor  g08832(.dina(n8895), .dinb(n8887), .dout(n8896));
  jxor g08833(.dina(n8660), .dinb(n8659), .dout(n8897));
  jnot g08834(.din(n8897), .dout(n8898));
  jor  g08835(.dina(n6988), .dinb(n5694), .dout(n8899));
  jor  g08836(.dina(n5692), .dinb(n3085), .dout(n8900));
  jor  g08837(.dina(n6208), .dinb(n2953), .dout(n8901));
  jor  g08838(.dina(n6132), .dinb(n2990), .dout(n8902));
  jand g08839(.dina(n8902), .dinb(n8901), .dout(n8903));
  jand g08840(.dina(n8903), .dinb(n8900), .dout(n8904));
  jand g08841(.dina(n8904), .dinb(n8899), .dout(n8905));
  jxor g08842(.dina(n8905), .dinb(\a[20] ), .dout(n8906));
  jor  g08843(.dina(n8906), .dinb(n8898), .dout(n8907));
  jxor g08844(.dina(n8657), .dinb(n8656), .dout(n8908));
  jnot g08845(.din(n8908), .dout(n8909));
  jor  g08846(.dina(n6681), .dinb(n5694), .dout(n8910));
  jor  g08847(.dina(n6132), .dinb(n3085), .dout(n8911));
  jor  g08848(.dina(n6208), .dinb(n2990), .dout(n8912));
  jor  g08849(.dina(n5692), .dinb(n3182), .dout(n8913));
  jand g08850(.dina(n8913), .dinb(n8912), .dout(n8914));
  jand g08851(.dina(n8914), .dinb(n8911), .dout(n8915));
  jand g08852(.dina(n8915), .dinb(n8910), .dout(n8916));
  jxor g08853(.dina(n8916), .dinb(\a[20] ), .dout(n8917));
  jor  g08854(.dina(n8917), .dinb(n8909), .dout(n8918));
  jor  g08855(.dina(n7031), .dinb(n5694), .dout(n8919));
  jor  g08856(.dina(n6208), .dinb(n3085), .dout(n8920));
  jor  g08857(.dina(n5692), .dinb(n7962), .dout(n8921));
  jor  g08858(.dina(n6132), .dinb(n3182), .dout(n8922));
  jand g08859(.dina(n8922), .dinb(n8921), .dout(n8923));
  jand g08860(.dina(n8923), .dinb(n8920), .dout(n8924));
  jand g08861(.dina(n8924), .dinb(n8919), .dout(n8925));
  jxor g08862(.dina(n8925), .dinb(\a[20] ), .dout(n8926));
  jnot g08863(.din(n8926), .dout(n8927));
  jxor g08864(.dina(n8654), .dinb(n8653), .dout(n8928));
  jand g08865(.dina(n8928), .dinb(n8927), .dout(n8929));
  jor  g08866(.dina(n7076), .dinb(n5694), .dout(n8930));
  jor  g08867(.dina(n6132), .dinb(n7962), .dout(n8931));
  jor  g08868(.dina(n6208), .dinb(n3182), .dout(n8932));
  jor  g08869(.dina(n5692), .dinb(n3684), .dout(n8933));
  jand g08870(.dina(n8933), .dinb(n8932), .dout(n8934));
  jand g08871(.dina(n8934), .dinb(n8931), .dout(n8935));
  jand g08872(.dina(n8935), .dinb(n8930), .dout(n8936));
  jxor g08873(.dina(n8936), .dinb(\a[20] ), .dout(n8937));
  jnot g08874(.din(n8937), .dout(n8938));
  jxor g08875(.dina(n8651), .dinb(n8650), .dout(n8939));
  jand g08876(.dina(n8939), .dinb(n8938), .dout(n8940));
  jor  g08877(.dina(n7131), .dinb(n5694), .dout(n8941));
  jor  g08878(.dina(n6208), .dinb(n7962), .dout(n8942));
  jor  g08879(.dina(n5692), .dinb(n3414), .dout(n8943));
  jor  g08880(.dina(n6132), .dinb(n3684), .dout(n8944));
  jand g08881(.dina(n8944), .dinb(n8943), .dout(n8945));
  jand g08882(.dina(n8945), .dinb(n8942), .dout(n8946));
  jand g08883(.dina(n8946), .dinb(n8941), .dout(n8947));
  jxor g08884(.dina(n8947), .dinb(\a[20] ), .dout(n8948));
  jnot g08885(.din(n8948), .dout(n8949));
  jor  g08886(.dina(n8631), .dinb(n72), .dout(n8950));
  jxor g08887(.dina(n8950), .dinb(n8639), .dout(n8951));
  jand g08888(.dina(n8951), .dinb(n8949), .dout(n8952));
  jor  g08889(.dina(n7177), .dinb(n5694), .dout(n8953));
  jor  g08890(.dina(n5692), .dinb(n3516), .dout(n8954));
  jor  g08891(.dina(n6208), .dinb(n3684), .dout(n8955));
  jor  g08892(.dina(n6132), .dinb(n3414), .dout(n8956));
  jand g08893(.dina(n8956), .dinb(n8955), .dout(n8957));
  jand g08894(.dina(n8957), .dinb(n8954), .dout(n8958));
  jand g08895(.dina(n8958), .dinb(n8953), .dout(n8959));
  jxor g08896(.dina(n8959), .dinb(\a[20] ), .dout(n8960));
  jnot g08897(.din(n8960), .dout(n8961));
  jand g08898(.dina(n8628), .dinb(\a[23] ), .dout(n8962));
  jxor g08899(.dina(n8962), .dinb(n8626), .dout(n8963));
  jand g08900(.dina(n8963), .dinb(n8961), .dout(n8964));
  jand g08901(.dina(n8004), .dinb(n5693), .dout(n8965));
  jand g08902(.dina(n6131), .dinb(n7411), .dout(n8966));
  jand g08903(.dina(n6209), .dinb(n7405), .dout(n8967));
  jor  g08904(.dina(n8967), .dinb(n8966), .dout(n8968));
  jor  g08905(.dina(n8968), .dinb(n8965), .dout(n8969));
  jnot g08906(.din(n8969), .dout(n8970));
  jand g08907(.dina(n5687), .dinb(n7411), .dout(n8971));
  jnot g08908(.din(n8971), .dout(n8972));
  jand g08909(.dina(n8972), .dinb(\a[20] ), .dout(n8973));
  jand g08910(.dina(n8973), .dinb(n8970), .dout(n8974));
  jand g08911(.dina(n7407), .dinb(n5693), .dout(n8975));
  jand g08912(.dina(n6209), .dinb(n7326), .dout(n8976));
  jand g08913(.dina(n5691), .dinb(n7411), .dout(n8977));
  jand g08914(.dina(n6131), .dinb(n7405), .dout(n8978));
  jor  g08915(.dina(n8978), .dinb(n8977), .dout(n8979));
  jor  g08916(.dina(n8979), .dinb(n8976), .dout(n8980));
  jor  g08917(.dina(n8980), .dinb(n8975), .dout(n8981));
  jnot g08918(.din(n8981), .dout(n8982));
  jand g08919(.dina(n8982), .dinb(n8974), .dout(n8983));
  jand g08920(.dina(n8983), .dinb(n8628), .dout(n8984));
  jor  g08921(.dina(n7466), .dinb(n5694), .dout(n8985));
  jor  g08922(.dina(n6132), .dinb(n3516), .dout(n8986));
  jor  g08923(.dina(n6208), .dinb(n3414), .dout(n8987));
  jor  g08924(.dina(n5692), .dinb(n3677), .dout(n8988));
  jand g08925(.dina(n8988), .dinb(n8987), .dout(n8989));
  jand g08926(.dina(n8989), .dinb(n8986), .dout(n8990));
  jand g08927(.dina(n8990), .dinb(n8985), .dout(n8991));
  jxor g08928(.dina(n8991), .dinb(\a[20] ), .dout(n8992));
  jnot g08929(.din(n8992), .dout(n8993));
  jxor g08930(.dina(n8983), .dinb(n8628), .dout(n8994));
  jand g08931(.dina(n8994), .dinb(n8993), .dout(n8995));
  jor  g08932(.dina(n8995), .dinb(n8984), .dout(n8996));
  jxor g08933(.dina(n8963), .dinb(n8961), .dout(n8997));
  jand g08934(.dina(n8997), .dinb(n8996), .dout(n8998));
  jor  g08935(.dina(n8998), .dinb(n8964), .dout(n8999));
  jxor g08936(.dina(n8951), .dinb(n8949), .dout(n9000));
  jand g08937(.dina(n9000), .dinb(n8999), .dout(n9001));
  jor  g08938(.dina(n9001), .dinb(n8952), .dout(n9002));
  jxor g08939(.dina(n8939), .dinb(n8938), .dout(n9003));
  jand g08940(.dina(n9003), .dinb(n9002), .dout(n9004));
  jor  g08941(.dina(n9004), .dinb(n8940), .dout(n9005));
  jxor g08942(.dina(n8928), .dinb(n8927), .dout(n9006));
  jand g08943(.dina(n9006), .dinb(n9005), .dout(n9007));
  jor  g08944(.dina(n9007), .dinb(n8929), .dout(n9008));
  jxor g08945(.dina(n8917), .dinb(n8909), .dout(n9009));
  jand g08946(.dina(n9009), .dinb(n9008), .dout(n9010));
  jnot g08947(.din(n9010), .dout(n9011));
  jand g08948(.dina(n9011), .dinb(n8918), .dout(n9012));
  jnot g08949(.din(n9012), .dout(n9013));
  jxor g08950(.dina(n8906), .dinb(n8898), .dout(n9014));
  jand g08951(.dina(n9014), .dinb(n9013), .dout(n9015));
  jnot g08952(.din(n9015), .dout(n9016));
  jand g08953(.dina(n9016), .dinb(n8907), .dout(n9017));
  jnot g08954(.din(n9017), .dout(n9018));
  jxor g08955(.dina(n8895), .dinb(n8887), .dout(n9019));
  jand g08956(.dina(n9019), .dinb(n9018), .dout(n9020));
  jnot g08957(.din(n9020), .dout(n9021));
  jand g08958(.dina(n9021), .dinb(n8896), .dout(n9022));
  jnot g08959(.din(n9022), .dout(n9023));
  jxor g08960(.dina(n8884), .dinb(n8883), .dout(n9024));
  jand g08961(.dina(n9024), .dinb(n9023), .dout(n9025));
  jor  g08962(.dina(n9025), .dinb(n8885), .dout(n9026));
  jxor g08963(.dina(n8873), .dinb(n8872), .dout(n9027));
  jand g08964(.dina(n9027), .dinb(n9026), .dout(n9028));
  jor  g08965(.dina(n9028), .dinb(n8874), .dout(n9029));
  jxor g08966(.dina(n8862), .dinb(n8854), .dout(n9030));
  jand g08967(.dina(n9030), .dinb(n9029), .dout(n9031));
  jnot g08968(.din(n9031), .dout(n9032));
  jand g08969(.dina(n9032), .dinb(n8863), .dout(n9033));
  jnot g08970(.din(n9033), .dout(n9034));
  jxor g08971(.dina(n8851), .dinb(n8843), .dout(n9035));
  jand g08972(.dina(n9035), .dinb(n9034), .dout(n9036));
  jnot g08973(.din(n9036), .dout(n9037));
  jand g08974(.dina(n9037), .dinb(n8852), .dout(n9038));
  jnot g08975(.din(n9038), .dout(n9039));
  jxor g08976(.dina(n8840), .dinb(n8832), .dout(n9040));
  jand g08977(.dina(n9040), .dinb(n9039), .dout(n9041));
  jnot g08978(.din(n9041), .dout(n9042));
  jand g08979(.dina(n9042), .dinb(n8841), .dout(n9043));
  jnot g08980(.din(n9043), .dout(n9044));
  jxor g08981(.dina(n8829), .dinb(n8821), .dout(n9045));
  jand g08982(.dina(n9045), .dinb(n9044), .dout(n9046));
  jnot g08983(.din(n9046), .dout(n9047));
  jand g08984(.dina(n9047), .dinb(n8830), .dout(n9048));
  jnot g08985(.din(n9048), .dout(n9049));
  jxor g08986(.dina(n8818), .dinb(n8810), .dout(n9050));
  jand g08987(.dina(n9050), .dinb(n9049), .dout(n9051));
  jnot g08988(.din(n9051), .dout(n9052));
  jand g08989(.dina(n9052), .dinb(n8819), .dout(n9053));
  jnot g08990(.din(n9053), .dout(n9054));
  jxor g08991(.dina(n8807), .dinb(n8799), .dout(n9055));
  jand g08992(.dina(n9055), .dinb(n9054), .dout(n9056));
  jnot g08993(.din(n9056), .dout(n9057));
  jand g08994(.dina(n9057), .dinb(n8808), .dout(n9058));
  jnot g08995(.din(n9058), .dout(n9059));
  jxor g08996(.dina(n8796), .dinb(n8788), .dout(n9060));
  jand g08997(.dina(n9060), .dinb(n9059), .dout(n9061));
  jnot g08998(.din(n9061), .dout(n9062));
  jand g08999(.dina(n9062), .dinb(n8797), .dout(n9063));
  jnot g09000(.din(n9063), .dout(n9064));
  jxor g09001(.dina(n8708), .dinb(n8707), .dout(n9065));
  jand g09002(.dina(n9065), .dinb(n9064), .dout(n9066));
  jand g09003(.dina(n6340), .dinb(n5092), .dout(n9067));
  jand g09004(.dina(n6798), .dinb(n1776), .dout(n9068));
  jand g09005(.dina(n6556), .dinb(n1862), .dout(n9069));
  jand g09006(.dina(n6338), .dinb(n1956), .dout(n9070));
  jor  g09007(.dina(n9070), .dinb(n9069), .dout(n9071));
  jor  g09008(.dina(n9071), .dinb(n9068), .dout(n9072));
  jor  g09009(.dina(n9072), .dinb(n9067), .dout(n9073));
  jxor g09010(.dina(n9073), .dinb(n5064), .dout(n9074));
  jnot g09011(.din(n9074), .dout(n9075));
  jxor g09012(.dina(n9065), .dinb(n9064), .dout(n9076));
  jand g09013(.dina(n9076), .dinb(n9075), .dout(n9077));
  jor  g09014(.dina(n9077), .dinb(n9066), .dout(n9078));
  jxor g09015(.dina(n8723), .dinb(n8715), .dout(n9079));
  jand g09016(.dina(n9079), .dinb(n9078), .dout(n9080));
  jnot g09017(.din(n9080), .dout(n9081));
  jxor g09018(.dina(n9079), .dinb(n9078), .dout(n9082));
  jnot g09019(.din(n9082), .dout(n9083));
  jand g09020(.dina(n6936), .dinb(n4258), .dout(n9084));
  jand g09021(.dina(n7741), .dinb(n1343), .dout(n9085));
  jand g09022(.dina(n7613), .dinb(n1445), .dout(n9086));
  jand g09023(.dina(n6934), .dinb(n1560), .dout(n9087));
  jor  g09024(.dina(n9087), .dinb(n9086), .dout(n9088));
  jor  g09025(.dina(n9088), .dinb(n9085), .dout(n9089));
  jor  g09026(.dina(n9089), .dinb(n9084), .dout(n9090));
  jxor g09027(.dina(n9090), .dinb(n5292), .dout(n9091));
  jor  g09028(.dina(n9091), .dinb(n9083), .dout(n9092));
  jand g09029(.dina(n9092), .dinb(n9081), .dout(n9093));
  jnot g09030(.din(n9093), .dout(n9094));
  jxor g09031(.dina(n8739), .dinb(n8731), .dout(n9095));
  jand g09032(.dina(n9095), .dinb(n9094), .dout(n9096));
  jnot g09033(.din(n9096), .dout(n9097));
  jxor g09034(.dina(n9095), .dinb(n9094), .dout(n9098));
  jnot g09035(.din(n9098), .dout(n9099));
  jand g09036(.dina(n7890), .dinb(n3848), .dout(n9100));
  jand g09037(.dina(n8154), .dinb(n922), .dout(n9101));
  jand g09038(.dina(n8441), .dinb(n3853), .dout(n9102));
  jand g09039(.dina(n7888), .dinb(n1076), .dout(n9103));
  jor  g09040(.dina(n9103), .dinb(n9102), .dout(n9104));
  jor  g09041(.dina(n9104), .dinb(n9101), .dout(n9105));
  jor  g09042(.dina(n9105), .dinb(n9100), .dout(n9106));
  jxor g09043(.dina(n9106), .dinb(n5833), .dout(n9107));
  jor  g09044(.dina(n9107), .dinb(n9099), .dout(n9108));
  jand g09045(.dina(n9108), .dinb(n9097), .dout(n9109));
  jand g09046(.dina(n7890), .dinb(n4545), .dout(n9110));
  jand g09047(.dina(n7888), .dinb(n922), .dout(n9111));
  jand g09048(.dina(n8154), .dinb(n3853), .dout(n9112));
  jand g09049(.dina(n8441), .dinb(n4358), .dout(n9113));
  jor  g09050(.dina(n9113), .dinb(n9112), .dout(n9114));
  jor  g09051(.dina(n9114), .dinb(n9111), .dout(n9115));
  jor  g09052(.dina(n9115), .dinb(n9110), .dout(n9116));
  jxor g09053(.dina(n9116), .dinb(n5833), .dout(n9117));
  jor  g09054(.dina(n9117), .dinb(n9109), .dout(n9118));
  jxor g09055(.dina(n9117), .dinb(n9109), .dout(n9119));
  jxor g09056(.dina(n8743), .dinb(n8742), .dout(n9120));
  jand g09057(.dina(n9120), .dinb(n9119), .dout(n9121));
  jnot g09058(.din(n9121), .dout(n9122));
  jand g09059(.dina(n9122), .dinb(n9118), .dout(n9123));
  jor  g09060(.dina(n8772), .dinb(n4731), .dout(n9124));
  jor  g09061(.dina(n8770), .dinb(n4597), .dout(n9125));
  jand g09062(.dina(n8766), .dinb(n8763), .dout(n9126));
  jnot g09063(.din(n9126), .dout(n9127));
  jor  g09064(.dina(n9127), .dinb(n4630), .dout(n9128));
  jand g09065(.dina(n9128), .dinb(n9125), .dout(n9129));
  jand g09066(.dina(n9129), .dinb(n9124), .dout(n9130));
  jxor g09067(.dina(n9130), .dinb(\a[8] ), .dout(n9131));
  jor  g09068(.dina(n9131), .dinb(n9123), .dout(n9132));
  jxor g09069(.dina(n9131), .dinb(n9123), .dout(n9133));
  jxor g09070(.dina(n8760), .dinb(n8752), .dout(n9134));
  jand g09071(.dina(n9134), .dinb(n9133), .dout(n9135));
  jnot g09072(.din(n9135), .dout(n9136));
  jand g09073(.dina(n9136), .dinb(n9132), .dout(n9137));
  jnot g09074(.din(n9137), .dout(n9138));
  jxor g09075(.dina(n8779), .dinb(n8778), .dout(n9139));
  jand g09076(.dina(n9139), .dinb(n9138), .dout(n9140));
  jxor g09077(.dina(n9139), .dinb(n9138), .dout(n9141));
  jand g09078(.dina(n6340), .dinb(n5440), .dout(n9142));
  jand g09079(.dina(n6556), .dinb(n1956), .dout(n9143));
  jand g09080(.dina(n6798), .dinb(n1862), .dout(n9144));
  jand g09081(.dina(n6338), .dinb(n2067), .dout(n9145));
  jor  g09082(.dina(n9145), .dinb(n9144), .dout(n9146));
  jor  g09083(.dina(n9146), .dinb(n9143), .dout(n9147));
  jor  g09084(.dina(n9147), .dinb(n9142), .dout(n9148));
  jxor g09085(.dina(n9148), .dinb(n5064), .dout(n9149));
  jnot g09086(.din(n9149), .dout(n9150));
  jxor g09087(.dina(n9060), .dinb(n9059), .dout(n9151));
  jand g09088(.dina(n9151), .dinb(n9150), .dout(n9152));
  jand g09089(.dina(n6340), .dinb(n5303), .dout(n9153));
  jand g09090(.dina(n6556), .dinb(n2067), .dout(n9154));
  jand g09091(.dina(n6798), .dinb(n1956), .dout(n9155));
  jand g09092(.dina(n6338), .dinb(n2128), .dout(n9156));
  jor  g09093(.dina(n9156), .dinb(n9155), .dout(n9157));
  jor  g09094(.dina(n9157), .dinb(n9154), .dout(n9158));
  jor  g09095(.dina(n9158), .dinb(n9153), .dout(n9159));
  jxor g09096(.dina(n9159), .dinb(n5064), .dout(n9160));
  jnot g09097(.din(n9160), .dout(n9161));
  jxor g09098(.dina(n9055), .dinb(n9054), .dout(n9162));
  jand g09099(.dina(n9162), .dinb(n9161), .dout(n9163));
  jand g09100(.dina(n6340), .dinb(n5624), .dout(n9164));
  jand g09101(.dina(n6338), .dinb(n2237), .dout(n9165));
  jand g09102(.dina(n6556), .dinb(n2128), .dout(n9166));
  jand g09103(.dina(n6798), .dinb(n2067), .dout(n9167));
  jor  g09104(.dina(n9167), .dinb(n9166), .dout(n9168));
  jor  g09105(.dina(n9168), .dinb(n9165), .dout(n9169));
  jor  g09106(.dina(n9169), .dinb(n9164), .dout(n9170));
  jxor g09107(.dina(n9170), .dinb(n5064), .dout(n9171));
  jnot g09108(.din(n9171), .dout(n9172));
  jxor g09109(.dina(n9050), .dinb(n9049), .dout(n9173));
  jand g09110(.dina(n9173), .dinb(n9172), .dout(n9174));
  jand g09111(.dina(n6340), .dinb(n5607), .dout(n9175));
  jand g09112(.dina(n6556), .dinb(n2237), .dout(n9176));
  jand g09113(.dina(n6338), .dinb(n2343), .dout(n9177));
  jand g09114(.dina(n6798), .dinb(n2128), .dout(n9178));
  jor  g09115(.dina(n9178), .dinb(n9177), .dout(n9179));
  jor  g09116(.dina(n9179), .dinb(n9176), .dout(n9180));
  jor  g09117(.dina(n9180), .dinb(n9175), .dout(n9181));
  jxor g09118(.dina(n9181), .dinb(n5064), .dout(n9182));
  jnot g09119(.din(n9182), .dout(n9183));
  jxor g09120(.dina(n9045), .dinb(n9044), .dout(n9184));
  jand g09121(.dina(n9184), .dinb(n9183), .dout(n9185));
  jand g09122(.dina(n6340), .dinb(n5844), .dout(n9186));
  jand g09123(.dina(n6338), .dinb(n2411), .dout(n9187));
  jand g09124(.dina(n6798), .dinb(n2237), .dout(n9188));
  jand g09125(.dina(n6556), .dinb(n2343), .dout(n9189));
  jor  g09126(.dina(n9189), .dinb(n9188), .dout(n9190));
  jor  g09127(.dina(n9190), .dinb(n9187), .dout(n9191));
  jor  g09128(.dina(n9191), .dinb(n9186), .dout(n9192));
  jxor g09129(.dina(n9192), .dinb(n5064), .dout(n9193));
  jnot g09130(.din(n9193), .dout(n9194));
  jxor g09131(.dina(n9040), .dinb(n9039), .dout(n9195));
  jand g09132(.dina(n9195), .dinb(n9194), .dout(n9196));
  jand g09133(.dina(n6340), .dinb(n5861), .dout(n9197));
  jand g09134(.dina(n6556), .dinb(n2411), .dout(n9198));
  jand g09135(.dina(n6798), .dinb(n2343), .dout(n9199));
  jand g09136(.dina(n6338), .dinb(n2497), .dout(n9200));
  jor  g09137(.dina(n9200), .dinb(n9199), .dout(n9201));
  jor  g09138(.dina(n9201), .dinb(n9198), .dout(n9202));
  jor  g09139(.dina(n9202), .dinb(n9197), .dout(n9203));
  jxor g09140(.dina(n9203), .dinb(n5064), .dout(n9204));
  jnot g09141(.din(n9204), .dout(n9205));
  jxor g09142(.dina(n9035), .dinb(n9034), .dout(n9206));
  jand g09143(.dina(n9206), .dinb(n9205), .dout(n9207));
  jand g09144(.dina(n6340), .dinb(n6247), .dout(n9208));
  jand g09145(.dina(n6798), .dinb(n2411), .dout(n9209));
  jand g09146(.dina(n6338), .dinb(n2602), .dout(n9210));
  jand g09147(.dina(n6556), .dinb(n2497), .dout(n9211));
  jor  g09148(.dina(n9211), .dinb(n9210), .dout(n9212));
  jor  g09149(.dina(n9212), .dinb(n9209), .dout(n9213));
  jor  g09150(.dina(n9213), .dinb(n9208), .dout(n9214));
  jxor g09151(.dina(n9214), .dinb(n5064), .dout(n9215));
  jnot g09152(.din(n9215), .dout(n9216));
  jxor g09153(.dina(n9030), .dinb(n9029), .dout(n9217));
  jand g09154(.dina(n9217), .dinb(n9216), .dout(n9218));
  jxor g09155(.dina(n9027), .dinb(n9026), .dout(n9219));
  jnot g09156(.din(n9219), .dout(n9220));
  jand g09157(.dina(n6340), .dinb(n6050), .dout(n9221));
  jand g09158(.dina(n6556), .dinb(n2602), .dout(n9222));
  jand g09159(.dina(n6338), .dinb(n2695), .dout(n9223));
  jand g09160(.dina(n6798), .dinb(n2497), .dout(n9224));
  jor  g09161(.dina(n9224), .dinb(n9223), .dout(n9225));
  jor  g09162(.dina(n9225), .dinb(n9222), .dout(n9226));
  jor  g09163(.dina(n9226), .dinb(n9221), .dout(n9227));
  jxor g09164(.dina(n9227), .dinb(n5064), .dout(n9228));
  jor  g09165(.dina(n9228), .dinb(n9220), .dout(n9229));
  jxor g09166(.dina(n9024), .dinb(n9023), .dout(n9230));
  jnot g09167(.din(n9230), .dout(n9231));
  jor  g09168(.dina(n6464), .dinb(n6341), .dout(n9232));
  jor  g09169(.dina(n6797), .dinb(n2601), .dout(n9233));
  jor  g09170(.dina(n6557), .dinb(n2694), .dout(n9234));
  jor  g09171(.dina(n6339), .dinb(n2731), .dout(n9235));
  jand g09172(.dina(n9235), .dinb(n9234), .dout(n9236));
  jand g09173(.dina(n9236), .dinb(n9233), .dout(n9237));
  jand g09174(.dina(n9237), .dinb(n9232), .dout(n9238));
  jxor g09175(.dina(n9238), .dinb(\a[17] ), .dout(n9239));
  jor  g09176(.dina(n9239), .dinb(n9231), .dout(n9240));
  jand g09177(.dina(n6591), .dinb(n6340), .dout(n9241));
  jand g09178(.dina(n6798), .dinb(n2695), .dout(n9242));
  jand g09179(.dina(n6338), .dinb(n2808), .dout(n9243));
  jand g09180(.dina(n6556), .dinb(n2732), .dout(n9244));
  jor  g09181(.dina(n9244), .dinb(n9243), .dout(n9245));
  jor  g09182(.dina(n9245), .dinb(n9242), .dout(n9246));
  jor  g09183(.dina(n9246), .dinb(n9241), .dout(n9247));
  jxor g09184(.dina(n9247), .dinb(n5064), .dout(n9248));
  jnot g09185(.din(n9248), .dout(n9249));
  jxor g09186(.dina(n9019), .dinb(n9018), .dout(n9250));
  jand g09187(.dina(n9250), .dinb(n9249), .dout(n9251));
  jand g09188(.dina(n6439), .dinb(n6340), .dout(n9252));
  jand g09189(.dina(n6556), .dinb(n2808), .dout(n9253));
  jand g09190(.dina(n6798), .dinb(n2732), .dout(n9254));
  jand g09191(.dina(n6338), .dinb(n2867), .dout(n9255));
  jor  g09192(.dina(n9255), .dinb(n9254), .dout(n9256));
  jor  g09193(.dina(n9256), .dinb(n9253), .dout(n9257));
  jor  g09194(.dina(n9257), .dinb(n9252), .dout(n9258));
  jxor g09195(.dina(n9258), .dinb(n5064), .dout(n9259));
  jnot g09196(.din(n9259), .dout(n9260));
  jxor g09197(.dina(n9014), .dinb(n9013), .dout(n9261));
  jand g09198(.dina(n9261), .dinb(n9260), .dout(n9262));
  jand g09199(.dina(n6706), .dinb(n6340), .dout(n9263));
  jand g09200(.dina(n6798), .dinb(n2808), .dout(n9264));
  jand g09201(.dina(n6338), .dinb(n2954), .dout(n9265));
  jand g09202(.dina(n6556), .dinb(n2867), .dout(n9266));
  jor  g09203(.dina(n9266), .dinb(n9265), .dout(n9267));
  jor  g09204(.dina(n9267), .dinb(n9264), .dout(n9268));
  jor  g09205(.dina(n9268), .dinb(n9263), .dout(n9269));
  jxor g09206(.dina(n9269), .dinb(n5064), .dout(n9270));
  jnot g09207(.din(n9270), .dout(n9271));
  jxor g09208(.dina(n9009), .dinb(n9008), .dout(n9272));
  jand g09209(.dina(n9272), .dinb(n9271), .dout(n9273));
  jxor g09210(.dina(n9006), .dinb(n9005), .dout(n9274));
  jnot g09211(.din(n9274), .dout(n9275));
  jor  g09212(.dina(n6976), .dinb(n6341), .dout(n9276));
  jor  g09213(.dina(n6557), .dinb(n2953), .dout(n9277));
  jor  g09214(.dina(n6339), .dinb(n2990), .dout(n9278));
  jor  g09215(.dina(n6797), .dinb(n2866), .dout(n9279));
  jand g09216(.dina(n9279), .dinb(n9278), .dout(n9280));
  jand g09217(.dina(n9280), .dinb(n9277), .dout(n9281));
  jand g09218(.dina(n9281), .dinb(n9276), .dout(n9282));
  jxor g09219(.dina(n9282), .dinb(\a[17] ), .dout(n9283));
  jor  g09220(.dina(n9283), .dinb(n9275), .dout(n9284));
  jxor g09221(.dina(n9003), .dinb(n9002), .dout(n9285));
  jnot g09222(.din(n9285), .dout(n9286));
  jor  g09223(.dina(n6988), .dinb(n6341), .dout(n9287));
  jor  g09224(.dina(n6339), .dinb(n3085), .dout(n9288));
  jor  g09225(.dina(n6797), .dinb(n2953), .dout(n9289));
  jor  g09226(.dina(n6557), .dinb(n2990), .dout(n9290));
  jand g09227(.dina(n9290), .dinb(n9289), .dout(n9291));
  jand g09228(.dina(n9291), .dinb(n9288), .dout(n9292));
  jand g09229(.dina(n9292), .dinb(n9287), .dout(n9293));
  jxor g09230(.dina(n9293), .dinb(\a[17] ), .dout(n9294));
  jor  g09231(.dina(n9294), .dinb(n9286), .dout(n9295));
  jxor g09232(.dina(n9000), .dinb(n8999), .dout(n9296));
  jnot g09233(.din(n9296), .dout(n9297));
  jor  g09234(.dina(n6681), .dinb(n6341), .dout(n9298));
  jor  g09235(.dina(n6557), .dinb(n3085), .dout(n9299));
  jor  g09236(.dina(n6797), .dinb(n2990), .dout(n9300));
  jor  g09237(.dina(n6339), .dinb(n3182), .dout(n9301));
  jand g09238(.dina(n9301), .dinb(n9300), .dout(n9302));
  jand g09239(.dina(n9302), .dinb(n9299), .dout(n9303));
  jand g09240(.dina(n9303), .dinb(n9298), .dout(n9304));
  jxor g09241(.dina(n9304), .dinb(\a[17] ), .dout(n9305));
  jor  g09242(.dina(n9305), .dinb(n9297), .dout(n9306));
  jor  g09243(.dina(n7031), .dinb(n6341), .dout(n9307));
  jor  g09244(.dina(n6797), .dinb(n3085), .dout(n9308));
  jor  g09245(.dina(n6339), .dinb(n7962), .dout(n9309));
  jor  g09246(.dina(n6557), .dinb(n3182), .dout(n9310));
  jand g09247(.dina(n9310), .dinb(n9309), .dout(n9311));
  jand g09248(.dina(n9311), .dinb(n9308), .dout(n9312));
  jand g09249(.dina(n9312), .dinb(n9307), .dout(n9313));
  jxor g09250(.dina(n9313), .dinb(\a[17] ), .dout(n9314));
  jnot g09251(.din(n9314), .dout(n9315));
  jxor g09252(.dina(n8997), .dinb(n8996), .dout(n9316));
  jand g09253(.dina(n9316), .dinb(n9315), .dout(n9317));
  jor  g09254(.dina(n7076), .dinb(n6341), .dout(n9318));
  jor  g09255(.dina(n6557), .dinb(n7962), .dout(n9319));
  jor  g09256(.dina(n6797), .dinb(n3182), .dout(n9320));
  jor  g09257(.dina(n6339), .dinb(n3684), .dout(n9321));
  jand g09258(.dina(n9321), .dinb(n9320), .dout(n9322));
  jand g09259(.dina(n9322), .dinb(n9319), .dout(n9323));
  jand g09260(.dina(n9323), .dinb(n9318), .dout(n9324));
  jxor g09261(.dina(n9324), .dinb(\a[17] ), .dout(n9325));
  jnot g09262(.din(n9325), .dout(n9326));
  jxor g09263(.dina(n8994), .dinb(n8993), .dout(n9327));
  jand g09264(.dina(n9327), .dinb(n9326), .dout(n9328));
  jor  g09265(.dina(n7131), .dinb(n6341), .dout(n9329));
  jor  g09266(.dina(n6797), .dinb(n7962), .dout(n9330));
  jor  g09267(.dina(n6339), .dinb(n3414), .dout(n9331));
  jor  g09268(.dina(n6557), .dinb(n3684), .dout(n9332));
  jand g09269(.dina(n9332), .dinb(n9331), .dout(n9333));
  jand g09270(.dina(n9333), .dinb(n9330), .dout(n9334));
  jand g09271(.dina(n9334), .dinb(n9329), .dout(n9335));
  jxor g09272(.dina(n9335), .dinb(\a[17] ), .dout(n9336));
  jnot g09273(.din(n9336), .dout(n9337));
  jor  g09274(.dina(n8974), .dinb(n4247), .dout(n9338));
  jxor g09275(.dina(n9338), .dinb(n8982), .dout(n9339));
  jand g09276(.dina(n9339), .dinb(n9337), .dout(n9340));
  jor  g09277(.dina(n7177), .dinb(n6341), .dout(n9341));
  jor  g09278(.dina(n6339), .dinb(n3516), .dout(n9342));
  jor  g09279(.dina(n6797), .dinb(n3684), .dout(n9343));
  jor  g09280(.dina(n6557), .dinb(n3414), .dout(n9344));
  jand g09281(.dina(n9344), .dinb(n9343), .dout(n9345));
  jand g09282(.dina(n9345), .dinb(n9342), .dout(n9346));
  jand g09283(.dina(n9346), .dinb(n9341), .dout(n9347));
  jxor g09284(.dina(n9347), .dinb(\a[17] ), .dout(n9348));
  jnot g09285(.din(n9348), .dout(n9349));
  jand g09286(.dina(n8971), .dinb(\a[20] ), .dout(n9350));
  jxor g09287(.dina(n9350), .dinb(n8969), .dout(n9351));
  jand g09288(.dina(n9351), .dinb(n9349), .dout(n9352));
  jand g09289(.dina(n8004), .dinb(n6340), .dout(n9353));
  jand g09290(.dina(n6556), .dinb(n7411), .dout(n9354));
  jand g09291(.dina(n6798), .dinb(n7405), .dout(n9355));
  jor  g09292(.dina(n9355), .dinb(n9354), .dout(n9356));
  jor  g09293(.dina(n9356), .dinb(n9353), .dout(n9357));
  jnot g09294(.din(n9357), .dout(n9358));
  jand g09295(.dina(n6334), .dinb(n7411), .dout(n9359));
  jnot g09296(.din(n9359), .dout(n9360));
  jand g09297(.dina(n9360), .dinb(\a[17] ), .dout(n9361));
  jand g09298(.dina(n9361), .dinb(n9358), .dout(n9362));
  jand g09299(.dina(n7407), .dinb(n6340), .dout(n9363));
  jand g09300(.dina(n6798), .dinb(n7326), .dout(n9364));
  jand g09301(.dina(n6338), .dinb(n7411), .dout(n9365));
  jand g09302(.dina(n6556), .dinb(n7405), .dout(n9366));
  jor  g09303(.dina(n9366), .dinb(n9365), .dout(n9367));
  jor  g09304(.dina(n9367), .dinb(n9364), .dout(n9368));
  jor  g09305(.dina(n9368), .dinb(n9363), .dout(n9369));
  jnot g09306(.din(n9369), .dout(n9370));
  jand g09307(.dina(n9370), .dinb(n9362), .dout(n9371));
  jand g09308(.dina(n9371), .dinb(n8971), .dout(n9372));
  jor  g09309(.dina(n7466), .dinb(n6341), .dout(n9373));
  jor  g09310(.dina(n6557), .dinb(n3516), .dout(n9374));
  jor  g09311(.dina(n6797), .dinb(n3414), .dout(n9375));
  jor  g09312(.dina(n6339), .dinb(n3677), .dout(n9376));
  jand g09313(.dina(n9376), .dinb(n9375), .dout(n9377));
  jand g09314(.dina(n9377), .dinb(n9374), .dout(n9378));
  jand g09315(.dina(n9378), .dinb(n9373), .dout(n9379));
  jxor g09316(.dina(n9379), .dinb(\a[17] ), .dout(n9380));
  jnot g09317(.din(n9380), .dout(n9381));
  jxor g09318(.dina(n9371), .dinb(n8971), .dout(n9382));
  jand g09319(.dina(n9382), .dinb(n9381), .dout(n9383));
  jor  g09320(.dina(n9383), .dinb(n9372), .dout(n9384));
  jxor g09321(.dina(n9351), .dinb(n9349), .dout(n9385));
  jand g09322(.dina(n9385), .dinb(n9384), .dout(n9386));
  jor  g09323(.dina(n9386), .dinb(n9352), .dout(n9387));
  jxor g09324(.dina(n9339), .dinb(n9337), .dout(n9388));
  jand g09325(.dina(n9388), .dinb(n9387), .dout(n9389));
  jor  g09326(.dina(n9389), .dinb(n9340), .dout(n9390));
  jxor g09327(.dina(n9327), .dinb(n9326), .dout(n9391));
  jand g09328(.dina(n9391), .dinb(n9390), .dout(n9392));
  jor  g09329(.dina(n9392), .dinb(n9328), .dout(n9393));
  jxor g09330(.dina(n9316), .dinb(n9315), .dout(n9394));
  jand g09331(.dina(n9394), .dinb(n9393), .dout(n9395));
  jor  g09332(.dina(n9395), .dinb(n9317), .dout(n9396));
  jxor g09333(.dina(n9305), .dinb(n9297), .dout(n9397));
  jand g09334(.dina(n9397), .dinb(n9396), .dout(n9398));
  jnot g09335(.din(n9398), .dout(n9399));
  jand g09336(.dina(n9399), .dinb(n9306), .dout(n9400));
  jnot g09337(.din(n9400), .dout(n9401));
  jxor g09338(.dina(n9294), .dinb(n9286), .dout(n9402));
  jand g09339(.dina(n9402), .dinb(n9401), .dout(n9403));
  jnot g09340(.din(n9403), .dout(n9404));
  jand g09341(.dina(n9404), .dinb(n9295), .dout(n9405));
  jnot g09342(.din(n9405), .dout(n9406));
  jxor g09343(.dina(n9283), .dinb(n9275), .dout(n9407));
  jand g09344(.dina(n9407), .dinb(n9406), .dout(n9408));
  jnot g09345(.din(n9408), .dout(n9409));
  jand g09346(.dina(n9409), .dinb(n9284), .dout(n9410));
  jnot g09347(.din(n9410), .dout(n9411));
  jxor g09348(.dina(n9272), .dinb(n9271), .dout(n9412));
  jand g09349(.dina(n9412), .dinb(n9411), .dout(n9413));
  jor  g09350(.dina(n9413), .dinb(n9273), .dout(n9414));
  jxor g09351(.dina(n9261), .dinb(n9260), .dout(n9415));
  jand g09352(.dina(n9415), .dinb(n9414), .dout(n9416));
  jor  g09353(.dina(n9416), .dinb(n9262), .dout(n9417));
  jxor g09354(.dina(n9250), .dinb(n9249), .dout(n9418));
  jand g09355(.dina(n9418), .dinb(n9417), .dout(n9419));
  jor  g09356(.dina(n9419), .dinb(n9251), .dout(n9420));
  jxor g09357(.dina(n9239), .dinb(n9231), .dout(n9421));
  jand g09358(.dina(n9421), .dinb(n9420), .dout(n9422));
  jnot g09359(.din(n9422), .dout(n9423));
  jand g09360(.dina(n9423), .dinb(n9240), .dout(n9424));
  jnot g09361(.din(n9424), .dout(n9425));
  jxor g09362(.dina(n9228), .dinb(n9220), .dout(n9426));
  jand g09363(.dina(n9426), .dinb(n9425), .dout(n9427));
  jnot g09364(.din(n9427), .dout(n9428));
  jand g09365(.dina(n9428), .dinb(n9229), .dout(n9429));
  jnot g09366(.din(n9429), .dout(n9430));
  jxor g09367(.dina(n9217), .dinb(n9216), .dout(n9431));
  jand g09368(.dina(n9431), .dinb(n9430), .dout(n9432));
  jor  g09369(.dina(n9432), .dinb(n9218), .dout(n9433));
  jxor g09370(.dina(n9206), .dinb(n9205), .dout(n9434));
  jand g09371(.dina(n9434), .dinb(n9433), .dout(n9435));
  jor  g09372(.dina(n9435), .dinb(n9207), .dout(n9436));
  jxor g09373(.dina(n9195), .dinb(n9194), .dout(n9437));
  jand g09374(.dina(n9437), .dinb(n9436), .dout(n9438));
  jor  g09375(.dina(n9438), .dinb(n9196), .dout(n9439));
  jxor g09376(.dina(n9184), .dinb(n9183), .dout(n9440));
  jand g09377(.dina(n9440), .dinb(n9439), .dout(n9441));
  jor  g09378(.dina(n9441), .dinb(n9185), .dout(n9442));
  jxor g09379(.dina(n9173), .dinb(n9172), .dout(n9443));
  jand g09380(.dina(n9443), .dinb(n9442), .dout(n9444));
  jor  g09381(.dina(n9444), .dinb(n9174), .dout(n9445));
  jxor g09382(.dina(n9162), .dinb(n9161), .dout(n9446));
  jand g09383(.dina(n9446), .dinb(n9445), .dout(n9447));
  jor  g09384(.dina(n9447), .dinb(n9163), .dout(n9448));
  jxor g09385(.dina(n9151), .dinb(n9150), .dout(n9449));
  jand g09386(.dina(n9449), .dinb(n9448), .dout(n9450));
  jor  g09387(.dina(n9450), .dinb(n9152), .dout(n9451));
  jxor g09388(.dina(n9076), .dinb(n9075), .dout(n9452));
  jand g09389(.dina(n9452), .dinb(n9451), .dout(n9453));
  jand g09390(.dina(n6936), .dinb(n4866), .dout(n9454));
  jand g09391(.dina(n7741), .dinb(n1445), .dout(n9455));
  jand g09392(.dina(n7613), .dinb(n1560), .dout(n9456));
  jand g09393(.dina(n6934), .dinb(n1624), .dout(n9457));
  jor  g09394(.dina(n9457), .dinb(n9456), .dout(n9458));
  jor  g09395(.dina(n9458), .dinb(n9455), .dout(n9459));
  jor  g09396(.dina(n9459), .dinb(n9454), .dout(n9460));
  jxor g09397(.dina(n9460), .dinb(n5292), .dout(n9461));
  jnot g09398(.din(n9461), .dout(n9462));
  jxor g09399(.dina(n9452), .dinb(n9451), .dout(n9463));
  jand g09400(.dina(n9463), .dinb(n9462), .dout(n9464));
  jor  g09401(.dina(n9464), .dinb(n9453), .dout(n9465));
  jxor g09402(.dina(n9091), .dinb(n9083), .dout(n9466));
  jand g09403(.dina(n9466), .dinb(n9465), .dout(n9467));
  jnot g09404(.din(n9467), .dout(n9468));
  jxor g09405(.dina(n9466), .dinb(n9465), .dout(n9469));
  jnot g09406(.din(n9469), .dout(n9470));
  jand g09407(.dina(n7890), .dinb(n4026), .dout(n9471));
  jand g09408(.dina(n8154), .dinb(n1076), .dout(n9472));
  jand g09409(.dina(n8441), .dinb(n922), .dout(n9473));
  jand g09410(.dina(n7888), .dinb(n1213), .dout(n9474));
  jor  g09411(.dina(n9474), .dinb(n9473), .dout(n9475));
  jor  g09412(.dina(n9475), .dinb(n9472), .dout(n9476));
  jor  g09413(.dina(n9476), .dinb(n9471), .dout(n9477));
  jxor g09414(.dina(n9477), .dinb(n5833), .dout(n9478));
  jor  g09415(.dina(n9478), .dinb(n9470), .dout(n9479));
  jand g09416(.dina(n9479), .dinb(n9468), .dout(n9480));
  jnot g09417(.din(n9480), .dout(n9481));
  jxor g09418(.dina(n9107), .dinb(n9099), .dout(n9482));
  jand g09419(.dina(n9482), .dinb(n9481), .dout(n9483));
  jnot g09420(.din(n9483), .dout(n9484));
  jxor g09421(.dina(n9482), .dinb(n9481), .dout(n9485));
  jnot g09422(.din(n9485), .dout(n9486));
  jand g09423(.dina(n8771), .dinb(n4752), .dout(n9487));
  jand g09424(.dina(n9126), .dinb(n4451), .dout(n9488));
  jand g09425(.dina(n8769), .dinb(n4358), .dout(n9489));
  jor  g09426(.dina(n8768), .dinb(n8766), .dout(n9490));
  jnot g09427(.din(n9490), .dout(n9491));
  jand g09428(.dina(n9491), .dinb(n4598), .dout(n9492));
  jor  g09429(.dina(n9492), .dinb(n9489), .dout(n9493));
  jor  g09430(.dina(n9493), .dinb(n9488), .dout(n9494));
  jor  g09431(.dina(n9494), .dinb(n9487), .dout(n9495));
  jxor g09432(.dina(n9495), .dinb(n6039), .dout(n9496));
  jor  g09433(.dina(n9496), .dinb(n9486), .dout(n9497));
  jand g09434(.dina(n9497), .dinb(n9484), .dout(n9498));
  jand g09435(.dina(n8771), .dinb(n4636), .dout(n9499));
  jand g09436(.dina(n8769), .dinb(n4451), .dout(n9500));
  jand g09437(.dina(n9126), .dinb(n4598), .dout(n9501));
  jand g09438(.dina(n9491), .dinb(n4631), .dout(n9502));
  jor  g09439(.dina(n9502), .dinb(n9501), .dout(n9503));
  jor  g09440(.dina(n9503), .dinb(n9500), .dout(n9504));
  jor  g09441(.dina(n9504), .dinb(n9499), .dout(n9505));
  jxor g09442(.dina(n9505), .dinb(n6039), .dout(n9506));
  jor  g09443(.dina(n9506), .dinb(n9498), .dout(n9507));
  jxor g09444(.dina(n9120), .dinb(n9119), .dout(n9508));
  jxor g09445(.dina(n9506), .dinb(n9498), .dout(n9509));
  jand g09446(.dina(n9509), .dinb(n9508), .dout(n9510));
  jnot g09447(.din(n9510), .dout(n9511));
  jand g09448(.dina(n9511), .dinb(n9507), .dout(n9512));
  jnot g09449(.din(n9512), .dout(n9513));
  jxor g09450(.dina(n9134), .dinb(n9133), .dout(n9514));
  jand g09451(.dina(n9514), .dinb(n9513), .dout(n9515));
  jxor g09452(.dina(n9449), .dinb(n9448), .dout(n9516));
  jnot g09453(.din(n9516), .dout(n9517));
  jand g09454(.dina(n6936), .dinb(n4849), .dout(n9518));
  jand g09455(.dina(n7613), .dinb(n1624), .dout(n9519));
  jand g09456(.dina(n6934), .dinb(n1776), .dout(n9520));
  jand g09457(.dina(n7741), .dinb(n1560), .dout(n9521));
  jor  g09458(.dina(n9521), .dinb(n9520), .dout(n9522));
  jor  g09459(.dina(n9522), .dinb(n9519), .dout(n9523));
  jor  g09460(.dina(n9523), .dinb(n9518), .dout(n9524));
  jxor g09461(.dina(n9524), .dinb(n5292), .dout(n9525));
  jor  g09462(.dina(n9525), .dinb(n9517), .dout(n9526));
  jxor g09463(.dina(n9446), .dinb(n9445), .dout(n9527));
  jnot g09464(.din(n9527), .dout(n9528));
  jand g09465(.dina(n6936), .dinb(n5075), .dout(n9529));
  jand g09466(.dina(n7613), .dinb(n1776), .dout(n9530));
  jand g09467(.dina(n6934), .dinb(n1862), .dout(n9531));
  jand g09468(.dina(n7741), .dinb(n1624), .dout(n9532));
  jor  g09469(.dina(n9532), .dinb(n9531), .dout(n9533));
  jor  g09470(.dina(n9533), .dinb(n9530), .dout(n9534));
  jor  g09471(.dina(n9534), .dinb(n9529), .dout(n9535));
  jxor g09472(.dina(n9535), .dinb(n5292), .dout(n9536));
  jor  g09473(.dina(n9536), .dinb(n9528), .dout(n9537));
  jxor g09474(.dina(n9443), .dinb(n9442), .dout(n9538));
  jnot g09475(.din(n9538), .dout(n9539));
  jand g09476(.dina(n6936), .dinb(n5092), .dout(n9540));
  jand g09477(.dina(n7613), .dinb(n1862), .dout(n9541));
  jand g09478(.dina(n6934), .dinb(n1956), .dout(n9542));
  jand g09479(.dina(n7741), .dinb(n1776), .dout(n9543));
  jor  g09480(.dina(n9543), .dinb(n9542), .dout(n9544));
  jor  g09481(.dina(n9544), .dinb(n9541), .dout(n9545));
  jor  g09482(.dina(n9545), .dinb(n9540), .dout(n9546));
  jxor g09483(.dina(n9546), .dinb(n5292), .dout(n9547));
  jor  g09484(.dina(n9547), .dinb(n9539), .dout(n9548));
  jxor g09485(.dina(n9440), .dinb(n9439), .dout(n9549));
  jnot g09486(.din(n9549), .dout(n9550));
  jand g09487(.dina(n6936), .dinb(n5440), .dout(n9551));
  jand g09488(.dina(n6934), .dinb(n2067), .dout(n9552));
  jand g09489(.dina(n7613), .dinb(n1956), .dout(n9553));
  jand g09490(.dina(n7741), .dinb(n1862), .dout(n9554));
  jor  g09491(.dina(n9554), .dinb(n9553), .dout(n9555));
  jor  g09492(.dina(n9555), .dinb(n9552), .dout(n9556));
  jor  g09493(.dina(n9556), .dinb(n9551), .dout(n9557));
  jxor g09494(.dina(n9557), .dinb(n5292), .dout(n9558));
  jor  g09495(.dina(n9558), .dinb(n9550), .dout(n9559));
  jxor g09496(.dina(n9437), .dinb(n9436), .dout(n9560));
  jnot g09497(.din(n9560), .dout(n9561));
  jand g09498(.dina(n6936), .dinb(n5303), .dout(n9562));
  jand g09499(.dina(n6934), .dinb(n2128), .dout(n9563));
  jand g09500(.dina(n7613), .dinb(n2067), .dout(n9564));
  jand g09501(.dina(n7741), .dinb(n1956), .dout(n9565));
  jor  g09502(.dina(n9565), .dinb(n9564), .dout(n9566));
  jor  g09503(.dina(n9566), .dinb(n9563), .dout(n9567));
  jor  g09504(.dina(n9567), .dinb(n9562), .dout(n9568));
  jxor g09505(.dina(n9568), .dinb(n5292), .dout(n9569));
  jor  g09506(.dina(n9569), .dinb(n9561), .dout(n9570));
  jxor g09507(.dina(n9434), .dinb(n9433), .dout(n9571));
  jnot g09508(.din(n9571), .dout(n9572));
  jand g09509(.dina(n6936), .dinb(n5624), .dout(n9573));
  jand g09510(.dina(n6934), .dinb(n2237), .dout(n9574));
  jand g09511(.dina(n7613), .dinb(n2128), .dout(n9575));
  jand g09512(.dina(n7741), .dinb(n2067), .dout(n9576));
  jor  g09513(.dina(n9576), .dinb(n9575), .dout(n9577));
  jor  g09514(.dina(n9577), .dinb(n9574), .dout(n9578));
  jor  g09515(.dina(n9578), .dinb(n9573), .dout(n9579));
  jxor g09516(.dina(n9579), .dinb(n5292), .dout(n9580));
  jor  g09517(.dina(n9580), .dinb(n9572), .dout(n9581));
  jxor g09518(.dina(n9431), .dinb(n9430), .dout(n9582));
  jnot g09519(.din(n9582), .dout(n9583));
  jand g09520(.dina(n6936), .dinb(n5607), .dout(n9584));
  jand g09521(.dina(n7613), .dinb(n2237), .dout(n9585));
  jand g09522(.dina(n6934), .dinb(n2343), .dout(n9586));
  jand g09523(.dina(n7741), .dinb(n2128), .dout(n9587));
  jor  g09524(.dina(n9587), .dinb(n9586), .dout(n9588));
  jor  g09525(.dina(n9588), .dinb(n9585), .dout(n9589));
  jor  g09526(.dina(n9589), .dinb(n9584), .dout(n9590));
  jxor g09527(.dina(n9590), .dinb(n5292), .dout(n9591));
  jor  g09528(.dina(n9591), .dinb(n9583), .dout(n9592));
  jand g09529(.dina(n6936), .dinb(n5844), .dout(n9593));
  jand g09530(.dina(n6934), .dinb(n2411), .dout(n9594));
  jand g09531(.dina(n7741), .dinb(n2237), .dout(n9595));
  jand g09532(.dina(n7613), .dinb(n2343), .dout(n9596));
  jor  g09533(.dina(n9596), .dinb(n9595), .dout(n9597));
  jor  g09534(.dina(n9597), .dinb(n9594), .dout(n9598));
  jor  g09535(.dina(n9598), .dinb(n9593), .dout(n9599));
  jxor g09536(.dina(n9599), .dinb(n5292), .dout(n9600));
  jnot g09537(.din(n9600), .dout(n9601));
  jxor g09538(.dina(n9426), .dinb(n9425), .dout(n9602));
  jand g09539(.dina(n9602), .dinb(n9601), .dout(n9603));
  jand g09540(.dina(n6936), .dinb(n5861), .dout(n9604));
  jand g09541(.dina(n7613), .dinb(n2411), .dout(n9605));
  jand g09542(.dina(n7741), .dinb(n2343), .dout(n9606));
  jand g09543(.dina(n6934), .dinb(n2497), .dout(n9607));
  jor  g09544(.dina(n9607), .dinb(n9606), .dout(n9608));
  jor  g09545(.dina(n9608), .dinb(n9605), .dout(n9609));
  jor  g09546(.dina(n9609), .dinb(n9604), .dout(n9610));
  jxor g09547(.dina(n9610), .dinb(n5292), .dout(n9611));
  jnot g09548(.din(n9611), .dout(n9612));
  jxor g09549(.dina(n9421), .dinb(n9420), .dout(n9613));
  jand g09550(.dina(n9613), .dinb(n9612), .dout(n9614));
  jxor g09551(.dina(n9418), .dinb(n9417), .dout(n9615));
  jnot g09552(.din(n9615), .dout(n9616));
  jand g09553(.dina(n6936), .dinb(n6247), .dout(n9617));
  jand g09554(.dina(n7741), .dinb(n2411), .dout(n9618));
  jand g09555(.dina(n6934), .dinb(n2602), .dout(n9619));
  jand g09556(.dina(n7613), .dinb(n2497), .dout(n9620));
  jor  g09557(.dina(n9620), .dinb(n9619), .dout(n9621));
  jor  g09558(.dina(n9621), .dinb(n9618), .dout(n9622));
  jor  g09559(.dina(n9622), .dinb(n9617), .dout(n9623));
  jxor g09560(.dina(n9623), .dinb(n5292), .dout(n9624));
  jor  g09561(.dina(n9624), .dinb(n9616), .dout(n9625));
  jxor g09562(.dina(n9415), .dinb(n9414), .dout(n9626));
  jnot g09563(.din(n9626), .dout(n9627));
  jand g09564(.dina(n6936), .dinb(n6050), .dout(n9628));
  jand g09565(.dina(n7613), .dinb(n2602), .dout(n9629));
  jand g09566(.dina(n6934), .dinb(n2695), .dout(n9630));
  jand g09567(.dina(n7741), .dinb(n2497), .dout(n9631));
  jor  g09568(.dina(n9631), .dinb(n9630), .dout(n9632));
  jor  g09569(.dina(n9632), .dinb(n9629), .dout(n9633));
  jor  g09570(.dina(n9633), .dinb(n9628), .dout(n9634));
  jxor g09571(.dina(n9634), .dinb(n5292), .dout(n9635));
  jor  g09572(.dina(n9635), .dinb(n9627), .dout(n9636));
  jxor g09573(.dina(n9412), .dinb(n9411), .dout(n9637));
  jnot g09574(.din(n9637), .dout(n9638));
  jor  g09575(.dina(n6937), .dinb(n6464), .dout(n9639));
  jor  g09576(.dina(n7740), .dinb(n2601), .dout(n9640));
  jor  g09577(.dina(n7614), .dinb(n2694), .dout(n9641));
  jor  g09578(.dina(n6935), .dinb(n2731), .dout(n9642));
  jand g09579(.dina(n9642), .dinb(n9641), .dout(n9643));
  jand g09580(.dina(n9643), .dinb(n9640), .dout(n9644));
  jand g09581(.dina(n9644), .dinb(n9639), .dout(n9645));
  jxor g09582(.dina(n9645), .dinb(\a[14] ), .dout(n9646));
  jor  g09583(.dina(n9646), .dinb(n9638), .dout(n9647));
  jand g09584(.dina(n6936), .dinb(n6591), .dout(n9648));
  jand g09585(.dina(n7741), .dinb(n2695), .dout(n9649));
  jand g09586(.dina(n6934), .dinb(n2808), .dout(n9650));
  jand g09587(.dina(n7613), .dinb(n2732), .dout(n9651));
  jor  g09588(.dina(n9651), .dinb(n9650), .dout(n9652));
  jor  g09589(.dina(n9652), .dinb(n9649), .dout(n9653));
  jor  g09590(.dina(n9653), .dinb(n9648), .dout(n9654));
  jxor g09591(.dina(n9654), .dinb(n5292), .dout(n9655));
  jnot g09592(.din(n9655), .dout(n9656));
  jxor g09593(.dina(n9407), .dinb(n9406), .dout(n9657));
  jand g09594(.dina(n9657), .dinb(n9656), .dout(n9658));
  jand g09595(.dina(n6936), .dinb(n6439), .dout(n9659));
  jand g09596(.dina(n7613), .dinb(n2808), .dout(n9660));
  jand g09597(.dina(n7741), .dinb(n2732), .dout(n9661));
  jand g09598(.dina(n6934), .dinb(n2867), .dout(n9662));
  jor  g09599(.dina(n9662), .dinb(n9661), .dout(n9663));
  jor  g09600(.dina(n9663), .dinb(n9660), .dout(n9664));
  jor  g09601(.dina(n9664), .dinb(n9659), .dout(n9665));
  jxor g09602(.dina(n9665), .dinb(n5292), .dout(n9666));
  jnot g09603(.din(n9666), .dout(n9667));
  jxor g09604(.dina(n9402), .dinb(n9401), .dout(n9668));
  jand g09605(.dina(n9668), .dinb(n9667), .dout(n9669));
  jand g09606(.dina(n6936), .dinb(n6706), .dout(n9670));
  jand g09607(.dina(n7741), .dinb(n2808), .dout(n9671));
  jand g09608(.dina(n6934), .dinb(n2954), .dout(n9672));
  jand g09609(.dina(n7613), .dinb(n2867), .dout(n9673));
  jor  g09610(.dina(n9673), .dinb(n9672), .dout(n9674));
  jor  g09611(.dina(n9674), .dinb(n9671), .dout(n9675));
  jor  g09612(.dina(n9675), .dinb(n9670), .dout(n9676));
  jxor g09613(.dina(n9676), .dinb(n5292), .dout(n9677));
  jnot g09614(.din(n9677), .dout(n9678));
  jxor g09615(.dina(n9397), .dinb(n9396), .dout(n9679));
  jand g09616(.dina(n9679), .dinb(n9678), .dout(n9680));
  jxor g09617(.dina(n9394), .dinb(n9393), .dout(n9681));
  jnot g09618(.din(n9681), .dout(n9682));
  jor  g09619(.dina(n6976), .dinb(n6937), .dout(n9683));
  jor  g09620(.dina(n7614), .dinb(n2953), .dout(n9684));
  jor  g09621(.dina(n6935), .dinb(n2990), .dout(n9685));
  jor  g09622(.dina(n7740), .dinb(n2866), .dout(n9686));
  jand g09623(.dina(n9686), .dinb(n9685), .dout(n9687));
  jand g09624(.dina(n9687), .dinb(n9684), .dout(n9688));
  jand g09625(.dina(n9688), .dinb(n9683), .dout(n9689));
  jxor g09626(.dina(n9689), .dinb(\a[14] ), .dout(n9690));
  jor  g09627(.dina(n9690), .dinb(n9682), .dout(n9691));
  jxor g09628(.dina(n9391), .dinb(n9390), .dout(n9692));
  jnot g09629(.din(n9692), .dout(n9693));
  jor  g09630(.dina(n6988), .dinb(n6937), .dout(n9694));
  jor  g09631(.dina(n6935), .dinb(n3085), .dout(n9695));
  jor  g09632(.dina(n7740), .dinb(n2953), .dout(n9696));
  jor  g09633(.dina(n7614), .dinb(n2990), .dout(n9697));
  jand g09634(.dina(n9697), .dinb(n9696), .dout(n9698));
  jand g09635(.dina(n9698), .dinb(n9695), .dout(n9699));
  jand g09636(.dina(n9699), .dinb(n9694), .dout(n9700));
  jxor g09637(.dina(n9700), .dinb(\a[14] ), .dout(n9701));
  jor  g09638(.dina(n9701), .dinb(n9693), .dout(n9702));
  jxor g09639(.dina(n9388), .dinb(n9387), .dout(n9703));
  jnot g09640(.din(n9703), .dout(n9704));
  jor  g09641(.dina(n6937), .dinb(n6681), .dout(n9705));
  jor  g09642(.dina(n7614), .dinb(n3085), .dout(n9706));
  jor  g09643(.dina(n7740), .dinb(n2990), .dout(n9707));
  jor  g09644(.dina(n6935), .dinb(n3182), .dout(n9708));
  jand g09645(.dina(n9708), .dinb(n9707), .dout(n9709));
  jand g09646(.dina(n9709), .dinb(n9706), .dout(n9710));
  jand g09647(.dina(n9710), .dinb(n9705), .dout(n9711));
  jxor g09648(.dina(n9711), .dinb(\a[14] ), .dout(n9712));
  jor  g09649(.dina(n9712), .dinb(n9704), .dout(n9713));
  jor  g09650(.dina(n7031), .dinb(n6937), .dout(n9714));
  jor  g09651(.dina(n7740), .dinb(n3085), .dout(n9715));
  jor  g09652(.dina(n6935), .dinb(n7962), .dout(n9716));
  jor  g09653(.dina(n7614), .dinb(n3182), .dout(n9717));
  jand g09654(.dina(n9717), .dinb(n9716), .dout(n9718));
  jand g09655(.dina(n9718), .dinb(n9715), .dout(n9719));
  jand g09656(.dina(n9719), .dinb(n9714), .dout(n9720));
  jxor g09657(.dina(n9720), .dinb(\a[14] ), .dout(n9721));
  jnot g09658(.din(n9721), .dout(n9722));
  jxor g09659(.dina(n9385), .dinb(n9384), .dout(n9723));
  jand g09660(.dina(n9723), .dinb(n9722), .dout(n9724));
  jor  g09661(.dina(n7076), .dinb(n6937), .dout(n9725));
  jor  g09662(.dina(n7614), .dinb(n7962), .dout(n9726));
  jor  g09663(.dina(n7740), .dinb(n3182), .dout(n9727));
  jor  g09664(.dina(n6935), .dinb(n3684), .dout(n9728));
  jand g09665(.dina(n9728), .dinb(n9727), .dout(n9729));
  jand g09666(.dina(n9729), .dinb(n9726), .dout(n9730));
  jand g09667(.dina(n9730), .dinb(n9725), .dout(n9731));
  jxor g09668(.dina(n9731), .dinb(\a[14] ), .dout(n9732));
  jnot g09669(.din(n9732), .dout(n9733));
  jxor g09670(.dina(n9382), .dinb(n9381), .dout(n9734));
  jand g09671(.dina(n9734), .dinb(n9733), .dout(n9735));
  jor  g09672(.dina(n7131), .dinb(n6937), .dout(n9736));
  jor  g09673(.dina(n7740), .dinb(n7962), .dout(n9737));
  jor  g09674(.dina(n6935), .dinb(n3414), .dout(n9738));
  jor  g09675(.dina(n7614), .dinb(n3684), .dout(n9739));
  jand g09676(.dina(n9739), .dinb(n9738), .dout(n9740));
  jand g09677(.dina(n9740), .dinb(n9737), .dout(n9741));
  jand g09678(.dina(n9741), .dinb(n9736), .dout(n9742));
  jxor g09679(.dina(n9742), .dinb(\a[14] ), .dout(n9743));
  jnot g09680(.din(n9743), .dout(n9744));
  jor  g09681(.dina(n9362), .dinb(n5064), .dout(n9745));
  jxor g09682(.dina(n9745), .dinb(n9370), .dout(n9746));
  jand g09683(.dina(n9746), .dinb(n9744), .dout(n9747));
  jor  g09684(.dina(n7177), .dinb(n6937), .dout(n9748));
  jor  g09685(.dina(n6935), .dinb(n3516), .dout(n9749));
  jor  g09686(.dina(n7740), .dinb(n3684), .dout(n9750));
  jor  g09687(.dina(n7614), .dinb(n3414), .dout(n9751));
  jand g09688(.dina(n9751), .dinb(n9750), .dout(n9752));
  jand g09689(.dina(n9752), .dinb(n9749), .dout(n9753));
  jand g09690(.dina(n9753), .dinb(n9748), .dout(n9754));
  jxor g09691(.dina(n9754), .dinb(\a[14] ), .dout(n9755));
  jnot g09692(.din(n9755), .dout(n9756));
  jand g09693(.dina(n9359), .dinb(\a[17] ), .dout(n9757));
  jxor g09694(.dina(n9757), .dinb(n9357), .dout(n9758));
  jand g09695(.dina(n9758), .dinb(n9756), .dout(n9759));
  jand g09696(.dina(n8004), .dinb(n6936), .dout(n9760));
  jand g09697(.dina(n7613), .dinb(n7411), .dout(n9761));
  jand g09698(.dina(n7741), .dinb(n7405), .dout(n9762));
  jor  g09699(.dina(n9762), .dinb(n9761), .dout(n9763));
  jor  g09700(.dina(n9763), .dinb(n9760), .dout(n9764));
  jnot g09701(.din(n9764), .dout(n9765));
  jand g09702(.dina(n6928), .dinb(n7411), .dout(n9766));
  jnot g09703(.din(n9766), .dout(n9767));
  jand g09704(.dina(n9767), .dinb(\a[14] ), .dout(n9768));
  jand g09705(.dina(n9768), .dinb(n9765), .dout(n9769));
  jand g09706(.dina(n7407), .dinb(n6936), .dout(n9770));
  jand g09707(.dina(n7741), .dinb(n7326), .dout(n9771));
  jand g09708(.dina(n6934), .dinb(n7411), .dout(n9772));
  jand g09709(.dina(n7613), .dinb(n7405), .dout(n9773));
  jor  g09710(.dina(n9773), .dinb(n9772), .dout(n9774));
  jor  g09711(.dina(n9774), .dinb(n9771), .dout(n9775));
  jor  g09712(.dina(n9775), .dinb(n9770), .dout(n9776));
  jnot g09713(.din(n9776), .dout(n9777));
  jand g09714(.dina(n9777), .dinb(n9769), .dout(n9778));
  jand g09715(.dina(n9778), .dinb(n9359), .dout(n9779));
  jor  g09716(.dina(n7466), .dinb(n6937), .dout(n9780));
  jor  g09717(.dina(n7614), .dinb(n3516), .dout(n9781));
  jor  g09718(.dina(n7740), .dinb(n3414), .dout(n9782));
  jor  g09719(.dina(n6935), .dinb(n3677), .dout(n9783));
  jand g09720(.dina(n9783), .dinb(n9782), .dout(n9784));
  jand g09721(.dina(n9784), .dinb(n9781), .dout(n9785));
  jand g09722(.dina(n9785), .dinb(n9780), .dout(n9786));
  jxor g09723(.dina(n9786), .dinb(\a[14] ), .dout(n9787));
  jnot g09724(.din(n9787), .dout(n9788));
  jxor g09725(.dina(n9778), .dinb(n9359), .dout(n9789));
  jand g09726(.dina(n9789), .dinb(n9788), .dout(n9790));
  jor  g09727(.dina(n9790), .dinb(n9779), .dout(n9791));
  jxor g09728(.dina(n9758), .dinb(n9756), .dout(n9792));
  jand g09729(.dina(n9792), .dinb(n9791), .dout(n9793));
  jor  g09730(.dina(n9793), .dinb(n9759), .dout(n9794));
  jxor g09731(.dina(n9746), .dinb(n9744), .dout(n9795));
  jand g09732(.dina(n9795), .dinb(n9794), .dout(n9796));
  jor  g09733(.dina(n9796), .dinb(n9747), .dout(n9797));
  jxor g09734(.dina(n9734), .dinb(n9733), .dout(n9798));
  jand g09735(.dina(n9798), .dinb(n9797), .dout(n9799));
  jor  g09736(.dina(n9799), .dinb(n9735), .dout(n9800));
  jxor g09737(.dina(n9723), .dinb(n9722), .dout(n9801));
  jand g09738(.dina(n9801), .dinb(n9800), .dout(n9802));
  jor  g09739(.dina(n9802), .dinb(n9724), .dout(n9803));
  jxor g09740(.dina(n9712), .dinb(n9704), .dout(n9804));
  jand g09741(.dina(n9804), .dinb(n9803), .dout(n9805));
  jnot g09742(.din(n9805), .dout(n9806));
  jand g09743(.dina(n9806), .dinb(n9713), .dout(n9807));
  jnot g09744(.din(n9807), .dout(n9808));
  jxor g09745(.dina(n9701), .dinb(n9693), .dout(n9809));
  jand g09746(.dina(n9809), .dinb(n9808), .dout(n9810));
  jnot g09747(.din(n9810), .dout(n9811));
  jand g09748(.dina(n9811), .dinb(n9702), .dout(n9812));
  jnot g09749(.din(n9812), .dout(n9813));
  jxor g09750(.dina(n9690), .dinb(n9682), .dout(n9814));
  jand g09751(.dina(n9814), .dinb(n9813), .dout(n9815));
  jnot g09752(.din(n9815), .dout(n9816));
  jand g09753(.dina(n9816), .dinb(n9691), .dout(n9817));
  jnot g09754(.din(n9817), .dout(n9818));
  jxor g09755(.dina(n9679), .dinb(n9678), .dout(n9819));
  jand g09756(.dina(n9819), .dinb(n9818), .dout(n9820));
  jor  g09757(.dina(n9820), .dinb(n9680), .dout(n9821));
  jxor g09758(.dina(n9668), .dinb(n9667), .dout(n9822));
  jand g09759(.dina(n9822), .dinb(n9821), .dout(n9823));
  jor  g09760(.dina(n9823), .dinb(n9669), .dout(n9824));
  jxor g09761(.dina(n9657), .dinb(n9656), .dout(n9825));
  jand g09762(.dina(n9825), .dinb(n9824), .dout(n9826));
  jor  g09763(.dina(n9826), .dinb(n9658), .dout(n9827));
  jxor g09764(.dina(n9646), .dinb(n9638), .dout(n9828));
  jand g09765(.dina(n9828), .dinb(n9827), .dout(n9829));
  jnot g09766(.din(n9829), .dout(n9830));
  jand g09767(.dina(n9830), .dinb(n9647), .dout(n9831));
  jnot g09768(.din(n9831), .dout(n9832));
  jxor g09769(.dina(n9635), .dinb(n9627), .dout(n9833));
  jand g09770(.dina(n9833), .dinb(n9832), .dout(n9834));
  jnot g09771(.din(n9834), .dout(n9835));
  jand g09772(.dina(n9835), .dinb(n9636), .dout(n9836));
  jnot g09773(.din(n9836), .dout(n9837));
  jxor g09774(.dina(n9624), .dinb(n9616), .dout(n9838));
  jand g09775(.dina(n9838), .dinb(n9837), .dout(n9839));
  jnot g09776(.din(n9839), .dout(n9840));
  jand g09777(.dina(n9840), .dinb(n9625), .dout(n9841));
  jnot g09778(.din(n9841), .dout(n9842));
  jxor g09779(.dina(n9613), .dinb(n9612), .dout(n9843));
  jand g09780(.dina(n9843), .dinb(n9842), .dout(n9844));
  jor  g09781(.dina(n9844), .dinb(n9614), .dout(n9845));
  jxor g09782(.dina(n9602), .dinb(n9601), .dout(n9846));
  jand g09783(.dina(n9846), .dinb(n9845), .dout(n9847));
  jor  g09784(.dina(n9847), .dinb(n9603), .dout(n9848));
  jxor g09785(.dina(n9591), .dinb(n9583), .dout(n9849));
  jand g09786(.dina(n9849), .dinb(n9848), .dout(n9850));
  jnot g09787(.din(n9850), .dout(n9851));
  jand g09788(.dina(n9851), .dinb(n9592), .dout(n9852));
  jnot g09789(.din(n9852), .dout(n9853));
  jxor g09790(.dina(n9580), .dinb(n9572), .dout(n9854));
  jand g09791(.dina(n9854), .dinb(n9853), .dout(n9855));
  jnot g09792(.din(n9855), .dout(n9856));
  jand g09793(.dina(n9856), .dinb(n9581), .dout(n9857));
  jnot g09794(.din(n9857), .dout(n9858));
  jxor g09795(.dina(n9569), .dinb(n9561), .dout(n9859));
  jand g09796(.dina(n9859), .dinb(n9858), .dout(n9860));
  jnot g09797(.din(n9860), .dout(n9861));
  jand g09798(.dina(n9861), .dinb(n9570), .dout(n9862));
  jnot g09799(.din(n9862), .dout(n9863));
  jxor g09800(.dina(n9558), .dinb(n9550), .dout(n9864));
  jand g09801(.dina(n9864), .dinb(n9863), .dout(n9865));
  jnot g09802(.din(n9865), .dout(n9866));
  jand g09803(.dina(n9866), .dinb(n9559), .dout(n9867));
  jnot g09804(.din(n9867), .dout(n9868));
  jxor g09805(.dina(n9547), .dinb(n9539), .dout(n9869));
  jand g09806(.dina(n9869), .dinb(n9868), .dout(n9870));
  jnot g09807(.din(n9870), .dout(n9871));
  jand g09808(.dina(n9871), .dinb(n9548), .dout(n9872));
  jnot g09809(.din(n9872), .dout(n9873));
  jxor g09810(.dina(n9536), .dinb(n9528), .dout(n9874));
  jand g09811(.dina(n9874), .dinb(n9873), .dout(n9875));
  jnot g09812(.din(n9875), .dout(n9876));
  jand g09813(.dina(n9876), .dinb(n9537), .dout(n9877));
  jnot g09814(.din(n9877), .dout(n9878));
  jxor g09815(.dina(n9525), .dinb(n9517), .dout(n9879));
  jand g09816(.dina(n9879), .dinb(n9878), .dout(n9880));
  jnot g09817(.din(n9880), .dout(n9881));
  jand g09818(.dina(n9881), .dinb(n9526), .dout(n9882));
  jnot g09819(.din(n9882), .dout(n9883));
  jxor g09820(.dina(n9463), .dinb(n9462), .dout(n9884));
  jand g09821(.dina(n9884), .dinb(n9883), .dout(n9885));
  jand g09822(.dina(n7890), .dinb(n4043), .dout(n9886));
  jand g09823(.dina(n8441), .dinb(n1076), .dout(n9887));
  jand g09824(.dina(n8154), .dinb(n1213), .dout(n9888));
  jand g09825(.dina(n7888), .dinb(n1343), .dout(n9889));
  jor  g09826(.dina(n9889), .dinb(n9888), .dout(n9890));
  jor  g09827(.dina(n9890), .dinb(n9887), .dout(n9891));
  jor  g09828(.dina(n9891), .dinb(n9886), .dout(n9892));
  jxor g09829(.dina(n9892), .dinb(n5833), .dout(n9893));
  jnot g09830(.din(n9893), .dout(n9894));
  jxor g09831(.dina(n9884), .dinb(n9883), .dout(n9895));
  jand g09832(.dina(n9895), .dinb(n9894), .dout(n9896));
  jor  g09833(.dina(n9896), .dinb(n9885), .dout(n9897));
  jxor g09834(.dina(n9478), .dinb(n9470), .dout(n9898));
  jand g09835(.dina(n9898), .dinb(n9897), .dout(n9899));
  jnot g09836(.din(n9899), .dout(n9900));
  jxor g09837(.dina(n9898), .dinb(n9897), .dout(n9901));
  jnot g09838(.din(n9901), .dout(n9902));
  jand g09839(.dina(n8771), .dinb(n4446), .dout(n9903));
  jand g09840(.dina(n9491), .dinb(n4451), .dout(n9904));
  jand g09841(.dina(n9126), .dinb(n4358), .dout(n9905));
  jand g09842(.dina(n8769), .dinb(n3853), .dout(n9906));
  jor  g09843(.dina(n9906), .dinb(n9905), .dout(n9907));
  jor  g09844(.dina(n9907), .dinb(n9904), .dout(n9908));
  jor  g09845(.dina(n9908), .dinb(n9903), .dout(n9909));
  jxor g09846(.dina(n9909), .dinb(n6039), .dout(n9910));
  jor  g09847(.dina(n9910), .dinb(n9902), .dout(n9911));
  jand g09848(.dina(n9911), .dinb(n9900), .dout(n9912));
  jnot g09849(.din(n65), .dout(n9913));
  jxor g09850(.dina(\a[4] ), .dinb(\a[3] ), .dout(n9914));
  jnot g09851(.din(n9914), .dout(n9915));
  jand g09852(.dina(n9915), .dinb(n9913), .dout(n9916));
  jand g09853(.dina(n9916), .dinb(n66), .dout(n9917));
  jnot g09854(.din(n9917), .dout(n9918));
  jnot g09855(.din(n67), .dout(n9919));
  jor  g09856(.dina(n4728), .dinb(n9919), .dout(n9920));
  jand g09857(.dina(n9920), .dinb(n9918), .dout(n9921));
  jor  g09858(.dina(n9921), .dinb(n4630), .dout(n9922));
  jxor g09859(.dina(n9922), .dinb(\a[5] ), .dout(n9923));
  jor  g09860(.dina(n9923), .dinb(n9912), .dout(n9924));
  jxor g09861(.dina(n9923), .dinb(n9912), .dout(n9925));
  jxor g09862(.dina(n9496), .dinb(n9486), .dout(n9926));
  jand g09863(.dina(n9926), .dinb(n9925), .dout(n9927));
  jnot g09864(.din(n9927), .dout(n9928));
  jand g09865(.dina(n9928), .dinb(n9924), .dout(n9929));
  jnot g09866(.din(n9929), .dout(n9930));
  jxor g09867(.dina(n9509), .dinb(n9508), .dout(n9931));
  jand g09868(.dina(n9931), .dinb(n9930), .dout(n9932));
  jand g09869(.dina(n7890), .dinb(n4772), .dout(n9933));
  jand g09870(.dina(n8441), .dinb(n1213), .dout(n9934));
  jand g09871(.dina(n8154), .dinb(n1343), .dout(n9935));
  jand g09872(.dina(n7888), .dinb(n1445), .dout(n9936));
  jor  g09873(.dina(n9936), .dinb(n9935), .dout(n9937));
  jor  g09874(.dina(n9937), .dinb(n9934), .dout(n9938));
  jor  g09875(.dina(n9938), .dinb(n9933), .dout(n9939));
  jxor g09876(.dina(n9939), .dinb(n5833), .dout(n9940));
  jnot g09877(.din(n9940), .dout(n9941));
  jxor g09878(.dina(n9879), .dinb(n9878), .dout(n9942));
  jand g09879(.dina(n9942), .dinb(n9941), .dout(n9943));
  jand g09880(.dina(n7890), .dinb(n4258), .dout(n9944));
  jand g09881(.dina(n8441), .dinb(n1343), .dout(n9945));
  jand g09882(.dina(n8154), .dinb(n1445), .dout(n9946));
  jand g09883(.dina(n7888), .dinb(n1560), .dout(n9947));
  jor  g09884(.dina(n9947), .dinb(n9946), .dout(n9948));
  jor  g09885(.dina(n9948), .dinb(n9945), .dout(n9949));
  jor  g09886(.dina(n9949), .dinb(n9944), .dout(n9950));
  jxor g09887(.dina(n9950), .dinb(n5833), .dout(n9951));
  jnot g09888(.din(n9951), .dout(n9952));
  jxor g09889(.dina(n9874), .dinb(n9873), .dout(n9953));
  jand g09890(.dina(n9953), .dinb(n9952), .dout(n9954));
  jand g09891(.dina(n7890), .dinb(n4866), .dout(n9955));
  jand g09892(.dina(n8441), .dinb(n1445), .dout(n9956));
  jand g09893(.dina(n8154), .dinb(n1560), .dout(n9957));
  jand g09894(.dina(n7888), .dinb(n1624), .dout(n9958));
  jor  g09895(.dina(n9958), .dinb(n9957), .dout(n9959));
  jor  g09896(.dina(n9959), .dinb(n9956), .dout(n9960));
  jor  g09897(.dina(n9960), .dinb(n9955), .dout(n9961));
  jxor g09898(.dina(n9961), .dinb(n5833), .dout(n9962));
  jnot g09899(.din(n9962), .dout(n9963));
  jxor g09900(.dina(n9869), .dinb(n9868), .dout(n9964));
  jand g09901(.dina(n9964), .dinb(n9963), .dout(n9965));
  jand g09902(.dina(n7890), .dinb(n4849), .dout(n9966));
  jand g09903(.dina(n8441), .dinb(n1560), .dout(n9967));
  jand g09904(.dina(n8154), .dinb(n1624), .dout(n9968));
  jand g09905(.dina(n7888), .dinb(n1776), .dout(n9969));
  jor  g09906(.dina(n9969), .dinb(n9968), .dout(n9970));
  jor  g09907(.dina(n9970), .dinb(n9967), .dout(n9971));
  jor  g09908(.dina(n9971), .dinb(n9966), .dout(n9972));
  jxor g09909(.dina(n9972), .dinb(n5833), .dout(n9973));
  jnot g09910(.din(n9973), .dout(n9974));
  jxor g09911(.dina(n9864), .dinb(n9863), .dout(n9975));
  jand g09912(.dina(n9975), .dinb(n9974), .dout(n9976));
  jand g09913(.dina(n7890), .dinb(n5075), .dout(n9977));
  jand g09914(.dina(n8441), .dinb(n1624), .dout(n9978));
  jand g09915(.dina(n8154), .dinb(n1776), .dout(n9979));
  jand g09916(.dina(n7888), .dinb(n1862), .dout(n9980));
  jor  g09917(.dina(n9980), .dinb(n9979), .dout(n9981));
  jor  g09918(.dina(n9981), .dinb(n9978), .dout(n9982));
  jor  g09919(.dina(n9982), .dinb(n9977), .dout(n9983));
  jxor g09920(.dina(n9983), .dinb(n5833), .dout(n9984));
  jnot g09921(.din(n9984), .dout(n9985));
  jxor g09922(.dina(n9859), .dinb(n9858), .dout(n9986));
  jand g09923(.dina(n9986), .dinb(n9985), .dout(n9987));
  jand g09924(.dina(n7890), .dinb(n5092), .dout(n9988));
  jand g09925(.dina(n8441), .dinb(n1776), .dout(n9989));
  jand g09926(.dina(n8154), .dinb(n1862), .dout(n9990));
  jand g09927(.dina(n7888), .dinb(n1956), .dout(n9991));
  jor  g09928(.dina(n9991), .dinb(n9990), .dout(n9992));
  jor  g09929(.dina(n9992), .dinb(n9989), .dout(n9993));
  jor  g09930(.dina(n9993), .dinb(n9988), .dout(n9994));
  jxor g09931(.dina(n9994), .dinb(n5833), .dout(n9995));
  jnot g09932(.din(n9995), .dout(n9996));
  jxor g09933(.dina(n9854), .dinb(n9853), .dout(n9997));
  jand g09934(.dina(n9997), .dinb(n9996), .dout(n9998));
  jand g09935(.dina(n7890), .dinb(n5440), .dout(n9999));
  jand g09936(.dina(n8154), .dinb(n1956), .dout(n10000));
  jand g09937(.dina(n8441), .dinb(n1862), .dout(n10001));
  jand g09938(.dina(n7888), .dinb(n2067), .dout(n10002));
  jor  g09939(.dina(n10002), .dinb(n10001), .dout(n10003));
  jor  g09940(.dina(n10003), .dinb(n10000), .dout(n10004));
  jor  g09941(.dina(n10004), .dinb(n9999), .dout(n10005));
  jxor g09942(.dina(n10005), .dinb(n5833), .dout(n10006));
  jnot g09943(.din(n10006), .dout(n10007));
  jxor g09944(.dina(n9849), .dinb(n9848), .dout(n10008));
  jand g09945(.dina(n10008), .dinb(n10007), .dout(n10009));
  jxor g09946(.dina(n9846), .dinb(n9845), .dout(n10010));
  jnot g09947(.din(n10010), .dout(n10011));
  jand g09948(.dina(n7890), .dinb(n5303), .dout(n10012));
  jand g09949(.dina(n7888), .dinb(n2128), .dout(n10013));
  jand g09950(.dina(n8154), .dinb(n2067), .dout(n10014));
  jand g09951(.dina(n8441), .dinb(n1956), .dout(n10015));
  jor  g09952(.dina(n10015), .dinb(n10014), .dout(n10016));
  jor  g09953(.dina(n10016), .dinb(n10013), .dout(n10017));
  jor  g09954(.dina(n10017), .dinb(n10012), .dout(n10018));
  jxor g09955(.dina(n10018), .dinb(n5833), .dout(n10019));
  jor  g09956(.dina(n10019), .dinb(n10011), .dout(n10020));
  jxor g09957(.dina(n9843), .dinb(n9842), .dout(n10021));
  jnot g09958(.din(n10021), .dout(n10022));
  jand g09959(.dina(n7890), .dinb(n5624), .dout(n10023));
  jand g09960(.dina(n7888), .dinb(n2237), .dout(n10024));
  jand g09961(.dina(n8154), .dinb(n2128), .dout(n10025));
  jand g09962(.dina(n8441), .dinb(n2067), .dout(n10026));
  jor  g09963(.dina(n10026), .dinb(n10025), .dout(n10027));
  jor  g09964(.dina(n10027), .dinb(n10024), .dout(n10028));
  jor  g09965(.dina(n10028), .dinb(n10023), .dout(n10029));
  jxor g09966(.dina(n10029), .dinb(n5833), .dout(n10030));
  jor  g09967(.dina(n10030), .dinb(n10022), .dout(n10031));
  jand g09968(.dina(n7890), .dinb(n5607), .dout(n10032));
  jand g09969(.dina(n8154), .dinb(n2237), .dout(n10033));
  jand g09970(.dina(n7888), .dinb(n2343), .dout(n10034));
  jand g09971(.dina(n8441), .dinb(n2128), .dout(n10035));
  jor  g09972(.dina(n10035), .dinb(n10034), .dout(n10036));
  jor  g09973(.dina(n10036), .dinb(n10033), .dout(n10037));
  jor  g09974(.dina(n10037), .dinb(n10032), .dout(n10038));
  jxor g09975(.dina(n10038), .dinb(n5833), .dout(n10039));
  jnot g09976(.din(n10039), .dout(n10040));
  jxor g09977(.dina(n9838), .dinb(n9837), .dout(n10041));
  jand g09978(.dina(n10041), .dinb(n10040), .dout(n10042));
  jand g09979(.dina(n7890), .dinb(n5844), .dout(n10043));
  jand g09980(.dina(n7888), .dinb(n2411), .dout(n10044));
  jand g09981(.dina(n8441), .dinb(n2237), .dout(n10045));
  jand g09982(.dina(n8154), .dinb(n2343), .dout(n10046));
  jor  g09983(.dina(n10046), .dinb(n10045), .dout(n10047));
  jor  g09984(.dina(n10047), .dinb(n10044), .dout(n10048));
  jor  g09985(.dina(n10048), .dinb(n10043), .dout(n10049));
  jxor g09986(.dina(n10049), .dinb(n5833), .dout(n10050));
  jnot g09987(.din(n10050), .dout(n10051));
  jxor g09988(.dina(n9833), .dinb(n9832), .dout(n10052));
  jand g09989(.dina(n10052), .dinb(n10051), .dout(n10053));
  jand g09990(.dina(n7890), .dinb(n5861), .dout(n10054));
  jand g09991(.dina(n8154), .dinb(n2411), .dout(n10055));
  jand g09992(.dina(n8441), .dinb(n2343), .dout(n10056));
  jand g09993(.dina(n7888), .dinb(n2497), .dout(n10057));
  jor  g09994(.dina(n10057), .dinb(n10056), .dout(n10058));
  jor  g09995(.dina(n10058), .dinb(n10055), .dout(n10059));
  jor  g09996(.dina(n10059), .dinb(n10054), .dout(n10060));
  jxor g09997(.dina(n10060), .dinb(n5833), .dout(n10061));
  jnot g09998(.din(n10061), .dout(n10062));
  jxor g09999(.dina(n9828), .dinb(n9827), .dout(n10063));
  jand g10000(.dina(n10063), .dinb(n10062), .dout(n10064));
  jxor g10001(.dina(n9825), .dinb(n9824), .dout(n10065));
  jnot g10002(.din(n10065), .dout(n10066));
  jand g10003(.dina(n7890), .dinb(n6247), .dout(n10067));
  jand g10004(.dina(n8441), .dinb(n2411), .dout(n10068));
  jand g10005(.dina(n7888), .dinb(n2602), .dout(n10069));
  jand g10006(.dina(n8154), .dinb(n2497), .dout(n10070));
  jor  g10007(.dina(n10070), .dinb(n10069), .dout(n10071));
  jor  g10008(.dina(n10071), .dinb(n10068), .dout(n10072));
  jor  g10009(.dina(n10072), .dinb(n10067), .dout(n10073));
  jxor g10010(.dina(n10073), .dinb(n5833), .dout(n10074));
  jor  g10011(.dina(n10074), .dinb(n10066), .dout(n10075));
  jxor g10012(.dina(n9822), .dinb(n9821), .dout(n10076));
  jnot g10013(.din(n10076), .dout(n10077));
  jand g10014(.dina(n7890), .dinb(n6050), .dout(n10078));
  jand g10015(.dina(n8154), .dinb(n2602), .dout(n10079));
  jand g10016(.dina(n7888), .dinb(n2695), .dout(n10080));
  jand g10017(.dina(n8441), .dinb(n2497), .dout(n10081));
  jor  g10018(.dina(n10081), .dinb(n10080), .dout(n10082));
  jor  g10019(.dina(n10082), .dinb(n10079), .dout(n10083));
  jor  g10020(.dina(n10083), .dinb(n10078), .dout(n10084));
  jxor g10021(.dina(n10084), .dinb(n5833), .dout(n10085));
  jor  g10022(.dina(n10085), .dinb(n10077), .dout(n10086));
  jxor g10023(.dina(n9819), .dinb(n9818), .dout(n10087));
  jnot g10024(.din(n10087), .dout(n10088));
  jor  g10025(.dina(n7891), .dinb(n6464), .dout(n10089));
  jor  g10026(.dina(n8440), .dinb(n2601), .dout(n10090));
  jor  g10027(.dina(n8155), .dinb(n2694), .dout(n10091));
  jor  g10028(.dina(n7889), .dinb(n2731), .dout(n10092));
  jand g10029(.dina(n10092), .dinb(n10091), .dout(n10093));
  jand g10030(.dina(n10093), .dinb(n10090), .dout(n10094));
  jand g10031(.dina(n10094), .dinb(n10089), .dout(n10095));
  jxor g10032(.dina(n10095), .dinb(\a[11] ), .dout(n10096));
  jor  g10033(.dina(n10096), .dinb(n10088), .dout(n10097));
  jand g10034(.dina(n7890), .dinb(n6591), .dout(n10098));
  jand g10035(.dina(n8441), .dinb(n2695), .dout(n10099));
  jand g10036(.dina(n7888), .dinb(n2808), .dout(n10100));
  jand g10037(.dina(n8154), .dinb(n2732), .dout(n10101));
  jor  g10038(.dina(n10101), .dinb(n10100), .dout(n10102));
  jor  g10039(.dina(n10102), .dinb(n10099), .dout(n10103));
  jor  g10040(.dina(n10103), .dinb(n10098), .dout(n10104));
  jxor g10041(.dina(n10104), .dinb(n5833), .dout(n10105));
  jnot g10042(.din(n10105), .dout(n10106));
  jxor g10043(.dina(n9814), .dinb(n9813), .dout(n10107));
  jand g10044(.dina(n10107), .dinb(n10106), .dout(n10108));
  jand g10045(.dina(n7890), .dinb(n6439), .dout(n10109));
  jand g10046(.dina(n8154), .dinb(n2808), .dout(n10110));
  jand g10047(.dina(n8441), .dinb(n2732), .dout(n10111));
  jand g10048(.dina(n7888), .dinb(n2867), .dout(n10112));
  jor  g10049(.dina(n10112), .dinb(n10111), .dout(n10113));
  jor  g10050(.dina(n10113), .dinb(n10110), .dout(n10114));
  jor  g10051(.dina(n10114), .dinb(n10109), .dout(n10115));
  jxor g10052(.dina(n10115), .dinb(n5833), .dout(n10116));
  jnot g10053(.din(n10116), .dout(n10117));
  jxor g10054(.dina(n9809), .dinb(n9808), .dout(n10118));
  jand g10055(.dina(n10118), .dinb(n10117), .dout(n10119));
  jand g10056(.dina(n7890), .dinb(n6706), .dout(n10120));
  jand g10057(.dina(n8441), .dinb(n2808), .dout(n10121));
  jand g10058(.dina(n7888), .dinb(n2954), .dout(n10122));
  jand g10059(.dina(n8154), .dinb(n2867), .dout(n10123));
  jor  g10060(.dina(n10123), .dinb(n10122), .dout(n10124));
  jor  g10061(.dina(n10124), .dinb(n10121), .dout(n10125));
  jor  g10062(.dina(n10125), .dinb(n10120), .dout(n10126));
  jxor g10063(.dina(n10126), .dinb(n5833), .dout(n10127));
  jnot g10064(.din(n10127), .dout(n10128));
  jxor g10065(.dina(n9804), .dinb(n9803), .dout(n10129));
  jand g10066(.dina(n10129), .dinb(n10128), .dout(n10130));
  jxor g10067(.dina(n9801), .dinb(n9800), .dout(n10131));
  jnot g10068(.din(n10131), .dout(n10132));
  jor  g10069(.dina(n7891), .dinb(n6976), .dout(n10133));
  jor  g10070(.dina(n8155), .dinb(n2953), .dout(n10134));
  jor  g10071(.dina(n7889), .dinb(n2990), .dout(n10135));
  jor  g10072(.dina(n8440), .dinb(n2866), .dout(n10136));
  jand g10073(.dina(n10136), .dinb(n10135), .dout(n10137));
  jand g10074(.dina(n10137), .dinb(n10134), .dout(n10138));
  jand g10075(.dina(n10138), .dinb(n10133), .dout(n10139));
  jxor g10076(.dina(n10139), .dinb(\a[11] ), .dout(n10140));
  jor  g10077(.dina(n10140), .dinb(n10132), .dout(n10141));
  jxor g10078(.dina(n9798), .dinb(n9797), .dout(n10142));
  jnot g10079(.din(n10142), .dout(n10143));
  jor  g10080(.dina(n7891), .dinb(n6988), .dout(n10144));
  jor  g10081(.dina(n7889), .dinb(n3085), .dout(n10145));
  jor  g10082(.dina(n8440), .dinb(n2953), .dout(n10146));
  jor  g10083(.dina(n8155), .dinb(n2990), .dout(n10147));
  jand g10084(.dina(n10147), .dinb(n10146), .dout(n10148));
  jand g10085(.dina(n10148), .dinb(n10145), .dout(n10149));
  jand g10086(.dina(n10149), .dinb(n10144), .dout(n10150));
  jxor g10087(.dina(n10150), .dinb(\a[11] ), .dout(n10151));
  jor  g10088(.dina(n10151), .dinb(n10143), .dout(n10152));
  jxor g10089(.dina(n9795), .dinb(n9794), .dout(n10153));
  jnot g10090(.din(n10153), .dout(n10154));
  jor  g10091(.dina(n7891), .dinb(n6681), .dout(n10155));
  jor  g10092(.dina(n8155), .dinb(n3085), .dout(n10156));
  jor  g10093(.dina(n8440), .dinb(n2990), .dout(n10157));
  jor  g10094(.dina(n7889), .dinb(n3182), .dout(n10158));
  jand g10095(.dina(n10158), .dinb(n10157), .dout(n10159));
  jand g10096(.dina(n10159), .dinb(n10156), .dout(n10160));
  jand g10097(.dina(n10160), .dinb(n10155), .dout(n10161));
  jxor g10098(.dina(n10161), .dinb(\a[11] ), .dout(n10162));
  jor  g10099(.dina(n10162), .dinb(n10154), .dout(n10163));
  jor  g10100(.dina(n7891), .dinb(n7031), .dout(n10164));
  jor  g10101(.dina(n8440), .dinb(n3085), .dout(n10165));
  jor  g10102(.dina(n7889), .dinb(n7962), .dout(n10166));
  jor  g10103(.dina(n8155), .dinb(n3182), .dout(n10167));
  jand g10104(.dina(n10167), .dinb(n10166), .dout(n10168));
  jand g10105(.dina(n10168), .dinb(n10165), .dout(n10169));
  jand g10106(.dina(n10169), .dinb(n10164), .dout(n10170));
  jxor g10107(.dina(n10170), .dinb(\a[11] ), .dout(n10171));
  jnot g10108(.din(n10171), .dout(n10172));
  jxor g10109(.dina(n9792), .dinb(n9791), .dout(n10173));
  jand g10110(.dina(n10173), .dinb(n10172), .dout(n10174));
  jor  g10111(.dina(n7891), .dinb(n7076), .dout(n10175));
  jor  g10112(.dina(n8155), .dinb(n7962), .dout(n10176));
  jor  g10113(.dina(n8440), .dinb(n3182), .dout(n10177));
  jor  g10114(.dina(n7889), .dinb(n3684), .dout(n10178));
  jand g10115(.dina(n10178), .dinb(n10177), .dout(n10179));
  jand g10116(.dina(n10179), .dinb(n10176), .dout(n10180));
  jand g10117(.dina(n10180), .dinb(n10175), .dout(n10181));
  jxor g10118(.dina(n10181), .dinb(\a[11] ), .dout(n10182));
  jnot g10119(.din(n10182), .dout(n10183));
  jxor g10120(.dina(n9789), .dinb(n9788), .dout(n10184));
  jand g10121(.dina(n10184), .dinb(n10183), .dout(n10185));
  jor  g10122(.dina(n7891), .dinb(n7131), .dout(n10186));
  jor  g10123(.dina(n8440), .dinb(n7962), .dout(n10187));
  jor  g10124(.dina(n7889), .dinb(n3414), .dout(n10188));
  jor  g10125(.dina(n8155), .dinb(n3684), .dout(n10189));
  jand g10126(.dina(n10189), .dinb(n10188), .dout(n10190));
  jand g10127(.dina(n10190), .dinb(n10187), .dout(n10191));
  jand g10128(.dina(n10191), .dinb(n10186), .dout(n10192));
  jxor g10129(.dina(n10192), .dinb(\a[11] ), .dout(n10193));
  jnot g10130(.din(n10193), .dout(n10194));
  jor  g10131(.dina(n9769), .dinb(n5292), .dout(n10195));
  jxor g10132(.dina(n10195), .dinb(n9777), .dout(n10196));
  jand g10133(.dina(n10196), .dinb(n10194), .dout(n10197));
  jor  g10134(.dina(n7891), .dinb(n7177), .dout(n10198));
  jor  g10135(.dina(n7889), .dinb(n3516), .dout(n10199));
  jor  g10136(.dina(n8440), .dinb(n3684), .dout(n10200));
  jor  g10137(.dina(n8155), .dinb(n3414), .dout(n10201));
  jand g10138(.dina(n10201), .dinb(n10200), .dout(n10202));
  jand g10139(.dina(n10202), .dinb(n10199), .dout(n10203));
  jand g10140(.dina(n10203), .dinb(n10198), .dout(n10204));
  jxor g10141(.dina(n10204), .dinb(\a[11] ), .dout(n10205));
  jnot g10142(.din(n10205), .dout(n10206));
  jand g10143(.dina(n9766), .dinb(\a[14] ), .dout(n10207));
  jxor g10144(.dina(n10207), .dinb(n9764), .dout(n10208));
  jand g10145(.dina(n10208), .dinb(n10206), .dout(n10209));
  jand g10146(.dina(n8004), .dinb(n7890), .dout(n10210));
  jand g10147(.dina(n8154), .dinb(n7411), .dout(n10211));
  jand g10148(.dina(n8441), .dinb(n7405), .dout(n10212));
  jor  g10149(.dina(n10212), .dinb(n10211), .dout(n10213));
  jor  g10150(.dina(n10213), .dinb(n10210), .dout(n10214));
  jnot g10151(.din(n10214), .dout(n10215));
  jand g10152(.dina(n7884), .dinb(n7411), .dout(n10216));
  jnot g10153(.din(n10216), .dout(n10217));
  jand g10154(.dina(n10217), .dinb(\a[11] ), .dout(n10218));
  jand g10155(.dina(n10218), .dinb(n10215), .dout(n10219));
  jand g10156(.dina(n7890), .dinb(n7407), .dout(n10220));
  jand g10157(.dina(n8441), .dinb(n7326), .dout(n10221));
  jand g10158(.dina(n7888), .dinb(n7411), .dout(n10222));
  jand g10159(.dina(n8154), .dinb(n7405), .dout(n10223));
  jor  g10160(.dina(n10223), .dinb(n10222), .dout(n10224));
  jor  g10161(.dina(n10224), .dinb(n10221), .dout(n10225));
  jor  g10162(.dina(n10225), .dinb(n10220), .dout(n10226));
  jnot g10163(.din(n10226), .dout(n10227));
  jand g10164(.dina(n10227), .dinb(n10219), .dout(n10228));
  jand g10165(.dina(n10228), .dinb(n9766), .dout(n10229));
  jor  g10166(.dina(n7891), .dinb(n7466), .dout(n10230));
  jor  g10167(.dina(n8155), .dinb(n3516), .dout(n10231));
  jor  g10168(.dina(n8440), .dinb(n3414), .dout(n10232));
  jor  g10169(.dina(n7889), .dinb(n3677), .dout(n10233));
  jand g10170(.dina(n10233), .dinb(n10232), .dout(n10234));
  jand g10171(.dina(n10234), .dinb(n10231), .dout(n10235));
  jand g10172(.dina(n10235), .dinb(n10230), .dout(n10236));
  jxor g10173(.dina(n10236), .dinb(\a[11] ), .dout(n10237));
  jnot g10174(.din(n10237), .dout(n10238));
  jxor g10175(.dina(n10228), .dinb(n9766), .dout(n10239));
  jand g10176(.dina(n10239), .dinb(n10238), .dout(n10240));
  jor  g10177(.dina(n10240), .dinb(n10229), .dout(n10241));
  jxor g10178(.dina(n10208), .dinb(n10206), .dout(n10242));
  jand g10179(.dina(n10242), .dinb(n10241), .dout(n10243));
  jor  g10180(.dina(n10243), .dinb(n10209), .dout(n10244));
  jxor g10181(.dina(n10196), .dinb(n10194), .dout(n10245));
  jand g10182(.dina(n10245), .dinb(n10244), .dout(n10246));
  jor  g10183(.dina(n10246), .dinb(n10197), .dout(n10247));
  jxor g10184(.dina(n10184), .dinb(n10183), .dout(n10248));
  jand g10185(.dina(n10248), .dinb(n10247), .dout(n10249));
  jor  g10186(.dina(n10249), .dinb(n10185), .dout(n10250));
  jxor g10187(.dina(n10173), .dinb(n10172), .dout(n10251));
  jand g10188(.dina(n10251), .dinb(n10250), .dout(n10252));
  jor  g10189(.dina(n10252), .dinb(n10174), .dout(n10253));
  jxor g10190(.dina(n10162), .dinb(n10154), .dout(n10254));
  jand g10191(.dina(n10254), .dinb(n10253), .dout(n10255));
  jnot g10192(.din(n10255), .dout(n10256));
  jand g10193(.dina(n10256), .dinb(n10163), .dout(n10257));
  jnot g10194(.din(n10257), .dout(n10258));
  jxor g10195(.dina(n10151), .dinb(n10143), .dout(n10259));
  jand g10196(.dina(n10259), .dinb(n10258), .dout(n10260));
  jnot g10197(.din(n10260), .dout(n10261));
  jand g10198(.dina(n10261), .dinb(n10152), .dout(n10262));
  jnot g10199(.din(n10262), .dout(n10263));
  jxor g10200(.dina(n10140), .dinb(n10132), .dout(n10264));
  jand g10201(.dina(n10264), .dinb(n10263), .dout(n10265));
  jnot g10202(.din(n10265), .dout(n10266));
  jand g10203(.dina(n10266), .dinb(n10141), .dout(n10267));
  jnot g10204(.din(n10267), .dout(n10268));
  jxor g10205(.dina(n10129), .dinb(n10128), .dout(n10269));
  jand g10206(.dina(n10269), .dinb(n10268), .dout(n10270));
  jor  g10207(.dina(n10270), .dinb(n10130), .dout(n10271));
  jxor g10208(.dina(n10118), .dinb(n10117), .dout(n10272));
  jand g10209(.dina(n10272), .dinb(n10271), .dout(n10273));
  jor  g10210(.dina(n10273), .dinb(n10119), .dout(n10274));
  jxor g10211(.dina(n10107), .dinb(n10106), .dout(n10275));
  jand g10212(.dina(n10275), .dinb(n10274), .dout(n10276));
  jor  g10213(.dina(n10276), .dinb(n10108), .dout(n10277));
  jxor g10214(.dina(n10096), .dinb(n10088), .dout(n10278));
  jand g10215(.dina(n10278), .dinb(n10277), .dout(n10279));
  jnot g10216(.din(n10279), .dout(n10280));
  jand g10217(.dina(n10280), .dinb(n10097), .dout(n10281));
  jnot g10218(.din(n10281), .dout(n10282));
  jxor g10219(.dina(n10085), .dinb(n10077), .dout(n10283));
  jand g10220(.dina(n10283), .dinb(n10282), .dout(n10284));
  jnot g10221(.din(n10284), .dout(n10285));
  jand g10222(.dina(n10285), .dinb(n10086), .dout(n10286));
  jnot g10223(.din(n10286), .dout(n10287));
  jxor g10224(.dina(n10074), .dinb(n10066), .dout(n10288));
  jand g10225(.dina(n10288), .dinb(n10287), .dout(n10289));
  jnot g10226(.din(n10289), .dout(n10290));
  jand g10227(.dina(n10290), .dinb(n10075), .dout(n10291));
  jnot g10228(.din(n10291), .dout(n10292));
  jxor g10229(.dina(n10063), .dinb(n10062), .dout(n10293));
  jand g10230(.dina(n10293), .dinb(n10292), .dout(n10294));
  jor  g10231(.dina(n10294), .dinb(n10064), .dout(n10295));
  jxor g10232(.dina(n10052), .dinb(n10051), .dout(n10296));
  jand g10233(.dina(n10296), .dinb(n10295), .dout(n10297));
  jor  g10234(.dina(n10297), .dinb(n10053), .dout(n10298));
  jxor g10235(.dina(n10041), .dinb(n10040), .dout(n10299));
  jand g10236(.dina(n10299), .dinb(n10298), .dout(n10300));
  jor  g10237(.dina(n10300), .dinb(n10042), .dout(n10301));
  jxor g10238(.dina(n10030), .dinb(n10022), .dout(n10302));
  jand g10239(.dina(n10302), .dinb(n10301), .dout(n10303));
  jnot g10240(.din(n10303), .dout(n10304));
  jand g10241(.dina(n10304), .dinb(n10031), .dout(n10305));
  jnot g10242(.din(n10305), .dout(n10306));
  jxor g10243(.dina(n10019), .dinb(n10011), .dout(n10307));
  jand g10244(.dina(n10307), .dinb(n10306), .dout(n10308));
  jnot g10245(.din(n10308), .dout(n10309));
  jand g10246(.dina(n10309), .dinb(n10020), .dout(n10310));
  jnot g10247(.din(n10310), .dout(n10311));
  jxor g10248(.dina(n10008), .dinb(n10007), .dout(n10312));
  jand g10249(.dina(n10312), .dinb(n10311), .dout(n10313));
  jor  g10250(.dina(n10313), .dinb(n10009), .dout(n10314));
  jxor g10251(.dina(n9997), .dinb(n9996), .dout(n10315));
  jand g10252(.dina(n10315), .dinb(n10314), .dout(n10316));
  jor  g10253(.dina(n10316), .dinb(n9998), .dout(n10317));
  jxor g10254(.dina(n9986), .dinb(n9985), .dout(n10318));
  jand g10255(.dina(n10318), .dinb(n10317), .dout(n10319));
  jor  g10256(.dina(n10319), .dinb(n9987), .dout(n10320));
  jxor g10257(.dina(n9975), .dinb(n9974), .dout(n10321));
  jand g10258(.dina(n10321), .dinb(n10320), .dout(n10322));
  jor  g10259(.dina(n10322), .dinb(n9976), .dout(n10323));
  jxor g10260(.dina(n9964), .dinb(n9963), .dout(n10324));
  jand g10261(.dina(n10324), .dinb(n10323), .dout(n10325));
  jor  g10262(.dina(n10325), .dinb(n9965), .dout(n10326));
  jxor g10263(.dina(n9953), .dinb(n9952), .dout(n10327));
  jand g10264(.dina(n10327), .dinb(n10326), .dout(n10328));
  jor  g10265(.dina(n10328), .dinb(n9954), .dout(n10329));
  jxor g10266(.dina(n9942), .dinb(n9941), .dout(n10330));
  jand g10267(.dina(n10330), .dinb(n10329), .dout(n10331));
  jor  g10268(.dina(n10331), .dinb(n9943), .dout(n10332));
  jxor g10269(.dina(n9895), .dinb(n9894), .dout(n10333));
  jand g10270(.dina(n10333), .dinb(n10332), .dout(n10334));
  jand g10271(.dina(n8771), .dinb(n4545), .dout(n10335));
  jand g10272(.dina(n9126), .dinb(n3853), .dout(n10336));
  jand g10273(.dina(n9491), .dinb(n4358), .dout(n10337));
  jand g10274(.dina(n8769), .dinb(n922), .dout(n10338));
  jor  g10275(.dina(n10338), .dinb(n10337), .dout(n10339));
  jor  g10276(.dina(n10339), .dinb(n10336), .dout(n10340));
  jor  g10277(.dina(n10340), .dinb(n10335), .dout(n10341));
  jxor g10278(.dina(n10341), .dinb(n6039), .dout(n10342));
  jnot g10279(.din(n10342), .dout(n10343));
  jxor g10280(.dina(n10333), .dinb(n10332), .dout(n10344));
  jand g10281(.dina(n10344), .dinb(n10343), .dout(n10345));
  jor  g10282(.dina(n10345), .dinb(n10334), .dout(n10346));
  jnot g10283(.din(n10346), .dout(n10347));
  jor  g10284(.dina(n4731), .dinb(n9919), .dout(n10348));
  jor  g10285(.dina(n9918), .dinb(n4597), .dout(n10349));
  jand g10286(.dina(n9914), .dinb(n9913), .dout(n10350));
  jnot g10287(.din(n10350), .dout(n10351));
  jor  g10288(.dina(n10351), .dinb(n4630), .dout(n10352));
  jand g10289(.dina(n10352), .dinb(n10349), .dout(n10353));
  jand g10290(.dina(n10353), .dinb(n10348), .dout(n10354));
  jxor g10291(.dina(n10354), .dinb(\a[5] ), .dout(n10355));
  jor  g10292(.dina(n10355), .dinb(n10347), .dout(n10356));
  jxor g10293(.dina(n10355), .dinb(n10347), .dout(n10357));
  jxor g10294(.dina(n9910), .dinb(n9902), .dout(n10358));
  jand g10295(.dina(n10358), .dinb(n10357), .dout(n10359));
  jnot g10296(.din(n10359), .dout(n10360));
  jand g10297(.dina(n10360), .dinb(n10356), .dout(n10361));
  jnot g10298(.din(n10361), .dout(n10362));
  jxor g10299(.dina(n9926), .dinb(n9925), .dout(n10363));
  jand g10300(.dina(n10363), .dinb(n10362), .dout(n10364));
  jnot g10301(.din(n10364), .dout(n10365));
  jxor g10302(.dina(n10363), .dinb(n10362), .dout(n10366));
  jnot g10303(.din(n10366), .dout(n10367));
  jxor g10304(.dina(n10330), .dinb(n10329), .dout(n10368));
  jnot g10305(.din(n10368), .dout(n10369));
  jand g10306(.dina(n8771), .dinb(n3848), .dout(n10370));
  jand g10307(.dina(n8769), .dinb(n1076), .dout(n10371));
  jand g10308(.dina(n9126), .dinb(n922), .dout(n10372));
  jand g10309(.dina(n9491), .dinb(n3853), .dout(n10373));
  jor  g10310(.dina(n10373), .dinb(n10372), .dout(n10374));
  jor  g10311(.dina(n10374), .dinb(n10371), .dout(n10375));
  jor  g10312(.dina(n10375), .dinb(n10370), .dout(n10376));
  jxor g10313(.dina(n10376), .dinb(n6039), .dout(n10377));
  jor  g10314(.dina(n10377), .dinb(n10369), .dout(n10378));
  jxor g10315(.dina(n10327), .dinb(n10326), .dout(n10379));
  jnot g10316(.din(n10379), .dout(n10380));
  jand g10317(.dina(n8771), .dinb(n4026), .dout(n10381));
  jand g10318(.dina(n8769), .dinb(n1213), .dout(n10382));
  jand g10319(.dina(n9126), .dinb(n1076), .dout(n10383));
  jand g10320(.dina(n9491), .dinb(n922), .dout(n10384));
  jor  g10321(.dina(n10384), .dinb(n10383), .dout(n10385));
  jor  g10322(.dina(n10385), .dinb(n10382), .dout(n10386));
  jor  g10323(.dina(n10386), .dinb(n10381), .dout(n10387));
  jxor g10324(.dina(n10387), .dinb(n6039), .dout(n10388));
  jor  g10325(.dina(n10388), .dinb(n10380), .dout(n10389));
  jxor g10326(.dina(n10324), .dinb(n10323), .dout(n10390));
  jnot g10327(.din(n10390), .dout(n10391));
  jand g10328(.dina(n8771), .dinb(n4043), .dout(n10392));
  jand g10329(.dina(n9126), .dinb(n1213), .dout(n10393));
  jand g10330(.dina(n8769), .dinb(n1343), .dout(n10394));
  jand g10331(.dina(n9491), .dinb(n1076), .dout(n10395));
  jor  g10332(.dina(n10395), .dinb(n10394), .dout(n10396));
  jor  g10333(.dina(n10396), .dinb(n10393), .dout(n10397));
  jor  g10334(.dina(n10397), .dinb(n10392), .dout(n10398));
  jxor g10335(.dina(n10398), .dinb(n6039), .dout(n10399));
  jor  g10336(.dina(n10399), .dinb(n10391), .dout(n10400));
  jnot g10337(.din(n10400), .dout(n10401));
  jxor g10338(.dina(n10321), .dinb(n10320), .dout(n10402));
  jnot g10339(.din(n10402), .dout(n10403));
  jand g10340(.dina(n8771), .dinb(n4772), .dout(n10404));
  jand g10341(.dina(n9126), .dinb(n1343), .dout(n10405));
  jand g10342(.dina(n8769), .dinb(n1445), .dout(n10406));
  jand g10343(.dina(n9491), .dinb(n1213), .dout(n10407));
  jor  g10344(.dina(n10407), .dinb(n10406), .dout(n10408));
  jor  g10345(.dina(n10408), .dinb(n10405), .dout(n10409));
  jor  g10346(.dina(n10409), .dinb(n10404), .dout(n10410));
  jxor g10347(.dina(n10410), .dinb(n6039), .dout(n10411));
  jor  g10348(.dina(n10411), .dinb(n10403), .dout(n10412));
  jnot g10349(.din(n10412), .dout(n10413));
  jxor g10350(.dina(n10318), .dinb(n10317), .dout(n10414));
  jnot g10351(.din(n10414), .dout(n10415));
  jand g10352(.dina(n8771), .dinb(n4258), .dout(n10416));
  jand g10353(.dina(n9126), .dinb(n1445), .dout(n10417));
  jand g10354(.dina(n8769), .dinb(n1560), .dout(n10418));
  jand g10355(.dina(n9491), .dinb(n1343), .dout(n10419));
  jor  g10356(.dina(n10419), .dinb(n10418), .dout(n10420));
  jor  g10357(.dina(n10420), .dinb(n10417), .dout(n10421));
  jor  g10358(.dina(n10421), .dinb(n10416), .dout(n10422));
  jxor g10359(.dina(n10422), .dinb(n6039), .dout(n10423));
  jor  g10360(.dina(n10423), .dinb(n10415), .dout(n10424));
  jnot g10361(.din(n10424), .dout(n10425));
  jxor g10362(.dina(n10315), .dinb(n10314), .dout(n10426));
  jnot g10363(.din(n10426), .dout(n10427));
  jand g10364(.dina(n8771), .dinb(n4866), .dout(n10428));
  jand g10365(.dina(n9126), .dinb(n1560), .dout(n10429));
  jand g10366(.dina(n8769), .dinb(n1624), .dout(n10430));
  jand g10367(.dina(n9491), .dinb(n1445), .dout(n10431));
  jor  g10368(.dina(n10431), .dinb(n10430), .dout(n10432));
  jor  g10369(.dina(n10432), .dinb(n10429), .dout(n10433));
  jor  g10370(.dina(n10433), .dinb(n10428), .dout(n10434));
  jxor g10371(.dina(n10434), .dinb(n6039), .dout(n10435));
  jor  g10372(.dina(n10435), .dinb(n10427), .dout(n10436));
  jnot g10373(.din(n10436), .dout(n10437));
  jxor g10374(.dina(n10312), .dinb(n10311), .dout(n10438));
  jnot g10375(.din(n10438), .dout(n10439));
  jand g10376(.dina(n8771), .dinb(n4849), .dout(n10440));
  jand g10377(.dina(n9126), .dinb(n1624), .dout(n10441));
  jand g10378(.dina(n8769), .dinb(n1776), .dout(n10442));
  jand g10379(.dina(n9491), .dinb(n1560), .dout(n10443));
  jor  g10380(.dina(n10443), .dinb(n10442), .dout(n10444));
  jor  g10381(.dina(n10444), .dinb(n10441), .dout(n10445));
  jor  g10382(.dina(n10445), .dinb(n10440), .dout(n10446));
  jxor g10383(.dina(n10446), .dinb(n6039), .dout(n10447));
  jor  g10384(.dina(n10447), .dinb(n10439), .dout(n10448));
  jnot g10385(.din(n10448), .dout(n10449));
  jand g10386(.dina(n8771), .dinb(n5075), .dout(n10450));
  jand g10387(.dina(n9491), .dinb(n1624), .dout(n10451));
  jand g10388(.dina(n9126), .dinb(n1776), .dout(n10452));
  jand g10389(.dina(n8769), .dinb(n1862), .dout(n10453));
  jor  g10390(.dina(n10453), .dinb(n10452), .dout(n10454));
  jor  g10391(.dina(n10454), .dinb(n10451), .dout(n10455));
  jor  g10392(.dina(n10455), .dinb(n10450), .dout(n10456));
  jxor g10393(.dina(n10456), .dinb(n6039), .dout(n10457));
  jnot g10394(.din(n10457), .dout(n10458));
  jxor g10395(.dina(n10307), .dinb(n10306), .dout(n10459));
  jand g10396(.dina(n10459), .dinb(n10458), .dout(n10460));
  jand g10397(.dina(n8771), .dinb(n5092), .dout(n10461));
  jand g10398(.dina(n9491), .dinb(n1776), .dout(n10462));
  jand g10399(.dina(n9126), .dinb(n1862), .dout(n10463));
  jand g10400(.dina(n8769), .dinb(n1956), .dout(n10464));
  jor  g10401(.dina(n10464), .dinb(n10463), .dout(n10465));
  jor  g10402(.dina(n10465), .dinb(n10462), .dout(n10466));
  jor  g10403(.dina(n10466), .dinb(n10461), .dout(n10467));
  jxor g10404(.dina(n10467), .dinb(n6039), .dout(n10468));
  jnot g10405(.din(n10468), .dout(n10469));
  jxor g10406(.dina(n10302), .dinb(n10301), .dout(n10470));
  jand g10407(.dina(n10470), .dinb(n10469), .dout(n10471));
  jxor g10408(.dina(n10299), .dinb(n10298), .dout(n10472));
  jnot g10409(.din(n10472), .dout(n10473));
  jand g10410(.dina(n8771), .dinb(n5440), .dout(n10474));
  jand g10411(.dina(n8769), .dinb(n2067), .dout(n10475));
  jand g10412(.dina(n9126), .dinb(n1956), .dout(n10476));
  jand g10413(.dina(n9491), .dinb(n1862), .dout(n10477));
  jor  g10414(.dina(n10477), .dinb(n10476), .dout(n10478));
  jor  g10415(.dina(n10478), .dinb(n10475), .dout(n10479));
  jor  g10416(.dina(n10479), .dinb(n10474), .dout(n10480));
  jxor g10417(.dina(n10480), .dinb(n6039), .dout(n10481));
  jor  g10418(.dina(n10481), .dinb(n10473), .dout(n10482));
  jxor g10419(.dina(n10296), .dinb(n10295), .dout(n10483));
  jnot g10420(.din(n10483), .dout(n10484));
  jand g10421(.dina(n8771), .dinb(n5303), .dout(n10485));
  jand g10422(.dina(n8769), .dinb(n2128), .dout(n10486));
  jand g10423(.dina(n9126), .dinb(n2067), .dout(n10487));
  jand g10424(.dina(n9491), .dinb(n1956), .dout(n10488));
  jor  g10425(.dina(n10488), .dinb(n10487), .dout(n10489));
  jor  g10426(.dina(n10489), .dinb(n10486), .dout(n10490));
  jor  g10427(.dina(n10490), .dinb(n10485), .dout(n10491));
  jxor g10428(.dina(n10491), .dinb(n6039), .dout(n10492));
  jor  g10429(.dina(n10492), .dinb(n10484), .dout(n10493));
  jxor g10430(.dina(n10293), .dinb(n10292), .dout(n10494));
  jnot g10431(.din(n10494), .dout(n10495));
  jand g10432(.dina(n8771), .dinb(n5624), .dout(n10496));
  jand g10433(.dina(n8769), .dinb(n2237), .dout(n10497));
  jand g10434(.dina(n9126), .dinb(n2128), .dout(n10498));
  jand g10435(.dina(n9491), .dinb(n2067), .dout(n10499));
  jor  g10436(.dina(n10499), .dinb(n10498), .dout(n10500));
  jor  g10437(.dina(n10500), .dinb(n10497), .dout(n10501));
  jor  g10438(.dina(n10501), .dinb(n10496), .dout(n10502));
  jxor g10439(.dina(n10502), .dinb(n6039), .dout(n10503));
  jor  g10440(.dina(n10503), .dinb(n10495), .dout(n10504));
  jand g10441(.dina(n8771), .dinb(n5607), .dout(n10505));
  jand g10442(.dina(n9126), .dinb(n2237), .dout(n10506));
  jand g10443(.dina(n8769), .dinb(n2343), .dout(n10507));
  jand g10444(.dina(n9491), .dinb(n2128), .dout(n10508));
  jor  g10445(.dina(n10508), .dinb(n10507), .dout(n10509));
  jor  g10446(.dina(n10509), .dinb(n10506), .dout(n10510));
  jor  g10447(.dina(n10510), .dinb(n10505), .dout(n10511));
  jxor g10448(.dina(n10511), .dinb(n6039), .dout(n10512));
  jnot g10449(.din(n10512), .dout(n10513));
  jxor g10450(.dina(n10288), .dinb(n10287), .dout(n10514));
  jand g10451(.dina(n10514), .dinb(n10513), .dout(n10515));
  jand g10452(.dina(n8771), .dinb(n5844), .dout(n10516));
  jand g10453(.dina(n8769), .dinb(n2411), .dout(n10517));
  jand g10454(.dina(n9491), .dinb(n2237), .dout(n10518));
  jand g10455(.dina(n9126), .dinb(n2343), .dout(n10519));
  jor  g10456(.dina(n10519), .dinb(n10518), .dout(n10520));
  jor  g10457(.dina(n10520), .dinb(n10517), .dout(n10521));
  jor  g10458(.dina(n10521), .dinb(n10516), .dout(n10522));
  jxor g10459(.dina(n10522), .dinb(n6039), .dout(n10523));
  jnot g10460(.din(n10523), .dout(n10524));
  jxor g10461(.dina(n10283), .dinb(n10282), .dout(n10525));
  jand g10462(.dina(n10525), .dinb(n10524), .dout(n10526));
  jand g10463(.dina(n8771), .dinb(n5861), .dout(n10527));
  jand g10464(.dina(n9126), .dinb(n2411), .dout(n10528));
  jand g10465(.dina(n9491), .dinb(n2343), .dout(n10529));
  jand g10466(.dina(n8769), .dinb(n2497), .dout(n10530));
  jor  g10467(.dina(n10530), .dinb(n10529), .dout(n10531));
  jor  g10468(.dina(n10531), .dinb(n10528), .dout(n10532));
  jor  g10469(.dina(n10532), .dinb(n10527), .dout(n10533));
  jxor g10470(.dina(n10533), .dinb(n6039), .dout(n10534));
  jnot g10471(.din(n10534), .dout(n10535));
  jxor g10472(.dina(n10278), .dinb(n10277), .dout(n10536));
  jand g10473(.dina(n10536), .dinb(n10535), .dout(n10537));
  jxor g10474(.dina(n10275), .dinb(n10274), .dout(n10538));
  jnot g10475(.din(n10538), .dout(n10539));
  jand g10476(.dina(n8771), .dinb(n6247), .dout(n10540));
  jand g10477(.dina(n9491), .dinb(n2411), .dout(n10541));
  jand g10478(.dina(n8769), .dinb(n2602), .dout(n10542));
  jand g10479(.dina(n9126), .dinb(n2497), .dout(n10543));
  jor  g10480(.dina(n10543), .dinb(n10542), .dout(n10544));
  jor  g10481(.dina(n10544), .dinb(n10541), .dout(n10545));
  jor  g10482(.dina(n10545), .dinb(n10540), .dout(n10546));
  jxor g10483(.dina(n10546), .dinb(n6039), .dout(n10547));
  jor  g10484(.dina(n10547), .dinb(n10539), .dout(n10548));
  jxor g10485(.dina(n10272), .dinb(n10271), .dout(n10549));
  jnot g10486(.din(n10549), .dout(n10550));
  jand g10487(.dina(n8771), .dinb(n6050), .dout(n10551));
  jand g10488(.dina(n9126), .dinb(n2602), .dout(n10552));
  jand g10489(.dina(n8769), .dinb(n2695), .dout(n10553));
  jand g10490(.dina(n9491), .dinb(n2497), .dout(n10554));
  jor  g10491(.dina(n10554), .dinb(n10553), .dout(n10555));
  jor  g10492(.dina(n10555), .dinb(n10552), .dout(n10556));
  jor  g10493(.dina(n10556), .dinb(n10551), .dout(n10557));
  jxor g10494(.dina(n10557), .dinb(n6039), .dout(n10558));
  jor  g10495(.dina(n10558), .dinb(n10550), .dout(n10559));
  jxor g10496(.dina(n10269), .dinb(n10268), .dout(n10560));
  jnot g10497(.din(n10560), .dout(n10561));
  jor  g10498(.dina(n8772), .dinb(n6464), .dout(n10562));
  jor  g10499(.dina(n9490), .dinb(n2601), .dout(n10563));
  jor  g10500(.dina(n9127), .dinb(n2694), .dout(n10564));
  jor  g10501(.dina(n8770), .dinb(n2731), .dout(n10565));
  jand g10502(.dina(n10565), .dinb(n10564), .dout(n10566));
  jand g10503(.dina(n10566), .dinb(n10563), .dout(n10567));
  jand g10504(.dina(n10567), .dinb(n10562), .dout(n10568));
  jxor g10505(.dina(n10568), .dinb(\a[8] ), .dout(n10569));
  jor  g10506(.dina(n10569), .dinb(n10561), .dout(n10570));
  jand g10507(.dina(n8771), .dinb(n6591), .dout(n10571));
  jand g10508(.dina(n9491), .dinb(n2695), .dout(n10572));
  jand g10509(.dina(n8769), .dinb(n2808), .dout(n10573));
  jand g10510(.dina(n9126), .dinb(n2732), .dout(n10574));
  jor  g10511(.dina(n10574), .dinb(n10573), .dout(n10575));
  jor  g10512(.dina(n10575), .dinb(n10572), .dout(n10576));
  jor  g10513(.dina(n10576), .dinb(n10571), .dout(n10577));
  jxor g10514(.dina(n10577), .dinb(n6039), .dout(n10578));
  jnot g10515(.din(n10578), .dout(n10579));
  jxor g10516(.dina(n10264), .dinb(n10263), .dout(n10580));
  jand g10517(.dina(n10580), .dinb(n10579), .dout(n10581));
  jand g10518(.dina(n8771), .dinb(n6439), .dout(n10582));
  jand g10519(.dina(n9126), .dinb(n2808), .dout(n10583));
  jand g10520(.dina(n9491), .dinb(n2732), .dout(n10584));
  jand g10521(.dina(n8769), .dinb(n2867), .dout(n10585));
  jor  g10522(.dina(n10585), .dinb(n10584), .dout(n10586));
  jor  g10523(.dina(n10586), .dinb(n10583), .dout(n10587));
  jor  g10524(.dina(n10587), .dinb(n10582), .dout(n10588));
  jxor g10525(.dina(n10588), .dinb(n6039), .dout(n10589));
  jnot g10526(.din(n10589), .dout(n10590));
  jxor g10527(.dina(n10259), .dinb(n10258), .dout(n10591));
  jand g10528(.dina(n10591), .dinb(n10590), .dout(n10592));
  jand g10529(.dina(n8771), .dinb(n6706), .dout(n10593));
  jand g10530(.dina(n9491), .dinb(n2808), .dout(n10594));
  jand g10531(.dina(n8769), .dinb(n2954), .dout(n10595));
  jand g10532(.dina(n9126), .dinb(n2867), .dout(n10596));
  jor  g10533(.dina(n10596), .dinb(n10595), .dout(n10597));
  jor  g10534(.dina(n10597), .dinb(n10594), .dout(n10598));
  jor  g10535(.dina(n10598), .dinb(n10593), .dout(n10599));
  jxor g10536(.dina(n10599), .dinb(n6039), .dout(n10600));
  jnot g10537(.din(n10600), .dout(n10601));
  jxor g10538(.dina(n10254), .dinb(n10253), .dout(n10602));
  jand g10539(.dina(n10602), .dinb(n10601), .dout(n10603));
  jxor g10540(.dina(n10251), .dinb(n10250), .dout(n10604));
  jnot g10541(.din(n10604), .dout(n10605));
  jor  g10542(.dina(n8772), .dinb(n6976), .dout(n10606));
  jor  g10543(.dina(n9127), .dinb(n2953), .dout(n10607));
  jor  g10544(.dina(n8770), .dinb(n2990), .dout(n10608));
  jor  g10545(.dina(n9490), .dinb(n2866), .dout(n10609));
  jand g10546(.dina(n10609), .dinb(n10608), .dout(n10610));
  jand g10547(.dina(n10610), .dinb(n10607), .dout(n10611));
  jand g10548(.dina(n10611), .dinb(n10606), .dout(n10612));
  jxor g10549(.dina(n10612), .dinb(\a[8] ), .dout(n10613));
  jor  g10550(.dina(n10613), .dinb(n10605), .dout(n10614));
  jxor g10551(.dina(n10248), .dinb(n10247), .dout(n10615));
  jnot g10552(.din(n10615), .dout(n10616));
  jor  g10553(.dina(n8772), .dinb(n6988), .dout(n10617));
  jor  g10554(.dina(n8770), .dinb(n3085), .dout(n10618));
  jor  g10555(.dina(n9490), .dinb(n2953), .dout(n10619));
  jor  g10556(.dina(n9127), .dinb(n2990), .dout(n10620));
  jand g10557(.dina(n10620), .dinb(n10619), .dout(n10621));
  jand g10558(.dina(n10621), .dinb(n10618), .dout(n10622));
  jand g10559(.dina(n10622), .dinb(n10617), .dout(n10623));
  jxor g10560(.dina(n10623), .dinb(\a[8] ), .dout(n10624));
  jor  g10561(.dina(n10624), .dinb(n10616), .dout(n10625));
  jxor g10562(.dina(n10245), .dinb(n10244), .dout(n10626));
  jnot g10563(.din(n10626), .dout(n10627));
  jor  g10564(.dina(n8772), .dinb(n6681), .dout(n10628));
  jor  g10565(.dina(n9127), .dinb(n3085), .dout(n10629));
  jor  g10566(.dina(n9490), .dinb(n2990), .dout(n10630));
  jor  g10567(.dina(n8770), .dinb(n3182), .dout(n10631));
  jand g10568(.dina(n10631), .dinb(n10630), .dout(n10632));
  jand g10569(.dina(n10632), .dinb(n10629), .dout(n10633));
  jand g10570(.dina(n10633), .dinb(n10628), .dout(n10634));
  jxor g10571(.dina(n10634), .dinb(\a[8] ), .dout(n10635));
  jor  g10572(.dina(n10635), .dinb(n10627), .dout(n10636));
  jor  g10573(.dina(n8772), .dinb(n7031), .dout(n10637));
  jor  g10574(.dina(n9490), .dinb(n3085), .dout(n10638));
  jor  g10575(.dina(n8770), .dinb(n7962), .dout(n10639));
  jor  g10576(.dina(n9127), .dinb(n3182), .dout(n10640));
  jand g10577(.dina(n10640), .dinb(n10639), .dout(n10641));
  jand g10578(.dina(n10641), .dinb(n10638), .dout(n10642));
  jand g10579(.dina(n10642), .dinb(n10637), .dout(n10643));
  jxor g10580(.dina(n10643), .dinb(\a[8] ), .dout(n10644));
  jnot g10581(.din(n10644), .dout(n10645));
  jxor g10582(.dina(n10242), .dinb(n10241), .dout(n10646));
  jand g10583(.dina(n10646), .dinb(n10645), .dout(n10647));
  jor  g10584(.dina(n8772), .dinb(n7076), .dout(n10648));
  jor  g10585(.dina(n9127), .dinb(n7962), .dout(n10649));
  jor  g10586(.dina(n9490), .dinb(n3182), .dout(n10650));
  jor  g10587(.dina(n8770), .dinb(n3684), .dout(n10651));
  jand g10588(.dina(n10651), .dinb(n10650), .dout(n10652));
  jand g10589(.dina(n10652), .dinb(n10649), .dout(n10653));
  jand g10590(.dina(n10653), .dinb(n10648), .dout(n10654));
  jxor g10591(.dina(n10654), .dinb(\a[8] ), .dout(n10655));
  jnot g10592(.din(n10655), .dout(n10656));
  jxor g10593(.dina(n10239), .dinb(n10238), .dout(n10657));
  jand g10594(.dina(n10657), .dinb(n10656), .dout(n10658));
  jor  g10595(.dina(n8772), .dinb(n7131), .dout(n10659));
  jor  g10596(.dina(n9490), .dinb(n7962), .dout(n10660));
  jor  g10597(.dina(n8770), .dinb(n3414), .dout(n10661));
  jor  g10598(.dina(n9127), .dinb(n3684), .dout(n10662));
  jand g10599(.dina(n10662), .dinb(n10661), .dout(n10663));
  jand g10600(.dina(n10663), .dinb(n10660), .dout(n10664));
  jand g10601(.dina(n10664), .dinb(n10659), .dout(n10665));
  jxor g10602(.dina(n10665), .dinb(\a[8] ), .dout(n10666));
  jnot g10603(.din(n10666), .dout(n10667));
  jor  g10604(.dina(n10219), .dinb(n5833), .dout(n10668));
  jxor g10605(.dina(n10668), .dinb(n10227), .dout(n10669));
  jand g10606(.dina(n10669), .dinb(n10667), .dout(n10670));
  jor  g10607(.dina(n8772), .dinb(n7177), .dout(n10671));
  jor  g10608(.dina(n8770), .dinb(n3516), .dout(n10672));
  jor  g10609(.dina(n9490), .dinb(n3684), .dout(n10673));
  jor  g10610(.dina(n9127), .dinb(n3414), .dout(n10674));
  jand g10611(.dina(n10674), .dinb(n10673), .dout(n10675));
  jand g10612(.dina(n10675), .dinb(n10672), .dout(n10676));
  jand g10613(.dina(n10676), .dinb(n10671), .dout(n10677));
  jxor g10614(.dina(n10677), .dinb(\a[8] ), .dout(n10678));
  jnot g10615(.din(n10678), .dout(n10679));
  jand g10616(.dina(n10216), .dinb(\a[11] ), .dout(n10680));
  jxor g10617(.dina(n10680), .dinb(n10214), .dout(n10681));
  jand g10618(.dina(n10681), .dinb(n10679), .dout(n10682));
  jand g10619(.dina(n8771), .dinb(n8004), .dout(n10683));
  jand g10620(.dina(n9126), .dinb(n7411), .dout(n10684));
  jand g10621(.dina(n9491), .dinb(n7405), .dout(n10685));
  jor  g10622(.dina(n10685), .dinb(n10684), .dout(n10686));
  jor  g10623(.dina(n10686), .dinb(n10683), .dout(n10687));
  jnot g10624(.din(n10687), .dout(n10688));
  jand g10625(.dina(n8765), .dinb(n7411), .dout(n10689));
  jnot g10626(.din(n10689), .dout(n10690));
  jand g10627(.dina(n10690), .dinb(\a[8] ), .dout(n10691));
  jand g10628(.dina(n10691), .dinb(n10688), .dout(n10692));
  jand g10629(.dina(n8771), .dinb(n7407), .dout(n10693));
  jand g10630(.dina(n9491), .dinb(n7326), .dout(n10694));
  jand g10631(.dina(n8769), .dinb(n7411), .dout(n10695));
  jand g10632(.dina(n9126), .dinb(n7405), .dout(n10696));
  jor  g10633(.dina(n10696), .dinb(n10695), .dout(n10697));
  jor  g10634(.dina(n10697), .dinb(n10694), .dout(n10698));
  jor  g10635(.dina(n10698), .dinb(n10693), .dout(n10699));
  jnot g10636(.din(n10699), .dout(n10700));
  jand g10637(.dina(n10700), .dinb(n10692), .dout(n10701));
  jand g10638(.dina(n10701), .dinb(n10216), .dout(n10702));
  jor  g10639(.dina(n8772), .dinb(n7466), .dout(n10703));
  jor  g10640(.dina(n9127), .dinb(n3516), .dout(n10704));
  jor  g10641(.dina(n9490), .dinb(n3414), .dout(n10705));
  jor  g10642(.dina(n8770), .dinb(n3677), .dout(n10706));
  jand g10643(.dina(n10706), .dinb(n10705), .dout(n10707));
  jand g10644(.dina(n10707), .dinb(n10704), .dout(n10708));
  jand g10645(.dina(n10708), .dinb(n10703), .dout(n10709));
  jxor g10646(.dina(n10709), .dinb(\a[8] ), .dout(n10710));
  jnot g10647(.din(n10710), .dout(n10711));
  jxor g10648(.dina(n10701), .dinb(n10216), .dout(n10712));
  jand g10649(.dina(n10712), .dinb(n10711), .dout(n10713));
  jor  g10650(.dina(n10713), .dinb(n10702), .dout(n10714));
  jxor g10651(.dina(n10681), .dinb(n10679), .dout(n10715));
  jand g10652(.dina(n10715), .dinb(n10714), .dout(n10716));
  jor  g10653(.dina(n10716), .dinb(n10682), .dout(n10717));
  jxor g10654(.dina(n10669), .dinb(n10667), .dout(n10718));
  jand g10655(.dina(n10718), .dinb(n10717), .dout(n10719));
  jor  g10656(.dina(n10719), .dinb(n10670), .dout(n10720));
  jxor g10657(.dina(n10657), .dinb(n10656), .dout(n10721));
  jand g10658(.dina(n10721), .dinb(n10720), .dout(n10722));
  jor  g10659(.dina(n10722), .dinb(n10658), .dout(n10723));
  jxor g10660(.dina(n10646), .dinb(n10645), .dout(n10724));
  jand g10661(.dina(n10724), .dinb(n10723), .dout(n10725));
  jor  g10662(.dina(n10725), .dinb(n10647), .dout(n10726));
  jxor g10663(.dina(n10635), .dinb(n10627), .dout(n10727));
  jand g10664(.dina(n10727), .dinb(n10726), .dout(n10728));
  jnot g10665(.din(n10728), .dout(n10729));
  jand g10666(.dina(n10729), .dinb(n10636), .dout(n10730));
  jnot g10667(.din(n10730), .dout(n10731));
  jxor g10668(.dina(n10624), .dinb(n10616), .dout(n10732));
  jand g10669(.dina(n10732), .dinb(n10731), .dout(n10733));
  jnot g10670(.din(n10733), .dout(n10734));
  jand g10671(.dina(n10734), .dinb(n10625), .dout(n10735));
  jnot g10672(.din(n10735), .dout(n10736));
  jxor g10673(.dina(n10613), .dinb(n10605), .dout(n10737));
  jand g10674(.dina(n10737), .dinb(n10736), .dout(n10738));
  jnot g10675(.din(n10738), .dout(n10739));
  jand g10676(.dina(n10739), .dinb(n10614), .dout(n10740));
  jnot g10677(.din(n10740), .dout(n10741));
  jxor g10678(.dina(n10602), .dinb(n10601), .dout(n10742));
  jand g10679(.dina(n10742), .dinb(n10741), .dout(n10743));
  jor  g10680(.dina(n10743), .dinb(n10603), .dout(n10744));
  jxor g10681(.dina(n10591), .dinb(n10590), .dout(n10745));
  jand g10682(.dina(n10745), .dinb(n10744), .dout(n10746));
  jor  g10683(.dina(n10746), .dinb(n10592), .dout(n10747));
  jxor g10684(.dina(n10580), .dinb(n10579), .dout(n10748));
  jand g10685(.dina(n10748), .dinb(n10747), .dout(n10749));
  jor  g10686(.dina(n10749), .dinb(n10581), .dout(n10750));
  jxor g10687(.dina(n10569), .dinb(n10561), .dout(n10751));
  jand g10688(.dina(n10751), .dinb(n10750), .dout(n10752));
  jnot g10689(.din(n10752), .dout(n10753));
  jand g10690(.dina(n10753), .dinb(n10570), .dout(n10754));
  jnot g10691(.din(n10754), .dout(n10755));
  jxor g10692(.dina(n10558), .dinb(n10550), .dout(n10756));
  jand g10693(.dina(n10756), .dinb(n10755), .dout(n10757));
  jnot g10694(.din(n10757), .dout(n10758));
  jand g10695(.dina(n10758), .dinb(n10559), .dout(n10759));
  jnot g10696(.din(n10759), .dout(n10760));
  jxor g10697(.dina(n10547), .dinb(n10539), .dout(n10761));
  jand g10698(.dina(n10761), .dinb(n10760), .dout(n10762));
  jnot g10699(.din(n10762), .dout(n10763));
  jand g10700(.dina(n10763), .dinb(n10548), .dout(n10764));
  jnot g10701(.din(n10764), .dout(n10765));
  jxor g10702(.dina(n10536), .dinb(n10535), .dout(n10766));
  jand g10703(.dina(n10766), .dinb(n10765), .dout(n10767));
  jor  g10704(.dina(n10767), .dinb(n10537), .dout(n10768));
  jxor g10705(.dina(n10525), .dinb(n10524), .dout(n10769));
  jand g10706(.dina(n10769), .dinb(n10768), .dout(n10770));
  jor  g10707(.dina(n10770), .dinb(n10526), .dout(n10771));
  jxor g10708(.dina(n10514), .dinb(n10513), .dout(n10772));
  jand g10709(.dina(n10772), .dinb(n10771), .dout(n10773));
  jor  g10710(.dina(n10773), .dinb(n10515), .dout(n10774));
  jxor g10711(.dina(n10503), .dinb(n10495), .dout(n10775));
  jand g10712(.dina(n10775), .dinb(n10774), .dout(n10776));
  jnot g10713(.din(n10776), .dout(n10777));
  jand g10714(.dina(n10777), .dinb(n10504), .dout(n10778));
  jnot g10715(.din(n10778), .dout(n10779));
  jxor g10716(.dina(n10492), .dinb(n10484), .dout(n10780));
  jand g10717(.dina(n10780), .dinb(n10779), .dout(n10781));
  jnot g10718(.din(n10781), .dout(n10782));
  jand g10719(.dina(n10782), .dinb(n10493), .dout(n10783));
  jnot g10720(.din(n10783), .dout(n10784));
  jxor g10721(.dina(n10481), .dinb(n10473), .dout(n10785));
  jand g10722(.dina(n10785), .dinb(n10784), .dout(n10786));
  jnot g10723(.din(n10786), .dout(n10787));
  jand g10724(.dina(n10787), .dinb(n10482), .dout(n10788));
  jnot g10725(.din(n10788), .dout(n10789));
  jxor g10726(.dina(n10470), .dinb(n10469), .dout(n10790));
  jand g10727(.dina(n10790), .dinb(n10789), .dout(n10791));
  jor  g10728(.dina(n10791), .dinb(n10471), .dout(n10792));
  jxor g10729(.dina(n10459), .dinb(n10458), .dout(n10793));
  jand g10730(.dina(n10793), .dinb(n10792), .dout(n10794));
  jor  g10731(.dina(n10794), .dinb(n10460), .dout(n10795));
  jxor g10732(.dina(n10447), .dinb(n10439), .dout(n10796));
  jand g10733(.dina(n10796), .dinb(n10795), .dout(n10797));
  jor  g10734(.dina(n10797), .dinb(n10449), .dout(n10798));
  jxor g10735(.dina(n10435), .dinb(n10427), .dout(n10799));
  jand g10736(.dina(n10799), .dinb(n10798), .dout(n10800));
  jor  g10737(.dina(n10800), .dinb(n10437), .dout(n10801));
  jxor g10738(.dina(n10423), .dinb(n10415), .dout(n10802));
  jand g10739(.dina(n10802), .dinb(n10801), .dout(n10803));
  jor  g10740(.dina(n10803), .dinb(n10425), .dout(n10804));
  jxor g10741(.dina(n10411), .dinb(n10403), .dout(n10805));
  jand g10742(.dina(n10805), .dinb(n10804), .dout(n10806));
  jor  g10743(.dina(n10806), .dinb(n10413), .dout(n10807));
  jxor g10744(.dina(n10399), .dinb(n10391), .dout(n10808));
  jand g10745(.dina(n10808), .dinb(n10807), .dout(n10809));
  jor  g10746(.dina(n10809), .dinb(n10401), .dout(n10810));
  jxor g10747(.dina(n10388), .dinb(n10380), .dout(n10811));
  jand g10748(.dina(n10811), .dinb(n10810), .dout(n10812));
  jnot g10749(.din(n10812), .dout(n10813));
  jand g10750(.dina(n10813), .dinb(n10389), .dout(n10814));
  jnot g10751(.din(n10814), .dout(n10815));
  jxor g10752(.dina(n10377), .dinb(n10369), .dout(n10816));
  jand g10753(.dina(n10816), .dinb(n10815), .dout(n10817));
  jnot g10754(.din(n10817), .dout(n10818));
  jand g10755(.dina(n10818), .dinb(n10378), .dout(n10819));
  jnot g10756(.din(n10819), .dout(n10820));
  jxor g10757(.dina(n10344), .dinb(n10343), .dout(n10821));
  jand g10758(.dina(n10821), .dinb(n10820), .dout(n10822));
  jand g10759(.dina(n4636), .dinb(n67), .dout(n10823));
  jand g10760(.dina(n9917), .dinb(n4451), .dout(n10824));
  jand g10761(.dina(n10350), .dinb(n4598), .dout(n10825));
  jor  g10762(.dina(n66), .dinb(n9913), .dout(n10826));
  jnot g10763(.din(n10826), .dout(n10827));
  jand g10764(.dina(n10827), .dinb(n4631), .dout(n10828));
  jor  g10765(.dina(n10828), .dinb(n10825), .dout(n10829));
  jor  g10766(.dina(n10829), .dinb(n10824), .dout(n10830));
  jor  g10767(.dina(n10830), .dinb(n10823), .dout(n10831));
  jxor g10768(.dina(n10831), .dinb(n64), .dout(n10832));
  jnot g10769(.din(n10832), .dout(n10833));
  jxor g10770(.dina(n10821), .dinb(n10820), .dout(n10834));
  jand g10771(.dina(n10834), .dinb(n10833), .dout(n10835));
  jor  g10772(.dina(n10835), .dinb(n10822), .dout(n10836));
  jxor g10773(.dina(n10358), .dinb(n10357), .dout(n10837));
  jand g10774(.dina(n10837), .dinb(n10836), .dout(n10838));
  jnot g10775(.din(n10838), .dout(n10839));
  jnot g10776(.din(\a[0] ), .dout(n10840));
  jnot g10777(.din(\a[1] ), .dout(n10841));
  jand g10778(.dina(n10841), .dinb(n10840), .dout(n10842));
  jxor g10779(.dina(\a[2] ), .dinb(\a[1] ), .dout(n10843));
  jand g10780(.dina(n10843), .dinb(n10842), .dout(n10844));
  jnot g10781(.din(n10844), .dout(n10845));
  jand g10782(.dina(n10843), .dinb(\a[0] ), .dout(n10846));
  jnot g10783(.din(n10846), .dout(n10847));
  jor  g10784(.dina(n10847), .dinb(n4728), .dout(n10848));
  jand g10785(.dina(n10848), .dinb(n10845), .dout(n10849));
  jor  g10786(.dina(n10849), .dinb(n4630), .dout(n10850));
  jxor g10787(.dina(n10850), .dinb(\a[2] ), .dout(n10851));
  jand g10788(.dina(n4752), .dinb(n67), .dout(n10852));
  jand g10789(.dina(n10350), .dinb(n4451), .dout(n10853));
  jand g10790(.dina(n9917), .dinb(n4358), .dout(n10854));
  jand g10791(.dina(n10827), .dinb(n4598), .dout(n10855));
  jor  g10792(.dina(n10855), .dinb(n10854), .dout(n10856));
  jor  g10793(.dina(n10856), .dinb(n10853), .dout(n10857));
  jor  g10794(.dina(n10857), .dinb(n10852), .dout(n10858));
  jxor g10795(.dina(n10858), .dinb(n64), .dout(n10859));
  jor  g10796(.dina(n10859), .dinb(n10851), .dout(n10860));
  jxor g10797(.dina(n10859), .dinb(n10851), .dout(n10861));
  jxor g10798(.dina(n10816), .dinb(n10815), .dout(n10862));
  jand g10799(.dina(n10862), .dinb(n10861), .dout(n10863));
  jnot g10800(.din(n10863), .dout(n10864));
  jand g10801(.dina(n10864), .dinb(n10860), .dout(n10865));
  jnot g10802(.din(n10865), .dout(n10866));
  jxor g10803(.dina(n10834), .dinb(n10833), .dout(n10867));
  jand g10804(.dina(n10867), .dinb(n10866), .dout(n10868));
  jnot g10805(.din(n10868), .dout(n10869));
  jand g10806(.dina(n4446), .dinb(n67), .dout(n10870));
  jand g10807(.dina(n10827), .dinb(n4451), .dout(n10871));
  jand g10808(.dina(n10350), .dinb(n4358), .dout(n10872));
  jand g10809(.dina(n9917), .dinb(n3853), .dout(n10873));
  jor  g10810(.dina(n10873), .dinb(n10872), .dout(n10874));
  jor  g10811(.dina(n10874), .dinb(n10871), .dout(n10875));
  jor  g10812(.dina(n10875), .dinb(n10870), .dout(n10876));
  jxor g10813(.dina(n10876), .dinb(n64), .dout(n10877));
  jnot g10814(.din(n10877), .dout(n10878));
  jxor g10815(.dina(n10811), .dinb(n10810), .dout(n10879));
  jand g10816(.dina(n10879), .dinb(n10878), .dout(n10880));
  jand g10817(.dina(n4545), .dinb(n67), .dout(n10881));
  jand g10818(.dina(n10350), .dinb(n3853), .dout(n10882));
  jand g10819(.dina(n10827), .dinb(n4358), .dout(n10883));
  jand g10820(.dina(n9917), .dinb(n922), .dout(n10884));
  jor  g10821(.dina(n10884), .dinb(n10883), .dout(n10885));
  jor  g10822(.dina(n10885), .dinb(n10882), .dout(n10886));
  jor  g10823(.dina(n10886), .dinb(n10881), .dout(n10887));
  jxor g10824(.dina(n10887), .dinb(n64), .dout(n10888));
  jnot g10825(.din(n10888), .dout(n10889));
  jxor g10826(.dina(n10808), .dinb(n10807), .dout(n10890));
  jand g10827(.dina(n10890), .dinb(n10889), .dout(n10891));
  jnot g10828(.din(n10891), .dout(n10892));
  jand g10829(.dina(n3848), .dinb(n67), .dout(n10893));
  jand g10830(.dina(n10350), .dinb(n922), .dout(n10894));
  jand g10831(.dina(n10827), .dinb(n3853), .dout(n10895));
  jand g10832(.dina(n9917), .dinb(n1076), .dout(n10896));
  jor  g10833(.dina(n10896), .dinb(n10895), .dout(n10897));
  jor  g10834(.dina(n10897), .dinb(n10894), .dout(n10898));
  jor  g10835(.dina(n10898), .dinb(n10893), .dout(n10899));
  jxor g10836(.dina(n10899), .dinb(n64), .dout(n10900));
  jnot g10837(.din(n10900), .dout(n10901));
  jxor g10838(.dina(n10805), .dinb(n10804), .dout(n10902));
  jand g10839(.dina(n10902), .dinb(n10901), .dout(n10903));
  jnot g10840(.din(n10903), .dout(n10904));
  jand g10841(.dina(n4026), .dinb(n67), .dout(n10905));
  jand g10842(.dina(n10350), .dinb(n1076), .dout(n10906));
  jand g10843(.dina(n10827), .dinb(n922), .dout(n10907));
  jand g10844(.dina(n9917), .dinb(n1213), .dout(n10908));
  jor  g10845(.dina(n10908), .dinb(n10907), .dout(n10909));
  jor  g10846(.dina(n10909), .dinb(n10906), .dout(n10910));
  jor  g10847(.dina(n10910), .dinb(n10905), .dout(n10911));
  jxor g10848(.dina(n10911), .dinb(n64), .dout(n10912));
  jnot g10849(.din(n10912), .dout(n10913));
  jxor g10850(.dina(n10802), .dinb(n10801), .dout(n10914));
  jand g10851(.dina(n10914), .dinb(n10913), .dout(n10915));
  jnot g10852(.din(n10915), .dout(n10916));
  jand g10853(.dina(n4043), .dinb(n67), .dout(n10917));
  jand g10854(.dina(n10827), .dinb(n1076), .dout(n10918));
  jand g10855(.dina(n10350), .dinb(n1213), .dout(n10919));
  jand g10856(.dina(n9917), .dinb(n1343), .dout(n10920));
  jor  g10857(.dina(n10920), .dinb(n10919), .dout(n10921));
  jor  g10858(.dina(n10921), .dinb(n10918), .dout(n10922));
  jor  g10859(.dina(n10922), .dinb(n10917), .dout(n10923));
  jxor g10860(.dina(n10923), .dinb(n64), .dout(n10924));
  jnot g10861(.din(n10924), .dout(n10925));
  jxor g10862(.dina(n10799), .dinb(n10798), .dout(n10926));
  jand g10863(.dina(n10926), .dinb(n10925), .dout(n10927));
  jnot g10864(.din(n10927), .dout(n10928));
  jand g10865(.dina(n4772), .dinb(n67), .dout(n10929));
  jand g10866(.dina(n10827), .dinb(n1213), .dout(n10930));
  jand g10867(.dina(n10350), .dinb(n1343), .dout(n10931));
  jand g10868(.dina(n9917), .dinb(n1445), .dout(n10932));
  jor  g10869(.dina(n10932), .dinb(n10931), .dout(n10933));
  jor  g10870(.dina(n10933), .dinb(n10930), .dout(n10934));
  jor  g10871(.dina(n10934), .dinb(n10929), .dout(n10935));
  jxor g10872(.dina(n10935), .dinb(n64), .dout(n10936));
  jnot g10873(.din(n10936), .dout(n10937));
  jxor g10874(.dina(n10796), .dinb(n10795), .dout(n10938));
  jand g10875(.dina(n10938), .dinb(n10937), .dout(n10939));
  jnot g10876(.din(n10939), .dout(n10940));
  jxor g10877(.dina(n10793), .dinb(n10792), .dout(n10941));
  jnot g10878(.din(n10941), .dout(n10942));
  jand g10879(.dina(n4258), .dinb(n67), .dout(n10943));
  jand g10880(.dina(n10350), .dinb(n1445), .dout(n10944));
  jand g10881(.dina(n9917), .dinb(n1560), .dout(n10945));
  jand g10882(.dina(n10827), .dinb(n1343), .dout(n10946));
  jor  g10883(.dina(n10946), .dinb(n10945), .dout(n10947));
  jor  g10884(.dina(n10947), .dinb(n10944), .dout(n10948));
  jor  g10885(.dina(n10948), .dinb(n10943), .dout(n10949));
  jxor g10886(.dina(n10949), .dinb(n64), .dout(n10950));
  jor  g10887(.dina(n10950), .dinb(n10942), .dout(n10951));
  jxor g10888(.dina(n10790), .dinb(n10789), .dout(n10952));
  jnot g10889(.din(n10952), .dout(n10953));
  jand g10890(.dina(n4866), .dinb(n67), .dout(n10954));
  jand g10891(.dina(n10350), .dinb(n1560), .dout(n10955));
  jand g10892(.dina(n9917), .dinb(n1624), .dout(n10956));
  jand g10893(.dina(n10827), .dinb(n1445), .dout(n10957));
  jor  g10894(.dina(n10957), .dinb(n10956), .dout(n10958));
  jor  g10895(.dina(n10958), .dinb(n10955), .dout(n10959));
  jor  g10896(.dina(n10959), .dinb(n10954), .dout(n10960));
  jxor g10897(.dina(n10960), .dinb(n64), .dout(n10961));
  jor  g10898(.dina(n10961), .dinb(n10953), .dout(n10962));
  jand g10899(.dina(n4849), .dinb(n67), .dout(n10963));
  jand g10900(.dina(n10827), .dinb(n1560), .dout(n10964));
  jand g10901(.dina(n10350), .dinb(n1624), .dout(n10965));
  jand g10902(.dina(n9917), .dinb(n1776), .dout(n10966));
  jor  g10903(.dina(n10966), .dinb(n10965), .dout(n10967));
  jor  g10904(.dina(n10967), .dinb(n10964), .dout(n10968));
  jor  g10905(.dina(n10968), .dinb(n10963), .dout(n10969));
  jxor g10906(.dina(n10969), .dinb(n64), .dout(n10970));
  jnot g10907(.din(n10970), .dout(n10971));
  jxor g10908(.dina(n10785), .dinb(n10784), .dout(n10972));
  jand g10909(.dina(n10972), .dinb(n10971), .dout(n10973));
  jand g10910(.dina(n5075), .dinb(n67), .dout(n10974));
  jand g10911(.dina(n10827), .dinb(n1624), .dout(n10975));
  jand g10912(.dina(n10350), .dinb(n1776), .dout(n10976));
  jand g10913(.dina(n9917), .dinb(n1862), .dout(n10977));
  jor  g10914(.dina(n10977), .dinb(n10976), .dout(n10978));
  jor  g10915(.dina(n10978), .dinb(n10975), .dout(n10979));
  jor  g10916(.dina(n10979), .dinb(n10974), .dout(n10980));
  jxor g10917(.dina(n10980), .dinb(n64), .dout(n10981));
  jnot g10918(.din(n10981), .dout(n10982));
  jxor g10919(.dina(n10780), .dinb(n10779), .dout(n10983));
  jand g10920(.dina(n10983), .dinb(n10982), .dout(n10984));
  jand g10921(.dina(n5092), .dinb(n67), .dout(n10985));
  jand g10922(.dina(n10827), .dinb(n1776), .dout(n10986));
  jand g10923(.dina(n10350), .dinb(n1862), .dout(n10987));
  jand g10924(.dina(n9917), .dinb(n1956), .dout(n10988));
  jor  g10925(.dina(n10988), .dinb(n10987), .dout(n10989));
  jor  g10926(.dina(n10989), .dinb(n10986), .dout(n10990));
  jor  g10927(.dina(n10990), .dinb(n10985), .dout(n10991));
  jxor g10928(.dina(n10991), .dinb(n64), .dout(n10992));
  jnot g10929(.din(n10992), .dout(n10993));
  jxor g10930(.dina(n10775), .dinb(n10774), .dout(n10994));
  jand g10931(.dina(n10994), .dinb(n10993), .dout(n10995));
  jxor g10932(.dina(n10772), .dinb(n10771), .dout(n10996));
  jnot g10933(.din(n10996), .dout(n10997));
  jand g10934(.dina(n5440), .dinb(n67), .dout(n10998));
  jand g10935(.dina(n9917), .dinb(n2067), .dout(n10999));
  jand g10936(.dina(n10350), .dinb(n1956), .dout(n11000));
  jand g10937(.dina(n10827), .dinb(n1862), .dout(n11001));
  jor  g10938(.dina(n11001), .dinb(n11000), .dout(n11002));
  jor  g10939(.dina(n11002), .dinb(n10999), .dout(n11003));
  jor  g10940(.dina(n11003), .dinb(n10998), .dout(n11004));
  jxor g10941(.dina(n11004), .dinb(n64), .dout(n11005));
  jor  g10942(.dina(n11005), .dinb(n10997), .dout(n11006));
  jxor g10943(.dina(n10769), .dinb(n10768), .dout(n11007));
  jnot g10944(.din(n11007), .dout(n11008));
  jand g10945(.dina(n5303), .dinb(n67), .dout(n11009));
  jand g10946(.dina(n9917), .dinb(n2128), .dout(n11010));
  jand g10947(.dina(n10350), .dinb(n2067), .dout(n11011));
  jand g10948(.dina(n10827), .dinb(n1956), .dout(n11012));
  jor  g10949(.dina(n11012), .dinb(n11011), .dout(n11013));
  jor  g10950(.dina(n11013), .dinb(n11010), .dout(n11014));
  jor  g10951(.dina(n11014), .dinb(n11009), .dout(n11015));
  jxor g10952(.dina(n11015), .dinb(n64), .dout(n11016));
  jor  g10953(.dina(n11016), .dinb(n11008), .dout(n11017));
  jxor g10954(.dina(n10766), .dinb(n10765), .dout(n11018));
  jnot g10955(.din(n11018), .dout(n11019));
  jand g10956(.dina(n5624), .dinb(n67), .dout(n11020));
  jand g10957(.dina(n9917), .dinb(n2237), .dout(n11021));
  jand g10958(.dina(n10350), .dinb(n2128), .dout(n11022));
  jand g10959(.dina(n10827), .dinb(n2067), .dout(n11023));
  jor  g10960(.dina(n11023), .dinb(n11022), .dout(n11024));
  jor  g10961(.dina(n11024), .dinb(n11021), .dout(n11025));
  jor  g10962(.dina(n11025), .dinb(n11020), .dout(n11026));
  jxor g10963(.dina(n11026), .dinb(n64), .dout(n11027));
  jor  g10964(.dina(n11027), .dinb(n11019), .dout(n11028));
  jand g10965(.dina(n5607), .dinb(n67), .dout(n11029));
  jand g10966(.dina(n10350), .dinb(n2237), .dout(n11030));
  jand g10967(.dina(n9917), .dinb(n2343), .dout(n11031));
  jand g10968(.dina(n10827), .dinb(n2128), .dout(n11032));
  jor  g10969(.dina(n11032), .dinb(n11031), .dout(n11033));
  jor  g10970(.dina(n11033), .dinb(n11030), .dout(n11034));
  jor  g10971(.dina(n11034), .dinb(n11029), .dout(n11035));
  jxor g10972(.dina(n11035), .dinb(n64), .dout(n11036));
  jnot g10973(.din(n11036), .dout(n11037));
  jxor g10974(.dina(n10761), .dinb(n10760), .dout(n11038));
  jand g10975(.dina(n11038), .dinb(n11037), .dout(n11039));
  jand g10976(.dina(n5844), .dinb(n67), .dout(n11040));
  jand g10977(.dina(n9917), .dinb(n2411), .dout(n11041));
  jand g10978(.dina(n10827), .dinb(n2237), .dout(n11042));
  jand g10979(.dina(n10350), .dinb(n2343), .dout(n11043));
  jor  g10980(.dina(n11043), .dinb(n11042), .dout(n11044));
  jor  g10981(.dina(n11044), .dinb(n11041), .dout(n11045));
  jor  g10982(.dina(n11045), .dinb(n11040), .dout(n11046));
  jxor g10983(.dina(n11046), .dinb(n64), .dout(n11047));
  jnot g10984(.din(n11047), .dout(n11048));
  jxor g10985(.dina(n10756), .dinb(n10755), .dout(n11049));
  jand g10986(.dina(n11049), .dinb(n11048), .dout(n11050));
  jand g10987(.dina(n5861), .dinb(n67), .dout(n11051));
  jand g10988(.dina(n10350), .dinb(n2411), .dout(n11052));
  jand g10989(.dina(n10827), .dinb(n2343), .dout(n11053));
  jand g10990(.dina(n9917), .dinb(n2497), .dout(n11054));
  jor  g10991(.dina(n11054), .dinb(n11053), .dout(n11055));
  jor  g10992(.dina(n11055), .dinb(n11052), .dout(n11056));
  jor  g10993(.dina(n11056), .dinb(n11051), .dout(n11057));
  jxor g10994(.dina(n11057), .dinb(n64), .dout(n11058));
  jnot g10995(.din(n11058), .dout(n11059));
  jxor g10996(.dina(n10751), .dinb(n10750), .dout(n11060));
  jand g10997(.dina(n11060), .dinb(n11059), .dout(n11061));
  jxor g10998(.dina(n10748), .dinb(n10747), .dout(n11062));
  jnot g10999(.din(n11062), .dout(n11063));
  jand g11000(.dina(n6247), .dinb(n67), .dout(n11064));
  jand g11001(.dina(n10827), .dinb(n2411), .dout(n11065));
  jand g11002(.dina(n9917), .dinb(n2602), .dout(n11066));
  jand g11003(.dina(n10350), .dinb(n2497), .dout(n11067));
  jor  g11004(.dina(n11067), .dinb(n11066), .dout(n11068));
  jor  g11005(.dina(n11068), .dinb(n11065), .dout(n11069));
  jor  g11006(.dina(n11069), .dinb(n11064), .dout(n11070));
  jxor g11007(.dina(n11070), .dinb(n64), .dout(n11071));
  jor  g11008(.dina(n11071), .dinb(n11063), .dout(n11072));
  jxor g11009(.dina(n10745), .dinb(n10744), .dout(n11073));
  jnot g11010(.din(n11073), .dout(n11074));
  jand g11011(.dina(n6050), .dinb(n67), .dout(n11075));
  jand g11012(.dina(n10350), .dinb(n2602), .dout(n11076));
  jand g11013(.dina(n9917), .dinb(n2695), .dout(n11077));
  jand g11014(.dina(n10827), .dinb(n2497), .dout(n11078));
  jor  g11015(.dina(n11078), .dinb(n11077), .dout(n11079));
  jor  g11016(.dina(n11079), .dinb(n11076), .dout(n11080));
  jor  g11017(.dina(n11080), .dinb(n11075), .dout(n11081));
  jxor g11018(.dina(n11081), .dinb(n64), .dout(n11082));
  jor  g11019(.dina(n11082), .dinb(n11074), .dout(n11083));
  jxor g11020(.dina(n10742), .dinb(n10741), .dout(n11084));
  jnot g11021(.din(n11084), .dout(n11085));
  jor  g11022(.dina(n6464), .dinb(n9919), .dout(n11086));
  jor  g11023(.dina(n10826), .dinb(n2601), .dout(n11087));
  jor  g11024(.dina(n10351), .dinb(n2694), .dout(n11088));
  jor  g11025(.dina(n9918), .dinb(n2731), .dout(n11089));
  jand g11026(.dina(n11089), .dinb(n11088), .dout(n11090));
  jand g11027(.dina(n11090), .dinb(n11087), .dout(n11091));
  jand g11028(.dina(n11091), .dinb(n11086), .dout(n11092));
  jxor g11029(.dina(n11092), .dinb(\a[5] ), .dout(n11093));
  jor  g11030(.dina(n11093), .dinb(n11085), .dout(n11094));
  jand g11031(.dina(n6591), .dinb(n67), .dout(n11095));
  jand g11032(.dina(n10827), .dinb(n2695), .dout(n11096));
  jand g11033(.dina(n9917), .dinb(n2808), .dout(n11097));
  jand g11034(.dina(n10350), .dinb(n2732), .dout(n11098));
  jor  g11035(.dina(n11098), .dinb(n11097), .dout(n11099));
  jor  g11036(.dina(n11099), .dinb(n11096), .dout(n11100));
  jor  g11037(.dina(n11100), .dinb(n11095), .dout(n11101));
  jxor g11038(.dina(n11101), .dinb(n64), .dout(n11102));
  jnot g11039(.din(n11102), .dout(n11103));
  jxor g11040(.dina(n10737), .dinb(n10736), .dout(n11104));
  jand g11041(.dina(n11104), .dinb(n11103), .dout(n11105));
  jand g11042(.dina(n6439), .dinb(n67), .dout(n11106));
  jand g11043(.dina(n10350), .dinb(n2808), .dout(n11107));
  jand g11044(.dina(n10827), .dinb(n2732), .dout(n11108));
  jand g11045(.dina(n9917), .dinb(n2867), .dout(n11109));
  jor  g11046(.dina(n11109), .dinb(n11108), .dout(n11110));
  jor  g11047(.dina(n11110), .dinb(n11107), .dout(n11111));
  jor  g11048(.dina(n11111), .dinb(n11106), .dout(n11112));
  jxor g11049(.dina(n11112), .dinb(n64), .dout(n11113));
  jnot g11050(.din(n11113), .dout(n11114));
  jxor g11051(.dina(n10732), .dinb(n10731), .dout(n11115));
  jand g11052(.dina(n11115), .dinb(n11114), .dout(n11116));
  jand g11053(.dina(n6706), .dinb(n67), .dout(n11117));
  jand g11054(.dina(n10827), .dinb(n2808), .dout(n11118));
  jand g11055(.dina(n9917), .dinb(n2954), .dout(n11119));
  jand g11056(.dina(n10350), .dinb(n2867), .dout(n11120));
  jor  g11057(.dina(n11120), .dinb(n11119), .dout(n11121));
  jor  g11058(.dina(n11121), .dinb(n11118), .dout(n11122));
  jor  g11059(.dina(n11122), .dinb(n11117), .dout(n11123));
  jxor g11060(.dina(n11123), .dinb(n64), .dout(n11124));
  jnot g11061(.din(n11124), .dout(n11125));
  jxor g11062(.dina(n10727), .dinb(n10726), .dout(n11126));
  jand g11063(.dina(n11126), .dinb(n11125), .dout(n11127));
  jxor g11064(.dina(n10724), .dinb(n10723), .dout(n11128));
  jnot g11065(.din(n11128), .dout(n11129));
  jor  g11066(.dina(n6976), .dinb(n9919), .dout(n11130));
  jor  g11067(.dina(n10351), .dinb(n2953), .dout(n11131));
  jor  g11068(.dina(n9918), .dinb(n2990), .dout(n11132));
  jor  g11069(.dina(n10826), .dinb(n2866), .dout(n11133));
  jand g11070(.dina(n11133), .dinb(n11132), .dout(n11134));
  jand g11071(.dina(n11134), .dinb(n11131), .dout(n11135));
  jand g11072(.dina(n11135), .dinb(n11130), .dout(n11136));
  jxor g11073(.dina(n11136), .dinb(\a[5] ), .dout(n11137));
  jor  g11074(.dina(n11137), .dinb(n11129), .dout(n11138));
  jxor g11075(.dina(n10721), .dinb(n10720), .dout(n11139));
  jnot g11076(.din(n11139), .dout(n11140));
  jor  g11077(.dina(n6988), .dinb(n9919), .dout(n11141));
  jor  g11078(.dina(n9918), .dinb(n3085), .dout(n11142));
  jor  g11079(.dina(n10826), .dinb(n2953), .dout(n11143));
  jor  g11080(.dina(n10351), .dinb(n2990), .dout(n11144));
  jand g11081(.dina(n11144), .dinb(n11143), .dout(n11145));
  jand g11082(.dina(n11145), .dinb(n11142), .dout(n11146));
  jand g11083(.dina(n11146), .dinb(n11141), .dout(n11147));
  jxor g11084(.dina(n11147), .dinb(\a[5] ), .dout(n11148));
  jor  g11085(.dina(n11148), .dinb(n11140), .dout(n11149));
  jxor g11086(.dina(n10718), .dinb(n10717), .dout(n11150));
  jnot g11087(.din(n11150), .dout(n11151));
  jor  g11088(.dina(n6681), .dinb(n9919), .dout(n11152));
  jor  g11089(.dina(n10351), .dinb(n3085), .dout(n11153));
  jor  g11090(.dina(n10826), .dinb(n2990), .dout(n11154));
  jor  g11091(.dina(n9918), .dinb(n3182), .dout(n11155));
  jand g11092(.dina(n11155), .dinb(n11154), .dout(n11156));
  jand g11093(.dina(n11156), .dinb(n11153), .dout(n11157));
  jand g11094(.dina(n11157), .dinb(n11152), .dout(n11158));
  jxor g11095(.dina(n11158), .dinb(\a[5] ), .dout(n11159));
  jor  g11096(.dina(n11159), .dinb(n11151), .dout(n11160));
  jor  g11097(.dina(n7031), .dinb(n9919), .dout(n11161));
  jor  g11098(.dina(n10826), .dinb(n3085), .dout(n11162));
  jor  g11099(.dina(n9918), .dinb(n7962), .dout(n11163));
  jor  g11100(.dina(n10351), .dinb(n3182), .dout(n11164));
  jand g11101(.dina(n11164), .dinb(n11163), .dout(n11165));
  jand g11102(.dina(n11165), .dinb(n11162), .dout(n11166));
  jand g11103(.dina(n11166), .dinb(n11161), .dout(n11167));
  jxor g11104(.dina(n11167), .dinb(\a[5] ), .dout(n11168));
  jnot g11105(.din(n11168), .dout(n11169));
  jxor g11106(.dina(n10715), .dinb(n10714), .dout(n11170));
  jand g11107(.dina(n11170), .dinb(n11169), .dout(n11171));
  jor  g11108(.dina(n7076), .dinb(n9919), .dout(n11172));
  jor  g11109(.dina(n10351), .dinb(n7962), .dout(n11173));
  jor  g11110(.dina(n10826), .dinb(n3182), .dout(n11174));
  jor  g11111(.dina(n9918), .dinb(n3684), .dout(n11175));
  jand g11112(.dina(n11175), .dinb(n11174), .dout(n11176));
  jand g11113(.dina(n11176), .dinb(n11173), .dout(n11177));
  jand g11114(.dina(n11177), .dinb(n11172), .dout(n11178));
  jxor g11115(.dina(n11178), .dinb(\a[5] ), .dout(n11179));
  jnot g11116(.din(n11179), .dout(n11180));
  jxor g11117(.dina(n10712), .dinb(n10711), .dout(n11181));
  jand g11118(.dina(n11181), .dinb(n11180), .dout(n11182));
  jor  g11119(.dina(n7131), .dinb(n9919), .dout(n11183));
  jor  g11120(.dina(n10826), .dinb(n7962), .dout(n11184));
  jor  g11121(.dina(n9918), .dinb(n3414), .dout(n11185));
  jor  g11122(.dina(n10351), .dinb(n3684), .dout(n11186));
  jand g11123(.dina(n11186), .dinb(n11185), .dout(n11187));
  jand g11124(.dina(n11187), .dinb(n11184), .dout(n11188));
  jand g11125(.dina(n11188), .dinb(n11183), .dout(n11189));
  jxor g11126(.dina(n11189), .dinb(n64), .dout(n11190));
  jor  g11127(.dina(n10692), .dinb(n6039), .dout(n11191));
  jxor g11128(.dina(n11191), .dinb(n10700), .dout(n11192));
  jand g11129(.dina(n11192), .dinb(n11190), .dout(n11193));
  jor  g11130(.dina(n7177), .dinb(n9919), .dout(n11194));
  jor  g11131(.dina(n9918), .dinb(n3516), .dout(n11195));
  jor  g11132(.dina(n10826), .dinb(n3684), .dout(n11196));
  jor  g11133(.dina(n10351), .dinb(n3414), .dout(n11197));
  jand g11134(.dina(n11197), .dinb(n11196), .dout(n11198));
  jand g11135(.dina(n11198), .dinb(n11195), .dout(n11199));
  jand g11136(.dina(n11199), .dinb(n11194), .dout(n11200));
  jxor g11137(.dina(n11200), .dinb(\a[5] ), .dout(n11201));
  jand g11138(.dina(n10689), .dinb(\a[8] ), .dout(n11202));
  jxor g11139(.dina(n11202), .dinb(n10687), .dout(n11203));
  jnot g11140(.din(n11203), .dout(n11204));
  jor  g11141(.dina(n11204), .dinb(n11201), .dout(n11205));
  jand g11142(.dina(n8004), .dinb(n67), .dout(n11206));
  jand g11143(.dina(n10350), .dinb(n7411), .dout(n11207));
  jand g11144(.dina(n10827), .dinb(n7405), .dout(n11208));
  jor  g11145(.dina(n11208), .dinb(n11207), .dout(n11209));
  jor  g11146(.dina(n11209), .dinb(n11206), .dout(n11210));
  jnot g11147(.din(n11210), .dout(n11211));
  jand g11148(.dina(n7411), .dinb(n65), .dout(n11212));
  jnot g11149(.din(n11212), .dout(n11213));
  jand g11150(.dina(n11213), .dinb(\a[5] ), .dout(n11214));
  jand g11151(.dina(n11214), .dinb(n11211), .dout(n11215));
  jand g11152(.dina(n7407), .dinb(n67), .dout(n11216));
  jand g11153(.dina(n10827), .dinb(n7326), .dout(n11217));
  jand g11154(.dina(n9917), .dinb(n7411), .dout(n11218));
  jand g11155(.dina(n10350), .dinb(n7405), .dout(n11219));
  jor  g11156(.dina(n11219), .dinb(n11218), .dout(n11220));
  jor  g11157(.dina(n11220), .dinb(n11217), .dout(n11221));
  jor  g11158(.dina(n11221), .dinb(n11216), .dout(n11222));
  jnot g11159(.din(n11222), .dout(n11223));
  jand g11160(.dina(n11223), .dinb(n11215), .dout(n11224));
  jand g11161(.dina(n11224), .dinb(n10689), .dout(n11225));
  jnot g11162(.din(n11225), .dout(n11226));
  jor  g11163(.dina(n7466), .dinb(n9919), .dout(n11227));
  jor  g11164(.dina(n10351), .dinb(n3516), .dout(n11228));
  jor  g11165(.dina(n10826), .dinb(n3414), .dout(n11229));
  jor  g11166(.dina(n9918), .dinb(n3677), .dout(n11230));
  jand g11167(.dina(n11230), .dinb(n11229), .dout(n11231));
  jand g11168(.dina(n11231), .dinb(n11228), .dout(n11232));
  jand g11169(.dina(n11232), .dinb(n11227), .dout(n11233));
  jxor g11170(.dina(n11233), .dinb(\a[5] ), .dout(n11234));
  jxor g11171(.dina(n11224), .dinb(n10689), .dout(n11235));
  jnot g11172(.din(n11235), .dout(n11236));
  jor  g11173(.dina(n11236), .dinb(n11234), .dout(n11237));
  jand g11174(.dina(n11237), .dinb(n11226), .dout(n11238));
  jxor g11175(.dina(n11203), .dinb(n11201), .dout(n11239));
  jor  g11176(.dina(n11239), .dinb(n11238), .dout(n11240));
  jand g11177(.dina(n11240), .dinb(n11205), .dout(n11241));
  jnot g11178(.din(n11241), .dout(n11242));
  jxor g11179(.dina(n11192), .dinb(n11190), .dout(n11243));
  jand g11180(.dina(n11243), .dinb(n11242), .dout(n11244));
  jor  g11181(.dina(n11244), .dinb(n11193), .dout(n11245));
  jxor g11182(.dina(n11181), .dinb(n11180), .dout(n11246));
  jand g11183(.dina(n11246), .dinb(n11245), .dout(n11247));
  jor  g11184(.dina(n11247), .dinb(n11182), .dout(n11248));
  jxor g11185(.dina(n11170), .dinb(n11169), .dout(n11249));
  jand g11186(.dina(n11249), .dinb(n11248), .dout(n11250));
  jor  g11187(.dina(n11250), .dinb(n11171), .dout(n11251));
  jxor g11188(.dina(n11159), .dinb(n11151), .dout(n11252));
  jand g11189(.dina(n11252), .dinb(n11251), .dout(n11253));
  jnot g11190(.din(n11253), .dout(n11254));
  jand g11191(.dina(n11254), .dinb(n11160), .dout(n11255));
  jnot g11192(.din(n11255), .dout(n11256));
  jxor g11193(.dina(n11148), .dinb(n11140), .dout(n11257));
  jand g11194(.dina(n11257), .dinb(n11256), .dout(n11258));
  jnot g11195(.din(n11258), .dout(n11259));
  jand g11196(.dina(n11259), .dinb(n11149), .dout(n11260));
  jxor g11197(.dina(n11137), .dinb(n11129), .dout(n11261));
  jnot g11198(.din(n11261), .dout(n11262));
  jor  g11199(.dina(n11262), .dinb(n11260), .dout(n11263));
  jand g11200(.dina(n11263), .dinb(n11138), .dout(n11264));
  jnot g11201(.din(n11264), .dout(n11265));
  jxor g11202(.dina(n11126), .dinb(n11125), .dout(n11266));
  jand g11203(.dina(n11266), .dinb(n11265), .dout(n11267));
  jor  g11204(.dina(n11267), .dinb(n11127), .dout(n11268));
  jxor g11205(.dina(n11115), .dinb(n11114), .dout(n11269));
  jand g11206(.dina(n11269), .dinb(n11268), .dout(n11270));
  jor  g11207(.dina(n11270), .dinb(n11116), .dout(n11271));
  jxor g11208(.dina(n11104), .dinb(n11103), .dout(n11272));
  jand g11209(.dina(n11272), .dinb(n11271), .dout(n11273));
  jor  g11210(.dina(n11273), .dinb(n11105), .dout(n11274));
  jxor g11211(.dina(n11093), .dinb(n11085), .dout(n11275));
  jand g11212(.dina(n11275), .dinb(n11274), .dout(n11276));
  jnot g11213(.din(n11276), .dout(n11277));
  jand g11214(.dina(n11277), .dinb(n11094), .dout(n11278));
  jnot g11215(.din(n11278), .dout(n11279));
  jxor g11216(.dina(n11082), .dinb(n11074), .dout(n11280));
  jand g11217(.dina(n11280), .dinb(n11279), .dout(n11281));
  jnot g11218(.din(n11281), .dout(n11282));
  jand g11219(.dina(n11282), .dinb(n11083), .dout(n11283));
  jxor g11220(.dina(n11071), .dinb(n11063), .dout(n11284));
  jnot g11221(.din(n11284), .dout(n11285));
  jor  g11222(.dina(n11285), .dinb(n11283), .dout(n11286));
  jand g11223(.dina(n11286), .dinb(n11072), .dout(n11287));
  jnot g11224(.din(n11287), .dout(n11288));
  jxor g11225(.dina(n11060), .dinb(n11059), .dout(n11289));
  jand g11226(.dina(n11289), .dinb(n11288), .dout(n11290));
  jor  g11227(.dina(n11290), .dinb(n11061), .dout(n11291));
  jxor g11228(.dina(n11049), .dinb(n11048), .dout(n11292));
  jand g11229(.dina(n11292), .dinb(n11291), .dout(n11293));
  jor  g11230(.dina(n11293), .dinb(n11050), .dout(n11294));
  jxor g11231(.dina(n11038), .dinb(n11037), .dout(n11295));
  jand g11232(.dina(n11295), .dinb(n11294), .dout(n11296));
  jor  g11233(.dina(n11296), .dinb(n11039), .dout(n11297));
  jxor g11234(.dina(n11027), .dinb(n11019), .dout(n11298));
  jand g11235(.dina(n11298), .dinb(n11297), .dout(n11299));
  jnot g11236(.din(n11299), .dout(n11300));
  jand g11237(.dina(n11300), .dinb(n11028), .dout(n11301));
  jxor g11238(.dina(n11016), .dinb(n11008), .dout(n11302));
  jnot g11239(.din(n11302), .dout(n11303));
  jor  g11240(.dina(n11303), .dinb(n11301), .dout(n11304));
  jand g11241(.dina(n11304), .dinb(n11017), .dout(n11305));
  jxor g11242(.dina(n11005), .dinb(n10997), .dout(n11306));
  jnot g11243(.din(n11306), .dout(n11307));
  jor  g11244(.dina(n11307), .dinb(n11305), .dout(n11308));
  jand g11245(.dina(n11308), .dinb(n11006), .dout(n11309));
  jnot g11246(.din(n11309), .dout(n11310));
  jxor g11247(.dina(n10994), .dinb(n10993), .dout(n11311));
  jand g11248(.dina(n11311), .dinb(n11310), .dout(n11312));
  jor  g11249(.dina(n11312), .dinb(n10995), .dout(n11313));
  jxor g11250(.dina(n10983), .dinb(n10982), .dout(n11314));
  jand g11251(.dina(n11314), .dinb(n11313), .dout(n11315));
  jor  g11252(.dina(n11315), .dinb(n10984), .dout(n11316));
  jxor g11253(.dina(n10972), .dinb(n10971), .dout(n11317));
  jand g11254(.dina(n11317), .dinb(n11316), .dout(n11318));
  jor  g11255(.dina(n11318), .dinb(n10973), .dout(n11319));
  jnot g11256(.din(n11319), .dout(n11320));
  jxor g11257(.dina(n10961), .dinb(n10952), .dout(n11321));
  jor  g11258(.dina(n11321), .dinb(n11320), .dout(n11322));
  jand g11259(.dina(n11322), .dinb(n10962), .dout(n11323));
  jxor g11260(.dina(n10950), .dinb(n10941), .dout(n11324));
  jor  g11261(.dina(n11324), .dinb(n11323), .dout(n11325));
  jand g11262(.dina(n11325), .dinb(n10951), .dout(n11326));
  jxor g11263(.dina(n10938), .dinb(n10937), .dout(n11327));
  jnot g11264(.din(n11327), .dout(n11328));
  jor  g11265(.dina(n11328), .dinb(n11326), .dout(n11329));
  jand g11266(.dina(n11329), .dinb(n10940), .dout(n11330));
  jxor g11267(.dina(n10926), .dinb(n10925), .dout(n11331));
  jnot g11268(.din(n11331), .dout(n11332));
  jor  g11269(.dina(n11332), .dinb(n11330), .dout(n11333));
  jand g11270(.dina(n11333), .dinb(n10928), .dout(n11334));
  jxor g11271(.dina(n10914), .dinb(n10913), .dout(n11335));
  jnot g11272(.din(n11335), .dout(n11336));
  jor  g11273(.dina(n11336), .dinb(n11334), .dout(n11337));
  jand g11274(.dina(n11337), .dinb(n10916), .dout(n11338));
  jxor g11275(.dina(n10902), .dinb(n10901), .dout(n11339));
  jnot g11276(.din(n11339), .dout(n11340));
  jor  g11277(.dina(n11340), .dinb(n11338), .dout(n11341));
  jand g11278(.dina(n11341), .dinb(n10904), .dout(n11342));
  jxor g11279(.dina(n10890), .dinb(n10889), .dout(n11343));
  jnot g11280(.din(n11343), .dout(n11344));
  jor  g11281(.dina(n11344), .dinb(n11342), .dout(n11345));
  jand g11282(.dina(n11345), .dinb(n10892), .dout(n11346));
  jnot g11283(.din(n11346), .dout(n11347));
  jxor g11284(.dina(n10879), .dinb(n10878), .dout(n11348));
  jand g11285(.dina(n11348), .dinb(n11347), .dout(n11349));
  jor  g11286(.dina(n11349), .dinb(n10880), .dout(n11350));
  jxor g11287(.dina(n10862), .dinb(n10861), .dout(n11351));
  jand g11288(.dina(n11351), .dinb(n11350), .dout(n11352));
  jnot g11289(.din(n11352), .dout(n11353));
  jxor g11290(.dina(n11351), .dinb(n11350), .dout(n11354));
  jnot g11291(.din(n11354), .dout(n11355));
  jxor g11292(.dina(n11348), .dinb(n11346), .dout(n11356));
  jor  g11293(.dina(n10847), .dinb(n4731), .dout(n11357));
  jor  g11294(.dina(n10845), .dinb(n4597), .dout(n11358));
  jand g11295(.dina(\a[1] ), .dinb(n10840), .dout(n11359));
  jnot g11296(.din(n11359), .dout(n11360));
  jor  g11297(.dina(n11360), .dinb(n4630), .dout(n11361));
  jand g11298(.dina(n11361), .dinb(n11358), .dout(n11362));
  jand g11299(.dina(n11362), .dinb(n11357), .dout(n11363));
  jxor g11300(.dina(n11363), .dinb(\a[2] ), .dout(n11364));
  jor  g11301(.dina(n11364), .dinb(n11356), .dout(n11365));
  jxor g11302(.dina(n11344), .dinb(n11342), .dout(n11366));
  jnot g11303(.din(n11366), .dout(n11367));
  jand g11304(.dina(n10846), .dinb(n4636), .dout(n11368));
  jand g11305(.dina(n10844), .dinb(n4451), .dout(n11369));
  jand g11306(.dina(n11359), .dinb(n4598), .dout(n11370));
  jnot g11307(.din(n10843), .dout(n11371));
  jand g11308(.dina(n11371), .dinb(\a[0] ), .dout(n11372));
  jand g11309(.dina(n11372), .dinb(n4631), .dout(n11373));
  jor  g11310(.dina(n11373), .dinb(n11370), .dout(n11374));
  jor  g11311(.dina(n11374), .dinb(n11369), .dout(n11375));
  jor  g11312(.dina(n11375), .dinb(n11368), .dout(n11376));
  jxor g11313(.dina(n11376), .dinb(n6600), .dout(n11377));
  jor  g11314(.dina(n11377), .dinb(n11367), .dout(n11378));
  jxor g11315(.dina(n11340), .dinb(n11338), .dout(n11379));
  jnot g11316(.din(n11379), .dout(n11380));
  jand g11317(.dina(n10846), .dinb(n4752), .dout(n11381));
  jand g11318(.dina(n11359), .dinb(n4451), .dout(n11382));
  jand g11319(.dina(n10844), .dinb(n4358), .dout(n11383));
  jand g11320(.dina(n11372), .dinb(n4598), .dout(n11384));
  jor  g11321(.dina(n11384), .dinb(n11383), .dout(n11385));
  jor  g11322(.dina(n11385), .dinb(n11382), .dout(n11386));
  jor  g11323(.dina(n11386), .dinb(n11381), .dout(n11387));
  jxor g11324(.dina(n11387), .dinb(n6600), .dout(n11388));
  jor  g11325(.dina(n11388), .dinb(n11380), .dout(n11389));
  jxor g11326(.dina(n11336), .dinb(n11334), .dout(n11390));
  jnot g11327(.din(n11390), .dout(n11391));
  jand g11328(.dina(n10846), .dinb(n4446), .dout(n11392));
  jand g11329(.dina(n11372), .dinb(n4451), .dout(n11393));
  jand g11330(.dina(n11359), .dinb(n4358), .dout(n11394));
  jand g11331(.dina(n10844), .dinb(n3853), .dout(n11395));
  jor  g11332(.dina(n11395), .dinb(n11394), .dout(n11396));
  jor  g11333(.dina(n11396), .dinb(n11393), .dout(n11397));
  jor  g11334(.dina(n11397), .dinb(n11392), .dout(n11398));
  jxor g11335(.dina(n11398), .dinb(n6600), .dout(n11399));
  jor  g11336(.dina(n11399), .dinb(n11391), .dout(n11400));
  jxor g11337(.dina(n11332), .dinb(n11330), .dout(n11401));
  jnot g11338(.din(n11401), .dout(n11402));
  jand g11339(.dina(n10846), .dinb(n4545), .dout(n11403));
  jand g11340(.dina(n10844), .dinb(n922), .dout(n11404));
  jand g11341(.dina(n11359), .dinb(n3853), .dout(n11405));
  jand g11342(.dina(n11372), .dinb(n4358), .dout(n11406));
  jor  g11343(.dina(n11406), .dinb(n11405), .dout(n11407));
  jor  g11344(.dina(n11407), .dinb(n11404), .dout(n11408));
  jor  g11345(.dina(n11408), .dinb(n11403), .dout(n11409));
  jxor g11346(.dina(n11409), .dinb(n6600), .dout(n11410));
  jor  g11347(.dina(n11410), .dinb(n11402), .dout(n11411));
  jxor g11348(.dina(n11410), .dinb(n11401), .dout(n11412));
  jxor g11349(.dina(n11324), .dinb(n11323), .dout(n11413));
  jnot g11350(.din(n11413), .dout(n11414));
  jxor g11351(.dina(n11321), .dinb(n11320), .dout(n11415));
  jnot g11352(.din(n11415), .dout(n11416));
  jxor g11353(.dina(n11317), .dinb(n11316), .dout(n11417));
  jnot g11354(.din(n11417), .dout(n11418));
  jxor g11355(.dina(n11314), .dinb(n11313), .dout(n11419));
  jnot g11356(.din(n11419), .dout(n11420));
  jxor g11357(.dina(n11307), .dinb(n11305), .dout(n11421));
  jnot g11358(.din(n11421), .dout(n11422));
  jxor g11359(.dina(n11303), .dinb(n11301), .dout(n11423));
  jnot g11360(.din(n11423), .dout(n11424));
  jxor g11361(.dina(n11298), .dinb(n11297), .dout(n11425));
  jnot g11362(.din(n11425), .dout(n11426));
  jxor g11363(.dina(n11295), .dinb(n11294), .dout(n11427));
  jnot g11364(.din(n11427), .dout(n11428));
  jxor g11365(.dina(n11292), .dinb(n11291), .dout(n11429));
  jnot g11366(.din(n11429), .dout(n11430));
  jxor g11367(.dina(n11285), .dinb(n11283), .dout(n11431));
  jnot g11368(.din(n11431), .dout(n11432));
  jxor g11369(.dina(n11280), .dinb(n11279), .dout(n11433));
  jnot g11370(.din(n11433), .dout(n11434));
  jxor g11371(.dina(n11275), .dinb(n11274), .dout(n11435));
  jnot g11372(.din(n11435), .dout(n11436));
  jxor g11373(.dina(n11272), .dinb(n11271), .dout(n11437));
  jnot g11374(.din(n11437), .dout(n11438));
  jxor g11375(.dina(n11269), .dinb(n11268), .dout(n11439));
  jnot g11376(.din(n11439), .dout(n11440));
  jxor g11377(.dina(n11262), .dinb(n11260), .dout(n11441));
  jnot g11378(.din(n11441), .dout(n11442));
  jxor g11379(.dina(n11257), .dinb(n11256), .dout(n11443));
  jnot g11380(.din(n11443), .dout(n11444));
  jxor g11381(.dina(n11252), .dinb(n11251), .dout(n11445));
  jnot g11382(.din(n11445), .dout(n11446));
  jxor g11383(.dina(n11249), .dinb(n11248), .dout(n11447));
  jnot g11384(.din(n11447), .dout(n11448));
  jxor g11385(.dina(n11246), .dinb(n11245), .dout(n11449));
  jnot g11386(.din(n11449), .dout(n11450));
  jxor g11387(.dina(n11239), .dinb(n11238), .dout(n11451));
  jnot g11388(.din(n11451), .dout(n11452));
  jnot g11389(.din(n11215), .dout(n11453));
  jand g11390(.dina(n11453), .dinb(\a[5] ), .dout(n11454));
  jxor g11391(.dina(n11454), .dinb(n11223), .dout(n11455));
  jor  g11392(.dina(n10847), .dinb(n7177), .dout(n11456));
  jor  g11393(.dina(n10845), .dinb(n3516), .dout(n11457));
  jnot g11394(.din(n11372), .dout(n11458));
  jor  g11395(.dina(n11458), .dinb(n3684), .dout(n11459));
  jor  g11396(.dina(n11360), .dinb(n3414), .dout(n11460));
  jand g11397(.dina(n11460), .dinb(n11459), .dout(n11461));
  jand g11398(.dina(n11461), .dinb(n11457), .dout(n11462));
  jand g11399(.dina(n11462), .dinb(n11456), .dout(n11463));
  jxor g11400(.dina(n11463), .dinb(\a[2] ), .dout(n11464));
  jand g11401(.dina(n11371), .dinb(n10842), .dout(n11465));
  jnot g11402(.din(n11465), .dout(n11466));
  jand g11403(.dina(n11372), .dinb(n7326), .dout(n11467));
  jor  g11404(.dina(n11467), .dinb(n7405), .dout(n11468));
  jand g11405(.dina(n11458), .dinb(n11360), .dout(n11469));
  jnot g11406(.din(n11469), .dout(n11470));
  jand g11407(.dina(n11470), .dinb(n11468), .dout(n11471));
  jand g11408(.dina(n10846), .dinb(n7405), .dout(n11472));
  jor  g11409(.dina(n11472), .dinb(n7411), .dout(n11473));
  jor  g11410(.dina(n11473), .dinb(n11471), .dout(n11474));
  jand g11411(.dina(n11474), .dinb(n11466), .dout(n11475));
  jand g11412(.dina(n10846), .dinb(n7407), .dout(n11476));
  jor  g11413(.dina(n11476), .dinb(n6600), .dout(n11477));
  jor  g11414(.dina(n11477), .dinb(n11475), .dout(n11478));
  jand g11415(.dina(n11478), .dinb(n11213), .dout(n11479));
  jor  g11416(.dina(n10847), .dinb(n7466), .dout(n11481));
  jor  g11417(.dina(n11360), .dinb(n3516), .dout(n11482));
  jor  g11418(.dina(n11458), .dinb(n3414), .dout(n11483));
  jor  g11419(.dina(n10845), .dinb(n3677), .dout(n11484));
  jand g11420(.dina(n11484), .dinb(n11483), .dout(n11485));
  jand g11421(.dina(n11485), .dinb(n11482), .dout(n11486));
  jand g11422(.dina(n11486), .dinb(n11481), .dout(n11487));
  jxor g11423(.dina(n11487), .dinb(\a[2] ), .dout(n11488));
  jor  g11424(.dina(n11488), .dinb(n11479), .dout(n11490));
  jor  g11425(.dina(n11490), .dinb(n11464), .dout(n11491));
  jand g11426(.dina(n11490), .dinb(n11464), .dout(n11492));
  jand g11427(.dina(n11212), .dinb(\a[5] ), .dout(n11493));
  jxor g11428(.dina(n11493), .dinb(n11210), .dout(n11494));
  jnot g11429(.din(n11494), .dout(n11495));
  jor  g11430(.dina(n11495), .dinb(n11492), .dout(n11496));
  jand g11431(.dina(n11496), .dinb(n11491), .dout(n11497));
  jand g11432(.dina(n11497), .dinb(n11455), .dout(n11498));
  jor  g11433(.dina(n10847), .dinb(n7131), .dout(n11499));
  jor  g11434(.dina(n11458), .dinb(n7962), .dout(n11500));
  jor  g11435(.dina(n10845), .dinb(n3414), .dout(n11501));
  jor  g11436(.dina(n11360), .dinb(n3684), .dout(n11502));
  jand g11437(.dina(n11502), .dinb(n11501), .dout(n11503));
  jand g11438(.dina(n11503), .dinb(n11500), .dout(n11504));
  jand g11439(.dina(n11504), .dinb(n11499), .dout(n11505));
  jxor g11440(.dina(n11505), .dinb(n6600), .dout(n11506));
  jnot g11441(.din(n11506), .dout(n11507));
  jor  g11442(.dina(n11507), .dinb(n11498), .dout(n11508));
  jor  g11443(.dina(n11497), .dinb(n11455), .dout(n11509));
  jor  g11444(.dina(n10847), .dinb(n7076), .dout(n11510));
  jor  g11445(.dina(n11360), .dinb(n7962), .dout(n11511));
  jor  g11446(.dina(n11458), .dinb(n3182), .dout(n11512));
  jor  g11447(.dina(n10845), .dinb(n3684), .dout(n11513));
  jand g11448(.dina(n11513), .dinb(n11512), .dout(n11514));
  jand g11449(.dina(n11514), .dinb(n11511), .dout(n11515));
  jand g11450(.dina(n11515), .dinb(n11510), .dout(n11516));
  jxor g11451(.dina(n11516), .dinb(\a[2] ), .dout(n11517));
  jxor g11452(.dina(n11235), .dinb(n11234), .dout(n11518));
  jor  g11453(.dina(n11518), .dinb(n11517), .dout(n11519));
  jand g11454(.dina(n11519), .dinb(n11509), .dout(n11520));
  jand g11455(.dina(n11520), .dinb(n11508), .dout(n11521));
  jand g11456(.dina(n11518), .dinb(n11517), .dout(n11522));
  jor  g11457(.dina(n11522), .dinb(n11521), .dout(n11523));
  jand g11458(.dina(n11523), .dinb(n11452), .dout(n11524));
  jor  g11459(.dina(n10847), .dinb(n7031), .dout(n11525));
  jor  g11460(.dina(n11458), .dinb(n3085), .dout(n11526));
  jor  g11461(.dina(n10845), .dinb(n7962), .dout(n11527));
  jor  g11462(.dina(n11360), .dinb(n3182), .dout(n11528));
  jand g11463(.dina(n11528), .dinb(n11527), .dout(n11529));
  jand g11464(.dina(n11529), .dinb(n11526), .dout(n11530));
  jand g11465(.dina(n11530), .dinb(n11525), .dout(n11531));
  jxor g11466(.dina(n11531), .dinb(n6600), .dout(n11532));
  jnot g11467(.din(n11532), .dout(n11533));
  jor  g11468(.dina(n11533), .dinb(n11524), .dout(n11534));
  jor  g11469(.dina(n11523), .dinb(n11452), .dout(n11535));
  jor  g11470(.dina(n10847), .dinb(n6681), .dout(n11536));
  jor  g11471(.dina(n11360), .dinb(n3085), .dout(n11537));
  jor  g11472(.dina(n11458), .dinb(n2990), .dout(n11538));
  jor  g11473(.dina(n10845), .dinb(n3182), .dout(n11539));
  jand g11474(.dina(n11539), .dinb(n11538), .dout(n11540));
  jand g11475(.dina(n11540), .dinb(n11537), .dout(n11541));
  jand g11476(.dina(n11541), .dinb(n11536), .dout(n11542));
  jxor g11477(.dina(n11542), .dinb(\a[2] ), .dout(n11543));
  jxor g11478(.dina(n11243), .dinb(n11241), .dout(n11544));
  jor  g11479(.dina(n11544), .dinb(n11543), .dout(n11545));
  jand g11480(.dina(n11545), .dinb(n11535), .dout(n11546));
  jand g11481(.dina(n11546), .dinb(n11534), .dout(n11547));
  jand g11482(.dina(n11544), .dinb(n11543), .dout(n11548));
  jor  g11483(.dina(n11548), .dinb(n11547), .dout(n11549));
  jor  g11484(.dina(n11549), .dinb(n11450), .dout(n11550));
  jor  g11485(.dina(n10847), .dinb(n6988), .dout(n11551));
  jor  g11486(.dina(n10845), .dinb(n3085), .dout(n11552));
  jor  g11487(.dina(n11458), .dinb(n2953), .dout(n11553));
  jor  g11488(.dina(n11360), .dinb(n2990), .dout(n11554));
  jand g11489(.dina(n11554), .dinb(n11553), .dout(n11555));
  jand g11490(.dina(n11555), .dinb(n11552), .dout(n11556));
  jand g11491(.dina(n11556), .dinb(n11551), .dout(n11557));
  jxor g11492(.dina(n11557), .dinb(\a[2] ), .dout(n11558));
  jand g11493(.dina(n11558), .dinb(n11550), .dout(n11559));
  jand g11494(.dina(n11549), .dinb(n11450), .dout(n11560));
  jor  g11495(.dina(n11560), .dinb(n11559), .dout(n11561));
  jor  g11496(.dina(n11561), .dinb(n11448), .dout(n11562));
  jor  g11497(.dina(n10847), .dinb(n6976), .dout(n11563));
  jor  g11498(.dina(n11360), .dinb(n2953), .dout(n11564));
  jor  g11499(.dina(n10845), .dinb(n2990), .dout(n11565));
  jor  g11500(.dina(n11458), .dinb(n2866), .dout(n11566));
  jand g11501(.dina(n11566), .dinb(n11565), .dout(n11567));
  jand g11502(.dina(n11567), .dinb(n11564), .dout(n11568));
  jand g11503(.dina(n11568), .dinb(n11563), .dout(n11569));
  jxor g11504(.dina(n11569), .dinb(\a[2] ), .dout(n11570));
  jand g11505(.dina(n11570), .dinb(n11562), .dout(n11571));
  jand g11506(.dina(n11561), .dinb(n11448), .dout(n11572));
  jor  g11507(.dina(n11572), .dinb(n11571), .dout(n11573));
  jor  g11508(.dina(n11573), .dinb(n11446), .dout(n11574));
  jand g11509(.dina(n11573), .dinb(n11446), .dout(n11575));
  jnot g11510(.din(n6706), .dout(n11576));
  jor  g11511(.dina(n10847), .dinb(n11576), .dout(n11577));
  jor  g11512(.dina(n11458), .dinb(n2807), .dout(n11578));
  jor  g11513(.dina(n10845), .dinb(n2953), .dout(n11579));
  jor  g11514(.dina(n11360), .dinb(n2866), .dout(n11580));
  jand g11515(.dina(n11580), .dinb(n11579), .dout(n11581));
  jand g11516(.dina(n11581), .dinb(n11578), .dout(n11582));
  jand g11517(.dina(n11582), .dinb(n11577), .dout(n11583));
  jxor g11518(.dina(n11583), .dinb(\a[2] ), .dout(n11584));
  jor  g11519(.dina(n11584), .dinb(n11575), .dout(n11585));
  jand g11520(.dina(n11585), .dinb(n11574), .dout(n11586));
  jor  g11521(.dina(n11586), .dinb(n11444), .dout(n11587));
  jand g11522(.dina(n11586), .dinb(n11444), .dout(n11588));
  jnot g11523(.din(n6439), .dout(n11589));
  jor  g11524(.dina(n10847), .dinb(n11589), .dout(n11590));
  jor  g11525(.dina(n11360), .dinb(n2807), .dout(n11591));
  jor  g11526(.dina(n11458), .dinb(n2731), .dout(n11592));
  jor  g11527(.dina(n10845), .dinb(n2866), .dout(n11593));
  jand g11528(.dina(n11593), .dinb(n11592), .dout(n11594));
  jand g11529(.dina(n11594), .dinb(n11591), .dout(n11595));
  jand g11530(.dina(n11595), .dinb(n11590), .dout(n11596));
  jxor g11531(.dina(n11596), .dinb(n6600), .dout(n11597));
  jnot g11532(.din(n11597), .dout(n11598));
  jor  g11533(.dina(n11598), .dinb(n11588), .dout(n11599));
  jand g11534(.dina(n11599), .dinb(n11587), .dout(n11600));
  jand g11535(.dina(n11600), .dinb(n11442), .dout(n11601));
  jnot g11536(.din(n6591), .dout(n11602));
  jor  g11537(.dina(n10847), .dinb(n11602), .dout(n11603));
  jor  g11538(.dina(n11458), .dinb(n2694), .dout(n11604));
  jor  g11539(.dina(n10845), .dinb(n2807), .dout(n11605));
  jor  g11540(.dina(n11360), .dinb(n2731), .dout(n11606));
  jand g11541(.dina(n11606), .dinb(n11605), .dout(n11607));
  jand g11542(.dina(n11607), .dinb(n11604), .dout(n11608));
  jand g11543(.dina(n11608), .dinb(n11603), .dout(n11609));
  jxor g11544(.dina(n11609), .dinb(n6600), .dout(n11610));
  jnot g11545(.din(n11610), .dout(n11611));
  jor  g11546(.dina(n11611), .dinb(n11601), .dout(n11612));
  jor  g11547(.dina(n11600), .dinb(n11442), .dout(n11613));
  jor  g11548(.dina(n10847), .dinb(n6464), .dout(n11614));
  jor  g11549(.dina(n11458), .dinb(n2601), .dout(n11615));
  jor  g11550(.dina(n11360), .dinb(n2694), .dout(n11616));
  jor  g11551(.dina(n10845), .dinb(n2731), .dout(n11617));
  jand g11552(.dina(n11617), .dinb(n11616), .dout(n11618));
  jand g11553(.dina(n11618), .dinb(n11615), .dout(n11619));
  jand g11554(.dina(n11619), .dinb(n11614), .dout(n11620));
  jxor g11555(.dina(n11620), .dinb(\a[2] ), .dout(n11621));
  jxor g11556(.dina(n11266), .dinb(n11264), .dout(n11622));
  jor  g11557(.dina(n11622), .dinb(n11621), .dout(n11623));
  jand g11558(.dina(n11623), .dinb(n11613), .dout(n11624));
  jand g11559(.dina(n11624), .dinb(n11612), .dout(n11625));
  jand g11560(.dina(n11622), .dinb(n11621), .dout(n11626));
  jor  g11561(.dina(n11626), .dinb(n11625), .dout(n11627));
  jor  g11562(.dina(n11627), .dinb(n11440), .dout(n11628));
  jnot g11563(.din(n6050), .dout(n11629));
  jor  g11564(.dina(n10847), .dinb(n11629), .dout(n11630));
  jor  g11565(.dina(n11360), .dinb(n2601), .dout(n11631));
  jor  g11566(.dina(n10845), .dinb(n2694), .dout(n11632));
  jor  g11567(.dina(n11458), .dinb(n2496), .dout(n11633));
  jand g11568(.dina(n11633), .dinb(n11632), .dout(n11634));
  jand g11569(.dina(n11634), .dinb(n11631), .dout(n11635));
  jand g11570(.dina(n11635), .dinb(n11630), .dout(n11636));
  jxor g11571(.dina(n11636), .dinb(\a[2] ), .dout(n11637));
  jand g11572(.dina(n11637), .dinb(n11628), .dout(n11638));
  jand g11573(.dina(n11627), .dinb(n11440), .dout(n11639));
  jor  g11574(.dina(n11639), .dinb(n11638), .dout(n11640));
  jor  g11575(.dina(n11640), .dinb(n11438), .dout(n11641));
  jnot g11576(.din(n6247), .dout(n11642));
  jor  g11577(.dina(n10847), .dinb(n11642), .dout(n11643));
  jor  g11578(.dina(n11458), .dinb(n2410), .dout(n11644));
  jor  g11579(.dina(n10845), .dinb(n2601), .dout(n11645));
  jor  g11580(.dina(n11360), .dinb(n2496), .dout(n11646));
  jand g11581(.dina(n11646), .dinb(n11645), .dout(n11647));
  jand g11582(.dina(n11647), .dinb(n11644), .dout(n11648));
  jand g11583(.dina(n11648), .dinb(n11643), .dout(n11649));
  jxor g11584(.dina(n11649), .dinb(\a[2] ), .dout(n11650));
  jand g11585(.dina(n11650), .dinb(n11641), .dout(n11651));
  jand g11586(.dina(n11640), .dinb(n11438), .dout(n11652));
  jor  g11587(.dina(n11652), .dinb(n11651), .dout(n11653));
  jor  g11588(.dina(n11653), .dinb(n11436), .dout(n11654));
  jand g11589(.dina(n11653), .dinb(n11436), .dout(n11655));
  jnot g11590(.din(n5861), .dout(n11656));
  jor  g11591(.dina(n10847), .dinb(n11656), .dout(n11657));
  jor  g11592(.dina(n11360), .dinb(n2410), .dout(n11658));
  jor  g11593(.dina(n11458), .dinb(n2342), .dout(n11659));
  jor  g11594(.dina(n10845), .dinb(n2496), .dout(n11660));
  jand g11595(.dina(n11660), .dinb(n11659), .dout(n11661));
  jand g11596(.dina(n11661), .dinb(n11658), .dout(n11662));
  jand g11597(.dina(n11662), .dinb(n11657), .dout(n11663));
  jxor g11598(.dina(n11663), .dinb(n6600), .dout(n11664));
  jnot g11599(.din(n11664), .dout(n11665));
  jor  g11600(.dina(n11665), .dinb(n11655), .dout(n11666));
  jand g11601(.dina(n11666), .dinb(n11654), .dout(n11667));
  jor  g11602(.dina(n11667), .dinb(n11434), .dout(n11668));
  jand g11603(.dina(n11667), .dinb(n11434), .dout(n11669));
  jnot g11604(.din(n5844), .dout(n11670));
  jor  g11605(.dina(n10847), .dinb(n11670), .dout(n11671));
  jor  g11606(.dina(n10845), .dinb(n2410), .dout(n11672));
  jor  g11607(.dina(n11458), .dinb(n2236), .dout(n11673));
  jor  g11608(.dina(n11360), .dinb(n2342), .dout(n11674));
  jand g11609(.dina(n11674), .dinb(n11673), .dout(n11675));
  jand g11610(.dina(n11675), .dinb(n11672), .dout(n11676));
  jand g11611(.dina(n11676), .dinb(n11671), .dout(n11677));
  jxor g11612(.dina(n11677), .dinb(n6600), .dout(n11678));
  jnot g11613(.din(n11678), .dout(n11679));
  jor  g11614(.dina(n11679), .dinb(n11669), .dout(n11680));
  jand g11615(.dina(n11680), .dinb(n11668), .dout(n11681));
  jand g11616(.dina(n11681), .dinb(n11432), .dout(n11682));
  jnot g11617(.din(n5607), .dout(n11683));
  jor  g11618(.dina(n10847), .dinb(n11683), .dout(n11684));
  jor  g11619(.dina(n11360), .dinb(n2236), .dout(n11685));
  jor  g11620(.dina(n10845), .dinb(n2342), .dout(n11686));
  jor  g11621(.dina(n11458), .dinb(n2127), .dout(n11687));
  jand g11622(.dina(n11687), .dinb(n11686), .dout(n11688));
  jand g11623(.dina(n11688), .dinb(n11685), .dout(n11689));
  jand g11624(.dina(n11689), .dinb(n11684), .dout(n11690));
  jxor g11625(.dina(n11690), .dinb(n6600), .dout(n11691));
  jnot g11626(.din(n11691), .dout(n11692));
  jor  g11627(.dina(n11692), .dinb(n11682), .dout(n11693));
  jor  g11628(.dina(n11681), .dinb(n11432), .dout(n11694));
  jand g11629(.dina(n10846), .dinb(n5624), .dout(n11695));
  jand g11630(.dina(n10844), .dinb(n2237), .dout(n11696));
  jand g11631(.dina(n11359), .dinb(n2128), .dout(n11697));
  jand g11632(.dina(n11372), .dinb(n2067), .dout(n11698));
  jor  g11633(.dina(n11698), .dinb(n11697), .dout(n11699));
  jor  g11634(.dina(n11699), .dinb(n11696), .dout(n11700));
  jor  g11635(.dina(n11700), .dinb(n11695), .dout(n11701));
  jxor g11636(.dina(n11701), .dinb(n6600), .dout(n11702));
  jxor g11637(.dina(n11289), .dinb(n11287), .dout(n11703));
  jor  g11638(.dina(n11703), .dinb(n11702), .dout(n11704));
  jand g11639(.dina(n11704), .dinb(n11694), .dout(n11705));
  jand g11640(.dina(n11705), .dinb(n11693), .dout(n11706));
  jand g11641(.dina(n11703), .dinb(n11702), .dout(n11707));
  jor  g11642(.dina(n11707), .dinb(n11706), .dout(n11708));
  jor  g11643(.dina(n11708), .dinb(n11430), .dout(n11709));
  jnot g11644(.din(n5303), .dout(n11710));
  jor  g11645(.dina(n10847), .dinb(n11710), .dout(n11711));
  jor  g11646(.dina(n10845), .dinb(n2127), .dout(n11712));
  jor  g11647(.dina(n11360), .dinb(n2066), .dout(n11713));
  jor  g11648(.dina(n11458), .dinb(n1955), .dout(n11714));
  jand g11649(.dina(n11714), .dinb(n11713), .dout(n11715));
  jand g11650(.dina(n11715), .dinb(n11712), .dout(n11716));
  jand g11651(.dina(n11716), .dinb(n11711), .dout(n11717));
  jxor g11652(.dina(n11717), .dinb(\a[2] ), .dout(n11718));
  jand g11653(.dina(n11718), .dinb(n11709), .dout(n11719));
  jand g11654(.dina(n11708), .dinb(n11430), .dout(n11720));
  jor  g11655(.dina(n11720), .dinb(n11719), .dout(n11721));
  jor  g11656(.dina(n11721), .dinb(n11428), .dout(n11722));
  jnot g11657(.din(n5440), .dout(n11723));
  jor  g11658(.dina(n10847), .dinb(n11723), .dout(n11724));
  jor  g11659(.dina(n10845), .dinb(n2066), .dout(n11725));
  jor  g11660(.dina(n11360), .dinb(n1955), .dout(n11726));
  jor  g11661(.dina(n11458), .dinb(n1861), .dout(n11727));
  jand g11662(.dina(n11727), .dinb(n11726), .dout(n11728));
  jand g11663(.dina(n11728), .dinb(n11725), .dout(n11729));
  jand g11664(.dina(n11729), .dinb(n11724), .dout(n11730));
  jxor g11665(.dina(n11730), .dinb(\a[2] ), .dout(n11731));
  jand g11666(.dina(n11731), .dinb(n11722), .dout(n11732));
  jand g11667(.dina(n11721), .dinb(n11428), .dout(n11733));
  jor  g11668(.dina(n11733), .dinb(n11732), .dout(n11734));
  jor  g11669(.dina(n11734), .dinb(n11426), .dout(n11735));
  jand g11670(.dina(n11734), .dinb(n11426), .dout(n11736));
  jnot g11671(.din(n5092), .dout(n11737));
  jor  g11672(.dina(n10847), .dinb(n11737), .dout(n11738));
  jor  g11673(.dina(n11458), .dinb(n1775), .dout(n11739));
  jor  g11674(.dina(n11360), .dinb(n1861), .dout(n11740));
  jor  g11675(.dina(n10845), .dinb(n1955), .dout(n11741));
  jand g11676(.dina(n11741), .dinb(n11740), .dout(n11742));
  jand g11677(.dina(n11742), .dinb(n11739), .dout(n11743));
  jand g11678(.dina(n11743), .dinb(n11738), .dout(n11744));
  jxor g11679(.dina(n11744), .dinb(n6600), .dout(n11745));
  jnot g11680(.din(n11745), .dout(n11746));
  jor  g11681(.dina(n11746), .dinb(n11736), .dout(n11747));
  jand g11682(.dina(n11747), .dinb(n11735), .dout(n11748));
  jor  g11683(.dina(n11748), .dinb(n11424), .dout(n11749));
  jand g11684(.dina(n11748), .dinb(n11424), .dout(n11750));
  jnot g11685(.din(n5075), .dout(n11751));
  jor  g11686(.dina(n10847), .dinb(n11751), .dout(n11752));
  jor  g11687(.dina(n11458), .dinb(n1623), .dout(n11753));
  jor  g11688(.dina(n11360), .dinb(n1775), .dout(n11754));
  jor  g11689(.dina(n10845), .dinb(n1861), .dout(n11755));
  jand g11690(.dina(n11755), .dinb(n11754), .dout(n11756));
  jand g11691(.dina(n11756), .dinb(n11753), .dout(n11757));
  jand g11692(.dina(n11757), .dinb(n11752), .dout(n11758));
  jxor g11693(.dina(n11758), .dinb(n6600), .dout(n11759));
  jnot g11694(.din(n11759), .dout(n11760));
  jor  g11695(.dina(n11760), .dinb(n11750), .dout(n11761));
  jand g11696(.dina(n11761), .dinb(n11749), .dout(n11762));
  jand g11697(.dina(n11762), .dinb(n11422), .dout(n11763));
  jnot g11698(.din(n4849), .dout(n11764));
  jor  g11699(.dina(n10847), .dinb(n11764), .dout(n11765));
  jor  g11700(.dina(n11458), .dinb(n1559), .dout(n11766));
  jor  g11701(.dina(n11360), .dinb(n1623), .dout(n11767));
  jor  g11702(.dina(n10845), .dinb(n1775), .dout(n11768));
  jand g11703(.dina(n11768), .dinb(n11767), .dout(n11769));
  jand g11704(.dina(n11769), .dinb(n11766), .dout(n11770));
  jand g11705(.dina(n11770), .dinb(n11765), .dout(n11771));
  jxor g11706(.dina(n11771), .dinb(n6600), .dout(n11772));
  jnot g11707(.din(n11772), .dout(n11773));
  jor  g11708(.dina(n11773), .dinb(n11763), .dout(n11774));
  jor  g11709(.dina(n11762), .dinb(n11422), .dout(n11775));
  jand g11710(.dina(n10846), .dinb(n4866), .dout(n11776));
  jand g11711(.dina(n11359), .dinb(n1560), .dout(n11777));
  jand g11712(.dina(n10844), .dinb(n1624), .dout(n11778));
  jand g11713(.dina(n11372), .dinb(n1445), .dout(n11779));
  jor  g11714(.dina(n11779), .dinb(n11778), .dout(n11780));
  jor  g11715(.dina(n11780), .dinb(n11777), .dout(n11781));
  jor  g11716(.dina(n11781), .dinb(n11776), .dout(n11782));
  jxor g11717(.dina(n11782), .dinb(n6600), .dout(n11783));
  jxor g11718(.dina(n11311), .dinb(n11309), .dout(n11784));
  jor  g11719(.dina(n11784), .dinb(n11783), .dout(n11785));
  jand g11720(.dina(n11785), .dinb(n11775), .dout(n11786));
  jand g11721(.dina(n11786), .dinb(n11774), .dout(n11787));
  jand g11722(.dina(n11784), .dinb(n11783), .dout(n11788));
  jor  g11723(.dina(n11788), .dinb(n11787), .dout(n11789));
  jor  g11724(.dina(n11789), .dinb(n11420), .dout(n11790));
  jnot g11725(.din(n4258), .dout(n11791));
  jor  g11726(.dina(n10847), .dinb(n11791), .dout(n11792));
  jor  g11727(.dina(n11360), .dinb(n1444), .dout(n11793));
  jor  g11728(.dina(n10845), .dinb(n1559), .dout(n11794));
  jor  g11729(.dina(n11458), .dinb(n1342), .dout(n11795));
  jand g11730(.dina(n11795), .dinb(n11794), .dout(n11796));
  jand g11731(.dina(n11796), .dinb(n11793), .dout(n11797));
  jand g11732(.dina(n11797), .dinb(n11792), .dout(n11798));
  jxor g11733(.dina(n11798), .dinb(\a[2] ), .dout(n11799));
  jand g11734(.dina(n11799), .dinb(n11790), .dout(n11800));
  jand g11735(.dina(n11789), .dinb(n11420), .dout(n11801));
  jor  g11736(.dina(n11801), .dinb(n11800), .dout(n11802));
  jor  g11737(.dina(n11802), .dinb(n11418), .dout(n11803));
  jnot g11738(.din(n4772), .dout(n11804));
  jor  g11739(.dina(n10847), .dinb(n11804), .dout(n11805));
  jor  g11740(.dina(n11360), .dinb(n1342), .dout(n11806));
  jor  g11741(.dina(n10845), .dinb(n1444), .dout(n11807));
  jor  g11742(.dina(n11458), .dinb(n1212), .dout(n11808));
  jand g11743(.dina(n11808), .dinb(n11807), .dout(n11809));
  jand g11744(.dina(n11809), .dinb(n11806), .dout(n11810));
  jand g11745(.dina(n11810), .dinb(n11805), .dout(n11811));
  jxor g11746(.dina(n11811), .dinb(\a[2] ), .dout(n11812));
  jand g11747(.dina(n11812), .dinb(n11803), .dout(n11813));
  jand g11748(.dina(n11802), .dinb(n11418), .dout(n11814));
  jor  g11749(.dina(n11814), .dinb(n11813), .dout(n11815));
  jor  g11750(.dina(n11815), .dinb(n11416), .dout(n11816));
  jand g11751(.dina(n11815), .dinb(n11416), .dout(n11817));
  jnot g11752(.din(n4043), .dout(n11818));
  jor  g11753(.dina(n10847), .dinb(n11818), .dout(n11819));
  jor  g11754(.dina(n11458), .dinb(n1075), .dout(n11820));
  jor  g11755(.dina(n11360), .dinb(n1212), .dout(n11821));
  jor  g11756(.dina(n10845), .dinb(n1342), .dout(n11822));
  jand g11757(.dina(n11822), .dinb(n11821), .dout(n11823));
  jand g11758(.dina(n11823), .dinb(n11820), .dout(n11824));
  jand g11759(.dina(n11824), .dinb(n11819), .dout(n11825));
  jxor g11760(.dina(n11825), .dinb(n6600), .dout(n11826));
  jnot g11761(.din(n11826), .dout(n11827));
  jor  g11762(.dina(n11827), .dinb(n11817), .dout(n11828));
  jand g11763(.dina(n11828), .dinb(n11816), .dout(n11829));
  jand g11764(.dina(n11829), .dinb(n11414), .dout(n11830));
  jnot g11765(.din(n4026), .dout(n11831));
  jor  g11766(.dina(n10847), .dinb(n11831), .dout(n11832));
  jor  g11767(.dina(n11360), .dinb(n1075), .dout(n11833));
  jor  g11768(.dina(n11458), .dinb(n921), .dout(n11834));
  jor  g11769(.dina(n10845), .dinb(n1212), .dout(n11835));
  jand g11770(.dina(n11835), .dinb(n11834), .dout(n11836));
  jand g11771(.dina(n11836), .dinb(n11833), .dout(n11837));
  jand g11772(.dina(n11837), .dinb(n11832), .dout(n11838));
  jxor g11773(.dina(n11838), .dinb(n6600), .dout(n11839));
  jnot g11774(.din(n11839), .dout(n11840));
  jor  g11775(.dina(n11840), .dinb(n11830), .dout(n11841));
  jor  g11776(.dina(n11829), .dinb(n11414), .dout(n11842));
  jand g11777(.dina(n10846), .dinb(n3848), .dout(n11843));
  jand g11778(.dina(n10844), .dinb(n1076), .dout(n11844));
  jand g11779(.dina(n11359), .dinb(n922), .dout(n11845));
  jand g11780(.dina(n11372), .dinb(n3853), .dout(n11846));
  jor  g11781(.dina(n11846), .dinb(n11845), .dout(n11847));
  jor  g11782(.dina(n11847), .dinb(n11844), .dout(n11848));
  jor  g11783(.dina(n11848), .dinb(n11843), .dout(n11849));
  jxor g11784(.dina(n11849), .dinb(n6600), .dout(n11850));
  jxor g11785(.dina(n11327), .dinb(n11326), .dout(n11851));
  jor  g11786(.dina(n11851), .dinb(n11850), .dout(n11852));
  jand g11787(.dina(n11852), .dinb(n11842), .dout(n11853));
  jand g11788(.dina(n11853), .dinb(n11841), .dout(n11854));
  jand g11789(.dina(n11851), .dinb(n11850), .dout(n11855));
  jor  g11790(.dina(n11855), .dinb(n11854), .dout(n11856));
  jor  g11791(.dina(n11856), .dinb(n11412), .dout(n11857));
  jand g11792(.dina(n11857), .dinb(n11411), .dout(n11858));
  jxor g11793(.dina(n11399), .dinb(n11390), .dout(n11859));
  jor  g11794(.dina(n11859), .dinb(n11858), .dout(n11860));
  jand g11795(.dina(n11860), .dinb(n11400), .dout(n11861));
  jxor g11796(.dina(n11388), .dinb(n11379), .dout(n11862));
  jor  g11797(.dina(n11862), .dinb(n11861), .dout(n11863));
  jand g11798(.dina(n11863), .dinb(n11389), .dout(n11864));
  jxor g11799(.dina(n11377), .dinb(n11367), .dout(n11865));
  jnot g11800(.din(n11865), .dout(n11866));
  jor  g11801(.dina(n11866), .dinb(n11864), .dout(n11867));
  jand g11802(.dina(n11867), .dinb(n11378), .dout(n11868));
  jxor g11803(.dina(n11364), .dinb(n11356), .dout(n11869));
  jnot g11804(.din(n11869), .dout(n11870));
  jor  g11805(.dina(n11870), .dinb(n11868), .dout(n11871));
  jand g11806(.dina(n11871), .dinb(n11365), .dout(n11872));
  jor  g11807(.dina(n11872), .dinb(n11355), .dout(n11873));
  jand g11808(.dina(n11873), .dinb(n11353), .dout(n11874));
  jxor g11809(.dina(n10867), .dinb(n10866), .dout(n11875));
  jnot g11810(.din(n11875), .dout(n11876));
  jor  g11811(.dina(n11876), .dinb(n11874), .dout(n11877));
  jand g11812(.dina(n11877), .dinb(n10869), .dout(n11878));
  jxor g11813(.dina(n10837), .dinb(n10836), .dout(n11879));
  jnot g11814(.din(n11879), .dout(n11880));
  jor  g11815(.dina(n11880), .dinb(n11878), .dout(n11881));
  jand g11816(.dina(n11881), .dinb(n10839), .dout(n11882));
  jor  g11817(.dina(n11882), .dinb(n10367), .dout(n11883));
  jand g11818(.dina(n11883), .dinb(n10365), .dout(n11884));
  jnot g11819(.din(n11884), .dout(n11885));
  jxor g11820(.dina(n9931), .dinb(n9930), .dout(n11886));
  jand g11821(.dina(n11886), .dinb(n11885), .dout(n11887));
  jor  g11822(.dina(n11887), .dinb(n9932), .dout(n11888));
  jxor g11823(.dina(n9514), .dinb(n9513), .dout(n11889));
  jand g11824(.dina(n11889), .dinb(n11888), .dout(n11890));
  jor  g11825(.dina(n11890), .dinb(n9515), .dout(n11891));
  jand g11826(.dina(n11891), .dinb(n9141), .dout(n11892));
  jor  g11827(.dina(n11892), .dinb(n9140), .dout(n11893));
  jand g11828(.dina(n11893), .dinb(n8786), .dout(n11894));
  jor  g11829(.dina(n11894), .dinb(n8785), .dout(n11895));
  jxor g11830(.dina(n8464), .dinb(n8463), .dout(n11896));
  jand g11831(.dina(n11896), .dinb(n11895), .dout(n11897));
  jor  g11832(.dina(n11897), .dinb(n8465), .dout(n11898));
  jand g11833(.dina(n11898), .dinb(n8169), .dout(n11899));
  jor  g11834(.dina(n11899), .dinb(n8168), .dout(n11900));
  jxor g11835(.dina(n7903), .dinb(n7902), .dout(n11901));
  jand g11836(.dina(n11901), .dinb(n11900), .dout(n11902));
  jor  g11837(.dina(n11902), .dinb(n7904), .dout(n11903));
  jxor g11838(.dina(n7764), .dinb(n7763), .dout(n11904));
  jand g11839(.dina(n11904), .dinb(n11903), .dout(n11905));
  jor  g11840(.dina(n11905), .dinb(n7765), .dout(n11906));
  jand g11841(.dina(n11906), .dinb(n7628), .dout(n11907));
  jor  g11842(.dina(n11907), .dinb(n7627), .dout(n11908));
  jand g11843(.dina(n11908), .dinb(n6951), .dout(n11909));
  jor  g11844(.dina(n11909), .dinb(n6950), .dout(n11910));
  jand g11845(.dina(n11910), .dinb(n6823), .dout(n11911));
  jor  g11846(.dina(n11911), .dinb(n6822), .dout(n11912));
  jand g11847(.dina(n11912), .dinb(n6567), .dout(n11913));
  jor  g11848(.dina(n11913), .dinb(n6566), .dout(n11914));
  jxor g11849(.dina(n6353), .dinb(n6352), .dout(n11915));
  jand g11850(.dina(n11915), .dinb(n11914), .dout(n11916));
  jor  g11851(.dina(n11916), .dinb(n6354), .dout(n11917));
  jand g11852(.dina(n11917), .dinb(n6234), .dout(n11918));
  jor  g11853(.dina(n11918), .dinb(n6233), .dout(n11919));
  jand g11854(.dina(n11919), .dinb(n6142), .dout(n11920));
  jor  g11855(.dina(n11920), .dinb(n6141), .dout(n11921));
  jand g11856(.dina(n11921), .dinb(n5708), .dout(n11922));
  jor  g11857(.dina(n11922), .dinb(n5707), .dout(n11923));
  jxor g11858(.dina(n5523), .dinb(n5522), .dout(n11924));
  jand g11859(.dina(n11924), .dinb(n11923), .dout(n11925));
  jor  g11860(.dina(n11925), .dinb(n5524), .dout(n11926));
  jand g11861(.dina(n11926), .dinb(n5438), .dout(n11927));
  jor  g11862(.dina(n11927), .dinb(n5437), .dout(n11928));
  jxor g11863(.dina(n5377), .dinb(n4979), .dout(n11929));
  jand g11864(.dina(n11929), .dinb(n11928), .dout(n11930));
  jor  g11865(.dina(n11930), .dinb(n5378), .dout(n11931));
  jxor g11866(.dina(n4977), .dinb(n4976), .dout(n11932));
  jand g11867(.dina(n11932), .dinb(n11931), .dout(n11933));
  jor  g11868(.dina(n11933), .dinb(n4978), .dout(n11934));
  jxor g11869(.dina(n4928), .dinb(n4927), .dout(n11935));
  jand g11870(.dina(n11935), .dinb(n11934), .dout(n11936));
  jor  g11871(.dina(n11936), .dinb(n4929), .dout(n11937));
  jxor g11872(.dina(n4768), .dinb(n4767), .dout(n11938));
  jand g11873(.dina(n11938), .dinb(n11937), .dout(n11939));
  jor  g11874(.dina(n11939), .dinb(n4769), .dout(n11940));
  jxor g11875(.dina(n11940), .dinb(n4741), .dout(n11941));
  jxor g11876(.dina(n11938), .dinb(n11937), .dout(n11942));
  jand g11877(.dina(n11942), .dinb(n11941), .dout(n11943));
  jxor g11878(.dina(n11935), .dinb(n11934), .dout(n11944));
  jand g11879(.dina(n11944), .dinb(n11942), .dout(n11945));
  jxor g11880(.dina(n11932), .dinb(n11931), .dout(n11946));
  jand g11881(.dina(n11946), .dinb(n11944), .dout(n11947));
  jxor g11882(.dina(n11929), .dinb(n11928), .dout(n11948));
  jand g11883(.dina(n11948), .dinb(n11946), .dout(n11949));
  jxor g11884(.dina(n11926), .dinb(n5438), .dout(n11950));
  jand g11885(.dina(n11950), .dinb(n11948), .dout(n11951));
  jxor g11886(.dina(n11924), .dinb(n11923), .dout(n11952));
  jand g11887(.dina(n11952), .dinb(n11950), .dout(n11953));
  jxor g11888(.dina(n11921), .dinb(n5708), .dout(n11954));
  jand g11889(.dina(n11954), .dinb(n11952), .dout(n11955));
  jxor g11890(.dina(n11919), .dinb(n6142), .dout(n11956));
  jand g11891(.dina(n11956), .dinb(n11954), .dout(n11957));
  jxor g11892(.dina(n11917), .dinb(n6234), .dout(n11958));
  jand g11893(.dina(n11958), .dinb(n11956), .dout(n11959));
  jxor g11894(.dina(n11915), .dinb(n11914), .dout(n11960));
  jand g11895(.dina(n11960), .dinb(n11958), .dout(n11961));
  jxor g11896(.dina(n11912), .dinb(n6567), .dout(n11962));
  jand g11897(.dina(n11962), .dinb(n11960), .dout(n11963));
  jxor g11898(.dina(n11910), .dinb(n6823), .dout(n11964));
  jand g11899(.dina(n11964), .dinb(n11962), .dout(n11965));
  jxor g11900(.dina(n11908), .dinb(n6951), .dout(n11966));
  jand g11901(.dina(n11966), .dinb(n11964), .dout(n11967));
  jxor g11902(.dina(n11906), .dinb(n7628), .dout(n11968));
  jand g11903(.dina(n11968), .dinb(n11966), .dout(n11969));
  jxor g11904(.dina(n11904), .dinb(n11903), .dout(n11970));
  jand g11905(.dina(n11970), .dinb(n11968), .dout(n11971));
  jxor g11906(.dina(n11901), .dinb(n11900), .dout(n11972));
  jand g11907(.dina(n11972), .dinb(n11970), .dout(n11973));
  jxor g11908(.dina(n11898), .dinb(n8169), .dout(n11974));
  jand g11909(.dina(n11974), .dinb(n11972), .dout(n11975));
  jxor g11910(.dina(n11896), .dinb(n11895), .dout(n11976));
  jand g11911(.dina(n11976), .dinb(n11974), .dout(n11977));
  jxor g11912(.dina(n11893), .dinb(n8786), .dout(n11978));
  jand g11913(.dina(n11978), .dinb(n11976), .dout(n11979));
  jxor g11914(.dina(n11891), .dinb(n9141), .dout(n11980));
  jand g11915(.dina(n11980), .dinb(n11978), .dout(n11981));
  jxor g11916(.dina(n11889), .dinb(n11888), .dout(n11982));
  jand g11917(.dina(n11982), .dinb(n11980), .dout(n11983));
  jxor g11918(.dina(n11886), .dinb(n11884), .dout(n11984));
  jnot g11919(.din(n11984), .dout(n11985));
  jand g11920(.dina(n11985), .dinb(n11982), .dout(n11986));
  jxor g11921(.dina(n11882), .dinb(n10366), .dout(n11987));
  jnot g11922(.din(n11987), .dout(n11988));
  jand g11923(.dina(n11988), .dinb(n11985), .dout(n11989));
  jnot g11924(.din(n11989), .dout(n11990));
  jxor g11925(.dina(n11879), .dinb(n11878), .dout(n11991));
  jnot g11926(.din(n11991), .dout(n11992));
  jand g11927(.dina(n11992), .dinb(n11988), .dout(n11993));
  jnot g11928(.din(n11993), .dout(n11994));
  jxor g11929(.dina(n11875), .dinb(n11874), .dout(n11995));
  jor  g11930(.dina(n11995), .dinb(n11991), .dout(n11996));
  jxor g11931(.dina(n11872), .dinb(n11354), .dout(n11997));
  jor  g11932(.dina(n11997), .dinb(n11995), .dout(n11998));
  jxor g11933(.dina(n11869), .dinb(n11868), .dout(n11999));
  jor  g11934(.dina(n11999), .dinb(n11997), .dout(n12000));
  jxor g11935(.dina(n11865), .dinb(n11864), .dout(n12001));
  jor  g11936(.dina(n12001), .dinb(n11999), .dout(n12002));
  jnot g11937(.din(n11862), .dout(n12003));
  jxor g11938(.dina(n12003), .dinb(n11861), .dout(n12004));
  jor  g11939(.dina(n12004), .dinb(n12001), .dout(n12005));
  jxor g11940(.dina(n11862), .dinb(n11861), .dout(n12006));
  jxor g11941(.dina(n12006), .dinb(n12001), .dout(n12007));
  jxor g11942(.dina(n11859), .dinb(n11858), .dout(n12008));
  jnot g11943(.din(n12008), .dout(n12009));
  jxor g11944(.dina(n11856), .dinb(n11412), .dout(n12010));
  jnot g11945(.din(n12010), .dout(n12011));
  jand g11946(.dina(n12011), .dinb(n12004), .dout(n12012));
  jor  g11947(.dina(n12012), .dinb(n12009), .dout(n12013));
  jor  g11948(.dina(n12013), .dinb(n12007), .dout(n12014));
  jand g11949(.dina(n12014), .dinb(n12005), .dout(n12015));
  jxor g11950(.dina(n12001), .dinb(n11999), .dout(n12016));
  jnot g11951(.din(n12016), .dout(n12017));
  jor  g11952(.dina(n12017), .dinb(n12015), .dout(n12018));
  jand g11953(.dina(n12018), .dinb(n12002), .dout(n12019));
  jxor g11954(.dina(n11999), .dinb(n11997), .dout(n12020));
  jnot g11955(.din(n12020), .dout(n12021));
  jor  g11956(.dina(n12021), .dinb(n12019), .dout(n12022));
  jand g11957(.dina(n12022), .dinb(n12000), .dout(n12023));
  jxor g11958(.dina(n11997), .dinb(n11995), .dout(n12024));
  jnot g11959(.din(n12024), .dout(n12025));
  jor  g11960(.dina(n12025), .dinb(n12023), .dout(n12026));
  jand g11961(.dina(n12026), .dinb(n11998), .dout(n12027));
  jxor g11962(.dina(n11995), .dinb(n11991), .dout(n12028));
  jnot g11963(.din(n12028), .dout(n12029));
  jor  g11964(.dina(n12029), .dinb(n12027), .dout(n12030));
  jand g11965(.dina(n12030), .dinb(n11996), .dout(n12031));
  jxor g11966(.dina(n11991), .dinb(n11987), .dout(n12032));
  jnot g11967(.din(n12032), .dout(n12033));
  jor  g11968(.dina(n12033), .dinb(n12031), .dout(n12034));
  jand g11969(.dina(n12034), .dinb(n11994), .dout(n12035));
  jxor g11970(.dina(n11987), .dinb(n11984), .dout(n12036));
  jnot g11971(.din(n12036), .dout(n12037));
  jor  g11972(.dina(n12037), .dinb(n12035), .dout(n12038));
  jand g11973(.dina(n12038), .dinb(n11990), .dout(n12039));
  jnot g11974(.din(n12039), .dout(n12040));
  jxor g11975(.dina(n11985), .dinb(n11982), .dout(n12041));
  jand g11976(.dina(n12041), .dinb(n12040), .dout(n12042));
  jor  g11977(.dina(n12042), .dinb(n11986), .dout(n12043));
  jxor g11978(.dina(n11982), .dinb(n11980), .dout(n12044));
  jand g11979(.dina(n12044), .dinb(n12043), .dout(n12045));
  jor  g11980(.dina(n12045), .dinb(n11983), .dout(n12046));
  jxor g11981(.dina(n11980), .dinb(n11978), .dout(n12047));
  jand g11982(.dina(n12047), .dinb(n12046), .dout(n12048));
  jor  g11983(.dina(n12048), .dinb(n11981), .dout(n12049));
  jxor g11984(.dina(n11978), .dinb(n11976), .dout(n12050));
  jand g11985(.dina(n12050), .dinb(n12049), .dout(n12051));
  jor  g11986(.dina(n12051), .dinb(n11979), .dout(n12052));
  jxor g11987(.dina(n11976), .dinb(n11974), .dout(n12053));
  jand g11988(.dina(n12053), .dinb(n12052), .dout(n12054));
  jor  g11989(.dina(n12054), .dinb(n11977), .dout(n12055));
  jxor g11990(.dina(n11974), .dinb(n11972), .dout(n12056));
  jand g11991(.dina(n12056), .dinb(n12055), .dout(n12057));
  jor  g11992(.dina(n12057), .dinb(n11975), .dout(n12058));
  jxor g11993(.dina(n11972), .dinb(n11970), .dout(n12059));
  jand g11994(.dina(n12059), .dinb(n12058), .dout(n12060));
  jor  g11995(.dina(n12060), .dinb(n11973), .dout(n12061));
  jxor g11996(.dina(n11970), .dinb(n11968), .dout(n12062));
  jand g11997(.dina(n12062), .dinb(n12061), .dout(n12063));
  jor  g11998(.dina(n12063), .dinb(n11971), .dout(n12064));
  jxor g11999(.dina(n11968), .dinb(n11966), .dout(n12065));
  jand g12000(.dina(n12065), .dinb(n12064), .dout(n12066));
  jor  g12001(.dina(n12066), .dinb(n11969), .dout(n12067));
  jxor g12002(.dina(n11966), .dinb(n11964), .dout(n12068));
  jand g12003(.dina(n12068), .dinb(n12067), .dout(n12069));
  jor  g12004(.dina(n12069), .dinb(n11967), .dout(n12070));
  jxor g12005(.dina(n11964), .dinb(n11962), .dout(n12071));
  jand g12006(.dina(n12071), .dinb(n12070), .dout(n12072));
  jor  g12007(.dina(n12072), .dinb(n11965), .dout(n12073));
  jxor g12008(.dina(n11962), .dinb(n11960), .dout(n12074));
  jand g12009(.dina(n12074), .dinb(n12073), .dout(n12075));
  jor  g12010(.dina(n12075), .dinb(n11963), .dout(n12076));
  jxor g12011(.dina(n11960), .dinb(n11958), .dout(n12077));
  jand g12012(.dina(n12077), .dinb(n12076), .dout(n12078));
  jor  g12013(.dina(n12078), .dinb(n11961), .dout(n12079));
  jxor g12014(.dina(n11958), .dinb(n11956), .dout(n12080));
  jand g12015(.dina(n12080), .dinb(n12079), .dout(n12081));
  jor  g12016(.dina(n12081), .dinb(n11959), .dout(n12082));
  jxor g12017(.dina(n11956), .dinb(n11954), .dout(n12083));
  jand g12018(.dina(n12083), .dinb(n12082), .dout(n12084));
  jor  g12019(.dina(n12084), .dinb(n11957), .dout(n12085));
  jxor g12020(.dina(n11954), .dinb(n11952), .dout(n12086));
  jand g12021(.dina(n12086), .dinb(n12085), .dout(n12087));
  jor  g12022(.dina(n12087), .dinb(n11955), .dout(n12088));
  jxor g12023(.dina(n11952), .dinb(n11950), .dout(n12089));
  jand g12024(.dina(n12089), .dinb(n12088), .dout(n12090));
  jor  g12025(.dina(n12090), .dinb(n11953), .dout(n12091));
  jxor g12026(.dina(n11950), .dinb(n11948), .dout(n12092));
  jand g12027(.dina(n12092), .dinb(n12091), .dout(n12093));
  jor  g12028(.dina(n12093), .dinb(n11951), .dout(n12094));
  jxor g12029(.dina(n11948), .dinb(n11946), .dout(n12095));
  jand g12030(.dina(n12095), .dinb(n12094), .dout(n12096));
  jor  g12031(.dina(n12096), .dinb(n11949), .dout(n12097));
  jxor g12032(.dina(n11946), .dinb(n11944), .dout(n12098));
  jand g12033(.dina(n12098), .dinb(n12097), .dout(n12099));
  jor  g12034(.dina(n12099), .dinb(n11947), .dout(n12100));
  jxor g12035(.dina(n11944), .dinb(n11942), .dout(n12101));
  jand g12036(.dina(n12101), .dinb(n12100), .dout(n12102));
  jor  g12037(.dina(n12102), .dinb(n11945), .dout(n12103));
  jxor g12038(.dina(n11942), .dinb(n11941), .dout(n12104));
  jand g12039(.dina(n12104), .dinb(n12103), .dout(n12105));
  jor  g12040(.dina(n12105), .dinb(n11943), .dout(n12106));
  jand g12041(.dina(n4740), .dinb(n4648), .dout(n12107));
  jand g12042(.dina(n11940), .dinb(n4741), .dout(n12108));
  jor  g12043(.dina(n12108), .dinb(n12107), .dout(n12109));
  jand g12044(.dina(n4721), .dinb(n4653), .dout(n12110));
  jnot g12045(.din(n12110), .dout(n12111));
  jor  g12046(.dina(n4739), .dinb(n4723), .dout(n12112));
  jand g12047(.dina(n12112), .dinb(n12111), .dout(n12113));
  jnot g12048(.din(n12113), .dout(n12114));
  jnot g12049(.din(n4719), .dout(n12115));
  jand g12050(.dina(n2766), .dinb(n2301), .dout(n12116));
  jand g12051(.dina(n12116), .dinb(n3585), .dout(n12117));
  jand g12052(.dina(n3363), .dinb(n1281), .dout(n12118));
  jand g12053(.dina(n2130), .dinb(n880), .dout(n12119));
  jand g12054(.dina(n12119), .dinb(n12118), .dout(n12120));
  jand g12055(.dina(n12120), .dinb(n12117), .dout(n12121));
  jand g12056(.dina(n12121), .dinb(n2563), .dout(n12122));
  jand g12057(.dina(n4670), .dinb(n1984), .dout(n12123));
  jand g12058(.dina(n3989), .dinb(n1287), .dout(n12124));
  jand g12059(.dina(n12124), .dinb(n12123), .dout(n12125));
  jand g12060(.dina(n707), .dinb(n778), .dout(n12126));
  jand g12061(.dina(n12126), .dinb(n1178), .dout(n12127));
  jand g12062(.dina(n874), .dinb(n161), .dout(n12128));
  jand g12063(.dina(n667), .dinb(n245), .dout(n12129));
  jand g12064(.dina(n12129), .dinb(n12128), .dout(n12130));
  jand g12065(.dina(n12130), .dinb(n12127), .dout(n12131));
  jand g12066(.dina(n12131), .dinb(n12125), .dout(n12132));
  jand g12067(.dina(n913), .dinb(n197), .dout(n12133));
  jand g12068(.dina(n1346), .dinb(n1314), .dout(n12134));
  jand g12069(.dina(n12134), .dinb(n12133), .dout(n12135));
  jand g12070(.dina(n12135), .dinb(n3467), .dout(n12136));
  jand g12071(.dina(n5815), .dinb(n1988), .dout(n12137));
  jand g12072(.dina(n12137), .dinb(n12136), .dout(n12138));
  jand g12073(.dina(n12138), .dinb(n12132), .dout(n12139));
  jand g12074(.dina(n12139), .dinb(n1650), .dout(n12140));
  jand g12075(.dina(n12140), .dinb(n12122), .dout(n12141));
  jand g12076(.dina(n1205), .dinb(n869), .dout(n12142));
  jand g12077(.dina(n12142), .dinb(n3789), .dout(n12143));
  jand g12078(.dina(n997), .dinb(n751), .dout(n12144));
  jand g12079(.dina(n692), .dinb(n383), .dout(n12145));
  jand g12080(.dina(n12145), .dinb(n12144), .dout(n12146));
  jand g12081(.dina(n2304), .dinb(n2282), .dout(n12147));
  jand g12082(.dina(n12147), .dinb(n12146), .dout(n12148));
  jand g12083(.dina(n12148), .dinb(n932), .dout(n12149));
  jand g12084(.dina(n12149), .dinb(n12143), .dout(n12150));
  jand g12085(.dina(n1032), .dinb(n305), .dout(n12151));
  jand g12086(.dina(n12151), .dinb(n12150), .dout(n12152));
  jand g12087(.dina(n12152), .dinb(n2095), .dout(n12153));
  jand g12088(.dina(n12153), .dinb(n12141), .dout(n12154));
  jxor g12089(.dina(n12154), .dinb(n12115), .dout(n12155));
  jand g12090(.dina(n4719), .dinb(n4539), .dout(n12156));
  jand g12091(.dina(n12115), .dinb(n4540), .dout(n12157));
  jnot g12092(.din(n12157), .dout(n12158));
  jand g12093(.dina(n12158), .dinb(n4660), .dout(n12159));
  jor  g12094(.dina(n12159), .dinb(n12156), .dout(n12160));
  jxor g12095(.dina(n12160), .dinb(n12155), .dout(n12161));
  jor  g12096(.dina(n4728), .dinb(n4724), .dout(n12162));
  jand g12097(.dina(n12162), .dinb(n4733), .dout(n12163));
  jor  g12098(.dina(n12163), .dinb(n4630), .dout(n12164));
  jxor g12099(.dina(n12164), .dinb(\a[29] ), .dout(n12165));
  jnot g12100(.din(n12165), .dout(n12166));
  jand g12101(.dina(n4752), .dinb(n732), .dout(n12167));
  jand g12102(.dina(n4451), .dinb(n3858), .dout(n12168));
  jand g12103(.dina(n4358), .dinb(n3851), .dout(n12169));
  jand g12104(.dina(n4598), .dinb(n3855), .dout(n12170));
  jor  g12105(.dina(n12170), .dinb(n12169), .dout(n12171));
  jor  g12106(.dina(n12171), .dinb(n12168), .dout(n12172));
  jor  g12107(.dina(n12172), .dinb(n12167), .dout(n12173));
  jxor g12108(.dina(n12173), .dinb(n12166), .dout(n12174));
  jxor g12109(.dina(n12174), .dinb(n12161), .dout(n12175));
  jxor g12110(.dina(n12175), .dinb(n12114), .dout(n12176));
  jxor g12111(.dina(n12176), .dinb(n12109), .dout(n12177));
  jxor g12112(.dina(n12177), .dinb(n11941), .dout(n12178));
  jxor g12113(.dina(n12178), .dinb(n12106), .dout(n12179));
  jand g12114(.dina(n12179), .dinb(n75), .dout(n12180));
  jand g12115(.dina(n12177), .dinb(n4933), .dout(n12181));
  jand g12116(.dina(n11941), .dinb(n4918), .dout(n12182));
  jand g12117(.dina(n11942), .dinb(n4745), .dout(n12183));
  jor  g12118(.dina(n12183), .dinb(n12182), .dout(n12184));
  jor  g12119(.dina(n12184), .dinb(n12181), .dout(n12185));
  jor  g12120(.dina(n12185), .dinb(n12180), .dout(n12186));
  jxor g12121(.dina(n12186), .dinb(n68), .dout(n12187));
  jnot g12122(.din(n12187), .dout(n12188));
  jxor g12123(.dina(n12098), .dinb(n12097), .dout(n12189));
  jand g12124(.dina(n12189), .dinb(n4449), .dout(n12190));
  jand g12125(.dina(n11944), .dinb(n4453), .dout(n12191));
  jand g12126(.dina(n11946), .dinb(n4457), .dout(n12192));
  jand g12127(.dina(n11948), .dinb(n4461), .dout(n12193));
  jor  g12128(.dina(n12193), .dinb(n12192), .dout(n12194));
  jor  g12129(.dina(n12194), .dinb(n12191), .dout(n12195));
  jor  g12130(.dina(n12195), .dinb(n12190), .dout(n12196));
  jxor g12131(.dina(n12196), .dinb(n88), .dout(n12197));
  jnot g12132(.din(n12197), .dout(n12198));
  jand g12133(.dina(n907), .dinb(n346), .dout(n12199));
  jand g12134(.dina(n12199), .dinb(n4163), .dout(n12200));
  jand g12135(.dina(n12200), .dinb(n2301), .dout(n12201));
  jand g12136(.dina(n703), .dinb(n511), .dout(n12202));
  jand g12137(.dina(n434), .dinb(n292), .dout(n12203));
  jand g12138(.dina(n12203), .dinb(n12202), .dout(n12204));
  jand g12139(.dina(n635), .dinb(n194), .dout(n12205));
  jnot g12140(.din(n12205), .dout(n12206));
  jor  g12141(.dina(n12206), .dinb(n3383), .dout(n12207));
  jnot g12142(.din(n12207), .dout(n12208));
  jand g12143(.dina(n12208), .dinb(n12204), .dout(n12209));
  jand g12144(.dina(n12209), .dinb(n12201), .dout(n12210));
  jand g12145(.dina(n786), .dinb(n336), .dout(n12211));
  jand g12146(.dina(n687), .dinb(n778), .dout(n12212));
  jand g12147(.dina(n12212), .dinb(n12211), .dout(n12213));
  jand g12148(.dina(n12213), .dinb(n4301), .dout(n12214));
  jand g12149(.dina(n12214), .dinb(n6604), .dout(n12215));
  jand g12150(.dina(n12215), .dinb(n12210), .dout(n12216));
  jand g12151(.dina(n12216), .dinb(n5194), .dout(n12217));
  jnot g12152(.din(n3611), .dout(n12218));
  jand g12153(.dina(n12218), .dinb(n311), .dout(n12219));
  jand g12154(.dina(n12219), .dinb(n12217), .dout(n12220));
  jand g12155(.dina(n1454), .dinb(n1216), .dout(n12221));
  jand g12156(.dina(n1405), .dinb(n538), .dout(n12222));
  jand g12157(.dina(n12222), .dinb(n12221), .dout(n12223));
  jand g12158(.dina(n641), .dinb(n221), .dout(n12224));
  jand g12159(.dina(n12224), .dinb(n413), .dout(n12225));
  jand g12160(.dina(n3550), .dinb(n2135), .dout(n12226));
  jand g12161(.dina(n12226), .dinb(n12225), .dout(n12227));
  jand g12162(.dina(n12227), .dinb(n12223), .dout(n12228));
  jand g12163(.dina(n1409), .dinb(n228), .dout(n12229));
  jand g12164(.dina(n12229), .dinb(n177), .dout(n12230));
  jand g12165(.dina(n12230), .dinb(n2751), .dout(n12231));
  jand g12166(.dina(n3471), .dinb(n2483), .dout(n12232));
  jand g12167(.dina(n12232), .dinb(n2190), .dout(n12233));
  jand g12168(.dina(n12233), .dinb(n12231), .dout(n12234));
  jand g12169(.dina(n888), .dinb(n1597), .dout(n12235));
  jand g12170(.dina(n12235), .dinb(n1728), .dout(n12236));
  jand g12171(.dina(n1986), .dinb(n693), .dout(n12237));
  jand g12172(.dina(n12237), .dinb(n12236), .dout(n12238));
  jand g12173(.dina(n12238), .dinb(n380), .dout(n12239));
  jand g12174(.dina(n12239), .dinb(n12234), .dout(n12240));
  jand g12175(.dina(n12240), .dinb(n12228), .dout(n12241));
  jand g12176(.dina(n12241), .dinb(n3541), .dout(n12242));
  jand g12177(.dina(n12242), .dinb(n12220), .dout(n12243));
  jnot g12178(.din(n12243), .dout(n12244));
  jnot g12179(.din(n2089), .dout(n12245));
  jand g12180(.dina(n5807), .dinb(n12245), .dout(n12246));
  jand g12181(.dina(n607), .dinb(n286), .dout(n12247));
  jand g12182(.dina(n336), .dinb(n161), .dout(n12248));
  jand g12183(.dina(n12248), .dinb(n12247), .dout(n12249));
  jand g12184(.dina(n3496), .dinb(n1792), .dout(n12250));
  jand g12185(.dina(n4514), .dinb(n4076), .dout(n12251));
  jand g12186(.dina(n12251), .dinb(n12250), .dout(n12252));
  jand g12187(.dina(n12252), .dinb(n12249), .dout(n12253));
  jand g12188(.dina(n12253), .dinb(n5983), .dout(n12254));
  jand g12189(.dina(n3659), .dinb(n2029), .dout(n12255));
  jand g12190(.dina(n12255), .dinb(n12254), .dout(n12256));
  jand g12191(.dina(n12256), .dinb(n1173), .dout(n12257));
  jand g12192(.dina(n12257), .dinb(n12246), .dout(n12258));
  jand g12193(.dina(n542), .dinb(n441), .dout(n12259));
  jand g12194(.dina(n12259), .dinb(n2580), .dout(n12260));
  jand g12195(.dina(n719), .dinb(n249), .dout(n12261));
  jand g12196(.dina(n12261), .dinb(n2222), .dout(n12262));
  jand g12197(.dina(n12262), .dinb(n12260), .dout(n12263));
  jand g12198(.dina(n12263), .dinb(n1449), .dout(n12264));
  jand g12199(.dina(n842), .dinb(n337), .dout(n12265));
  jand g12200(.dina(n12265), .dinb(n2301), .dout(n12266));
  jand g12201(.dina(n217), .dinb(n134), .dout(n12267));
  jand g12202(.dina(n12267), .dinb(n1474), .dout(n12268));
  jand g12203(.dina(n12268), .dinb(n12266), .dout(n12269));
  jand g12204(.dina(n12269), .dinb(n4067), .dout(n12270));
  jand g12205(.dina(n12270), .dinb(n12264), .dout(n12271));
  jand g12206(.dina(n1991), .dinb(n178), .dout(n12272));
  jand g12207(.dina(n511), .dinb(n371), .dout(n12273));
  jand g12208(.dina(n12273), .dinb(n322), .dout(n12274));
  jand g12209(.dina(n12274), .dinb(n5168), .dout(n12275));
  jand g12210(.dina(n12275), .dinb(n12272), .dout(n12276));
  jand g12211(.dina(n12276), .dinb(n2615), .dout(n12277));
  jand g12212(.dina(n12277), .dinb(n12271), .dout(n12278));
  jand g12213(.dina(n12278), .dinb(n2658), .dout(n12279));
  jand g12214(.dina(n12279), .dinb(n7028), .dout(n12280));
  jor  g12215(.dina(n12280), .dinb(n12258), .dout(n12281));
  jand g12216(.dina(n4431), .dinb(n1167), .dout(n12282));
  jand g12217(.dina(n12282), .dinb(n1488), .dout(n12283));
  jand g12218(.dina(n12283), .dinb(n4580), .dout(n12284));
  jand g12219(.dina(n2583), .dinb(n607), .dout(n12285));
  jand g12220(.dina(n352), .dinb(n154), .dout(n12286));
  jand g12221(.dina(n12286), .dinb(n1584), .dout(n12287));
  jand g12222(.dina(n12287), .dinb(n12285), .dout(n12288));
  jand g12223(.dina(n12288), .dinb(n4350), .dout(n12289));
  jand g12224(.dina(n12289), .dinb(n4618), .dout(n12290));
  jand g12225(.dina(n12290), .dinb(n12284), .dout(n12291));
  jand g12226(.dina(n12291), .dinb(n4566), .dout(n12292));
  jnot g12227(.din(n12292), .dout(n12293));
  jand g12228(.dina(n3445), .dinb(n1268), .dout(n12294));
  jand g12229(.dina(n12294), .dinb(n4332), .dout(n12295));
  jand g12230(.dina(n4314), .dinb(n3032), .dout(n12296));
  jand g12231(.dina(n12296), .dinb(n12295), .dout(n12297));
  jand g12232(.dina(n12297), .dinb(n4563), .dout(n12298));
  jand g12233(.dina(n5919), .dinb(n4614), .dout(n12299));
  jand g12234(.dina(n12299), .dinb(n12298), .dout(n12300));
  jand g12235(.dina(n1615), .dinb(n180), .dout(n12301));
  jand g12236(.dina(n12301), .dinb(n2672), .dout(n12302));
  jand g12237(.dina(n12302), .dinb(n1078), .dout(n12303));
  jand g12238(.dina(n12303), .dinb(n4412), .dout(n12304));
  jand g12239(.dina(n12304), .dinb(n948), .dout(n12305));
  jand g12240(.dina(n12305), .dinb(n12300), .dout(n12306));
  jand g12241(.dina(n12306), .dinb(n4406), .dout(n12307));
  jand g12242(.dina(n12307), .dinb(n12293), .dout(n12308));
  jxor g12243(.dina(n12307), .dinb(n12293), .dout(n12309));
  jnot g12244(.din(n12308), .dout(n12315));
  jand g12245(.dina(n4314), .dinb(n946), .dout(n12316));
  jand g12246(.dina(n888), .dinb(n82), .dout(n12317));
  jand g12247(.dina(n12317), .dinb(n330), .dout(n12318));
  jand g12248(.dina(n12318), .dinb(n4431), .dout(n12319));
  jand g12249(.dina(n12319), .dinb(n12316), .dout(n12320));
  jand g12250(.dina(n12320), .dinb(n4579), .dout(n12321));
  jand g12251(.dina(n12321), .dinb(n4416), .dout(n12322));
  jxor g12252(.dina(n12322), .dinb(n12307), .dout(n12323));
  jnot g12253(.din(n12309), .dout(n12326));
  jnot g12254(.din(n12154), .dout(n12327));
  jand g12255(.dina(n7425), .dinb(n5790), .dout(n12328));
  jand g12256(.dina(n12328), .dinb(n4323), .dout(n12329));
  jand g12257(.dina(n2547), .dinb(n202), .dout(n12330));
  jand g12258(.dina(n888), .dinb(n276), .dout(n12331));
  jand g12259(.dina(n12331), .dinb(n2164), .dout(n12332));
  jand g12260(.dina(n2239), .dinb(n1142), .dout(n12333));
  jand g12261(.dina(n12333), .dinb(n12332), .dout(n12334));
  jand g12262(.dina(n12334), .dinb(n12330), .dout(n12335));
  jand g12263(.dina(n12335), .dinb(n12284), .dout(n12336));
  jand g12264(.dina(n12336), .dinb(n4398), .dout(n12337));
  jand g12265(.dina(n12304), .dinb(n4331), .dout(n12338));
  jand g12266(.dina(n12338), .dinb(n12337), .dout(n12339));
  jand g12267(.dina(n12339), .dinb(n12329), .dout(n12340));
  jnot g12268(.din(n12340), .dout(n12341));
  jand g12269(.dina(n12341), .dinb(n12327), .dout(n12342));
  jnot g12270(.din(n12342), .dout(n12343));
  jand g12271(.dina(n12340), .dinb(n12154), .dout(n12344));
  jnot g12272(.din(n12344), .dout(n12345));
  jand g12273(.dina(n12345), .dinb(n88), .dout(n12346));
  jand g12274(.dina(n12346), .dinb(n12343), .dout(n12347));
  jnot g12275(.din(n12347), .dout(n12348));
  jand g12276(.dina(n12348), .dinb(n12343), .dout(n12349));
  jnot g12277(.din(n12349), .dout(n12350));
  jand g12278(.dina(n12350), .dinb(n12307), .dout(n12351));
  jnot g12279(.din(n12351), .dout(n12352));
  jnot g12280(.din(n12307), .dout(n12353));
  jand g12281(.dina(n12349), .dinb(n12353), .dout(n12354));
  jor  g12282(.dina(n4731), .dinb(n6463), .dout(n12355));
  jand g12283(.dina(n4631), .dinb(n3858), .dout(n12357));
  jnot g12284(.din(n12357), .dout(n12359));
  jand g12285(.dina(n12359), .dinb(n12355), .dout(n12360));
  jor  g12286(.dina(n12360), .dinb(n12354), .dout(n12361));
  jand g12287(.dina(n12361), .dinb(n12352), .dout(n12362));
  jor  g12288(.dina(n12362), .dinb(n12326), .dout(n12363));
  jxor g12289(.dina(n12362), .dinb(n12326), .dout(n12364));
  jand g12290(.dina(n12154), .dinb(n12115), .dout(n12365));
  jand g12291(.dina(n12160), .dinb(n12155), .dout(n12366));
  jor  g12292(.dina(n12366), .dinb(n12365), .dout(n12367));
  jand g12293(.dina(n12348), .dinb(n88), .dout(n12368));
  jand g12294(.dina(n12349), .dinb(n12345), .dout(n12369));
  jor  g12295(.dina(n12369), .dinb(n12368), .dout(n12370));
  jand g12296(.dina(n12370), .dinb(n12367), .dout(n12371));
  jxor g12297(.dina(n12370), .dinb(n12367), .dout(n12372));
  jand g12298(.dina(n4636), .dinb(n732), .dout(n12373));
  jand g12299(.dina(n4451), .dinb(n3851), .dout(n12374));
  jand g12300(.dina(n4598), .dinb(n3858), .dout(n12375));
  jor  g12301(.dina(n12375), .dinb(n12374), .dout(n12378));
  jor  g12302(.dina(n12378), .dinb(n12373), .dout(n12379));
  jand g12303(.dina(n12379), .dinb(n12372), .dout(n12380));
  jor  g12304(.dina(n12380), .dinb(n12371), .dout(n12381));
  jxor g12305(.dina(n12349), .dinb(n12353), .dout(n12382));
  jxor g12306(.dina(n12382), .dinb(n12360), .dout(n12383));
  jnot g12307(.din(n12383), .dout(n12384));
  jand g12308(.dina(n12384), .dinb(n12381), .dout(n12385));
  jxor g12309(.dina(n12384), .dinb(n12381), .dout(n12386));
  jand g12310(.dina(n12173), .dinb(n12166), .dout(n12387));
  jand g12311(.dina(n12174), .dinb(n12161), .dout(n12388));
  jor  g12312(.dina(n12388), .dinb(n12387), .dout(n12389));
  jxor g12313(.dina(n12379), .dinb(n12372), .dout(n12390));
  jand g12314(.dina(n12390), .dinb(n12389), .dout(n12391));
  jand g12315(.dina(n12175), .dinb(n12114), .dout(n12392));
  jand g12316(.dina(n12176), .dinb(n12109), .dout(n12393));
  jor  g12317(.dina(n12393), .dinb(n12392), .dout(n12394));
  jxor g12318(.dina(n12390), .dinb(n12389), .dout(n12395));
  jand g12319(.dina(n12395), .dinb(n12394), .dout(n12396));
  jor  g12320(.dina(n12396), .dinb(n12391), .dout(n12397));
  jand g12321(.dina(n12397), .dinb(n12386), .dout(n12398));
  jor  g12322(.dina(n12398), .dinb(n12385), .dout(n12399));
  jand g12323(.dina(n12399), .dinb(n12364), .dout(n12400));
  jnot g12324(.din(n12400), .dout(n12401));
  jand g12325(.dina(n12401), .dinb(n12363), .dout(n12402));
  jnot g12326(.din(n12402), .dout(n12403));
  jxor g12327(.dina(n12323), .dinb(n12315), .dout(n12404));
  jand g12328(.dina(n12404), .dinb(n12403), .dout(n12405));
  jnot g12329(.din(n12405), .dout(n12406));
  jand g12330(.dina(n12406), .dinb(n12315), .dout(n12407));
  jnot g12331(.din(n12407), .dout(n12408));
  jand g12332(.dina(n12322), .dinb(n12307), .dout(n12409));
  jnot g12333(.din(n12409), .dout(n12410));
  jand g12334(.dina(n1264), .dinb(n959), .dout(n12411));
  jand g12335(.dina(n1184), .dinb(n505), .dout(n12412));
  jand g12336(.dina(n12412), .dinb(n12411), .dout(n12413));
  jand g12337(.dina(n3144), .dinb(n2150), .dout(n12414));
  jand g12338(.dina(n12414), .dinb(n12413), .dout(n12415));
  jand g12339(.dina(n184), .dinb(n177), .dout(n12416));
  jand g12340(.dina(n12416), .dinb(n197), .dout(n12417));
  jand g12341(.dina(n414), .dinb(n357), .dout(n12418));
  jand g12342(.dina(n12418), .dinb(n736), .dout(n12419));
  jand g12343(.dina(n12419), .dinb(n12417), .dout(n12420));
  jand g12344(.dina(n12420), .dinb(n12415), .dout(n12421));
  jand g12345(.dina(n965), .dinb(n449), .dout(n12422));
  jand g12346(.dina(n12422), .dinb(n417), .dout(n12423));
  jand g12347(.dina(n12423), .dinb(n1405), .dout(n12424));
  jand g12348(.dina(n2606), .dinb(n2514), .dout(n12425));
  jand g12349(.dina(n12425), .dinb(n425), .dout(n12426));
  jand g12350(.dina(n12426), .dinb(n12424), .dout(n12427));
  jand g12351(.dina(n12427), .dinb(n12421), .dout(n12428));
  jand g12352(.dina(n12428), .dinb(n3522), .dout(n12429));
  jand g12353(.dina(n12429), .dinb(n591), .dout(n12430));
  jand g12354(.dina(n12430), .dinb(n2376), .dout(n12431));
  jand g12355(.dina(n5026), .dinb(n1204), .dout(n12432));
  jand g12356(.dina(n12432), .dinb(n1780), .dout(n12433));
  jand g12357(.dina(n4161), .dinb(n276), .dout(n12434));
  jand g12358(.dina(n913), .dinb(n1031), .dout(n12435));
  jand g12359(.dina(n12435), .dinb(n1243), .dout(n12436));
  jand g12360(.dina(n12436), .dinb(n12434), .dout(n12437));
  jand g12361(.dina(n12437), .dinb(n5041), .dout(n12438));
  jand g12362(.dina(n12438), .dinb(n12433), .dout(n12439));
  jand g12363(.dina(n690), .dinb(n483), .dout(n12455));
  jand g12364(.dina(n12455), .dinb(n4587), .dout(n12456));
  jand g12365(.dina(n12456), .dinb(n24127), .dout(n12457));
  jnot g12366(.din(n12457), .dout(n12458));
  jand g12367(.dina(n12458), .dinb(n12410), .dout(n12459));
  jand g12368(.dina(n12459), .dinb(n12408), .dout(n12460));
  jnot g12369(.din(n12460), .dout(n12461));
  jnot g12370(.din(n6932), .dout(n12462));
  jor  g12371(.dina(n6933), .dinb(n12462), .dout(n12463));
  jand g12372(.dina(n12463), .dinb(n12461), .dout(n12464));
  jxor g12373(.dina(n12464), .dinb(n5292), .dout(n12465));
  jxor g12374(.dina(n12280), .dinb(n12258), .dout(n12466));
  jand g12375(.dina(n12466), .dinb(n12465), .dout(n12467));
  jnot g12376(.din(n12467), .dout(n12468));
  jand g12377(.dina(n12468), .dinb(n12281), .dout(n12469));
  jor  g12378(.dina(n12469), .dinb(n12244), .dout(n12470));
  jxor g12379(.dina(n12469), .dinb(n12244), .dout(n12471));
  jxor g12380(.dina(n12083), .dinb(n12082), .dout(n12472));
  jand g12381(.dina(n12472), .dinb(n732), .dout(n12473));
  jand g12382(.dina(n11954), .dinb(n3855), .dout(n12474));
  jand g12383(.dina(n11958), .dinb(n3851), .dout(n12475));
  jand g12384(.dina(n11956), .dinb(n3858), .dout(n12476));
  jor  g12385(.dina(n12476), .dinb(n12475), .dout(n12477));
  jor  g12386(.dina(n12477), .dinb(n12474), .dout(n12478));
  jor  g12387(.dina(n12478), .dinb(n12473), .dout(n12479));
  jand g12388(.dina(n12479), .dinb(n12471), .dout(n12480));
  jnot g12389(.din(n12480), .dout(n12481));
  jand g12390(.dina(n12481), .dinb(n12470), .dout(n12482));
  jnot g12391(.din(n12482), .dout(n12483));
  jand g12392(.dina(n1047), .dinb(n716), .dout(n12484));
  jand g12393(.dina(n658), .dinb(n622), .dout(n12485));
  jand g12394(.dina(n12485), .dinb(n12484), .dout(n12486));
  jand g12395(.dina(n3590), .dinb(n2262), .dout(n12487));
  jand g12396(.dina(n12487), .dinb(n12486), .dout(n12488));
  jand g12397(.dina(n1727), .dinb(n1088), .dout(n12489));
  jand g12398(.dina(n3445), .dinb(n2620), .dout(n12490));
  jand g12399(.dina(n12490), .dinb(n12489), .dout(n12491));
  jand g12400(.dina(n508), .dinb(n340), .dout(n12492));
  jand g12401(.dina(n12492), .dinb(n429), .dout(n12493));
  jand g12402(.dina(n843), .dinb(n626), .dout(n12494));
  jand g12403(.dina(n12494), .dinb(n1281), .dout(n12495));
  jand g12404(.dina(n12495), .dinb(n12493), .dout(n12496));
  jand g12405(.dina(n12496), .dinb(n12491), .dout(n12497));
  jand g12406(.dina(n12497), .dinb(n12488), .dout(n12498));
  jand g12407(.dina(n472), .dinb(n92), .dout(n12499));
  jand g12408(.dina(n824), .dinb(n304), .dout(n12500));
  jand g12409(.dina(n12500), .dinb(n12499), .dout(n12501));
  jand g12410(.dina(n12501), .dinb(n3289), .dout(n12502));
  jand g12411(.dina(n12502), .dinb(n2251), .dout(n12503));
  jand g12412(.dina(n12503), .dinb(n5996), .dout(n12504));
  jand g12413(.dina(n12504), .dinb(n12498), .dout(n12505));
  jand g12414(.dina(n12505), .dinb(n4139), .dout(n12506));
  jand g12415(.dina(n12506), .dinb(n3153), .dout(n12507));
  jxor g12416(.dina(n12507), .dinb(n12244), .dout(n12508));
  jxor g12417(.dina(n12508), .dinb(n12483), .dout(n12509));
  jxor g12418(.dina(n12086), .dinb(n12085), .dout(n12510));
  jand g12419(.dina(n12510), .dinb(n732), .dout(n12511));
  jand g12420(.dina(n11952), .dinb(n3855), .dout(n12512));
  jand g12421(.dina(n11954), .dinb(n3858), .dout(n12513));
  jand g12422(.dina(n11956), .dinb(n3851), .dout(n12514));
  jor  g12423(.dina(n12514), .dinb(n12513), .dout(n12515));
  jor  g12424(.dina(n12515), .dinb(n12512), .dout(n12516));
  jor  g12425(.dina(n12516), .dinb(n12511), .dout(n12517));
  jand g12426(.dina(n12517), .dinb(n12509), .dout(n12518));
  jxor g12427(.dina(n12095), .dinb(n12094), .dout(n12519));
  jand g12428(.dina(n12519), .dinb(n4449), .dout(n12520));
  jand g12429(.dina(n11946), .dinb(n4453), .dout(n12521));
  jand g12430(.dina(n11948), .dinb(n4457), .dout(n12522));
  jand g12431(.dina(n11950), .dinb(n4461), .dout(n12523));
  jor  g12432(.dina(n12523), .dinb(n12522), .dout(n12524));
  jor  g12433(.dina(n12524), .dinb(n12521), .dout(n12525));
  jor  g12434(.dina(n12525), .dinb(n12520), .dout(n12526));
  jxor g12435(.dina(n12526), .dinb(n88), .dout(n12527));
  jnot g12436(.din(n12527), .dout(n12528));
  jxor g12437(.dina(n12517), .dinb(n12509), .dout(n12529));
  jand g12438(.dina(n12529), .dinb(n12528), .dout(n12530));
  jor  g12439(.dina(n12530), .dinb(n12518), .dout(n12531));
  jand g12440(.dina(n12507), .dinb(n12244), .dout(n12532));
  jand g12441(.dina(n12508), .dinb(n12483), .dout(n12533));
  jor  g12442(.dina(n12533), .dinb(n12532), .dout(n12534));
  jnot g12443(.din(n6336), .dout(n12535));
  jor  g12444(.dina(n6337), .dinb(n12535), .dout(n12536));
  jand g12445(.dina(n12536), .dinb(n12461), .dout(n12537));
  jxor g12446(.dina(n12537), .dinb(n5064), .dout(n12538));
  jand g12447(.dina(n605), .dinb(n214), .dout(n12539));
  jand g12448(.dina(n1066), .dinb(n671), .dout(n12540));
  jand g12449(.dina(n12540), .dinb(n12539), .dout(n12541));
  jand g12450(.dina(n3608), .dinb(n473), .dout(n12542));
  jand g12451(.dina(n12542), .dinb(n12541), .dout(n12543));
  jand g12452(.dina(n3911), .dinb(n1410), .dout(n12544));
  jand g12453(.dina(n12544), .dinb(n5196), .dout(n12545));
  jand g12454(.dina(n12545), .dinb(n12543), .dout(n12546));
  jand g12455(.dina(n234), .dinb(n136), .dout(n12547));
  jand g12456(.dina(n12547), .dinb(n1024), .dout(n12548));
  jand g12457(.dina(n12548), .dinb(n3566), .dout(n12549));
  jand g12458(.dina(n12549), .dinb(n7152), .dout(n12550));
  jand g12459(.dina(n3250), .dinb(n2292), .dout(n12551));
  jand g12460(.dina(n2483), .dinb(n647), .dout(n12552));
  jand g12461(.dina(n12552), .dinb(n12551), .dout(n12553));
  jand g12462(.dina(n893), .dinb(n92), .dout(n12554));
  jand g12463(.dina(n865), .dinb(n290), .dout(n12555));
  jand g12464(.dina(n12555), .dinb(n12554), .dout(n12556));
  jand g12465(.dina(n515), .dinb(n377), .dout(n12557));
  jand g12466(.dina(n1144), .dinb(n509), .dout(n12558));
  jand g12467(.dina(n12558), .dinb(n12557), .dout(n12559));
  jand g12468(.dina(n12559), .dinb(n12556), .dout(n12560));
  jand g12469(.dina(n12560), .dinb(n12553), .dout(n12561));
  jand g12470(.dina(n12561), .dinb(n12550), .dout(n12562));
  jand g12471(.dina(n12562), .dinb(n12546), .dout(n12563));
  jand g12472(.dina(n12563), .dinb(n3429), .dout(n12564));
  jand g12473(.dina(n12152), .dinb(n5584), .dout(n12565));
  jand g12474(.dina(n12565), .dinb(n12564), .dout(n12566));
  jxor g12475(.dina(n12566), .dinb(n12507), .dout(n12567));
  jxor g12476(.dina(n12567), .dinb(n12538), .dout(n12568));
  jxor g12477(.dina(n12089), .dinb(n12088), .dout(n12569));
  jand g12478(.dina(n12569), .dinb(n732), .dout(n12570));
  jand g12479(.dina(n11950), .dinb(n3855), .dout(n12571));
  jand g12480(.dina(n11952), .dinb(n3858), .dout(n12572));
  jand g12481(.dina(n11954), .dinb(n3851), .dout(n12573));
  jor  g12482(.dina(n12573), .dinb(n12572), .dout(n12574));
  jor  g12483(.dina(n12574), .dinb(n12571), .dout(n12575));
  jor  g12484(.dina(n12575), .dinb(n12570), .dout(n12576));
  jxor g12485(.dina(n12576), .dinb(n12568), .dout(n12577));
  jxor g12486(.dina(n12577), .dinb(n12534), .dout(n12578));
  jxor g12487(.dina(n12578), .dinb(n12531), .dout(n12579));
  jxor g12488(.dina(n12579), .dinb(n12198), .dout(n12580));
  jand g12489(.dina(n12580), .dinb(n12188), .dout(n12581));
  jnot g12490(.din(n12258), .dout(n12582));
  jand g12491(.dina(n1175), .dinb(n333), .dout(n12583));
  jand g12492(.dina(n1964), .dinb(n1852), .dout(n12584));
  jand g12493(.dina(n12584), .dinb(n12583), .dout(n12585));
  jand g12494(.dina(n757), .dinb(n385), .dout(n12586));
  jand g12495(.dina(n12586), .dinb(n1907), .dout(n12587));
  jand g12496(.dina(n12587), .dinb(n4422), .dout(n12588));
  jand g12497(.dina(n4109), .dinb(n501), .dout(n12589));
  jand g12498(.dina(n12589), .dinb(n558), .dout(n12590));
  jand g12499(.dina(n1221), .dinb(n407), .dout(n12591));
  jand g12500(.dina(n12591), .dinb(n1847), .dout(n12592));
  jand g12501(.dina(n2580), .dinb(n1119), .dout(n12593));
  jand g12502(.dina(n12593), .dinb(n12592), .dout(n12594));
  jand g12503(.dina(n12594), .dinb(n12590), .dout(n12595));
  jand g12504(.dina(n12595), .dinb(n12588), .dout(n12596));
  jand g12505(.dina(n12596), .dinb(n12585), .dout(n12597));
  jand g12506(.dina(n5003), .dinb(n263), .dout(n12598));
  jand g12507(.dina(n377), .dinb(n305), .dout(n12599));
  jand g12508(.dina(n465), .dinb(n441), .dout(n12600));
  jand g12509(.dina(n12600), .dinb(n12599), .dout(n12601));
  jand g12510(.dina(n12601), .dinb(n1511), .dout(n12602));
  jand g12511(.dina(n12602), .dinb(n12598), .dout(n12603));
  jand g12512(.dina(n483), .dinb(n413), .dout(n12604));
  jand g12513(.dina(n12604), .dinb(n5741), .dout(n12605));
  jand g12514(.dina(n1475), .dinb(n771), .dout(n12606));
  jand g12515(.dina(n12606), .dinb(n12605), .dout(n12607));
  jand g12516(.dina(n12607), .dinb(n3157), .dout(n12608));
  jand g12517(.dina(n12608), .dinb(n12603), .dout(n12609));
  jand g12518(.dina(n2660), .dinb(n1889), .dout(n12610));
  jand g12519(.dina(n3236), .dinb(n547), .dout(n12611));
  jand g12520(.dina(n12611), .dinb(n12610), .dout(n12612));
  jand g12521(.dina(n708), .dinb(n197), .dout(n12613));
  jand g12522(.dina(n926), .dinb(n805), .dout(n12614));
  jand g12523(.dina(n12614), .dinb(n12613), .dout(n12615));
  jand g12524(.dina(n12615), .dinb(n4168), .dout(n12616));
  jand g12525(.dina(n12616), .dinb(n12612), .dout(n12617));
  jand g12526(.dina(n12617), .dinb(n3926), .dout(n12618));
  jand g12527(.dina(n12618), .dinb(n12609), .dout(n12619));
  jand g12528(.dina(n12619), .dinb(n2951), .dout(n12620));
  jand g12529(.dina(n12620), .dinb(n12597), .dout(n12621));
  jor  g12530(.dina(n12621), .dinb(n12582), .dout(n12622));
  jxor g12531(.dina(n12621), .dinb(n12582), .dout(n12623));
  jxor g12532(.dina(n12077), .dinb(n12076), .dout(n12624));
  jand g12533(.dina(n12624), .dinb(n732), .dout(n12625));
  jand g12534(.dina(n11958), .dinb(n3855), .dout(n12626));
  jand g12535(.dina(n11960), .dinb(n3858), .dout(n12627));
  jand g12536(.dina(n11962), .dinb(n3851), .dout(n12628));
  jor  g12537(.dina(n12628), .dinb(n12627), .dout(n12629));
  jor  g12538(.dina(n12629), .dinb(n12626), .dout(n12630));
  jor  g12539(.dina(n12630), .dinb(n12625), .dout(n12631));
  jand g12540(.dina(n12631), .dinb(n12623), .dout(n12632));
  jnot g12541(.din(n12632), .dout(n12633));
  jand g12542(.dina(n12633), .dinb(n12622), .dout(n12634));
  jnot g12543(.din(n12634), .dout(n12635));
  jxor g12544(.dina(n12466), .dinb(n12465), .dout(n12636));
  jand g12545(.dina(n12636), .dinb(n12635), .dout(n12637));
  jxor g12546(.dina(n12636), .dinb(n12635), .dout(n12638));
  jxor g12547(.dina(n12080), .dinb(n12079), .dout(n12639));
  jand g12548(.dina(n12639), .dinb(n732), .dout(n12640));
  jand g12549(.dina(n11956), .dinb(n3855), .dout(n12641));
  jand g12550(.dina(n11958), .dinb(n3858), .dout(n12642));
  jand g12551(.dina(n11960), .dinb(n3851), .dout(n12643));
  jor  g12552(.dina(n12643), .dinb(n12642), .dout(n12644));
  jor  g12553(.dina(n12644), .dinb(n12641), .dout(n12645));
  jor  g12554(.dina(n12645), .dinb(n12640), .dout(n12646));
  jand g12555(.dina(n12646), .dinb(n12638), .dout(n12647));
  jor  g12556(.dina(n12647), .dinb(n12637), .dout(n12648));
  jxor g12557(.dina(n12479), .dinb(n12471), .dout(n12649));
  jand g12558(.dina(n12649), .dinb(n12648), .dout(n12650));
  jnot g12559(.din(n12650), .dout(n12651));
  jxor g12560(.dina(n12649), .dinb(n12648), .dout(n12652));
  jnot g12561(.din(n12652), .dout(n12653));
  jxor g12562(.dina(n12092), .dinb(n12091), .dout(n12654));
  jand g12563(.dina(n12654), .dinb(n4449), .dout(n12655));
  jand g12564(.dina(n11948), .dinb(n4453), .dout(n12656));
  jand g12565(.dina(n11950), .dinb(n4457), .dout(n12657));
  jand g12566(.dina(n11952), .dinb(n4461), .dout(n12658));
  jor  g12567(.dina(n12658), .dinb(n12657), .dout(n12659));
  jor  g12568(.dina(n12659), .dinb(n12656), .dout(n12660));
  jor  g12569(.dina(n12660), .dinb(n12655), .dout(n12661));
  jxor g12570(.dina(n12661), .dinb(n88), .dout(n12662));
  jor  g12571(.dina(n12662), .dinb(n12653), .dout(n12663));
  jand g12572(.dina(n12663), .dinb(n12651), .dout(n12664));
  jnot g12573(.din(n12664), .dout(n12665));
  jxor g12574(.dina(n12529), .dinb(n12528), .dout(n12666));
  jand g12575(.dina(n12666), .dinb(n12665), .dout(n12667));
  jnot g12576(.din(n12667), .dout(n12668));
  jxor g12577(.dina(n12666), .dinb(n12665), .dout(n12669));
  jnot g12578(.din(n12669), .dout(n12670));
  jxor g12579(.dina(n12104), .dinb(n12103), .dout(n12671));
  jand g12580(.dina(n12671), .dinb(n75), .dout(n12672));
  jand g12581(.dina(n11941), .dinb(n4933), .dout(n12673));
  jand g12582(.dina(n11942), .dinb(n4918), .dout(n12674));
  jand g12583(.dina(n11944), .dinb(n4745), .dout(n12675));
  jor  g12584(.dina(n12675), .dinb(n12674), .dout(n12676));
  jor  g12585(.dina(n12676), .dinb(n12673), .dout(n12677));
  jor  g12586(.dina(n12677), .dinb(n12672), .dout(n12678));
  jxor g12587(.dina(n12678), .dinb(n68), .dout(n12679));
  jor  g12588(.dina(n12679), .dinb(n12670), .dout(n12680));
  jand g12589(.dina(n12680), .dinb(n12668), .dout(n12681));
  jnot g12590(.din(n12681), .dout(n12682));
  jxor g12591(.dina(n12580), .dinb(n12188), .dout(n12683));
  jand g12592(.dina(n12683), .dinb(n12682), .dout(n12684));
  jor  g12593(.dina(n12684), .dinb(n12581), .dout(n12685));
  jand g12594(.dina(n12578), .dinb(n12531), .dout(n12686));
  jand g12595(.dina(n12579), .dinb(n12198), .dout(n12687));
  jor  g12596(.dina(n12687), .dinb(n12686), .dout(n12688));
  jand g12597(.dina(n12576), .dinb(n12568), .dout(n12689));
  jand g12598(.dina(n12577), .dinb(n12534), .dout(n12690));
  jor  g12599(.dina(n12690), .dinb(n12689), .dout(n12691));
  jor  g12600(.dina(n12566), .dinb(n12507), .dout(n12692));
  jand g12601(.dina(n12567), .dinb(n12538), .dout(n12693));
  jnot g12602(.din(n12693), .dout(n12694));
  jand g12603(.dina(n12694), .dinb(n12692), .dout(n12695));
  jand g12604(.dina(n503), .dinb(n314), .dout(n12696));
  jand g12605(.dina(n12696), .dinb(n2812), .dout(n12697));
  jand g12606(.dina(n12697), .dinb(n2660), .dout(n12698));
  jand g12607(.dina(n1144), .dinb(n224), .dout(n12699));
  jand g12608(.dina(n12699), .dinb(n5033), .dout(n12700));
  jand g12609(.dina(n12700), .dinb(n6999), .dout(n12701));
  jand g12610(.dina(n12701), .dinb(n12698), .dout(n12702));
  jand g12611(.dina(n3068), .dinb(n377), .dout(n12703));
  jand g12612(.dina(n12703), .dinb(n548), .dout(n12704));
  jand g12613(.dina(n12704), .dinb(n3261), .dout(n12705));
  jand g12614(.dina(n1231), .dinb(n641), .dout(n12706));
  jand g12615(.dina(n12706), .dinb(n154), .dout(n12707));
  jand g12616(.dina(n12331), .dinb(n2872), .dout(n12708));
  jand g12617(.dina(n12708), .dinb(n12707), .dout(n12709));
  jand g12618(.dina(n12709), .dinb(n5740), .dout(n12710));
  jand g12619(.dina(n12710), .dinb(n12705), .dout(n12711));
  jand g12620(.dina(n12711), .dinb(n12702), .dout(n12712));
  jand g12621(.dina(n1314), .dinb(n626), .dout(n12713));
  jand g12622(.dina(n1184), .dinb(n817), .dout(n12714));
  jand g12623(.dina(n12714), .dinb(n12713), .dout(n12715));
  jand g12624(.dina(n5122), .dinb(n544), .dout(n12716));
  jand g12625(.dina(n12716), .dinb(n12715), .dout(n12717));
  jand g12626(.dina(n12717), .dinb(n5166), .dout(n12718));
  jand g12627(.dina(n1167), .dinb(n174), .dout(n12719));
  jand g12628(.dina(n238), .dinb(n157), .dout(n12720));
  jand g12629(.dina(n12720), .dinb(n12719), .dout(n12721));
  jand g12630(.dina(n950), .dinb(n418), .dout(n12722));
  jand g12631(.dina(n708), .dinb(n635), .dout(n12723));
  jand g12632(.dina(n12723), .dinb(n12722), .dout(n12724));
  jand g12633(.dina(n12724), .dinb(n12721), .dout(n12725));
  jand g12634(.dina(n2164), .dinb(n1280), .dout(n12726));
  jand g12635(.dina(n12726), .dinb(n271), .dout(n12727));
  jand g12636(.dina(n12727), .dinb(n12725), .dout(n12728));
  jand g12637(.dina(n12728), .dinb(n12718), .dout(n12729));
  jand g12638(.dina(n926), .dinb(n500), .dout(n12730));
  jand g12639(.dina(n12730), .dinb(n551), .dout(n12731));
  jand g12640(.dina(n1519), .dinb(n393), .dout(n12732));
  jand g12641(.dina(n12732), .dinb(n1385), .dout(n12733));
  jand g12642(.dina(n12733), .dinb(n12731), .dout(n12734));
  jand g12643(.dina(n12734), .dinb(n12546), .dout(n12735));
  jand g12644(.dina(n12735), .dinb(n12729), .dout(n12736));
  jand g12645(.dina(n12736), .dinb(n12712), .dout(n12737));
  jand g12646(.dina(n12737), .dinb(n3456), .dout(n12738));
  jnot g12647(.din(n12738), .dout(n12739));
  jxor g12648(.dina(n12739), .dinb(n12695), .dout(n12740));
  jand g12649(.dina(n12654), .dinb(n732), .dout(n12741));
  jand g12650(.dina(n11948), .dinb(n3855), .dout(n12742));
  jand g12651(.dina(n11952), .dinb(n3851), .dout(n12743));
  jand g12652(.dina(n11950), .dinb(n3858), .dout(n12744));
  jor  g12653(.dina(n12744), .dinb(n12743), .dout(n12745));
  jor  g12654(.dina(n12745), .dinb(n12742), .dout(n12746));
  jor  g12655(.dina(n12746), .dinb(n12741), .dout(n12747));
  jxor g12656(.dina(n12747), .dinb(n12740), .dout(n12748));
  jxor g12657(.dina(n12748), .dinb(n12691), .dout(n12749));
  jnot g12658(.din(n12749), .dout(n12750));
  jxor g12659(.dina(n12101), .dinb(n12100), .dout(n12751));
  jand g12660(.dina(n12751), .dinb(n4449), .dout(n12752));
  jand g12661(.dina(n11942), .dinb(n4453), .dout(n12753));
  jand g12662(.dina(n11944), .dinb(n4457), .dout(n12754));
  jand g12663(.dina(n11946), .dinb(n4461), .dout(n12755));
  jor  g12664(.dina(n12755), .dinb(n12754), .dout(n12756));
  jor  g12665(.dina(n12756), .dinb(n12753), .dout(n12757));
  jor  g12666(.dina(n12757), .dinb(n12752), .dout(n12758));
  jxor g12667(.dina(n12758), .dinb(n88), .dout(n12759));
  jxor g12668(.dina(n12759), .dinb(n12750), .dout(n12760));
  jxor g12669(.dina(n12760), .dinb(n12688), .dout(n12761));
  jnot g12670(.din(n12761), .dout(n12762));
  jand g12671(.dina(n12177), .dinb(n11941), .dout(n12763));
  jand g12672(.dina(n12178), .dinb(n12106), .dout(n12764));
  jor  g12673(.dina(n12764), .dinb(n12763), .dout(n12765));
  jxor g12674(.dina(n12395), .dinb(n12394), .dout(n12766));
  jxor g12675(.dina(n12766), .dinb(n12177), .dout(n12767));
  jxor g12676(.dina(n12767), .dinb(n12765), .dout(n12768));
  jand g12677(.dina(n12768), .dinb(n75), .dout(n12769));
  jand g12678(.dina(n12766), .dinb(n4933), .dout(n12770));
  jand g12679(.dina(n12177), .dinb(n4918), .dout(n12771));
  jand g12680(.dina(n11941), .dinb(n4745), .dout(n12772));
  jor  g12681(.dina(n12772), .dinb(n12771), .dout(n12773));
  jor  g12682(.dina(n12773), .dinb(n12770), .dout(n12774));
  jor  g12683(.dina(n12774), .dinb(n12769), .dout(n12775));
  jxor g12684(.dina(n12775), .dinb(n68), .dout(n12776));
  jxor g12685(.dina(n12776), .dinb(n12762), .dout(n12777));
  jand g12686(.dina(n12777), .dinb(n12685), .dout(n12778));
  jnot g12687(.din(n12778), .dout(n12779));
  jxor g12688(.dina(n12777), .dinb(n12685), .dout(n12780));
  jnot g12689(.din(n12780), .dout(n12781));
  jxor g12690(.dina(n12399), .dinb(n12364), .dout(n12782));
  jxor g12691(.dina(n12397), .dinb(n12386), .dout(n12783));
  jand g12692(.dina(n12783), .dinb(n12782), .dout(n12784));
  jand g12693(.dina(n12783), .dinb(n12766), .dout(n12785));
  jand g12694(.dina(n12766), .dinb(n12177), .dout(n12786));
  jand g12695(.dina(n12767), .dinb(n12765), .dout(n12787));
  jor  g12696(.dina(n12787), .dinb(n12786), .dout(n12788));
  jxor g12697(.dina(n12783), .dinb(n12766), .dout(n12789));
  jand g12698(.dina(n12789), .dinb(n12788), .dout(n12790));
  jor  g12699(.dina(n12790), .dinb(n12785), .dout(n12791));
  jxor g12700(.dina(n12783), .dinb(n12782), .dout(n12792));
  jand g12701(.dina(n12792), .dinb(n12791), .dout(n12793));
  jor  g12702(.dina(n12793), .dinb(n12784), .dout(n12794));
  jxor g12703(.dina(n12404), .dinb(n12403), .dout(n12795));
  jxor g12704(.dina(n12795), .dinb(n12782), .dout(n12796));
  jxor g12705(.dina(n12796), .dinb(n12794), .dout(n12797));
  jand g12706(.dina(n12797), .dinb(n5365), .dout(n12798));
  jand g12707(.dina(n12795), .dinb(n5500), .dout(n12799));
  jand g12708(.dina(n12782), .dinb(n5424), .dout(n12800));
  jand g12709(.dina(n12783), .dinb(n5363), .dout(n12801));
  jor  g12710(.dina(n12801), .dinb(n12800), .dout(n12802));
  jor  g12711(.dina(n12802), .dinb(n12799), .dout(n12803));
  jor  g12712(.dina(n12803), .dinb(n12798), .dout(n12804));
  jxor g12713(.dina(n12804), .dinb(n72), .dout(n12805));
  jor  g12714(.dina(n12805), .dinb(n12781), .dout(n12806));
  jand g12715(.dina(n12806), .dinb(n12779), .dout(n12807));
  jand g12716(.dina(n12457), .dinb(n12409), .dout(n12808));
  jand g12717(.dina(n12808), .dinb(n12407), .dout(n12809));
  jnot g12718(.din(n12809), .dout(n12810));
  jand g12719(.dina(n12810), .dinb(n12461), .dout(n12811));
  jxor g12720(.dina(n12457), .dinb(n12409), .dout(n12813));
  jxor g12721(.dina(n12813), .dinb(n12408), .dout(n12814));
  jnot g12722(.din(n12814), .dout(n12815));
  jand g12723(.dina(n12815), .dinb(n12795), .dout(n12816));
  jand g12724(.dina(n12795), .dinb(n12782), .dout(n12817));
  jand g12725(.dina(n12796), .dinb(n12794), .dout(n12818));
  jor  g12726(.dina(n12818), .dinb(n12817), .dout(n12819));
  jnot g12727(.din(n12795), .dout(n12820));
  jxor g12728(.dina(n12814), .dinb(n12820), .dout(n12821));
  jand g12729(.dina(n12821), .dinb(n12819), .dout(n12822));
  jor  g12730(.dina(n12822), .dinb(n12816), .dout(n12823));
  jand g12731(.dina(n12823), .dinb(n12809), .dout(n12824));
  jnot g12732(.din(n12824), .dout(n12825));
  jand g12733(.dina(n6208), .dinb(n6132), .dout(n12829));
  jor  g12734(.dina(n12961), .dinb(n12807), .dout(n12834));
  jxor g12735(.dina(n12961), .dinb(n12807), .dout(n12835));
  jand g12736(.dina(n12760), .dinb(n12688), .dout(n12836));
  jnot g12737(.din(n12836), .dout(n12837));
  jor  g12738(.dina(n12776), .dinb(n12762), .dout(n12838));
  jand g12739(.dina(n12838), .dinb(n12837), .dout(n12839));
  jnot g12740(.din(n12839), .dout(n12840));
  jxor g12741(.dina(n12789), .dinb(n12788), .dout(n12841));
  jand g12742(.dina(n12841), .dinb(n75), .dout(n12842));
  jand g12743(.dina(n12783), .dinb(n4933), .dout(n12843));
  jand g12744(.dina(n12766), .dinb(n4918), .dout(n12844));
  jand g12745(.dina(n12177), .dinb(n4745), .dout(n12845));
  jor  g12746(.dina(n12845), .dinb(n12844), .dout(n12846));
  jor  g12747(.dina(n12846), .dinb(n12843), .dout(n12847));
  jor  g12748(.dina(n12847), .dinb(n12842), .dout(n12848));
  jxor g12749(.dina(n12848), .dinb(n68), .dout(n12849));
  jnot g12750(.din(n12849), .dout(n12850));
  jnot g12751(.din(n12695), .dout(n12851));
  jand g12752(.dina(n12738), .dinb(n12851), .dout(n12852));
  jand g12753(.dina(n12747), .dinb(n12740), .dout(n12853));
  jor  g12754(.dina(n12853), .dinb(n12852), .dout(n12854));
  jand g12755(.dina(n1519), .dinb(n500), .dout(n12855));
  jand g12756(.dina(n12855), .dinb(n874), .dout(n12856));
  jand g12757(.dina(n314), .dinb(n190), .dout(n12857));
  jand g12758(.dina(n12857), .dinb(n253), .dout(n12858));
  jand g12759(.dina(n12858), .dinb(n12856), .dout(n12859));
  jand g12760(.dina(n12859), .dinb(n5208), .dout(n12860));
  jand g12761(.dina(n331), .dinb(n165), .dout(n12861));
  jand g12762(.dina(n12861), .dinb(n586), .dout(n12862));
  jand g12763(.dina(n12862), .dinb(n2152), .dout(n12863));
  jand g12764(.dina(n292), .dinb(n134), .dout(n12864));
  jand g12765(.dina(n12864), .dinb(n3462), .dout(n12865));
  jand g12766(.dina(n4691), .dinb(n4382), .dout(n12866));
  jand g12767(.dina(n12866), .dinb(n12865), .dout(n12867));
  jand g12768(.dina(n12867), .dinb(n12863), .dout(n12868));
  jand g12769(.dina(n4184), .dinb(n2110), .dout(n12869));
  jand g12770(.dina(n12869), .dinb(n12868), .dout(n12870));
  jand g12771(.dina(n12870), .dinb(n12860), .dout(n12871));
  jand g12772(.dina(n12871), .dinb(n2775), .dout(n12872));
  jand g12773(.dina(n1205), .dinb(n883), .dout(n12873));
  jand g12774(.dina(n2606), .dinb(n1196), .dout(n12874));
  jand g12775(.dina(n12874), .dinb(n12873), .dout(n12875));
  jand g12776(.dina(n553), .dinb(n542), .dout(n12876));
  jand g12777(.dina(n1066), .dinb(n197), .dout(n12877));
  jand g12778(.dina(n12877), .dinb(n12876), .dout(n12878));
  jand g12779(.dina(n1986), .dinb(n1760), .dout(n12879));
  jand g12780(.dina(n12879), .dinb(n12878), .dout(n12880));
  jand g12781(.dina(n595), .dinb(n757), .dout(n12881));
  jand g12782(.dina(n404), .dinb(n382), .dout(n12882));
  jand g12783(.dina(n12882), .dinb(n12881), .dout(n12883));
  jand g12784(.dina(n12883), .dinb(n5147), .dout(n12884));
  jand g12785(.dina(n12884), .dinb(n12880), .dout(n12885));
  jand g12786(.dina(n12885), .dinb(n12875), .dout(n12886));
  jand g12787(.dina(n12886), .dinb(n2783), .dout(n12887));
  jand g12788(.dina(n12887), .dinb(n5954), .dout(n12888));
  jand g12789(.dina(n12888), .dinb(n12872), .dout(n12889));
  jxor g12790(.dina(n12889), .dinb(n12739), .dout(n12890));
  jand g12791(.dina(n12519), .dinb(n732), .dout(n12891));
  jand g12792(.dina(n11946), .dinb(n3855), .dout(n12892));
  jand g12793(.dina(n11948), .dinb(n3858), .dout(n12893));
  jand g12794(.dina(n11950), .dinb(n3851), .dout(n12894));
  jor  g12795(.dina(n12894), .dinb(n12893), .dout(n12895));
  jor  g12796(.dina(n12895), .dinb(n12892), .dout(n12896));
  jor  g12797(.dina(n12896), .dinb(n12891), .dout(n12897));
  jxor g12798(.dina(n12897), .dinb(n12890), .dout(n12898));
  jxor g12799(.dina(n12898), .dinb(n12854), .dout(n12899));
  jnot g12800(.din(n12899), .dout(n12900));
  jand g12801(.dina(n12748), .dinb(n12691), .dout(n12901));
  jnot g12802(.din(n12901), .dout(n12902));
  jor  g12803(.dina(n12759), .dinb(n12750), .dout(n12903));
  jand g12804(.dina(n12903), .dinb(n12902), .dout(n12904));
  jxor g12805(.dina(n12904), .dinb(n12900), .dout(n12905));
  jnot g12806(.din(n12905), .dout(n12906));
  jand g12807(.dina(n12671), .dinb(n4449), .dout(n12907));
  jand g12808(.dina(n11941), .dinb(n4453), .dout(n12908));
  jand g12809(.dina(n11942), .dinb(n4457), .dout(n12909));
  jand g12810(.dina(n11944), .dinb(n4461), .dout(n12910));
  jor  g12811(.dina(n12910), .dinb(n12909), .dout(n12911));
  jor  g12812(.dina(n12911), .dinb(n12908), .dout(n12912));
  jor  g12813(.dina(n12912), .dinb(n12907), .dout(n12913));
  jxor g12814(.dina(n12913), .dinb(n88), .dout(n12914));
  jxor g12815(.dina(n12914), .dinb(n12906), .dout(n12915));
  jxor g12816(.dina(n12915), .dinb(n12850), .dout(n12916));
  jxor g12817(.dina(n12916), .dinb(n12840), .dout(n12917));
  jnot g12818(.din(n12917), .dout(n12918));
  jxor g12819(.dina(n12821), .dinb(n12819), .dout(n12919));
  jand g12820(.dina(n12919), .dinb(n5365), .dout(n12920));
  jand g12821(.dina(n12815), .dinb(n5500), .dout(n12921));
  jand g12822(.dina(n12795), .dinb(n5424), .dout(n12922));
  jand g12823(.dina(n12782), .dinb(n5363), .dout(n12923));
  jor  g12824(.dina(n12923), .dinb(n12922), .dout(n12924));
  jor  g12825(.dina(n12924), .dinb(n12921), .dout(n12925));
  jor  g12826(.dina(n12925), .dinb(n12920), .dout(n12926));
  jxor g12827(.dina(n12926), .dinb(n72), .dout(n12927));
  jxor g12828(.dina(n12927), .dinb(n12918), .dout(n12928));
  jand g12829(.dina(n12928), .dinb(n12835), .dout(n12929));
  jnot g12830(.din(n12929), .dout(n12930));
  jand g12831(.dina(n12930), .dinb(n12834), .dout(n12931));
  jnot g12832(.din(n12931), .dout(n12932));
  jor  g12833(.dina(n12914), .dinb(n12906), .dout(n12933));
  jand g12834(.dina(n12915), .dinb(n12850), .dout(n12934));
  jnot g12835(.din(n12934), .dout(n12935));
  jand g12836(.dina(n12935), .dinb(n12933), .dout(n12936));
  jnot g12837(.din(n12936), .dout(n12937));
  jxor g12838(.dina(n12792), .dinb(n12791), .dout(n12938));
  jand g12839(.dina(n12938), .dinb(n75), .dout(n12939));
  jand g12840(.dina(n12782), .dinb(n4933), .dout(n12940));
  jand g12841(.dina(n12783), .dinb(n4918), .dout(n12941));
  jand g12842(.dina(n12766), .dinb(n4745), .dout(n12942));
  jor  g12843(.dina(n12942), .dinb(n12941), .dout(n12943));
  jor  g12844(.dina(n12943), .dinb(n12940), .dout(n12944));
  jor  g12845(.dina(n12944), .dinb(n12939), .dout(n12945));
  jxor g12846(.dina(n12945), .dinb(n68), .dout(n12946));
  jnot g12847(.din(n12946), .dout(n12947));
  jand g12848(.dina(n12898), .dinb(n12854), .dout(n12948));
  jnot g12849(.din(n12948), .dout(n12949));
  jor  g12850(.dina(n12904), .dinb(n12900), .dout(n12950));
  jand g12851(.dina(n12950), .dinb(n12949), .dout(n12951));
  jnot g12852(.din(n12951), .dout(n12952));
  jor  g12853(.dina(n12889), .dinb(n12739), .dout(n12953));
  jand g12854(.dina(n12897), .dinb(n12890), .dout(n12954));
  jnot g12855(.din(n12954), .dout(n12955));
  jand g12856(.dina(n12955), .dinb(n12953), .dout(n12956));
  jnot g12857(.din(n12956), .dout(n12957));
  jnot g12858(.din(n5689), .dout(n12958));
  jor  g12859(.dina(n5690), .dinb(n12958), .dout(n12959));
  jxor g12860(.dina(n12959), .dinb(n4247), .dout(n12961));
  jand g12861(.dina(n712), .dinb(n574), .dout(n12962));
  jand g12862(.dina(n12962), .dinb(n511), .dout(n12963));
  jand g12863(.dina(n1409), .dinb(n262), .dout(n12964));
  jand g12864(.dina(n12964), .dinb(n1435), .dout(n12965));
  jand g12865(.dina(n12965), .dinb(n12963), .dout(n12966));
  jand g12866(.dina(n2130), .dinb(n1412), .dout(n12967));
  jand g12867(.dina(n12967), .dinb(n845), .dout(n12968));
  jand g12868(.dina(n12968), .dinb(n12966), .dout(n12969));
  jand g12869(.dina(n5768), .dinb(n2840), .dout(n12970));
  jand g12870(.dina(n2697), .dinb(n858), .dout(n12971));
  jand g12871(.dina(n12971), .dinb(n12970), .dout(n12972));
  jand g12872(.dina(n12972), .dinb(n3416), .dout(n12973));
  jand g12873(.dina(n12973), .dinb(n12969), .dout(n12974));
  jand g12874(.dina(n12974), .dinb(n2215), .dout(n12975));
  jand g12875(.dina(n4667), .dinb(n1475), .dout(n12976));
  jand g12876(.dina(n12976), .dinb(n2239), .dout(n12977));
  jand g12877(.dina(n715), .dinb(n578), .dout(n12978));
  jand g12878(.dina(n700), .dinb(n622), .dout(n12979));
  jand g12879(.dina(n12979), .dinb(n12978), .dout(n12980));
  jand g12880(.dina(n1846), .dinb(n1600), .dout(n12981));
  jand g12881(.dina(n12981), .dinb(n12980), .dout(n12982));
  jand g12882(.dina(n3057), .dinb(n431), .dout(n12983));
  jand g12883(.dina(n12983), .dinb(n4190), .dout(n12984));
  jand g12884(.dina(n12984), .dinb(n12982), .dout(n12985));
  jand g12885(.dina(n12985), .dinb(n12977), .dout(n12986));
  jand g12886(.dina(n3582), .dinb(n1871), .dout(n12987));
  jand g12887(.dina(n12987), .dinb(n12986), .dout(n12988));
  jand g12888(.dina(n12988), .dinb(n12975), .dout(n12989));
  jand g12889(.dina(n12989), .dinb(n2532), .dout(n12990));
  jxor g12890(.dina(n12990), .dinb(n12738), .dout(n12991));
  jxor g12891(.dina(n12991), .dinb(n12961), .dout(n12992));
  jxor g12892(.dina(n12992), .dinb(n12957), .dout(n12993));
  jand g12893(.dina(n12189), .dinb(n732), .dout(n12994));
  jand g12894(.dina(n11944), .dinb(n3855), .dout(n12995));
  jand g12895(.dina(n11946), .dinb(n3858), .dout(n12996));
  jand g12896(.dina(n11948), .dinb(n3851), .dout(n12997));
  jor  g12897(.dina(n12997), .dinb(n12996), .dout(n12998));
  jor  g12898(.dina(n12998), .dinb(n12995), .dout(n12999));
  jor  g12899(.dina(n12999), .dinb(n12994), .dout(n13000));
  jxor g12900(.dina(n13000), .dinb(n12993), .dout(n13001));
  jxor g12901(.dina(n13001), .dinb(n12952), .dout(n13002));
  jnot g12902(.din(n13002), .dout(n13003));
  jand g12903(.dina(n12179), .dinb(n4449), .dout(n13004));
  jand g12904(.dina(n12177), .dinb(n4453), .dout(n13005));
  jand g12905(.dina(n11941), .dinb(n4457), .dout(n13006));
  jand g12906(.dina(n11942), .dinb(n4461), .dout(n13007));
  jor  g12907(.dina(n13007), .dinb(n13006), .dout(n13008));
  jor  g12908(.dina(n13008), .dinb(n13005), .dout(n13009));
  jor  g12909(.dina(n13009), .dinb(n13004), .dout(n13010));
  jxor g12910(.dina(n13010), .dinb(n88), .dout(n13011));
  jxor g12911(.dina(n13011), .dinb(n13003), .dout(n13012));
  jxor g12912(.dina(n13012), .dinb(n12947), .dout(n13013));
  jxor g12913(.dina(n13013), .dinb(n12937), .dout(n13014));
  jand g12914(.dina(n12916), .dinb(n12840), .dout(n13015));
  jnot g12915(.din(n13015), .dout(n13016));
  jor  g12916(.dina(n12927), .dinb(n12918), .dout(n13017));
  jand g12917(.dina(n13017), .dinb(n13016), .dout(n13018));
  jand g12918(.dina(n12407), .dinb(n12813), .dout(n13021));
  jxor g12919(.dina(n13021), .dinb(n12823), .dout(n13022));
  jand g12920(.dina(n13022), .dinb(n5365), .dout(n13023));
  jand g12921(.dina(n12815), .dinb(n5424), .dout(n13025));
  jand g12922(.dina(n12795), .dinb(n5363), .dout(n13026));
  jor  g12923(.dina(n13026), .dinb(n13025), .dout(n13027));
  jor  g12924(.dina(n13027), .dinb(n5500), .dout(n13028));
  jor  g12925(.dina(n13028), .dinb(n13023), .dout(n13029));
  jxor g12926(.dina(n13029), .dinb(n72), .dout(n13030));
  jxor g12927(.dina(n13030), .dinb(n13018), .dout(n13031));
  jxor g12928(.dina(n13031), .dinb(n13014), .dout(n13032));
  jand g12929(.dina(n13032), .dinb(n12932), .dout(n13033));
  jxor g12930(.dina(n12683), .dinb(n12682), .dout(n13034));
  jnot g12931(.din(n13034), .dout(n13035));
  jand g12932(.dina(n12938), .dinb(n5365), .dout(n13036));
  jand g12933(.dina(n12782), .dinb(n5500), .dout(n13037));
  jand g12934(.dina(n12783), .dinb(n5424), .dout(n13038));
  jand g12935(.dina(n12766), .dinb(n5363), .dout(n13039));
  jor  g12936(.dina(n13039), .dinb(n13038), .dout(n13040));
  jor  g12937(.dina(n13040), .dinb(n13037), .dout(n13041));
  jor  g12938(.dina(n13041), .dinb(n13036), .dout(n13042));
  jxor g12939(.dina(n13042), .dinb(n72), .dout(n13043));
  jor  g12940(.dina(n13043), .dinb(n13035), .dout(n13044));
  jand g12941(.dina(n12569), .dinb(n4449), .dout(n13045));
  jand g12942(.dina(n11950), .dinb(n4453), .dout(n13046));
  jand g12943(.dina(n11952), .dinb(n4457), .dout(n13047));
  jand g12944(.dina(n11954), .dinb(n4461), .dout(n13048));
  jor  g12945(.dina(n13048), .dinb(n13047), .dout(n13049));
  jor  g12946(.dina(n13049), .dinb(n13046), .dout(n13050));
  jor  g12947(.dina(n13050), .dinb(n13045), .dout(n13051));
  jxor g12948(.dina(n13051), .dinb(n88), .dout(n13052));
  jnot g12949(.din(n13052), .dout(n13053));
  jxor g12950(.dina(n12646), .dinb(n12638), .dout(n13054));
  jand g12951(.dina(n13054), .dinb(n13053), .dout(n13055));
  jand g12952(.dina(n532), .dinb(n529), .dout(n13056));
  jand g12953(.dina(n13056), .dinb(n1264), .dout(n13057));
  jand g12954(.dina(n826), .dinb(n667), .dout(n13058));
  jand g12955(.dina(n13058), .dinb(n5790), .dout(n13059));
  jand g12956(.dina(n13059), .dinb(n13057), .dout(n13060));
  jand g12957(.dina(n331), .dinb(n255), .dout(n13061));
  jand g12958(.dina(n13061), .dinb(n2315), .dout(n13062));
  jand g12959(.dina(n5165), .dinb(n3445), .dout(n13063));
  jand g12960(.dina(n13063), .dinb(n13062), .dout(n13064));
  jand g12961(.dina(n13064), .dinb(n5024), .dout(n13065));
  jand g12962(.dina(n13065), .dinb(n13060), .dout(n13066));
  jand g12963(.dina(n3662), .dinb(n3077), .dout(n13067));
  jand g12964(.dina(n2420), .dinb(n816), .dout(n13068));
  jand g12965(.dina(n13068), .dinb(n13067), .dout(n13069));
  jand g12966(.dina(n1346), .dinb(n441), .dout(n13070));
  jand g12967(.dina(n860), .dinb(n756), .dout(n13071));
  jand g12968(.dina(n13071), .dinb(n13070), .dout(n13072));
  jand g12969(.dina(n13072), .dinb(n2145), .dout(n13073));
  jand g12970(.dina(n13073), .dinb(n13069), .dout(n13074));
  jand g12971(.dina(n1305), .dinb(n1119), .dout(n13075));
  jand g12972(.dina(n913), .dinb(n434), .dout(n13076));
  jand g12973(.dina(n509), .dinb(n476), .dout(n13077));
  jand g12974(.dina(n13077), .dinb(n13076), .dout(n13078));
  jand g12975(.dina(n13078), .dinb(n13075), .dout(n13079));
  jand g12976(.dina(n12127), .dinb(n2816), .dout(n13080));
  jand g12977(.dina(n13080), .dinb(n13079), .dout(n13081));
  jand g12978(.dina(n13081), .dinb(n13074), .dout(n13082));
  jand g12979(.dina(n13082), .dinb(n13066), .dout(n13083));
  jand g12980(.dina(n13083), .dinb(n3573), .dout(n13084));
  jand g12981(.dina(n13084), .dinb(n6659), .dout(n13085));
  jand g12982(.dina(n6405), .dinb(n1420), .dout(n13086));
  jand g12983(.dina(n13086), .dinb(n1972), .dout(n13087));
  jand g12984(.dina(n553), .dinb(n161), .dout(n13088));
  jand g12985(.dina(n13088), .dinb(n692), .dout(n13089));
  jand g12986(.dina(n13089), .dinb(n3074), .dout(n13090));
  jand g12987(.dina(n13090), .dinb(n2042), .dout(n13091));
  jand g12988(.dina(n1793), .dinb(n1169), .dout(n13092));
  jand g12989(.dina(n13092), .dinb(n3104), .dout(n13093));
  jand g12990(.dina(n609), .dinb(n481), .dout(n13094));
  jand g12991(.dina(n13094), .dinb(n1840), .dout(n13095));
  jand g12992(.dina(n13095), .dinb(n2015), .dout(n13096));
  jand g12993(.dina(n893), .dinb(n311), .dout(n13097));
  jand g12994(.dina(n13097), .dinb(n3363), .dout(n13098));
  jand g12995(.dina(n13098), .dinb(n5166), .dout(n13099));
  jand g12996(.dina(n13099), .dinb(n13096), .dout(n13100));
  jand g12997(.dina(n13100), .dinb(n13093), .dout(n13101));
  jand g12998(.dina(n13101), .dinb(n13091), .dout(n13102));
  jand g12999(.dina(n13102), .dinb(n784), .dout(n13103));
  jand g13000(.dina(n13103), .dinb(n13087), .dout(n13104));
  jor  g13001(.dina(n13104), .dinb(n13085), .dout(n13105));
  jnot g13002(.din(n7886), .dout(n13106));
  jor  g13003(.dina(n7887), .dinb(n13106), .dout(n13107));
  jand g13004(.dina(n13107), .dinb(n12461), .dout(n13108));
  jxor g13005(.dina(n13108), .dinb(n5833), .dout(n13109));
  jxor g13006(.dina(n13104), .dinb(n13085), .dout(n13110));
  jand g13007(.dina(n13110), .dinb(n13109), .dout(n13111));
  jnot g13008(.din(n13111), .dout(n13112));
  jand g13009(.dina(n13112), .dinb(n13105), .dout(n13113));
  jor  g13010(.dina(n13113), .dinb(n12582), .dout(n13114));
  jxor g13011(.dina(n13113), .dinb(n12582), .dout(n13115));
  jxor g13012(.dina(n12074), .dinb(n12073), .dout(n13116));
  jand g13013(.dina(n13116), .dinb(n732), .dout(n13117));
  jand g13014(.dina(n11960), .dinb(n3855), .dout(n13118));
  jand g13015(.dina(n11964), .dinb(n3851), .dout(n13119));
  jand g13016(.dina(n11962), .dinb(n3858), .dout(n13120));
  jor  g13017(.dina(n13120), .dinb(n13119), .dout(n13121));
  jor  g13018(.dina(n13121), .dinb(n13118), .dout(n13122));
  jor  g13019(.dina(n13122), .dinb(n13117), .dout(n13123));
  jand g13020(.dina(n13123), .dinb(n13115), .dout(n13124));
  jnot g13021(.din(n13124), .dout(n13125));
  jand g13022(.dina(n13125), .dinb(n13114), .dout(n13126));
  jnot g13023(.din(n13126), .dout(n13127));
  jxor g13024(.dina(n12631), .dinb(n12623), .dout(n13128));
  jand g13025(.dina(n13128), .dinb(n13127), .dout(n13129));
  jnot g13026(.din(n13129), .dout(n13130));
  jxor g13027(.dina(n13128), .dinb(n13127), .dout(n13131));
  jnot g13028(.din(n13131), .dout(n13132));
  jxor g13029(.dina(n13110), .dinb(n13109), .dout(n13133));
  jxor g13030(.dina(n12071), .dinb(n12070), .dout(n13134));
  jand g13031(.dina(n13134), .dinb(n732), .dout(n13135));
  jand g13032(.dina(n11962), .dinb(n3855), .dout(n13136));
  jand g13033(.dina(n11964), .dinb(n3858), .dout(n13137));
  jand g13034(.dina(n11966), .dinb(n3851), .dout(n13138));
  jor  g13035(.dina(n13138), .dinb(n13137), .dout(n13139));
  jor  g13036(.dina(n13139), .dinb(n13136), .dout(n13140));
  jor  g13037(.dina(n13140), .dinb(n13135), .dout(n13141));
  jand g13038(.dina(n13141), .dinb(n13133), .dout(n13142));
  jnot g13039(.din(n13085), .dout(n13143));
  jand g13040(.dina(n392), .dinb(n161), .dout(n13144));
  jand g13041(.dina(n13144), .dinb(n354), .dout(n13145));
  jand g13042(.dina(n1264), .dinb(n424), .dout(n13146));
  jand g13043(.dina(n13146), .dinb(n1082), .dout(n13147));
  jand g13044(.dina(n13147), .dinb(n13145), .dout(n13148));
  jand g13045(.dina(n801), .dinb(n154), .dout(n13149));
  jand g13046(.dina(n515), .dinb(n418), .dout(n13150));
  jand g13047(.dina(n13150), .dinb(n13149), .dout(n13151));
  jand g13048(.dina(n13151), .dinb(n5248), .dout(n13152));
  jand g13049(.dina(n13152), .dinb(n13148), .dout(n13153));
  jand g13050(.dina(n2239), .dinb(n2228), .dout(n13154));
  jand g13051(.dina(n2292), .dinb(n1025), .dout(n13155));
  jand g13052(.dina(n13155), .dinb(n13154), .dout(n13156));
  jand g13053(.dina(n13156), .dinb(n3508), .dout(n13157));
  jand g13054(.dina(n865), .dinb(n716), .dout(n13158));
  jand g13055(.dina(n13158), .dinb(n562), .dout(n13159));
  jand g13056(.dina(n13159), .dinb(n1506), .dout(n13160));
  jand g13057(.dina(n13160), .dinb(n1061), .dout(n13161));
  jand g13058(.dina(n13161), .dinb(n13157), .dout(n13162));
  jand g13059(.dina(n13162), .dinb(n13153), .dout(n13163));
  jand g13060(.dina(n13163), .dinb(n2747), .dout(n13164));
  jand g13061(.dina(n12723), .dinb(n2118), .dout(n13165));
  jand g13062(.dina(n13165), .dinb(n1584), .dout(n13166));
  jand g13063(.dina(n860), .dinb(n396), .dout(n13167));
  jand g13064(.dina(n13167), .dinb(n417), .dout(n13168));
  jand g13065(.dina(n5760), .dinb(n659), .dout(n13169));
  jand g13066(.dina(n13169), .dinb(n13168), .dout(n13170));
  jand g13067(.dina(n13170), .dinb(n13166), .dout(n13171));
  jand g13068(.dina(n4382), .dinb(n558), .dout(n13172));
  jand g13069(.dina(n1409), .dinb(n529), .dout(n13173));
  jand g13070(.dina(n13173), .dinb(n914), .dout(n13174));
  jand g13071(.dina(n13174), .dinb(n13172), .dout(n13175));
  jand g13072(.dina(n492), .dinb(n348), .dout(n13176));
  jand g13073(.dina(n449), .dinb(n190), .dout(n13177));
  jand g13074(.dina(n13177), .dinb(n13176), .dout(n13178));
  jand g13075(.dina(n3550), .dinb(n501), .dout(n13179));
  jand g13076(.dina(n13179), .dinb(n13178), .dout(n13180));
  jand g13077(.dina(n2490), .dinb(n1049), .dout(n13181));
  jand g13078(.dina(n13181), .dinb(n13180), .dout(n13182));
  jand g13079(.dina(n13182), .dinb(n13175), .dout(n13183));
  jand g13080(.dina(n13183), .dinb(n13171), .dout(n13184));
  jand g13081(.dina(n13184), .dinb(n5136), .dout(n13185));
  jand g13082(.dina(n13185), .dinb(n13164), .dout(n13186));
  jor  g13083(.dina(n13186), .dinb(n13143), .dout(n13187));
  jand g13084(.dina(n3462), .dinb(n501), .dout(n13188));
  jand g13085(.dina(n13188), .dinb(n802), .dout(n13189));
  jand g13086(.dina(n701), .dinb(n161), .dout(n13190));
  jand g13087(.dina(n13190), .dinb(n409), .dout(n13191));
  jand g13088(.dina(n2859), .dinb(n1249), .dout(n13192));
  jand g13089(.dina(n13192), .dinb(n13191), .dout(n13193));
  jand g13090(.dina(n13193), .dinb(n13189), .dout(n13194));
  jand g13091(.dina(n13194), .dinb(n4153), .dout(n13195));
  jand g13092(.dina(n515), .dinb(n470), .dout(n13196));
  jand g13093(.dina(n1135), .dinb(n923), .dout(n13197));
  jand g13094(.dina(n13197), .dinb(n13196), .dout(n13198));
  jand g13095(.dina(n1031), .dinb(n450), .dout(n13199));
  jand g13096(.dina(n13199), .dinb(n1295), .dout(n13200));
  jand g13097(.dina(n979), .dinb(n708), .dout(n13201));
  jand g13098(.dina(n13201), .dinb(n543), .dout(n13202));
  jand g13099(.dina(n13202), .dinb(n13200), .dout(n13203));
  jand g13100(.dina(n13203), .dinb(n13198), .dout(n13204));
  jand g13101(.dina(n3261), .dinb(n1124), .dout(n13205));
  jand g13102(.dina(n13205), .dinb(n1336), .dout(n13206));
  jand g13103(.dina(n13206), .dinb(n13204), .dout(n13207));
  jand g13104(.dina(n13207), .dinb(n13195), .dout(n13208));
  jand g13105(.dina(n6667), .dinb(n818), .dout(n13209));
  jand g13106(.dina(n13209), .dinb(n2022), .dout(n13210));
  jnot g13107(.din(n1373), .dout(n13211));
  jand g13108(.dina(n805), .dinb(n465), .dout(n13212));
  jand g13109(.dina(n865), .dinb(n607), .dout(n13213));
  jand g13110(.dina(n13213), .dinb(n13212), .dout(n13214));
  jand g13111(.dina(n13214), .dinb(n13211), .dout(n13215));
  jand g13112(.dina(n13215), .dinb(n12548), .dout(n13216));
  jand g13113(.dina(n13216), .dinb(n13210), .dout(n13217));
  jand g13114(.dina(n1475), .dinb(n384), .dout(n13218));
  jand g13115(.dina(n13218), .dinb(n1537), .dout(n13219));
  jand g13116(.dina(n230), .dinb(n165), .dout(n13220));
  jand g13117(.dina(n13220), .dinb(n190), .dout(n13221));
  jand g13118(.dina(n3041), .dinb(n2962), .dout(n13222));
  jand g13119(.dina(n13222), .dinb(n13221), .dout(n13223));
  jand g13120(.dina(n5019), .dinb(n2201), .dout(n13224));
  jand g13121(.dina(n13224), .dinb(n13223), .dout(n13225));
  jand g13122(.dina(n13225), .dinb(n13219), .dout(n13226));
  jand g13123(.dina(n13226), .dinb(n13217), .dout(n13227));
  jand g13124(.dina(n13227), .dinb(n13208), .dout(n13228));
  jand g13125(.dina(n13228), .dinb(n3180), .dout(n13229));
  jand g13126(.dina(n687), .dinb(n434), .dout(n13230));
  jand g13127(.dina(n13230), .dinb(n2420), .dout(n13231));
  jand g13128(.dina(n1730), .dinb(n868), .dout(n13232));
  jand g13129(.dina(n13232), .dinb(n13231), .dout(n13233));
  jand g13130(.dina(n13233), .dinb(n2516), .dout(n13234));
  jand g13131(.dina(n13234), .dinb(n2842), .dout(n13235));
  jand g13132(.dina(n759), .dinb(n208), .dout(n13236));
  jand g13133(.dina(n1034), .dinb(n609), .dout(n13237));
  jand g13134(.dina(n13237), .dinb(n13236), .dout(n13238));
  jand g13135(.dina(n392), .dinb(n357), .dout(n13239));
  jand g13136(.dina(n13239), .dinb(n109), .dout(n13240));
  jand g13137(.dina(n13240), .dinb(n13238), .dout(n13241));
  jand g13138(.dina(n5734), .dinb(n1613), .dout(n13242));
  jand g13139(.dina(n13242), .dinb(n13241), .dout(n13243));
  jand g13140(.dina(n805), .dinb(n280), .dout(n13244));
  jand g13141(.dina(n13244), .dinb(n979), .dout(n13245));
  jand g13142(.dina(n508), .dinb(n386), .dout(n13246));
  jand g13143(.dina(n13246), .dinb(n5268), .dout(n13247));
  jand g13144(.dina(n13247), .dinb(n13245), .dout(n13248));
  jand g13145(.dina(n2526), .dinb(n451), .dout(n13249));
  jand g13146(.dina(n13249), .dinb(n3154), .dout(n13250));
  jand g13147(.dina(n13250), .dinb(n2699), .dout(n13251));
  jand g13148(.dina(n13251), .dinb(n13248), .dout(n13252));
  jand g13149(.dina(n13252), .dinb(n13243), .dout(n13253));
  jand g13150(.dina(n13253), .dinb(n13235), .dout(n13254));
  jand g13151(.dina(n4499), .dinb(n2040), .dout(n13255));
  jand g13152(.dina(n13255), .dinb(n13254), .dout(n13256));
  jor  g13153(.dina(n13256), .dinb(n13229), .dout(n13257));
  jnot g13154(.din(n8767), .dout(n13258));
  jor  g13155(.dina(n8768), .dinb(n13258), .dout(n13259));
  jand g13156(.dina(n13259), .dinb(n12461), .dout(n13260));
  jxor g13157(.dina(n13260), .dinb(n6039), .dout(n13261));
  jxor g13158(.dina(n13256), .dinb(n13229), .dout(n13262));
  jand g13159(.dina(n13262), .dinb(n13261), .dout(n13263));
  jnot g13160(.din(n13263), .dout(n13264));
  jand g13161(.dina(n13264), .dinb(n13257), .dout(n13265));
  jor  g13162(.dina(n13265), .dinb(n13143), .dout(n13266));
  jxor g13163(.dina(n13265), .dinb(n13143), .dout(n13267));
  jxor g13164(.dina(n12065), .dinb(n12064), .dout(n13268));
  jand g13165(.dina(n13268), .dinb(n732), .dout(n13269));
  jand g13166(.dina(n11966), .dinb(n3855), .dout(n13270));
  jand g13167(.dina(n11970), .dinb(n3851), .dout(n13271));
  jand g13168(.dina(n11968), .dinb(n3858), .dout(n13272));
  jor  g13169(.dina(n13272), .dinb(n13271), .dout(n13273));
  jor  g13170(.dina(n13273), .dinb(n13270), .dout(n13274));
  jor  g13171(.dina(n13274), .dinb(n13269), .dout(n13275));
  jand g13172(.dina(n13275), .dinb(n13267), .dout(n13276));
  jnot g13173(.din(n13276), .dout(n13277));
  jand g13174(.dina(n13277), .dinb(n13266), .dout(n13278));
  jnot g13175(.din(n13278), .dout(n13279));
  jxor g13176(.dina(n13186), .dinb(n13143), .dout(n13280));
  jand g13177(.dina(n13280), .dinb(n13279), .dout(n13281));
  jnot g13178(.din(n13281), .dout(n13282));
  jand g13179(.dina(n13282), .dinb(n13187), .dout(n13283));
  jnot g13180(.din(n13283), .dout(n13284));
  jxor g13181(.dina(n13141), .dinb(n13133), .dout(n13285));
  jand g13182(.dina(n13285), .dinb(n13284), .dout(n13286));
  jor  g13183(.dina(n13286), .dinb(n13142), .dout(n13287));
  jxor g13184(.dina(n13123), .dinb(n13115), .dout(n13288));
  jand g13185(.dina(n13288), .dinb(n13287), .dout(n13289));
  jnot g13186(.din(n13289), .dout(n13290));
  jxor g13187(.dina(n13288), .dinb(n13287), .dout(n13291));
  jnot g13188(.din(n13291), .dout(n13292));
  jand g13189(.dina(n12472), .dinb(n4449), .dout(n13293));
  jand g13190(.dina(n11954), .dinb(n4453), .dout(n13294));
  jand g13191(.dina(n11956), .dinb(n4457), .dout(n13295));
  jand g13192(.dina(n11958), .dinb(n4461), .dout(n13296));
  jor  g13193(.dina(n13296), .dinb(n13295), .dout(n13297));
  jor  g13194(.dina(n13297), .dinb(n13294), .dout(n13298));
  jor  g13195(.dina(n13298), .dinb(n13293), .dout(n13299));
  jxor g13196(.dina(n13299), .dinb(n88), .dout(n13300));
  jor  g13197(.dina(n13300), .dinb(n13292), .dout(n13301));
  jand g13198(.dina(n13301), .dinb(n13290), .dout(n13302));
  jor  g13199(.dina(n13302), .dinb(n13132), .dout(n13303));
  jand g13200(.dina(n13303), .dinb(n13130), .dout(n13304));
  jnot g13201(.din(n13304), .dout(n13305));
  jxor g13202(.dina(n13054), .dinb(n13053), .dout(n13306));
  jand g13203(.dina(n13306), .dinb(n13305), .dout(n13307));
  jor  g13204(.dina(n13307), .dinb(n13055), .dout(n13308));
  jxor g13205(.dina(n12662), .dinb(n12653), .dout(n13309));
  jand g13206(.dina(n13309), .dinb(n13308), .dout(n13310));
  jnot g13207(.din(n13310), .dout(n13311));
  jxor g13208(.dina(n13309), .dinb(n13308), .dout(n13312));
  jnot g13209(.din(n13312), .dout(n13313));
  jand g13210(.dina(n12751), .dinb(n75), .dout(n13314));
  jand g13211(.dina(n11942), .dinb(n4933), .dout(n13315));
  jand g13212(.dina(n11944), .dinb(n4918), .dout(n13316));
  jand g13213(.dina(n11946), .dinb(n4745), .dout(n13317));
  jor  g13214(.dina(n13317), .dinb(n13316), .dout(n13318));
  jor  g13215(.dina(n13318), .dinb(n13315), .dout(n13319));
  jor  g13216(.dina(n13319), .dinb(n13314), .dout(n13320));
  jxor g13217(.dina(n13320), .dinb(n68), .dout(n13321));
  jor  g13218(.dina(n13321), .dinb(n13313), .dout(n13322));
  jand g13219(.dina(n13322), .dinb(n13311), .dout(n13323));
  jnot g13220(.din(n13323), .dout(n13324));
  jxor g13221(.dina(n12679), .dinb(n12670), .dout(n13325));
  jand g13222(.dina(n13325), .dinb(n13324), .dout(n13326));
  jnot g13223(.din(n13326), .dout(n13327));
  jxor g13224(.dina(n13325), .dinb(n13324), .dout(n13328));
  jnot g13225(.din(n13328), .dout(n13329));
  jand g13226(.dina(n12841), .dinb(n5365), .dout(n13330));
  jand g13227(.dina(n12783), .dinb(n5500), .dout(n13331));
  jand g13228(.dina(n12766), .dinb(n5424), .dout(n13332));
  jand g13229(.dina(n12177), .dinb(n5363), .dout(n13333));
  jor  g13230(.dina(n13333), .dinb(n13332), .dout(n13334));
  jor  g13231(.dina(n13334), .dinb(n13331), .dout(n13335));
  jor  g13232(.dina(n13335), .dinb(n13330), .dout(n13336));
  jxor g13233(.dina(n13336), .dinb(n72), .dout(n13337));
  jor  g13234(.dina(n13337), .dinb(n13329), .dout(n13338));
  jand g13235(.dina(n13338), .dinb(n13327), .dout(n13339));
  jnot g13236(.din(n13339), .dout(n13340));
  jxor g13237(.dina(n13043), .dinb(n13035), .dout(n13341));
  jand g13238(.dina(n13341), .dinb(n13340), .dout(n13342));
  jnot g13239(.din(n13342), .dout(n13343));
  jand g13240(.dina(n13343), .dinb(n13044), .dout(n13344));
  jnot g13241(.din(n13344), .dout(n13345));
  jxor g13242(.dina(n12805), .dinb(n12781), .dout(n13346));
  jand g13243(.dina(n13346), .dinb(n13345), .dout(n13347));
  jnot g13244(.din(n13347), .dout(n13348));
  jxor g13245(.dina(n13346), .dinb(n13345), .dout(n13349));
  jnot g13246(.din(n13349), .dout(n13350));
  jor  g13247(.dina(n13021), .dinb(n12815), .dout(n13352));
  jand g13248(.dina(n13352), .dinb(n12825), .dout(n13353));
  jnot g13249(.din(n13353), .dout(n13354));
  jor  g13250(.dina(n12814), .dinb(n5692), .dout(n13356));
  jand g13251(.dina(n12829), .dinb(n13356), .dout(n13360));
  jand g13252(.dina(n13360), .dinb(n5694), .dout(n13361));
  jxor g13253(.dina(n13361), .dinb(\a[20] ), .dout(n13362));
  jor  g13254(.dina(n13362), .dinb(n13350), .dout(n13363));
  jand g13255(.dina(n13363), .dinb(n13348), .dout(n13364));
  jnot g13256(.din(n13364), .dout(n13365));
  jxor g13257(.dina(n12928), .dinb(n12835), .dout(n13366));
  jand g13258(.dina(n13366), .dinb(n13365), .dout(n13367));
  jxor g13259(.dina(n13366), .dinb(n13365), .dout(n13368));
  jxor g13260(.dina(n13306), .dinb(n13305), .dout(n13369));
  jnot g13261(.din(n13369), .dout(n13370));
  jand g13262(.dina(n12189), .dinb(n75), .dout(n13371));
  jand g13263(.dina(n11944), .dinb(n4933), .dout(n13372));
  jand g13264(.dina(n11946), .dinb(n4918), .dout(n13373));
  jand g13265(.dina(n11948), .dinb(n4745), .dout(n13374));
  jor  g13266(.dina(n13374), .dinb(n13373), .dout(n13375));
  jor  g13267(.dina(n13375), .dinb(n13372), .dout(n13376));
  jor  g13268(.dina(n13376), .dinb(n13371), .dout(n13377));
  jxor g13269(.dina(n13377), .dinb(n68), .dout(n13378));
  jor  g13270(.dina(n13378), .dinb(n13370), .dout(n13379));
  jxor g13271(.dina(n13302), .dinb(n13132), .dout(n13380));
  jnot g13272(.din(n13380), .dout(n13381));
  jand g13273(.dina(n12510), .dinb(n4449), .dout(n13382));
  jand g13274(.dina(n11952), .dinb(n4453), .dout(n13383));
  jand g13275(.dina(n11954), .dinb(n4457), .dout(n13384));
  jand g13276(.dina(n11956), .dinb(n4461), .dout(n13385));
  jor  g13277(.dina(n13385), .dinb(n13384), .dout(n13386));
  jor  g13278(.dina(n13386), .dinb(n13383), .dout(n13387));
  jor  g13279(.dina(n13387), .dinb(n13382), .dout(n13388));
  jxor g13280(.dina(n13388), .dinb(n88), .dout(n13389));
  jor  g13281(.dina(n13389), .dinb(n13381), .dout(n13390));
  jand g13282(.dina(n12519), .dinb(n75), .dout(n13391));
  jand g13283(.dina(n11946), .dinb(n4933), .dout(n13392));
  jand g13284(.dina(n11948), .dinb(n4918), .dout(n13393));
  jand g13285(.dina(n11950), .dinb(n4745), .dout(n13394));
  jor  g13286(.dina(n13394), .dinb(n13393), .dout(n13395));
  jor  g13287(.dina(n13395), .dinb(n13392), .dout(n13396));
  jor  g13288(.dina(n13396), .dinb(n13391), .dout(n13397));
  jxor g13289(.dina(n13397), .dinb(n68), .dout(n13398));
  jnot g13290(.din(n13398), .dout(n13399));
  jxor g13291(.dina(n13389), .dinb(n13381), .dout(n13400));
  jand g13292(.dina(n13400), .dinb(n13399), .dout(n13401));
  jnot g13293(.din(n13401), .dout(n13402));
  jand g13294(.dina(n13402), .dinb(n13390), .dout(n13403));
  jnot g13295(.din(n13403), .dout(n13404));
  jxor g13296(.dina(n13378), .dinb(n13370), .dout(n13405));
  jand g13297(.dina(n13405), .dinb(n13404), .dout(n13406));
  jnot g13298(.din(n13406), .dout(n13407));
  jand g13299(.dina(n13407), .dinb(n13379), .dout(n13408));
  jnot g13300(.din(n13408), .dout(n13409));
  jxor g13301(.dina(n13321), .dinb(n13313), .dout(n13410));
  jand g13302(.dina(n13410), .dinb(n13409), .dout(n13411));
  jnot g13303(.din(n13411), .dout(n13412));
  jxor g13304(.dina(n13410), .dinb(n13409), .dout(n13413));
  jnot g13305(.din(n13413), .dout(n13414));
  jand g13306(.dina(n12768), .dinb(n5365), .dout(n13415));
  jand g13307(.dina(n12766), .dinb(n5500), .dout(n13416));
  jand g13308(.dina(n12177), .dinb(n5424), .dout(n13417));
  jand g13309(.dina(n11941), .dinb(n5363), .dout(n13418));
  jor  g13310(.dina(n13418), .dinb(n13417), .dout(n13419));
  jor  g13311(.dina(n13419), .dinb(n13416), .dout(n13420));
  jor  g13312(.dina(n13420), .dinb(n13415), .dout(n13421));
  jxor g13313(.dina(n13421), .dinb(n72), .dout(n13422));
  jor  g13314(.dina(n13422), .dinb(n13414), .dout(n13423));
  jand g13315(.dina(n13423), .dinb(n13412), .dout(n13424));
  jnot g13316(.din(n13424), .dout(n13425));
  jxor g13317(.dina(n13337), .dinb(n13329), .dout(n13426));
  jand g13318(.dina(n13426), .dinb(n13425), .dout(n13427));
  jnot g13319(.din(n13427), .dout(n13428));
  jxor g13320(.dina(n13426), .dinb(n13425), .dout(n13429));
  jnot g13321(.din(n13429), .dout(n13430));
  jand g13322(.dina(n12919), .dinb(n5693), .dout(n13431));
  jand g13323(.dina(n12815), .dinb(n6209), .dout(n13432));
  jand g13324(.dina(n12795), .dinb(n6131), .dout(n13433));
  jand g13325(.dina(n12782), .dinb(n5691), .dout(n13434));
  jor  g13326(.dina(n13434), .dinb(n13433), .dout(n13435));
  jor  g13327(.dina(n13435), .dinb(n13432), .dout(n13436));
  jor  g13328(.dina(n13436), .dinb(n13431), .dout(n13437));
  jxor g13329(.dina(n13437), .dinb(n4247), .dout(n13438));
  jor  g13330(.dina(n13438), .dinb(n13430), .dout(n13439));
  jand g13331(.dina(n13439), .dinb(n13428), .dout(n13440));
  jand g13332(.dina(n13022), .dinb(n5693), .dout(n13441));
  jand g13333(.dina(n12811), .dinb(n6209), .dout(n13442));
  jand g13334(.dina(n12815), .dinb(n6131), .dout(n13443));
  jand g13335(.dina(n12795), .dinb(n5691), .dout(n13444));
  jor  g13336(.dina(n13444), .dinb(n13443), .dout(n13445));
  jor  g13337(.dina(n13445), .dinb(n13442), .dout(n13446));
  jor  g13338(.dina(n13446), .dinb(n13441), .dout(n13447));
  jxor g13339(.dina(n13447), .dinb(n4247), .dout(n13448));
  jor  g13340(.dina(n13448), .dinb(n13440), .dout(n13449));
  jxor g13341(.dina(n13341), .dinb(n13340), .dout(n13450));
  jxor g13342(.dina(n13448), .dinb(n13440), .dout(n13451));
  jand g13343(.dina(n13451), .dinb(n13450), .dout(n13452));
  jnot g13344(.din(n13452), .dout(n13453));
  jand g13345(.dina(n13453), .dinb(n13449), .dout(n13454));
  jnot g13346(.din(n13454), .dout(n13455));
  jxor g13347(.dina(n13362), .dinb(n13350), .dout(n13456));
  jand g13348(.dina(n13456), .dinb(n13455), .dout(n13457));
  jxor g13349(.dina(n13405), .dinb(n13404), .dout(n13458));
  jnot g13350(.din(n13458), .dout(n13459));
  jand g13351(.dina(n12179), .dinb(n5365), .dout(n13460));
  jand g13352(.dina(n12177), .dinb(n5500), .dout(n13461));
  jand g13353(.dina(n11941), .dinb(n5424), .dout(n13462));
  jand g13354(.dina(n11942), .dinb(n5363), .dout(n13463));
  jor  g13355(.dina(n13463), .dinb(n13462), .dout(n13464));
  jor  g13356(.dina(n13464), .dinb(n13461), .dout(n13465));
  jor  g13357(.dina(n13465), .dinb(n13460), .dout(n13466));
  jxor g13358(.dina(n13466), .dinb(n72), .dout(n13467));
  jor  g13359(.dina(n13467), .dinb(n13459), .dout(n13468));
  jxor g13360(.dina(n13280), .dinb(n13279), .dout(n13469));
  jxor g13361(.dina(n12068), .dinb(n12067), .dout(n13470));
  jand g13362(.dina(n13470), .dinb(n732), .dout(n13471));
  jand g13363(.dina(n11964), .dinb(n3855), .dout(n13472));
  jand g13364(.dina(n11966), .dinb(n3858), .dout(n13473));
  jand g13365(.dina(n11968), .dinb(n3851), .dout(n13474));
  jor  g13366(.dina(n13474), .dinb(n13473), .dout(n13475));
  jor  g13367(.dina(n13475), .dinb(n13472), .dout(n13476));
  jor  g13368(.dina(n13476), .dinb(n13471), .dout(n13477));
  jand g13369(.dina(n13477), .dinb(n13469), .dout(n13478));
  jand g13370(.dina(n12624), .dinb(n4449), .dout(n13479));
  jand g13371(.dina(n11958), .dinb(n4453), .dout(n13480));
  jand g13372(.dina(n11960), .dinb(n4457), .dout(n13481));
  jand g13373(.dina(n11962), .dinb(n4461), .dout(n13482));
  jor  g13374(.dina(n13482), .dinb(n13481), .dout(n13483));
  jor  g13375(.dina(n13483), .dinb(n13480), .dout(n13484));
  jor  g13376(.dina(n13484), .dinb(n13479), .dout(n13485));
  jxor g13377(.dina(n13485), .dinb(n88), .dout(n13486));
  jnot g13378(.din(n13486), .dout(n13487));
  jxor g13379(.dina(n13477), .dinb(n13469), .dout(n13488));
  jand g13380(.dina(n13488), .dinb(n13487), .dout(n13489));
  jor  g13381(.dina(n13489), .dinb(n13478), .dout(n13490));
  jxor g13382(.dina(n13285), .dinb(n13284), .dout(n13491));
  jand g13383(.dina(n13491), .dinb(n13490), .dout(n13492));
  jand g13384(.dina(n12639), .dinb(n4449), .dout(n13493));
  jand g13385(.dina(n11956), .dinb(n4453), .dout(n13494));
  jand g13386(.dina(n11958), .dinb(n4457), .dout(n13495));
  jand g13387(.dina(n11960), .dinb(n4461), .dout(n13496));
  jor  g13388(.dina(n13496), .dinb(n13495), .dout(n13497));
  jor  g13389(.dina(n13497), .dinb(n13494), .dout(n13498));
  jor  g13390(.dina(n13498), .dinb(n13493), .dout(n13499));
  jxor g13391(.dina(n13499), .dinb(n88), .dout(n13500));
  jnot g13392(.din(n13500), .dout(n13501));
  jxor g13393(.dina(n13491), .dinb(n13490), .dout(n13502));
  jand g13394(.dina(n13502), .dinb(n13501), .dout(n13503));
  jor  g13395(.dina(n13503), .dinb(n13492), .dout(n13504));
  jxor g13396(.dina(n13300), .dinb(n13292), .dout(n13505));
  jand g13397(.dina(n13505), .dinb(n13504), .dout(n13506));
  jnot g13398(.din(n13506), .dout(n13507));
  jxor g13399(.dina(n13505), .dinb(n13504), .dout(n13508));
  jnot g13400(.din(n13508), .dout(n13509));
  jand g13401(.dina(n12654), .dinb(n75), .dout(n13510));
  jand g13402(.dina(n11948), .dinb(n4933), .dout(n13511));
  jand g13403(.dina(n11950), .dinb(n4918), .dout(n13512));
  jand g13404(.dina(n11952), .dinb(n4745), .dout(n13513));
  jor  g13405(.dina(n13513), .dinb(n13512), .dout(n13514));
  jor  g13406(.dina(n13514), .dinb(n13511), .dout(n13515));
  jor  g13407(.dina(n13515), .dinb(n13510), .dout(n13516));
  jxor g13408(.dina(n13516), .dinb(n68), .dout(n13517));
  jor  g13409(.dina(n13517), .dinb(n13509), .dout(n13518));
  jand g13410(.dina(n13518), .dinb(n13507), .dout(n13519));
  jnot g13411(.din(n13519), .dout(n13520));
  jxor g13412(.dina(n13400), .dinb(n13399), .dout(n13521));
  jand g13413(.dina(n13521), .dinb(n13520), .dout(n13522));
  jnot g13414(.din(n13522), .dout(n13523));
  jxor g13415(.dina(n13521), .dinb(n13520), .dout(n13524));
  jnot g13416(.din(n13524), .dout(n13525));
  jand g13417(.dina(n12671), .dinb(n5365), .dout(n13526));
  jand g13418(.dina(n11941), .dinb(n5500), .dout(n13527));
  jand g13419(.dina(n11942), .dinb(n5424), .dout(n13528));
  jand g13420(.dina(n11944), .dinb(n5363), .dout(n13529));
  jor  g13421(.dina(n13529), .dinb(n13528), .dout(n13530));
  jor  g13422(.dina(n13530), .dinb(n13527), .dout(n13531));
  jor  g13423(.dina(n13531), .dinb(n13526), .dout(n13532));
  jxor g13424(.dina(n13532), .dinb(n72), .dout(n13533));
  jor  g13425(.dina(n13533), .dinb(n13525), .dout(n13534));
  jand g13426(.dina(n13534), .dinb(n13523), .dout(n13535));
  jnot g13427(.din(n13535), .dout(n13536));
  jxor g13428(.dina(n13467), .dinb(n13459), .dout(n13537));
  jand g13429(.dina(n13537), .dinb(n13536), .dout(n13538));
  jnot g13430(.din(n13538), .dout(n13539));
  jand g13431(.dina(n13539), .dinb(n13468), .dout(n13540));
  jnot g13432(.din(n13540), .dout(n13541));
  jxor g13433(.dina(n13422), .dinb(n13414), .dout(n13542));
  jand g13434(.dina(n13542), .dinb(n13541), .dout(n13543));
  jnot g13435(.din(n13543), .dout(n13544));
  jxor g13436(.dina(n13542), .dinb(n13541), .dout(n13545));
  jnot g13437(.din(n13545), .dout(n13546));
  jand g13438(.dina(n12797), .dinb(n5693), .dout(n13547));
  jand g13439(.dina(n12795), .dinb(n6209), .dout(n13548));
  jand g13440(.dina(n12782), .dinb(n6131), .dout(n13549));
  jand g13441(.dina(n12783), .dinb(n5691), .dout(n13550));
  jor  g13442(.dina(n13550), .dinb(n13549), .dout(n13551));
  jor  g13443(.dina(n13551), .dinb(n13548), .dout(n13552));
  jor  g13444(.dina(n13552), .dinb(n13547), .dout(n13553));
  jxor g13445(.dina(n13553), .dinb(n4247), .dout(n13554));
  jor  g13446(.dina(n13554), .dinb(n13546), .dout(n13555));
  jand g13447(.dina(n13555), .dinb(n13544), .dout(n13556));
  jand g13448(.dina(n6797), .dinb(n6557), .dout(n13559));
  jor  g13449(.dina(n12538), .dinb(n13556), .dout(n13564));
  jxor g13450(.dina(n12538), .dinb(n13556), .dout(n13565));
  jxor g13451(.dina(n13438), .dinb(n13430), .dout(n13566));
  jand g13452(.dina(n13566), .dinb(n13565), .dout(n13567));
  jnot g13453(.din(n13567), .dout(n13568));
  jand g13454(.dina(n13568), .dinb(n13564), .dout(n13569));
  jnot g13455(.din(n13569), .dout(n13570));
  jxor g13456(.dina(n13451), .dinb(n13450), .dout(n13571));
  jand g13457(.dina(n13571), .dinb(n13570), .dout(n13572));
  jxor g13458(.dina(n13537), .dinb(n13536), .dout(n13573));
  jnot g13459(.din(n13573), .dout(n13574));
  jand g13460(.dina(n12938), .dinb(n5693), .dout(n13575));
  jand g13461(.dina(n12782), .dinb(n6209), .dout(n13576));
  jand g13462(.dina(n12783), .dinb(n6131), .dout(n13577));
  jand g13463(.dina(n12766), .dinb(n5691), .dout(n13578));
  jor  g13464(.dina(n13578), .dinb(n13577), .dout(n13579));
  jor  g13465(.dina(n13579), .dinb(n13576), .dout(n13580));
  jor  g13466(.dina(n13580), .dinb(n13575), .dout(n13581));
  jxor g13467(.dina(n13581), .dinb(n4247), .dout(n13582));
  jor  g13468(.dina(n13582), .dinb(n13574), .dout(n13583));
  jand g13469(.dina(n12569), .dinb(n75), .dout(n13584));
  jand g13470(.dina(n11950), .dinb(n4933), .dout(n13585));
  jand g13471(.dina(n11952), .dinb(n4918), .dout(n13586));
  jand g13472(.dina(n11954), .dinb(n4745), .dout(n13587));
  jor  g13473(.dina(n13587), .dinb(n13586), .dout(n13588));
  jor  g13474(.dina(n13588), .dinb(n13585), .dout(n13589));
  jor  g13475(.dina(n13589), .dinb(n13584), .dout(n13590));
  jxor g13476(.dina(n13590), .dinb(n68), .dout(n13591));
  jnot g13477(.din(n13591), .dout(n13592));
  jxor g13478(.dina(n13502), .dinb(n13501), .dout(n13593));
  jand g13479(.dina(n13593), .dinb(n13592), .dout(n13594));
  jnot g13480(.din(n13229), .dout(n13595));
  jand g13481(.dina(n331), .dinb(n190), .dout(n13596));
  jand g13482(.dina(n13596), .dinb(n5230), .dout(n13597));
  jand g13483(.dina(n3544), .dinb(n2870), .dout(n13598));
  jand g13484(.dina(n13598), .dinb(n13597), .dout(n13599));
  jand g13485(.dina(n12205), .dinb(n2041), .dout(n13600));
  jand g13486(.dina(n13600), .dinb(n5956), .dout(n13601));
  jand g13487(.dina(n13601), .dinb(n13599), .dout(n13602));
  jand g13488(.dina(n827), .dinb(n596), .dout(n13603));
  jand g13489(.dina(n4567), .dinb(n1416), .dout(n13604));
  jand g13490(.dina(n13604), .dinb(n13603), .dout(n13605));
  jand g13491(.dina(n13605), .dinb(n956), .dout(n13606));
  jand g13492(.dina(n13606), .dinb(n13602), .dout(n13607));
  jand g13493(.dina(n13607), .dinb(n1046), .dout(n13608));
  jand g13494(.dina(n13608), .dinb(n2765), .dout(n13609));
  jand g13495(.dina(n13609), .dinb(n2636), .dout(n13610));
  jor  g13496(.dina(n13610), .dinb(n13595), .dout(n13611));
  jand g13497(.dina(n470), .dinb(n290), .dout(n13612));
  jand g13498(.dina(n13612), .dinb(n302), .dout(n13613));
  jand g13499(.dina(n671), .dinb(n311), .dout(n13614));
  jand g13500(.dina(n13614), .dinb(n2022), .dout(n13615));
  jand g13501(.dina(n1296), .dinb(n258), .dout(n13616));
  jand g13502(.dina(n13616), .dinb(n13615), .dout(n13617));
  jand g13503(.dina(n13617), .dinb(n13613), .dout(n13618));
  jand g13504(.dina(n1034), .dinb(n997), .dout(n13619));
  jand g13505(.dina(n13619), .dinb(n3896), .dout(n13620));
  jand g13506(.dina(n13620), .dinb(n2565), .dout(n13621));
  jand g13507(.dina(n13621), .dinb(n1018), .dout(n13622));
  jand g13508(.dina(n13622), .dinb(n13618), .dout(n13623));
  jand g13509(.dina(n1409), .dinb(n739), .dout(n13624));
  jand g13510(.dina(n13624), .dinb(n1185), .dout(n13625));
  jand g13511(.dina(n13625), .dinb(n13151), .dout(n13626));
  jand g13512(.dina(n4192), .dinb(n2672), .dout(n13627));
  jand g13513(.dina(n13627), .dinb(n639), .dout(n13628));
  jand g13514(.dina(n13628), .dinb(n13626), .dout(n13629));
  jand g13515(.dina(n12272), .dinb(n1878), .dout(n13630));
  jand g13516(.dina(n3010), .dinb(n1389), .dout(n13631));
  jand g13517(.dina(n13631), .dinb(n13630), .dout(n13632));
  jand g13518(.dina(n13632), .dinb(n3437), .dout(n13633));
  jand g13519(.dina(n13633), .dinb(n13629), .dout(n13634));
  jand g13520(.dina(n13634), .dinb(n13623), .dout(n13635));
  jand g13521(.dina(n3865), .dinb(n1350), .dout(n13636));
  jand g13522(.dina(n3448), .dinb(n253), .dout(n13637));
  jand g13523(.dina(n13637), .dinb(n13636), .dout(n13638));
  jand g13524(.dina(n439), .dinb(n348), .dout(n13639));
  jand g13525(.dina(n13639), .dinb(n877), .dout(n13640));
  jand g13526(.dina(n13640), .dinb(n4190), .dout(n13641));
  jand g13527(.dina(n13641), .dinb(n13638), .dout(n13642));
  jand g13528(.dina(n7163), .dinb(n6669), .dout(n13643));
  jand g13529(.dina(n13643), .dinb(n13642), .dout(n13644));
  jand g13530(.dina(n13074), .dinb(n3992), .dout(n13645));
  jand g13531(.dina(n13645), .dinb(n13644), .dout(n13646));
  jand g13532(.dina(n13646), .dinb(n13635), .dout(n13647));
  jnot g13533(.din(n13647), .dout(n13648));
  jand g13534(.dina(n11466), .dinb(n6600), .dout(n13649));
  jnot g13535(.din(n13649), .dout(n13650));
  jand g13536(.dina(n13650), .dinb(n12461), .dout(n13651));
  jand g13537(.dina(n12460), .dinb(n6600), .dout(n13652));
  jor  g13538(.dina(n13652), .dinb(n13651), .dout(n13653));
  jand g13539(.dina(n13653), .dinb(n13648), .dout(n13654));
  jnot g13540(.din(n9916), .dout(n13655));
  jor  g13541(.dina(n13655), .dinb(n66), .dout(n13656));
  jand g13542(.dina(n13656), .dinb(n12461), .dout(n13657));
  jxor g13543(.dina(n13657), .dinb(n64), .dout(n13658));
  jxor g13544(.dina(n13653), .dinb(n13648), .dout(n13659));
  jand g13545(.dina(n13659), .dinb(n13658), .dout(n13660));
  jor  g13546(.dina(n13660), .dinb(n13654), .dout(n13661));
  jand g13547(.dina(n13661), .dinb(n13229), .dout(n13662));
  jxor g13548(.dina(n13661), .dinb(n13229), .dout(n13663));
  jxor g13549(.dina(n12056), .dinb(n12055), .dout(n13664));
  jand g13550(.dina(n13664), .dinb(n732), .dout(n13665));
  jand g13551(.dina(n11972), .dinb(n3855), .dout(n13666));
  jand g13552(.dina(n11976), .dinb(n3851), .dout(n13667));
  jand g13553(.dina(n11974), .dinb(n3858), .dout(n13668));
  jor  g13554(.dina(n13668), .dinb(n13667), .dout(n13669));
  jor  g13555(.dina(n13669), .dinb(n13666), .dout(n13670));
  jor  g13556(.dina(n13670), .dinb(n13665), .dout(n13671));
  jand g13557(.dina(n13671), .dinb(n13663), .dout(n13672));
  jor  g13558(.dina(n13672), .dinb(n13662), .dout(n13673));
  jxor g13559(.dina(n13610), .dinb(n13595), .dout(n13674));
  jand g13560(.dina(n13674), .dinb(n13673), .dout(n13675));
  jnot g13561(.din(n13675), .dout(n13676));
  jand g13562(.dina(n13676), .dinb(n13611), .dout(n13677));
  jnot g13563(.din(n13677), .dout(n13678));
  jxor g13564(.dina(n13262), .dinb(n13261), .dout(n13679));
  jand g13565(.dina(n13679), .dinb(n13678), .dout(n13680));
  jxor g13566(.dina(n13679), .dinb(n13678), .dout(n13681));
  jxor g13567(.dina(n12062), .dinb(n12061), .dout(n13682));
  jand g13568(.dina(n13682), .dinb(n732), .dout(n13683));
  jand g13569(.dina(n11968), .dinb(n3855), .dout(n13684));
  jand g13570(.dina(n11970), .dinb(n3858), .dout(n13685));
  jand g13571(.dina(n11972), .dinb(n3851), .dout(n13686));
  jor  g13572(.dina(n13686), .dinb(n13685), .dout(n13687));
  jor  g13573(.dina(n13687), .dinb(n13684), .dout(n13688));
  jor  g13574(.dina(n13688), .dinb(n13683), .dout(n13689));
  jand g13575(.dina(n13689), .dinb(n13681), .dout(n13690));
  jor  g13576(.dina(n13690), .dinb(n13680), .dout(n13691));
  jxor g13577(.dina(n13275), .dinb(n13267), .dout(n13692));
  jand g13578(.dina(n13692), .dinb(n13691), .dout(n13693));
  jnot g13579(.din(n13693), .dout(n13694));
  jxor g13580(.dina(n13692), .dinb(n13691), .dout(n13695));
  jnot g13581(.din(n13695), .dout(n13696));
  jand g13582(.dina(n13116), .dinb(n4449), .dout(n13697));
  jand g13583(.dina(n11960), .dinb(n4453), .dout(n13698));
  jand g13584(.dina(n11962), .dinb(n4457), .dout(n13699));
  jand g13585(.dina(n11964), .dinb(n4461), .dout(n13700));
  jor  g13586(.dina(n13700), .dinb(n13699), .dout(n13701));
  jor  g13587(.dina(n13701), .dinb(n13698), .dout(n13702));
  jor  g13588(.dina(n13702), .dinb(n13697), .dout(n13703));
  jxor g13589(.dina(n13703), .dinb(n88), .dout(n13704));
  jor  g13590(.dina(n13704), .dinb(n13696), .dout(n13705));
  jand g13591(.dina(n13705), .dinb(n13694), .dout(n13706));
  jnot g13592(.din(n13706), .dout(n13707));
  jxor g13593(.dina(n13488), .dinb(n13487), .dout(n13708));
  jand g13594(.dina(n13708), .dinb(n13707), .dout(n13709));
  jnot g13595(.din(n13709), .dout(n13710));
  jxor g13596(.dina(n13708), .dinb(n13707), .dout(n13711));
  jnot g13597(.din(n13711), .dout(n13712));
  jand g13598(.dina(n12510), .dinb(n75), .dout(n13713));
  jand g13599(.dina(n11952), .dinb(n4933), .dout(n13714));
  jand g13600(.dina(n11954), .dinb(n4918), .dout(n13715));
  jand g13601(.dina(n11956), .dinb(n4745), .dout(n13716));
  jor  g13602(.dina(n13716), .dinb(n13715), .dout(n13717));
  jor  g13603(.dina(n13717), .dinb(n13714), .dout(n13718));
  jor  g13604(.dina(n13718), .dinb(n13713), .dout(n13719));
  jxor g13605(.dina(n13719), .dinb(n68), .dout(n13720));
  jor  g13606(.dina(n13720), .dinb(n13712), .dout(n13721));
  jand g13607(.dina(n13721), .dinb(n13710), .dout(n13722));
  jnot g13608(.din(n13722), .dout(n13723));
  jxor g13609(.dina(n13593), .dinb(n13592), .dout(n13724));
  jand g13610(.dina(n13724), .dinb(n13723), .dout(n13725));
  jor  g13611(.dina(n13725), .dinb(n13594), .dout(n13726));
  jxor g13612(.dina(n13517), .dinb(n13509), .dout(n13727));
  jand g13613(.dina(n13727), .dinb(n13726), .dout(n13728));
  jnot g13614(.din(n13728), .dout(n13729));
  jxor g13615(.dina(n13727), .dinb(n13726), .dout(n13730));
  jnot g13616(.din(n13730), .dout(n13731));
  jand g13617(.dina(n12751), .dinb(n5365), .dout(n13732));
  jand g13618(.dina(n11942), .dinb(n5500), .dout(n13733));
  jand g13619(.dina(n11944), .dinb(n5424), .dout(n13734));
  jand g13620(.dina(n11946), .dinb(n5363), .dout(n13735));
  jor  g13621(.dina(n13735), .dinb(n13734), .dout(n13736));
  jor  g13622(.dina(n13736), .dinb(n13733), .dout(n13737));
  jor  g13623(.dina(n13737), .dinb(n13732), .dout(n13738));
  jxor g13624(.dina(n13738), .dinb(n72), .dout(n13739));
  jor  g13625(.dina(n13739), .dinb(n13731), .dout(n13740));
  jand g13626(.dina(n13740), .dinb(n13729), .dout(n13741));
  jnot g13627(.din(n13741), .dout(n13742));
  jxor g13628(.dina(n13533), .dinb(n13525), .dout(n13743));
  jand g13629(.dina(n13743), .dinb(n13742), .dout(n13744));
  jnot g13630(.din(n13744), .dout(n13745));
  jxor g13631(.dina(n13743), .dinb(n13742), .dout(n13746));
  jnot g13632(.din(n13746), .dout(n13747));
  jand g13633(.dina(n12841), .dinb(n5693), .dout(n13748));
  jand g13634(.dina(n12783), .dinb(n6209), .dout(n13749));
  jand g13635(.dina(n12766), .dinb(n6131), .dout(n13750));
  jand g13636(.dina(n12177), .dinb(n5691), .dout(n13751));
  jor  g13637(.dina(n13751), .dinb(n13750), .dout(n13752));
  jor  g13638(.dina(n13752), .dinb(n13749), .dout(n13753));
  jor  g13639(.dina(n13753), .dinb(n13748), .dout(n13754));
  jxor g13640(.dina(n13754), .dinb(n4247), .dout(n13755));
  jor  g13641(.dina(n13755), .dinb(n13747), .dout(n13756));
  jand g13642(.dina(n13756), .dinb(n13745), .dout(n13757));
  jnot g13643(.din(n13757), .dout(n13758));
  jxor g13644(.dina(n13582), .dinb(n13574), .dout(n13759));
  jand g13645(.dina(n13759), .dinb(n13758), .dout(n13760));
  jnot g13646(.din(n13760), .dout(n13761));
  jand g13647(.dina(n13761), .dinb(n13583), .dout(n13762));
  jnot g13648(.din(n13762), .dout(n13763));
  jxor g13649(.dina(n13554), .dinb(n13546), .dout(n13764));
  jand g13650(.dina(n13764), .dinb(n13763), .dout(n13765));
  jnot g13651(.din(n13765), .dout(n13766));
  jxor g13652(.dina(n13764), .dinb(n13763), .dout(n13767));
  jnot g13653(.din(n13767), .dout(n13768));
  jor  g13654(.dina(n13354), .dinb(n6341), .dout(n13769));
  jor  g13655(.dina(n12814), .dinb(n6339), .dout(n13770));
  jand g13656(.dina(n12809), .dinb(n6797), .dout(n13771));
  jor  g13657(.dina(n13559), .dinb(n12460), .dout(n13772));
  jor  g13658(.dina(n13772), .dinb(n13771), .dout(n13773));
  jand g13659(.dina(n13773), .dinb(n13770), .dout(n13774));
  jand g13660(.dina(n13774), .dinb(n13769), .dout(n13775));
  jxor g13661(.dina(n13775), .dinb(\a[17] ), .dout(n13776));
  jor  g13662(.dina(n13776), .dinb(n13768), .dout(n13777));
  jand g13663(.dina(n13777), .dinb(n13766), .dout(n13778));
  jnot g13664(.din(n13778), .dout(n13779));
  jxor g13665(.dina(n13566), .dinb(n13565), .dout(n13780));
  jand g13666(.dina(n13780), .dinb(n13779), .dout(n13781));
  jxor g13667(.dina(n13780), .dinb(n13779), .dout(n13782));
  jxor g13668(.dina(n13724), .dinb(n13723), .dout(n13783));
  jnot g13669(.din(n13783), .dout(n13784));
  jand g13670(.dina(n12189), .dinb(n5365), .dout(n13785));
  jand g13671(.dina(n11944), .dinb(n5500), .dout(n13786));
  jand g13672(.dina(n11946), .dinb(n5424), .dout(n13787));
  jand g13673(.dina(n11948), .dinb(n5363), .dout(n13788));
  jor  g13674(.dina(n13788), .dinb(n13787), .dout(n13789));
  jor  g13675(.dina(n13789), .dinb(n13786), .dout(n13790));
  jor  g13676(.dina(n13790), .dinb(n13785), .dout(n13791));
  jxor g13677(.dina(n13791), .dinb(n72), .dout(n13792));
  jor  g13678(.dina(n13792), .dinb(n13784), .dout(n13793));
  jand g13679(.dina(n13134), .dinb(n4449), .dout(n13794));
  jand g13680(.dina(n11962), .dinb(n4453), .dout(n13795));
  jand g13681(.dina(n11964), .dinb(n4457), .dout(n13796));
  jand g13682(.dina(n11966), .dinb(n4461), .dout(n13797));
  jor  g13683(.dina(n13797), .dinb(n13796), .dout(n13798));
  jor  g13684(.dina(n13798), .dinb(n13795), .dout(n13799));
  jor  g13685(.dina(n13799), .dinb(n13794), .dout(n13800));
  jxor g13686(.dina(n13800), .dinb(n88), .dout(n13801));
  jnot g13687(.din(n13801), .dout(n13802));
  jxor g13688(.dina(n13689), .dinb(n13681), .dout(n13803));
  jand g13689(.dina(n13803), .dinb(n13802), .dout(n13804));
  jxor g13690(.dina(n13674), .dinb(n13673), .dout(n13805));
  jxor g13691(.dina(n12059), .dinb(n12058), .dout(n13806));
  jand g13692(.dina(n13806), .dinb(n732), .dout(n13807));
  jand g13693(.dina(n11970), .dinb(n3855), .dout(n13808));
  jand g13694(.dina(n11972), .dinb(n3858), .dout(n13809));
  jand g13695(.dina(n11974), .dinb(n3851), .dout(n13810));
  jor  g13696(.dina(n13810), .dinb(n13809), .dout(n13811));
  jor  g13697(.dina(n13811), .dinb(n13808), .dout(n13812));
  jor  g13698(.dina(n13812), .dinb(n13807), .dout(n13813));
  jand g13699(.dina(n13813), .dinb(n13805), .dout(n13814));
  jand g13700(.dina(n3097), .dinb(n2697), .dout(n13815));
  jand g13701(.dina(n12261), .dinb(n1249), .dout(n13816));
  jand g13702(.dina(n13816), .dinb(n13815), .dout(n13817));
  jand g13703(.dina(n756), .dinb(n202), .dout(n13818));
  jand g13704(.dina(n692), .dinb(n270), .dout(n13819));
  jand g13705(.dina(n13819), .dinb(n13818), .dout(n13820));
  jand g13706(.dina(n418), .dinb(n234), .dout(n13821));
  jand g13707(.dina(n815), .dinb(n243), .dout(n13822));
  jand g13708(.dina(n13822), .dinb(n13821), .dout(n13823));
  jand g13709(.dina(n13823), .dinb(n13820), .dout(n13824));
  jand g13710(.dina(n13824), .dinb(n13817), .dout(n13825));
  jnot g13711(.din(n2073), .dout(n13826));
  jand g13712(.dina(n3536), .dinb(n13826), .dout(n13827));
  jand g13713(.dina(n13827), .dinb(n13825), .dout(n13828));
  jand g13714(.dina(n13828), .dinb(n335), .dout(n13829));
  jand g13715(.dina(n13829), .dinb(n3775), .dout(n13830));
  jand g13716(.dina(n13830), .dinb(n3903), .dout(n13831));
  jor  g13717(.dina(n13831), .dinb(n13653), .dout(n13832));
  jand g13718(.dina(n563), .dinb(n330), .dout(n13833));
  jand g13719(.dina(n13833), .dinb(n12199), .dout(n13834));
  jand g13720(.dina(n2784), .dinb(n647), .dout(n13835));
  jand g13721(.dina(n2538), .dinb(n1424), .dout(n13836));
  jand g13722(.dina(n13836), .dinb(n13835), .dout(n13837));
  jand g13723(.dina(n13837), .dinb(n13834), .dout(n13838));
  jand g13724(.dina(n13838), .dinb(n12424), .dout(n13839));
  jand g13725(.dina(n431), .dinb(n194), .dout(n13840));
  jand g13726(.dina(n641), .dinb(n605), .dout(n13841));
  jand g13727(.dina(n13841), .dinb(n13840), .dout(n13842));
  jand g13728(.dina(n696), .dinb(n483), .dout(n13843));
  jand g13729(.dina(n13843), .dinb(n5003), .dout(n13844));
  jand g13730(.dina(n13844), .dinb(n13842), .dout(n13845));
  jand g13731(.dina(n4401), .dinb(n2770), .dout(n13846));
  jand g13732(.dina(n13846), .dinb(n13845), .dout(n13847));
  jand g13733(.dina(n13847), .dinb(n1540), .dout(n13848));
  jand g13734(.dina(n13848), .dinb(n1650), .dout(n13849));
  jand g13735(.dina(n13849), .dinb(n13839), .dout(n13850));
  jand g13736(.dina(n13850), .dinb(n13635), .dout(n13851));
  jor  g13737(.dina(n13851), .dinb(n13653), .dout(n13852));
  jand g13738(.dina(n5122), .dinb(n3092), .dout(n13853));
  jand g13739(.dina(n13853), .dinb(n2183), .dout(n13854));
  jand g13740(.dina(n435), .dinb(n257), .dout(n13855));
  jand g13741(.dina(n13855), .dinb(n527), .dout(n13856));
  jand g13742(.dina(n7043), .dinb(n1390), .dout(n13857));
  jand g13743(.dina(n13857), .dinb(n13856), .dout(n13858));
  jand g13744(.dina(n5815), .dinb(n4001), .dout(n13859));
  jand g13745(.dina(n13859), .dinb(n13858), .dout(n13860));
  jand g13746(.dina(n13860), .dinb(n13854), .dout(n13861));
  jand g13747(.dina(n1264), .dinb(n715), .dout(n13862));
  jand g13748(.dina(n13862), .dinb(n703), .dout(n13863));
  jand g13749(.dina(n1615), .dinb(n476), .dout(n13864));
  jand g13750(.dina(n13864), .dinb(n2378), .dout(n13865));
  jand g13751(.dina(n13865), .dinb(n3075), .dout(n13866));
  jand g13752(.dina(n13866), .dinb(n13863), .dout(n13867));
  jand g13753(.dina(n13867), .dinb(n2577), .dout(n13868));
  jand g13754(.dina(n13868), .dinb(n13861), .dout(n13869));
  jand g13755(.dina(n439), .dinb(n311), .dout(n13870));
  jand g13756(.dina(n13870), .dinb(n243), .dout(n13871));
  jand g13757(.dina(n2526), .dinb(n2291), .dout(n13872));
  jand g13758(.dina(n13872), .dinb(n13871), .dout(n13873));
  jand g13759(.dina(n13873), .dinb(n13869), .dout(n13874));
  jand g13760(.dina(n876), .dinb(n395), .dout(n13875));
  jand g13761(.dina(n13875), .dinb(n696), .dout(n13876));
  jand g13762(.dina(n511), .dinb(n329), .dout(n13877));
  jand g13763(.dina(n778), .dinb(n367), .dout(n13878));
  jand g13764(.dina(n13878), .dinb(n13877), .dout(n13879));
  jand g13765(.dina(n13879), .dinb(n13876), .dout(n13880));
  jand g13766(.dina(n13880), .dinb(n734), .dout(n13881));
  jand g13767(.dina(n543), .dinb(n450), .dout(n13882));
  jand g13768(.dina(n13882), .dinb(n234), .dout(n13883));
  jand g13769(.dina(n763), .dinb(n687), .dout(n13884));
  jand g13770(.dina(n533), .dinb(n503), .dout(n13885));
  jand g13771(.dina(n13885), .dinb(n13884), .dout(n13886));
  jand g13772(.dina(n13886), .dinb(n13883), .dout(n13887));
  jand g13773(.dina(n13151), .dinb(n186), .dout(n13888));
  jand g13774(.dina(n13888), .dinb(n13887), .dout(n13889));
  jand g13775(.dina(n1470), .dinb(n393), .dout(n13890));
  jand g13776(.dina(n13890), .dinb(n3590), .dout(n13891));
  jand g13777(.dina(n13891), .dinb(n2594), .dout(n13892));
  jand g13778(.dina(n13892), .dinb(n13889), .dout(n13893));
  jand g13779(.dina(n13893), .dinb(n13881), .dout(n13894));
  jand g13780(.dina(n13894), .dinb(n12887), .dout(n13895));
  jand g13781(.dina(n13895), .dinb(n13874), .dout(n13896));
  jor  g13782(.dina(n13896), .dinb(n13653), .dout(n13897));
  jxor g13783(.dina(n13896), .dinb(n13653), .dout(n13898));
  jxor g13784(.dina(n12044), .dinb(n12043), .dout(n13899));
  jand g13785(.dina(n13899), .dinb(n732), .dout(n13900));
  jand g13786(.dina(n11980), .dinb(n3855), .dout(n13901));
  jand g13787(.dina(n11982), .dinb(n3858), .dout(n13902));
  jand g13788(.dina(n11985), .dinb(n3851), .dout(n13903));
  jor  g13789(.dina(n13903), .dinb(n13902), .dout(n13904));
  jor  g13790(.dina(n13904), .dinb(n13901), .dout(n13905));
  jor  g13791(.dina(n13905), .dinb(n13900), .dout(n13906));
  jand g13792(.dina(n13906), .dinb(n13898), .dout(n13907));
  jnot g13793(.din(n13907), .dout(n13908));
  jand g13794(.dina(n13908), .dinb(n13897), .dout(n13909));
  jnot g13795(.din(n13909), .dout(n13910));
  jxor g13796(.dina(n13851), .dinb(n13653), .dout(n13911));
  jand g13797(.dina(n13911), .dinb(n13910), .dout(n13912));
  jnot g13798(.din(n13912), .dout(n13913));
  jand g13799(.dina(n13913), .dinb(n13852), .dout(n13914));
  jnot g13800(.din(n13914), .dout(n13915));
  jxor g13801(.dina(n13831), .dinb(n13653), .dout(n13916));
  jand g13802(.dina(n13916), .dinb(n13915), .dout(n13917));
  jnot g13803(.din(n13917), .dout(n13918));
  jand g13804(.dina(n13918), .dinb(n13832), .dout(n13919));
  jnot g13805(.din(n13919), .dout(n13920));
  jxor g13806(.dina(n13659), .dinb(n13658), .dout(n13921));
  jand g13807(.dina(n13921), .dinb(n13920), .dout(n13922));
  jxor g13808(.dina(n13921), .dinb(n13920), .dout(n13923));
  jxor g13809(.dina(n12053), .dinb(n12052), .dout(n13924));
  jand g13810(.dina(n13924), .dinb(n732), .dout(n13925));
  jand g13811(.dina(n11974), .dinb(n3855), .dout(n13926));
  jand g13812(.dina(n11976), .dinb(n3858), .dout(n13927));
  jand g13813(.dina(n11978), .dinb(n3851), .dout(n13928));
  jor  g13814(.dina(n13928), .dinb(n13927), .dout(n13929));
  jor  g13815(.dina(n13929), .dinb(n13926), .dout(n13930));
  jor  g13816(.dina(n13930), .dinb(n13925), .dout(n13931));
  jand g13817(.dina(n13931), .dinb(n13923), .dout(n13932));
  jor  g13818(.dina(n13932), .dinb(n13922), .dout(n13933));
  jxor g13819(.dina(n13671), .dinb(n13663), .dout(n13934));
  jand g13820(.dina(n13934), .dinb(n13933), .dout(n13935));
  jnot g13821(.din(n13935), .dout(n13936));
  jxor g13822(.dina(n13934), .dinb(n13933), .dout(n13937));
  jnot g13823(.din(n13937), .dout(n13938));
  jand g13824(.dina(n13268), .dinb(n4449), .dout(n13939));
  jand g13825(.dina(n11966), .dinb(n4453), .dout(n13940));
  jand g13826(.dina(n11968), .dinb(n4457), .dout(n13941));
  jand g13827(.dina(n11970), .dinb(n4461), .dout(n13942));
  jor  g13828(.dina(n13942), .dinb(n13941), .dout(n13943));
  jor  g13829(.dina(n13943), .dinb(n13940), .dout(n13944));
  jor  g13830(.dina(n13944), .dinb(n13939), .dout(n13945));
  jxor g13831(.dina(n13945), .dinb(n88), .dout(n13946));
  jor  g13832(.dina(n13946), .dinb(n13938), .dout(n13947));
  jand g13833(.dina(n13947), .dinb(n13936), .dout(n13948));
  jnot g13834(.din(n13948), .dout(n13949));
  jxor g13835(.dina(n13813), .dinb(n13805), .dout(n13950));
  jand g13836(.dina(n13950), .dinb(n13949), .dout(n13951));
  jor  g13837(.dina(n13951), .dinb(n13814), .dout(n13952));
  jxor g13838(.dina(n13803), .dinb(n13802), .dout(n13953));
  jand g13839(.dina(n13953), .dinb(n13952), .dout(n13954));
  jor  g13840(.dina(n13954), .dinb(n13804), .dout(n13955));
  jxor g13841(.dina(n13704), .dinb(n13696), .dout(n13956));
  jand g13842(.dina(n13956), .dinb(n13955), .dout(n13957));
  jnot g13843(.din(n13957), .dout(n13958));
  jxor g13844(.dina(n13956), .dinb(n13955), .dout(n13959));
  jnot g13845(.din(n13959), .dout(n13960));
  jand g13846(.dina(n12472), .dinb(n75), .dout(n13961));
  jand g13847(.dina(n11954), .dinb(n4933), .dout(n13962));
  jand g13848(.dina(n11956), .dinb(n4918), .dout(n13963));
  jand g13849(.dina(n11958), .dinb(n4745), .dout(n13964));
  jor  g13850(.dina(n13964), .dinb(n13963), .dout(n13965));
  jor  g13851(.dina(n13965), .dinb(n13962), .dout(n13966));
  jor  g13852(.dina(n13966), .dinb(n13961), .dout(n13967));
  jxor g13853(.dina(n13967), .dinb(n68), .dout(n13968));
  jor  g13854(.dina(n13968), .dinb(n13960), .dout(n13969));
  jand g13855(.dina(n13969), .dinb(n13958), .dout(n13970));
  jnot g13856(.din(n13970), .dout(n13971));
  jxor g13857(.dina(n13720), .dinb(n13712), .dout(n13972));
  jand g13858(.dina(n13972), .dinb(n13971), .dout(n13973));
  jnot g13859(.din(n13973), .dout(n13974));
  jxor g13860(.dina(n13972), .dinb(n13971), .dout(n13975));
  jnot g13861(.din(n13975), .dout(n13976));
  jand g13862(.dina(n12519), .dinb(n5365), .dout(n13977));
  jand g13863(.dina(n11946), .dinb(n5500), .dout(n13978));
  jand g13864(.dina(n11948), .dinb(n5424), .dout(n13979));
  jand g13865(.dina(n11950), .dinb(n5363), .dout(n13980));
  jor  g13866(.dina(n13980), .dinb(n13979), .dout(n13981));
  jor  g13867(.dina(n13981), .dinb(n13978), .dout(n13982));
  jor  g13868(.dina(n13982), .dinb(n13977), .dout(n13983));
  jxor g13869(.dina(n13983), .dinb(n72), .dout(n13984));
  jor  g13870(.dina(n13984), .dinb(n13976), .dout(n13985));
  jand g13871(.dina(n13985), .dinb(n13974), .dout(n13986));
  jnot g13872(.din(n13986), .dout(n13987));
  jxor g13873(.dina(n13792), .dinb(n13784), .dout(n13988));
  jand g13874(.dina(n13988), .dinb(n13987), .dout(n13989));
  jnot g13875(.din(n13989), .dout(n13990));
  jand g13876(.dina(n13990), .dinb(n13793), .dout(n13991));
  jnot g13877(.din(n13991), .dout(n13992));
  jxor g13878(.dina(n13739), .dinb(n13731), .dout(n13993));
  jand g13879(.dina(n13993), .dinb(n13992), .dout(n13994));
  jnot g13880(.din(n13994), .dout(n13995));
  jxor g13881(.dina(n13993), .dinb(n13992), .dout(n13996));
  jnot g13882(.din(n13996), .dout(n13997));
  jand g13883(.dina(n12768), .dinb(n5693), .dout(n13998));
  jand g13884(.dina(n12766), .dinb(n6209), .dout(n13999));
  jand g13885(.dina(n12177), .dinb(n6131), .dout(n14000));
  jand g13886(.dina(n11941), .dinb(n5691), .dout(n14001));
  jor  g13887(.dina(n14001), .dinb(n14000), .dout(n14002));
  jor  g13888(.dina(n14002), .dinb(n13999), .dout(n14003));
  jor  g13889(.dina(n14003), .dinb(n13998), .dout(n14004));
  jxor g13890(.dina(n14004), .dinb(n4247), .dout(n14005));
  jor  g13891(.dina(n14005), .dinb(n13997), .dout(n14006));
  jand g13892(.dina(n14006), .dinb(n13995), .dout(n14007));
  jnot g13893(.din(n14007), .dout(n14008));
  jxor g13894(.dina(n13755), .dinb(n13747), .dout(n14009));
  jand g13895(.dina(n14009), .dinb(n14008), .dout(n14010));
  jnot g13896(.din(n14010), .dout(n14011));
  jxor g13897(.dina(n14009), .dinb(n14008), .dout(n14012));
  jnot g13898(.din(n14012), .dout(n14013));
  jand g13899(.dina(n12919), .dinb(n6340), .dout(n14014));
  jand g13900(.dina(n12815), .dinb(n6798), .dout(n14015));
  jand g13901(.dina(n12795), .dinb(n6556), .dout(n14016));
  jand g13902(.dina(n12782), .dinb(n6338), .dout(n14017));
  jor  g13903(.dina(n14017), .dinb(n14016), .dout(n14018));
  jor  g13904(.dina(n14018), .dinb(n14015), .dout(n14019));
  jor  g13905(.dina(n14019), .dinb(n14014), .dout(n14020));
  jxor g13906(.dina(n14020), .dinb(n5064), .dout(n14021));
  jor  g13907(.dina(n14021), .dinb(n14013), .dout(n14022));
  jand g13908(.dina(n14022), .dinb(n14011), .dout(n14023));
  jand g13909(.dina(n13022), .dinb(n6340), .dout(n14024));
  jand g13910(.dina(n12815), .dinb(n6556), .dout(n14026));
  jand g13911(.dina(n12795), .dinb(n6338), .dout(n14027));
  jor  g13912(.dina(n14027), .dinb(n14026), .dout(n14028));
  jor  g13913(.dina(n14028), .dinb(n6798), .dout(n14029));
  jor  g13914(.dina(n14029), .dinb(n14024), .dout(n14030));
  jxor g13915(.dina(n14030), .dinb(n5064), .dout(n14031));
  jor  g13916(.dina(n14031), .dinb(n14023), .dout(n14032));
  jxor g13917(.dina(n13759), .dinb(n13758), .dout(n14033));
  jxor g13918(.dina(n14031), .dinb(n14023), .dout(n14034));
  jand g13919(.dina(n14034), .dinb(n14033), .dout(n14035));
  jnot g13920(.din(n14035), .dout(n14036));
  jand g13921(.dina(n14036), .dinb(n14032), .dout(n14037));
  jnot g13922(.din(n14037), .dout(n14038));
  jxor g13923(.dina(n13776), .dinb(n13768), .dout(n14039));
  jand g13924(.dina(n14039), .dinb(n14038), .dout(n14040));
  jxor g13925(.dina(n13988), .dinb(n13987), .dout(n14041));
  jnot g13926(.din(n14041), .dout(n14042));
  jand g13927(.dina(n12179), .dinb(n5693), .dout(n14043));
  jand g13928(.dina(n12177), .dinb(n6209), .dout(n14044));
  jand g13929(.dina(n11941), .dinb(n6131), .dout(n14045));
  jand g13930(.dina(n11942), .dinb(n5691), .dout(n14046));
  jor  g13931(.dina(n14046), .dinb(n14045), .dout(n14047));
  jor  g13932(.dina(n14047), .dinb(n14044), .dout(n14048));
  jor  g13933(.dina(n14048), .dinb(n14043), .dout(n14049));
  jxor g13934(.dina(n14049), .dinb(n4247), .dout(n14050));
  jor  g13935(.dina(n14050), .dinb(n14042), .dout(n14051));
  jxor g13936(.dina(n13953), .dinb(n13952), .dout(n14052));
  jnot g13937(.din(n14052), .dout(n14053));
  jand g13938(.dina(n12639), .dinb(n75), .dout(n14054));
  jand g13939(.dina(n11956), .dinb(n4933), .dout(n14055));
  jand g13940(.dina(n11958), .dinb(n4918), .dout(n14056));
  jand g13941(.dina(n11960), .dinb(n4745), .dout(n14057));
  jor  g13942(.dina(n14057), .dinb(n14056), .dout(n14058));
  jor  g13943(.dina(n14058), .dinb(n14055), .dout(n14059));
  jor  g13944(.dina(n14059), .dinb(n14054), .dout(n14060));
  jxor g13945(.dina(n14060), .dinb(n68), .dout(n14061));
  jor  g13946(.dina(n14061), .dinb(n14053), .dout(n14062));
  jxor g13947(.dina(n13950), .dinb(n13949), .dout(n14063));
  jnot g13948(.din(n14063), .dout(n14064));
  jand g13949(.dina(n13470), .dinb(n4449), .dout(n14065));
  jand g13950(.dina(n11964), .dinb(n4453), .dout(n14066));
  jand g13951(.dina(n11966), .dinb(n4457), .dout(n14067));
  jand g13952(.dina(n11968), .dinb(n4461), .dout(n14068));
  jor  g13953(.dina(n14068), .dinb(n14067), .dout(n14069));
  jor  g13954(.dina(n14069), .dinb(n14066), .dout(n14070));
  jor  g13955(.dina(n14070), .dinb(n14065), .dout(n14071));
  jxor g13956(.dina(n14071), .dinb(n88), .dout(n14072));
  jor  g13957(.dina(n14072), .dinb(n14064), .dout(n14073));
  jand g13958(.dina(n12624), .dinb(n75), .dout(n14074));
  jand g13959(.dina(n11958), .dinb(n4933), .dout(n14075));
  jand g13960(.dina(n11960), .dinb(n4918), .dout(n14076));
  jand g13961(.dina(n11962), .dinb(n4745), .dout(n14077));
  jor  g13962(.dina(n14077), .dinb(n14076), .dout(n14078));
  jor  g13963(.dina(n14078), .dinb(n14075), .dout(n14079));
  jor  g13964(.dina(n14079), .dinb(n14074), .dout(n14080));
  jxor g13965(.dina(n14080), .dinb(n68), .dout(n14081));
  jnot g13966(.din(n14081), .dout(n14082));
  jxor g13967(.dina(n14072), .dinb(n14064), .dout(n14083));
  jand g13968(.dina(n14083), .dinb(n14082), .dout(n14084));
  jnot g13969(.din(n14084), .dout(n14085));
  jand g13970(.dina(n14085), .dinb(n14073), .dout(n14086));
  jnot g13971(.din(n14086), .dout(n14087));
  jxor g13972(.dina(n14061), .dinb(n14053), .dout(n14088));
  jand g13973(.dina(n14088), .dinb(n14087), .dout(n14089));
  jnot g13974(.din(n14089), .dout(n14090));
  jand g13975(.dina(n14090), .dinb(n14062), .dout(n14091));
  jnot g13976(.din(n14091), .dout(n14092));
  jxor g13977(.dina(n13968), .dinb(n13960), .dout(n14093));
  jand g13978(.dina(n14093), .dinb(n14092), .dout(n14094));
  jnot g13979(.din(n14094), .dout(n14095));
  jxor g13980(.dina(n14093), .dinb(n14092), .dout(n14096));
  jnot g13981(.din(n14096), .dout(n14097));
  jand g13982(.dina(n12654), .dinb(n5365), .dout(n14098));
  jand g13983(.dina(n11948), .dinb(n5500), .dout(n14099));
  jand g13984(.dina(n11950), .dinb(n5424), .dout(n14100));
  jand g13985(.dina(n11952), .dinb(n5363), .dout(n14101));
  jor  g13986(.dina(n14101), .dinb(n14100), .dout(n14102));
  jor  g13987(.dina(n14102), .dinb(n14099), .dout(n14103));
  jor  g13988(.dina(n14103), .dinb(n14098), .dout(n14104));
  jxor g13989(.dina(n14104), .dinb(n72), .dout(n14105));
  jor  g13990(.dina(n14105), .dinb(n14097), .dout(n14106));
  jand g13991(.dina(n14106), .dinb(n14095), .dout(n14107));
  jnot g13992(.din(n14107), .dout(n14108));
  jxor g13993(.dina(n13984), .dinb(n13976), .dout(n14109));
  jand g13994(.dina(n14109), .dinb(n14108), .dout(n14110));
  jnot g13995(.din(n14110), .dout(n14111));
  jxor g13996(.dina(n14109), .dinb(n14108), .dout(n14112));
  jnot g13997(.din(n14112), .dout(n14113));
  jand g13998(.dina(n12671), .dinb(n5693), .dout(n14114));
  jand g13999(.dina(n11941), .dinb(n6209), .dout(n14115));
  jand g14000(.dina(n11942), .dinb(n6131), .dout(n14116));
  jand g14001(.dina(n11944), .dinb(n5691), .dout(n14117));
  jor  g14002(.dina(n14117), .dinb(n14116), .dout(n14118));
  jor  g14003(.dina(n14118), .dinb(n14115), .dout(n14119));
  jor  g14004(.dina(n14119), .dinb(n14114), .dout(n14120));
  jxor g14005(.dina(n14120), .dinb(n4247), .dout(n14121));
  jor  g14006(.dina(n14121), .dinb(n14113), .dout(n14122));
  jand g14007(.dina(n14122), .dinb(n14111), .dout(n14123));
  jnot g14008(.din(n14123), .dout(n14124));
  jxor g14009(.dina(n14050), .dinb(n14042), .dout(n14125));
  jand g14010(.dina(n14125), .dinb(n14124), .dout(n14126));
  jnot g14011(.din(n14126), .dout(n14127));
  jand g14012(.dina(n14127), .dinb(n14051), .dout(n14128));
  jnot g14013(.din(n14128), .dout(n14129));
  jxor g14014(.dina(n14005), .dinb(n13997), .dout(n14130));
  jand g14015(.dina(n14130), .dinb(n14129), .dout(n14131));
  jnot g14016(.din(n14131), .dout(n14132));
  jxor g14017(.dina(n14130), .dinb(n14129), .dout(n14133));
  jnot g14018(.din(n14133), .dout(n14134));
  jand g14019(.dina(n12797), .dinb(n6340), .dout(n14135));
  jand g14020(.dina(n12795), .dinb(n6798), .dout(n14136));
  jand g14021(.dina(n12782), .dinb(n6556), .dout(n14137));
  jand g14022(.dina(n12783), .dinb(n6338), .dout(n14138));
  jor  g14023(.dina(n14138), .dinb(n14137), .dout(n14139));
  jor  g14024(.dina(n14139), .dinb(n14136), .dout(n14140));
  jor  g14025(.dina(n14140), .dinb(n14135), .dout(n14141));
  jxor g14026(.dina(n14141), .dinb(n5064), .dout(n14142));
  jor  g14027(.dina(n14142), .dinb(n14134), .dout(n14143));
  jand g14028(.dina(n14143), .dinb(n14132), .dout(n14144));
  jand g14029(.dina(n7740), .dinb(n7614), .dout(n14147));
  jor  g14030(.dina(n12465), .dinb(n14144), .dout(n14152));
  jxor g14031(.dina(n12465), .dinb(n14144), .dout(n14153));
  jxor g14032(.dina(n14021), .dinb(n14013), .dout(n14154));
  jand g14033(.dina(n14154), .dinb(n14153), .dout(n14155));
  jnot g14034(.din(n14155), .dout(n14156));
  jand g14035(.dina(n14156), .dinb(n14152), .dout(n14157));
  jnot g14036(.din(n14157), .dout(n14158));
  jxor g14037(.dina(n14034), .dinb(n14033), .dout(n14159));
  jand g14038(.dina(n14159), .dinb(n14158), .dout(n14160));
  jxor g14039(.dina(n14125), .dinb(n14124), .dout(n14161));
  jnot g14040(.din(n14161), .dout(n14162));
  jand g14041(.dina(n12938), .dinb(n6340), .dout(n14163));
  jand g14042(.dina(n12782), .dinb(n6798), .dout(n14164));
  jand g14043(.dina(n12783), .dinb(n6556), .dout(n14165));
  jand g14044(.dina(n12766), .dinb(n6338), .dout(n14166));
  jor  g14045(.dina(n14166), .dinb(n14165), .dout(n14167));
  jor  g14046(.dina(n14167), .dinb(n14164), .dout(n14168));
  jor  g14047(.dina(n14168), .dinb(n14163), .dout(n14169));
  jxor g14048(.dina(n14169), .dinb(n5064), .dout(n14170));
  jor  g14049(.dina(n14170), .dinb(n14162), .dout(n14171));
  jxor g14050(.dina(n14088), .dinb(n14087), .dout(n14172));
  jnot g14051(.din(n14172), .dout(n14173));
  jand g14052(.dina(n12569), .dinb(n5365), .dout(n14174));
  jand g14053(.dina(n11950), .dinb(n5500), .dout(n14175));
  jand g14054(.dina(n11952), .dinb(n5424), .dout(n14176));
  jand g14055(.dina(n11954), .dinb(n5363), .dout(n14177));
  jor  g14056(.dina(n14177), .dinb(n14176), .dout(n14178));
  jor  g14057(.dina(n14178), .dinb(n14175), .dout(n14179));
  jor  g14058(.dina(n14179), .dinb(n14174), .dout(n14180));
  jxor g14059(.dina(n14180), .dinb(n72), .dout(n14181));
  jor  g14060(.dina(n14181), .dinb(n14173), .dout(n14182));
  jxor g14061(.dina(n13916), .dinb(n13915), .dout(n14183));
  jxor g14062(.dina(n12050), .dinb(n12049), .dout(n14184));
  jand g14063(.dina(n14184), .dinb(n732), .dout(n14185));
  jand g14064(.dina(n11976), .dinb(n3855), .dout(n14186));
  jand g14065(.dina(n11978), .dinb(n3858), .dout(n14187));
  jand g14066(.dina(n11980), .dinb(n3851), .dout(n14188));
  jor  g14067(.dina(n14188), .dinb(n14187), .dout(n14189));
  jor  g14068(.dina(n14189), .dinb(n14186), .dout(n14190));
  jor  g14069(.dina(n14190), .dinb(n14185), .dout(n14191));
  jand g14070(.dina(n14191), .dinb(n14183), .dout(n14192));
  jxor g14071(.dina(n13911), .dinb(n13910), .dout(n14193));
  jxor g14072(.dina(n12047), .dinb(n12046), .dout(n14194));
  jand g14073(.dina(n14194), .dinb(n732), .dout(n14195));
  jand g14074(.dina(n11978), .dinb(n3855), .dout(n14196));
  jand g14075(.dina(n11980), .dinb(n3858), .dout(n14197));
  jand g14076(.dina(n11982), .dinb(n3851), .dout(n14198));
  jor  g14077(.dina(n14198), .dinb(n14197), .dout(n14199));
  jor  g14078(.dina(n14199), .dinb(n14196), .dout(n14200));
  jor  g14079(.dina(n14200), .dinb(n14195), .dout(n14201));
  jand g14080(.dina(n14201), .dinb(n14193), .dout(n14202));
  jand g14081(.dina(n1285), .dinb(n1150), .dout(n14203));
  jand g14082(.dina(n3595), .dinb(n1242), .dout(n14204));
  jand g14083(.dina(n14204), .dinb(n14203), .dout(n14205));
  jand g14084(.dina(n14205), .dinb(n13060), .dout(n14206));
  jand g14085(.dina(n14206), .dinb(n3063), .dout(n14207));
  jand g14086(.dina(n751), .dinb(n230), .dout(n14208));
  jand g14087(.dina(n14208), .dinb(n721), .dout(n14209));
  jand g14088(.dina(n14209), .dinb(n2361), .dout(n14210));
  jand g14089(.dina(n14210), .dinb(n705), .dout(n14211));
  jand g14090(.dina(n288), .dinb(n174), .dout(n14212));
  jand g14091(.dina(n14212), .dinb(n190), .dout(n14213));
  jand g14092(.dina(n14213), .dinb(n507), .dout(n14214));
  jand g14093(.dina(n4166), .dinb(n3528), .dout(n14215));
  jand g14094(.dina(n14215), .dinb(n14214), .dout(n14216));
  jand g14095(.dina(n14216), .dinb(n14211), .dout(n14217));
  jand g14096(.dina(n14217), .dinb(n14207), .dout(n14218));
  jand g14097(.dina(n14218), .dinb(n1590), .dout(n14219));
  jand g14098(.dina(n14219), .dinb(n5584), .dout(n14220));
  jxor g14099(.dina(n12041), .dinb(n12039), .dout(n14221));
  jor  g14100(.dina(n14221), .dinb(n6463), .dout(n14222));
  jand g14101(.dina(n11982), .dinb(n3855), .dout(n14223));
  jand g14102(.dina(n11988), .dinb(n3851), .dout(n14224));
  jand g14103(.dina(n11985), .dinb(n3858), .dout(n14225));
  jor  g14104(.dina(n14225), .dinb(n14224), .dout(n14226));
  jor  g14105(.dina(n14226), .dinb(n14223), .dout(n14227));
  jnot g14106(.din(n14227), .dout(n14228));
  jand g14107(.dina(n14228), .dinb(n14222), .dout(n14229));
  jor  g14108(.dina(n14229), .dinb(n14220), .dout(n14230));
  jand g14109(.dina(n643), .dinb(n280), .dout(n14231));
  jand g14110(.dina(n418), .dinb(n304), .dout(n14232));
  jand g14111(.dina(n14232), .dinb(n14231), .dout(n14233));
  jand g14112(.dina(n739), .dinb(n352), .dout(n14234));
  jand g14113(.dina(n14234), .dinb(n1295), .dout(n14235));
  jand g14114(.dina(n3594), .dinb(n1410), .dout(n14236));
  jand g14115(.dina(n14236), .dinb(n14235), .dout(n14237));
  jand g14116(.dina(n14237), .dinb(n14233), .dout(n14238));
  jnot g14117(.din(n3214), .dout(n14239));
  jand g14118(.dina(n4084), .dinb(n3644), .dout(n14240));
  jand g14119(.dina(n14240), .dinb(n2026), .dout(n14241));
  jand g14120(.dina(n14241), .dinb(n14239), .dout(n14242));
  jand g14121(.dina(n14242), .dinb(n14238), .dout(n14243));
  jand g14122(.dina(n6614), .dinb(n4715), .dout(n14244));
  jand g14123(.dina(n14244), .dinb(n14243), .dout(n14245));
  jand g14124(.dina(n14245), .dinb(n1921), .dout(n14246));
  jand g14125(.dina(n14246), .dinb(n1517), .dout(n14247));
  jxor g14126(.dina(n12036), .dinb(n12035), .dout(n14248));
  jor  g14127(.dina(n14248), .dinb(n6463), .dout(n14249));
  jand g14128(.dina(n11985), .dinb(n3855), .dout(n14250));
  jand g14129(.dina(n11992), .dinb(n3851), .dout(n14251));
  jand g14130(.dina(n11988), .dinb(n3858), .dout(n14252));
  jor  g14131(.dina(n14252), .dinb(n14251), .dout(n14253));
  jor  g14132(.dina(n14253), .dinb(n14250), .dout(n14254));
  jnot g14133(.din(n14254), .dout(n14255));
  jand g14134(.dina(n14255), .dinb(n14249), .dout(n14256));
  jor  g14135(.dina(n14256), .dinb(n14247), .dout(n14257));
  jand g14136(.dina(n5166), .dinb(n3439), .dout(n14258));
  jand g14137(.dina(n14258), .dinb(n2383), .dout(n14259));
  jand g14138(.dina(n13619), .dinb(n1847), .dout(n14260));
  jand g14139(.dina(n2413), .dinb(n1924), .dout(n14261));
  jand g14140(.dina(n14261), .dinb(n14260), .dout(n14262));
  jand g14141(.dina(n770), .dinb(n331), .dout(n14263));
  jand g14142(.dina(n14263), .dinb(n413), .dout(n14264));
  jand g14143(.dina(n14264), .dinb(n4383), .dout(n14265));
  jand g14144(.dina(n14265), .dinb(n14262), .dout(n14266));
  jand g14145(.dina(n14266), .dinb(n14259), .dout(n14267));
  jand g14146(.dina(n14267), .dinb(n3380), .dout(n14268));
  jand g14147(.dina(n14268), .dinb(n2571), .dout(n14269));
  jand g14148(.dina(n14269), .dinb(n13874), .dout(n14270));
  jxor g14149(.dina(n12032), .dinb(n12031), .dout(n14271));
  jor  g14150(.dina(n14271), .dinb(n6463), .dout(n14272));
  jand g14151(.dina(n11988), .dinb(n3855), .dout(n14273));
  jnot g14152(.din(n11995), .dout(n14274));
  jand g14153(.dina(n14274), .dinb(n3851), .dout(n14275));
  jand g14154(.dina(n11992), .dinb(n3858), .dout(n14276));
  jor  g14155(.dina(n14276), .dinb(n14275), .dout(n14277));
  jor  g14156(.dina(n14277), .dinb(n14273), .dout(n14278));
  jnot g14157(.din(n14278), .dout(n14279));
  jand g14158(.dina(n14279), .dinb(n14272), .dout(n14280));
  jor  g14159(.dina(n14280), .dinb(n14270), .dout(n14281));
  jand g14160(.dina(n165), .dinb(n120), .dout(n14282));
  jand g14161(.dina(n843), .dinb(n352), .dout(n14283));
  jand g14162(.dina(n14283), .dinb(n14282), .dout(n14284));
  jand g14163(.dina(n2151), .dinb(n1287), .dout(n14285));
  jand g14164(.dina(n14285), .dinb(n14284), .dout(n14286));
  jand g14165(.dina(n4692), .dinb(n2383), .dout(n14287));
  jand g14166(.dina(n14287), .dinb(n14286), .dout(n14288));
  jand g14167(.dina(n325), .dinb(n205), .dout(n14289));
  jand g14168(.dina(n382), .dinb(n357), .dout(n14290));
  jand g14169(.dina(n14290), .dinb(n14289), .dout(n14291));
  jand g14170(.dina(n1829), .dinb(n647), .dout(n14292));
  jand g14171(.dina(n14292), .dinb(n14291), .dout(n14293));
  jand g14172(.dina(n5212), .dinb(n1197), .dout(n14294));
  jand g14173(.dina(n14294), .dinb(n277), .dout(n14295));
  jand g14174(.dina(n14295), .dinb(n14293), .dout(n14296));
  jand g14175(.dina(n14296), .dinb(n14288), .dout(n14297));
  jand g14176(.dina(n4221), .dinb(n823), .dout(n14298));
  jand g14177(.dina(n14298), .dinb(n14297), .dout(n14299));
  jand g14178(.dina(n14299), .dinb(n3973), .dout(n14300));
  jxor g14179(.dina(n12028), .dinb(n12027), .dout(n14301));
  jor  g14180(.dina(n14301), .dinb(n6463), .dout(n14302));
  jand g14181(.dina(n11992), .dinb(n3855), .dout(n14303));
  jnot g14182(.din(n11997), .dout(n14304));
  jand g14183(.dina(n14304), .dinb(n3851), .dout(n14305));
  jand g14184(.dina(n14274), .dinb(n3858), .dout(n14306));
  jor  g14185(.dina(n14306), .dinb(n14305), .dout(n14307));
  jor  g14186(.dina(n14307), .dinb(n14303), .dout(n14308));
  jnot g14187(.din(n14308), .dout(n14309));
  jand g14188(.dina(n14309), .dinb(n14302), .dout(n14310));
  jor  g14189(.dina(n14310), .dinb(n14300), .dout(n14311));
  jand g14190(.dina(n13200), .dinb(n5897), .dout(n14312));
  jand g14191(.dina(n4692), .dinb(n4400), .dout(n14313));
  jand g14192(.dina(n14313), .dinb(n14312), .dout(n14314));
  jand g14193(.dina(n7159), .dinb(n1057), .dout(n14315));
  jand g14194(.dina(n14315), .dinb(n433), .dout(n14316));
  jand g14195(.dina(n607), .dinb(n322), .dout(n14317));
  jand g14196(.dina(n14317), .dinb(n717), .dout(n14318));
  jand g14197(.dina(n3075), .dinb(n771), .dout(n14319));
  jand g14198(.dina(n14319), .dinb(n14318), .dout(n14320));
  jand g14199(.dina(n14320), .dinb(n14316), .dout(n14321));
  jand g14200(.dina(n14321), .dinb(n4386), .dout(n14322));
  jand g14201(.dina(n14322), .dinb(n14314), .dout(n14323));
  jand g14202(.dina(n443), .dinb(n336), .dout(n14324));
  jand g14203(.dina(n14324), .dinb(n641), .dout(n14325));
  jand g14204(.dina(n14325), .dinb(n2277), .dout(n14326));
  jand g14205(.dina(n1641), .dinb(n208), .dout(n14327));
  jand g14206(.dina(n14327), .dinb(n435), .dout(n14328));
  jand g14207(.dina(n14328), .dinb(n12598), .dout(n14329));
  jand g14208(.dina(n14329), .dinb(n14326), .dout(n14330));
  jand g14209(.dina(n857), .dinb(n288), .dout(n14331));
  jand g14210(.dina(n719), .dinb(n707), .dout(n14332));
  jand g14211(.dina(n14332), .dinb(n14331), .dout(n14333));
  jand g14212(.dina(n14333), .dinb(n1603), .dout(n14334));
  jand g14213(.dina(n14334), .dinb(n4174), .dout(n14335));
  jand g14214(.dina(n14335), .dinb(n14330), .dout(n14336));
  jand g14215(.dina(n14336), .dinb(n7104), .dout(n14337));
  jand g14216(.dina(n12864), .dinb(n2784), .dout(n14338));
  jand g14217(.dina(n3445), .dinb(n2473), .dout(n14339));
  jand g14218(.dina(n14339), .dinb(n14338), .dout(n14340));
  jand g14219(.dina(n7069), .dinb(n512), .dout(n14341));
  jand g14220(.dina(n3503), .dinb(n177), .dout(n14342));
  jand g14221(.dina(n14342), .dinb(n14341), .dout(n14343));
  jand g14222(.dina(n14343), .dinb(n14340), .dout(n14344));
  jand g14223(.dina(n7003), .dinb(n3641), .dout(n14345));
  jand g14224(.dina(n14345), .dinb(n14344), .dout(n14346));
  jand g14225(.dina(n5982), .dinb(n2147), .dout(n14347));
  jand g14226(.dina(n14347), .dinb(n3556), .dout(n14348));
  jand g14227(.dina(n14348), .dinb(n12617), .dout(n14349));
  jand g14228(.dina(n14349), .dinb(n14346), .dout(n14350));
  jand g14229(.dina(n14350), .dinb(n14337), .dout(n14351));
  jand g14230(.dina(n14351), .dinb(n14323), .dout(n14352));
  jxor g14231(.dina(n12024), .dinb(n12023), .dout(n14353));
  jor  g14232(.dina(n14353), .dinb(n6463), .dout(n14354));
  jand g14233(.dina(n14274), .dinb(n3855), .dout(n14355));
  jnot g14234(.din(n11999), .dout(n14356));
  jand g14235(.dina(n14356), .dinb(n3851), .dout(n14357));
  jand g14236(.dina(n14304), .dinb(n3858), .dout(n14358));
  jor  g14237(.dina(n14358), .dinb(n14357), .dout(n14359));
  jor  g14238(.dina(n14359), .dinb(n14355), .dout(n14360));
  jnot g14239(.din(n14360), .dout(n14361));
  jand g14240(.dina(n14361), .dinb(n14354), .dout(n14362));
  jor  g14241(.dina(n14362), .dinb(n14352), .dout(n14363));
  jand g14242(.dina(n500), .dinb(n404), .dout(n14364));
  jand g14243(.dina(n1014), .dinb(n736), .dout(n14365));
  jand g14244(.dina(n14365), .dinb(n14364), .dout(n14366));
  jand g14245(.dina(n14366), .dinb(n669), .dout(n14367));
  jand g14246(.dina(n14367), .dinb(n4483), .dout(n14368));
  jand g14247(.dina(n2769), .dinb(n558), .dout(n14369));
  jand g14248(.dina(n14369), .dinb(n4231), .dout(n14370));
  jand g14249(.dina(n2672), .dinb(n2014), .dout(n14371));
  jand g14250(.dina(n877), .dinb(n563), .dout(n14372));
  jand g14251(.dina(n14372), .dinb(n14371), .dout(n14373));
  jand g14252(.dina(n14373), .dinb(n14370), .dout(n14374));
  jand g14253(.dina(n14374), .dinb(n14368), .dout(n14375));
  jand g14254(.dina(n14375), .dinb(n13235), .dout(n14376));
  jand g14255(.dina(n14376), .dinb(n2140), .dout(n14377));
  jand g14256(.dina(n1663), .dinb(n1119), .dout(n14378));
  jand g14257(.dina(n3260), .dinb(n880), .dout(n14379));
  jand g14258(.dina(n14379), .dinb(n14378), .dout(n14380));
  jand g14259(.dina(n424), .dinb(n336), .dout(n14381));
  jand g14260(.dina(n14381), .dinb(n967), .dout(n14382));
  jand g14261(.dina(n2160), .dinb(n484), .dout(n14383));
  jand g14262(.dina(n14383), .dinb(n14382), .dout(n14384));
  jand g14263(.dina(n14384), .dinb(n14380), .dout(n14385));
  jand g14264(.dina(n14385), .dinb(n2651), .dout(n14386));
  jand g14265(.dina(n14386), .dinb(n12439), .dout(n14387));
  jand g14266(.dina(n14387), .dinb(n631), .dout(n14388));
  jand g14267(.dina(n14388), .dinb(n14377), .dout(n14389));
  jxor g14268(.dina(n12020), .dinb(n12019), .dout(n14390));
  jor  g14269(.dina(n14390), .dinb(n6463), .dout(n14391));
  jand g14270(.dina(n14304), .dinb(n3855), .dout(n14392));
  jxor g14271(.dina(n11866), .dinb(n11864), .dout(n14393));
  jand g14272(.dina(n14393), .dinb(n3851), .dout(n14394));
  jand g14273(.dina(n14356), .dinb(n3858), .dout(n14395));
  jor  g14274(.dina(n14395), .dinb(n14394), .dout(n14396));
  jor  g14275(.dina(n14396), .dinb(n14392), .dout(n14397));
  jnot g14276(.din(n14397), .dout(n14398));
  jand g14277(.dina(n14398), .dinb(n14391), .dout(n14399));
  jor  g14278(.dina(n14399), .dinb(n14389), .dout(n14400));
  jand g14279(.dina(n445), .dinb(n366), .dout(n14401));
  jand g14280(.dina(n696), .dinb(n527), .dout(n14402));
  jand g14281(.dina(n14402), .dinb(n14401), .dout(n14403));
  jand g14282(.dina(n14403), .dinb(n4558), .dout(n14404));
  jand g14283(.dina(n14404), .dinb(n3261), .dout(n14405));
  jand g14284(.dina(n12494), .dinb(n1039), .dout(n14406));
  jand g14285(.dina(n14406), .dinb(n1704), .dout(n14407));
  jand g14286(.dina(n12259), .dinb(n3878), .dout(n14408));
  jand g14287(.dina(n14408), .dinb(n1299), .dout(n14409));
  jand g14288(.dina(n14409), .dinb(n14407), .dout(n14410));
  jand g14289(.dina(n14410), .dinb(n14405), .dout(n14411));
  jand g14290(.dina(n472), .dinb(n311), .dout(n14412));
  jand g14291(.dina(n14412), .dinb(n926), .dout(n14413));
  jand g14292(.dina(n14413), .dinb(n4163), .dout(n14414));
  jand g14293(.dina(n14414), .dinb(n761), .dout(n14415));
  jand g14294(.dina(n14415), .dinb(n13171), .dout(n14416));
  jand g14295(.dina(n14416), .dinb(n14411), .dout(n14417));
  jand g14296(.dina(n694), .dinb(n770), .dout(n14418));
  jand g14297(.dina(n14418), .dinb(n461), .dout(n14419));
  jand g14298(.dina(n536), .dinb(n478), .dout(n14420));
  jand g14299(.dina(n14420), .dinb(n806), .dout(n14421));
  jand g14300(.dina(n14421), .dinb(n14419), .dout(n14422));
  jand g14301(.dina(n14422), .dinb(n2050), .dout(n14423));
  jand g14302(.dina(n3041), .dinb(n2135), .dout(n14424));
  jand g14303(.dina(n14424), .dinb(n2514), .dout(n14425));
  jand g14304(.dina(n14425), .dinb(n5539), .dout(n14426));
  jand g14305(.dina(n14426), .dinb(n1469), .dout(n14427));
  jand g14306(.dina(n14427), .dinb(n14423), .dout(n14428));
  jand g14307(.dina(n14428), .dinb(n3102), .dout(n14429));
  jand g14308(.dina(n14429), .dinb(n14417), .dout(n14430));
  jand g14309(.dina(n14430), .dinb(n299), .dout(n14431));
  jxor g14310(.dina(n12016), .dinb(n12015), .dout(n14432));
  jor  g14311(.dina(n14432), .dinb(n6463), .dout(n14433));
  jand g14312(.dina(n14356), .dinb(n3855), .dout(n14434));
  jand g14313(.dina(n12006), .dinb(n3851), .dout(n14435));
  jand g14314(.dina(n14393), .dinb(n3858), .dout(n14436));
  jor  g14315(.dina(n14436), .dinb(n14435), .dout(n14437));
  jor  g14316(.dina(n14437), .dinb(n14434), .dout(n14438));
  jnot g14317(.din(n14438), .dout(n14439));
  jand g14318(.dina(n14439), .dinb(n14433), .dout(n14440));
  jor  g14319(.dina(n14440), .dinb(n14431), .dout(n14441));
  jand g14320(.dina(n4310), .dinb(n3478), .dout(n14442));
  jand g14321(.dina(n14442), .dinb(n7042), .dout(n14443));
  jand g14322(.dina(n1287), .dinb(n788), .dout(n14444));
  jand g14323(.dina(n14444), .dinb(n1591), .dout(n14445));
  jand g14324(.dina(n909), .dinb(n533), .dout(n14446));
  jand g14325(.dina(n494), .dinb(n280), .dout(n14447));
  jand g14326(.dina(n14447), .dinb(n14446), .dout(n14448));
  jand g14327(.dina(n14448), .dinb(n4235), .dout(n14449));
  jand g14328(.dina(n14449), .dinb(n14445), .dout(n14450));
  jand g14329(.dina(n14450), .dinb(n6031), .dout(n14451));
  jand g14330(.dina(n14451), .dinb(n14443), .dout(n14452));
  jand g14331(.dina(n12150), .dinb(n4690), .dout(n14453));
  jand g14332(.dina(n14453), .dinb(n14452), .dout(n14454));
  jand g14333(.dina(n14454), .dinb(n4207), .dout(n14455));
  jnot g14334(.din(n14455), .dout(n14456));
  jxor g14335(.dina(n12013), .dinb(n12007), .dout(n14457));
  jand g14336(.dina(n14457), .dinb(n732), .dout(n14458));
  jand g14337(.dina(n14393), .dinb(n3855), .dout(n14459));
  jand g14338(.dina(n12008), .dinb(n3851), .dout(n14460));
  jand g14339(.dina(n12006), .dinb(n3858), .dout(n14461));
  jor  g14340(.dina(n14461), .dinb(n14460), .dout(n14462));
  jor  g14341(.dina(n14462), .dinb(n14459), .dout(n14463));
  jor  g14342(.dina(n14463), .dinb(n14458), .dout(n14464));
  jand g14343(.dina(n14464), .dinb(n14456), .dout(n14465));
  jand g14344(.dina(n4523), .dinb(n4298), .dout(n14466));
  jand g14345(.dina(n14466), .dinb(n14293), .dout(n14467));
  jand g14346(.dina(n786), .dinb(n641), .dout(n14468));
  jand g14347(.dina(n14468), .dinb(n689), .dout(n14469));
  jand g14348(.dina(n407), .dinb(n286), .dout(n14470));
  jand g14349(.dina(n14470), .dinb(n3046), .dout(n14471));
  jand g14350(.dina(n14471), .dinb(n14469), .dout(n14472));
  jand g14351(.dina(n14472), .dinb(n1985), .dout(n14473));
  jand g14352(.dina(n983), .dinb(n615), .dout(n14474));
  jand g14353(.dina(n2261), .dinb(n1019), .dout(n14475));
  jand g14354(.dina(n14475), .dinb(n14474), .dout(n14476));
  jand g14355(.dina(n763), .dinb(n184), .dout(n14477));
  jand g14356(.dina(n14477), .dinb(n6417), .dout(n14478));
  jand g14357(.dina(n14478), .dinb(n4101), .dout(n14479));
  jand g14358(.dina(n14479), .dinb(n14476), .dout(n14480));
  jand g14359(.dina(n14480), .dinb(n14473), .dout(n14481));
  jand g14360(.dina(n14481), .dinb(n14467), .dout(n14482));
  jand g14361(.dina(n1314), .dinb(n696), .dout(n14483));
  jand g14362(.dina(n14483), .dinb(n143), .dout(n14484));
  jand g14363(.dina(n3092), .dinb(n2484), .dout(n14485));
  jand g14364(.dina(n2327), .dinb(n1868), .dout(n14486));
  jand g14365(.dina(n14486), .dinb(n14485), .dout(n14487));
  jand g14366(.dina(n14487), .dinb(n14484), .dout(n14488));
  jand g14367(.dina(n3813), .dinb(n2914), .dout(n14489));
  jand g14368(.dina(n2971), .dinb(n2926), .dout(n14490));
  jand g14369(.dina(n14490), .dinb(n14489), .dout(n14491));
  jand g14370(.dina(n14491), .dinb(n14488), .dout(n14492));
  jand g14371(.dina(n14492), .dinb(n7150), .dout(n14493));
  jand g14372(.dina(n14493), .dinb(n14482), .dout(n14494));
  jand g14373(.dina(n14494), .dinb(n3227), .dout(n14495));
  jnot g14374(.din(n14495), .dout(n14496));
  jxor g14375(.dina(n12010), .dinb(n12008), .dout(n14497));
  jand g14376(.dina(n14497), .dinb(n732), .dout(n14498));
  jand g14377(.dina(n12008), .dinb(n3855), .dout(n14499));
  jand g14378(.dina(n12010), .dinb(n3858), .dout(n14500));
  jor  g14379(.dina(n14500), .dinb(n14499), .dout(n14501));
  jor  g14380(.dina(n14501), .dinb(n14498), .dout(n14502));
  jand g14381(.dina(n14502), .dinb(n14496), .dout(n14503));
  jnot g14382(.din(n14503), .dout(n14504));
  jand g14383(.dina(n643), .dinb(n324), .dout(n14505));
  jand g14384(.dina(n14505), .dinb(n1829), .dout(n14506));
  jand g14385(.dina(n2327), .dinb(n1959), .dout(n14507));
  jand g14386(.dina(n14507), .dinb(n14506), .dout(n14508));
  jand g14387(.dina(n1144), .dinb(n503), .dout(n14509));
  jand g14388(.dina(n14509), .dinb(n276), .dout(n14510));
  jand g14389(.dina(n14510), .dinb(n2461), .dout(n14511));
  jand g14390(.dina(n793), .dinb(n533), .dout(n14512));
  jand g14391(.dina(n14512), .dinb(n1615), .dout(n14513));
  jand g14392(.dina(n14513), .dinb(n3012), .dout(n14514));
  jand g14393(.dina(n14514), .dinb(n14511), .dout(n14515));
  jand g14394(.dina(n14515), .dinb(n14508), .dout(n14516));
  jand g14395(.dina(n815), .dinb(n143), .dout(n14517));
  jand g14396(.dina(n14517), .dinb(n330), .dout(n14518));
  jand g14397(.dina(n14518), .dinb(n1333), .dout(n14519));
  jand g14398(.dina(n5815), .dinb(n585), .dout(n14520));
  jand g14399(.dina(n14520), .dinb(n14519), .dout(n14521));
  jand g14400(.dina(n1581), .dinb(n818), .dout(n14522));
  jand g14401(.dina(n14522), .dinb(n1160), .dout(n14523));
  jand g14402(.dina(n721), .dinb(n280), .dout(n14524));
  jand g14403(.dina(n1314), .dinb(n217), .dout(n14525));
  jand g14404(.dina(n14525), .dinb(n14524), .dout(n14526));
  jand g14405(.dina(n3793), .dinb(n601), .dout(n14527));
  jand g14406(.dina(n14527), .dinb(n14526), .dout(n14528));
  jand g14407(.dina(n14528), .dinb(n14523), .dout(n14529));
  jand g14408(.dina(n14529), .dinb(n14521), .dout(n14530));
  jand g14409(.dina(n14530), .dinb(n13881), .dout(n14531));
  jand g14410(.dina(n14531), .dinb(n14516), .dout(n14532));
  jand g14411(.dina(n14532), .dinb(n13164), .dout(n14533));
  jor  g14412(.dina(n14533), .dinb(n14504), .dout(n14534));
  jxor g14413(.dina(n14533), .dinb(n14504), .dout(n14535));
  jand g14414(.dina(n12011), .dinb(n12008), .dout(n14536));
  jxor g14415(.dina(n14536), .dinb(n12006), .dout(n14537));
  jand g14416(.dina(n14537), .dinb(n732), .dout(n14538));
  jand g14417(.dina(n12006), .dinb(n3855), .dout(n14539));
  jand g14418(.dina(n12008), .dinb(n3858), .dout(n14540));
  jand g14419(.dina(n12010), .dinb(n3851), .dout(n14541));
  jor  g14420(.dina(n14541), .dinb(n14540), .dout(n14542));
  jor  g14421(.dina(n14542), .dinb(n14539), .dout(n14543));
  jor  g14422(.dina(n14543), .dinb(n14538), .dout(n14544));
  jand g14423(.dina(n14544), .dinb(n14535), .dout(n14545));
  jnot g14424(.din(n14545), .dout(n14546));
  jand g14425(.dina(n14546), .dinb(n14534), .dout(n14547));
  jnot g14426(.din(n14547), .dout(n14548));
  jxor g14427(.dina(n14464), .dinb(n14456), .dout(n14549));
  jand g14428(.dina(n14549), .dinb(n14548), .dout(n14550));
  jor  g14429(.dina(n14550), .dinb(n14465), .dout(n14551));
  jxor g14430(.dina(n14440), .dinb(n14431), .dout(n14552));
  jand g14431(.dina(n14552), .dinb(n14551), .dout(n14553));
  jnot g14432(.din(n14553), .dout(n14554));
  jand g14433(.dina(n14554), .dinb(n14441), .dout(n14555));
  jnot g14434(.din(n14555), .dout(n14556));
  jxor g14435(.dina(n14399), .dinb(n14389), .dout(n14557));
  jand g14436(.dina(n14557), .dinb(n14556), .dout(n14558));
  jnot g14437(.din(n14558), .dout(n14559));
  jand g14438(.dina(n14559), .dinb(n14400), .dout(n14560));
  jnot g14439(.din(n14560), .dout(n14561));
  jxor g14440(.dina(n14362), .dinb(n14352), .dout(n14562));
  jand g14441(.dina(n14562), .dinb(n14561), .dout(n14563));
  jnot g14442(.din(n14563), .dout(n14564));
  jand g14443(.dina(n14564), .dinb(n14363), .dout(n14565));
  jnot g14444(.din(n14565), .dout(n14566));
  jxor g14445(.dina(n14310), .dinb(n14300), .dout(n14567));
  jand g14446(.dina(n14567), .dinb(n14566), .dout(n14568));
  jnot g14447(.din(n14568), .dout(n14569));
  jand g14448(.dina(n14569), .dinb(n14311), .dout(n14570));
  jnot g14449(.din(n14570), .dout(n14571));
  jxor g14450(.dina(n14280), .dinb(n14270), .dout(n14572));
  jand g14451(.dina(n14572), .dinb(n14571), .dout(n14573));
  jnot g14452(.din(n14573), .dout(n14574));
  jand g14453(.dina(n14574), .dinb(n14281), .dout(n14575));
  jnot g14454(.din(n14575), .dout(n14576));
  jxor g14455(.dina(n14256), .dinb(n14247), .dout(n14577));
  jand g14456(.dina(n14577), .dinb(n14576), .dout(n14578));
  jnot g14457(.din(n14578), .dout(n14579));
  jand g14458(.dina(n14579), .dinb(n14257), .dout(n14580));
  jnot g14459(.din(n14580), .dout(n14581));
  jxor g14460(.dina(n14229), .dinb(n14220), .dout(n14582));
  jand g14461(.dina(n14582), .dinb(n14581), .dout(n14583));
  jnot g14462(.din(n14583), .dout(n14584));
  jand g14463(.dina(n14584), .dinb(n14230), .dout(n14585));
  jnot g14464(.din(n14585), .dout(n14586));
  jxor g14465(.dina(n13906), .dinb(n13898), .dout(n14587));
  jand g14466(.dina(n14587), .dinb(n14586), .dout(n14588));
  jnot g14467(.din(n14588), .dout(n14589));
  jxor g14468(.dina(n14587), .dinb(n14586), .dout(n14590));
  jnot g14469(.din(n14590), .dout(n14591));
  jand g14470(.dina(n13924), .dinb(n4449), .dout(n14592));
  jand g14471(.dina(n11974), .dinb(n4453), .dout(n14593));
  jand g14472(.dina(n11976), .dinb(n4457), .dout(n14594));
  jand g14473(.dina(n11978), .dinb(n4461), .dout(n14595));
  jor  g14474(.dina(n14595), .dinb(n14594), .dout(n14596));
  jor  g14475(.dina(n14596), .dinb(n14593), .dout(n14597));
  jor  g14476(.dina(n14597), .dinb(n14592), .dout(n14598));
  jxor g14477(.dina(n14598), .dinb(n88), .dout(n14599));
  jor  g14478(.dina(n14599), .dinb(n14591), .dout(n14600));
  jand g14479(.dina(n14600), .dinb(n14589), .dout(n14601));
  jnot g14480(.din(n14601), .dout(n14602));
  jxor g14481(.dina(n14201), .dinb(n14193), .dout(n14603));
  jand g14482(.dina(n14603), .dinb(n14602), .dout(n14604));
  jor  g14483(.dina(n14604), .dinb(n14202), .dout(n14605));
  jxor g14484(.dina(n14191), .dinb(n14183), .dout(n14606));
  jand g14485(.dina(n14606), .dinb(n14605), .dout(n14607));
  jor  g14486(.dina(n14607), .dinb(n14192), .dout(n14608));
  jxor g14487(.dina(n13931), .dinb(n13923), .dout(n14609));
  jand g14488(.dina(n14609), .dinb(n14608), .dout(n14610));
  jnot g14489(.din(n14610), .dout(n14611));
  jxor g14490(.dina(n14609), .dinb(n14608), .dout(n14612));
  jnot g14491(.din(n14612), .dout(n14613));
  jand g14492(.dina(n13682), .dinb(n4449), .dout(n14614));
  jand g14493(.dina(n11968), .dinb(n4453), .dout(n14615));
  jand g14494(.dina(n11970), .dinb(n4457), .dout(n14616));
  jand g14495(.dina(n11972), .dinb(n4461), .dout(n14617));
  jor  g14496(.dina(n14617), .dinb(n14616), .dout(n14618));
  jor  g14497(.dina(n14618), .dinb(n14615), .dout(n14619));
  jor  g14498(.dina(n14619), .dinb(n14614), .dout(n14620));
  jxor g14499(.dina(n14620), .dinb(n88), .dout(n14621));
  jor  g14500(.dina(n14621), .dinb(n14613), .dout(n14622));
  jand g14501(.dina(n14622), .dinb(n14611), .dout(n14623));
  jnot g14502(.din(n14623), .dout(n14624));
  jxor g14503(.dina(n13946), .dinb(n13938), .dout(n14625));
  jand g14504(.dina(n14625), .dinb(n14624), .dout(n14626));
  jnot g14505(.din(n14626), .dout(n14627));
  jxor g14506(.dina(n14625), .dinb(n14624), .dout(n14628));
  jnot g14507(.din(n14628), .dout(n14629));
  jand g14508(.dina(n13116), .dinb(n75), .dout(n14630));
  jand g14509(.dina(n11960), .dinb(n4933), .dout(n14631));
  jand g14510(.dina(n11962), .dinb(n4918), .dout(n14632));
  jand g14511(.dina(n11964), .dinb(n4745), .dout(n14633));
  jor  g14512(.dina(n14633), .dinb(n14632), .dout(n14634));
  jor  g14513(.dina(n14634), .dinb(n14631), .dout(n14635));
  jor  g14514(.dina(n14635), .dinb(n14630), .dout(n14636));
  jxor g14515(.dina(n14636), .dinb(n68), .dout(n14637));
  jor  g14516(.dina(n14637), .dinb(n14629), .dout(n14638));
  jand g14517(.dina(n14638), .dinb(n14627), .dout(n14639));
  jnot g14518(.din(n14639), .dout(n14640));
  jxor g14519(.dina(n14083), .dinb(n14082), .dout(n14641));
  jand g14520(.dina(n14641), .dinb(n14640), .dout(n14642));
  jnot g14521(.din(n14642), .dout(n14643));
  jxor g14522(.dina(n14641), .dinb(n14640), .dout(n14644));
  jnot g14523(.din(n14644), .dout(n14645));
  jand g14524(.dina(n12510), .dinb(n5365), .dout(n14646));
  jand g14525(.dina(n11952), .dinb(n5500), .dout(n14647));
  jand g14526(.dina(n11954), .dinb(n5424), .dout(n14648));
  jand g14527(.dina(n11956), .dinb(n5363), .dout(n14649));
  jor  g14528(.dina(n14649), .dinb(n14648), .dout(n14650));
  jor  g14529(.dina(n14650), .dinb(n14647), .dout(n14651));
  jor  g14530(.dina(n14651), .dinb(n14646), .dout(n14652));
  jxor g14531(.dina(n14652), .dinb(n72), .dout(n14653));
  jor  g14532(.dina(n14653), .dinb(n14645), .dout(n14654));
  jand g14533(.dina(n14654), .dinb(n14643), .dout(n14655));
  jnot g14534(.din(n14655), .dout(n14656));
  jxor g14535(.dina(n14181), .dinb(n14173), .dout(n14657));
  jand g14536(.dina(n14657), .dinb(n14656), .dout(n14658));
  jnot g14537(.din(n14658), .dout(n14659));
  jand g14538(.dina(n14659), .dinb(n14182), .dout(n14660));
  jnot g14539(.din(n14660), .dout(n14661));
  jxor g14540(.dina(n14105), .dinb(n14097), .dout(n14662));
  jand g14541(.dina(n14662), .dinb(n14661), .dout(n14663));
  jnot g14542(.din(n14663), .dout(n14664));
  jxor g14543(.dina(n14662), .dinb(n14661), .dout(n14665));
  jnot g14544(.din(n14665), .dout(n14666));
  jand g14545(.dina(n12751), .dinb(n5693), .dout(n14667));
  jand g14546(.dina(n11942), .dinb(n6209), .dout(n14668));
  jand g14547(.dina(n11944), .dinb(n6131), .dout(n14669));
  jand g14548(.dina(n11946), .dinb(n5691), .dout(n14670));
  jor  g14549(.dina(n14670), .dinb(n14669), .dout(n14671));
  jor  g14550(.dina(n14671), .dinb(n14668), .dout(n14672));
  jor  g14551(.dina(n14672), .dinb(n14667), .dout(n14673));
  jxor g14552(.dina(n14673), .dinb(n4247), .dout(n14674));
  jor  g14553(.dina(n14674), .dinb(n14666), .dout(n14675));
  jand g14554(.dina(n14675), .dinb(n14664), .dout(n14676));
  jnot g14555(.din(n14676), .dout(n14677));
  jxor g14556(.dina(n14121), .dinb(n14113), .dout(n14678));
  jand g14557(.dina(n14678), .dinb(n14677), .dout(n14679));
  jnot g14558(.din(n14679), .dout(n14680));
  jxor g14559(.dina(n14678), .dinb(n14677), .dout(n14681));
  jnot g14560(.din(n14681), .dout(n14682));
  jand g14561(.dina(n12841), .dinb(n6340), .dout(n14683));
  jand g14562(.dina(n12783), .dinb(n6798), .dout(n14684));
  jand g14563(.dina(n12766), .dinb(n6556), .dout(n14685));
  jand g14564(.dina(n12177), .dinb(n6338), .dout(n14686));
  jor  g14565(.dina(n14686), .dinb(n14685), .dout(n14687));
  jor  g14566(.dina(n14687), .dinb(n14684), .dout(n14688));
  jor  g14567(.dina(n14688), .dinb(n14683), .dout(n14689));
  jxor g14568(.dina(n14689), .dinb(n5064), .dout(n14690));
  jor  g14569(.dina(n14690), .dinb(n14682), .dout(n14691));
  jand g14570(.dina(n14691), .dinb(n14680), .dout(n14692));
  jnot g14571(.din(n14692), .dout(n14693));
  jxor g14572(.dina(n14170), .dinb(n14162), .dout(n14694));
  jand g14573(.dina(n14694), .dinb(n14693), .dout(n14695));
  jnot g14574(.din(n14695), .dout(n14696));
  jand g14575(.dina(n14696), .dinb(n14171), .dout(n14697));
  jnot g14576(.din(n14697), .dout(n14698));
  jxor g14577(.dina(n14142), .dinb(n14134), .dout(n14699));
  jand g14578(.dina(n14699), .dinb(n14698), .dout(n14700));
  jnot g14579(.din(n14700), .dout(n14701));
  jxor g14580(.dina(n14699), .dinb(n14698), .dout(n14702));
  jnot g14581(.din(n14702), .dout(n14703));
  jor  g14582(.dina(n12814), .dinb(n6935), .dout(n14705));
  jand g14583(.dina(n14147), .dinb(n14705), .dout(n14709));
  jand g14584(.dina(n14709), .dinb(n6937), .dout(n14710));
  jxor g14585(.dina(n14710), .dinb(\a[14] ), .dout(n14711));
  jor  g14586(.dina(n14711), .dinb(n14703), .dout(n14712));
  jand g14587(.dina(n14712), .dinb(n14701), .dout(n14713));
  jnot g14588(.din(n14713), .dout(n14714));
  jxor g14589(.dina(n14154), .dinb(n14153), .dout(n14715));
  jand g14590(.dina(n14715), .dinb(n14714), .dout(n14716));
  jxor g14591(.dina(n14715), .dinb(n14714), .dout(n14717));
  jxor g14592(.dina(n14657), .dinb(n14656), .dout(n14718));
  jnot g14593(.din(n14718), .dout(n14719));
  jand g14594(.dina(n12189), .dinb(n5693), .dout(n14720));
  jand g14595(.dina(n11944), .dinb(n6209), .dout(n14721));
  jand g14596(.dina(n11946), .dinb(n6131), .dout(n14722));
  jand g14597(.dina(n11948), .dinb(n5691), .dout(n14723));
  jor  g14598(.dina(n14723), .dinb(n14722), .dout(n14724));
  jor  g14599(.dina(n14724), .dinb(n14721), .dout(n14725));
  jor  g14600(.dina(n14725), .dinb(n14720), .dout(n14726));
  jxor g14601(.dina(n14726), .dinb(n4247), .dout(n14727));
  jor  g14602(.dina(n14727), .dinb(n14719), .dout(n14728));
  jand g14603(.dina(n13134), .dinb(n75), .dout(n14729));
  jand g14604(.dina(n11962), .dinb(n4933), .dout(n14730));
  jand g14605(.dina(n11964), .dinb(n4918), .dout(n14731));
  jand g14606(.dina(n11966), .dinb(n4745), .dout(n14732));
  jor  g14607(.dina(n14732), .dinb(n14731), .dout(n14733));
  jor  g14608(.dina(n14733), .dinb(n14730), .dout(n14734));
  jor  g14609(.dina(n14734), .dinb(n14729), .dout(n14735));
  jxor g14610(.dina(n14735), .dinb(n68), .dout(n14736));
  jnot g14611(.din(n14736), .dout(n14737));
  jxor g14612(.dina(n14621), .dinb(n14613), .dout(n14738));
  jand g14613(.dina(n14738), .dinb(n14737), .dout(n14739));
  jxor g14614(.dina(n14606), .dinb(n14605), .dout(n14740));
  jnot g14615(.din(n14740), .dout(n14741));
  jand g14616(.dina(n13806), .dinb(n4449), .dout(n14742));
  jand g14617(.dina(n11970), .dinb(n4453), .dout(n14743));
  jand g14618(.dina(n11972), .dinb(n4457), .dout(n14744));
  jand g14619(.dina(n11974), .dinb(n4461), .dout(n14745));
  jor  g14620(.dina(n14745), .dinb(n14744), .dout(n14746));
  jor  g14621(.dina(n14746), .dinb(n14743), .dout(n14747));
  jor  g14622(.dina(n14747), .dinb(n14742), .dout(n14748));
  jxor g14623(.dina(n14748), .dinb(n88), .dout(n14749));
  jor  g14624(.dina(n14749), .dinb(n14741), .dout(n14750));
  jand g14625(.dina(n13470), .dinb(n75), .dout(n14751));
  jand g14626(.dina(n11964), .dinb(n4933), .dout(n14752));
  jand g14627(.dina(n11966), .dinb(n4918), .dout(n14753));
  jand g14628(.dina(n11968), .dinb(n4745), .dout(n14754));
  jor  g14629(.dina(n14754), .dinb(n14753), .dout(n14755));
  jor  g14630(.dina(n14755), .dinb(n14752), .dout(n14756));
  jor  g14631(.dina(n14756), .dinb(n14751), .dout(n14757));
  jxor g14632(.dina(n14757), .dinb(n68), .dout(n14758));
  jnot g14633(.din(n14758), .dout(n14759));
  jxor g14634(.dina(n14749), .dinb(n14741), .dout(n14760));
  jand g14635(.dina(n14760), .dinb(n14759), .dout(n14761));
  jnot g14636(.din(n14761), .dout(n14762));
  jand g14637(.dina(n14762), .dinb(n14750), .dout(n14763));
  jnot g14638(.din(n14763), .dout(n14764));
  jxor g14639(.dina(n14738), .dinb(n14737), .dout(n14765));
  jand g14640(.dina(n14765), .dinb(n14764), .dout(n14766));
  jor  g14641(.dina(n14766), .dinb(n14739), .dout(n14767));
  jxor g14642(.dina(n14637), .dinb(n14629), .dout(n14768));
  jand g14643(.dina(n14768), .dinb(n14767), .dout(n14769));
  jnot g14644(.din(n14769), .dout(n14770));
  jxor g14645(.dina(n14768), .dinb(n14767), .dout(n14771));
  jnot g14646(.din(n14771), .dout(n14772));
  jand g14647(.dina(n12472), .dinb(n5365), .dout(n14773));
  jand g14648(.dina(n11954), .dinb(n5500), .dout(n14774));
  jand g14649(.dina(n11956), .dinb(n5424), .dout(n14775));
  jand g14650(.dina(n11958), .dinb(n5363), .dout(n14776));
  jor  g14651(.dina(n14776), .dinb(n14775), .dout(n14777));
  jor  g14652(.dina(n14777), .dinb(n14774), .dout(n14778));
  jor  g14653(.dina(n14778), .dinb(n14773), .dout(n14779));
  jxor g14654(.dina(n14779), .dinb(n72), .dout(n14780));
  jor  g14655(.dina(n14780), .dinb(n14772), .dout(n14781));
  jand g14656(.dina(n14781), .dinb(n14770), .dout(n14782));
  jnot g14657(.din(n14782), .dout(n14783));
  jxor g14658(.dina(n14653), .dinb(n14645), .dout(n14784));
  jand g14659(.dina(n14784), .dinb(n14783), .dout(n14785));
  jnot g14660(.din(n14785), .dout(n14786));
  jxor g14661(.dina(n14784), .dinb(n14783), .dout(n14787));
  jnot g14662(.din(n14787), .dout(n14788));
  jand g14663(.dina(n12519), .dinb(n5693), .dout(n14789));
  jand g14664(.dina(n11946), .dinb(n6209), .dout(n14790));
  jand g14665(.dina(n11948), .dinb(n6131), .dout(n14791));
  jand g14666(.dina(n11950), .dinb(n5691), .dout(n14792));
  jor  g14667(.dina(n14792), .dinb(n14791), .dout(n14793));
  jor  g14668(.dina(n14793), .dinb(n14790), .dout(n14794));
  jor  g14669(.dina(n14794), .dinb(n14789), .dout(n14795));
  jxor g14670(.dina(n14795), .dinb(n4247), .dout(n14796));
  jor  g14671(.dina(n14796), .dinb(n14788), .dout(n14797));
  jand g14672(.dina(n14797), .dinb(n14786), .dout(n14798));
  jnot g14673(.din(n14798), .dout(n14799));
  jxor g14674(.dina(n14727), .dinb(n14719), .dout(n14800));
  jand g14675(.dina(n14800), .dinb(n14799), .dout(n14801));
  jnot g14676(.din(n14801), .dout(n14802));
  jand g14677(.dina(n14802), .dinb(n14728), .dout(n14803));
  jnot g14678(.din(n14803), .dout(n14804));
  jxor g14679(.dina(n14674), .dinb(n14666), .dout(n14805));
  jand g14680(.dina(n14805), .dinb(n14804), .dout(n14806));
  jnot g14681(.din(n14806), .dout(n14807));
  jxor g14682(.dina(n14805), .dinb(n14804), .dout(n14808));
  jnot g14683(.din(n14808), .dout(n14809));
  jand g14684(.dina(n12768), .dinb(n6340), .dout(n14810));
  jand g14685(.dina(n12766), .dinb(n6798), .dout(n14811));
  jand g14686(.dina(n12177), .dinb(n6556), .dout(n14812));
  jand g14687(.dina(n11941), .dinb(n6338), .dout(n14813));
  jor  g14688(.dina(n14813), .dinb(n14812), .dout(n14814));
  jor  g14689(.dina(n14814), .dinb(n14811), .dout(n14815));
  jor  g14690(.dina(n14815), .dinb(n14810), .dout(n14816));
  jxor g14691(.dina(n14816), .dinb(n5064), .dout(n14817));
  jor  g14692(.dina(n14817), .dinb(n14809), .dout(n14818));
  jand g14693(.dina(n14818), .dinb(n14807), .dout(n14819));
  jnot g14694(.din(n14819), .dout(n14820));
  jxor g14695(.dina(n14690), .dinb(n14682), .dout(n14821));
  jand g14696(.dina(n14821), .dinb(n14820), .dout(n14822));
  jnot g14697(.din(n14822), .dout(n14823));
  jxor g14698(.dina(n14821), .dinb(n14820), .dout(n14824));
  jnot g14699(.din(n14824), .dout(n14825));
  jand g14700(.dina(n12919), .dinb(n6936), .dout(n14826));
  jand g14701(.dina(n12815), .dinb(n7741), .dout(n14827));
  jand g14702(.dina(n12795), .dinb(n7613), .dout(n14828));
  jand g14703(.dina(n12782), .dinb(n6934), .dout(n14829));
  jor  g14704(.dina(n14829), .dinb(n14828), .dout(n14830));
  jor  g14705(.dina(n14830), .dinb(n14827), .dout(n14831));
  jor  g14706(.dina(n14831), .dinb(n14826), .dout(n14832));
  jxor g14707(.dina(n14832), .dinb(n5292), .dout(n14833));
  jor  g14708(.dina(n14833), .dinb(n14825), .dout(n14834));
  jand g14709(.dina(n14834), .dinb(n14823), .dout(n14835));
  jand g14710(.dina(n13022), .dinb(n6936), .dout(n14836));
  jand g14711(.dina(n12815), .dinb(n7613), .dout(n14838));
  jand g14712(.dina(n12795), .dinb(n6934), .dout(n14839));
  jor  g14713(.dina(n14839), .dinb(n14838), .dout(n14840));
  jor  g14714(.dina(n14840), .dinb(n7741), .dout(n14841));
  jor  g14715(.dina(n14841), .dinb(n14836), .dout(n14842));
  jxor g14716(.dina(n14842), .dinb(n5292), .dout(n14843));
  jor  g14717(.dina(n14843), .dinb(n14835), .dout(n14844));
  jxor g14718(.dina(n14694), .dinb(n14693), .dout(n14845));
  jxor g14719(.dina(n14843), .dinb(n14835), .dout(n14846));
  jand g14720(.dina(n14846), .dinb(n14845), .dout(n14847));
  jnot g14721(.din(n14847), .dout(n14848));
  jand g14722(.dina(n14848), .dinb(n14844), .dout(n14849));
  jnot g14723(.din(n14849), .dout(n14850));
  jxor g14724(.dina(n14711), .dinb(n14703), .dout(n14851));
  jand g14725(.dina(n14851), .dinb(n14850), .dout(n14852));
  jxor g14726(.dina(n14800), .dinb(n14799), .dout(n14853));
  jnot g14727(.din(n14853), .dout(n14854));
  jand g14728(.dina(n12179), .dinb(n6340), .dout(n14855));
  jand g14729(.dina(n12177), .dinb(n6798), .dout(n14856));
  jand g14730(.dina(n11941), .dinb(n6556), .dout(n14857));
  jand g14731(.dina(n11942), .dinb(n6338), .dout(n14858));
  jor  g14732(.dina(n14858), .dinb(n14857), .dout(n14859));
  jor  g14733(.dina(n14859), .dinb(n14856), .dout(n14860));
  jor  g14734(.dina(n14860), .dinb(n14855), .dout(n14861));
  jxor g14735(.dina(n14861), .dinb(n5064), .dout(n14862));
  jor  g14736(.dina(n14862), .dinb(n14854), .dout(n14863));
  jxor g14737(.dina(n14765), .dinb(n14764), .dout(n14864));
  jnot g14738(.din(n14864), .dout(n14865));
  jand g14739(.dina(n12639), .dinb(n5365), .dout(n14866));
  jand g14740(.dina(n11956), .dinb(n5500), .dout(n14867));
  jand g14741(.dina(n11958), .dinb(n5424), .dout(n14868));
  jand g14742(.dina(n11960), .dinb(n5363), .dout(n14869));
  jor  g14743(.dina(n14869), .dinb(n14868), .dout(n14870));
  jor  g14744(.dina(n14870), .dinb(n14867), .dout(n14871));
  jor  g14745(.dina(n14871), .dinb(n14866), .dout(n14872));
  jxor g14746(.dina(n14872), .dinb(n72), .dout(n14873));
  jor  g14747(.dina(n14873), .dinb(n14865), .dout(n14874));
  jxor g14748(.dina(n14603), .dinb(n14602), .dout(n14875));
  jnot g14749(.din(n14875), .dout(n14876));
  jand g14750(.dina(n13664), .dinb(n4449), .dout(n14877));
  jand g14751(.dina(n11972), .dinb(n4453), .dout(n14878));
  jand g14752(.dina(n11974), .dinb(n4457), .dout(n14879));
  jand g14753(.dina(n11976), .dinb(n4461), .dout(n14880));
  jor  g14754(.dina(n14880), .dinb(n14879), .dout(n14881));
  jor  g14755(.dina(n14881), .dinb(n14878), .dout(n14882));
  jor  g14756(.dina(n14882), .dinb(n14877), .dout(n14883));
  jxor g14757(.dina(n14883), .dinb(n88), .dout(n14884));
  jor  g14758(.dina(n14884), .dinb(n14876), .dout(n14885));
  jand g14759(.dina(n13268), .dinb(n75), .dout(n14886));
  jand g14760(.dina(n11966), .dinb(n4933), .dout(n14887));
  jand g14761(.dina(n11970), .dinb(n4745), .dout(n14888));
  jand g14762(.dina(n11968), .dinb(n4918), .dout(n14889));
  jor  g14763(.dina(n14889), .dinb(n14888), .dout(n14890));
  jor  g14764(.dina(n14890), .dinb(n14887), .dout(n14891));
  jor  g14765(.dina(n14891), .dinb(n14886), .dout(n14892));
  jxor g14766(.dina(n14892), .dinb(n68), .dout(n14893));
  jnot g14767(.din(n14893), .dout(n14894));
  jxor g14768(.dina(n14884), .dinb(n14876), .dout(n14895));
  jand g14769(.dina(n14895), .dinb(n14894), .dout(n14896));
  jnot g14770(.din(n14896), .dout(n14897));
  jand g14771(.dina(n14897), .dinb(n14885), .dout(n14898));
  jnot g14772(.din(n14898), .dout(n14899));
  jxor g14773(.dina(n14760), .dinb(n14759), .dout(n14900));
  jand g14774(.dina(n14900), .dinb(n14899), .dout(n14901));
  jnot g14775(.din(n14901), .dout(n14902));
  jxor g14776(.dina(n14900), .dinb(n14899), .dout(n14903));
  jnot g14777(.din(n14903), .dout(n14904));
  jand g14778(.dina(n12624), .dinb(n5365), .dout(n14905));
  jand g14779(.dina(n11958), .dinb(n5500), .dout(n14906));
  jand g14780(.dina(n11960), .dinb(n5424), .dout(n14907));
  jand g14781(.dina(n11962), .dinb(n5363), .dout(n14908));
  jor  g14782(.dina(n14908), .dinb(n14907), .dout(n14909));
  jor  g14783(.dina(n14909), .dinb(n14906), .dout(n14910));
  jor  g14784(.dina(n14910), .dinb(n14905), .dout(n14911));
  jxor g14785(.dina(n14911), .dinb(n72), .dout(n14912));
  jor  g14786(.dina(n14912), .dinb(n14904), .dout(n14913));
  jand g14787(.dina(n14913), .dinb(n14902), .dout(n14914));
  jnot g14788(.din(n14914), .dout(n14915));
  jxor g14789(.dina(n14873), .dinb(n14865), .dout(n14916));
  jand g14790(.dina(n14916), .dinb(n14915), .dout(n14917));
  jnot g14791(.din(n14917), .dout(n14918));
  jand g14792(.dina(n14918), .dinb(n14874), .dout(n14919));
  jnot g14793(.din(n14919), .dout(n14920));
  jxor g14794(.dina(n14780), .dinb(n14772), .dout(n14921));
  jand g14795(.dina(n14921), .dinb(n14920), .dout(n14922));
  jnot g14796(.din(n14922), .dout(n14923));
  jxor g14797(.dina(n14921), .dinb(n14920), .dout(n14924));
  jnot g14798(.din(n14924), .dout(n14925));
  jand g14799(.dina(n12654), .dinb(n5693), .dout(n14926));
  jand g14800(.dina(n11948), .dinb(n6209), .dout(n14927));
  jand g14801(.dina(n11950), .dinb(n6131), .dout(n14928));
  jand g14802(.dina(n11952), .dinb(n5691), .dout(n14929));
  jor  g14803(.dina(n14929), .dinb(n14928), .dout(n14930));
  jor  g14804(.dina(n14930), .dinb(n14927), .dout(n14931));
  jor  g14805(.dina(n14931), .dinb(n14926), .dout(n14932));
  jxor g14806(.dina(n14932), .dinb(n4247), .dout(n14933));
  jor  g14807(.dina(n14933), .dinb(n14925), .dout(n14934));
  jand g14808(.dina(n14934), .dinb(n14923), .dout(n14935));
  jnot g14809(.din(n14935), .dout(n14936));
  jxor g14810(.dina(n14796), .dinb(n14788), .dout(n14937));
  jand g14811(.dina(n14937), .dinb(n14936), .dout(n14938));
  jnot g14812(.din(n14938), .dout(n14939));
  jxor g14813(.dina(n14937), .dinb(n14936), .dout(n14940));
  jnot g14814(.din(n14940), .dout(n14941));
  jand g14815(.dina(n12671), .dinb(n6340), .dout(n14942));
  jand g14816(.dina(n11941), .dinb(n6798), .dout(n14943));
  jand g14817(.dina(n11942), .dinb(n6556), .dout(n14944));
  jand g14818(.dina(n11944), .dinb(n6338), .dout(n14945));
  jor  g14819(.dina(n14945), .dinb(n14944), .dout(n14946));
  jor  g14820(.dina(n14946), .dinb(n14943), .dout(n14947));
  jor  g14821(.dina(n14947), .dinb(n14942), .dout(n14948));
  jxor g14822(.dina(n14948), .dinb(n5064), .dout(n14949));
  jor  g14823(.dina(n14949), .dinb(n14941), .dout(n14950));
  jand g14824(.dina(n14950), .dinb(n14939), .dout(n14951));
  jnot g14825(.din(n14951), .dout(n14952));
  jxor g14826(.dina(n14862), .dinb(n14854), .dout(n14953));
  jand g14827(.dina(n14953), .dinb(n14952), .dout(n14954));
  jnot g14828(.din(n14954), .dout(n14955));
  jand g14829(.dina(n14955), .dinb(n14863), .dout(n14956));
  jnot g14830(.din(n14956), .dout(n14957));
  jxor g14831(.dina(n14817), .dinb(n14809), .dout(n14958));
  jand g14832(.dina(n14958), .dinb(n14957), .dout(n14959));
  jnot g14833(.din(n14959), .dout(n14960));
  jxor g14834(.dina(n14958), .dinb(n14957), .dout(n14961));
  jnot g14835(.din(n14961), .dout(n14962));
  jand g14836(.dina(n12797), .dinb(n6936), .dout(n14963));
  jand g14837(.dina(n12795), .dinb(n7741), .dout(n14964));
  jand g14838(.dina(n12782), .dinb(n7613), .dout(n14965));
  jand g14839(.dina(n12783), .dinb(n6934), .dout(n14966));
  jor  g14840(.dina(n14966), .dinb(n14965), .dout(n14967));
  jor  g14841(.dina(n14967), .dinb(n14964), .dout(n14968));
  jor  g14842(.dina(n14968), .dinb(n14963), .dout(n14969));
  jxor g14843(.dina(n14969), .dinb(n5292), .dout(n14970));
  jor  g14844(.dina(n14970), .dinb(n14962), .dout(n14971));
  jand g14845(.dina(n14971), .dinb(n14960), .dout(n14972));
  jand g14846(.dina(n8440), .dinb(n8155), .dout(n14975));
  jor  g14847(.dina(n13109), .dinb(n14972), .dout(n14980));
  jxor g14848(.dina(n13109), .dinb(n14972), .dout(n14981));
  jxor g14849(.dina(n14833), .dinb(n14825), .dout(n14982));
  jand g14850(.dina(n14982), .dinb(n14981), .dout(n14983));
  jnot g14851(.din(n14983), .dout(n14984));
  jand g14852(.dina(n14984), .dinb(n14980), .dout(n14985));
  jnot g14853(.din(n14985), .dout(n14986));
  jxor g14854(.dina(n14846), .dinb(n14845), .dout(n14987));
  jand g14855(.dina(n14987), .dinb(n14986), .dout(n14988));
  jxor g14856(.dina(n14953), .dinb(n14952), .dout(n14989));
  jnot g14857(.din(n14989), .dout(n14990));
  jand g14858(.dina(n12938), .dinb(n6936), .dout(n14991));
  jand g14859(.dina(n12782), .dinb(n7741), .dout(n14992));
  jand g14860(.dina(n12783), .dinb(n7613), .dout(n14993));
  jand g14861(.dina(n12766), .dinb(n6934), .dout(n14994));
  jor  g14862(.dina(n14994), .dinb(n14993), .dout(n14995));
  jor  g14863(.dina(n14995), .dinb(n14992), .dout(n14996));
  jor  g14864(.dina(n14996), .dinb(n14991), .dout(n14997));
  jxor g14865(.dina(n14997), .dinb(n5292), .dout(n14998));
  jor  g14866(.dina(n14998), .dinb(n14990), .dout(n14999));
  jxor g14867(.dina(n14916), .dinb(n14915), .dout(n15000));
  jnot g14868(.din(n15000), .dout(n15001));
  jand g14869(.dina(n12569), .dinb(n5693), .dout(n15002));
  jand g14870(.dina(n11950), .dinb(n6209), .dout(n15003));
  jand g14871(.dina(n11952), .dinb(n6131), .dout(n15004));
  jand g14872(.dina(n11954), .dinb(n5691), .dout(n15005));
  jor  g14873(.dina(n15005), .dinb(n15004), .dout(n15006));
  jor  g14874(.dina(n15006), .dinb(n15003), .dout(n15007));
  jor  g14875(.dina(n15007), .dinb(n15002), .dout(n15008));
  jxor g14876(.dina(n15008), .dinb(n4247), .dout(n15009));
  jor  g14877(.dina(n15009), .dinb(n15001), .dout(n15010));
  jand g14878(.dina(n14184), .dinb(n4449), .dout(n15011));
  jand g14879(.dina(n11976), .dinb(n4453), .dout(n15012));
  jand g14880(.dina(n11978), .dinb(n4457), .dout(n15013));
  jand g14881(.dina(n11980), .dinb(n4461), .dout(n15014));
  jor  g14882(.dina(n15014), .dinb(n15013), .dout(n15015));
  jor  g14883(.dina(n15015), .dinb(n15012), .dout(n15016));
  jor  g14884(.dina(n15016), .dinb(n15011), .dout(n15017));
  jxor g14885(.dina(n15017), .dinb(n88), .dout(n15018));
  jnot g14886(.din(n15018), .dout(n15019));
  jxor g14887(.dina(n14582), .dinb(n14581), .dout(n15020));
  jand g14888(.dina(n15020), .dinb(n15019), .dout(n15021));
  jand g14889(.dina(n14194), .dinb(n4449), .dout(n15022));
  jand g14890(.dina(n11978), .dinb(n4453), .dout(n15023));
  jand g14891(.dina(n11980), .dinb(n4457), .dout(n15024));
  jand g14892(.dina(n11982), .dinb(n4461), .dout(n15025));
  jor  g14893(.dina(n15025), .dinb(n15024), .dout(n15026));
  jor  g14894(.dina(n15026), .dinb(n15023), .dout(n15027));
  jor  g14895(.dina(n15027), .dinb(n15022), .dout(n15028));
  jxor g14896(.dina(n15028), .dinb(n88), .dout(n15029));
  jnot g14897(.din(n15029), .dout(n15030));
  jxor g14898(.dina(n14577), .dinb(n14576), .dout(n15031));
  jand g14899(.dina(n15031), .dinb(n15030), .dout(n15032));
  jand g14900(.dina(n13899), .dinb(n4449), .dout(n15033));
  jand g14901(.dina(n11980), .dinb(n4453), .dout(n15034));
  jand g14902(.dina(n11982), .dinb(n4457), .dout(n15035));
  jand g14903(.dina(n11985), .dinb(n4461), .dout(n15036));
  jor  g14904(.dina(n15036), .dinb(n15035), .dout(n15037));
  jor  g14905(.dina(n15037), .dinb(n15034), .dout(n15038));
  jor  g14906(.dina(n15038), .dinb(n15033), .dout(n15039));
  jxor g14907(.dina(n15039), .dinb(n88), .dout(n15040));
  jnot g14908(.din(n15040), .dout(n15041));
  jxor g14909(.dina(n14572), .dinb(n14571), .dout(n15042));
  jand g14910(.dina(n15042), .dinb(n15041), .dout(n15043));
  jor  g14911(.dina(n14221), .dinb(n4724), .dout(n15044));
  jnot g14912(.din(n11982), .dout(n15045));
  jor  g14913(.dina(n15045), .dinb(n4905), .dout(n15046));
  jor  g14914(.dina(n11984), .dinb(n4735), .dout(n15047));
  jor  g14915(.dina(n11987), .dinb(n4733), .dout(n15048));
  jand g14916(.dina(n15048), .dinb(n15047), .dout(n15049));
  jand g14917(.dina(n15049), .dinb(n15046), .dout(n15050));
  jand g14918(.dina(n15050), .dinb(n15044), .dout(n15051));
  jxor g14919(.dina(n15051), .dinb(\a[29] ), .dout(n15052));
  jnot g14920(.din(n15052), .dout(n15053));
  jxor g14921(.dina(n14567), .dinb(n14566), .dout(n15054));
  jand g14922(.dina(n15054), .dinb(n15053), .dout(n15055));
  jor  g14923(.dina(n14248), .dinb(n4724), .dout(n15056));
  jor  g14924(.dina(n11984), .dinb(n4905), .dout(n15057));
  jor  g14925(.dina(n11987), .dinb(n4735), .dout(n15058));
  jor  g14926(.dina(n11991), .dinb(n4733), .dout(n15059));
  jand g14927(.dina(n15059), .dinb(n15058), .dout(n15060));
  jand g14928(.dina(n15060), .dinb(n15057), .dout(n15061));
  jand g14929(.dina(n15061), .dinb(n15056), .dout(n15062));
  jxor g14930(.dina(n15062), .dinb(\a[29] ), .dout(n15063));
  jnot g14931(.din(n15063), .dout(n15064));
  jxor g14932(.dina(n14562), .dinb(n14561), .dout(n15065));
  jand g14933(.dina(n15065), .dinb(n15064), .dout(n15066));
  jor  g14934(.dina(n14271), .dinb(n4724), .dout(n15067));
  jor  g14935(.dina(n11987), .dinb(n4905), .dout(n15068));
  jor  g14936(.dina(n11991), .dinb(n4735), .dout(n15069));
  jor  g14937(.dina(n11995), .dinb(n4733), .dout(n15070));
  jand g14938(.dina(n15070), .dinb(n15069), .dout(n15071));
  jand g14939(.dina(n15071), .dinb(n15068), .dout(n15072));
  jand g14940(.dina(n15072), .dinb(n15067), .dout(n15073));
  jxor g14941(.dina(n15073), .dinb(\a[29] ), .dout(n15074));
  jnot g14942(.din(n15074), .dout(n15075));
  jxor g14943(.dina(n14557), .dinb(n14556), .dout(n15076));
  jand g14944(.dina(n15076), .dinb(n15075), .dout(n15077));
  jor  g14945(.dina(n14301), .dinb(n4724), .dout(n15078));
  jor  g14946(.dina(n11991), .dinb(n4905), .dout(n15079));
  jor  g14947(.dina(n11995), .dinb(n4735), .dout(n15080));
  jor  g14948(.dina(n11997), .dinb(n4733), .dout(n15081));
  jand g14949(.dina(n15081), .dinb(n15080), .dout(n15082));
  jand g14950(.dina(n15082), .dinb(n15079), .dout(n15083));
  jand g14951(.dina(n15083), .dinb(n15078), .dout(n15084));
  jxor g14952(.dina(n15084), .dinb(\a[29] ), .dout(n15085));
  jnot g14953(.din(n15085), .dout(n15086));
  jxor g14954(.dina(n14552), .dinb(n14551), .dout(n15087));
  jand g14955(.dina(n15087), .dinb(n15086), .dout(n15088));
  jor  g14956(.dina(n14353), .dinb(n4724), .dout(n15089));
  jor  g14957(.dina(n11995), .dinb(n4905), .dout(n15090));
  jor  g14958(.dina(n11997), .dinb(n4735), .dout(n15091));
  jor  g14959(.dina(n11999), .dinb(n4733), .dout(n15092));
  jand g14960(.dina(n15092), .dinb(n15091), .dout(n15093));
  jand g14961(.dina(n15093), .dinb(n15090), .dout(n15094));
  jand g14962(.dina(n15094), .dinb(n15089), .dout(n15095));
  jxor g14963(.dina(n15095), .dinb(\a[29] ), .dout(n15096));
  jnot g14964(.din(n15096), .dout(n15097));
  jxor g14965(.dina(n14549), .dinb(n14548), .dout(n15098));
  jand g14966(.dina(n15098), .dinb(n15097), .dout(n15099));
  jor  g14967(.dina(n14390), .dinb(n4724), .dout(n15100));
  jor  g14968(.dina(n11997), .dinb(n4905), .dout(n15101));
  jor  g14969(.dina(n11999), .dinb(n4735), .dout(n15102));
  jor  g14970(.dina(n12001), .dinb(n4733), .dout(n15103));
  jand g14971(.dina(n15103), .dinb(n15102), .dout(n15104));
  jand g14972(.dina(n15104), .dinb(n15101), .dout(n15105));
  jand g14973(.dina(n15105), .dinb(n15100), .dout(n15106));
  jxor g14974(.dina(n15106), .dinb(\a[29] ), .dout(n15107));
  jnot g14975(.din(n15107), .dout(n15108));
  jxor g14976(.dina(n14544), .dinb(n14535), .dout(n15109));
  jand g14977(.dina(n15109), .dinb(n15108), .dout(n15110));
  jor  g14978(.dina(n14432), .dinb(n4724), .dout(n15111));
  jor  g14979(.dina(n11999), .dinb(n4905), .dout(n15112));
  jor  g14980(.dina(n12001), .dinb(n4735), .dout(n15113));
  jor  g14981(.dina(n12004), .dinb(n4733), .dout(n15114));
  jand g14982(.dina(n15114), .dinb(n15113), .dout(n15115));
  jand g14983(.dina(n15115), .dinb(n15112), .dout(n15116));
  jand g14984(.dina(n15116), .dinb(n15111), .dout(n15117));
  jxor g14985(.dina(n15117), .dinb(\a[29] ), .dout(n15118));
  jnot g14986(.din(n15118), .dout(n15119));
  jxor g14987(.dina(n14502), .dinb(n14496), .dout(n15120));
  jand g14988(.dina(n15120), .dinb(n15119), .dout(n15121));
  jand g14989(.dina(n12010), .dinb(n731), .dout(n15122));
  jand g14990(.dina(n14497), .dinb(n4449), .dout(n15123));
  jand g14991(.dina(n12010), .dinb(n4457), .dout(n15124));
  jand g14992(.dina(n12008), .dinb(n4453), .dout(n15125));
  jor  g14993(.dina(n15125), .dinb(n15124), .dout(n15126));
  jor  g14994(.dina(n15126), .dinb(n15123), .dout(n15127));
  jnot g14995(.din(n15127), .dout(n15128));
  jand g14996(.dina(n12010), .dinb(n4447), .dout(n15129));
  jnot g14997(.din(n15129), .dout(n15130));
  jand g14998(.dina(n15130), .dinb(\a[29] ), .dout(n15131));
  jand g14999(.dina(n15131), .dinb(n15128), .dout(n15132));
  jand g15000(.dina(n14537), .dinb(n4449), .dout(n15133));
  jand g15001(.dina(n12006), .dinb(n4453), .dout(n15134));
  jand g15002(.dina(n12008), .dinb(n4457), .dout(n15135));
  jand g15003(.dina(n12010), .dinb(n4461), .dout(n15136));
  jor  g15004(.dina(n15136), .dinb(n15135), .dout(n15137));
  jor  g15005(.dina(n15137), .dinb(n15134), .dout(n15138));
  jor  g15006(.dina(n15138), .dinb(n15133), .dout(n15139));
  jnot g15007(.din(n15139), .dout(n15140));
  jand g15008(.dina(n15140), .dinb(n15132), .dout(n15141));
  jand g15009(.dina(n15141), .dinb(n15122), .dout(n15142));
  jxor g15010(.dina(n12004), .dinb(n12001), .dout(n15143));
  jxor g15011(.dina(n12013), .dinb(n15143), .dout(n15144));
  jor  g15012(.dina(n15144), .dinb(n4724), .dout(n15145));
  jor  g15013(.dina(n12001), .dinb(n4905), .dout(n15146));
  jor  g15014(.dina(n12004), .dinb(n4735), .dout(n15147));
  jor  g15015(.dina(n12009), .dinb(n4733), .dout(n15148));
  jand g15016(.dina(n15148), .dinb(n15147), .dout(n15149));
  jand g15017(.dina(n15149), .dinb(n15146), .dout(n15150));
  jand g15018(.dina(n15150), .dinb(n15145), .dout(n15151));
  jxor g15019(.dina(n15151), .dinb(\a[29] ), .dout(n15152));
  jnot g15020(.din(n15152), .dout(n15153));
  jxor g15021(.dina(n15141), .dinb(n15122), .dout(n15154));
  jand g15022(.dina(n15154), .dinb(n15153), .dout(n15155));
  jor  g15023(.dina(n15155), .dinb(n15142), .dout(n15156));
  jxor g15024(.dina(n15120), .dinb(n15119), .dout(n15157));
  jand g15025(.dina(n15157), .dinb(n15156), .dout(n15158));
  jor  g15026(.dina(n15158), .dinb(n15121), .dout(n15159));
  jxor g15027(.dina(n15109), .dinb(n15108), .dout(n15160));
  jand g15028(.dina(n15160), .dinb(n15159), .dout(n15161));
  jor  g15029(.dina(n15161), .dinb(n15110), .dout(n15162));
  jxor g15030(.dina(n15098), .dinb(n15097), .dout(n15163));
  jand g15031(.dina(n15163), .dinb(n15162), .dout(n15164));
  jor  g15032(.dina(n15164), .dinb(n15099), .dout(n15165));
  jxor g15033(.dina(n15087), .dinb(n15086), .dout(n15166));
  jand g15034(.dina(n15166), .dinb(n15165), .dout(n15167));
  jor  g15035(.dina(n15167), .dinb(n15088), .dout(n15168));
  jxor g15036(.dina(n15076), .dinb(n15075), .dout(n15169));
  jand g15037(.dina(n15169), .dinb(n15168), .dout(n15170));
  jor  g15038(.dina(n15170), .dinb(n15077), .dout(n15171));
  jxor g15039(.dina(n15065), .dinb(n15064), .dout(n15172));
  jand g15040(.dina(n15172), .dinb(n15171), .dout(n15173));
  jor  g15041(.dina(n15173), .dinb(n15066), .dout(n15174));
  jxor g15042(.dina(n15054), .dinb(n15053), .dout(n15175));
  jand g15043(.dina(n15175), .dinb(n15174), .dout(n15176));
  jor  g15044(.dina(n15176), .dinb(n15055), .dout(n15177));
  jxor g15045(.dina(n15042), .dinb(n15041), .dout(n15178));
  jand g15046(.dina(n15178), .dinb(n15177), .dout(n15179));
  jor  g15047(.dina(n15179), .dinb(n15043), .dout(n15180));
  jxor g15048(.dina(n15031), .dinb(n15030), .dout(n15181));
  jand g15049(.dina(n15181), .dinb(n15180), .dout(n15182));
  jor  g15050(.dina(n15182), .dinb(n15032), .dout(n15183));
  jxor g15051(.dina(n15020), .dinb(n15019), .dout(n15184));
  jand g15052(.dina(n15184), .dinb(n15183), .dout(n15185));
  jor  g15053(.dina(n15185), .dinb(n15021), .dout(n15186));
  jxor g15054(.dina(n14599), .dinb(n14591), .dout(n15187));
  jand g15055(.dina(n15187), .dinb(n15186), .dout(n15188));
  jnot g15056(.din(n15188), .dout(n15189));
  jxor g15057(.dina(n15187), .dinb(n15186), .dout(n15190));
  jnot g15058(.din(n15190), .dout(n15191));
  jand g15059(.dina(n13682), .dinb(n75), .dout(n15192));
  jand g15060(.dina(n11968), .dinb(n4933), .dout(n15193));
  jand g15061(.dina(n11970), .dinb(n4918), .dout(n15194));
  jand g15062(.dina(n11972), .dinb(n4745), .dout(n15195));
  jor  g15063(.dina(n15195), .dinb(n15194), .dout(n15196));
  jor  g15064(.dina(n15196), .dinb(n15193), .dout(n15197));
  jor  g15065(.dina(n15197), .dinb(n15192), .dout(n15198));
  jxor g15066(.dina(n15198), .dinb(n68), .dout(n15199));
  jor  g15067(.dina(n15199), .dinb(n15191), .dout(n15200));
  jand g15068(.dina(n15200), .dinb(n15189), .dout(n15201));
  jnot g15069(.din(n15201), .dout(n15202));
  jxor g15070(.dina(n14895), .dinb(n14894), .dout(n15203));
  jand g15071(.dina(n15203), .dinb(n15202), .dout(n15204));
  jnot g15072(.din(n15204), .dout(n15205));
  jxor g15073(.dina(n15203), .dinb(n15202), .dout(n15206));
  jnot g15074(.din(n15206), .dout(n15207));
  jand g15075(.dina(n13116), .dinb(n5365), .dout(n15208));
  jand g15076(.dina(n11960), .dinb(n5500), .dout(n15209));
  jand g15077(.dina(n11962), .dinb(n5424), .dout(n15210));
  jand g15078(.dina(n11964), .dinb(n5363), .dout(n15211));
  jor  g15079(.dina(n15211), .dinb(n15210), .dout(n15212));
  jor  g15080(.dina(n15212), .dinb(n15209), .dout(n15213));
  jor  g15081(.dina(n15213), .dinb(n15208), .dout(n15214));
  jxor g15082(.dina(n15214), .dinb(n72), .dout(n15215));
  jor  g15083(.dina(n15215), .dinb(n15207), .dout(n15216));
  jand g15084(.dina(n15216), .dinb(n15205), .dout(n15217));
  jnot g15085(.din(n15217), .dout(n15218));
  jxor g15086(.dina(n14912), .dinb(n14904), .dout(n15219));
  jand g15087(.dina(n15219), .dinb(n15218), .dout(n15220));
  jnot g15088(.din(n15220), .dout(n15221));
  jxor g15089(.dina(n15219), .dinb(n15218), .dout(n15222));
  jnot g15090(.din(n15222), .dout(n15223));
  jand g15091(.dina(n12510), .dinb(n5693), .dout(n15224));
  jand g15092(.dina(n11952), .dinb(n6209), .dout(n15225));
  jand g15093(.dina(n11954), .dinb(n6131), .dout(n15226));
  jand g15094(.dina(n11956), .dinb(n5691), .dout(n15227));
  jor  g15095(.dina(n15227), .dinb(n15226), .dout(n15228));
  jor  g15096(.dina(n15228), .dinb(n15225), .dout(n15229));
  jor  g15097(.dina(n15229), .dinb(n15224), .dout(n15230));
  jxor g15098(.dina(n15230), .dinb(n4247), .dout(n15231));
  jor  g15099(.dina(n15231), .dinb(n15223), .dout(n15232));
  jand g15100(.dina(n15232), .dinb(n15221), .dout(n15233));
  jnot g15101(.din(n15233), .dout(n15234));
  jxor g15102(.dina(n15009), .dinb(n15001), .dout(n15235));
  jand g15103(.dina(n15235), .dinb(n15234), .dout(n15236));
  jnot g15104(.din(n15236), .dout(n15237));
  jand g15105(.dina(n15237), .dinb(n15010), .dout(n15238));
  jnot g15106(.din(n15238), .dout(n15239));
  jxor g15107(.dina(n14933), .dinb(n14925), .dout(n15240));
  jand g15108(.dina(n15240), .dinb(n15239), .dout(n15241));
  jnot g15109(.din(n15241), .dout(n15242));
  jxor g15110(.dina(n15240), .dinb(n15239), .dout(n15243));
  jnot g15111(.din(n15243), .dout(n15244));
  jand g15112(.dina(n12751), .dinb(n6340), .dout(n15245));
  jand g15113(.dina(n11942), .dinb(n6798), .dout(n15246));
  jand g15114(.dina(n11944), .dinb(n6556), .dout(n15247));
  jand g15115(.dina(n11946), .dinb(n6338), .dout(n15248));
  jor  g15116(.dina(n15248), .dinb(n15247), .dout(n15249));
  jor  g15117(.dina(n15249), .dinb(n15246), .dout(n15250));
  jor  g15118(.dina(n15250), .dinb(n15245), .dout(n15251));
  jxor g15119(.dina(n15251), .dinb(n5064), .dout(n15252));
  jor  g15120(.dina(n15252), .dinb(n15244), .dout(n15253));
  jand g15121(.dina(n15253), .dinb(n15242), .dout(n15254));
  jnot g15122(.din(n15254), .dout(n15255));
  jxor g15123(.dina(n14949), .dinb(n14941), .dout(n15256));
  jand g15124(.dina(n15256), .dinb(n15255), .dout(n15257));
  jnot g15125(.din(n15257), .dout(n15258));
  jxor g15126(.dina(n15256), .dinb(n15255), .dout(n15259));
  jnot g15127(.din(n15259), .dout(n15260));
  jand g15128(.dina(n12841), .dinb(n6936), .dout(n15261));
  jand g15129(.dina(n12783), .dinb(n7741), .dout(n15262));
  jand g15130(.dina(n12766), .dinb(n7613), .dout(n15263));
  jand g15131(.dina(n12177), .dinb(n6934), .dout(n15264));
  jor  g15132(.dina(n15264), .dinb(n15263), .dout(n15265));
  jor  g15133(.dina(n15265), .dinb(n15262), .dout(n15266));
  jor  g15134(.dina(n15266), .dinb(n15261), .dout(n15267));
  jxor g15135(.dina(n15267), .dinb(n5292), .dout(n15268));
  jor  g15136(.dina(n15268), .dinb(n15260), .dout(n15269));
  jand g15137(.dina(n15269), .dinb(n15258), .dout(n15270));
  jnot g15138(.din(n15270), .dout(n15271));
  jxor g15139(.dina(n14998), .dinb(n14990), .dout(n15272));
  jand g15140(.dina(n15272), .dinb(n15271), .dout(n15273));
  jnot g15141(.din(n15273), .dout(n15274));
  jand g15142(.dina(n15274), .dinb(n14999), .dout(n15275));
  jnot g15143(.din(n15275), .dout(n15276));
  jxor g15144(.dina(n14970), .dinb(n14962), .dout(n15277));
  jand g15145(.dina(n15277), .dinb(n15276), .dout(n15278));
  jnot g15146(.din(n15278), .dout(n15279));
  jxor g15147(.dina(n15277), .dinb(n15276), .dout(n15280));
  jnot g15148(.din(n15280), .dout(n15281));
  jor  g15149(.dina(n12814), .dinb(n7889), .dout(n15283));
  jand g15150(.dina(n14975), .dinb(n15283), .dout(n15287));
  jand g15151(.dina(n15287), .dinb(n7891), .dout(n15288));
  jxor g15152(.dina(n15288), .dinb(\a[11] ), .dout(n15289));
  jor  g15153(.dina(n15289), .dinb(n15281), .dout(n15290));
  jand g15154(.dina(n15290), .dinb(n15279), .dout(n15291));
  jnot g15155(.din(n15291), .dout(n15292));
  jxor g15156(.dina(n14982), .dinb(n14981), .dout(n15293));
  jand g15157(.dina(n15293), .dinb(n15292), .dout(n15294));
  jxor g15158(.dina(n15293), .dinb(n15292), .dout(n15295));
  jxor g15159(.dina(n15235), .dinb(n15234), .dout(n15296));
  jnot g15160(.din(n15296), .dout(n15297));
  jand g15161(.dina(n12189), .dinb(n6340), .dout(n15298));
  jand g15162(.dina(n11944), .dinb(n6798), .dout(n15299));
  jand g15163(.dina(n11946), .dinb(n6556), .dout(n15300));
  jand g15164(.dina(n11948), .dinb(n6338), .dout(n15301));
  jor  g15165(.dina(n15301), .dinb(n15300), .dout(n15302));
  jor  g15166(.dina(n15302), .dinb(n15299), .dout(n15303));
  jor  g15167(.dina(n15303), .dinb(n15298), .dout(n15304));
  jxor g15168(.dina(n15304), .dinb(n5064), .dout(n15305));
  jor  g15169(.dina(n15305), .dinb(n15297), .dout(n15306));
  jxor g15170(.dina(n15184), .dinb(n15183), .dout(n15307));
  jnot g15171(.din(n15307), .dout(n15308));
  jand g15172(.dina(n13806), .dinb(n75), .dout(n15309));
  jand g15173(.dina(n11970), .dinb(n4933), .dout(n15310));
  jand g15174(.dina(n11972), .dinb(n4918), .dout(n15311));
  jand g15175(.dina(n11974), .dinb(n4745), .dout(n15312));
  jor  g15176(.dina(n15312), .dinb(n15311), .dout(n15313));
  jor  g15177(.dina(n15313), .dinb(n15310), .dout(n15314));
  jor  g15178(.dina(n15314), .dinb(n15309), .dout(n15315));
  jxor g15179(.dina(n15315), .dinb(n68), .dout(n15316));
  jor  g15180(.dina(n15316), .dinb(n15308), .dout(n15317));
  jxor g15181(.dina(n15181), .dinb(n15180), .dout(n15318));
  jnot g15182(.din(n15318), .dout(n15319));
  jand g15183(.dina(n13664), .dinb(n75), .dout(n15320));
  jand g15184(.dina(n11972), .dinb(n4933), .dout(n15321));
  jand g15185(.dina(n11974), .dinb(n4918), .dout(n15322));
  jand g15186(.dina(n11976), .dinb(n4745), .dout(n15323));
  jor  g15187(.dina(n15323), .dinb(n15322), .dout(n15324));
  jor  g15188(.dina(n15324), .dinb(n15321), .dout(n15325));
  jor  g15189(.dina(n15325), .dinb(n15320), .dout(n15326));
  jxor g15190(.dina(n15326), .dinb(n68), .dout(n15327));
  jor  g15191(.dina(n15327), .dinb(n15319), .dout(n15328));
  jxor g15192(.dina(n15178), .dinb(n15177), .dout(n15329));
  jnot g15193(.din(n15329), .dout(n15330));
  jand g15194(.dina(n13924), .dinb(n75), .dout(n15331));
  jand g15195(.dina(n11974), .dinb(n4933), .dout(n15332));
  jand g15196(.dina(n11976), .dinb(n4918), .dout(n15333));
  jand g15197(.dina(n11978), .dinb(n4745), .dout(n15334));
  jor  g15198(.dina(n15334), .dinb(n15333), .dout(n15335));
  jor  g15199(.dina(n15335), .dinb(n15332), .dout(n15336));
  jor  g15200(.dina(n15336), .dinb(n15331), .dout(n15337));
  jxor g15201(.dina(n15337), .dinb(n68), .dout(n15338));
  jor  g15202(.dina(n15338), .dinb(n15330), .dout(n15339));
  jxor g15203(.dina(n15175), .dinb(n15174), .dout(n15340));
  jnot g15204(.din(n15340), .dout(n15341));
  jand g15205(.dina(n14184), .dinb(n75), .dout(n15342));
  jand g15206(.dina(n11976), .dinb(n4933), .dout(n15343));
  jand g15207(.dina(n11978), .dinb(n4918), .dout(n15344));
  jand g15208(.dina(n11980), .dinb(n4745), .dout(n15345));
  jor  g15209(.dina(n15345), .dinb(n15344), .dout(n15346));
  jor  g15210(.dina(n15346), .dinb(n15343), .dout(n15347));
  jor  g15211(.dina(n15347), .dinb(n15342), .dout(n15348));
  jxor g15212(.dina(n15348), .dinb(n68), .dout(n15349));
  jor  g15213(.dina(n15349), .dinb(n15341), .dout(n15350));
  jxor g15214(.dina(n15172), .dinb(n15171), .dout(n15351));
  jnot g15215(.din(n15351), .dout(n15352));
  jand g15216(.dina(n14194), .dinb(n75), .dout(n15353));
  jand g15217(.dina(n11978), .dinb(n4933), .dout(n15354));
  jand g15218(.dina(n11980), .dinb(n4918), .dout(n15355));
  jand g15219(.dina(n11982), .dinb(n4745), .dout(n15356));
  jor  g15220(.dina(n15356), .dinb(n15355), .dout(n15357));
  jor  g15221(.dina(n15357), .dinb(n15354), .dout(n15358));
  jor  g15222(.dina(n15358), .dinb(n15353), .dout(n15359));
  jxor g15223(.dina(n15359), .dinb(n68), .dout(n15360));
  jor  g15224(.dina(n15360), .dinb(n15352), .dout(n15361));
  jxor g15225(.dina(n15169), .dinb(n15168), .dout(n15362));
  jnot g15226(.din(n15362), .dout(n15363));
  jand g15227(.dina(n13899), .dinb(n75), .dout(n15364));
  jand g15228(.dina(n11980), .dinb(n4933), .dout(n15365));
  jand g15229(.dina(n11982), .dinb(n4918), .dout(n15366));
  jand g15230(.dina(n11985), .dinb(n4745), .dout(n15367));
  jor  g15231(.dina(n15367), .dinb(n15366), .dout(n15368));
  jor  g15232(.dina(n15368), .dinb(n15365), .dout(n15369));
  jor  g15233(.dina(n15369), .dinb(n15364), .dout(n15370));
  jxor g15234(.dina(n15370), .dinb(n68), .dout(n15371));
  jor  g15235(.dina(n15371), .dinb(n15363), .dout(n15372));
  jxor g15236(.dina(n15166), .dinb(n15165), .dout(n15373));
  jnot g15237(.din(n15373), .dout(n15374));
  jor  g15238(.dina(n14221), .dinb(n4747), .dout(n15375));
  jor  g15239(.dina(n15045), .dinb(n4959), .dout(n15376));
  jor  g15240(.dina(n11984), .dinb(n4919), .dout(n15377));
  jor  g15241(.dina(n11987), .dinb(n4746), .dout(n15378));
  jand g15242(.dina(n15378), .dinb(n15377), .dout(n15379));
  jand g15243(.dina(n15379), .dinb(n15376), .dout(n15380));
  jand g15244(.dina(n15380), .dinb(n15375), .dout(n15381));
  jxor g15245(.dina(n15381), .dinb(\a[26] ), .dout(n15382));
  jor  g15246(.dina(n15382), .dinb(n15374), .dout(n15383));
  jxor g15247(.dina(n15163), .dinb(n15162), .dout(n15384));
  jnot g15248(.din(n15384), .dout(n15385));
  jor  g15249(.dina(n14248), .dinb(n4747), .dout(n15386));
  jor  g15250(.dina(n11984), .dinb(n4959), .dout(n15387));
  jor  g15251(.dina(n11987), .dinb(n4919), .dout(n15388));
  jor  g15252(.dina(n11991), .dinb(n4746), .dout(n15389));
  jand g15253(.dina(n15389), .dinb(n15388), .dout(n15390));
  jand g15254(.dina(n15390), .dinb(n15387), .dout(n15391));
  jand g15255(.dina(n15391), .dinb(n15386), .dout(n15392));
  jxor g15256(.dina(n15392), .dinb(\a[26] ), .dout(n15393));
  jor  g15257(.dina(n15393), .dinb(n15385), .dout(n15394));
  jxor g15258(.dina(n15160), .dinb(n15159), .dout(n15395));
  jnot g15259(.din(n15395), .dout(n15396));
  jor  g15260(.dina(n14271), .dinb(n4747), .dout(n15397));
  jor  g15261(.dina(n11987), .dinb(n4959), .dout(n15398));
  jor  g15262(.dina(n11995), .dinb(n4746), .dout(n15399));
  jor  g15263(.dina(n11991), .dinb(n4919), .dout(n15400));
  jand g15264(.dina(n15400), .dinb(n15399), .dout(n15401));
  jand g15265(.dina(n15401), .dinb(n15398), .dout(n15402));
  jand g15266(.dina(n15402), .dinb(n15397), .dout(n15403));
  jxor g15267(.dina(n15403), .dinb(\a[26] ), .dout(n15404));
  jor  g15268(.dina(n15404), .dinb(n15396), .dout(n15405));
  jor  g15269(.dina(n14301), .dinb(n4747), .dout(n15406));
  jor  g15270(.dina(n11991), .dinb(n4959), .dout(n15407));
  jor  g15271(.dina(n11995), .dinb(n4919), .dout(n15408));
  jor  g15272(.dina(n11997), .dinb(n4746), .dout(n15409));
  jand g15273(.dina(n15409), .dinb(n15408), .dout(n15410));
  jand g15274(.dina(n15410), .dinb(n15407), .dout(n15411));
  jand g15275(.dina(n15411), .dinb(n15406), .dout(n15412));
  jxor g15276(.dina(n15412), .dinb(\a[26] ), .dout(n15413));
  jnot g15277(.din(n15413), .dout(n15414));
  jxor g15278(.dina(n15157), .dinb(n15156), .dout(n15415));
  jand g15279(.dina(n15415), .dinb(n15414), .dout(n15416));
  jor  g15280(.dina(n14353), .dinb(n4747), .dout(n15417));
  jor  g15281(.dina(n11995), .dinb(n4959), .dout(n15418));
  jor  g15282(.dina(n11999), .dinb(n4746), .dout(n15419));
  jor  g15283(.dina(n11997), .dinb(n4919), .dout(n15420));
  jand g15284(.dina(n15420), .dinb(n15419), .dout(n15421));
  jand g15285(.dina(n15421), .dinb(n15418), .dout(n15422));
  jand g15286(.dina(n15422), .dinb(n15417), .dout(n15423));
  jxor g15287(.dina(n15423), .dinb(\a[26] ), .dout(n15424));
  jnot g15288(.din(n15424), .dout(n15425));
  jxor g15289(.dina(n15154), .dinb(n15153), .dout(n15426));
  jand g15290(.dina(n15426), .dinb(n15425), .dout(n15427));
  jor  g15291(.dina(n14390), .dinb(n4747), .dout(n15428));
  jor  g15292(.dina(n11997), .dinb(n4959), .dout(n15429));
  jor  g15293(.dina(n11999), .dinb(n4919), .dout(n15430));
  jor  g15294(.dina(n12001), .dinb(n4746), .dout(n15431));
  jand g15295(.dina(n15431), .dinb(n15430), .dout(n15432));
  jand g15296(.dina(n15432), .dinb(n15429), .dout(n15433));
  jand g15297(.dina(n15433), .dinb(n15428), .dout(n15434));
  jxor g15298(.dina(n15434), .dinb(\a[26] ), .dout(n15435));
  jnot g15299(.din(n15435), .dout(n15436));
  jor  g15300(.dina(n15132), .dinb(n88), .dout(n15437));
  jxor g15301(.dina(n15437), .dinb(n15140), .dout(n15438));
  jand g15302(.dina(n15438), .dinb(n15436), .dout(n15439));
  jor  g15303(.dina(n14432), .dinb(n4747), .dout(n15440));
  jor  g15304(.dina(n11999), .dinb(n4959), .dout(n15441));
  jor  g15305(.dina(n12001), .dinb(n4919), .dout(n15442));
  jor  g15306(.dina(n12004), .dinb(n4746), .dout(n15443));
  jand g15307(.dina(n15443), .dinb(n15442), .dout(n15444));
  jand g15308(.dina(n15444), .dinb(n15441), .dout(n15445));
  jand g15309(.dina(n15445), .dinb(n15440), .dout(n15446));
  jxor g15310(.dina(n15446), .dinb(\a[26] ), .dout(n15447));
  jnot g15311(.din(n15447), .dout(n15448));
  jand g15312(.dina(n15129), .dinb(\a[29] ), .dout(n15449));
  jxor g15313(.dina(n15449), .dinb(n15127), .dout(n15450));
  jand g15314(.dina(n15450), .dinb(n15448), .dout(n15451));
  jand g15315(.dina(n14497), .dinb(n75), .dout(n15452));
  jand g15316(.dina(n12008), .dinb(n4933), .dout(n15453));
  jand g15317(.dina(n12010), .dinb(n4918), .dout(n15454));
  jor  g15318(.dina(n15454), .dinb(n15453), .dout(n15455));
  jor  g15319(.dina(n15455), .dinb(n15452), .dout(n15456));
  jnot g15320(.din(n15456), .dout(n15457));
  jand g15321(.dina(n12010), .dinb(n74), .dout(n15458));
  jnot g15322(.din(n15458), .dout(n15459));
  jand g15323(.dina(n15459), .dinb(\a[26] ), .dout(n15460));
  jand g15324(.dina(n15460), .dinb(n15457), .dout(n15461));
  jand g15325(.dina(n14537), .dinb(n75), .dout(n15462));
  jand g15326(.dina(n12006), .dinb(n4933), .dout(n15463));
  jand g15327(.dina(n12008), .dinb(n4918), .dout(n15464));
  jand g15328(.dina(n12010), .dinb(n4745), .dout(n15465));
  jor  g15329(.dina(n15465), .dinb(n15464), .dout(n15466));
  jor  g15330(.dina(n15466), .dinb(n15463), .dout(n15467));
  jor  g15331(.dina(n15467), .dinb(n15462), .dout(n15468));
  jnot g15332(.din(n15468), .dout(n15469));
  jand g15333(.dina(n15469), .dinb(n15461), .dout(n15470));
  jand g15334(.dina(n15470), .dinb(n15129), .dout(n15471));
  jor  g15335(.dina(n15144), .dinb(n4747), .dout(n15472));
  jor  g15336(.dina(n12001), .dinb(n4959), .dout(n15473));
  jor  g15337(.dina(n12004), .dinb(n4919), .dout(n15474));
  jor  g15338(.dina(n12009), .dinb(n4746), .dout(n15475));
  jand g15339(.dina(n15475), .dinb(n15474), .dout(n15476));
  jand g15340(.dina(n15476), .dinb(n15473), .dout(n15477));
  jand g15341(.dina(n15477), .dinb(n15472), .dout(n15478));
  jxor g15342(.dina(n15478), .dinb(\a[26] ), .dout(n15479));
  jnot g15343(.din(n15479), .dout(n15480));
  jxor g15344(.dina(n15470), .dinb(n15129), .dout(n15481));
  jand g15345(.dina(n15481), .dinb(n15480), .dout(n15482));
  jor  g15346(.dina(n15482), .dinb(n15471), .dout(n15483));
  jxor g15347(.dina(n15450), .dinb(n15448), .dout(n15484));
  jand g15348(.dina(n15484), .dinb(n15483), .dout(n15485));
  jor  g15349(.dina(n15485), .dinb(n15451), .dout(n15486));
  jxor g15350(.dina(n15438), .dinb(n15436), .dout(n15487));
  jand g15351(.dina(n15487), .dinb(n15486), .dout(n15488));
  jor  g15352(.dina(n15488), .dinb(n15439), .dout(n15489));
  jxor g15353(.dina(n15426), .dinb(n15425), .dout(n15490));
  jand g15354(.dina(n15490), .dinb(n15489), .dout(n15491));
  jor  g15355(.dina(n15491), .dinb(n15427), .dout(n15492));
  jxor g15356(.dina(n15415), .dinb(n15414), .dout(n15493));
  jand g15357(.dina(n15493), .dinb(n15492), .dout(n15494));
  jor  g15358(.dina(n15494), .dinb(n15416), .dout(n15495));
  jxor g15359(.dina(n15404), .dinb(n15396), .dout(n15496));
  jand g15360(.dina(n15496), .dinb(n15495), .dout(n15497));
  jnot g15361(.din(n15497), .dout(n15498));
  jand g15362(.dina(n15498), .dinb(n15405), .dout(n15499));
  jnot g15363(.din(n15499), .dout(n15500));
  jxor g15364(.dina(n15393), .dinb(n15385), .dout(n15501));
  jand g15365(.dina(n15501), .dinb(n15500), .dout(n15502));
  jnot g15366(.din(n15502), .dout(n15503));
  jand g15367(.dina(n15503), .dinb(n15394), .dout(n15504));
  jnot g15368(.din(n15504), .dout(n15505));
  jxor g15369(.dina(n15382), .dinb(n15374), .dout(n15506));
  jand g15370(.dina(n15506), .dinb(n15505), .dout(n15507));
  jnot g15371(.din(n15507), .dout(n15508));
  jand g15372(.dina(n15508), .dinb(n15383), .dout(n15509));
  jnot g15373(.din(n15509), .dout(n15510));
  jxor g15374(.dina(n15371), .dinb(n15363), .dout(n15511));
  jand g15375(.dina(n15511), .dinb(n15510), .dout(n15512));
  jnot g15376(.din(n15512), .dout(n15513));
  jand g15377(.dina(n15513), .dinb(n15372), .dout(n15514));
  jnot g15378(.din(n15514), .dout(n15515));
  jxor g15379(.dina(n15360), .dinb(n15352), .dout(n15516));
  jand g15380(.dina(n15516), .dinb(n15515), .dout(n15517));
  jnot g15381(.din(n15517), .dout(n15518));
  jand g15382(.dina(n15518), .dinb(n15361), .dout(n15519));
  jnot g15383(.din(n15519), .dout(n15520));
  jxor g15384(.dina(n15349), .dinb(n15341), .dout(n15521));
  jand g15385(.dina(n15521), .dinb(n15520), .dout(n15522));
  jnot g15386(.din(n15522), .dout(n15523));
  jand g15387(.dina(n15523), .dinb(n15350), .dout(n15524));
  jnot g15388(.din(n15524), .dout(n15525));
  jxor g15389(.dina(n15338), .dinb(n15330), .dout(n15526));
  jand g15390(.dina(n15526), .dinb(n15525), .dout(n15527));
  jnot g15391(.din(n15527), .dout(n15528));
  jand g15392(.dina(n15528), .dinb(n15339), .dout(n15529));
  jnot g15393(.din(n15529), .dout(n15530));
  jxor g15394(.dina(n15327), .dinb(n15319), .dout(n15531));
  jand g15395(.dina(n15531), .dinb(n15530), .dout(n15532));
  jnot g15396(.din(n15532), .dout(n15533));
  jand g15397(.dina(n15533), .dinb(n15328), .dout(n15534));
  jnot g15398(.din(n15534), .dout(n15535));
  jxor g15399(.dina(n15316), .dinb(n15308), .dout(n15536));
  jand g15400(.dina(n15536), .dinb(n15535), .dout(n15537));
  jnot g15401(.din(n15537), .dout(n15538));
  jand g15402(.dina(n15538), .dinb(n15317), .dout(n15539));
  jnot g15403(.din(n15539), .dout(n15540));
  jxor g15404(.dina(n15199), .dinb(n15191), .dout(n15541));
  jand g15405(.dina(n15541), .dinb(n15540), .dout(n15542));
  jnot g15406(.din(n15542), .dout(n15543));
  jxor g15407(.dina(n15541), .dinb(n15540), .dout(n15544));
  jnot g15408(.din(n15544), .dout(n15545));
  jand g15409(.dina(n13134), .dinb(n5365), .dout(n15546));
  jand g15410(.dina(n11962), .dinb(n5500), .dout(n15547));
  jand g15411(.dina(n11964), .dinb(n5424), .dout(n15548));
  jand g15412(.dina(n11966), .dinb(n5363), .dout(n15549));
  jor  g15413(.dina(n15549), .dinb(n15548), .dout(n15550));
  jor  g15414(.dina(n15550), .dinb(n15547), .dout(n15551));
  jor  g15415(.dina(n15551), .dinb(n15546), .dout(n15552));
  jxor g15416(.dina(n15552), .dinb(n72), .dout(n15553));
  jor  g15417(.dina(n15553), .dinb(n15545), .dout(n15554));
  jand g15418(.dina(n15554), .dinb(n15543), .dout(n15555));
  jnot g15419(.din(n15555), .dout(n15556));
  jxor g15420(.dina(n15215), .dinb(n15207), .dout(n15557));
  jand g15421(.dina(n15557), .dinb(n15556), .dout(n15558));
  jnot g15422(.din(n15558), .dout(n15559));
  jxor g15423(.dina(n15557), .dinb(n15556), .dout(n15560));
  jnot g15424(.din(n15560), .dout(n15561));
  jand g15425(.dina(n12472), .dinb(n5693), .dout(n15562));
  jand g15426(.dina(n11954), .dinb(n6209), .dout(n15563));
  jand g15427(.dina(n11956), .dinb(n6131), .dout(n15564));
  jand g15428(.dina(n11958), .dinb(n5691), .dout(n15565));
  jor  g15429(.dina(n15565), .dinb(n15564), .dout(n15566));
  jor  g15430(.dina(n15566), .dinb(n15563), .dout(n15567));
  jor  g15431(.dina(n15567), .dinb(n15562), .dout(n15568));
  jxor g15432(.dina(n15568), .dinb(n4247), .dout(n15569));
  jor  g15433(.dina(n15569), .dinb(n15561), .dout(n15570));
  jand g15434(.dina(n15570), .dinb(n15559), .dout(n15571));
  jnot g15435(.din(n15571), .dout(n15572));
  jxor g15436(.dina(n15231), .dinb(n15223), .dout(n15573));
  jand g15437(.dina(n15573), .dinb(n15572), .dout(n15574));
  jnot g15438(.din(n15574), .dout(n15575));
  jxor g15439(.dina(n15573), .dinb(n15572), .dout(n15576));
  jnot g15440(.din(n15576), .dout(n15577));
  jand g15441(.dina(n12519), .dinb(n6340), .dout(n15578));
  jand g15442(.dina(n11946), .dinb(n6798), .dout(n15579));
  jand g15443(.dina(n11948), .dinb(n6556), .dout(n15580));
  jand g15444(.dina(n11950), .dinb(n6338), .dout(n15581));
  jor  g15445(.dina(n15581), .dinb(n15580), .dout(n15582));
  jor  g15446(.dina(n15582), .dinb(n15579), .dout(n15583));
  jor  g15447(.dina(n15583), .dinb(n15578), .dout(n15584));
  jxor g15448(.dina(n15584), .dinb(n5064), .dout(n15585));
  jor  g15449(.dina(n15585), .dinb(n15577), .dout(n15586));
  jand g15450(.dina(n15586), .dinb(n15575), .dout(n15587));
  jnot g15451(.din(n15587), .dout(n15588));
  jxor g15452(.dina(n15305), .dinb(n15297), .dout(n15589));
  jand g15453(.dina(n15589), .dinb(n15588), .dout(n15590));
  jnot g15454(.din(n15590), .dout(n15591));
  jand g15455(.dina(n15591), .dinb(n15306), .dout(n15592));
  jnot g15456(.din(n15592), .dout(n15593));
  jxor g15457(.dina(n15252), .dinb(n15244), .dout(n15594));
  jand g15458(.dina(n15594), .dinb(n15593), .dout(n15595));
  jnot g15459(.din(n15595), .dout(n15596));
  jxor g15460(.dina(n15594), .dinb(n15593), .dout(n15597));
  jnot g15461(.din(n15597), .dout(n15598));
  jand g15462(.dina(n12768), .dinb(n6936), .dout(n15599));
  jand g15463(.dina(n12766), .dinb(n7741), .dout(n15600));
  jand g15464(.dina(n12177), .dinb(n7613), .dout(n15601));
  jand g15465(.dina(n11941), .dinb(n6934), .dout(n15602));
  jor  g15466(.dina(n15602), .dinb(n15601), .dout(n15603));
  jor  g15467(.dina(n15603), .dinb(n15600), .dout(n15604));
  jor  g15468(.dina(n15604), .dinb(n15599), .dout(n15605));
  jxor g15469(.dina(n15605), .dinb(n5292), .dout(n15606));
  jor  g15470(.dina(n15606), .dinb(n15598), .dout(n15607));
  jand g15471(.dina(n15607), .dinb(n15596), .dout(n15608));
  jnot g15472(.din(n15608), .dout(n15609));
  jxor g15473(.dina(n15268), .dinb(n15260), .dout(n15610));
  jand g15474(.dina(n15610), .dinb(n15609), .dout(n15611));
  jnot g15475(.din(n15611), .dout(n15612));
  jxor g15476(.dina(n15610), .dinb(n15609), .dout(n15613));
  jnot g15477(.din(n15613), .dout(n15614));
  jand g15478(.dina(n12919), .dinb(n7890), .dout(n15615));
  jand g15479(.dina(n12815), .dinb(n8441), .dout(n15616));
  jand g15480(.dina(n12795), .dinb(n8154), .dout(n15617));
  jand g15481(.dina(n12782), .dinb(n7888), .dout(n15618));
  jor  g15482(.dina(n15618), .dinb(n15617), .dout(n15619));
  jor  g15483(.dina(n15619), .dinb(n15616), .dout(n15620));
  jor  g15484(.dina(n15620), .dinb(n15615), .dout(n15621));
  jxor g15485(.dina(n15621), .dinb(n5833), .dout(n15622));
  jor  g15486(.dina(n15622), .dinb(n15614), .dout(n15623));
  jand g15487(.dina(n15623), .dinb(n15612), .dout(n15624));
  jand g15488(.dina(n13022), .dinb(n7890), .dout(n15625));
  jand g15489(.dina(n12815), .dinb(n8154), .dout(n15627));
  jand g15490(.dina(n12795), .dinb(n7888), .dout(n15628));
  jor  g15491(.dina(n15628), .dinb(n15627), .dout(n15629));
  jor  g15492(.dina(n15629), .dinb(n8441), .dout(n15630));
  jor  g15493(.dina(n15630), .dinb(n15625), .dout(n15631));
  jxor g15494(.dina(n15631), .dinb(n5833), .dout(n15632));
  jor  g15495(.dina(n15632), .dinb(n15624), .dout(n15633));
  jxor g15496(.dina(n15272), .dinb(n15271), .dout(n15634));
  jxor g15497(.dina(n15632), .dinb(n15624), .dout(n15635));
  jand g15498(.dina(n15635), .dinb(n15634), .dout(n15636));
  jnot g15499(.din(n15636), .dout(n15637));
  jand g15500(.dina(n15637), .dinb(n15633), .dout(n15638));
  jnot g15501(.din(n15638), .dout(n15639));
  jxor g15502(.dina(n15289), .dinb(n15281), .dout(n15640));
  jand g15503(.dina(n15640), .dinb(n15639), .dout(n15641));
  jxor g15504(.dina(n15589), .dinb(n15588), .dout(n15642));
  jnot g15505(.din(n15642), .dout(n15643));
  jand g15506(.dina(n12179), .dinb(n6936), .dout(n15644));
  jand g15507(.dina(n12177), .dinb(n7741), .dout(n15645));
  jand g15508(.dina(n11941), .dinb(n7613), .dout(n15646));
  jand g15509(.dina(n11942), .dinb(n6934), .dout(n15647));
  jor  g15510(.dina(n15647), .dinb(n15646), .dout(n15648));
  jor  g15511(.dina(n15648), .dinb(n15645), .dout(n15649));
  jor  g15512(.dina(n15649), .dinb(n15644), .dout(n15650));
  jxor g15513(.dina(n15650), .dinb(n5292), .dout(n15651));
  jor  g15514(.dina(n15651), .dinb(n15643), .dout(n15652));
  jand g15515(.dina(n13470), .dinb(n5365), .dout(n15653));
  jand g15516(.dina(n11964), .dinb(n5500), .dout(n15654));
  jand g15517(.dina(n11966), .dinb(n5424), .dout(n15655));
  jand g15518(.dina(n11968), .dinb(n5363), .dout(n15656));
  jor  g15519(.dina(n15656), .dinb(n15655), .dout(n15657));
  jor  g15520(.dina(n15657), .dinb(n15654), .dout(n15658));
  jor  g15521(.dina(n15658), .dinb(n15653), .dout(n15659));
  jxor g15522(.dina(n15659), .dinb(n72), .dout(n15660));
  jnot g15523(.din(n15660), .dout(n15661));
  jxor g15524(.dina(n15536), .dinb(n15535), .dout(n15662));
  jand g15525(.dina(n15662), .dinb(n15661), .dout(n15663));
  jand g15526(.dina(n13268), .dinb(n5365), .dout(n15664));
  jand g15527(.dina(n11966), .dinb(n5500), .dout(n15665));
  jand g15528(.dina(n11968), .dinb(n5424), .dout(n15666));
  jand g15529(.dina(n11970), .dinb(n5363), .dout(n15667));
  jor  g15530(.dina(n15667), .dinb(n15666), .dout(n15668));
  jor  g15531(.dina(n15668), .dinb(n15665), .dout(n15669));
  jor  g15532(.dina(n15669), .dinb(n15664), .dout(n15670));
  jxor g15533(.dina(n15670), .dinb(n72), .dout(n15671));
  jnot g15534(.din(n15671), .dout(n15672));
  jxor g15535(.dina(n15531), .dinb(n15530), .dout(n15673));
  jand g15536(.dina(n15673), .dinb(n15672), .dout(n15674));
  jand g15537(.dina(n13682), .dinb(n5365), .dout(n15675));
  jand g15538(.dina(n11968), .dinb(n5500), .dout(n15676));
  jand g15539(.dina(n11970), .dinb(n5424), .dout(n15677));
  jand g15540(.dina(n11972), .dinb(n5363), .dout(n15678));
  jor  g15541(.dina(n15678), .dinb(n15677), .dout(n15679));
  jor  g15542(.dina(n15679), .dinb(n15676), .dout(n15680));
  jor  g15543(.dina(n15680), .dinb(n15675), .dout(n15681));
  jxor g15544(.dina(n15681), .dinb(n72), .dout(n15682));
  jnot g15545(.din(n15682), .dout(n15683));
  jxor g15546(.dina(n15526), .dinb(n15525), .dout(n15684));
  jand g15547(.dina(n15684), .dinb(n15683), .dout(n15685));
  jand g15548(.dina(n13806), .dinb(n5365), .dout(n15686));
  jand g15549(.dina(n11970), .dinb(n5500), .dout(n15687));
  jand g15550(.dina(n11972), .dinb(n5424), .dout(n15688));
  jand g15551(.dina(n11974), .dinb(n5363), .dout(n15689));
  jor  g15552(.dina(n15689), .dinb(n15688), .dout(n15690));
  jor  g15553(.dina(n15690), .dinb(n15687), .dout(n15691));
  jor  g15554(.dina(n15691), .dinb(n15686), .dout(n15692));
  jxor g15555(.dina(n15692), .dinb(n72), .dout(n15693));
  jnot g15556(.din(n15693), .dout(n15694));
  jxor g15557(.dina(n15521), .dinb(n15520), .dout(n15695));
  jand g15558(.dina(n15695), .dinb(n15694), .dout(n15696));
  jand g15559(.dina(n13664), .dinb(n5365), .dout(n15697));
  jand g15560(.dina(n11972), .dinb(n5500), .dout(n15698));
  jand g15561(.dina(n11974), .dinb(n5424), .dout(n15699));
  jand g15562(.dina(n11976), .dinb(n5363), .dout(n15700));
  jor  g15563(.dina(n15700), .dinb(n15699), .dout(n15701));
  jor  g15564(.dina(n15701), .dinb(n15698), .dout(n15702));
  jor  g15565(.dina(n15702), .dinb(n15697), .dout(n15703));
  jxor g15566(.dina(n15703), .dinb(n72), .dout(n15704));
  jnot g15567(.din(n15704), .dout(n15705));
  jxor g15568(.dina(n15516), .dinb(n15515), .dout(n15706));
  jand g15569(.dina(n15706), .dinb(n15705), .dout(n15707));
  jand g15570(.dina(n13924), .dinb(n5365), .dout(n15708));
  jand g15571(.dina(n11974), .dinb(n5500), .dout(n15709));
  jand g15572(.dina(n11976), .dinb(n5424), .dout(n15710));
  jand g15573(.dina(n11978), .dinb(n5363), .dout(n15711));
  jor  g15574(.dina(n15711), .dinb(n15710), .dout(n15712));
  jor  g15575(.dina(n15712), .dinb(n15709), .dout(n15713));
  jor  g15576(.dina(n15713), .dinb(n15708), .dout(n15714));
  jxor g15577(.dina(n15714), .dinb(n72), .dout(n15715));
  jnot g15578(.din(n15715), .dout(n15716));
  jxor g15579(.dina(n15511), .dinb(n15510), .dout(n15717));
  jand g15580(.dina(n15717), .dinb(n15716), .dout(n15718));
  jand g15581(.dina(n14184), .dinb(n5365), .dout(n15719));
  jand g15582(.dina(n11976), .dinb(n5500), .dout(n15720));
  jand g15583(.dina(n11978), .dinb(n5424), .dout(n15721));
  jand g15584(.dina(n11980), .dinb(n5363), .dout(n15722));
  jor  g15585(.dina(n15722), .dinb(n15721), .dout(n15723));
  jor  g15586(.dina(n15723), .dinb(n15720), .dout(n15724));
  jor  g15587(.dina(n15724), .dinb(n15719), .dout(n15725));
  jxor g15588(.dina(n15725), .dinb(n72), .dout(n15726));
  jnot g15589(.din(n15726), .dout(n15727));
  jxor g15590(.dina(n15506), .dinb(n15505), .dout(n15728));
  jand g15591(.dina(n15728), .dinb(n15727), .dout(n15729));
  jand g15592(.dina(n14194), .dinb(n5365), .dout(n15730));
  jand g15593(.dina(n11978), .dinb(n5500), .dout(n15731));
  jand g15594(.dina(n11980), .dinb(n5424), .dout(n15732));
  jand g15595(.dina(n11982), .dinb(n5363), .dout(n15733));
  jor  g15596(.dina(n15733), .dinb(n15732), .dout(n15734));
  jor  g15597(.dina(n15734), .dinb(n15731), .dout(n15735));
  jor  g15598(.dina(n15735), .dinb(n15730), .dout(n15736));
  jxor g15599(.dina(n15736), .dinb(n72), .dout(n15737));
  jnot g15600(.din(n15737), .dout(n15738));
  jxor g15601(.dina(n15501), .dinb(n15500), .dout(n15739));
  jand g15602(.dina(n15739), .dinb(n15738), .dout(n15740));
  jand g15603(.dina(n13899), .dinb(n5365), .dout(n15741));
  jand g15604(.dina(n11980), .dinb(n5500), .dout(n15742));
  jand g15605(.dina(n11982), .dinb(n5424), .dout(n15743));
  jand g15606(.dina(n11985), .dinb(n5363), .dout(n15744));
  jor  g15607(.dina(n15744), .dinb(n15743), .dout(n15745));
  jor  g15608(.dina(n15745), .dinb(n15742), .dout(n15746));
  jor  g15609(.dina(n15746), .dinb(n15741), .dout(n15747));
  jxor g15610(.dina(n15747), .dinb(n72), .dout(n15748));
  jnot g15611(.din(n15748), .dout(n15749));
  jxor g15612(.dina(n15496), .dinb(n15495), .dout(n15750));
  jand g15613(.dina(n15750), .dinb(n15749), .dout(n15751));
  jor  g15614(.dina(n14221), .dinb(n5366), .dout(n15752));
  jor  g15615(.dina(n15045), .dinb(n5499), .dout(n15753));
  jor  g15616(.dina(n11984), .dinb(n5425), .dout(n15754));
  jor  g15617(.dina(n11987), .dinb(n5364), .dout(n15755));
  jand g15618(.dina(n15755), .dinb(n15754), .dout(n15756));
  jand g15619(.dina(n15756), .dinb(n15753), .dout(n15757));
  jand g15620(.dina(n15757), .dinb(n15752), .dout(n15758));
  jxor g15621(.dina(n15758), .dinb(\a[23] ), .dout(n15759));
  jnot g15622(.din(n15759), .dout(n15760));
  jxor g15623(.dina(n15493), .dinb(n15492), .dout(n15761));
  jand g15624(.dina(n15761), .dinb(n15760), .dout(n15762));
  jxor g15625(.dina(n15490), .dinb(n15489), .dout(n15763));
  jnot g15626(.din(n15763), .dout(n15764));
  jor  g15627(.dina(n14248), .dinb(n5366), .dout(n15765));
  jor  g15628(.dina(n11984), .dinb(n5499), .dout(n15766));
  jor  g15629(.dina(n11987), .dinb(n5425), .dout(n15767));
  jor  g15630(.dina(n11991), .dinb(n5364), .dout(n15768));
  jand g15631(.dina(n15768), .dinb(n15767), .dout(n15769));
  jand g15632(.dina(n15769), .dinb(n15766), .dout(n15770));
  jand g15633(.dina(n15770), .dinb(n15765), .dout(n15771));
  jxor g15634(.dina(n15771), .dinb(\a[23] ), .dout(n15772));
  jor  g15635(.dina(n15772), .dinb(n15764), .dout(n15773));
  jxor g15636(.dina(n15487), .dinb(n15486), .dout(n15774));
  jnot g15637(.din(n15774), .dout(n15775));
  jor  g15638(.dina(n14271), .dinb(n5366), .dout(n15776));
  jor  g15639(.dina(n11987), .dinb(n5499), .dout(n15777));
  jor  g15640(.dina(n11991), .dinb(n5425), .dout(n15778));
  jor  g15641(.dina(n11995), .dinb(n5364), .dout(n15779));
  jand g15642(.dina(n15779), .dinb(n15778), .dout(n15780));
  jand g15643(.dina(n15780), .dinb(n15777), .dout(n15781));
  jand g15644(.dina(n15781), .dinb(n15776), .dout(n15782));
  jxor g15645(.dina(n15782), .dinb(\a[23] ), .dout(n15783));
  jor  g15646(.dina(n15783), .dinb(n15775), .dout(n15784));
  jor  g15647(.dina(n14301), .dinb(n5366), .dout(n15785));
  jor  g15648(.dina(n11991), .dinb(n5499), .dout(n15786));
  jor  g15649(.dina(n11995), .dinb(n5425), .dout(n15787));
  jor  g15650(.dina(n11997), .dinb(n5364), .dout(n15788));
  jand g15651(.dina(n15788), .dinb(n15787), .dout(n15789));
  jand g15652(.dina(n15789), .dinb(n15786), .dout(n15790));
  jand g15653(.dina(n15790), .dinb(n15785), .dout(n15791));
  jxor g15654(.dina(n15791), .dinb(\a[23] ), .dout(n15792));
  jnot g15655(.din(n15792), .dout(n15793));
  jxor g15656(.dina(n15484), .dinb(n15483), .dout(n15794));
  jand g15657(.dina(n15794), .dinb(n15793), .dout(n15795));
  jor  g15658(.dina(n14353), .dinb(n5366), .dout(n15796));
  jor  g15659(.dina(n11995), .dinb(n5499), .dout(n15797));
  jor  g15660(.dina(n11997), .dinb(n5425), .dout(n15798));
  jor  g15661(.dina(n11999), .dinb(n5364), .dout(n15799));
  jand g15662(.dina(n15799), .dinb(n15798), .dout(n15800));
  jand g15663(.dina(n15800), .dinb(n15797), .dout(n15801));
  jand g15664(.dina(n15801), .dinb(n15796), .dout(n15802));
  jxor g15665(.dina(n15802), .dinb(\a[23] ), .dout(n15803));
  jnot g15666(.din(n15803), .dout(n15804));
  jxor g15667(.dina(n15481), .dinb(n15480), .dout(n15805));
  jand g15668(.dina(n15805), .dinb(n15804), .dout(n15806));
  jor  g15669(.dina(n14390), .dinb(n5366), .dout(n15807));
  jor  g15670(.dina(n11997), .dinb(n5499), .dout(n15808));
  jor  g15671(.dina(n11999), .dinb(n5425), .dout(n15809));
  jor  g15672(.dina(n12001), .dinb(n5364), .dout(n15810));
  jand g15673(.dina(n15810), .dinb(n15809), .dout(n15811));
  jand g15674(.dina(n15811), .dinb(n15808), .dout(n15812));
  jand g15675(.dina(n15812), .dinb(n15807), .dout(n15813));
  jxor g15676(.dina(n15813), .dinb(\a[23] ), .dout(n15814));
  jnot g15677(.din(n15814), .dout(n15815));
  jor  g15678(.dina(n15461), .dinb(n68), .dout(n15816));
  jxor g15679(.dina(n15816), .dinb(n15469), .dout(n15817));
  jand g15680(.dina(n15817), .dinb(n15815), .dout(n15818));
  jor  g15681(.dina(n14432), .dinb(n5366), .dout(n15819));
  jor  g15682(.dina(n11999), .dinb(n5499), .dout(n15820));
  jor  g15683(.dina(n12001), .dinb(n5425), .dout(n15821));
  jor  g15684(.dina(n12004), .dinb(n5364), .dout(n15822));
  jand g15685(.dina(n15822), .dinb(n15821), .dout(n15823));
  jand g15686(.dina(n15823), .dinb(n15820), .dout(n15824));
  jand g15687(.dina(n15824), .dinb(n15819), .dout(n15825));
  jxor g15688(.dina(n15825), .dinb(\a[23] ), .dout(n15826));
  jnot g15689(.din(n15826), .dout(n15827));
  jand g15690(.dina(n15458), .dinb(\a[26] ), .dout(n15828));
  jxor g15691(.dina(n15828), .dinb(n15456), .dout(n15829));
  jand g15692(.dina(n15829), .dinb(n15827), .dout(n15830));
  jand g15693(.dina(n14497), .dinb(n5365), .dout(n15831));
  jand g15694(.dina(n12010), .dinb(n5424), .dout(n15832));
  jand g15695(.dina(n12008), .dinb(n5500), .dout(n15833));
  jor  g15696(.dina(n15833), .dinb(n15832), .dout(n15834));
  jor  g15697(.dina(n15834), .dinb(n15831), .dout(n15835));
  jnot g15698(.din(n15835), .dout(n15836));
  jand g15699(.dina(n12010), .dinb(n5358), .dout(n15837));
  jnot g15700(.din(n15837), .dout(n15838));
  jand g15701(.dina(n15838), .dinb(\a[23] ), .dout(n15839));
  jand g15702(.dina(n15839), .dinb(n15836), .dout(n15840));
  jand g15703(.dina(n14537), .dinb(n5365), .dout(n15841));
  jand g15704(.dina(n12006), .dinb(n5500), .dout(n15842));
  jand g15705(.dina(n12008), .dinb(n5424), .dout(n15843));
  jand g15706(.dina(n12010), .dinb(n5363), .dout(n15844));
  jor  g15707(.dina(n15844), .dinb(n15843), .dout(n15845));
  jor  g15708(.dina(n15845), .dinb(n15842), .dout(n15846));
  jor  g15709(.dina(n15846), .dinb(n15841), .dout(n15847));
  jnot g15710(.din(n15847), .dout(n15848));
  jand g15711(.dina(n15848), .dinb(n15840), .dout(n15849));
  jand g15712(.dina(n15849), .dinb(n15458), .dout(n15850));
  jor  g15713(.dina(n15144), .dinb(n5366), .dout(n15851));
  jor  g15714(.dina(n12001), .dinb(n5499), .dout(n15852));
  jor  g15715(.dina(n12004), .dinb(n5425), .dout(n15853));
  jor  g15716(.dina(n12009), .dinb(n5364), .dout(n15854));
  jand g15717(.dina(n15854), .dinb(n15853), .dout(n15855));
  jand g15718(.dina(n15855), .dinb(n15852), .dout(n15856));
  jand g15719(.dina(n15856), .dinb(n15851), .dout(n15857));
  jxor g15720(.dina(n15857), .dinb(\a[23] ), .dout(n15858));
  jnot g15721(.din(n15858), .dout(n15859));
  jxor g15722(.dina(n15849), .dinb(n15458), .dout(n15860));
  jand g15723(.dina(n15860), .dinb(n15859), .dout(n15861));
  jor  g15724(.dina(n15861), .dinb(n15850), .dout(n15862));
  jxor g15725(.dina(n15829), .dinb(n15827), .dout(n15863));
  jand g15726(.dina(n15863), .dinb(n15862), .dout(n15864));
  jor  g15727(.dina(n15864), .dinb(n15830), .dout(n15865));
  jxor g15728(.dina(n15817), .dinb(n15815), .dout(n15866));
  jand g15729(.dina(n15866), .dinb(n15865), .dout(n15867));
  jor  g15730(.dina(n15867), .dinb(n15818), .dout(n15868));
  jxor g15731(.dina(n15805), .dinb(n15804), .dout(n15869));
  jand g15732(.dina(n15869), .dinb(n15868), .dout(n15870));
  jor  g15733(.dina(n15870), .dinb(n15806), .dout(n15871));
  jxor g15734(.dina(n15794), .dinb(n15793), .dout(n15872));
  jand g15735(.dina(n15872), .dinb(n15871), .dout(n15873));
  jor  g15736(.dina(n15873), .dinb(n15795), .dout(n15874));
  jxor g15737(.dina(n15783), .dinb(n15775), .dout(n15875));
  jand g15738(.dina(n15875), .dinb(n15874), .dout(n15876));
  jnot g15739(.din(n15876), .dout(n15877));
  jand g15740(.dina(n15877), .dinb(n15784), .dout(n15878));
  jnot g15741(.din(n15878), .dout(n15879));
  jxor g15742(.dina(n15772), .dinb(n15764), .dout(n15880));
  jand g15743(.dina(n15880), .dinb(n15879), .dout(n15881));
  jnot g15744(.din(n15881), .dout(n15882));
  jand g15745(.dina(n15882), .dinb(n15773), .dout(n15883));
  jnot g15746(.din(n15883), .dout(n15884));
  jxor g15747(.dina(n15761), .dinb(n15760), .dout(n15885));
  jand g15748(.dina(n15885), .dinb(n15884), .dout(n15886));
  jor  g15749(.dina(n15886), .dinb(n15762), .dout(n15887));
  jxor g15750(.dina(n15750), .dinb(n15749), .dout(n15888));
  jand g15751(.dina(n15888), .dinb(n15887), .dout(n15889));
  jor  g15752(.dina(n15889), .dinb(n15751), .dout(n15890));
  jxor g15753(.dina(n15739), .dinb(n15738), .dout(n15891));
  jand g15754(.dina(n15891), .dinb(n15890), .dout(n15892));
  jor  g15755(.dina(n15892), .dinb(n15740), .dout(n15893));
  jxor g15756(.dina(n15728), .dinb(n15727), .dout(n15894));
  jand g15757(.dina(n15894), .dinb(n15893), .dout(n15895));
  jor  g15758(.dina(n15895), .dinb(n15729), .dout(n15896));
  jxor g15759(.dina(n15717), .dinb(n15716), .dout(n15897));
  jand g15760(.dina(n15897), .dinb(n15896), .dout(n15898));
  jor  g15761(.dina(n15898), .dinb(n15718), .dout(n15899));
  jxor g15762(.dina(n15706), .dinb(n15705), .dout(n15900));
  jand g15763(.dina(n15900), .dinb(n15899), .dout(n15901));
  jor  g15764(.dina(n15901), .dinb(n15707), .dout(n15902));
  jxor g15765(.dina(n15695), .dinb(n15694), .dout(n15903));
  jand g15766(.dina(n15903), .dinb(n15902), .dout(n15904));
  jor  g15767(.dina(n15904), .dinb(n15696), .dout(n15905));
  jxor g15768(.dina(n15684), .dinb(n15683), .dout(n15906));
  jand g15769(.dina(n15906), .dinb(n15905), .dout(n15907));
  jor  g15770(.dina(n15907), .dinb(n15685), .dout(n15908));
  jxor g15771(.dina(n15673), .dinb(n15672), .dout(n15909));
  jand g15772(.dina(n15909), .dinb(n15908), .dout(n15910));
  jor  g15773(.dina(n15910), .dinb(n15674), .dout(n15911));
  jxor g15774(.dina(n15662), .dinb(n15661), .dout(n15912));
  jand g15775(.dina(n15912), .dinb(n15911), .dout(n15913));
  jor  g15776(.dina(n15913), .dinb(n15663), .dout(n15914));
  jxor g15777(.dina(n15553), .dinb(n15545), .dout(n15915));
  jand g15778(.dina(n15915), .dinb(n15914), .dout(n15916));
  jnot g15779(.din(n15916), .dout(n15917));
  jxor g15780(.dina(n15915), .dinb(n15914), .dout(n15918));
  jnot g15781(.din(n15918), .dout(n15919));
  jand g15782(.dina(n12639), .dinb(n5693), .dout(n15920));
  jand g15783(.dina(n11956), .dinb(n6209), .dout(n15921));
  jand g15784(.dina(n11958), .dinb(n6131), .dout(n15922));
  jand g15785(.dina(n11960), .dinb(n5691), .dout(n15923));
  jor  g15786(.dina(n15923), .dinb(n15922), .dout(n15924));
  jor  g15787(.dina(n15924), .dinb(n15921), .dout(n15925));
  jor  g15788(.dina(n15925), .dinb(n15920), .dout(n15926));
  jxor g15789(.dina(n15926), .dinb(n4247), .dout(n15927));
  jor  g15790(.dina(n15927), .dinb(n15919), .dout(n15928));
  jand g15791(.dina(n15928), .dinb(n15917), .dout(n15929));
  jnot g15792(.din(n15929), .dout(n15930));
  jxor g15793(.dina(n15569), .dinb(n15561), .dout(n15931));
  jand g15794(.dina(n15931), .dinb(n15930), .dout(n15932));
  jnot g15795(.din(n15932), .dout(n15933));
  jxor g15796(.dina(n15931), .dinb(n15930), .dout(n15934));
  jnot g15797(.din(n15934), .dout(n15935));
  jand g15798(.dina(n12654), .dinb(n6340), .dout(n15936));
  jand g15799(.dina(n11948), .dinb(n6798), .dout(n15937));
  jand g15800(.dina(n11950), .dinb(n6556), .dout(n15938));
  jand g15801(.dina(n11952), .dinb(n6338), .dout(n15939));
  jor  g15802(.dina(n15939), .dinb(n15938), .dout(n15940));
  jor  g15803(.dina(n15940), .dinb(n15937), .dout(n15941));
  jor  g15804(.dina(n15941), .dinb(n15936), .dout(n15942));
  jxor g15805(.dina(n15942), .dinb(n5064), .dout(n15943));
  jor  g15806(.dina(n15943), .dinb(n15935), .dout(n15944));
  jand g15807(.dina(n15944), .dinb(n15933), .dout(n15945));
  jnot g15808(.din(n15945), .dout(n15946));
  jxor g15809(.dina(n15585), .dinb(n15577), .dout(n15947));
  jand g15810(.dina(n15947), .dinb(n15946), .dout(n15948));
  jnot g15811(.din(n15948), .dout(n15949));
  jxor g15812(.dina(n15947), .dinb(n15946), .dout(n15950));
  jnot g15813(.din(n15950), .dout(n15951));
  jand g15814(.dina(n12671), .dinb(n6936), .dout(n15952));
  jand g15815(.dina(n11941), .dinb(n7741), .dout(n15953));
  jand g15816(.dina(n11942), .dinb(n7613), .dout(n15954));
  jand g15817(.dina(n11944), .dinb(n6934), .dout(n15955));
  jor  g15818(.dina(n15955), .dinb(n15954), .dout(n15956));
  jor  g15819(.dina(n15956), .dinb(n15953), .dout(n15957));
  jor  g15820(.dina(n15957), .dinb(n15952), .dout(n15958));
  jxor g15821(.dina(n15958), .dinb(n5292), .dout(n15959));
  jor  g15822(.dina(n15959), .dinb(n15951), .dout(n15960));
  jand g15823(.dina(n15960), .dinb(n15949), .dout(n15961));
  jnot g15824(.din(n15961), .dout(n15962));
  jxor g15825(.dina(n15651), .dinb(n15643), .dout(n15963));
  jand g15826(.dina(n15963), .dinb(n15962), .dout(n15964));
  jnot g15827(.din(n15964), .dout(n15965));
  jand g15828(.dina(n15965), .dinb(n15652), .dout(n15966));
  jnot g15829(.din(n15966), .dout(n15967));
  jxor g15830(.dina(n15606), .dinb(n15598), .dout(n15968));
  jand g15831(.dina(n15968), .dinb(n15967), .dout(n15969));
  jnot g15832(.din(n15969), .dout(n15970));
  jxor g15833(.dina(n15968), .dinb(n15967), .dout(n15971));
  jnot g15834(.din(n15971), .dout(n15972));
  jand g15835(.dina(n12797), .dinb(n7890), .dout(n15973));
  jand g15836(.dina(n12795), .dinb(n8441), .dout(n15974));
  jand g15837(.dina(n12782), .dinb(n8154), .dout(n15975));
  jand g15838(.dina(n12783), .dinb(n7888), .dout(n15976));
  jor  g15839(.dina(n15976), .dinb(n15975), .dout(n15977));
  jor  g15840(.dina(n15977), .dinb(n15974), .dout(n15978));
  jor  g15841(.dina(n15978), .dinb(n15973), .dout(n15979));
  jxor g15842(.dina(n15979), .dinb(n5833), .dout(n15980));
  jor  g15843(.dina(n15980), .dinb(n15972), .dout(n15981));
  jand g15844(.dina(n15981), .dinb(n15970), .dout(n15982));
  jand g15845(.dina(n9490), .dinb(n9127), .dout(n15985));
  jor  g15846(.dina(n13261), .dinb(n15982), .dout(n15990));
  jxor g15847(.dina(n13261), .dinb(n15982), .dout(n15991));
  jxor g15848(.dina(n15622), .dinb(n15614), .dout(n15992));
  jand g15849(.dina(n15992), .dinb(n15991), .dout(n15993));
  jnot g15850(.din(n15993), .dout(n15994));
  jand g15851(.dina(n15994), .dinb(n15990), .dout(n15995));
  jnot g15852(.din(n15995), .dout(n15996));
  jxor g15853(.dina(n15635), .dinb(n15634), .dout(n15997));
  jand g15854(.dina(n15997), .dinb(n15996), .dout(n15998));
  jxor g15855(.dina(n15963), .dinb(n15962), .dout(n15999));
  jnot g15856(.din(n15999), .dout(n16000));
  jand g15857(.dina(n12938), .dinb(n7890), .dout(n16001));
  jand g15858(.dina(n12782), .dinb(n8441), .dout(n16002));
  jand g15859(.dina(n12783), .dinb(n8154), .dout(n16003));
  jand g15860(.dina(n12766), .dinb(n7888), .dout(n16004));
  jor  g15861(.dina(n16004), .dinb(n16003), .dout(n16005));
  jor  g15862(.dina(n16005), .dinb(n16002), .dout(n16006));
  jor  g15863(.dina(n16006), .dinb(n16001), .dout(n16007));
  jxor g15864(.dina(n16007), .dinb(n5833), .dout(n16008));
  jor  g15865(.dina(n16008), .dinb(n16000), .dout(n16009));
  jxor g15866(.dina(n15912), .dinb(n15911), .dout(n16010));
  jnot g15867(.din(n16010), .dout(n16011));
  jand g15868(.dina(n12624), .dinb(n5693), .dout(n16012));
  jand g15869(.dina(n11958), .dinb(n6209), .dout(n16013));
  jand g15870(.dina(n11960), .dinb(n6131), .dout(n16014));
  jand g15871(.dina(n11962), .dinb(n5691), .dout(n16015));
  jor  g15872(.dina(n16015), .dinb(n16014), .dout(n16016));
  jor  g15873(.dina(n16016), .dinb(n16013), .dout(n16017));
  jor  g15874(.dina(n16017), .dinb(n16012), .dout(n16018));
  jxor g15875(.dina(n16018), .dinb(n4247), .dout(n16019));
  jor  g15876(.dina(n16019), .dinb(n16011), .dout(n16020));
  jxor g15877(.dina(n15909), .dinb(n15908), .dout(n16021));
  jnot g15878(.din(n16021), .dout(n16022));
  jand g15879(.dina(n13116), .dinb(n5693), .dout(n16023));
  jand g15880(.dina(n11960), .dinb(n6209), .dout(n16024));
  jand g15881(.dina(n11962), .dinb(n6131), .dout(n16025));
  jand g15882(.dina(n11964), .dinb(n5691), .dout(n16026));
  jor  g15883(.dina(n16026), .dinb(n16025), .dout(n16027));
  jor  g15884(.dina(n16027), .dinb(n16024), .dout(n16028));
  jor  g15885(.dina(n16028), .dinb(n16023), .dout(n16029));
  jxor g15886(.dina(n16029), .dinb(n4247), .dout(n16030));
  jor  g15887(.dina(n16030), .dinb(n16022), .dout(n16031));
  jxor g15888(.dina(n15906), .dinb(n15905), .dout(n16032));
  jnot g15889(.din(n16032), .dout(n16033));
  jand g15890(.dina(n13134), .dinb(n5693), .dout(n16034));
  jand g15891(.dina(n11962), .dinb(n6209), .dout(n16035));
  jand g15892(.dina(n11964), .dinb(n6131), .dout(n16036));
  jand g15893(.dina(n11966), .dinb(n5691), .dout(n16037));
  jor  g15894(.dina(n16037), .dinb(n16036), .dout(n16038));
  jor  g15895(.dina(n16038), .dinb(n16035), .dout(n16039));
  jor  g15896(.dina(n16039), .dinb(n16034), .dout(n16040));
  jxor g15897(.dina(n16040), .dinb(n4247), .dout(n16041));
  jor  g15898(.dina(n16041), .dinb(n16033), .dout(n16042));
  jxor g15899(.dina(n15903), .dinb(n15902), .dout(n16043));
  jnot g15900(.din(n16043), .dout(n16044));
  jand g15901(.dina(n13470), .dinb(n5693), .dout(n16045));
  jand g15902(.dina(n11964), .dinb(n6209), .dout(n16046));
  jand g15903(.dina(n11966), .dinb(n6131), .dout(n16047));
  jand g15904(.dina(n11968), .dinb(n5691), .dout(n16048));
  jor  g15905(.dina(n16048), .dinb(n16047), .dout(n16049));
  jor  g15906(.dina(n16049), .dinb(n16046), .dout(n16050));
  jor  g15907(.dina(n16050), .dinb(n16045), .dout(n16051));
  jxor g15908(.dina(n16051), .dinb(n4247), .dout(n16052));
  jor  g15909(.dina(n16052), .dinb(n16044), .dout(n16053));
  jxor g15910(.dina(n15900), .dinb(n15899), .dout(n16054));
  jnot g15911(.din(n16054), .dout(n16055));
  jand g15912(.dina(n13268), .dinb(n5693), .dout(n16056));
  jand g15913(.dina(n11966), .dinb(n6209), .dout(n16057));
  jand g15914(.dina(n11968), .dinb(n6131), .dout(n16058));
  jand g15915(.dina(n11970), .dinb(n5691), .dout(n16059));
  jor  g15916(.dina(n16059), .dinb(n16058), .dout(n16060));
  jor  g15917(.dina(n16060), .dinb(n16057), .dout(n16061));
  jor  g15918(.dina(n16061), .dinb(n16056), .dout(n16062));
  jxor g15919(.dina(n16062), .dinb(n4247), .dout(n16063));
  jor  g15920(.dina(n16063), .dinb(n16055), .dout(n16064));
  jxor g15921(.dina(n15897), .dinb(n15896), .dout(n16065));
  jnot g15922(.din(n16065), .dout(n16066));
  jand g15923(.dina(n13682), .dinb(n5693), .dout(n16067));
  jand g15924(.dina(n11968), .dinb(n6209), .dout(n16068));
  jand g15925(.dina(n11970), .dinb(n6131), .dout(n16069));
  jand g15926(.dina(n11972), .dinb(n5691), .dout(n16070));
  jor  g15927(.dina(n16070), .dinb(n16069), .dout(n16071));
  jor  g15928(.dina(n16071), .dinb(n16068), .dout(n16072));
  jor  g15929(.dina(n16072), .dinb(n16067), .dout(n16073));
  jxor g15930(.dina(n16073), .dinb(n4247), .dout(n16074));
  jor  g15931(.dina(n16074), .dinb(n16066), .dout(n16075));
  jxor g15932(.dina(n15894), .dinb(n15893), .dout(n16076));
  jnot g15933(.din(n16076), .dout(n16077));
  jand g15934(.dina(n13806), .dinb(n5693), .dout(n16078));
  jand g15935(.dina(n11970), .dinb(n6209), .dout(n16079));
  jand g15936(.dina(n11972), .dinb(n6131), .dout(n16080));
  jand g15937(.dina(n11974), .dinb(n5691), .dout(n16081));
  jor  g15938(.dina(n16081), .dinb(n16080), .dout(n16082));
  jor  g15939(.dina(n16082), .dinb(n16079), .dout(n16083));
  jor  g15940(.dina(n16083), .dinb(n16078), .dout(n16084));
  jxor g15941(.dina(n16084), .dinb(n4247), .dout(n16085));
  jor  g15942(.dina(n16085), .dinb(n16077), .dout(n16086));
  jxor g15943(.dina(n15891), .dinb(n15890), .dout(n16087));
  jnot g15944(.din(n16087), .dout(n16088));
  jand g15945(.dina(n13664), .dinb(n5693), .dout(n16089));
  jand g15946(.dina(n11972), .dinb(n6209), .dout(n16090));
  jand g15947(.dina(n11974), .dinb(n6131), .dout(n16091));
  jand g15948(.dina(n11976), .dinb(n5691), .dout(n16092));
  jor  g15949(.dina(n16092), .dinb(n16091), .dout(n16093));
  jor  g15950(.dina(n16093), .dinb(n16090), .dout(n16094));
  jor  g15951(.dina(n16094), .dinb(n16089), .dout(n16095));
  jxor g15952(.dina(n16095), .dinb(n4247), .dout(n16096));
  jor  g15953(.dina(n16096), .dinb(n16088), .dout(n16097));
  jxor g15954(.dina(n15888), .dinb(n15887), .dout(n16098));
  jnot g15955(.din(n16098), .dout(n16099));
  jand g15956(.dina(n13924), .dinb(n5693), .dout(n16100));
  jand g15957(.dina(n11974), .dinb(n6209), .dout(n16101));
  jand g15958(.dina(n11976), .dinb(n6131), .dout(n16102));
  jand g15959(.dina(n11978), .dinb(n5691), .dout(n16103));
  jor  g15960(.dina(n16103), .dinb(n16102), .dout(n16104));
  jor  g15961(.dina(n16104), .dinb(n16101), .dout(n16105));
  jor  g15962(.dina(n16105), .dinb(n16100), .dout(n16106));
  jxor g15963(.dina(n16106), .dinb(n4247), .dout(n16107));
  jor  g15964(.dina(n16107), .dinb(n16099), .dout(n16108));
  jxor g15965(.dina(n15885), .dinb(n15884), .dout(n16109));
  jnot g15966(.din(n16109), .dout(n16110));
  jand g15967(.dina(n14184), .dinb(n5693), .dout(n16111));
  jand g15968(.dina(n11976), .dinb(n6209), .dout(n16112));
  jand g15969(.dina(n11978), .dinb(n6131), .dout(n16113));
  jand g15970(.dina(n11980), .dinb(n5691), .dout(n16114));
  jor  g15971(.dina(n16114), .dinb(n16113), .dout(n16115));
  jor  g15972(.dina(n16115), .dinb(n16112), .dout(n16116));
  jor  g15973(.dina(n16116), .dinb(n16111), .dout(n16117));
  jxor g15974(.dina(n16117), .dinb(n4247), .dout(n16118));
  jor  g15975(.dina(n16118), .dinb(n16110), .dout(n16119));
  jand g15976(.dina(n14194), .dinb(n5693), .dout(n16120));
  jand g15977(.dina(n11978), .dinb(n6209), .dout(n16121));
  jand g15978(.dina(n11980), .dinb(n6131), .dout(n16122));
  jand g15979(.dina(n11982), .dinb(n5691), .dout(n16123));
  jor  g15980(.dina(n16123), .dinb(n16122), .dout(n16124));
  jor  g15981(.dina(n16124), .dinb(n16121), .dout(n16125));
  jor  g15982(.dina(n16125), .dinb(n16120), .dout(n16126));
  jxor g15983(.dina(n16126), .dinb(n4247), .dout(n16127));
  jnot g15984(.din(n16127), .dout(n16128));
  jxor g15985(.dina(n15880), .dinb(n15879), .dout(n16129));
  jand g15986(.dina(n16129), .dinb(n16128), .dout(n16130));
  jand g15987(.dina(n13899), .dinb(n5693), .dout(n16131));
  jand g15988(.dina(n11980), .dinb(n6209), .dout(n16132));
  jand g15989(.dina(n11982), .dinb(n6131), .dout(n16133));
  jand g15990(.dina(n11985), .dinb(n5691), .dout(n16134));
  jor  g15991(.dina(n16134), .dinb(n16133), .dout(n16135));
  jor  g15992(.dina(n16135), .dinb(n16132), .dout(n16136));
  jor  g15993(.dina(n16136), .dinb(n16131), .dout(n16137));
  jxor g15994(.dina(n16137), .dinb(n4247), .dout(n16138));
  jnot g15995(.din(n16138), .dout(n16139));
  jxor g15996(.dina(n15875), .dinb(n15874), .dout(n16140));
  jand g15997(.dina(n16140), .dinb(n16139), .dout(n16141));
  jxor g15998(.dina(n15872), .dinb(n15871), .dout(n16142));
  jnot g15999(.din(n16142), .dout(n16143));
  jor  g16000(.dina(n14221), .dinb(n5694), .dout(n16144));
  jor  g16001(.dina(n15045), .dinb(n6208), .dout(n16145));
  jor  g16002(.dina(n11984), .dinb(n6132), .dout(n16146));
  jor  g16003(.dina(n11987), .dinb(n5692), .dout(n16147));
  jand g16004(.dina(n16147), .dinb(n16146), .dout(n16148));
  jand g16005(.dina(n16148), .dinb(n16145), .dout(n16149));
  jand g16006(.dina(n16149), .dinb(n16144), .dout(n16150));
  jxor g16007(.dina(n16150), .dinb(\a[20] ), .dout(n16151));
  jor  g16008(.dina(n16151), .dinb(n16143), .dout(n16152));
  jxor g16009(.dina(n15869), .dinb(n15868), .dout(n16153));
  jnot g16010(.din(n16153), .dout(n16154));
  jor  g16011(.dina(n14248), .dinb(n5694), .dout(n16155));
  jor  g16012(.dina(n11984), .dinb(n6208), .dout(n16156));
  jor  g16013(.dina(n11987), .dinb(n6132), .dout(n16157));
  jor  g16014(.dina(n11991), .dinb(n5692), .dout(n16158));
  jand g16015(.dina(n16158), .dinb(n16157), .dout(n16159));
  jand g16016(.dina(n16159), .dinb(n16156), .dout(n16160));
  jand g16017(.dina(n16160), .dinb(n16155), .dout(n16161));
  jxor g16018(.dina(n16161), .dinb(\a[20] ), .dout(n16162));
  jor  g16019(.dina(n16162), .dinb(n16154), .dout(n16163));
  jxor g16020(.dina(n15866), .dinb(n15865), .dout(n16164));
  jnot g16021(.din(n16164), .dout(n16165));
  jor  g16022(.dina(n14271), .dinb(n5694), .dout(n16166));
  jor  g16023(.dina(n11987), .dinb(n6208), .dout(n16167));
  jor  g16024(.dina(n11991), .dinb(n6132), .dout(n16168));
  jor  g16025(.dina(n11995), .dinb(n5692), .dout(n16169));
  jand g16026(.dina(n16169), .dinb(n16168), .dout(n16170));
  jand g16027(.dina(n16170), .dinb(n16167), .dout(n16171));
  jand g16028(.dina(n16171), .dinb(n16166), .dout(n16172));
  jxor g16029(.dina(n16172), .dinb(\a[20] ), .dout(n16173));
  jor  g16030(.dina(n16173), .dinb(n16165), .dout(n16174));
  jor  g16031(.dina(n14301), .dinb(n5694), .dout(n16175));
  jor  g16032(.dina(n11991), .dinb(n6208), .dout(n16176));
  jor  g16033(.dina(n11995), .dinb(n6132), .dout(n16177));
  jor  g16034(.dina(n11997), .dinb(n5692), .dout(n16178));
  jand g16035(.dina(n16178), .dinb(n16177), .dout(n16179));
  jand g16036(.dina(n16179), .dinb(n16176), .dout(n16180));
  jand g16037(.dina(n16180), .dinb(n16175), .dout(n16181));
  jxor g16038(.dina(n16181), .dinb(\a[20] ), .dout(n16182));
  jnot g16039(.din(n16182), .dout(n16183));
  jxor g16040(.dina(n15863), .dinb(n15862), .dout(n16184));
  jand g16041(.dina(n16184), .dinb(n16183), .dout(n16185));
  jor  g16042(.dina(n14353), .dinb(n5694), .dout(n16186));
  jor  g16043(.dina(n11995), .dinb(n6208), .dout(n16187));
  jor  g16044(.dina(n11997), .dinb(n6132), .dout(n16188));
  jor  g16045(.dina(n11999), .dinb(n5692), .dout(n16189));
  jand g16046(.dina(n16189), .dinb(n16188), .dout(n16190));
  jand g16047(.dina(n16190), .dinb(n16187), .dout(n16191));
  jand g16048(.dina(n16191), .dinb(n16186), .dout(n16192));
  jxor g16049(.dina(n16192), .dinb(\a[20] ), .dout(n16193));
  jnot g16050(.din(n16193), .dout(n16194));
  jxor g16051(.dina(n15860), .dinb(n15859), .dout(n16195));
  jand g16052(.dina(n16195), .dinb(n16194), .dout(n16196));
  jor  g16053(.dina(n14390), .dinb(n5694), .dout(n16197));
  jor  g16054(.dina(n11997), .dinb(n6208), .dout(n16198));
  jor  g16055(.dina(n11999), .dinb(n6132), .dout(n16199));
  jor  g16056(.dina(n12001), .dinb(n5692), .dout(n16200));
  jand g16057(.dina(n16200), .dinb(n16199), .dout(n16201));
  jand g16058(.dina(n16201), .dinb(n16198), .dout(n16202));
  jand g16059(.dina(n16202), .dinb(n16197), .dout(n16203));
  jxor g16060(.dina(n16203), .dinb(\a[20] ), .dout(n16204));
  jnot g16061(.din(n16204), .dout(n16205));
  jor  g16062(.dina(n15840), .dinb(n72), .dout(n16206));
  jxor g16063(.dina(n16206), .dinb(n15848), .dout(n16207));
  jand g16064(.dina(n16207), .dinb(n16205), .dout(n16208));
  jor  g16065(.dina(n14432), .dinb(n5694), .dout(n16209));
  jor  g16066(.dina(n11999), .dinb(n6208), .dout(n16210));
  jor  g16067(.dina(n12001), .dinb(n6132), .dout(n16211));
  jor  g16068(.dina(n12004), .dinb(n5692), .dout(n16212));
  jand g16069(.dina(n16212), .dinb(n16211), .dout(n16213));
  jand g16070(.dina(n16213), .dinb(n16210), .dout(n16214));
  jand g16071(.dina(n16214), .dinb(n16209), .dout(n16215));
  jxor g16072(.dina(n16215), .dinb(\a[20] ), .dout(n16216));
  jnot g16073(.din(n16216), .dout(n16217));
  jand g16074(.dina(n15837), .dinb(\a[23] ), .dout(n16218));
  jxor g16075(.dina(n16218), .dinb(n15835), .dout(n16219));
  jand g16076(.dina(n16219), .dinb(n16217), .dout(n16220));
  jand g16077(.dina(n14497), .dinb(n5693), .dout(n16221));
  jand g16078(.dina(n12010), .dinb(n6131), .dout(n16222));
  jand g16079(.dina(n12008), .dinb(n6209), .dout(n16223));
  jor  g16080(.dina(n16223), .dinb(n16222), .dout(n16224));
  jor  g16081(.dina(n16224), .dinb(n16221), .dout(n16225));
  jnot g16082(.din(n16225), .dout(n16226));
  jand g16083(.dina(n12010), .dinb(n5687), .dout(n16227));
  jnot g16084(.din(n16227), .dout(n16228));
  jand g16085(.dina(n16228), .dinb(\a[20] ), .dout(n16229));
  jand g16086(.dina(n16229), .dinb(n16226), .dout(n16230));
  jand g16087(.dina(n14537), .dinb(n5693), .dout(n16231));
  jand g16088(.dina(n12006), .dinb(n6209), .dout(n16232));
  jand g16089(.dina(n12008), .dinb(n6131), .dout(n16233));
  jand g16090(.dina(n12010), .dinb(n5691), .dout(n16234));
  jor  g16091(.dina(n16234), .dinb(n16233), .dout(n16235));
  jor  g16092(.dina(n16235), .dinb(n16232), .dout(n16236));
  jor  g16093(.dina(n16236), .dinb(n16231), .dout(n16237));
  jnot g16094(.din(n16237), .dout(n16238));
  jand g16095(.dina(n16238), .dinb(n16230), .dout(n16239));
  jand g16096(.dina(n16239), .dinb(n15837), .dout(n16240));
  jor  g16097(.dina(n15144), .dinb(n5694), .dout(n16241));
  jor  g16098(.dina(n12001), .dinb(n6208), .dout(n16242));
  jor  g16099(.dina(n12004), .dinb(n6132), .dout(n16243));
  jor  g16100(.dina(n12009), .dinb(n5692), .dout(n16244));
  jand g16101(.dina(n16244), .dinb(n16243), .dout(n16245));
  jand g16102(.dina(n16245), .dinb(n16242), .dout(n16246));
  jand g16103(.dina(n16246), .dinb(n16241), .dout(n16247));
  jxor g16104(.dina(n16247), .dinb(\a[20] ), .dout(n16248));
  jnot g16105(.din(n16248), .dout(n16249));
  jxor g16106(.dina(n16239), .dinb(n15837), .dout(n16250));
  jand g16107(.dina(n16250), .dinb(n16249), .dout(n16251));
  jor  g16108(.dina(n16251), .dinb(n16240), .dout(n16252));
  jxor g16109(.dina(n16219), .dinb(n16217), .dout(n16253));
  jand g16110(.dina(n16253), .dinb(n16252), .dout(n16254));
  jor  g16111(.dina(n16254), .dinb(n16220), .dout(n16255));
  jxor g16112(.dina(n16207), .dinb(n16205), .dout(n16256));
  jand g16113(.dina(n16256), .dinb(n16255), .dout(n16257));
  jor  g16114(.dina(n16257), .dinb(n16208), .dout(n16258));
  jxor g16115(.dina(n16195), .dinb(n16194), .dout(n16259));
  jand g16116(.dina(n16259), .dinb(n16258), .dout(n16260));
  jor  g16117(.dina(n16260), .dinb(n16196), .dout(n16261));
  jxor g16118(.dina(n16184), .dinb(n16183), .dout(n16262));
  jand g16119(.dina(n16262), .dinb(n16261), .dout(n16263));
  jor  g16120(.dina(n16263), .dinb(n16185), .dout(n16264));
  jxor g16121(.dina(n16173), .dinb(n16165), .dout(n16265));
  jand g16122(.dina(n16265), .dinb(n16264), .dout(n16266));
  jnot g16123(.din(n16266), .dout(n16267));
  jand g16124(.dina(n16267), .dinb(n16174), .dout(n16268));
  jnot g16125(.din(n16268), .dout(n16269));
  jxor g16126(.dina(n16162), .dinb(n16154), .dout(n16270));
  jand g16127(.dina(n16270), .dinb(n16269), .dout(n16271));
  jnot g16128(.din(n16271), .dout(n16272));
  jand g16129(.dina(n16272), .dinb(n16163), .dout(n16273));
  jnot g16130(.din(n16273), .dout(n16274));
  jxor g16131(.dina(n16151), .dinb(n16143), .dout(n16275));
  jand g16132(.dina(n16275), .dinb(n16274), .dout(n16276));
  jnot g16133(.din(n16276), .dout(n16277));
  jand g16134(.dina(n16277), .dinb(n16152), .dout(n16278));
  jnot g16135(.din(n16278), .dout(n16279));
  jxor g16136(.dina(n16140), .dinb(n16139), .dout(n16280));
  jand g16137(.dina(n16280), .dinb(n16279), .dout(n16281));
  jor  g16138(.dina(n16281), .dinb(n16141), .dout(n16282));
  jxor g16139(.dina(n16129), .dinb(n16128), .dout(n16283));
  jand g16140(.dina(n16283), .dinb(n16282), .dout(n16284));
  jor  g16141(.dina(n16284), .dinb(n16130), .dout(n16285));
  jxor g16142(.dina(n16118), .dinb(n16110), .dout(n16286));
  jand g16143(.dina(n16286), .dinb(n16285), .dout(n16287));
  jnot g16144(.din(n16287), .dout(n16288));
  jand g16145(.dina(n16288), .dinb(n16119), .dout(n16289));
  jnot g16146(.din(n16289), .dout(n16290));
  jxor g16147(.dina(n16107), .dinb(n16099), .dout(n16291));
  jand g16148(.dina(n16291), .dinb(n16290), .dout(n16292));
  jnot g16149(.din(n16292), .dout(n16293));
  jand g16150(.dina(n16293), .dinb(n16108), .dout(n16294));
  jnot g16151(.din(n16294), .dout(n16295));
  jxor g16152(.dina(n16096), .dinb(n16088), .dout(n16296));
  jand g16153(.dina(n16296), .dinb(n16295), .dout(n16297));
  jnot g16154(.din(n16297), .dout(n16298));
  jand g16155(.dina(n16298), .dinb(n16097), .dout(n16299));
  jnot g16156(.din(n16299), .dout(n16300));
  jxor g16157(.dina(n16085), .dinb(n16077), .dout(n16301));
  jand g16158(.dina(n16301), .dinb(n16300), .dout(n16302));
  jnot g16159(.din(n16302), .dout(n16303));
  jand g16160(.dina(n16303), .dinb(n16086), .dout(n16304));
  jnot g16161(.din(n16304), .dout(n16305));
  jxor g16162(.dina(n16074), .dinb(n16066), .dout(n16306));
  jand g16163(.dina(n16306), .dinb(n16305), .dout(n16307));
  jnot g16164(.din(n16307), .dout(n16308));
  jand g16165(.dina(n16308), .dinb(n16075), .dout(n16309));
  jnot g16166(.din(n16309), .dout(n16310));
  jxor g16167(.dina(n16063), .dinb(n16055), .dout(n16311));
  jand g16168(.dina(n16311), .dinb(n16310), .dout(n16312));
  jnot g16169(.din(n16312), .dout(n16313));
  jand g16170(.dina(n16313), .dinb(n16064), .dout(n16314));
  jnot g16171(.din(n16314), .dout(n16315));
  jxor g16172(.dina(n16052), .dinb(n16044), .dout(n16316));
  jand g16173(.dina(n16316), .dinb(n16315), .dout(n16317));
  jnot g16174(.din(n16317), .dout(n16318));
  jand g16175(.dina(n16318), .dinb(n16053), .dout(n16319));
  jnot g16176(.din(n16319), .dout(n16320));
  jxor g16177(.dina(n16041), .dinb(n16033), .dout(n16321));
  jand g16178(.dina(n16321), .dinb(n16320), .dout(n16322));
  jnot g16179(.din(n16322), .dout(n16323));
  jand g16180(.dina(n16323), .dinb(n16042), .dout(n16324));
  jnot g16181(.din(n16324), .dout(n16325));
  jxor g16182(.dina(n16030), .dinb(n16022), .dout(n16326));
  jand g16183(.dina(n16326), .dinb(n16325), .dout(n16327));
  jnot g16184(.din(n16327), .dout(n16328));
  jand g16185(.dina(n16328), .dinb(n16031), .dout(n16329));
  jnot g16186(.din(n16329), .dout(n16330));
  jxor g16187(.dina(n16019), .dinb(n16011), .dout(n16331));
  jand g16188(.dina(n16331), .dinb(n16330), .dout(n16332));
  jnot g16189(.din(n16332), .dout(n16333));
  jand g16190(.dina(n16333), .dinb(n16020), .dout(n16334));
  jnot g16191(.din(n16334), .dout(n16335));
  jxor g16192(.dina(n15927), .dinb(n15919), .dout(n16336));
  jand g16193(.dina(n16336), .dinb(n16335), .dout(n16337));
  jnot g16194(.din(n16337), .dout(n16338));
  jxor g16195(.dina(n16336), .dinb(n16335), .dout(n16339));
  jnot g16196(.din(n16339), .dout(n16340));
  jand g16197(.dina(n12569), .dinb(n6340), .dout(n16341));
  jand g16198(.dina(n11950), .dinb(n6798), .dout(n16342));
  jand g16199(.dina(n11952), .dinb(n6556), .dout(n16343));
  jand g16200(.dina(n11954), .dinb(n6338), .dout(n16344));
  jor  g16201(.dina(n16344), .dinb(n16343), .dout(n16345));
  jor  g16202(.dina(n16345), .dinb(n16342), .dout(n16346));
  jor  g16203(.dina(n16346), .dinb(n16341), .dout(n16347));
  jxor g16204(.dina(n16347), .dinb(n5064), .dout(n16348));
  jor  g16205(.dina(n16348), .dinb(n16340), .dout(n16349));
  jand g16206(.dina(n16349), .dinb(n16338), .dout(n16350));
  jnot g16207(.din(n16350), .dout(n16351));
  jxor g16208(.dina(n15943), .dinb(n15935), .dout(n16352));
  jand g16209(.dina(n16352), .dinb(n16351), .dout(n16353));
  jnot g16210(.din(n16353), .dout(n16354));
  jxor g16211(.dina(n16352), .dinb(n16351), .dout(n16355));
  jnot g16212(.din(n16355), .dout(n16356));
  jand g16213(.dina(n12751), .dinb(n6936), .dout(n16357));
  jand g16214(.dina(n11942), .dinb(n7741), .dout(n16358));
  jand g16215(.dina(n11944), .dinb(n7613), .dout(n16359));
  jand g16216(.dina(n11946), .dinb(n6934), .dout(n16360));
  jor  g16217(.dina(n16360), .dinb(n16359), .dout(n16361));
  jor  g16218(.dina(n16361), .dinb(n16358), .dout(n16362));
  jor  g16219(.dina(n16362), .dinb(n16357), .dout(n16363));
  jxor g16220(.dina(n16363), .dinb(n5292), .dout(n16364));
  jor  g16221(.dina(n16364), .dinb(n16356), .dout(n16365));
  jand g16222(.dina(n16365), .dinb(n16354), .dout(n16366));
  jnot g16223(.din(n16366), .dout(n16367));
  jxor g16224(.dina(n15959), .dinb(n15951), .dout(n16368));
  jand g16225(.dina(n16368), .dinb(n16367), .dout(n16369));
  jnot g16226(.din(n16369), .dout(n16370));
  jxor g16227(.dina(n16368), .dinb(n16367), .dout(n16371));
  jnot g16228(.din(n16371), .dout(n16372));
  jand g16229(.dina(n12841), .dinb(n7890), .dout(n16373));
  jand g16230(.dina(n12783), .dinb(n8441), .dout(n16374));
  jand g16231(.dina(n12766), .dinb(n8154), .dout(n16375));
  jand g16232(.dina(n12177), .dinb(n7888), .dout(n16376));
  jor  g16233(.dina(n16376), .dinb(n16375), .dout(n16377));
  jor  g16234(.dina(n16377), .dinb(n16374), .dout(n16378));
  jor  g16235(.dina(n16378), .dinb(n16373), .dout(n16379));
  jxor g16236(.dina(n16379), .dinb(n5833), .dout(n16380));
  jor  g16237(.dina(n16380), .dinb(n16372), .dout(n16381));
  jand g16238(.dina(n16381), .dinb(n16370), .dout(n16382));
  jnot g16239(.din(n16382), .dout(n16383));
  jxor g16240(.dina(n16008), .dinb(n16000), .dout(n16384));
  jand g16241(.dina(n16384), .dinb(n16383), .dout(n16385));
  jnot g16242(.din(n16385), .dout(n16386));
  jand g16243(.dina(n16386), .dinb(n16009), .dout(n16387));
  jnot g16244(.din(n16387), .dout(n16388));
  jxor g16245(.dina(n15980), .dinb(n15972), .dout(n16389));
  jand g16246(.dina(n16389), .dinb(n16388), .dout(n16390));
  jnot g16247(.din(n16390), .dout(n16391));
  jxor g16248(.dina(n16389), .dinb(n16388), .dout(n16392));
  jnot g16249(.din(n16392), .dout(n16393));
  jor  g16250(.dina(n12814), .dinb(n8770), .dout(n16395));
  jand g16251(.dina(n15985), .dinb(n16395), .dout(n16399));
  jand g16252(.dina(n16399), .dinb(n8772), .dout(n16400));
  jxor g16253(.dina(n16400), .dinb(\a[8] ), .dout(n16401));
  jor  g16254(.dina(n16401), .dinb(n16393), .dout(n16402));
  jand g16255(.dina(n16402), .dinb(n16391), .dout(n16403));
  jnot g16256(.din(n16403), .dout(n16404));
  jxor g16257(.dina(n15992), .dinb(n15991), .dout(n16405));
  jand g16258(.dina(n16405), .dinb(n16404), .dout(n16406));
  jxor g16259(.dina(n16405), .dinb(n16404), .dout(n16407));
  jand g16260(.dina(n12510), .dinb(n6340), .dout(n16408));
  jand g16261(.dina(n11952), .dinb(n6798), .dout(n16409));
  jand g16262(.dina(n11954), .dinb(n6556), .dout(n16410));
  jand g16263(.dina(n11956), .dinb(n6338), .dout(n16411));
  jor  g16264(.dina(n16411), .dinb(n16410), .dout(n16412));
  jor  g16265(.dina(n16412), .dinb(n16409), .dout(n16413));
  jor  g16266(.dina(n16413), .dinb(n16408), .dout(n16414));
  jxor g16267(.dina(n16414), .dinb(n5064), .dout(n16415));
  jnot g16268(.din(n16415), .dout(n16416));
  jxor g16269(.dina(n16331), .dinb(n16330), .dout(n16417));
  jand g16270(.dina(n16417), .dinb(n16416), .dout(n16418));
  jand g16271(.dina(n12472), .dinb(n6340), .dout(n16419));
  jand g16272(.dina(n11954), .dinb(n6798), .dout(n16420));
  jand g16273(.dina(n11956), .dinb(n6556), .dout(n16421));
  jand g16274(.dina(n11958), .dinb(n6338), .dout(n16422));
  jor  g16275(.dina(n16422), .dinb(n16421), .dout(n16423));
  jor  g16276(.dina(n16423), .dinb(n16420), .dout(n16424));
  jor  g16277(.dina(n16424), .dinb(n16419), .dout(n16425));
  jxor g16278(.dina(n16425), .dinb(n5064), .dout(n16426));
  jnot g16279(.din(n16426), .dout(n16427));
  jxor g16280(.dina(n16326), .dinb(n16325), .dout(n16428));
  jand g16281(.dina(n16428), .dinb(n16427), .dout(n16429));
  jand g16282(.dina(n12639), .dinb(n6340), .dout(n16430));
  jand g16283(.dina(n11956), .dinb(n6798), .dout(n16431));
  jand g16284(.dina(n11958), .dinb(n6556), .dout(n16432));
  jand g16285(.dina(n11960), .dinb(n6338), .dout(n16433));
  jor  g16286(.dina(n16433), .dinb(n16432), .dout(n16434));
  jor  g16287(.dina(n16434), .dinb(n16431), .dout(n16435));
  jor  g16288(.dina(n16435), .dinb(n16430), .dout(n16436));
  jxor g16289(.dina(n16436), .dinb(n5064), .dout(n16437));
  jnot g16290(.din(n16437), .dout(n16438));
  jxor g16291(.dina(n16321), .dinb(n16320), .dout(n16439));
  jand g16292(.dina(n16439), .dinb(n16438), .dout(n16440));
  jand g16293(.dina(n12624), .dinb(n6340), .dout(n16441));
  jand g16294(.dina(n11958), .dinb(n6798), .dout(n16442));
  jand g16295(.dina(n11960), .dinb(n6556), .dout(n16443));
  jand g16296(.dina(n11962), .dinb(n6338), .dout(n16444));
  jor  g16297(.dina(n16444), .dinb(n16443), .dout(n16445));
  jor  g16298(.dina(n16445), .dinb(n16442), .dout(n16446));
  jor  g16299(.dina(n16446), .dinb(n16441), .dout(n16447));
  jxor g16300(.dina(n16447), .dinb(n5064), .dout(n16448));
  jnot g16301(.din(n16448), .dout(n16449));
  jxor g16302(.dina(n16316), .dinb(n16315), .dout(n16450));
  jand g16303(.dina(n16450), .dinb(n16449), .dout(n16451));
  jand g16304(.dina(n13116), .dinb(n6340), .dout(n16452));
  jand g16305(.dina(n11960), .dinb(n6798), .dout(n16453));
  jand g16306(.dina(n11962), .dinb(n6556), .dout(n16454));
  jand g16307(.dina(n11964), .dinb(n6338), .dout(n16455));
  jor  g16308(.dina(n16455), .dinb(n16454), .dout(n16456));
  jor  g16309(.dina(n16456), .dinb(n16453), .dout(n16457));
  jor  g16310(.dina(n16457), .dinb(n16452), .dout(n16458));
  jxor g16311(.dina(n16458), .dinb(n5064), .dout(n16459));
  jnot g16312(.din(n16459), .dout(n16460));
  jxor g16313(.dina(n16311), .dinb(n16310), .dout(n16461));
  jand g16314(.dina(n16461), .dinb(n16460), .dout(n16462));
  jand g16315(.dina(n13134), .dinb(n6340), .dout(n16463));
  jand g16316(.dina(n11962), .dinb(n6798), .dout(n16464));
  jand g16317(.dina(n11964), .dinb(n6556), .dout(n16465));
  jand g16318(.dina(n11966), .dinb(n6338), .dout(n16466));
  jor  g16319(.dina(n16466), .dinb(n16465), .dout(n16467));
  jor  g16320(.dina(n16467), .dinb(n16464), .dout(n16468));
  jor  g16321(.dina(n16468), .dinb(n16463), .dout(n16469));
  jxor g16322(.dina(n16469), .dinb(n5064), .dout(n16470));
  jnot g16323(.din(n16470), .dout(n16471));
  jxor g16324(.dina(n16306), .dinb(n16305), .dout(n16472));
  jand g16325(.dina(n16472), .dinb(n16471), .dout(n16473));
  jand g16326(.dina(n13470), .dinb(n6340), .dout(n16474));
  jand g16327(.dina(n11964), .dinb(n6798), .dout(n16475));
  jand g16328(.dina(n11966), .dinb(n6556), .dout(n16476));
  jand g16329(.dina(n11968), .dinb(n6338), .dout(n16477));
  jor  g16330(.dina(n16477), .dinb(n16476), .dout(n16478));
  jor  g16331(.dina(n16478), .dinb(n16475), .dout(n16479));
  jor  g16332(.dina(n16479), .dinb(n16474), .dout(n16480));
  jxor g16333(.dina(n16480), .dinb(n5064), .dout(n16481));
  jnot g16334(.din(n16481), .dout(n16482));
  jxor g16335(.dina(n16301), .dinb(n16300), .dout(n16483));
  jand g16336(.dina(n16483), .dinb(n16482), .dout(n16484));
  jand g16337(.dina(n13268), .dinb(n6340), .dout(n16485));
  jand g16338(.dina(n11966), .dinb(n6798), .dout(n16486));
  jand g16339(.dina(n11968), .dinb(n6556), .dout(n16487));
  jand g16340(.dina(n11970), .dinb(n6338), .dout(n16488));
  jor  g16341(.dina(n16488), .dinb(n16487), .dout(n16489));
  jor  g16342(.dina(n16489), .dinb(n16486), .dout(n16490));
  jor  g16343(.dina(n16490), .dinb(n16485), .dout(n16491));
  jxor g16344(.dina(n16491), .dinb(n5064), .dout(n16492));
  jnot g16345(.din(n16492), .dout(n16493));
  jxor g16346(.dina(n16296), .dinb(n16295), .dout(n16494));
  jand g16347(.dina(n16494), .dinb(n16493), .dout(n16495));
  jand g16348(.dina(n13682), .dinb(n6340), .dout(n16496));
  jand g16349(.dina(n11968), .dinb(n6798), .dout(n16497));
  jand g16350(.dina(n11970), .dinb(n6556), .dout(n16498));
  jand g16351(.dina(n11972), .dinb(n6338), .dout(n16499));
  jor  g16352(.dina(n16499), .dinb(n16498), .dout(n16500));
  jor  g16353(.dina(n16500), .dinb(n16497), .dout(n16501));
  jor  g16354(.dina(n16501), .dinb(n16496), .dout(n16502));
  jxor g16355(.dina(n16502), .dinb(n5064), .dout(n16503));
  jnot g16356(.din(n16503), .dout(n16504));
  jxor g16357(.dina(n16291), .dinb(n16290), .dout(n16505));
  jand g16358(.dina(n16505), .dinb(n16504), .dout(n16506));
  jand g16359(.dina(n13806), .dinb(n6340), .dout(n16507));
  jand g16360(.dina(n11970), .dinb(n6798), .dout(n16508));
  jand g16361(.dina(n11972), .dinb(n6556), .dout(n16509));
  jand g16362(.dina(n11974), .dinb(n6338), .dout(n16510));
  jor  g16363(.dina(n16510), .dinb(n16509), .dout(n16511));
  jor  g16364(.dina(n16511), .dinb(n16508), .dout(n16512));
  jor  g16365(.dina(n16512), .dinb(n16507), .dout(n16513));
  jxor g16366(.dina(n16513), .dinb(n5064), .dout(n16514));
  jnot g16367(.din(n16514), .dout(n16515));
  jxor g16368(.dina(n16286), .dinb(n16285), .dout(n16516));
  jand g16369(.dina(n16516), .dinb(n16515), .dout(n16517));
  jxor g16370(.dina(n16283), .dinb(n16282), .dout(n16518));
  jnot g16371(.din(n16518), .dout(n16519));
  jand g16372(.dina(n13664), .dinb(n6340), .dout(n16520));
  jand g16373(.dina(n11972), .dinb(n6798), .dout(n16521));
  jand g16374(.dina(n11974), .dinb(n6556), .dout(n16522));
  jand g16375(.dina(n11976), .dinb(n6338), .dout(n16523));
  jor  g16376(.dina(n16523), .dinb(n16522), .dout(n16524));
  jor  g16377(.dina(n16524), .dinb(n16521), .dout(n16525));
  jor  g16378(.dina(n16525), .dinb(n16520), .dout(n16526));
  jxor g16379(.dina(n16526), .dinb(n5064), .dout(n16527));
  jor  g16380(.dina(n16527), .dinb(n16519), .dout(n16528));
  jxor g16381(.dina(n16280), .dinb(n16279), .dout(n16529));
  jnot g16382(.din(n16529), .dout(n16530));
  jand g16383(.dina(n13924), .dinb(n6340), .dout(n16531));
  jand g16384(.dina(n11974), .dinb(n6798), .dout(n16532));
  jand g16385(.dina(n11976), .dinb(n6556), .dout(n16533));
  jand g16386(.dina(n11978), .dinb(n6338), .dout(n16534));
  jor  g16387(.dina(n16534), .dinb(n16533), .dout(n16535));
  jor  g16388(.dina(n16535), .dinb(n16532), .dout(n16536));
  jor  g16389(.dina(n16536), .dinb(n16531), .dout(n16537));
  jxor g16390(.dina(n16537), .dinb(n5064), .dout(n16538));
  jor  g16391(.dina(n16538), .dinb(n16530), .dout(n16539));
  jand g16392(.dina(n14184), .dinb(n6340), .dout(n16540));
  jand g16393(.dina(n11976), .dinb(n6798), .dout(n16541));
  jand g16394(.dina(n11978), .dinb(n6556), .dout(n16542));
  jand g16395(.dina(n11980), .dinb(n6338), .dout(n16543));
  jor  g16396(.dina(n16543), .dinb(n16542), .dout(n16544));
  jor  g16397(.dina(n16544), .dinb(n16541), .dout(n16545));
  jor  g16398(.dina(n16545), .dinb(n16540), .dout(n16546));
  jxor g16399(.dina(n16546), .dinb(n5064), .dout(n16547));
  jnot g16400(.din(n16547), .dout(n16548));
  jxor g16401(.dina(n16275), .dinb(n16274), .dout(n16549));
  jand g16402(.dina(n16549), .dinb(n16548), .dout(n16550));
  jand g16403(.dina(n14194), .dinb(n6340), .dout(n16551));
  jand g16404(.dina(n11978), .dinb(n6798), .dout(n16552));
  jand g16405(.dina(n11980), .dinb(n6556), .dout(n16553));
  jand g16406(.dina(n11982), .dinb(n6338), .dout(n16554));
  jor  g16407(.dina(n16554), .dinb(n16553), .dout(n16555));
  jor  g16408(.dina(n16555), .dinb(n16552), .dout(n16556));
  jor  g16409(.dina(n16556), .dinb(n16551), .dout(n16557));
  jxor g16410(.dina(n16557), .dinb(n5064), .dout(n16558));
  jnot g16411(.din(n16558), .dout(n16559));
  jxor g16412(.dina(n16270), .dinb(n16269), .dout(n16560));
  jand g16413(.dina(n16560), .dinb(n16559), .dout(n16561));
  jand g16414(.dina(n13899), .dinb(n6340), .dout(n16562));
  jand g16415(.dina(n11980), .dinb(n6798), .dout(n16563));
  jand g16416(.dina(n11982), .dinb(n6556), .dout(n16564));
  jand g16417(.dina(n11985), .dinb(n6338), .dout(n16565));
  jor  g16418(.dina(n16565), .dinb(n16564), .dout(n16566));
  jor  g16419(.dina(n16566), .dinb(n16563), .dout(n16567));
  jor  g16420(.dina(n16567), .dinb(n16562), .dout(n16568));
  jxor g16421(.dina(n16568), .dinb(n5064), .dout(n16569));
  jnot g16422(.din(n16569), .dout(n16570));
  jxor g16423(.dina(n16265), .dinb(n16264), .dout(n16571));
  jand g16424(.dina(n16571), .dinb(n16570), .dout(n16572));
  jxor g16425(.dina(n16262), .dinb(n16261), .dout(n16573));
  jnot g16426(.din(n16573), .dout(n16574));
  jor  g16427(.dina(n14221), .dinb(n6341), .dout(n16575));
  jor  g16428(.dina(n15045), .dinb(n6797), .dout(n16576));
  jor  g16429(.dina(n11984), .dinb(n6557), .dout(n16577));
  jor  g16430(.dina(n11987), .dinb(n6339), .dout(n16578));
  jand g16431(.dina(n16578), .dinb(n16577), .dout(n16579));
  jand g16432(.dina(n16579), .dinb(n16576), .dout(n16580));
  jand g16433(.dina(n16580), .dinb(n16575), .dout(n16581));
  jxor g16434(.dina(n16581), .dinb(\a[17] ), .dout(n16582));
  jor  g16435(.dina(n16582), .dinb(n16574), .dout(n16583));
  jxor g16436(.dina(n16259), .dinb(n16258), .dout(n16584));
  jnot g16437(.din(n16584), .dout(n16585));
  jor  g16438(.dina(n14248), .dinb(n6341), .dout(n16586));
  jor  g16439(.dina(n11984), .dinb(n6797), .dout(n16587));
  jor  g16440(.dina(n11987), .dinb(n6557), .dout(n16588));
  jor  g16441(.dina(n11991), .dinb(n6339), .dout(n16589));
  jand g16442(.dina(n16589), .dinb(n16588), .dout(n16590));
  jand g16443(.dina(n16590), .dinb(n16587), .dout(n16591));
  jand g16444(.dina(n16591), .dinb(n16586), .dout(n16592));
  jxor g16445(.dina(n16592), .dinb(\a[17] ), .dout(n16593));
  jor  g16446(.dina(n16593), .dinb(n16585), .dout(n16594));
  jxor g16447(.dina(n16256), .dinb(n16255), .dout(n16595));
  jnot g16448(.din(n16595), .dout(n16596));
  jor  g16449(.dina(n14271), .dinb(n6341), .dout(n16597));
  jor  g16450(.dina(n11987), .dinb(n6797), .dout(n16598));
  jor  g16451(.dina(n11991), .dinb(n6557), .dout(n16599));
  jor  g16452(.dina(n11995), .dinb(n6339), .dout(n16600));
  jand g16453(.dina(n16600), .dinb(n16599), .dout(n16601));
  jand g16454(.dina(n16601), .dinb(n16598), .dout(n16602));
  jand g16455(.dina(n16602), .dinb(n16597), .dout(n16603));
  jxor g16456(.dina(n16603), .dinb(\a[17] ), .dout(n16604));
  jor  g16457(.dina(n16604), .dinb(n16596), .dout(n16605));
  jor  g16458(.dina(n14301), .dinb(n6341), .dout(n16606));
  jor  g16459(.dina(n11991), .dinb(n6797), .dout(n16607));
  jor  g16460(.dina(n11995), .dinb(n6557), .dout(n16608));
  jor  g16461(.dina(n11997), .dinb(n6339), .dout(n16609));
  jand g16462(.dina(n16609), .dinb(n16608), .dout(n16610));
  jand g16463(.dina(n16610), .dinb(n16607), .dout(n16611));
  jand g16464(.dina(n16611), .dinb(n16606), .dout(n16612));
  jxor g16465(.dina(n16612), .dinb(\a[17] ), .dout(n16613));
  jnot g16466(.din(n16613), .dout(n16614));
  jxor g16467(.dina(n16253), .dinb(n16252), .dout(n16615));
  jand g16468(.dina(n16615), .dinb(n16614), .dout(n16616));
  jor  g16469(.dina(n14353), .dinb(n6341), .dout(n16617));
  jor  g16470(.dina(n11995), .dinb(n6797), .dout(n16618));
  jor  g16471(.dina(n11997), .dinb(n6557), .dout(n16619));
  jor  g16472(.dina(n11999), .dinb(n6339), .dout(n16620));
  jand g16473(.dina(n16620), .dinb(n16619), .dout(n16621));
  jand g16474(.dina(n16621), .dinb(n16618), .dout(n16622));
  jand g16475(.dina(n16622), .dinb(n16617), .dout(n16623));
  jxor g16476(.dina(n16623), .dinb(\a[17] ), .dout(n16624));
  jnot g16477(.din(n16624), .dout(n16625));
  jxor g16478(.dina(n16250), .dinb(n16249), .dout(n16626));
  jand g16479(.dina(n16626), .dinb(n16625), .dout(n16627));
  jor  g16480(.dina(n14390), .dinb(n6341), .dout(n16628));
  jor  g16481(.dina(n11997), .dinb(n6797), .dout(n16629));
  jor  g16482(.dina(n11999), .dinb(n6557), .dout(n16630));
  jor  g16483(.dina(n12001), .dinb(n6339), .dout(n16631));
  jand g16484(.dina(n16631), .dinb(n16630), .dout(n16632));
  jand g16485(.dina(n16632), .dinb(n16629), .dout(n16633));
  jand g16486(.dina(n16633), .dinb(n16628), .dout(n16634));
  jxor g16487(.dina(n16634), .dinb(\a[17] ), .dout(n16635));
  jnot g16488(.din(n16635), .dout(n16636));
  jor  g16489(.dina(n16230), .dinb(n4247), .dout(n16637));
  jxor g16490(.dina(n16637), .dinb(n16238), .dout(n16638));
  jand g16491(.dina(n16638), .dinb(n16636), .dout(n16639));
  jor  g16492(.dina(n14432), .dinb(n6341), .dout(n16640));
  jor  g16493(.dina(n11999), .dinb(n6797), .dout(n16641));
  jor  g16494(.dina(n12001), .dinb(n6557), .dout(n16642));
  jor  g16495(.dina(n12004), .dinb(n6339), .dout(n16643));
  jand g16496(.dina(n16643), .dinb(n16642), .dout(n16644));
  jand g16497(.dina(n16644), .dinb(n16641), .dout(n16645));
  jand g16498(.dina(n16645), .dinb(n16640), .dout(n16646));
  jxor g16499(.dina(n16646), .dinb(\a[17] ), .dout(n16647));
  jnot g16500(.din(n16647), .dout(n16648));
  jand g16501(.dina(n16227), .dinb(\a[20] ), .dout(n16649));
  jxor g16502(.dina(n16649), .dinb(n16225), .dout(n16650));
  jand g16503(.dina(n16650), .dinb(n16648), .dout(n16651));
  jand g16504(.dina(n14497), .dinb(n6340), .dout(n16652));
  jand g16505(.dina(n12010), .dinb(n6556), .dout(n16653));
  jand g16506(.dina(n12008), .dinb(n6798), .dout(n16654));
  jor  g16507(.dina(n16654), .dinb(n16653), .dout(n16655));
  jor  g16508(.dina(n16655), .dinb(n16652), .dout(n16656));
  jnot g16509(.din(n16656), .dout(n16657));
  jand g16510(.dina(n12010), .dinb(n6334), .dout(n16658));
  jnot g16511(.din(n16658), .dout(n16659));
  jand g16512(.dina(n16659), .dinb(\a[17] ), .dout(n16660));
  jand g16513(.dina(n16660), .dinb(n16657), .dout(n16661));
  jand g16514(.dina(n14537), .dinb(n6340), .dout(n16662));
  jand g16515(.dina(n12006), .dinb(n6798), .dout(n16663));
  jand g16516(.dina(n12008), .dinb(n6556), .dout(n16664));
  jand g16517(.dina(n12010), .dinb(n6338), .dout(n16665));
  jor  g16518(.dina(n16665), .dinb(n16664), .dout(n16666));
  jor  g16519(.dina(n16666), .dinb(n16663), .dout(n16667));
  jor  g16520(.dina(n16667), .dinb(n16662), .dout(n16668));
  jnot g16521(.din(n16668), .dout(n16669));
  jand g16522(.dina(n16669), .dinb(n16661), .dout(n16670));
  jand g16523(.dina(n16670), .dinb(n16227), .dout(n16671));
  jor  g16524(.dina(n15144), .dinb(n6341), .dout(n16672));
  jor  g16525(.dina(n12001), .dinb(n6797), .dout(n16673));
  jor  g16526(.dina(n12004), .dinb(n6557), .dout(n16674));
  jor  g16527(.dina(n12009), .dinb(n6339), .dout(n16675));
  jand g16528(.dina(n16675), .dinb(n16674), .dout(n16676));
  jand g16529(.dina(n16676), .dinb(n16673), .dout(n16677));
  jand g16530(.dina(n16677), .dinb(n16672), .dout(n16678));
  jxor g16531(.dina(n16678), .dinb(\a[17] ), .dout(n16679));
  jnot g16532(.din(n16679), .dout(n16680));
  jxor g16533(.dina(n16670), .dinb(n16227), .dout(n16681));
  jand g16534(.dina(n16681), .dinb(n16680), .dout(n16682));
  jor  g16535(.dina(n16682), .dinb(n16671), .dout(n16683));
  jxor g16536(.dina(n16650), .dinb(n16648), .dout(n16684));
  jand g16537(.dina(n16684), .dinb(n16683), .dout(n16685));
  jor  g16538(.dina(n16685), .dinb(n16651), .dout(n16686));
  jxor g16539(.dina(n16638), .dinb(n16636), .dout(n16687));
  jand g16540(.dina(n16687), .dinb(n16686), .dout(n16688));
  jor  g16541(.dina(n16688), .dinb(n16639), .dout(n16689));
  jxor g16542(.dina(n16626), .dinb(n16625), .dout(n16690));
  jand g16543(.dina(n16690), .dinb(n16689), .dout(n16691));
  jor  g16544(.dina(n16691), .dinb(n16627), .dout(n16692));
  jxor g16545(.dina(n16615), .dinb(n16614), .dout(n16693));
  jand g16546(.dina(n16693), .dinb(n16692), .dout(n16694));
  jor  g16547(.dina(n16694), .dinb(n16616), .dout(n16695));
  jxor g16548(.dina(n16604), .dinb(n16596), .dout(n16696));
  jand g16549(.dina(n16696), .dinb(n16695), .dout(n16697));
  jnot g16550(.din(n16697), .dout(n16698));
  jand g16551(.dina(n16698), .dinb(n16605), .dout(n16699));
  jnot g16552(.din(n16699), .dout(n16700));
  jxor g16553(.dina(n16593), .dinb(n16585), .dout(n16701));
  jand g16554(.dina(n16701), .dinb(n16700), .dout(n16702));
  jnot g16555(.din(n16702), .dout(n16703));
  jand g16556(.dina(n16703), .dinb(n16594), .dout(n16704));
  jnot g16557(.din(n16704), .dout(n16705));
  jxor g16558(.dina(n16582), .dinb(n16574), .dout(n16706));
  jand g16559(.dina(n16706), .dinb(n16705), .dout(n16707));
  jnot g16560(.din(n16707), .dout(n16708));
  jand g16561(.dina(n16708), .dinb(n16583), .dout(n16709));
  jnot g16562(.din(n16709), .dout(n16710));
  jxor g16563(.dina(n16571), .dinb(n16570), .dout(n16711));
  jand g16564(.dina(n16711), .dinb(n16710), .dout(n16712));
  jor  g16565(.dina(n16712), .dinb(n16572), .dout(n16713));
  jxor g16566(.dina(n16560), .dinb(n16559), .dout(n16714));
  jand g16567(.dina(n16714), .dinb(n16713), .dout(n16715));
  jor  g16568(.dina(n16715), .dinb(n16561), .dout(n16716));
  jxor g16569(.dina(n16549), .dinb(n16548), .dout(n16717));
  jand g16570(.dina(n16717), .dinb(n16716), .dout(n16718));
  jor  g16571(.dina(n16718), .dinb(n16550), .dout(n16719));
  jxor g16572(.dina(n16538), .dinb(n16530), .dout(n16720));
  jand g16573(.dina(n16720), .dinb(n16719), .dout(n16721));
  jnot g16574(.din(n16721), .dout(n16722));
  jand g16575(.dina(n16722), .dinb(n16539), .dout(n16723));
  jnot g16576(.din(n16723), .dout(n16724));
  jxor g16577(.dina(n16527), .dinb(n16519), .dout(n16725));
  jand g16578(.dina(n16725), .dinb(n16724), .dout(n16726));
  jnot g16579(.din(n16726), .dout(n16727));
  jand g16580(.dina(n16727), .dinb(n16528), .dout(n16728));
  jnot g16581(.din(n16728), .dout(n16729));
  jxor g16582(.dina(n16516), .dinb(n16515), .dout(n16730));
  jand g16583(.dina(n16730), .dinb(n16729), .dout(n16731));
  jor  g16584(.dina(n16731), .dinb(n16517), .dout(n16732));
  jxor g16585(.dina(n16505), .dinb(n16504), .dout(n16733));
  jand g16586(.dina(n16733), .dinb(n16732), .dout(n16734));
  jor  g16587(.dina(n16734), .dinb(n16506), .dout(n16735));
  jxor g16588(.dina(n16494), .dinb(n16493), .dout(n16736));
  jand g16589(.dina(n16736), .dinb(n16735), .dout(n16737));
  jor  g16590(.dina(n16737), .dinb(n16495), .dout(n16738));
  jxor g16591(.dina(n16483), .dinb(n16482), .dout(n16739));
  jand g16592(.dina(n16739), .dinb(n16738), .dout(n16740));
  jor  g16593(.dina(n16740), .dinb(n16484), .dout(n16741));
  jxor g16594(.dina(n16472), .dinb(n16471), .dout(n16742));
  jand g16595(.dina(n16742), .dinb(n16741), .dout(n16743));
  jor  g16596(.dina(n16743), .dinb(n16473), .dout(n16744));
  jxor g16597(.dina(n16461), .dinb(n16460), .dout(n16745));
  jand g16598(.dina(n16745), .dinb(n16744), .dout(n16746));
  jor  g16599(.dina(n16746), .dinb(n16462), .dout(n16747));
  jxor g16600(.dina(n16450), .dinb(n16449), .dout(n16748));
  jand g16601(.dina(n16748), .dinb(n16747), .dout(n16749));
  jor  g16602(.dina(n16749), .dinb(n16451), .dout(n16750));
  jxor g16603(.dina(n16439), .dinb(n16438), .dout(n16751));
  jand g16604(.dina(n16751), .dinb(n16750), .dout(n16752));
  jor  g16605(.dina(n16752), .dinb(n16440), .dout(n16753));
  jxor g16606(.dina(n16428), .dinb(n16427), .dout(n16754));
  jand g16607(.dina(n16754), .dinb(n16753), .dout(n16755));
  jor  g16608(.dina(n16755), .dinb(n16429), .dout(n16756));
  jxor g16609(.dina(n16417), .dinb(n16416), .dout(n16757));
  jand g16610(.dina(n16757), .dinb(n16756), .dout(n16758));
  jor  g16611(.dina(n16758), .dinb(n16418), .dout(n16759));
  jxor g16612(.dina(n16348), .dinb(n16340), .dout(n16760));
  jand g16613(.dina(n16760), .dinb(n16759), .dout(n16761));
  jnot g16614(.din(n16761), .dout(n16762));
  jxor g16615(.dina(n16760), .dinb(n16759), .dout(n16763));
  jnot g16616(.din(n16763), .dout(n16764));
  jand g16617(.dina(n12189), .dinb(n6936), .dout(n16765));
  jand g16618(.dina(n11944), .dinb(n7741), .dout(n16766));
  jand g16619(.dina(n11946), .dinb(n7613), .dout(n16767));
  jand g16620(.dina(n11948), .dinb(n6934), .dout(n16768));
  jor  g16621(.dina(n16768), .dinb(n16767), .dout(n16769));
  jor  g16622(.dina(n16769), .dinb(n16766), .dout(n16770));
  jor  g16623(.dina(n16770), .dinb(n16765), .dout(n16771));
  jxor g16624(.dina(n16771), .dinb(n5292), .dout(n16772));
  jor  g16625(.dina(n16772), .dinb(n16764), .dout(n16773));
  jand g16626(.dina(n16773), .dinb(n16762), .dout(n16774));
  jnot g16627(.din(n16774), .dout(n16775));
  jxor g16628(.dina(n16364), .dinb(n16356), .dout(n16776));
  jand g16629(.dina(n16776), .dinb(n16775), .dout(n16777));
  jnot g16630(.din(n16777), .dout(n16778));
  jxor g16631(.dina(n16776), .dinb(n16775), .dout(n16779));
  jnot g16632(.din(n16779), .dout(n16780));
  jand g16633(.dina(n12768), .dinb(n7890), .dout(n16781));
  jand g16634(.dina(n12766), .dinb(n8441), .dout(n16782));
  jand g16635(.dina(n12177), .dinb(n8154), .dout(n16783));
  jand g16636(.dina(n11941), .dinb(n7888), .dout(n16784));
  jor  g16637(.dina(n16784), .dinb(n16783), .dout(n16785));
  jor  g16638(.dina(n16785), .dinb(n16782), .dout(n16786));
  jor  g16639(.dina(n16786), .dinb(n16781), .dout(n16787));
  jxor g16640(.dina(n16787), .dinb(n5833), .dout(n16788));
  jor  g16641(.dina(n16788), .dinb(n16780), .dout(n16789));
  jand g16642(.dina(n16789), .dinb(n16778), .dout(n16790));
  jnot g16643(.din(n16790), .dout(n16791));
  jxor g16644(.dina(n16380), .dinb(n16372), .dout(n16792));
  jand g16645(.dina(n16792), .dinb(n16791), .dout(n16793));
  jnot g16646(.din(n16793), .dout(n16794));
  jxor g16647(.dina(n16792), .dinb(n16791), .dout(n16795));
  jnot g16648(.din(n16795), .dout(n16796));
  jand g16649(.dina(n12919), .dinb(n8771), .dout(n16797));
  jand g16650(.dina(n12815), .dinb(n9491), .dout(n16798));
  jand g16651(.dina(n12795), .dinb(n9126), .dout(n16799));
  jand g16652(.dina(n12782), .dinb(n8769), .dout(n16800));
  jor  g16653(.dina(n16800), .dinb(n16799), .dout(n16801));
  jor  g16654(.dina(n16801), .dinb(n16798), .dout(n16802));
  jor  g16655(.dina(n16802), .dinb(n16797), .dout(n16803));
  jxor g16656(.dina(n16803), .dinb(n6039), .dout(n16804));
  jor  g16657(.dina(n16804), .dinb(n16796), .dout(n16805));
  jand g16658(.dina(n16805), .dinb(n16794), .dout(n16806));
  jand g16659(.dina(n13022), .dinb(n8771), .dout(n16807));
  jand g16660(.dina(n12815), .dinb(n9126), .dout(n16809));
  jand g16661(.dina(n12795), .dinb(n8769), .dout(n16810));
  jor  g16662(.dina(n16810), .dinb(n16809), .dout(n16811));
  jor  g16663(.dina(n16811), .dinb(n9491), .dout(n16812));
  jor  g16664(.dina(n16812), .dinb(n16807), .dout(n16813));
  jxor g16665(.dina(n16813), .dinb(n6039), .dout(n16814));
  jor  g16666(.dina(n16814), .dinb(n16806), .dout(n16815));
  jxor g16667(.dina(n16384), .dinb(n16383), .dout(n16816));
  jxor g16668(.dina(n16814), .dinb(n16806), .dout(n16817));
  jand g16669(.dina(n16817), .dinb(n16816), .dout(n16818));
  jnot g16670(.din(n16818), .dout(n16819));
  jand g16671(.dina(n16819), .dinb(n16815), .dout(n16820));
  jnot g16672(.din(n16820), .dout(n16821));
  jxor g16673(.dina(n16401), .dinb(n16393), .dout(n16822));
  jand g16674(.dina(n16822), .dinb(n16821), .dout(n16823));
  jxor g16675(.dina(n16757), .dinb(n16756), .dout(n16824));
  jnot g16676(.din(n16824), .dout(n16825));
  jand g16677(.dina(n12519), .dinb(n6936), .dout(n16826));
  jand g16678(.dina(n11946), .dinb(n7741), .dout(n16827));
  jand g16679(.dina(n11948), .dinb(n7613), .dout(n16828));
  jand g16680(.dina(n11950), .dinb(n6934), .dout(n16829));
  jor  g16681(.dina(n16829), .dinb(n16828), .dout(n16830));
  jor  g16682(.dina(n16830), .dinb(n16827), .dout(n16831));
  jor  g16683(.dina(n16831), .dinb(n16826), .dout(n16832));
  jxor g16684(.dina(n16832), .dinb(n5292), .dout(n16833));
  jor  g16685(.dina(n16833), .dinb(n16825), .dout(n16834));
  jxor g16686(.dina(n16754), .dinb(n16753), .dout(n16835));
  jnot g16687(.din(n16835), .dout(n16836));
  jand g16688(.dina(n12654), .dinb(n6936), .dout(n16837));
  jand g16689(.dina(n11948), .dinb(n7741), .dout(n16838));
  jand g16690(.dina(n11950), .dinb(n7613), .dout(n16839));
  jand g16691(.dina(n11952), .dinb(n6934), .dout(n16840));
  jor  g16692(.dina(n16840), .dinb(n16839), .dout(n16841));
  jor  g16693(.dina(n16841), .dinb(n16838), .dout(n16842));
  jor  g16694(.dina(n16842), .dinb(n16837), .dout(n16843));
  jxor g16695(.dina(n16843), .dinb(n5292), .dout(n16844));
  jor  g16696(.dina(n16844), .dinb(n16836), .dout(n16845));
  jxor g16697(.dina(n16751), .dinb(n16750), .dout(n16846));
  jnot g16698(.din(n16846), .dout(n16847));
  jand g16699(.dina(n12569), .dinb(n6936), .dout(n16848));
  jand g16700(.dina(n11950), .dinb(n7741), .dout(n16849));
  jand g16701(.dina(n11952), .dinb(n7613), .dout(n16850));
  jand g16702(.dina(n11954), .dinb(n6934), .dout(n16851));
  jor  g16703(.dina(n16851), .dinb(n16850), .dout(n16852));
  jor  g16704(.dina(n16852), .dinb(n16849), .dout(n16853));
  jor  g16705(.dina(n16853), .dinb(n16848), .dout(n16854));
  jxor g16706(.dina(n16854), .dinb(n5292), .dout(n16855));
  jor  g16707(.dina(n16855), .dinb(n16847), .dout(n16856));
  jxor g16708(.dina(n16748), .dinb(n16747), .dout(n16857));
  jnot g16709(.din(n16857), .dout(n16858));
  jand g16710(.dina(n12510), .dinb(n6936), .dout(n16859));
  jand g16711(.dina(n11952), .dinb(n7741), .dout(n16860));
  jand g16712(.dina(n11954), .dinb(n7613), .dout(n16861));
  jand g16713(.dina(n11956), .dinb(n6934), .dout(n16862));
  jor  g16714(.dina(n16862), .dinb(n16861), .dout(n16863));
  jor  g16715(.dina(n16863), .dinb(n16860), .dout(n16864));
  jor  g16716(.dina(n16864), .dinb(n16859), .dout(n16865));
  jxor g16717(.dina(n16865), .dinb(n5292), .dout(n16866));
  jor  g16718(.dina(n16866), .dinb(n16858), .dout(n16867));
  jxor g16719(.dina(n16745), .dinb(n16744), .dout(n16868));
  jnot g16720(.din(n16868), .dout(n16869));
  jand g16721(.dina(n12472), .dinb(n6936), .dout(n16870));
  jand g16722(.dina(n11954), .dinb(n7741), .dout(n16871));
  jand g16723(.dina(n11956), .dinb(n7613), .dout(n16872));
  jand g16724(.dina(n11958), .dinb(n6934), .dout(n16873));
  jor  g16725(.dina(n16873), .dinb(n16872), .dout(n16874));
  jor  g16726(.dina(n16874), .dinb(n16871), .dout(n16875));
  jor  g16727(.dina(n16875), .dinb(n16870), .dout(n16876));
  jxor g16728(.dina(n16876), .dinb(n5292), .dout(n16877));
  jor  g16729(.dina(n16877), .dinb(n16869), .dout(n16878));
  jxor g16730(.dina(n16742), .dinb(n16741), .dout(n16879));
  jnot g16731(.din(n16879), .dout(n16880));
  jand g16732(.dina(n12639), .dinb(n6936), .dout(n16881));
  jand g16733(.dina(n11956), .dinb(n7741), .dout(n16882));
  jand g16734(.dina(n11958), .dinb(n7613), .dout(n16883));
  jand g16735(.dina(n11960), .dinb(n6934), .dout(n16884));
  jor  g16736(.dina(n16884), .dinb(n16883), .dout(n16885));
  jor  g16737(.dina(n16885), .dinb(n16882), .dout(n16886));
  jor  g16738(.dina(n16886), .dinb(n16881), .dout(n16887));
  jxor g16739(.dina(n16887), .dinb(n5292), .dout(n16888));
  jor  g16740(.dina(n16888), .dinb(n16880), .dout(n16889));
  jxor g16741(.dina(n16739), .dinb(n16738), .dout(n16890));
  jnot g16742(.din(n16890), .dout(n16891));
  jand g16743(.dina(n12624), .dinb(n6936), .dout(n16892));
  jand g16744(.dina(n11958), .dinb(n7741), .dout(n16893));
  jand g16745(.dina(n11960), .dinb(n7613), .dout(n16894));
  jand g16746(.dina(n11962), .dinb(n6934), .dout(n16895));
  jor  g16747(.dina(n16895), .dinb(n16894), .dout(n16896));
  jor  g16748(.dina(n16896), .dinb(n16893), .dout(n16897));
  jor  g16749(.dina(n16897), .dinb(n16892), .dout(n16898));
  jxor g16750(.dina(n16898), .dinb(n5292), .dout(n16899));
  jor  g16751(.dina(n16899), .dinb(n16891), .dout(n16900));
  jxor g16752(.dina(n16736), .dinb(n16735), .dout(n16901));
  jnot g16753(.din(n16901), .dout(n16902));
  jand g16754(.dina(n13116), .dinb(n6936), .dout(n16903));
  jand g16755(.dina(n11960), .dinb(n7741), .dout(n16904));
  jand g16756(.dina(n11962), .dinb(n7613), .dout(n16905));
  jand g16757(.dina(n11964), .dinb(n6934), .dout(n16906));
  jor  g16758(.dina(n16906), .dinb(n16905), .dout(n16907));
  jor  g16759(.dina(n16907), .dinb(n16904), .dout(n16908));
  jor  g16760(.dina(n16908), .dinb(n16903), .dout(n16909));
  jxor g16761(.dina(n16909), .dinb(n5292), .dout(n16910));
  jor  g16762(.dina(n16910), .dinb(n16902), .dout(n16911));
  jxor g16763(.dina(n16733), .dinb(n16732), .dout(n16912));
  jnot g16764(.din(n16912), .dout(n16913));
  jand g16765(.dina(n13134), .dinb(n6936), .dout(n16914));
  jand g16766(.dina(n11962), .dinb(n7741), .dout(n16915));
  jand g16767(.dina(n11964), .dinb(n7613), .dout(n16916));
  jand g16768(.dina(n11966), .dinb(n6934), .dout(n16917));
  jor  g16769(.dina(n16917), .dinb(n16916), .dout(n16918));
  jor  g16770(.dina(n16918), .dinb(n16915), .dout(n16919));
  jor  g16771(.dina(n16919), .dinb(n16914), .dout(n16920));
  jxor g16772(.dina(n16920), .dinb(n5292), .dout(n16921));
  jor  g16773(.dina(n16921), .dinb(n16913), .dout(n16922));
  jxor g16774(.dina(n16730), .dinb(n16729), .dout(n16923));
  jnot g16775(.din(n16923), .dout(n16924));
  jand g16776(.dina(n13470), .dinb(n6936), .dout(n16925));
  jand g16777(.dina(n11964), .dinb(n7741), .dout(n16926));
  jand g16778(.dina(n11966), .dinb(n7613), .dout(n16927));
  jand g16779(.dina(n11968), .dinb(n6934), .dout(n16928));
  jor  g16780(.dina(n16928), .dinb(n16927), .dout(n16929));
  jor  g16781(.dina(n16929), .dinb(n16926), .dout(n16930));
  jor  g16782(.dina(n16930), .dinb(n16925), .dout(n16931));
  jxor g16783(.dina(n16931), .dinb(n5292), .dout(n16932));
  jor  g16784(.dina(n16932), .dinb(n16924), .dout(n16933));
  jand g16785(.dina(n13268), .dinb(n6936), .dout(n16934));
  jand g16786(.dina(n11966), .dinb(n7741), .dout(n16935));
  jand g16787(.dina(n11968), .dinb(n7613), .dout(n16936));
  jand g16788(.dina(n11970), .dinb(n6934), .dout(n16937));
  jor  g16789(.dina(n16937), .dinb(n16936), .dout(n16938));
  jor  g16790(.dina(n16938), .dinb(n16935), .dout(n16939));
  jor  g16791(.dina(n16939), .dinb(n16934), .dout(n16940));
  jxor g16792(.dina(n16940), .dinb(n5292), .dout(n16941));
  jnot g16793(.din(n16941), .dout(n16942));
  jxor g16794(.dina(n16725), .dinb(n16724), .dout(n16943));
  jand g16795(.dina(n16943), .dinb(n16942), .dout(n16944));
  jand g16796(.dina(n13682), .dinb(n6936), .dout(n16945));
  jand g16797(.dina(n11968), .dinb(n7741), .dout(n16946));
  jand g16798(.dina(n11970), .dinb(n7613), .dout(n16947));
  jand g16799(.dina(n11972), .dinb(n6934), .dout(n16948));
  jor  g16800(.dina(n16948), .dinb(n16947), .dout(n16949));
  jor  g16801(.dina(n16949), .dinb(n16946), .dout(n16950));
  jor  g16802(.dina(n16950), .dinb(n16945), .dout(n16951));
  jxor g16803(.dina(n16951), .dinb(n5292), .dout(n16952));
  jnot g16804(.din(n16952), .dout(n16953));
  jxor g16805(.dina(n16720), .dinb(n16719), .dout(n16954));
  jand g16806(.dina(n16954), .dinb(n16953), .dout(n16955));
  jxor g16807(.dina(n16717), .dinb(n16716), .dout(n16956));
  jnot g16808(.din(n16956), .dout(n16957));
  jand g16809(.dina(n13806), .dinb(n6936), .dout(n16958));
  jand g16810(.dina(n11970), .dinb(n7741), .dout(n16959));
  jand g16811(.dina(n11972), .dinb(n7613), .dout(n16960));
  jand g16812(.dina(n11974), .dinb(n6934), .dout(n16961));
  jor  g16813(.dina(n16961), .dinb(n16960), .dout(n16962));
  jor  g16814(.dina(n16962), .dinb(n16959), .dout(n16963));
  jor  g16815(.dina(n16963), .dinb(n16958), .dout(n16964));
  jxor g16816(.dina(n16964), .dinb(n5292), .dout(n16965));
  jor  g16817(.dina(n16965), .dinb(n16957), .dout(n16966));
  jxor g16818(.dina(n16714), .dinb(n16713), .dout(n16967));
  jnot g16819(.din(n16967), .dout(n16968));
  jand g16820(.dina(n13664), .dinb(n6936), .dout(n16969));
  jand g16821(.dina(n11972), .dinb(n7741), .dout(n16970));
  jand g16822(.dina(n11974), .dinb(n7613), .dout(n16971));
  jand g16823(.dina(n11976), .dinb(n6934), .dout(n16972));
  jor  g16824(.dina(n16972), .dinb(n16971), .dout(n16973));
  jor  g16825(.dina(n16973), .dinb(n16970), .dout(n16974));
  jor  g16826(.dina(n16974), .dinb(n16969), .dout(n16975));
  jxor g16827(.dina(n16975), .dinb(n5292), .dout(n16976));
  jor  g16828(.dina(n16976), .dinb(n16968), .dout(n16977));
  jxor g16829(.dina(n16711), .dinb(n16710), .dout(n16978));
  jnot g16830(.din(n16978), .dout(n16979));
  jand g16831(.dina(n13924), .dinb(n6936), .dout(n16980));
  jand g16832(.dina(n11974), .dinb(n7741), .dout(n16981));
  jand g16833(.dina(n11976), .dinb(n7613), .dout(n16982));
  jand g16834(.dina(n11978), .dinb(n6934), .dout(n16983));
  jor  g16835(.dina(n16983), .dinb(n16982), .dout(n16984));
  jor  g16836(.dina(n16984), .dinb(n16981), .dout(n16985));
  jor  g16837(.dina(n16985), .dinb(n16980), .dout(n16986));
  jxor g16838(.dina(n16986), .dinb(n5292), .dout(n16987));
  jor  g16839(.dina(n16987), .dinb(n16979), .dout(n16988));
  jand g16840(.dina(n14184), .dinb(n6936), .dout(n16989));
  jand g16841(.dina(n11976), .dinb(n7741), .dout(n16990));
  jand g16842(.dina(n11978), .dinb(n7613), .dout(n16991));
  jand g16843(.dina(n11980), .dinb(n6934), .dout(n16992));
  jor  g16844(.dina(n16992), .dinb(n16991), .dout(n16993));
  jor  g16845(.dina(n16993), .dinb(n16990), .dout(n16994));
  jor  g16846(.dina(n16994), .dinb(n16989), .dout(n16995));
  jxor g16847(.dina(n16995), .dinb(n5292), .dout(n16996));
  jnot g16848(.din(n16996), .dout(n16997));
  jxor g16849(.dina(n16706), .dinb(n16705), .dout(n16998));
  jand g16850(.dina(n16998), .dinb(n16997), .dout(n16999));
  jand g16851(.dina(n14194), .dinb(n6936), .dout(n17000));
  jand g16852(.dina(n11978), .dinb(n7741), .dout(n17001));
  jand g16853(.dina(n11980), .dinb(n7613), .dout(n17002));
  jand g16854(.dina(n11982), .dinb(n6934), .dout(n17003));
  jor  g16855(.dina(n17003), .dinb(n17002), .dout(n17004));
  jor  g16856(.dina(n17004), .dinb(n17001), .dout(n17005));
  jor  g16857(.dina(n17005), .dinb(n17000), .dout(n17006));
  jxor g16858(.dina(n17006), .dinb(n5292), .dout(n17007));
  jnot g16859(.din(n17007), .dout(n17008));
  jxor g16860(.dina(n16701), .dinb(n16700), .dout(n17009));
  jand g16861(.dina(n17009), .dinb(n17008), .dout(n17010));
  jand g16862(.dina(n13899), .dinb(n6936), .dout(n17011));
  jand g16863(.dina(n11980), .dinb(n7741), .dout(n17012));
  jand g16864(.dina(n11982), .dinb(n7613), .dout(n17013));
  jand g16865(.dina(n11985), .dinb(n6934), .dout(n17014));
  jor  g16866(.dina(n17014), .dinb(n17013), .dout(n17015));
  jor  g16867(.dina(n17015), .dinb(n17012), .dout(n17016));
  jor  g16868(.dina(n17016), .dinb(n17011), .dout(n17017));
  jxor g16869(.dina(n17017), .dinb(n5292), .dout(n17018));
  jnot g16870(.din(n17018), .dout(n17019));
  jxor g16871(.dina(n16696), .dinb(n16695), .dout(n17020));
  jand g16872(.dina(n17020), .dinb(n17019), .dout(n17021));
  jxor g16873(.dina(n16693), .dinb(n16692), .dout(n17022));
  jnot g16874(.din(n17022), .dout(n17023));
  jor  g16875(.dina(n14221), .dinb(n6937), .dout(n17024));
  jor  g16876(.dina(n15045), .dinb(n7740), .dout(n17025));
  jor  g16877(.dina(n11984), .dinb(n7614), .dout(n17026));
  jor  g16878(.dina(n11987), .dinb(n6935), .dout(n17027));
  jand g16879(.dina(n17027), .dinb(n17026), .dout(n17028));
  jand g16880(.dina(n17028), .dinb(n17025), .dout(n17029));
  jand g16881(.dina(n17029), .dinb(n17024), .dout(n17030));
  jxor g16882(.dina(n17030), .dinb(\a[14] ), .dout(n17031));
  jor  g16883(.dina(n17031), .dinb(n17023), .dout(n17032));
  jxor g16884(.dina(n16690), .dinb(n16689), .dout(n17033));
  jnot g16885(.din(n17033), .dout(n17034));
  jor  g16886(.dina(n14248), .dinb(n6937), .dout(n17035));
  jor  g16887(.dina(n11984), .dinb(n7740), .dout(n17036));
  jor  g16888(.dina(n11987), .dinb(n7614), .dout(n17037));
  jor  g16889(.dina(n11991), .dinb(n6935), .dout(n17038));
  jand g16890(.dina(n17038), .dinb(n17037), .dout(n17039));
  jand g16891(.dina(n17039), .dinb(n17036), .dout(n17040));
  jand g16892(.dina(n17040), .dinb(n17035), .dout(n17041));
  jxor g16893(.dina(n17041), .dinb(\a[14] ), .dout(n17042));
  jor  g16894(.dina(n17042), .dinb(n17034), .dout(n17043));
  jxor g16895(.dina(n16687), .dinb(n16686), .dout(n17044));
  jnot g16896(.din(n17044), .dout(n17045));
  jor  g16897(.dina(n14271), .dinb(n6937), .dout(n17046));
  jor  g16898(.dina(n11987), .dinb(n7740), .dout(n17047));
  jor  g16899(.dina(n11991), .dinb(n7614), .dout(n17048));
  jor  g16900(.dina(n11995), .dinb(n6935), .dout(n17049));
  jand g16901(.dina(n17049), .dinb(n17048), .dout(n17050));
  jand g16902(.dina(n17050), .dinb(n17047), .dout(n17051));
  jand g16903(.dina(n17051), .dinb(n17046), .dout(n17052));
  jxor g16904(.dina(n17052), .dinb(\a[14] ), .dout(n17053));
  jor  g16905(.dina(n17053), .dinb(n17045), .dout(n17054));
  jor  g16906(.dina(n14301), .dinb(n6937), .dout(n17055));
  jor  g16907(.dina(n11991), .dinb(n7740), .dout(n17056));
  jor  g16908(.dina(n11995), .dinb(n7614), .dout(n17057));
  jor  g16909(.dina(n11997), .dinb(n6935), .dout(n17058));
  jand g16910(.dina(n17058), .dinb(n17057), .dout(n17059));
  jand g16911(.dina(n17059), .dinb(n17056), .dout(n17060));
  jand g16912(.dina(n17060), .dinb(n17055), .dout(n17061));
  jxor g16913(.dina(n17061), .dinb(\a[14] ), .dout(n17062));
  jnot g16914(.din(n17062), .dout(n17063));
  jxor g16915(.dina(n16684), .dinb(n16683), .dout(n17064));
  jand g16916(.dina(n17064), .dinb(n17063), .dout(n17065));
  jor  g16917(.dina(n14353), .dinb(n6937), .dout(n17066));
  jor  g16918(.dina(n11995), .dinb(n7740), .dout(n17067));
  jor  g16919(.dina(n11997), .dinb(n7614), .dout(n17068));
  jor  g16920(.dina(n11999), .dinb(n6935), .dout(n17069));
  jand g16921(.dina(n17069), .dinb(n17068), .dout(n17070));
  jand g16922(.dina(n17070), .dinb(n17067), .dout(n17071));
  jand g16923(.dina(n17071), .dinb(n17066), .dout(n17072));
  jxor g16924(.dina(n17072), .dinb(\a[14] ), .dout(n17073));
  jnot g16925(.din(n17073), .dout(n17074));
  jxor g16926(.dina(n16681), .dinb(n16680), .dout(n17075));
  jand g16927(.dina(n17075), .dinb(n17074), .dout(n17076));
  jor  g16928(.dina(n14390), .dinb(n6937), .dout(n17077));
  jor  g16929(.dina(n11997), .dinb(n7740), .dout(n17078));
  jor  g16930(.dina(n11999), .dinb(n7614), .dout(n17079));
  jor  g16931(.dina(n12001), .dinb(n6935), .dout(n17080));
  jand g16932(.dina(n17080), .dinb(n17079), .dout(n17081));
  jand g16933(.dina(n17081), .dinb(n17078), .dout(n17082));
  jand g16934(.dina(n17082), .dinb(n17077), .dout(n17083));
  jxor g16935(.dina(n17083), .dinb(\a[14] ), .dout(n17084));
  jnot g16936(.din(n17084), .dout(n17085));
  jor  g16937(.dina(n16661), .dinb(n5064), .dout(n17086));
  jxor g16938(.dina(n17086), .dinb(n16669), .dout(n17087));
  jand g16939(.dina(n17087), .dinb(n17085), .dout(n17088));
  jor  g16940(.dina(n14432), .dinb(n6937), .dout(n17089));
  jor  g16941(.dina(n11999), .dinb(n7740), .dout(n17090));
  jor  g16942(.dina(n12001), .dinb(n7614), .dout(n17091));
  jor  g16943(.dina(n12004), .dinb(n6935), .dout(n17092));
  jand g16944(.dina(n17092), .dinb(n17091), .dout(n17093));
  jand g16945(.dina(n17093), .dinb(n17090), .dout(n17094));
  jand g16946(.dina(n17094), .dinb(n17089), .dout(n17095));
  jxor g16947(.dina(n17095), .dinb(\a[14] ), .dout(n17096));
  jnot g16948(.din(n17096), .dout(n17097));
  jand g16949(.dina(n16658), .dinb(\a[17] ), .dout(n17098));
  jxor g16950(.dina(n17098), .dinb(n16656), .dout(n17099));
  jand g16951(.dina(n17099), .dinb(n17097), .dout(n17100));
  jand g16952(.dina(n14497), .dinb(n6936), .dout(n17101));
  jand g16953(.dina(n12010), .dinb(n7613), .dout(n17102));
  jand g16954(.dina(n12008), .dinb(n7741), .dout(n17103));
  jor  g16955(.dina(n17103), .dinb(n17102), .dout(n17104));
  jor  g16956(.dina(n17104), .dinb(n17101), .dout(n17105));
  jnot g16957(.din(n17105), .dout(n17106));
  jand g16958(.dina(n12010), .dinb(n6928), .dout(n17107));
  jnot g16959(.din(n17107), .dout(n17108));
  jand g16960(.dina(n17108), .dinb(\a[14] ), .dout(n17109));
  jand g16961(.dina(n17109), .dinb(n17106), .dout(n17110));
  jand g16962(.dina(n14537), .dinb(n6936), .dout(n17111));
  jand g16963(.dina(n12006), .dinb(n7741), .dout(n17112));
  jand g16964(.dina(n12008), .dinb(n7613), .dout(n17113));
  jand g16965(.dina(n12010), .dinb(n6934), .dout(n17114));
  jor  g16966(.dina(n17114), .dinb(n17113), .dout(n17115));
  jor  g16967(.dina(n17115), .dinb(n17112), .dout(n17116));
  jor  g16968(.dina(n17116), .dinb(n17111), .dout(n17117));
  jnot g16969(.din(n17117), .dout(n17118));
  jand g16970(.dina(n17118), .dinb(n17110), .dout(n17119));
  jand g16971(.dina(n17119), .dinb(n16658), .dout(n17120));
  jor  g16972(.dina(n15144), .dinb(n6937), .dout(n17121));
  jor  g16973(.dina(n12001), .dinb(n7740), .dout(n17122));
  jor  g16974(.dina(n12004), .dinb(n7614), .dout(n17123));
  jor  g16975(.dina(n12009), .dinb(n6935), .dout(n17124));
  jand g16976(.dina(n17124), .dinb(n17123), .dout(n17125));
  jand g16977(.dina(n17125), .dinb(n17122), .dout(n17126));
  jand g16978(.dina(n17126), .dinb(n17121), .dout(n17127));
  jxor g16979(.dina(n17127), .dinb(\a[14] ), .dout(n17128));
  jnot g16980(.din(n17128), .dout(n17129));
  jxor g16981(.dina(n17119), .dinb(n16658), .dout(n17130));
  jand g16982(.dina(n17130), .dinb(n17129), .dout(n17131));
  jor  g16983(.dina(n17131), .dinb(n17120), .dout(n17132));
  jxor g16984(.dina(n17099), .dinb(n17097), .dout(n17133));
  jand g16985(.dina(n17133), .dinb(n17132), .dout(n17134));
  jor  g16986(.dina(n17134), .dinb(n17100), .dout(n17135));
  jxor g16987(.dina(n17087), .dinb(n17085), .dout(n17136));
  jand g16988(.dina(n17136), .dinb(n17135), .dout(n17137));
  jor  g16989(.dina(n17137), .dinb(n17088), .dout(n17138));
  jxor g16990(.dina(n17075), .dinb(n17074), .dout(n17139));
  jand g16991(.dina(n17139), .dinb(n17138), .dout(n17140));
  jor  g16992(.dina(n17140), .dinb(n17076), .dout(n17141));
  jxor g16993(.dina(n17064), .dinb(n17063), .dout(n17142));
  jand g16994(.dina(n17142), .dinb(n17141), .dout(n17143));
  jor  g16995(.dina(n17143), .dinb(n17065), .dout(n17144));
  jxor g16996(.dina(n17053), .dinb(n17045), .dout(n17145));
  jand g16997(.dina(n17145), .dinb(n17144), .dout(n17146));
  jnot g16998(.din(n17146), .dout(n17147));
  jand g16999(.dina(n17147), .dinb(n17054), .dout(n17148));
  jnot g17000(.din(n17148), .dout(n17149));
  jxor g17001(.dina(n17042), .dinb(n17034), .dout(n17150));
  jand g17002(.dina(n17150), .dinb(n17149), .dout(n17151));
  jnot g17003(.din(n17151), .dout(n17152));
  jand g17004(.dina(n17152), .dinb(n17043), .dout(n17153));
  jnot g17005(.din(n17153), .dout(n17154));
  jxor g17006(.dina(n17031), .dinb(n17023), .dout(n17155));
  jand g17007(.dina(n17155), .dinb(n17154), .dout(n17156));
  jnot g17008(.din(n17156), .dout(n17157));
  jand g17009(.dina(n17157), .dinb(n17032), .dout(n17158));
  jnot g17010(.din(n17158), .dout(n17159));
  jxor g17011(.dina(n17020), .dinb(n17019), .dout(n17160));
  jand g17012(.dina(n17160), .dinb(n17159), .dout(n17161));
  jor  g17013(.dina(n17161), .dinb(n17021), .dout(n17162));
  jxor g17014(.dina(n17009), .dinb(n17008), .dout(n17163));
  jand g17015(.dina(n17163), .dinb(n17162), .dout(n17164));
  jor  g17016(.dina(n17164), .dinb(n17010), .dout(n17165));
  jxor g17017(.dina(n16998), .dinb(n16997), .dout(n17166));
  jand g17018(.dina(n17166), .dinb(n17165), .dout(n17167));
  jor  g17019(.dina(n17167), .dinb(n16999), .dout(n17168));
  jxor g17020(.dina(n16987), .dinb(n16979), .dout(n17169));
  jand g17021(.dina(n17169), .dinb(n17168), .dout(n17170));
  jnot g17022(.din(n17170), .dout(n17171));
  jand g17023(.dina(n17171), .dinb(n16988), .dout(n17172));
  jnot g17024(.din(n17172), .dout(n17173));
  jxor g17025(.dina(n16976), .dinb(n16968), .dout(n17174));
  jand g17026(.dina(n17174), .dinb(n17173), .dout(n17175));
  jnot g17027(.din(n17175), .dout(n17176));
  jand g17028(.dina(n17176), .dinb(n16977), .dout(n17177));
  jnot g17029(.din(n17177), .dout(n17178));
  jxor g17030(.dina(n16965), .dinb(n16957), .dout(n17179));
  jand g17031(.dina(n17179), .dinb(n17178), .dout(n17180));
  jnot g17032(.din(n17180), .dout(n17181));
  jand g17033(.dina(n17181), .dinb(n16966), .dout(n17182));
  jnot g17034(.din(n17182), .dout(n17183));
  jxor g17035(.dina(n16954), .dinb(n16953), .dout(n17184));
  jand g17036(.dina(n17184), .dinb(n17183), .dout(n17185));
  jor  g17037(.dina(n17185), .dinb(n16955), .dout(n17186));
  jxor g17038(.dina(n16943), .dinb(n16942), .dout(n17187));
  jand g17039(.dina(n17187), .dinb(n17186), .dout(n17188));
  jor  g17040(.dina(n17188), .dinb(n16944), .dout(n17189));
  jxor g17041(.dina(n16932), .dinb(n16924), .dout(n17190));
  jand g17042(.dina(n17190), .dinb(n17189), .dout(n17191));
  jnot g17043(.din(n17191), .dout(n17192));
  jand g17044(.dina(n17192), .dinb(n16933), .dout(n17193));
  jnot g17045(.din(n17193), .dout(n17194));
  jxor g17046(.dina(n16921), .dinb(n16913), .dout(n17195));
  jand g17047(.dina(n17195), .dinb(n17194), .dout(n17196));
  jnot g17048(.din(n17196), .dout(n17197));
  jand g17049(.dina(n17197), .dinb(n16922), .dout(n17198));
  jnot g17050(.din(n17198), .dout(n17199));
  jxor g17051(.dina(n16910), .dinb(n16902), .dout(n17200));
  jand g17052(.dina(n17200), .dinb(n17199), .dout(n17201));
  jnot g17053(.din(n17201), .dout(n17202));
  jand g17054(.dina(n17202), .dinb(n16911), .dout(n17203));
  jnot g17055(.din(n17203), .dout(n17204));
  jxor g17056(.dina(n16899), .dinb(n16891), .dout(n17205));
  jand g17057(.dina(n17205), .dinb(n17204), .dout(n17206));
  jnot g17058(.din(n17206), .dout(n17207));
  jand g17059(.dina(n17207), .dinb(n16900), .dout(n17208));
  jnot g17060(.din(n17208), .dout(n17209));
  jxor g17061(.dina(n16888), .dinb(n16880), .dout(n17210));
  jand g17062(.dina(n17210), .dinb(n17209), .dout(n17211));
  jnot g17063(.din(n17211), .dout(n17212));
  jand g17064(.dina(n17212), .dinb(n16889), .dout(n17213));
  jnot g17065(.din(n17213), .dout(n17214));
  jxor g17066(.dina(n16877), .dinb(n16869), .dout(n17215));
  jand g17067(.dina(n17215), .dinb(n17214), .dout(n17216));
  jnot g17068(.din(n17216), .dout(n17217));
  jand g17069(.dina(n17217), .dinb(n16878), .dout(n17218));
  jnot g17070(.din(n17218), .dout(n17219));
  jxor g17071(.dina(n16866), .dinb(n16858), .dout(n17220));
  jand g17072(.dina(n17220), .dinb(n17219), .dout(n17221));
  jnot g17073(.din(n17221), .dout(n17222));
  jand g17074(.dina(n17222), .dinb(n16867), .dout(n17223));
  jnot g17075(.din(n17223), .dout(n17224));
  jxor g17076(.dina(n16855), .dinb(n16847), .dout(n17225));
  jand g17077(.dina(n17225), .dinb(n17224), .dout(n17226));
  jnot g17078(.din(n17226), .dout(n17227));
  jand g17079(.dina(n17227), .dinb(n16856), .dout(n17228));
  jnot g17080(.din(n17228), .dout(n17229));
  jxor g17081(.dina(n16844), .dinb(n16836), .dout(n17230));
  jand g17082(.dina(n17230), .dinb(n17229), .dout(n17231));
  jnot g17083(.din(n17231), .dout(n17232));
  jand g17084(.dina(n17232), .dinb(n16845), .dout(n17233));
  jnot g17085(.din(n17233), .dout(n17234));
  jxor g17086(.dina(n16833), .dinb(n16825), .dout(n17235));
  jand g17087(.dina(n17235), .dinb(n17234), .dout(n17236));
  jnot g17088(.din(n17236), .dout(n17237));
  jand g17089(.dina(n17237), .dinb(n16834), .dout(n17238));
  jnot g17090(.din(n17238), .dout(n17239));
  jxor g17091(.dina(n16772), .dinb(n16764), .dout(n17240));
  jand g17092(.dina(n17240), .dinb(n17239), .dout(n17241));
  jnot g17093(.din(n17241), .dout(n17242));
  jxor g17094(.dina(n17240), .dinb(n17239), .dout(n17243));
  jnot g17095(.din(n17243), .dout(n17244));
  jand g17096(.dina(n12179), .dinb(n7890), .dout(n17245));
  jand g17097(.dina(n12177), .dinb(n8441), .dout(n17246));
  jand g17098(.dina(n11941), .dinb(n8154), .dout(n17247));
  jand g17099(.dina(n11942), .dinb(n7888), .dout(n17248));
  jor  g17100(.dina(n17248), .dinb(n17247), .dout(n17249));
  jor  g17101(.dina(n17249), .dinb(n17246), .dout(n17250));
  jor  g17102(.dina(n17250), .dinb(n17245), .dout(n17251));
  jxor g17103(.dina(n17251), .dinb(n5833), .dout(n17252));
  jor  g17104(.dina(n17252), .dinb(n17244), .dout(n17253));
  jand g17105(.dina(n17253), .dinb(n17242), .dout(n17254));
  jnot g17106(.din(n17254), .dout(n17255));
  jxor g17107(.dina(n16788), .dinb(n16780), .dout(n17256));
  jand g17108(.dina(n17256), .dinb(n17255), .dout(n17257));
  jnot g17109(.din(n17257), .dout(n17258));
  jxor g17110(.dina(n17256), .dinb(n17255), .dout(n17259));
  jnot g17111(.din(n17259), .dout(n17260));
  jand g17112(.dina(n12797), .dinb(n8771), .dout(n17261));
  jand g17113(.dina(n12795), .dinb(n9491), .dout(n17262));
  jand g17114(.dina(n12782), .dinb(n9126), .dout(n17263));
  jand g17115(.dina(n12783), .dinb(n8769), .dout(n17264));
  jor  g17116(.dina(n17264), .dinb(n17263), .dout(n17265));
  jor  g17117(.dina(n17265), .dinb(n17262), .dout(n17266));
  jor  g17118(.dina(n17266), .dinb(n17261), .dout(n17267));
  jxor g17119(.dina(n17267), .dinb(n6039), .dout(n17268));
  jor  g17120(.dina(n17268), .dinb(n17260), .dout(n17269));
  jand g17121(.dina(n17269), .dinb(n17258), .dout(n17270));
  jand g17122(.dina(n10826), .dinb(n10351), .dout(n17273));
  jor  g17123(.dina(n13658), .dinb(n17270), .dout(n17278));
  jxor g17124(.dina(n13658), .dinb(n17270), .dout(n17279));
  jxor g17125(.dina(n16804), .dinb(n16796), .dout(n17280));
  jand g17126(.dina(n17280), .dinb(n17279), .dout(n17281));
  jnot g17127(.din(n17281), .dout(n17282));
  jand g17128(.dina(n17282), .dinb(n17278), .dout(n17283));
  jnot g17129(.din(n17283), .dout(n17284));
  jxor g17130(.dina(n16817), .dinb(n16816), .dout(n17285));
  jand g17131(.dina(n17285), .dinb(n17284), .dout(n17286));
  jand g17132(.dina(n12671), .dinb(n7890), .dout(n17287));
  jand g17133(.dina(n11941), .dinb(n8441), .dout(n17288));
  jand g17134(.dina(n11942), .dinb(n8154), .dout(n17289));
  jand g17135(.dina(n11944), .dinb(n7888), .dout(n17290));
  jor  g17136(.dina(n17290), .dinb(n17289), .dout(n17291));
  jor  g17137(.dina(n17291), .dinb(n17288), .dout(n17292));
  jor  g17138(.dina(n17292), .dinb(n17287), .dout(n17293));
  jxor g17139(.dina(n17293), .dinb(n5833), .dout(n17294));
  jnot g17140(.din(n17294), .dout(n17295));
  jxor g17141(.dina(n17235), .dinb(n17234), .dout(n17296));
  jand g17142(.dina(n17296), .dinb(n17295), .dout(n17297));
  jand g17143(.dina(n12751), .dinb(n7890), .dout(n17298));
  jand g17144(.dina(n11942), .dinb(n8441), .dout(n17299));
  jand g17145(.dina(n11944), .dinb(n8154), .dout(n17300));
  jand g17146(.dina(n11946), .dinb(n7888), .dout(n17301));
  jor  g17147(.dina(n17301), .dinb(n17300), .dout(n17302));
  jor  g17148(.dina(n17302), .dinb(n17299), .dout(n17303));
  jor  g17149(.dina(n17303), .dinb(n17298), .dout(n17304));
  jxor g17150(.dina(n17304), .dinb(n5833), .dout(n17305));
  jnot g17151(.din(n17305), .dout(n17306));
  jxor g17152(.dina(n17230), .dinb(n17229), .dout(n17307));
  jand g17153(.dina(n17307), .dinb(n17306), .dout(n17308));
  jand g17154(.dina(n12189), .dinb(n7890), .dout(n17309));
  jand g17155(.dina(n11944), .dinb(n8441), .dout(n17310));
  jand g17156(.dina(n11946), .dinb(n8154), .dout(n17311));
  jand g17157(.dina(n11948), .dinb(n7888), .dout(n17312));
  jor  g17158(.dina(n17312), .dinb(n17311), .dout(n17313));
  jor  g17159(.dina(n17313), .dinb(n17310), .dout(n17314));
  jor  g17160(.dina(n17314), .dinb(n17309), .dout(n17315));
  jxor g17161(.dina(n17315), .dinb(n5833), .dout(n17316));
  jnot g17162(.din(n17316), .dout(n17317));
  jxor g17163(.dina(n17225), .dinb(n17224), .dout(n17318));
  jand g17164(.dina(n17318), .dinb(n17317), .dout(n17319));
  jand g17165(.dina(n12519), .dinb(n7890), .dout(n17320));
  jand g17166(.dina(n11946), .dinb(n8441), .dout(n17321));
  jand g17167(.dina(n11948), .dinb(n8154), .dout(n17322));
  jand g17168(.dina(n11950), .dinb(n7888), .dout(n17323));
  jor  g17169(.dina(n17323), .dinb(n17322), .dout(n17324));
  jor  g17170(.dina(n17324), .dinb(n17321), .dout(n17325));
  jor  g17171(.dina(n17325), .dinb(n17320), .dout(n17326));
  jxor g17172(.dina(n17326), .dinb(n5833), .dout(n17327));
  jnot g17173(.din(n17327), .dout(n17328));
  jxor g17174(.dina(n17220), .dinb(n17219), .dout(n17329));
  jand g17175(.dina(n17329), .dinb(n17328), .dout(n17330));
  jand g17176(.dina(n12654), .dinb(n7890), .dout(n17331));
  jand g17177(.dina(n11948), .dinb(n8441), .dout(n17332));
  jand g17178(.dina(n11950), .dinb(n8154), .dout(n17333));
  jand g17179(.dina(n11952), .dinb(n7888), .dout(n17334));
  jor  g17180(.dina(n17334), .dinb(n17333), .dout(n17335));
  jor  g17181(.dina(n17335), .dinb(n17332), .dout(n17336));
  jor  g17182(.dina(n17336), .dinb(n17331), .dout(n17337));
  jxor g17183(.dina(n17337), .dinb(n5833), .dout(n17338));
  jnot g17184(.din(n17338), .dout(n17339));
  jxor g17185(.dina(n17215), .dinb(n17214), .dout(n17340));
  jand g17186(.dina(n17340), .dinb(n17339), .dout(n17341));
  jand g17187(.dina(n12569), .dinb(n7890), .dout(n17342));
  jand g17188(.dina(n11950), .dinb(n8441), .dout(n17343));
  jand g17189(.dina(n11952), .dinb(n8154), .dout(n17344));
  jand g17190(.dina(n11954), .dinb(n7888), .dout(n17345));
  jor  g17191(.dina(n17345), .dinb(n17344), .dout(n17346));
  jor  g17192(.dina(n17346), .dinb(n17343), .dout(n17347));
  jor  g17193(.dina(n17347), .dinb(n17342), .dout(n17348));
  jxor g17194(.dina(n17348), .dinb(n5833), .dout(n17349));
  jnot g17195(.din(n17349), .dout(n17350));
  jxor g17196(.dina(n17210), .dinb(n17209), .dout(n17351));
  jand g17197(.dina(n17351), .dinb(n17350), .dout(n17352));
  jand g17198(.dina(n12510), .dinb(n7890), .dout(n17353));
  jand g17199(.dina(n11952), .dinb(n8441), .dout(n17354));
  jand g17200(.dina(n11954), .dinb(n8154), .dout(n17355));
  jand g17201(.dina(n11956), .dinb(n7888), .dout(n17356));
  jor  g17202(.dina(n17356), .dinb(n17355), .dout(n17357));
  jor  g17203(.dina(n17357), .dinb(n17354), .dout(n17358));
  jor  g17204(.dina(n17358), .dinb(n17353), .dout(n17359));
  jxor g17205(.dina(n17359), .dinb(n5833), .dout(n17360));
  jnot g17206(.din(n17360), .dout(n17361));
  jxor g17207(.dina(n17205), .dinb(n17204), .dout(n17362));
  jand g17208(.dina(n17362), .dinb(n17361), .dout(n17363));
  jand g17209(.dina(n12472), .dinb(n7890), .dout(n17364));
  jand g17210(.dina(n11954), .dinb(n8441), .dout(n17365));
  jand g17211(.dina(n11956), .dinb(n8154), .dout(n17366));
  jand g17212(.dina(n11958), .dinb(n7888), .dout(n17367));
  jor  g17213(.dina(n17367), .dinb(n17366), .dout(n17368));
  jor  g17214(.dina(n17368), .dinb(n17365), .dout(n17369));
  jor  g17215(.dina(n17369), .dinb(n17364), .dout(n17370));
  jxor g17216(.dina(n17370), .dinb(n5833), .dout(n17371));
  jnot g17217(.din(n17371), .dout(n17372));
  jxor g17218(.dina(n17200), .dinb(n17199), .dout(n17373));
  jand g17219(.dina(n17373), .dinb(n17372), .dout(n17374));
  jand g17220(.dina(n12639), .dinb(n7890), .dout(n17375));
  jand g17221(.dina(n11956), .dinb(n8441), .dout(n17376));
  jand g17222(.dina(n11958), .dinb(n8154), .dout(n17377));
  jand g17223(.dina(n11960), .dinb(n7888), .dout(n17378));
  jor  g17224(.dina(n17378), .dinb(n17377), .dout(n17379));
  jor  g17225(.dina(n17379), .dinb(n17376), .dout(n17380));
  jor  g17226(.dina(n17380), .dinb(n17375), .dout(n17381));
  jxor g17227(.dina(n17381), .dinb(n5833), .dout(n17382));
  jnot g17228(.din(n17382), .dout(n17383));
  jxor g17229(.dina(n17195), .dinb(n17194), .dout(n17384));
  jand g17230(.dina(n17384), .dinb(n17383), .dout(n17385));
  jand g17231(.dina(n12624), .dinb(n7890), .dout(n17386));
  jand g17232(.dina(n11958), .dinb(n8441), .dout(n17387));
  jand g17233(.dina(n11960), .dinb(n8154), .dout(n17388));
  jand g17234(.dina(n11962), .dinb(n7888), .dout(n17389));
  jor  g17235(.dina(n17389), .dinb(n17388), .dout(n17390));
  jor  g17236(.dina(n17390), .dinb(n17387), .dout(n17391));
  jor  g17237(.dina(n17391), .dinb(n17386), .dout(n17392));
  jxor g17238(.dina(n17392), .dinb(n5833), .dout(n17393));
  jnot g17239(.din(n17393), .dout(n17394));
  jxor g17240(.dina(n17190), .dinb(n17189), .dout(n17395));
  jand g17241(.dina(n17395), .dinb(n17394), .dout(n17396));
  jxor g17242(.dina(n17187), .dinb(n17186), .dout(n17397));
  jnot g17243(.din(n17397), .dout(n17398));
  jand g17244(.dina(n13116), .dinb(n7890), .dout(n17399));
  jand g17245(.dina(n11960), .dinb(n8441), .dout(n17400));
  jand g17246(.dina(n11962), .dinb(n8154), .dout(n17401));
  jand g17247(.dina(n11964), .dinb(n7888), .dout(n17402));
  jor  g17248(.dina(n17402), .dinb(n17401), .dout(n17403));
  jor  g17249(.dina(n17403), .dinb(n17400), .dout(n17404));
  jor  g17250(.dina(n17404), .dinb(n17399), .dout(n17405));
  jxor g17251(.dina(n17405), .dinb(n5833), .dout(n17406));
  jor  g17252(.dina(n17406), .dinb(n17398), .dout(n17407));
  jxor g17253(.dina(n17184), .dinb(n17183), .dout(n17408));
  jnot g17254(.din(n17408), .dout(n17409));
  jand g17255(.dina(n13134), .dinb(n7890), .dout(n17410));
  jand g17256(.dina(n11962), .dinb(n8441), .dout(n17411));
  jand g17257(.dina(n11964), .dinb(n8154), .dout(n17412));
  jand g17258(.dina(n11966), .dinb(n7888), .dout(n17413));
  jor  g17259(.dina(n17413), .dinb(n17412), .dout(n17414));
  jor  g17260(.dina(n17414), .dinb(n17411), .dout(n17415));
  jor  g17261(.dina(n17415), .dinb(n17410), .dout(n17416));
  jxor g17262(.dina(n17416), .dinb(n5833), .dout(n17417));
  jor  g17263(.dina(n17417), .dinb(n17409), .dout(n17418));
  jand g17264(.dina(n13470), .dinb(n7890), .dout(n17419));
  jand g17265(.dina(n11964), .dinb(n8441), .dout(n17420));
  jand g17266(.dina(n11966), .dinb(n8154), .dout(n17421));
  jand g17267(.dina(n11968), .dinb(n7888), .dout(n17422));
  jor  g17268(.dina(n17422), .dinb(n17421), .dout(n17423));
  jor  g17269(.dina(n17423), .dinb(n17420), .dout(n17424));
  jor  g17270(.dina(n17424), .dinb(n17419), .dout(n17425));
  jxor g17271(.dina(n17425), .dinb(n5833), .dout(n17426));
  jnot g17272(.din(n17426), .dout(n17427));
  jxor g17273(.dina(n17179), .dinb(n17178), .dout(n17428));
  jand g17274(.dina(n17428), .dinb(n17427), .dout(n17429));
  jand g17275(.dina(n13268), .dinb(n7890), .dout(n17430));
  jand g17276(.dina(n11966), .dinb(n8441), .dout(n17431));
  jand g17277(.dina(n11968), .dinb(n8154), .dout(n17432));
  jand g17278(.dina(n11970), .dinb(n7888), .dout(n17433));
  jor  g17279(.dina(n17433), .dinb(n17432), .dout(n17434));
  jor  g17280(.dina(n17434), .dinb(n17431), .dout(n17435));
  jor  g17281(.dina(n17435), .dinb(n17430), .dout(n17436));
  jxor g17282(.dina(n17436), .dinb(n5833), .dout(n17437));
  jnot g17283(.din(n17437), .dout(n17438));
  jxor g17284(.dina(n17174), .dinb(n17173), .dout(n17439));
  jand g17285(.dina(n17439), .dinb(n17438), .dout(n17440));
  jand g17286(.dina(n13682), .dinb(n7890), .dout(n17441));
  jand g17287(.dina(n11968), .dinb(n8441), .dout(n17442));
  jand g17288(.dina(n11970), .dinb(n8154), .dout(n17443));
  jand g17289(.dina(n11972), .dinb(n7888), .dout(n17444));
  jor  g17290(.dina(n17444), .dinb(n17443), .dout(n17445));
  jor  g17291(.dina(n17445), .dinb(n17442), .dout(n17446));
  jor  g17292(.dina(n17446), .dinb(n17441), .dout(n17447));
  jxor g17293(.dina(n17447), .dinb(n5833), .dout(n17448));
  jnot g17294(.din(n17448), .dout(n17449));
  jxor g17295(.dina(n17169), .dinb(n17168), .dout(n17450));
  jand g17296(.dina(n17450), .dinb(n17449), .dout(n17451));
  jxor g17297(.dina(n17166), .dinb(n17165), .dout(n17452));
  jnot g17298(.din(n17452), .dout(n17453));
  jand g17299(.dina(n13806), .dinb(n7890), .dout(n17454));
  jand g17300(.dina(n11970), .dinb(n8441), .dout(n17455));
  jand g17301(.dina(n11972), .dinb(n8154), .dout(n17456));
  jand g17302(.dina(n11974), .dinb(n7888), .dout(n17457));
  jor  g17303(.dina(n17457), .dinb(n17456), .dout(n17458));
  jor  g17304(.dina(n17458), .dinb(n17455), .dout(n17459));
  jor  g17305(.dina(n17459), .dinb(n17454), .dout(n17460));
  jxor g17306(.dina(n17460), .dinb(n5833), .dout(n17461));
  jor  g17307(.dina(n17461), .dinb(n17453), .dout(n17462));
  jxor g17308(.dina(n17163), .dinb(n17162), .dout(n17463));
  jnot g17309(.din(n17463), .dout(n17464));
  jand g17310(.dina(n13664), .dinb(n7890), .dout(n17465));
  jand g17311(.dina(n11972), .dinb(n8441), .dout(n17466));
  jand g17312(.dina(n11974), .dinb(n8154), .dout(n17467));
  jand g17313(.dina(n11976), .dinb(n7888), .dout(n17468));
  jor  g17314(.dina(n17468), .dinb(n17467), .dout(n17469));
  jor  g17315(.dina(n17469), .dinb(n17466), .dout(n17470));
  jor  g17316(.dina(n17470), .dinb(n17465), .dout(n17471));
  jxor g17317(.dina(n17471), .dinb(n5833), .dout(n17472));
  jor  g17318(.dina(n17472), .dinb(n17464), .dout(n17473));
  jxor g17319(.dina(n17160), .dinb(n17159), .dout(n17474));
  jnot g17320(.din(n17474), .dout(n17475));
  jand g17321(.dina(n13924), .dinb(n7890), .dout(n17476));
  jand g17322(.dina(n11974), .dinb(n8441), .dout(n17477));
  jand g17323(.dina(n11976), .dinb(n8154), .dout(n17478));
  jand g17324(.dina(n11978), .dinb(n7888), .dout(n17479));
  jor  g17325(.dina(n17479), .dinb(n17478), .dout(n17480));
  jor  g17326(.dina(n17480), .dinb(n17477), .dout(n17481));
  jor  g17327(.dina(n17481), .dinb(n17476), .dout(n17482));
  jxor g17328(.dina(n17482), .dinb(n5833), .dout(n17483));
  jor  g17329(.dina(n17483), .dinb(n17475), .dout(n17484));
  jand g17330(.dina(n14184), .dinb(n7890), .dout(n17485));
  jand g17331(.dina(n11976), .dinb(n8441), .dout(n17486));
  jand g17332(.dina(n11978), .dinb(n8154), .dout(n17487));
  jand g17333(.dina(n11980), .dinb(n7888), .dout(n17488));
  jor  g17334(.dina(n17488), .dinb(n17487), .dout(n17489));
  jor  g17335(.dina(n17489), .dinb(n17486), .dout(n17490));
  jor  g17336(.dina(n17490), .dinb(n17485), .dout(n17491));
  jxor g17337(.dina(n17491), .dinb(n5833), .dout(n17492));
  jnot g17338(.din(n17492), .dout(n17493));
  jxor g17339(.dina(n17155), .dinb(n17154), .dout(n17494));
  jand g17340(.dina(n17494), .dinb(n17493), .dout(n17495));
  jand g17341(.dina(n14194), .dinb(n7890), .dout(n17496));
  jand g17342(.dina(n11978), .dinb(n8441), .dout(n17497));
  jand g17343(.dina(n11980), .dinb(n8154), .dout(n17498));
  jand g17344(.dina(n11982), .dinb(n7888), .dout(n17499));
  jor  g17345(.dina(n17499), .dinb(n17498), .dout(n17500));
  jor  g17346(.dina(n17500), .dinb(n17497), .dout(n17501));
  jor  g17347(.dina(n17501), .dinb(n17496), .dout(n17502));
  jxor g17348(.dina(n17502), .dinb(n5833), .dout(n17503));
  jnot g17349(.din(n17503), .dout(n17504));
  jxor g17350(.dina(n17150), .dinb(n17149), .dout(n17505));
  jand g17351(.dina(n17505), .dinb(n17504), .dout(n17506));
  jand g17352(.dina(n13899), .dinb(n7890), .dout(n17507));
  jand g17353(.dina(n11980), .dinb(n8441), .dout(n17508));
  jand g17354(.dina(n11982), .dinb(n8154), .dout(n17509));
  jand g17355(.dina(n11985), .dinb(n7888), .dout(n17510));
  jor  g17356(.dina(n17510), .dinb(n17509), .dout(n17511));
  jor  g17357(.dina(n17511), .dinb(n17508), .dout(n17512));
  jor  g17358(.dina(n17512), .dinb(n17507), .dout(n17513));
  jxor g17359(.dina(n17513), .dinb(n5833), .dout(n17514));
  jnot g17360(.din(n17514), .dout(n17515));
  jxor g17361(.dina(n17145), .dinb(n17144), .dout(n17516));
  jand g17362(.dina(n17516), .dinb(n17515), .dout(n17517));
  jxor g17363(.dina(n17142), .dinb(n17141), .dout(n17518));
  jnot g17364(.din(n17518), .dout(n17519));
  jor  g17365(.dina(n14221), .dinb(n7891), .dout(n17520));
  jor  g17366(.dina(n15045), .dinb(n8440), .dout(n17521));
  jor  g17367(.dina(n11984), .dinb(n8155), .dout(n17522));
  jor  g17368(.dina(n11987), .dinb(n7889), .dout(n17523));
  jand g17369(.dina(n17523), .dinb(n17522), .dout(n17524));
  jand g17370(.dina(n17524), .dinb(n17521), .dout(n17525));
  jand g17371(.dina(n17525), .dinb(n17520), .dout(n17526));
  jxor g17372(.dina(n17526), .dinb(\a[11] ), .dout(n17527));
  jor  g17373(.dina(n17527), .dinb(n17519), .dout(n17528));
  jxor g17374(.dina(n17139), .dinb(n17138), .dout(n17529));
  jnot g17375(.din(n17529), .dout(n17530));
  jor  g17376(.dina(n14248), .dinb(n7891), .dout(n17531));
  jor  g17377(.dina(n11984), .dinb(n8440), .dout(n17532));
  jor  g17378(.dina(n11987), .dinb(n8155), .dout(n17533));
  jor  g17379(.dina(n11991), .dinb(n7889), .dout(n17534));
  jand g17380(.dina(n17534), .dinb(n17533), .dout(n17535));
  jand g17381(.dina(n17535), .dinb(n17532), .dout(n17536));
  jand g17382(.dina(n17536), .dinb(n17531), .dout(n17537));
  jxor g17383(.dina(n17537), .dinb(\a[11] ), .dout(n17538));
  jor  g17384(.dina(n17538), .dinb(n17530), .dout(n17539));
  jxor g17385(.dina(n17136), .dinb(n17135), .dout(n17540));
  jnot g17386(.din(n17540), .dout(n17541));
  jor  g17387(.dina(n14271), .dinb(n7891), .dout(n17542));
  jor  g17388(.dina(n11987), .dinb(n8440), .dout(n17543));
  jor  g17389(.dina(n11991), .dinb(n8155), .dout(n17544));
  jor  g17390(.dina(n11995), .dinb(n7889), .dout(n17545));
  jand g17391(.dina(n17545), .dinb(n17544), .dout(n17546));
  jand g17392(.dina(n17546), .dinb(n17543), .dout(n17547));
  jand g17393(.dina(n17547), .dinb(n17542), .dout(n17548));
  jxor g17394(.dina(n17548), .dinb(\a[11] ), .dout(n17549));
  jor  g17395(.dina(n17549), .dinb(n17541), .dout(n17550));
  jor  g17396(.dina(n14301), .dinb(n7891), .dout(n17551));
  jor  g17397(.dina(n11991), .dinb(n8440), .dout(n17552));
  jor  g17398(.dina(n11995), .dinb(n8155), .dout(n17553));
  jor  g17399(.dina(n11997), .dinb(n7889), .dout(n17554));
  jand g17400(.dina(n17554), .dinb(n17553), .dout(n17555));
  jand g17401(.dina(n17555), .dinb(n17552), .dout(n17556));
  jand g17402(.dina(n17556), .dinb(n17551), .dout(n17557));
  jxor g17403(.dina(n17557), .dinb(\a[11] ), .dout(n17558));
  jnot g17404(.din(n17558), .dout(n17559));
  jxor g17405(.dina(n17133), .dinb(n17132), .dout(n17560));
  jand g17406(.dina(n17560), .dinb(n17559), .dout(n17561));
  jor  g17407(.dina(n14353), .dinb(n7891), .dout(n17562));
  jor  g17408(.dina(n11995), .dinb(n8440), .dout(n17563));
  jor  g17409(.dina(n11997), .dinb(n8155), .dout(n17564));
  jor  g17410(.dina(n11999), .dinb(n7889), .dout(n17565));
  jand g17411(.dina(n17565), .dinb(n17564), .dout(n17566));
  jand g17412(.dina(n17566), .dinb(n17563), .dout(n17567));
  jand g17413(.dina(n17567), .dinb(n17562), .dout(n17568));
  jxor g17414(.dina(n17568), .dinb(\a[11] ), .dout(n17569));
  jnot g17415(.din(n17569), .dout(n17570));
  jxor g17416(.dina(n17130), .dinb(n17129), .dout(n17571));
  jand g17417(.dina(n17571), .dinb(n17570), .dout(n17572));
  jor  g17418(.dina(n14390), .dinb(n7891), .dout(n17573));
  jor  g17419(.dina(n11997), .dinb(n8440), .dout(n17574));
  jor  g17420(.dina(n11999), .dinb(n8155), .dout(n17575));
  jor  g17421(.dina(n12001), .dinb(n7889), .dout(n17576));
  jand g17422(.dina(n17576), .dinb(n17575), .dout(n17577));
  jand g17423(.dina(n17577), .dinb(n17574), .dout(n17578));
  jand g17424(.dina(n17578), .dinb(n17573), .dout(n17579));
  jxor g17425(.dina(n17579), .dinb(\a[11] ), .dout(n17580));
  jnot g17426(.din(n17580), .dout(n17581));
  jor  g17427(.dina(n17110), .dinb(n5292), .dout(n17582));
  jxor g17428(.dina(n17582), .dinb(n17118), .dout(n17583));
  jand g17429(.dina(n17583), .dinb(n17581), .dout(n17584));
  jor  g17430(.dina(n14432), .dinb(n7891), .dout(n17585));
  jor  g17431(.dina(n11999), .dinb(n8440), .dout(n17586));
  jor  g17432(.dina(n12001), .dinb(n8155), .dout(n17587));
  jor  g17433(.dina(n12004), .dinb(n7889), .dout(n17588));
  jand g17434(.dina(n17588), .dinb(n17587), .dout(n17589));
  jand g17435(.dina(n17589), .dinb(n17586), .dout(n17590));
  jand g17436(.dina(n17590), .dinb(n17585), .dout(n17591));
  jxor g17437(.dina(n17591), .dinb(\a[11] ), .dout(n17592));
  jnot g17438(.din(n17592), .dout(n17593));
  jand g17439(.dina(n17107), .dinb(\a[14] ), .dout(n17594));
  jxor g17440(.dina(n17594), .dinb(n17105), .dout(n17595));
  jand g17441(.dina(n17595), .dinb(n17593), .dout(n17596));
  jand g17442(.dina(n14497), .dinb(n7890), .dout(n17597));
  jand g17443(.dina(n12010), .dinb(n8154), .dout(n17598));
  jand g17444(.dina(n12008), .dinb(n8441), .dout(n17599));
  jor  g17445(.dina(n17599), .dinb(n17598), .dout(n17600));
  jor  g17446(.dina(n17600), .dinb(n17597), .dout(n17601));
  jnot g17447(.din(n17601), .dout(n17602));
  jand g17448(.dina(n12010), .dinb(n7884), .dout(n17603));
  jnot g17449(.din(n17603), .dout(n17604));
  jand g17450(.dina(n17604), .dinb(\a[11] ), .dout(n17605));
  jand g17451(.dina(n17605), .dinb(n17602), .dout(n17606));
  jand g17452(.dina(n14537), .dinb(n7890), .dout(n17607));
  jand g17453(.dina(n12006), .dinb(n8441), .dout(n17608));
  jand g17454(.dina(n12008), .dinb(n8154), .dout(n17609));
  jand g17455(.dina(n12010), .dinb(n7888), .dout(n17610));
  jor  g17456(.dina(n17610), .dinb(n17609), .dout(n17611));
  jor  g17457(.dina(n17611), .dinb(n17608), .dout(n17612));
  jor  g17458(.dina(n17612), .dinb(n17607), .dout(n17613));
  jnot g17459(.din(n17613), .dout(n17614));
  jand g17460(.dina(n17614), .dinb(n17606), .dout(n17615));
  jand g17461(.dina(n17615), .dinb(n17107), .dout(n17616));
  jor  g17462(.dina(n15144), .dinb(n7891), .dout(n17617));
  jor  g17463(.dina(n12001), .dinb(n8440), .dout(n17618));
  jor  g17464(.dina(n12004), .dinb(n8155), .dout(n17619));
  jor  g17465(.dina(n12009), .dinb(n7889), .dout(n17620));
  jand g17466(.dina(n17620), .dinb(n17619), .dout(n17621));
  jand g17467(.dina(n17621), .dinb(n17618), .dout(n17622));
  jand g17468(.dina(n17622), .dinb(n17617), .dout(n17623));
  jxor g17469(.dina(n17623), .dinb(\a[11] ), .dout(n17624));
  jnot g17470(.din(n17624), .dout(n17625));
  jxor g17471(.dina(n17615), .dinb(n17107), .dout(n17626));
  jand g17472(.dina(n17626), .dinb(n17625), .dout(n17627));
  jor  g17473(.dina(n17627), .dinb(n17616), .dout(n17628));
  jxor g17474(.dina(n17595), .dinb(n17593), .dout(n17629));
  jand g17475(.dina(n17629), .dinb(n17628), .dout(n17630));
  jor  g17476(.dina(n17630), .dinb(n17596), .dout(n17631));
  jxor g17477(.dina(n17583), .dinb(n17581), .dout(n17632));
  jand g17478(.dina(n17632), .dinb(n17631), .dout(n17633));
  jor  g17479(.dina(n17633), .dinb(n17584), .dout(n17634));
  jxor g17480(.dina(n17571), .dinb(n17570), .dout(n17635));
  jand g17481(.dina(n17635), .dinb(n17634), .dout(n17636));
  jor  g17482(.dina(n17636), .dinb(n17572), .dout(n17637));
  jxor g17483(.dina(n17560), .dinb(n17559), .dout(n17638));
  jand g17484(.dina(n17638), .dinb(n17637), .dout(n17639));
  jor  g17485(.dina(n17639), .dinb(n17561), .dout(n17640));
  jxor g17486(.dina(n17549), .dinb(n17541), .dout(n17641));
  jand g17487(.dina(n17641), .dinb(n17640), .dout(n17642));
  jnot g17488(.din(n17642), .dout(n17643));
  jand g17489(.dina(n17643), .dinb(n17550), .dout(n17644));
  jnot g17490(.din(n17644), .dout(n17645));
  jxor g17491(.dina(n17538), .dinb(n17530), .dout(n17646));
  jand g17492(.dina(n17646), .dinb(n17645), .dout(n17647));
  jnot g17493(.din(n17647), .dout(n17648));
  jand g17494(.dina(n17648), .dinb(n17539), .dout(n17649));
  jnot g17495(.din(n17649), .dout(n17650));
  jxor g17496(.dina(n17527), .dinb(n17519), .dout(n17651));
  jand g17497(.dina(n17651), .dinb(n17650), .dout(n17652));
  jnot g17498(.din(n17652), .dout(n17653));
  jand g17499(.dina(n17653), .dinb(n17528), .dout(n17654));
  jnot g17500(.din(n17654), .dout(n17655));
  jxor g17501(.dina(n17516), .dinb(n17515), .dout(n17656));
  jand g17502(.dina(n17656), .dinb(n17655), .dout(n17657));
  jor  g17503(.dina(n17657), .dinb(n17517), .dout(n17658));
  jxor g17504(.dina(n17505), .dinb(n17504), .dout(n17659));
  jand g17505(.dina(n17659), .dinb(n17658), .dout(n17660));
  jor  g17506(.dina(n17660), .dinb(n17506), .dout(n17661));
  jxor g17507(.dina(n17494), .dinb(n17493), .dout(n17662));
  jand g17508(.dina(n17662), .dinb(n17661), .dout(n17663));
  jor  g17509(.dina(n17663), .dinb(n17495), .dout(n17664));
  jxor g17510(.dina(n17483), .dinb(n17475), .dout(n17665));
  jand g17511(.dina(n17665), .dinb(n17664), .dout(n17666));
  jnot g17512(.din(n17666), .dout(n17667));
  jand g17513(.dina(n17667), .dinb(n17484), .dout(n17668));
  jnot g17514(.din(n17668), .dout(n17669));
  jxor g17515(.dina(n17472), .dinb(n17464), .dout(n17670));
  jand g17516(.dina(n17670), .dinb(n17669), .dout(n17671));
  jnot g17517(.din(n17671), .dout(n17672));
  jand g17518(.dina(n17672), .dinb(n17473), .dout(n17673));
  jnot g17519(.din(n17673), .dout(n17674));
  jxor g17520(.dina(n17461), .dinb(n17453), .dout(n17675));
  jand g17521(.dina(n17675), .dinb(n17674), .dout(n17676));
  jnot g17522(.din(n17676), .dout(n17677));
  jand g17523(.dina(n17677), .dinb(n17462), .dout(n17678));
  jnot g17524(.din(n17678), .dout(n17679));
  jxor g17525(.dina(n17450), .dinb(n17449), .dout(n17680));
  jand g17526(.dina(n17680), .dinb(n17679), .dout(n17681));
  jor  g17527(.dina(n17681), .dinb(n17451), .dout(n17682));
  jxor g17528(.dina(n17439), .dinb(n17438), .dout(n17683));
  jand g17529(.dina(n17683), .dinb(n17682), .dout(n17684));
  jor  g17530(.dina(n17684), .dinb(n17440), .dout(n17685));
  jxor g17531(.dina(n17428), .dinb(n17427), .dout(n17686));
  jand g17532(.dina(n17686), .dinb(n17685), .dout(n17687));
  jor  g17533(.dina(n17687), .dinb(n17429), .dout(n17688));
  jxor g17534(.dina(n17417), .dinb(n17409), .dout(n17689));
  jand g17535(.dina(n17689), .dinb(n17688), .dout(n17690));
  jnot g17536(.din(n17690), .dout(n17691));
  jand g17537(.dina(n17691), .dinb(n17418), .dout(n17692));
  jnot g17538(.din(n17692), .dout(n17693));
  jxor g17539(.dina(n17406), .dinb(n17398), .dout(n17694));
  jand g17540(.dina(n17694), .dinb(n17693), .dout(n17695));
  jnot g17541(.din(n17695), .dout(n17696));
  jand g17542(.dina(n17696), .dinb(n17407), .dout(n17697));
  jnot g17543(.din(n17697), .dout(n17698));
  jxor g17544(.dina(n17395), .dinb(n17394), .dout(n17699));
  jand g17545(.dina(n17699), .dinb(n17698), .dout(n17700));
  jor  g17546(.dina(n17700), .dinb(n17396), .dout(n17701));
  jxor g17547(.dina(n17384), .dinb(n17383), .dout(n17702));
  jand g17548(.dina(n17702), .dinb(n17701), .dout(n17703));
  jor  g17549(.dina(n17703), .dinb(n17385), .dout(n17704));
  jxor g17550(.dina(n17373), .dinb(n17372), .dout(n17705));
  jand g17551(.dina(n17705), .dinb(n17704), .dout(n17706));
  jor  g17552(.dina(n17706), .dinb(n17374), .dout(n17707));
  jxor g17553(.dina(n17362), .dinb(n17361), .dout(n17708));
  jand g17554(.dina(n17708), .dinb(n17707), .dout(n17709));
  jor  g17555(.dina(n17709), .dinb(n17363), .dout(n17710));
  jxor g17556(.dina(n17351), .dinb(n17350), .dout(n17711));
  jand g17557(.dina(n17711), .dinb(n17710), .dout(n17712));
  jor  g17558(.dina(n17712), .dinb(n17352), .dout(n17713));
  jxor g17559(.dina(n17340), .dinb(n17339), .dout(n17714));
  jand g17560(.dina(n17714), .dinb(n17713), .dout(n17715));
  jor  g17561(.dina(n17715), .dinb(n17341), .dout(n17716));
  jxor g17562(.dina(n17329), .dinb(n17328), .dout(n17717));
  jand g17563(.dina(n17717), .dinb(n17716), .dout(n17718));
  jor  g17564(.dina(n17718), .dinb(n17330), .dout(n17719));
  jxor g17565(.dina(n17318), .dinb(n17317), .dout(n17720));
  jand g17566(.dina(n17720), .dinb(n17719), .dout(n17721));
  jor  g17567(.dina(n17721), .dinb(n17319), .dout(n17722));
  jxor g17568(.dina(n17307), .dinb(n17306), .dout(n17723));
  jand g17569(.dina(n17723), .dinb(n17722), .dout(n17724));
  jor  g17570(.dina(n17724), .dinb(n17308), .dout(n17725));
  jxor g17571(.dina(n17296), .dinb(n17295), .dout(n17726));
  jand g17572(.dina(n17726), .dinb(n17725), .dout(n17727));
  jor  g17573(.dina(n17727), .dinb(n17297), .dout(n17728));
  jxor g17574(.dina(n17252), .dinb(n17244), .dout(n17729));
  jand g17575(.dina(n17729), .dinb(n17728), .dout(n17730));
  jnot g17576(.din(n17730), .dout(n17731));
  jxor g17577(.dina(n17729), .dinb(n17728), .dout(n17732));
  jnot g17578(.din(n17732), .dout(n17733));
  jand g17579(.dina(n12938), .dinb(n8771), .dout(n17734));
  jand g17580(.dina(n12782), .dinb(n9491), .dout(n17735));
  jand g17581(.dina(n12783), .dinb(n9126), .dout(n17736));
  jand g17582(.dina(n12766), .dinb(n8769), .dout(n17737));
  jor  g17583(.dina(n17737), .dinb(n17736), .dout(n17738));
  jor  g17584(.dina(n17738), .dinb(n17735), .dout(n17739));
  jor  g17585(.dina(n17739), .dinb(n17734), .dout(n17740));
  jxor g17586(.dina(n17740), .dinb(n6039), .dout(n17741));
  jor  g17587(.dina(n17741), .dinb(n17733), .dout(n17742));
  jand g17588(.dina(n17742), .dinb(n17731), .dout(n17743));
  jnot g17589(.din(n17743), .dout(n17744));
  jxor g17590(.dina(n17268), .dinb(n17260), .dout(n17745));
  jand g17591(.dina(n17745), .dinb(n17744), .dout(n17746));
  jnot g17592(.din(n17746), .dout(n17747));
  jxor g17593(.dina(n17745), .dinb(n17744), .dout(n17748));
  jnot g17594(.din(n17748), .dout(n17749));
  jor  g17595(.dina(n12814), .dinb(n9918), .dout(n17751));
  jand g17596(.dina(n17273), .dinb(n17751), .dout(n17755));
  jand g17597(.dina(n17755), .dinb(n9919), .dout(n17756));
  jxor g17598(.dina(n17756), .dinb(\a[5] ), .dout(n17757));
  jor  g17599(.dina(n17757), .dinb(n17749), .dout(n17758));
  jand g17600(.dina(n17758), .dinb(n17747), .dout(n17759));
  jnot g17601(.din(n17759), .dout(n17760));
  jxor g17602(.dina(n17280), .dinb(n17279), .dout(n17761));
  jand g17603(.dina(n17761), .dinb(n17760), .dout(n17762));
  jnot g17604(.din(n17762), .dout(n17763));
  jxor g17605(.dina(n17761), .dinb(n17760), .dout(n17764));
  jnot g17606(.din(n17764), .dout(n17765));
  jxor g17607(.dina(n17726), .dinb(n17725), .dout(n17766));
  jnot g17608(.din(n17766), .dout(n17767));
  jand g17609(.dina(n12841), .dinb(n8771), .dout(n17768));
  jand g17610(.dina(n12783), .dinb(n9491), .dout(n17769));
  jand g17611(.dina(n12766), .dinb(n9126), .dout(n17770));
  jand g17612(.dina(n12177), .dinb(n8769), .dout(n17771));
  jor  g17613(.dina(n17771), .dinb(n17770), .dout(n17772));
  jor  g17614(.dina(n17772), .dinb(n17769), .dout(n17773));
  jor  g17615(.dina(n17773), .dinb(n17768), .dout(n17774));
  jxor g17616(.dina(n17774), .dinb(n6039), .dout(n17775));
  jor  g17617(.dina(n17775), .dinb(n17767), .dout(n17776));
  jxor g17618(.dina(n17723), .dinb(n17722), .dout(n17777));
  jnot g17619(.din(n17777), .dout(n17778));
  jand g17620(.dina(n12768), .dinb(n8771), .dout(n17779));
  jand g17621(.dina(n12766), .dinb(n9491), .dout(n17780));
  jand g17622(.dina(n12177), .dinb(n9126), .dout(n17781));
  jand g17623(.dina(n11941), .dinb(n8769), .dout(n17782));
  jor  g17624(.dina(n17782), .dinb(n17781), .dout(n17783));
  jor  g17625(.dina(n17783), .dinb(n17780), .dout(n17784));
  jor  g17626(.dina(n17784), .dinb(n17779), .dout(n17785));
  jxor g17627(.dina(n17785), .dinb(n6039), .dout(n17786));
  jor  g17628(.dina(n17786), .dinb(n17778), .dout(n17787));
  jxor g17629(.dina(n17720), .dinb(n17719), .dout(n17788));
  jnot g17630(.din(n17788), .dout(n17789));
  jand g17631(.dina(n12179), .dinb(n8771), .dout(n17790));
  jand g17632(.dina(n12177), .dinb(n9491), .dout(n17791));
  jand g17633(.dina(n11941), .dinb(n9126), .dout(n17792));
  jand g17634(.dina(n11942), .dinb(n8769), .dout(n17793));
  jor  g17635(.dina(n17793), .dinb(n17792), .dout(n17794));
  jor  g17636(.dina(n17794), .dinb(n17791), .dout(n17795));
  jor  g17637(.dina(n17795), .dinb(n17790), .dout(n17796));
  jxor g17638(.dina(n17796), .dinb(n6039), .dout(n17797));
  jor  g17639(.dina(n17797), .dinb(n17789), .dout(n17798));
  jnot g17640(.din(n17798), .dout(n17799));
  jxor g17641(.dina(n17717), .dinb(n17716), .dout(n17800));
  jnot g17642(.din(n17800), .dout(n17801));
  jand g17643(.dina(n12671), .dinb(n8771), .dout(n17802));
  jand g17644(.dina(n11941), .dinb(n9491), .dout(n17803));
  jand g17645(.dina(n11942), .dinb(n9126), .dout(n17804));
  jand g17646(.dina(n11944), .dinb(n8769), .dout(n17805));
  jor  g17647(.dina(n17805), .dinb(n17804), .dout(n17806));
  jor  g17648(.dina(n17806), .dinb(n17803), .dout(n17807));
  jor  g17649(.dina(n17807), .dinb(n17802), .dout(n17808));
  jxor g17650(.dina(n17808), .dinb(n6039), .dout(n17809));
  jor  g17651(.dina(n17809), .dinb(n17801), .dout(n17810));
  jxor g17652(.dina(n17714), .dinb(n17713), .dout(n17811));
  jnot g17653(.din(n17811), .dout(n17812));
  jand g17654(.dina(n12751), .dinb(n8771), .dout(n17813));
  jand g17655(.dina(n11942), .dinb(n9491), .dout(n17814));
  jand g17656(.dina(n11944), .dinb(n9126), .dout(n17815));
  jand g17657(.dina(n11946), .dinb(n8769), .dout(n17816));
  jor  g17658(.dina(n17816), .dinb(n17815), .dout(n17817));
  jor  g17659(.dina(n17817), .dinb(n17814), .dout(n17818));
  jor  g17660(.dina(n17818), .dinb(n17813), .dout(n17819));
  jxor g17661(.dina(n17819), .dinb(n6039), .dout(n17820));
  jor  g17662(.dina(n17820), .dinb(n17812), .dout(n17821));
  jxor g17663(.dina(n17711), .dinb(n17710), .dout(n17822));
  jnot g17664(.din(n17822), .dout(n17823));
  jand g17665(.dina(n12189), .dinb(n8771), .dout(n17824));
  jand g17666(.dina(n11944), .dinb(n9491), .dout(n17825));
  jand g17667(.dina(n11946), .dinb(n9126), .dout(n17826));
  jand g17668(.dina(n11948), .dinb(n8769), .dout(n17827));
  jor  g17669(.dina(n17827), .dinb(n17826), .dout(n17828));
  jor  g17670(.dina(n17828), .dinb(n17825), .dout(n17829));
  jor  g17671(.dina(n17829), .dinb(n17824), .dout(n17830));
  jxor g17672(.dina(n17830), .dinb(n6039), .dout(n17831));
  jor  g17673(.dina(n17831), .dinb(n17823), .dout(n17832));
  jxor g17674(.dina(n17708), .dinb(n17707), .dout(n17833));
  jnot g17675(.din(n17833), .dout(n17834));
  jand g17676(.dina(n12519), .dinb(n8771), .dout(n17835));
  jand g17677(.dina(n11946), .dinb(n9491), .dout(n17836));
  jand g17678(.dina(n11948), .dinb(n9126), .dout(n17837));
  jand g17679(.dina(n11950), .dinb(n8769), .dout(n17838));
  jor  g17680(.dina(n17838), .dinb(n17837), .dout(n17839));
  jor  g17681(.dina(n17839), .dinb(n17836), .dout(n17840));
  jor  g17682(.dina(n17840), .dinb(n17835), .dout(n17841));
  jxor g17683(.dina(n17841), .dinb(n6039), .dout(n17842));
  jor  g17684(.dina(n17842), .dinb(n17834), .dout(n17843));
  jxor g17685(.dina(n17705), .dinb(n17704), .dout(n17844));
  jnot g17686(.din(n17844), .dout(n17845));
  jand g17687(.dina(n12654), .dinb(n8771), .dout(n17846));
  jand g17688(.dina(n11948), .dinb(n9491), .dout(n17847));
  jand g17689(.dina(n11950), .dinb(n9126), .dout(n17848));
  jand g17690(.dina(n11952), .dinb(n8769), .dout(n17849));
  jor  g17691(.dina(n17849), .dinb(n17848), .dout(n17850));
  jor  g17692(.dina(n17850), .dinb(n17847), .dout(n17851));
  jor  g17693(.dina(n17851), .dinb(n17846), .dout(n17852));
  jxor g17694(.dina(n17852), .dinb(n6039), .dout(n17853));
  jor  g17695(.dina(n17853), .dinb(n17845), .dout(n17854));
  jxor g17696(.dina(n17702), .dinb(n17701), .dout(n17855));
  jnot g17697(.din(n17855), .dout(n17856));
  jand g17698(.dina(n12569), .dinb(n8771), .dout(n17857));
  jand g17699(.dina(n11950), .dinb(n9491), .dout(n17858));
  jand g17700(.dina(n11952), .dinb(n9126), .dout(n17859));
  jand g17701(.dina(n11954), .dinb(n8769), .dout(n17860));
  jor  g17702(.dina(n17860), .dinb(n17859), .dout(n17861));
  jor  g17703(.dina(n17861), .dinb(n17858), .dout(n17862));
  jor  g17704(.dina(n17862), .dinb(n17857), .dout(n17863));
  jxor g17705(.dina(n17863), .dinb(n6039), .dout(n17864));
  jor  g17706(.dina(n17864), .dinb(n17856), .dout(n17865));
  jxor g17707(.dina(n17699), .dinb(n17698), .dout(n17866));
  jnot g17708(.din(n17866), .dout(n17867));
  jand g17709(.dina(n12510), .dinb(n8771), .dout(n17868));
  jand g17710(.dina(n11952), .dinb(n9491), .dout(n17869));
  jand g17711(.dina(n11954), .dinb(n9126), .dout(n17870));
  jand g17712(.dina(n11956), .dinb(n8769), .dout(n17871));
  jor  g17713(.dina(n17871), .dinb(n17870), .dout(n17872));
  jor  g17714(.dina(n17872), .dinb(n17869), .dout(n17873));
  jor  g17715(.dina(n17873), .dinb(n17868), .dout(n17874));
  jxor g17716(.dina(n17874), .dinb(n6039), .dout(n17875));
  jor  g17717(.dina(n17875), .dinb(n17867), .dout(n17876));
  jand g17718(.dina(n12472), .dinb(n8771), .dout(n17877));
  jand g17719(.dina(n11954), .dinb(n9491), .dout(n17878));
  jand g17720(.dina(n11956), .dinb(n9126), .dout(n17879));
  jand g17721(.dina(n11958), .dinb(n8769), .dout(n17880));
  jor  g17722(.dina(n17880), .dinb(n17879), .dout(n17881));
  jor  g17723(.dina(n17881), .dinb(n17878), .dout(n17882));
  jor  g17724(.dina(n17882), .dinb(n17877), .dout(n17883));
  jxor g17725(.dina(n17883), .dinb(n6039), .dout(n17884));
  jnot g17726(.din(n17884), .dout(n17885));
  jxor g17727(.dina(n17694), .dinb(n17693), .dout(n17886));
  jand g17728(.dina(n17886), .dinb(n17885), .dout(n17887));
  jand g17729(.dina(n12639), .dinb(n8771), .dout(n17888));
  jand g17730(.dina(n11956), .dinb(n9491), .dout(n17889));
  jand g17731(.dina(n11958), .dinb(n9126), .dout(n17890));
  jand g17732(.dina(n11960), .dinb(n8769), .dout(n17891));
  jor  g17733(.dina(n17891), .dinb(n17890), .dout(n17892));
  jor  g17734(.dina(n17892), .dinb(n17889), .dout(n17893));
  jor  g17735(.dina(n17893), .dinb(n17888), .dout(n17894));
  jxor g17736(.dina(n17894), .dinb(n6039), .dout(n17895));
  jnot g17737(.din(n17895), .dout(n17896));
  jxor g17738(.dina(n17689), .dinb(n17688), .dout(n17897));
  jand g17739(.dina(n17897), .dinb(n17896), .dout(n17898));
  jxor g17740(.dina(n17686), .dinb(n17685), .dout(n17899));
  jnot g17741(.din(n17899), .dout(n17900));
  jand g17742(.dina(n12624), .dinb(n8771), .dout(n17901));
  jand g17743(.dina(n11958), .dinb(n9491), .dout(n17902));
  jand g17744(.dina(n11960), .dinb(n9126), .dout(n17903));
  jand g17745(.dina(n11962), .dinb(n8769), .dout(n17904));
  jor  g17746(.dina(n17904), .dinb(n17903), .dout(n17905));
  jor  g17747(.dina(n17905), .dinb(n17902), .dout(n17906));
  jor  g17748(.dina(n17906), .dinb(n17901), .dout(n17907));
  jxor g17749(.dina(n17907), .dinb(n6039), .dout(n17908));
  jor  g17750(.dina(n17908), .dinb(n17900), .dout(n17909));
  jxor g17751(.dina(n17683), .dinb(n17682), .dout(n17910));
  jnot g17752(.din(n17910), .dout(n17911));
  jand g17753(.dina(n13116), .dinb(n8771), .dout(n17912));
  jand g17754(.dina(n11960), .dinb(n9491), .dout(n17913));
  jand g17755(.dina(n11962), .dinb(n9126), .dout(n17914));
  jand g17756(.dina(n11964), .dinb(n8769), .dout(n17915));
  jor  g17757(.dina(n17915), .dinb(n17914), .dout(n17916));
  jor  g17758(.dina(n17916), .dinb(n17913), .dout(n17917));
  jor  g17759(.dina(n17917), .dinb(n17912), .dout(n17918));
  jxor g17760(.dina(n17918), .dinb(n6039), .dout(n17919));
  jor  g17761(.dina(n17919), .dinb(n17911), .dout(n17920));
  jxor g17762(.dina(n17680), .dinb(n17679), .dout(n17921));
  jnot g17763(.din(n17921), .dout(n17922));
  jand g17764(.dina(n13134), .dinb(n8771), .dout(n17923));
  jand g17765(.dina(n11962), .dinb(n9491), .dout(n17924));
  jand g17766(.dina(n11964), .dinb(n9126), .dout(n17925));
  jand g17767(.dina(n11966), .dinb(n8769), .dout(n17926));
  jor  g17768(.dina(n17926), .dinb(n17925), .dout(n17927));
  jor  g17769(.dina(n17927), .dinb(n17924), .dout(n17928));
  jor  g17770(.dina(n17928), .dinb(n17923), .dout(n17929));
  jxor g17771(.dina(n17929), .dinb(n6039), .dout(n17930));
  jor  g17772(.dina(n17930), .dinb(n17922), .dout(n17931));
  jand g17773(.dina(n13470), .dinb(n8771), .dout(n17932));
  jand g17774(.dina(n11964), .dinb(n9491), .dout(n17933));
  jand g17775(.dina(n11966), .dinb(n9126), .dout(n17934));
  jand g17776(.dina(n11968), .dinb(n8769), .dout(n17935));
  jor  g17777(.dina(n17935), .dinb(n17934), .dout(n17936));
  jor  g17778(.dina(n17936), .dinb(n17933), .dout(n17937));
  jor  g17779(.dina(n17937), .dinb(n17932), .dout(n17938));
  jxor g17780(.dina(n17938), .dinb(n6039), .dout(n17939));
  jnot g17781(.din(n17939), .dout(n17940));
  jxor g17782(.dina(n17675), .dinb(n17674), .dout(n17941));
  jand g17783(.dina(n17941), .dinb(n17940), .dout(n17942));
  jand g17784(.dina(n13268), .dinb(n8771), .dout(n17943));
  jand g17785(.dina(n11966), .dinb(n9491), .dout(n17944));
  jand g17786(.dina(n11968), .dinb(n9126), .dout(n17945));
  jand g17787(.dina(n11970), .dinb(n8769), .dout(n17946));
  jor  g17788(.dina(n17946), .dinb(n17945), .dout(n17947));
  jor  g17789(.dina(n17947), .dinb(n17944), .dout(n17948));
  jor  g17790(.dina(n17948), .dinb(n17943), .dout(n17949));
  jxor g17791(.dina(n17949), .dinb(n6039), .dout(n17950));
  jnot g17792(.din(n17950), .dout(n17951));
  jxor g17793(.dina(n17670), .dinb(n17669), .dout(n17952));
  jand g17794(.dina(n17952), .dinb(n17951), .dout(n17953));
  jand g17795(.dina(n13682), .dinb(n8771), .dout(n17954));
  jand g17796(.dina(n11968), .dinb(n9491), .dout(n17955));
  jand g17797(.dina(n11970), .dinb(n9126), .dout(n17956));
  jand g17798(.dina(n11972), .dinb(n8769), .dout(n17957));
  jor  g17799(.dina(n17957), .dinb(n17956), .dout(n17958));
  jor  g17800(.dina(n17958), .dinb(n17955), .dout(n17959));
  jor  g17801(.dina(n17959), .dinb(n17954), .dout(n17960));
  jxor g17802(.dina(n17960), .dinb(n6039), .dout(n17961));
  jnot g17803(.din(n17961), .dout(n17962));
  jxor g17804(.dina(n17665), .dinb(n17664), .dout(n17963));
  jand g17805(.dina(n17963), .dinb(n17962), .dout(n17964));
  jxor g17806(.dina(n17662), .dinb(n17661), .dout(n17965));
  jnot g17807(.din(n17965), .dout(n17966));
  jand g17808(.dina(n13806), .dinb(n8771), .dout(n17967));
  jand g17809(.dina(n11970), .dinb(n9491), .dout(n17968));
  jand g17810(.dina(n11972), .dinb(n9126), .dout(n17969));
  jand g17811(.dina(n11974), .dinb(n8769), .dout(n17970));
  jor  g17812(.dina(n17970), .dinb(n17969), .dout(n17971));
  jor  g17813(.dina(n17971), .dinb(n17968), .dout(n17972));
  jor  g17814(.dina(n17972), .dinb(n17967), .dout(n17973));
  jxor g17815(.dina(n17973), .dinb(n6039), .dout(n17974));
  jor  g17816(.dina(n17974), .dinb(n17966), .dout(n17975));
  jxor g17817(.dina(n17659), .dinb(n17658), .dout(n17976));
  jnot g17818(.din(n17976), .dout(n17977));
  jand g17819(.dina(n13664), .dinb(n8771), .dout(n17978));
  jand g17820(.dina(n11972), .dinb(n9491), .dout(n17979));
  jand g17821(.dina(n11974), .dinb(n9126), .dout(n17980));
  jand g17822(.dina(n11976), .dinb(n8769), .dout(n17981));
  jor  g17823(.dina(n17981), .dinb(n17980), .dout(n17982));
  jor  g17824(.dina(n17982), .dinb(n17979), .dout(n17983));
  jor  g17825(.dina(n17983), .dinb(n17978), .dout(n17984));
  jxor g17826(.dina(n17984), .dinb(n6039), .dout(n17985));
  jor  g17827(.dina(n17985), .dinb(n17977), .dout(n17986));
  jxor g17828(.dina(n17656), .dinb(n17655), .dout(n17987));
  jnot g17829(.din(n17987), .dout(n17988));
  jand g17830(.dina(n13924), .dinb(n8771), .dout(n17989));
  jand g17831(.dina(n11974), .dinb(n9491), .dout(n17990));
  jand g17832(.dina(n11976), .dinb(n9126), .dout(n17991));
  jand g17833(.dina(n11978), .dinb(n8769), .dout(n17992));
  jor  g17834(.dina(n17992), .dinb(n17991), .dout(n17993));
  jor  g17835(.dina(n17993), .dinb(n17990), .dout(n17994));
  jor  g17836(.dina(n17994), .dinb(n17989), .dout(n17995));
  jxor g17837(.dina(n17995), .dinb(n6039), .dout(n17996));
  jor  g17838(.dina(n17996), .dinb(n17988), .dout(n17997));
  jand g17839(.dina(n14184), .dinb(n8771), .dout(n17998));
  jand g17840(.dina(n11976), .dinb(n9491), .dout(n17999));
  jand g17841(.dina(n11978), .dinb(n9126), .dout(n18000));
  jand g17842(.dina(n11980), .dinb(n8769), .dout(n18001));
  jor  g17843(.dina(n18001), .dinb(n18000), .dout(n18002));
  jor  g17844(.dina(n18002), .dinb(n17999), .dout(n18003));
  jor  g17845(.dina(n18003), .dinb(n17998), .dout(n18004));
  jxor g17846(.dina(n18004), .dinb(n6039), .dout(n18005));
  jnot g17847(.din(n18005), .dout(n18006));
  jxor g17848(.dina(n17651), .dinb(n17650), .dout(n18007));
  jand g17849(.dina(n18007), .dinb(n18006), .dout(n18008));
  jand g17850(.dina(n14194), .dinb(n8771), .dout(n18009));
  jand g17851(.dina(n11978), .dinb(n9491), .dout(n18010));
  jand g17852(.dina(n11980), .dinb(n9126), .dout(n18011));
  jand g17853(.dina(n11982), .dinb(n8769), .dout(n18012));
  jor  g17854(.dina(n18012), .dinb(n18011), .dout(n18013));
  jor  g17855(.dina(n18013), .dinb(n18010), .dout(n18014));
  jor  g17856(.dina(n18014), .dinb(n18009), .dout(n18015));
  jxor g17857(.dina(n18015), .dinb(n6039), .dout(n18016));
  jnot g17858(.din(n18016), .dout(n18017));
  jxor g17859(.dina(n17646), .dinb(n17645), .dout(n18018));
  jand g17860(.dina(n18018), .dinb(n18017), .dout(n18019));
  jand g17861(.dina(n13899), .dinb(n8771), .dout(n18020));
  jand g17862(.dina(n11980), .dinb(n9491), .dout(n18021));
  jand g17863(.dina(n11982), .dinb(n9126), .dout(n18022));
  jand g17864(.dina(n11985), .dinb(n8769), .dout(n18023));
  jor  g17865(.dina(n18023), .dinb(n18022), .dout(n18024));
  jor  g17866(.dina(n18024), .dinb(n18021), .dout(n18025));
  jor  g17867(.dina(n18025), .dinb(n18020), .dout(n18026));
  jxor g17868(.dina(n18026), .dinb(n6039), .dout(n18027));
  jnot g17869(.din(n18027), .dout(n18028));
  jxor g17870(.dina(n17641), .dinb(n17640), .dout(n18029));
  jand g17871(.dina(n18029), .dinb(n18028), .dout(n18030));
  jxor g17872(.dina(n17638), .dinb(n17637), .dout(n18031));
  jnot g17873(.din(n18031), .dout(n18032));
  jor  g17874(.dina(n14221), .dinb(n8772), .dout(n18033));
  jor  g17875(.dina(n15045), .dinb(n9490), .dout(n18034));
  jor  g17876(.dina(n11984), .dinb(n9127), .dout(n18035));
  jor  g17877(.dina(n11987), .dinb(n8770), .dout(n18036));
  jand g17878(.dina(n18036), .dinb(n18035), .dout(n18037));
  jand g17879(.dina(n18037), .dinb(n18034), .dout(n18038));
  jand g17880(.dina(n18038), .dinb(n18033), .dout(n18039));
  jxor g17881(.dina(n18039), .dinb(\a[8] ), .dout(n18040));
  jor  g17882(.dina(n18040), .dinb(n18032), .dout(n18041));
  jxor g17883(.dina(n17635), .dinb(n17634), .dout(n18042));
  jnot g17884(.din(n18042), .dout(n18043));
  jor  g17885(.dina(n14248), .dinb(n8772), .dout(n18044));
  jor  g17886(.dina(n11984), .dinb(n9490), .dout(n18045));
  jor  g17887(.dina(n11987), .dinb(n9127), .dout(n18046));
  jor  g17888(.dina(n11991), .dinb(n8770), .dout(n18047));
  jand g17889(.dina(n18047), .dinb(n18046), .dout(n18048));
  jand g17890(.dina(n18048), .dinb(n18045), .dout(n18049));
  jand g17891(.dina(n18049), .dinb(n18044), .dout(n18050));
  jxor g17892(.dina(n18050), .dinb(\a[8] ), .dout(n18051));
  jor  g17893(.dina(n18051), .dinb(n18043), .dout(n18052));
  jxor g17894(.dina(n17632), .dinb(n17631), .dout(n18053));
  jnot g17895(.din(n18053), .dout(n18054));
  jor  g17896(.dina(n14271), .dinb(n8772), .dout(n18055));
  jor  g17897(.dina(n11987), .dinb(n9490), .dout(n18056));
  jor  g17898(.dina(n11991), .dinb(n9127), .dout(n18057));
  jor  g17899(.dina(n11995), .dinb(n8770), .dout(n18058));
  jand g17900(.dina(n18058), .dinb(n18057), .dout(n18059));
  jand g17901(.dina(n18059), .dinb(n18056), .dout(n18060));
  jand g17902(.dina(n18060), .dinb(n18055), .dout(n18061));
  jxor g17903(.dina(n18061), .dinb(\a[8] ), .dout(n18062));
  jor  g17904(.dina(n18062), .dinb(n18054), .dout(n18063));
  jor  g17905(.dina(n14301), .dinb(n8772), .dout(n18064));
  jor  g17906(.dina(n11991), .dinb(n9490), .dout(n18065));
  jor  g17907(.dina(n11995), .dinb(n9127), .dout(n18066));
  jor  g17908(.dina(n11997), .dinb(n8770), .dout(n18067));
  jand g17909(.dina(n18067), .dinb(n18066), .dout(n18068));
  jand g17910(.dina(n18068), .dinb(n18065), .dout(n18069));
  jand g17911(.dina(n18069), .dinb(n18064), .dout(n18070));
  jxor g17912(.dina(n18070), .dinb(\a[8] ), .dout(n18071));
  jnot g17913(.din(n18071), .dout(n18072));
  jxor g17914(.dina(n17629), .dinb(n17628), .dout(n18073));
  jand g17915(.dina(n18073), .dinb(n18072), .dout(n18074));
  jor  g17916(.dina(n14353), .dinb(n8772), .dout(n18075));
  jor  g17917(.dina(n11995), .dinb(n9490), .dout(n18076));
  jor  g17918(.dina(n11997), .dinb(n9127), .dout(n18077));
  jor  g17919(.dina(n11999), .dinb(n8770), .dout(n18078));
  jand g17920(.dina(n18078), .dinb(n18077), .dout(n18079));
  jand g17921(.dina(n18079), .dinb(n18076), .dout(n18080));
  jand g17922(.dina(n18080), .dinb(n18075), .dout(n18081));
  jxor g17923(.dina(n18081), .dinb(\a[8] ), .dout(n18082));
  jnot g17924(.din(n18082), .dout(n18083));
  jxor g17925(.dina(n17626), .dinb(n17625), .dout(n18084));
  jand g17926(.dina(n18084), .dinb(n18083), .dout(n18085));
  jor  g17927(.dina(n14390), .dinb(n8772), .dout(n18086));
  jor  g17928(.dina(n11997), .dinb(n9490), .dout(n18087));
  jor  g17929(.dina(n11999), .dinb(n9127), .dout(n18088));
  jor  g17930(.dina(n12001), .dinb(n8770), .dout(n18089));
  jand g17931(.dina(n18089), .dinb(n18088), .dout(n18090));
  jand g17932(.dina(n18090), .dinb(n18087), .dout(n18091));
  jand g17933(.dina(n18091), .dinb(n18086), .dout(n18092));
  jxor g17934(.dina(n18092), .dinb(\a[8] ), .dout(n18093));
  jnot g17935(.din(n18093), .dout(n18094));
  jor  g17936(.dina(n17606), .dinb(n5833), .dout(n18095));
  jxor g17937(.dina(n18095), .dinb(n17614), .dout(n18096));
  jand g17938(.dina(n18096), .dinb(n18094), .dout(n18097));
  jor  g17939(.dina(n14432), .dinb(n8772), .dout(n18098));
  jor  g17940(.dina(n11999), .dinb(n9490), .dout(n18099));
  jor  g17941(.dina(n12001), .dinb(n9127), .dout(n18100));
  jor  g17942(.dina(n12004), .dinb(n8770), .dout(n18101));
  jand g17943(.dina(n18101), .dinb(n18100), .dout(n18102));
  jand g17944(.dina(n18102), .dinb(n18099), .dout(n18103));
  jand g17945(.dina(n18103), .dinb(n18098), .dout(n18104));
  jxor g17946(.dina(n18104), .dinb(\a[8] ), .dout(n18105));
  jnot g17947(.din(n18105), .dout(n18106));
  jand g17948(.dina(n17603), .dinb(\a[11] ), .dout(n18107));
  jxor g17949(.dina(n18107), .dinb(n17601), .dout(n18108));
  jand g17950(.dina(n18108), .dinb(n18106), .dout(n18109));
  jand g17951(.dina(n14497), .dinb(n8771), .dout(n18110));
  jand g17952(.dina(n12010), .dinb(n9126), .dout(n18111));
  jand g17953(.dina(n12008), .dinb(n9491), .dout(n18112));
  jor  g17954(.dina(n18112), .dinb(n18111), .dout(n18113));
  jor  g17955(.dina(n18113), .dinb(n18110), .dout(n18114));
  jnot g17956(.din(n18114), .dout(n18115));
  jand g17957(.dina(n12010), .dinb(n8765), .dout(n18116));
  jnot g17958(.din(n18116), .dout(n18117));
  jand g17959(.dina(n18117), .dinb(\a[8] ), .dout(n18118));
  jand g17960(.dina(n18118), .dinb(n18115), .dout(n18119));
  jand g17961(.dina(n14537), .dinb(n8771), .dout(n18120));
  jand g17962(.dina(n12006), .dinb(n9491), .dout(n18121));
  jand g17963(.dina(n12008), .dinb(n9126), .dout(n18122));
  jand g17964(.dina(n12010), .dinb(n8769), .dout(n18123));
  jor  g17965(.dina(n18123), .dinb(n18122), .dout(n18124));
  jor  g17966(.dina(n18124), .dinb(n18121), .dout(n18125));
  jor  g17967(.dina(n18125), .dinb(n18120), .dout(n18126));
  jnot g17968(.din(n18126), .dout(n18127));
  jand g17969(.dina(n18127), .dinb(n18119), .dout(n18128));
  jand g17970(.dina(n18128), .dinb(n17603), .dout(n18129));
  jor  g17971(.dina(n15144), .dinb(n8772), .dout(n18130));
  jor  g17972(.dina(n12001), .dinb(n9490), .dout(n18131));
  jor  g17973(.dina(n12004), .dinb(n9127), .dout(n18132));
  jor  g17974(.dina(n12009), .dinb(n8770), .dout(n18133));
  jand g17975(.dina(n18133), .dinb(n18132), .dout(n18134));
  jand g17976(.dina(n18134), .dinb(n18131), .dout(n18135));
  jand g17977(.dina(n18135), .dinb(n18130), .dout(n18136));
  jxor g17978(.dina(n18136), .dinb(\a[8] ), .dout(n18137));
  jnot g17979(.din(n18137), .dout(n18138));
  jxor g17980(.dina(n18128), .dinb(n17603), .dout(n18139));
  jand g17981(.dina(n18139), .dinb(n18138), .dout(n18140));
  jor  g17982(.dina(n18140), .dinb(n18129), .dout(n18141));
  jxor g17983(.dina(n18108), .dinb(n18106), .dout(n18142));
  jand g17984(.dina(n18142), .dinb(n18141), .dout(n18143));
  jor  g17985(.dina(n18143), .dinb(n18109), .dout(n18144));
  jxor g17986(.dina(n18096), .dinb(n18094), .dout(n18145));
  jand g17987(.dina(n18145), .dinb(n18144), .dout(n18146));
  jor  g17988(.dina(n18146), .dinb(n18097), .dout(n18147));
  jxor g17989(.dina(n18084), .dinb(n18083), .dout(n18148));
  jand g17990(.dina(n18148), .dinb(n18147), .dout(n18149));
  jor  g17991(.dina(n18149), .dinb(n18085), .dout(n18150));
  jxor g17992(.dina(n18073), .dinb(n18072), .dout(n18151));
  jand g17993(.dina(n18151), .dinb(n18150), .dout(n18152));
  jor  g17994(.dina(n18152), .dinb(n18074), .dout(n18153));
  jxor g17995(.dina(n18062), .dinb(n18054), .dout(n18154));
  jand g17996(.dina(n18154), .dinb(n18153), .dout(n18155));
  jnot g17997(.din(n18155), .dout(n18156));
  jand g17998(.dina(n18156), .dinb(n18063), .dout(n18157));
  jnot g17999(.din(n18157), .dout(n18158));
  jxor g18000(.dina(n18051), .dinb(n18043), .dout(n18159));
  jand g18001(.dina(n18159), .dinb(n18158), .dout(n18160));
  jnot g18002(.din(n18160), .dout(n18161));
  jand g18003(.dina(n18161), .dinb(n18052), .dout(n18162));
  jnot g18004(.din(n18162), .dout(n18163));
  jxor g18005(.dina(n18040), .dinb(n18032), .dout(n18164));
  jand g18006(.dina(n18164), .dinb(n18163), .dout(n18165));
  jnot g18007(.din(n18165), .dout(n18166));
  jand g18008(.dina(n18166), .dinb(n18041), .dout(n18167));
  jnot g18009(.din(n18167), .dout(n18168));
  jxor g18010(.dina(n18029), .dinb(n18028), .dout(n18169));
  jand g18011(.dina(n18169), .dinb(n18168), .dout(n18170));
  jor  g18012(.dina(n18170), .dinb(n18030), .dout(n18171));
  jxor g18013(.dina(n18018), .dinb(n18017), .dout(n18172));
  jand g18014(.dina(n18172), .dinb(n18171), .dout(n18173));
  jor  g18015(.dina(n18173), .dinb(n18019), .dout(n18174));
  jxor g18016(.dina(n18007), .dinb(n18006), .dout(n18175));
  jand g18017(.dina(n18175), .dinb(n18174), .dout(n18176));
  jor  g18018(.dina(n18176), .dinb(n18008), .dout(n18177));
  jxor g18019(.dina(n17996), .dinb(n17988), .dout(n18178));
  jand g18020(.dina(n18178), .dinb(n18177), .dout(n18179));
  jnot g18021(.din(n18179), .dout(n18180));
  jand g18022(.dina(n18180), .dinb(n17997), .dout(n18181));
  jnot g18023(.din(n18181), .dout(n18182));
  jxor g18024(.dina(n17985), .dinb(n17977), .dout(n18183));
  jand g18025(.dina(n18183), .dinb(n18182), .dout(n18184));
  jnot g18026(.din(n18184), .dout(n18185));
  jand g18027(.dina(n18185), .dinb(n17986), .dout(n18186));
  jnot g18028(.din(n18186), .dout(n18187));
  jxor g18029(.dina(n17974), .dinb(n17966), .dout(n18188));
  jand g18030(.dina(n18188), .dinb(n18187), .dout(n18189));
  jnot g18031(.din(n18189), .dout(n18190));
  jand g18032(.dina(n18190), .dinb(n17975), .dout(n18191));
  jnot g18033(.din(n18191), .dout(n18192));
  jxor g18034(.dina(n17963), .dinb(n17962), .dout(n18193));
  jand g18035(.dina(n18193), .dinb(n18192), .dout(n18194));
  jor  g18036(.dina(n18194), .dinb(n17964), .dout(n18195));
  jxor g18037(.dina(n17952), .dinb(n17951), .dout(n18196));
  jand g18038(.dina(n18196), .dinb(n18195), .dout(n18197));
  jor  g18039(.dina(n18197), .dinb(n17953), .dout(n18198));
  jxor g18040(.dina(n17941), .dinb(n17940), .dout(n18199));
  jand g18041(.dina(n18199), .dinb(n18198), .dout(n18200));
  jor  g18042(.dina(n18200), .dinb(n17942), .dout(n18201));
  jxor g18043(.dina(n17930), .dinb(n17922), .dout(n18202));
  jand g18044(.dina(n18202), .dinb(n18201), .dout(n18203));
  jnot g18045(.din(n18203), .dout(n18204));
  jand g18046(.dina(n18204), .dinb(n17931), .dout(n18205));
  jnot g18047(.din(n18205), .dout(n18206));
  jxor g18048(.dina(n17919), .dinb(n17911), .dout(n18207));
  jand g18049(.dina(n18207), .dinb(n18206), .dout(n18208));
  jnot g18050(.din(n18208), .dout(n18209));
  jand g18051(.dina(n18209), .dinb(n17920), .dout(n18210));
  jnot g18052(.din(n18210), .dout(n18211));
  jxor g18053(.dina(n17908), .dinb(n17900), .dout(n18212));
  jand g18054(.dina(n18212), .dinb(n18211), .dout(n18213));
  jnot g18055(.din(n18213), .dout(n18214));
  jand g18056(.dina(n18214), .dinb(n17909), .dout(n18215));
  jnot g18057(.din(n18215), .dout(n18216));
  jxor g18058(.dina(n17897), .dinb(n17896), .dout(n18217));
  jand g18059(.dina(n18217), .dinb(n18216), .dout(n18218));
  jor  g18060(.dina(n18218), .dinb(n17898), .dout(n18219));
  jxor g18061(.dina(n17886), .dinb(n17885), .dout(n18220));
  jand g18062(.dina(n18220), .dinb(n18219), .dout(n18221));
  jor  g18063(.dina(n18221), .dinb(n17887), .dout(n18222));
  jxor g18064(.dina(n17875), .dinb(n17867), .dout(n18223));
  jand g18065(.dina(n18223), .dinb(n18222), .dout(n18224));
  jnot g18066(.din(n18224), .dout(n18225));
  jand g18067(.dina(n18225), .dinb(n17876), .dout(n18226));
  jnot g18068(.din(n18226), .dout(n18227));
  jxor g18069(.dina(n17864), .dinb(n17856), .dout(n18228));
  jand g18070(.dina(n18228), .dinb(n18227), .dout(n18229));
  jnot g18071(.din(n18229), .dout(n18230));
  jand g18072(.dina(n18230), .dinb(n17865), .dout(n18231));
  jnot g18073(.din(n18231), .dout(n18232));
  jxor g18074(.dina(n17853), .dinb(n17845), .dout(n18233));
  jand g18075(.dina(n18233), .dinb(n18232), .dout(n18234));
  jnot g18076(.din(n18234), .dout(n18235));
  jand g18077(.dina(n18235), .dinb(n17854), .dout(n18236));
  jnot g18078(.din(n18236), .dout(n18237));
  jxor g18079(.dina(n17842), .dinb(n17834), .dout(n18238));
  jand g18080(.dina(n18238), .dinb(n18237), .dout(n18239));
  jnot g18081(.din(n18239), .dout(n18240));
  jand g18082(.dina(n18240), .dinb(n17843), .dout(n18241));
  jnot g18083(.din(n18241), .dout(n18242));
  jxor g18084(.dina(n17831), .dinb(n17823), .dout(n18243));
  jand g18085(.dina(n18243), .dinb(n18242), .dout(n18244));
  jnot g18086(.din(n18244), .dout(n18245));
  jand g18087(.dina(n18245), .dinb(n17832), .dout(n18246));
  jnot g18088(.din(n18246), .dout(n18247));
  jxor g18089(.dina(n17820), .dinb(n17812), .dout(n18248));
  jand g18090(.dina(n18248), .dinb(n18247), .dout(n18249));
  jnot g18091(.din(n18249), .dout(n18250));
  jand g18092(.dina(n18250), .dinb(n17821), .dout(n18251));
  jnot g18093(.din(n18251), .dout(n18252));
  jxor g18094(.dina(n17809), .dinb(n17801), .dout(n18253));
  jand g18095(.dina(n18253), .dinb(n18252), .dout(n18254));
  jnot g18096(.din(n18254), .dout(n18255));
  jand g18097(.dina(n18255), .dinb(n17810), .dout(n18256));
  jnot g18098(.din(n18256), .dout(n18257));
  jxor g18099(.dina(n17797), .dinb(n17789), .dout(n18258));
  jand g18100(.dina(n18258), .dinb(n18257), .dout(n18259));
  jor  g18101(.dina(n18259), .dinb(n17799), .dout(n18260));
  jxor g18102(.dina(n17786), .dinb(n17778), .dout(n18261));
  jand g18103(.dina(n18261), .dinb(n18260), .dout(n18262));
  jnot g18104(.din(n18262), .dout(n18263));
  jand g18105(.dina(n18263), .dinb(n17787), .dout(n18264));
  jnot g18106(.din(n18264), .dout(n18265));
  jxor g18107(.dina(n17775), .dinb(n17767), .dout(n18266));
  jand g18108(.dina(n18266), .dinb(n18265), .dout(n18267));
  jnot g18109(.din(n18267), .dout(n18268));
  jand g18110(.dina(n18268), .dinb(n17776), .dout(n18269));
  jnot g18111(.din(n18269), .dout(n18270));
  jxor g18112(.dina(n17741), .dinb(n17733), .dout(n18271));
  jand g18113(.dina(n18271), .dinb(n18270), .dout(n18272));
  jnot g18114(.din(n18272), .dout(n18273));
  jxor g18115(.dina(n18271), .dinb(n18269), .dout(n18274));
  jand g18116(.dina(n13022), .dinb(n67), .dout(n18275));
  jand g18117(.dina(n12815), .dinb(n10350), .dout(n18277));
  jand g18118(.dina(n12795), .dinb(n9917), .dout(n18278));
  jor  g18119(.dina(n18278), .dinb(n18277), .dout(n18279));
  jor  g18120(.dina(n18279), .dinb(n10827), .dout(n18280));
  jor  g18121(.dina(n18280), .dinb(n18275), .dout(n18281));
  jxor g18122(.dina(n18281), .dinb(n64), .dout(n18282));
  jor  g18123(.dina(n18282), .dinb(n18274), .dout(n18283));
  jand g18124(.dina(n18283), .dinb(n18273), .dout(n18284));
  jnot g18125(.din(n18284), .dout(n18285));
  jxor g18126(.dina(n17757), .dinb(n17749), .dout(n18286));
  jand g18127(.dina(n18286), .dinb(n18285), .dout(n18287));
  jnot g18128(.din(n18287), .dout(n18288));
  jxor g18129(.dina(n18286), .dinb(n18285), .dout(n18289));
  jnot g18130(.din(n18289), .dout(n18290));
  jand g18131(.dina(n12919), .dinb(n67), .dout(n18291));
  jand g18132(.dina(n12815), .dinb(n10827), .dout(n18292));
  jand g18133(.dina(n12795), .dinb(n10350), .dout(n18293));
  jand g18134(.dina(n12782), .dinb(n9917), .dout(n18294));
  jor  g18135(.dina(n18294), .dinb(n18293), .dout(n18295));
  jor  g18136(.dina(n18295), .dinb(n18292), .dout(n18296));
  jor  g18137(.dina(n18296), .dinb(n18291), .dout(n18297));
  jxor g18138(.dina(n18297), .dinb(n64), .dout(n18298));
  jnot g18139(.din(n18298), .dout(n18299));
  jxor g18140(.dina(n18266), .dinb(n18265), .dout(n18300));
  jand g18141(.dina(n18300), .dinb(n18299), .dout(n18301));
  jxor g18142(.dina(n18300), .dinb(n18299), .dout(n18309));
  jand g18143(.dina(n18309), .dinb(n13649), .dout(n18310));
  jor  g18144(.dina(n18310), .dinb(n18301), .dout(n18311));
  jxor g18145(.dina(n18282), .dinb(n18274), .dout(n18312));
  jand g18146(.dina(n18312), .dinb(n18311), .dout(n18313));
  jnot g18147(.din(n18313), .dout(n18314));
  jxor g18148(.dina(n18312), .dinb(n18311), .dout(n18315));
  jnot g18149(.din(n18315), .dout(n18316));
  jand g18150(.dina(n12797), .dinb(n67), .dout(n18317));
  jand g18151(.dina(n12795), .dinb(n10827), .dout(n18318));
  jand g18152(.dina(n12782), .dinb(n10350), .dout(n18319));
  jand g18153(.dina(n12783), .dinb(n9917), .dout(n18320));
  jor  g18154(.dina(n18320), .dinb(n18319), .dout(n18321));
  jor  g18155(.dina(n18321), .dinb(n18318), .dout(n18322));
  jor  g18156(.dina(n18322), .dinb(n18317), .dout(n18323));
  jxor g18157(.dina(n18323), .dinb(n64), .dout(n18324));
  jnot g18158(.din(n18324), .dout(n18325));
  jxor g18159(.dina(n18261), .dinb(n18260), .dout(n18326));
  jand g18160(.dina(n18326), .dinb(n18325), .dout(n18327));
  jand g18161(.dina(n12938), .dinb(n67), .dout(n18328));
  jand g18162(.dina(n12782), .dinb(n10827), .dout(n18329));
  jand g18163(.dina(n12783), .dinb(n10350), .dout(n18330));
  jand g18164(.dina(n12766), .dinb(n9917), .dout(n18331));
  jor  g18165(.dina(n18331), .dinb(n18330), .dout(n18332));
  jor  g18166(.dina(n18332), .dinb(n18329), .dout(n18333));
  jor  g18167(.dina(n18333), .dinb(n18328), .dout(n18334));
  jxor g18168(.dina(n18334), .dinb(n64), .dout(n18335));
  jnot g18169(.din(n18335), .dout(n18336));
  jxor g18170(.dina(n18258), .dinb(n18257), .dout(n18337));
  jand g18171(.dina(n18337), .dinb(n18336), .dout(n18338));
  jand g18172(.dina(n12841), .dinb(n67), .dout(n18339));
  jand g18173(.dina(n12783), .dinb(n10827), .dout(n18340));
  jand g18174(.dina(n12766), .dinb(n10350), .dout(n18341));
  jand g18175(.dina(n12177), .dinb(n9917), .dout(n18342));
  jor  g18176(.dina(n18342), .dinb(n18341), .dout(n18343));
  jor  g18177(.dina(n18343), .dinb(n18340), .dout(n18344));
  jor  g18178(.dina(n18344), .dinb(n18339), .dout(n18345));
  jxor g18179(.dina(n18345), .dinb(n64), .dout(n18346));
  jnot g18180(.din(n18346), .dout(n18347));
  jxor g18181(.dina(n18253), .dinb(n18252), .dout(n18348));
  jand g18182(.dina(n18348), .dinb(n18347), .dout(n18349));
  jand g18183(.dina(n12768), .dinb(n67), .dout(n18350));
  jand g18184(.dina(n12766), .dinb(n10827), .dout(n18351));
  jand g18185(.dina(n12177), .dinb(n10350), .dout(n18352));
  jand g18186(.dina(n11941), .dinb(n9917), .dout(n18353));
  jor  g18187(.dina(n18353), .dinb(n18352), .dout(n18354));
  jor  g18188(.dina(n18354), .dinb(n18351), .dout(n18355));
  jor  g18189(.dina(n18355), .dinb(n18350), .dout(n18356));
  jxor g18190(.dina(n18356), .dinb(n64), .dout(n18357));
  jnot g18191(.din(n18357), .dout(n18358));
  jxor g18192(.dina(n18248), .dinb(n18247), .dout(n18359));
  jand g18193(.dina(n18359), .dinb(n18358), .dout(n18360));
  jand g18194(.dina(n12179), .dinb(n67), .dout(n18361));
  jand g18195(.dina(n12177), .dinb(n10827), .dout(n18362));
  jand g18196(.dina(n11941), .dinb(n10350), .dout(n18363));
  jand g18197(.dina(n11942), .dinb(n9917), .dout(n18364));
  jor  g18198(.dina(n18364), .dinb(n18363), .dout(n18365));
  jor  g18199(.dina(n18365), .dinb(n18362), .dout(n18366));
  jor  g18200(.dina(n18366), .dinb(n18361), .dout(n18367));
  jxor g18201(.dina(n18367), .dinb(n64), .dout(n18368));
  jnot g18202(.din(n18368), .dout(n18369));
  jxor g18203(.dina(n18243), .dinb(n18242), .dout(n18370));
  jand g18204(.dina(n18370), .dinb(n18369), .dout(n18371));
  jand g18205(.dina(n12671), .dinb(n67), .dout(n18372));
  jand g18206(.dina(n11941), .dinb(n10827), .dout(n18373));
  jand g18207(.dina(n11942), .dinb(n10350), .dout(n18374));
  jand g18208(.dina(n11944), .dinb(n9917), .dout(n18375));
  jor  g18209(.dina(n18375), .dinb(n18374), .dout(n18376));
  jor  g18210(.dina(n18376), .dinb(n18373), .dout(n18377));
  jor  g18211(.dina(n18377), .dinb(n18372), .dout(n18378));
  jxor g18212(.dina(n18378), .dinb(n64), .dout(n18379));
  jnot g18213(.din(n18379), .dout(n18380));
  jxor g18214(.dina(n18238), .dinb(n18237), .dout(n18381));
  jand g18215(.dina(n18381), .dinb(n18380), .dout(n18382));
  jand g18216(.dina(n12751), .dinb(n67), .dout(n18383));
  jand g18217(.dina(n11942), .dinb(n10827), .dout(n18384));
  jand g18218(.dina(n11944), .dinb(n10350), .dout(n18385));
  jand g18219(.dina(n11946), .dinb(n9917), .dout(n18386));
  jor  g18220(.dina(n18386), .dinb(n18385), .dout(n18387));
  jor  g18221(.dina(n18387), .dinb(n18384), .dout(n18388));
  jor  g18222(.dina(n18388), .dinb(n18383), .dout(n18389));
  jxor g18223(.dina(n18389), .dinb(n64), .dout(n18390));
  jnot g18224(.din(n18390), .dout(n18391));
  jxor g18225(.dina(n18233), .dinb(n18232), .dout(n18392));
  jand g18226(.dina(n18392), .dinb(n18391), .dout(n18393));
  jand g18227(.dina(n12189), .dinb(n67), .dout(n18394));
  jand g18228(.dina(n11944), .dinb(n10827), .dout(n18395));
  jand g18229(.dina(n11946), .dinb(n10350), .dout(n18396));
  jand g18230(.dina(n11948), .dinb(n9917), .dout(n18397));
  jor  g18231(.dina(n18397), .dinb(n18396), .dout(n18398));
  jor  g18232(.dina(n18398), .dinb(n18395), .dout(n18399));
  jor  g18233(.dina(n18399), .dinb(n18394), .dout(n18400));
  jxor g18234(.dina(n18400), .dinb(n64), .dout(n18401));
  jnot g18235(.din(n18401), .dout(n18402));
  jxor g18236(.dina(n18228), .dinb(n18227), .dout(n18403));
  jand g18237(.dina(n18403), .dinb(n18402), .dout(n18404));
  jand g18238(.dina(n12519), .dinb(n67), .dout(n18405));
  jand g18239(.dina(n11946), .dinb(n10827), .dout(n18406));
  jand g18240(.dina(n11948), .dinb(n10350), .dout(n18407));
  jand g18241(.dina(n11950), .dinb(n9917), .dout(n18408));
  jor  g18242(.dina(n18408), .dinb(n18407), .dout(n18409));
  jor  g18243(.dina(n18409), .dinb(n18406), .dout(n18410));
  jor  g18244(.dina(n18410), .dinb(n18405), .dout(n18411));
  jxor g18245(.dina(n18411), .dinb(n64), .dout(n18412));
  jnot g18246(.din(n18412), .dout(n18413));
  jxor g18247(.dina(n18223), .dinb(n18222), .dout(n18414));
  jand g18248(.dina(n18414), .dinb(n18413), .dout(n18415));
  jxor g18249(.dina(n18220), .dinb(n18219), .dout(n18416));
  jnot g18250(.din(n18416), .dout(n18417));
  jand g18251(.dina(n12654), .dinb(n67), .dout(n18418));
  jand g18252(.dina(n11948), .dinb(n10827), .dout(n18419));
  jand g18253(.dina(n11950), .dinb(n10350), .dout(n18420));
  jand g18254(.dina(n11952), .dinb(n9917), .dout(n18421));
  jor  g18255(.dina(n18421), .dinb(n18420), .dout(n18422));
  jor  g18256(.dina(n18422), .dinb(n18419), .dout(n18423));
  jor  g18257(.dina(n18423), .dinb(n18418), .dout(n18424));
  jxor g18258(.dina(n18424), .dinb(n64), .dout(n18425));
  jor  g18259(.dina(n18425), .dinb(n18417), .dout(n18426));
  jxor g18260(.dina(n18217), .dinb(n18216), .dout(n18427));
  jnot g18261(.din(n18427), .dout(n18428));
  jand g18262(.dina(n12569), .dinb(n67), .dout(n18429));
  jand g18263(.dina(n11950), .dinb(n10827), .dout(n18430));
  jand g18264(.dina(n11952), .dinb(n10350), .dout(n18431));
  jand g18265(.dina(n11954), .dinb(n9917), .dout(n18432));
  jor  g18266(.dina(n18432), .dinb(n18431), .dout(n18433));
  jor  g18267(.dina(n18433), .dinb(n18430), .dout(n18434));
  jor  g18268(.dina(n18434), .dinb(n18429), .dout(n18435));
  jxor g18269(.dina(n18435), .dinb(n64), .dout(n18436));
  jor  g18270(.dina(n18436), .dinb(n18428), .dout(n18437));
  jand g18271(.dina(n12510), .dinb(n67), .dout(n18438));
  jand g18272(.dina(n11952), .dinb(n10827), .dout(n18439));
  jand g18273(.dina(n11954), .dinb(n10350), .dout(n18440));
  jand g18274(.dina(n11956), .dinb(n9917), .dout(n18441));
  jor  g18275(.dina(n18441), .dinb(n18440), .dout(n18442));
  jor  g18276(.dina(n18442), .dinb(n18439), .dout(n18443));
  jor  g18277(.dina(n18443), .dinb(n18438), .dout(n18444));
  jxor g18278(.dina(n18444), .dinb(n64), .dout(n18445));
  jnot g18279(.din(n18445), .dout(n18446));
  jxor g18280(.dina(n18212), .dinb(n18211), .dout(n18447));
  jand g18281(.dina(n18447), .dinb(n18446), .dout(n18448));
  jand g18282(.dina(n12472), .dinb(n67), .dout(n18449));
  jand g18283(.dina(n11954), .dinb(n10827), .dout(n18450));
  jand g18284(.dina(n11956), .dinb(n10350), .dout(n18451));
  jand g18285(.dina(n11958), .dinb(n9917), .dout(n18452));
  jor  g18286(.dina(n18452), .dinb(n18451), .dout(n18453));
  jor  g18287(.dina(n18453), .dinb(n18450), .dout(n18454));
  jor  g18288(.dina(n18454), .dinb(n18449), .dout(n18455));
  jxor g18289(.dina(n18455), .dinb(n64), .dout(n18456));
  jnot g18290(.din(n18456), .dout(n18457));
  jxor g18291(.dina(n18207), .dinb(n18206), .dout(n18458));
  jand g18292(.dina(n18458), .dinb(n18457), .dout(n18459));
  jand g18293(.dina(n12639), .dinb(n67), .dout(n18460));
  jand g18294(.dina(n11956), .dinb(n10827), .dout(n18461));
  jand g18295(.dina(n11958), .dinb(n10350), .dout(n18462));
  jand g18296(.dina(n11960), .dinb(n9917), .dout(n18463));
  jor  g18297(.dina(n18463), .dinb(n18462), .dout(n18464));
  jor  g18298(.dina(n18464), .dinb(n18461), .dout(n18465));
  jor  g18299(.dina(n18465), .dinb(n18460), .dout(n18466));
  jxor g18300(.dina(n18466), .dinb(n64), .dout(n18467));
  jnot g18301(.din(n18467), .dout(n18468));
  jxor g18302(.dina(n18202), .dinb(n18201), .dout(n18469));
  jand g18303(.dina(n18469), .dinb(n18468), .dout(n18470));
  jxor g18304(.dina(n18199), .dinb(n18198), .dout(n18471));
  jnot g18305(.din(n18471), .dout(n18472));
  jand g18306(.dina(n12624), .dinb(n67), .dout(n18473));
  jand g18307(.dina(n11958), .dinb(n10827), .dout(n18474));
  jand g18308(.dina(n11960), .dinb(n10350), .dout(n18475));
  jand g18309(.dina(n11962), .dinb(n9917), .dout(n18476));
  jor  g18310(.dina(n18476), .dinb(n18475), .dout(n18477));
  jor  g18311(.dina(n18477), .dinb(n18474), .dout(n18478));
  jor  g18312(.dina(n18478), .dinb(n18473), .dout(n18479));
  jxor g18313(.dina(n18479), .dinb(n64), .dout(n18480));
  jor  g18314(.dina(n18480), .dinb(n18472), .dout(n18481));
  jxor g18315(.dina(n18196), .dinb(n18195), .dout(n18482));
  jnot g18316(.din(n18482), .dout(n18483));
  jand g18317(.dina(n13116), .dinb(n67), .dout(n18484));
  jand g18318(.dina(n11960), .dinb(n10827), .dout(n18485));
  jand g18319(.dina(n11962), .dinb(n10350), .dout(n18486));
  jand g18320(.dina(n11964), .dinb(n9917), .dout(n18487));
  jor  g18321(.dina(n18487), .dinb(n18486), .dout(n18488));
  jor  g18322(.dina(n18488), .dinb(n18485), .dout(n18489));
  jor  g18323(.dina(n18489), .dinb(n18484), .dout(n18490));
  jxor g18324(.dina(n18490), .dinb(n64), .dout(n18491));
  jor  g18325(.dina(n18491), .dinb(n18483), .dout(n18492));
  jxor g18326(.dina(n18193), .dinb(n18192), .dout(n18493));
  jnot g18327(.din(n18493), .dout(n18494));
  jand g18328(.dina(n13134), .dinb(n67), .dout(n18495));
  jand g18329(.dina(n11962), .dinb(n10827), .dout(n18496));
  jand g18330(.dina(n11964), .dinb(n10350), .dout(n18497));
  jand g18331(.dina(n11966), .dinb(n9917), .dout(n18498));
  jor  g18332(.dina(n18498), .dinb(n18497), .dout(n18499));
  jor  g18333(.dina(n18499), .dinb(n18496), .dout(n18500));
  jor  g18334(.dina(n18500), .dinb(n18495), .dout(n18501));
  jxor g18335(.dina(n18501), .dinb(n64), .dout(n18502));
  jor  g18336(.dina(n18502), .dinb(n18494), .dout(n18503));
  jand g18337(.dina(n13470), .dinb(n67), .dout(n18504));
  jand g18338(.dina(n11964), .dinb(n10827), .dout(n18505));
  jand g18339(.dina(n11966), .dinb(n10350), .dout(n18506));
  jand g18340(.dina(n11968), .dinb(n9917), .dout(n18507));
  jor  g18341(.dina(n18507), .dinb(n18506), .dout(n18508));
  jor  g18342(.dina(n18508), .dinb(n18505), .dout(n18509));
  jor  g18343(.dina(n18509), .dinb(n18504), .dout(n18510));
  jxor g18344(.dina(n18510), .dinb(n64), .dout(n18511));
  jnot g18345(.din(n18511), .dout(n18512));
  jxor g18346(.dina(n18188), .dinb(n18187), .dout(n18513));
  jand g18347(.dina(n18513), .dinb(n18512), .dout(n18514));
  jand g18348(.dina(n13268), .dinb(n67), .dout(n18515));
  jand g18349(.dina(n11966), .dinb(n10827), .dout(n18516));
  jand g18350(.dina(n11968), .dinb(n10350), .dout(n18517));
  jand g18351(.dina(n11970), .dinb(n9917), .dout(n18518));
  jor  g18352(.dina(n18518), .dinb(n18517), .dout(n18519));
  jor  g18353(.dina(n18519), .dinb(n18516), .dout(n18520));
  jor  g18354(.dina(n18520), .dinb(n18515), .dout(n18521));
  jxor g18355(.dina(n18521), .dinb(n64), .dout(n18522));
  jnot g18356(.din(n18522), .dout(n18523));
  jxor g18357(.dina(n18183), .dinb(n18182), .dout(n18524));
  jand g18358(.dina(n18524), .dinb(n18523), .dout(n18525));
  jand g18359(.dina(n13682), .dinb(n67), .dout(n18526));
  jand g18360(.dina(n11968), .dinb(n10827), .dout(n18527));
  jand g18361(.dina(n11970), .dinb(n10350), .dout(n18528));
  jand g18362(.dina(n11972), .dinb(n9917), .dout(n18529));
  jor  g18363(.dina(n18529), .dinb(n18528), .dout(n18530));
  jor  g18364(.dina(n18530), .dinb(n18527), .dout(n18531));
  jor  g18365(.dina(n18531), .dinb(n18526), .dout(n18532));
  jxor g18366(.dina(n18532), .dinb(n64), .dout(n18533));
  jnot g18367(.din(n18533), .dout(n18534));
  jxor g18368(.dina(n18178), .dinb(n18177), .dout(n18535));
  jand g18369(.dina(n18535), .dinb(n18534), .dout(n18536));
  jxor g18370(.dina(n18175), .dinb(n18174), .dout(n18537));
  jnot g18371(.din(n18537), .dout(n18538));
  jand g18372(.dina(n13806), .dinb(n67), .dout(n18539));
  jand g18373(.dina(n11970), .dinb(n10827), .dout(n18540));
  jand g18374(.dina(n11972), .dinb(n10350), .dout(n18541));
  jand g18375(.dina(n11974), .dinb(n9917), .dout(n18542));
  jor  g18376(.dina(n18542), .dinb(n18541), .dout(n18543));
  jor  g18377(.dina(n18543), .dinb(n18540), .dout(n18544));
  jor  g18378(.dina(n18544), .dinb(n18539), .dout(n18545));
  jxor g18379(.dina(n18545), .dinb(n64), .dout(n18546));
  jor  g18380(.dina(n18546), .dinb(n18538), .dout(n18547));
  jxor g18381(.dina(n18172), .dinb(n18171), .dout(n18548));
  jnot g18382(.din(n18548), .dout(n18549));
  jand g18383(.dina(n13664), .dinb(n67), .dout(n18550));
  jand g18384(.dina(n11972), .dinb(n10827), .dout(n18551));
  jand g18385(.dina(n11974), .dinb(n10350), .dout(n18552));
  jand g18386(.dina(n11976), .dinb(n9917), .dout(n18553));
  jor  g18387(.dina(n18553), .dinb(n18552), .dout(n18554));
  jor  g18388(.dina(n18554), .dinb(n18551), .dout(n18555));
  jor  g18389(.dina(n18555), .dinb(n18550), .dout(n18556));
  jxor g18390(.dina(n18556), .dinb(n64), .dout(n18557));
  jor  g18391(.dina(n18557), .dinb(n18549), .dout(n18558));
  jxor g18392(.dina(n18169), .dinb(n18168), .dout(n18559));
  jnot g18393(.din(n18559), .dout(n18560));
  jand g18394(.dina(n13924), .dinb(n67), .dout(n18561));
  jand g18395(.dina(n11974), .dinb(n10827), .dout(n18562));
  jand g18396(.dina(n11976), .dinb(n10350), .dout(n18563));
  jand g18397(.dina(n11978), .dinb(n9917), .dout(n18564));
  jor  g18398(.dina(n18564), .dinb(n18563), .dout(n18565));
  jor  g18399(.dina(n18565), .dinb(n18562), .dout(n18566));
  jor  g18400(.dina(n18566), .dinb(n18561), .dout(n18567));
  jxor g18401(.dina(n18567), .dinb(n64), .dout(n18568));
  jor  g18402(.dina(n18568), .dinb(n18560), .dout(n18569));
  jand g18403(.dina(n14184), .dinb(n67), .dout(n18570));
  jand g18404(.dina(n11976), .dinb(n10827), .dout(n18571));
  jand g18405(.dina(n11978), .dinb(n10350), .dout(n18572));
  jand g18406(.dina(n11980), .dinb(n9917), .dout(n18573));
  jor  g18407(.dina(n18573), .dinb(n18572), .dout(n18574));
  jor  g18408(.dina(n18574), .dinb(n18571), .dout(n18575));
  jor  g18409(.dina(n18575), .dinb(n18570), .dout(n18576));
  jxor g18410(.dina(n18576), .dinb(n64), .dout(n18577));
  jnot g18411(.din(n18577), .dout(n18578));
  jxor g18412(.dina(n18164), .dinb(n18163), .dout(n18579));
  jand g18413(.dina(n18579), .dinb(n18578), .dout(n18580));
  jand g18414(.dina(n14194), .dinb(n67), .dout(n18581));
  jand g18415(.dina(n11978), .dinb(n10827), .dout(n18582));
  jand g18416(.dina(n11980), .dinb(n10350), .dout(n18583));
  jand g18417(.dina(n11982), .dinb(n9917), .dout(n18584));
  jor  g18418(.dina(n18584), .dinb(n18583), .dout(n18585));
  jor  g18419(.dina(n18585), .dinb(n18582), .dout(n18586));
  jor  g18420(.dina(n18586), .dinb(n18581), .dout(n18587));
  jxor g18421(.dina(n18587), .dinb(n64), .dout(n18588));
  jnot g18422(.din(n18588), .dout(n18589));
  jxor g18423(.dina(n18159), .dinb(n18158), .dout(n18590));
  jand g18424(.dina(n18590), .dinb(n18589), .dout(n18591));
  jand g18425(.dina(n13899), .dinb(n67), .dout(n18592));
  jand g18426(.dina(n11980), .dinb(n10827), .dout(n18593));
  jand g18427(.dina(n11982), .dinb(n10350), .dout(n18594));
  jand g18428(.dina(n11985), .dinb(n9917), .dout(n18595));
  jor  g18429(.dina(n18595), .dinb(n18594), .dout(n18596));
  jor  g18430(.dina(n18596), .dinb(n18593), .dout(n18597));
  jor  g18431(.dina(n18597), .dinb(n18592), .dout(n18598));
  jxor g18432(.dina(n18598), .dinb(n64), .dout(n18599));
  jnot g18433(.din(n18599), .dout(n18600));
  jxor g18434(.dina(n18154), .dinb(n18153), .dout(n18601));
  jand g18435(.dina(n18601), .dinb(n18600), .dout(n18602));
  jxor g18436(.dina(n18151), .dinb(n18150), .dout(n18603));
  jnot g18437(.din(n18603), .dout(n18604));
  jor  g18438(.dina(n14221), .dinb(n9919), .dout(n18605));
  jor  g18439(.dina(n15045), .dinb(n10826), .dout(n18606));
  jor  g18440(.dina(n11984), .dinb(n10351), .dout(n18607));
  jor  g18441(.dina(n11987), .dinb(n9918), .dout(n18608));
  jand g18442(.dina(n18608), .dinb(n18607), .dout(n18609));
  jand g18443(.dina(n18609), .dinb(n18606), .dout(n18610));
  jand g18444(.dina(n18610), .dinb(n18605), .dout(n18611));
  jxor g18445(.dina(n18611), .dinb(\a[5] ), .dout(n18612));
  jor  g18446(.dina(n18612), .dinb(n18604), .dout(n18613));
  jxor g18447(.dina(n18148), .dinb(n18147), .dout(n18614));
  jnot g18448(.din(n18614), .dout(n18615));
  jor  g18449(.dina(n14248), .dinb(n9919), .dout(n18616));
  jor  g18450(.dina(n11984), .dinb(n10826), .dout(n18617));
  jor  g18451(.dina(n11987), .dinb(n10351), .dout(n18618));
  jor  g18452(.dina(n11991), .dinb(n9918), .dout(n18619));
  jand g18453(.dina(n18619), .dinb(n18618), .dout(n18620));
  jand g18454(.dina(n18620), .dinb(n18617), .dout(n18621));
  jand g18455(.dina(n18621), .dinb(n18616), .dout(n18622));
  jxor g18456(.dina(n18622), .dinb(\a[5] ), .dout(n18623));
  jor  g18457(.dina(n18623), .dinb(n18615), .dout(n18624));
  jxor g18458(.dina(n18145), .dinb(n18144), .dout(n18625));
  jnot g18459(.din(n18625), .dout(n18626));
  jor  g18460(.dina(n14271), .dinb(n9919), .dout(n18627));
  jor  g18461(.dina(n11987), .dinb(n10826), .dout(n18628));
  jor  g18462(.dina(n11991), .dinb(n10351), .dout(n18629));
  jor  g18463(.dina(n11995), .dinb(n9918), .dout(n18630));
  jand g18464(.dina(n18630), .dinb(n18629), .dout(n18631));
  jand g18465(.dina(n18631), .dinb(n18628), .dout(n18632));
  jand g18466(.dina(n18632), .dinb(n18627), .dout(n18633));
  jxor g18467(.dina(n18633), .dinb(\a[5] ), .dout(n18634));
  jor  g18468(.dina(n18634), .dinb(n18626), .dout(n18635));
  jor  g18469(.dina(n14301), .dinb(n9919), .dout(n18636));
  jor  g18470(.dina(n11991), .dinb(n10826), .dout(n18637));
  jor  g18471(.dina(n11995), .dinb(n10351), .dout(n18638));
  jor  g18472(.dina(n11997), .dinb(n9918), .dout(n18639));
  jand g18473(.dina(n18639), .dinb(n18638), .dout(n18640));
  jand g18474(.dina(n18640), .dinb(n18637), .dout(n18641));
  jand g18475(.dina(n18641), .dinb(n18636), .dout(n18642));
  jxor g18476(.dina(n18642), .dinb(\a[5] ), .dout(n18643));
  jnot g18477(.din(n18643), .dout(n18644));
  jxor g18478(.dina(n18142), .dinb(n18141), .dout(n18645));
  jand g18479(.dina(n18645), .dinb(n18644), .dout(n18646));
  jor  g18480(.dina(n14353), .dinb(n9919), .dout(n18647));
  jor  g18481(.dina(n11995), .dinb(n10826), .dout(n18648));
  jor  g18482(.dina(n11997), .dinb(n10351), .dout(n18649));
  jor  g18483(.dina(n11999), .dinb(n9918), .dout(n18650));
  jand g18484(.dina(n18650), .dinb(n18649), .dout(n18651));
  jand g18485(.dina(n18651), .dinb(n18648), .dout(n18652));
  jand g18486(.dina(n18652), .dinb(n18647), .dout(n18653));
  jxor g18487(.dina(n18653), .dinb(\a[5] ), .dout(n18654));
  jnot g18488(.din(n18654), .dout(n18655));
  jxor g18489(.dina(n18139), .dinb(n18138), .dout(n18656));
  jand g18490(.dina(n18656), .dinb(n18655), .dout(n18657));
  jor  g18491(.dina(n14390), .dinb(n9919), .dout(n18658));
  jor  g18492(.dina(n11997), .dinb(n10826), .dout(n18659));
  jor  g18493(.dina(n11999), .dinb(n10351), .dout(n18660));
  jor  g18494(.dina(n12001), .dinb(n9918), .dout(n18661));
  jand g18495(.dina(n18661), .dinb(n18660), .dout(n18662));
  jand g18496(.dina(n18662), .dinb(n18659), .dout(n18663));
  jand g18497(.dina(n18663), .dinb(n18658), .dout(n18664));
  jxor g18498(.dina(n18664), .dinb(\a[5] ), .dout(n18665));
  jnot g18499(.din(n18665), .dout(n18666));
  jor  g18500(.dina(n18119), .dinb(n6039), .dout(n18667));
  jxor g18501(.dina(n18667), .dinb(n18127), .dout(n18668));
  jand g18502(.dina(n18668), .dinb(n18666), .dout(n18669));
  jor  g18503(.dina(n14432), .dinb(n9919), .dout(n18670));
  jor  g18504(.dina(n11999), .dinb(n10826), .dout(n18671));
  jor  g18505(.dina(n12001), .dinb(n10351), .dout(n18672));
  jor  g18506(.dina(n12004), .dinb(n9918), .dout(n18673));
  jand g18507(.dina(n18673), .dinb(n18672), .dout(n18674));
  jand g18508(.dina(n18674), .dinb(n18671), .dout(n18675));
  jand g18509(.dina(n18675), .dinb(n18670), .dout(n18676));
  jxor g18510(.dina(n18676), .dinb(\a[5] ), .dout(n18677));
  jnot g18511(.din(n18677), .dout(n18678));
  jand g18512(.dina(n18116), .dinb(\a[8] ), .dout(n18679));
  jxor g18513(.dina(n18679), .dinb(n18114), .dout(n18680));
  jand g18514(.dina(n18680), .dinb(n18678), .dout(n18681));
  jand g18515(.dina(n14497), .dinb(n67), .dout(n18682));
  jand g18516(.dina(n12010), .dinb(n10350), .dout(n18683));
  jand g18517(.dina(n12008), .dinb(n10827), .dout(n18684));
  jor  g18518(.dina(n18684), .dinb(n18683), .dout(n18685));
  jor  g18519(.dina(n18685), .dinb(n18682), .dout(n18686));
  jnot g18520(.din(n18686), .dout(n18687));
  jand g18521(.dina(n12010), .dinb(n65), .dout(n18688));
  jnot g18522(.din(n18688), .dout(n18689));
  jand g18523(.dina(n18689), .dinb(\a[5] ), .dout(n18690));
  jand g18524(.dina(n18690), .dinb(n18687), .dout(n18691));
  jand g18525(.dina(n14537), .dinb(n67), .dout(n18692));
  jand g18526(.dina(n12006), .dinb(n10827), .dout(n18693));
  jand g18527(.dina(n12008), .dinb(n10350), .dout(n18694));
  jand g18528(.dina(n12010), .dinb(n9917), .dout(n18695));
  jor  g18529(.dina(n18695), .dinb(n18694), .dout(n18696));
  jor  g18530(.dina(n18696), .dinb(n18693), .dout(n18697));
  jor  g18531(.dina(n18697), .dinb(n18692), .dout(n18698));
  jnot g18532(.din(n18698), .dout(n18699));
  jand g18533(.dina(n18699), .dinb(n18691), .dout(n18700));
  jand g18534(.dina(n18700), .dinb(n18116), .dout(n18701));
  jor  g18535(.dina(n15144), .dinb(n9919), .dout(n18702));
  jor  g18536(.dina(n12001), .dinb(n10826), .dout(n18703));
  jor  g18537(.dina(n12004), .dinb(n10351), .dout(n18704));
  jor  g18538(.dina(n12009), .dinb(n9918), .dout(n18705));
  jand g18539(.dina(n18705), .dinb(n18704), .dout(n18706));
  jand g18540(.dina(n18706), .dinb(n18703), .dout(n18707));
  jand g18541(.dina(n18707), .dinb(n18702), .dout(n18708));
  jxor g18542(.dina(n18708), .dinb(\a[5] ), .dout(n18709));
  jnot g18543(.din(n18709), .dout(n18710));
  jxor g18544(.dina(n18700), .dinb(n18116), .dout(n18711));
  jand g18545(.dina(n18711), .dinb(n18710), .dout(n18712));
  jor  g18546(.dina(n18712), .dinb(n18701), .dout(n18713));
  jxor g18547(.dina(n18680), .dinb(n18678), .dout(n18714));
  jand g18548(.dina(n18714), .dinb(n18713), .dout(n18715));
  jor  g18549(.dina(n18715), .dinb(n18681), .dout(n18716));
  jxor g18550(.dina(n18668), .dinb(n18666), .dout(n18717));
  jand g18551(.dina(n18717), .dinb(n18716), .dout(n18718));
  jor  g18552(.dina(n18718), .dinb(n18669), .dout(n18719));
  jxor g18553(.dina(n18656), .dinb(n18655), .dout(n18720));
  jand g18554(.dina(n18720), .dinb(n18719), .dout(n18721));
  jor  g18555(.dina(n18721), .dinb(n18657), .dout(n18722));
  jxor g18556(.dina(n18645), .dinb(n18644), .dout(n18723));
  jand g18557(.dina(n18723), .dinb(n18722), .dout(n18724));
  jor  g18558(.dina(n18724), .dinb(n18646), .dout(n18725));
  jxor g18559(.dina(n18634), .dinb(n18626), .dout(n18726));
  jand g18560(.dina(n18726), .dinb(n18725), .dout(n18727));
  jnot g18561(.din(n18727), .dout(n18728));
  jand g18562(.dina(n18728), .dinb(n18635), .dout(n18729));
  jnot g18563(.din(n18729), .dout(n18730));
  jxor g18564(.dina(n18623), .dinb(n18615), .dout(n18731));
  jand g18565(.dina(n18731), .dinb(n18730), .dout(n18732));
  jnot g18566(.din(n18732), .dout(n18733));
  jand g18567(.dina(n18733), .dinb(n18624), .dout(n18734));
  jnot g18568(.din(n18734), .dout(n18735));
  jxor g18569(.dina(n18612), .dinb(n18604), .dout(n18736));
  jand g18570(.dina(n18736), .dinb(n18735), .dout(n18737));
  jnot g18571(.din(n18737), .dout(n18738));
  jand g18572(.dina(n18738), .dinb(n18613), .dout(n18739));
  jnot g18573(.din(n18739), .dout(n18740));
  jxor g18574(.dina(n18601), .dinb(n18600), .dout(n18741));
  jand g18575(.dina(n18741), .dinb(n18740), .dout(n18742));
  jor  g18576(.dina(n18742), .dinb(n18602), .dout(n18743));
  jxor g18577(.dina(n18590), .dinb(n18589), .dout(n18744));
  jand g18578(.dina(n18744), .dinb(n18743), .dout(n18745));
  jor  g18579(.dina(n18745), .dinb(n18591), .dout(n18746));
  jxor g18580(.dina(n18579), .dinb(n18578), .dout(n18747));
  jand g18581(.dina(n18747), .dinb(n18746), .dout(n18748));
  jor  g18582(.dina(n18748), .dinb(n18580), .dout(n18749));
  jxor g18583(.dina(n18568), .dinb(n18560), .dout(n18750));
  jand g18584(.dina(n18750), .dinb(n18749), .dout(n18751));
  jnot g18585(.din(n18751), .dout(n18752));
  jand g18586(.dina(n18752), .dinb(n18569), .dout(n18753));
  jnot g18587(.din(n18753), .dout(n18754));
  jxor g18588(.dina(n18557), .dinb(n18549), .dout(n18755));
  jand g18589(.dina(n18755), .dinb(n18754), .dout(n18756));
  jnot g18590(.din(n18756), .dout(n18757));
  jand g18591(.dina(n18757), .dinb(n18558), .dout(n18758));
  jnot g18592(.din(n18758), .dout(n18759));
  jxor g18593(.dina(n18546), .dinb(n18538), .dout(n18760));
  jand g18594(.dina(n18760), .dinb(n18759), .dout(n18761));
  jnot g18595(.din(n18761), .dout(n18762));
  jand g18596(.dina(n18762), .dinb(n18547), .dout(n18763));
  jnot g18597(.din(n18763), .dout(n18764));
  jxor g18598(.dina(n18535), .dinb(n18534), .dout(n18765));
  jand g18599(.dina(n18765), .dinb(n18764), .dout(n18766));
  jor  g18600(.dina(n18766), .dinb(n18536), .dout(n18767));
  jxor g18601(.dina(n18524), .dinb(n18523), .dout(n18768));
  jand g18602(.dina(n18768), .dinb(n18767), .dout(n18769));
  jor  g18603(.dina(n18769), .dinb(n18525), .dout(n18770));
  jxor g18604(.dina(n18513), .dinb(n18512), .dout(n18771));
  jand g18605(.dina(n18771), .dinb(n18770), .dout(n18772));
  jor  g18606(.dina(n18772), .dinb(n18514), .dout(n18773));
  jxor g18607(.dina(n18502), .dinb(n18494), .dout(n18774));
  jand g18608(.dina(n18774), .dinb(n18773), .dout(n18775));
  jnot g18609(.din(n18775), .dout(n18776));
  jand g18610(.dina(n18776), .dinb(n18503), .dout(n18777));
  jnot g18611(.din(n18777), .dout(n18778));
  jxor g18612(.dina(n18491), .dinb(n18483), .dout(n18779));
  jand g18613(.dina(n18779), .dinb(n18778), .dout(n18780));
  jnot g18614(.din(n18780), .dout(n18781));
  jand g18615(.dina(n18781), .dinb(n18492), .dout(n18782));
  jnot g18616(.din(n18782), .dout(n18783));
  jxor g18617(.dina(n18480), .dinb(n18472), .dout(n18784));
  jand g18618(.dina(n18784), .dinb(n18783), .dout(n18785));
  jnot g18619(.din(n18785), .dout(n18786));
  jand g18620(.dina(n18786), .dinb(n18481), .dout(n18787));
  jnot g18621(.din(n18787), .dout(n18788));
  jxor g18622(.dina(n18469), .dinb(n18468), .dout(n18789));
  jand g18623(.dina(n18789), .dinb(n18788), .dout(n18790));
  jor  g18624(.dina(n18790), .dinb(n18470), .dout(n18791));
  jxor g18625(.dina(n18458), .dinb(n18457), .dout(n18792));
  jand g18626(.dina(n18792), .dinb(n18791), .dout(n18793));
  jor  g18627(.dina(n18793), .dinb(n18459), .dout(n18794));
  jxor g18628(.dina(n18447), .dinb(n18446), .dout(n18795));
  jand g18629(.dina(n18795), .dinb(n18794), .dout(n18796));
  jor  g18630(.dina(n18796), .dinb(n18448), .dout(n18797));
  jxor g18631(.dina(n18436), .dinb(n18428), .dout(n18798));
  jand g18632(.dina(n18798), .dinb(n18797), .dout(n18799));
  jnot g18633(.din(n18799), .dout(n18800));
  jand g18634(.dina(n18800), .dinb(n18437), .dout(n18801));
  jnot g18635(.din(n18801), .dout(n18802));
  jxor g18636(.dina(n18425), .dinb(n18417), .dout(n18803));
  jand g18637(.dina(n18803), .dinb(n18802), .dout(n18804));
  jnot g18638(.din(n18804), .dout(n18805));
  jand g18639(.dina(n18805), .dinb(n18426), .dout(n18806));
  jnot g18640(.din(n18806), .dout(n18807));
  jxor g18641(.dina(n18414), .dinb(n18413), .dout(n18808));
  jand g18642(.dina(n18808), .dinb(n18807), .dout(n18809));
  jor  g18643(.dina(n18809), .dinb(n18415), .dout(n18810));
  jxor g18644(.dina(n18403), .dinb(n18402), .dout(n18811));
  jand g18645(.dina(n18811), .dinb(n18810), .dout(n18812));
  jor  g18646(.dina(n18812), .dinb(n18404), .dout(n18813));
  jxor g18647(.dina(n18392), .dinb(n18391), .dout(n18814));
  jand g18648(.dina(n18814), .dinb(n18813), .dout(n18815));
  jor  g18649(.dina(n18815), .dinb(n18393), .dout(n18816));
  jxor g18650(.dina(n18381), .dinb(n18380), .dout(n18817));
  jand g18651(.dina(n18817), .dinb(n18816), .dout(n18818));
  jor  g18652(.dina(n18818), .dinb(n18382), .dout(n18819));
  jxor g18653(.dina(n18370), .dinb(n18369), .dout(n18820));
  jand g18654(.dina(n18820), .dinb(n18819), .dout(n18821));
  jor  g18655(.dina(n18821), .dinb(n18371), .dout(n18822));
  jxor g18656(.dina(n18359), .dinb(n18358), .dout(n18823));
  jand g18657(.dina(n18823), .dinb(n18822), .dout(n18824));
  jor  g18658(.dina(n18824), .dinb(n18360), .dout(n18825));
  jxor g18659(.dina(n18348), .dinb(n18347), .dout(n18826));
  jand g18660(.dina(n18826), .dinb(n18825), .dout(n18827));
  jor  g18661(.dina(n18827), .dinb(n18349), .dout(n18828));
  jxor g18662(.dina(n18337), .dinb(n18336), .dout(n18829));
  jand g18663(.dina(n18829), .dinb(n18828), .dout(n18830));
  jor  g18664(.dina(n18830), .dinb(n18338), .dout(n18831));
  jxor g18665(.dina(n18326), .dinb(n18325), .dout(n18832));
  jand g18666(.dina(n18832), .dinb(n18831), .dout(n18833));
  jor  g18667(.dina(n18833), .dinb(n18327), .dout(n18834));
  jxor g18668(.dina(n18309), .dinb(n13649), .dout(n18835));
  jand g18669(.dina(n18835), .dinb(n18834), .dout(n18836));
  jnot g18670(.din(n18836), .dout(n18837));
  jxor g18671(.dina(n18835), .dinb(n18834), .dout(n18838));
  jnot g18672(.din(n18838), .dout(n18839));
  jxor g18673(.dina(n18832), .dinb(n18831), .dout(n18840));
  jnot g18674(.din(n18840), .dout(n18841));
  jand g18675(.dina(n12815), .dinb(n10844), .dout(n18843));
  jor  g18676(.dina(n11470), .dinb(n18843), .dout(n18847));
  jor  g18677(.dina(n18847), .dinb(n10846), .dout(n18848));
  jxor g18678(.dina(n18848), .dinb(n6600), .dout(n18849));
  jor  g18679(.dina(n18849), .dinb(n18841), .dout(n18850));
  jxor g18680(.dina(n18829), .dinb(n18828), .dout(n18851));
  jnot g18681(.din(n18851), .dout(n18852));
  jand g18682(.dina(n13022), .dinb(n10846), .dout(n18853));
  jand g18683(.dina(n12815), .dinb(n11359), .dout(n18855));
  jand g18684(.dina(n12795), .dinb(n10844), .dout(n18856));
  jor  g18685(.dina(n18856), .dinb(n18855), .dout(n18857));
  jor  g18686(.dina(n18857), .dinb(n11372), .dout(n18858));
  jor  g18687(.dina(n18858), .dinb(n18853), .dout(n18859));
  jxor g18688(.dina(n18859), .dinb(n6600), .dout(n18860));
  jor  g18689(.dina(n18860), .dinb(n18852), .dout(n18861));
  jxor g18690(.dina(n18826), .dinb(n18825), .dout(n18862));
  jnot g18691(.din(n18862), .dout(n18863));
  jand g18692(.dina(n12919), .dinb(n10846), .dout(n18864));
  jand g18693(.dina(n12815), .dinb(n11372), .dout(n18865));
  jand g18694(.dina(n12795), .dinb(n11359), .dout(n18866));
  jand g18695(.dina(n12782), .dinb(n10844), .dout(n18867));
  jor  g18696(.dina(n18867), .dinb(n18866), .dout(n18868));
  jor  g18697(.dina(n18868), .dinb(n18865), .dout(n18869));
  jor  g18698(.dina(n18869), .dinb(n18864), .dout(n18870));
  jxor g18699(.dina(n18870), .dinb(n6600), .dout(n18871));
  jor  g18700(.dina(n18871), .dinb(n18863), .dout(n18872));
  jxor g18701(.dina(n18823), .dinb(n18822), .dout(n18873));
  jnot g18702(.din(n18873), .dout(n18874));
  jand g18703(.dina(n12797), .dinb(n10846), .dout(n18875));
  jand g18704(.dina(n12795), .dinb(n11372), .dout(n18876));
  jand g18705(.dina(n12782), .dinb(n11359), .dout(n18877));
  jand g18706(.dina(n12783), .dinb(n10844), .dout(n18878));
  jor  g18707(.dina(n18878), .dinb(n18877), .dout(n18879));
  jor  g18708(.dina(n18879), .dinb(n18876), .dout(n18880));
  jor  g18709(.dina(n18880), .dinb(n18875), .dout(n18881));
  jxor g18710(.dina(n18881), .dinb(n6600), .dout(n18882));
  jor  g18711(.dina(n18882), .dinb(n18874), .dout(n18883));
  jxor g18712(.dina(n18820), .dinb(n18819), .dout(n18884));
  jnot g18713(.din(n18884), .dout(n18885));
  jand g18714(.dina(n12938), .dinb(n10846), .dout(n18886));
  jand g18715(.dina(n12782), .dinb(n11372), .dout(n18887));
  jand g18716(.dina(n12783), .dinb(n11359), .dout(n18888));
  jand g18717(.dina(n12766), .dinb(n10844), .dout(n18889));
  jor  g18718(.dina(n18889), .dinb(n18888), .dout(n18890));
  jor  g18719(.dina(n18890), .dinb(n18887), .dout(n18891));
  jor  g18720(.dina(n18891), .dinb(n18886), .dout(n18892));
  jxor g18721(.dina(n18892), .dinb(n6600), .dout(n18893));
  jor  g18722(.dina(n18893), .dinb(n18885), .dout(n18894));
  jxor g18723(.dina(n18817), .dinb(n18816), .dout(n18895));
  jnot g18724(.din(n18895), .dout(n18896));
  jand g18725(.dina(n12841), .dinb(n10846), .dout(n18897));
  jand g18726(.dina(n12783), .dinb(n11372), .dout(n18898));
  jand g18727(.dina(n12766), .dinb(n11359), .dout(n18899));
  jand g18728(.dina(n12177), .dinb(n10844), .dout(n18900));
  jor  g18729(.dina(n18900), .dinb(n18899), .dout(n18901));
  jor  g18730(.dina(n18901), .dinb(n18898), .dout(n18902));
  jor  g18731(.dina(n18902), .dinb(n18897), .dout(n18903));
  jxor g18732(.dina(n18903), .dinb(n6600), .dout(n18904));
  jor  g18733(.dina(n18904), .dinb(n18896), .dout(n18905));
  jxor g18734(.dina(n18814), .dinb(n18813), .dout(n18906));
  jnot g18735(.din(n18906), .dout(n18907));
  jand g18736(.dina(n12768), .dinb(n10846), .dout(n18908));
  jand g18737(.dina(n12766), .dinb(n11372), .dout(n18909));
  jand g18738(.dina(n12177), .dinb(n11359), .dout(n18910));
  jand g18739(.dina(n11941), .dinb(n10844), .dout(n18911));
  jor  g18740(.dina(n18911), .dinb(n18910), .dout(n18912));
  jor  g18741(.dina(n18912), .dinb(n18909), .dout(n18913));
  jor  g18742(.dina(n18913), .dinb(n18908), .dout(n18914));
  jxor g18743(.dina(n18914), .dinb(n6600), .dout(n18915));
  jor  g18744(.dina(n18915), .dinb(n18907), .dout(n18916));
  jxor g18745(.dina(n18811), .dinb(n18810), .dout(n18917));
  jnot g18746(.din(n18917), .dout(n18918));
  jand g18747(.dina(n12179), .dinb(n10846), .dout(n18919));
  jand g18748(.dina(n12177), .dinb(n11372), .dout(n18920));
  jand g18749(.dina(n11941), .dinb(n11359), .dout(n18921));
  jand g18750(.dina(n11942), .dinb(n10844), .dout(n18922));
  jor  g18751(.dina(n18922), .dinb(n18921), .dout(n18923));
  jor  g18752(.dina(n18923), .dinb(n18920), .dout(n18924));
  jor  g18753(.dina(n18924), .dinb(n18919), .dout(n18925));
  jxor g18754(.dina(n18925), .dinb(n6600), .dout(n18926));
  jor  g18755(.dina(n18926), .dinb(n18918), .dout(n18927));
  jxor g18756(.dina(n18808), .dinb(n18807), .dout(n18928));
  jnot g18757(.din(n18928), .dout(n18929));
  jand g18758(.dina(n12671), .dinb(n10846), .dout(n18930));
  jand g18759(.dina(n11941), .dinb(n11372), .dout(n18931));
  jand g18760(.dina(n11942), .dinb(n11359), .dout(n18932));
  jand g18761(.dina(n11944), .dinb(n10844), .dout(n18933));
  jor  g18762(.dina(n18933), .dinb(n18932), .dout(n18934));
  jor  g18763(.dina(n18934), .dinb(n18931), .dout(n18935));
  jor  g18764(.dina(n18935), .dinb(n18930), .dout(n18936));
  jxor g18765(.dina(n18936), .dinb(n6600), .dout(n18937));
  jor  g18766(.dina(n18937), .dinb(n18929), .dout(n18938));
  jxor g18767(.dina(n18937), .dinb(n18929), .dout(n18939));
  jnot g18768(.din(n18939), .dout(n18940));
  jxor g18769(.dina(n18803), .dinb(n18802), .dout(n18941));
  jnot g18770(.din(n18941), .dout(n18942));
  jxor g18771(.dina(n18798), .dinb(n18797), .dout(n18943));
  jnot g18772(.din(n18943), .dout(n18944));
  jand g18773(.dina(n12519), .dinb(n10846), .dout(n18945));
  jand g18774(.dina(n11946), .dinb(n11372), .dout(n18946));
  jand g18775(.dina(n11948), .dinb(n11359), .dout(n18947));
  jand g18776(.dina(n11950), .dinb(n10844), .dout(n18948));
  jor  g18777(.dina(n18948), .dinb(n18947), .dout(n18949));
  jor  g18778(.dina(n18949), .dinb(n18946), .dout(n18950));
  jor  g18779(.dina(n18950), .dinb(n18945), .dout(n18951));
  jxor g18780(.dina(n18951), .dinb(n6600), .dout(n18952));
  jand g18781(.dina(n12654), .dinb(n10846), .dout(n18953));
  jand g18782(.dina(n11948), .dinb(n11372), .dout(n18954));
  jand g18783(.dina(n11950), .dinb(n11359), .dout(n18955));
  jand g18784(.dina(n11952), .dinb(n10844), .dout(n18956));
  jor  g18785(.dina(n18956), .dinb(n18955), .dout(n18957));
  jor  g18786(.dina(n18957), .dinb(n18954), .dout(n18958));
  jor  g18787(.dina(n18958), .dinb(n18953), .dout(n18959));
  jxor g18788(.dina(n18959), .dinb(n6600), .dout(n18960));
  jand g18789(.dina(n12569), .dinb(n10846), .dout(n18961));
  jand g18790(.dina(n11950), .dinb(n11372), .dout(n18962));
  jand g18791(.dina(n11952), .dinb(n11359), .dout(n18963));
  jand g18792(.dina(n11954), .dinb(n10844), .dout(n18964));
  jor  g18793(.dina(n18964), .dinb(n18963), .dout(n18965));
  jor  g18794(.dina(n18965), .dinb(n18962), .dout(n18966));
  jor  g18795(.dina(n18966), .dinb(n18961), .dout(n18967));
  jxor g18796(.dina(n18967), .dinb(n6600), .dout(n18968));
  jxor g18797(.dina(n18784), .dinb(n18783), .dout(n18969));
  jnot g18798(.din(n18969), .dout(n18970));
  jxor g18799(.dina(n18779), .dinb(n18778), .dout(n18971));
  jnot g18800(.din(n18971), .dout(n18972));
  jxor g18801(.dina(n18774), .dinb(n18773), .dout(n18973));
  jnot g18802(.din(n18973), .dout(n18974));
  jand g18803(.dina(n12624), .dinb(n10846), .dout(n18975));
  jand g18804(.dina(n11958), .dinb(n11372), .dout(n18976));
  jand g18805(.dina(n11960), .dinb(n11359), .dout(n18977));
  jand g18806(.dina(n11962), .dinb(n10844), .dout(n18978));
  jor  g18807(.dina(n18978), .dinb(n18977), .dout(n18979));
  jor  g18808(.dina(n18979), .dinb(n18976), .dout(n18980));
  jor  g18809(.dina(n18980), .dinb(n18975), .dout(n18981));
  jxor g18810(.dina(n18981), .dinb(n6600), .dout(n18982));
  jand g18811(.dina(n13116), .dinb(n10846), .dout(n18983));
  jand g18812(.dina(n11960), .dinb(n11372), .dout(n18984));
  jand g18813(.dina(n11962), .dinb(n11359), .dout(n18985));
  jand g18814(.dina(n11964), .dinb(n10844), .dout(n18986));
  jor  g18815(.dina(n18986), .dinb(n18985), .dout(n18987));
  jor  g18816(.dina(n18987), .dinb(n18984), .dout(n18988));
  jor  g18817(.dina(n18988), .dinb(n18983), .dout(n18989));
  jxor g18818(.dina(n18989), .dinb(n6600), .dout(n18990));
  jand g18819(.dina(n13134), .dinb(n10846), .dout(n18991));
  jand g18820(.dina(n11962), .dinb(n11372), .dout(n18992));
  jand g18821(.dina(n11964), .dinb(n11359), .dout(n18993));
  jand g18822(.dina(n11966), .dinb(n10844), .dout(n18994));
  jor  g18823(.dina(n18994), .dinb(n18993), .dout(n18995));
  jor  g18824(.dina(n18995), .dinb(n18992), .dout(n18996));
  jor  g18825(.dina(n18996), .dinb(n18991), .dout(n18997));
  jxor g18826(.dina(n18997), .dinb(n6600), .dout(n18998));
  jxor g18827(.dina(n18760), .dinb(n18759), .dout(n18999));
  jnot g18828(.din(n18999), .dout(n19000));
  jxor g18829(.dina(n18755), .dinb(n18754), .dout(n19001));
  jnot g18830(.din(n19001), .dout(n19002));
  jxor g18831(.dina(n18750), .dinb(n18749), .dout(n19003));
  jnot g18832(.din(n19003), .dout(n19004));
  jand g18833(.dina(n13806), .dinb(n10846), .dout(n19005));
  jand g18834(.dina(n11970), .dinb(n11372), .dout(n19006));
  jand g18835(.dina(n11972), .dinb(n11359), .dout(n19007));
  jand g18836(.dina(n11974), .dinb(n10844), .dout(n19008));
  jor  g18837(.dina(n19008), .dinb(n19007), .dout(n19009));
  jor  g18838(.dina(n19009), .dinb(n19006), .dout(n19010));
  jor  g18839(.dina(n19010), .dinb(n19005), .dout(n19011));
  jxor g18840(.dina(n19011), .dinb(n6600), .dout(n19012));
  jand g18841(.dina(n13664), .dinb(n10846), .dout(n19013));
  jand g18842(.dina(n11972), .dinb(n11372), .dout(n19014));
  jand g18843(.dina(n11974), .dinb(n11359), .dout(n19015));
  jand g18844(.dina(n11976), .dinb(n10844), .dout(n19016));
  jor  g18845(.dina(n19016), .dinb(n19015), .dout(n19017));
  jor  g18846(.dina(n19017), .dinb(n19014), .dout(n19018));
  jor  g18847(.dina(n19018), .dinb(n19013), .dout(n19019));
  jxor g18848(.dina(n19019), .dinb(n6600), .dout(n19020));
  jand g18849(.dina(n13924), .dinb(n10846), .dout(n19021));
  jand g18850(.dina(n11974), .dinb(n11372), .dout(n19022));
  jand g18851(.dina(n11976), .dinb(n11359), .dout(n19023));
  jand g18852(.dina(n11978), .dinb(n10844), .dout(n19024));
  jor  g18853(.dina(n19024), .dinb(n19023), .dout(n19025));
  jor  g18854(.dina(n19025), .dinb(n19022), .dout(n19026));
  jor  g18855(.dina(n19026), .dinb(n19021), .dout(n19027));
  jxor g18856(.dina(n19027), .dinb(n6600), .dout(n19028));
  jxor g18857(.dina(n18736), .dinb(n18735), .dout(n19029));
  jnot g18858(.din(n19029), .dout(n19030));
  jxor g18859(.dina(n18731), .dinb(n18730), .dout(n19031));
  jnot g18860(.din(n19031), .dout(n19032));
  jxor g18861(.dina(n18726), .dinb(n18725), .dout(n19033));
  jnot g18862(.din(n19033), .dout(n19034));
  jor  g18863(.dina(n14221), .dinb(n10847), .dout(n19035));
  jor  g18864(.dina(n15045), .dinb(n11458), .dout(n19036));
  jor  g18865(.dina(n11984), .dinb(n11360), .dout(n19037));
  jor  g18866(.dina(n11987), .dinb(n10845), .dout(n19038));
  jand g18867(.dina(n19038), .dinb(n19037), .dout(n19039));
  jand g18868(.dina(n19039), .dinb(n19036), .dout(n19040));
  jand g18869(.dina(n19040), .dinb(n19035), .dout(n19041));
  jxor g18870(.dina(n19041), .dinb(\a[2] ), .dout(n19042));
  jor  g18871(.dina(n14248), .dinb(n10847), .dout(n19043));
  jor  g18872(.dina(n11984), .dinb(n11458), .dout(n19044));
  jor  g18873(.dina(n11987), .dinb(n11360), .dout(n19045));
  jor  g18874(.dina(n11991), .dinb(n10845), .dout(n19046));
  jand g18875(.dina(n19046), .dinb(n19045), .dout(n19047));
  jand g18876(.dina(n19047), .dinb(n19044), .dout(n19048));
  jand g18877(.dina(n19048), .dinb(n19043), .dout(n19049));
  jxor g18878(.dina(n19049), .dinb(\a[2] ), .dout(n19050));
  jor  g18879(.dina(n14271), .dinb(n10847), .dout(n19051));
  jor  g18880(.dina(n11987), .dinb(n11458), .dout(n19052));
  jor  g18881(.dina(n11991), .dinb(n11360), .dout(n19053));
  jor  g18882(.dina(n11995), .dinb(n10845), .dout(n19054));
  jand g18883(.dina(n19054), .dinb(n19053), .dout(n19055));
  jand g18884(.dina(n19055), .dinb(n19052), .dout(n19056));
  jand g18885(.dina(n19056), .dinb(n19051), .dout(n19057));
  jxor g18886(.dina(n19057), .dinb(\a[2] ), .dout(n19058));
  jxor g18887(.dina(n18714), .dinb(n18713), .dout(n19059));
  jnot g18888(.din(n19059), .dout(n19060));
  jor  g18889(.dina(n14353), .dinb(n10847), .dout(n19061));
  jor  g18890(.dina(n11995), .dinb(n11458), .dout(n19062));
  jor  g18891(.dina(n11997), .dinb(n11360), .dout(n19063));
  jor  g18892(.dina(n11999), .dinb(n10845), .dout(n19064));
  jand g18893(.dina(n19064), .dinb(n19063), .dout(n19065));
  jand g18894(.dina(n19065), .dinb(n19062), .dout(n19066));
  jand g18895(.dina(n19066), .dinb(n19061), .dout(n19067));
  jxor g18896(.dina(n19067), .dinb(\a[2] ), .dout(n19068));
  jor  g18897(.dina(n18691), .dinb(n64), .dout(n19069));
  jxor g18898(.dina(n19069), .dinb(n18699), .dout(n19070));
  jnot g18899(.din(n19070), .dout(n19071));
  jor  g18900(.dina(n14432), .dinb(n10847), .dout(n19072));
  jor  g18901(.dina(n11999), .dinb(n11458), .dout(n19073));
  jor  g18902(.dina(n12001), .dinb(n11360), .dout(n19074));
  jor  g18903(.dina(n12004), .dinb(n10845), .dout(n19075));
  jand g18904(.dina(n19075), .dinb(n19074), .dout(n19076));
  jand g18905(.dina(n19076), .dinb(n19073), .dout(n19077));
  jand g18906(.dina(n19077), .dinb(n19072), .dout(n19078));
  jxor g18907(.dina(n19078), .dinb(\a[2] ), .dout(n19079));
  jand g18908(.dina(n14457), .dinb(n10846), .dout(n19080));
  jand g18909(.dina(n14393), .dinb(n11372), .dout(n19081));
  jand g18910(.dina(n12006), .dinb(n11359), .dout(n19082));
  jand g18911(.dina(n12008), .dinb(n10844), .dout(n19083));
  jor  g18912(.dina(n19083), .dinb(n19082), .dout(n19084));
  jor  g18913(.dina(n19084), .dinb(n19081), .dout(n19085));
  jor  g18914(.dina(n19085), .dinb(n19080), .dout(n19086));
  jor  g18915(.dina(n19086), .dinb(n18689), .dout(n19087));
  jor  g18916(.dina(n12006), .dinb(n10843), .dout(n19088));
  jand g18917(.dina(n19088), .dinb(\a[0] ), .dout(n19089));
  jnot g18918(.din(n10842), .dout(n19090));
  jand g18919(.dina(n12008), .dinb(n19090), .dout(n19091));
  jor  g18920(.dina(n19091), .dinb(n19089), .dout(n19092));
  jor  g18921(.dina(n14497), .dinb(n10847), .dout(n19093));
  jor  g18922(.dina(n19093), .dinb(n14537), .dout(n19094));
  jand g18923(.dina(n19094), .dinb(n19092), .dout(n19095));
  jor  g18924(.dina(n19095), .dinb(n12010), .dout(n19096));
  jand g18925(.dina(n19096), .dinb(\a[2] ), .dout(n19097));
  jand g18926(.dina(n19097), .dinb(n19087), .dout(n19098));
  jor  g18927(.dina(n15144), .dinb(n10847), .dout(n19099));
  jor  g18928(.dina(n12001), .dinb(n11458), .dout(n19100));
  jnot g18929(.din(n19084), .dout(n19101));
  jand g18930(.dina(n19101), .dinb(n19100), .dout(n19102));
  jand g18931(.dina(n19102), .dinb(n19099), .dout(n19103));
  jand g18932(.dina(n19103), .dinb(n6600), .dout(n19104));
  jand g18933(.dina(n19086), .dinb(n18689), .dout(n19105));
  jor  g18934(.dina(n19105), .dinb(n19104), .dout(n19106));
  jor  g18935(.dina(n19106), .dinb(n19098), .dout(n19107));
  jor  g18936(.dina(n19107), .dinb(n19079), .dout(n19108));
  jand g18937(.dina(n19107), .dinb(n19079), .dout(n19109));
  jand g18938(.dina(n18688), .dinb(\a[5] ), .dout(n19110));
  jxor g18939(.dina(n19110), .dinb(n18686), .dout(n19111));
  jnot g18940(.din(n19111), .dout(n19112));
  jor  g18941(.dina(n19112), .dinb(n19109), .dout(n19113));
  jand g18942(.dina(n19113), .dinb(n19108), .dout(n19114));
  jor  g18943(.dina(n19114), .dinb(n19071), .dout(n19115));
  jand g18944(.dina(n19114), .dinb(n19071), .dout(n19116));
  jor  g18945(.dina(n14390), .dinb(n10847), .dout(n19117));
  jor  g18946(.dina(n11997), .dinb(n11458), .dout(n19118));
  jor  g18947(.dina(n11999), .dinb(n11360), .dout(n19119));
  jor  g18948(.dina(n12001), .dinb(n10845), .dout(n19120));
  jand g18949(.dina(n19120), .dinb(n19119), .dout(n19121));
  jand g18950(.dina(n19121), .dinb(n19118), .dout(n19122));
  jand g18951(.dina(n19122), .dinb(n19117), .dout(n19123));
  jxor g18952(.dina(n19123), .dinb(\a[2] ), .dout(n19124));
  jor  g18953(.dina(n19124), .dinb(n19116), .dout(n19125));
  jand g18954(.dina(n19125), .dinb(n19115), .dout(n19126));
  jor  g18955(.dina(n19126), .dinb(n19068), .dout(n19127));
  jand g18956(.dina(n19126), .dinb(n19068), .dout(n19128));
  jxor g18957(.dina(n18711), .dinb(n18710), .dout(n19129));
  jnot g18958(.din(n19129), .dout(n19130));
  jor  g18959(.dina(n19130), .dinb(n19128), .dout(n19131));
  jand g18960(.dina(n19131), .dinb(n19127), .dout(n19132));
  jor  g18961(.dina(n19132), .dinb(n19060), .dout(n19133));
  jand g18962(.dina(n19132), .dinb(n19060), .dout(n19134));
  jor  g18963(.dina(n14301), .dinb(n10847), .dout(n19135));
  jor  g18964(.dina(n11991), .dinb(n11458), .dout(n19136));
  jor  g18965(.dina(n11995), .dinb(n11360), .dout(n19137));
  jor  g18966(.dina(n11997), .dinb(n10845), .dout(n19138));
  jand g18967(.dina(n19138), .dinb(n19137), .dout(n19139));
  jand g18968(.dina(n19139), .dinb(n19136), .dout(n19140));
  jand g18969(.dina(n19140), .dinb(n19135), .dout(n19141));
  jxor g18970(.dina(n19141), .dinb(\a[2] ), .dout(n19142));
  jor  g18971(.dina(n19142), .dinb(n19134), .dout(n19143));
  jand g18972(.dina(n19143), .dinb(n19133), .dout(n19144));
  jor  g18973(.dina(n19144), .dinb(n19058), .dout(n19145));
  jand g18974(.dina(n19144), .dinb(n19058), .dout(n19146));
  jxor g18975(.dina(n18717), .dinb(n18716), .dout(n19147));
  jnot g18976(.din(n19147), .dout(n19148));
  jor  g18977(.dina(n19148), .dinb(n19146), .dout(n19149));
  jand g18978(.dina(n19149), .dinb(n19145), .dout(n19150));
  jor  g18979(.dina(n19150), .dinb(n19050), .dout(n19151));
  jand g18980(.dina(n19150), .dinb(n19050), .dout(n19152));
  jxor g18981(.dina(n18720), .dinb(n18719), .dout(n19153));
  jnot g18982(.din(n19153), .dout(n19154));
  jor  g18983(.dina(n19154), .dinb(n19152), .dout(n19155));
  jand g18984(.dina(n19155), .dinb(n19151), .dout(n19156));
  jor  g18985(.dina(n19156), .dinb(n19042), .dout(n19157));
  jand g18986(.dina(n19156), .dinb(n19042), .dout(n19158));
  jxor g18987(.dina(n18723), .dinb(n18722), .dout(n19159));
  jnot g18988(.din(n19159), .dout(n19160));
  jor  g18989(.dina(n19160), .dinb(n19158), .dout(n19161));
  jand g18990(.dina(n19161), .dinb(n19157), .dout(n19162));
  jor  g18991(.dina(n19162), .dinb(n19034), .dout(n19163));
  jand g18992(.dina(n19162), .dinb(n19034), .dout(n19164));
  jand g18993(.dina(n13899), .dinb(n10846), .dout(n19165));
  jand g18994(.dina(n11980), .dinb(n11372), .dout(n19166));
  jand g18995(.dina(n11982), .dinb(n11359), .dout(n19167));
  jand g18996(.dina(n11985), .dinb(n10844), .dout(n19168));
  jor  g18997(.dina(n19168), .dinb(n19167), .dout(n19169));
  jor  g18998(.dina(n19169), .dinb(n19166), .dout(n19170));
  jor  g18999(.dina(n19170), .dinb(n19165), .dout(n19171));
  jxor g19000(.dina(n19171), .dinb(\a[2] ), .dout(n19172));
  jnot g19001(.din(n19172), .dout(n19173));
  jor  g19002(.dina(n19173), .dinb(n19164), .dout(n19174));
  jand g19003(.dina(n19174), .dinb(n19163), .dout(n19175));
  jor  g19004(.dina(n19175), .dinb(n19032), .dout(n19176));
  jand g19005(.dina(n19175), .dinb(n19032), .dout(n19177));
  jand g19006(.dina(n14194), .dinb(n10846), .dout(n19178));
  jand g19007(.dina(n11978), .dinb(n11372), .dout(n19179));
  jand g19008(.dina(n11980), .dinb(n11359), .dout(n19180));
  jand g19009(.dina(n11982), .dinb(n10844), .dout(n19181));
  jor  g19010(.dina(n19181), .dinb(n19180), .dout(n19182));
  jor  g19011(.dina(n19182), .dinb(n19179), .dout(n19183));
  jor  g19012(.dina(n19183), .dinb(n19178), .dout(n19184));
  jxor g19013(.dina(n19184), .dinb(\a[2] ), .dout(n19185));
  jnot g19014(.din(n19185), .dout(n19186));
  jor  g19015(.dina(n19186), .dinb(n19177), .dout(n19187));
  jand g19016(.dina(n19187), .dinb(n19176), .dout(n19188));
  jor  g19017(.dina(n19188), .dinb(n19030), .dout(n19189));
  jand g19018(.dina(n19188), .dinb(n19030), .dout(n19190));
  jand g19019(.dina(n14184), .dinb(n10846), .dout(n19191));
  jand g19020(.dina(n11976), .dinb(n11372), .dout(n19192));
  jand g19021(.dina(n11978), .dinb(n11359), .dout(n19193));
  jand g19022(.dina(n11980), .dinb(n10844), .dout(n19194));
  jor  g19023(.dina(n19194), .dinb(n19193), .dout(n19195));
  jor  g19024(.dina(n19195), .dinb(n19192), .dout(n19196));
  jor  g19025(.dina(n19196), .dinb(n19191), .dout(n19197));
  jxor g19026(.dina(n19197), .dinb(\a[2] ), .dout(n19198));
  jnot g19027(.din(n19198), .dout(n19199));
  jor  g19028(.dina(n19199), .dinb(n19190), .dout(n19200));
  jand g19029(.dina(n19200), .dinb(n19189), .dout(n19201));
  jor  g19030(.dina(n19201), .dinb(n19028), .dout(n19202));
  jand g19031(.dina(n19201), .dinb(n19028), .dout(n19203));
  jxor g19032(.dina(n18741), .dinb(n18740), .dout(n19204));
  jnot g19033(.din(n19204), .dout(n19205));
  jor  g19034(.dina(n19205), .dinb(n19203), .dout(n19206));
  jand g19035(.dina(n19206), .dinb(n19202), .dout(n19207));
  jor  g19036(.dina(n19207), .dinb(n19020), .dout(n19208));
  jand g19037(.dina(n19207), .dinb(n19020), .dout(n19209));
  jxor g19038(.dina(n18744), .dinb(n18743), .dout(n19210));
  jnot g19039(.din(n19210), .dout(n19211));
  jor  g19040(.dina(n19211), .dinb(n19209), .dout(n19212));
  jand g19041(.dina(n19212), .dinb(n19208), .dout(n19213));
  jor  g19042(.dina(n19213), .dinb(n19012), .dout(n19214));
  jand g19043(.dina(n19213), .dinb(n19012), .dout(n19215));
  jxor g19044(.dina(n18747), .dinb(n18746), .dout(n19216));
  jnot g19045(.din(n19216), .dout(n19217));
  jor  g19046(.dina(n19217), .dinb(n19215), .dout(n19218));
  jand g19047(.dina(n19218), .dinb(n19214), .dout(n19219));
  jor  g19048(.dina(n19219), .dinb(n19004), .dout(n19220));
  jand g19049(.dina(n19219), .dinb(n19004), .dout(n19221));
  jand g19050(.dina(n13682), .dinb(n10846), .dout(n19222));
  jand g19051(.dina(n11968), .dinb(n11372), .dout(n19223));
  jand g19052(.dina(n11970), .dinb(n11359), .dout(n19224));
  jand g19053(.dina(n11972), .dinb(n10844), .dout(n19225));
  jor  g19054(.dina(n19225), .dinb(n19224), .dout(n19226));
  jor  g19055(.dina(n19226), .dinb(n19223), .dout(n19227));
  jor  g19056(.dina(n19227), .dinb(n19222), .dout(n19228));
  jxor g19057(.dina(n19228), .dinb(\a[2] ), .dout(n19229));
  jnot g19058(.din(n19229), .dout(n19230));
  jor  g19059(.dina(n19230), .dinb(n19221), .dout(n19231));
  jand g19060(.dina(n19231), .dinb(n19220), .dout(n19232));
  jor  g19061(.dina(n19232), .dinb(n19002), .dout(n19233));
  jand g19062(.dina(n19232), .dinb(n19002), .dout(n19234));
  jand g19063(.dina(n13268), .dinb(n10846), .dout(n19235));
  jand g19064(.dina(n11966), .dinb(n11372), .dout(n19236));
  jand g19065(.dina(n11968), .dinb(n11359), .dout(n19237));
  jand g19066(.dina(n11970), .dinb(n10844), .dout(n19238));
  jor  g19067(.dina(n19238), .dinb(n19237), .dout(n19239));
  jor  g19068(.dina(n19239), .dinb(n19236), .dout(n19240));
  jor  g19069(.dina(n19240), .dinb(n19235), .dout(n19241));
  jxor g19070(.dina(n19241), .dinb(\a[2] ), .dout(n19242));
  jnot g19071(.din(n19242), .dout(n19243));
  jor  g19072(.dina(n19243), .dinb(n19234), .dout(n19244));
  jand g19073(.dina(n19244), .dinb(n19233), .dout(n19245));
  jor  g19074(.dina(n19245), .dinb(n19000), .dout(n19246));
  jand g19075(.dina(n19245), .dinb(n19000), .dout(n19247));
  jand g19076(.dina(n13470), .dinb(n10846), .dout(n19248));
  jand g19077(.dina(n11964), .dinb(n11372), .dout(n19249));
  jand g19078(.dina(n11966), .dinb(n11359), .dout(n19250));
  jand g19079(.dina(n11968), .dinb(n10844), .dout(n19251));
  jor  g19080(.dina(n19251), .dinb(n19250), .dout(n19252));
  jor  g19081(.dina(n19252), .dinb(n19249), .dout(n19253));
  jor  g19082(.dina(n19253), .dinb(n19248), .dout(n19254));
  jxor g19083(.dina(n19254), .dinb(\a[2] ), .dout(n19255));
  jnot g19084(.din(n19255), .dout(n19256));
  jor  g19085(.dina(n19256), .dinb(n19247), .dout(n19257));
  jand g19086(.dina(n19257), .dinb(n19246), .dout(n19258));
  jor  g19087(.dina(n19258), .dinb(n18998), .dout(n19259));
  jand g19088(.dina(n19258), .dinb(n18998), .dout(n19260));
  jxor g19089(.dina(n18765), .dinb(n18764), .dout(n19261));
  jnot g19090(.din(n19261), .dout(n19262));
  jor  g19091(.dina(n19262), .dinb(n19260), .dout(n19263));
  jand g19092(.dina(n19263), .dinb(n19259), .dout(n19264));
  jor  g19093(.dina(n19264), .dinb(n18990), .dout(n19265));
  jand g19094(.dina(n19264), .dinb(n18990), .dout(n19266));
  jxor g19095(.dina(n18768), .dinb(n18767), .dout(n19267));
  jnot g19096(.din(n19267), .dout(n19268));
  jor  g19097(.dina(n19268), .dinb(n19266), .dout(n19269));
  jand g19098(.dina(n19269), .dinb(n19265), .dout(n19270));
  jor  g19099(.dina(n19270), .dinb(n18982), .dout(n19271));
  jand g19100(.dina(n19270), .dinb(n18982), .dout(n19272));
  jxor g19101(.dina(n18771), .dinb(n18770), .dout(n19273));
  jnot g19102(.din(n19273), .dout(n19274));
  jor  g19103(.dina(n19274), .dinb(n19272), .dout(n19275));
  jand g19104(.dina(n19275), .dinb(n19271), .dout(n19276));
  jor  g19105(.dina(n19276), .dinb(n18974), .dout(n19277));
  jand g19106(.dina(n19276), .dinb(n18974), .dout(n19278));
  jand g19107(.dina(n12639), .dinb(n10846), .dout(n19279));
  jand g19108(.dina(n11956), .dinb(n11372), .dout(n19280));
  jand g19109(.dina(n11958), .dinb(n11359), .dout(n19281));
  jand g19110(.dina(n11960), .dinb(n10844), .dout(n19282));
  jor  g19111(.dina(n19282), .dinb(n19281), .dout(n19283));
  jor  g19112(.dina(n19283), .dinb(n19280), .dout(n19284));
  jor  g19113(.dina(n19284), .dinb(n19279), .dout(n19285));
  jxor g19114(.dina(n19285), .dinb(\a[2] ), .dout(n19286));
  jnot g19115(.din(n19286), .dout(n19287));
  jor  g19116(.dina(n19287), .dinb(n19278), .dout(n19288));
  jand g19117(.dina(n19288), .dinb(n19277), .dout(n19289));
  jor  g19118(.dina(n19289), .dinb(n18972), .dout(n19290));
  jand g19119(.dina(n19289), .dinb(n18972), .dout(n19291));
  jand g19120(.dina(n12472), .dinb(n10846), .dout(n19292));
  jand g19121(.dina(n11954), .dinb(n11372), .dout(n19293));
  jand g19122(.dina(n11956), .dinb(n11359), .dout(n19294));
  jand g19123(.dina(n11958), .dinb(n10844), .dout(n19295));
  jor  g19124(.dina(n19295), .dinb(n19294), .dout(n19296));
  jor  g19125(.dina(n19296), .dinb(n19293), .dout(n19297));
  jor  g19126(.dina(n19297), .dinb(n19292), .dout(n19298));
  jxor g19127(.dina(n19298), .dinb(\a[2] ), .dout(n19299));
  jnot g19128(.din(n19299), .dout(n19300));
  jor  g19129(.dina(n19300), .dinb(n19291), .dout(n19301));
  jand g19130(.dina(n19301), .dinb(n19290), .dout(n19302));
  jor  g19131(.dina(n19302), .dinb(n18970), .dout(n19303));
  jand g19132(.dina(n19302), .dinb(n18970), .dout(n19304));
  jand g19133(.dina(n12510), .dinb(n10846), .dout(n19305));
  jand g19134(.dina(n11952), .dinb(n11372), .dout(n19306));
  jand g19135(.dina(n11954), .dinb(n11359), .dout(n19307));
  jand g19136(.dina(n11956), .dinb(n10844), .dout(n19308));
  jor  g19137(.dina(n19308), .dinb(n19307), .dout(n19309));
  jor  g19138(.dina(n19309), .dinb(n19306), .dout(n19310));
  jor  g19139(.dina(n19310), .dinb(n19305), .dout(n19311));
  jxor g19140(.dina(n19311), .dinb(\a[2] ), .dout(n19312));
  jnot g19141(.din(n19312), .dout(n19313));
  jor  g19142(.dina(n19313), .dinb(n19304), .dout(n19314));
  jand g19143(.dina(n19314), .dinb(n19303), .dout(n19315));
  jor  g19144(.dina(n19315), .dinb(n18968), .dout(n19316));
  jand g19145(.dina(n19315), .dinb(n18968), .dout(n19317));
  jxor g19146(.dina(n18789), .dinb(n18788), .dout(n19318));
  jnot g19147(.din(n19318), .dout(n19319));
  jor  g19148(.dina(n19319), .dinb(n19317), .dout(n19320));
  jand g19149(.dina(n19320), .dinb(n19316), .dout(n19321));
  jor  g19150(.dina(n19321), .dinb(n18960), .dout(n19322));
  jand g19151(.dina(n19321), .dinb(n18960), .dout(n19323));
  jxor g19152(.dina(n18792), .dinb(n18791), .dout(n19324));
  jnot g19153(.din(n19324), .dout(n19325));
  jor  g19154(.dina(n19325), .dinb(n19323), .dout(n19326));
  jand g19155(.dina(n19326), .dinb(n19322), .dout(n19327));
  jor  g19156(.dina(n19327), .dinb(n18952), .dout(n19328));
  jand g19157(.dina(n19327), .dinb(n18952), .dout(n19329));
  jxor g19158(.dina(n18795), .dinb(n18794), .dout(n19330));
  jnot g19159(.din(n19330), .dout(n19331));
  jor  g19160(.dina(n19331), .dinb(n19329), .dout(n19332));
  jand g19161(.dina(n19332), .dinb(n19328), .dout(n19333));
  jor  g19162(.dina(n19333), .dinb(n18944), .dout(n19334));
  jand g19163(.dina(n19333), .dinb(n18944), .dout(n19335));
  jand g19164(.dina(n12189), .dinb(n10846), .dout(n19336));
  jand g19165(.dina(n11944), .dinb(n11372), .dout(n19337));
  jand g19166(.dina(n11946), .dinb(n11359), .dout(n19338));
  jand g19167(.dina(n11948), .dinb(n10844), .dout(n19339));
  jor  g19168(.dina(n19339), .dinb(n19338), .dout(n19340));
  jor  g19169(.dina(n19340), .dinb(n19337), .dout(n19341));
  jor  g19170(.dina(n19341), .dinb(n19336), .dout(n19342));
  jxor g19171(.dina(n19342), .dinb(\a[2] ), .dout(n19343));
  jnot g19172(.din(n19343), .dout(n19344));
  jor  g19173(.dina(n19344), .dinb(n19335), .dout(n19345));
  jand g19174(.dina(n19345), .dinb(n19334), .dout(n19346));
  jor  g19175(.dina(n19346), .dinb(n18942), .dout(n19347));
  jand g19176(.dina(n19346), .dinb(n18942), .dout(n19348));
  jand g19177(.dina(n12751), .dinb(n10846), .dout(n19349));
  jand g19178(.dina(n11942), .dinb(n11372), .dout(n19350));
  jand g19179(.dina(n11944), .dinb(n11359), .dout(n19351));
  jand g19180(.dina(n11946), .dinb(n10844), .dout(n19352));
  jor  g19181(.dina(n19352), .dinb(n19351), .dout(n19353));
  jor  g19182(.dina(n19353), .dinb(n19350), .dout(n19354));
  jor  g19183(.dina(n19354), .dinb(n19349), .dout(n19355));
  jxor g19184(.dina(n19355), .dinb(\a[2] ), .dout(n19356));
  jnot g19185(.din(n19356), .dout(n19357));
  jor  g19186(.dina(n19357), .dinb(n19348), .dout(n19358));
  jand g19187(.dina(n19358), .dinb(n19347), .dout(n19359));
  jor  g19188(.dina(n19359), .dinb(n18940), .dout(n19360));
  jand g19189(.dina(n19360), .dinb(n18938), .dout(n19361));
  jxor g19190(.dina(n18926), .dinb(n18918), .dout(n19362));
  jnot g19191(.din(n19362), .dout(n19363));
  jor  g19192(.dina(n19363), .dinb(n19361), .dout(n19364));
  jand g19193(.dina(n19364), .dinb(n18927), .dout(n19365));
  jxor g19194(.dina(n18915), .dinb(n18907), .dout(n19366));
  jnot g19195(.din(n19366), .dout(n19367));
  jor  g19196(.dina(n19367), .dinb(n19365), .dout(n19368));
  jand g19197(.dina(n19368), .dinb(n18916), .dout(n19369));
  jxor g19198(.dina(n18904), .dinb(n18896), .dout(n19370));
  jnot g19199(.din(n19370), .dout(n19371));
  jor  g19200(.dina(n19371), .dinb(n19369), .dout(n19372));
  jand g19201(.dina(n19372), .dinb(n18905), .dout(n19373));
  jxor g19202(.dina(n18893), .dinb(n18885), .dout(n19374));
  jnot g19203(.din(n19374), .dout(n19375));
  jor  g19204(.dina(n19375), .dinb(n19373), .dout(n19376));
  jand g19205(.dina(n19376), .dinb(n18894), .dout(n19377));
  jxor g19206(.dina(n18882), .dinb(n18874), .dout(n19378));
  jnot g19207(.din(n19378), .dout(n19379));
  jor  g19208(.dina(n19379), .dinb(n19377), .dout(n19380));
  jand g19209(.dina(n19380), .dinb(n18883), .dout(n19381));
  jxor g19210(.dina(n18871), .dinb(n18863), .dout(n19382));
  jnot g19211(.din(n19382), .dout(n19383));
  jor  g19212(.dina(n19383), .dinb(n19381), .dout(n19384));
  jand g19213(.dina(n19384), .dinb(n18872), .dout(n19385));
  jxor g19214(.dina(n18860), .dinb(n18851), .dout(n19386));
  jor  g19215(.dina(n19386), .dinb(n19385), .dout(n19387));
  jand g19216(.dina(n19387), .dinb(n18861), .dout(n19388));
  jxor g19217(.dina(n18849), .dinb(n18841), .dout(n19389));
  jnot g19218(.din(n19389), .dout(n19390));
  jor  g19219(.dina(n19390), .dinb(n19388), .dout(n19391));
  jand g19220(.dina(n19391), .dinb(n18850), .dout(n19392));
  jor  g19221(.dina(n19392), .dinb(n18839), .dout(n19393));
  jand g19222(.dina(n19393), .dinb(n18837), .dout(n19394));
  jor  g19223(.dina(n19394), .dinb(n18316), .dout(n19395));
  jand g19224(.dina(n19395), .dinb(n18314), .dout(n19396));
  jor  g19225(.dina(n19396), .dinb(n18290), .dout(n19397));
  jand g19226(.dina(n19397), .dinb(n18288), .dout(n19398));
  jor  g19227(.dina(n19398), .dinb(n17765), .dout(n19399));
  jand g19228(.dina(n19399), .dinb(n17763), .dout(n19400));
  jnot g19229(.din(n19400), .dout(n19401));
  jxor g19230(.dina(n17285), .dinb(n17284), .dout(n19402));
  jand g19231(.dina(n19402), .dinb(n19401), .dout(n19403));
  jor  g19232(.dina(n19403), .dinb(n17286), .dout(n19404));
  jxor g19233(.dina(n16822), .dinb(n16821), .dout(n19405));
  jand g19234(.dina(n19405), .dinb(n19404), .dout(n19406));
  jor  g19235(.dina(n19406), .dinb(n16823), .dout(n19407));
  jand g19236(.dina(n19407), .dinb(n16407), .dout(n19408));
  jor  g19237(.dina(n19408), .dinb(n16406), .dout(n19409));
  jxor g19238(.dina(n15997), .dinb(n15996), .dout(n19410));
  jand g19239(.dina(n19410), .dinb(n19409), .dout(n19411));
  jor  g19240(.dina(n19411), .dinb(n15998), .dout(n19412));
  jxor g19241(.dina(n15640), .dinb(n15639), .dout(n19413));
  jand g19242(.dina(n19413), .dinb(n19412), .dout(n19414));
  jor  g19243(.dina(n19414), .dinb(n15641), .dout(n19415));
  jand g19244(.dina(n19415), .dinb(n15295), .dout(n19416));
  jor  g19245(.dina(n19416), .dinb(n15294), .dout(n19417));
  jxor g19246(.dina(n14987), .dinb(n14986), .dout(n19418));
  jand g19247(.dina(n19418), .dinb(n19417), .dout(n19419));
  jor  g19248(.dina(n19419), .dinb(n14988), .dout(n19420));
  jxor g19249(.dina(n14851), .dinb(n14850), .dout(n19421));
  jand g19250(.dina(n19421), .dinb(n19420), .dout(n19422));
  jor  g19251(.dina(n19422), .dinb(n14852), .dout(n19423));
  jand g19252(.dina(n19423), .dinb(n14717), .dout(n19424));
  jor  g19253(.dina(n19424), .dinb(n14716), .dout(n19425));
  jxor g19254(.dina(n14159), .dinb(n14158), .dout(n19426));
  jand g19255(.dina(n19426), .dinb(n19425), .dout(n19427));
  jor  g19256(.dina(n19427), .dinb(n14160), .dout(n19428));
  jxor g19257(.dina(n14039), .dinb(n14038), .dout(n19429));
  jand g19258(.dina(n19429), .dinb(n19428), .dout(n19430));
  jor  g19259(.dina(n19430), .dinb(n14040), .dout(n19431));
  jand g19260(.dina(n19431), .dinb(n13782), .dout(n19432));
  jor  g19261(.dina(n19432), .dinb(n13781), .dout(n19433));
  jxor g19262(.dina(n13571), .dinb(n13570), .dout(n19434));
  jand g19263(.dina(n19434), .dinb(n19433), .dout(n19435));
  jor  g19264(.dina(n19435), .dinb(n13572), .dout(n19436));
  jxor g19265(.dina(n13456), .dinb(n13455), .dout(n19437));
  jand g19266(.dina(n19437), .dinb(n19436), .dout(n19438));
  jor  g19267(.dina(n19438), .dinb(n13457), .dout(n19439));
  jand g19268(.dina(n19439), .dinb(n13368), .dout(n19440));
  jor  g19269(.dina(n19440), .dinb(n13367), .dout(n19441));
  jxor g19270(.dina(n13032), .dinb(n12932), .dout(n19442));
  jand g19271(.dina(n19442), .dinb(n19441), .dout(n19443));
  jor  g19272(.dina(n19443), .dinb(n13033), .dout(n19444));
  jor  g19273(.dina(n13030), .dinb(n13018), .dout(n19445));
  jand g19274(.dina(n13031), .dinb(n13014), .dout(n19446));
  jnot g19275(.din(n19446), .dout(n19447));
  jand g19276(.dina(n19447), .dinb(n19445), .dout(n19448));
  jnot g19277(.din(n19448), .dout(n19449));
  jor  g19278(.dina(n5424), .dinb(n5500), .dout(n19452));
  jand g19279(.dina(n12815), .dinb(n5363), .dout(n19454));
  jor  g19280(.dina(n19454), .dinb(n19452), .dout(n19455));
  jor  g19281(.dina(n19455), .dinb(n5365), .dout(n19456));
  jxor g19282(.dina(n19456), .dinb(n72), .dout(n19457));
  jnot g19283(.din(n19457), .dout(n19458));
  jand g19284(.dina(n13012), .dinb(n12947), .dout(n19459));
  jand g19285(.dina(n13013), .dinb(n12937), .dout(n19460));
  jor  g19286(.dina(n19460), .dinb(n19459), .dout(n19461));
  jand g19287(.dina(n12797), .dinb(n75), .dout(n19462));
  jand g19288(.dina(n12795), .dinb(n4933), .dout(n19463));
  jand g19289(.dina(n12782), .dinb(n4918), .dout(n19464));
  jand g19290(.dina(n12783), .dinb(n4745), .dout(n19465));
  jor  g19291(.dina(n19465), .dinb(n19464), .dout(n19466));
  jor  g19292(.dina(n19466), .dinb(n19463), .dout(n19467));
  jor  g19293(.dina(n19467), .dinb(n19462), .dout(n19468));
  jxor g19294(.dina(n19468), .dinb(n68), .dout(n19469));
  jnot g19295(.din(n19469), .dout(n19470));
  jand g19296(.dina(n13001), .dinb(n12952), .dout(n19471));
  jnot g19297(.din(n19471), .dout(n19472));
  jor  g19298(.dina(n13011), .dinb(n13003), .dout(n19473));
  jand g19299(.dina(n19473), .dinb(n19472), .dout(n19474));
  jnot g19300(.din(n12431), .dout(n19475));
  jor  g19301(.dina(n12990), .dinb(n12738), .dout(n19476));
  jand g19302(.dina(n12991), .dinb(n12961), .dout(n19477));
  jnot g19303(.din(n19477), .dout(n19478));
  jand g19304(.dina(n19478), .dinb(n19476), .dout(n19479));
  jxor g19305(.dina(n19479), .dinb(n19475), .dout(n19480));
  jand g19306(.dina(n12751), .dinb(n732), .dout(n19481));
  jand g19307(.dina(n11942), .dinb(n3855), .dout(n19482));
  jand g19308(.dina(n11946), .dinb(n3851), .dout(n19483));
  jand g19309(.dina(n11944), .dinb(n3858), .dout(n19484));
  jor  g19310(.dina(n19484), .dinb(n19483), .dout(n19485));
  jor  g19311(.dina(n19485), .dinb(n19482), .dout(n19486));
  jor  g19312(.dina(n19486), .dinb(n19481), .dout(n19487));
  jxor g19313(.dina(n19487), .dinb(n19480), .dout(n19488));
  jor  g19314(.dina(n12992), .dinb(n12957), .dout(n19489));
  jand g19315(.dina(n12992), .dinb(n12957), .dout(n19490));
  jor  g19316(.dina(n13000), .dinb(n19490), .dout(n19491));
  jand g19317(.dina(n19491), .dinb(n19489), .dout(n19492));
  jxor g19318(.dina(n19492), .dinb(n19488), .dout(n19493));
  jnot g19319(.din(n19493), .dout(n19494));
  jand g19320(.dina(n12768), .dinb(n4449), .dout(n19495));
  jand g19321(.dina(n12766), .dinb(n4453), .dout(n19496));
  jand g19322(.dina(n12177), .dinb(n4457), .dout(n19497));
  jand g19323(.dina(n11941), .dinb(n4461), .dout(n19498));
  jor  g19324(.dina(n19498), .dinb(n19497), .dout(n19499));
  jor  g19325(.dina(n19499), .dinb(n19496), .dout(n19500));
  jor  g19326(.dina(n19500), .dinb(n19495), .dout(n19501));
  jxor g19327(.dina(n19501), .dinb(n88), .dout(n19502));
  jxor g19328(.dina(n19502), .dinb(n19494), .dout(n19503));
  jnot g19329(.din(n19503), .dout(n19504));
  jxor g19330(.dina(n19504), .dinb(n19474), .dout(n19505));
  jxor g19331(.dina(n19505), .dinb(n19470), .dout(n19506));
  jxor g19332(.dina(n19506), .dinb(n19461), .dout(n19507));
  jxor g19333(.dina(n19507), .dinb(n19458), .dout(n19508));
  jxor g19334(.dina(n19508), .dinb(n19449), .dout(n19509));
  jxor g19335(.dina(n19509), .dinb(n19444), .dout(n19510));
  jxor g19336(.dina(n19442), .dinb(n19441), .dout(n19511));
  jand g19337(.dina(n19511), .dinb(n19510), .dout(n19512));
  jxor g19338(.dina(n19439), .dinb(n13368), .dout(n19513));
  jand g19339(.dina(n19513), .dinb(n19511), .dout(n19514));
  jxor g19340(.dina(n19437), .dinb(n19436), .dout(n19515));
  jand g19341(.dina(n19515), .dinb(n19513), .dout(n19516));
  jxor g19342(.dina(n19434), .dinb(n19433), .dout(n19517));
  jand g19343(.dina(n19517), .dinb(n19515), .dout(n19518));
  jxor g19344(.dina(n19431), .dinb(n13782), .dout(n19519));
  jand g19345(.dina(n19519), .dinb(n19517), .dout(n19520));
  jxor g19346(.dina(n19429), .dinb(n19428), .dout(n19521));
  jand g19347(.dina(n19521), .dinb(n19519), .dout(n19522));
  jxor g19348(.dina(n19426), .dinb(n19425), .dout(n19523));
  jand g19349(.dina(n19523), .dinb(n19521), .dout(n19524));
  jxor g19350(.dina(n19423), .dinb(n14717), .dout(n19525));
  jand g19351(.dina(n19525), .dinb(n19523), .dout(n19526));
  jxor g19352(.dina(n19421), .dinb(n19420), .dout(n19527));
  jand g19353(.dina(n19527), .dinb(n19525), .dout(n19528));
  jxor g19354(.dina(n19418), .dinb(n19417), .dout(n19529));
  jand g19355(.dina(n19529), .dinb(n19527), .dout(n19530));
  jxor g19356(.dina(n19415), .dinb(n15295), .dout(n19531));
  jand g19357(.dina(n19531), .dinb(n19529), .dout(n19532));
  jxor g19358(.dina(n19413), .dinb(n19412), .dout(n19533));
  jand g19359(.dina(n19533), .dinb(n19531), .dout(n19534));
  jxor g19360(.dina(n19410), .dinb(n19409), .dout(n19535));
  jand g19361(.dina(n19535), .dinb(n19533), .dout(n19536));
  jxor g19362(.dina(n19407), .dinb(n16407), .dout(n19537));
  jand g19363(.dina(n19537), .dinb(n19535), .dout(n19538));
  jxor g19364(.dina(n19405), .dinb(n19404), .dout(n19539));
  jand g19365(.dina(n19539), .dinb(n19537), .dout(n19540));
  jxor g19366(.dina(n19402), .dinb(n19401), .dout(n19541));
  jand g19367(.dina(n19541), .dinb(n19539), .dout(n19542));
  jxor g19368(.dina(n19398), .dinb(n17765), .dout(n19543));
  jand g19369(.dina(n19543), .dinb(n19541), .dout(n19544));
  jxor g19370(.dina(n19396), .dinb(n18290), .dout(n19545));
  jand g19371(.dina(n19545), .dinb(n19543), .dout(n19546));
  jxor g19372(.dina(n19394), .dinb(n18315), .dout(n19547));
  jnot g19373(.din(n19547), .dout(n19548));
  jand g19374(.dina(n19548), .dinb(n19545), .dout(n19549));
  jxor g19375(.dina(n19392), .dinb(n18838), .dout(n19550));
  jnot g19376(.din(n19550), .dout(n19551));
  jand g19377(.dina(n19551), .dinb(n19548), .dout(n19552));
  jxor g19378(.dina(n19389), .dinb(n19388), .dout(n19553));
  jnot g19379(.din(n19553), .dout(n19554));
  jand g19380(.dina(n19554), .dinb(n19551), .dout(n19555));
  jnot g19381(.din(n19555), .dout(n19556));
  jnot g19382(.din(n19386), .dout(n19557));
  jxor g19383(.dina(n19557), .dinb(n19385), .dout(n19558));
  jnot g19384(.din(n19558), .dout(n19559));
  jand g19385(.dina(n19559), .dinb(n19554), .dout(n19560));
  jnot g19386(.din(n19560), .dout(n19561));
  jxor g19387(.dina(n19382), .dinb(n19381), .dout(n19562));
  jor  g19388(.dina(n19562), .dinb(n19558), .dout(n19563));
  jxor g19389(.dina(n19378), .dinb(n19377), .dout(n19564));
  jor  g19390(.dina(n19564), .dinb(n19562), .dout(n19565));
  jxor g19391(.dina(n19374), .dinb(n19373), .dout(n19566));
  jor  g19392(.dina(n19566), .dinb(n19564), .dout(n19567));
  jxor g19393(.dina(n19370), .dinb(n19369), .dout(n19568));
  jor  g19394(.dina(n19568), .dinb(n19566), .dout(n19569));
  jxor g19395(.dina(n19366), .dinb(n19365), .dout(n19570));
  jor  g19396(.dina(n19570), .dinb(n19568), .dout(n19571));
  jxor g19397(.dina(n19367), .dinb(n19365), .dout(n19572));
  jxor g19398(.dina(n19572), .dinb(n19568), .dout(n19573));
  jxor g19399(.dina(n19363), .dinb(n19361), .dout(n19574));
  jnot g19400(.din(n19574), .dout(n19575));
  jxor g19401(.dina(n19359), .dinb(n18940), .dout(n19576));
  jnot g19402(.din(n19576), .dout(n19577));
  jand g19403(.dina(n19577), .dinb(n19570), .dout(n19578));
  jor  g19404(.dina(n19578), .dinb(n19575), .dout(n19579));
  jor  g19405(.dina(n19579), .dinb(n19573), .dout(n19580));
  jand g19406(.dina(n19580), .dinb(n19571), .dout(n19581));
  jxor g19407(.dina(n19568), .dinb(n19566), .dout(n19582));
  jnot g19408(.din(n19582), .dout(n19583));
  jor  g19409(.dina(n19583), .dinb(n19581), .dout(n19584));
  jand g19410(.dina(n19584), .dinb(n19569), .dout(n19585));
  jxor g19411(.dina(n19566), .dinb(n19564), .dout(n19586));
  jnot g19412(.din(n19586), .dout(n19587));
  jor  g19413(.dina(n19587), .dinb(n19585), .dout(n19588));
  jand g19414(.dina(n19588), .dinb(n19567), .dout(n19589));
  jxor g19415(.dina(n19564), .dinb(n19562), .dout(n19590));
  jnot g19416(.din(n19590), .dout(n19591));
  jor  g19417(.dina(n19591), .dinb(n19589), .dout(n19592));
  jand g19418(.dina(n19592), .dinb(n19565), .dout(n19593));
  jxor g19419(.dina(n19562), .dinb(n19558), .dout(n19594));
  jnot g19420(.din(n19594), .dout(n19595));
  jor  g19421(.dina(n19595), .dinb(n19593), .dout(n19596));
  jand g19422(.dina(n19596), .dinb(n19563), .dout(n19597));
  jxor g19423(.dina(n19558), .dinb(n19553), .dout(n19598));
  jnot g19424(.din(n19598), .dout(n19599));
  jor  g19425(.dina(n19599), .dinb(n19597), .dout(n19600));
  jand g19426(.dina(n19600), .dinb(n19561), .dout(n19601));
  jxor g19427(.dina(n19553), .dinb(n19550), .dout(n19602));
  jnot g19428(.din(n19602), .dout(n19603));
  jor  g19429(.dina(n19603), .dinb(n19601), .dout(n19604));
  jand g19430(.dina(n19604), .dinb(n19556), .dout(n19605));
  jnot g19431(.din(n19605), .dout(n19606));
  jxor g19432(.dina(n19550), .dinb(n19547), .dout(n19607));
  jand g19433(.dina(n19607), .dinb(n19606), .dout(n19608));
  jor  g19434(.dina(n19608), .dinb(n19552), .dout(n19609));
  jxor g19435(.dina(n19548), .dinb(n19545), .dout(n19610));
  jand g19436(.dina(n19610), .dinb(n19609), .dout(n19611));
  jor  g19437(.dina(n19611), .dinb(n19549), .dout(n19612));
  jxor g19438(.dina(n19545), .dinb(n19543), .dout(n19613));
  jand g19439(.dina(n19613), .dinb(n19612), .dout(n19614));
  jor  g19440(.dina(n19614), .dinb(n19546), .dout(n19615));
  jxor g19441(.dina(n19543), .dinb(n19541), .dout(n19616));
  jand g19442(.dina(n19616), .dinb(n19615), .dout(n19617));
  jor  g19443(.dina(n19617), .dinb(n19544), .dout(n19618));
  jxor g19444(.dina(n19541), .dinb(n19539), .dout(n19619));
  jand g19445(.dina(n19619), .dinb(n19618), .dout(n19620));
  jor  g19446(.dina(n19620), .dinb(n19542), .dout(n19621));
  jxor g19447(.dina(n19539), .dinb(n19537), .dout(n19622));
  jand g19448(.dina(n19622), .dinb(n19621), .dout(n19623));
  jor  g19449(.dina(n19623), .dinb(n19540), .dout(n19624));
  jxor g19450(.dina(n19537), .dinb(n19535), .dout(n19625));
  jand g19451(.dina(n19625), .dinb(n19624), .dout(n19626));
  jor  g19452(.dina(n19626), .dinb(n19538), .dout(n19627));
  jxor g19453(.dina(n19535), .dinb(n19533), .dout(n19628));
  jand g19454(.dina(n19628), .dinb(n19627), .dout(n19629));
  jor  g19455(.dina(n19629), .dinb(n19536), .dout(n19630));
  jxor g19456(.dina(n19533), .dinb(n19531), .dout(n19631));
  jand g19457(.dina(n19631), .dinb(n19630), .dout(n19632));
  jor  g19458(.dina(n19632), .dinb(n19534), .dout(n19633));
  jxor g19459(.dina(n19531), .dinb(n19529), .dout(n19634));
  jand g19460(.dina(n19634), .dinb(n19633), .dout(n19635));
  jor  g19461(.dina(n19635), .dinb(n19532), .dout(n19636));
  jxor g19462(.dina(n19529), .dinb(n19527), .dout(n19637));
  jand g19463(.dina(n19637), .dinb(n19636), .dout(n19638));
  jor  g19464(.dina(n19638), .dinb(n19530), .dout(n19639));
  jxor g19465(.dina(n19527), .dinb(n19525), .dout(n19640));
  jand g19466(.dina(n19640), .dinb(n19639), .dout(n19641));
  jor  g19467(.dina(n19641), .dinb(n19528), .dout(n19642));
  jxor g19468(.dina(n19525), .dinb(n19523), .dout(n19643));
  jand g19469(.dina(n19643), .dinb(n19642), .dout(n19644));
  jor  g19470(.dina(n19644), .dinb(n19526), .dout(n19645));
  jxor g19471(.dina(n19523), .dinb(n19521), .dout(n19646));
  jand g19472(.dina(n19646), .dinb(n19645), .dout(n19647));
  jor  g19473(.dina(n19647), .dinb(n19524), .dout(n19648));
  jxor g19474(.dina(n19521), .dinb(n19519), .dout(n19649));
  jand g19475(.dina(n19649), .dinb(n19648), .dout(n19650));
  jor  g19476(.dina(n19650), .dinb(n19522), .dout(n19651));
  jxor g19477(.dina(n19519), .dinb(n19517), .dout(n19652));
  jand g19478(.dina(n19652), .dinb(n19651), .dout(n19653));
  jor  g19479(.dina(n19653), .dinb(n19520), .dout(n19654));
  jxor g19480(.dina(n19517), .dinb(n19515), .dout(n19655));
  jand g19481(.dina(n19655), .dinb(n19654), .dout(n19656));
  jor  g19482(.dina(n19656), .dinb(n19518), .dout(n19657));
  jxor g19483(.dina(n19515), .dinb(n19513), .dout(n19658));
  jand g19484(.dina(n19658), .dinb(n19657), .dout(n19659));
  jor  g19485(.dina(n19659), .dinb(n19516), .dout(n19660));
  jxor g19486(.dina(n19513), .dinb(n19511), .dout(n19661));
  jand g19487(.dina(n19661), .dinb(n19660), .dout(n19662));
  jor  g19488(.dina(n19662), .dinb(n19514), .dout(n19663));
  jxor g19489(.dina(n19511), .dinb(n19510), .dout(n19664));
  jand g19490(.dina(n19664), .dinb(n19663), .dout(n19665));
  jor  g19491(.dina(n19665), .dinb(n19512), .dout(n19666));
  jnot g19492(.din(n22204), .dout(n19674));
  jand g19493(.dina(n19504), .dinb(n19474), .dout(n19675));
  jnot g19494(.din(n19675), .dout(n19676));
  jnot g19495(.din(n19474), .dout(n19677));
  jand g19496(.dina(n19503), .dinb(n19677), .dout(n19678));
  jor  g19497(.dina(n19678), .dinb(n19470), .dout(n19679));
  jand g19498(.dina(n19679), .dinb(n19676), .dout(n19680));
  jxor g19499(.dina(n19680), .dinb(n19674), .dout(n19681));
  jand g19500(.dina(n19492), .dinb(n19488), .dout(n19682));
  jnot g19501(.din(n19682), .dout(n19683));
  jor  g19502(.dina(n19502), .dinb(n19494), .dout(n19684));
  jand g19503(.dina(n19684), .dinb(n19683), .dout(n19685));
  jnot g19504(.din(n19685), .dout(n19686));
  jand g19505(.dina(n12841), .dinb(n4449), .dout(n19687));
  jand g19506(.dina(n12783), .dinb(n4453), .dout(n19688));
  jand g19507(.dina(n12766), .dinb(n4457), .dout(n19689));
  jand g19508(.dina(n12177), .dinb(n4461), .dout(n19690));
  jor  g19509(.dina(n19690), .dinb(n19689), .dout(n19691));
  jor  g19510(.dina(n19691), .dinb(n19688), .dout(n19692));
  jor  g19511(.dina(n19692), .dinb(n19687), .dout(n19693));
  jxor g19512(.dina(n19693), .dinb(n88), .dout(n19694));
  jnot g19513(.din(n19694), .dout(n19695));
  jor  g19514(.dina(n19479), .dinb(n19475), .dout(n19696));
  jand g19515(.dina(n19487), .dinb(n19480), .dout(n19697));
  jnot g19516(.din(n19697), .dout(n19698));
  jand g19517(.dina(n19698), .dinb(n19696), .dout(n19699));
  jnot g19518(.din(n19699), .dout(n19700));
  jand g19519(.dina(n3988), .dinb(n1023), .dout(n19701));
  jand g19520(.dina(n19701), .dinb(n3117), .dout(n19702));
  jand g19521(.dina(n566), .dinb(n465), .dout(n19703));
  jand g19522(.dina(n19703), .dinb(n13088), .dout(n19704));
  jand g19523(.dina(n1889), .dinb(n1424), .dout(n19705));
  jand g19524(.dina(n19705), .dinb(n19704), .dout(n19706));
  jand g19525(.dina(n3823), .dinb(n654), .dout(n19707));
  jand g19526(.dina(n19707), .dinb(n19706), .dout(n19708));
  jand g19527(.dina(n19708), .dinb(n19702), .dout(n19709));
  jand g19528(.dina(n1787), .dinb(n1025), .dout(n19710));
  jand g19529(.dina(n19710), .dinb(n1085), .dout(n19711));
  jand g19530(.dina(n687), .dinb(n494), .dout(n19712));
  jand g19531(.dina(n19712), .dinb(n897), .dout(n19713));
  jand g19532(.dina(n557), .dinb(n197), .dout(n19714));
  jand g19533(.dina(n19714), .dinb(n4287), .dout(n19715));
  jand g19534(.dina(n19715), .dinb(n19713), .dout(n19716));
  jand g19535(.dina(n19716), .dinb(n19711), .dout(n19717));
  jand g19536(.dina(n3978), .dinb(n781), .dout(n19718));
  jand g19537(.dina(n19718), .dinb(n6401), .dout(n19719));
  jand g19538(.dina(n19719), .dinb(n19717), .dout(n19720));
  jand g19539(.dina(n19720), .dinb(n19709), .dout(n19721));
  jand g19540(.dina(n19721), .dinb(n12712), .dout(n19722));
  jand g19541(.dina(n19722), .dinb(n5164), .dout(n19723));
  jxor g19542(.dina(n19723), .dinb(n19475), .dout(n19724));
  jxor g19543(.dina(n19724), .dinb(n19700), .dout(n19725));
  jand g19544(.dina(n12671), .dinb(n732), .dout(n19726));
  jand g19545(.dina(n11941), .dinb(n3855), .dout(n19727));
  jand g19546(.dina(n11942), .dinb(n3858), .dout(n19728));
  jand g19547(.dina(n11944), .dinb(n3851), .dout(n19729));
  jor  g19548(.dina(n19729), .dinb(n19728), .dout(n19730));
  jor  g19549(.dina(n19730), .dinb(n19727), .dout(n19731));
  jor  g19550(.dina(n19731), .dinb(n19726), .dout(n19732));
  jxor g19551(.dina(n19732), .dinb(n19725), .dout(n19733));
  jxor g19552(.dina(n19733), .dinb(n19695), .dout(n19734));
  jxor g19553(.dina(n19734), .dinb(n19686), .dout(n19735));
  jand g19554(.dina(n12919), .dinb(n75), .dout(n19736));
  jand g19555(.dina(n12815), .dinb(n4933), .dout(n19737));
  jand g19556(.dina(n12795), .dinb(n4918), .dout(n19738));
  jand g19557(.dina(n12782), .dinb(n4745), .dout(n19739));
  jor  g19558(.dina(n19739), .dinb(n19738), .dout(n19740));
  jor  g19559(.dina(n19740), .dinb(n19737), .dout(n19741));
  jor  g19560(.dina(n19741), .dinb(n19736), .dout(n19742));
  jxor g19561(.dina(n19742), .dinb(n68), .dout(n19743));
  jnot g19562(.din(n19743), .dout(n19744));
  jxor g19563(.dina(n19744), .dinb(n19735), .dout(n19745));
  jxor g19564(.dina(n19745), .dinb(n19681), .dout(n19746));
  jnot g19565(.din(n19461), .dout(n19747));
  jnot g19566(.din(n19506), .dout(n19748));
  jand g19567(.dina(n19748), .dinb(n19747), .dout(n19749));
  jnot g19568(.din(n19749), .dout(n19750));
  jand g19569(.dina(n19506), .dinb(n19461), .dout(n19751));
  jor  g19570(.dina(n19751), .dinb(n19458), .dout(n19752));
  jand g19571(.dina(n19752), .dinb(n19750), .dout(n19753));
  jxor g19572(.dina(n19753), .dinb(n19746), .dout(n19754));
  jand g19573(.dina(n19508), .dinb(n19449), .dout(n19755));
  jand g19574(.dina(n19509), .dinb(n19444), .dout(n19756));
  jor  g19575(.dina(n19756), .dinb(n19755), .dout(n19757));
  jxor g19576(.dina(n19757), .dinb(n19754), .dout(n19758));
  jxor g19577(.dina(n19758), .dinb(n19510), .dout(n19759));
  jxor g19578(.dina(n19759), .dinb(n19666), .dout(n19760));
  jand g19579(.dina(n19760), .dinb(n67), .dout(n19761));
  jand g19580(.dina(n19758), .dinb(n10827), .dout(n19762));
  jand g19581(.dina(n19510), .dinb(n10350), .dout(n19763));
  jand g19582(.dina(n19511), .dinb(n9917), .dout(n19764));
  jor  g19583(.dina(n19764), .dinb(n19763), .dout(n19765));
  jor  g19584(.dina(n19765), .dinb(n19762), .dout(n19766));
  jor  g19585(.dina(n19766), .dinb(n19761), .dout(n19767));
  jxor g19586(.dina(n19767), .dinb(n64), .dout(n19768));
  jnot g19587(.din(n19768), .dout(n19769));
  jxor g19588(.dina(n19643), .dinb(n19642), .dout(n19770));
  jand g19589(.dina(n19770), .dinb(n7890), .dout(n19771));
  jand g19590(.dina(n19523), .dinb(n8441), .dout(n19772));
  jand g19591(.dina(n19525), .dinb(n8154), .dout(n19773));
  jand g19592(.dina(n19527), .dinb(n7888), .dout(n19774));
  jor  g19593(.dina(n19774), .dinb(n19773), .dout(n19775));
  jor  g19594(.dina(n19775), .dinb(n19772), .dout(n19776));
  jor  g19595(.dina(n19776), .dinb(n19771), .dout(n19777));
  jxor g19596(.dina(n19777), .dinb(n5833), .dout(n19778));
  jnot g19597(.din(n19778), .dout(n19779));
  jxor g19598(.dina(n19631), .dinb(n19630), .dout(n19780));
  jand g19599(.dina(n19780), .dinb(n6936), .dout(n19781));
  jand g19600(.dina(n19531), .dinb(n7741), .dout(n19782));
  jand g19601(.dina(n19533), .dinb(n7613), .dout(n19783));
  jand g19602(.dina(n19535), .dinb(n6934), .dout(n19784));
  jor  g19603(.dina(n19784), .dinb(n19783), .dout(n19785));
  jor  g19604(.dina(n19785), .dinb(n19782), .dout(n19786));
  jor  g19605(.dina(n19786), .dinb(n19781), .dout(n19787));
  jxor g19606(.dina(n19787), .dinb(n5292), .dout(n19788));
  jnot g19607(.din(n19788), .dout(n19789));
  jxor g19608(.dina(n19590), .dinb(n19589), .dout(n19790));
  jor  g19609(.dina(n19790), .dinb(n5366), .dout(n19791));
  jor  g19610(.dina(n19562), .dinb(n5499), .dout(n19792));
  jor  g19611(.dina(n19564), .dinb(n5425), .dout(n19793));
  jor  g19612(.dina(n19566), .dinb(n5364), .dout(n19794));
  jand g19613(.dina(n19794), .dinb(n19793), .dout(n19795));
  jand g19614(.dina(n19795), .dinb(n19792), .dout(n19796));
  jand g19615(.dina(n19796), .dinb(n19791), .dout(n19797));
  jxor g19616(.dina(n19797), .dinb(\a[23] ), .dout(n19798));
  jnot g19617(.din(n19798), .dout(n19799));
  jxor g19618(.dina(n19570), .dinb(n19568), .dout(n19800));
  jxor g19619(.dina(n19579), .dinb(n19800), .dout(n19801));
  jor  g19620(.dina(n19801), .dinb(n4747), .dout(n19802));
  jor  g19621(.dina(n19568), .dinb(n4959), .dout(n19803));
  jor  g19622(.dina(n19570), .dinb(n4919), .dout(n19804));
  jor  g19623(.dina(n19575), .dinb(n4746), .dout(n19805));
  jand g19624(.dina(n19805), .dinb(n19804), .dout(n19806));
  jand g19625(.dina(n19806), .dinb(n19803), .dout(n19807));
  jand g19626(.dina(n19807), .dinb(n19802), .dout(n19808));
  jxor g19627(.dina(n19808), .dinb(\a[26] ), .dout(n19809));
  jnot g19628(.din(n19809), .dout(n19810));
  jand g19629(.dina(n19576), .dinb(n4447), .dout(n19811));
  jxor g19630(.dina(n19577), .dinb(n19574), .dout(n19812));
  jnot g19631(.din(n19812), .dout(n19813));
  jand g19632(.dina(n19813), .dinb(n75), .dout(n19814));
  jand g19633(.dina(n19576), .dinb(n4918), .dout(n19815));
  jand g19634(.dina(n19574), .dinb(n4933), .dout(n19816));
  jor  g19635(.dina(n19816), .dinb(n19815), .dout(n19817));
  jor  g19636(.dina(n19817), .dinb(n19814), .dout(n19818));
  jnot g19637(.din(n19818), .dout(n19819));
  jand g19638(.dina(n19576), .dinb(n74), .dout(n19820));
  jnot g19639(.din(n19820), .dout(n19821));
  jand g19640(.dina(n19821), .dinb(\a[26] ), .dout(n19822));
  jand g19641(.dina(n19822), .dinb(n19819), .dout(n19823));
  jand g19642(.dina(n19577), .dinb(n19574), .dout(n19824));
  jxor g19643(.dina(n19824), .dinb(n19570), .dout(n19825));
  jnot g19644(.din(n19825), .dout(n19826));
  jand g19645(.dina(n19826), .dinb(n75), .dout(n19827));
  jand g19646(.dina(n19572), .dinb(n4933), .dout(n19828));
  jand g19647(.dina(n19574), .dinb(n4918), .dout(n19829));
  jand g19648(.dina(n19576), .dinb(n4745), .dout(n19830));
  jor  g19649(.dina(n19830), .dinb(n19829), .dout(n19831));
  jor  g19650(.dina(n19831), .dinb(n19828), .dout(n19832));
  jor  g19651(.dina(n19832), .dinb(n19827), .dout(n19833));
  jnot g19652(.din(n19833), .dout(n19834));
  jand g19653(.dina(n19834), .dinb(n19823), .dout(n19835));
  jxor g19654(.dina(n19835), .dinb(n19811), .dout(n19836));
  jxor g19655(.dina(n19836), .dinb(n19810), .dout(n19837));
  jand g19656(.dina(n19837), .dinb(n19799), .dout(n19838));
  jxor g19657(.dina(n19586), .dinb(n19585), .dout(n19839));
  jor  g19658(.dina(n19839), .dinb(n5366), .dout(n19840));
  jor  g19659(.dina(n19564), .dinb(n5499), .dout(n19841));
  jor  g19660(.dina(n19566), .dinb(n5425), .dout(n19842));
  jor  g19661(.dina(n19568), .dinb(n5364), .dout(n19843));
  jand g19662(.dina(n19843), .dinb(n19842), .dout(n19844));
  jand g19663(.dina(n19844), .dinb(n19841), .dout(n19845));
  jand g19664(.dina(n19845), .dinb(n19840), .dout(n19846));
  jxor g19665(.dina(n19846), .dinb(\a[23] ), .dout(n19847));
  jnot g19666(.din(n19847), .dout(n19848));
  jor  g19667(.dina(n19823), .dinb(n68), .dout(n19849));
  jxor g19668(.dina(n19849), .dinb(n19834), .dout(n19850));
  jand g19669(.dina(n19850), .dinb(n19848), .dout(n19851));
  jxor g19670(.dina(n19582), .dinb(n19581), .dout(n19852));
  jor  g19671(.dina(n19852), .dinb(n5366), .dout(n19853));
  jor  g19672(.dina(n19566), .dinb(n5499), .dout(n19854));
  jor  g19673(.dina(n19568), .dinb(n5425), .dout(n19855));
  jor  g19674(.dina(n19570), .dinb(n5364), .dout(n19856));
  jand g19675(.dina(n19856), .dinb(n19855), .dout(n19857));
  jand g19676(.dina(n19857), .dinb(n19854), .dout(n19858));
  jand g19677(.dina(n19858), .dinb(n19853), .dout(n19859));
  jxor g19678(.dina(n19859), .dinb(\a[23] ), .dout(n19860));
  jnot g19679(.din(n19860), .dout(n19861));
  jand g19680(.dina(n19820), .dinb(\a[26] ), .dout(n19862));
  jxor g19681(.dina(n19862), .dinb(n19818), .dout(n19863));
  jand g19682(.dina(n19863), .dinb(n19861), .dout(n19864));
  jand g19683(.dina(n19813), .dinb(n5365), .dout(n19865));
  jand g19684(.dina(n19576), .dinb(n5424), .dout(n19866));
  jand g19685(.dina(n19574), .dinb(n5500), .dout(n19867));
  jor  g19686(.dina(n19867), .dinb(n19866), .dout(n19868));
  jor  g19687(.dina(n19868), .dinb(n19865), .dout(n19869));
  jnot g19688(.din(n19869), .dout(n19870));
  jand g19689(.dina(n19576), .dinb(n5358), .dout(n19871));
  jnot g19690(.din(n19871), .dout(n19872));
  jand g19691(.dina(n19872), .dinb(\a[23] ), .dout(n19873));
  jand g19692(.dina(n19873), .dinb(n19870), .dout(n19874));
  jand g19693(.dina(n19826), .dinb(n5365), .dout(n19875));
  jand g19694(.dina(n19572), .dinb(n5500), .dout(n19876));
  jand g19695(.dina(n19574), .dinb(n5424), .dout(n19877));
  jand g19696(.dina(n19576), .dinb(n5363), .dout(n19878));
  jor  g19697(.dina(n19878), .dinb(n19877), .dout(n19879));
  jor  g19698(.dina(n19879), .dinb(n19876), .dout(n19880));
  jor  g19699(.dina(n19880), .dinb(n19875), .dout(n19881));
  jnot g19700(.din(n19881), .dout(n19882));
  jand g19701(.dina(n19882), .dinb(n19874), .dout(n19883));
  jand g19702(.dina(n19883), .dinb(n19820), .dout(n19884));
  jor  g19703(.dina(n19801), .dinb(n5366), .dout(n19885));
  jor  g19704(.dina(n19568), .dinb(n5499), .dout(n19886));
  jor  g19705(.dina(n19570), .dinb(n5425), .dout(n19887));
  jor  g19706(.dina(n19575), .dinb(n5364), .dout(n19888));
  jand g19707(.dina(n19888), .dinb(n19887), .dout(n19889));
  jand g19708(.dina(n19889), .dinb(n19886), .dout(n19890));
  jand g19709(.dina(n19890), .dinb(n19885), .dout(n19891));
  jxor g19710(.dina(n19891), .dinb(\a[23] ), .dout(n19892));
  jnot g19711(.din(n19892), .dout(n19893));
  jxor g19712(.dina(n19883), .dinb(n19820), .dout(n19894));
  jand g19713(.dina(n19894), .dinb(n19893), .dout(n19895));
  jor  g19714(.dina(n19895), .dinb(n19884), .dout(n19896));
  jxor g19715(.dina(n19863), .dinb(n19861), .dout(n19897));
  jand g19716(.dina(n19897), .dinb(n19896), .dout(n19898));
  jor  g19717(.dina(n19898), .dinb(n19864), .dout(n19899));
  jxor g19718(.dina(n19850), .dinb(n19848), .dout(n19900));
  jand g19719(.dina(n19900), .dinb(n19899), .dout(n19901));
  jor  g19720(.dina(n19901), .dinb(n19851), .dout(n19902));
  jxor g19721(.dina(n19837), .dinb(n19799), .dout(n19903));
  jand g19722(.dina(n19903), .dinb(n19902), .dout(n19904));
  jor  g19723(.dina(n19904), .dinb(n19838), .dout(n19905));
  jxor g19724(.dina(n19594), .dinb(n19593), .dout(n19906));
  jor  g19725(.dina(n19906), .dinb(n5366), .dout(n19907));
  jor  g19726(.dina(n19558), .dinb(n5499), .dout(n19908));
  jor  g19727(.dina(n19562), .dinb(n5425), .dout(n19909));
  jor  g19728(.dina(n19564), .dinb(n5364), .dout(n19910));
  jand g19729(.dina(n19910), .dinb(n19909), .dout(n19911));
  jand g19730(.dina(n19911), .dinb(n19908), .dout(n19912));
  jand g19731(.dina(n19912), .dinb(n19907), .dout(n19913));
  jxor g19732(.dina(n19913), .dinb(\a[23] ), .dout(n19914));
  jnot g19733(.din(n19914), .dout(n19915));
  jand g19734(.dina(n19835), .dinb(n19811), .dout(n19916));
  jand g19735(.dina(n19836), .dinb(n19810), .dout(n19917));
  jor  g19736(.dina(n19917), .dinb(n19916), .dout(n19918));
  jor  g19737(.dina(n19852), .dinb(n4747), .dout(n19919));
  jor  g19738(.dina(n19566), .dinb(n4959), .dout(n19920));
  jor  g19739(.dina(n19568), .dinb(n4919), .dout(n19921));
  jor  g19740(.dina(n19570), .dinb(n4746), .dout(n19922));
  jand g19741(.dina(n19922), .dinb(n19921), .dout(n19923));
  jand g19742(.dina(n19923), .dinb(n19920), .dout(n19924));
  jand g19743(.dina(n19924), .dinb(n19919), .dout(n19925));
  jxor g19744(.dina(n19925), .dinb(\a[26] ), .dout(n19926));
  jnot g19745(.din(n19926), .dout(n19927));
  jand g19746(.dina(n19811), .dinb(\a[29] ), .dout(n19928));
  jand g19747(.dina(n19813), .dinb(n4449), .dout(n19929));
  jand g19748(.dina(n19576), .dinb(n4457), .dout(n19930));
  jand g19749(.dina(n19574), .dinb(n4453), .dout(n19931));
  jor  g19750(.dina(n19931), .dinb(n19930), .dout(n19932));
  jor  g19751(.dina(n19932), .dinb(n19929), .dout(n19933));
  jxor g19752(.dina(n19933), .dinb(n19928), .dout(n19934));
  jxor g19753(.dina(n19934), .dinb(n19927), .dout(n19935));
  jxor g19754(.dina(n19935), .dinb(n19918), .dout(n19936));
  jxor g19755(.dina(n19936), .dinb(n19915), .dout(n19937));
  jxor g19756(.dina(n19937), .dinb(n19905), .dout(n19938));
  jnot g19757(.din(n19938), .dout(n19939));
  jxor g19758(.dina(n19607), .dinb(n19605), .dout(n19940));
  jor  g19759(.dina(n19940), .dinb(n5694), .dout(n19941));
  jor  g19760(.dina(n19547), .dinb(n6208), .dout(n19942));
  jor  g19761(.dina(n19550), .dinb(n6132), .dout(n19943));
  jor  g19762(.dina(n19553), .dinb(n5692), .dout(n19944));
  jand g19763(.dina(n19944), .dinb(n19943), .dout(n19945));
  jand g19764(.dina(n19945), .dinb(n19942), .dout(n19946));
  jand g19765(.dina(n19946), .dinb(n19941), .dout(n19947));
  jxor g19766(.dina(n19947), .dinb(\a[20] ), .dout(n19948));
  jor  g19767(.dina(n19948), .dinb(n19939), .dout(n19949));
  jxor g19768(.dina(n19903), .dinb(n19902), .dout(n19950));
  jnot g19769(.din(n19950), .dout(n19951));
  jxor g19770(.dina(n19602), .dinb(n19601), .dout(n19952));
  jor  g19771(.dina(n19952), .dinb(n5694), .dout(n19953));
  jor  g19772(.dina(n19550), .dinb(n6208), .dout(n19954));
  jor  g19773(.dina(n19553), .dinb(n6132), .dout(n19955));
  jor  g19774(.dina(n19558), .dinb(n5692), .dout(n19956));
  jand g19775(.dina(n19956), .dinb(n19955), .dout(n19957));
  jand g19776(.dina(n19957), .dinb(n19954), .dout(n19958));
  jand g19777(.dina(n19958), .dinb(n19953), .dout(n19959));
  jxor g19778(.dina(n19959), .dinb(\a[20] ), .dout(n19960));
  jor  g19779(.dina(n19960), .dinb(n19951), .dout(n19961));
  jxor g19780(.dina(n19900), .dinb(n19899), .dout(n19962));
  jnot g19781(.din(n19962), .dout(n19963));
  jxor g19782(.dina(n19598), .dinb(n19597), .dout(n19964));
  jor  g19783(.dina(n19964), .dinb(n5694), .dout(n19965));
  jor  g19784(.dina(n19553), .dinb(n6208), .dout(n19966));
  jor  g19785(.dina(n19558), .dinb(n6132), .dout(n19967));
  jor  g19786(.dina(n19562), .dinb(n5692), .dout(n19968));
  jand g19787(.dina(n19968), .dinb(n19967), .dout(n19969));
  jand g19788(.dina(n19969), .dinb(n19966), .dout(n19970));
  jand g19789(.dina(n19970), .dinb(n19965), .dout(n19971));
  jxor g19790(.dina(n19971), .dinb(\a[20] ), .dout(n19972));
  jor  g19791(.dina(n19972), .dinb(n19963), .dout(n19973));
  jor  g19792(.dina(n19906), .dinb(n5694), .dout(n19974));
  jor  g19793(.dina(n19558), .dinb(n6208), .dout(n19975));
  jor  g19794(.dina(n19562), .dinb(n6132), .dout(n19976));
  jor  g19795(.dina(n19564), .dinb(n5692), .dout(n19977));
  jand g19796(.dina(n19977), .dinb(n19976), .dout(n19978));
  jand g19797(.dina(n19978), .dinb(n19975), .dout(n19979));
  jand g19798(.dina(n19979), .dinb(n19974), .dout(n19980));
  jxor g19799(.dina(n19980), .dinb(\a[20] ), .dout(n19981));
  jnot g19800(.din(n19981), .dout(n19982));
  jxor g19801(.dina(n19897), .dinb(n19896), .dout(n19983));
  jand g19802(.dina(n19983), .dinb(n19982), .dout(n19984));
  jor  g19803(.dina(n19790), .dinb(n5694), .dout(n19985));
  jor  g19804(.dina(n19562), .dinb(n6208), .dout(n19986));
  jor  g19805(.dina(n19564), .dinb(n6132), .dout(n19987));
  jor  g19806(.dina(n19566), .dinb(n5692), .dout(n19988));
  jand g19807(.dina(n19988), .dinb(n19987), .dout(n19989));
  jand g19808(.dina(n19989), .dinb(n19986), .dout(n19990));
  jand g19809(.dina(n19990), .dinb(n19985), .dout(n19991));
  jxor g19810(.dina(n19991), .dinb(\a[20] ), .dout(n19992));
  jnot g19811(.din(n19992), .dout(n19993));
  jxor g19812(.dina(n19894), .dinb(n19893), .dout(n19994));
  jand g19813(.dina(n19994), .dinb(n19993), .dout(n19995));
  jor  g19814(.dina(n19839), .dinb(n5694), .dout(n19996));
  jor  g19815(.dina(n19564), .dinb(n6208), .dout(n19997));
  jor  g19816(.dina(n19566), .dinb(n6132), .dout(n19998));
  jor  g19817(.dina(n19568), .dinb(n5692), .dout(n19999));
  jand g19818(.dina(n19999), .dinb(n19998), .dout(n20000));
  jand g19819(.dina(n20000), .dinb(n19997), .dout(n20001));
  jand g19820(.dina(n20001), .dinb(n19996), .dout(n20002));
  jxor g19821(.dina(n20002), .dinb(\a[20] ), .dout(n20003));
  jnot g19822(.din(n20003), .dout(n20004));
  jor  g19823(.dina(n19874), .dinb(n72), .dout(n20005));
  jxor g19824(.dina(n20005), .dinb(n19882), .dout(n20006));
  jand g19825(.dina(n20006), .dinb(n20004), .dout(n20007));
  jor  g19826(.dina(n19852), .dinb(n5694), .dout(n20008));
  jor  g19827(.dina(n19566), .dinb(n6208), .dout(n20009));
  jor  g19828(.dina(n19568), .dinb(n6132), .dout(n20010));
  jor  g19829(.dina(n19570), .dinb(n5692), .dout(n20011));
  jand g19830(.dina(n20011), .dinb(n20010), .dout(n20012));
  jand g19831(.dina(n20012), .dinb(n20009), .dout(n20013));
  jand g19832(.dina(n20013), .dinb(n20008), .dout(n20014));
  jxor g19833(.dina(n20014), .dinb(\a[20] ), .dout(n20015));
  jnot g19834(.din(n20015), .dout(n20016));
  jand g19835(.dina(n19871), .dinb(\a[23] ), .dout(n20017));
  jxor g19836(.dina(n20017), .dinb(n19869), .dout(n20018));
  jand g19837(.dina(n20018), .dinb(n20016), .dout(n20019));
  jand g19838(.dina(n19813), .dinb(n5693), .dout(n20020));
  jand g19839(.dina(n19576), .dinb(n6131), .dout(n20021));
  jand g19840(.dina(n19574), .dinb(n6209), .dout(n20022));
  jor  g19841(.dina(n20022), .dinb(n20021), .dout(n20023));
  jor  g19842(.dina(n20023), .dinb(n20020), .dout(n20024));
  jnot g19843(.din(n20024), .dout(n20025));
  jand g19844(.dina(n19576), .dinb(n5687), .dout(n20026));
  jnot g19845(.din(n20026), .dout(n20027));
  jand g19846(.dina(n20027), .dinb(\a[20] ), .dout(n20028));
  jand g19847(.dina(n20028), .dinb(n20025), .dout(n20029));
  jand g19848(.dina(n19826), .dinb(n5693), .dout(n20030));
  jand g19849(.dina(n19572), .dinb(n6209), .dout(n20031));
  jand g19850(.dina(n19574), .dinb(n6131), .dout(n20032));
  jand g19851(.dina(n19576), .dinb(n5691), .dout(n20033));
  jor  g19852(.dina(n20033), .dinb(n20032), .dout(n20034));
  jor  g19853(.dina(n20034), .dinb(n20031), .dout(n20035));
  jor  g19854(.dina(n20035), .dinb(n20030), .dout(n20036));
  jnot g19855(.din(n20036), .dout(n20037));
  jand g19856(.dina(n20037), .dinb(n20029), .dout(n20038));
  jand g19857(.dina(n20038), .dinb(n19871), .dout(n20039));
  jor  g19858(.dina(n19801), .dinb(n5694), .dout(n20040));
  jor  g19859(.dina(n19568), .dinb(n6208), .dout(n20041));
  jor  g19860(.dina(n19570), .dinb(n6132), .dout(n20042));
  jor  g19861(.dina(n19575), .dinb(n5692), .dout(n20043));
  jand g19862(.dina(n20043), .dinb(n20042), .dout(n20044));
  jand g19863(.dina(n20044), .dinb(n20041), .dout(n20045));
  jand g19864(.dina(n20045), .dinb(n20040), .dout(n20046));
  jxor g19865(.dina(n20046), .dinb(\a[20] ), .dout(n20047));
  jnot g19866(.din(n20047), .dout(n20048));
  jxor g19867(.dina(n20038), .dinb(n19871), .dout(n20049));
  jand g19868(.dina(n20049), .dinb(n20048), .dout(n20050));
  jor  g19869(.dina(n20050), .dinb(n20039), .dout(n20051));
  jxor g19870(.dina(n20018), .dinb(n20016), .dout(n20052));
  jand g19871(.dina(n20052), .dinb(n20051), .dout(n20053));
  jor  g19872(.dina(n20053), .dinb(n20019), .dout(n20054));
  jxor g19873(.dina(n20006), .dinb(n20004), .dout(n20055));
  jand g19874(.dina(n20055), .dinb(n20054), .dout(n20056));
  jor  g19875(.dina(n20056), .dinb(n20007), .dout(n20057));
  jxor g19876(.dina(n19994), .dinb(n19993), .dout(n20058));
  jand g19877(.dina(n20058), .dinb(n20057), .dout(n20059));
  jor  g19878(.dina(n20059), .dinb(n19995), .dout(n20060));
  jxor g19879(.dina(n19983), .dinb(n19982), .dout(n20061));
  jand g19880(.dina(n20061), .dinb(n20060), .dout(n20062));
  jor  g19881(.dina(n20062), .dinb(n19984), .dout(n20063));
  jxor g19882(.dina(n19972), .dinb(n19963), .dout(n20064));
  jand g19883(.dina(n20064), .dinb(n20063), .dout(n20065));
  jnot g19884(.din(n20065), .dout(n20066));
  jand g19885(.dina(n20066), .dinb(n19973), .dout(n20067));
  jnot g19886(.din(n20067), .dout(n20068));
  jxor g19887(.dina(n19960), .dinb(n19951), .dout(n20069));
  jand g19888(.dina(n20069), .dinb(n20068), .dout(n20070));
  jnot g19889(.din(n20070), .dout(n20071));
  jand g19890(.dina(n20071), .dinb(n19961), .dout(n20072));
  jnot g19891(.din(n20072), .dout(n20073));
  jxor g19892(.dina(n19948), .dinb(n19939), .dout(n20074));
  jand g19893(.dina(n20074), .dinb(n20073), .dout(n20075));
  jnot g19894(.din(n20075), .dout(n20076));
  jand g19895(.dina(n20076), .dinb(n19949), .dout(n20077));
  jnot g19896(.din(n20077), .dout(n20078));
  jxor g19897(.dina(n19610), .dinb(n19609), .dout(n20079));
  jand g19898(.dina(n20079), .dinb(n5693), .dout(n20080));
  jand g19899(.dina(n19545), .dinb(n6209), .dout(n20081));
  jand g19900(.dina(n19548), .dinb(n6131), .dout(n20082));
  jand g19901(.dina(n19551), .dinb(n5691), .dout(n20083));
  jor  g19902(.dina(n20083), .dinb(n20082), .dout(n20084));
  jor  g19903(.dina(n20084), .dinb(n20081), .dout(n20085));
  jor  g19904(.dina(n20085), .dinb(n20080), .dout(n20086));
  jxor g19905(.dina(n20086), .dinb(n4247), .dout(n20087));
  jnot g19906(.din(n20087), .dout(n20088));
  jand g19907(.dina(n19936), .dinb(n19915), .dout(n20089));
  jand g19908(.dina(n19937), .dinb(n19905), .dout(n20090));
  jor  g19909(.dina(n20090), .dinb(n20089), .dout(n20091));
  jand g19910(.dina(n19934), .dinb(n19927), .dout(n20092));
  jand g19911(.dina(n19935), .dinb(n19918), .dout(n20093));
  jor  g19912(.dina(n20093), .dinb(n20092), .dout(n20094));
  jor  g19913(.dina(n19839), .dinb(n4747), .dout(n20095));
  jor  g19914(.dina(n19564), .dinb(n4959), .dout(n20096));
  jor  g19915(.dina(n19566), .dinb(n4919), .dout(n20097));
  jor  g19916(.dina(n19568), .dinb(n4746), .dout(n20098));
  jand g19917(.dina(n20098), .dinb(n20097), .dout(n20099));
  jand g19918(.dina(n20099), .dinb(n20096), .dout(n20100));
  jand g19919(.dina(n20100), .dinb(n20095), .dout(n20101));
  jxor g19920(.dina(n20101), .dinb(\a[26] ), .dout(n20102));
  jnot g19921(.din(n20102), .dout(n20103));
  jor  g19922(.dina(n19811), .dinb(n88), .dout(n20104));
  jor  g19923(.dina(n20104), .dinb(n19933), .dout(n20105));
  jand g19924(.dina(n20105), .dinb(\a[29] ), .dout(n20106));
  jand g19925(.dina(n19826), .dinb(n4449), .dout(n20107));
  jand g19926(.dina(n19572), .dinb(n4453), .dout(n20108));
  jand g19927(.dina(n19574), .dinb(n4457), .dout(n20109));
  jand g19928(.dina(n19576), .dinb(n4461), .dout(n20110));
  jor  g19929(.dina(n20110), .dinb(n20109), .dout(n20111));
  jor  g19930(.dina(n20111), .dinb(n20108), .dout(n20112));
  jor  g19931(.dina(n20112), .dinb(n20107), .dout(n20113));
  jxor g19932(.dina(n20113), .dinb(n20106), .dout(n20114));
  jxor g19933(.dina(n20114), .dinb(n20103), .dout(n20115));
  jxor g19934(.dina(n20115), .dinb(n20094), .dout(n20116));
  jnot g19935(.din(n20116), .dout(n20117));
  jor  g19936(.dina(n19964), .dinb(n5366), .dout(n20118));
  jor  g19937(.dina(n19553), .dinb(n5499), .dout(n20119));
  jor  g19938(.dina(n19558), .dinb(n5425), .dout(n20120));
  jor  g19939(.dina(n19562), .dinb(n5364), .dout(n20121));
  jand g19940(.dina(n20121), .dinb(n20120), .dout(n20122));
  jand g19941(.dina(n20122), .dinb(n20119), .dout(n20123));
  jand g19942(.dina(n20123), .dinb(n20118), .dout(n20124));
  jxor g19943(.dina(n20124), .dinb(\a[23] ), .dout(n20125));
  jxor g19944(.dina(n20125), .dinb(n20117), .dout(n20126));
  jxor g19945(.dina(n20126), .dinb(n20091), .dout(n20127));
  jxor g19946(.dina(n20127), .dinb(n20088), .dout(n20128));
  jxor g19947(.dina(n20128), .dinb(n20078), .dout(n20129));
  jnot g19948(.din(n20129), .dout(n20130));
  jxor g19949(.dina(n19619), .dinb(n19618), .dout(n20131));
  jand g19950(.dina(n20131), .dinb(n6340), .dout(n20132));
  jand g19951(.dina(n19539), .dinb(n6798), .dout(n20133));
  jand g19952(.dina(n19541), .dinb(n6556), .dout(n20134));
  jand g19953(.dina(n19543), .dinb(n6338), .dout(n20135));
  jor  g19954(.dina(n20135), .dinb(n20134), .dout(n20136));
  jor  g19955(.dina(n20136), .dinb(n20133), .dout(n20137));
  jor  g19956(.dina(n20137), .dinb(n20132), .dout(n20138));
  jxor g19957(.dina(n20138), .dinb(n5064), .dout(n20139));
  jor  g19958(.dina(n20139), .dinb(n20130), .dout(n20140));
  jxor g19959(.dina(n19616), .dinb(n19615), .dout(n20141));
  jand g19960(.dina(n20141), .dinb(n6340), .dout(n20142));
  jand g19961(.dina(n19541), .dinb(n6798), .dout(n20143));
  jand g19962(.dina(n19543), .dinb(n6556), .dout(n20144));
  jand g19963(.dina(n19545), .dinb(n6338), .dout(n20145));
  jor  g19964(.dina(n20145), .dinb(n20144), .dout(n20146));
  jor  g19965(.dina(n20146), .dinb(n20143), .dout(n20147));
  jor  g19966(.dina(n20147), .dinb(n20142), .dout(n20148));
  jxor g19967(.dina(n20148), .dinb(n5064), .dout(n20149));
  jnot g19968(.din(n20149), .dout(n20150));
  jxor g19969(.dina(n20074), .dinb(n20073), .dout(n20151));
  jand g19970(.dina(n20151), .dinb(n20150), .dout(n20152));
  jxor g19971(.dina(n19613), .dinb(n19612), .dout(n20153));
  jand g19972(.dina(n20153), .dinb(n6340), .dout(n20154));
  jand g19973(.dina(n19543), .dinb(n6798), .dout(n20155));
  jand g19974(.dina(n19545), .dinb(n6556), .dout(n20156));
  jand g19975(.dina(n19548), .dinb(n6338), .dout(n20157));
  jor  g19976(.dina(n20157), .dinb(n20156), .dout(n20158));
  jor  g19977(.dina(n20158), .dinb(n20155), .dout(n20159));
  jor  g19978(.dina(n20159), .dinb(n20154), .dout(n20160));
  jxor g19979(.dina(n20160), .dinb(n5064), .dout(n20161));
  jnot g19980(.din(n20161), .dout(n20162));
  jxor g19981(.dina(n20069), .dinb(n20068), .dout(n20163));
  jand g19982(.dina(n20163), .dinb(n20162), .dout(n20164));
  jand g19983(.dina(n20079), .dinb(n6340), .dout(n20165));
  jand g19984(.dina(n19545), .dinb(n6798), .dout(n20166));
  jand g19985(.dina(n19548), .dinb(n6556), .dout(n20167));
  jand g19986(.dina(n19551), .dinb(n6338), .dout(n20168));
  jor  g19987(.dina(n20168), .dinb(n20167), .dout(n20169));
  jor  g19988(.dina(n20169), .dinb(n20166), .dout(n20170));
  jor  g19989(.dina(n20170), .dinb(n20165), .dout(n20171));
  jxor g19990(.dina(n20171), .dinb(n5064), .dout(n20172));
  jnot g19991(.din(n20172), .dout(n20173));
  jxor g19992(.dina(n20064), .dinb(n20063), .dout(n20174));
  jand g19993(.dina(n20174), .dinb(n20173), .dout(n20175));
  jxor g19994(.dina(n20061), .dinb(n20060), .dout(n20176));
  jnot g19995(.din(n20176), .dout(n20177));
  jor  g19996(.dina(n19940), .dinb(n6341), .dout(n20178));
  jor  g19997(.dina(n19547), .dinb(n6797), .dout(n20179));
  jor  g19998(.dina(n19550), .dinb(n6557), .dout(n20180));
  jor  g19999(.dina(n19553), .dinb(n6339), .dout(n20181));
  jand g20000(.dina(n20181), .dinb(n20180), .dout(n20182));
  jand g20001(.dina(n20182), .dinb(n20179), .dout(n20183));
  jand g20002(.dina(n20183), .dinb(n20178), .dout(n20184));
  jxor g20003(.dina(n20184), .dinb(\a[17] ), .dout(n20185));
  jor  g20004(.dina(n20185), .dinb(n20177), .dout(n20186));
  jxor g20005(.dina(n20058), .dinb(n20057), .dout(n20187));
  jnot g20006(.din(n20187), .dout(n20188));
  jor  g20007(.dina(n19952), .dinb(n6341), .dout(n20189));
  jor  g20008(.dina(n19550), .dinb(n6797), .dout(n20190));
  jor  g20009(.dina(n19553), .dinb(n6557), .dout(n20191));
  jor  g20010(.dina(n19558), .dinb(n6339), .dout(n20192));
  jand g20011(.dina(n20192), .dinb(n20191), .dout(n20193));
  jand g20012(.dina(n20193), .dinb(n20190), .dout(n20194));
  jand g20013(.dina(n20194), .dinb(n20189), .dout(n20195));
  jxor g20014(.dina(n20195), .dinb(\a[17] ), .dout(n20196));
  jor  g20015(.dina(n20196), .dinb(n20188), .dout(n20197));
  jxor g20016(.dina(n20055), .dinb(n20054), .dout(n20198));
  jnot g20017(.din(n20198), .dout(n20199));
  jor  g20018(.dina(n19964), .dinb(n6341), .dout(n20200));
  jor  g20019(.dina(n19553), .dinb(n6797), .dout(n20201));
  jor  g20020(.dina(n19558), .dinb(n6557), .dout(n20202));
  jor  g20021(.dina(n19562), .dinb(n6339), .dout(n20203));
  jand g20022(.dina(n20203), .dinb(n20202), .dout(n20204));
  jand g20023(.dina(n20204), .dinb(n20201), .dout(n20205));
  jand g20024(.dina(n20205), .dinb(n20200), .dout(n20206));
  jxor g20025(.dina(n20206), .dinb(\a[17] ), .dout(n20207));
  jor  g20026(.dina(n20207), .dinb(n20199), .dout(n20208));
  jor  g20027(.dina(n19906), .dinb(n6341), .dout(n20209));
  jor  g20028(.dina(n19558), .dinb(n6797), .dout(n20210));
  jor  g20029(.dina(n19562), .dinb(n6557), .dout(n20211));
  jor  g20030(.dina(n19564), .dinb(n6339), .dout(n20212));
  jand g20031(.dina(n20212), .dinb(n20211), .dout(n20213));
  jand g20032(.dina(n20213), .dinb(n20210), .dout(n20214));
  jand g20033(.dina(n20214), .dinb(n20209), .dout(n20215));
  jxor g20034(.dina(n20215), .dinb(\a[17] ), .dout(n20216));
  jnot g20035(.din(n20216), .dout(n20217));
  jxor g20036(.dina(n20052), .dinb(n20051), .dout(n20218));
  jand g20037(.dina(n20218), .dinb(n20217), .dout(n20219));
  jor  g20038(.dina(n19790), .dinb(n6341), .dout(n20220));
  jor  g20039(.dina(n19562), .dinb(n6797), .dout(n20221));
  jor  g20040(.dina(n19564), .dinb(n6557), .dout(n20222));
  jor  g20041(.dina(n19566), .dinb(n6339), .dout(n20223));
  jand g20042(.dina(n20223), .dinb(n20222), .dout(n20224));
  jand g20043(.dina(n20224), .dinb(n20221), .dout(n20225));
  jand g20044(.dina(n20225), .dinb(n20220), .dout(n20226));
  jxor g20045(.dina(n20226), .dinb(\a[17] ), .dout(n20227));
  jnot g20046(.din(n20227), .dout(n20228));
  jxor g20047(.dina(n20049), .dinb(n20048), .dout(n20229));
  jand g20048(.dina(n20229), .dinb(n20228), .dout(n20230));
  jor  g20049(.dina(n19839), .dinb(n6341), .dout(n20231));
  jor  g20050(.dina(n19564), .dinb(n6797), .dout(n20232));
  jor  g20051(.dina(n19566), .dinb(n6557), .dout(n20233));
  jor  g20052(.dina(n19568), .dinb(n6339), .dout(n20234));
  jand g20053(.dina(n20234), .dinb(n20233), .dout(n20235));
  jand g20054(.dina(n20235), .dinb(n20232), .dout(n20236));
  jand g20055(.dina(n20236), .dinb(n20231), .dout(n20237));
  jxor g20056(.dina(n20237), .dinb(\a[17] ), .dout(n20238));
  jnot g20057(.din(n20238), .dout(n20239));
  jor  g20058(.dina(n20029), .dinb(n4247), .dout(n20240));
  jxor g20059(.dina(n20240), .dinb(n20037), .dout(n20241));
  jand g20060(.dina(n20241), .dinb(n20239), .dout(n20242));
  jor  g20061(.dina(n19852), .dinb(n6341), .dout(n20243));
  jor  g20062(.dina(n19566), .dinb(n6797), .dout(n20244));
  jor  g20063(.dina(n19568), .dinb(n6557), .dout(n20245));
  jor  g20064(.dina(n19570), .dinb(n6339), .dout(n20246));
  jand g20065(.dina(n20246), .dinb(n20245), .dout(n20247));
  jand g20066(.dina(n20247), .dinb(n20244), .dout(n20248));
  jand g20067(.dina(n20248), .dinb(n20243), .dout(n20249));
  jxor g20068(.dina(n20249), .dinb(\a[17] ), .dout(n20250));
  jnot g20069(.din(n20250), .dout(n20251));
  jand g20070(.dina(n20026), .dinb(\a[20] ), .dout(n20252));
  jxor g20071(.dina(n20252), .dinb(n20024), .dout(n20253));
  jand g20072(.dina(n20253), .dinb(n20251), .dout(n20254));
  jand g20073(.dina(n19813), .dinb(n6340), .dout(n20255));
  jand g20074(.dina(n19576), .dinb(n6556), .dout(n20256));
  jand g20075(.dina(n19574), .dinb(n6798), .dout(n20257));
  jor  g20076(.dina(n20257), .dinb(n20256), .dout(n20258));
  jor  g20077(.dina(n20258), .dinb(n20255), .dout(n20259));
  jnot g20078(.din(n20259), .dout(n20260));
  jand g20079(.dina(n19576), .dinb(n6334), .dout(n20261));
  jnot g20080(.din(n20261), .dout(n20262));
  jand g20081(.dina(n20262), .dinb(\a[17] ), .dout(n20263));
  jand g20082(.dina(n20263), .dinb(n20260), .dout(n20264));
  jand g20083(.dina(n19826), .dinb(n6340), .dout(n20265));
  jand g20084(.dina(n19572), .dinb(n6798), .dout(n20266));
  jand g20085(.dina(n19574), .dinb(n6556), .dout(n20267));
  jand g20086(.dina(n19576), .dinb(n6338), .dout(n20268));
  jor  g20087(.dina(n20268), .dinb(n20267), .dout(n20269));
  jor  g20088(.dina(n20269), .dinb(n20266), .dout(n20270));
  jor  g20089(.dina(n20270), .dinb(n20265), .dout(n20271));
  jnot g20090(.din(n20271), .dout(n20272));
  jand g20091(.dina(n20272), .dinb(n20264), .dout(n20273));
  jand g20092(.dina(n20273), .dinb(n20026), .dout(n20274));
  jor  g20093(.dina(n19801), .dinb(n6341), .dout(n20275));
  jor  g20094(.dina(n19568), .dinb(n6797), .dout(n20276));
  jor  g20095(.dina(n19570), .dinb(n6557), .dout(n20277));
  jor  g20096(.dina(n19575), .dinb(n6339), .dout(n20278));
  jand g20097(.dina(n20278), .dinb(n20277), .dout(n20279));
  jand g20098(.dina(n20279), .dinb(n20276), .dout(n20280));
  jand g20099(.dina(n20280), .dinb(n20275), .dout(n20281));
  jxor g20100(.dina(n20281), .dinb(\a[17] ), .dout(n20282));
  jnot g20101(.din(n20282), .dout(n20283));
  jxor g20102(.dina(n20273), .dinb(n20026), .dout(n20284));
  jand g20103(.dina(n20284), .dinb(n20283), .dout(n20285));
  jor  g20104(.dina(n20285), .dinb(n20274), .dout(n20286));
  jxor g20105(.dina(n20253), .dinb(n20251), .dout(n20287));
  jand g20106(.dina(n20287), .dinb(n20286), .dout(n20288));
  jor  g20107(.dina(n20288), .dinb(n20254), .dout(n20289));
  jxor g20108(.dina(n20241), .dinb(n20239), .dout(n20290));
  jand g20109(.dina(n20290), .dinb(n20289), .dout(n20291));
  jor  g20110(.dina(n20291), .dinb(n20242), .dout(n20292));
  jxor g20111(.dina(n20229), .dinb(n20228), .dout(n20293));
  jand g20112(.dina(n20293), .dinb(n20292), .dout(n20294));
  jor  g20113(.dina(n20294), .dinb(n20230), .dout(n20295));
  jxor g20114(.dina(n20218), .dinb(n20217), .dout(n20296));
  jand g20115(.dina(n20296), .dinb(n20295), .dout(n20297));
  jor  g20116(.dina(n20297), .dinb(n20219), .dout(n20298));
  jxor g20117(.dina(n20207), .dinb(n20199), .dout(n20299));
  jand g20118(.dina(n20299), .dinb(n20298), .dout(n20300));
  jnot g20119(.din(n20300), .dout(n20301));
  jand g20120(.dina(n20301), .dinb(n20208), .dout(n20302));
  jnot g20121(.din(n20302), .dout(n20303));
  jxor g20122(.dina(n20196), .dinb(n20188), .dout(n20304));
  jand g20123(.dina(n20304), .dinb(n20303), .dout(n20305));
  jnot g20124(.din(n20305), .dout(n20306));
  jand g20125(.dina(n20306), .dinb(n20197), .dout(n20307));
  jnot g20126(.din(n20307), .dout(n20308));
  jxor g20127(.dina(n20185), .dinb(n20177), .dout(n20309));
  jand g20128(.dina(n20309), .dinb(n20308), .dout(n20310));
  jnot g20129(.din(n20310), .dout(n20311));
  jand g20130(.dina(n20311), .dinb(n20186), .dout(n20312));
  jnot g20131(.din(n20312), .dout(n20313));
  jxor g20132(.dina(n20174), .dinb(n20173), .dout(n20314));
  jand g20133(.dina(n20314), .dinb(n20313), .dout(n20315));
  jor  g20134(.dina(n20315), .dinb(n20175), .dout(n20316));
  jxor g20135(.dina(n20163), .dinb(n20162), .dout(n20317));
  jand g20136(.dina(n20317), .dinb(n20316), .dout(n20318));
  jor  g20137(.dina(n20318), .dinb(n20164), .dout(n20319));
  jxor g20138(.dina(n20151), .dinb(n20150), .dout(n20320));
  jand g20139(.dina(n20320), .dinb(n20319), .dout(n20321));
  jor  g20140(.dina(n20321), .dinb(n20152), .dout(n20322));
  jxor g20141(.dina(n20139), .dinb(n20130), .dout(n20323));
  jand g20142(.dina(n20323), .dinb(n20322), .dout(n20324));
  jnot g20143(.din(n20324), .dout(n20325));
  jand g20144(.dina(n20325), .dinb(n20140), .dout(n20326));
  jnot g20145(.din(n20326), .dout(n20327));
  jand g20146(.dina(n20127), .dinb(n20088), .dout(n20328));
  jand g20147(.dina(n20128), .dinb(n20078), .dout(n20329));
  jor  g20148(.dina(n20329), .dinb(n20328), .dout(n20330));
  jand g20149(.dina(n20153), .dinb(n5693), .dout(n20331));
  jand g20150(.dina(n19543), .dinb(n6209), .dout(n20332));
  jand g20151(.dina(n19545), .dinb(n6131), .dout(n20333));
  jand g20152(.dina(n19548), .dinb(n5691), .dout(n20334));
  jor  g20153(.dina(n20334), .dinb(n20333), .dout(n20335));
  jor  g20154(.dina(n20335), .dinb(n20332), .dout(n20336));
  jor  g20155(.dina(n20336), .dinb(n20331), .dout(n20337));
  jxor g20156(.dina(n20337), .dinb(n4247), .dout(n20338));
  jnot g20157(.din(n20338), .dout(n20339));
  jor  g20158(.dina(n20125), .dinb(n20117), .dout(n20340));
  jand g20159(.dina(n20126), .dinb(n20091), .dout(n20341));
  jnot g20160(.din(n20341), .dout(n20342));
  jand g20161(.dina(n20342), .dinb(n20340), .dout(n20343));
  jnot g20162(.din(n20343), .dout(n20344));
  jand g20163(.dina(n20114), .dinb(n20103), .dout(n20345));
  jand g20164(.dina(n20115), .dinb(n20094), .dout(n20346));
  jor  g20165(.dina(n20346), .dinb(n20345), .dout(n20347));
  jor  g20166(.dina(n19790), .dinb(n4747), .dout(n20348));
  jor  g20167(.dina(n19562), .dinb(n4959), .dout(n20349));
  jor  g20168(.dina(n19564), .dinb(n4919), .dout(n20350));
  jor  g20169(.dina(n19566), .dinb(n4746), .dout(n20351));
  jand g20170(.dina(n20351), .dinb(n20350), .dout(n20352));
  jand g20171(.dina(n20352), .dinb(n20349), .dout(n20353));
  jand g20172(.dina(n20353), .dinb(n20348), .dout(n20354));
  jxor g20173(.dina(n20354), .dinb(\a[26] ), .dout(n20355));
  jnot g20174(.din(n20355), .dout(n20356));
  jor  g20175(.dina(n19801), .dinb(n4724), .dout(n20357));
  jor  g20176(.dina(n19568), .dinb(n4905), .dout(n20358));
  jor  g20177(.dina(n19570), .dinb(n4735), .dout(n20359));
  jor  g20178(.dina(n19575), .dinb(n4733), .dout(n20360));
  jand g20179(.dina(n20360), .dinb(n20359), .dout(n20361));
  jand g20180(.dina(n20361), .dinb(n20358), .dout(n20362));
  jand g20181(.dina(n20362), .dinb(n20357), .dout(n20363));
  jxor g20182(.dina(n20363), .dinb(\a[29] ), .dout(n20364));
  jnot g20183(.din(n20364), .dout(n20365));
  jor  g20184(.dina(n20113), .dinb(n20105), .dout(n20366));
  jnot g20185(.din(n20366), .dout(n20367));
  jand g20186(.dina(n19576), .dinb(n731), .dout(n20368));
  jxor g20187(.dina(n20368), .dinb(n20367), .dout(n20369));
  jxor g20188(.dina(n20369), .dinb(n20365), .dout(n20370));
  jxor g20189(.dina(n20370), .dinb(n20356), .dout(n20371));
  jxor g20190(.dina(n20371), .dinb(n20347), .dout(n20372));
  jnot g20191(.din(n20372), .dout(n20373));
  jor  g20192(.dina(n19952), .dinb(n5366), .dout(n20374));
  jor  g20193(.dina(n19550), .dinb(n5499), .dout(n20375));
  jor  g20194(.dina(n19553), .dinb(n5425), .dout(n20376));
  jor  g20195(.dina(n19558), .dinb(n5364), .dout(n20377));
  jand g20196(.dina(n20377), .dinb(n20376), .dout(n20378));
  jand g20197(.dina(n20378), .dinb(n20375), .dout(n20379));
  jand g20198(.dina(n20379), .dinb(n20374), .dout(n20380));
  jxor g20199(.dina(n20380), .dinb(\a[23] ), .dout(n20381));
  jxor g20200(.dina(n20381), .dinb(n20373), .dout(n20382));
  jxor g20201(.dina(n20382), .dinb(n20344), .dout(n20383));
  jxor g20202(.dina(n20383), .dinb(n20339), .dout(n20384));
  jxor g20203(.dina(n20384), .dinb(n20330), .dout(n20385));
  jnot g20204(.din(n20385), .dout(n20386));
  jxor g20205(.dina(n19622), .dinb(n19621), .dout(n20387));
  jand g20206(.dina(n20387), .dinb(n6340), .dout(n20388));
  jand g20207(.dina(n19537), .dinb(n6798), .dout(n20389));
  jand g20208(.dina(n19539), .dinb(n6556), .dout(n20390));
  jand g20209(.dina(n19541), .dinb(n6338), .dout(n20391));
  jor  g20210(.dina(n20391), .dinb(n20390), .dout(n20392));
  jor  g20211(.dina(n20392), .dinb(n20389), .dout(n20393));
  jor  g20212(.dina(n20393), .dinb(n20388), .dout(n20394));
  jxor g20213(.dina(n20394), .dinb(n5064), .dout(n20395));
  jxor g20214(.dina(n20395), .dinb(n20386), .dout(n20396));
  jxor g20215(.dina(n20396), .dinb(n20327), .dout(n20397));
  jand g20216(.dina(n20397), .dinb(n19789), .dout(n20398));
  jxor g20217(.dina(n19628), .dinb(n19627), .dout(n20399));
  jand g20218(.dina(n20399), .dinb(n6936), .dout(n20400));
  jand g20219(.dina(n19533), .dinb(n7741), .dout(n20401));
  jand g20220(.dina(n19535), .dinb(n7613), .dout(n20402));
  jand g20221(.dina(n19537), .dinb(n6934), .dout(n20403));
  jor  g20222(.dina(n20403), .dinb(n20402), .dout(n20404));
  jor  g20223(.dina(n20404), .dinb(n20401), .dout(n20405));
  jor  g20224(.dina(n20405), .dinb(n20400), .dout(n20406));
  jxor g20225(.dina(n20406), .dinb(n5292), .dout(n20407));
  jnot g20226(.din(n20407), .dout(n20408));
  jxor g20227(.dina(n20323), .dinb(n20322), .dout(n20409));
  jand g20228(.dina(n20409), .dinb(n20408), .dout(n20410));
  jxor g20229(.dina(n20320), .dinb(n20319), .dout(n20411));
  jnot g20230(.din(n20411), .dout(n20412));
  jxor g20231(.dina(n19625), .dinb(n19624), .dout(n20413));
  jand g20232(.dina(n20413), .dinb(n6936), .dout(n20414));
  jand g20233(.dina(n19535), .dinb(n7741), .dout(n20415));
  jand g20234(.dina(n19537), .dinb(n7613), .dout(n20416));
  jand g20235(.dina(n19539), .dinb(n6934), .dout(n20417));
  jor  g20236(.dina(n20417), .dinb(n20416), .dout(n20418));
  jor  g20237(.dina(n20418), .dinb(n20415), .dout(n20419));
  jor  g20238(.dina(n20419), .dinb(n20414), .dout(n20420));
  jxor g20239(.dina(n20420), .dinb(n5292), .dout(n20421));
  jor  g20240(.dina(n20421), .dinb(n20412), .dout(n20422));
  jxor g20241(.dina(n20317), .dinb(n20316), .dout(n20423));
  jnot g20242(.din(n20423), .dout(n20424));
  jand g20243(.dina(n20387), .dinb(n6936), .dout(n20425));
  jand g20244(.dina(n19537), .dinb(n7741), .dout(n20426));
  jand g20245(.dina(n19539), .dinb(n7613), .dout(n20427));
  jand g20246(.dina(n19541), .dinb(n6934), .dout(n20428));
  jor  g20247(.dina(n20428), .dinb(n20427), .dout(n20429));
  jor  g20248(.dina(n20429), .dinb(n20426), .dout(n20430));
  jor  g20249(.dina(n20430), .dinb(n20425), .dout(n20431));
  jxor g20250(.dina(n20431), .dinb(n5292), .dout(n20432));
  jor  g20251(.dina(n20432), .dinb(n20424), .dout(n20433));
  jxor g20252(.dina(n20314), .dinb(n20313), .dout(n20434));
  jnot g20253(.din(n20434), .dout(n20435));
  jand g20254(.dina(n20131), .dinb(n6936), .dout(n20436));
  jand g20255(.dina(n19539), .dinb(n7741), .dout(n20437));
  jand g20256(.dina(n19541), .dinb(n7613), .dout(n20438));
  jand g20257(.dina(n19543), .dinb(n6934), .dout(n20439));
  jor  g20258(.dina(n20439), .dinb(n20438), .dout(n20440));
  jor  g20259(.dina(n20440), .dinb(n20437), .dout(n20441));
  jor  g20260(.dina(n20441), .dinb(n20436), .dout(n20442));
  jxor g20261(.dina(n20442), .dinb(n5292), .dout(n20443));
  jor  g20262(.dina(n20443), .dinb(n20435), .dout(n20444));
  jand g20263(.dina(n20141), .dinb(n6936), .dout(n20445));
  jand g20264(.dina(n19541), .dinb(n7741), .dout(n20446));
  jand g20265(.dina(n19543), .dinb(n7613), .dout(n20447));
  jand g20266(.dina(n19545), .dinb(n6934), .dout(n20448));
  jor  g20267(.dina(n20448), .dinb(n20447), .dout(n20449));
  jor  g20268(.dina(n20449), .dinb(n20446), .dout(n20450));
  jor  g20269(.dina(n20450), .dinb(n20445), .dout(n20451));
  jxor g20270(.dina(n20451), .dinb(n5292), .dout(n20452));
  jnot g20271(.din(n20452), .dout(n20453));
  jxor g20272(.dina(n20309), .dinb(n20308), .dout(n20454));
  jand g20273(.dina(n20454), .dinb(n20453), .dout(n20455));
  jand g20274(.dina(n20153), .dinb(n6936), .dout(n20456));
  jand g20275(.dina(n19543), .dinb(n7741), .dout(n20457));
  jand g20276(.dina(n19545), .dinb(n7613), .dout(n20458));
  jand g20277(.dina(n19548), .dinb(n6934), .dout(n20459));
  jor  g20278(.dina(n20459), .dinb(n20458), .dout(n20460));
  jor  g20279(.dina(n20460), .dinb(n20457), .dout(n20461));
  jor  g20280(.dina(n20461), .dinb(n20456), .dout(n20462));
  jxor g20281(.dina(n20462), .dinb(n5292), .dout(n20463));
  jnot g20282(.din(n20463), .dout(n20464));
  jxor g20283(.dina(n20304), .dinb(n20303), .dout(n20465));
  jand g20284(.dina(n20465), .dinb(n20464), .dout(n20466));
  jand g20285(.dina(n20079), .dinb(n6936), .dout(n20467));
  jand g20286(.dina(n19545), .dinb(n7741), .dout(n20468));
  jand g20287(.dina(n19548), .dinb(n7613), .dout(n20469));
  jand g20288(.dina(n19551), .dinb(n6934), .dout(n20470));
  jor  g20289(.dina(n20470), .dinb(n20469), .dout(n20471));
  jor  g20290(.dina(n20471), .dinb(n20468), .dout(n20472));
  jor  g20291(.dina(n20472), .dinb(n20467), .dout(n20473));
  jxor g20292(.dina(n20473), .dinb(n5292), .dout(n20474));
  jnot g20293(.din(n20474), .dout(n20475));
  jxor g20294(.dina(n20299), .dinb(n20298), .dout(n20476));
  jand g20295(.dina(n20476), .dinb(n20475), .dout(n20477));
  jxor g20296(.dina(n20296), .dinb(n20295), .dout(n20478));
  jnot g20297(.din(n20478), .dout(n20479));
  jor  g20298(.dina(n19940), .dinb(n6937), .dout(n20480));
  jor  g20299(.dina(n19547), .dinb(n7740), .dout(n20481));
  jor  g20300(.dina(n19550), .dinb(n7614), .dout(n20482));
  jor  g20301(.dina(n19553), .dinb(n6935), .dout(n20483));
  jand g20302(.dina(n20483), .dinb(n20482), .dout(n20484));
  jand g20303(.dina(n20484), .dinb(n20481), .dout(n20485));
  jand g20304(.dina(n20485), .dinb(n20480), .dout(n20486));
  jxor g20305(.dina(n20486), .dinb(\a[14] ), .dout(n20487));
  jor  g20306(.dina(n20487), .dinb(n20479), .dout(n20488));
  jxor g20307(.dina(n20293), .dinb(n20292), .dout(n20489));
  jnot g20308(.din(n20489), .dout(n20490));
  jor  g20309(.dina(n19952), .dinb(n6937), .dout(n20491));
  jor  g20310(.dina(n19550), .dinb(n7740), .dout(n20492));
  jor  g20311(.dina(n19553), .dinb(n7614), .dout(n20493));
  jor  g20312(.dina(n19558), .dinb(n6935), .dout(n20494));
  jand g20313(.dina(n20494), .dinb(n20493), .dout(n20495));
  jand g20314(.dina(n20495), .dinb(n20492), .dout(n20496));
  jand g20315(.dina(n20496), .dinb(n20491), .dout(n20497));
  jxor g20316(.dina(n20497), .dinb(\a[14] ), .dout(n20498));
  jor  g20317(.dina(n20498), .dinb(n20490), .dout(n20499));
  jxor g20318(.dina(n20290), .dinb(n20289), .dout(n20500));
  jnot g20319(.din(n20500), .dout(n20501));
  jor  g20320(.dina(n19964), .dinb(n6937), .dout(n20502));
  jor  g20321(.dina(n19553), .dinb(n7740), .dout(n20503));
  jor  g20322(.dina(n19558), .dinb(n7614), .dout(n20504));
  jor  g20323(.dina(n19562), .dinb(n6935), .dout(n20505));
  jand g20324(.dina(n20505), .dinb(n20504), .dout(n20506));
  jand g20325(.dina(n20506), .dinb(n20503), .dout(n20507));
  jand g20326(.dina(n20507), .dinb(n20502), .dout(n20508));
  jxor g20327(.dina(n20508), .dinb(\a[14] ), .dout(n20509));
  jor  g20328(.dina(n20509), .dinb(n20501), .dout(n20510));
  jor  g20329(.dina(n19906), .dinb(n6937), .dout(n20511));
  jor  g20330(.dina(n19558), .dinb(n7740), .dout(n20512));
  jor  g20331(.dina(n19562), .dinb(n7614), .dout(n20513));
  jor  g20332(.dina(n19564), .dinb(n6935), .dout(n20514));
  jand g20333(.dina(n20514), .dinb(n20513), .dout(n20515));
  jand g20334(.dina(n20515), .dinb(n20512), .dout(n20516));
  jand g20335(.dina(n20516), .dinb(n20511), .dout(n20517));
  jxor g20336(.dina(n20517), .dinb(\a[14] ), .dout(n20518));
  jnot g20337(.din(n20518), .dout(n20519));
  jxor g20338(.dina(n20287), .dinb(n20286), .dout(n20520));
  jand g20339(.dina(n20520), .dinb(n20519), .dout(n20521));
  jor  g20340(.dina(n19790), .dinb(n6937), .dout(n20522));
  jor  g20341(.dina(n19562), .dinb(n7740), .dout(n20523));
  jor  g20342(.dina(n19564), .dinb(n7614), .dout(n20524));
  jor  g20343(.dina(n19566), .dinb(n6935), .dout(n20525));
  jand g20344(.dina(n20525), .dinb(n20524), .dout(n20526));
  jand g20345(.dina(n20526), .dinb(n20523), .dout(n20527));
  jand g20346(.dina(n20527), .dinb(n20522), .dout(n20528));
  jxor g20347(.dina(n20528), .dinb(\a[14] ), .dout(n20529));
  jnot g20348(.din(n20529), .dout(n20530));
  jxor g20349(.dina(n20284), .dinb(n20283), .dout(n20531));
  jand g20350(.dina(n20531), .dinb(n20530), .dout(n20532));
  jor  g20351(.dina(n19839), .dinb(n6937), .dout(n20533));
  jor  g20352(.dina(n19564), .dinb(n7740), .dout(n20534));
  jor  g20353(.dina(n19566), .dinb(n7614), .dout(n20535));
  jor  g20354(.dina(n19568), .dinb(n6935), .dout(n20536));
  jand g20355(.dina(n20536), .dinb(n20535), .dout(n20537));
  jand g20356(.dina(n20537), .dinb(n20534), .dout(n20538));
  jand g20357(.dina(n20538), .dinb(n20533), .dout(n20539));
  jxor g20358(.dina(n20539), .dinb(\a[14] ), .dout(n20540));
  jnot g20359(.din(n20540), .dout(n20541));
  jor  g20360(.dina(n20264), .dinb(n5064), .dout(n20542));
  jxor g20361(.dina(n20542), .dinb(n20272), .dout(n20543));
  jand g20362(.dina(n20543), .dinb(n20541), .dout(n20544));
  jor  g20363(.dina(n19852), .dinb(n6937), .dout(n20545));
  jor  g20364(.dina(n19566), .dinb(n7740), .dout(n20546));
  jor  g20365(.dina(n19568), .dinb(n7614), .dout(n20547));
  jor  g20366(.dina(n19570), .dinb(n6935), .dout(n20548));
  jand g20367(.dina(n20548), .dinb(n20547), .dout(n20549));
  jand g20368(.dina(n20549), .dinb(n20546), .dout(n20550));
  jand g20369(.dina(n20550), .dinb(n20545), .dout(n20551));
  jxor g20370(.dina(n20551), .dinb(\a[14] ), .dout(n20552));
  jnot g20371(.din(n20552), .dout(n20553));
  jand g20372(.dina(n20261), .dinb(\a[17] ), .dout(n20554));
  jxor g20373(.dina(n20554), .dinb(n20259), .dout(n20555));
  jand g20374(.dina(n20555), .dinb(n20553), .dout(n20556));
  jand g20375(.dina(n19813), .dinb(n6936), .dout(n20557));
  jand g20376(.dina(n19576), .dinb(n7613), .dout(n20558));
  jand g20377(.dina(n19574), .dinb(n7741), .dout(n20559));
  jor  g20378(.dina(n20559), .dinb(n20558), .dout(n20560));
  jor  g20379(.dina(n20560), .dinb(n20557), .dout(n20561));
  jnot g20380(.din(n20561), .dout(n20562));
  jand g20381(.dina(n19576), .dinb(n6928), .dout(n20563));
  jnot g20382(.din(n20563), .dout(n20564));
  jand g20383(.dina(n20564), .dinb(\a[14] ), .dout(n20565));
  jand g20384(.dina(n20565), .dinb(n20562), .dout(n20566));
  jand g20385(.dina(n19826), .dinb(n6936), .dout(n20567));
  jand g20386(.dina(n19572), .dinb(n7741), .dout(n20568));
  jand g20387(.dina(n19574), .dinb(n7613), .dout(n20569));
  jand g20388(.dina(n19576), .dinb(n6934), .dout(n20570));
  jor  g20389(.dina(n20570), .dinb(n20569), .dout(n20571));
  jor  g20390(.dina(n20571), .dinb(n20568), .dout(n20572));
  jor  g20391(.dina(n20572), .dinb(n20567), .dout(n20573));
  jnot g20392(.din(n20573), .dout(n20574));
  jand g20393(.dina(n20574), .dinb(n20566), .dout(n20575));
  jand g20394(.dina(n20575), .dinb(n20261), .dout(n20576));
  jor  g20395(.dina(n19801), .dinb(n6937), .dout(n20577));
  jor  g20396(.dina(n19568), .dinb(n7740), .dout(n20578));
  jor  g20397(.dina(n19570), .dinb(n7614), .dout(n20579));
  jor  g20398(.dina(n19575), .dinb(n6935), .dout(n20580));
  jand g20399(.dina(n20580), .dinb(n20579), .dout(n20581));
  jand g20400(.dina(n20581), .dinb(n20578), .dout(n20582));
  jand g20401(.dina(n20582), .dinb(n20577), .dout(n20583));
  jxor g20402(.dina(n20583), .dinb(\a[14] ), .dout(n20584));
  jnot g20403(.din(n20584), .dout(n20585));
  jxor g20404(.dina(n20575), .dinb(n20261), .dout(n20586));
  jand g20405(.dina(n20586), .dinb(n20585), .dout(n20587));
  jor  g20406(.dina(n20587), .dinb(n20576), .dout(n20588));
  jxor g20407(.dina(n20555), .dinb(n20553), .dout(n20589));
  jand g20408(.dina(n20589), .dinb(n20588), .dout(n20590));
  jor  g20409(.dina(n20590), .dinb(n20556), .dout(n20591));
  jxor g20410(.dina(n20543), .dinb(n20541), .dout(n20592));
  jand g20411(.dina(n20592), .dinb(n20591), .dout(n20593));
  jor  g20412(.dina(n20593), .dinb(n20544), .dout(n20594));
  jxor g20413(.dina(n20531), .dinb(n20530), .dout(n20595));
  jand g20414(.dina(n20595), .dinb(n20594), .dout(n20596));
  jor  g20415(.dina(n20596), .dinb(n20532), .dout(n20597));
  jxor g20416(.dina(n20520), .dinb(n20519), .dout(n20598));
  jand g20417(.dina(n20598), .dinb(n20597), .dout(n20599));
  jor  g20418(.dina(n20599), .dinb(n20521), .dout(n20600));
  jxor g20419(.dina(n20509), .dinb(n20501), .dout(n20601));
  jand g20420(.dina(n20601), .dinb(n20600), .dout(n20602));
  jnot g20421(.din(n20602), .dout(n20603));
  jand g20422(.dina(n20603), .dinb(n20510), .dout(n20604));
  jnot g20423(.din(n20604), .dout(n20605));
  jxor g20424(.dina(n20498), .dinb(n20490), .dout(n20606));
  jand g20425(.dina(n20606), .dinb(n20605), .dout(n20607));
  jnot g20426(.din(n20607), .dout(n20608));
  jand g20427(.dina(n20608), .dinb(n20499), .dout(n20609));
  jnot g20428(.din(n20609), .dout(n20610));
  jxor g20429(.dina(n20487), .dinb(n20479), .dout(n20611));
  jand g20430(.dina(n20611), .dinb(n20610), .dout(n20612));
  jnot g20431(.din(n20612), .dout(n20613));
  jand g20432(.dina(n20613), .dinb(n20488), .dout(n20614));
  jnot g20433(.din(n20614), .dout(n20615));
  jxor g20434(.dina(n20476), .dinb(n20475), .dout(n20616));
  jand g20435(.dina(n20616), .dinb(n20615), .dout(n20617));
  jor  g20436(.dina(n20617), .dinb(n20477), .dout(n20618));
  jxor g20437(.dina(n20465), .dinb(n20464), .dout(n20619));
  jand g20438(.dina(n20619), .dinb(n20618), .dout(n20620));
  jor  g20439(.dina(n20620), .dinb(n20466), .dout(n20621));
  jxor g20440(.dina(n20454), .dinb(n20453), .dout(n20622));
  jand g20441(.dina(n20622), .dinb(n20621), .dout(n20623));
  jor  g20442(.dina(n20623), .dinb(n20455), .dout(n20624));
  jxor g20443(.dina(n20443), .dinb(n20435), .dout(n20625));
  jand g20444(.dina(n20625), .dinb(n20624), .dout(n20626));
  jnot g20445(.din(n20626), .dout(n20627));
  jand g20446(.dina(n20627), .dinb(n20444), .dout(n20628));
  jnot g20447(.din(n20628), .dout(n20629));
  jxor g20448(.dina(n20432), .dinb(n20424), .dout(n20630));
  jand g20449(.dina(n20630), .dinb(n20629), .dout(n20631));
  jnot g20450(.din(n20631), .dout(n20632));
  jand g20451(.dina(n20632), .dinb(n20433), .dout(n20633));
  jnot g20452(.din(n20633), .dout(n20634));
  jxor g20453(.dina(n20421), .dinb(n20412), .dout(n20635));
  jand g20454(.dina(n20635), .dinb(n20634), .dout(n20636));
  jnot g20455(.din(n20636), .dout(n20637));
  jand g20456(.dina(n20637), .dinb(n20422), .dout(n20638));
  jnot g20457(.din(n20638), .dout(n20639));
  jxor g20458(.dina(n20409), .dinb(n20408), .dout(n20640));
  jand g20459(.dina(n20640), .dinb(n20639), .dout(n20641));
  jor  g20460(.dina(n20641), .dinb(n20410), .dout(n20642));
  jxor g20461(.dina(n20397), .dinb(n19789), .dout(n20643));
  jand g20462(.dina(n20643), .dinb(n20642), .dout(n20644));
  jor  g20463(.dina(n20644), .dinb(n20398), .dout(n20645));
  jor  g20464(.dina(n20395), .dinb(n20386), .dout(n20646));
  jand g20465(.dina(n20396), .dinb(n20327), .dout(n20647));
  jnot g20466(.din(n20647), .dout(n20648));
  jand g20467(.dina(n20648), .dinb(n20646), .dout(n20649));
  jnot g20468(.din(n20649), .dout(n20650));
  jand g20469(.dina(n20413), .dinb(n6340), .dout(n20651));
  jand g20470(.dina(n19535), .dinb(n6798), .dout(n20652));
  jand g20471(.dina(n19537), .dinb(n6556), .dout(n20653));
  jand g20472(.dina(n19539), .dinb(n6338), .dout(n20654));
  jor  g20473(.dina(n20654), .dinb(n20653), .dout(n20655));
  jor  g20474(.dina(n20655), .dinb(n20652), .dout(n20656));
  jor  g20475(.dina(n20656), .dinb(n20651), .dout(n20657));
  jxor g20476(.dina(n20657), .dinb(n5064), .dout(n20658));
  jnot g20477(.din(n20658), .dout(n20659));
  jand g20478(.dina(n20383), .dinb(n20339), .dout(n20660));
  jand g20479(.dina(n20384), .dinb(n20330), .dout(n20661));
  jor  g20480(.dina(n20661), .dinb(n20660), .dout(n20662));
  jor  g20481(.dina(n20381), .dinb(n20373), .dout(n20663));
  jand g20482(.dina(n20382), .dinb(n20344), .dout(n20664));
  jnot g20483(.din(n20664), .dout(n20665));
  jand g20484(.dina(n20665), .dinb(n20663), .dout(n20666));
  jnot g20485(.din(n20666), .dout(n20667));
  jor  g20486(.dina(n19940), .dinb(n5366), .dout(n20668));
  jor  g20487(.dina(n19547), .dinb(n5499), .dout(n20669));
  jor  g20488(.dina(n19550), .dinb(n5425), .dout(n20670));
  jor  g20489(.dina(n19553), .dinb(n5364), .dout(n20671));
  jand g20490(.dina(n20671), .dinb(n20670), .dout(n20672));
  jand g20491(.dina(n20672), .dinb(n20669), .dout(n20673));
  jand g20492(.dina(n20673), .dinb(n20668), .dout(n20674));
  jxor g20493(.dina(n20674), .dinb(\a[23] ), .dout(n20675));
  jnot g20494(.din(n20675), .dout(n20676));
  jand g20495(.dina(n20370), .dinb(n20356), .dout(n20677));
  jand g20496(.dina(n20371), .dinb(n20347), .dout(n20678));
  jor  g20497(.dina(n20678), .dinb(n20677), .dout(n20679));
  jor  g20498(.dina(n19906), .dinb(n4747), .dout(n20680));
  jor  g20499(.dina(n19558), .dinb(n4959), .dout(n20681));
  jor  g20500(.dina(n19562), .dinb(n4919), .dout(n20682));
  jor  g20501(.dina(n19564), .dinb(n4746), .dout(n20683));
  jand g20502(.dina(n20683), .dinb(n20682), .dout(n20684));
  jand g20503(.dina(n20684), .dinb(n20681), .dout(n20685));
  jand g20504(.dina(n20685), .dinb(n20680), .dout(n20686));
  jxor g20505(.dina(n20686), .dinb(\a[26] ), .dout(n20687));
  jnot g20506(.din(n20687), .dout(n20688));
  jand g20507(.dina(n20368), .dinb(n20367), .dout(n20689));
  jand g20508(.dina(n20369), .dinb(n20365), .dout(n20690));
  jor  g20509(.dina(n20690), .dinb(n20689), .dout(n20691));
  jor  g20510(.dina(n19852), .dinb(n4724), .dout(n20692));
  jor  g20511(.dina(n19566), .dinb(n4905), .dout(n20693));
  jor  g20512(.dina(n19568), .dinb(n4735), .dout(n20694));
  jor  g20513(.dina(n19570), .dinb(n4733), .dout(n20695));
  jand g20514(.dina(n20695), .dinb(n20694), .dout(n20696));
  jand g20515(.dina(n20696), .dinb(n20693), .dout(n20697));
  jand g20516(.dina(n20697), .dinb(n20692), .dout(n20698));
  jxor g20517(.dina(n20698), .dinb(\a[29] ), .dout(n20699));
  jnot g20518(.din(n20699), .dout(n20700));
  jand g20519(.dina(n1785), .dinb(n1383), .dout(n20701));
  jand g20520(.dina(n20701), .dinb(n2315), .dout(n20702));
  jand g20521(.dina(n574), .dinb(n252), .dout(n20703));
  jand g20522(.dina(n492), .dinb(n371), .dout(n20704));
  jand g20523(.dina(n20704), .dinb(n20703), .dout(n20705));
  jand g20524(.dina(n1275), .dinb(n1137), .dout(n20706));
  jand g20525(.dina(n20706), .dinb(n20705), .dout(n20707));
  jand g20526(.dina(n20707), .dinb(n1151), .dout(n20708));
  jand g20527(.dina(n20708), .dinb(n20702), .dout(n20709));
  jand g20528(.dina(n392), .dinb(n340), .dout(n20710));
  jand g20529(.dina(n20710), .dinb(n1082), .dout(n20711));
  jand g20530(.dina(n868), .dinb(n93), .dout(n20712));
  jand g20531(.dina(n20712), .dinb(n20711), .dout(n20713));
  jand g20532(.dina(n826), .dinb(n805), .dout(n20714));
  jand g20533(.dina(n20714), .dinb(n346), .dout(n20715));
  jand g20534(.dina(n20715), .dinb(n2946), .dout(n20716));
  jand g20535(.dina(n20716), .dinb(n20713), .dout(n20717));
  jand g20536(.dina(n2053), .dinb(n2963), .dout(n20718));
  jand g20537(.dina(n1986), .dinb(n1249), .dout(n20719));
  jand g20538(.dina(n20719), .dinb(n20718), .dout(n20720));
  jand g20539(.dina(n20720), .dinb(n14407), .dout(n20721));
  jand g20540(.dina(n20721), .dinb(n1926), .dout(n20722));
  jand g20541(.dina(n20722), .dinb(n20717), .dout(n20723));
  jand g20542(.dina(n20723), .dinb(n20709), .dout(n20724));
  jand g20543(.dina(n4576), .dinb(n3591), .dout(n20725));
  jand g20544(.dina(n20725), .dinb(n4998), .dout(n20726));
  jand g20545(.dina(n4211), .dinb(n4004), .dout(n20727));
  jand g20546(.dina(n1711), .dinb(n563), .dout(n20728));
  jand g20547(.dina(n20728), .dinb(n20727), .dout(n20729));
  jand g20548(.dina(n1615), .dinb(n365), .dout(n20730));
  jand g20549(.dina(n860), .dinb(n423), .dout(n20731));
  jand g20550(.dina(n20731), .dinb(n20730), .dout(n20732));
  jand g20551(.dina(n1487), .dinb(n1160), .dout(n20733));
  jand g20552(.dina(n20733), .dinb(n20732), .dout(n20734));
  jand g20553(.dina(n20734), .dinb(n20729), .dout(n20735));
  jand g20554(.dina(n20735), .dinb(n12588), .dout(n20736));
  jand g20555(.dina(n20736), .dinb(n20726), .dout(n20737));
  jand g20556(.dina(n20737), .dinb(n14337), .dout(n20738));
  jand g20557(.dina(n20738), .dinb(n20724), .dout(n20739));
  jnot g20558(.din(n20739), .dout(n20740));
  jand g20559(.dina(n19813), .dinb(n732), .dout(n20741));
  jand g20560(.dina(n19574), .dinb(n3855), .dout(n20742));
  jand g20561(.dina(n19576), .dinb(n3858), .dout(n20743));
  jor  g20562(.dina(n20743), .dinb(n20742), .dout(n20744));
  jor  g20563(.dina(n20744), .dinb(n20741), .dout(n20745));
  jxor g20564(.dina(n20745), .dinb(n20740), .dout(n20746));
  jxor g20565(.dina(n20746), .dinb(n20700), .dout(n20747));
  jxor g20566(.dina(n20747), .dinb(n20691), .dout(n20748));
  jxor g20567(.dina(n20748), .dinb(n20688), .dout(n20749));
  jxor g20568(.dina(n20749), .dinb(n20679), .dout(n20750));
  jxor g20569(.dina(n20750), .dinb(n20676), .dout(n20751));
  jxor g20570(.dina(n20751), .dinb(n20667), .dout(n20752));
  jnot g20571(.din(n20752), .dout(n20753));
  jand g20572(.dina(n20141), .dinb(n5693), .dout(n20754));
  jand g20573(.dina(n19541), .dinb(n6209), .dout(n20755));
  jand g20574(.dina(n19543), .dinb(n6131), .dout(n20756));
  jand g20575(.dina(n19545), .dinb(n5691), .dout(n20757));
  jor  g20576(.dina(n20757), .dinb(n20756), .dout(n20758));
  jor  g20577(.dina(n20758), .dinb(n20755), .dout(n20759));
  jor  g20578(.dina(n20759), .dinb(n20754), .dout(n20760));
  jxor g20579(.dina(n20760), .dinb(n4247), .dout(n20761));
  jxor g20580(.dina(n20761), .dinb(n20753), .dout(n20762));
  jxor g20581(.dina(n20762), .dinb(n20662), .dout(n20763));
  jxor g20582(.dina(n20763), .dinb(n20659), .dout(n20764));
  jxor g20583(.dina(n20764), .dinb(n20650), .dout(n20765));
  jnot g20584(.din(n20765), .dout(n20766));
  jxor g20585(.dina(n19634), .dinb(n19633), .dout(n20767));
  jand g20586(.dina(n20767), .dinb(n6936), .dout(n20768));
  jand g20587(.dina(n19529), .dinb(n7741), .dout(n20769));
  jand g20588(.dina(n19531), .dinb(n7613), .dout(n20770));
  jand g20589(.dina(n19533), .dinb(n6934), .dout(n20771));
  jor  g20590(.dina(n20771), .dinb(n20770), .dout(n20772));
  jor  g20591(.dina(n20772), .dinb(n20769), .dout(n20773));
  jor  g20592(.dina(n20773), .dinb(n20768), .dout(n20774));
  jxor g20593(.dina(n20774), .dinb(n5292), .dout(n20775));
  jxor g20594(.dina(n20775), .dinb(n20766), .dout(n20776));
  jxor g20595(.dina(n20776), .dinb(n20645), .dout(n20777));
  jand g20596(.dina(n20777), .dinb(n19779), .dout(n20778));
  jxor g20597(.dina(n20643), .dinb(n20642), .dout(n20779));
  jnot g20598(.din(n20779), .dout(n20780));
  jxor g20599(.dina(n19640), .dinb(n19639), .dout(n20781));
  jand g20600(.dina(n20781), .dinb(n7890), .dout(n20782));
  jand g20601(.dina(n19525), .dinb(n8441), .dout(n20783));
  jand g20602(.dina(n19527), .dinb(n8154), .dout(n20784));
  jand g20603(.dina(n19529), .dinb(n7888), .dout(n20785));
  jor  g20604(.dina(n20785), .dinb(n20784), .dout(n20786));
  jor  g20605(.dina(n20786), .dinb(n20783), .dout(n20787));
  jor  g20606(.dina(n20787), .dinb(n20782), .dout(n20788));
  jxor g20607(.dina(n20788), .dinb(n5833), .dout(n20789));
  jor  g20608(.dina(n20789), .dinb(n20780), .dout(n20790));
  jxor g20609(.dina(n20640), .dinb(n20639), .dout(n20791));
  jnot g20610(.din(n20791), .dout(n20792));
  jxor g20611(.dina(n19637), .dinb(n19636), .dout(n20793));
  jand g20612(.dina(n20793), .dinb(n7890), .dout(n20794));
  jand g20613(.dina(n19527), .dinb(n8441), .dout(n20795));
  jand g20614(.dina(n19529), .dinb(n8154), .dout(n20796));
  jand g20615(.dina(n19531), .dinb(n7888), .dout(n20797));
  jor  g20616(.dina(n20797), .dinb(n20796), .dout(n20798));
  jor  g20617(.dina(n20798), .dinb(n20795), .dout(n20799));
  jor  g20618(.dina(n20799), .dinb(n20794), .dout(n20800));
  jxor g20619(.dina(n20800), .dinb(n5833), .dout(n20801));
  jor  g20620(.dina(n20801), .dinb(n20792), .dout(n20802));
  jand g20621(.dina(n20767), .dinb(n7890), .dout(n20803));
  jand g20622(.dina(n19529), .dinb(n8441), .dout(n20804));
  jand g20623(.dina(n19531), .dinb(n8154), .dout(n20805));
  jand g20624(.dina(n19533), .dinb(n7888), .dout(n20806));
  jor  g20625(.dina(n20806), .dinb(n20805), .dout(n20807));
  jor  g20626(.dina(n20807), .dinb(n20804), .dout(n20808));
  jor  g20627(.dina(n20808), .dinb(n20803), .dout(n20809));
  jxor g20628(.dina(n20809), .dinb(n5833), .dout(n20810));
  jnot g20629(.din(n20810), .dout(n20811));
  jxor g20630(.dina(n20635), .dinb(n20634), .dout(n20812));
  jand g20631(.dina(n20812), .dinb(n20811), .dout(n20813));
  jand g20632(.dina(n19780), .dinb(n7890), .dout(n20814));
  jand g20633(.dina(n19531), .dinb(n8441), .dout(n20815));
  jand g20634(.dina(n19533), .dinb(n8154), .dout(n20816));
  jand g20635(.dina(n19535), .dinb(n7888), .dout(n20817));
  jor  g20636(.dina(n20817), .dinb(n20816), .dout(n20818));
  jor  g20637(.dina(n20818), .dinb(n20815), .dout(n20819));
  jor  g20638(.dina(n20819), .dinb(n20814), .dout(n20820));
  jxor g20639(.dina(n20820), .dinb(n5833), .dout(n20821));
  jnot g20640(.din(n20821), .dout(n20822));
  jxor g20641(.dina(n20630), .dinb(n20629), .dout(n20823));
  jand g20642(.dina(n20823), .dinb(n20822), .dout(n20824));
  jand g20643(.dina(n20399), .dinb(n7890), .dout(n20825));
  jand g20644(.dina(n19533), .dinb(n8441), .dout(n20826));
  jand g20645(.dina(n19535), .dinb(n8154), .dout(n20827));
  jand g20646(.dina(n19537), .dinb(n7888), .dout(n20828));
  jor  g20647(.dina(n20828), .dinb(n20827), .dout(n20829));
  jor  g20648(.dina(n20829), .dinb(n20826), .dout(n20830));
  jor  g20649(.dina(n20830), .dinb(n20825), .dout(n20831));
  jxor g20650(.dina(n20831), .dinb(n5833), .dout(n20832));
  jnot g20651(.din(n20832), .dout(n20833));
  jxor g20652(.dina(n20625), .dinb(n20624), .dout(n20834));
  jand g20653(.dina(n20834), .dinb(n20833), .dout(n20835));
  jxor g20654(.dina(n20622), .dinb(n20621), .dout(n20836));
  jnot g20655(.din(n20836), .dout(n20837));
  jand g20656(.dina(n20413), .dinb(n7890), .dout(n20838));
  jand g20657(.dina(n19535), .dinb(n8441), .dout(n20839));
  jand g20658(.dina(n19537), .dinb(n8154), .dout(n20840));
  jand g20659(.dina(n19539), .dinb(n7888), .dout(n20841));
  jor  g20660(.dina(n20841), .dinb(n20840), .dout(n20842));
  jor  g20661(.dina(n20842), .dinb(n20839), .dout(n20843));
  jor  g20662(.dina(n20843), .dinb(n20838), .dout(n20844));
  jxor g20663(.dina(n20844), .dinb(n5833), .dout(n20845));
  jor  g20664(.dina(n20845), .dinb(n20837), .dout(n20846));
  jxor g20665(.dina(n20619), .dinb(n20618), .dout(n20847));
  jnot g20666(.din(n20847), .dout(n20848));
  jand g20667(.dina(n20387), .dinb(n7890), .dout(n20849));
  jand g20668(.dina(n19537), .dinb(n8441), .dout(n20850));
  jand g20669(.dina(n19539), .dinb(n8154), .dout(n20851));
  jand g20670(.dina(n19541), .dinb(n7888), .dout(n20852));
  jor  g20671(.dina(n20852), .dinb(n20851), .dout(n20853));
  jor  g20672(.dina(n20853), .dinb(n20850), .dout(n20854));
  jor  g20673(.dina(n20854), .dinb(n20849), .dout(n20855));
  jxor g20674(.dina(n20855), .dinb(n5833), .dout(n20856));
  jor  g20675(.dina(n20856), .dinb(n20848), .dout(n20857));
  jxor g20676(.dina(n20616), .dinb(n20615), .dout(n20858));
  jnot g20677(.din(n20858), .dout(n20859));
  jand g20678(.dina(n20131), .dinb(n7890), .dout(n20860));
  jand g20679(.dina(n19539), .dinb(n8441), .dout(n20861));
  jand g20680(.dina(n19541), .dinb(n8154), .dout(n20862));
  jand g20681(.dina(n19543), .dinb(n7888), .dout(n20863));
  jor  g20682(.dina(n20863), .dinb(n20862), .dout(n20864));
  jor  g20683(.dina(n20864), .dinb(n20861), .dout(n20865));
  jor  g20684(.dina(n20865), .dinb(n20860), .dout(n20866));
  jxor g20685(.dina(n20866), .dinb(n5833), .dout(n20867));
  jor  g20686(.dina(n20867), .dinb(n20859), .dout(n20868));
  jand g20687(.dina(n20141), .dinb(n7890), .dout(n20869));
  jand g20688(.dina(n19541), .dinb(n8441), .dout(n20870));
  jand g20689(.dina(n19543), .dinb(n8154), .dout(n20871));
  jand g20690(.dina(n19545), .dinb(n7888), .dout(n20872));
  jor  g20691(.dina(n20872), .dinb(n20871), .dout(n20873));
  jor  g20692(.dina(n20873), .dinb(n20870), .dout(n20874));
  jor  g20693(.dina(n20874), .dinb(n20869), .dout(n20875));
  jxor g20694(.dina(n20875), .dinb(n5833), .dout(n20876));
  jnot g20695(.din(n20876), .dout(n20877));
  jxor g20696(.dina(n20611), .dinb(n20610), .dout(n20878));
  jand g20697(.dina(n20878), .dinb(n20877), .dout(n20879));
  jand g20698(.dina(n20153), .dinb(n7890), .dout(n20880));
  jand g20699(.dina(n19543), .dinb(n8441), .dout(n20881));
  jand g20700(.dina(n19545), .dinb(n8154), .dout(n20882));
  jand g20701(.dina(n19548), .dinb(n7888), .dout(n20883));
  jor  g20702(.dina(n20883), .dinb(n20882), .dout(n20884));
  jor  g20703(.dina(n20884), .dinb(n20881), .dout(n20885));
  jor  g20704(.dina(n20885), .dinb(n20880), .dout(n20886));
  jxor g20705(.dina(n20886), .dinb(n5833), .dout(n20887));
  jnot g20706(.din(n20887), .dout(n20888));
  jxor g20707(.dina(n20606), .dinb(n20605), .dout(n20889));
  jand g20708(.dina(n20889), .dinb(n20888), .dout(n20890));
  jand g20709(.dina(n20079), .dinb(n7890), .dout(n20891));
  jand g20710(.dina(n19545), .dinb(n8441), .dout(n20892));
  jand g20711(.dina(n19548), .dinb(n8154), .dout(n20893));
  jand g20712(.dina(n19551), .dinb(n7888), .dout(n20894));
  jor  g20713(.dina(n20894), .dinb(n20893), .dout(n20895));
  jor  g20714(.dina(n20895), .dinb(n20892), .dout(n20896));
  jor  g20715(.dina(n20896), .dinb(n20891), .dout(n20897));
  jxor g20716(.dina(n20897), .dinb(n5833), .dout(n20898));
  jnot g20717(.din(n20898), .dout(n20899));
  jxor g20718(.dina(n20601), .dinb(n20600), .dout(n20900));
  jand g20719(.dina(n20900), .dinb(n20899), .dout(n20901));
  jxor g20720(.dina(n20598), .dinb(n20597), .dout(n20902));
  jnot g20721(.din(n20902), .dout(n20903));
  jor  g20722(.dina(n19940), .dinb(n7891), .dout(n20904));
  jor  g20723(.dina(n19547), .dinb(n8440), .dout(n20905));
  jor  g20724(.dina(n19550), .dinb(n8155), .dout(n20906));
  jor  g20725(.dina(n19553), .dinb(n7889), .dout(n20907));
  jand g20726(.dina(n20907), .dinb(n20906), .dout(n20908));
  jand g20727(.dina(n20908), .dinb(n20905), .dout(n20909));
  jand g20728(.dina(n20909), .dinb(n20904), .dout(n20910));
  jxor g20729(.dina(n20910), .dinb(\a[11] ), .dout(n20911));
  jor  g20730(.dina(n20911), .dinb(n20903), .dout(n20912));
  jxor g20731(.dina(n20595), .dinb(n20594), .dout(n20913));
  jnot g20732(.din(n20913), .dout(n20914));
  jor  g20733(.dina(n19952), .dinb(n7891), .dout(n20915));
  jor  g20734(.dina(n19550), .dinb(n8440), .dout(n20916));
  jor  g20735(.dina(n19553), .dinb(n8155), .dout(n20917));
  jor  g20736(.dina(n19558), .dinb(n7889), .dout(n20918));
  jand g20737(.dina(n20918), .dinb(n20917), .dout(n20919));
  jand g20738(.dina(n20919), .dinb(n20916), .dout(n20920));
  jand g20739(.dina(n20920), .dinb(n20915), .dout(n20921));
  jxor g20740(.dina(n20921), .dinb(\a[11] ), .dout(n20922));
  jor  g20741(.dina(n20922), .dinb(n20914), .dout(n20923));
  jxor g20742(.dina(n20592), .dinb(n20591), .dout(n20924));
  jnot g20743(.din(n20924), .dout(n20925));
  jor  g20744(.dina(n19964), .dinb(n7891), .dout(n20926));
  jor  g20745(.dina(n19553), .dinb(n8440), .dout(n20927));
  jor  g20746(.dina(n19558), .dinb(n8155), .dout(n20928));
  jor  g20747(.dina(n19562), .dinb(n7889), .dout(n20929));
  jand g20748(.dina(n20929), .dinb(n20928), .dout(n20930));
  jand g20749(.dina(n20930), .dinb(n20927), .dout(n20931));
  jand g20750(.dina(n20931), .dinb(n20926), .dout(n20932));
  jxor g20751(.dina(n20932), .dinb(\a[11] ), .dout(n20933));
  jor  g20752(.dina(n20933), .dinb(n20925), .dout(n20934));
  jor  g20753(.dina(n19906), .dinb(n7891), .dout(n20935));
  jor  g20754(.dina(n19558), .dinb(n8440), .dout(n20936));
  jor  g20755(.dina(n19562), .dinb(n8155), .dout(n20937));
  jor  g20756(.dina(n19564), .dinb(n7889), .dout(n20938));
  jand g20757(.dina(n20938), .dinb(n20937), .dout(n20939));
  jand g20758(.dina(n20939), .dinb(n20936), .dout(n20940));
  jand g20759(.dina(n20940), .dinb(n20935), .dout(n20941));
  jxor g20760(.dina(n20941), .dinb(\a[11] ), .dout(n20942));
  jnot g20761(.din(n20942), .dout(n20943));
  jxor g20762(.dina(n20589), .dinb(n20588), .dout(n20944));
  jand g20763(.dina(n20944), .dinb(n20943), .dout(n20945));
  jor  g20764(.dina(n19790), .dinb(n7891), .dout(n20946));
  jor  g20765(.dina(n19562), .dinb(n8440), .dout(n20947));
  jor  g20766(.dina(n19564), .dinb(n8155), .dout(n20948));
  jor  g20767(.dina(n19566), .dinb(n7889), .dout(n20949));
  jand g20768(.dina(n20949), .dinb(n20948), .dout(n20950));
  jand g20769(.dina(n20950), .dinb(n20947), .dout(n20951));
  jand g20770(.dina(n20951), .dinb(n20946), .dout(n20952));
  jxor g20771(.dina(n20952), .dinb(\a[11] ), .dout(n20953));
  jnot g20772(.din(n20953), .dout(n20954));
  jxor g20773(.dina(n20586), .dinb(n20585), .dout(n20955));
  jand g20774(.dina(n20955), .dinb(n20954), .dout(n20956));
  jor  g20775(.dina(n19839), .dinb(n7891), .dout(n20957));
  jor  g20776(.dina(n19564), .dinb(n8440), .dout(n20958));
  jor  g20777(.dina(n19566), .dinb(n8155), .dout(n20959));
  jor  g20778(.dina(n19568), .dinb(n7889), .dout(n20960));
  jand g20779(.dina(n20960), .dinb(n20959), .dout(n20961));
  jand g20780(.dina(n20961), .dinb(n20958), .dout(n20962));
  jand g20781(.dina(n20962), .dinb(n20957), .dout(n20963));
  jxor g20782(.dina(n20963), .dinb(\a[11] ), .dout(n20964));
  jnot g20783(.din(n20964), .dout(n20965));
  jor  g20784(.dina(n20566), .dinb(n5292), .dout(n20966));
  jxor g20785(.dina(n20966), .dinb(n20574), .dout(n20967));
  jand g20786(.dina(n20967), .dinb(n20965), .dout(n20968));
  jor  g20787(.dina(n19852), .dinb(n7891), .dout(n20969));
  jor  g20788(.dina(n19566), .dinb(n8440), .dout(n20970));
  jor  g20789(.dina(n19568), .dinb(n8155), .dout(n20971));
  jor  g20790(.dina(n19570), .dinb(n7889), .dout(n20972));
  jand g20791(.dina(n20972), .dinb(n20971), .dout(n20973));
  jand g20792(.dina(n20973), .dinb(n20970), .dout(n20974));
  jand g20793(.dina(n20974), .dinb(n20969), .dout(n20975));
  jxor g20794(.dina(n20975), .dinb(\a[11] ), .dout(n20976));
  jnot g20795(.din(n20976), .dout(n20977));
  jand g20796(.dina(n20563), .dinb(\a[14] ), .dout(n20978));
  jxor g20797(.dina(n20978), .dinb(n20561), .dout(n20979));
  jand g20798(.dina(n20979), .dinb(n20977), .dout(n20980));
  jand g20799(.dina(n19813), .dinb(n7890), .dout(n20981));
  jand g20800(.dina(n19576), .dinb(n8154), .dout(n20982));
  jand g20801(.dina(n19574), .dinb(n8441), .dout(n20983));
  jor  g20802(.dina(n20983), .dinb(n20982), .dout(n20984));
  jor  g20803(.dina(n20984), .dinb(n20981), .dout(n20985));
  jnot g20804(.din(n20985), .dout(n20986));
  jand g20805(.dina(n19576), .dinb(n7884), .dout(n20987));
  jnot g20806(.din(n20987), .dout(n20988));
  jand g20807(.dina(n20988), .dinb(\a[11] ), .dout(n20989));
  jand g20808(.dina(n20989), .dinb(n20986), .dout(n20990));
  jand g20809(.dina(n19826), .dinb(n7890), .dout(n20991));
  jand g20810(.dina(n19572), .dinb(n8441), .dout(n20992));
  jand g20811(.dina(n19574), .dinb(n8154), .dout(n20993));
  jand g20812(.dina(n19576), .dinb(n7888), .dout(n20994));
  jor  g20813(.dina(n20994), .dinb(n20993), .dout(n20995));
  jor  g20814(.dina(n20995), .dinb(n20992), .dout(n20996));
  jor  g20815(.dina(n20996), .dinb(n20991), .dout(n20997));
  jnot g20816(.din(n20997), .dout(n20998));
  jand g20817(.dina(n20998), .dinb(n20990), .dout(n20999));
  jand g20818(.dina(n20999), .dinb(n20563), .dout(n21000));
  jor  g20819(.dina(n19801), .dinb(n7891), .dout(n21001));
  jor  g20820(.dina(n19568), .dinb(n8440), .dout(n21002));
  jor  g20821(.dina(n19570), .dinb(n8155), .dout(n21003));
  jor  g20822(.dina(n19575), .dinb(n7889), .dout(n21004));
  jand g20823(.dina(n21004), .dinb(n21003), .dout(n21005));
  jand g20824(.dina(n21005), .dinb(n21002), .dout(n21006));
  jand g20825(.dina(n21006), .dinb(n21001), .dout(n21007));
  jxor g20826(.dina(n21007), .dinb(\a[11] ), .dout(n21008));
  jnot g20827(.din(n21008), .dout(n21009));
  jxor g20828(.dina(n20999), .dinb(n20563), .dout(n21010));
  jand g20829(.dina(n21010), .dinb(n21009), .dout(n21011));
  jor  g20830(.dina(n21011), .dinb(n21000), .dout(n21012));
  jxor g20831(.dina(n20979), .dinb(n20977), .dout(n21013));
  jand g20832(.dina(n21013), .dinb(n21012), .dout(n21014));
  jor  g20833(.dina(n21014), .dinb(n20980), .dout(n21015));
  jxor g20834(.dina(n20967), .dinb(n20965), .dout(n21016));
  jand g20835(.dina(n21016), .dinb(n21015), .dout(n21017));
  jor  g20836(.dina(n21017), .dinb(n20968), .dout(n21018));
  jxor g20837(.dina(n20955), .dinb(n20954), .dout(n21019));
  jand g20838(.dina(n21019), .dinb(n21018), .dout(n21020));
  jor  g20839(.dina(n21020), .dinb(n20956), .dout(n21021));
  jxor g20840(.dina(n20944), .dinb(n20943), .dout(n21022));
  jand g20841(.dina(n21022), .dinb(n21021), .dout(n21023));
  jor  g20842(.dina(n21023), .dinb(n20945), .dout(n21024));
  jxor g20843(.dina(n20933), .dinb(n20925), .dout(n21025));
  jand g20844(.dina(n21025), .dinb(n21024), .dout(n21026));
  jnot g20845(.din(n21026), .dout(n21027));
  jand g20846(.dina(n21027), .dinb(n20934), .dout(n21028));
  jnot g20847(.din(n21028), .dout(n21029));
  jxor g20848(.dina(n20922), .dinb(n20914), .dout(n21030));
  jand g20849(.dina(n21030), .dinb(n21029), .dout(n21031));
  jnot g20850(.din(n21031), .dout(n21032));
  jand g20851(.dina(n21032), .dinb(n20923), .dout(n21033));
  jnot g20852(.din(n21033), .dout(n21034));
  jxor g20853(.dina(n20911), .dinb(n20903), .dout(n21035));
  jand g20854(.dina(n21035), .dinb(n21034), .dout(n21036));
  jnot g20855(.din(n21036), .dout(n21037));
  jand g20856(.dina(n21037), .dinb(n20912), .dout(n21038));
  jnot g20857(.din(n21038), .dout(n21039));
  jxor g20858(.dina(n20900), .dinb(n20899), .dout(n21040));
  jand g20859(.dina(n21040), .dinb(n21039), .dout(n21041));
  jor  g20860(.dina(n21041), .dinb(n20901), .dout(n21042));
  jxor g20861(.dina(n20889), .dinb(n20888), .dout(n21043));
  jand g20862(.dina(n21043), .dinb(n21042), .dout(n21044));
  jor  g20863(.dina(n21044), .dinb(n20890), .dout(n21045));
  jxor g20864(.dina(n20878), .dinb(n20877), .dout(n21046));
  jand g20865(.dina(n21046), .dinb(n21045), .dout(n21047));
  jor  g20866(.dina(n21047), .dinb(n20879), .dout(n21048));
  jxor g20867(.dina(n20867), .dinb(n20859), .dout(n21049));
  jand g20868(.dina(n21049), .dinb(n21048), .dout(n21050));
  jnot g20869(.din(n21050), .dout(n21051));
  jand g20870(.dina(n21051), .dinb(n20868), .dout(n21052));
  jnot g20871(.din(n21052), .dout(n21053));
  jxor g20872(.dina(n20856), .dinb(n20848), .dout(n21054));
  jand g20873(.dina(n21054), .dinb(n21053), .dout(n21055));
  jnot g20874(.din(n21055), .dout(n21056));
  jand g20875(.dina(n21056), .dinb(n20857), .dout(n21057));
  jnot g20876(.din(n21057), .dout(n21058));
  jxor g20877(.dina(n20845), .dinb(n20837), .dout(n21059));
  jand g20878(.dina(n21059), .dinb(n21058), .dout(n21060));
  jnot g20879(.din(n21060), .dout(n21061));
  jand g20880(.dina(n21061), .dinb(n20846), .dout(n21062));
  jnot g20881(.din(n21062), .dout(n21063));
  jxor g20882(.dina(n20834), .dinb(n20833), .dout(n21064));
  jand g20883(.dina(n21064), .dinb(n21063), .dout(n21065));
  jor  g20884(.dina(n21065), .dinb(n20835), .dout(n21066));
  jxor g20885(.dina(n20823), .dinb(n20822), .dout(n21067));
  jand g20886(.dina(n21067), .dinb(n21066), .dout(n21068));
  jor  g20887(.dina(n21068), .dinb(n20824), .dout(n21069));
  jxor g20888(.dina(n20812), .dinb(n20811), .dout(n21070));
  jand g20889(.dina(n21070), .dinb(n21069), .dout(n21071));
  jor  g20890(.dina(n21071), .dinb(n20813), .dout(n21072));
  jxor g20891(.dina(n20801), .dinb(n20792), .dout(n21073));
  jand g20892(.dina(n21073), .dinb(n21072), .dout(n21074));
  jnot g20893(.din(n21074), .dout(n21075));
  jand g20894(.dina(n21075), .dinb(n20802), .dout(n21076));
  jnot g20895(.din(n21076), .dout(n21077));
  jxor g20896(.dina(n20789), .dinb(n20780), .dout(n21078));
  jand g20897(.dina(n21078), .dinb(n21077), .dout(n21079));
  jnot g20898(.din(n21079), .dout(n21080));
  jand g20899(.dina(n21080), .dinb(n20790), .dout(n21081));
  jnot g20900(.din(n21081), .dout(n21082));
  jxor g20901(.dina(n20777), .dinb(n19779), .dout(n21083));
  jand g20902(.dina(n21083), .dinb(n21082), .dout(n21084));
  jor  g20903(.dina(n21084), .dinb(n20778), .dout(n21085));
  jxor g20904(.dina(n19646), .dinb(n19645), .dout(n21086));
  jand g20905(.dina(n21086), .dinb(n7890), .dout(n21087));
  jand g20906(.dina(n19521), .dinb(n8441), .dout(n21088));
  jand g20907(.dina(n19523), .dinb(n8154), .dout(n21089));
  jand g20908(.dina(n19525), .dinb(n7888), .dout(n21090));
  jor  g20909(.dina(n21090), .dinb(n21089), .dout(n21091));
  jor  g20910(.dina(n21091), .dinb(n21088), .dout(n21092));
  jor  g20911(.dina(n21092), .dinb(n21087), .dout(n21093));
  jxor g20912(.dina(n21093), .dinb(n5833), .dout(n21094));
  jnot g20913(.din(n21094), .dout(n21095));
  jor  g20914(.dina(n20775), .dinb(n20766), .dout(n21096));
  jand g20915(.dina(n20776), .dinb(n20645), .dout(n21097));
  jnot g20916(.din(n21097), .dout(n21098));
  jand g20917(.dina(n21098), .dinb(n21096), .dout(n21099));
  jnot g20918(.din(n21099), .dout(n21100));
  jand g20919(.dina(n20763), .dinb(n20659), .dout(n21101));
  jand g20920(.dina(n20764), .dinb(n20650), .dout(n21102));
  jor  g20921(.dina(n21102), .dinb(n21101), .dout(n21103));
  jand g20922(.dina(n20399), .dinb(n6340), .dout(n21104));
  jand g20923(.dina(n19533), .dinb(n6798), .dout(n21105));
  jand g20924(.dina(n19535), .dinb(n6556), .dout(n21106));
  jand g20925(.dina(n19537), .dinb(n6338), .dout(n21107));
  jor  g20926(.dina(n21107), .dinb(n21106), .dout(n21108));
  jor  g20927(.dina(n21108), .dinb(n21105), .dout(n21109));
  jor  g20928(.dina(n21109), .dinb(n21104), .dout(n21110));
  jxor g20929(.dina(n21110), .dinb(n5064), .dout(n21111));
  jnot g20930(.din(n21111), .dout(n21112));
  jor  g20931(.dina(n20761), .dinb(n20753), .dout(n21113));
  jand g20932(.dina(n20762), .dinb(n20662), .dout(n21114));
  jnot g20933(.din(n21114), .dout(n21115));
  jand g20934(.dina(n21115), .dinb(n21113), .dout(n21116));
  jnot g20935(.din(n21116), .dout(n21117));
  jand g20936(.dina(n20750), .dinb(n20676), .dout(n21118));
  jand g20937(.dina(n20751), .dinb(n20667), .dout(n21119));
  jor  g20938(.dina(n21119), .dinb(n21118), .dout(n21120));
  jand g20939(.dina(n20079), .dinb(n5365), .dout(n21121));
  jand g20940(.dina(n19545), .dinb(n5500), .dout(n21122));
  jand g20941(.dina(n19548), .dinb(n5424), .dout(n21123));
  jand g20942(.dina(n19551), .dinb(n5363), .dout(n21124));
  jor  g20943(.dina(n21124), .dinb(n21123), .dout(n21125));
  jor  g20944(.dina(n21125), .dinb(n21122), .dout(n21126));
  jor  g20945(.dina(n21126), .dinb(n21121), .dout(n21127));
  jxor g20946(.dina(n21127), .dinb(n72), .dout(n21128));
  jnot g20947(.din(n21128), .dout(n21129));
  jand g20948(.dina(n20748), .dinb(n20688), .dout(n21130));
  jand g20949(.dina(n20749), .dinb(n20679), .dout(n21131));
  jor  g20950(.dina(n21131), .dinb(n21130), .dout(n21132));
  jand g20951(.dina(n20746), .dinb(n20700), .dout(n21133));
  jand g20952(.dina(n20747), .dinb(n20691), .dout(n21134));
  jor  g20953(.dina(n21134), .dinb(n21133), .dout(n21135));
  jor  g20954(.dina(n19839), .dinb(n4724), .dout(n21136));
  jor  g20955(.dina(n19564), .dinb(n4905), .dout(n21137));
  jor  g20956(.dina(n19566), .dinb(n4735), .dout(n21138));
  jor  g20957(.dina(n19568), .dinb(n4733), .dout(n21139));
  jand g20958(.dina(n21139), .dinb(n21138), .dout(n21140));
  jand g20959(.dina(n21140), .dinb(n21137), .dout(n21141));
  jand g20960(.dina(n21141), .dinb(n21136), .dout(n21142));
  jxor g20961(.dina(n21142), .dinb(\a[29] ), .dout(n21143));
  jnot g20962(.din(n21143), .dout(n21144));
  jand g20963(.dina(n20745), .dinb(n20740), .dout(n21145));
  jand g20964(.dina(n1663), .dinb(n938), .dout(n21146));
  jand g20965(.dina(n21146), .dinb(n1435), .dout(n21147));
  jand g20966(.dina(n21147), .dinb(n3975), .dout(n21148));
  jand g20967(.dina(n4788), .dinb(n1932), .dout(n21149));
  jand g20968(.dina(n21149), .dinb(n21148), .dout(n21150));
  jand g20969(.dina(n476), .dinb(n371), .dout(n21151));
  jand g20970(.dina(n21151), .dinb(n4076), .dout(n21152));
  jand g20971(.dina(n12199), .dinb(n271), .dout(n21153));
  jand g20972(.dina(n21153), .dinb(n21152), .dout(n21154));
  jand g20973(.dina(n757), .dinb(n655), .dout(n21155));
  jand g20974(.dina(n21155), .dinb(n304), .dout(n21156));
  jand g20975(.dina(n614), .dinb(n607), .dout(n21157));
  jand g20976(.dina(n888), .dinb(n595), .dout(n21158));
  jand g20977(.dina(n21158), .dinb(n21157), .dout(n21159));
  jand g20978(.dina(n21159), .dinb(n21156), .dout(n21160));
  jand g20979(.dina(n21160), .dinb(n21154), .dout(n21161));
  jand g20980(.dina(n21161), .dinb(n5952), .dout(n21162));
  jand g20981(.dina(n21162), .dinb(n21150), .dout(n21163));
  jand g20982(.dina(n21163), .dinb(n7127), .dout(n21164));
  jand g20983(.dina(n21164), .dinb(n14337), .dout(n21165));
  jnot g20984(.din(n21165), .dout(n21166));
  jxor g20985(.dina(n21166), .dinb(n21145), .dout(n21167));
  jand g20986(.dina(n19826), .dinb(n732), .dout(n21168));
  jand g20987(.dina(n19572), .dinb(n3855), .dout(n21169));
  jand g20988(.dina(n19574), .dinb(n3858), .dout(n21170));
  jand g20989(.dina(n19576), .dinb(n3851), .dout(n21171));
  jor  g20990(.dina(n21171), .dinb(n21170), .dout(n21172));
  jor  g20991(.dina(n21172), .dinb(n21169), .dout(n21173));
  jor  g20992(.dina(n21173), .dinb(n21168), .dout(n21174));
  jxor g20993(.dina(n21174), .dinb(n21167), .dout(n21175));
  jxor g20994(.dina(n21175), .dinb(n21144), .dout(n21176));
  jxor g20995(.dina(n21176), .dinb(n21135), .dout(n21177));
  jnot g20996(.din(n21177), .dout(n21178));
  jor  g20997(.dina(n19964), .dinb(n4747), .dout(n21179));
  jor  g20998(.dina(n19553), .dinb(n4959), .dout(n21180));
  jor  g20999(.dina(n19558), .dinb(n4919), .dout(n21181));
  jor  g21000(.dina(n19562), .dinb(n4746), .dout(n21182));
  jand g21001(.dina(n21182), .dinb(n21181), .dout(n21183));
  jand g21002(.dina(n21183), .dinb(n21180), .dout(n21184));
  jand g21003(.dina(n21184), .dinb(n21179), .dout(n21185));
  jxor g21004(.dina(n21185), .dinb(\a[26] ), .dout(n21186));
  jxor g21005(.dina(n21186), .dinb(n21178), .dout(n21187));
  jxor g21006(.dina(n21187), .dinb(n21132), .dout(n21188));
  jxor g21007(.dina(n21188), .dinb(n21129), .dout(n21189));
  jxor g21008(.dina(n21189), .dinb(n21120), .dout(n21190));
  jnot g21009(.din(n21190), .dout(n21191));
  jand g21010(.dina(n20131), .dinb(n5693), .dout(n21192));
  jand g21011(.dina(n19539), .dinb(n6209), .dout(n21193));
  jand g21012(.dina(n19541), .dinb(n6131), .dout(n21194));
  jand g21013(.dina(n19543), .dinb(n5691), .dout(n21195));
  jor  g21014(.dina(n21195), .dinb(n21194), .dout(n21196));
  jor  g21015(.dina(n21196), .dinb(n21193), .dout(n21197));
  jor  g21016(.dina(n21197), .dinb(n21192), .dout(n21198));
  jxor g21017(.dina(n21198), .dinb(n4247), .dout(n21199));
  jxor g21018(.dina(n21199), .dinb(n21191), .dout(n21200));
  jxor g21019(.dina(n21200), .dinb(n21117), .dout(n21201));
  jxor g21020(.dina(n21201), .dinb(n21112), .dout(n21202));
  jxor g21021(.dina(n21202), .dinb(n21103), .dout(n21203));
  jnot g21022(.din(n21203), .dout(n21204));
  jand g21023(.dina(n20793), .dinb(n6936), .dout(n21205));
  jand g21024(.dina(n19527), .dinb(n7741), .dout(n21206));
  jand g21025(.dina(n19529), .dinb(n7613), .dout(n21207));
  jand g21026(.dina(n19531), .dinb(n6934), .dout(n21208));
  jor  g21027(.dina(n21208), .dinb(n21207), .dout(n21209));
  jor  g21028(.dina(n21209), .dinb(n21206), .dout(n21210));
  jor  g21029(.dina(n21210), .dinb(n21205), .dout(n21211));
  jxor g21030(.dina(n21211), .dinb(n5292), .dout(n21212));
  jxor g21031(.dina(n21212), .dinb(n21204), .dout(n21213));
  jxor g21032(.dina(n21213), .dinb(n21100), .dout(n21214));
  jxor g21033(.dina(n21214), .dinb(n21095), .dout(n21215));
  jxor g21034(.dina(n21215), .dinb(n21085), .dout(n21216));
  jnot g21035(.din(n21216), .dout(n21217));
  jxor g21036(.dina(n19655), .dinb(n19654), .dout(n21218));
  jand g21037(.dina(n21218), .dinb(n8771), .dout(n21219));
  jand g21038(.dina(n19515), .dinb(n9491), .dout(n21220));
  jand g21039(.dina(n19517), .dinb(n9126), .dout(n21221));
  jand g21040(.dina(n19519), .dinb(n8769), .dout(n21222));
  jor  g21041(.dina(n21222), .dinb(n21221), .dout(n21223));
  jor  g21042(.dina(n21223), .dinb(n21220), .dout(n21224));
  jor  g21043(.dina(n21224), .dinb(n21219), .dout(n21225));
  jxor g21044(.dina(n21225), .dinb(n6039), .dout(n21226));
  jor  g21045(.dina(n21226), .dinb(n21217), .dout(n21227));
  jxor g21046(.dina(n21083), .dinb(n21082), .dout(n21228));
  jnot g21047(.din(n21228), .dout(n21229));
  jxor g21048(.dina(n19652), .dinb(n19651), .dout(n21230));
  jand g21049(.dina(n21230), .dinb(n8771), .dout(n21231));
  jand g21050(.dina(n19517), .dinb(n9491), .dout(n21232));
  jand g21051(.dina(n19519), .dinb(n9126), .dout(n21233));
  jand g21052(.dina(n19521), .dinb(n8769), .dout(n21234));
  jor  g21053(.dina(n21234), .dinb(n21233), .dout(n21235));
  jor  g21054(.dina(n21235), .dinb(n21232), .dout(n21236));
  jor  g21055(.dina(n21236), .dinb(n21231), .dout(n21237));
  jxor g21056(.dina(n21237), .dinb(n6039), .dout(n21238));
  jor  g21057(.dina(n21238), .dinb(n21229), .dout(n21239));
  jxor g21058(.dina(n19649), .dinb(n19648), .dout(n21240));
  jand g21059(.dina(n21240), .dinb(n8771), .dout(n21241));
  jand g21060(.dina(n19519), .dinb(n9491), .dout(n21242));
  jand g21061(.dina(n19521), .dinb(n9126), .dout(n21243));
  jand g21062(.dina(n19523), .dinb(n8769), .dout(n21244));
  jor  g21063(.dina(n21244), .dinb(n21243), .dout(n21245));
  jor  g21064(.dina(n21245), .dinb(n21242), .dout(n21246));
  jor  g21065(.dina(n21246), .dinb(n21241), .dout(n21247));
  jxor g21066(.dina(n21247), .dinb(n6039), .dout(n21248));
  jnot g21067(.din(n21248), .dout(n21249));
  jxor g21068(.dina(n21078), .dinb(n21077), .dout(n21250));
  jand g21069(.dina(n21250), .dinb(n21249), .dout(n21251));
  jand g21070(.dina(n21086), .dinb(n8771), .dout(n21252));
  jand g21071(.dina(n19521), .dinb(n9491), .dout(n21253));
  jand g21072(.dina(n19523), .dinb(n9126), .dout(n21254));
  jand g21073(.dina(n19525), .dinb(n8769), .dout(n21255));
  jor  g21074(.dina(n21255), .dinb(n21254), .dout(n21256));
  jor  g21075(.dina(n21256), .dinb(n21253), .dout(n21257));
  jor  g21076(.dina(n21257), .dinb(n21252), .dout(n21258));
  jxor g21077(.dina(n21258), .dinb(n6039), .dout(n21259));
  jnot g21078(.din(n21259), .dout(n21260));
  jxor g21079(.dina(n21073), .dinb(n21072), .dout(n21261));
  jand g21080(.dina(n21261), .dinb(n21260), .dout(n21262));
  jxor g21081(.dina(n21070), .dinb(n21069), .dout(n21263));
  jnot g21082(.din(n21263), .dout(n21264));
  jand g21083(.dina(n19770), .dinb(n8771), .dout(n21265));
  jand g21084(.dina(n19523), .dinb(n9491), .dout(n21266));
  jand g21085(.dina(n19525), .dinb(n9126), .dout(n21267));
  jand g21086(.dina(n19527), .dinb(n8769), .dout(n21268));
  jor  g21087(.dina(n21268), .dinb(n21267), .dout(n21269));
  jor  g21088(.dina(n21269), .dinb(n21266), .dout(n21270));
  jor  g21089(.dina(n21270), .dinb(n21265), .dout(n21271));
  jxor g21090(.dina(n21271), .dinb(n6039), .dout(n21272));
  jor  g21091(.dina(n21272), .dinb(n21264), .dout(n21273));
  jxor g21092(.dina(n21067), .dinb(n21066), .dout(n21274));
  jnot g21093(.din(n21274), .dout(n21275));
  jand g21094(.dina(n20781), .dinb(n8771), .dout(n21276));
  jand g21095(.dina(n19525), .dinb(n9491), .dout(n21277));
  jand g21096(.dina(n19527), .dinb(n9126), .dout(n21278));
  jand g21097(.dina(n19529), .dinb(n8769), .dout(n21279));
  jor  g21098(.dina(n21279), .dinb(n21278), .dout(n21280));
  jor  g21099(.dina(n21280), .dinb(n21277), .dout(n21281));
  jor  g21100(.dina(n21281), .dinb(n21276), .dout(n21282));
  jxor g21101(.dina(n21282), .dinb(n6039), .dout(n21283));
  jor  g21102(.dina(n21283), .dinb(n21275), .dout(n21284));
  jxor g21103(.dina(n21064), .dinb(n21063), .dout(n21285));
  jnot g21104(.din(n21285), .dout(n21286));
  jand g21105(.dina(n20793), .dinb(n8771), .dout(n21287));
  jand g21106(.dina(n19527), .dinb(n9491), .dout(n21288));
  jand g21107(.dina(n19529), .dinb(n9126), .dout(n21289));
  jand g21108(.dina(n19531), .dinb(n8769), .dout(n21290));
  jor  g21109(.dina(n21290), .dinb(n21289), .dout(n21291));
  jor  g21110(.dina(n21291), .dinb(n21288), .dout(n21292));
  jor  g21111(.dina(n21292), .dinb(n21287), .dout(n21293));
  jxor g21112(.dina(n21293), .dinb(n6039), .dout(n21294));
  jor  g21113(.dina(n21294), .dinb(n21286), .dout(n21295));
  jand g21114(.dina(n20767), .dinb(n8771), .dout(n21296));
  jand g21115(.dina(n19529), .dinb(n9491), .dout(n21297));
  jand g21116(.dina(n19531), .dinb(n9126), .dout(n21298));
  jand g21117(.dina(n19533), .dinb(n8769), .dout(n21299));
  jor  g21118(.dina(n21299), .dinb(n21298), .dout(n21300));
  jor  g21119(.dina(n21300), .dinb(n21297), .dout(n21301));
  jor  g21120(.dina(n21301), .dinb(n21296), .dout(n21302));
  jxor g21121(.dina(n21302), .dinb(n6039), .dout(n21303));
  jnot g21122(.din(n21303), .dout(n21304));
  jxor g21123(.dina(n21059), .dinb(n21058), .dout(n21305));
  jand g21124(.dina(n21305), .dinb(n21304), .dout(n21306));
  jand g21125(.dina(n19780), .dinb(n8771), .dout(n21307));
  jand g21126(.dina(n19531), .dinb(n9491), .dout(n21308));
  jand g21127(.dina(n19533), .dinb(n9126), .dout(n21309));
  jand g21128(.dina(n19535), .dinb(n8769), .dout(n21310));
  jor  g21129(.dina(n21310), .dinb(n21309), .dout(n21311));
  jor  g21130(.dina(n21311), .dinb(n21308), .dout(n21312));
  jor  g21131(.dina(n21312), .dinb(n21307), .dout(n21313));
  jxor g21132(.dina(n21313), .dinb(n6039), .dout(n21314));
  jnot g21133(.din(n21314), .dout(n21315));
  jxor g21134(.dina(n21054), .dinb(n21053), .dout(n21316));
  jand g21135(.dina(n21316), .dinb(n21315), .dout(n21317));
  jand g21136(.dina(n20399), .dinb(n8771), .dout(n21318));
  jand g21137(.dina(n19533), .dinb(n9491), .dout(n21319));
  jand g21138(.dina(n19535), .dinb(n9126), .dout(n21320));
  jand g21139(.dina(n19537), .dinb(n8769), .dout(n21321));
  jor  g21140(.dina(n21321), .dinb(n21320), .dout(n21322));
  jor  g21141(.dina(n21322), .dinb(n21319), .dout(n21323));
  jor  g21142(.dina(n21323), .dinb(n21318), .dout(n21324));
  jxor g21143(.dina(n21324), .dinb(n6039), .dout(n21325));
  jnot g21144(.din(n21325), .dout(n21326));
  jxor g21145(.dina(n21049), .dinb(n21048), .dout(n21327));
  jand g21146(.dina(n21327), .dinb(n21326), .dout(n21328));
  jxor g21147(.dina(n21046), .dinb(n21045), .dout(n21329));
  jnot g21148(.din(n21329), .dout(n21330));
  jand g21149(.dina(n20413), .dinb(n8771), .dout(n21331));
  jand g21150(.dina(n19535), .dinb(n9491), .dout(n21332));
  jand g21151(.dina(n19537), .dinb(n9126), .dout(n21333));
  jand g21152(.dina(n19539), .dinb(n8769), .dout(n21334));
  jor  g21153(.dina(n21334), .dinb(n21333), .dout(n21335));
  jor  g21154(.dina(n21335), .dinb(n21332), .dout(n21336));
  jor  g21155(.dina(n21336), .dinb(n21331), .dout(n21337));
  jxor g21156(.dina(n21337), .dinb(n6039), .dout(n21338));
  jor  g21157(.dina(n21338), .dinb(n21330), .dout(n21339));
  jxor g21158(.dina(n21043), .dinb(n21042), .dout(n21340));
  jnot g21159(.din(n21340), .dout(n21341));
  jand g21160(.dina(n20387), .dinb(n8771), .dout(n21342));
  jand g21161(.dina(n19537), .dinb(n9491), .dout(n21343));
  jand g21162(.dina(n19539), .dinb(n9126), .dout(n21344));
  jand g21163(.dina(n19541), .dinb(n8769), .dout(n21345));
  jor  g21164(.dina(n21345), .dinb(n21344), .dout(n21346));
  jor  g21165(.dina(n21346), .dinb(n21343), .dout(n21347));
  jor  g21166(.dina(n21347), .dinb(n21342), .dout(n21348));
  jxor g21167(.dina(n21348), .dinb(n6039), .dout(n21349));
  jor  g21168(.dina(n21349), .dinb(n21341), .dout(n21350));
  jxor g21169(.dina(n21040), .dinb(n21039), .dout(n21351));
  jnot g21170(.din(n21351), .dout(n21352));
  jand g21171(.dina(n20131), .dinb(n8771), .dout(n21353));
  jand g21172(.dina(n19539), .dinb(n9491), .dout(n21354));
  jand g21173(.dina(n19541), .dinb(n9126), .dout(n21355));
  jand g21174(.dina(n19543), .dinb(n8769), .dout(n21356));
  jor  g21175(.dina(n21356), .dinb(n21355), .dout(n21357));
  jor  g21176(.dina(n21357), .dinb(n21354), .dout(n21358));
  jor  g21177(.dina(n21358), .dinb(n21353), .dout(n21359));
  jxor g21178(.dina(n21359), .dinb(n6039), .dout(n21360));
  jor  g21179(.dina(n21360), .dinb(n21352), .dout(n21361));
  jand g21180(.dina(n20141), .dinb(n8771), .dout(n21362));
  jand g21181(.dina(n19541), .dinb(n9491), .dout(n21363));
  jand g21182(.dina(n19543), .dinb(n9126), .dout(n21364));
  jand g21183(.dina(n19545), .dinb(n8769), .dout(n21365));
  jor  g21184(.dina(n21365), .dinb(n21364), .dout(n21366));
  jor  g21185(.dina(n21366), .dinb(n21363), .dout(n21367));
  jor  g21186(.dina(n21367), .dinb(n21362), .dout(n21368));
  jxor g21187(.dina(n21368), .dinb(n6039), .dout(n21369));
  jnot g21188(.din(n21369), .dout(n21370));
  jxor g21189(.dina(n21035), .dinb(n21034), .dout(n21371));
  jand g21190(.dina(n21371), .dinb(n21370), .dout(n21372));
  jand g21191(.dina(n20153), .dinb(n8771), .dout(n21373));
  jand g21192(.dina(n19543), .dinb(n9491), .dout(n21374));
  jand g21193(.dina(n19545), .dinb(n9126), .dout(n21375));
  jand g21194(.dina(n19548), .dinb(n8769), .dout(n21376));
  jor  g21195(.dina(n21376), .dinb(n21375), .dout(n21377));
  jor  g21196(.dina(n21377), .dinb(n21374), .dout(n21378));
  jor  g21197(.dina(n21378), .dinb(n21373), .dout(n21379));
  jxor g21198(.dina(n21379), .dinb(n6039), .dout(n21380));
  jnot g21199(.din(n21380), .dout(n21381));
  jxor g21200(.dina(n21030), .dinb(n21029), .dout(n21382));
  jand g21201(.dina(n21382), .dinb(n21381), .dout(n21383));
  jand g21202(.dina(n20079), .dinb(n8771), .dout(n21384));
  jand g21203(.dina(n19545), .dinb(n9491), .dout(n21385));
  jand g21204(.dina(n19548), .dinb(n9126), .dout(n21386));
  jand g21205(.dina(n19551), .dinb(n8769), .dout(n21387));
  jor  g21206(.dina(n21387), .dinb(n21386), .dout(n21388));
  jor  g21207(.dina(n21388), .dinb(n21385), .dout(n21389));
  jor  g21208(.dina(n21389), .dinb(n21384), .dout(n21390));
  jxor g21209(.dina(n21390), .dinb(n6039), .dout(n21391));
  jnot g21210(.din(n21391), .dout(n21392));
  jxor g21211(.dina(n21025), .dinb(n21024), .dout(n21393));
  jand g21212(.dina(n21393), .dinb(n21392), .dout(n21394));
  jxor g21213(.dina(n21022), .dinb(n21021), .dout(n21395));
  jnot g21214(.din(n21395), .dout(n21396));
  jor  g21215(.dina(n19940), .dinb(n8772), .dout(n21397));
  jor  g21216(.dina(n19547), .dinb(n9490), .dout(n21398));
  jor  g21217(.dina(n19550), .dinb(n9127), .dout(n21399));
  jor  g21218(.dina(n19553), .dinb(n8770), .dout(n21400));
  jand g21219(.dina(n21400), .dinb(n21399), .dout(n21401));
  jand g21220(.dina(n21401), .dinb(n21398), .dout(n21402));
  jand g21221(.dina(n21402), .dinb(n21397), .dout(n21403));
  jxor g21222(.dina(n21403), .dinb(\a[8] ), .dout(n21404));
  jor  g21223(.dina(n21404), .dinb(n21396), .dout(n21405));
  jxor g21224(.dina(n21019), .dinb(n21018), .dout(n21406));
  jnot g21225(.din(n21406), .dout(n21407));
  jor  g21226(.dina(n19952), .dinb(n8772), .dout(n21408));
  jor  g21227(.dina(n19550), .dinb(n9490), .dout(n21409));
  jor  g21228(.dina(n19553), .dinb(n9127), .dout(n21410));
  jor  g21229(.dina(n19558), .dinb(n8770), .dout(n21411));
  jand g21230(.dina(n21411), .dinb(n21410), .dout(n21412));
  jand g21231(.dina(n21412), .dinb(n21409), .dout(n21413));
  jand g21232(.dina(n21413), .dinb(n21408), .dout(n21414));
  jxor g21233(.dina(n21414), .dinb(\a[8] ), .dout(n21415));
  jor  g21234(.dina(n21415), .dinb(n21407), .dout(n21416));
  jxor g21235(.dina(n21016), .dinb(n21015), .dout(n21417));
  jnot g21236(.din(n21417), .dout(n21418));
  jor  g21237(.dina(n19964), .dinb(n8772), .dout(n21419));
  jor  g21238(.dina(n19553), .dinb(n9490), .dout(n21420));
  jor  g21239(.dina(n19558), .dinb(n9127), .dout(n21421));
  jor  g21240(.dina(n19562), .dinb(n8770), .dout(n21422));
  jand g21241(.dina(n21422), .dinb(n21421), .dout(n21423));
  jand g21242(.dina(n21423), .dinb(n21420), .dout(n21424));
  jand g21243(.dina(n21424), .dinb(n21419), .dout(n21425));
  jxor g21244(.dina(n21425), .dinb(\a[8] ), .dout(n21426));
  jor  g21245(.dina(n21426), .dinb(n21418), .dout(n21427));
  jor  g21246(.dina(n19906), .dinb(n8772), .dout(n21428));
  jor  g21247(.dina(n19558), .dinb(n9490), .dout(n21429));
  jor  g21248(.dina(n19562), .dinb(n9127), .dout(n21430));
  jor  g21249(.dina(n19564), .dinb(n8770), .dout(n21431));
  jand g21250(.dina(n21431), .dinb(n21430), .dout(n21432));
  jand g21251(.dina(n21432), .dinb(n21429), .dout(n21433));
  jand g21252(.dina(n21433), .dinb(n21428), .dout(n21434));
  jxor g21253(.dina(n21434), .dinb(\a[8] ), .dout(n21435));
  jnot g21254(.din(n21435), .dout(n21436));
  jxor g21255(.dina(n21013), .dinb(n21012), .dout(n21437));
  jand g21256(.dina(n21437), .dinb(n21436), .dout(n21438));
  jor  g21257(.dina(n19790), .dinb(n8772), .dout(n21439));
  jor  g21258(.dina(n19562), .dinb(n9490), .dout(n21440));
  jor  g21259(.dina(n19564), .dinb(n9127), .dout(n21441));
  jor  g21260(.dina(n19566), .dinb(n8770), .dout(n21442));
  jand g21261(.dina(n21442), .dinb(n21441), .dout(n21443));
  jand g21262(.dina(n21443), .dinb(n21440), .dout(n21444));
  jand g21263(.dina(n21444), .dinb(n21439), .dout(n21445));
  jxor g21264(.dina(n21445), .dinb(\a[8] ), .dout(n21446));
  jnot g21265(.din(n21446), .dout(n21447));
  jxor g21266(.dina(n21010), .dinb(n21009), .dout(n21448));
  jand g21267(.dina(n21448), .dinb(n21447), .dout(n21449));
  jor  g21268(.dina(n19839), .dinb(n8772), .dout(n21450));
  jor  g21269(.dina(n19564), .dinb(n9490), .dout(n21451));
  jor  g21270(.dina(n19566), .dinb(n9127), .dout(n21452));
  jor  g21271(.dina(n19568), .dinb(n8770), .dout(n21453));
  jand g21272(.dina(n21453), .dinb(n21452), .dout(n21454));
  jand g21273(.dina(n21454), .dinb(n21451), .dout(n21455));
  jand g21274(.dina(n21455), .dinb(n21450), .dout(n21456));
  jxor g21275(.dina(n21456), .dinb(\a[8] ), .dout(n21457));
  jnot g21276(.din(n21457), .dout(n21458));
  jor  g21277(.dina(n20990), .dinb(n5833), .dout(n21459));
  jxor g21278(.dina(n21459), .dinb(n20998), .dout(n21460));
  jand g21279(.dina(n21460), .dinb(n21458), .dout(n21461));
  jor  g21280(.dina(n19852), .dinb(n8772), .dout(n21462));
  jor  g21281(.dina(n19566), .dinb(n9490), .dout(n21463));
  jor  g21282(.dina(n19568), .dinb(n9127), .dout(n21464));
  jor  g21283(.dina(n19570), .dinb(n8770), .dout(n21465));
  jand g21284(.dina(n21465), .dinb(n21464), .dout(n21466));
  jand g21285(.dina(n21466), .dinb(n21463), .dout(n21467));
  jand g21286(.dina(n21467), .dinb(n21462), .dout(n21468));
  jxor g21287(.dina(n21468), .dinb(\a[8] ), .dout(n21469));
  jnot g21288(.din(n21469), .dout(n21470));
  jand g21289(.dina(n20987), .dinb(\a[11] ), .dout(n21471));
  jxor g21290(.dina(n21471), .dinb(n20985), .dout(n21472));
  jand g21291(.dina(n21472), .dinb(n21470), .dout(n21473));
  jand g21292(.dina(n19813), .dinb(n8771), .dout(n21474));
  jand g21293(.dina(n19576), .dinb(n9126), .dout(n21475));
  jand g21294(.dina(n19574), .dinb(n9491), .dout(n21476));
  jor  g21295(.dina(n21476), .dinb(n21475), .dout(n21477));
  jor  g21296(.dina(n21477), .dinb(n21474), .dout(n21478));
  jnot g21297(.din(n21478), .dout(n21479));
  jand g21298(.dina(n19576), .dinb(n8765), .dout(n21480));
  jnot g21299(.din(n21480), .dout(n21481));
  jand g21300(.dina(n21481), .dinb(\a[8] ), .dout(n21482));
  jand g21301(.dina(n21482), .dinb(n21479), .dout(n21483));
  jand g21302(.dina(n19826), .dinb(n8771), .dout(n21484));
  jand g21303(.dina(n19572), .dinb(n9491), .dout(n21485));
  jand g21304(.dina(n19574), .dinb(n9126), .dout(n21486));
  jand g21305(.dina(n19576), .dinb(n8769), .dout(n21487));
  jor  g21306(.dina(n21487), .dinb(n21486), .dout(n21488));
  jor  g21307(.dina(n21488), .dinb(n21485), .dout(n21489));
  jor  g21308(.dina(n21489), .dinb(n21484), .dout(n21490));
  jnot g21309(.din(n21490), .dout(n21491));
  jand g21310(.dina(n21491), .dinb(n21483), .dout(n21492));
  jand g21311(.dina(n21492), .dinb(n20987), .dout(n21493));
  jor  g21312(.dina(n19801), .dinb(n8772), .dout(n21494));
  jor  g21313(.dina(n19568), .dinb(n9490), .dout(n21495));
  jor  g21314(.dina(n19570), .dinb(n9127), .dout(n21496));
  jor  g21315(.dina(n19575), .dinb(n8770), .dout(n21497));
  jand g21316(.dina(n21497), .dinb(n21496), .dout(n21498));
  jand g21317(.dina(n21498), .dinb(n21495), .dout(n21499));
  jand g21318(.dina(n21499), .dinb(n21494), .dout(n21500));
  jxor g21319(.dina(n21500), .dinb(\a[8] ), .dout(n21501));
  jnot g21320(.din(n21501), .dout(n21502));
  jxor g21321(.dina(n21492), .dinb(n20987), .dout(n21503));
  jand g21322(.dina(n21503), .dinb(n21502), .dout(n21504));
  jor  g21323(.dina(n21504), .dinb(n21493), .dout(n21505));
  jxor g21324(.dina(n21472), .dinb(n21470), .dout(n21506));
  jand g21325(.dina(n21506), .dinb(n21505), .dout(n21507));
  jor  g21326(.dina(n21507), .dinb(n21473), .dout(n21508));
  jxor g21327(.dina(n21460), .dinb(n21458), .dout(n21509));
  jand g21328(.dina(n21509), .dinb(n21508), .dout(n21510));
  jor  g21329(.dina(n21510), .dinb(n21461), .dout(n21511));
  jxor g21330(.dina(n21448), .dinb(n21447), .dout(n21512));
  jand g21331(.dina(n21512), .dinb(n21511), .dout(n21513));
  jor  g21332(.dina(n21513), .dinb(n21449), .dout(n21514));
  jxor g21333(.dina(n21437), .dinb(n21436), .dout(n21515));
  jand g21334(.dina(n21515), .dinb(n21514), .dout(n21516));
  jor  g21335(.dina(n21516), .dinb(n21438), .dout(n21517));
  jxor g21336(.dina(n21426), .dinb(n21418), .dout(n21518));
  jand g21337(.dina(n21518), .dinb(n21517), .dout(n21519));
  jnot g21338(.din(n21519), .dout(n21520));
  jand g21339(.dina(n21520), .dinb(n21427), .dout(n21521));
  jnot g21340(.din(n21521), .dout(n21522));
  jxor g21341(.dina(n21415), .dinb(n21407), .dout(n21523));
  jand g21342(.dina(n21523), .dinb(n21522), .dout(n21524));
  jnot g21343(.din(n21524), .dout(n21525));
  jand g21344(.dina(n21525), .dinb(n21416), .dout(n21526));
  jnot g21345(.din(n21526), .dout(n21527));
  jxor g21346(.dina(n21404), .dinb(n21396), .dout(n21528));
  jand g21347(.dina(n21528), .dinb(n21527), .dout(n21529));
  jnot g21348(.din(n21529), .dout(n21530));
  jand g21349(.dina(n21530), .dinb(n21405), .dout(n21531));
  jnot g21350(.din(n21531), .dout(n21532));
  jxor g21351(.dina(n21393), .dinb(n21392), .dout(n21533));
  jand g21352(.dina(n21533), .dinb(n21532), .dout(n21534));
  jor  g21353(.dina(n21534), .dinb(n21394), .dout(n21535));
  jxor g21354(.dina(n21382), .dinb(n21381), .dout(n21536));
  jand g21355(.dina(n21536), .dinb(n21535), .dout(n21537));
  jor  g21356(.dina(n21537), .dinb(n21383), .dout(n21538));
  jxor g21357(.dina(n21371), .dinb(n21370), .dout(n21539));
  jand g21358(.dina(n21539), .dinb(n21538), .dout(n21540));
  jor  g21359(.dina(n21540), .dinb(n21372), .dout(n21541));
  jxor g21360(.dina(n21360), .dinb(n21352), .dout(n21542));
  jand g21361(.dina(n21542), .dinb(n21541), .dout(n21543));
  jnot g21362(.din(n21543), .dout(n21544));
  jand g21363(.dina(n21544), .dinb(n21361), .dout(n21545));
  jnot g21364(.din(n21545), .dout(n21546));
  jxor g21365(.dina(n21349), .dinb(n21341), .dout(n21547));
  jand g21366(.dina(n21547), .dinb(n21546), .dout(n21548));
  jnot g21367(.din(n21548), .dout(n21549));
  jand g21368(.dina(n21549), .dinb(n21350), .dout(n21550));
  jnot g21369(.din(n21550), .dout(n21551));
  jxor g21370(.dina(n21338), .dinb(n21330), .dout(n21552));
  jand g21371(.dina(n21552), .dinb(n21551), .dout(n21553));
  jnot g21372(.din(n21553), .dout(n21554));
  jand g21373(.dina(n21554), .dinb(n21339), .dout(n21555));
  jnot g21374(.din(n21555), .dout(n21556));
  jxor g21375(.dina(n21327), .dinb(n21326), .dout(n21557));
  jand g21376(.dina(n21557), .dinb(n21556), .dout(n21558));
  jor  g21377(.dina(n21558), .dinb(n21328), .dout(n21559));
  jxor g21378(.dina(n21316), .dinb(n21315), .dout(n21560));
  jand g21379(.dina(n21560), .dinb(n21559), .dout(n21561));
  jor  g21380(.dina(n21561), .dinb(n21317), .dout(n21562));
  jxor g21381(.dina(n21305), .dinb(n21304), .dout(n21563));
  jand g21382(.dina(n21563), .dinb(n21562), .dout(n21564));
  jor  g21383(.dina(n21564), .dinb(n21306), .dout(n21565));
  jxor g21384(.dina(n21294), .dinb(n21286), .dout(n21566));
  jand g21385(.dina(n21566), .dinb(n21565), .dout(n21567));
  jnot g21386(.din(n21567), .dout(n21568));
  jand g21387(.dina(n21568), .dinb(n21295), .dout(n21569));
  jnot g21388(.din(n21569), .dout(n21570));
  jxor g21389(.dina(n21283), .dinb(n21275), .dout(n21571));
  jand g21390(.dina(n21571), .dinb(n21570), .dout(n21572));
  jnot g21391(.din(n21572), .dout(n21573));
  jand g21392(.dina(n21573), .dinb(n21284), .dout(n21574));
  jnot g21393(.din(n21574), .dout(n21575));
  jxor g21394(.dina(n21272), .dinb(n21264), .dout(n21576));
  jand g21395(.dina(n21576), .dinb(n21575), .dout(n21577));
  jnot g21396(.din(n21577), .dout(n21578));
  jand g21397(.dina(n21578), .dinb(n21273), .dout(n21579));
  jnot g21398(.din(n21579), .dout(n21580));
  jxor g21399(.dina(n21261), .dinb(n21260), .dout(n21581));
  jand g21400(.dina(n21581), .dinb(n21580), .dout(n21582));
  jor  g21401(.dina(n21582), .dinb(n21262), .dout(n21583));
  jxor g21402(.dina(n21250), .dinb(n21249), .dout(n21584));
  jand g21403(.dina(n21584), .dinb(n21583), .dout(n21585));
  jor  g21404(.dina(n21585), .dinb(n21251), .dout(n21586));
  jxor g21405(.dina(n21238), .dinb(n21229), .dout(n21587));
  jand g21406(.dina(n21587), .dinb(n21586), .dout(n21588));
  jnot g21407(.din(n21588), .dout(n21589));
  jand g21408(.dina(n21589), .dinb(n21239), .dout(n21590));
  jnot g21409(.din(n21590), .dout(n21591));
  jxor g21410(.dina(n21226), .dinb(n21217), .dout(n21592));
  jand g21411(.dina(n21592), .dinb(n21591), .dout(n21593));
  jnot g21412(.din(n21593), .dout(n21594));
  jand g21413(.dina(n21594), .dinb(n21227), .dout(n21595));
  jnot g21414(.din(n21595), .dout(n21596));
  jand g21415(.dina(n21214), .dinb(n21095), .dout(n21597));
  jand g21416(.dina(n21215), .dinb(n21085), .dout(n21598));
  jor  g21417(.dina(n21598), .dinb(n21597), .dout(n21599));
  jand g21418(.dina(n21240), .dinb(n7890), .dout(n21600));
  jand g21419(.dina(n19519), .dinb(n8441), .dout(n21601));
  jand g21420(.dina(n19521), .dinb(n8154), .dout(n21602));
  jand g21421(.dina(n19523), .dinb(n7888), .dout(n21603));
  jor  g21422(.dina(n21603), .dinb(n21602), .dout(n21604));
  jor  g21423(.dina(n21604), .dinb(n21601), .dout(n21605));
  jor  g21424(.dina(n21605), .dinb(n21600), .dout(n21606));
  jxor g21425(.dina(n21606), .dinb(n5833), .dout(n21607));
  jnot g21426(.din(n21607), .dout(n21608));
  jor  g21427(.dina(n21212), .dinb(n21204), .dout(n21609));
  jand g21428(.dina(n21213), .dinb(n21100), .dout(n21610));
  jnot g21429(.din(n21610), .dout(n21611));
  jand g21430(.dina(n21611), .dinb(n21609), .dout(n21612));
  jnot g21431(.din(n21612), .dout(n21613));
  jand g21432(.dina(n21201), .dinb(n21112), .dout(n21614));
  jand g21433(.dina(n21202), .dinb(n21103), .dout(n21615));
  jor  g21434(.dina(n21615), .dinb(n21614), .dout(n21616));
  jand g21435(.dina(n19780), .dinb(n6340), .dout(n21617));
  jand g21436(.dina(n19531), .dinb(n6798), .dout(n21618));
  jand g21437(.dina(n19533), .dinb(n6556), .dout(n21619));
  jand g21438(.dina(n19535), .dinb(n6338), .dout(n21620));
  jor  g21439(.dina(n21620), .dinb(n21619), .dout(n21621));
  jor  g21440(.dina(n21621), .dinb(n21618), .dout(n21622));
  jor  g21441(.dina(n21622), .dinb(n21617), .dout(n21623));
  jxor g21442(.dina(n21623), .dinb(n5064), .dout(n21624));
  jnot g21443(.din(n21624), .dout(n21625));
  jor  g21444(.dina(n21199), .dinb(n21191), .dout(n21626));
  jand g21445(.dina(n21200), .dinb(n21117), .dout(n21627));
  jnot g21446(.din(n21627), .dout(n21628));
  jand g21447(.dina(n21628), .dinb(n21626), .dout(n21629));
  jnot g21448(.din(n21629), .dout(n21630));
  jand g21449(.dina(n21188), .dinb(n21129), .dout(n21631));
  jand g21450(.dina(n21189), .dinb(n21120), .dout(n21632));
  jor  g21451(.dina(n21632), .dinb(n21631), .dout(n21633));
  jand g21452(.dina(n20153), .dinb(n5365), .dout(n21634));
  jand g21453(.dina(n19543), .dinb(n5500), .dout(n21635));
  jand g21454(.dina(n19545), .dinb(n5424), .dout(n21636));
  jand g21455(.dina(n19548), .dinb(n5363), .dout(n21637));
  jor  g21456(.dina(n21637), .dinb(n21636), .dout(n21638));
  jor  g21457(.dina(n21638), .dinb(n21635), .dout(n21639));
  jor  g21458(.dina(n21639), .dinb(n21634), .dout(n21640));
  jxor g21459(.dina(n21640), .dinb(n72), .dout(n21641));
  jnot g21460(.din(n21641), .dout(n21642));
  jor  g21461(.dina(n21186), .dinb(n21178), .dout(n21643));
  jand g21462(.dina(n21187), .dinb(n21132), .dout(n21644));
  jnot g21463(.din(n21644), .dout(n21645));
  jand g21464(.dina(n21645), .dinb(n21643), .dout(n21646));
  jnot g21465(.din(n21646), .dout(n21647));
  jand g21466(.dina(n21175), .dinb(n21144), .dout(n21648));
  jand g21467(.dina(n21176), .dinb(n21135), .dout(n21649));
  jor  g21468(.dina(n21649), .dinb(n21648), .dout(n21650));
  jor  g21469(.dina(n19790), .dinb(n4724), .dout(n21651));
  jor  g21470(.dina(n19562), .dinb(n4905), .dout(n21652));
  jor  g21471(.dina(n19564), .dinb(n4735), .dout(n21653));
  jor  g21472(.dina(n19566), .dinb(n4733), .dout(n21654));
  jand g21473(.dina(n21654), .dinb(n21653), .dout(n21655));
  jand g21474(.dina(n21655), .dinb(n21652), .dout(n21656));
  jand g21475(.dina(n21656), .dinb(n21651), .dout(n21657));
  jxor g21476(.dina(n21657), .dinb(\a[29] ), .dout(n21658));
  jnot g21477(.din(n21658), .dout(n21659));
  jand g21478(.dina(n21166), .dinb(n21145), .dout(n21660));
  jnot g21479(.din(n21145), .dout(n21661));
  jand g21480(.dina(n21165), .dinb(n21661), .dout(n21662));
  jnot g21481(.din(n21662), .dout(n21663));
  jand g21482(.dina(n21174), .dinb(n21663), .dout(n21664));
  jor  g21483(.dina(n21664), .dinb(n21660), .dout(n21665));
  jand g21484(.dina(n1500), .dinb(n752), .dout(n21666));
  jand g21485(.dina(n827), .dinb(n277), .dout(n21667));
  jand g21486(.dina(n21667), .dinb(n21666), .dout(n21668));
  jand g21487(.dina(n965), .dinb(n372), .dout(n21669));
  jand g21488(.dina(n21669), .dinb(n506), .dout(n21670));
  jand g21489(.dina(n450), .dinb(n382), .dout(n21671));
  jand g21490(.dina(n1014), .dinb(n517), .dout(n21672));
  jand g21491(.dina(n21672), .dinb(n21671), .dout(n21673));
  jand g21492(.dina(n21673), .dinb(n21670), .dout(n21674));
  jand g21493(.dina(n21674), .dinb(n21668), .dout(n21675));
  jand g21494(.dina(n5768), .dinb(n4670), .dout(n21676));
  jand g21495(.dina(n21676), .dinb(n3092), .dout(n21677));
  jand g21496(.dina(n21677), .dinb(n2440), .dout(n21678));
  jand g21497(.dina(n21678), .dinb(n21675), .dout(n21679));
  jand g21498(.dina(n6025), .dinb(n4815), .dout(n21680));
  jand g21499(.dina(n21680), .dinb(n21679), .dout(n21681));
  jand g21500(.dina(n21681), .dinb(n2735), .dout(n21682));
  jand g21501(.dina(n21682), .dinb(n1810), .dout(n21683));
  jnot g21502(.din(n21683), .dout(n21684));
  jxor g21503(.dina(n19579), .dinb(n19573), .dout(n21685));
  jand g21504(.dina(n21685), .dinb(n732), .dout(n21686));
  jxor g21505(.dina(n19371), .dinb(n19369), .dout(n21687));
  jand g21506(.dina(n21687), .dinb(n3855), .dout(n21688));
  jand g21507(.dina(n19574), .dinb(n3851), .dout(n21689));
  jand g21508(.dina(n19572), .dinb(n3858), .dout(n21690));
  jor  g21509(.dina(n21690), .dinb(n21689), .dout(n21691));
  jor  g21510(.dina(n21691), .dinb(n21688), .dout(n21692));
  jor  g21511(.dina(n21692), .dinb(n21686), .dout(n21693));
  jxor g21512(.dina(n21693), .dinb(n21684), .dout(n21694));
  jxor g21513(.dina(n21694), .dinb(n21665), .dout(n21695));
  jxor g21514(.dina(n21695), .dinb(n21659), .dout(n21696));
  jxor g21515(.dina(n21696), .dinb(n21650), .dout(n21697));
  jnot g21516(.din(n21697), .dout(n21698));
  jor  g21517(.dina(n19952), .dinb(n4747), .dout(n21699));
  jor  g21518(.dina(n19550), .dinb(n4959), .dout(n21700));
  jor  g21519(.dina(n19553), .dinb(n4919), .dout(n21701));
  jor  g21520(.dina(n19558), .dinb(n4746), .dout(n21702));
  jand g21521(.dina(n21702), .dinb(n21701), .dout(n21703));
  jand g21522(.dina(n21703), .dinb(n21700), .dout(n21704));
  jand g21523(.dina(n21704), .dinb(n21699), .dout(n21705));
  jxor g21524(.dina(n21705), .dinb(\a[26] ), .dout(n21706));
  jxor g21525(.dina(n21706), .dinb(n21698), .dout(n21707));
  jxor g21526(.dina(n21707), .dinb(n21647), .dout(n21708));
  jxor g21527(.dina(n21708), .dinb(n21642), .dout(n21709));
  jxor g21528(.dina(n21709), .dinb(n21633), .dout(n21710));
  jnot g21529(.din(n21710), .dout(n21711));
  jand g21530(.dina(n20387), .dinb(n5693), .dout(n21712));
  jand g21531(.dina(n19537), .dinb(n6209), .dout(n21713));
  jand g21532(.dina(n19539), .dinb(n6131), .dout(n21714));
  jand g21533(.dina(n19541), .dinb(n5691), .dout(n21715));
  jor  g21534(.dina(n21715), .dinb(n21714), .dout(n21716));
  jor  g21535(.dina(n21716), .dinb(n21713), .dout(n21717));
  jor  g21536(.dina(n21717), .dinb(n21712), .dout(n21718));
  jxor g21537(.dina(n21718), .dinb(n4247), .dout(n21719));
  jxor g21538(.dina(n21719), .dinb(n21711), .dout(n21720));
  jxor g21539(.dina(n21720), .dinb(n21630), .dout(n21721));
  jxor g21540(.dina(n21721), .dinb(n21625), .dout(n21722));
  jxor g21541(.dina(n21722), .dinb(n21616), .dout(n21723));
  jnot g21542(.din(n21723), .dout(n21724));
  jand g21543(.dina(n20781), .dinb(n6936), .dout(n21725));
  jand g21544(.dina(n19525), .dinb(n7741), .dout(n21726));
  jand g21545(.dina(n19527), .dinb(n7613), .dout(n21727));
  jand g21546(.dina(n19529), .dinb(n6934), .dout(n21728));
  jor  g21547(.dina(n21728), .dinb(n21727), .dout(n21729));
  jor  g21548(.dina(n21729), .dinb(n21726), .dout(n21730));
  jor  g21549(.dina(n21730), .dinb(n21725), .dout(n21731));
  jxor g21550(.dina(n21731), .dinb(n5292), .dout(n21732));
  jxor g21551(.dina(n21732), .dinb(n21724), .dout(n21733));
  jxor g21552(.dina(n21733), .dinb(n21613), .dout(n21734));
  jxor g21553(.dina(n21734), .dinb(n21608), .dout(n21735));
  jxor g21554(.dina(n21735), .dinb(n21599), .dout(n21736));
  jnot g21555(.din(n21736), .dout(n21737));
  jxor g21556(.dina(n19658), .dinb(n19657), .dout(n21738));
  jand g21557(.dina(n21738), .dinb(n8771), .dout(n21739));
  jand g21558(.dina(n19513), .dinb(n9491), .dout(n21740));
  jand g21559(.dina(n19515), .dinb(n9126), .dout(n21741));
  jand g21560(.dina(n19517), .dinb(n8769), .dout(n21742));
  jor  g21561(.dina(n21742), .dinb(n21741), .dout(n21743));
  jor  g21562(.dina(n21743), .dinb(n21740), .dout(n21744));
  jor  g21563(.dina(n21744), .dinb(n21739), .dout(n21745));
  jxor g21564(.dina(n21745), .dinb(n6039), .dout(n21746));
  jxor g21565(.dina(n21746), .dinb(n21737), .dout(n21747));
  jxor g21566(.dina(n21747), .dinb(n21596), .dout(n21748));
  jand g21567(.dina(n21748), .dinb(n19769), .dout(n21749));
  jxor g21568(.dina(n19664), .dinb(n19663), .dout(n21750));
  jand g21569(.dina(n21750), .dinb(n67), .dout(n21751));
  jand g21570(.dina(n19510), .dinb(n10827), .dout(n21752));
  jand g21571(.dina(n19511), .dinb(n10350), .dout(n21753));
  jand g21572(.dina(n19513), .dinb(n9917), .dout(n21754));
  jor  g21573(.dina(n21754), .dinb(n21753), .dout(n21755));
  jor  g21574(.dina(n21755), .dinb(n21752), .dout(n21756));
  jor  g21575(.dina(n21756), .dinb(n21751), .dout(n21757));
  jxor g21576(.dina(n21757), .dinb(n64), .dout(n21758));
  jnot g21577(.din(n21758), .dout(n21759));
  jxor g21578(.dina(n21592), .dinb(n21591), .dout(n21760));
  jand g21579(.dina(n21760), .dinb(n21759), .dout(n21761));
  jxor g21580(.dina(n19661), .dinb(n19660), .dout(n21762));
  jand g21581(.dina(n21762), .dinb(n67), .dout(n21763));
  jand g21582(.dina(n19511), .dinb(n10827), .dout(n21764));
  jand g21583(.dina(n19513), .dinb(n10350), .dout(n21765));
  jand g21584(.dina(n19515), .dinb(n9917), .dout(n21766));
  jor  g21585(.dina(n21766), .dinb(n21765), .dout(n21767));
  jor  g21586(.dina(n21767), .dinb(n21764), .dout(n21768));
  jor  g21587(.dina(n21768), .dinb(n21763), .dout(n21769));
  jxor g21588(.dina(n21769), .dinb(n64), .dout(n21770));
  jnot g21589(.din(n21770), .dout(n21771));
  jxor g21590(.dina(n21587), .dinb(n21586), .dout(n21772));
  jand g21591(.dina(n21772), .dinb(n21771), .dout(n21773));
  jxor g21592(.dina(n21584), .dinb(n21583), .dout(n21774));
  jnot g21593(.din(n21774), .dout(n21775));
  jand g21594(.dina(n21738), .dinb(n67), .dout(n21776));
  jand g21595(.dina(n19513), .dinb(n10827), .dout(n21777));
  jand g21596(.dina(n19515), .dinb(n10350), .dout(n21778));
  jand g21597(.dina(n19517), .dinb(n9917), .dout(n21779));
  jor  g21598(.dina(n21779), .dinb(n21778), .dout(n21780));
  jor  g21599(.dina(n21780), .dinb(n21777), .dout(n21781));
  jor  g21600(.dina(n21781), .dinb(n21776), .dout(n21782));
  jxor g21601(.dina(n21782), .dinb(n64), .dout(n21783));
  jor  g21602(.dina(n21783), .dinb(n21775), .dout(n21784));
  jxor g21603(.dina(n21581), .dinb(n21580), .dout(n21785));
  jnot g21604(.din(n21785), .dout(n21786));
  jand g21605(.dina(n21218), .dinb(n67), .dout(n21787));
  jand g21606(.dina(n19515), .dinb(n10827), .dout(n21788));
  jand g21607(.dina(n19517), .dinb(n10350), .dout(n21789));
  jand g21608(.dina(n19519), .dinb(n9917), .dout(n21790));
  jor  g21609(.dina(n21790), .dinb(n21789), .dout(n21791));
  jor  g21610(.dina(n21791), .dinb(n21788), .dout(n21792));
  jor  g21611(.dina(n21792), .dinb(n21787), .dout(n21793));
  jxor g21612(.dina(n21793), .dinb(n64), .dout(n21794));
  jor  g21613(.dina(n21794), .dinb(n21786), .dout(n21795));
  jand g21614(.dina(n21230), .dinb(n67), .dout(n21796));
  jand g21615(.dina(n19517), .dinb(n10827), .dout(n21797));
  jand g21616(.dina(n19519), .dinb(n10350), .dout(n21798));
  jand g21617(.dina(n19521), .dinb(n9917), .dout(n21799));
  jor  g21618(.dina(n21799), .dinb(n21798), .dout(n21800));
  jor  g21619(.dina(n21800), .dinb(n21797), .dout(n21801));
  jor  g21620(.dina(n21801), .dinb(n21796), .dout(n21802));
  jxor g21621(.dina(n21802), .dinb(n64), .dout(n21803));
  jnot g21622(.din(n21803), .dout(n21804));
  jxor g21623(.dina(n21576), .dinb(n21575), .dout(n21805));
  jand g21624(.dina(n21805), .dinb(n21804), .dout(n21806));
  jand g21625(.dina(n21240), .dinb(n67), .dout(n21807));
  jand g21626(.dina(n19519), .dinb(n10827), .dout(n21808));
  jand g21627(.dina(n19521), .dinb(n10350), .dout(n21809));
  jand g21628(.dina(n19523), .dinb(n9917), .dout(n21810));
  jor  g21629(.dina(n21810), .dinb(n21809), .dout(n21811));
  jor  g21630(.dina(n21811), .dinb(n21808), .dout(n21812));
  jor  g21631(.dina(n21812), .dinb(n21807), .dout(n21813));
  jxor g21632(.dina(n21813), .dinb(n64), .dout(n21814));
  jnot g21633(.din(n21814), .dout(n21815));
  jxor g21634(.dina(n21571), .dinb(n21570), .dout(n21816));
  jand g21635(.dina(n21816), .dinb(n21815), .dout(n21817));
  jand g21636(.dina(n21086), .dinb(n67), .dout(n21818));
  jand g21637(.dina(n19521), .dinb(n10827), .dout(n21819));
  jand g21638(.dina(n19523), .dinb(n10350), .dout(n21820));
  jand g21639(.dina(n19525), .dinb(n9917), .dout(n21821));
  jor  g21640(.dina(n21821), .dinb(n21820), .dout(n21822));
  jor  g21641(.dina(n21822), .dinb(n21819), .dout(n21823));
  jor  g21642(.dina(n21823), .dinb(n21818), .dout(n21824));
  jxor g21643(.dina(n21824), .dinb(n64), .dout(n21825));
  jnot g21644(.din(n21825), .dout(n21826));
  jxor g21645(.dina(n21566), .dinb(n21565), .dout(n21827));
  jand g21646(.dina(n21827), .dinb(n21826), .dout(n21828));
  jxor g21647(.dina(n21563), .dinb(n21562), .dout(n21829));
  jnot g21648(.din(n21829), .dout(n21830));
  jand g21649(.dina(n19770), .dinb(n67), .dout(n21831));
  jand g21650(.dina(n19523), .dinb(n10827), .dout(n21832));
  jand g21651(.dina(n19525), .dinb(n10350), .dout(n21833));
  jand g21652(.dina(n19527), .dinb(n9917), .dout(n21834));
  jor  g21653(.dina(n21834), .dinb(n21833), .dout(n21835));
  jor  g21654(.dina(n21835), .dinb(n21832), .dout(n21836));
  jor  g21655(.dina(n21836), .dinb(n21831), .dout(n21837));
  jxor g21656(.dina(n21837), .dinb(n64), .dout(n21838));
  jor  g21657(.dina(n21838), .dinb(n21830), .dout(n21839));
  jxor g21658(.dina(n21560), .dinb(n21559), .dout(n21840));
  jnot g21659(.din(n21840), .dout(n21841));
  jand g21660(.dina(n20781), .dinb(n67), .dout(n21842));
  jand g21661(.dina(n19525), .dinb(n10827), .dout(n21843));
  jand g21662(.dina(n19527), .dinb(n10350), .dout(n21844));
  jand g21663(.dina(n19529), .dinb(n9917), .dout(n21845));
  jor  g21664(.dina(n21845), .dinb(n21844), .dout(n21846));
  jor  g21665(.dina(n21846), .dinb(n21843), .dout(n21847));
  jor  g21666(.dina(n21847), .dinb(n21842), .dout(n21848));
  jxor g21667(.dina(n21848), .dinb(n64), .dout(n21849));
  jor  g21668(.dina(n21849), .dinb(n21841), .dout(n21850));
  jxor g21669(.dina(n21557), .dinb(n21556), .dout(n21851));
  jnot g21670(.din(n21851), .dout(n21852));
  jand g21671(.dina(n20793), .dinb(n67), .dout(n21853));
  jand g21672(.dina(n19527), .dinb(n10827), .dout(n21854));
  jand g21673(.dina(n19529), .dinb(n10350), .dout(n21855));
  jand g21674(.dina(n19531), .dinb(n9917), .dout(n21856));
  jor  g21675(.dina(n21856), .dinb(n21855), .dout(n21857));
  jor  g21676(.dina(n21857), .dinb(n21854), .dout(n21858));
  jor  g21677(.dina(n21858), .dinb(n21853), .dout(n21859));
  jxor g21678(.dina(n21859), .dinb(n64), .dout(n21860));
  jor  g21679(.dina(n21860), .dinb(n21852), .dout(n21861));
  jand g21680(.dina(n20767), .dinb(n67), .dout(n21862));
  jand g21681(.dina(n19529), .dinb(n10827), .dout(n21863));
  jand g21682(.dina(n19531), .dinb(n10350), .dout(n21864));
  jand g21683(.dina(n19533), .dinb(n9917), .dout(n21865));
  jor  g21684(.dina(n21865), .dinb(n21864), .dout(n21866));
  jor  g21685(.dina(n21866), .dinb(n21863), .dout(n21867));
  jor  g21686(.dina(n21867), .dinb(n21862), .dout(n21868));
  jxor g21687(.dina(n21868), .dinb(n64), .dout(n21869));
  jnot g21688(.din(n21869), .dout(n21870));
  jxor g21689(.dina(n21552), .dinb(n21551), .dout(n21871));
  jand g21690(.dina(n21871), .dinb(n21870), .dout(n21872));
  jand g21691(.dina(n19780), .dinb(n67), .dout(n21873));
  jand g21692(.dina(n19531), .dinb(n10827), .dout(n21874));
  jand g21693(.dina(n19533), .dinb(n10350), .dout(n21875));
  jand g21694(.dina(n19535), .dinb(n9917), .dout(n21876));
  jor  g21695(.dina(n21876), .dinb(n21875), .dout(n21877));
  jor  g21696(.dina(n21877), .dinb(n21874), .dout(n21878));
  jor  g21697(.dina(n21878), .dinb(n21873), .dout(n21879));
  jxor g21698(.dina(n21879), .dinb(n64), .dout(n21880));
  jnot g21699(.din(n21880), .dout(n21881));
  jxor g21700(.dina(n21547), .dinb(n21546), .dout(n21882));
  jand g21701(.dina(n21882), .dinb(n21881), .dout(n21883));
  jand g21702(.dina(n20399), .dinb(n67), .dout(n21884));
  jand g21703(.dina(n19533), .dinb(n10827), .dout(n21885));
  jand g21704(.dina(n19535), .dinb(n10350), .dout(n21886));
  jand g21705(.dina(n19537), .dinb(n9917), .dout(n21887));
  jor  g21706(.dina(n21887), .dinb(n21886), .dout(n21888));
  jor  g21707(.dina(n21888), .dinb(n21885), .dout(n21889));
  jor  g21708(.dina(n21889), .dinb(n21884), .dout(n21890));
  jxor g21709(.dina(n21890), .dinb(n64), .dout(n21891));
  jnot g21710(.din(n21891), .dout(n21892));
  jxor g21711(.dina(n21542), .dinb(n21541), .dout(n21893));
  jand g21712(.dina(n21893), .dinb(n21892), .dout(n21894));
  jxor g21713(.dina(n21539), .dinb(n21538), .dout(n21895));
  jnot g21714(.din(n21895), .dout(n21896));
  jand g21715(.dina(n20413), .dinb(n67), .dout(n21897));
  jand g21716(.dina(n19535), .dinb(n10827), .dout(n21898));
  jand g21717(.dina(n19537), .dinb(n10350), .dout(n21899));
  jand g21718(.dina(n19539), .dinb(n9917), .dout(n21900));
  jor  g21719(.dina(n21900), .dinb(n21899), .dout(n21901));
  jor  g21720(.dina(n21901), .dinb(n21898), .dout(n21902));
  jor  g21721(.dina(n21902), .dinb(n21897), .dout(n21903));
  jxor g21722(.dina(n21903), .dinb(n64), .dout(n21904));
  jor  g21723(.dina(n21904), .dinb(n21896), .dout(n21905));
  jxor g21724(.dina(n21536), .dinb(n21535), .dout(n21906));
  jnot g21725(.din(n21906), .dout(n21907));
  jand g21726(.dina(n20387), .dinb(n67), .dout(n21908));
  jand g21727(.dina(n19537), .dinb(n10827), .dout(n21909));
  jand g21728(.dina(n19539), .dinb(n10350), .dout(n21910));
  jand g21729(.dina(n19541), .dinb(n9917), .dout(n21911));
  jor  g21730(.dina(n21911), .dinb(n21910), .dout(n21912));
  jor  g21731(.dina(n21912), .dinb(n21909), .dout(n21913));
  jor  g21732(.dina(n21913), .dinb(n21908), .dout(n21914));
  jxor g21733(.dina(n21914), .dinb(n64), .dout(n21915));
  jor  g21734(.dina(n21915), .dinb(n21907), .dout(n21916));
  jxor g21735(.dina(n21533), .dinb(n21532), .dout(n21917));
  jnot g21736(.din(n21917), .dout(n21918));
  jand g21737(.dina(n20131), .dinb(n67), .dout(n21919));
  jand g21738(.dina(n19539), .dinb(n10827), .dout(n21920));
  jand g21739(.dina(n19541), .dinb(n10350), .dout(n21921));
  jand g21740(.dina(n19543), .dinb(n9917), .dout(n21922));
  jor  g21741(.dina(n21922), .dinb(n21921), .dout(n21923));
  jor  g21742(.dina(n21923), .dinb(n21920), .dout(n21924));
  jor  g21743(.dina(n21924), .dinb(n21919), .dout(n21925));
  jxor g21744(.dina(n21925), .dinb(n64), .dout(n21926));
  jor  g21745(.dina(n21926), .dinb(n21918), .dout(n21927));
  jand g21746(.dina(n20141), .dinb(n67), .dout(n21928));
  jand g21747(.dina(n19541), .dinb(n10827), .dout(n21929));
  jand g21748(.dina(n19543), .dinb(n10350), .dout(n21930));
  jand g21749(.dina(n19545), .dinb(n9917), .dout(n21931));
  jor  g21750(.dina(n21931), .dinb(n21930), .dout(n21932));
  jor  g21751(.dina(n21932), .dinb(n21929), .dout(n21933));
  jor  g21752(.dina(n21933), .dinb(n21928), .dout(n21934));
  jxor g21753(.dina(n21934), .dinb(n64), .dout(n21935));
  jnot g21754(.din(n21935), .dout(n21936));
  jxor g21755(.dina(n21528), .dinb(n21527), .dout(n21937));
  jand g21756(.dina(n21937), .dinb(n21936), .dout(n21938));
  jand g21757(.dina(n20153), .dinb(n67), .dout(n21939));
  jand g21758(.dina(n19543), .dinb(n10827), .dout(n21940));
  jand g21759(.dina(n19545), .dinb(n10350), .dout(n21941));
  jand g21760(.dina(n19548), .dinb(n9917), .dout(n21942));
  jor  g21761(.dina(n21942), .dinb(n21941), .dout(n21943));
  jor  g21762(.dina(n21943), .dinb(n21940), .dout(n21944));
  jor  g21763(.dina(n21944), .dinb(n21939), .dout(n21945));
  jxor g21764(.dina(n21945), .dinb(n64), .dout(n21946));
  jnot g21765(.din(n21946), .dout(n21947));
  jxor g21766(.dina(n21523), .dinb(n21522), .dout(n21948));
  jand g21767(.dina(n21948), .dinb(n21947), .dout(n21949));
  jand g21768(.dina(n20079), .dinb(n67), .dout(n21950));
  jand g21769(.dina(n19545), .dinb(n10827), .dout(n21951));
  jand g21770(.dina(n19548), .dinb(n10350), .dout(n21952));
  jand g21771(.dina(n19551), .dinb(n9917), .dout(n21953));
  jor  g21772(.dina(n21953), .dinb(n21952), .dout(n21954));
  jor  g21773(.dina(n21954), .dinb(n21951), .dout(n21955));
  jor  g21774(.dina(n21955), .dinb(n21950), .dout(n21956));
  jxor g21775(.dina(n21956), .dinb(n64), .dout(n21957));
  jnot g21776(.din(n21957), .dout(n21958));
  jxor g21777(.dina(n21518), .dinb(n21517), .dout(n21959));
  jand g21778(.dina(n21959), .dinb(n21958), .dout(n21960));
  jxor g21779(.dina(n21515), .dinb(n21514), .dout(n21961));
  jnot g21780(.din(n21961), .dout(n21962));
  jor  g21781(.dina(n19940), .dinb(n9919), .dout(n21963));
  jor  g21782(.dina(n19547), .dinb(n10826), .dout(n21964));
  jor  g21783(.dina(n19550), .dinb(n10351), .dout(n21965));
  jor  g21784(.dina(n19553), .dinb(n9918), .dout(n21966));
  jand g21785(.dina(n21966), .dinb(n21965), .dout(n21967));
  jand g21786(.dina(n21967), .dinb(n21964), .dout(n21968));
  jand g21787(.dina(n21968), .dinb(n21963), .dout(n21969));
  jxor g21788(.dina(n21969), .dinb(\a[5] ), .dout(n21970));
  jor  g21789(.dina(n21970), .dinb(n21962), .dout(n21971));
  jxor g21790(.dina(n21512), .dinb(n21511), .dout(n21972));
  jnot g21791(.din(n21972), .dout(n21973));
  jor  g21792(.dina(n19952), .dinb(n9919), .dout(n21974));
  jor  g21793(.dina(n19550), .dinb(n10826), .dout(n21975));
  jor  g21794(.dina(n19553), .dinb(n10351), .dout(n21976));
  jor  g21795(.dina(n19558), .dinb(n9918), .dout(n21977));
  jand g21796(.dina(n21977), .dinb(n21976), .dout(n21978));
  jand g21797(.dina(n21978), .dinb(n21975), .dout(n21979));
  jand g21798(.dina(n21979), .dinb(n21974), .dout(n21980));
  jxor g21799(.dina(n21980), .dinb(\a[5] ), .dout(n21981));
  jor  g21800(.dina(n21981), .dinb(n21973), .dout(n21982));
  jxor g21801(.dina(n21509), .dinb(n21508), .dout(n21983));
  jnot g21802(.din(n21983), .dout(n21984));
  jor  g21803(.dina(n19964), .dinb(n9919), .dout(n21985));
  jor  g21804(.dina(n19553), .dinb(n10826), .dout(n21986));
  jor  g21805(.dina(n19558), .dinb(n10351), .dout(n21987));
  jor  g21806(.dina(n19562), .dinb(n9918), .dout(n21988));
  jand g21807(.dina(n21988), .dinb(n21987), .dout(n21989));
  jand g21808(.dina(n21989), .dinb(n21986), .dout(n21990));
  jand g21809(.dina(n21990), .dinb(n21985), .dout(n21991));
  jxor g21810(.dina(n21991), .dinb(\a[5] ), .dout(n21992));
  jor  g21811(.dina(n21992), .dinb(n21984), .dout(n21993));
  jor  g21812(.dina(n19906), .dinb(n9919), .dout(n21994));
  jor  g21813(.dina(n19558), .dinb(n10826), .dout(n21995));
  jor  g21814(.dina(n19562), .dinb(n10351), .dout(n21996));
  jor  g21815(.dina(n19564), .dinb(n9918), .dout(n21997));
  jand g21816(.dina(n21997), .dinb(n21996), .dout(n21998));
  jand g21817(.dina(n21998), .dinb(n21995), .dout(n21999));
  jand g21818(.dina(n21999), .dinb(n21994), .dout(n22000));
  jxor g21819(.dina(n22000), .dinb(\a[5] ), .dout(n22001));
  jnot g21820(.din(n22001), .dout(n22002));
  jxor g21821(.dina(n21506), .dinb(n21505), .dout(n22003));
  jand g21822(.dina(n22003), .dinb(n22002), .dout(n22004));
  jor  g21823(.dina(n19790), .dinb(n9919), .dout(n22005));
  jor  g21824(.dina(n19562), .dinb(n10826), .dout(n22006));
  jor  g21825(.dina(n19564), .dinb(n10351), .dout(n22007));
  jor  g21826(.dina(n19566), .dinb(n9918), .dout(n22008));
  jand g21827(.dina(n22008), .dinb(n22007), .dout(n22009));
  jand g21828(.dina(n22009), .dinb(n22006), .dout(n22010));
  jand g21829(.dina(n22010), .dinb(n22005), .dout(n22011));
  jxor g21830(.dina(n22011), .dinb(\a[5] ), .dout(n22012));
  jnot g21831(.din(n22012), .dout(n22013));
  jxor g21832(.dina(n21503), .dinb(n21502), .dout(n22014));
  jand g21833(.dina(n22014), .dinb(n22013), .dout(n22015));
  jor  g21834(.dina(n19839), .dinb(n9919), .dout(n22016));
  jor  g21835(.dina(n19564), .dinb(n10826), .dout(n22017));
  jor  g21836(.dina(n19566), .dinb(n10351), .dout(n22018));
  jor  g21837(.dina(n19568), .dinb(n9918), .dout(n22019));
  jand g21838(.dina(n22019), .dinb(n22018), .dout(n22020));
  jand g21839(.dina(n22020), .dinb(n22017), .dout(n22021));
  jand g21840(.dina(n22021), .dinb(n22016), .dout(n22022));
  jxor g21841(.dina(n22022), .dinb(\a[5] ), .dout(n22023));
  jnot g21842(.din(n22023), .dout(n22024));
  jor  g21843(.dina(n21483), .dinb(n6039), .dout(n22025));
  jxor g21844(.dina(n22025), .dinb(n21491), .dout(n22026));
  jand g21845(.dina(n22026), .dinb(n22024), .dout(n22027));
  jor  g21846(.dina(n19852), .dinb(n9919), .dout(n22028));
  jor  g21847(.dina(n19566), .dinb(n10826), .dout(n22029));
  jor  g21848(.dina(n19568), .dinb(n10351), .dout(n22030));
  jor  g21849(.dina(n19570), .dinb(n9918), .dout(n22031));
  jand g21850(.dina(n22031), .dinb(n22030), .dout(n22032));
  jand g21851(.dina(n22032), .dinb(n22029), .dout(n22033));
  jand g21852(.dina(n22033), .dinb(n22028), .dout(n22034));
  jxor g21853(.dina(n22034), .dinb(\a[5] ), .dout(n22035));
  jnot g21854(.din(n22035), .dout(n22036));
  jand g21855(.dina(n21480), .dinb(\a[8] ), .dout(n22037));
  jxor g21856(.dina(n22037), .dinb(n21478), .dout(n22038));
  jand g21857(.dina(n22038), .dinb(n22036), .dout(n22039));
  jand g21858(.dina(n19813), .dinb(n67), .dout(n22040));
  jand g21859(.dina(n19576), .dinb(n10350), .dout(n22041));
  jand g21860(.dina(n19574), .dinb(n10827), .dout(n22042));
  jor  g21861(.dina(n22042), .dinb(n22041), .dout(n22043));
  jor  g21862(.dina(n22043), .dinb(n22040), .dout(n22044));
  jnot g21863(.din(n22044), .dout(n22045));
  jand g21864(.dina(n19576), .dinb(n65), .dout(n22046));
  jnot g21865(.din(n22046), .dout(n22047));
  jand g21866(.dina(n22047), .dinb(\a[5] ), .dout(n22048));
  jand g21867(.dina(n22048), .dinb(n22045), .dout(n22049));
  jand g21868(.dina(n19826), .dinb(n67), .dout(n22050));
  jand g21869(.dina(n19572), .dinb(n10827), .dout(n22051));
  jand g21870(.dina(n19574), .dinb(n10350), .dout(n22052));
  jand g21871(.dina(n19576), .dinb(n9917), .dout(n22053));
  jor  g21872(.dina(n22053), .dinb(n22052), .dout(n22054));
  jor  g21873(.dina(n22054), .dinb(n22051), .dout(n22055));
  jor  g21874(.dina(n22055), .dinb(n22050), .dout(n22056));
  jnot g21875(.din(n22056), .dout(n22057));
  jand g21876(.dina(n22057), .dinb(n22049), .dout(n22058));
  jand g21877(.dina(n22058), .dinb(n21480), .dout(n22059));
  jor  g21878(.dina(n19801), .dinb(n9919), .dout(n22060));
  jor  g21879(.dina(n19568), .dinb(n10826), .dout(n22061));
  jor  g21880(.dina(n19570), .dinb(n10351), .dout(n22062));
  jor  g21881(.dina(n19575), .dinb(n9918), .dout(n22063));
  jand g21882(.dina(n22063), .dinb(n22062), .dout(n22064));
  jand g21883(.dina(n22064), .dinb(n22061), .dout(n22065));
  jand g21884(.dina(n22065), .dinb(n22060), .dout(n22066));
  jxor g21885(.dina(n22066), .dinb(\a[5] ), .dout(n22067));
  jnot g21886(.din(n22067), .dout(n22068));
  jxor g21887(.dina(n22058), .dinb(n21480), .dout(n22069));
  jand g21888(.dina(n22069), .dinb(n22068), .dout(n22070));
  jor  g21889(.dina(n22070), .dinb(n22059), .dout(n22071));
  jxor g21890(.dina(n22038), .dinb(n22036), .dout(n22072));
  jand g21891(.dina(n22072), .dinb(n22071), .dout(n22073));
  jor  g21892(.dina(n22073), .dinb(n22039), .dout(n22074));
  jxor g21893(.dina(n22026), .dinb(n22024), .dout(n22075));
  jand g21894(.dina(n22075), .dinb(n22074), .dout(n22076));
  jor  g21895(.dina(n22076), .dinb(n22027), .dout(n22077));
  jxor g21896(.dina(n22014), .dinb(n22013), .dout(n22078));
  jand g21897(.dina(n22078), .dinb(n22077), .dout(n22079));
  jor  g21898(.dina(n22079), .dinb(n22015), .dout(n22080));
  jxor g21899(.dina(n22003), .dinb(n22002), .dout(n22081));
  jand g21900(.dina(n22081), .dinb(n22080), .dout(n22082));
  jor  g21901(.dina(n22082), .dinb(n22004), .dout(n22083));
  jxor g21902(.dina(n21992), .dinb(n21984), .dout(n22084));
  jand g21903(.dina(n22084), .dinb(n22083), .dout(n22085));
  jnot g21904(.din(n22085), .dout(n22086));
  jand g21905(.dina(n22086), .dinb(n21993), .dout(n22087));
  jnot g21906(.din(n22087), .dout(n22088));
  jxor g21907(.dina(n21981), .dinb(n21973), .dout(n22089));
  jand g21908(.dina(n22089), .dinb(n22088), .dout(n22090));
  jnot g21909(.din(n22090), .dout(n22091));
  jand g21910(.dina(n22091), .dinb(n21982), .dout(n22092));
  jnot g21911(.din(n22092), .dout(n22093));
  jxor g21912(.dina(n21970), .dinb(n21962), .dout(n22094));
  jand g21913(.dina(n22094), .dinb(n22093), .dout(n22095));
  jnot g21914(.din(n22095), .dout(n22096));
  jand g21915(.dina(n22096), .dinb(n21971), .dout(n22097));
  jnot g21916(.din(n22097), .dout(n22098));
  jxor g21917(.dina(n21959), .dinb(n21958), .dout(n22099));
  jand g21918(.dina(n22099), .dinb(n22098), .dout(n22100));
  jor  g21919(.dina(n22100), .dinb(n21960), .dout(n22101));
  jxor g21920(.dina(n21948), .dinb(n21947), .dout(n22102));
  jand g21921(.dina(n22102), .dinb(n22101), .dout(n22103));
  jor  g21922(.dina(n22103), .dinb(n21949), .dout(n22104));
  jxor g21923(.dina(n21937), .dinb(n21936), .dout(n22105));
  jand g21924(.dina(n22105), .dinb(n22104), .dout(n22106));
  jor  g21925(.dina(n22106), .dinb(n21938), .dout(n22107));
  jxor g21926(.dina(n21926), .dinb(n21918), .dout(n22108));
  jand g21927(.dina(n22108), .dinb(n22107), .dout(n22109));
  jnot g21928(.din(n22109), .dout(n22110));
  jand g21929(.dina(n22110), .dinb(n21927), .dout(n22111));
  jnot g21930(.din(n22111), .dout(n22112));
  jxor g21931(.dina(n21915), .dinb(n21907), .dout(n22113));
  jand g21932(.dina(n22113), .dinb(n22112), .dout(n22114));
  jnot g21933(.din(n22114), .dout(n22115));
  jand g21934(.dina(n22115), .dinb(n21916), .dout(n22116));
  jnot g21935(.din(n22116), .dout(n22117));
  jxor g21936(.dina(n21904), .dinb(n21896), .dout(n22118));
  jand g21937(.dina(n22118), .dinb(n22117), .dout(n22119));
  jnot g21938(.din(n22119), .dout(n22120));
  jand g21939(.dina(n22120), .dinb(n21905), .dout(n22121));
  jnot g21940(.din(n22121), .dout(n22122));
  jxor g21941(.dina(n21893), .dinb(n21892), .dout(n22123));
  jand g21942(.dina(n22123), .dinb(n22122), .dout(n22124));
  jor  g21943(.dina(n22124), .dinb(n21894), .dout(n22125));
  jxor g21944(.dina(n21882), .dinb(n21881), .dout(n22126));
  jand g21945(.dina(n22126), .dinb(n22125), .dout(n22127));
  jor  g21946(.dina(n22127), .dinb(n21883), .dout(n22128));
  jxor g21947(.dina(n21871), .dinb(n21870), .dout(n22129));
  jand g21948(.dina(n22129), .dinb(n22128), .dout(n22130));
  jor  g21949(.dina(n22130), .dinb(n21872), .dout(n22131));
  jxor g21950(.dina(n21860), .dinb(n21852), .dout(n22132));
  jand g21951(.dina(n22132), .dinb(n22131), .dout(n22133));
  jnot g21952(.din(n22133), .dout(n22134));
  jand g21953(.dina(n22134), .dinb(n21861), .dout(n22135));
  jnot g21954(.din(n22135), .dout(n22136));
  jxor g21955(.dina(n21849), .dinb(n21841), .dout(n22137));
  jand g21956(.dina(n22137), .dinb(n22136), .dout(n22138));
  jnot g21957(.din(n22138), .dout(n22139));
  jand g21958(.dina(n22139), .dinb(n21850), .dout(n22140));
  jnot g21959(.din(n22140), .dout(n22141));
  jxor g21960(.dina(n21838), .dinb(n21830), .dout(n22142));
  jand g21961(.dina(n22142), .dinb(n22141), .dout(n22143));
  jnot g21962(.din(n22143), .dout(n22144));
  jand g21963(.dina(n22144), .dinb(n21839), .dout(n22145));
  jnot g21964(.din(n22145), .dout(n22146));
  jxor g21965(.dina(n21827), .dinb(n21826), .dout(n22147));
  jand g21966(.dina(n22147), .dinb(n22146), .dout(n22148));
  jor  g21967(.dina(n22148), .dinb(n21828), .dout(n22149));
  jxor g21968(.dina(n21816), .dinb(n21815), .dout(n22150));
  jand g21969(.dina(n22150), .dinb(n22149), .dout(n22151));
  jor  g21970(.dina(n22151), .dinb(n21817), .dout(n22152));
  jxor g21971(.dina(n21805), .dinb(n21804), .dout(n22153));
  jand g21972(.dina(n22153), .dinb(n22152), .dout(n22154));
  jor  g21973(.dina(n22154), .dinb(n21806), .dout(n22155));
  jxor g21974(.dina(n21794), .dinb(n21786), .dout(n22156));
  jand g21975(.dina(n22156), .dinb(n22155), .dout(n22157));
  jnot g21976(.din(n22157), .dout(n22158));
  jand g21977(.dina(n22158), .dinb(n21795), .dout(n22159));
  jnot g21978(.din(n22159), .dout(n22160));
  jxor g21979(.dina(n21783), .dinb(n21775), .dout(n22161));
  jand g21980(.dina(n22161), .dinb(n22160), .dout(n22162));
  jnot g21981(.din(n22162), .dout(n22163));
  jand g21982(.dina(n22163), .dinb(n21784), .dout(n22164));
  jnot g21983(.din(n22164), .dout(n22165));
  jxor g21984(.dina(n21772), .dinb(n21771), .dout(n22166));
  jand g21985(.dina(n22166), .dinb(n22165), .dout(n22167));
  jor  g21986(.dina(n22167), .dinb(n21773), .dout(n22168));
  jxor g21987(.dina(n21760), .dinb(n21759), .dout(n22169));
  jand g21988(.dina(n22169), .dinb(n22168), .dout(n22170));
  jor  g21989(.dina(n22170), .dinb(n21761), .dout(n22171));
  jxor g21990(.dina(n21748), .dinb(n19769), .dout(n22172));
  jand g21991(.dina(n22172), .dinb(n22171), .dout(n22173));
  jor  g21992(.dina(n22173), .dinb(n21749), .dout(n22174));
  jand g21993(.dina(n19758), .dinb(n19510), .dout(n22175));
  jand g21994(.dina(n19759), .dinb(n19666), .dout(n22176));
  jor  g21995(.dina(n22176), .dinb(n22175), .dout(n22177));
  jand g21996(.dina(n19753), .dinb(n19746), .dout(n22178));
  jand g21997(.dina(n19757), .dinb(n19754), .dout(n22179));
  jor  g21998(.dina(n22179), .dinb(n22178), .dout(n22180));
  jand g21999(.dina(n13022), .dinb(n75), .dout(n22181));
  jand g22000(.dina(n12815), .dinb(n4918), .dout(n22183));
  jand g22001(.dina(n12795), .dinb(n4745), .dout(n22184));
  jor  g22002(.dina(n22184), .dinb(n22183), .dout(n22185));
  jor  g22003(.dina(n22185), .dinb(n4933), .dout(n22186));
  jor  g22004(.dina(n22186), .dinb(n22181), .dout(n22187));
  jxor g22005(.dina(n22187), .dinb(n68), .dout(n22188));
  jnot g22006(.din(n22188), .dout(n22189));
  jor  g22007(.dina(n19734), .dinb(n19686), .dout(n22190));
  jand g22008(.dina(n19734), .dinb(n19686), .dout(n22191));
  jor  g22009(.dina(n19744), .dinb(n22191), .dout(n22192));
  jand g22010(.dina(n22192), .dinb(n22190), .dout(n22193));
  jxor g22011(.dina(n22193), .dinb(n22189), .dout(n22194));
  jand g22012(.dina(n19732), .dinb(n19725), .dout(n22195));
  jand g22013(.dina(n19733), .dinb(n19695), .dout(n22196));
  jor  g22014(.dina(n22196), .dinb(n22195), .dout(n22197));
  jand g22015(.dina(n19723), .dinb(n19475), .dout(n22198));
  jand g22016(.dina(n19724), .dinb(n19700), .dout(n22199));
  jor  g22017(.dina(n22199), .dinb(n22198), .dout(n22200));
  jnot g22018(.din(n5362), .dout(n22201));
  jor  g22019(.dina(n22201), .dinb(n5357), .dout(n22202));
  jxor g22020(.dina(n22202), .dinb(n72), .dout(n22204));
  jand g22021(.dina(n515), .dinb(n197), .dout(n22205));
  jand g22022(.dina(n427), .dinb(n383), .dout(n22206));
  jand g22023(.dina(n22206), .dinb(n22205), .dout(n22207));
  jand g22024(.dina(n7161), .dinb(n1082), .dout(n22208));
  jand g22025(.dina(n22208), .dinb(n22207), .dout(n22209));
  jand g22026(.dina(n22209), .dinb(n7055), .dout(n22210));
  jand g22027(.dina(n2580), .dinb(n827), .dout(n22211));
  jand g22028(.dina(n4084), .dinb(n982), .dout(n22212));
  jand g22029(.dina(n22212), .dinb(n22211), .dout(n22213));
  jand g22030(.dina(n22213), .dinb(n3791), .dout(n22214));
  jand g22031(.dina(n22214), .dinb(n22210), .dout(n22215));
  jand g22032(.dina(n22215), .dinb(n14516), .dout(n22216));
  jand g22033(.dina(n13217), .dinb(n5548), .dout(n22217));
  jand g22034(.dina(n22217), .dinb(n22216), .dout(n22218));
  jand g22035(.dina(n22218), .dinb(n12217), .dout(n22219));
  jxor g22036(.dina(n22219), .dinb(n19723), .dout(n22220));
  jxor g22037(.dina(n22220), .dinb(n22204), .dout(n22221));
  jxor g22038(.dina(n22221), .dinb(n22200), .dout(n22222));
  jand g22039(.dina(n12179), .dinb(n732), .dout(n22223));
  jand g22040(.dina(n12177), .dinb(n3855), .dout(n22224));
  jand g22041(.dina(n11941), .dinb(n3858), .dout(n22225));
  jand g22042(.dina(n11942), .dinb(n3851), .dout(n22226));
  jor  g22043(.dina(n22226), .dinb(n22225), .dout(n22227));
  jor  g22044(.dina(n22227), .dinb(n22224), .dout(n22228));
  jor  g22045(.dina(n22228), .dinb(n22223), .dout(n22229));
  jxor g22046(.dina(n22229), .dinb(n22222), .dout(n22230));
  jxor g22047(.dina(n22230), .dinb(n22197), .dout(n22231));
  jand g22048(.dina(n12938), .dinb(n4449), .dout(n22232));
  jand g22049(.dina(n12782), .dinb(n4453), .dout(n22233));
  jand g22050(.dina(n12783), .dinb(n4457), .dout(n22234));
  jand g22051(.dina(n12766), .dinb(n4461), .dout(n22235));
  jor  g22052(.dina(n22235), .dinb(n22234), .dout(n22236));
  jor  g22053(.dina(n22236), .dinb(n22233), .dout(n22237));
  jor  g22054(.dina(n22237), .dinb(n22232), .dout(n22238));
  jxor g22055(.dina(n22238), .dinb(n88), .dout(n22239));
  jnot g22056(.din(n22239), .dout(n22240));
  jxor g22057(.dina(n22240), .dinb(n22231), .dout(n22241));
  jxor g22058(.dina(n22241), .dinb(n22194), .dout(n22242));
  jor  g22059(.dina(n19680), .dinb(n19674), .dout(n22243));
  jand g22060(.dina(n19680), .dinb(n19674), .dout(n22244));
  jor  g22061(.dina(n19745), .dinb(n22244), .dout(n22245));
  jand g22062(.dina(n22245), .dinb(n22243), .dout(n22246));
  jxor g22063(.dina(n22246), .dinb(n22242), .dout(n22247));
  jxor g22064(.dina(n22247), .dinb(n22180), .dout(n22248));
  jxor g22065(.dina(n22248), .dinb(n19758), .dout(n22249));
  jxor g22066(.dina(n22249), .dinb(n22177), .dout(n22250));
  jand g22067(.dina(n22250), .dinb(n67), .dout(n22251));
  jand g22068(.dina(n22248), .dinb(n10827), .dout(n22252));
  jand g22069(.dina(n19758), .dinb(n10350), .dout(n22253));
  jand g22070(.dina(n19510), .dinb(n9917), .dout(n22254));
  jor  g22071(.dina(n22254), .dinb(n22253), .dout(n22255));
  jor  g22072(.dina(n22255), .dinb(n22252), .dout(n22256));
  jor  g22073(.dina(n22256), .dinb(n22251), .dout(n22257));
  jxor g22074(.dina(n22257), .dinb(n64), .dout(n22258));
  jnot g22075(.din(n22258), .dout(n22259));
  jor  g22076(.dina(n21746), .dinb(n21737), .dout(n22260));
  jand g22077(.dina(n21747), .dinb(n21596), .dout(n22261));
  jnot g22078(.din(n22261), .dout(n22262));
  jand g22079(.dina(n22262), .dinb(n22260), .dout(n22263));
  jnot g22080(.din(n22263), .dout(n22264));
  jand g22081(.dina(n21734), .dinb(n21608), .dout(n22265));
  jand g22082(.dina(n21735), .dinb(n21599), .dout(n22266));
  jor  g22083(.dina(n22266), .dinb(n22265), .dout(n22267));
  jand g22084(.dina(n21230), .dinb(n7890), .dout(n22268));
  jand g22085(.dina(n19517), .dinb(n8441), .dout(n22269));
  jand g22086(.dina(n19519), .dinb(n8154), .dout(n22270));
  jand g22087(.dina(n19521), .dinb(n7888), .dout(n22271));
  jor  g22088(.dina(n22271), .dinb(n22270), .dout(n22272));
  jor  g22089(.dina(n22272), .dinb(n22269), .dout(n22273));
  jor  g22090(.dina(n22273), .dinb(n22268), .dout(n22274));
  jxor g22091(.dina(n22274), .dinb(n5833), .dout(n22275));
  jnot g22092(.din(n22275), .dout(n22276));
  jor  g22093(.dina(n21732), .dinb(n21724), .dout(n22277));
  jand g22094(.dina(n21733), .dinb(n21613), .dout(n22278));
  jnot g22095(.din(n22278), .dout(n22279));
  jand g22096(.dina(n22279), .dinb(n22277), .dout(n22280));
  jnot g22097(.din(n22280), .dout(n22281));
  jand g22098(.dina(n21721), .dinb(n21625), .dout(n22282));
  jand g22099(.dina(n21722), .dinb(n21616), .dout(n22283));
  jor  g22100(.dina(n22283), .dinb(n22282), .dout(n22284));
  jand g22101(.dina(n20767), .dinb(n6340), .dout(n22285));
  jand g22102(.dina(n19529), .dinb(n6798), .dout(n22286));
  jand g22103(.dina(n19531), .dinb(n6556), .dout(n22287));
  jand g22104(.dina(n19533), .dinb(n6338), .dout(n22288));
  jor  g22105(.dina(n22288), .dinb(n22287), .dout(n22289));
  jor  g22106(.dina(n22289), .dinb(n22286), .dout(n22290));
  jor  g22107(.dina(n22290), .dinb(n22285), .dout(n22291));
  jxor g22108(.dina(n22291), .dinb(n5064), .dout(n22292));
  jnot g22109(.din(n22292), .dout(n22293));
  jor  g22110(.dina(n21719), .dinb(n21711), .dout(n22294));
  jand g22111(.dina(n21720), .dinb(n21630), .dout(n22295));
  jnot g22112(.din(n22295), .dout(n22296));
  jand g22113(.dina(n22296), .dinb(n22294), .dout(n22297));
  jnot g22114(.din(n22297), .dout(n22298));
  jand g22115(.dina(n21708), .dinb(n21642), .dout(n22299));
  jand g22116(.dina(n21709), .dinb(n21633), .dout(n22300));
  jor  g22117(.dina(n22300), .dinb(n22299), .dout(n22301));
  jand g22118(.dina(n20141), .dinb(n5365), .dout(n22302));
  jand g22119(.dina(n19541), .dinb(n5500), .dout(n22303));
  jand g22120(.dina(n19543), .dinb(n5424), .dout(n22304));
  jand g22121(.dina(n19545), .dinb(n5363), .dout(n22305));
  jor  g22122(.dina(n22305), .dinb(n22304), .dout(n22306));
  jor  g22123(.dina(n22306), .dinb(n22303), .dout(n22307));
  jor  g22124(.dina(n22307), .dinb(n22302), .dout(n22308));
  jxor g22125(.dina(n22308), .dinb(n72), .dout(n22309));
  jnot g22126(.din(n22309), .dout(n22310));
  jor  g22127(.dina(n21706), .dinb(n21698), .dout(n22311));
  jand g22128(.dina(n21707), .dinb(n21647), .dout(n22312));
  jnot g22129(.din(n22312), .dout(n22313));
  jand g22130(.dina(n22313), .dinb(n22311), .dout(n22314));
  jnot g22131(.din(n22314), .dout(n22315));
  jand g22132(.dina(n21695), .dinb(n21659), .dout(n22316));
  jand g22133(.dina(n21696), .dinb(n21650), .dout(n22317));
  jor  g22134(.dina(n22317), .dinb(n22316), .dout(n22318));
  jor  g22135(.dina(n19906), .dinb(n4724), .dout(n22319));
  jor  g22136(.dina(n19558), .dinb(n4905), .dout(n22320));
  jor  g22137(.dina(n19562), .dinb(n4735), .dout(n22321));
  jor  g22138(.dina(n19564), .dinb(n4733), .dout(n22322));
  jand g22139(.dina(n22322), .dinb(n22321), .dout(n22323));
  jand g22140(.dina(n22323), .dinb(n22320), .dout(n22324));
  jand g22141(.dina(n22324), .dinb(n22319), .dout(n22325));
  jxor g22142(.dina(n22325), .dinb(\a[29] ), .dout(n22326));
  jnot g22143(.din(n22326), .dout(n22327));
  jand g22144(.dina(n21693), .dinb(n21684), .dout(n22328));
  jand g22145(.dina(n21694), .dinb(n21665), .dout(n22329));
  jor  g22146(.dina(n22329), .dinb(n22328), .dout(n22330));
  jand g22147(.dina(n1264), .dinb(n382), .dout(n22331));
  jand g22148(.dina(n22331), .dinb(n536), .dout(n22332));
  jand g22149(.dina(n805), .dinb(n716), .dout(n22333));
  jand g22150(.dina(n22333), .dinb(n473), .dout(n22334));
  jand g22151(.dina(n22334), .dinb(n22332), .dout(n22335));
  jand g22152(.dina(n6378), .dinb(n1050), .dout(n22336));
  jand g22153(.dina(n22336), .dinb(n22335), .dout(n22337));
  jand g22154(.dina(n5153), .dinb(n1598), .dout(n22338));
  jand g22155(.dina(n22338), .dinb(n833), .dout(n22339));
  jand g22156(.dina(n22339), .dinb(n12725), .dout(n22340));
  jand g22157(.dina(n22340), .dinb(n22337), .dout(n22341));
  jand g22158(.dina(n22341), .dinb(n12702), .dout(n22342));
  jand g22159(.dina(n22342), .dinb(n19709), .dout(n22343));
  jand g22160(.dina(n22343), .dinb(n14377), .dout(n22344));
  jor  g22161(.dina(n19852), .dinb(n6463), .dout(n22345));
  jnot g22162(.din(n19566), .dout(n22346));
  jand g22163(.dina(n22346), .dinb(n3855), .dout(n22347));
  jand g22164(.dina(n19572), .dinb(n3851), .dout(n22348));
  jand g22165(.dina(n21687), .dinb(n3858), .dout(n22349));
  jor  g22166(.dina(n22349), .dinb(n22348), .dout(n22350));
  jor  g22167(.dina(n22350), .dinb(n22347), .dout(n22351));
  jnot g22168(.din(n22351), .dout(n22352));
  jand g22169(.dina(n22352), .dinb(n22345), .dout(n22353));
  jxor g22170(.dina(n22353), .dinb(n22344), .dout(n22354));
  jxor g22171(.dina(n22354), .dinb(n22330), .dout(n22355));
  jxor g22172(.dina(n22355), .dinb(n22327), .dout(n22356));
  jxor g22173(.dina(n22356), .dinb(n22318), .dout(n22357));
  jnot g22174(.din(n22357), .dout(n22358));
  jor  g22175(.dina(n19940), .dinb(n4747), .dout(n22359));
  jor  g22176(.dina(n19547), .dinb(n4959), .dout(n22360));
  jor  g22177(.dina(n19550), .dinb(n4919), .dout(n22361));
  jor  g22178(.dina(n19553), .dinb(n4746), .dout(n22362));
  jand g22179(.dina(n22362), .dinb(n22361), .dout(n22363));
  jand g22180(.dina(n22363), .dinb(n22360), .dout(n22364));
  jand g22181(.dina(n22364), .dinb(n22359), .dout(n22365));
  jxor g22182(.dina(n22365), .dinb(\a[26] ), .dout(n22366));
  jxor g22183(.dina(n22366), .dinb(n22358), .dout(n22367));
  jxor g22184(.dina(n22367), .dinb(n22315), .dout(n22368));
  jxor g22185(.dina(n22368), .dinb(n22310), .dout(n22369));
  jxor g22186(.dina(n22369), .dinb(n22301), .dout(n22370));
  jnot g22187(.din(n22370), .dout(n22371));
  jand g22188(.dina(n20413), .dinb(n5693), .dout(n22372));
  jand g22189(.dina(n19535), .dinb(n6209), .dout(n22373));
  jand g22190(.dina(n19537), .dinb(n6131), .dout(n22374));
  jand g22191(.dina(n19539), .dinb(n5691), .dout(n22375));
  jor  g22192(.dina(n22375), .dinb(n22374), .dout(n22376));
  jor  g22193(.dina(n22376), .dinb(n22373), .dout(n22377));
  jor  g22194(.dina(n22377), .dinb(n22372), .dout(n22378));
  jxor g22195(.dina(n22378), .dinb(n4247), .dout(n22379));
  jxor g22196(.dina(n22379), .dinb(n22371), .dout(n22380));
  jxor g22197(.dina(n22380), .dinb(n22298), .dout(n22381));
  jxor g22198(.dina(n22381), .dinb(n22293), .dout(n22382));
  jxor g22199(.dina(n22382), .dinb(n22284), .dout(n22383));
  jnot g22200(.din(n22383), .dout(n22384));
  jand g22201(.dina(n19770), .dinb(n6936), .dout(n22385));
  jand g22202(.dina(n19523), .dinb(n7741), .dout(n22386));
  jand g22203(.dina(n19525), .dinb(n7613), .dout(n22387));
  jand g22204(.dina(n19527), .dinb(n6934), .dout(n22388));
  jor  g22205(.dina(n22388), .dinb(n22387), .dout(n22389));
  jor  g22206(.dina(n22389), .dinb(n22386), .dout(n22390));
  jor  g22207(.dina(n22390), .dinb(n22385), .dout(n22391));
  jxor g22208(.dina(n22391), .dinb(n5292), .dout(n22392));
  jxor g22209(.dina(n22392), .dinb(n22384), .dout(n22393));
  jxor g22210(.dina(n22393), .dinb(n22281), .dout(n22394));
  jxor g22211(.dina(n22394), .dinb(n22276), .dout(n22395));
  jxor g22212(.dina(n22395), .dinb(n22267), .dout(n22396));
  jnot g22213(.din(n22396), .dout(n22397));
  jand g22214(.dina(n21762), .dinb(n8771), .dout(n22398));
  jand g22215(.dina(n19511), .dinb(n9491), .dout(n22399));
  jand g22216(.dina(n19513), .dinb(n9126), .dout(n22400));
  jand g22217(.dina(n19515), .dinb(n8769), .dout(n22401));
  jor  g22218(.dina(n22401), .dinb(n22400), .dout(n22402));
  jor  g22219(.dina(n22402), .dinb(n22399), .dout(n22403));
  jor  g22220(.dina(n22403), .dinb(n22398), .dout(n22404));
  jxor g22221(.dina(n22404), .dinb(n6039), .dout(n22405));
  jxor g22222(.dina(n22405), .dinb(n22397), .dout(n22406));
  jxor g22223(.dina(n22406), .dinb(n22264), .dout(n22407));
  jxor g22224(.dina(n22407), .dinb(n22259), .dout(n22408));
  jxor g22225(.dina(n22408), .dinb(n22174), .dout(n22409));
  jnot g22226(.din(n22409), .dout(n22410));
  jand g22227(.dina(n22193), .dinb(n22189), .dout(n22411));
  jand g22228(.dina(n22241), .dinb(n22194), .dout(n22412));
  jor  g22229(.dina(n22412), .dinb(n22411), .dout(n22413));
  jor  g22230(.dina(n4918), .dinb(n4933), .dout(n22416));
  jand g22231(.dina(n12815), .dinb(n4745), .dout(n22418));
  jor  g22232(.dina(n22418), .dinb(n22416), .dout(n22419));
  jor  g22233(.dina(n22419), .dinb(n75), .dout(n22420));
  jxor g22234(.dina(n22420), .dinb(n68), .dout(n22421));
  jnot g22235(.din(n22421), .dout(n22422));
  jor  g22236(.dina(n22219), .dinb(n19723), .dout(n22423));
  jand g22237(.dina(n22220), .dinb(n22204), .dout(n22424));
  jnot g22238(.din(n22424), .dout(n22425));
  jand g22239(.dina(n22425), .dinb(n22423), .dout(n22426));
  jand g22240(.dina(n689), .dinb(n190), .dout(n22427));
  jand g22241(.dina(n553), .dinb(n435), .dout(n22428));
  jand g22242(.dina(n22428), .dinb(n22427), .dout(n22429));
  jand g22243(.dina(n22429), .dinb(n2580), .dout(n22430));
  jand g22244(.dina(n7447), .dinb(n4288), .dout(n22431));
  jand g22245(.dina(n22431), .dinb(n22430), .dout(n22432));
  jand g22246(.dina(n1768), .dinb(n325), .dout(n22433));
  jand g22247(.dina(n2132), .dinb(n1128), .dout(n22434));
  jand g22248(.dina(n3054), .dinb(n2315), .dout(n22435));
  jand g22249(.dina(n22435), .dinb(n22434), .dout(n22436));
  jand g22250(.dina(n22436), .dinb(n22433), .dout(n22437));
  jand g22251(.dina(n22437), .dinb(n22432), .dout(n22438));
  jand g22252(.dina(n22438), .dinb(n3842), .dout(n22439));
  jand g22253(.dina(n22439), .dinb(n12304), .dout(n22440));
  jand g22254(.dina(n22440), .dinb(n840), .dout(n22441));
  jnot g22255(.din(n22441), .dout(n22442));
  jxor g22256(.dina(n22442), .dinb(n22426), .dout(n22443));
  jand g22257(.dina(n12768), .dinb(n732), .dout(n22444));
  jand g22258(.dina(n12766), .dinb(n3855), .dout(n22445));
  jand g22259(.dina(n11941), .dinb(n3851), .dout(n22446));
  jand g22260(.dina(n12177), .dinb(n3858), .dout(n22447));
  jor  g22261(.dina(n22447), .dinb(n22446), .dout(n22448));
  jor  g22262(.dina(n22448), .dinb(n22445), .dout(n22449));
  jor  g22263(.dina(n22449), .dinb(n22444), .dout(n22450));
  jxor g22264(.dina(n22450), .dinb(n22443), .dout(n22451));
  jor  g22265(.dina(n22221), .dinb(n22200), .dout(n22452));
  jand g22266(.dina(n22221), .dinb(n22200), .dout(n22453));
  jor  g22267(.dina(n22229), .dinb(n22453), .dout(n22454));
  jand g22268(.dina(n22454), .dinb(n22452), .dout(n22455));
  jxor g22269(.dina(n22455), .dinb(n22451), .dout(n22456));
  jnot g22270(.din(n22456), .dout(n22457));
  jand g22271(.dina(n12797), .dinb(n4449), .dout(n22458));
  jand g22272(.dina(n12795), .dinb(n4453), .dout(n22459));
  jand g22273(.dina(n12782), .dinb(n4457), .dout(n22460));
  jand g22274(.dina(n12783), .dinb(n4461), .dout(n22461));
  jor  g22275(.dina(n22461), .dinb(n22460), .dout(n22462));
  jor  g22276(.dina(n22462), .dinb(n22459), .dout(n22463));
  jor  g22277(.dina(n22463), .dinb(n22458), .dout(n22464));
  jxor g22278(.dina(n22464), .dinb(n88), .dout(n22465));
  jxor g22279(.dina(n22465), .dinb(n22457), .dout(n22466));
  jnot g22280(.din(n22197), .dout(n22467));
  jnot g22281(.din(n22230), .dout(n22468));
  jand g22282(.dina(n22468), .dinb(n22467), .dout(n22469));
  jnot g22283(.din(n22469), .dout(n22470));
  jand g22284(.dina(n22230), .dinb(n22197), .dout(n22471));
  jor  g22285(.dina(n22240), .dinb(n22471), .dout(n22472));
  jand g22286(.dina(n22472), .dinb(n22470), .dout(n22473));
  jxor g22287(.dina(n22473), .dinb(n22466), .dout(n22474));
  jxor g22288(.dina(n22474), .dinb(n22422), .dout(n22475));
  jand g22289(.dina(n22475), .dinb(n22413), .dout(n22476));
  jand g22290(.dina(n22246), .dinb(n22242), .dout(n22477));
  jand g22291(.dina(n22247), .dinb(n22180), .dout(n22478));
  jor  g22292(.dina(n22478), .dinb(n22477), .dout(n22479));
  jxor g22293(.dina(n22475), .dinb(n22413), .dout(n22480));
  jand g22294(.dina(n22480), .dinb(n22479), .dout(n22481));
  jor  g22295(.dina(n22481), .dinb(n22476), .dout(n22482));
  jnot g22296(.din(n22426), .dout(n22483));
  jand g22297(.dina(n22441), .dinb(n22483), .dout(n22484));
  jand g22298(.dina(n22450), .dinb(n22443), .dout(n22485));
  jor  g22299(.dina(n22485), .dinb(n22484), .dout(n22486));
  jand g22300(.dina(n1153), .dinb(n696), .dout(n22487));
  jand g22301(.dina(n22487), .dinb(n6385), .dout(n22488));
  jand g22302(.dina(n4336), .dinb(n596), .dout(n22489));
  jand g22303(.dina(n22489), .dinb(n22488), .dout(n22490));
  jand g22304(.dina(n1946), .dinb(n1460), .dout(n22491));
  jand g22305(.dina(n22491), .dinb(n22490), .dout(n22492));
  jand g22306(.dina(n22492), .dinb(n2559), .dout(n22493));
  jand g22307(.dina(n22493), .dinb(n4435), .dout(n22494));
  jand g22308(.dina(n22494), .dinb(n12304), .dout(n22495));
  jand g22309(.dina(n22495), .dinb(n3818), .dout(n22496));
  jand g22310(.dina(n22496), .dinb(n3799), .dout(n22497));
  jxor g22311(.dina(n22497), .dinb(n22442), .dout(n22498));
  jand g22312(.dina(n12841), .dinb(n732), .dout(n22499));
  jand g22313(.dina(n12783), .dinb(n3855), .dout(n22500));
  jand g22314(.dina(n12766), .dinb(n3858), .dout(n22501));
  jand g22315(.dina(n12177), .dinb(n3851), .dout(n22502));
  jor  g22316(.dina(n22502), .dinb(n22501), .dout(n22503));
  jor  g22317(.dina(n22503), .dinb(n22500), .dout(n22504));
  jor  g22318(.dina(n22504), .dinb(n22499), .dout(n22505));
  jxor g22319(.dina(n22505), .dinb(n22498), .dout(n22506));
  jxor g22320(.dina(n22506), .dinb(n22486), .dout(n22507));
  jnot g22321(.din(n22507), .dout(n22508));
  jand g22322(.dina(n22455), .dinb(n22451), .dout(n22509));
  jnot g22323(.din(n22509), .dout(n22510));
  jor  g22324(.dina(n22465), .dinb(n22457), .dout(n22511));
  jand g22325(.dina(n22511), .dinb(n22510), .dout(n22512));
  jxor g22326(.dina(n22512), .dinb(n22508), .dout(n22513));
  jand g22327(.dina(n12919), .dinb(n4449), .dout(n22521));
  jand g22328(.dina(n12815), .dinb(n4453), .dout(n22522));
  jand g22329(.dina(n12795), .dinb(n4457), .dout(n22523));
  jand g22330(.dina(n12782), .dinb(n4461), .dout(n22524));
  jor  g22331(.dina(n22524), .dinb(n22523), .dout(n22525));
  jor  g22332(.dina(n22525), .dinb(n22522), .dout(n22526));
  jor  g22333(.dina(n22526), .dinb(n22521), .dout(n22527));
  jxor g22334(.dina(n22527), .dinb(n88), .dout(n22528));
  jxor g22335(.dina(n22528), .dinb(n22577), .dout(n22529));
  jxor g22336(.dina(n22529), .dinb(n22513), .dout(n22530));
  jnot g22337(.din(n22466), .dout(n22531));
  jnot g22338(.din(n22473), .dout(n22532));
  jand g22339(.dina(n22532), .dinb(n22531), .dout(n22533));
  jnot g22340(.din(n22533), .dout(n22534));
  jand g22341(.dina(n22473), .dinb(n22466), .dout(n22535));
  jor  g22342(.dina(n22535), .dinb(n22422), .dout(n22536));
  jand g22343(.dina(n22536), .dinb(n22534), .dout(n22537));
  jxor g22344(.dina(n22537), .dinb(n22530), .dout(n22538));
  jxor g22345(.dina(n22538), .dinb(n22482), .dout(n22539));
  jxor g22346(.dina(n22480), .dinb(n22479), .dout(n22540));
  jand g22347(.dina(n22540), .dinb(n22539), .dout(n22541));
  jand g22348(.dina(n22540), .dinb(n22248), .dout(n22542));
  jand g22349(.dina(n22248), .dinb(n19758), .dout(n22543));
  jand g22350(.dina(n22249), .dinb(n22177), .dout(n22544));
  jor  g22351(.dina(n22544), .dinb(n22543), .dout(n22545));
  jxor g22352(.dina(n22540), .dinb(n22248), .dout(n22546));
  jand g22353(.dina(n22546), .dinb(n22545), .dout(n22547));
  jor  g22354(.dina(n22547), .dinb(n22542), .dout(n22548));
  jxor g22355(.dina(n22540), .dinb(n22539), .dout(n22549));
  jand g22356(.dina(n22549), .dinb(n22548), .dout(n22550));
  jor  g22357(.dina(n22550), .dinb(n22541), .dout(n22551));
  jand g22358(.dina(n22537), .dinb(n22530), .dout(n22552));
  jand g22359(.dina(n22538), .dinb(n22482), .dout(n22553));
  jor  g22360(.dina(n22553), .dinb(n22552), .dout(n22554));
  jand g22361(.dina(n22506), .dinb(n22486), .dout(n22555));
  jnot g22362(.din(n22555), .dout(n22556));
  jor  g22363(.dina(n22512), .dinb(n22508), .dout(n22557));
  jand g22364(.dina(n22557), .dinb(n22556), .dout(n22558));
  jnot g22365(.din(n22558), .dout(n22559));
  jand g22366(.dina(n13022), .dinb(n4449), .dout(n22560));
  jand g22367(.dina(n12815), .dinb(n4457), .dout(n22562));
  jand g22368(.dina(n12795), .dinb(n4461), .dout(n22563));
  jor  g22369(.dina(n22563), .dinb(n22562), .dout(n22564));
  jor  g22370(.dina(n22564), .dinb(n4453), .dout(n22565));
  jor  g22371(.dina(n22565), .dinb(n22560), .dout(n22566));
  jxor g22372(.dina(n22566), .dinb(n88), .dout(n22567));
  jnot g22373(.din(n22567), .dout(n22568));
  jor  g22374(.dina(n22497), .dinb(n22442), .dout(n22569));
  jand g22375(.dina(n22505), .dinb(n22498), .dout(n22570));
  jnot g22376(.din(n22570), .dout(n22571));
  jand g22377(.dina(n22571), .dinb(n22569), .dout(n22572));
  jnot g22378(.din(n22572), .dout(n22573));
  jnot g22379(.din(n4744), .dout(n22574));
  jor  g22380(.dina(n22574), .dinb(n71), .dout(n22575));
  jxor g22381(.dina(n22575), .dinb(n68), .dout(n22577));
  jand g22382(.dina(n4606), .dinb(n4582), .dout(n22578));
  jand g22383(.dina(n330), .dinb(n154), .dout(n22579));
  jand g22384(.dina(n22579), .dinb(n869), .dout(n22580));
  jand g22385(.dina(n22580), .dinb(n4427), .dout(n22581));
  jand g22386(.dina(n22581), .dinb(n4406), .dout(n22582));
  jand g22387(.dina(n22582), .dinb(n22578), .dout(n22583));
  jxor g22388(.dina(n22583), .dinb(n22441), .dout(n22584));
  jxor g22389(.dina(n22584), .dinb(n22577), .dout(n22585));
  jxor g22390(.dina(n22585), .dinb(n22573), .dout(n22586));
  jand g22391(.dina(n12938), .dinb(n732), .dout(n22587));
  jand g22392(.dina(n12782), .dinb(n3855), .dout(n22588));
  jand g22393(.dina(n12783), .dinb(n3858), .dout(n22589));
  jand g22394(.dina(n12766), .dinb(n3851), .dout(n22590));
  jor  g22395(.dina(n22590), .dinb(n22589), .dout(n22591));
  jor  g22396(.dina(n22591), .dinb(n22588), .dout(n22592));
  jor  g22397(.dina(n22592), .dinb(n22587), .dout(n22593));
  jxor g22398(.dina(n22593), .dinb(n22586), .dout(n22594));
  jxor g22399(.dina(n22594), .dinb(n22568), .dout(n22595));
  jxor g22400(.dina(n22595), .dinb(n22559), .dout(n22596));
  jnot g22401(.din(n22596), .dout(n22597));
  jor  g22402(.dina(n22528), .dinb(n22577), .dout(n22598));
  jand g22403(.dina(n22529), .dinb(n22513), .dout(n22599));
  jnot g22404(.din(n22599), .dout(n22600));
  jand g22405(.dina(n22600), .dinb(n22598), .dout(n22601));
  jxor g22406(.dina(n22601), .dinb(n22597), .dout(n22602));
  jxor g22407(.dina(n22602), .dinb(n22554), .dout(n22603));
  jxor g22408(.dina(n22603), .dinb(n22539), .dout(n22604));
  jxor g22409(.dina(n22604), .dinb(n22551), .dout(n22605));
  jand g22410(.dina(n22605), .dinb(n10846), .dout(n22606));
  jand g22411(.dina(n22603), .dinb(n11372), .dout(n22607));
  jand g22412(.dina(n22539), .dinb(n11359), .dout(n22608));
  jand g22413(.dina(n22540), .dinb(n10844), .dout(n22609));
  jor  g22414(.dina(n22609), .dinb(n22608), .dout(n22610));
  jor  g22415(.dina(n22610), .dinb(n22607), .dout(n22611));
  jor  g22416(.dina(n22611), .dinb(n22606), .dout(n22612));
  jxor g22417(.dina(n22612), .dinb(n6600), .dout(n22613));
  jor  g22418(.dina(n22613), .dinb(n22410), .dout(n22614));
  jnot g22419(.din(n22614), .dout(n22615));
  jxor g22420(.dina(n22613), .dinb(n22410), .dout(n22616));
  jxor g22421(.dina(n22549), .dinb(n22548), .dout(n22617));
  jand g22422(.dina(n22617), .dinb(n10846), .dout(n22618));
  jand g22423(.dina(n22539), .dinb(n11372), .dout(n22619));
  jand g22424(.dina(n22540), .dinb(n11359), .dout(n22620));
  jand g22425(.dina(n22248), .dinb(n10844), .dout(n22621));
  jor  g22426(.dina(n22621), .dinb(n22620), .dout(n22622));
  jor  g22427(.dina(n22622), .dinb(n22619), .dout(n22623));
  jor  g22428(.dina(n22623), .dinb(n22618), .dout(n22624));
  jxor g22429(.dina(n22624), .dinb(n6600), .dout(n22625));
  jnot g22430(.din(n22625), .dout(n22626));
  jxor g22431(.dina(n22546), .dinb(n22545), .dout(n22627));
  jand g22432(.dina(n22627), .dinb(n10846), .dout(n22628));
  jand g22433(.dina(n22540), .dinb(n11372), .dout(n22629));
  jand g22434(.dina(n22248), .dinb(n11359), .dout(n22630));
  jand g22435(.dina(n19758), .dinb(n10844), .dout(n22631));
  jor  g22436(.dina(n22631), .dinb(n22630), .dout(n22632));
  jor  g22437(.dina(n22632), .dinb(n22629), .dout(n22633));
  jor  g22438(.dina(n22633), .dinb(n22628), .dout(n22634));
  jxor g22439(.dina(n22634), .dinb(n6600), .dout(n22635));
  jnot g22440(.din(n22635), .dout(n22636));
  jand g22441(.dina(n22250), .dinb(n10846), .dout(n22637));
  jand g22442(.dina(n22248), .dinb(n11372), .dout(n22638));
  jand g22443(.dina(n19758), .dinb(n11359), .dout(n22639));
  jand g22444(.dina(n19510), .dinb(n10844), .dout(n22640));
  jor  g22445(.dina(n22640), .dinb(n22639), .dout(n22641));
  jor  g22446(.dina(n22641), .dinb(n22638), .dout(n22642));
  jor  g22447(.dina(n22642), .dinb(n22637), .dout(n22643));
  jxor g22448(.dina(n22643), .dinb(n6600), .dout(n22644));
  jnot g22449(.din(n22644), .dout(n22645));
  jxor g22450(.dina(n22161), .dinb(n22160), .dout(n22646));
  jxor g22451(.dina(n22156), .dinb(n22155), .dout(n22647));
  jand g22452(.dina(n21762), .dinb(n10846), .dout(n22648));
  jand g22453(.dina(n19511), .dinb(n11372), .dout(n22649));
  jand g22454(.dina(n19513), .dinb(n11359), .dout(n22650));
  jand g22455(.dina(n19515), .dinb(n10844), .dout(n22651));
  jor  g22456(.dina(n22651), .dinb(n22650), .dout(n22652));
  jor  g22457(.dina(n22652), .dinb(n22649), .dout(n22653));
  jor  g22458(.dina(n22653), .dinb(n22648), .dout(n22654));
  jxor g22459(.dina(n22654), .dinb(n6600), .dout(n22655));
  jnot g22460(.din(n22655), .dout(n22656));
  jand g22461(.dina(n21738), .dinb(n10846), .dout(n22657));
  jand g22462(.dina(n19513), .dinb(n11372), .dout(n22658));
  jand g22463(.dina(n19515), .dinb(n11359), .dout(n22659));
  jand g22464(.dina(n19517), .dinb(n10844), .dout(n22660));
  jor  g22465(.dina(n22660), .dinb(n22659), .dout(n22661));
  jor  g22466(.dina(n22661), .dinb(n22658), .dout(n22662));
  jor  g22467(.dina(n22662), .dinb(n22657), .dout(n22663));
  jxor g22468(.dina(n22663), .dinb(n6600), .dout(n22664));
  jnot g22469(.din(n22664), .dout(n22665));
  jand g22470(.dina(n21218), .dinb(n10846), .dout(n22666));
  jand g22471(.dina(n19515), .dinb(n11372), .dout(n22667));
  jand g22472(.dina(n19517), .dinb(n11359), .dout(n22668));
  jand g22473(.dina(n19519), .dinb(n10844), .dout(n22669));
  jor  g22474(.dina(n22669), .dinb(n22668), .dout(n22670));
  jor  g22475(.dina(n22670), .dinb(n22667), .dout(n22671));
  jor  g22476(.dina(n22671), .dinb(n22666), .dout(n22672));
  jxor g22477(.dina(n22672), .dinb(n6600), .dout(n22673));
  jnot g22478(.din(n22673), .dout(n22674));
  jxor g22479(.dina(n22142), .dinb(n22141), .dout(n22675));
  jxor g22480(.dina(n22137), .dinb(n22136), .dout(n22676));
  jxor g22481(.dina(n22132), .dinb(n22131), .dout(n22677));
  jand g22482(.dina(n19770), .dinb(n10846), .dout(n22678));
  jand g22483(.dina(n19523), .dinb(n11372), .dout(n22679));
  jand g22484(.dina(n19525), .dinb(n11359), .dout(n22680));
  jand g22485(.dina(n19527), .dinb(n10844), .dout(n22681));
  jor  g22486(.dina(n22681), .dinb(n22680), .dout(n22682));
  jor  g22487(.dina(n22682), .dinb(n22679), .dout(n22683));
  jor  g22488(.dina(n22683), .dinb(n22678), .dout(n22684));
  jxor g22489(.dina(n22684), .dinb(n6600), .dout(n22685));
  jnot g22490(.din(n22685), .dout(n22686));
  jand g22491(.dina(n20781), .dinb(n10846), .dout(n22687));
  jand g22492(.dina(n19525), .dinb(n11372), .dout(n22688));
  jand g22493(.dina(n19527), .dinb(n11359), .dout(n22689));
  jand g22494(.dina(n19529), .dinb(n10844), .dout(n22690));
  jor  g22495(.dina(n22690), .dinb(n22689), .dout(n22691));
  jor  g22496(.dina(n22691), .dinb(n22688), .dout(n22692));
  jor  g22497(.dina(n22692), .dinb(n22687), .dout(n22693));
  jxor g22498(.dina(n22693), .dinb(n6600), .dout(n22694));
  jnot g22499(.din(n22694), .dout(n22695));
  jand g22500(.dina(n20793), .dinb(n10846), .dout(n22696));
  jand g22501(.dina(n19527), .dinb(n11372), .dout(n22697));
  jand g22502(.dina(n19529), .dinb(n11359), .dout(n22698));
  jand g22503(.dina(n19531), .dinb(n10844), .dout(n22699));
  jor  g22504(.dina(n22699), .dinb(n22698), .dout(n22700));
  jor  g22505(.dina(n22700), .dinb(n22697), .dout(n22701));
  jor  g22506(.dina(n22701), .dinb(n22696), .dout(n22702));
  jxor g22507(.dina(n22702), .dinb(n6600), .dout(n22703));
  jnot g22508(.din(n22703), .dout(n22704));
  jxor g22509(.dina(n22118), .dinb(n22117), .dout(n22705));
  jxor g22510(.dina(n22113), .dinb(n22112), .dout(n22706));
  jxor g22511(.dina(n22108), .dinb(n22107), .dout(n22707));
  jand g22512(.dina(n20413), .dinb(n10846), .dout(n22708));
  jand g22513(.dina(n19535), .dinb(n11372), .dout(n22709));
  jand g22514(.dina(n19537), .dinb(n11359), .dout(n22710));
  jand g22515(.dina(n19539), .dinb(n10844), .dout(n22711));
  jor  g22516(.dina(n22711), .dinb(n22710), .dout(n22712));
  jor  g22517(.dina(n22712), .dinb(n22709), .dout(n22713));
  jor  g22518(.dina(n22713), .dinb(n22708), .dout(n22714));
  jxor g22519(.dina(n22714), .dinb(n6600), .dout(n22715));
  jnot g22520(.din(n22715), .dout(n22716));
  jand g22521(.dina(n20387), .dinb(n10846), .dout(n22717));
  jand g22522(.dina(n19537), .dinb(n11372), .dout(n22718));
  jand g22523(.dina(n19539), .dinb(n11359), .dout(n22719));
  jand g22524(.dina(n19541), .dinb(n10844), .dout(n22720));
  jor  g22525(.dina(n22720), .dinb(n22719), .dout(n22721));
  jor  g22526(.dina(n22721), .dinb(n22718), .dout(n22722));
  jor  g22527(.dina(n22722), .dinb(n22717), .dout(n22723));
  jxor g22528(.dina(n22723), .dinb(n6600), .dout(n22724));
  jnot g22529(.din(n22724), .dout(n22725));
  jand g22530(.dina(n20131), .dinb(n10846), .dout(n22726));
  jand g22531(.dina(n19539), .dinb(n11372), .dout(n22727));
  jand g22532(.dina(n19541), .dinb(n11359), .dout(n22728));
  jand g22533(.dina(n19543), .dinb(n10844), .dout(n22729));
  jor  g22534(.dina(n22729), .dinb(n22728), .dout(n22730));
  jor  g22535(.dina(n22730), .dinb(n22727), .dout(n22731));
  jor  g22536(.dina(n22731), .dinb(n22726), .dout(n22732));
  jxor g22537(.dina(n22732), .dinb(n6600), .dout(n22733));
  jnot g22538(.din(n22733), .dout(n22734));
  jxor g22539(.dina(n22094), .dinb(n22093), .dout(n22735));
  jxor g22540(.dina(n22089), .dinb(n22088), .dout(n22736));
  jxor g22541(.dina(n22084), .dinb(n22083), .dout(n22737));
  jor  g22542(.dina(n19940), .dinb(n10847), .dout(n22738));
  jor  g22543(.dina(n19547), .dinb(n11458), .dout(n22739));
  jor  g22544(.dina(n19550), .dinb(n11360), .dout(n22740));
  jor  g22545(.dina(n19553), .dinb(n10845), .dout(n22741));
  jand g22546(.dina(n22741), .dinb(n22740), .dout(n22742));
  jand g22547(.dina(n22742), .dinb(n22739), .dout(n22743));
  jand g22548(.dina(n22743), .dinb(n22738), .dout(n22744));
  jxor g22549(.dina(n22744), .dinb(n6600), .dout(n22745));
  jor  g22550(.dina(n19952), .dinb(n10847), .dout(n22746));
  jor  g22551(.dina(n19550), .dinb(n11458), .dout(n22747));
  jor  g22552(.dina(n19553), .dinb(n11360), .dout(n22748));
  jor  g22553(.dina(n19558), .dinb(n10845), .dout(n22749));
  jand g22554(.dina(n22749), .dinb(n22748), .dout(n22750));
  jand g22555(.dina(n22750), .dinb(n22747), .dout(n22751));
  jand g22556(.dina(n22751), .dinb(n22746), .dout(n22752));
  jxor g22557(.dina(n22752), .dinb(n6600), .dout(n22753));
  jor  g22558(.dina(n19964), .dinb(n10847), .dout(n22754));
  jor  g22559(.dina(n19553), .dinb(n11458), .dout(n22755));
  jor  g22560(.dina(n19558), .dinb(n11360), .dout(n22756));
  jor  g22561(.dina(n19562), .dinb(n10845), .dout(n22757));
  jand g22562(.dina(n22757), .dinb(n22756), .dout(n22758));
  jand g22563(.dina(n22758), .dinb(n22755), .dout(n22759));
  jand g22564(.dina(n22759), .dinb(n22754), .dout(n22760));
  jxor g22565(.dina(n22760), .dinb(n6600), .dout(n22761));
  jxor g22566(.dina(n22072), .dinb(n22071), .dout(n22762));
  jor  g22567(.dina(n19790), .dinb(n10847), .dout(n22763));
  jor  g22568(.dina(n19562), .dinb(n11458), .dout(n22764));
  jor  g22569(.dina(n19564), .dinb(n11360), .dout(n22765));
  jor  g22570(.dina(n19566), .dinb(n10845), .dout(n22766));
  jand g22571(.dina(n22766), .dinb(n22765), .dout(n22767));
  jand g22572(.dina(n22767), .dinb(n22764), .dout(n22768));
  jand g22573(.dina(n22768), .dinb(n22763), .dout(n22769));
  jxor g22574(.dina(n22769), .dinb(n6600), .dout(n22770));
  jor  g22575(.dina(n22049), .dinb(n64), .dout(n22771));
  jxor g22576(.dina(n22771), .dinb(n22057), .dout(n22772));
  jor  g22577(.dina(n19852), .dinb(n10847), .dout(n22773));
  jor  g22578(.dina(n19566), .dinb(n11458), .dout(n22774));
  jor  g22579(.dina(n19568), .dinb(n11360), .dout(n22775));
  jor  g22580(.dina(n19570), .dinb(n10845), .dout(n22776));
  jand g22581(.dina(n22776), .dinb(n22775), .dout(n22777));
  jand g22582(.dina(n22777), .dinb(n22774), .dout(n22778));
  jand g22583(.dina(n22778), .dinb(n22773), .dout(n22779));
  jxor g22584(.dina(n22779), .dinb(n6600), .dout(n22780));
  jor  g22585(.dina(n19801), .dinb(n10847), .dout(n22781));
  jor  g22586(.dina(n19568), .dinb(n11458), .dout(n22782));
  jand g22587(.dina(n19572), .dinb(n11359), .dout(n22783));
  jand g22588(.dina(n19574), .dinb(n10844), .dout(n22784));
  jor  g22589(.dina(n22784), .dinb(n22783), .dout(n22785));
  jnot g22590(.din(n22785), .dout(n22786));
  jand g22591(.dina(n22786), .dinb(n22782), .dout(n22787));
  jand g22592(.dina(n22787), .dinb(n22781), .dout(n22788));
  jand g22593(.dina(n22788), .dinb(n22046), .dout(n22789));
  jand g22594(.dina(n19570), .dinb(n11371), .dout(n22790));
  jor  g22595(.dina(n22790), .dinb(n10840), .dout(n22791));
  jor  g22596(.dina(n19575), .dinb(n10842), .dout(n22792));
  jand g22597(.dina(n22792), .dinb(n22791), .dout(n22793));
  jand g22598(.dina(n19812), .dinb(n10846), .dout(n22794));
  jand g22599(.dina(n22794), .dinb(n19825), .dout(n22795));
  jor  g22600(.dina(n22795), .dinb(n22793), .dout(n22796));
  jand g22601(.dina(n22796), .dinb(n19577), .dout(n22797));
  jor  g22602(.dina(n22797), .dinb(n6600), .dout(n22798));
  jor  g22603(.dina(n22798), .dinb(n22789), .dout(n22799));
  jand g22604(.dina(n21685), .dinb(n10846), .dout(n22800));
  jand g22605(.dina(n21687), .dinb(n11372), .dout(n22801));
  jor  g22606(.dina(n22785), .dinb(n22801), .dout(n22802));
  jor  g22607(.dina(n22802), .dinb(n22800), .dout(n22803));
  jor  g22608(.dina(n22803), .dinb(\a[2] ), .dout(n22804));
  jor  g22609(.dina(n22788), .dinb(n22046), .dout(n22805));
  jand g22610(.dina(n22805), .dinb(n22804), .dout(n22806));
  jand g22611(.dina(n22806), .dinb(n22799), .dout(n22807));
  jand g22612(.dina(n22807), .dinb(n22780), .dout(n22808));
  jor  g22613(.dina(n22807), .dinb(n22780), .dout(n22809));
  jand g22614(.dina(n22046), .dinb(\a[5] ), .dout(n22810));
  jxor g22615(.dina(n22810), .dinb(n22044), .dout(n22811));
  jand g22616(.dina(n22811), .dinb(n22809), .dout(n22812));
  jor  g22617(.dina(n22812), .dinb(n22808), .dout(n22813));
  jand g22618(.dina(n22813), .dinb(n22772), .dout(n22814));
  jor  g22619(.dina(n22813), .dinb(n22772), .dout(n22815));
  jor  g22620(.dina(n19839), .dinb(n10847), .dout(n22816));
  jor  g22621(.dina(n19564), .dinb(n11458), .dout(n22817));
  jor  g22622(.dina(n19566), .dinb(n11360), .dout(n22818));
  jor  g22623(.dina(n19568), .dinb(n10845), .dout(n22819));
  jand g22624(.dina(n22819), .dinb(n22818), .dout(n22820));
  jand g22625(.dina(n22820), .dinb(n22817), .dout(n22821));
  jand g22626(.dina(n22821), .dinb(n22816), .dout(n22822));
  jxor g22627(.dina(n22822), .dinb(n6600), .dout(n22823));
  jand g22628(.dina(n22823), .dinb(n22815), .dout(n22824));
  jor  g22629(.dina(n22824), .dinb(n22814), .dout(n22825));
  jand g22630(.dina(n22825), .dinb(n22770), .dout(n22826));
  jor  g22631(.dina(n22825), .dinb(n22770), .dout(n22827));
  jxor g22632(.dina(n22069), .dinb(n22068), .dout(n22828));
  jand g22633(.dina(n22828), .dinb(n22827), .dout(n22829));
  jor  g22634(.dina(n22829), .dinb(n22826), .dout(n22830));
  jand g22635(.dina(n22830), .dinb(n22762), .dout(n22831));
  jor  g22636(.dina(n22830), .dinb(n22762), .dout(n22832));
  jor  g22637(.dina(n19906), .dinb(n10847), .dout(n22833));
  jor  g22638(.dina(n19558), .dinb(n11458), .dout(n22834));
  jor  g22639(.dina(n19562), .dinb(n11360), .dout(n22835));
  jor  g22640(.dina(n19564), .dinb(n10845), .dout(n22836));
  jand g22641(.dina(n22836), .dinb(n22835), .dout(n22837));
  jand g22642(.dina(n22837), .dinb(n22834), .dout(n22838));
  jand g22643(.dina(n22838), .dinb(n22833), .dout(n22839));
  jxor g22644(.dina(n22839), .dinb(n6600), .dout(n22840));
  jand g22645(.dina(n22840), .dinb(n22832), .dout(n22841));
  jor  g22646(.dina(n22841), .dinb(n22831), .dout(n22842));
  jand g22647(.dina(n22842), .dinb(n22761), .dout(n22843));
  jor  g22648(.dina(n22842), .dinb(n22761), .dout(n22844));
  jxor g22649(.dina(n22075), .dinb(n22074), .dout(n22845));
  jand g22650(.dina(n22845), .dinb(n22844), .dout(n22846));
  jor  g22651(.dina(n22846), .dinb(n22843), .dout(n22847));
  jand g22652(.dina(n22847), .dinb(n22753), .dout(n22848));
  jor  g22653(.dina(n22847), .dinb(n22753), .dout(n22849));
  jxor g22654(.dina(n22078), .dinb(n22077), .dout(n22850));
  jand g22655(.dina(n22850), .dinb(n22849), .dout(n22851));
  jor  g22656(.dina(n22851), .dinb(n22848), .dout(n22852));
  jand g22657(.dina(n22852), .dinb(n22745), .dout(n22853));
  jor  g22658(.dina(n22852), .dinb(n22745), .dout(n22854));
  jxor g22659(.dina(n22081), .dinb(n22080), .dout(n22855));
  jand g22660(.dina(n22855), .dinb(n22854), .dout(n22856));
  jor  g22661(.dina(n22856), .dinb(n22853), .dout(n22857));
  jand g22662(.dina(n22857), .dinb(n22737), .dout(n22858));
  jor  g22663(.dina(n22857), .dinb(n22737), .dout(n22859));
  jand g22664(.dina(n20079), .dinb(n10846), .dout(n22860));
  jand g22665(.dina(n19545), .dinb(n11372), .dout(n22861));
  jand g22666(.dina(n19548), .dinb(n11359), .dout(n22862));
  jand g22667(.dina(n19551), .dinb(n10844), .dout(n22863));
  jor  g22668(.dina(n22863), .dinb(n22862), .dout(n22864));
  jor  g22669(.dina(n22864), .dinb(n22861), .dout(n22865));
  jor  g22670(.dina(n22865), .dinb(n22860), .dout(n22866));
  jxor g22671(.dina(n22866), .dinb(\a[2] ), .dout(n22867));
  jand g22672(.dina(n22867), .dinb(n22859), .dout(n22868));
  jor  g22673(.dina(n22868), .dinb(n22858), .dout(n22869));
  jand g22674(.dina(n22869), .dinb(n22736), .dout(n22870));
  jor  g22675(.dina(n22869), .dinb(n22736), .dout(n22871));
  jand g22676(.dina(n20153), .dinb(n10846), .dout(n22872));
  jand g22677(.dina(n19543), .dinb(n11372), .dout(n22873));
  jand g22678(.dina(n19545), .dinb(n11359), .dout(n22874));
  jand g22679(.dina(n19548), .dinb(n10844), .dout(n22875));
  jor  g22680(.dina(n22875), .dinb(n22874), .dout(n22876));
  jor  g22681(.dina(n22876), .dinb(n22873), .dout(n22877));
  jor  g22682(.dina(n22877), .dinb(n22872), .dout(n22878));
  jxor g22683(.dina(n22878), .dinb(\a[2] ), .dout(n22879));
  jand g22684(.dina(n22879), .dinb(n22871), .dout(n22880));
  jor  g22685(.dina(n22880), .dinb(n22870), .dout(n22881));
  jand g22686(.dina(n22881), .dinb(n22735), .dout(n22882));
  jor  g22687(.dina(n22881), .dinb(n22735), .dout(n22883));
  jand g22688(.dina(n20141), .dinb(n10846), .dout(n22884));
  jand g22689(.dina(n19541), .dinb(n11372), .dout(n22885));
  jand g22690(.dina(n19543), .dinb(n11359), .dout(n22886));
  jand g22691(.dina(n19545), .dinb(n10844), .dout(n22887));
  jor  g22692(.dina(n22887), .dinb(n22886), .dout(n22888));
  jor  g22693(.dina(n22888), .dinb(n22885), .dout(n22889));
  jor  g22694(.dina(n22889), .dinb(n22884), .dout(n22890));
  jxor g22695(.dina(n22890), .dinb(\a[2] ), .dout(n22891));
  jand g22696(.dina(n22891), .dinb(n22883), .dout(n22892));
  jor  g22697(.dina(n22892), .dinb(n22882), .dout(n22893));
  jand g22698(.dina(n22893), .dinb(n22734), .dout(n22894));
  jor  g22699(.dina(n22893), .dinb(n22734), .dout(n22895));
  jxor g22700(.dina(n22099), .dinb(n22098), .dout(n22896));
  jand g22701(.dina(n22896), .dinb(n22895), .dout(n22897));
  jor  g22702(.dina(n22897), .dinb(n22894), .dout(n22898));
  jand g22703(.dina(n22898), .dinb(n22725), .dout(n22899));
  jor  g22704(.dina(n22898), .dinb(n22725), .dout(n22900));
  jxor g22705(.dina(n22102), .dinb(n22101), .dout(n22901));
  jand g22706(.dina(n22901), .dinb(n22900), .dout(n22902));
  jor  g22707(.dina(n22902), .dinb(n22899), .dout(n22903));
  jand g22708(.dina(n22903), .dinb(n22716), .dout(n22904));
  jor  g22709(.dina(n22903), .dinb(n22716), .dout(n22905));
  jxor g22710(.dina(n22105), .dinb(n22104), .dout(n22906));
  jand g22711(.dina(n22906), .dinb(n22905), .dout(n22907));
  jor  g22712(.dina(n22907), .dinb(n22904), .dout(n22908));
  jand g22713(.dina(n22908), .dinb(n22707), .dout(n22909));
  jor  g22714(.dina(n22908), .dinb(n22707), .dout(n22910));
  jand g22715(.dina(n20399), .dinb(n10846), .dout(n22911));
  jand g22716(.dina(n19533), .dinb(n11372), .dout(n22912));
  jand g22717(.dina(n19535), .dinb(n11359), .dout(n22913));
  jand g22718(.dina(n19537), .dinb(n10844), .dout(n22914));
  jor  g22719(.dina(n22914), .dinb(n22913), .dout(n22915));
  jor  g22720(.dina(n22915), .dinb(n22912), .dout(n22916));
  jor  g22721(.dina(n22916), .dinb(n22911), .dout(n22917));
  jxor g22722(.dina(n22917), .dinb(\a[2] ), .dout(n22918));
  jand g22723(.dina(n22918), .dinb(n22910), .dout(n22919));
  jor  g22724(.dina(n22919), .dinb(n22909), .dout(n22920));
  jand g22725(.dina(n22920), .dinb(n22706), .dout(n22921));
  jor  g22726(.dina(n22920), .dinb(n22706), .dout(n22922));
  jand g22727(.dina(n19780), .dinb(n10846), .dout(n22923));
  jand g22728(.dina(n19531), .dinb(n11372), .dout(n22924));
  jand g22729(.dina(n19533), .dinb(n11359), .dout(n22925));
  jand g22730(.dina(n19535), .dinb(n10844), .dout(n22926));
  jor  g22731(.dina(n22926), .dinb(n22925), .dout(n22927));
  jor  g22732(.dina(n22927), .dinb(n22924), .dout(n22928));
  jor  g22733(.dina(n22928), .dinb(n22923), .dout(n22929));
  jxor g22734(.dina(n22929), .dinb(\a[2] ), .dout(n22930));
  jand g22735(.dina(n22930), .dinb(n22922), .dout(n22931));
  jor  g22736(.dina(n22931), .dinb(n22921), .dout(n22932));
  jand g22737(.dina(n22932), .dinb(n22705), .dout(n22933));
  jor  g22738(.dina(n22932), .dinb(n22705), .dout(n22934));
  jand g22739(.dina(n20767), .dinb(n10846), .dout(n22935));
  jand g22740(.dina(n19529), .dinb(n11372), .dout(n22936));
  jand g22741(.dina(n19531), .dinb(n11359), .dout(n22937));
  jand g22742(.dina(n19533), .dinb(n10844), .dout(n22938));
  jor  g22743(.dina(n22938), .dinb(n22937), .dout(n22939));
  jor  g22744(.dina(n22939), .dinb(n22936), .dout(n22940));
  jor  g22745(.dina(n22940), .dinb(n22935), .dout(n22941));
  jxor g22746(.dina(n22941), .dinb(\a[2] ), .dout(n22942));
  jand g22747(.dina(n22942), .dinb(n22934), .dout(n22943));
  jor  g22748(.dina(n22943), .dinb(n22933), .dout(n22944));
  jand g22749(.dina(n22944), .dinb(n22704), .dout(n22945));
  jor  g22750(.dina(n22944), .dinb(n22704), .dout(n22946));
  jxor g22751(.dina(n22123), .dinb(n22122), .dout(n22947));
  jand g22752(.dina(n22947), .dinb(n22946), .dout(n22948));
  jor  g22753(.dina(n22948), .dinb(n22945), .dout(n22949));
  jand g22754(.dina(n22949), .dinb(n22695), .dout(n22950));
  jor  g22755(.dina(n22949), .dinb(n22695), .dout(n22951));
  jxor g22756(.dina(n22126), .dinb(n22125), .dout(n22952));
  jand g22757(.dina(n22952), .dinb(n22951), .dout(n22953));
  jor  g22758(.dina(n22953), .dinb(n22950), .dout(n22954));
  jand g22759(.dina(n22954), .dinb(n22686), .dout(n22955));
  jor  g22760(.dina(n22954), .dinb(n22686), .dout(n22956));
  jxor g22761(.dina(n22129), .dinb(n22128), .dout(n22957));
  jand g22762(.dina(n22957), .dinb(n22956), .dout(n22958));
  jor  g22763(.dina(n22958), .dinb(n22955), .dout(n22959));
  jand g22764(.dina(n22959), .dinb(n22677), .dout(n22960));
  jor  g22765(.dina(n22959), .dinb(n22677), .dout(n22961));
  jand g22766(.dina(n21086), .dinb(n10846), .dout(n22962));
  jand g22767(.dina(n19521), .dinb(n11372), .dout(n22963));
  jand g22768(.dina(n19523), .dinb(n11359), .dout(n22964));
  jand g22769(.dina(n19525), .dinb(n10844), .dout(n22965));
  jor  g22770(.dina(n22965), .dinb(n22964), .dout(n22966));
  jor  g22771(.dina(n22966), .dinb(n22963), .dout(n22967));
  jor  g22772(.dina(n22967), .dinb(n22962), .dout(n22968));
  jxor g22773(.dina(n22968), .dinb(\a[2] ), .dout(n22969));
  jand g22774(.dina(n22969), .dinb(n22961), .dout(n22970));
  jor  g22775(.dina(n22970), .dinb(n22960), .dout(n22971));
  jand g22776(.dina(n22971), .dinb(n22676), .dout(n22972));
  jor  g22777(.dina(n22971), .dinb(n22676), .dout(n22973));
  jand g22778(.dina(n21240), .dinb(n10846), .dout(n22974));
  jand g22779(.dina(n19519), .dinb(n11372), .dout(n22975));
  jand g22780(.dina(n19521), .dinb(n11359), .dout(n22976));
  jand g22781(.dina(n19523), .dinb(n10844), .dout(n22977));
  jor  g22782(.dina(n22977), .dinb(n22976), .dout(n22978));
  jor  g22783(.dina(n22978), .dinb(n22975), .dout(n22979));
  jor  g22784(.dina(n22979), .dinb(n22974), .dout(n22980));
  jxor g22785(.dina(n22980), .dinb(\a[2] ), .dout(n22981));
  jand g22786(.dina(n22981), .dinb(n22973), .dout(n22982));
  jor  g22787(.dina(n22982), .dinb(n22972), .dout(n22983));
  jand g22788(.dina(n22983), .dinb(n22675), .dout(n22984));
  jor  g22789(.dina(n22983), .dinb(n22675), .dout(n22985));
  jand g22790(.dina(n21230), .dinb(n10846), .dout(n22986));
  jand g22791(.dina(n19517), .dinb(n11372), .dout(n22987));
  jand g22792(.dina(n19519), .dinb(n11359), .dout(n22988));
  jand g22793(.dina(n19521), .dinb(n10844), .dout(n22989));
  jor  g22794(.dina(n22989), .dinb(n22988), .dout(n22990));
  jor  g22795(.dina(n22990), .dinb(n22987), .dout(n22991));
  jor  g22796(.dina(n22991), .dinb(n22986), .dout(n22992));
  jxor g22797(.dina(n22992), .dinb(\a[2] ), .dout(n22993));
  jand g22798(.dina(n22993), .dinb(n22985), .dout(n22994));
  jor  g22799(.dina(n22994), .dinb(n22984), .dout(n22995));
  jand g22800(.dina(n22995), .dinb(n22674), .dout(n22996));
  jor  g22801(.dina(n22995), .dinb(n22674), .dout(n22997));
  jxor g22802(.dina(n22147), .dinb(n22146), .dout(n22998));
  jand g22803(.dina(n22998), .dinb(n22997), .dout(n22999));
  jor  g22804(.dina(n22999), .dinb(n22996), .dout(n23000));
  jand g22805(.dina(n23000), .dinb(n22665), .dout(n23001));
  jor  g22806(.dina(n23000), .dinb(n22665), .dout(n23002));
  jxor g22807(.dina(n22150), .dinb(n22149), .dout(n23003));
  jand g22808(.dina(n23003), .dinb(n23002), .dout(n23004));
  jor  g22809(.dina(n23004), .dinb(n23001), .dout(n23005));
  jand g22810(.dina(n23005), .dinb(n22656), .dout(n23006));
  jor  g22811(.dina(n23005), .dinb(n22656), .dout(n23007));
  jxor g22812(.dina(n22153), .dinb(n22152), .dout(n23008));
  jand g22813(.dina(n23008), .dinb(n23007), .dout(n23009));
  jor  g22814(.dina(n23009), .dinb(n23006), .dout(n23010));
  jand g22815(.dina(n23010), .dinb(n22647), .dout(n23011));
  jor  g22816(.dina(n23010), .dinb(n22647), .dout(n23012));
  jand g22817(.dina(n21750), .dinb(n10846), .dout(n23013));
  jand g22818(.dina(n19510), .dinb(n11372), .dout(n23014));
  jand g22819(.dina(n19511), .dinb(n11359), .dout(n23015));
  jand g22820(.dina(n19513), .dinb(n10844), .dout(n23016));
  jor  g22821(.dina(n23016), .dinb(n23015), .dout(n23017));
  jor  g22822(.dina(n23017), .dinb(n23014), .dout(n23018));
  jor  g22823(.dina(n23018), .dinb(n23013), .dout(n23019));
  jxor g22824(.dina(n23019), .dinb(\a[2] ), .dout(n23020));
  jand g22825(.dina(n23020), .dinb(n23012), .dout(n23021));
  jor  g22826(.dina(n23021), .dinb(n23011), .dout(n23022));
  jand g22827(.dina(n23022), .dinb(n22646), .dout(n23023));
  jor  g22828(.dina(n23022), .dinb(n22646), .dout(n23024));
  jand g22829(.dina(n19760), .dinb(n10846), .dout(n23025));
  jand g22830(.dina(n19758), .dinb(n11372), .dout(n23026));
  jand g22831(.dina(n19510), .dinb(n11359), .dout(n23027));
  jand g22832(.dina(n19511), .dinb(n10844), .dout(n23028));
  jor  g22833(.dina(n23028), .dinb(n23027), .dout(n23029));
  jor  g22834(.dina(n23029), .dinb(n23026), .dout(n23030));
  jor  g22835(.dina(n23030), .dinb(n23025), .dout(n23031));
  jxor g22836(.dina(n23031), .dinb(\a[2] ), .dout(n23032));
  jand g22837(.dina(n23032), .dinb(n23024), .dout(n23033));
  jor  g22838(.dina(n23033), .dinb(n23023), .dout(n23034));
  jand g22839(.dina(n23034), .dinb(n22645), .dout(n23035));
  jor  g22840(.dina(n23034), .dinb(n22645), .dout(n23036));
  jxor g22841(.dina(n22166), .dinb(n22165), .dout(n23037));
  jand g22842(.dina(n23037), .dinb(n23036), .dout(n23038));
  jor  g22843(.dina(n23038), .dinb(n23035), .dout(n23039));
  jand g22844(.dina(n23039), .dinb(n22636), .dout(n23040));
  jor  g22845(.dina(n23039), .dinb(n22636), .dout(n23041));
  jxor g22846(.dina(n22169), .dinb(n22168), .dout(n23042));
  jand g22847(.dina(n23042), .dinb(n23041), .dout(n23043));
  jor  g22848(.dina(n23043), .dinb(n23040), .dout(n23044));
  jand g22849(.dina(n23044), .dinb(n22626), .dout(n23045));
  jor  g22850(.dina(n23044), .dinb(n22626), .dout(n23046));
  jxor g22851(.dina(n22172), .dinb(n22171), .dout(n23047));
  jand g22852(.dina(n23047), .dinb(n23046), .dout(n23048));
  jor  g22853(.dina(n23048), .dinb(n23045), .dout(n23049));
  jand g22854(.dina(n23049), .dinb(n22616), .dout(n23050));
  jor  g22855(.dina(n23050), .dinb(n22615), .dout(n23051));
  jand g22856(.dina(n22407), .dinb(n22259), .dout(n23052));
  jand g22857(.dina(n22408), .dinb(n22174), .dout(n23053));
  jor  g22858(.dina(n23053), .dinb(n23052), .dout(n23054));
  jand g22859(.dina(n22627), .dinb(n67), .dout(n23055));
  jand g22860(.dina(n22540), .dinb(n10827), .dout(n23056));
  jand g22861(.dina(n22248), .dinb(n10350), .dout(n23057));
  jand g22862(.dina(n19758), .dinb(n9917), .dout(n23058));
  jor  g22863(.dina(n23058), .dinb(n23057), .dout(n23059));
  jor  g22864(.dina(n23059), .dinb(n23056), .dout(n23060));
  jor  g22865(.dina(n23060), .dinb(n23055), .dout(n23061));
  jxor g22866(.dina(n23061), .dinb(n64), .dout(n23062));
  jnot g22867(.din(n23062), .dout(n23063));
  jor  g22868(.dina(n22405), .dinb(n22397), .dout(n23064));
  jand g22869(.dina(n22406), .dinb(n22264), .dout(n23065));
  jnot g22870(.din(n23065), .dout(n23066));
  jand g22871(.dina(n23066), .dinb(n23064), .dout(n23067));
  jnot g22872(.din(n23067), .dout(n23068));
  jand g22873(.dina(n22394), .dinb(n22276), .dout(n23069));
  jand g22874(.dina(n22395), .dinb(n22267), .dout(n23070));
  jor  g22875(.dina(n23070), .dinb(n23069), .dout(n23071));
  jand g22876(.dina(n21218), .dinb(n7890), .dout(n23072));
  jand g22877(.dina(n19515), .dinb(n8441), .dout(n23073));
  jand g22878(.dina(n19517), .dinb(n8154), .dout(n23074));
  jand g22879(.dina(n19519), .dinb(n7888), .dout(n23075));
  jor  g22880(.dina(n23075), .dinb(n23074), .dout(n23076));
  jor  g22881(.dina(n23076), .dinb(n23073), .dout(n23077));
  jor  g22882(.dina(n23077), .dinb(n23072), .dout(n23078));
  jxor g22883(.dina(n23078), .dinb(n5833), .dout(n23079));
  jnot g22884(.din(n23079), .dout(n23080));
  jor  g22885(.dina(n22392), .dinb(n22384), .dout(n23081));
  jand g22886(.dina(n22393), .dinb(n22281), .dout(n23082));
  jnot g22887(.din(n23082), .dout(n23083));
  jand g22888(.dina(n23083), .dinb(n23081), .dout(n23084));
  jnot g22889(.din(n23084), .dout(n23085));
  jand g22890(.dina(n22381), .dinb(n22293), .dout(n23086));
  jand g22891(.dina(n22382), .dinb(n22284), .dout(n23087));
  jor  g22892(.dina(n23087), .dinb(n23086), .dout(n23088));
  jand g22893(.dina(n20793), .dinb(n6340), .dout(n23089));
  jand g22894(.dina(n19527), .dinb(n6798), .dout(n23090));
  jand g22895(.dina(n19529), .dinb(n6556), .dout(n23091));
  jand g22896(.dina(n19531), .dinb(n6338), .dout(n23092));
  jor  g22897(.dina(n23092), .dinb(n23091), .dout(n23093));
  jor  g22898(.dina(n23093), .dinb(n23090), .dout(n23094));
  jor  g22899(.dina(n23094), .dinb(n23089), .dout(n23095));
  jxor g22900(.dina(n23095), .dinb(n5064), .dout(n23096));
  jnot g22901(.din(n23096), .dout(n23097));
  jor  g22902(.dina(n22379), .dinb(n22371), .dout(n23098));
  jand g22903(.dina(n22380), .dinb(n22298), .dout(n23099));
  jnot g22904(.din(n23099), .dout(n23100));
  jand g22905(.dina(n23100), .dinb(n23098), .dout(n23101));
  jnot g22906(.din(n23101), .dout(n23102));
  jand g22907(.dina(n22368), .dinb(n22310), .dout(n23103));
  jand g22908(.dina(n22369), .dinb(n22301), .dout(n23104));
  jor  g22909(.dina(n23104), .dinb(n23103), .dout(n23105));
  jand g22910(.dina(n20131), .dinb(n5365), .dout(n23106));
  jand g22911(.dina(n19539), .dinb(n5500), .dout(n23107));
  jand g22912(.dina(n19541), .dinb(n5424), .dout(n23108));
  jand g22913(.dina(n19543), .dinb(n5363), .dout(n23109));
  jor  g22914(.dina(n23109), .dinb(n23108), .dout(n23110));
  jor  g22915(.dina(n23110), .dinb(n23107), .dout(n23111));
  jor  g22916(.dina(n23111), .dinb(n23106), .dout(n23112));
  jxor g22917(.dina(n23112), .dinb(n72), .dout(n23113));
  jnot g22918(.din(n23113), .dout(n23114));
  jor  g22919(.dina(n22366), .dinb(n22358), .dout(n23115));
  jand g22920(.dina(n22367), .dinb(n22315), .dout(n23116));
  jnot g22921(.din(n23116), .dout(n23117));
  jand g22922(.dina(n23117), .dinb(n23115), .dout(n23118));
  jnot g22923(.din(n23118), .dout(n23119));
  jand g22924(.dina(n22355), .dinb(n22327), .dout(n23120));
  jand g22925(.dina(n22356), .dinb(n22318), .dout(n23121));
  jor  g22926(.dina(n23121), .dinb(n23120), .dout(n23122));
  jor  g22927(.dina(n19964), .dinb(n4724), .dout(n23123));
  jor  g22928(.dina(n19553), .dinb(n4905), .dout(n23124));
  jor  g22929(.dina(n19558), .dinb(n4735), .dout(n23125));
  jor  g22930(.dina(n19562), .dinb(n4733), .dout(n23126));
  jand g22931(.dina(n23126), .dinb(n23125), .dout(n23127));
  jand g22932(.dina(n23127), .dinb(n23124), .dout(n23128));
  jand g22933(.dina(n23128), .dinb(n23123), .dout(n23129));
  jxor g22934(.dina(n23129), .dinb(\a[29] ), .dout(n23130));
  jnot g22935(.din(n23130), .dout(n23131));
  jor  g22936(.dina(n22353), .dinb(n22344), .dout(n23132));
  jand g22937(.dina(n22354), .dinb(n22330), .dout(n23133));
  jnot g22938(.din(n23133), .dout(n23134));
  jand g22939(.dina(n23134), .dinb(n23132), .dout(n23135));
  jnot g22940(.din(n23135), .dout(n23136));
  jand g22941(.dina(n1840), .dinb(n393), .dout(n23137));
  jand g22942(.dina(n3989), .dinb(n1306), .dout(n23138));
  jand g22943(.dina(n23138), .dinb(n23137), .dout(n23139));
  jand g22944(.dina(n23139), .dinb(n5596), .dout(n23140));
  jand g22945(.dina(n23140), .dinb(n12488), .dout(n23141));
  jand g22946(.dina(n12722), .dinb(n2507), .dout(n23142));
  jand g22947(.dina(n983), .dinb(n506), .dout(n23143));
  jand g22948(.dina(n23143), .dinb(n23142), .dout(n23144));
  jand g22949(.dina(n23144), .dinb(n2702), .dout(n23145));
  jand g22950(.dina(n23145), .dinb(n4239), .dout(n23146));
  jand g22951(.dina(n23146), .dinb(n23141), .dout(n23147));
  jand g22952(.dina(n23147), .dinb(n5181), .dout(n23148));
  jand g22953(.dina(n23148), .dinb(n12220), .dout(n23149));
  jor  g22954(.dina(n19839), .dinb(n6463), .dout(n23150));
  jnot g22955(.din(n19564), .dout(n23151));
  jand g22956(.dina(n23151), .dinb(n3855), .dout(n23152));
  jand g22957(.dina(n21687), .dinb(n3851), .dout(n23153));
  jand g22958(.dina(n22346), .dinb(n3858), .dout(n23154));
  jor  g22959(.dina(n23154), .dinb(n23153), .dout(n23155));
  jor  g22960(.dina(n23155), .dinb(n23152), .dout(n23156));
  jnot g22961(.din(n23156), .dout(n23157));
  jand g22962(.dina(n23157), .dinb(n23150), .dout(n23158));
  jxor g22963(.dina(n23158), .dinb(n23149), .dout(n23159));
  jxor g22964(.dina(n23159), .dinb(n23136), .dout(n23160));
  jxor g22965(.dina(n23160), .dinb(n23131), .dout(n23161));
  jxor g22966(.dina(n23161), .dinb(n23122), .dout(n23162));
  jnot g22967(.din(n23162), .dout(n23163));
  jand g22968(.dina(n20079), .dinb(n75), .dout(n23164));
  jand g22969(.dina(n19545), .dinb(n4933), .dout(n23165));
  jand g22970(.dina(n19548), .dinb(n4918), .dout(n23166));
  jand g22971(.dina(n19551), .dinb(n4745), .dout(n23167));
  jor  g22972(.dina(n23167), .dinb(n23166), .dout(n23168));
  jor  g22973(.dina(n23168), .dinb(n23165), .dout(n23169));
  jor  g22974(.dina(n23169), .dinb(n23164), .dout(n23170));
  jxor g22975(.dina(n23170), .dinb(n68), .dout(n23171));
  jxor g22976(.dina(n23171), .dinb(n23163), .dout(n23172));
  jxor g22977(.dina(n23172), .dinb(n23119), .dout(n23173));
  jxor g22978(.dina(n23173), .dinb(n23114), .dout(n23174));
  jxor g22979(.dina(n23174), .dinb(n23105), .dout(n23175));
  jnot g22980(.din(n23175), .dout(n23176));
  jand g22981(.dina(n20399), .dinb(n5693), .dout(n23177));
  jand g22982(.dina(n19533), .dinb(n6209), .dout(n23178));
  jand g22983(.dina(n19535), .dinb(n6131), .dout(n23179));
  jand g22984(.dina(n19537), .dinb(n5691), .dout(n23180));
  jor  g22985(.dina(n23180), .dinb(n23179), .dout(n23181));
  jor  g22986(.dina(n23181), .dinb(n23178), .dout(n23182));
  jor  g22987(.dina(n23182), .dinb(n23177), .dout(n23183));
  jxor g22988(.dina(n23183), .dinb(n4247), .dout(n23184));
  jxor g22989(.dina(n23184), .dinb(n23176), .dout(n23185));
  jxor g22990(.dina(n23185), .dinb(n23102), .dout(n23186));
  jxor g22991(.dina(n23186), .dinb(n23097), .dout(n23187));
  jxor g22992(.dina(n23187), .dinb(n23088), .dout(n23188));
  jnot g22993(.din(n23188), .dout(n23189));
  jand g22994(.dina(n21086), .dinb(n6936), .dout(n23190));
  jand g22995(.dina(n19521), .dinb(n7741), .dout(n23191));
  jand g22996(.dina(n19523), .dinb(n7613), .dout(n23192));
  jand g22997(.dina(n19525), .dinb(n6934), .dout(n23193));
  jor  g22998(.dina(n23193), .dinb(n23192), .dout(n23194));
  jor  g22999(.dina(n23194), .dinb(n23191), .dout(n23195));
  jor  g23000(.dina(n23195), .dinb(n23190), .dout(n23196));
  jxor g23001(.dina(n23196), .dinb(n5292), .dout(n23197));
  jxor g23002(.dina(n23197), .dinb(n23189), .dout(n23198));
  jxor g23003(.dina(n23198), .dinb(n23085), .dout(n23199));
  jxor g23004(.dina(n23199), .dinb(n23080), .dout(n23200));
  jxor g23005(.dina(n23200), .dinb(n23071), .dout(n23201));
  jnot g23006(.din(n23201), .dout(n23202));
  jand g23007(.dina(n21750), .dinb(n8771), .dout(n23203));
  jand g23008(.dina(n19510), .dinb(n9491), .dout(n23204));
  jand g23009(.dina(n19511), .dinb(n9126), .dout(n23205));
  jand g23010(.dina(n19513), .dinb(n8769), .dout(n23206));
  jor  g23011(.dina(n23206), .dinb(n23205), .dout(n23207));
  jor  g23012(.dina(n23207), .dinb(n23204), .dout(n23208));
  jor  g23013(.dina(n23208), .dinb(n23203), .dout(n23209));
  jxor g23014(.dina(n23209), .dinb(n6039), .dout(n23210));
  jxor g23015(.dina(n23210), .dinb(n23202), .dout(n23211));
  jxor g23016(.dina(n23211), .dinb(n23068), .dout(n23212));
  jxor g23017(.dina(n23212), .dinb(n23063), .dout(n23213));
  jxor g23018(.dina(n23213), .dinb(n23054), .dout(n23214));
  jnot g23019(.din(n23214), .dout(n23215));
  jand g23020(.dina(n22603), .dinb(n22539), .dout(n23216));
  jand g23021(.dina(n22604), .dinb(n22551), .dout(n23217));
  jor  g23022(.dina(n23217), .dinb(n23216), .dout(n23218));
  jor  g23023(.dina(n22601), .dinb(n22597), .dout(n23219));
  jand g23024(.dina(n22602), .dinb(n22554), .dout(n23220));
  jnot g23025(.din(n23220), .dout(n23221));
  jand g23026(.dina(n23221), .dinb(n23219), .dout(n23222));
  jnot g23027(.din(n23222), .dout(n23223));
  jand g23028(.dina(n22594), .dinb(n22568), .dout(n23224));
  jand g23029(.dina(n22595), .dinb(n22559), .dout(n23225));
  jor  g23030(.dina(n23225), .dinb(n23224), .dout(n23226));
  jor  g23031(.dina(n22583), .dinb(n22441), .dout(n23227));
  jand g23032(.dina(n22584), .dinb(n22577), .dout(n23228));
  jnot g23033(.din(n23228), .dout(n23229));
  jand g23034(.dina(n23229), .dinb(n23227), .dout(n23230));
  jand g23035(.dina(n4627), .dinb(n330), .dout(n23231));
  jand g23036(.dina(n23231), .dinb(n4376), .dout(n23232));
  jand g23037(.dina(n23232), .dinb(n22578), .dout(n23233));
  jnot g23038(.din(n23233), .dout(n23234));
  jxor g23039(.dina(n23234), .dinb(n23230), .dout(n23235));
  jand g23040(.dina(n12797), .dinb(n732), .dout(n23236));
  jand g23041(.dina(n12795), .dinb(n3855), .dout(n23237));
  jand g23042(.dina(n12782), .dinb(n3858), .dout(n23238));
  jor  g23043(.dina(n22590), .dinb(n23238), .dout(n23240));
  jor  g23044(.dina(n23240), .dinb(n23237), .dout(n23241));
  jor  g23045(.dina(n23241), .dinb(n23236), .dout(n23242));
  jxor g23046(.dina(n23242), .dinb(n23235), .dout(n23243));
  jor  g23047(.dina(n22585), .dinb(n22573), .dout(n23244));
  jand g23048(.dina(n22585), .dinb(n22573), .dout(n23245));
  jor  g23049(.dina(n22593), .dinb(n23245), .dout(n23246));
  jand g23050(.dina(n23246), .dinb(n23244), .dout(n23247));
  jxor g23051(.dina(n23247), .dinb(n23243), .dout(n23248));
  jnot g23052(.din(n23248), .dout(n23249));
  jxor g23053(.dina(n23693), .dinb(n23249), .dout(n23258));
  jxor g23054(.dina(n23258), .dinb(n23226), .dout(n23259));
  jxor g23055(.dina(n23259), .dinb(n23223), .dout(n23260));
  jxor g23056(.dina(n23260), .dinb(n22603), .dout(n23261));
  jxor g23057(.dina(n23261), .dinb(n23218), .dout(n23262));
  jand g23058(.dina(n23262), .dinb(n10846), .dout(n23263));
  jand g23059(.dina(n23260), .dinb(n11372), .dout(n23264));
  jand g23060(.dina(n22603), .dinb(n11359), .dout(n23265));
  jand g23061(.dina(n22539), .dinb(n10844), .dout(n23266));
  jor  g23062(.dina(n23266), .dinb(n23265), .dout(n23267));
  jor  g23063(.dina(n23267), .dinb(n23264), .dout(n23268));
  jor  g23064(.dina(n23268), .dinb(n23263), .dout(n23269));
  jxor g23065(.dina(n23269), .dinb(n6600), .dout(n23270));
  jxor g23066(.dina(n23270), .dinb(n23215), .dout(n23271));
  jxor g23067(.dina(n23271), .dinb(n23051), .dout(n23272));
  jxor g23068(.dina(n23049), .dinb(n22616), .dout(n23273));
  jxor g23069(.dina(n23273), .dinb(n23272), .dout(\result[0] ));
  jand g23070(.dina(n23273), .dinb(n23272), .dout(n23275));
  jor  g23071(.dina(n23270), .dinb(n23215), .dout(n23276));
  jnot g23072(.din(n23276), .dout(n23277));
  jand g23073(.dina(n23271), .dinb(n23051), .dout(n23278));
  jor  g23074(.dina(n23278), .dinb(n23277), .dout(n23279));
  jand g23075(.dina(n23212), .dinb(n23063), .dout(n23280));
  jand g23076(.dina(n23213), .dinb(n23054), .dout(n23281));
  jor  g23077(.dina(n23281), .dinb(n23280), .dout(n23282));
  jand g23078(.dina(n22617), .dinb(n67), .dout(n23283));
  jand g23079(.dina(n22539), .dinb(n10827), .dout(n23284));
  jand g23080(.dina(n22540), .dinb(n10350), .dout(n23285));
  jand g23081(.dina(n22248), .dinb(n9917), .dout(n23286));
  jor  g23082(.dina(n23286), .dinb(n23285), .dout(n23287));
  jor  g23083(.dina(n23287), .dinb(n23284), .dout(n23288));
  jor  g23084(.dina(n23288), .dinb(n23283), .dout(n23289));
  jxor g23085(.dina(n23289), .dinb(n64), .dout(n23290));
  jnot g23086(.din(n23290), .dout(n23291));
  jor  g23087(.dina(n23210), .dinb(n23202), .dout(n23292));
  jand g23088(.dina(n23211), .dinb(n23068), .dout(n23293));
  jnot g23089(.din(n23293), .dout(n23294));
  jand g23090(.dina(n23294), .dinb(n23292), .dout(n23295));
  jnot g23091(.din(n23295), .dout(n23296));
  jand g23092(.dina(n23199), .dinb(n23080), .dout(n23297));
  jand g23093(.dina(n23200), .dinb(n23071), .dout(n23298));
  jor  g23094(.dina(n23298), .dinb(n23297), .dout(n23299));
  jand g23095(.dina(n21738), .dinb(n7890), .dout(n23300));
  jand g23096(.dina(n19513), .dinb(n8441), .dout(n23301));
  jand g23097(.dina(n19515), .dinb(n8154), .dout(n23302));
  jand g23098(.dina(n19517), .dinb(n7888), .dout(n23303));
  jor  g23099(.dina(n23303), .dinb(n23302), .dout(n23304));
  jor  g23100(.dina(n23304), .dinb(n23301), .dout(n23305));
  jor  g23101(.dina(n23305), .dinb(n23300), .dout(n23306));
  jxor g23102(.dina(n23306), .dinb(n5833), .dout(n23307));
  jnot g23103(.din(n23307), .dout(n23308));
  jor  g23104(.dina(n23197), .dinb(n23189), .dout(n23309));
  jand g23105(.dina(n23198), .dinb(n23085), .dout(n23310));
  jnot g23106(.din(n23310), .dout(n23311));
  jand g23107(.dina(n23311), .dinb(n23309), .dout(n23312));
  jnot g23108(.din(n23312), .dout(n23313));
  jand g23109(.dina(n23186), .dinb(n23097), .dout(n23314));
  jand g23110(.dina(n23187), .dinb(n23088), .dout(n23315));
  jor  g23111(.dina(n23315), .dinb(n23314), .dout(n23316));
  jand g23112(.dina(n20781), .dinb(n6340), .dout(n23317));
  jand g23113(.dina(n19525), .dinb(n6798), .dout(n23318));
  jand g23114(.dina(n19527), .dinb(n6556), .dout(n23319));
  jand g23115(.dina(n19529), .dinb(n6338), .dout(n23320));
  jor  g23116(.dina(n23320), .dinb(n23319), .dout(n23321));
  jor  g23117(.dina(n23321), .dinb(n23318), .dout(n23322));
  jor  g23118(.dina(n23322), .dinb(n23317), .dout(n23323));
  jxor g23119(.dina(n23323), .dinb(n5064), .dout(n23324));
  jnot g23120(.din(n23324), .dout(n23325));
  jor  g23121(.dina(n23184), .dinb(n23176), .dout(n23326));
  jand g23122(.dina(n23185), .dinb(n23102), .dout(n23327));
  jnot g23123(.din(n23327), .dout(n23328));
  jand g23124(.dina(n23328), .dinb(n23326), .dout(n23329));
  jnot g23125(.din(n23329), .dout(n23330));
  jand g23126(.dina(n23173), .dinb(n23114), .dout(n23331));
  jand g23127(.dina(n23174), .dinb(n23105), .dout(n23332));
  jor  g23128(.dina(n23332), .dinb(n23331), .dout(n23333));
  jand g23129(.dina(n20387), .dinb(n5365), .dout(n23334));
  jand g23130(.dina(n19537), .dinb(n5500), .dout(n23335));
  jand g23131(.dina(n19539), .dinb(n5424), .dout(n23336));
  jand g23132(.dina(n19541), .dinb(n5363), .dout(n23337));
  jor  g23133(.dina(n23337), .dinb(n23336), .dout(n23338));
  jor  g23134(.dina(n23338), .dinb(n23335), .dout(n23339));
  jor  g23135(.dina(n23339), .dinb(n23334), .dout(n23340));
  jxor g23136(.dina(n23340), .dinb(n72), .dout(n23341));
  jnot g23137(.din(n23341), .dout(n23342));
  jor  g23138(.dina(n23171), .dinb(n23163), .dout(n23343));
  jand g23139(.dina(n23172), .dinb(n23119), .dout(n23344));
  jnot g23140(.din(n23344), .dout(n23345));
  jand g23141(.dina(n23345), .dinb(n23343), .dout(n23346));
  jnot g23142(.din(n23346), .dout(n23347));
  jand g23143(.dina(n23160), .dinb(n23131), .dout(n23348));
  jand g23144(.dina(n23161), .dinb(n23122), .dout(n23349));
  jor  g23145(.dina(n23349), .dinb(n23348), .dout(n23350));
  jor  g23146(.dina(n19952), .dinb(n4724), .dout(n23351));
  jor  g23147(.dina(n19550), .dinb(n4905), .dout(n23352));
  jor  g23148(.dina(n19553), .dinb(n4735), .dout(n23353));
  jor  g23149(.dina(n19558), .dinb(n4733), .dout(n23354));
  jand g23150(.dina(n23354), .dinb(n23353), .dout(n23355));
  jand g23151(.dina(n23355), .dinb(n23352), .dout(n23356));
  jand g23152(.dina(n23356), .dinb(n23351), .dout(n23357));
  jxor g23153(.dina(n23357), .dinb(\a[29] ), .dout(n23358));
  jnot g23154(.din(n23358), .dout(n23359));
  jor  g23155(.dina(n23158), .dinb(n23149), .dout(n23360));
  jand g23156(.dina(n23159), .dinb(n23136), .dout(n23361));
  jnot g23157(.din(n23361), .dout(n23362));
  jand g23158(.dina(n23362), .dinb(n23360), .dout(n23363));
  jnot g23159(.din(n23363), .dout(n23364));
  jand g23160(.dina(n2483), .dinb(n263), .dout(n23365));
  jand g23161(.dina(n23365), .dinb(n393), .dout(n23366));
  jand g23162(.dina(n756), .dinb(n367), .dout(n23367));
  jand g23163(.dina(n23367), .dinb(n1023), .dout(n23368));
  jand g23164(.dina(n3445), .dinb(n2416), .dout(n23369));
  jand g23165(.dina(n23369), .dinb(n23368), .dout(n23370));
  jand g23166(.dina(n23370), .dinb(n23366), .dout(n23371));
  jand g23167(.dina(n23371), .dinb(n7088), .dout(n23372));
  jand g23168(.dina(n1153), .dinb(n626), .dout(n23373));
  jand g23169(.dina(n997), .dinb(n424), .dout(n23374));
  jand g23170(.dina(n23374), .dinb(n23373), .dout(n23375));
  jand g23171(.dina(n23375), .dinb(n2849), .dout(n23376));
  jand g23172(.dina(n23376), .dinb(n1122), .dout(n23377));
  jand g23173(.dina(n23377), .dinb(n7341), .dout(n23378));
  jand g23174(.dina(n23378), .dinb(n23372), .dout(n23379));
  jand g23175(.dina(n13226), .dinb(n3245), .dout(n23380));
  jand g23176(.dina(n23380), .dinb(n23379), .dout(n23381));
  jand g23177(.dina(n23381), .dinb(n1292), .dout(n23382));
  jor  g23178(.dina(n19790), .dinb(n6463), .dout(n23383));
  jnot g23179(.din(n19562), .dout(n23384));
  jand g23180(.dina(n23384), .dinb(n3855), .dout(n23385));
  jand g23181(.dina(n22346), .dinb(n3851), .dout(n23386));
  jand g23182(.dina(n23151), .dinb(n3858), .dout(n23387));
  jor  g23183(.dina(n23387), .dinb(n23386), .dout(n23388));
  jor  g23184(.dina(n23388), .dinb(n23385), .dout(n23389));
  jnot g23185(.din(n23389), .dout(n23390));
  jand g23186(.dina(n23390), .dinb(n23383), .dout(n23391));
  jxor g23187(.dina(n23391), .dinb(n23382), .dout(n23392));
  jxor g23188(.dina(n23392), .dinb(n23364), .dout(n23393));
  jxor g23189(.dina(n23393), .dinb(n23359), .dout(n23394));
  jxor g23190(.dina(n23394), .dinb(n23350), .dout(n23395));
  jnot g23191(.din(n23395), .dout(n23396));
  jand g23192(.dina(n20153), .dinb(n75), .dout(n23397));
  jand g23193(.dina(n19543), .dinb(n4933), .dout(n23398));
  jand g23194(.dina(n19545), .dinb(n4918), .dout(n23399));
  jand g23195(.dina(n19548), .dinb(n4745), .dout(n23400));
  jor  g23196(.dina(n23400), .dinb(n23399), .dout(n23401));
  jor  g23197(.dina(n23401), .dinb(n23398), .dout(n23402));
  jor  g23198(.dina(n23402), .dinb(n23397), .dout(n23403));
  jxor g23199(.dina(n23403), .dinb(n68), .dout(n23404));
  jxor g23200(.dina(n23404), .dinb(n23396), .dout(n23405));
  jxor g23201(.dina(n23405), .dinb(n23347), .dout(n23406));
  jxor g23202(.dina(n23406), .dinb(n23342), .dout(n23407));
  jxor g23203(.dina(n23407), .dinb(n23333), .dout(n23408));
  jnot g23204(.din(n23408), .dout(n23409));
  jand g23205(.dina(n19780), .dinb(n5693), .dout(n23410));
  jand g23206(.dina(n19531), .dinb(n6209), .dout(n23411));
  jand g23207(.dina(n19533), .dinb(n6131), .dout(n23412));
  jand g23208(.dina(n19535), .dinb(n5691), .dout(n23413));
  jor  g23209(.dina(n23413), .dinb(n23412), .dout(n23414));
  jor  g23210(.dina(n23414), .dinb(n23411), .dout(n23415));
  jor  g23211(.dina(n23415), .dinb(n23410), .dout(n23416));
  jxor g23212(.dina(n23416), .dinb(n4247), .dout(n23417));
  jxor g23213(.dina(n23417), .dinb(n23409), .dout(n23418));
  jxor g23214(.dina(n23418), .dinb(n23330), .dout(n23419));
  jxor g23215(.dina(n23419), .dinb(n23325), .dout(n23420));
  jxor g23216(.dina(n23420), .dinb(n23316), .dout(n23421));
  jnot g23217(.din(n23421), .dout(n23422));
  jand g23218(.dina(n21240), .dinb(n6936), .dout(n23423));
  jand g23219(.dina(n19519), .dinb(n7741), .dout(n23424));
  jand g23220(.dina(n19521), .dinb(n7613), .dout(n23425));
  jand g23221(.dina(n19523), .dinb(n6934), .dout(n23426));
  jor  g23222(.dina(n23426), .dinb(n23425), .dout(n23427));
  jor  g23223(.dina(n23427), .dinb(n23424), .dout(n23428));
  jor  g23224(.dina(n23428), .dinb(n23423), .dout(n23429));
  jxor g23225(.dina(n23429), .dinb(n5292), .dout(n23430));
  jxor g23226(.dina(n23430), .dinb(n23422), .dout(n23431));
  jxor g23227(.dina(n23431), .dinb(n23313), .dout(n23432));
  jxor g23228(.dina(n23432), .dinb(n23308), .dout(n23433));
  jxor g23229(.dina(n23433), .dinb(n23299), .dout(n23434));
  jnot g23230(.din(n23434), .dout(n23435));
  jand g23231(.dina(n19760), .dinb(n8771), .dout(n23436));
  jand g23232(.dina(n19758), .dinb(n9491), .dout(n23437));
  jand g23233(.dina(n19510), .dinb(n9126), .dout(n23438));
  jand g23234(.dina(n19511), .dinb(n8769), .dout(n23439));
  jor  g23235(.dina(n23439), .dinb(n23438), .dout(n23440));
  jor  g23236(.dina(n23440), .dinb(n23437), .dout(n23441));
  jor  g23237(.dina(n23441), .dinb(n23436), .dout(n23442));
  jxor g23238(.dina(n23442), .dinb(n6039), .dout(n23443));
  jxor g23239(.dina(n23443), .dinb(n23435), .dout(n23444));
  jxor g23240(.dina(n23444), .dinb(n23296), .dout(n23445));
  jxor g23241(.dina(n23445), .dinb(n23291), .dout(n23446));
  jxor g23242(.dina(n23446), .dinb(n23282), .dout(n23447));
  jnot g23243(.din(n23447), .dout(n23448));
  jnot g23244(.din(n22603), .dout(n23449));
  jnot g23245(.din(n23260), .dout(n23450));
  jor  g23246(.dina(n23450), .dinb(n23449), .dout(n23451));
  jnot g23247(.din(n23218), .dout(n23452));
  jnot g23248(.din(n23261), .dout(n23453));
  jor  g23249(.dina(n23453), .dinb(n23452), .dout(n23454));
  jand g23250(.dina(n23454), .dinb(n23451), .dout(n23455));
  jand g23251(.dina(n23258), .dinb(n23226), .dout(n23456));
  jand g23252(.dina(n23259), .dinb(n23223), .dout(n23457));
  jor  g23253(.dina(n23457), .dinb(n23456), .dout(n23458));
  jand g23254(.dina(n23247), .dinb(n23243), .dout(n23459));
  jnot g23255(.din(n23459), .dout(n23460));
  jor  g23256(.dina(n23693), .dinb(n23249), .dout(n23461));
  jand g23257(.dina(n23461), .dinb(n23460), .dout(n23462));
  jnot g23258(.din(n23462), .dout(n23463));
  jand g23259(.dina(n4629), .dinb(n4566), .dout(n23464));
  jnot g23260(.din(n23464), .dout(n23465));
  jxor g23261(.dina(n23465), .dinb(n23233), .dout(n23466));
  jand g23262(.dina(n23234), .dinb(n23230), .dout(n23467));
  jnot g23263(.din(n23467), .dout(n23468));
  jnot g23264(.din(n23230), .dout(n23469));
  jand g23265(.dina(n23233), .dinb(n23469), .dout(n23470));
  jor  g23266(.dina(n23242), .dinb(n23470), .dout(n23471));
  jand g23267(.dina(n23471), .dinb(n23468), .dout(n23472));
  jxor g23268(.dina(n23472), .dinb(n23466), .dout(n23473));
  jnot g23269(.din(n23693), .dout(n23481));
  jand g23270(.dina(n12919), .dinb(n732), .dout(n23482));
  jand g23271(.dina(n12795), .dinb(n3858), .dout(n23484));
  jand g23272(.dina(n12782), .dinb(n3851), .dout(n23485));
  jor  g23273(.dina(n23485), .dinb(n23484), .dout(n23486));
  jor  g23274(.dina(n23486), .dinb(n3855), .dout(n23487));
  jor  g23275(.dina(n23487), .dinb(n23482), .dout(n23488));
  jxor g23276(.dina(n23488), .dinb(n23481), .dout(n23489));
  jxor g23277(.dina(n23489), .dinb(n23473), .dout(n23490));
  jxor g23278(.dina(n23490), .dinb(n23463), .dout(n23491));
  jxor g23279(.dina(n23491), .dinb(n23458), .dout(n23492));
  jxor g23280(.dina(n23492), .dinb(n23260), .dout(n23493));
  jxor g23281(.dina(n23493), .dinb(n23455), .dout(n23494));
  jor  g23282(.dina(n23494), .dinb(n10847), .dout(n23495));
  jnot g23283(.din(n23492), .dout(n23496));
  jor  g23284(.dina(n23496), .dinb(n11458), .dout(n23497));
  jor  g23285(.dina(n23450), .dinb(n11360), .dout(n23498));
  jor  g23286(.dina(n23449), .dinb(n10845), .dout(n23499));
  jand g23287(.dina(n23499), .dinb(n23498), .dout(n23500));
  jand g23288(.dina(n23500), .dinb(n23497), .dout(n23501));
  jand g23289(.dina(n23501), .dinb(n23495), .dout(n23502));
  jxor g23290(.dina(n23502), .dinb(\a[2] ), .dout(n23503));
  jxor g23291(.dina(n23503), .dinb(n23448), .dout(n23504));
  jxor g23292(.dina(n23504), .dinb(n23279), .dout(n23505));
  jxor g23293(.dina(n23505), .dinb(n23275), .dout(\result[1] ));
  jand g23294(.dina(n23505), .dinb(n23275), .dout(n23507));
  jor  g23295(.dina(n23503), .dinb(n23448), .dout(n23508));
  jnot g23296(.din(n23508), .dout(n23509));
  jand g23297(.dina(n23504), .dinb(n23279), .dout(n23510));
  jor  g23298(.dina(n23510), .dinb(n23509), .dout(n23511));
  jand g23299(.dina(n23445), .dinb(n23291), .dout(n23512));
  jand g23300(.dina(n23446), .dinb(n23282), .dout(n23513));
  jor  g23301(.dina(n23513), .dinb(n23512), .dout(n23514));
  jand g23302(.dina(n22605), .dinb(n67), .dout(n23515));
  jand g23303(.dina(n22603), .dinb(n10827), .dout(n23516));
  jand g23304(.dina(n22539), .dinb(n10350), .dout(n23517));
  jand g23305(.dina(n22540), .dinb(n9917), .dout(n23518));
  jor  g23306(.dina(n23518), .dinb(n23517), .dout(n23519));
  jor  g23307(.dina(n23519), .dinb(n23516), .dout(n23520));
  jor  g23308(.dina(n23520), .dinb(n23515), .dout(n23521));
  jxor g23309(.dina(n23521), .dinb(n64), .dout(n23522));
  jnot g23310(.din(n23522), .dout(n23523));
  jor  g23311(.dina(n23443), .dinb(n23435), .dout(n23524));
  jand g23312(.dina(n23444), .dinb(n23296), .dout(n23525));
  jnot g23313(.din(n23525), .dout(n23526));
  jand g23314(.dina(n23526), .dinb(n23524), .dout(n23527));
  jnot g23315(.din(n23527), .dout(n23528));
  jand g23316(.dina(n23432), .dinb(n23308), .dout(n23529));
  jand g23317(.dina(n23433), .dinb(n23299), .dout(n23530));
  jor  g23318(.dina(n23530), .dinb(n23529), .dout(n23531));
  jand g23319(.dina(n21762), .dinb(n7890), .dout(n23532));
  jand g23320(.dina(n19511), .dinb(n8441), .dout(n23533));
  jand g23321(.dina(n19513), .dinb(n8154), .dout(n23534));
  jand g23322(.dina(n19515), .dinb(n7888), .dout(n23535));
  jor  g23323(.dina(n23535), .dinb(n23534), .dout(n23536));
  jor  g23324(.dina(n23536), .dinb(n23533), .dout(n23537));
  jor  g23325(.dina(n23537), .dinb(n23532), .dout(n23538));
  jxor g23326(.dina(n23538), .dinb(n5833), .dout(n23539));
  jnot g23327(.din(n23539), .dout(n23540));
  jor  g23328(.dina(n23430), .dinb(n23422), .dout(n23541));
  jand g23329(.dina(n23431), .dinb(n23313), .dout(n23542));
  jnot g23330(.din(n23542), .dout(n23543));
  jand g23331(.dina(n23543), .dinb(n23541), .dout(n23544));
  jnot g23332(.din(n23544), .dout(n23545));
  jand g23333(.dina(n23419), .dinb(n23325), .dout(n23546));
  jand g23334(.dina(n23420), .dinb(n23316), .dout(n23547));
  jor  g23335(.dina(n23547), .dinb(n23546), .dout(n23548));
  jand g23336(.dina(n19770), .dinb(n6340), .dout(n23549));
  jand g23337(.dina(n19523), .dinb(n6798), .dout(n23550));
  jand g23338(.dina(n19525), .dinb(n6556), .dout(n23551));
  jand g23339(.dina(n19527), .dinb(n6338), .dout(n23552));
  jor  g23340(.dina(n23552), .dinb(n23551), .dout(n23553));
  jor  g23341(.dina(n23553), .dinb(n23550), .dout(n23554));
  jor  g23342(.dina(n23554), .dinb(n23549), .dout(n23555));
  jxor g23343(.dina(n23555), .dinb(n5064), .dout(n23556));
  jnot g23344(.din(n23556), .dout(n23557));
  jor  g23345(.dina(n23417), .dinb(n23409), .dout(n23558));
  jand g23346(.dina(n23418), .dinb(n23330), .dout(n23559));
  jnot g23347(.din(n23559), .dout(n23560));
  jand g23348(.dina(n23560), .dinb(n23558), .dout(n23561));
  jnot g23349(.din(n23561), .dout(n23562));
  jand g23350(.dina(n23406), .dinb(n23342), .dout(n23563));
  jand g23351(.dina(n23407), .dinb(n23333), .dout(n23564));
  jor  g23352(.dina(n23564), .dinb(n23563), .dout(n23565));
  jand g23353(.dina(n20413), .dinb(n5365), .dout(n23566));
  jand g23354(.dina(n19535), .dinb(n5500), .dout(n23567));
  jand g23355(.dina(n19537), .dinb(n5424), .dout(n23568));
  jand g23356(.dina(n19539), .dinb(n5363), .dout(n23569));
  jor  g23357(.dina(n23569), .dinb(n23568), .dout(n23570));
  jor  g23358(.dina(n23570), .dinb(n23567), .dout(n23571));
  jor  g23359(.dina(n23571), .dinb(n23566), .dout(n23572));
  jxor g23360(.dina(n23572), .dinb(n72), .dout(n23573));
  jnot g23361(.din(n23573), .dout(n23574));
  jor  g23362(.dina(n23404), .dinb(n23396), .dout(n23575));
  jand g23363(.dina(n23405), .dinb(n23347), .dout(n23576));
  jnot g23364(.din(n23576), .dout(n23577));
  jand g23365(.dina(n23577), .dinb(n23575), .dout(n23578));
  jnot g23366(.din(n23578), .dout(n23579));
  jand g23367(.dina(n23393), .dinb(n23359), .dout(n23580));
  jand g23368(.dina(n23394), .dinb(n23350), .dout(n23581));
  jor  g23369(.dina(n23581), .dinb(n23580), .dout(n23582));
  jor  g23370(.dina(n19940), .dinb(n4724), .dout(n23583));
  jor  g23371(.dina(n19547), .dinb(n4905), .dout(n23584));
  jor  g23372(.dina(n19550), .dinb(n4735), .dout(n23585));
  jor  g23373(.dina(n19553), .dinb(n4733), .dout(n23586));
  jand g23374(.dina(n23586), .dinb(n23585), .dout(n23587));
  jand g23375(.dina(n23587), .dinb(n23584), .dout(n23588));
  jand g23376(.dina(n23588), .dinb(n23583), .dout(n23589));
  jxor g23377(.dina(n23589), .dinb(\a[29] ), .dout(n23590));
  jnot g23378(.din(n23590), .dout(n23591));
  jor  g23379(.dina(n23391), .dinb(n23382), .dout(n23592));
  jand g23380(.dina(n23392), .dinb(n23364), .dout(n23593));
  jnot g23381(.din(n23593), .dout(n23594));
  jand g23382(.dina(n23594), .dinb(n23592), .dout(n23595));
  jnot g23383(.din(n23595), .dout(n23596));
  jand g23384(.dina(n13884), .dinb(n833), .dout(n23597));
  jand g23385(.dina(n3189), .dinb(n1082), .dout(n23598));
  jand g23386(.dina(n23598), .dinb(n23597), .dout(n23599));
  jand g23387(.dina(n876), .dinb(n824), .dout(n23600));
  jand g23388(.dina(n23600), .dinb(n860), .dout(n23601));
  jand g23389(.dina(n2564), .dinb(n697), .dout(n23602));
  jand g23390(.dina(n23602), .dinb(n23601), .dout(n23603));
  jand g23391(.dina(n23603), .dinb(n23599), .dout(n23604));
  jand g23392(.dina(n7453), .dinb(n2631), .dout(n23605));
  jand g23393(.dina(n23605), .dinb(n23604), .dout(n23606));
  jand g23394(.dina(n13245), .dinb(n1611), .dout(n23607));
  jand g23395(.dina(n23607), .dinb(n12272), .dout(n23608));
  jand g23396(.dina(n23608), .dinb(n4205), .dout(n23609));
  jand g23397(.dina(n23609), .dinb(n23606), .dout(n23610));
  jand g23398(.dina(n23610), .dinb(n2465), .dout(n23611));
  jand g23399(.dina(n23611), .dinb(n4182), .dout(n23612));
  jor  g23400(.dina(n19906), .dinb(n6463), .dout(n23613));
  jand g23401(.dina(n19559), .dinb(n3855), .dout(n23614));
  jand g23402(.dina(n23151), .dinb(n3851), .dout(n23615));
  jand g23403(.dina(n23384), .dinb(n3858), .dout(n23616));
  jor  g23404(.dina(n23616), .dinb(n23615), .dout(n23617));
  jor  g23405(.dina(n23617), .dinb(n23614), .dout(n23618));
  jnot g23406(.din(n23618), .dout(n23619));
  jand g23407(.dina(n23619), .dinb(n23613), .dout(n23620));
  jxor g23408(.dina(n23620), .dinb(n23612), .dout(n23621));
  jxor g23409(.dina(n23621), .dinb(n23596), .dout(n23622));
  jxor g23410(.dina(n23622), .dinb(n23591), .dout(n23623));
  jxor g23411(.dina(n23623), .dinb(n23582), .dout(n23624));
  jnot g23412(.din(n23624), .dout(n23625));
  jand g23413(.dina(n20141), .dinb(n75), .dout(n23626));
  jand g23414(.dina(n19541), .dinb(n4933), .dout(n23627));
  jand g23415(.dina(n19543), .dinb(n4918), .dout(n23628));
  jand g23416(.dina(n19545), .dinb(n4745), .dout(n23629));
  jor  g23417(.dina(n23629), .dinb(n23628), .dout(n23630));
  jor  g23418(.dina(n23630), .dinb(n23627), .dout(n23631));
  jor  g23419(.dina(n23631), .dinb(n23626), .dout(n23632));
  jxor g23420(.dina(n23632), .dinb(n68), .dout(n23633));
  jxor g23421(.dina(n23633), .dinb(n23625), .dout(n23634));
  jxor g23422(.dina(n23634), .dinb(n23579), .dout(n23635));
  jxor g23423(.dina(n23635), .dinb(n23574), .dout(n23636));
  jxor g23424(.dina(n23636), .dinb(n23565), .dout(n23637));
  jnot g23425(.din(n23637), .dout(n23638));
  jand g23426(.dina(n20767), .dinb(n5693), .dout(n23639));
  jand g23427(.dina(n19529), .dinb(n6209), .dout(n23640));
  jand g23428(.dina(n19531), .dinb(n6131), .dout(n23641));
  jand g23429(.dina(n19533), .dinb(n5691), .dout(n23642));
  jor  g23430(.dina(n23642), .dinb(n23641), .dout(n23643));
  jor  g23431(.dina(n23643), .dinb(n23640), .dout(n23644));
  jor  g23432(.dina(n23644), .dinb(n23639), .dout(n23645));
  jxor g23433(.dina(n23645), .dinb(n4247), .dout(n23646));
  jxor g23434(.dina(n23646), .dinb(n23638), .dout(n23647));
  jxor g23435(.dina(n23647), .dinb(n23562), .dout(n23648));
  jxor g23436(.dina(n23648), .dinb(n23557), .dout(n23649));
  jxor g23437(.dina(n23649), .dinb(n23548), .dout(n23650));
  jnot g23438(.din(n23650), .dout(n23651));
  jand g23439(.dina(n21230), .dinb(n6936), .dout(n23652));
  jand g23440(.dina(n19517), .dinb(n7741), .dout(n23653));
  jand g23441(.dina(n19519), .dinb(n7613), .dout(n23654));
  jand g23442(.dina(n19521), .dinb(n6934), .dout(n23655));
  jor  g23443(.dina(n23655), .dinb(n23654), .dout(n23656));
  jor  g23444(.dina(n23656), .dinb(n23653), .dout(n23657));
  jor  g23445(.dina(n23657), .dinb(n23652), .dout(n23658));
  jxor g23446(.dina(n23658), .dinb(n5292), .dout(n23659));
  jxor g23447(.dina(n23659), .dinb(n23651), .dout(n23660));
  jxor g23448(.dina(n23660), .dinb(n23545), .dout(n23661));
  jxor g23449(.dina(n23661), .dinb(n23540), .dout(n23662));
  jxor g23450(.dina(n23662), .dinb(n23531), .dout(n23663));
  jnot g23451(.din(n23663), .dout(n23664));
  jand g23452(.dina(n22250), .dinb(n8771), .dout(n23665));
  jand g23453(.dina(n22248), .dinb(n9491), .dout(n23666));
  jand g23454(.dina(n19758), .dinb(n9126), .dout(n23667));
  jand g23455(.dina(n19510), .dinb(n8769), .dout(n23668));
  jor  g23456(.dina(n23668), .dinb(n23667), .dout(n23669));
  jor  g23457(.dina(n23669), .dinb(n23666), .dout(n23670));
  jor  g23458(.dina(n23670), .dinb(n23665), .dout(n23671));
  jxor g23459(.dina(n23671), .dinb(n6039), .dout(n23672));
  jxor g23460(.dina(n23672), .dinb(n23664), .dout(n23673));
  jxor g23461(.dina(n23673), .dinb(n23528), .dout(n23674));
  jxor g23462(.dina(n23674), .dinb(n23523), .dout(n23675));
  jxor g23463(.dina(n23675), .dinb(n23514), .dout(n23676));
  jnot g23464(.din(n23676), .dout(n23677));
  jor  g23465(.dina(n23496), .dinb(n23450), .dout(n23678));
  jnot g23466(.din(n23493), .dout(n23679));
  jor  g23467(.dina(n23679), .dinb(n23455), .dout(n23680));
  jand g23468(.dina(n23680), .dinb(n23678), .dout(n23681));
  jand g23469(.dina(n23490), .dinb(n23463), .dout(n23682));
  jand g23470(.dina(n23491), .dinb(n23458), .dout(n23683));
  jor  g23471(.dina(n23683), .dinb(n23682), .dout(n23684));
  jand g23472(.dina(n23488), .dinb(n23481), .dout(n23685));
  jand g23473(.dina(n23489), .dinb(n23473), .dout(n23686));
  jor  g23474(.dina(n23686), .dinb(n23685), .dout(n23687));
  jand g23475(.dina(n23464), .dinb(n23234), .dout(n23688));
  jand g23476(.dina(n23472), .dinb(n23466), .dout(n23689));
  jor  g23477(.dina(n23689), .dinb(n23688), .dout(n23690));
  jand g23478(.dina(n4460), .dinb(n4452), .dout(n23691));
  jxor g23479(.dina(n23691), .dinb(\a[29] ), .dout(n23693));
  jxor g23480(.dina(n23464), .dinb(n24127), .dout(n23694));
  jxor g23481(.dina(n23694), .dinb(n23693), .dout(n23695));
  jand g23482(.dina(n13022), .dinb(n732), .dout(n23696));
  jand g23483(.dina(n12815), .dinb(n3858), .dout(n23697));
  jor  g23484(.dina(n23909), .dinb(n23697), .dout(n23701));
  jor  g23485(.dina(n23701), .dinb(n23696), .dout(n23702));
  jxor g23486(.dina(n23702), .dinb(n23695), .dout(n23703));
  jxor g23487(.dina(n23703), .dinb(n23690), .dout(n23704));
  jxor g23488(.dina(n23704), .dinb(n23687), .dout(n23705));
  jxor g23489(.dina(n23705), .dinb(n23684), .dout(n23706));
  jxor g23490(.dina(n23706), .dinb(n23492), .dout(n23707));
  jxor g23491(.dina(n23707), .dinb(n23681), .dout(n23708));
  jor  g23492(.dina(n23708), .dinb(n10847), .dout(n23709));
  jnot g23493(.din(n23706), .dout(n23710));
  jor  g23494(.dina(n23710), .dinb(n11458), .dout(n23711));
  jor  g23495(.dina(n23496), .dinb(n11360), .dout(n23712));
  jor  g23496(.dina(n23450), .dinb(n10845), .dout(n23713));
  jand g23497(.dina(n23713), .dinb(n23712), .dout(n23714));
  jand g23498(.dina(n23714), .dinb(n23711), .dout(n23715));
  jand g23499(.dina(n23715), .dinb(n23709), .dout(n23716));
  jxor g23500(.dina(n23716), .dinb(\a[2] ), .dout(n23717));
  jxor g23501(.dina(n23717), .dinb(n23677), .dout(n23718));
  jxor g23502(.dina(n23718), .dinb(n23511), .dout(n23719));
  jxor g23503(.dina(n23719), .dinb(n23507), .dout(\result[2] ));
  jand g23504(.dina(n23719), .dinb(n23507), .dout(n23721));
  jor  g23505(.dina(n23717), .dinb(n23677), .dout(n23722));
  jnot g23506(.din(n23722), .dout(n23723));
  jand g23507(.dina(n23718), .dinb(n23511), .dout(n23724));
  jor  g23508(.dina(n23724), .dinb(n23723), .dout(n23725));
  jand g23509(.dina(n23674), .dinb(n23523), .dout(n23726));
  jand g23510(.dina(n23675), .dinb(n23514), .dout(n23727));
  jor  g23511(.dina(n23727), .dinb(n23726), .dout(n23728));
  jnot g23512(.din(n23728), .dout(n23729));
  jnot g23513(.din(n23262), .dout(n23730));
  jor  g23514(.dina(n23730), .dinb(n9919), .dout(n23731));
  jor  g23515(.dina(n23450), .dinb(n10826), .dout(n23732));
  jor  g23516(.dina(n23449), .dinb(n10351), .dout(n23733));
  jnot g23517(.din(n22539), .dout(n23734));
  jor  g23518(.dina(n23734), .dinb(n9918), .dout(n23735));
  jand g23519(.dina(n23735), .dinb(n23733), .dout(n23736));
  jand g23520(.dina(n23736), .dinb(n23732), .dout(n23737));
  jand g23521(.dina(n23737), .dinb(n23731), .dout(n23738));
  jxor g23522(.dina(n23738), .dinb(\a[5] ), .dout(n23739));
  jnot g23523(.din(n23739), .dout(n23740));
  jor  g23524(.dina(n23672), .dinb(n23664), .dout(n23741));
  jand g23525(.dina(n23673), .dinb(n23528), .dout(n23742));
  jnot g23526(.din(n23742), .dout(n23743));
  jand g23527(.dina(n23743), .dinb(n23741), .dout(n23744));
  jnot g23528(.din(n23744), .dout(n23745));
  jand g23529(.dina(n23661), .dinb(n23540), .dout(n23746));
  jand g23530(.dina(n23662), .dinb(n23531), .dout(n23747));
  jor  g23531(.dina(n23747), .dinb(n23746), .dout(n23748));
  jand g23532(.dina(n21750), .dinb(n7890), .dout(n23749));
  jand g23533(.dina(n19510), .dinb(n8441), .dout(n23750));
  jand g23534(.dina(n19511), .dinb(n8154), .dout(n23751));
  jand g23535(.dina(n19513), .dinb(n7888), .dout(n23752));
  jor  g23536(.dina(n23752), .dinb(n23751), .dout(n23753));
  jor  g23537(.dina(n23753), .dinb(n23750), .dout(n23754));
  jor  g23538(.dina(n23754), .dinb(n23749), .dout(n23755));
  jxor g23539(.dina(n23755), .dinb(n5833), .dout(n23756));
  jnot g23540(.din(n23756), .dout(n23757));
  jor  g23541(.dina(n23659), .dinb(n23651), .dout(n23758));
  jand g23542(.dina(n23660), .dinb(n23545), .dout(n23759));
  jnot g23543(.din(n23759), .dout(n23760));
  jand g23544(.dina(n23760), .dinb(n23758), .dout(n23761));
  jnot g23545(.din(n23761), .dout(n23762));
  jand g23546(.dina(n23648), .dinb(n23557), .dout(n23763));
  jand g23547(.dina(n23649), .dinb(n23548), .dout(n23764));
  jor  g23548(.dina(n23764), .dinb(n23763), .dout(n23765));
  jand g23549(.dina(n21086), .dinb(n6340), .dout(n23766));
  jand g23550(.dina(n19521), .dinb(n6798), .dout(n23767));
  jand g23551(.dina(n19523), .dinb(n6556), .dout(n23768));
  jand g23552(.dina(n19525), .dinb(n6338), .dout(n23769));
  jor  g23553(.dina(n23769), .dinb(n23768), .dout(n23770));
  jor  g23554(.dina(n23770), .dinb(n23767), .dout(n23771));
  jor  g23555(.dina(n23771), .dinb(n23766), .dout(n23772));
  jxor g23556(.dina(n23772), .dinb(n5064), .dout(n23773));
  jnot g23557(.din(n23773), .dout(n23774));
  jor  g23558(.dina(n23646), .dinb(n23638), .dout(n23775));
  jand g23559(.dina(n23647), .dinb(n23562), .dout(n23776));
  jnot g23560(.din(n23776), .dout(n23777));
  jand g23561(.dina(n23777), .dinb(n23775), .dout(n23778));
  jnot g23562(.din(n23778), .dout(n23779));
  jand g23563(.dina(n23635), .dinb(n23574), .dout(n23780));
  jand g23564(.dina(n23636), .dinb(n23565), .dout(n23781));
  jor  g23565(.dina(n23781), .dinb(n23780), .dout(n23782));
  jand g23566(.dina(n20399), .dinb(n5365), .dout(n23783));
  jand g23567(.dina(n19533), .dinb(n5500), .dout(n23784));
  jand g23568(.dina(n19535), .dinb(n5424), .dout(n23785));
  jand g23569(.dina(n19537), .dinb(n5363), .dout(n23786));
  jor  g23570(.dina(n23786), .dinb(n23785), .dout(n23787));
  jor  g23571(.dina(n23787), .dinb(n23784), .dout(n23788));
  jor  g23572(.dina(n23788), .dinb(n23783), .dout(n23789));
  jxor g23573(.dina(n23789), .dinb(n72), .dout(n23790));
  jnot g23574(.din(n23790), .dout(n23791));
  jor  g23575(.dina(n23633), .dinb(n23625), .dout(n23792));
  jand g23576(.dina(n23634), .dinb(n23579), .dout(n23793));
  jnot g23577(.din(n23793), .dout(n23794));
  jand g23578(.dina(n23794), .dinb(n23792), .dout(n23795));
  jnot g23579(.din(n23795), .dout(n23796));
  jand g23580(.dina(n23622), .dinb(n23591), .dout(n23797));
  jand g23581(.dina(n23623), .dinb(n23582), .dout(n23798));
  jor  g23582(.dina(n23798), .dinb(n23797), .dout(n23799));
  jand g23583(.dina(n20079), .dinb(n4449), .dout(n23800));
  jand g23584(.dina(n19545), .dinb(n4453), .dout(n23801));
  jand g23585(.dina(n19548), .dinb(n4457), .dout(n23802));
  jand g23586(.dina(n19551), .dinb(n4461), .dout(n23803));
  jor  g23587(.dina(n23803), .dinb(n23802), .dout(n23804));
  jor  g23588(.dina(n23804), .dinb(n23801), .dout(n23805));
  jor  g23589(.dina(n23805), .dinb(n23800), .dout(n23806));
  jxor g23590(.dina(n23806), .dinb(n88), .dout(n23807));
  jnot g23591(.din(n23807), .dout(n23808));
  jor  g23592(.dina(n23620), .dinb(n23612), .dout(n23809));
  jand g23593(.dina(n23621), .dinb(n23596), .dout(n23810));
  jnot g23594(.din(n23810), .dout(n23811));
  jand g23595(.dina(n23811), .dinb(n23809), .dout(n23812));
  jnot g23596(.din(n23812), .dout(n23813));
  jand g23597(.dina(n924), .dinb(n146), .dout(n23814));
  jand g23598(.dina(n23814), .dinb(n1506), .dout(n23815));
  jand g23599(.dina(n23815), .dinb(n2573), .dout(n23816));
  jand g23600(.dina(n5589), .dinb(n2552), .dout(n23817));
  jand g23601(.dina(n23817), .dinb(n23816), .dout(n23818));
  jand g23602(.dina(n1281), .dinb(n1067), .dout(n23819));
  jand g23603(.dina(n23819), .dinb(n1334), .dout(n23820));
  jand g23604(.dina(n3189), .dinb(n960), .dout(n23821));
  jand g23605(.dina(n23821), .dinb(n798), .dout(n23822));
  jand g23606(.dina(n23822), .dinb(n23820), .dout(n23823));
  jand g23607(.dina(n23823), .dinb(n23818), .dout(n23824));
  jand g23608(.dina(n23824), .dinb(n14211), .dout(n23825));
  jand g23609(.dina(n23825), .dinb(n3001), .dout(n23826));
  jand g23610(.dina(n7459), .dinb(n3949), .dout(n23827));
  jand g23611(.dina(n23827), .dinb(n23826), .dout(n23828));
  jor  g23612(.dina(n19964), .dinb(n6463), .dout(n23829));
  jand g23613(.dina(n19554), .dinb(n3855), .dout(n23830));
  jand g23614(.dina(n23384), .dinb(n3851), .dout(n23831));
  jand g23615(.dina(n19559), .dinb(n3858), .dout(n23832));
  jor  g23616(.dina(n23832), .dinb(n23831), .dout(n23833));
  jor  g23617(.dina(n23833), .dinb(n23830), .dout(n23834));
  jnot g23618(.din(n23834), .dout(n23835));
  jand g23619(.dina(n23835), .dinb(n23829), .dout(n23836));
  jxor g23620(.dina(n23836), .dinb(n23828), .dout(n23837));
  jxor g23621(.dina(n23837), .dinb(n23813), .dout(n23838));
  jxor g23622(.dina(n23838), .dinb(n23808), .dout(n23839));
  jxor g23623(.dina(n23839), .dinb(n23799), .dout(n23840));
  jnot g23624(.din(n23840), .dout(n23841));
  jand g23625(.dina(n20131), .dinb(n75), .dout(n23842));
  jand g23626(.dina(n19539), .dinb(n4933), .dout(n23843));
  jand g23627(.dina(n19541), .dinb(n4918), .dout(n23844));
  jand g23628(.dina(n19543), .dinb(n4745), .dout(n23845));
  jor  g23629(.dina(n23845), .dinb(n23844), .dout(n23846));
  jor  g23630(.dina(n23846), .dinb(n23843), .dout(n23847));
  jor  g23631(.dina(n23847), .dinb(n23842), .dout(n23848));
  jxor g23632(.dina(n23848), .dinb(n68), .dout(n23849));
  jxor g23633(.dina(n23849), .dinb(n23841), .dout(n23850));
  jxor g23634(.dina(n23850), .dinb(n23796), .dout(n23851));
  jxor g23635(.dina(n23851), .dinb(n23791), .dout(n23852));
  jxor g23636(.dina(n23852), .dinb(n23782), .dout(n23853));
  jnot g23637(.din(n23853), .dout(n23854));
  jand g23638(.dina(n20793), .dinb(n5693), .dout(n23855));
  jand g23639(.dina(n19527), .dinb(n6209), .dout(n23856));
  jand g23640(.dina(n19529), .dinb(n6131), .dout(n23857));
  jand g23641(.dina(n19531), .dinb(n5691), .dout(n23858));
  jor  g23642(.dina(n23858), .dinb(n23857), .dout(n23859));
  jor  g23643(.dina(n23859), .dinb(n23856), .dout(n23860));
  jor  g23644(.dina(n23860), .dinb(n23855), .dout(n23861));
  jxor g23645(.dina(n23861), .dinb(n4247), .dout(n23862));
  jxor g23646(.dina(n23862), .dinb(n23854), .dout(n23863));
  jxor g23647(.dina(n23863), .dinb(n23779), .dout(n23864));
  jxor g23648(.dina(n23864), .dinb(n23774), .dout(n23865));
  jxor g23649(.dina(n23865), .dinb(n23765), .dout(n23866));
  jnot g23650(.din(n23866), .dout(n23867));
  jand g23651(.dina(n21218), .dinb(n6936), .dout(n23868));
  jand g23652(.dina(n19515), .dinb(n7741), .dout(n23869));
  jand g23653(.dina(n19517), .dinb(n7613), .dout(n23870));
  jand g23654(.dina(n19519), .dinb(n6934), .dout(n23871));
  jor  g23655(.dina(n23871), .dinb(n23870), .dout(n23872));
  jor  g23656(.dina(n23872), .dinb(n23869), .dout(n23873));
  jor  g23657(.dina(n23873), .dinb(n23868), .dout(n23874));
  jxor g23658(.dina(n23874), .dinb(n5292), .dout(n23875));
  jxor g23659(.dina(n23875), .dinb(n23867), .dout(n23876));
  jxor g23660(.dina(n23876), .dinb(n23762), .dout(n23877));
  jxor g23661(.dina(n23877), .dinb(n23757), .dout(n23878));
  jxor g23662(.dina(n23878), .dinb(n23748), .dout(n23879));
  jnot g23663(.din(n23879), .dout(n23880));
  jand g23664(.dina(n22627), .dinb(n8771), .dout(n23881));
  jand g23665(.dina(n22540), .dinb(n9491), .dout(n23882));
  jand g23666(.dina(n22248), .dinb(n9126), .dout(n23883));
  jand g23667(.dina(n19758), .dinb(n8769), .dout(n23884));
  jor  g23668(.dina(n23884), .dinb(n23883), .dout(n23885));
  jor  g23669(.dina(n23885), .dinb(n23882), .dout(n23886));
  jor  g23670(.dina(n23886), .dinb(n23881), .dout(n23887));
  jxor g23671(.dina(n23887), .dinb(n6039), .dout(n23888));
  jxor g23672(.dina(n23888), .dinb(n23880), .dout(n23889));
  jxor g23673(.dina(n23889), .dinb(n23745), .dout(n23890));
  jxor g23674(.dina(n23890), .dinb(n23740), .dout(n23891));
  jxor g23675(.dina(n23891), .dinb(n23729), .dout(n23892));
  jor  g23676(.dina(n23710), .dinb(n23496), .dout(n23893));
  jnot g23677(.din(n23707), .dout(n23894));
  jor  g23678(.dina(n23894), .dinb(n23681), .dout(n23895));
  jand g23679(.dina(n23895), .dinb(n23893), .dout(n23896));
  jand g23680(.dina(n23702), .dinb(n23695), .dout(n23897));
  jand g23681(.dina(n23703), .dinb(n23690), .dout(n23898));
  jor  g23682(.dina(n23898), .dinb(n23897), .dout(n23899));
  jand g23683(.dina(n23694), .dinb(n23693), .dout(n23902));
  jor  g23684(.dina(n23902), .dinb(n23465), .dout(n23903));
  jxor g23685(.dina(n23903), .dinb(n4594), .dout(n23904));
  jor  g23686(.dina(n3855), .dinb(n3851), .dout(n23909));
  jor  g23687(.dina(n23909), .dinb(n3858), .dout(n23910));
  jor  g23688(.dina(n23910), .dinb(n732), .dout(n23911));
  jxor g23689(.dina(n23911), .dinb(n23904), .dout(n23912));
  jxor g23690(.dina(n23912), .dinb(n23899), .dout(n23913));
  jand g23691(.dina(n23704), .dinb(n23687), .dout(n23914));
  jand g23692(.dina(n23705), .dinb(n23684), .dout(n23915));
  jor  g23693(.dina(n23915), .dinb(n23914), .dout(n23916));
  jxor g23694(.dina(n23916), .dinb(n23913), .dout(n23917));
  jxor g23695(.dina(n23917), .dinb(n23706), .dout(n23918));
  jxor g23696(.dina(n23918), .dinb(n23896), .dout(n23919));
  jor  g23697(.dina(n23919), .dinb(n10847), .dout(n23920));
  jnot g23698(.din(n23917), .dout(n23921));
  jor  g23699(.dina(n23921), .dinb(n11458), .dout(n23922));
  jor  g23700(.dina(n23710), .dinb(n11360), .dout(n23923));
  jor  g23701(.dina(n23496), .dinb(n10845), .dout(n23924));
  jand g23702(.dina(n23924), .dinb(n23923), .dout(n23925));
  jand g23703(.dina(n23925), .dinb(n23922), .dout(n23926));
  jand g23704(.dina(n23926), .dinb(n23920), .dout(n23927));
  jxor g23705(.dina(n23927), .dinb(\a[2] ), .dout(n23928));
  jxor g23706(.dina(n23928), .dinb(n23892), .dout(n23929));
  jxor g23707(.dina(n23929), .dinb(n23725), .dout(n23930));
  jxor g23708(.dina(n23930), .dinb(n23721), .dout(\result[3] ));
  jand g23709(.dina(n23930), .dinb(n23721), .dout(n23932));
  jor  g23710(.dina(n23928), .dinb(n23892), .dout(n23933));
  jnot g23711(.din(n23933), .dout(n23934));
  jand g23712(.dina(n23929), .dinb(n23725), .dout(n23935));
  jor  g23713(.dina(n23935), .dinb(n23934), .dout(n23936));
  jand g23714(.dina(n23890), .dinb(n23740), .dout(n23937));
  jnot g23715(.din(n23937), .dout(n23938));
  jnot g23716(.din(n23891), .dout(n23939));
  jor  g23717(.dina(n23939), .dinb(n23729), .dout(n23940));
  jand g23718(.dina(n23940), .dinb(n23938), .dout(n23941));
  jor  g23719(.dina(n23494), .dinb(n9919), .dout(n23942));
  jor  g23720(.dina(n23496), .dinb(n10826), .dout(n23943));
  jor  g23721(.dina(n23450), .dinb(n10351), .dout(n23944));
  jor  g23722(.dina(n23449), .dinb(n9918), .dout(n23945));
  jand g23723(.dina(n23945), .dinb(n23944), .dout(n23946));
  jand g23724(.dina(n23946), .dinb(n23943), .dout(n23947));
  jand g23725(.dina(n23947), .dinb(n23942), .dout(n23948));
  jxor g23726(.dina(n23948), .dinb(\a[5] ), .dout(n23949));
  jnot g23727(.din(n23949), .dout(n23950));
  jor  g23728(.dina(n23888), .dinb(n23880), .dout(n23951));
  jnot g23729(.din(n23951), .dout(n23952));
  jand g23730(.dina(n23889), .dinb(n23745), .dout(n23953));
  jor  g23731(.dina(n23953), .dinb(n23952), .dout(n23954));
  jand g23732(.dina(n23877), .dinb(n23757), .dout(n23955));
  jand g23733(.dina(n23878), .dinb(n23748), .dout(n23956));
  jor  g23734(.dina(n23956), .dinb(n23955), .dout(n23957));
  jand g23735(.dina(n19760), .dinb(n7890), .dout(n23958));
  jand g23736(.dina(n19758), .dinb(n8441), .dout(n23959));
  jand g23737(.dina(n19510), .dinb(n8154), .dout(n23960));
  jand g23738(.dina(n19511), .dinb(n7888), .dout(n23961));
  jor  g23739(.dina(n23961), .dinb(n23960), .dout(n23962));
  jor  g23740(.dina(n23962), .dinb(n23959), .dout(n23963));
  jor  g23741(.dina(n23963), .dinb(n23958), .dout(n23964));
  jxor g23742(.dina(n23964), .dinb(n5833), .dout(n23965));
  jnot g23743(.din(n23965), .dout(n23966));
  jor  g23744(.dina(n23875), .dinb(n23867), .dout(n23967));
  jand g23745(.dina(n23876), .dinb(n23762), .dout(n23968));
  jnot g23746(.din(n23968), .dout(n23969));
  jand g23747(.dina(n23969), .dinb(n23967), .dout(n23970));
  jnot g23748(.din(n23970), .dout(n23971));
  jand g23749(.dina(n23864), .dinb(n23774), .dout(n23972));
  jand g23750(.dina(n23865), .dinb(n23765), .dout(n23973));
  jor  g23751(.dina(n23973), .dinb(n23972), .dout(n23974));
  jand g23752(.dina(n21240), .dinb(n6340), .dout(n23975));
  jand g23753(.dina(n19519), .dinb(n6798), .dout(n23976));
  jand g23754(.dina(n19521), .dinb(n6556), .dout(n23977));
  jand g23755(.dina(n19523), .dinb(n6338), .dout(n23978));
  jor  g23756(.dina(n23978), .dinb(n23977), .dout(n23979));
  jor  g23757(.dina(n23979), .dinb(n23976), .dout(n23980));
  jor  g23758(.dina(n23980), .dinb(n23975), .dout(n23981));
  jxor g23759(.dina(n23981), .dinb(n5064), .dout(n23982));
  jnot g23760(.din(n23982), .dout(n23983));
  jor  g23761(.dina(n23862), .dinb(n23854), .dout(n23984));
  jand g23762(.dina(n23863), .dinb(n23779), .dout(n23985));
  jnot g23763(.din(n23985), .dout(n23986));
  jand g23764(.dina(n23986), .dinb(n23984), .dout(n23987));
  jnot g23765(.din(n23987), .dout(n23988));
  jand g23766(.dina(n23851), .dinb(n23791), .dout(n23989));
  jand g23767(.dina(n23852), .dinb(n23782), .dout(n23990));
  jor  g23768(.dina(n23990), .dinb(n23989), .dout(n23991));
  jand g23769(.dina(n19780), .dinb(n5365), .dout(n23992));
  jand g23770(.dina(n19531), .dinb(n5500), .dout(n23993));
  jand g23771(.dina(n19533), .dinb(n5424), .dout(n23994));
  jand g23772(.dina(n19535), .dinb(n5363), .dout(n23995));
  jor  g23773(.dina(n23995), .dinb(n23994), .dout(n23996));
  jor  g23774(.dina(n23996), .dinb(n23993), .dout(n23997));
  jor  g23775(.dina(n23997), .dinb(n23992), .dout(n23998));
  jxor g23776(.dina(n23998), .dinb(n72), .dout(n23999));
  jnot g23777(.din(n23999), .dout(n24000));
  jor  g23778(.dina(n23849), .dinb(n23841), .dout(n24001));
  jand g23779(.dina(n23850), .dinb(n23796), .dout(n24002));
  jnot g23780(.din(n24002), .dout(n24003));
  jand g23781(.dina(n24003), .dinb(n24001), .dout(n24004));
  jnot g23782(.din(n24004), .dout(n24005));
  jand g23783(.dina(n23838), .dinb(n23808), .dout(n24006));
  jand g23784(.dina(n23839), .dinb(n23799), .dout(n24007));
  jor  g23785(.dina(n24007), .dinb(n24006), .dout(n24008));
  jand g23786(.dina(n20153), .dinb(n4449), .dout(n24009));
  jand g23787(.dina(n19543), .dinb(n4453), .dout(n24010));
  jand g23788(.dina(n19545), .dinb(n4457), .dout(n24011));
  jand g23789(.dina(n19548), .dinb(n4461), .dout(n24012));
  jor  g23790(.dina(n24012), .dinb(n24011), .dout(n24013));
  jor  g23791(.dina(n24013), .dinb(n24010), .dout(n24014));
  jor  g23792(.dina(n24014), .dinb(n24009), .dout(n24015));
  jxor g23793(.dina(n24015), .dinb(n88), .dout(n24016));
  jnot g23794(.din(n24016), .dout(n24017));
  jor  g23795(.dina(n23836), .dinb(n23828), .dout(n24018));
  jand g23796(.dina(n23837), .dinb(n23813), .dout(n24019));
  jnot g23797(.din(n24019), .dout(n24020));
  jand g23798(.dina(n24020), .dinb(n24018), .dout(n24021));
  jnot g23799(.din(n24021), .dout(n24022));
  jand g23800(.dina(n2538), .dinb(n880), .dout(n24023));
  jand g23801(.dina(n939), .dinb(n717), .dout(n24024));
  jand g23802(.dina(n24024), .dinb(n24023), .dout(n24025));
  jand g23803(.dina(n5902), .dinb(n2872), .dout(n24026));
  jand g23804(.dina(n3819), .dinb(n451), .dout(n24027));
  jand g23805(.dina(n24027), .dinb(n24026), .dout(n24028));
  jand g23806(.dina(n24028), .dinb(n24025), .dout(n24029));
  jand g23807(.dina(n24029), .dinb(n2842), .dout(n24030));
  jand g23808(.dina(n13094), .dinb(n6627), .dout(n24031));
  jand g23809(.dina(n2483), .dinb(n1259), .dout(n24032));
  jand g23810(.dina(n24032), .dinb(n24031), .dout(n24033));
  jand g23811(.dina(n503), .dinb(n383), .dout(n24034));
  jand g23812(.dina(n860), .dinb(n1031), .dout(n24035));
  jand g23813(.dina(n24035), .dinb(n24034), .dout(n24036));
  jand g23814(.dina(n2870), .dinb(n1023), .dout(n24037));
  jand g23815(.dina(n24037), .dinb(n24036), .dout(n24038));
  jand g23816(.dina(n24038), .dinb(n24033), .dout(n24039));
  jand g23817(.dina(n876), .dinb(n763), .dout(n24040));
  jand g23818(.dina(n24040), .dinb(n626), .dout(n24041));
  jand g23819(.dina(n24041), .dinb(n2210), .dout(n24042));
  jand g23820(.dina(n2042), .dinb(n977), .dout(n24043));
  jand g23821(.dina(n24043), .dinb(n24042), .dout(n24044));
  jand g23822(.dina(n24044), .dinb(n24039), .dout(n24045));
  jand g23823(.dina(n24045), .dinb(n24030), .dout(n24046));
  jand g23824(.dina(n24046), .dinb(n4156), .dout(n24047));
  jand g23825(.dina(n24047), .dinb(n5241), .dout(n24048));
  jor  g23826(.dina(n19952), .dinb(n6463), .dout(n24049));
  jand g23827(.dina(n19551), .dinb(n3855), .dout(n24050));
  jand g23828(.dina(n19559), .dinb(n3851), .dout(n24051));
  jand g23829(.dina(n19554), .dinb(n3858), .dout(n24052));
  jor  g23830(.dina(n24052), .dinb(n24051), .dout(n24053));
  jor  g23831(.dina(n24053), .dinb(n24050), .dout(n24054));
  jnot g23832(.din(n24054), .dout(n24055));
  jand g23833(.dina(n24055), .dinb(n24049), .dout(n24056));
  jxor g23834(.dina(n24056), .dinb(n24048), .dout(n24057));
  jxor g23835(.dina(n24057), .dinb(n24022), .dout(n24058));
  jxor g23836(.dina(n24058), .dinb(n24017), .dout(n24059));
  jxor g23837(.dina(n24059), .dinb(n24008), .dout(n24060));
  jnot g23838(.din(n24060), .dout(n24061));
  jand g23839(.dina(n20387), .dinb(n75), .dout(n24062));
  jand g23840(.dina(n19537), .dinb(n4933), .dout(n24063));
  jand g23841(.dina(n19539), .dinb(n4918), .dout(n24064));
  jand g23842(.dina(n19541), .dinb(n4745), .dout(n24065));
  jor  g23843(.dina(n24065), .dinb(n24064), .dout(n24066));
  jor  g23844(.dina(n24066), .dinb(n24063), .dout(n24067));
  jor  g23845(.dina(n24067), .dinb(n24062), .dout(n24068));
  jxor g23846(.dina(n24068), .dinb(n68), .dout(n24069));
  jxor g23847(.dina(n24069), .dinb(n24061), .dout(n24070));
  jxor g23848(.dina(n24070), .dinb(n24005), .dout(n24071));
  jxor g23849(.dina(n24071), .dinb(n24000), .dout(n24072));
  jxor g23850(.dina(n24072), .dinb(n23991), .dout(n24073));
  jnot g23851(.din(n24073), .dout(n24074));
  jand g23852(.dina(n20781), .dinb(n5693), .dout(n24075));
  jand g23853(.dina(n19525), .dinb(n6209), .dout(n24076));
  jand g23854(.dina(n19527), .dinb(n6131), .dout(n24077));
  jand g23855(.dina(n19529), .dinb(n5691), .dout(n24078));
  jor  g23856(.dina(n24078), .dinb(n24077), .dout(n24079));
  jor  g23857(.dina(n24079), .dinb(n24076), .dout(n24080));
  jor  g23858(.dina(n24080), .dinb(n24075), .dout(n24081));
  jxor g23859(.dina(n24081), .dinb(n4247), .dout(n24082));
  jxor g23860(.dina(n24082), .dinb(n24074), .dout(n24083));
  jxor g23861(.dina(n24083), .dinb(n23988), .dout(n24084));
  jxor g23862(.dina(n24084), .dinb(n23983), .dout(n24085));
  jxor g23863(.dina(n24085), .dinb(n23974), .dout(n24086));
  jnot g23864(.din(n24086), .dout(n24087));
  jand g23865(.dina(n21738), .dinb(n6936), .dout(n24088));
  jand g23866(.dina(n19513), .dinb(n7741), .dout(n24089));
  jand g23867(.dina(n19515), .dinb(n7613), .dout(n24090));
  jand g23868(.dina(n19517), .dinb(n6934), .dout(n24091));
  jor  g23869(.dina(n24091), .dinb(n24090), .dout(n24092));
  jor  g23870(.dina(n24092), .dinb(n24089), .dout(n24093));
  jor  g23871(.dina(n24093), .dinb(n24088), .dout(n24094));
  jxor g23872(.dina(n24094), .dinb(n5292), .dout(n24095));
  jxor g23873(.dina(n24095), .dinb(n24087), .dout(n24096));
  jxor g23874(.dina(n24096), .dinb(n23971), .dout(n24097));
  jxor g23875(.dina(n24097), .dinb(n23966), .dout(n24098));
  jxor g23876(.dina(n24098), .dinb(n23957), .dout(n24099));
  jnot g23877(.din(n24099), .dout(n24100));
  jand g23878(.dina(n22617), .dinb(n8771), .dout(n24101));
  jand g23879(.dina(n22539), .dinb(n9491), .dout(n24102));
  jand g23880(.dina(n22540), .dinb(n9126), .dout(n24103));
  jand g23881(.dina(n22248), .dinb(n8769), .dout(n24104));
  jor  g23882(.dina(n24104), .dinb(n24103), .dout(n24105));
  jor  g23883(.dina(n24105), .dinb(n24102), .dout(n24106));
  jor  g23884(.dina(n24106), .dinb(n24101), .dout(n24107));
  jxor g23885(.dina(n24107), .dinb(n6039), .dout(n24108));
  jxor g23886(.dina(n24108), .dinb(n24100), .dout(n24109));
  jxor g23887(.dina(n24109), .dinb(n23954), .dout(n24110));
  jxor g23888(.dina(n24110), .dinb(n23950), .dout(n24111));
  jxor g23889(.dina(n24111), .dinb(n23941), .dout(n24112));
  jor  g23890(.dina(n23921), .dinb(n23710), .dout(n24113));
  jnot g23891(.din(n23918), .dout(n24114));
  jor  g23892(.dina(n24114), .dinb(n23896), .dout(n24115));
  jand g23893(.dina(n24115), .dinb(n24113), .dout(n24116));
  jnot g23894(.din(n3858), .dout(n24120));
  jand g23895(.dina(n24120), .dinb(n3854), .dout(n24121));
  jand g23896(.dina(n24121), .dinb(n27660), .dout(n24122));
  jor  g23897(.dina(n24122), .dinb(n12460), .dout(n24123));
  jand g23898(.dina(n24123), .dinb(n6463), .dout(n24124));
  jxor g23899(.dina(n24124), .dinb(n4594), .dout(n24125));
  jnot g23900(.din(n24125), .dout(n24126));
  jnot g23901(.din(n4594), .dout(n24127));
  jxor g23902(.dina(n4594), .dinb(n24126), .dout(n24134));
  jand g23903(.dina(n23912), .dinb(n23899), .dout(n24135));
  jand g23904(.dina(n23916), .dinb(n23913), .dout(n24136));
  jor  g23905(.dina(n24136), .dinb(n24135), .dout(n24137));
  jxor g23906(.dina(n24137), .dinb(n24134), .dout(n24138));
  jxor g23907(.dina(n24138), .dinb(n23917), .dout(n24139));
  jxor g23908(.dina(n24139), .dinb(n24116), .dout(n24140));
  jor  g23909(.dina(n24140), .dinb(n10847), .dout(n24141));
  jnot g23910(.din(n24138), .dout(n24142));
  jor  g23911(.dina(n24142), .dinb(n11458), .dout(n24143));
  jor  g23912(.dina(n23921), .dinb(n11360), .dout(n24144));
  jor  g23913(.dina(n23710), .dinb(n10845), .dout(n24145));
  jand g23914(.dina(n24145), .dinb(n24144), .dout(n24146));
  jand g23915(.dina(n24146), .dinb(n24143), .dout(n24147));
  jand g23916(.dina(n24147), .dinb(n24141), .dout(n24148));
  jxor g23917(.dina(n24148), .dinb(\a[2] ), .dout(n24149));
  jxor g23918(.dina(n24149), .dinb(n24112), .dout(n24150));
  jxor g23919(.dina(n24150), .dinb(n23936), .dout(n24151));
  jxor g23920(.dina(n24151), .dinb(n23932), .dout(\result[4] ));
  jand g23921(.dina(n24151), .dinb(n23932), .dout(n24153));
  jor  g23922(.dina(n24149), .dinb(n24112), .dout(n24154));
  jnot g23923(.din(n24154), .dout(n24155));
  jand g23924(.dina(n24150), .dinb(n23936), .dout(n24156));
  jor  g23925(.dina(n24156), .dinb(n24155), .dout(n24157));
  jand g23926(.dina(n24110), .dinb(n23950), .dout(n24158));
  jnot g23927(.din(n24158), .dout(n24159));
  jnot g23928(.din(n24111), .dout(n24160));
  jor  g23929(.dina(n24160), .dinb(n23941), .dout(n24161));
  jand g23930(.dina(n24161), .dinb(n24159), .dout(n24162));
  jor  g23931(.dina(n23708), .dinb(n9919), .dout(n24163));
  jor  g23932(.dina(n23710), .dinb(n10826), .dout(n24164));
  jor  g23933(.dina(n23496), .dinb(n10351), .dout(n24165));
  jor  g23934(.dina(n23450), .dinb(n9918), .dout(n24166));
  jand g23935(.dina(n24166), .dinb(n24165), .dout(n24167));
  jand g23936(.dina(n24167), .dinb(n24164), .dout(n24168));
  jand g23937(.dina(n24168), .dinb(n24163), .dout(n24169));
  jxor g23938(.dina(n24169), .dinb(\a[5] ), .dout(n24170));
  jnot g23939(.din(n24170), .dout(n24171));
  jor  g23940(.dina(n24108), .dinb(n24100), .dout(n24172));
  jnot g23941(.din(n24172), .dout(n24173));
  jand g23942(.dina(n24109), .dinb(n23954), .dout(n24174));
  jor  g23943(.dina(n24174), .dinb(n24173), .dout(n24175));
  jand g23944(.dina(n24097), .dinb(n23966), .dout(n24176));
  jand g23945(.dina(n24098), .dinb(n23957), .dout(n24177));
  jor  g23946(.dina(n24177), .dinb(n24176), .dout(n24178));
  jand g23947(.dina(n22250), .dinb(n7890), .dout(n24179));
  jand g23948(.dina(n22248), .dinb(n8441), .dout(n24180));
  jand g23949(.dina(n19758), .dinb(n8154), .dout(n24181));
  jand g23950(.dina(n19510), .dinb(n7888), .dout(n24182));
  jor  g23951(.dina(n24182), .dinb(n24181), .dout(n24183));
  jor  g23952(.dina(n24183), .dinb(n24180), .dout(n24184));
  jor  g23953(.dina(n24184), .dinb(n24179), .dout(n24185));
  jxor g23954(.dina(n24185), .dinb(n5833), .dout(n24186));
  jnot g23955(.din(n24186), .dout(n24187));
  jor  g23956(.dina(n24095), .dinb(n24087), .dout(n24188));
  jand g23957(.dina(n24096), .dinb(n23971), .dout(n24189));
  jnot g23958(.din(n24189), .dout(n24190));
  jand g23959(.dina(n24190), .dinb(n24188), .dout(n24191));
  jnot g23960(.din(n24191), .dout(n24192));
  jand g23961(.dina(n24084), .dinb(n23983), .dout(n24193));
  jand g23962(.dina(n24085), .dinb(n23974), .dout(n24194));
  jor  g23963(.dina(n24194), .dinb(n24193), .dout(n24195));
  jand g23964(.dina(n21230), .dinb(n6340), .dout(n24196));
  jand g23965(.dina(n19517), .dinb(n6798), .dout(n24197));
  jand g23966(.dina(n19519), .dinb(n6556), .dout(n24198));
  jand g23967(.dina(n19521), .dinb(n6338), .dout(n24199));
  jor  g23968(.dina(n24199), .dinb(n24198), .dout(n24200));
  jor  g23969(.dina(n24200), .dinb(n24197), .dout(n24201));
  jor  g23970(.dina(n24201), .dinb(n24196), .dout(n24202));
  jxor g23971(.dina(n24202), .dinb(n5064), .dout(n24203));
  jnot g23972(.din(n24203), .dout(n24204));
  jor  g23973(.dina(n24082), .dinb(n24074), .dout(n24205));
  jand g23974(.dina(n24083), .dinb(n23988), .dout(n24206));
  jnot g23975(.din(n24206), .dout(n24207));
  jand g23976(.dina(n24207), .dinb(n24205), .dout(n24208));
  jnot g23977(.din(n24208), .dout(n24209));
  jand g23978(.dina(n24071), .dinb(n24000), .dout(n24210));
  jand g23979(.dina(n24072), .dinb(n23991), .dout(n24211));
  jor  g23980(.dina(n24211), .dinb(n24210), .dout(n24212));
  jand g23981(.dina(n20767), .dinb(n5365), .dout(n24213));
  jand g23982(.dina(n19529), .dinb(n5500), .dout(n24214));
  jand g23983(.dina(n19531), .dinb(n5424), .dout(n24215));
  jand g23984(.dina(n19533), .dinb(n5363), .dout(n24216));
  jor  g23985(.dina(n24216), .dinb(n24215), .dout(n24217));
  jor  g23986(.dina(n24217), .dinb(n24214), .dout(n24218));
  jor  g23987(.dina(n24218), .dinb(n24213), .dout(n24219));
  jxor g23988(.dina(n24219), .dinb(n72), .dout(n24220));
  jnot g23989(.din(n24220), .dout(n24221));
  jor  g23990(.dina(n24069), .dinb(n24061), .dout(n24222));
  jand g23991(.dina(n24070), .dinb(n24005), .dout(n24223));
  jnot g23992(.din(n24223), .dout(n24224));
  jand g23993(.dina(n24224), .dinb(n24222), .dout(n24225));
  jnot g23994(.din(n24225), .dout(n24226));
  jand g23995(.dina(n24058), .dinb(n24017), .dout(n24227));
  jand g23996(.dina(n24059), .dinb(n24008), .dout(n24228));
  jor  g23997(.dina(n24228), .dinb(n24227), .dout(n24229));
  jand g23998(.dina(n20141), .dinb(n4449), .dout(n24230));
  jand g23999(.dina(n19541), .dinb(n4453), .dout(n24231));
  jand g24000(.dina(n19543), .dinb(n4457), .dout(n24232));
  jand g24001(.dina(n19545), .dinb(n4461), .dout(n24233));
  jor  g24002(.dina(n24233), .dinb(n24232), .dout(n24234));
  jor  g24003(.dina(n24234), .dinb(n24231), .dout(n24235));
  jor  g24004(.dina(n24235), .dinb(n24230), .dout(n24236));
  jxor g24005(.dina(n24236), .dinb(n88), .dout(n24237));
  jnot g24006(.din(n24237), .dout(n24238));
  jor  g24007(.dina(n24056), .dinb(n24048), .dout(n24239));
  jand g24008(.dina(n24057), .dinb(n24022), .dout(n24240));
  jnot g24009(.din(n24240), .dout(n24241));
  jand g24010(.dina(n24241), .dinb(n24239), .dout(n24242));
  jnot g24011(.din(n24242), .dout(n24243));
  jand g24012(.dina(n1142), .dinb(n1048), .dout(n24244));
  jand g24013(.dina(n24244), .dinb(n13149), .dout(n24245));
  jand g24014(.dina(n24245), .dinb(n3954), .dout(n24246));
  jand g24015(.dina(n24246), .dinb(n962), .dout(n24247));
  jand g24016(.dina(n551), .dinb(n270), .dout(n24248));
  jand g24017(.dina(n24248), .dinb(n305), .dout(n24249));
  jand g24018(.dina(n407), .dinb(n357), .dout(n24250));
  jand g24019(.dina(n24250), .dinb(n12267), .dout(n24251));
  jand g24020(.dina(n12696), .dinb(n1603), .dout(n24252));
  jand g24021(.dina(n24252), .dinb(n24251), .dout(n24253));
  jand g24022(.dina(n24253), .dinb(n24249), .dout(n24254));
  jand g24023(.dina(n24254), .dinb(n3893), .dout(n24255));
  jand g24024(.dina(n24255), .dinb(n24247), .dout(n24256));
  jand g24025(.dina(n24256), .dinb(n6004), .dout(n24257));
  jand g24026(.dina(n24257), .dinb(n14417), .dout(n24258));
  jor  g24027(.dina(n19940), .dinb(n6463), .dout(n24259));
  jand g24028(.dina(n19548), .dinb(n3855), .dout(n24260));
  jand g24029(.dina(n19554), .dinb(n3851), .dout(n24261));
  jand g24030(.dina(n19551), .dinb(n3858), .dout(n24262));
  jor  g24031(.dina(n24262), .dinb(n24261), .dout(n24263));
  jor  g24032(.dina(n24263), .dinb(n24260), .dout(n24264));
  jnot g24033(.din(n24264), .dout(n24265));
  jand g24034(.dina(n24265), .dinb(n24259), .dout(n24266));
  jxor g24035(.dina(n24266), .dinb(n24258), .dout(n24267));
  jxor g24036(.dina(n24267), .dinb(n24243), .dout(n24268));
  jxor g24037(.dina(n24268), .dinb(n24238), .dout(n24269));
  jxor g24038(.dina(n24269), .dinb(n24229), .dout(n24270));
  jnot g24039(.din(n24270), .dout(n24271));
  jand g24040(.dina(n20413), .dinb(n75), .dout(n24272));
  jand g24041(.dina(n19535), .dinb(n4933), .dout(n24273));
  jand g24042(.dina(n19537), .dinb(n4918), .dout(n24274));
  jand g24043(.dina(n19539), .dinb(n4745), .dout(n24275));
  jor  g24044(.dina(n24275), .dinb(n24274), .dout(n24276));
  jor  g24045(.dina(n24276), .dinb(n24273), .dout(n24277));
  jor  g24046(.dina(n24277), .dinb(n24272), .dout(n24278));
  jxor g24047(.dina(n24278), .dinb(n68), .dout(n24279));
  jxor g24048(.dina(n24279), .dinb(n24271), .dout(n24280));
  jxor g24049(.dina(n24280), .dinb(n24226), .dout(n24281));
  jxor g24050(.dina(n24281), .dinb(n24221), .dout(n24282));
  jxor g24051(.dina(n24282), .dinb(n24212), .dout(n24283));
  jnot g24052(.din(n24283), .dout(n24284));
  jand g24053(.dina(n19770), .dinb(n5693), .dout(n24285));
  jand g24054(.dina(n19523), .dinb(n6209), .dout(n24286));
  jand g24055(.dina(n19525), .dinb(n6131), .dout(n24287));
  jand g24056(.dina(n19527), .dinb(n5691), .dout(n24288));
  jor  g24057(.dina(n24288), .dinb(n24287), .dout(n24289));
  jor  g24058(.dina(n24289), .dinb(n24286), .dout(n24290));
  jor  g24059(.dina(n24290), .dinb(n24285), .dout(n24291));
  jxor g24060(.dina(n24291), .dinb(n4247), .dout(n24292));
  jxor g24061(.dina(n24292), .dinb(n24284), .dout(n24293));
  jxor g24062(.dina(n24293), .dinb(n24209), .dout(n24294));
  jxor g24063(.dina(n24294), .dinb(n24204), .dout(n24295));
  jxor g24064(.dina(n24295), .dinb(n24195), .dout(n24296));
  jnot g24065(.din(n24296), .dout(n24297));
  jand g24066(.dina(n21762), .dinb(n6936), .dout(n24298));
  jand g24067(.dina(n19511), .dinb(n7741), .dout(n24299));
  jand g24068(.dina(n19513), .dinb(n7613), .dout(n24300));
  jand g24069(.dina(n19515), .dinb(n6934), .dout(n24301));
  jor  g24070(.dina(n24301), .dinb(n24300), .dout(n24302));
  jor  g24071(.dina(n24302), .dinb(n24299), .dout(n24303));
  jor  g24072(.dina(n24303), .dinb(n24298), .dout(n24304));
  jxor g24073(.dina(n24304), .dinb(n5292), .dout(n24305));
  jxor g24074(.dina(n24305), .dinb(n24297), .dout(n24306));
  jxor g24075(.dina(n24306), .dinb(n24192), .dout(n24307));
  jxor g24076(.dina(n24307), .dinb(n24187), .dout(n24308));
  jxor g24077(.dina(n24308), .dinb(n24178), .dout(n24309));
  jnot g24078(.din(n24309), .dout(n24310));
  jand g24079(.dina(n22605), .dinb(n8771), .dout(n24311));
  jand g24080(.dina(n22603), .dinb(n9491), .dout(n24312));
  jand g24081(.dina(n22539), .dinb(n9126), .dout(n24313));
  jand g24082(.dina(n22540), .dinb(n8769), .dout(n24314));
  jor  g24083(.dina(n24314), .dinb(n24313), .dout(n24315));
  jor  g24084(.dina(n24315), .dinb(n24312), .dout(n24316));
  jor  g24085(.dina(n24316), .dinb(n24311), .dout(n24317));
  jxor g24086(.dina(n24317), .dinb(n6039), .dout(n24318));
  jxor g24087(.dina(n24318), .dinb(n24310), .dout(n24319));
  jxor g24088(.dina(n24319), .dinb(n24175), .dout(n24320));
  jxor g24089(.dina(n24320), .dinb(n24171), .dout(n24321));
  jxor g24090(.dina(n24321), .dinb(n24162), .dout(n24322));
  jor  g24091(.dina(n24142), .dinb(n23921), .dout(n24323));
  jnot g24092(.din(n24139), .dout(n24324));
  jor  g24093(.dina(n24324), .dinb(n24116), .dout(n24325));
  jand g24094(.dina(n24325), .dinb(n24323), .dout(n24326));
  jand g24095(.dina(n24137), .dinb(n24134), .dout(n24328));
  jor  g24096(.dina(n24328), .dinb(n24330), .dout(n24329));
  jand g24097(.dina(n24124), .dinb(n4594), .dout(n24330));
  jnot g24098(.din(\a[31] ), .dout(n24331));
  jand g24099(.dina(n126), .dinb(n24331), .dout(n24332));
  jor  g24100(.dina(n24332), .dinb(n12460), .dout(n24333));
  jxor g24101(.dina(n24333), .dinb(n24330), .dout(n24334));
  jxor g24102(.dina(n24334), .dinb(n24329), .dout(n24335));
  jxor g24103(.dina(n24335), .dinb(n24142), .dout(n24336));
  jxor g24104(.dina(n24336), .dinb(n24326), .dout(n24337));
  jor  g24105(.dina(n24337), .dinb(n10847), .dout(n24338));
  jor  g24106(.dina(n24335), .dinb(n11458), .dout(n24339));
  jor  g24107(.dina(n24142), .dinb(n11360), .dout(n24340));
  jor  g24108(.dina(n23921), .dinb(n10845), .dout(n24341));
  jand g24109(.dina(n24341), .dinb(n24340), .dout(n24342));
  jand g24110(.dina(n24342), .dinb(n24339), .dout(n24343));
  jand g24111(.dina(n24343), .dinb(n24338), .dout(n24344));
  jxor g24112(.dina(n24344), .dinb(\a[2] ), .dout(n24345));
  jxor g24113(.dina(n24345), .dinb(n24322), .dout(n24346));
  jxor g24114(.dina(n24346), .dinb(n24157), .dout(n24347));
  jxor g24115(.dina(n24347), .dinb(n24153), .dout(\result[5] ));
  jand g24116(.dina(n24347), .dinb(n24153), .dout(n24349));
  jand g24117(.dina(n24320), .dinb(n24171), .dout(n24350));
  jnot g24118(.din(n24162), .dout(n24351));
  jand g24119(.dina(n24321), .dinb(n24351), .dout(n24352));
  jor  g24120(.dina(n24352), .dinb(n24350), .dout(n24353));
  jor  g24121(.dina(n24335), .dinb(n24142), .dout(n24354));
  jnot g24122(.din(n24336), .dout(n24355));
  jor  g24123(.dina(n24355), .dinb(n24326), .dout(n24356));
  jand g24124(.dina(n24356), .dinb(n24354), .dout(n24357));
  jor  g24125(.dina(n24357), .dinb(n10847), .dout(n24358));
  jor  g24126(.dina(n24335), .dinb(n11469), .dout(n24359));
  jor  g24127(.dina(n24142), .dinb(n10845), .dout(n24360));
  jand g24128(.dina(n24360), .dinb(n24359), .dout(n24361));
  jand g24129(.dina(n24361), .dinb(n24358), .dout(n24362));
  jxor g24130(.dina(n24362), .dinb(\a[2] ), .dout(n24363));
  jnot g24131(.din(n24363), .dout(n24364));
  jor  g24132(.dina(n23919), .dinb(n9919), .dout(n24365));
  jor  g24133(.dina(n23921), .dinb(n10826), .dout(n24366));
  jor  g24134(.dina(n23710), .dinb(n10351), .dout(n24367));
  jor  g24135(.dina(n23496), .dinb(n9918), .dout(n24368));
  jand g24136(.dina(n24368), .dinb(n24367), .dout(n24369));
  jand g24137(.dina(n24369), .dinb(n24366), .dout(n24370));
  jand g24138(.dina(n24370), .dinb(n24365), .dout(n24371));
  jxor g24139(.dina(n24371), .dinb(\a[5] ), .dout(n24372));
  jnot g24140(.din(n24372), .dout(n24373));
  jor  g24141(.dina(n24318), .dinb(n24310), .dout(n24374));
  jnot g24142(.din(n24374), .dout(n24375));
  jand g24143(.dina(n24319), .dinb(n24175), .dout(n24376));
  jor  g24144(.dina(n24376), .dinb(n24375), .dout(n24377));
  jand g24145(.dina(n24307), .dinb(n24187), .dout(n24378));
  jand g24146(.dina(n24308), .dinb(n24178), .dout(n24379));
  jor  g24147(.dina(n24379), .dinb(n24378), .dout(n24380));
  jand g24148(.dina(n22627), .dinb(n7890), .dout(n24381));
  jand g24149(.dina(n22540), .dinb(n8441), .dout(n24382));
  jand g24150(.dina(n22248), .dinb(n8154), .dout(n24383));
  jand g24151(.dina(n19758), .dinb(n7888), .dout(n24384));
  jor  g24152(.dina(n24384), .dinb(n24383), .dout(n24385));
  jor  g24153(.dina(n24385), .dinb(n24382), .dout(n24386));
  jor  g24154(.dina(n24386), .dinb(n24381), .dout(n24387));
  jxor g24155(.dina(n24387), .dinb(n5833), .dout(n24388));
  jnot g24156(.din(n24388), .dout(n24389));
  jor  g24157(.dina(n24305), .dinb(n24297), .dout(n24390));
  jand g24158(.dina(n24306), .dinb(n24192), .dout(n24391));
  jnot g24159(.din(n24391), .dout(n24392));
  jand g24160(.dina(n24392), .dinb(n24390), .dout(n24393));
  jnot g24161(.din(n24393), .dout(n24394));
  jand g24162(.dina(n24294), .dinb(n24204), .dout(n24395));
  jand g24163(.dina(n24295), .dinb(n24195), .dout(n24396));
  jor  g24164(.dina(n24396), .dinb(n24395), .dout(n24397));
  jand g24165(.dina(n21218), .dinb(n6340), .dout(n24398));
  jand g24166(.dina(n19515), .dinb(n6798), .dout(n24399));
  jand g24167(.dina(n19517), .dinb(n6556), .dout(n24400));
  jand g24168(.dina(n19519), .dinb(n6338), .dout(n24401));
  jor  g24169(.dina(n24401), .dinb(n24400), .dout(n24402));
  jor  g24170(.dina(n24402), .dinb(n24399), .dout(n24403));
  jor  g24171(.dina(n24403), .dinb(n24398), .dout(n24404));
  jxor g24172(.dina(n24404), .dinb(n5064), .dout(n24405));
  jnot g24173(.din(n24405), .dout(n24406));
  jor  g24174(.dina(n24292), .dinb(n24284), .dout(n24407));
  jand g24175(.dina(n24293), .dinb(n24209), .dout(n24408));
  jnot g24176(.din(n24408), .dout(n24409));
  jand g24177(.dina(n24409), .dinb(n24407), .dout(n24410));
  jnot g24178(.din(n24410), .dout(n24411));
  jand g24179(.dina(n24281), .dinb(n24221), .dout(n24412));
  jand g24180(.dina(n24282), .dinb(n24212), .dout(n24413));
  jor  g24181(.dina(n24413), .dinb(n24412), .dout(n24414));
  jand g24182(.dina(n20793), .dinb(n5365), .dout(n24415));
  jand g24183(.dina(n19527), .dinb(n5500), .dout(n24416));
  jand g24184(.dina(n19529), .dinb(n5424), .dout(n24417));
  jand g24185(.dina(n19531), .dinb(n5363), .dout(n24418));
  jor  g24186(.dina(n24418), .dinb(n24417), .dout(n24419));
  jor  g24187(.dina(n24419), .dinb(n24416), .dout(n24420));
  jor  g24188(.dina(n24420), .dinb(n24415), .dout(n24421));
  jxor g24189(.dina(n24421), .dinb(n72), .dout(n24422));
  jnot g24190(.din(n24422), .dout(n24423));
  jor  g24191(.dina(n24279), .dinb(n24271), .dout(n24424));
  jand g24192(.dina(n24280), .dinb(n24226), .dout(n24425));
  jnot g24193(.din(n24425), .dout(n24426));
  jand g24194(.dina(n24426), .dinb(n24424), .dout(n24427));
  jnot g24195(.din(n24427), .dout(n24428));
  jand g24196(.dina(n24268), .dinb(n24238), .dout(n24429));
  jand g24197(.dina(n24269), .dinb(n24229), .dout(n24430));
  jor  g24198(.dina(n24430), .dinb(n24429), .dout(n24431));
  jand g24199(.dina(n20131), .dinb(n4449), .dout(n24432));
  jand g24200(.dina(n19539), .dinb(n4453), .dout(n24433));
  jand g24201(.dina(n19541), .dinb(n4457), .dout(n24434));
  jand g24202(.dina(n19543), .dinb(n4461), .dout(n24435));
  jor  g24203(.dina(n24435), .dinb(n24434), .dout(n24436));
  jor  g24204(.dina(n24436), .dinb(n24433), .dout(n24437));
  jor  g24205(.dina(n24437), .dinb(n24432), .dout(n24438));
  jxor g24206(.dina(n24438), .dinb(n88), .dout(n24439));
  jnot g24207(.din(n24439), .dout(n24440));
  jor  g24208(.dina(n24266), .dinb(n24258), .dout(n24441));
  jand g24209(.dina(n24267), .dinb(n24243), .dout(n24442));
  jnot g24210(.din(n24442), .dout(n24443));
  jand g24211(.dina(n24443), .dinb(n24441), .dout(n24444));
  jnot g24212(.din(n24444), .dout(n24445));
  jand g24213(.dina(n2322), .dinb(n1492), .dout(n24446));
  jand g24214(.dina(n24446), .dinb(n506), .dout(n24447));
  jand g24215(.dina(n24447), .dinb(n23820), .dout(n24448));
  jand g24216(.dina(n24448), .dinb(n13248), .dout(n24449));
  jand g24217(.dina(n3491), .dinb(n2401), .dout(n24450));
  jand g24218(.dina(n5755), .dinb(n2514), .dout(n24451));
  jand g24219(.dina(n24451), .dinb(n3788), .dout(n24452));
  jand g24220(.dina(n24452), .dinb(n24450), .dout(n24453));
  jand g24221(.dina(n5198), .dinb(n1137), .dout(n24454));
  jand g24222(.dina(n3819), .dinb(n2653), .dout(n24455));
  jand g24223(.dina(n24455), .dinb(n24454), .dout(n24456));
  jand g24224(.dina(n354), .dinb(n268), .dout(n24457));
  jand g24225(.dina(n24457), .dinb(n1422), .dout(n24458));
  jand g24226(.dina(n24458), .dinb(n1877), .dout(n24459));
  jand g24227(.dina(n24459), .dinb(n24456), .dout(n24460));
  jand g24228(.dina(n24460), .dinb(n24453), .dout(n24461));
  jand g24229(.dina(n24461), .dinb(n24449), .dout(n24462));
  jand g24230(.dina(n13623), .dinb(n5776), .dout(n24463));
  jand g24231(.dina(n24463), .dinb(n3245), .dout(n24464));
  jand g24232(.dina(n24464), .dinb(n24462), .dout(n24465));
  jnot g24233(.din(n24465), .dout(n24466));
  jand g24234(.dina(n20079), .dinb(n732), .dout(n24467));
  jand g24235(.dina(n19545), .dinb(n3855), .dout(n24468));
  jand g24236(.dina(n19551), .dinb(n3851), .dout(n24469));
  jand g24237(.dina(n19548), .dinb(n3858), .dout(n24470));
  jor  g24238(.dina(n24470), .dinb(n24469), .dout(n24471));
  jor  g24239(.dina(n24471), .dinb(n24468), .dout(n24472));
  jor  g24240(.dina(n24472), .dinb(n24467), .dout(n24473));
  jxor g24241(.dina(n24473), .dinb(n24466), .dout(n24474));
  jxor g24242(.dina(n24474), .dinb(n24445), .dout(n24475));
  jxor g24243(.dina(n24475), .dinb(n24440), .dout(n24476));
  jxor g24244(.dina(n24476), .dinb(n24431), .dout(n24477));
  jnot g24245(.din(n24477), .dout(n24478));
  jand g24246(.dina(n20399), .dinb(n75), .dout(n24479));
  jand g24247(.dina(n19533), .dinb(n4933), .dout(n24480));
  jand g24248(.dina(n19535), .dinb(n4918), .dout(n24481));
  jand g24249(.dina(n19537), .dinb(n4745), .dout(n24482));
  jor  g24250(.dina(n24482), .dinb(n24481), .dout(n24483));
  jor  g24251(.dina(n24483), .dinb(n24480), .dout(n24484));
  jor  g24252(.dina(n24484), .dinb(n24479), .dout(n24485));
  jxor g24253(.dina(n24485), .dinb(n68), .dout(n24486));
  jxor g24254(.dina(n24486), .dinb(n24478), .dout(n24487));
  jxor g24255(.dina(n24487), .dinb(n24428), .dout(n24488));
  jxor g24256(.dina(n24488), .dinb(n24423), .dout(n24489));
  jxor g24257(.dina(n24489), .dinb(n24414), .dout(n24490));
  jnot g24258(.din(n24490), .dout(n24491));
  jand g24259(.dina(n21086), .dinb(n5693), .dout(n24492));
  jand g24260(.dina(n19521), .dinb(n6209), .dout(n24493));
  jand g24261(.dina(n19523), .dinb(n6131), .dout(n24494));
  jand g24262(.dina(n19525), .dinb(n5691), .dout(n24495));
  jor  g24263(.dina(n24495), .dinb(n24494), .dout(n24496));
  jor  g24264(.dina(n24496), .dinb(n24493), .dout(n24497));
  jor  g24265(.dina(n24497), .dinb(n24492), .dout(n24498));
  jxor g24266(.dina(n24498), .dinb(n4247), .dout(n24499));
  jxor g24267(.dina(n24499), .dinb(n24491), .dout(n24500));
  jxor g24268(.dina(n24500), .dinb(n24411), .dout(n24501));
  jxor g24269(.dina(n24501), .dinb(n24406), .dout(n24502));
  jxor g24270(.dina(n24502), .dinb(n24397), .dout(n24503));
  jnot g24271(.din(n24503), .dout(n24504));
  jand g24272(.dina(n21750), .dinb(n6936), .dout(n24505));
  jand g24273(.dina(n19510), .dinb(n7741), .dout(n24506));
  jand g24274(.dina(n19511), .dinb(n7613), .dout(n24507));
  jand g24275(.dina(n19513), .dinb(n6934), .dout(n24508));
  jor  g24276(.dina(n24508), .dinb(n24507), .dout(n24509));
  jor  g24277(.dina(n24509), .dinb(n24506), .dout(n24510));
  jor  g24278(.dina(n24510), .dinb(n24505), .dout(n24511));
  jxor g24279(.dina(n24511), .dinb(n5292), .dout(n24512));
  jxor g24280(.dina(n24512), .dinb(n24504), .dout(n24513));
  jxor g24281(.dina(n24513), .dinb(n24394), .dout(n24514));
  jxor g24282(.dina(n24514), .dinb(n24389), .dout(n24515));
  jxor g24283(.dina(n24515), .dinb(n24380), .dout(n24516));
  jnot g24284(.din(n24516), .dout(n24517));
  jand g24285(.dina(n23262), .dinb(n8771), .dout(n24518));
  jand g24286(.dina(n23260), .dinb(n9491), .dout(n24519));
  jand g24287(.dina(n22603), .dinb(n9126), .dout(n24520));
  jand g24288(.dina(n22539), .dinb(n8769), .dout(n24521));
  jor  g24289(.dina(n24521), .dinb(n24520), .dout(n24522));
  jor  g24290(.dina(n24522), .dinb(n24519), .dout(n24523));
  jor  g24291(.dina(n24523), .dinb(n24518), .dout(n24524));
  jxor g24292(.dina(n24524), .dinb(n6039), .dout(n24525));
  jxor g24293(.dina(n24525), .dinb(n24517), .dout(n24526));
  jxor g24294(.dina(n24526), .dinb(n24377), .dout(n24527));
  jxor g24295(.dina(n24527), .dinb(n24373), .dout(n24528));
  jxor g24296(.dina(n24528), .dinb(n24364), .dout(n24529));
  jxor g24297(.dina(n24529), .dinb(n24353), .dout(n24530));
  jor  g24298(.dina(n24345), .dinb(n24322), .dout(n24531));
  jnot g24299(.din(n24531), .dout(n24532));
  jand g24300(.dina(n24346), .dinb(n24157), .dout(n24533));
  jor  g24301(.dina(n24533), .dinb(n24532), .dout(n24534));
  jxor g24302(.dina(n24534), .dinb(n24530), .dout(n24535));
  jxor g24303(.dina(n24535), .dinb(n24349), .dout(\result[6] ));
  jand g24304(.dina(n24535), .dinb(n24349), .dout(n24537));
  jand g24305(.dina(n24527), .dinb(n24373), .dout(n24538));
  jand g24306(.dina(n24528), .dinb(n24364), .dout(n24539));
  jor  g24307(.dina(n24539), .dinb(n24538), .dout(n24540));
  jor  g24308(.dina(n24525), .dinb(n24517), .dout(n24541));
  jand g24309(.dina(n24526), .dinb(n24377), .dout(n24542));
  jnot g24310(.din(n24542), .dout(n24543));
  jand g24311(.dina(n24543), .dinb(n24541), .dout(n24544));
  jand g24312(.dina(n24514), .dinb(n24389), .dout(n24545));
  jand g24313(.dina(n24515), .dinb(n24380), .dout(n24546));
  jor  g24314(.dina(n24546), .dinb(n24545), .dout(n24547));
  jor  g24315(.dina(n24512), .dinb(n24504), .dout(n24548));
  jand g24316(.dina(n24513), .dinb(n24394), .dout(n24549));
  jnot g24317(.din(n24549), .dout(n24550));
  jand g24318(.dina(n24550), .dinb(n24548), .dout(n24551));
  jnot g24319(.din(n24551), .dout(n24552));
  jand g24320(.dina(n24501), .dinb(n24406), .dout(n24553));
  jand g24321(.dina(n24502), .dinb(n24397), .dout(n24554));
  jor  g24322(.dina(n24554), .dinb(n24553), .dout(n24555));
  jor  g24323(.dina(n24499), .dinb(n24491), .dout(n24556));
  jand g24324(.dina(n24500), .dinb(n24411), .dout(n24557));
  jnot g24325(.din(n24557), .dout(n24558));
  jand g24326(.dina(n24558), .dinb(n24556), .dout(n24559));
  jnot g24327(.din(n24559), .dout(n24560));
  jand g24328(.dina(n24488), .dinb(n24423), .dout(n24561));
  jand g24329(.dina(n24489), .dinb(n24414), .dout(n24562));
  jor  g24330(.dina(n24562), .dinb(n24561), .dout(n24563));
  jor  g24331(.dina(n24486), .dinb(n24478), .dout(n24564));
  jand g24332(.dina(n24487), .dinb(n24428), .dout(n24565));
  jnot g24333(.din(n24565), .dout(n24566));
  jand g24334(.dina(n24566), .dinb(n24564), .dout(n24567));
  jnot g24335(.din(n24567), .dout(n24568));
  jand g24336(.dina(n24475), .dinb(n24440), .dout(n24569));
  jand g24337(.dina(n24476), .dinb(n24431), .dout(n24570));
  jor  g24338(.dina(n24570), .dinb(n24569), .dout(n24571));
  jand g24339(.dina(n24473), .dinb(n24466), .dout(n24572));
  jand g24340(.dina(n24474), .dinb(n24445), .dout(n24573));
  jor  g24341(.dina(n24573), .dinb(n24572), .dout(n24574));
  jnot g24342(.din(n3357), .dout(n24575));
  jand g24343(.dina(n612), .dinb(n553), .dout(n24576));
  jand g24344(.dina(n692), .dinb(n197), .dout(n24577));
  jand g24345(.dina(n24577), .dinb(n24576), .dout(n24578));
  jand g24346(.dina(n24578), .dinb(n12556), .dout(n24579));
  jand g24347(.dina(n13075), .dinb(n2905), .dout(n24580));
  jand g24348(.dina(n24580), .dinb(n24579), .dout(n24581));
  jand g24349(.dina(n842), .dinb(n154), .dout(n24582));
  jand g24350(.dina(n24582), .dinb(n1009), .dout(n24583));
  jand g24351(.dina(n5898), .dinb(n436), .dout(n24584));
  jand g24352(.dina(n24584), .dinb(n24583), .dout(n24585));
  jand g24353(.dina(n24585), .dinb(n7426), .dout(n24586));
  jand g24354(.dina(n24586), .dinb(n24581), .dout(n24587));
  jand g24355(.dina(n4412), .dinb(n2716), .dout(n24588));
  jand g24356(.dina(n24588), .dinb(n12734), .dout(n24589));
  jand g24357(.dina(n24589), .dinb(n24587), .dout(n24590));
  jand g24358(.dina(n24590), .dinb(n24575), .dout(n24591));
  jand g24359(.dina(n24591), .dinb(n3799), .dout(n24592));
  jnot g24360(.din(n24335), .dout(n24593));
  jand g24361(.dina(n24593), .dinb(n13650), .dout(n24594));
  jand g24362(.dina(n24335), .dinb(n6600), .dout(n24595));
  jor  g24363(.dina(n24595), .dinb(n24594), .dout(n24596));
  jxor g24364(.dina(n24596), .dinb(n24592), .dout(n24597));
  jand g24365(.dina(n20153), .dinb(n732), .dout(n24598));
  jand g24366(.dina(n19543), .dinb(n3855), .dout(n24599));
  jand g24367(.dina(n19545), .dinb(n3858), .dout(n24600));
  jand g24368(.dina(n19548), .dinb(n3851), .dout(n24601));
  jor  g24369(.dina(n24601), .dinb(n24600), .dout(n24602));
  jor  g24370(.dina(n24602), .dinb(n24599), .dout(n24603));
  jor  g24371(.dina(n24603), .dinb(n24598), .dout(n24604));
  jxor g24372(.dina(n24604), .dinb(n24597), .dout(n24605));
  jxor g24373(.dina(n24605), .dinb(n24574), .dout(n24606));
  jnot g24374(.din(n24606), .dout(n24607));
  jand g24375(.dina(n20387), .dinb(n4449), .dout(n24608));
  jand g24376(.dina(n19537), .dinb(n4453), .dout(n24609));
  jand g24377(.dina(n19539), .dinb(n4457), .dout(n24610));
  jand g24378(.dina(n19541), .dinb(n4461), .dout(n24611));
  jor  g24379(.dina(n24611), .dinb(n24610), .dout(n24612));
  jor  g24380(.dina(n24612), .dinb(n24609), .dout(n24613));
  jor  g24381(.dina(n24613), .dinb(n24608), .dout(n24614));
  jxor g24382(.dina(n24614), .dinb(n88), .dout(n24615));
  jxor g24383(.dina(n24615), .dinb(n24607), .dout(n24616));
  jxor g24384(.dina(n24616), .dinb(n24571), .dout(n24617));
  jand g24385(.dina(n19780), .dinb(n75), .dout(n24618));
  jand g24386(.dina(n19531), .dinb(n4933), .dout(n24619));
  jand g24387(.dina(n19533), .dinb(n4918), .dout(n24620));
  jand g24388(.dina(n19535), .dinb(n4745), .dout(n24621));
  jor  g24389(.dina(n24621), .dinb(n24620), .dout(n24622));
  jor  g24390(.dina(n24622), .dinb(n24619), .dout(n24623));
  jor  g24391(.dina(n24623), .dinb(n24618), .dout(n24624));
  jxor g24392(.dina(n24624), .dinb(n68), .dout(n24625));
  jnot g24393(.din(n24625), .dout(n24626));
  jxor g24394(.dina(n24626), .dinb(n24617), .dout(n24627));
  jxor g24395(.dina(n24627), .dinb(n24568), .dout(n24628));
  jand g24396(.dina(n20781), .dinb(n5365), .dout(n24629));
  jand g24397(.dina(n19525), .dinb(n5500), .dout(n24630));
  jand g24398(.dina(n19527), .dinb(n5424), .dout(n24631));
  jand g24399(.dina(n19529), .dinb(n5363), .dout(n24632));
  jor  g24400(.dina(n24632), .dinb(n24631), .dout(n24633));
  jor  g24401(.dina(n24633), .dinb(n24630), .dout(n24634));
  jor  g24402(.dina(n24634), .dinb(n24629), .dout(n24635));
  jxor g24403(.dina(n24635), .dinb(n72), .dout(n24636));
  jnot g24404(.din(n24636), .dout(n24637));
  jxor g24405(.dina(n24637), .dinb(n24628), .dout(n24638));
  jxor g24406(.dina(n24638), .dinb(n24563), .dout(n24639));
  jand g24407(.dina(n21240), .dinb(n5693), .dout(n24640));
  jand g24408(.dina(n19519), .dinb(n6209), .dout(n24641));
  jand g24409(.dina(n19521), .dinb(n6131), .dout(n24642));
  jand g24410(.dina(n19523), .dinb(n5691), .dout(n24643));
  jor  g24411(.dina(n24643), .dinb(n24642), .dout(n24644));
  jor  g24412(.dina(n24644), .dinb(n24641), .dout(n24645));
  jor  g24413(.dina(n24645), .dinb(n24640), .dout(n24646));
  jxor g24414(.dina(n24646), .dinb(n4247), .dout(n24647));
  jnot g24415(.din(n24647), .dout(n24648));
  jxor g24416(.dina(n24648), .dinb(n24639), .dout(n24649));
  jxor g24417(.dina(n24649), .dinb(n24560), .dout(n24650));
  jand g24418(.dina(n21738), .dinb(n6340), .dout(n24651));
  jand g24419(.dina(n19513), .dinb(n6798), .dout(n24652));
  jand g24420(.dina(n19515), .dinb(n6556), .dout(n24653));
  jand g24421(.dina(n19517), .dinb(n6338), .dout(n24654));
  jor  g24422(.dina(n24654), .dinb(n24653), .dout(n24655));
  jor  g24423(.dina(n24655), .dinb(n24652), .dout(n24656));
  jor  g24424(.dina(n24656), .dinb(n24651), .dout(n24657));
  jxor g24425(.dina(n24657), .dinb(n5064), .dout(n24658));
  jnot g24426(.din(n24658), .dout(n24659));
  jxor g24427(.dina(n24659), .dinb(n24650), .dout(n24660));
  jxor g24428(.dina(n24660), .dinb(n24555), .dout(n24661));
  jand g24429(.dina(n19760), .dinb(n6936), .dout(n24662));
  jand g24430(.dina(n19758), .dinb(n7741), .dout(n24663));
  jand g24431(.dina(n19510), .dinb(n7613), .dout(n24664));
  jand g24432(.dina(n19511), .dinb(n6934), .dout(n24665));
  jor  g24433(.dina(n24665), .dinb(n24664), .dout(n24666));
  jor  g24434(.dina(n24666), .dinb(n24663), .dout(n24667));
  jor  g24435(.dina(n24667), .dinb(n24662), .dout(n24668));
  jxor g24436(.dina(n24668), .dinb(n5292), .dout(n24669));
  jnot g24437(.din(n24669), .dout(n24670));
  jxor g24438(.dina(n24670), .dinb(n24661), .dout(n24671));
  jxor g24439(.dina(n24671), .dinb(n24552), .dout(n24672));
  jand g24440(.dina(n22617), .dinb(n7890), .dout(n24673));
  jand g24441(.dina(n22539), .dinb(n8441), .dout(n24674));
  jand g24442(.dina(n22540), .dinb(n8154), .dout(n24675));
  jand g24443(.dina(n22248), .dinb(n7888), .dout(n24676));
  jor  g24444(.dina(n24676), .dinb(n24675), .dout(n24677));
  jor  g24445(.dina(n24677), .dinb(n24674), .dout(n24678));
  jor  g24446(.dina(n24678), .dinb(n24673), .dout(n24679));
  jxor g24447(.dina(n24679), .dinb(n5833), .dout(n24680));
  jnot g24448(.din(n24680), .dout(n24681));
  jxor g24449(.dina(n24681), .dinb(n24672), .dout(n24682));
  jxor g24450(.dina(n24682), .dinb(n24547), .dout(n24683));
  jor  g24451(.dina(n23494), .dinb(n8772), .dout(n24684));
  jor  g24452(.dina(n23496), .dinb(n9490), .dout(n24685));
  jor  g24453(.dina(n23450), .dinb(n9127), .dout(n24686));
  jor  g24454(.dina(n23449), .dinb(n8770), .dout(n24687));
  jand g24455(.dina(n24687), .dinb(n24686), .dout(n24688));
  jand g24456(.dina(n24688), .dinb(n24685), .dout(n24689));
  jand g24457(.dina(n24689), .dinb(n24684), .dout(n24690));
  jxor g24458(.dina(n24690), .dinb(\a[8] ), .dout(n24691));
  jnot g24459(.din(n24691), .dout(n24692));
  jxor g24460(.dina(n24692), .dinb(n24683), .dout(n24693));
  jxor g24461(.dina(n24693), .dinb(n24544), .dout(n24694));
  jor  g24462(.dina(n24140), .dinb(n9919), .dout(n24695));
  jor  g24463(.dina(n24142), .dinb(n10826), .dout(n24696));
  jor  g24464(.dina(n23921), .dinb(n10351), .dout(n24697));
  jor  g24465(.dina(n23710), .dinb(n9918), .dout(n24698));
  jand g24466(.dina(n24698), .dinb(n24697), .dout(n24699));
  jand g24467(.dina(n24699), .dinb(n24696), .dout(n24700));
  jand g24468(.dina(n24700), .dinb(n24695), .dout(n24701));
  jxor g24469(.dina(n24701), .dinb(\a[5] ), .dout(n24702));
  jxor g24470(.dina(n24702), .dinb(n24694), .dout(n24703));
  jxor g24471(.dina(n24703), .dinb(n24540), .dout(n24704));
  jand g24472(.dina(n24529), .dinb(n24353), .dout(n24705));
  jand g24473(.dina(n24534), .dinb(n24530), .dout(n24706));
  jor  g24474(.dina(n24706), .dinb(n24705), .dout(n24707));
  jxor g24475(.dina(n24707), .dinb(n24704), .dout(n24708));
  jxor g24476(.dina(n24708), .dinb(n24537), .dout(\result[7] ));
  jand g24477(.dina(n24708), .dinb(n24537), .dout(n24710));
  jand g24478(.dina(n20767), .dinb(n75), .dout(n24711));
  jand g24479(.dina(n19529), .dinb(n4933), .dout(n24712));
  jand g24480(.dina(n19531), .dinb(n4918), .dout(n24713));
  jand g24481(.dina(n19533), .dinb(n4745), .dout(n24714));
  jor  g24482(.dina(n24714), .dinb(n24713), .dout(n24715));
  jor  g24483(.dina(n24715), .dinb(n24712), .dout(n24716));
  jor  g24484(.dina(n24716), .dinb(n24711), .dout(n24717));
  jxor g24485(.dina(n24717), .dinb(n68), .dout(n24718));
  jnot g24486(.din(n24718), .dout(n24719));
  jand g24487(.dina(n24605), .dinb(n24574), .dout(n24720));
  jnot g24488(.din(n24720), .dout(n24721));
  jor  g24489(.dina(n24615), .dinb(n24607), .dout(n24722));
  jand g24490(.dina(n24722), .dinb(n24721), .dout(n24723));
  jnot g24491(.din(n24723), .dout(n24724));
  jand g24492(.dina(n1178), .dinb(n366), .dout(n24725));
  jand g24493(.dina(n24725), .dinb(n1546), .dout(n24726));
  jand g24494(.dina(n24726), .dinb(n21156), .dout(n24727));
  jand g24495(.dina(n24727), .dinb(n3617), .dout(n24728));
  jand g24496(.dina(n2660), .dinb(n2240), .dout(n24729));
  jand g24497(.dina(n4004), .dinb(n1432), .dout(n24730));
  jand g24498(.dina(n24730), .dinb(n24729), .dout(n24731));
  jand g24499(.dina(n3189), .dinb(n2046), .dout(n24732));
  jand g24500(.dina(n2227), .dinb(n1846), .dout(n24733));
  jand g24501(.dina(n24733), .dinb(n24732), .dout(n24734));
  jand g24502(.dina(n24734), .dinb(n24731), .dout(n24735));
  jand g24503(.dina(n24735), .dinb(n24728), .dout(n24736));
  jand g24504(.dina(n739), .dinb(n194), .dout(n24737));
  jand g24505(.dina(n24737), .dinb(n543), .dout(n24738));
  jand g24506(.dina(n24738), .dinb(n802), .dout(n24739));
  jand g24507(.dina(n24739), .dinb(n14513), .dout(n24740));
  jand g24508(.dina(n24740), .dinb(n2195), .dout(n24741));
  jand g24509(.dina(n24741), .dinb(n24736), .dout(n24742));
  jand g24510(.dina(n24742), .dinb(n14482), .dout(n24743));
  jand g24511(.dina(n24743), .dinb(n2951), .dout(n24744));
  jxor g24512(.dina(n24744), .dinb(n24596), .dout(n24745));
  jand g24513(.dina(n24596), .dinb(n24592), .dout(n24746));
  jnot g24514(.din(n24746), .dout(n24747));
  jnot g24515(.din(n24592), .dout(n24748));
  jnot g24516(.din(n24596), .dout(n24749));
  jand g24517(.dina(n24749), .dinb(n24748), .dout(n24750));
  jor  g24518(.dina(n24604), .dinb(n24750), .dout(n24751));
  jand g24519(.dina(n24751), .dinb(n24747), .dout(n24752));
  jxor g24520(.dina(n24752), .dinb(n24745), .dout(n24753));
  jand g24521(.dina(n20141), .dinb(n732), .dout(n24754));
  jand g24522(.dina(n19541), .dinb(n3855), .dout(n24755));
  jand g24523(.dina(n19543), .dinb(n3858), .dout(n24756));
  jand g24524(.dina(n19545), .dinb(n3851), .dout(n24757));
  jor  g24525(.dina(n24757), .dinb(n24756), .dout(n24758));
  jor  g24526(.dina(n24758), .dinb(n24755), .dout(n24759));
  jor  g24527(.dina(n24759), .dinb(n24754), .dout(n24760));
  jxor g24528(.dina(n24760), .dinb(n24753), .dout(n24761));
  jxor g24529(.dina(n24761), .dinb(n24724), .dout(n24762));
  jnot g24530(.din(n24762), .dout(n24763));
  jand g24531(.dina(n20413), .dinb(n4449), .dout(n24764));
  jand g24532(.dina(n19535), .dinb(n4453), .dout(n24765));
  jand g24533(.dina(n19537), .dinb(n4457), .dout(n24766));
  jand g24534(.dina(n19539), .dinb(n4461), .dout(n24767));
  jor  g24535(.dina(n24767), .dinb(n24766), .dout(n24768));
  jor  g24536(.dina(n24768), .dinb(n24765), .dout(n24769));
  jor  g24537(.dina(n24769), .dinb(n24764), .dout(n24770));
  jxor g24538(.dina(n24770), .dinb(n88), .dout(n24771));
  jxor g24539(.dina(n24771), .dinb(n24763), .dout(n24772));
  jxor g24540(.dina(n24772), .dinb(n24719), .dout(n24773));
  jor  g24541(.dina(n24616), .dinb(n24571), .dout(n24774));
  jand g24542(.dina(n24616), .dinb(n24571), .dout(n24775));
  jor  g24543(.dina(n24626), .dinb(n24775), .dout(n24776));
  jand g24544(.dina(n24776), .dinb(n24774), .dout(n24777));
  jxor g24545(.dina(n24777), .dinb(n24773), .dout(n24778));
  jand g24546(.dina(n19770), .dinb(n5365), .dout(n24779));
  jand g24547(.dina(n19523), .dinb(n5500), .dout(n24780));
  jand g24548(.dina(n19525), .dinb(n5424), .dout(n24781));
  jand g24549(.dina(n19527), .dinb(n5363), .dout(n24782));
  jor  g24550(.dina(n24782), .dinb(n24781), .dout(n24783));
  jor  g24551(.dina(n24783), .dinb(n24780), .dout(n24784));
  jor  g24552(.dina(n24784), .dinb(n24779), .dout(n24785));
  jxor g24553(.dina(n24785), .dinb(n72), .dout(n24786));
  jnot g24554(.din(n24786), .dout(n24787));
  jxor g24555(.dina(n24787), .dinb(n24778), .dout(n24788));
  jnot g24556(.din(n24627), .dout(n24789));
  jand g24557(.dina(n24789), .dinb(n24567), .dout(n24790));
  jnot g24558(.din(n24790), .dout(n24791));
  jand g24559(.dina(n24627), .dinb(n24568), .dout(n24792));
  jor  g24560(.dina(n24637), .dinb(n24792), .dout(n24793));
  jand g24561(.dina(n24793), .dinb(n24791), .dout(n24794));
  jxor g24562(.dina(n24794), .dinb(n24788), .dout(n24795));
  jand g24563(.dina(n21230), .dinb(n5693), .dout(n24796));
  jand g24564(.dina(n19517), .dinb(n6209), .dout(n24797));
  jand g24565(.dina(n19519), .dinb(n6131), .dout(n24798));
  jand g24566(.dina(n19521), .dinb(n5691), .dout(n24799));
  jor  g24567(.dina(n24799), .dinb(n24798), .dout(n24800));
  jor  g24568(.dina(n24800), .dinb(n24797), .dout(n24801));
  jor  g24569(.dina(n24801), .dinb(n24796), .dout(n24802));
  jxor g24570(.dina(n24802), .dinb(n4247), .dout(n24803));
  jnot g24571(.din(n24803), .dout(n24804));
  jxor g24572(.dina(n24804), .dinb(n24795), .dout(n24805));
  jnot g24573(.din(n24563), .dout(n24806));
  jnot g24574(.din(n24638), .dout(n24807));
  jand g24575(.dina(n24807), .dinb(n24806), .dout(n24808));
  jnot g24576(.din(n24808), .dout(n24809));
  jand g24577(.dina(n24638), .dinb(n24563), .dout(n24810));
  jor  g24578(.dina(n24648), .dinb(n24810), .dout(n24811));
  jand g24579(.dina(n24811), .dinb(n24809), .dout(n24812));
  jxor g24580(.dina(n24812), .dinb(n24805), .dout(n24813));
  jand g24581(.dina(n21762), .dinb(n6340), .dout(n24814));
  jand g24582(.dina(n19511), .dinb(n6798), .dout(n24815));
  jand g24583(.dina(n19513), .dinb(n6556), .dout(n24816));
  jand g24584(.dina(n19515), .dinb(n6338), .dout(n24817));
  jor  g24585(.dina(n24817), .dinb(n24816), .dout(n24818));
  jor  g24586(.dina(n24818), .dinb(n24815), .dout(n24819));
  jor  g24587(.dina(n24819), .dinb(n24814), .dout(n24820));
  jxor g24588(.dina(n24820), .dinb(n5064), .dout(n24821));
  jnot g24589(.din(n24821), .dout(n24822));
  jxor g24590(.dina(n24822), .dinb(n24813), .dout(n24823));
  jnot g24591(.din(n24649), .dout(n24824));
  jand g24592(.dina(n24824), .dinb(n24559), .dout(n24825));
  jnot g24593(.din(n24825), .dout(n24826));
  jand g24594(.dina(n24649), .dinb(n24560), .dout(n24827));
  jor  g24595(.dina(n24659), .dinb(n24827), .dout(n24828));
  jand g24596(.dina(n24828), .dinb(n24826), .dout(n24829));
  jxor g24597(.dina(n24829), .dinb(n24823), .dout(n24830));
  jand g24598(.dina(n22250), .dinb(n6936), .dout(n24831));
  jand g24599(.dina(n22248), .dinb(n7741), .dout(n24832));
  jand g24600(.dina(n19758), .dinb(n7613), .dout(n24833));
  jand g24601(.dina(n19510), .dinb(n6934), .dout(n24834));
  jor  g24602(.dina(n24834), .dinb(n24833), .dout(n24835));
  jor  g24603(.dina(n24835), .dinb(n24832), .dout(n24836));
  jor  g24604(.dina(n24836), .dinb(n24831), .dout(n24837));
  jxor g24605(.dina(n24837), .dinb(n5292), .dout(n24838));
  jnot g24606(.din(n24838), .dout(n24839));
  jxor g24607(.dina(n24839), .dinb(n24830), .dout(n24840));
  jnot g24608(.din(n24555), .dout(n24841));
  jnot g24609(.din(n24660), .dout(n24842));
  jand g24610(.dina(n24842), .dinb(n24841), .dout(n24843));
  jnot g24611(.din(n24843), .dout(n24844));
  jand g24612(.dina(n24660), .dinb(n24555), .dout(n24845));
  jor  g24613(.dina(n24670), .dinb(n24845), .dout(n24846));
  jand g24614(.dina(n24846), .dinb(n24844), .dout(n24847));
  jxor g24615(.dina(n24847), .dinb(n24840), .dout(n24848));
  jand g24616(.dina(n22605), .dinb(n7890), .dout(n24849));
  jand g24617(.dina(n22603), .dinb(n8441), .dout(n24850));
  jand g24618(.dina(n22539), .dinb(n8154), .dout(n24851));
  jand g24619(.dina(n22540), .dinb(n7888), .dout(n24852));
  jor  g24620(.dina(n24852), .dinb(n24851), .dout(n24853));
  jor  g24621(.dina(n24853), .dinb(n24850), .dout(n24854));
  jor  g24622(.dina(n24854), .dinb(n24849), .dout(n24855));
  jxor g24623(.dina(n24855), .dinb(n5833), .dout(n24856));
  jnot g24624(.din(n24856), .dout(n24857));
  jxor g24625(.dina(n24857), .dinb(n24848), .dout(n24858));
  jnot g24626(.din(n24671), .dout(n24859));
  jand g24627(.dina(n24859), .dinb(n24551), .dout(n24860));
  jnot g24628(.din(n24860), .dout(n24861));
  jand g24629(.dina(n24671), .dinb(n24552), .dout(n24862));
  jor  g24630(.dina(n24681), .dinb(n24862), .dout(n24863));
  jand g24631(.dina(n24863), .dinb(n24861), .dout(n24864));
  jxor g24632(.dina(n24864), .dinb(n24858), .dout(n24865));
  jor  g24633(.dina(n23708), .dinb(n8772), .dout(n24866));
  jor  g24634(.dina(n23710), .dinb(n9490), .dout(n24867));
  jor  g24635(.dina(n23496), .dinb(n9127), .dout(n24868));
  jor  g24636(.dina(n23450), .dinb(n8770), .dout(n24869));
  jand g24637(.dina(n24869), .dinb(n24868), .dout(n24870));
  jand g24638(.dina(n24870), .dinb(n24867), .dout(n24871));
  jand g24639(.dina(n24871), .dinb(n24866), .dout(n24872));
  jxor g24640(.dina(n24872), .dinb(\a[8] ), .dout(n24873));
  jnot g24641(.din(n24873), .dout(n24874));
  jxor g24642(.dina(n24874), .dinb(n24865), .dout(n24875));
  jnot g24643(.din(n24547), .dout(n24876));
  jnot g24644(.din(n24682), .dout(n24877));
  jand g24645(.dina(n24877), .dinb(n24876), .dout(n24878));
  jnot g24646(.din(n24878), .dout(n24879));
  jand g24647(.dina(n24682), .dinb(n24547), .dout(n24880));
  jor  g24648(.dina(n24692), .dinb(n24880), .dout(n24881));
  jand g24649(.dina(n24881), .dinb(n24879), .dout(n24882));
  jxor g24650(.dina(n24882), .dinb(n24875), .dout(n24883));
  jor  g24651(.dina(n24337), .dinb(n9919), .dout(n24884));
  jor  g24652(.dina(n24335), .dinb(n10826), .dout(n24885));
  jor  g24653(.dina(n24142), .dinb(n10351), .dout(n24886));
  jor  g24654(.dina(n23921), .dinb(n9918), .dout(n24887));
  jand g24655(.dina(n24887), .dinb(n24886), .dout(n24888));
  jand g24656(.dina(n24888), .dinb(n24885), .dout(n24889));
  jand g24657(.dina(n24889), .dinb(n24884), .dout(n24890));
  jxor g24658(.dina(n24890), .dinb(\a[5] ), .dout(n24891));
  jnot g24659(.din(n24891), .dout(n24892));
  jxor g24660(.dina(n24892), .dinb(n24883), .dout(n24893));
  jnot g24661(.din(n24693), .dout(n24894));
  jand g24662(.dina(n24894), .dinb(n24544), .dout(n24895));
  jnot g24663(.din(n24895), .dout(n24896));
  jnot g24664(.din(n24544), .dout(n24897));
  jand g24665(.dina(n24693), .dinb(n24897), .dout(n24898));
  jnot g24666(.din(n24702), .dout(n24899));
  jor  g24667(.dina(n24899), .dinb(n24898), .dout(n24900));
  jand g24668(.dina(n24900), .dinb(n24896), .dout(n24901));
  jxor g24669(.dina(n24901), .dinb(n24893), .dout(n24902));
  jand g24670(.dina(n24703), .dinb(n24540), .dout(n24903));
  jand g24671(.dina(n24707), .dinb(n24704), .dout(n24904));
  jor  g24672(.dina(n24904), .dinb(n24903), .dout(n24905));
  jxor g24673(.dina(n24905), .dinb(n24902), .dout(n24906));
  jxor g24674(.dina(n24906), .dinb(n24710), .dout(\result[8] ));
  jand g24675(.dina(n24906), .dinb(n24710), .dout(n24908));
  jor  g24676(.dina(n24357), .dinb(n9919), .dout(n24909));
  jor  g24677(.dina(n24335), .dinb(n17273), .dout(n24910));
  jor  g24678(.dina(n24142), .dinb(n9918), .dout(n24911));
  jand g24679(.dina(n24911), .dinb(n24910), .dout(n24912));
  jand g24680(.dina(n24912), .dinb(n24909), .dout(n24913));
  jxor g24681(.dina(n24913), .dinb(\a[5] ), .dout(n24914));
  jnot g24682(.din(n24914), .dout(n24915));
  jnot g24683(.din(n24858), .dout(n24916));
  jnot g24684(.din(n24864), .dout(n24917));
  jand g24685(.dina(n24917), .dinb(n24916), .dout(n24918));
  jnot g24686(.din(n24918), .dout(n24919));
  jand g24687(.dina(n24864), .dinb(n24858), .dout(n24920));
  jor  g24688(.dina(n24874), .dinb(n24920), .dout(n24921));
  jand g24689(.dina(n24921), .dinb(n24919), .dout(n24922));
  jxor g24690(.dina(n24922), .dinb(n24915), .dout(n24923));
  jor  g24691(.dina(n24771), .dinb(n24763), .dout(n24924));
  jand g24692(.dina(n24772), .dinb(n24719), .dout(n24925));
  jnot g24693(.din(n24925), .dout(n24926));
  jand g24694(.dina(n24926), .dinb(n24924), .dout(n24927));
  jnot g24695(.din(n24927), .dout(n24928));
  jand g24696(.dina(n20793), .dinb(n75), .dout(n24929));
  jand g24697(.dina(n19527), .dinb(n4933), .dout(n24930));
  jand g24698(.dina(n19529), .dinb(n4918), .dout(n24931));
  jand g24699(.dina(n19531), .dinb(n4745), .dout(n24932));
  jor  g24700(.dina(n24932), .dinb(n24931), .dout(n24933));
  jor  g24701(.dina(n24933), .dinb(n24930), .dout(n24934));
  jor  g24702(.dina(n24934), .dinb(n24929), .dout(n24935));
  jxor g24703(.dina(n24935), .dinb(n68), .dout(n24936));
  jnot g24704(.din(n24936), .dout(n24937));
  jand g24705(.dina(n24760), .dinb(n24753), .dout(n24938));
  jand g24706(.dina(n24761), .dinb(n24724), .dout(n24939));
  jor  g24707(.dina(n24939), .dinb(n24938), .dout(n24940));
  jor  g24708(.dina(n24744), .dinb(n24596), .dout(n24941));
  jand g24709(.dina(n24752), .dinb(n24745), .dout(n24942));
  jnot g24710(.din(n24942), .dout(n24943));
  jand g24711(.dina(n24943), .dinb(n24941), .dout(n24944));
  jnot g24712(.din(n24944), .dout(n24945));
  jand g24713(.dina(n3644), .dinb(n5989), .dout(n24946));
  jand g24714(.dina(n798), .dinb(n771), .dout(n24947));
  jand g24715(.dina(n24947), .dinb(n24946), .dout(n24948));
  jand g24716(.dina(n24948), .dinb(n13834), .dout(n24949));
  jand g24717(.dina(n24949), .dinb(n3914), .dout(n24950));
  jand g24718(.dina(n926), .dinb(n533), .dout(n24951));
  jand g24719(.dina(n24951), .dinb(n678), .dout(n24952));
  jand g24720(.dina(n719), .dinb(n238), .dout(n24953));
  jand g24721(.dina(n24953), .dinb(n1959), .dout(n24954));
  jand g24722(.dina(n24954), .dinb(n24952), .dout(n24955));
  jand g24723(.dina(n24955), .dinb(n3261), .dout(n24956));
  jand g24724(.dina(n24956), .dinb(n1555), .dout(n24957));
  jand g24725(.dina(n24957), .dinb(n5944), .dout(n24958));
  jand g24726(.dina(n24958), .dinb(n24950), .dout(n24959));
  jand g24727(.dina(n24959), .dinb(n2969), .dout(n24960));
  jand g24728(.dina(n24960), .dinb(n1674), .dout(n24961));
  jxor g24729(.dina(n24961), .dinb(n24596), .dout(n24962));
  jxor g24730(.dina(n24962), .dinb(n24945), .dout(n24963));
  jand g24731(.dina(n20131), .dinb(n732), .dout(n24964));
  jand g24732(.dina(n19539), .dinb(n3855), .dout(n24965));
  jand g24733(.dina(n19541), .dinb(n3858), .dout(n24966));
  jand g24734(.dina(n19543), .dinb(n3851), .dout(n24967));
  jor  g24735(.dina(n24967), .dinb(n24966), .dout(n24968));
  jor  g24736(.dina(n24968), .dinb(n24965), .dout(n24969));
  jor  g24737(.dina(n24969), .dinb(n24964), .dout(n24970));
  jxor g24738(.dina(n24970), .dinb(n24963), .dout(n24971));
  jxor g24739(.dina(n24971), .dinb(n24940), .dout(n24972));
  jnot g24740(.din(n24972), .dout(n24973));
  jand g24741(.dina(n20399), .dinb(n4449), .dout(n24974));
  jand g24742(.dina(n19533), .dinb(n4453), .dout(n24975));
  jand g24743(.dina(n19535), .dinb(n4457), .dout(n24976));
  jand g24744(.dina(n19537), .dinb(n4461), .dout(n24977));
  jor  g24745(.dina(n24977), .dinb(n24976), .dout(n24978));
  jor  g24746(.dina(n24978), .dinb(n24975), .dout(n24979));
  jor  g24747(.dina(n24979), .dinb(n24974), .dout(n24980));
  jxor g24748(.dina(n24980), .dinb(n88), .dout(n24981));
  jxor g24749(.dina(n24981), .dinb(n24973), .dout(n24982));
  jxor g24750(.dina(n24982), .dinb(n24937), .dout(n24983));
  jxor g24751(.dina(n24983), .dinb(n24928), .dout(n24984));
  jand g24752(.dina(n21086), .dinb(n5365), .dout(n24985));
  jand g24753(.dina(n19521), .dinb(n5500), .dout(n24986));
  jand g24754(.dina(n19523), .dinb(n5424), .dout(n24987));
  jand g24755(.dina(n19525), .dinb(n5363), .dout(n24988));
  jor  g24756(.dina(n24988), .dinb(n24987), .dout(n24989));
  jor  g24757(.dina(n24989), .dinb(n24986), .dout(n24990));
  jor  g24758(.dina(n24990), .dinb(n24985), .dout(n24991));
  jxor g24759(.dina(n24991), .dinb(n72), .dout(n24992));
  jnot g24760(.din(n24992), .dout(n24993));
  jxor g24761(.dina(n24993), .dinb(n24984), .dout(n24994));
  jnot g24762(.din(n24773), .dout(n24995));
  jnot g24763(.din(n24777), .dout(n24996));
  jand g24764(.dina(n24996), .dinb(n24995), .dout(n24997));
  jnot g24765(.din(n24997), .dout(n24998));
  jand g24766(.dina(n24777), .dinb(n24773), .dout(n24999));
  jor  g24767(.dina(n24787), .dinb(n24999), .dout(n25000));
  jand g24768(.dina(n25000), .dinb(n24998), .dout(n25001));
  jxor g24769(.dina(n25001), .dinb(n24994), .dout(n25002));
  jand g24770(.dina(n21218), .dinb(n5693), .dout(n25003));
  jand g24771(.dina(n19515), .dinb(n6209), .dout(n25004));
  jand g24772(.dina(n19517), .dinb(n6131), .dout(n25005));
  jand g24773(.dina(n19519), .dinb(n5691), .dout(n25006));
  jor  g24774(.dina(n25006), .dinb(n25005), .dout(n25007));
  jor  g24775(.dina(n25007), .dinb(n25004), .dout(n25008));
  jor  g24776(.dina(n25008), .dinb(n25003), .dout(n25009));
  jxor g24777(.dina(n25009), .dinb(n4247), .dout(n25010));
  jnot g24778(.din(n25010), .dout(n25011));
  jxor g24779(.dina(n25011), .dinb(n25002), .dout(n25012));
  jnot g24780(.din(n24788), .dout(n25013));
  jnot g24781(.din(n24794), .dout(n25014));
  jand g24782(.dina(n25014), .dinb(n25013), .dout(n25015));
  jnot g24783(.din(n25015), .dout(n25016));
  jand g24784(.dina(n24794), .dinb(n24788), .dout(n25017));
  jor  g24785(.dina(n24804), .dinb(n25017), .dout(n25018));
  jand g24786(.dina(n25018), .dinb(n25016), .dout(n25019));
  jxor g24787(.dina(n25019), .dinb(n25012), .dout(n25020));
  jand g24788(.dina(n21750), .dinb(n6340), .dout(n25021));
  jand g24789(.dina(n19510), .dinb(n6798), .dout(n25022));
  jand g24790(.dina(n19511), .dinb(n6556), .dout(n25023));
  jand g24791(.dina(n19513), .dinb(n6338), .dout(n25024));
  jor  g24792(.dina(n25024), .dinb(n25023), .dout(n25025));
  jor  g24793(.dina(n25025), .dinb(n25022), .dout(n25026));
  jor  g24794(.dina(n25026), .dinb(n25021), .dout(n25027));
  jxor g24795(.dina(n25027), .dinb(n5064), .dout(n25028));
  jnot g24796(.din(n25028), .dout(n25029));
  jxor g24797(.dina(n25029), .dinb(n25020), .dout(n25030));
  jnot g24798(.din(n24805), .dout(n25031));
  jnot g24799(.din(n24812), .dout(n25032));
  jand g24800(.dina(n25032), .dinb(n25031), .dout(n25033));
  jnot g24801(.din(n25033), .dout(n25034));
  jand g24802(.dina(n24812), .dinb(n24805), .dout(n25035));
  jor  g24803(.dina(n24822), .dinb(n25035), .dout(n25036));
  jand g24804(.dina(n25036), .dinb(n25034), .dout(n25037));
  jxor g24805(.dina(n25037), .dinb(n25030), .dout(n25038));
  jand g24806(.dina(n22627), .dinb(n6936), .dout(n25039));
  jand g24807(.dina(n22540), .dinb(n7741), .dout(n25040));
  jand g24808(.dina(n22248), .dinb(n7613), .dout(n25041));
  jand g24809(.dina(n19758), .dinb(n6934), .dout(n25042));
  jor  g24810(.dina(n25042), .dinb(n25041), .dout(n25043));
  jor  g24811(.dina(n25043), .dinb(n25040), .dout(n25044));
  jor  g24812(.dina(n25044), .dinb(n25039), .dout(n25045));
  jxor g24813(.dina(n25045), .dinb(n5292), .dout(n25046));
  jnot g24814(.din(n25046), .dout(n25047));
  jxor g24815(.dina(n25047), .dinb(n25038), .dout(n25048));
  jnot g24816(.din(n24823), .dout(n25049));
  jnot g24817(.din(n24829), .dout(n25050));
  jand g24818(.dina(n25050), .dinb(n25049), .dout(n25051));
  jnot g24819(.din(n25051), .dout(n25052));
  jand g24820(.dina(n24829), .dinb(n24823), .dout(n25053));
  jor  g24821(.dina(n24839), .dinb(n25053), .dout(n25054));
  jand g24822(.dina(n25054), .dinb(n25052), .dout(n25055));
  jxor g24823(.dina(n25055), .dinb(n25048), .dout(n25056));
  jand g24824(.dina(n23262), .dinb(n7890), .dout(n25057));
  jand g24825(.dina(n23260), .dinb(n8441), .dout(n25058));
  jand g24826(.dina(n22603), .dinb(n8154), .dout(n25059));
  jand g24827(.dina(n22539), .dinb(n7888), .dout(n25060));
  jor  g24828(.dina(n25060), .dinb(n25059), .dout(n25061));
  jor  g24829(.dina(n25061), .dinb(n25058), .dout(n25062));
  jor  g24830(.dina(n25062), .dinb(n25057), .dout(n25063));
  jxor g24831(.dina(n25063), .dinb(n5833), .dout(n25064));
  jnot g24832(.din(n25064), .dout(n25065));
  jxor g24833(.dina(n25065), .dinb(n25056), .dout(n25066));
  jnot g24834(.din(n24840), .dout(n25067));
  jnot g24835(.din(n24847), .dout(n25068));
  jand g24836(.dina(n25068), .dinb(n25067), .dout(n25069));
  jnot g24837(.din(n25069), .dout(n25070));
  jand g24838(.dina(n24847), .dinb(n24840), .dout(n25071));
  jor  g24839(.dina(n24857), .dinb(n25071), .dout(n25072));
  jand g24840(.dina(n25072), .dinb(n25070), .dout(n25073));
  jxor g24841(.dina(n25073), .dinb(n25066), .dout(n25074));
  jor  g24842(.dina(n23919), .dinb(n8772), .dout(n25075));
  jor  g24843(.dina(n23921), .dinb(n9490), .dout(n25076));
  jor  g24844(.dina(n23710), .dinb(n9127), .dout(n25077));
  jor  g24845(.dina(n23496), .dinb(n8770), .dout(n25078));
  jand g24846(.dina(n25078), .dinb(n25077), .dout(n25079));
  jand g24847(.dina(n25079), .dinb(n25076), .dout(n25080));
  jand g24848(.dina(n25080), .dinb(n25075), .dout(n25081));
  jxor g24849(.dina(n25081), .dinb(\a[8] ), .dout(n25082));
  jnot g24850(.din(n25082), .dout(n25083));
  jxor g24851(.dina(n25083), .dinb(n25074), .dout(n25084));
  jxor g24852(.dina(n25084), .dinb(n24923), .dout(n25085));
  jnot g24853(.din(n24875), .dout(n25086));
  jnot g24854(.din(n24882), .dout(n25087));
  jand g24855(.dina(n25087), .dinb(n25086), .dout(n25088));
  jnot g24856(.din(n25088), .dout(n25089));
  jand g24857(.dina(n24882), .dinb(n24875), .dout(n25090));
  jor  g24858(.dina(n24892), .dinb(n25090), .dout(n25091));
  jand g24859(.dina(n25091), .dinb(n25089), .dout(n25092));
  jxor g24860(.dina(n25092), .dinb(n25085), .dout(n25093));
  jand g24861(.dina(n24901), .dinb(n24893), .dout(n25094));
  jand g24862(.dina(n24905), .dinb(n24902), .dout(n25095));
  jor  g24863(.dina(n25095), .dinb(n25094), .dout(n25096));
  jxor g24864(.dina(n25096), .dinb(n25093), .dout(n25097));
  jxor g24865(.dina(n25097), .dinb(n24908), .dout(\result[9] ));
  jand g24866(.dina(n25097), .dinb(n24908), .dout(n25099));
  jand g24867(.dina(n25092), .dinb(n25085), .dout(n25100));
  jand g24868(.dina(n25096), .dinb(n25093), .dout(n25101));
  jor  g24869(.dina(n25101), .dinb(n25100), .dout(n25102));
  jor  g24870(.dina(n24981), .dinb(n24973), .dout(n25103));
  jand g24871(.dina(n24982), .dinb(n24937), .dout(n25104));
  jnot g24872(.din(n25104), .dout(n25105));
  jand g24873(.dina(n25105), .dinb(n25103), .dout(n25106));
  jnot g24874(.din(n25106), .dout(n25107));
  jand g24875(.dina(n20781), .dinb(n75), .dout(n25108));
  jand g24876(.dina(n19525), .dinb(n4933), .dout(n25109));
  jand g24877(.dina(n19527), .dinb(n4918), .dout(n25110));
  jand g24878(.dina(n19529), .dinb(n4745), .dout(n25111));
  jor  g24879(.dina(n25111), .dinb(n25110), .dout(n25112));
  jor  g24880(.dina(n25112), .dinb(n25109), .dout(n25113));
  jor  g24881(.dina(n25113), .dinb(n25108), .dout(n25114));
  jxor g24882(.dina(n25114), .dinb(n68), .dout(n25115));
  jnot g24883(.din(n25115), .dout(n25116));
  jand g24884(.dina(n24970), .dinb(n24963), .dout(n25117));
  jand g24885(.dina(n24971), .dinb(n24940), .dout(n25118));
  jor  g24886(.dina(n25118), .dinb(n25117), .dout(n25119));
  jor  g24887(.dina(n24961), .dinb(n24596), .dout(n25120));
  jand g24888(.dina(n24962), .dinb(n24945), .dout(n25121));
  jnot g24889(.din(n25121), .dout(n25122));
  jand g24890(.dina(n25122), .dinb(n25120), .dout(n25123));
  jnot g24891(.din(n25123), .dout(n25124));
  jand g24892(.dina(n778), .dinb(n449), .dout(n25125));
  jand g24893(.dina(n25125), .dinb(n4231), .dout(n25126));
  jand g24894(.dina(n5211), .dinb(n4287), .dout(n25127));
  jand g24895(.dina(n25127), .dinb(n25126), .dout(n25128));
  jand g24896(.dina(n696), .dinb(n103), .dout(n25129));
  jand g24897(.dina(n25129), .dinb(n614), .dout(n25130));
  jand g24898(.dina(n25130), .dinb(n12285), .dout(n25131));
  jand g24899(.dina(n25131), .dinb(n25128), .dout(n25132));
  jand g24900(.dina(n1930), .dinb(n939), .dout(n25133));
  jand g24901(.dina(n25133), .dinb(n2026), .dout(n25134));
  jand g24902(.dina(n25134), .dinb(n12269), .dout(n25135));
  jand g24903(.dina(n25135), .dinb(n25132), .dout(n25136));
  jand g24904(.dina(n25136), .dinb(n20709), .dout(n25137));
  jand g24905(.dina(n25137), .dinb(n4092), .dout(n25138));
  jand g24906(.dina(n25138), .dinb(n2638), .dout(n25139));
  jxor g24907(.dina(n25139), .dinb(n24749), .dout(n25140));
  jand g24908(.dina(n24593), .dinb(n13656), .dout(n25141));
  jxor g24909(.dina(n25141), .dinb(n64), .dout(n25142));
  jxor g24910(.dina(n25142), .dinb(n25140), .dout(n25143));
  jxor g24911(.dina(n25143), .dinb(n25124), .dout(n25144));
  jand g24912(.dina(n20387), .dinb(n732), .dout(n25145));
  jand g24913(.dina(n19537), .dinb(n3855), .dout(n25146));
  jand g24914(.dina(n19539), .dinb(n3858), .dout(n25147));
  jand g24915(.dina(n19541), .dinb(n3851), .dout(n25148));
  jor  g24916(.dina(n25148), .dinb(n25147), .dout(n25149));
  jor  g24917(.dina(n25149), .dinb(n25146), .dout(n25150));
  jor  g24918(.dina(n25150), .dinb(n25145), .dout(n25151));
  jxor g24919(.dina(n25151), .dinb(n25144), .dout(n25152));
  jxor g24920(.dina(n25152), .dinb(n25119), .dout(n25153));
  jand g24921(.dina(n19780), .dinb(n4449), .dout(n25154));
  jand g24922(.dina(n19531), .dinb(n4453), .dout(n25155));
  jand g24923(.dina(n19533), .dinb(n4457), .dout(n25156));
  jand g24924(.dina(n19535), .dinb(n4461), .dout(n25157));
  jor  g24925(.dina(n25157), .dinb(n25156), .dout(n25158));
  jor  g24926(.dina(n25158), .dinb(n25155), .dout(n25159));
  jor  g24927(.dina(n25159), .dinb(n25154), .dout(n25160));
  jxor g24928(.dina(n25160), .dinb(n88), .dout(n25161));
  jnot g24929(.din(n25161), .dout(n25162));
  jxor g24930(.dina(n25162), .dinb(n25153), .dout(n25163));
  jxor g24931(.dina(n25163), .dinb(n25116), .dout(n25164));
  jxor g24932(.dina(n25164), .dinb(n25107), .dout(n25165));
  jnot g24933(.din(n25165), .dout(n25166));
  jand g24934(.dina(n21240), .dinb(n5365), .dout(n25167));
  jand g24935(.dina(n19519), .dinb(n5500), .dout(n25168));
  jand g24936(.dina(n19521), .dinb(n5424), .dout(n25169));
  jand g24937(.dina(n19523), .dinb(n5363), .dout(n25170));
  jor  g24938(.dina(n25170), .dinb(n25169), .dout(n25171));
  jor  g24939(.dina(n25171), .dinb(n25168), .dout(n25172));
  jor  g24940(.dina(n25172), .dinb(n25167), .dout(n25173));
  jxor g24941(.dina(n25173), .dinb(n72), .dout(n25174));
  jxor g24942(.dina(n25174), .dinb(n25166), .dout(n25175));
  jnot g24943(.din(n24983), .dout(n25176));
  jand g24944(.dina(n25176), .dinb(n24927), .dout(n25177));
  jnot g24945(.din(n25177), .dout(n25178));
  jand g24946(.dina(n24983), .dinb(n24928), .dout(n25179));
  jor  g24947(.dina(n24993), .dinb(n25179), .dout(n25180));
  jand g24948(.dina(n25180), .dinb(n25178), .dout(n25181));
  jxor g24949(.dina(n25181), .dinb(n25175), .dout(n25182));
  jand g24950(.dina(n21738), .dinb(n5693), .dout(n25183));
  jand g24951(.dina(n19513), .dinb(n6209), .dout(n25184));
  jand g24952(.dina(n19515), .dinb(n6131), .dout(n25185));
  jand g24953(.dina(n19517), .dinb(n5691), .dout(n25186));
  jor  g24954(.dina(n25186), .dinb(n25185), .dout(n25187));
  jor  g24955(.dina(n25187), .dinb(n25184), .dout(n25188));
  jor  g24956(.dina(n25188), .dinb(n25183), .dout(n25189));
  jxor g24957(.dina(n25189), .dinb(n4247), .dout(n25190));
  jxor g24958(.dina(n25190), .dinb(n25182), .dout(n25191));
  jnot g24959(.din(n24994), .dout(n25192));
  jnot g24960(.din(n25001), .dout(n25193));
  jand g24961(.dina(n25193), .dinb(n25192), .dout(n25194));
  jnot g24962(.din(n25194), .dout(n25195));
  jand g24963(.dina(n25001), .dinb(n24994), .dout(n25196));
  jor  g24964(.dina(n25011), .dinb(n25196), .dout(n25197));
  jand g24965(.dina(n25197), .dinb(n25195), .dout(n25198));
  jnot g24966(.din(n25198), .dout(n25199));
  jxor g24967(.dina(n25199), .dinb(n25191), .dout(n25200));
  jand g24968(.dina(n19760), .dinb(n6340), .dout(n25201));
  jand g24969(.dina(n19758), .dinb(n6798), .dout(n25202));
  jand g24970(.dina(n19510), .dinb(n6556), .dout(n25203));
  jand g24971(.dina(n19511), .dinb(n6338), .dout(n25204));
  jor  g24972(.dina(n25204), .dinb(n25203), .dout(n25205));
  jor  g24973(.dina(n25205), .dinb(n25202), .dout(n25206));
  jor  g24974(.dina(n25206), .dinb(n25201), .dout(n25207));
  jxor g24975(.dina(n25207), .dinb(n5064), .dout(n25208));
  jxor g24976(.dina(n25208), .dinb(n25200), .dout(n25209));
  jnot g24977(.din(n25012), .dout(n25210));
  jnot g24978(.din(n25019), .dout(n25211));
  jand g24979(.dina(n25211), .dinb(n25210), .dout(n25212));
  jnot g24980(.din(n25212), .dout(n25213));
  jand g24981(.dina(n25019), .dinb(n25012), .dout(n25214));
  jor  g24982(.dina(n25029), .dinb(n25214), .dout(n25215));
  jand g24983(.dina(n25215), .dinb(n25213), .dout(n25216));
  jnot g24984(.din(n25216), .dout(n25217));
  jxor g24985(.dina(n25217), .dinb(n25209), .dout(n25218));
  jand g24986(.dina(n22617), .dinb(n6936), .dout(n25219));
  jand g24987(.dina(n22539), .dinb(n7741), .dout(n25220));
  jand g24988(.dina(n22540), .dinb(n7613), .dout(n25221));
  jand g24989(.dina(n22248), .dinb(n6934), .dout(n25222));
  jor  g24990(.dina(n25222), .dinb(n25221), .dout(n25223));
  jor  g24991(.dina(n25223), .dinb(n25220), .dout(n25224));
  jor  g24992(.dina(n25224), .dinb(n25219), .dout(n25225));
  jxor g24993(.dina(n25225), .dinb(n5292), .dout(n25226));
  jnot g24994(.din(n25226), .dout(n25227));
  jnot g24995(.din(n25030), .dout(n25228));
  jnot g24996(.din(n25037), .dout(n25229));
  jand g24997(.dina(n25229), .dinb(n25228), .dout(n25230));
  jnot g24998(.din(n25230), .dout(n25231));
  jand g24999(.dina(n25037), .dinb(n25030), .dout(n25232));
  jor  g25000(.dina(n25047), .dinb(n25232), .dout(n25233));
  jand g25001(.dina(n25233), .dinb(n25231), .dout(n25234));
  jxor g25002(.dina(n25234), .dinb(n25227), .dout(n25235));
  jxor g25003(.dina(n25235), .dinb(n25218), .dout(n25236));
  jnot g25004(.din(n25236), .dout(n25237));
  jor  g25005(.dina(n23494), .dinb(n7891), .dout(n25238));
  jor  g25006(.dina(n23496), .dinb(n8440), .dout(n25239));
  jor  g25007(.dina(n23450), .dinb(n8155), .dout(n25240));
  jor  g25008(.dina(n23449), .dinb(n7889), .dout(n25241));
  jand g25009(.dina(n25241), .dinb(n25240), .dout(n25242));
  jand g25010(.dina(n25242), .dinb(n25239), .dout(n25243));
  jand g25011(.dina(n25243), .dinb(n25238), .dout(n25244));
  jxor g25012(.dina(n25244), .dinb(\a[11] ), .dout(n25245));
  jxor g25013(.dina(n25245), .dinb(n25237), .dout(n25246));
  jnot g25014(.din(n25048), .dout(n25247));
  jnot g25015(.din(n25055), .dout(n25248));
  jand g25016(.dina(n25248), .dinb(n25247), .dout(n25249));
  jnot g25017(.din(n25249), .dout(n25250));
  jand g25018(.dina(n25055), .dinb(n25048), .dout(n25251));
  jor  g25019(.dina(n25065), .dinb(n25251), .dout(n25252));
  jand g25020(.dina(n25252), .dinb(n25250), .dout(n25253));
  jxor g25021(.dina(n25253), .dinb(n25246), .dout(n25254));
  jor  g25022(.dina(n24140), .dinb(n8772), .dout(n25255));
  jor  g25023(.dina(n24142), .dinb(n9490), .dout(n25256));
  jor  g25024(.dina(n23921), .dinb(n9127), .dout(n25257));
  jor  g25025(.dina(n23710), .dinb(n8770), .dout(n25258));
  jand g25026(.dina(n25258), .dinb(n25257), .dout(n25259));
  jand g25027(.dina(n25259), .dinb(n25256), .dout(n25260));
  jand g25028(.dina(n25260), .dinb(n25255), .dout(n25261));
  jxor g25029(.dina(n25261), .dinb(\a[8] ), .dout(n25262));
  jnot g25030(.din(n25262), .dout(n25263));
  jnot g25031(.din(n25066), .dout(n25264));
  jnot g25032(.din(n25073), .dout(n25265));
  jand g25033(.dina(n25265), .dinb(n25264), .dout(n25266));
  jnot g25034(.din(n25266), .dout(n25267));
  jand g25035(.dina(n25073), .dinb(n25066), .dout(n25268));
  jor  g25036(.dina(n25083), .dinb(n25268), .dout(n25269));
  jand g25037(.dina(n25269), .dinb(n25267), .dout(n25270));
  jxor g25038(.dina(n25270), .dinb(n25263), .dout(n25271));
  jxor g25039(.dina(n25271), .dinb(n25254), .dout(n25272));
  jor  g25040(.dina(n24922), .dinb(n24915), .dout(n25273));
  jand g25041(.dina(n24922), .dinb(n24915), .dout(n25274));
  jor  g25042(.dina(n25084), .dinb(n25274), .dout(n25275));
  jand g25043(.dina(n25275), .dinb(n25273), .dout(n25276));
  jxor g25044(.dina(n25276), .dinb(n25272), .dout(n25277));
  jxor g25045(.dina(n25277), .dinb(n25102), .dout(n25278));
  jxor g25046(.dina(n25278), .dinb(n25099), .dout(\result[10] ));
  jand g25047(.dina(n25278), .dinb(n25099), .dout(n25280));
  jand g25048(.dina(n25276), .dinb(n25272), .dout(n25281));
  jand g25049(.dina(n25277), .dinb(n25102), .dout(n25282));
  jor  g25050(.dina(n25282), .dinb(n25281), .dout(n25283));
  jand g25051(.dina(n25270), .dinb(n25263), .dout(n25284));
  jand g25052(.dina(n25271), .dinb(n25254), .dout(n25285));
  jor  g25053(.dina(n25285), .dinb(n25284), .dout(n25286));
  jor  g25054(.dina(n25245), .dinb(n25237), .dout(n25287));
  jand g25055(.dina(n25253), .dinb(n25246), .dout(n25288));
  jnot g25056(.din(n25288), .dout(n25289));
  jand g25057(.dina(n25289), .dinb(n25287), .dout(n25290));
  jor  g25058(.dina(n23708), .dinb(n7891), .dout(n25291));
  jor  g25059(.dina(n23710), .dinb(n8440), .dout(n25292));
  jor  g25060(.dina(n23496), .dinb(n8155), .dout(n25293));
  jor  g25061(.dina(n23450), .dinb(n7889), .dout(n25294));
  jand g25062(.dina(n25294), .dinb(n25293), .dout(n25295));
  jand g25063(.dina(n25295), .dinb(n25292), .dout(n25296));
  jand g25064(.dina(n25296), .dinb(n25291), .dout(n25297));
  jxor g25065(.dina(n25297), .dinb(\a[11] ), .dout(n25298));
  jnot g25066(.din(n25298), .dout(n25299));
  jand g25067(.dina(n25234), .dinb(n25227), .dout(n25300));
  jand g25068(.dina(n25235), .dinb(n25218), .dout(n25301));
  jor  g25069(.dina(n25301), .dinb(n25300), .dout(n25302));
  jnot g25070(.din(n25200), .dout(n25303));
  jor  g25071(.dina(n25208), .dinb(n25303), .dout(n25304));
  jor  g25072(.dina(n25217), .dinb(n25209), .dout(n25305));
  jand g25073(.dina(n25305), .dinb(n25304), .dout(n25306));
  jnot g25074(.din(n25182), .dout(n25307));
  jor  g25075(.dina(n25190), .dinb(n25307), .dout(n25308));
  jor  g25076(.dina(n25199), .dinb(n25191), .dout(n25309));
  jand g25077(.dina(n25309), .dinb(n25308), .dout(n25310));
  jor  g25078(.dina(n25174), .dinb(n25166), .dout(n25311));
  jand g25079(.dina(n25181), .dinb(n25175), .dout(n25312));
  jnot g25080(.din(n25312), .dout(n25313));
  jand g25081(.dina(n25313), .dinb(n25311), .dout(n25314));
  jand g25082(.dina(n25163), .dinb(n25116), .dout(n25315));
  jand g25083(.dina(n25164), .dinb(n25107), .dout(n25316));
  jor  g25084(.dina(n25316), .dinb(n25315), .dout(n25317));
  jand g25085(.dina(n25143), .dinb(n25124), .dout(n25318));
  jand g25086(.dina(n25151), .dinb(n25144), .dout(n25319));
  jor  g25087(.dina(n25319), .dinb(n25318), .dout(n25320));
  jor  g25088(.dina(n25139), .dinb(n24749), .dout(n25321));
  jand g25089(.dina(n25142), .dinb(n25140), .dout(n25322));
  jnot g25090(.din(n25322), .dout(n25323));
  jand g25091(.dina(n25323), .dinb(n25321), .dout(n25324));
  jand g25092(.dina(n858), .dinb(n807), .dout(n25325));
  jand g25093(.dina(n25325), .dinb(n2179), .dout(n25326));
  jand g25094(.dina(n25326), .dinb(n7430), .dout(n25327));
  jand g25095(.dina(n25327), .dinb(n6632), .dout(n25328));
  jand g25096(.dina(n13173), .dinb(n1846), .dout(n25329));
  jand g25097(.dina(n2222), .dinb(n1585), .dout(n25330));
  jand g25098(.dina(n25330), .dinb(n25329), .dout(n25331));
  jand g25099(.dina(n25331), .dinb(n2117), .dout(n25332));
  jand g25100(.dina(n25332), .dinb(n1159), .dout(n25333));
  jand g25101(.dina(n25333), .dinb(n25328), .dout(n25334));
  jand g25102(.dina(n2834), .dinb(n2560), .dout(n25335));
  jand g25103(.dina(n1299), .dinb(n1274), .dout(n25336));
  jand g25104(.dina(n25336), .dinb(n25335), .dout(n25337));
  jand g25105(.dina(n25337), .dinb(n1596), .dout(n25338));
  jand g25106(.dina(n25338), .dinb(n7352), .dout(n25339));
  jand g25107(.dina(n926), .dinb(n424), .dout(n25340));
  jand g25108(.dina(n25340), .dinb(n1278), .dout(n25341));
  jand g25109(.dina(n4163), .dinb(n263), .dout(n25342));
  jand g25110(.dina(n25342), .dinb(n25341), .dout(n25343));
  jand g25111(.dina(n375), .dinb(n108), .dout(n25344));
  jand g25112(.dina(n1221), .dinb(n357), .dout(n25345));
  jand g25113(.dina(n25345), .dinb(n25344), .dout(n25346));
  jand g25114(.dina(n25346), .dinb(n3628), .dout(n25347));
  jand g25115(.dina(n25347), .dinb(n25343), .dout(n25348));
  jand g25116(.dina(n25348), .dinb(n2326), .dout(n25349));
  jand g25117(.dina(n25349), .dinb(n25339), .dout(n25350));
  jand g25118(.dina(n25350), .dinb(n25334), .dout(n25351));
  jand g25119(.dina(n25351), .dinb(n1481), .dout(n25352));
  jnot g25120(.din(n25352), .dout(n25353));
  jxor g25121(.dina(n25353), .dinb(n25324), .dout(n25354));
  jand g25122(.dina(n20413), .dinb(n732), .dout(n25355));
  jand g25123(.dina(n19535), .dinb(n3855), .dout(n25356));
  jand g25124(.dina(n19537), .dinb(n3858), .dout(n25357));
  jand g25125(.dina(n19539), .dinb(n3851), .dout(n25358));
  jor  g25126(.dina(n25358), .dinb(n25357), .dout(n25359));
  jor  g25127(.dina(n25359), .dinb(n25356), .dout(n25360));
  jor  g25128(.dina(n25360), .dinb(n25355), .dout(n25361));
  jxor g25129(.dina(n25361), .dinb(n25354), .dout(n25362));
  jxor g25130(.dina(n25362), .dinb(n25320), .dout(n25363));
  jnot g25131(.din(n25363), .dout(n25364));
  jand g25132(.dina(n20767), .dinb(n4449), .dout(n25365));
  jand g25133(.dina(n19529), .dinb(n4453), .dout(n25366));
  jand g25134(.dina(n19531), .dinb(n4457), .dout(n25367));
  jand g25135(.dina(n19533), .dinb(n4461), .dout(n25368));
  jor  g25136(.dina(n25368), .dinb(n25367), .dout(n25369));
  jor  g25137(.dina(n25369), .dinb(n25366), .dout(n25370));
  jor  g25138(.dina(n25370), .dinb(n25365), .dout(n25371));
  jxor g25139(.dina(n25371), .dinb(n88), .dout(n25372));
  jxor g25140(.dina(n25372), .dinb(n25364), .dout(n25373));
  jnot g25141(.din(n25119), .dout(n25374));
  jnot g25142(.din(n25152), .dout(n25375));
  jand g25143(.dina(n25375), .dinb(n25374), .dout(n25376));
  jnot g25144(.din(n25376), .dout(n25377));
  jand g25145(.dina(n25152), .dinb(n25119), .dout(n25378));
  jor  g25146(.dina(n25162), .dinb(n25378), .dout(n25379));
  jand g25147(.dina(n25379), .dinb(n25377), .dout(n25380));
  jxor g25148(.dina(n25380), .dinb(n25373), .dout(n25381));
  jand g25149(.dina(n19770), .dinb(n75), .dout(n25382));
  jand g25150(.dina(n19523), .dinb(n4933), .dout(n25383));
  jand g25151(.dina(n19525), .dinb(n4918), .dout(n25384));
  jand g25152(.dina(n19527), .dinb(n4745), .dout(n25385));
  jor  g25153(.dina(n25385), .dinb(n25384), .dout(n25386));
  jor  g25154(.dina(n25386), .dinb(n25383), .dout(n25387));
  jor  g25155(.dina(n25387), .dinb(n25382), .dout(n25388));
  jxor g25156(.dina(n25388), .dinb(n68), .dout(n25389));
  jnot g25157(.din(n25389), .dout(n25390));
  jxor g25158(.dina(n25390), .dinb(n25381), .dout(n25391));
  jxor g25159(.dina(n25391), .dinb(n25317), .dout(n25392));
  jand g25160(.dina(n21230), .dinb(n5365), .dout(n25393));
  jand g25161(.dina(n19517), .dinb(n5500), .dout(n25394));
  jand g25162(.dina(n19519), .dinb(n5424), .dout(n25395));
  jand g25163(.dina(n19521), .dinb(n5363), .dout(n25396));
  jor  g25164(.dina(n25396), .dinb(n25395), .dout(n25397));
  jor  g25165(.dina(n25397), .dinb(n25394), .dout(n25398));
  jor  g25166(.dina(n25398), .dinb(n25393), .dout(n25399));
  jxor g25167(.dina(n25399), .dinb(n72), .dout(n25400));
  jnot g25168(.din(n25400), .dout(n25401));
  jxor g25169(.dina(n25401), .dinb(n25392), .dout(n25402));
  jxor g25170(.dina(n25402), .dinb(n25314), .dout(n25403));
  jnot g25171(.din(n21762), .dout(n25404));
  jor  g25172(.dina(n25404), .dinb(n5694), .dout(n25405));
  jnot g25173(.din(n19511), .dout(n25406));
  jor  g25174(.dina(n25406), .dinb(n6208), .dout(n25407));
  jnot g25175(.din(n19513), .dout(n25408));
  jor  g25176(.dina(n25408), .dinb(n6132), .dout(n25409));
  jnot g25177(.din(n19515), .dout(n25410));
  jor  g25178(.dina(n25410), .dinb(n5692), .dout(n25411));
  jand g25179(.dina(n25411), .dinb(n25409), .dout(n25412));
  jand g25180(.dina(n25412), .dinb(n25407), .dout(n25413));
  jand g25181(.dina(n25413), .dinb(n25405), .dout(n25414));
  jxor g25182(.dina(n25414), .dinb(\a[20] ), .dout(n25415));
  jxor g25183(.dina(n25415), .dinb(n25403), .dout(n25416));
  jxor g25184(.dina(n25416), .dinb(n25310), .dout(n25417));
  jand g25185(.dina(n22250), .dinb(n6340), .dout(n25418));
  jand g25186(.dina(n22248), .dinb(n6798), .dout(n25419));
  jand g25187(.dina(n19758), .dinb(n6556), .dout(n25420));
  jand g25188(.dina(n19510), .dinb(n6338), .dout(n25421));
  jor  g25189(.dina(n25421), .dinb(n25420), .dout(n25422));
  jor  g25190(.dina(n25422), .dinb(n25419), .dout(n25423));
  jor  g25191(.dina(n25423), .dinb(n25418), .dout(n25424));
  jxor g25192(.dina(n25424), .dinb(n5064), .dout(n25425));
  jxor g25193(.dina(n25425), .dinb(n25417), .dout(n25426));
  jxor g25194(.dina(n25426), .dinb(n25306), .dout(n25427));
  jand g25195(.dina(n22605), .dinb(n6936), .dout(n25428));
  jand g25196(.dina(n22603), .dinb(n7741), .dout(n25429));
  jand g25197(.dina(n22539), .dinb(n7613), .dout(n25430));
  jand g25198(.dina(n22540), .dinb(n6934), .dout(n25431));
  jor  g25199(.dina(n25431), .dinb(n25430), .dout(n25432));
  jor  g25200(.dina(n25432), .dinb(n25429), .dout(n25433));
  jor  g25201(.dina(n25433), .dinb(n25428), .dout(n25434));
  jxor g25202(.dina(n25434), .dinb(n5292), .dout(n25435));
  jxor g25203(.dina(n25435), .dinb(n25427), .dout(n25436));
  jxor g25204(.dina(n25436), .dinb(n25302), .dout(n25437));
  jxor g25205(.dina(n25437), .dinb(n25299), .dout(n25438));
  jxor g25206(.dina(n25438), .dinb(n25290), .dout(n25439));
  jor  g25207(.dina(n24337), .dinb(n8772), .dout(n25440));
  jor  g25208(.dina(n24335), .dinb(n9490), .dout(n25441));
  jor  g25209(.dina(n24142), .dinb(n9127), .dout(n25442));
  jor  g25210(.dina(n23921), .dinb(n8770), .dout(n25443));
  jand g25211(.dina(n25443), .dinb(n25442), .dout(n25444));
  jand g25212(.dina(n25444), .dinb(n25441), .dout(n25445));
  jand g25213(.dina(n25445), .dinb(n25440), .dout(n25446));
  jxor g25214(.dina(n25446), .dinb(\a[8] ), .dout(n25447));
  jxor g25215(.dina(n25447), .dinb(n25439), .dout(n25448));
  jxor g25216(.dina(n25448), .dinb(n25286), .dout(n25449));
  jxor g25217(.dina(n25449), .dinb(n25283), .dout(n25450));
  jxor g25218(.dina(n25450), .dinb(n25280), .dout(\result[11] ));
  jand g25219(.dina(n25450), .dinb(n25280), .dout(n25452));
  jand g25220(.dina(n25436), .dinb(n25302), .dout(n25453));
  jand g25221(.dina(n25437), .dinb(n25299), .dout(n25454));
  jor  g25222(.dina(n25454), .dinb(n25453), .dout(n25455));
  jor  g25223(.dina(n24357), .dinb(n8772), .dout(n25456));
  jor  g25224(.dina(n24335), .dinb(n15985), .dout(n25457));
  jor  g25225(.dina(n24142), .dinb(n8770), .dout(n25458));
  jand g25226(.dina(n25458), .dinb(n25457), .dout(n25459));
  jand g25227(.dina(n25459), .dinb(n25456), .dout(n25460));
  jxor g25228(.dina(n25460), .dinb(\a[8] ), .dout(n25461));
  jnot g25229(.din(n25461), .dout(n25462));
  jxor g25230(.dina(n25462), .dinb(n25455), .dout(n25463));
  jnot g25231(.din(n21086), .dout(n25464));
  jor  g25232(.dina(n25464), .dinb(n4747), .dout(n25465));
  jnot g25233(.din(n19521), .dout(n25466));
  jor  g25234(.dina(n25466), .dinb(n4959), .dout(n25467));
  jnot g25235(.din(n19523), .dout(n25468));
  jor  g25236(.dina(n25468), .dinb(n4919), .dout(n25469));
  jnot g25237(.din(n19525), .dout(n25470));
  jor  g25238(.dina(n25470), .dinb(n4746), .dout(n25471));
  jand g25239(.dina(n25471), .dinb(n25469), .dout(n25472));
  jand g25240(.dina(n25472), .dinb(n25467), .dout(n25473));
  jand g25241(.dina(n25473), .dinb(n25465), .dout(n25474));
  jxor g25242(.dina(n25474), .dinb(\a[26] ), .dout(n25475));
  jnot g25243(.din(n25475), .dout(n25476));
  jand g25244(.dina(n25362), .dinb(n25320), .dout(n25477));
  jnot g25245(.din(n25477), .dout(n25478));
  jor  g25246(.dina(n25372), .dinb(n25364), .dout(n25479));
  jand g25247(.dina(n25479), .dinb(n25478), .dout(n25480));
  jnot g25248(.din(n25480), .dout(n25481));
  jand g25249(.dina(n532), .dinb(n146), .dout(n25482));
  jand g25250(.dina(n25482), .dinb(n1066), .dout(n25483));
  jand g25251(.dina(n1785), .dinb(n1142), .dout(n25484));
  jand g25252(.dina(n25484), .dinb(n25483), .dout(n25485));
  jand g25253(.dina(n5166), .dinb(n513), .dout(n25486));
  jand g25254(.dina(n25486), .dinb(n25485), .dout(n25487));
  jand g25255(.dina(n3260), .dinb(n3250), .dout(n25488));
  jand g25256(.dina(n25488), .dinb(n2533), .dout(n25489));
  jand g25257(.dina(n25489), .dinb(n1835), .dout(n25490));
  jand g25258(.dina(n25490), .dinb(n25487), .dout(n25491));
  jand g25259(.dina(n25491), .dinb(n3192), .dout(n25492));
  jand g25260(.dina(n678), .dinb(n234), .dout(n25493));
  jand g25261(.dina(n25493), .dinb(n515), .dout(n25494));
  jand g25262(.dina(n819), .dinb(n472), .dout(n25495));
  jand g25263(.dina(n583), .dinb(n557), .dout(n25496));
  jand g25264(.dina(n25496), .dinb(n25495), .dout(n25497));
  jand g25265(.dina(n25497), .dinb(n12435), .dout(n25498));
  jand g25266(.dina(n25498), .dinb(n25494), .dout(n25499));
  jand g25267(.dina(n842), .dinb(n486), .dout(n25500));
  jand g25268(.dina(n757), .dinb(n432), .dout(n25501));
  jand g25269(.dina(n25501), .dinb(n25500), .dout(n25502));
  jand g25270(.dina(n703), .dinb(n409), .dout(n25503));
  jand g25271(.dina(n25503), .dinb(n3563), .dout(n25504));
  jand g25272(.dina(n25504), .dinb(n25502), .dout(n25505));
  jand g25273(.dina(n12544), .dinb(n7065), .dout(n25506));
  jand g25274(.dina(n25506), .dinb(n25505), .dout(n25507));
  jand g25275(.dina(n25507), .dinb(n25499), .dout(n25508));
  jand g25276(.dina(n25508), .dinb(n4057), .dout(n25509));
  jand g25277(.dina(n25509), .dinb(n3984), .dout(n25510));
  jand g25278(.dina(n25510), .dinb(n25492), .dout(n25511));
  jand g25279(.dina(n25511), .dinb(n12246), .dout(n25512));
  jxor g25280(.dina(n25512), .dinb(n25353), .dout(n25513));
  jand g25281(.dina(n25353), .dinb(n25324), .dout(n25514));
  jnot g25282(.din(n25514), .dout(n25515));
  jnot g25283(.din(n25324), .dout(n25516));
  jand g25284(.dina(n25352), .dinb(n25516), .dout(n25517));
  jor  g25285(.dina(n25361), .dinb(n25517), .dout(n25518));
  jand g25286(.dina(n25518), .dinb(n25515), .dout(n25519));
  jxor g25287(.dina(n25519), .dinb(n25513), .dout(n25520));
  jand g25288(.dina(n20399), .dinb(n732), .dout(n25521));
  jand g25289(.dina(n19533), .dinb(n3855), .dout(n25522));
  jand g25290(.dina(n19535), .dinb(n3858), .dout(n25523));
  jand g25291(.dina(n19537), .dinb(n3851), .dout(n25524));
  jor  g25292(.dina(n25524), .dinb(n25523), .dout(n25525));
  jor  g25293(.dina(n25525), .dinb(n25522), .dout(n25526));
  jor  g25294(.dina(n25526), .dinb(n25521), .dout(n25527));
  jxor g25295(.dina(n25527), .dinb(n25520), .dout(n25528));
  jxor g25296(.dina(n25528), .dinb(n25481), .dout(n25529));
  jnot g25297(.din(n25529), .dout(n25530));
  jand g25298(.dina(n20793), .dinb(n4449), .dout(n25531));
  jand g25299(.dina(n19527), .dinb(n4453), .dout(n25532));
  jand g25300(.dina(n19529), .dinb(n4457), .dout(n25533));
  jand g25301(.dina(n19531), .dinb(n4461), .dout(n25534));
  jor  g25302(.dina(n25534), .dinb(n25533), .dout(n25535));
  jor  g25303(.dina(n25535), .dinb(n25532), .dout(n25536));
  jor  g25304(.dina(n25536), .dinb(n25531), .dout(n25537));
  jxor g25305(.dina(n25537), .dinb(n88), .dout(n25538));
  jxor g25306(.dina(n25538), .dinb(n25530), .dout(n25539));
  jxor g25307(.dina(n25539), .dinb(n25476), .dout(n25540));
  jor  g25308(.dina(n25380), .dinb(n25373), .dout(n25541));
  jand g25309(.dina(n25380), .dinb(n25373), .dout(n25542));
  jor  g25310(.dina(n25390), .dinb(n25542), .dout(n25543));
  jand g25311(.dina(n25543), .dinb(n25541), .dout(n25544));
  jnot g25312(.din(n25544), .dout(n25545));
  jxor g25313(.dina(n25545), .dinb(n25540), .dout(n25546));
  jnot g25314(.din(n21218), .dout(n25547));
  jor  g25315(.dina(n25547), .dinb(n5366), .dout(n25548));
  jor  g25316(.dina(n25410), .dinb(n5499), .dout(n25549));
  jnot g25317(.din(n19517), .dout(n25550));
  jor  g25318(.dina(n25550), .dinb(n5425), .dout(n25551));
  jnot g25319(.din(n19519), .dout(n25552));
  jor  g25320(.dina(n25552), .dinb(n5364), .dout(n25553));
  jand g25321(.dina(n25553), .dinb(n25551), .dout(n25554));
  jand g25322(.dina(n25554), .dinb(n25549), .dout(n25555));
  jand g25323(.dina(n25555), .dinb(n25548), .dout(n25556));
  jxor g25324(.dina(n25556), .dinb(\a[23] ), .dout(n25557));
  jxor g25325(.dina(n25557), .dinb(n25546), .dout(n25558));
  jnot g25326(.din(n25317), .dout(n25559));
  jnot g25327(.din(n25391), .dout(n25560));
  jand g25328(.dina(n25560), .dinb(n25559), .dout(n25561));
  jnot g25329(.din(n25561), .dout(n25562));
  jand g25330(.dina(n25391), .dinb(n25317), .dout(n25563));
  jor  g25331(.dina(n25401), .dinb(n25563), .dout(n25564));
  jand g25332(.dina(n25564), .dinb(n25562), .dout(n25565));
  jnot g25333(.din(n25565), .dout(n25566));
  jxor g25334(.dina(n25566), .dinb(n25558), .dout(n25567));
  jnot g25335(.din(n21750), .dout(n25568));
  jor  g25336(.dina(n25568), .dinb(n5694), .dout(n25569));
  jnot g25337(.din(n19510), .dout(n25570));
  jor  g25338(.dina(n25570), .dinb(n6208), .dout(n25571));
  jor  g25339(.dina(n25406), .dinb(n6132), .dout(n25572));
  jor  g25340(.dina(n25408), .dinb(n5692), .dout(n25573));
  jand g25341(.dina(n25573), .dinb(n25572), .dout(n25574));
  jand g25342(.dina(n25574), .dinb(n25571), .dout(n25575));
  jand g25343(.dina(n25575), .dinb(n25569), .dout(n25576));
  jxor g25344(.dina(n25576), .dinb(\a[20] ), .dout(n25577));
  jxor g25345(.dina(n25577), .dinb(n25567), .dout(n25578));
  jnot g25346(.din(n25402), .dout(n25579));
  jand g25347(.dina(n25579), .dinb(n25314), .dout(n25580));
  jnot g25348(.din(n25580), .dout(n25581));
  jnot g25349(.din(n25314), .dout(n25582));
  jand g25350(.dina(n25402), .dinb(n25582), .dout(n25583));
  jnot g25351(.din(n25415), .dout(n25584));
  jor  g25352(.dina(n25584), .dinb(n25583), .dout(n25585));
  jand g25353(.dina(n25585), .dinb(n25581), .dout(n25586));
  jnot g25354(.din(n25586), .dout(n25587));
  jxor g25355(.dina(n25587), .dinb(n25578), .dout(n25588));
  jnot g25356(.din(n22627), .dout(n25589));
  jor  g25357(.dina(n25589), .dinb(n6341), .dout(n25590));
  jnot g25358(.din(n22540), .dout(n25591));
  jor  g25359(.dina(n25591), .dinb(n6797), .dout(n25592));
  jnot g25360(.din(n22248), .dout(n25593));
  jor  g25361(.dina(n25593), .dinb(n6557), .dout(n25594));
  jnot g25362(.din(n19758), .dout(n25595));
  jor  g25363(.dina(n25595), .dinb(n6339), .dout(n25596));
  jand g25364(.dina(n25596), .dinb(n25594), .dout(n25597));
  jand g25365(.dina(n25597), .dinb(n25592), .dout(n25598));
  jand g25366(.dina(n25598), .dinb(n25590), .dout(n25599));
  jxor g25367(.dina(n25599), .dinb(\a[17] ), .dout(n25600));
  jxor g25368(.dina(n25600), .dinb(n25588), .dout(n25601));
  jnot g25369(.din(n25416), .dout(n25602));
  jand g25370(.dina(n25602), .dinb(n25310), .dout(n25603));
  jnot g25371(.din(n25310), .dout(n25604));
  jand g25372(.dina(n25416), .dinb(n25604), .dout(n25605));
  jnot g25373(.din(n25605), .dout(n25606));
  jand g25374(.dina(n25425), .dinb(n25606), .dout(n25607));
  jor  g25375(.dina(n25607), .dinb(n25603), .dout(n25608));
  jxor g25376(.dina(n25608), .dinb(n25601), .dout(n25609));
  jor  g25377(.dina(n23730), .dinb(n6937), .dout(n25610));
  jor  g25378(.dina(n23450), .dinb(n7740), .dout(n25611));
  jor  g25379(.dina(n23449), .dinb(n7614), .dout(n25612));
  jor  g25380(.dina(n23734), .dinb(n6935), .dout(n25613));
  jand g25381(.dina(n25613), .dinb(n25612), .dout(n25614));
  jand g25382(.dina(n25614), .dinb(n25611), .dout(n25615));
  jand g25383(.dina(n25615), .dinb(n25610), .dout(n25616));
  jxor g25384(.dina(n25616), .dinb(\a[14] ), .dout(n25617));
  jxor g25385(.dina(n25617), .dinb(n25609), .dout(n25618));
  jnot g25386(.din(n25426), .dout(n25619));
  jand g25387(.dina(n25619), .dinb(n25306), .dout(n25620));
  jnot g25388(.din(n25306), .dout(n25621));
  jand g25389(.dina(n25426), .dinb(n25621), .dout(n25622));
  jnot g25390(.din(n25622), .dout(n25623));
  jand g25391(.dina(n25435), .dinb(n25623), .dout(n25624));
  jor  g25392(.dina(n25624), .dinb(n25620), .dout(n25625));
  jxor g25393(.dina(n25625), .dinb(n25618), .dout(n25626));
  jor  g25394(.dina(n23919), .dinb(n7891), .dout(n25627));
  jor  g25395(.dina(n23921), .dinb(n8440), .dout(n25628));
  jor  g25396(.dina(n23710), .dinb(n8155), .dout(n25629));
  jor  g25397(.dina(n23496), .dinb(n7889), .dout(n25630));
  jand g25398(.dina(n25630), .dinb(n25629), .dout(n25631));
  jand g25399(.dina(n25631), .dinb(n25628), .dout(n25632));
  jand g25400(.dina(n25632), .dinb(n25627), .dout(n25633));
  jxor g25401(.dina(n25633), .dinb(\a[11] ), .dout(n25634));
  jxor g25402(.dina(n25634), .dinb(n25626), .dout(n25635));
  jxor g25403(.dina(n25635), .dinb(n25463), .dout(n25636));
  jnot g25404(.din(n25438), .dout(n25637));
  jand g25405(.dina(n25637), .dinb(n25290), .dout(n25638));
  jnot g25406(.din(n25638), .dout(n25639));
  jnot g25407(.din(n25290), .dout(n25640));
  jand g25408(.dina(n25438), .dinb(n25640), .dout(n25641));
  jnot g25409(.din(n25447), .dout(n25642));
  jor  g25410(.dina(n25642), .dinb(n25641), .dout(n25643));
  jand g25411(.dina(n25643), .dinb(n25639), .dout(n25644));
  jxor g25412(.dina(n25644), .dinb(n25636), .dout(n25645));
  jand g25413(.dina(n25448), .dinb(n25286), .dout(n25646));
  jand g25414(.dina(n25449), .dinb(n25283), .dout(n25647));
  jor  g25415(.dina(n25647), .dinb(n25646), .dout(n25648));
  jxor g25416(.dina(n25648), .dinb(n25645), .dout(n25649));
  jxor g25417(.dina(n25649), .dinb(n25452), .dout(\result[12] ));
  jand g25418(.dina(n25649), .dinb(n25452), .dout(n25651));
  jand g25419(.dina(n25644), .dinb(n25636), .dout(n25652));
  jand g25420(.dina(n25648), .dinb(n25645), .dout(n25653));
  jor  g25421(.dina(n25653), .dinb(n25652), .dout(n25654));
  jor  g25422(.dina(n25538), .dinb(n25530), .dout(n25655));
  jand g25423(.dina(n25539), .dinb(n25476), .dout(n25656));
  jnot g25424(.din(n25656), .dout(n25657));
  jand g25425(.dina(n25657), .dinb(n25655), .dout(n25658));
  jand g25426(.dina(n25527), .dinb(n25520), .dout(n25659));
  jand g25427(.dina(n25528), .dinb(n25481), .dout(n25660));
  jor  g25428(.dina(n25660), .dinb(n25659), .dout(n25661));
  jand g25429(.dina(n20781), .dinb(n4449), .dout(n25662));
  jand g25430(.dina(n19525), .dinb(n4453), .dout(n25663));
  jand g25431(.dina(n19527), .dinb(n4457), .dout(n25664));
  jand g25432(.dina(n19529), .dinb(n4461), .dout(n25665));
  jor  g25433(.dina(n25665), .dinb(n25664), .dout(n25666));
  jor  g25434(.dina(n25666), .dinb(n25663), .dout(n25667));
  jor  g25435(.dina(n25667), .dinb(n25662), .dout(n25668));
  jxor g25436(.dina(n25668), .dinb(n88), .dout(n25669));
  jnot g25437(.din(n25669), .dout(n25670));
  jor  g25438(.dina(n25512), .dinb(n25353), .dout(n25671));
  jand g25439(.dina(n25519), .dinb(n25513), .dout(n25672));
  jnot g25440(.din(n25672), .dout(n25673));
  jand g25441(.dina(n25673), .dinb(n25671), .dout(n25674));
  jnot g25442(.din(n25674), .dout(n25675));
  jand g25443(.dina(n24593), .dinb(n13259), .dout(n25676));
  jxor g25444(.dina(n25676), .dinb(n6039), .dout(n25677));
  jand g25445(.dina(n1399), .dinb(n1162), .dout(n25678));
  jand g25446(.dina(n25678), .dinb(n2306), .dout(n25679));
  jand g25447(.dina(n1930), .dinb(n1067), .dout(n25680));
  jand g25448(.dina(n25680), .dinb(n596), .dout(n25681));
  jand g25449(.dina(n897), .dinb(n793), .dout(n25682));
  jand g25450(.dina(n25682), .dinb(n820), .dout(n25683));
  jand g25451(.dina(n25683), .dinb(n12232), .dout(n25684));
  jand g25452(.dina(n25684), .dinb(n25681), .dout(n25685));
  jand g25453(.dina(n25685), .dinb(n12214), .dout(n25686));
  jand g25454(.dina(n25686), .dinb(n25679), .dout(n25687));
  jand g25455(.dina(n25687), .dinb(n2822), .dout(n25688));
  jand g25456(.dina(n3626), .dinb(n1255), .dout(n25689));
  jand g25457(.dina(n25689), .dinb(n25688), .dout(n25690));
  jxor g25458(.dina(n25690), .dinb(n25352), .dout(n25691));
  jxor g25459(.dina(n25691), .dinb(n25677), .dout(n25692));
  jxor g25460(.dina(n25692), .dinb(n25675), .dout(n25693));
  jand g25461(.dina(n19780), .dinb(n732), .dout(n25694));
  jand g25462(.dina(n19531), .dinb(n3855), .dout(n25695));
  jand g25463(.dina(n19533), .dinb(n3858), .dout(n25696));
  jand g25464(.dina(n19535), .dinb(n3851), .dout(n25697));
  jor  g25465(.dina(n25697), .dinb(n25696), .dout(n25698));
  jor  g25466(.dina(n25698), .dinb(n25695), .dout(n25699));
  jor  g25467(.dina(n25699), .dinb(n25694), .dout(n25700));
  jxor g25468(.dina(n25700), .dinb(n25693), .dout(n25701));
  jxor g25469(.dina(n25701), .dinb(n25670), .dout(n25702));
  jxor g25470(.dina(n25702), .dinb(n25661), .dout(n25703));
  jnot g25471(.din(n25703), .dout(n25704));
  jand g25472(.dina(n21240), .dinb(n75), .dout(n25705));
  jand g25473(.dina(n19519), .dinb(n4933), .dout(n25706));
  jand g25474(.dina(n19521), .dinb(n4918), .dout(n25707));
  jand g25475(.dina(n19523), .dinb(n4745), .dout(n25708));
  jor  g25476(.dina(n25708), .dinb(n25707), .dout(n25709));
  jor  g25477(.dina(n25709), .dinb(n25706), .dout(n25710));
  jor  g25478(.dina(n25710), .dinb(n25705), .dout(n25711));
  jxor g25479(.dina(n25711), .dinb(n68), .dout(n25712));
  jxor g25480(.dina(n25712), .dinb(n25704), .dout(n25713));
  jnot g25481(.din(n25713), .dout(n25714));
  jxor g25482(.dina(n25714), .dinb(n25658), .dout(n25715));
  jand g25483(.dina(n21738), .dinb(n5365), .dout(n25716));
  jand g25484(.dina(n19513), .dinb(n5500), .dout(n25717));
  jand g25485(.dina(n19515), .dinb(n5424), .dout(n25718));
  jand g25486(.dina(n19517), .dinb(n5363), .dout(n25719));
  jor  g25487(.dina(n25719), .dinb(n25718), .dout(n25720));
  jor  g25488(.dina(n25720), .dinb(n25717), .dout(n25721));
  jor  g25489(.dina(n25721), .dinb(n25716), .dout(n25722));
  jxor g25490(.dina(n25722), .dinb(n72), .dout(n25723));
  jxor g25491(.dina(n25723), .dinb(n25715), .dout(n25724));
  jnot g25492(.din(n25540), .dout(n25725));
  jand g25493(.dina(n25545), .dinb(n25725), .dout(n25726));
  jnot g25494(.din(n25726), .dout(n25727));
  jand g25495(.dina(n25544), .dinb(n25540), .dout(n25728));
  jnot g25496(.din(n25557), .dout(n25729));
  jor  g25497(.dina(n25729), .dinb(n25728), .dout(n25730));
  jand g25498(.dina(n25730), .dinb(n25727), .dout(n25731));
  jnot g25499(.din(n25731), .dout(n25732));
  jxor g25500(.dina(n25732), .dinb(n25724), .dout(n25733));
  jand g25501(.dina(n19760), .dinb(n5693), .dout(n25734));
  jand g25502(.dina(n19758), .dinb(n6209), .dout(n25735));
  jand g25503(.dina(n19510), .dinb(n6131), .dout(n25736));
  jand g25504(.dina(n19511), .dinb(n5691), .dout(n25737));
  jor  g25505(.dina(n25737), .dinb(n25736), .dout(n25738));
  jor  g25506(.dina(n25738), .dinb(n25735), .dout(n25739));
  jor  g25507(.dina(n25739), .dinb(n25734), .dout(n25740));
  jxor g25508(.dina(n25740), .dinb(n4247), .dout(n25741));
  jxor g25509(.dina(n25741), .dinb(n25733), .dout(n25742));
  jnot g25510(.din(n25558), .dout(n25743));
  jand g25511(.dina(n25566), .dinb(n25743), .dout(n25744));
  jnot g25512(.din(n25744), .dout(n25745));
  jand g25513(.dina(n25565), .dinb(n25558), .dout(n25746));
  jnot g25514(.din(n25577), .dout(n25747));
  jor  g25515(.dina(n25747), .dinb(n25746), .dout(n25748));
  jand g25516(.dina(n25748), .dinb(n25745), .dout(n25749));
  jnot g25517(.din(n25749), .dout(n25750));
  jxor g25518(.dina(n25750), .dinb(n25742), .dout(n25751));
  jand g25519(.dina(n22617), .dinb(n6340), .dout(n25752));
  jand g25520(.dina(n22539), .dinb(n6798), .dout(n25753));
  jand g25521(.dina(n22540), .dinb(n6556), .dout(n25754));
  jand g25522(.dina(n22248), .dinb(n6338), .dout(n25755));
  jor  g25523(.dina(n25755), .dinb(n25754), .dout(n25756));
  jor  g25524(.dina(n25756), .dinb(n25753), .dout(n25757));
  jor  g25525(.dina(n25757), .dinb(n25752), .dout(n25758));
  jxor g25526(.dina(n25758), .dinb(n5064), .dout(n25759));
  jnot g25527(.din(n25759), .dout(n25760));
  jnot g25528(.din(n25578), .dout(n25761));
  jand g25529(.dina(n25587), .dinb(n25761), .dout(n25762));
  jnot g25530(.din(n25762), .dout(n25763));
  jand g25531(.dina(n25586), .dinb(n25578), .dout(n25764));
  jnot g25532(.din(n25600), .dout(n25765));
  jor  g25533(.dina(n25765), .dinb(n25764), .dout(n25766));
  jand g25534(.dina(n25766), .dinb(n25763), .dout(n25767));
  jxor g25535(.dina(n25767), .dinb(n25760), .dout(n25768));
  jxor g25536(.dina(n25768), .dinb(n25751), .dout(n25769));
  jor  g25537(.dina(n23494), .dinb(n6937), .dout(n25770));
  jor  g25538(.dina(n23496), .dinb(n7740), .dout(n25771));
  jor  g25539(.dina(n23450), .dinb(n7614), .dout(n25772));
  jor  g25540(.dina(n23449), .dinb(n6935), .dout(n25773));
  jand g25541(.dina(n25773), .dinb(n25772), .dout(n25774));
  jand g25542(.dina(n25774), .dinb(n25771), .dout(n25775));
  jand g25543(.dina(n25775), .dinb(n25770), .dout(n25776));
  jxor g25544(.dina(n25776), .dinb(\a[14] ), .dout(n25777));
  jxor g25545(.dina(n25777), .dinb(n25769), .dout(n25778));
  jnot g25546(.din(n25601), .dout(n25779));
  jand g25547(.dina(n25608), .dinb(n25779), .dout(n25780));
  jnot g25548(.din(n25780), .dout(n25781));
  jnot g25549(.din(n25608), .dout(n25782));
  jand g25550(.dina(n25782), .dinb(n25601), .dout(n25783));
  jnot g25551(.din(n25617), .dout(n25784));
  jor  g25552(.dina(n25784), .dinb(n25783), .dout(n25785));
  jand g25553(.dina(n25785), .dinb(n25781), .dout(n25786));
  jnot g25554(.din(n25786), .dout(n25787));
  jxor g25555(.dina(n25787), .dinb(n25778), .dout(n25788));
  jor  g25556(.dina(n24140), .dinb(n7891), .dout(n25789));
  jor  g25557(.dina(n24142), .dinb(n8440), .dout(n25790));
  jor  g25558(.dina(n23921), .dinb(n8155), .dout(n25791));
  jor  g25559(.dina(n23710), .dinb(n7889), .dout(n25792));
  jand g25560(.dina(n25792), .dinb(n25791), .dout(n25793));
  jand g25561(.dina(n25793), .dinb(n25790), .dout(n25794));
  jand g25562(.dina(n25794), .dinb(n25789), .dout(n25795));
  jxor g25563(.dina(n25795), .dinb(\a[11] ), .dout(n25796));
  jnot g25564(.din(n25796), .dout(n25797));
  jnot g25565(.din(n25618), .dout(n25798));
  jand g25566(.dina(n25625), .dinb(n25798), .dout(n25799));
  jnot g25567(.din(n25799), .dout(n25800));
  jnot g25568(.din(n25625), .dout(n25801));
  jand g25569(.dina(n25801), .dinb(n25618), .dout(n25802));
  jnot g25570(.din(n25634), .dout(n25803));
  jor  g25571(.dina(n25803), .dinb(n25802), .dout(n25804));
  jand g25572(.dina(n25804), .dinb(n25800), .dout(n25805));
  jxor g25573(.dina(n25805), .dinb(n25797), .dout(n25806));
  jxor g25574(.dina(n25806), .dinb(n25788), .dout(n25807));
  jnot g25575(.din(n25455), .dout(n25808));
  jand g25576(.dina(n25461), .dinb(n25808), .dout(n25809));
  jnot g25577(.din(n25809), .dout(n25810));
  jand g25578(.dina(n25462), .dinb(n25455), .dout(n25811));
  jor  g25579(.dina(n25635), .dinb(n25811), .dout(n25812));
  jand g25580(.dina(n25812), .dinb(n25810), .dout(n25813));
  jxor g25581(.dina(n25813), .dinb(n25807), .dout(n25814));
  jxor g25582(.dina(n25814), .dinb(n25654), .dout(n25815));
  jxor g25583(.dina(n25815), .dinb(n25651), .dout(\result[13] ));
  jand g25584(.dina(n25815), .dinb(n25651), .dout(n25817));
  jand g25585(.dina(n25813), .dinb(n25807), .dout(n25818));
  jand g25586(.dina(n25814), .dinb(n25654), .dout(n25819));
  jor  g25587(.dina(n25819), .dinb(n25818), .dout(n25820));
  jand g25588(.dina(n25805), .dinb(n25797), .dout(n25821));
  jand g25589(.dina(n25806), .dinb(n25788), .dout(n25822));
  jor  g25590(.dina(n25822), .dinb(n25821), .dout(n25823));
  jnot g25591(.din(n25769), .dout(n25824));
  jor  g25592(.dina(n25777), .dinb(n25824), .dout(n25825));
  jor  g25593(.dina(n25787), .dinb(n25778), .dout(n25826));
  jand g25594(.dina(n25826), .dinb(n25825), .dout(n25827));
  jor  g25595(.dina(n23708), .dinb(n6937), .dout(n25828));
  jor  g25596(.dina(n23710), .dinb(n7740), .dout(n25829));
  jor  g25597(.dina(n23496), .dinb(n7614), .dout(n25830));
  jor  g25598(.dina(n23450), .dinb(n6935), .dout(n25831));
  jand g25599(.dina(n25831), .dinb(n25830), .dout(n25832));
  jand g25600(.dina(n25832), .dinb(n25829), .dout(n25833));
  jand g25601(.dina(n25833), .dinb(n25828), .dout(n25834));
  jxor g25602(.dina(n25834), .dinb(\a[14] ), .dout(n25835));
  jnot g25603(.din(n25835), .dout(n25836));
  jand g25604(.dina(n25767), .dinb(n25760), .dout(n25837));
  jand g25605(.dina(n25768), .dinb(n25751), .dout(n25838));
  jor  g25606(.dina(n25838), .dinb(n25837), .dout(n25839));
  jnot g25607(.din(n25733), .dout(n25840));
  jor  g25608(.dina(n25741), .dinb(n25840), .dout(n25841));
  jor  g25609(.dina(n25750), .dinb(n25742), .dout(n25842));
  jand g25610(.dina(n25842), .dinb(n25841), .dout(n25843));
  jnot g25611(.din(n25715), .dout(n25844));
  jor  g25612(.dina(n25723), .dinb(n25844), .dout(n25845));
  jor  g25613(.dina(n25732), .dinb(n25724), .dout(n25846));
  jand g25614(.dina(n25846), .dinb(n25845), .dout(n25847));
  jor  g25615(.dina(n25712), .dinb(n25704), .dout(n25848));
  jor  g25616(.dina(n25714), .dinb(n25658), .dout(n25849));
  jand g25617(.dina(n25849), .dinb(n25848), .dout(n25850));
  jand g25618(.dina(n25701), .dinb(n25670), .dout(n25851));
  jand g25619(.dina(n25702), .dinb(n25661), .dout(n25852));
  jor  g25620(.dina(n25852), .dinb(n25851), .dout(n25853));
  jor  g25621(.dina(n25690), .dinb(n25352), .dout(n25854));
  jand g25622(.dina(n25691), .dinb(n25677), .dout(n25855));
  jnot g25623(.din(n25855), .dout(n25856));
  jand g25624(.dina(n25856), .dinb(n25854), .dout(n25857));
  jand g25625(.dina(n595), .dinb(n533), .dout(n25858));
  jand g25626(.dina(n25858), .dinb(n687), .dout(n25859));
  jand g25627(.dina(n25859), .dinb(n3467), .dout(n25860));
  jand g25628(.dina(n14328), .dinb(n2354), .dout(n25861));
  jand g25629(.dina(n25861), .dinb(n25860), .dout(n25862));
  jand g25630(.dina(n812), .dinb(n429), .dout(n25863));
  jand g25631(.dina(n13196), .dinb(n3483), .dout(n25864));
  jand g25632(.dina(n25864), .dinb(n25863), .dout(n25865));
  jand g25633(.dina(n25865), .dinb(n5559), .dout(n25866));
  jand g25634(.dina(n25866), .dinb(n25862), .dout(n25867));
  jand g25635(.dina(n25867), .dinb(n13091), .dout(n25868));
  jand g25636(.dina(n25868), .dinb(n1030), .dout(n25869));
  jand g25637(.dina(n25869), .dinb(n2543), .dout(n25870));
  jnot g25638(.din(n25870), .dout(n25871));
  jxor g25639(.dina(n25871), .dinb(n25857), .dout(n25872));
  jand g25640(.dina(n20767), .dinb(n732), .dout(n25873));
  jand g25641(.dina(n19529), .dinb(n3855), .dout(n25874));
  jand g25642(.dina(n19531), .dinb(n3858), .dout(n25875));
  jand g25643(.dina(n19533), .dinb(n3851), .dout(n25876));
  jor  g25644(.dina(n25876), .dinb(n25875), .dout(n25877));
  jor  g25645(.dina(n25877), .dinb(n25874), .dout(n25878));
  jor  g25646(.dina(n25878), .dinb(n25873), .dout(n25879));
  jxor g25647(.dina(n25879), .dinb(n25872), .dout(n25880));
  jor  g25648(.dina(n25692), .dinb(n25675), .dout(n25881));
  jand g25649(.dina(n25692), .dinb(n25675), .dout(n25882));
  jor  g25650(.dina(n25700), .dinb(n25882), .dout(n25883));
  jand g25651(.dina(n25883), .dinb(n25881), .dout(n25884));
  jxor g25652(.dina(n25884), .dinb(n25880), .dout(n25885));
  jnot g25653(.din(n25885), .dout(n25886));
  jand g25654(.dina(n19770), .dinb(n4449), .dout(n25887));
  jand g25655(.dina(n19523), .dinb(n4453), .dout(n25888));
  jand g25656(.dina(n19525), .dinb(n4457), .dout(n25889));
  jand g25657(.dina(n19527), .dinb(n4461), .dout(n25890));
  jor  g25658(.dina(n25890), .dinb(n25889), .dout(n25891));
  jor  g25659(.dina(n25891), .dinb(n25888), .dout(n25892));
  jor  g25660(.dina(n25892), .dinb(n25887), .dout(n25893));
  jxor g25661(.dina(n25893), .dinb(n88), .dout(n25894));
  jxor g25662(.dina(n25894), .dinb(n25886), .dout(n25895));
  jxor g25663(.dina(n25895), .dinb(n25853), .dout(n25896));
  jand g25664(.dina(n21230), .dinb(n75), .dout(n25897));
  jand g25665(.dina(n19517), .dinb(n4933), .dout(n25898));
  jand g25666(.dina(n19519), .dinb(n4918), .dout(n25899));
  jand g25667(.dina(n19521), .dinb(n4745), .dout(n25900));
  jor  g25668(.dina(n25900), .dinb(n25899), .dout(n25901));
  jor  g25669(.dina(n25901), .dinb(n25898), .dout(n25902));
  jor  g25670(.dina(n25902), .dinb(n25897), .dout(n25903));
  jxor g25671(.dina(n25903), .dinb(n68), .dout(n25904));
  jnot g25672(.din(n25904), .dout(n25905));
  jxor g25673(.dina(n25905), .dinb(n25896), .dout(n25906));
  jnot g25674(.din(n25906), .dout(n25907));
  jxor g25675(.dina(n25907), .dinb(n25850), .dout(n25908));
  jand g25676(.dina(n21762), .dinb(n5365), .dout(n25909));
  jand g25677(.dina(n19511), .dinb(n5500), .dout(n25910));
  jand g25678(.dina(n19513), .dinb(n5424), .dout(n25911));
  jand g25679(.dina(n19515), .dinb(n5363), .dout(n25912));
  jor  g25680(.dina(n25912), .dinb(n25911), .dout(n25913));
  jor  g25681(.dina(n25913), .dinb(n25910), .dout(n25914));
  jor  g25682(.dina(n25914), .dinb(n25909), .dout(n25915));
  jxor g25683(.dina(n25915), .dinb(n72), .dout(n25916));
  jnot g25684(.din(n25916), .dout(n25917));
  jxor g25685(.dina(n25917), .dinb(n25908), .dout(n25918));
  jxor g25686(.dina(n25918), .dinb(n25847), .dout(n25919));
  jand g25687(.dina(n22250), .dinb(n5693), .dout(n25920));
  jand g25688(.dina(n22248), .dinb(n6209), .dout(n25921));
  jand g25689(.dina(n19758), .dinb(n6131), .dout(n25922));
  jand g25690(.dina(n19510), .dinb(n5691), .dout(n25923));
  jor  g25691(.dina(n25923), .dinb(n25922), .dout(n25924));
  jor  g25692(.dina(n25924), .dinb(n25921), .dout(n25925));
  jor  g25693(.dina(n25925), .dinb(n25920), .dout(n25926));
  jxor g25694(.dina(n25926), .dinb(n4247), .dout(n25927));
  jxor g25695(.dina(n25927), .dinb(n25919), .dout(n25928));
  jxor g25696(.dina(n25928), .dinb(n25843), .dout(n25929));
  jand g25697(.dina(n22605), .dinb(n6340), .dout(n25930));
  jand g25698(.dina(n22603), .dinb(n6798), .dout(n25931));
  jand g25699(.dina(n22539), .dinb(n6556), .dout(n25932));
  jand g25700(.dina(n22540), .dinb(n6338), .dout(n25933));
  jor  g25701(.dina(n25933), .dinb(n25932), .dout(n25934));
  jor  g25702(.dina(n25934), .dinb(n25931), .dout(n25935));
  jor  g25703(.dina(n25935), .dinb(n25930), .dout(n25936));
  jxor g25704(.dina(n25936), .dinb(n5064), .dout(n25937));
  jxor g25705(.dina(n25937), .dinb(n25929), .dout(n25938));
  jxor g25706(.dina(n25938), .dinb(n25839), .dout(n25939));
  jxor g25707(.dina(n25939), .dinb(n25836), .dout(n25940));
  jxor g25708(.dina(n25940), .dinb(n25827), .dout(n25941));
  jor  g25709(.dina(n24337), .dinb(n7891), .dout(n25942));
  jor  g25710(.dina(n24335), .dinb(n8440), .dout(n25943));
  jor  g25711(.dina(n24142), .dinb(n8155), .dout(n25944));
  jor  g25712(.dina(n23921), .dinb(n7889), .dout(n25945));
  jand g25713(.dina(n25945), .dinb(n25944), .dout(n25946));
  jand g25714(.dina(n25946), .dinb(n25943), .dout(n25947));
  jand g25715(.dina(n25947), .dinb(n25942), .dout(n25948));
  jxor g25716(.dina(n25948), .dinb(\a[11] ), .dout(n25949));
  jxor g25717(.dina(n25949), .dinb(n25941), .dout(n25950));
  jxor g25718(.dina(n25950), .dinb(n25823), .dout(n25951));
  jxor g25719(.dina(n25951), .dinb(n25820), .dout(n25952));
  jxor g25720(.dina(n25952), .dinb(n25817), .dout(\result[14] ));
  jand g25721(.dina(n25952), .dinb(n25817), .dout(n25954));
  jand g25722(.dina(n25938), .dinb(n25839), .dout(n25955));
  jand g25723(.dina(n25939), .dinb(n25836), .dout(n25956));
  jor  g25724(.dina(n25956), .dinb(n25955), .dout(n25957));
  jor  g25725(.dina(n24357), .dinb(n7891), .dout(n25958));
  jor  g25726(.dina(n24335), .dinb(n14975), .dout(n25959));
  jor  g25727(.dina(n24142), .dinb(n7889), .dout(n25960));
  jand g25728(.dina(n25960), .dinb(n25959), .dout(n25961));
  jand g25729(.dina(n25961), .dinb(n25958), .dout(n25962));
  jxor g25730(.dina(n25962), .dinb(\a[11] ), .dout(n25963));
  jnot g25731(.din(n25963), .dout(n25964));
  jxor g25732(.dina(n25964), .dinb(n25957), .dout(n25965));
  jand g25733(.dina(n25884), .dinb(n25880), .dout(n25966));
  jnot g25734(.din(n25966), .dout(n25967));
  jor  g25735(.dina(n25894), .dinb(n25886), .dout(n25968));
  jand g25736(.dina(n25968), .dinb(n25967), .dout(n25969));
  jnot g25737(.din(n25969), .dout(n25970));
  jand g25738(.dina(n21086), .dinb(n4449), .dout(n25971));
  jand g25739(.dina(n19521), .dinb(n4453), .dout(n25972));
  jand g25740(.dina(n19523), .dinb(n4457), .dout(n25973));
  jand g25741(.dina(n19525), .dinb(n4461), .dout(n25974));
  jor  g25742(.dina(n25974), .dinb(n25973), .dout(n25975));
  jor  g25743(.dina(n25975), .dinb(n25972), .dout(n25976));
  jor  g25744(.dina(n25976), .dinb(n25971), .dout(n25977));
  jxor g25745(.dina(n25977), .dinb(n88), .dout(n25978));
  jnot g25746(.din(n25978), .dout(n25979));
  jand g25747(.dina(n612), .dinb(n517), .dout(n25980));
  jand g25748(.dina(n25980), .dinb(n950), .dout(n25981));
  jand g25749(.dina(n1829), .dinb(n1578), .dout(n25982));
  jand g25750(.dina(n25982), .dinb(n25981), .dout(n25983));
  jand g25751(.dina(n25983), .dinb(n3589), .dout(n25984));
  jand g25752(.dina(n1899), .dinb(n1019), .dout(n25985));
  jand g25753(.dina(n1663), .dinb(n198), .dout(n25986));
  jand g25754(.dina(n25986), .dinb(n25985), .dout(n25987));
  jand g25755(.dina(n4796), .dinb(n601), .dout(n25988));
  jand g25756(.dina(n1185), .dinb(n752), .dout(n25989));
  jand g25757(.dina(n25989), .dinb(n25988), .dout(n25990));
  jand g25758(.dina(n25990), .dinb(n25987), .dout(n25991));
  jand g25759(.dina(n25991), .dinb(n25984), .dout(n25992));
  jand g25760(.dina(n13867), .dinb(n12228), .dout(n25993));
  jand g25761(.dina(n25993), .dinb(n25992), .dout(n25994));
  jand g25762(.dina(n25994), .dinb(n25334), .dout(n25995));
  jand g25763(.dina(n25995), .dinb(n6004), .dout(n25996));
  jxor g25764(.dina(n25996), .dinb(n25871), .dout(n25997));
  jand g25765(.dina(n25871), .dinb(n25857), .dout(n25998));
  jnot g25766(.din(n25998), .dout(n25999));
  jnot g25767(.din(n25857), .dout(n26000));
  jand g25768(.dina(n25870), .dinb(n26000), .dout(n26001));
  jor  g25769(.dina(n25879), .dinb(n26001), .dout(n26002));
  jand g25770(.dina(n26002), .dinb(n25999), .dout(n26003));
  jxor g25771(.dina(n26003), .dinb(n25997), .dout(n26004));
  jand g25772(.dina(n20793), .dinb(n732), .dout(n26005));
  jand g25773(.dina(n19527), .dinb(n3855), .dout(n26006));
  jand g25774(.dina(n19529), .dinb(n3858), .dout(n26007));
  jand g25775(.dina(n19531), .dinb(n3851), .dout(n26008));
  jor  g25776(.dina(n26008), .dinb(n26007), .dout(n26009));
  jor  g25777(.dina(n26009), .dinb(n26006), .dout(n26010));
  jor  g25778(.dina(n26010), .dinb(n26005), .dout(n26011));
  jxor g25779(.dina(n26011), .dinb(n26004), .dout(n26012));
  jxor g25780(.dina(n26012), .dinb(n25979), .dout(n26013));
  jxor g25781(.dina(n26013), .dinb(n25970), .dout(n26014));
  jand g25782(.dina(n21218), .dinb(n75), .dout(n26015));
  jand g25783(.dina(n19515), .dinb(n4933), .dout(n26016));
  jand g25784(.dina(n19517), .dinb(n4918), .dout(n26017));
  jand g25785(.dina(n19519), .dinb(n4745), .dout(n26018));
  jor  g25786(.dina(n26018), .dinb(n26017), .dout(n26019));
  jor  g25787(.dina(n26019), .dinb(n26016), .dout(n26020));
  jor  g25788(.dina(n26020), .dinb(n26015), .dout(n26021));
  jxor g25789(.dina(n26021), .dinb(n68), .dout(n26022));
  jnot g25790(.din(n26022), .dout(n26023));
  jxor g25791(.dina(n26023), .dinb(n26014), .dout(n26024));
  jor  g25792(.dina(n25895), .dinb(n25853), .dout(n26025));
  jand g25793(.dina(n25895), .dinb(n25853), .dout(n26026));
  jor  g25794(.dina(n25905), .dinb(n26026), .dout(n26027));
  jand g25795(.dina(n26027), .dinb(n26025), .dout(n26028));
  jxor g25796(.dina(n26028), .dinb(n26024), .dout(n26029));
  jand g25797(.dina(n21750), .dinb(n5365), .dout(n26030));
  jand g25798(.dina(n19510), .dinb(n5500), .dout(n26031));
  jand g25799(.dina(n19511), .dinb(n5424), .dout(n26032));
  jand g25800(.dina(n19513), .dinb(n5363), .dout(n26033));
  jor  g25801(.dina(n26033), .dinb(n26032), .dout(n26034));
  jor  g25802(.dina(n26034), .dinb(n26031), .dout(n26035));
  jor  g25803(.dina(n26035), .dinb(n26030), .dout(n26036));
  jxor g25804(.dina(n26036), .dinb(n72), .dout(n26037));
  jnot g25805(.din(n26037), .dout(n26038));
  jxor g25806(.dina(n26038), .dinb(n26029), .dout(n26039));
  jand g25807(.dina(n25907), .dinb(n25850), .dout(n26040));
  jnot g25808(.din(n26040), .dout(n26041));
  jnot g25809(.din(n25850), .dout(n26042));
  jand g25810(.dina(n25906), .dinb(n26042), .dout(n26043));
  jor  g25811(.dina(n25917), .dinb(n26043), .dout(n26044));
  jand g25812(.dina(n26044), .dinb(n26041), .dout(n26045));
  jxor g25813(.dina(n26045), .dinb(n26039), .dout(n26046));
  jand g25814(.dina(n22627), .dinb(n5693), .dout(n26047));
  jand g25815(.dina(n22540), .dinb(n6209), .dout(n26048));
  jand g25816(.dina(n22248), .dinb(n6131), .dout(n26049));
  jand g25817(.dina(n19758), .dinb(n5691), .dout(n26050));
  jor  g25818(.dina(n26050), .dinb(n26049), .dout(n26051));
  jor  g25819(.dina(n26051), .dinb(n26048), .dout(n26052));
  jor  g25820(.dina(n26052), .dinb(n26047), .dout(n26053));
  jxor g25821(.dina(n26053), .dinb(n4247), .dout(n26054));
  jnot g25822(.din(n26054), .dout(n26055));
  jxor g25823(.dina(n26055), .dinb(n26046), .dout(n26056));
  jnot g25824(.din(n26056), .dout(n26057));
  jnot g25825(.din(n25918), .dout(n26058));
  jand g25826(.dina(n26058), .dinb(n25847), .dout(n26059));
  jnot g25827(.din(n25847), .dout(n26060));
  jand g25828(.dina(n25918), .dinb(n26060), .dout(n26061));
  jnot g25829(.din(n26061), .dout(n26062));
  jand g25830(.dina(n25927), .dinb(n26062), .dout(n26063));
  jor  g25831(.dina(n26063), .dinb(n26059), .dout(n26064));
  jxor g25832(.dina(n26064), .dinb(n26057), .dout(n26065));
  jand g25833(.dina(n23262), .dinb(n6340), .dout(n26066));
  jand g25834(.dina(n23260), .dinb(n6798), .dout(n26067));
  jand g25835(.dina(n22603), .dinb(n6556), .dout(n26068));
  jand g25836(.dina(n22539), .dinb(n6338), .dout(n26069));
  jor  g25837(.dina(n26069), .dinb(n26068), .dout(n26070));
  jor  g25838(.dina(n26070), .dinb(n26067), .dout(n26071));
  jor  g25839(.dina(n26071), .dinb(n26066), .dout(n26072));
  jxor g25840(.dina(n26072), .dinb(n5064), .dout(n26073));
  jnot g25841(.din(n26073), .dout(n26074));
  jxor g25842(.dina(n26074), .dinb(n26065), .dout(n26075));
  jnot g25843(.din(n25928), .dout(n26076));
  jand g25844(.dina(n26076), .dinb(n25843), .dout(n26077));
  jnot g25845(.din(n25843), .dout(n26078));
  jand g25846(.dina(n25928), .dinb(n26078), .dout(n26079));
  jnot g25847(.din(n26079), .dout(n26080));
  jand g25848(.dina(n25937), .dinb(n26080), .dout(n26081));
  jor  g25849(.dina(n26081), .dinb(n26077), .dout(n26082));
  jxor g25850(.dina(n26082), .dinb(n26075), .dout(n26083));
  jor  g25851(.dina(n23919), .dinb(n6937), .dout(n26084));
  jor  g25852(.dina(n23921), .dinb(n7740), .dout(n26085));
  jor  g25853(.dina(n23710), .dinb(n7614), .dout(n26086));
  jor  g25854(.dina(n23496), .dinb(n6935), .dout(n26087));
  jand g25855(.dina(n26087), .dinb(n26086), .dout(n26088));
  jand g25856(.dina(n26088), .dinb(n26085), .dout(n26089));
  jand g25857(.dina(n26089), .dinb(n26084), .dout(n26090));
  jxor g25858(.dina(n26090), .dinb(\a[14] ), .dout(n26091));
  jxor g25859(.dina(n26091), .dinb(n26083), .dout(n26092));
  jxor g25860(.dina(n26092), .dinb(n25965), .dout(n26093));
  jnot g25861(.din(n25940), .dout(n26094));
  jand g25862(.dina(n26094), .dinb(n25827), .dout(n26095));
  jnot g25863(.din(n26095), .dout(n26096));
  jnot g25864(.din(n25827), .dout(n26097));
  jand g25865(.dina(n25940), .dinb(n26097), .dout(n26098));
  jnot g25866(.din(n25949), .dout(n26099));
  jor  g25867(.dina(n26099), .dinb(n26098), .dout(n26100));
  jand g25868(.dina(n26100), .dinb(n26096), .dout(n26101));
  jxor g25869(.dina(n26101), .dinb(n26093), .dout(n26102));
  jand g25870(.dina(n25950), .dinb(n25823), .dout(n26103));
  jand g25871(.dina(n25951), .dinb(n25820), .dout(n26104));
  jor  g25872(.dina(n26104), .dinb(n26103), .dout(n26105));
  jxor g25873(.dina(n26105), .dinb(n26102), .dout(n26106));
  jxor g25874(.dina(n26106), .dinb(n25954), .dout(\result[15] ));
  jand g25875(.dina(n26106), .dinb(n25954), .dout(n26108));
  jand g25876(.dina(n26101), .dinb(n26093), .dout(n26109));
  jand g25877(.dina(n26105), .dinb(n26102), .dout(n26110));
  jor  g25878(.dina(n26110), .dinb(n26109), .dout(n26111));
  jand g25879(.dina(n21738), .dinb(n75), .dout(n26112));
  jand g25880(.dina(n19513), .dinb(n4933), .dout(n26113));
  jand g25881(.dina(n19515), .dinb(n4918), .dout(n26114));
  jand g25882(.dina(n19517), .dinb(n4745), .dout(n26115));
  jor  g25883(.dina(n26115), .dinb(n26114), .dout(n26116));
  jor  g25884(.dina(n26116), .dinb(n26113), .dout(n26117));
  jor  g25885(.dina(n26117), .dinb(n26112), .dout(n26118));
  jxor g25886(.dina(n26118), .dinb(n68), .dout(n26119));
  jnot g25887(.din(n26119), .dout(n26120));
  jand g25888(.dina(n21240), .dinb(n4449), .dout(n26121));
  jand g25889(.dina(n19519), .dinb(n4453), .dout(n26122));
  jand g25890(.dina(n19521), .dinb(n4457), .dout(n26123));
  jand g25891(.dina(n19523), .dinb(n4461), .dout(n26124));
  jor  g25892(.dina(n26124), .dinb(n26123), .dout(n26125));
  jor  g25893(.dina(n26125), .dinb(n26122), .dout(n26126));
  jor  g25894(.dina(n26126), .dinb(n26121), .dout(n26127));
  jxor g25895(.dina(n26127), .dinb(n88), .dout(n26128));
  jnot g25896(.din(n26128), .dout(n26129));
  jand g25897(.dina(n26011), .dinb(n26004), .dout(n26130));
  jand g25898(.dina(n26012), .dinb(n25979), .dout(n26131));
  jor  g25899(.dina(n26131), .dinb(n26130), .dout(n26132));
  jor  g25900(.dina(n25996), .dinb(n25871), .dout(n26133));
  jand g25901(.dina(n26003), .dinb(n25997), .dout(n26134));
  jnot g25902(.din(n26134), .dout(n26135));
  jand g25903(.dina(n26135), .dinb(n26133), .dout(n26136));
  jnot g25904(.din(n26136), .dout(n26137));
  jand g25905(.dina(n24593), .dinb(n13107), .dout(n26138));
  jxor g25906(.dina(n26138), .dinb(n5833), .dout(n26139));
  jand g25907(.dina(n366), .dinb(n314), .dout(n26140));
  jand g25908(.dina(n703), .dinb(n439), .dout(n26141));
  jand g25909(.dina(n26141), .dinb(n26140), .dout(n26142));
  jand g25910(.dina(n1569), .dinb(n218), .dout(n26143));
  jand g25911(.dina(n26143), .dinb(n26142), .dout(n26144));
  jand g25912(.dina(n12967), .dinb(n5736), .dout(n26145));
  jand g25913(.dina(n26145), .dinb(n26144), .dout(n26146));
  jand g25914(.dina(n3594), .dinb(n1135), .dout(n26147));
  jand g25915(.dina(n26147), .dinb(n4287), .dout(n26148));
  jand g25916(.dina(n26148), .dinb(n2985), .dout(n26149));
  jand g25917(.dina(n26149), .dinb(n5759), .dout(n26150));
  jand g25918(.dina(n26150), .dinb(n26146), .dout(n26151));
  jand g25919(.dina(n26151), .dinb(n2249), .dout(n26152));
  jand g25920(.dina(n2298), .dinb(n1116), .dout(n26153));
  jand g25921(.dina(n26153), .dinb(n26152), .dout(n26154));
  jxor g25922(.dina(n26154), .dinb(n25870), .dout(n26155));
  jxor g25923(.dina(n26155), .dinb(n26139), .dout(n26156));
  jand g25924(.dina(n20781), .dinb(n732), .dout(n26157));
  jand g25925(.dina(n19525), .dinb(n3855), .dout(n26158));
  jand g25926(.dina(n19527), .dinb(n3858), .dout(n26159));
  jand g25927(.dina(n19529), .dinb(n3851), .dout(n26160));
  jor  g25928(.dina(n26160), .dinb(n26159), .dout(n26161));
  jor  g25929(.dina(n26161), .dinb(n26158), .dout(n26162));
  jor  g25930(.dina(n26162), .dinb(n26157), .dout(n26163));
  jxor g25931(.dina(n26163), .dinb(n26156), .dout(n26164));
  jxor g25932(.dina(n26164), .dinb(n26137), .dout(n26165));
  jxor g25933(.dina(n26165), .dinb(n26132), .dout(n26166));
  jxor g25934(.dina(n26166), .dinb(n26129), .dout(n26167));
  jxor g25935(.dina(n26167), .dinb(n26120), .dout(n26168));
  jor  g25936(.dina(n26013), .dinb(n25970), .dout(n26169));
  jand g25937(.dina(n26013), .dinb(n25970), .dout(n26170));
  jor  g25938(.dina(n26023), .dinb(n26170), .dout(n26171));
  jand g25939(.dina(n26171), .dinb(n26169), .dout(n26172));
  jxor g25940(.dina(n26172), .dinb(n26168), .dout(n26173));
  jnot g25941(.din(n26173), .dout(n26174));
  jand g25942(.dina(n19760), .dinb(n5365), .dout(n26175));
  jand g25943(.dina(n19758), .dinb(n5500), .dout(n26176));
  jand g25944(.dina(n19510), .dinb(n5424), .dout(n26177));
  jand g25945(.dina(n19511), .dinb(n5363), .dout(n26178));
  jor  g25946(.dina(n26178), .dinb(n26177), .dout(n26179));
  jor  g25947(.dina(n26179), .dinb(n26176), .dout(n26180));
  jor  g25948(.dina(n26180), .dinb(n26175), .dout(n26181));
  jxor g25949(.dina(n26181), .dinb(n72), .dout(n26182));
  jxor g25950(.dina(n26182), .dinb(n26174), .dout(n26183));
  jnot g25951(.din(n26024), .dout(n26184));
  jnot g25952(.din(n26028), .dout(n26185));
  jand g25953(.dina(n26185), .dinb(n26184), .dout(n26186));
  jnot g25954(.din(n26186), .dout(n26187));
  jand g25955(.dina(n26028), .dinb(n26024), .dout(n26188));
  jor  g25956(.dina(n26038), .dinb(n26188), .dout(n26189));
  jand g25957(.dina(n26189), .dinb(n26187), .dout(n26190));
  jxor g25958(.dina(n26190), .dinb(n26183), .dout(n26191));
  jand g25959(.dina(n22617), .dinb(n5693), .dout(n26192));
  jand g25960(.dina(n22539), .dinb(n6209), .dout(n26193));
  jand g25961(.dina(n22540), .dinb(n6131), .dout(n26194));
  jand g25962(.dina(n22248), .dinb(n5691), .dout(n26195));
  jor  g25963(.dina(n26195), .dinb(n26194), .dout(n26196));
  jor  g25964(.dina(n26196), .dinb(n26193), .dout(n26197));
  jor  g25965(.dina(n26197), .dinb(n26192), .dout(n26198));
  jxor g25966(.dina(n26198), .dinb(n4247), .dout(n26199));
  jnot g25967(.din(n26199), .dout(n26200));
  jnot g25968(.din(n26039), .dout(n26201));
  jnot g25969(.din(n26045), .dout(n26202));
  jand g25970(.dina(n26202), .dinb(n26201), .dout(n26203));
  jnot g25971(.din(n26203), .dout(n26204));
  jand g25972(.dina(n26045), .dinb(n26039), .dout(n26205));
  jor  g25973(.dina(n26055), .dinb(n26205), .dout(n26206));
  jand g25974(.dina(n26206), .dinb(n26204), .dout(n26207));
  jxor g25975(.dina(n26207), .dinb(n26200), .dout(n26208));
  jxor g25976(.dina(n26208), .dinb(n26191), .dout(n26209));
  jnot g25977(.din(n26209), .dout(n26210));
  jor  g25978(.dina(n23494), .dinb(n6341), .dout(n26211));
  jor  g25979(.dina(n23496), .dinb(n6797), .dout(n26212));
  jor  g25980(.dina(n23450), .dinb(n6557), .dout(n26213));
  jor  g25981(.dina(n23449), .dinb(n6339), .dout(n26214));
  jand g25982(.dina(n26214), .dinb(n26213), .dout(n26215));
  jand g25983(.dina(n26215), .dinb(n26212), .dout(n26216));
  jand g25984(.dina(n26216), .dinb(n26211), .dout(n26217));
  jxor g25985(.dina(n26217), .dinb(\a[17] ), .dout(n26218));
  jxor g25986(.dina(n26218), .dinb(n26210), .dout(n26219));
  jand g25987(.dina(n26064), .dinb(n26057), .dout(n26220));
  jnot g25988(.din(n26220), .dout(n26221));
  jnot g25989(.din(n26064), .dout(n26222));
  jand g25990(.dina(n26222), .dinb(n26056), .dout(n26223));
  jor  g25991(.dina(n26074), .dinb(n26223), .dout(n26224));
  jand g25992(.dina(n26224), .dinb(n26221), .dout(n26225));
  jxor g25993(.dina(n26225), .dinb(n26219), .dout(n26226));
  jor  g25994(.dina(n24140), .dinb(n6937), .dout(n26227));
  jor  g25995(.dina(n24142), .dinb(n7740), .dout(n26228));
  jor  g25996(.dina(n23921), .dinb(n7614), .dout(n26229));
  jor  g25997(.dina(n23710), .dinb(n6935), .dout(n26230));
  jand g25998(.dina(n26230), .dinb(n26229), .dout(n26231));
  jand g25999(.dina(n26231), .dinb(n26228), .dout(n26232));
  jand g26000(.dina(n26232), .dinb(n26227), .dout(n26233));
  jxor g26001(.dina(n26233), .dinb(\a[14] ), .dout(n26234));
  jnot g26002(.din(n26234), .dout(n26235));
  jnot g26003(.din(n26075), .dout(n26236));
  jand g26004(.dina(n26082), .dinb(n26236), .dout(n26237));
  jnot g26005(.din(n26237), .dout(n26238));
  jnot g26006(.din(n26082), .dout(n26239));
  jand g26007(.dina(n26239), .dinb(n26075), .dout(n26240));
  jnot g26008(.din(n26091), .dout(n26241));
  jor  g26009(.dina(n26241), .dinb(n26240), .dout(n26242));
  jand g26010(.dina(n26242), .dinb(n26238), .dout(n26243));
  jxor g26011(.dina(n26243), .dinb(n26235), .dout(n26244));
  jxor g26012(.dina(n26244), .dinb(n26226), .dout(n26245));
  jnot g26013(.din(n25957), .dout(n26246));
  jand g26014(.dina(n25963), .dinb(n26246), .dout(n26247));
  jnot g26015(.din(n26247), .dout(n26248));
  jand g26016(.dina(n25964), .dinb(n25957), .dout(n26249));
  jor  g26017(.dina(n26092), .dinb(n26249), .dout(n26250));
  jand g26018(.dina(n26250), .dinb(n26248), .dout(n26251));
  jxor g26019(.dina(n26251), .dinb(n26245), .dout(n26252));
  jxor g26020(.dina(n26252), .dinb(n26111), .dout(n26253));
  jxor g26021(.dina(n26253), .dinb(n26108), .dout(\result[16] ));
  jand g26022(.dina(n26253), .dinb(n26108), .dout(n26255));
  jand g26023(.dina(n26251), .dinb(n26245), .dout(n26256));
  jand g26024(.dina(n26252), .dinb(n26111), .dout(n26257));
  jor  g26025(.dina(n26257), .dinb(n26256), .dout(n26258));
  jand g26026(.dina(n26243), .dinb(n26235), .dout(n26259));
  jand g26027(.dina(n26244), .dinb(n26226), .dout(n26260));
  jor  g26028(.dina(n26260), .dinb(n26259), .dout(n26261));
  jor  g26029(.dina(n26218), .dinb(n26210), .dout(n26262));
  jand g26030(.dina(n26225), .dinb(n26219), .dout(n26263));
  jnot g26031(.din(n26263), .dout(n26264));
  jand g26032(.dina(n26264), .dinb(n26262), .dout(n26265));
  jor  g26033(.dina(n23708), .dinb(n6341), .dout(n26266));
  jor  g26034(.dina(n23710), .dinb(n6797), .dout(n26267));
  jor  g26035(.dina(n23496), .dinb(n6557), .dout(n26268));
  jor  g26036(.dina(n23450), .dinb(n6339), .dout(n26269));
  jand g26037(.dina(n26269), .dinb(n26268), .dout(n26270));
  jand g26038(.dina(n26270), .dinb(n26267), .dout(n26271));
  jand g26039(.dina(n26271), .dinb(n26266), .dout(n26272));
  jxor g26040(.dina(n26272), .dinb(\a[17] ), .dout(n26273));
  jnot g26041(.din(n26273), .dout(n26274));
  jand g26042(.dina(n26207), .dinb(n26200), .dout(n26275));
  jand g26043(.dina(n26208), .dinb(n26191), .dout(n26276));
  jor  g26044(.dina(n26276), .dinb(n26275), .dout(n26277));
  jor  g26045(.dina(n26182), .dinb(n26174), .dout(n26278));
  jand g26046(.dina(n26190), .dinb(n26183), .dout(n26279));
  jnot g26047(.din(n26279), .dout(n26280));
  jand g26048(.dina(n26280), .dinb(n26278), .dout(n26281));
  jand g26049(.dina(n26167), .dinb(n26120), .dout(n26282));
  jand g26050(.dina(n26172), .dinb(n26168), .dout(n26283));
  jor  g26051(.dina(n26283), .dinb(n26282), .dout(n26284));
  jand g26052(.dina(n26163), .dinb(n26156), .dout(n26285));
  jand g26053(.dina(n26164), .dinb(n26137), .dout(n26286));
  jor  g26054(.dina(n26286), .dinb(n26285), .dout(n26287));
  jor  g26055(.dina(n26154), .dinb(n25870), .dout(n26288));
  jand g26056(.dina(n26155), .dinb(n26139), .dout(n26289));
  jnot g26057(.din(n26289), .dout(n26290));
  jand g26058(.dina(n26290), .dinb(n26288), .dout(n26291));
  jand g26059(.dina(n988), .dinb(n270), .dout(n26292));
  jand g26060(.dina(n26292), .dinb(n696), .dout(n26293));
  jand g26061(.dina(n2525), .dinb(n868), .dout(n26294));
  jand g26062(.dina(n26294), .dinb(n26293), .dout(n26295));
  jand g26063(.dina(n4101), .dinb(n2368), .dout(n26296));
  jand g26064(.dina(n26296), .dinb(n26295), .dout(n26297));
  jand g26065(.dina(n2940), .dinb(n2292), .dout(n26298));
  jand g26066(.dina(n26298), .dinb(n995), .dout(n26299));
  jand g26067(.dina(n26299), .dinb(n12863), .dout(n26300));
  jand g26068(.dina(n26300), .dinb(n26297), .dout(n26301));
  jand g26069(.dina(n24453), .dinb(n24039), .dout(n26302));
  jand g26070(.dina(n26302), .dinb(n26301), .dout(n26303));
  jand g26071(.dina(n26303), .dinb(n13869), .dout(n26304));
  jand g26072(.dina(n26304), .dinb(n12975), .dout(n26305));
  jnot g26073(.din(n26305), .dout(n26306));
  jxor g26074(.dina(n26306), .dinb(n26291), .dout(n26307));
  jand g26075(.dina(n19770), .dinb(n732), .dout(n26308));
  jand g26076(.dina(n19523), .dinb(n3855), .dout(n26309));
  jand g26077(.dina(n19525), .dinb(n3858), .dout(n26310));
  jand g26078(.dina(n19527), .dinb(n3851), .dout(n26311));
  jor  g26079(.dina(n26311), .dinb(n26310), .dout(n26312));
  jor  g26080(.dina(n26312), .dinb(n26309), .dout(n26313));
  jor  g26081(.dina(n26313), .dinb(n26308), .dout(n26314));
  jxor g26082(.dina(n26314), .dinb(n26307), .dout(n26315));
  jxor g26083(.dina(n26315), .dinb(n26287), .dout(n26316));
  jnot g26084(.din(n26316), .dout(n26317));
  jand g26085(.dina(n21230), .dinb(n4449), .dout(n26318));
  jand g26086(.dina(n19517), .dinb(n4453), .dout(n26319));
  jand g26087(.dina(n19519), .dinb(n4457), .dout(n26320));
  jand g26088(.dina(n19521), .dinb(n4461), .dout(n26321));
  jor  g26089(.dina(n26321), .dinb(n26320), .dout(n26322));
  jor  g26090(.dina(n26322), .dinb(n26319), .dout(n26323));
  jor  g26091(.dina(n26323), .dinb(n26318), .dout(n26324));
  jxor g26092(.dina(n26324), .dinb(n88), .dout(n26325));
  jxor g26093(.dina(n26325), .dinb(n26317), .dout(n26326));
  jor  g26094(.dina(n26165), .dinb(n26132), .dout(n26327));
  jand g26095(.dina(n26165), .dinb(n26132), .dout(n26328));
  jor  g26096(.dina(n26328), .dinb(n26129), .dout(n26329));
  jand g26097(.dina(n26329), .dinb(n26327), .dout(n26330));
  jxor g26098(.dina(n26330), .dinb(n26326), .dout(n26331));
  jand g26099(.dina(n21762), .dinb(n75), .dout(n26332));
  jand g26100(.dina(n19511), .dinb(n4933), .dout(n26333));
  jand g26101(.dina(n19513), .dinb(n4918), .dout(n26334));
  jand g26102(.dina(n19515), .dinb(n4745), .dout(n26335));
  jor  g26103(.dina(n26335), .dinb(n26334), .dout(n26336));
  jor  g26104(.dina(n26336), .dinb(n26333), .dout(n26337));
  jor  g26105(.dina(n26337), .dinb(n26332), .dout(n26338));
  jxor g26106(.dina(n26338), .dinb(n68), .dout(n26339));
  jnot g26107(.din(n26339), .dout(n26340));
  jxor g26108(.dina(n26340), .dinb(n26331), .dout(n26341));
  jxor g26109(.dina(n26341), .dinb(n26284), .dout(n26342));
  jand g26110(.dina(n22250), .dinb(n5365), .dout(n26343));
  jand g26111(.dina(n22248), .dinb(n5500), .dout(n26344));
  jand g26112(.dina(n19758), .dinb(n5424), .dout(n26345));
  jand g26113(.dina(n19510), .dinb(n5363), .dout(n26346));
  jor  g26114(.dina(n26346), .dinb(n26345), .dout(n26347));
  jor  g26115(.dina(n26347), .dinb(n26344), .dout(n26348));
  jor  g26116(.dina(n26348), .dinb(n26343), .dout(n26349));
  jxor g26117(.dina(n26349), .dinb(n72), .dout(n26350));
  jnot g26118(.din(n26350), .dout(n26351));
  jxor g26119(.dina(n26351), .dinb(n26342), .dout(n26352));
  jnot g26120(.din(n26352), .dout(n26353));
  jxor g26121(.dina(n26353), .dinb(n26281), .dout(n26354));
  jand g26122(.dina(n22605), .dinb(n5693), .dout(n26355));
  jand g26123(.dina(n22603), .dinb(n6209), .dout(n26356));
  jand g26124(.dina(n22539), .dinb(n6131), .dout(n26357));
  jand g26125(.dina(n22540), .dinb(n5691), .dout(n26358));
  jor  g26126(.dina(n26358), .dinb(n26357), .dout(n26359));
  jor  g26127(.dina(n26359), .dinb(n26356), .dout(n26360));
  jor  g26128(.dina(n26360), .dinb(n26355), .dout(n26361));
  jxor g26129(.dina(n26361), .dinb(n4247), .dout(n26362));
  jnot g26130(.din(n26362), .dout(n26363));
  jxor g26131(.dina(n26363), .dinb(n26354), .dout(n26364));
  jxor g26132(.dina(n26364), .dinb(n26277), .dout(n26365));
  jxor g26133(.dina(n26365), .dinb(n26274), .dout(n26366));
  jxor g26134(.dina(n26366), .dinb(n26265), .dout(n26367));
  jor  g26135(.dina(n24337), .dinb(n6937), .dout(n26368));
  jor  g26136(.dina(n24335), .dinb(n7740), .dout(n26369));
  jor  g26137(.dina(n24142), .dinb(n7614), .dout(n26370));
  jor  g26138(.dina(n23921), .dinb(n6935), .dout(n26371));
  jand g26139(.dina(n26371), .dinb(n26370), .dout(n26372));
  jand g26140(.dina(n26372), .dinb(n26369), .dout(n26373));
  jand g26141(.dina(n26373), .dinb(n26368), .dout(n26374));
  jxor g26142(.dina(n26374), .dinb(\a[14] ), .dout(n26375));
  jxor g26143(.dina(n26375), .dinb(n26367), .dout(n26376));
  jxor g26144(.dina(n26376), .dinb(n26261), .dout(n26377));
  jxor g26145(.dina(n26377), .dinb(n26258), .dout(n26378));
  jxor g26146(.dina(n26378), .dinb(n26255), .dout(\result[17] ));
  jand g26147(.dina(n26378), .dinb(n26255), .dout(n26380));
  jand g26148(.dina(n26364), .dinb(n26277), .dout(n26381));
  jand g26149(.dina(n26365), .dinb(n26274), .dout(n26382));
  jor  g26150(.dina(n26382), .dinb(n26381), .dout(n26383));
  jor  g26151(.dina(n24357), .dinb(n6937), .dout(n26384));
  jor  g26152(.dina(n24335), .dinb(n14147), .dout(n26385));
  jor  g26153(.dina(n24142), .dinb(n6935), .dout(n26386));
  jand g26154(.dina(n26386), .dinb(n26385), .dout(n26387));
  jand g26155(.dina(n26387), .dinb(n26384), .dout(n26388));
  jxor g26156(.dina(n26388), .dinb(\a[14] ), .dout(n26389));
  jnot g26157(.din(n26389), .dout(n26390));
  jxor g26158(.dina(n26390), .dinb(n26383), .dout(n26391));
  jand g26159(.dina(n21750), .dinb(n75), .dout(n26392));
  jand g26160(.dina(n19510), .dinb(n4933), .dout(n26393));
  jand g26161(.dina(n19511), .dinb(n4918), .dout(n26394));
  jand g26162(.dina(n19513), .dinb(n4745), .dout(n26395));
  jor  g26163(.dina(n26395), .dinb(n26394), .dout(n26396));
  jor  g26164(.dina(n26396), .dinb(n26393), .dout(n26397));
  jor  g26165(.dina(n26397), .dinb(n26392), .dout(n26398));
  jxor g26166(.dina(n26398), .dinb(n68), .dout(n26399));
  jnot g26167(.din(n26399), .dout(n26400));
  jand g26168(.dina(n12132), .dinb(n5952), .dout(n26401));
  jand g26169(.dina(n26401), .dinb(n744), .dout(n26402));
  jand g26170(.dina(n3550), .dinb(n1600), .dout(n26403));
  jand g26171(.dina(n26403), .dinb(n722), .dout(n26404));
  jand g26172(.dina(n113), .dinb(n108), .dout(n26405));
  jand g26173(.dina(n1066), .dinb(n988), .dout(n26406));
  jand g26174(.dina(n26406), .dinb(n26405), .dout(n26407));
  jand g26175(.dina(n1047), .dinb(n619), .dout(n26408));
  jand g26176(.dina(n26408), .dinb(n7004), .dout(n26409));
  jand g26177(.dina(n26409), .dinb(n26407), .dout(n26410));
  jand g26178(.dina(n26410), .dinb(n26404), .dout(n26411));
  jand g26179(.dina(n2983), .dinb(n421), .dout(n26412));
  jand g26180(.dina(n26412), .dinb(n26411), .dout(n26413));
  jand g26181(.dina(n26413), .dinb(n3293), .dout(n26414));
  jand g26182(.dina(n26414), .dinb(n26402), .dout(n26415));
  jand g26183(.dina(n26415), .dinb(n4139), .dout(n26416));
  jxor g26184(.dina(n26416), .dinb(n26306), .dout(n26417));
  jand g26185(.dina(n21086), .dinb(n732), .dout(n26418));
  jand g26186(.dina(n19521), .dinb(n3855), .dout(n26419));
  jand g26187(.dina(n19523), .dinb(n3858), .dout(n26420));
  jand g26188(.dina(n19525), .dinb(n3851), .dout(n26421));
  jor  g26189(.dina(n26421), .dinb(n26420), .dout(n26422));
  jor  g26190(.dina(n26422), .dinb(n26419), .dout(n26423));
  jor  g26191(.dina(n26423), .dinb(n26418), .dout(n26424));
  jxor g26192(.dina(n26424), .dinb(n26417), .dout(n26425));
  jand g26193(.dina(n26306), .dinb(n26291), .dout(n26426));
  jnot g26194(.din(n26426), .dout(n26427));
  jnot g26195(.din(n26291), .dout(n26428));
  jand g26196(.dina(n26305), .dinb(n26428), .dout(n26429));
  jor  g26197(.dina(n26314), .dinb(n26429), .dout(n26430));
  jand g26198(.dina(n26430), .dinb(n26427), .dout(n26431));
  jxor g26199(.dina(n26431), .dinb(n26425), .dout(n26432));
  jnot g26200(.din(n26432), .dout(n26433));
  jand g26201(.dina(n26315), .dinb(n26287), .dout(n26434));
  jnot g26202(.din(n26434), .dout(n26435));
  jor  g26203(.dina(n26325), .dinb(n26317), .dout(n26436));
  jand g26204(.dina(n26436), .dinb(n26435), .dout(n26437));
  jxor g26205(.dina(n26437), .dinb(n26433), .dout(n26438));
  jnot g26206(.din(n26438), .dout(n26439));
  jand g26207(.dina(n21218), .dinb(n4449), .dout(n26440));
  jand g26208(.dina(n19515), .dinb(n4453), .dout(n26441));
  jand g26209(.dina(n19517), .dinb(n4457), .dout(n26442));
  jand g26210(.dina(n19519), .dinb(n4461), .dout(n26443));
  jor  g26211(.dina(n26443), .dinb(n26442), .dout(n26444));
  jor  g26212(.dina(n26444), .dinb(n26441), .dout(n26445));
  jor  g26213(.dina(n26445), .dinb(n26440), .dout(n26446));
  jxor g26214(.dina(n26446), .dinb(n88), .dout(n26447));
  jxor g26215(.dina(n26447), .dinb(n26439), .dout(n26448));
  jxor g26216(.dina(n26448), .dinb(n26400), .dout(n26449));
  jor  g26217(.dina(n26330), .dinb(n26326), .dout(n26450));
  jand g26218(.dina(n26330), .dinb(n26326), .dout(n26451));
  jor  g26219(.dina(n26340), .dinb(n26451), .dout(n26452));
  jand g26220(.dina(n26452), .dinb(n26450), .dout(n26453));
  jxor g26221(.dina(n26453), .dinb(n26449), .dout(n26454));
  jand g26222(.dina(n22627), .dinb(n5365), .dout(n26455));
  jand g26223(.dina(n22540), .dinb(n5500), .dout(n26456));
  jand g26224(.dina(n22248), .dinb(n5424), .dout(n26457));
  jand g26225(.dina(n19758), .dinb(n5363), .dout(n26458));
  jor  g26226(.dina(n26458), .dinb(n26457), .dout(n26459));
  jor  g26227(.dina(n26459), .dinb(n26456), .dout(n26460));
  jor  g26228(.dina(n26460), .dinb(n26455), .dout(n26461));
  jxor g26229(.dina(n26461), .dinb(n72), .dout(n26462));
  jnot g26230(.din(n26462), .dout(n26463));
  jxor g26231(.dina(n26463), .dinb(n26454), .dout(n26464));
  jnot g26232(.din(n26284), .dout(n26465));
  jnot g26233(.din(n26341), .dout(n26466));
  jand g26234(.dina(n26466), .dinb(n26465), .dout(n26467));
  jnot g26235(.din(n26467), .dout(n26468));
  jand g26236(.dina(n26341), .dinb(n26284), .dout(n26469));
  jor  g26237(.dina(n26351), .dinb(n26469), .dout(n26470));
  jand g26238(.dina(n26470), .dinb(n26468), .dout(n26471));
  jxor g26239(.dina(n26471), .dinb(n26464), .dout(n26472));
  jand g26240(.dina(n23262), .dinb(n5693), .dout(n26473));
  jand g26241(.dina(n23260), .dinb(n6209), .dout(n26474));
  jand g26242(.dina(n22603), .dinb(n6131), .dout(n26475));
  jand g26243(.dina(n22539), .dinb(n5691), .dout(n26476));
  jor  g26244(.dina(n26476), .dinb(n26475), .dout(n26477));
  jor  g26245(.dina(n26477), .dinb(n26474), .dout(n26478));
  jor  g26246(.dina(n26478), .dinb(n26473), .dout(n26479));
  jxor g26247(.dina(n26479), .dinb(n4247), .dout(n26480));
  jnot g26248(.din(n26480), .dout(n26481));
  jxor g26249(.dina(n26481), .dinb(n26472), .dout(n26482));
  jand g26250(.dina(n26353), .dinb(n26281), .dout(n26483));
  jnot g26251(.din(n26483), .dout(n26484));
  jnot g26252(.din(n26281), .dout(n26485));
  jand g26253(.dina(n26352), .dinb(n26485), .dout(n26486));
  jor  g26254(.dina(n26363), .dinb(n26486), .dout(n26487));
  jand g26255(.dina(n26487), .dinb(n26484), .dout(n26488));
  jxor g26256(.dina(n26488), .dinb(n26482), .dout(n26489));
  jor  g26257(.dina(n23919), .dinb(n6341), .dout(n26490));
  jor  g26258(.dina(n23921), .dinb(n6797), .dout(n26491));
  jor  g26259(.dina(n23710), .dinb(n6557), .dout(n26492));
  jor  g26260(.dina(n23496), .dinb(n6339), .dout(n26493));
  jand g26261(.dina(n26493), .dinb(n26492), .dout(n26494));
  jand g26262(.dina(n26494), .dinb(n26491), .dout(n26495));
  jand g26263(.dina(n26495), .dinb(n26490), .dout(n26496));
  jxor g26264(.dina(n26496), .dinb(\a[17] ), .dout(n26497));
  jnot g26265(.din(n26497), .dout(n26498));
  jxor g26266(.dina(n26498), .dinb(n26489), .dout(n26499));
  jxor g26267(.dina(n26499), .dinb(n26391), .dout(n26500));
  jnot g26268(.din(n26366), .dout(n26501));
  jand g26269(.dina(n26501), .dinb(n26265), .dout(n26502));
  jnot g26270(.din(n26502), .dout(n26503));
  jnot g26271(.din(n26265), .dout(n26504));
  jand g26272(.dina(n26366), .dinb(n26504), .dout(n26505));
  jnot g26273(.din(n26375), .dout(n26506));
  jor  g26274(.dina(n26506), .dinb(n26505), .dout(n26507));
  jand g26275(.dina(n26507), .dinb(n26503), .dout(n26508));
  jxor g26276(.dina(n26508), .dinb(n26500), .dout(n26509));
  jand g26277(.dina(n26376), .dinb(n26261), .dout(n26510));
  jand g26278(.dina(n26377), .dinb(n26258), .dout(n26511));
  jor  g26279(.dina(n26511), .dinb(n26510), .dout(n26512));
  jxor g26280(.dina(n26512), .dinb(n26509), .dout(n26513));
  jxor g26281(.dina(n26513), .dinb(n26380), .dout(\result[18] ));
  jand g26282(.dina(n26513), .dinb(n26380), .dout(n26515));
  jand g26283(.dina(n26508), .dinb(n26500), .dout(n26516));
  jand g26284(.dina(n26512), .dinb(n26509), .dout(n26517));
  jor  g26285(.dina(n26517), .dinb(n26516), .dout(n26518));
  jor  g26286(.dina(n26447), .dinb(n26439), .dout(n26519));
  jand g26287(.dina(n26448), .dinb(n26400), .dout(n26520));
  jnot g26288(.din(n26520), .dout(n26521));
  jand g26289(.dina(n26521), .dinb(n26519), .dout(n26522));
  jnot g26290(.din(n26522), .dout(n26523));
  jand g26291(.dina(n26431), .dinb(n26425), .dout(n26524));
  jnot g26292(.din(n26524), .dout(n26525));
  jor  g26293(.dina(n26437), .dinb(n26433), .dout(n26526));
  jand g26294(.dina(n26526), .dinb(n26525), .dout(n26527));
  jnot g26295(.din(n26527), .dout(n26528));
  jand g26296(.dina(n21738), .dinb(n4449), .dout(n26529));
  jand g26297(.dina(n19513), .dinb(n4453), .dout(n26530));
  jand g26298(.dina(n19515), .dinb(n4457), .dout(n26531));
  jand g26299(.dina(n19517), .dinb(n4461), .dout(n26532));
  jor  g26300(.dina(n26532), .dinb(n26531), .dout(n26533));
  jor  g26301(.dina(n26533), .dinb(n26530), .dout(n26534));
  jor  g26302(.dina(n26534), .dinb(n26529), .dout(n26535));
  jxor g26303(.dina(n26535), .dinb(n88), .dout(n26536));
  jnot g26304(.din(n26536), .dout(n26537));
  jor  g26305(.dina(n26416), .dinb(n26306), .dout(n26538));
  jand g26306(.dina(n26424), .dinb(n26417), .dout(n26539));
  jnot g26307(.din(n26539), .dout(n26540));
  jand g26308(.dina(n26540), .dinb(n26538), .dout(n26541));
  jnot g26309(.din(n26541), .dout(n26542));
  jand g26310(.dina(n24593), .dinb(n12463), .dout(n26543));
  jxor g26311(.dina(n26543), .dinb(n5292), .dout(n26544));
  jand g26312(.dina(n4088), .dinb(n3386), .dout(n26545));
  jand g26313(.dina(n26545), .dinb(n1233), .dout(n26546));
  jand g26314(.dina(n689), .dinb(n184), .dout(n26547));
  jand g26315(.dina(n26547), .dinb(n108), .dout(n26548));
  jand g26316(.dina(n2697), .dinb(n2041), .dout(n26549));
  jand g26317(.dina(n26549), .dinb(n26548), .dout(n26550));
  jand g26318(.dina(n26550), .dinb(n13160), .dout(n26551));
  jand g26319(.dina(n26551), .dinb(n26546), .dout(n26552));
  jand g26320(.dina(n7441), .dinb(n1945), .dout(n26553));
  jand g26321(.dina(n26553), .dinb(n26552), .dout(n26554));
  jand g26322(.dina(n26554), .dinb(n12597), .dout(n26555));
  jand g26323(.dina(n26555), .dinb(n2170), .dout(n26556));
  jxor g26324(.dina(n26556), .dinb(n26305), .dout(n26557));
  jxor g26325(.dina(n26557), .dinb(n26544), .dout(n26558));
  jxor g26326(.dina(n26558), .dinb(n26542), .dout(n26559));
  jand g26327(.dina(n21240), .dinb(n732), .dout(n26560));
  jand g26328(.dina(n19519), .dinb(n3855), .dout(n26561));
  jand g26329(.dina(n19521), .dinb(n3858), .dout(n26562));
  jand g26330(.dina(n19523), .dinb(n3851), .dout(n26563));
  jor  g26331(.dina(n26563), .dinb(n26562), .dout(n26564));
  jor  g26332(.dina(n26564), .dinb(n26561), .dout(n26565));
  jor  g26333(.dina(n26565), .dinb(n26560), .dout(n26566));
  jxor g26334(.dina(n26566), .dinb(n26559), .dout(n26567));
  jxor g26335(.dina(n26567), .dinb(n26537), .dout(n26568));
  jxor g26336(.dina(n26568), .dinb(n26528), .dout(n26569));
  jnot g26337(.din(n26569), .dout(n26570));
  jand g26338(.dina(n19760), .dinb(n75), .dout(n26571));
  jand g26339(.dina(n19758), .dinb(n4933), .dout(n26572));
  jand g26340(.dina(n19510), .dinb(n4918), .dout(n26573));
  jand g26341(.dina(n19511), .dinb(n4745), .dout(n26574));
  jor  g26342(.dina(n26574), .dinb(n26573), .dout(n26575));
  jor  g26343(.dina(n26575), .dinb(n26572), .dout(n26576));
  jor  g26344(.dina(n26576), .dinb(n26571), .dout(n26577));
  jxor g26345(.dina(n26577), .dinb(n68), .dout(n26578));
  jxor g26346(.dina(n26578), .dinb(n26570), .dout(n26579));
  jxor g26347(.dina(n26579), .dinb(n26523), .dout(n26580));
  jand g26348(.dina(n22617), .dinb(n5365), .dout(n26581));
  jand g26349(.dina(n22539), .dinb(n5500), .dout(n26582));
  jand g26350(.dina(n22540), .dinb(n5424), .dout(n26583));
  jand g26351(.dina(n22248), .dinb(n5363), .dout(n26584));
  jor  g26352(.dina(n26584), .dinb(n26583), .dout(n26585));
  jor  g26353(.dina(n26585), .dinb(n26582), .dout(n26586));
  jor  g26354(.dina(n26586), .dinb(n26581), .dout(n26587));
  jxor g26355(.dina(n26587), .dinb(n72), .dout(n26588));
  jnot g26356(.din(n26588), .dout(n26589));
  jnot g26357(.din(n26449), .dout(n26590));
  jnot g26358(.din(n26453), .dout(n26591));
  jand g26359(.dina(n26591), .dinb(n26590), .dout(n26592));
  jnot g26360(.din(n26592), .dout(n26593));
  jand g26361(.dina(n26453), .dinb(n26449), .dout(n26594));
  jor  g26362(.dina(n26463), .dinb(n26594), .dout(n26595));
  jand g26363(.dina(n26595), .dinb(n26593), .dout(n26596));
  jxor g26364(.dina(n26596), .dinb(n26589), .dout(n26597));
  jxor g26365(.dina(n26597), .dinb(n26580), .dout(n26598));
  jnot g26366(.din(n26598), .dout(n26599));
  jor  g26367(.dina(n23494), .dinb(n5694), .dout(n26600));
  jor  g26368(.dina(n23496), .dinb(n6208), .dout(n26601));
  jor  g26369(.dina(n23450), .dinb(n6132), .dout(n26602));
  jor  g26370(.dina(n23449), .dinb(n5692), .dout(n26603));
  jand g26371(.dina(n26603), .dinb(n26602), .dout(n26604));
  jand g26372(.dina(n26604), .dinb(n26601), .dout(n26605));
  jand g26373(.dina(n26605), .dinb(n26600), .dout(n26606));
  jxor g26374(.dina(n26606), .dinb(\a[20] ), .dout(n26607));
  jxor g26375(.dina(n26607), .dinb(n26599), .dout(n26608));
  jnot g26376(.din(n26464), .dout(n26609));
  jnot g26377(.din(n26471), .dout(n26610));
  jand g26378(.dina(n26610), .dinb(n26609), .dout(n26611));
  jnot g26379(.din(n26611), .dout(n26612));
  jand g26380(.dina(n26471), .dinb(n26464), .dout(n26613));
  jor  g26381(.dina(n26481), .dinb(n26613), .dout(n26614));
  jand g26382(.dina(n26614), .dinb(n26612), .dout(n26615));
  jxor g26383(.dina(n26615), .dinb(n26608), .dout(n26616));
  jor  g26384(.dina(n24140), .dinb(n6341), .dout(n26617));
  jor  g26385(.dina(n24142), .dinb(n6797), .dout(n26618));
  jor  g26386(.dina(n23921), .dinb(n6557), .dout(n26619));
  jor  g26387(.dina(n23710), .dinb(n6339), .dout(n26620));
  jand g26388(.dina(n26620), .dinb(n26619), .dout(n26621));
  jand g26389(.dina(n26621), .dinb(n26618), .dout(n26622));
  jand g26390(.dina(n26622), .dinb(n26617), .dout(n26623));
  jxor g26391(.dina(n26623), .dinb(\a[17] ), .dout(n26624));
  jnot g26392(.din(n26624), .dout(n26625));
  jnot g26393(.din(n26482), .dout(n26626));
  jnot g26394(.din(n26488), .dout(n26627));
  jand g26395(.dina(n26627), .dinb(n26626), .dout(n26628));
  jnot g26396(.din(n26628), .dout(n26629));
  jand g26397(.dina(n26488), .dinb(n26482), .dout(n26630));
  jor  g26398(.dina(n26498), .dinb(n26630), .dout(n26631));
  jand g26399(.dina(n26631), .dinb(n26629), .dout(n26632));
  jxor g26400(.dina(n26632), .dinb(n26625), .dout(n26633));
  jxor g26401(.dina(n26633), .dinb(n26616), .dout(n26634));
  jnot g26402(.din(n26383), .dout(n26635));
  jand g26403(.dina(n26389), .dinb(n26635), .dout(n26636));
  jnot g26404(.din(n26636), .dout(n26637));
  jand g26405(.dina(n26390), .dinb(n26383), .dout(n26638));
  jor  g26406(.dina(n26499), .dinb(n26638), .dout(n26639));
  jand g26407(.dina(n26639), .dinb(n26637), .dout(n26640));
  jxor g26408(.dina(n26640), .dinb(n26634), .dout(n26641));
  jxor g26409(.dina(n26641), .dinb(n26518), .dout(n26642));
  jxor g26410(.dina(n26642), .dinb(n26515), .dout(\result[19] ));
  jand g26411(.dina(n26642), .dinb(n26515), .dout(n26644));
  jand g26412(.dina(n26640), .dinb(n26634), .dout(n26645));
  jand g26413(.dina(n26641), .dinb(n26518), .dout(n26646));
  jor  g26414(.dina(n26646), .dinb(n26645), .dout(n26647));
  jand g26415(.dina(n26632), .dinb(n26625), .dout(n26648));
  jand g26416(.dina(n26633), .dinb(n26616), .dout(n26649));
  jor  g26417(.dina(n26649), .dinb(n26648), .dout(n26650));
  jor  g26418(.dina(n26607), .dinb(n26599), .dout(n26651));
  jand g26419(.dina(n26615), .dinb(n26608), .dout(n26652));
  jnot g26420(.din(n26652), .dout(n26653));
  jand g26421(.dina(n26653), .dinb(n26651), .dout(n26654));
  jor  g26422(.dina(n23708), .dinb(n5694), .dout(n26655));
  jor  g26423(.dina(n23710), .dinb(n6208), .dout(n26656));
  jor  g26424(.dina(n23496), .dinb(n6132), .dout(n26657));
  jor  g26425(.dina(n23450), .dinb(n5692), .dout(n26658));
  jand g26426(.dina(n26658), .dinb(n26657), .dout(n26659));
  jand g26427(.dina(n26659), .dinb(n26656), .dout(n26660));
  jand g26428(.dina(n26660), .dinb(n26655), .dout(n26661));
  jxor g26429(.dina(n26661), .dinb(\a[20] ), .dout(n26662));
  jnot g26430(.din(n26662), .dout(n26663));
  jand g26431(.dina(n26596), .dinb(n26589), .dout(n26664));
  jand g26432(.dina(n26597), .dinb(n26580), .dout(n26665));
  jor  g26433(.dina(n26665), .dinb(n26664), .dout(n26666));
  jor  g26434(.dina(n26578), .dinb(n26570), .dout(n26667));
  jand g26435(.dina(n26579), .dinb(n26523), .dout(n26668));
  jnot g26436(.din(n26668), .dout(n26669));
  jand g26437(.dina(n26669), .dinb(n26667), .dout(n26670));
  jand g26438(.dina(n26567), .dinb(n26537), .dout(n26671));
  jand g26439(.dina(n26568), .dinb(n26528), .dout(n26672));
  jor  g26440(.dina(n26672), .dinb(n26671), .dout(n26673));
  jor  g26441(.dina(n26556), .dinb(n26305), .dout(n26674));
  jand g26442(.dina(n26557), .dinb(n26544), .dout(n26675));
  jnot g26443(.din(n26675), .dout(n26676));
  jand g26444(.dina(n26676), .dinb(n26674), .dout(n26677));
  jand g26445(.dina(n2660), .dinb(n442), .dout(n26678));
  jand g26446(.dina(n3092), .dinb(n861), .dout(n26679));
  jand g26447(.dina(n26679), .dinb(n26678), .dout(n26680));
  jand g26448(.dina(n391), .dinb(n103), .dout(n26681));
  jand g26449(.dina(n26681), .dinb(n1934), .dout(n26682));
  jand g26450(.dina(n26682), .dinb(n2321), .dout(n26683));
  jand g26451(.dina(n26683), .dinb(n26680), .dout(n26684));
  jand g26452(.dina(n14470), .dinb(n827), .dout(n26685));
  jand g26453(.dina(n26685), .dinb(n2769), .dout(n26686));
  jand g26454(.dina(n26686), .dinb(n773), .dout(n26687));
  jand g26455(.dina(n26687), .dinb(n26684), .dout(n26688));
  jand g26456(.dina(n13204), .dinb(n6427), .dout(n26689));
  jand g26457(.dina(n26689), .dinb(n26688), .dout(n26690));
  jand g26458(.dina(n26690), .dinb(n5765), .dout(n26691));
  jand g26459(.dina(n26691), .dinb(n3626), .dout(n26692));
  jnot g26460(.din(n26692), .dout(n26693));
  jxor g26461(.dina(n26693), .dinb(n26677), .dout(n26694));
  jand g26462(.dina(n21230), .dinb(n732), .dout(n26695));
  jand g26463(.dina(n19517), .dinb(n3855), .dout(n26696));
  jand g26464(.dina(n19519), .dinb(n3858), .dout(n26697));
  jand g26465(.dina(n19521), .dinb(n3851), .dout(n26698));
  jor  g26466(.dina(n26698), .dinb(n26697), .dout(n26699));
  jor  g26467(.dina(n26699), .dinb(n26696), .dout(n26700));
  jor  g26468(.dina(n26700), .dinb(n26695), .dout(n26701));
  jxor g26469(.dina(n26701), .dinb(n26694), .dout(n26702));
  jor  g26470(.dina(n26558), .dinb(n26542), .dout(n26703));
  jand g26471(.dina(n26558), .dinb(n26542), .dout(n26704));
  jor  g26472(.dina(n26566), .dinb(n26704), .dout(n26705));
  jand g26473(.dina(n26705), .dinb(n26703), .dout(n26706));
  jxor g26474(.dina(n26706), .dinb(n26702), .dout(n26707));
  jnot g26475(.din(n26707), .dout(n26708));
  jand g26476(.dina(n21762), .dinb(n4449), .dout(n26709));
  jand g26477(.dina(n19511), .dinb(n4453), .dout(n26710));
  jand g26478(.dina(n19513), .dinb(n4457), .dout(n26711));
  jand g26479(.dina(n19515), .dinb(n4461), .dout(n26712));
  jor  g26480(.dina(n26712), .dinb(n26711), .dout(n26713));
  jor  g26481(.dina(n26713), .dinb(n26710), .dout(n26714));
  jor  g26482(.dina(n26714), .dinb(n26709), .dout(n26715));
  jxor g26483(.dina(n26715), .dinb(n88), .dout(n26716));
  jxor g26484(.dina(n26716), .dinb(n26708), .dout(n26717));
  jxor g26485(.dina(n26717), .dinb(n26673), .dout(n26718));
  jand g26486(.dina(n22250), .dinb(n75), .dout(n26719));
  jand g26487(.dina(n22248), .dinb(n4933), .dout(n26720));
  jand g26488(.dina(n19758), .dinb(n4918), .dout(n26721));
  jand g26489(.dina(n19510), .dinb(n4745), .dout(n26722));
  jor  g26490(.dina(n26722), .dinb(n26721), .dout(n26723));
  jor  g26491(.dina(n26723), .dinb(n26720), .dout(n26724));
  jor  g26492(.dina(n26724), .dinb(n26719), .dout(n26725));
  jxor g26493(.dina(n26725), .dinb(n68), .dout(n26726));
  jnot g26494(.din(n26726), .dout(n26727));
  jxor g26495(.dina(n26727), .dinb(n26718), .dout(n26728));
  jnot g26496(.din(n26728), .dout(n26729));
  jxor g26497(.dina(n26729), .dinb(n26670), .dout(n26730));
  jand g26498(.dina(n22605), .dinb(n5365), .dout(n26731));
  jand g26499(.dina(n22603), .dinb(n5500), .dout(n26732));
  jand g26500(.dina(n22539), .dinb(n5424), .dout(n26733));
  jand g26501(.dina(n22540), .dinb(n5363), .dout(n26734));
  jor  g26502(.dina(n26734), .dinb(n26733), .dout(n26735));
  jor  g26503(.dina(n26735), .dinb(n26732), .dout(n26736));
  jor  g26504(.dina(n26736), .dinb(n26731), .dout(n26737));
  jxor g26505(.dina(n26737), .dinb(n72), .dout(n26738));
  jnot g26506(.din(n26738), .dout(n26739));
  jxor g26507(.dina(n26739), .dinb(n26730), .dout(n26740));
  jxor g26508(.dina(n26740), .dinb(n26666), .dout(n26741));
  jxor g26509(.dina(n26741), .dinb(n26663), .dout(n26742));
  jnot g26510(.din(n26742), .dout(n26743));
  jxor g26511(.dina(n26743), .dinb(n26654), .dout(n26744));
  jor  g26512(.dina(n24337), .dinb(n6341), .dout(n26745));
  jor  g26513(.dina(n24335), .dinb(n6797), .dout(n26746));
  jor  g26514(.dina(n24142), .dinb(n6557), .dout(n26747));
  jor  g26515(.dina(n23921), .dinb(n6339), .dout(n26748));
  jand g26516(.dina(n26748), .dinb(n26747), .dout(n26749));
  jand g26517(.dina(n26749), .dinb(n26746), .dout(n26750));
  jand g26518(.dina(n26750), .dinb(n26745), .dout(n26751));
  jxor g26519(.dina(n26751), .dinb(\a[17] ), .dout(n26752));
  jnot g26520(.din(n26752), .dout(n26753));
  jxor g26521(.dina(n26753), .dinb(n26744), .dout(n26754));
  jxor g26522(.dina(n26754), .dinb(n26650), .dout(n26755));
  jxor g26523(.dina(n26755), .dinb(n26647), .dout(n26756));
  jxor g26524(.dina(n26756), .dinb(n26644), .dout(\result[20] ));
  jand g26525(.dina(n26756), .dinb(n26644), .dout(n26758));
  jand g26526(.dina(n26740), .dinb(n26666), .dout(n26759));
  jand g26527(.dina(n26741), .dinb(n26663), .dout(n26760));
  jor  g26528(.dina(n26760), .dinb(n26759), .dout(n26761));
  jor  g26529(.dina(n24357), .dinb(n6341), .dout(n26762));
  jor  g26530(.dina(n24335), .dinb(n13559), .dout(n26763));
  jor  g26531(.dina(n24142), .dinb(n6339), .dout(n26764));
  jand g26532(.dina(n26764), .dinb(n26763), .dout(n26765));
  jand g26533(.dina(n26765), .dinb(n26762), .dout(n26766));
  jxor g26534(.dina(n26766), .dinb(\a[17] ), .dout(n26767));
  jnot g26535(.din(n26767), .dout(n26768));
  jxor g26536(.dina(n26768), .dinb(n26761), .dout(n26769));
  jand g26537(.dina(n26706), .dinb(n26702), .dout(n26770));
  jnot g26538(.din(n26770), .dout(n26771));
  jor  g26539(.dina(n26716), .dinb(n26708), .dout(n26772));
  jand g26540(.dina(n26772), .dinb(n26771), .dout(n26773));
  jnot g26541(.din(n26773), .dout(n26774));
  jand g26542(.dina(n21750), .dinb(n4449), .dout(n26775));
  jand g26543(.dina(n19510), .dinb(n4453), .dout(n26776));
  jand g26544(.dina(n19511), .dinb(n4457), .dout(n26777));
  jand g26545(.dina(n19513), .dinb(n4461), .dout(n26778));
  jor  g26546(.dina(n26778), .dinb(n26777), .dout(n26779));
  jor  g26547(.dina(n26779), .dinb(n26776), .dout(n26780));
  jor  g26548(.dina(n26780), .dinb(n26775), .dout(n26781));
  jxor g26549(.dina(n26781), .dinb(n88), .dout(n26782));
  jnot g26550(.din(n26782), .dout(n26783));
  jand g26551(.dina(n536), .dinb(n314), .dout(n26784));
  jand g26552(.dina(n26784), .dinb(n2135), .dout(n26785));
  jand g26553(.dina(n290), .dinb(n202), .dout(n26786));
  jand g26554(.dina(n1314), .dinb(n882), .dout(n26787));
  jand g26555(.dina(n26787), .dinb(n26786), .dout(n26788));
  jand g26556(.dina(n778), .dinb(n382), .dout(n26789));
  jand g26557(.dina(n26789), .dinb(n1359), .dout(n26790));
  jand g26558(.dina(n26790), .dinb(n26788), .dout(n26791));
  jand g26559(.dina(n26791), .dinb(n26785), .dout(n26792));
  jand g26560(.dina(n2859), .dinb(n1274), .dout(n26793));
  jand g26561(.dina(n2672), .dinb(n2292), .dout(n26794));
  jand g26562(.dina(n26794), .dinb(n26793), .dout(n26795));
  jand g26563(.dina(n26795), .dinb(n3299), .dout(n26796));
  jand g26564(.dina(n26796), .dinb(n3785), .dout(n26797));
  jand g26565(.dina(n26797), .dinb(n26792), .dout(n26798));
  jand g26566(.dina(n26798), .dinb(n4509), .dout(n26799));
  jand g26567(.dina(n5970), .dinb(n2040), .dout(n26800));
  jand g26568(.dina(n26800), .dinb(n26799), .dout(n26801));
  jxor g26569(.dina(n26801), .dinb(n26693), .dout(n26802));
  jand g26570(.dina(n26693), .dinb(n26677), .dout(n26803));
  jnot g26571(.din(n26803), .dout(n26804));
  jnot g26572(.din(n26677), .dout(n26805));
  jand g26573(.dina(n26692), .dinb(n26805), .dout(n26806));
  jor  g26574(.dina(n26701), .dinb(n26806), .dout(n26807));
  jand g26575(.dina(n26807), .dinb(n26804), .dout(n26808));
  jxor g26576(.dina(n26808), .dinb(n26802), .dout(n26809));
  jand g26577(.dina(n21218), .dinb(n732), .dout(n26810));
  jand g26578(.dina(n19515), .dinb(n3855), .dout(n26811));
  jand g26579(.dina(n19517), .dinb(n3858), .dout(n26812));
  jand g26580(.dina(n19519), .dinb(n3851), .dout(n26813));
  jor  g26581(.dina(n26813), .dinb(n26812), .dout(n26814));
  jor  g26582(.dina(n26814), .dinb(n26811), .dout(n26815));
  jor  g26583(.dina(n26815), .dinb(n26810), .dout(n26816));
  jxor g26584(.dina(n26816), .dinb(n26809), .dout(n26817));
  jxor g26585(.dina(n26817), .dinb(n26783), .dout(n26818));
  jxor g26586(.dina(n26818), .dinb(n26774), .dout(n26819));
  jand g26587(.dina(n22627), .dinb(n75), .dout(n26820));
  jand g26588(.dina(n22540), .dinb(n4933), .dout(n26821));
  jand g26589(.dina(n22248), .dinb(n4918), .dout(n26822));
  jand g26590(.dina(n19758), .dinb(n4745), .dout(n26823));
  jor  g26591(.dina(n26823), .dinb(n26822), .dout(n26824));
  jor  g26592(.dina(n26824), .dinb(n26821), .dout(n26825));
  jor  g26593(.dina(n26825), .dinb(n26820), .dout(n26826));
  jxor g26594(.dina(n26826), .dinb(n68), .dout(n26827));
  jnot g26595(.din(n26827), .dout(n26828));
  jxor g26596(.dina(n26828), .dinb(n26819), .dout(n26829));
  jor  g26597(.dina(n26717), .dinb(n26673), .dout(n26830));
  jand g26598(.dina(n26717), .dinb(n26673), .dout(n26831));
  jor  g26599(.dina(n26727), .dinb(n26831), .dout(n26832));
  jand g26600(.dina(n26832), .dinb(n26830), .dout(n26833));
  jxor g26601(.dina(n26833), .dinb(n26829), .dout(n26834));
  jand g26602(.dina(n23262), .dinb(n5365), .dout(n26835));
  jand g26603(.dina(n23260), .dinb(n5500), .dout(n26836));
  jand g26604(.dina(n22603), .dinb(n5424), .dout(n26837));
  jand g26605(.dina(n22539), .dinb(n5363), .dout(n26838));
  jor  g26606(.dina(n26838), .dinb(n26837), .dout(n26839));
  jor  g26607(.dina(n26839), .dinb(n26836), .dout(n26840));
  jor  g26608(.dina(n26840), .dinb(n26835), .dout(n26841));
  jxor g26609(.dina(n26841), .dinb(n72), .dout(n26842));
  jnot g26610(.din(n26842), .dout(n26843));
  jxor g26611(.dina(n26843), .dinb(n26834), .dout(n26844));
  jand g26612(.dina(n26729), .dinb(n26670), .dout(n26845));
  jnot g26613(.din(n26845), .dout(n26846));
  jnot g26614(.din(n26670), .dout(n26847));
  jand g26615(.dina(n26728), .dinb(n26847), .dout(n26848));
  jor  g26616(.dina(n26739), .dinb(n26848), .dout(n26849));
  jand g26617(.dina(n26849), .dinb(n26846), .dout(n26850));
  jxor g26618(.dina(n26850), .dinb(n26844), .dout(n26851));
  jor  g26619(.dina(n23919), .dinb(n5694), .dout(n26852));
  jor  g26620(.dina(n23921), .dinb(n6208), .dout(n26853));
  jor  g26621(.dina(n23710), .dinb(n6132), .dout(n26854));
  jor  g26622(.dina(n23496), .dinb(n5692), .dout(n26855));
  jand g26623(.dina(n26855), .dinb(n26854), .dout(n26856));
  jand g26624(.dina(n26856), .dinb(n26853), .dout(n26857));
  jand g26625(.dina(n26857), .dinb(n26852), .dout(n26858));
  jxor g26626(.dina(n26858), .dinb(\a[20] ), .dout(n26859));
  jnot g26627(.din(n26859), .dout(n26860));
  jxor g26628(.dina(n26860), .dinb(n26851), .dout(n26861));
  jxor g26629(.dina(n26861), .dinb(n26769), .dout(n26862));
  jand g26630(.dina(n26743), .dinb(n26654), .dout(n26863));
  jnot g26631(.din(n26863), .dout(n26864));
  jnot g26632(.din(n26654), .dout(n26865));
  jand g26633(.dina(n26742), .dinb(n26865), .dout(n26866));
  jor  g26634(.dina(n26753), .dinb(n26866), .dout(n26867));
  jand g26635(.dina(n26867), .dinb(n26864), .dout(n26868));
  jxor g26636(.dina(n26868), .dinb(n26862), .dout(n26869));
  jand g26637(.dina(n26754), .dinb(n26650), .dout(n26870));
  jand g26638(.dina(n26755), .dinb(n26647), .dout(n26871));
  jor  g26639(.dina(n26871), .dinb(n26870), .dout(n26872));
  jxor g26640(.dina(n26872), .dinb(n26869), .dout(n26873));
  jxor g26641(.dina(n26873), .dinb(n26758), .dout(\result[21] ));
  jand g26642(.dina(n26873), .dinb(n26758), .dout(n26875));
  jand g26643(.dina(n26868), .dinb(n26862), .dout(n26876));
  jand g26644(.dina(n26872), .dinb(n26869), .dout(n26877));
  jor  g26645(.dina(n26877), .dinb(n26876), .dout(n26878));
  jor  g26646(.dina(n23494), .dinb(n5366), .dout(n26879));
  jor  g26647(.dina(n23496), .dinb(n5499), .dout(n26880));
  jor  g26648(.dina(n23450), .dinb(n5425), .dout(n26881));
  jor  g26649(.dina(n23449), .dinb(n5364), .dout(n26882));
  jand g26650(.dina(n26882), .dinb(n26881), .dout(n26883));
  jand g26651(.dina(n26883), .dinb(n26880), .dout(n26884));
  jand g26652(.dina(n26884), .dinb(n26879), .dout(n26885));
  jxor g26653(.dina(n26885), .dinb(\a[23] ), .dout(n26886));
  jnot g26654(.din(n26886), .dout(n26887));
  jand g26655(.dina(n22617), .dinb(n75), .dout(n26888));
  jand g26656(.dina(n22539), .dinb(n4933), .dout(n26889));
  jand g26657(.dina(n22540), .dinb(n4918), .dout(n26890));
  jand g26658(.dina(n22248), .dinb(n4745), .dout(n26891));
  jor  g26659(.dina(n26891), .dinb(n26890), .dout(n26892));
  jor  g26660(.dina(n26892), .dinb(n26889), .dout(n26893));
  jor  g26661(.dina(n26893), .dinb(n26888), .dout(n26894));
  jxor g26662(.dina(n26894), .dinb(n68), .dout(n26895));
  jnot g26663(.din(n26895), .dout(n26896));
  jor  g26664(.dina(n26818), .dinb(n26774), .dout(n26897));
  jand g26665(.dina(n26818), .dinb(n26774), .dout(n26898));
  jor  g26666(.dina(n26828), .dinb(n26898), .dout(n26899));
  jand g26667(.dina(n26899), .dinb(n26897), .dout(n26900));
  jxor g26668(.dina(n26900), .dinb(n26896), .dout(n26901));
  jand g26669(.dina(n19760), .dinb(n4449), .dout(n26902));
  jand g26670(.dina(n19758), .dinb(n4453), .dout(n26903));
  jand g26671(.dina(n19510), .dinb(n4457), .dout(n26904));
  jand g26672(.dina(n19511), .dinb(n4461), .dout(n26905));
  jor  g26673(.dina(n26905), .dinb(n26904), .dout(n26906));
  jor  g26674(.dina(n26906), .dinb(n26903), .dout(n26907));
  jor  g26675(.dina(n26907), .dinb(n26902), .dout(n26908));
  jxor g26676(.dina(n26908), .dinb(n88), .dout(n26909));
  jnot g26677(.din(n26909), .dout(n26910));
  jand g26678(.dina(n26816), .dinb(n26809), .dout(n26911));
  jand g26679(.dina(n26817), .dinb(n26783), .dout(n26912));
  jor  g26680(.dina(n26912), .dinb(n26911), .dout(n26913));
  jand g26681(.dina(n26801), .dinb(n26693), .dout(n26914));
  jand g26682(.dina(n26808), .dinb(n26802), .dout(n26915));
  jor  g26683(.dina(n26915), .dinb(n26914), .dout(n26916));
  jand g26684(.dina(n24593), .dinb(n12536), .dout(n26917));
  jxor g26685(.dina(n26917), .dinb(n5064), .dout(n26918));
  jand g26686(.dina(n1409), .dinb(n819), .dout(n26919));
  jand g26687(.dina(n26919), .dinb(n202), .dout(n26920));
  jand g26688(.dina(n1821), .dinb(n1432), .dout(n26921));
  jand g26689(.dina(n26921), .dinb(n26920), .dout(n26922));
  jand g26690(.dina(n21670), .dinb(n2044), .dout(n26923));
  jand g26691(.dina(n26923), .dinb(n26922), .dout(n26924));
  jand g26692(.dina(n3633), .dinb(n1832), .dout(n26925));
  jand g26693(.dina(n26925), .dinb(n12709), .dout(n26926));
  jand g26694(.dina(n26926), .dinb(n26924), .dout(n26927));
  jand g26695(.dina(n26927), .dinb(n1458), .dout(n26928));
  jand g26696(.dina(n5602), .dinb(n4807), .dout(n26929));
  jand g26697(.dina(n26929), .dinb(n26928), .dout(n26930));
  jxor g26698(.dina(n26930), .dinb(n26801), .dout(n26931));
  jxor g26699(.dina(n26931), .dinb(n26918), .dout(n26932));
  jand g26700(.dina(n21738), .dinb(n732), .dout(n26933));
  jand g26701(.dina(n19513), .dinb(n3855), .dout(n26934));
  jand g26702(.dina(n19515), .dinb(n3858), .dout(n26935));
  jand g26703(.dina(n19517), .dinb(n3851), .dout(n26936));
  jor  g26704(.dina(n26936), .dinb(n26935), .dout(n26937));
  jor  g26705(.dina(n26937), .dinb(n26934), .dout(n26938));
  jor  g26706(.dina(n26938), .dinb(n26933), .dout(n26939));
  jxor g26707(.dina(n26939), .dinb(n26932), .dout(n26940));
  jxor g26708(.dina(n26940), .dinb(n26916), .dout(n26941));
  jxor g26709(.dina(n26941), .dinb(n26913), .dout(n26942));
  jxor g26710(.dina(n26942), .dinb(n26910), .dout(n26943));
  jxor g26711(.dina(n26943), .dinb(n26901), .dout(n26944));
  jxor g26712(.dina(n26944), .dinb(n26887), .dout(n26945));
  jnot g26713(.din(n26829), .dout(n26946));
  jnot g26714(.din(n26833), .dout(n26947));
  jand g26715(.dina(n26947), .dinb(n26946), .dout(n26948));
  jnot g26716(.din(n26948), .dout(n26949));
  jand g26717(.dina(n26833), .dinb(n26829), .dout(n26950));
  jor  g26718(.dina(n26843), .dinb(n26950), .dout(n26951));
  jand g26719(.dina(n26951), .dinb(n26949), .dout(n26952));
  jxor g26720(.dina(n26952), .dinb(n26945), .dout(n26953));
  jor  g26721(.dina(n24140), .dinb(n5694), .dout(n26954));
  jor  g26722(.dina(n24142), .dinb(n6208), .dout(n26955));
  jor  g26723(.dina(n23921), .dinb(n6132), .dout(n26956));
  jor  g26724(.dina(n23710), .dinb(n5692), .dout(n26957));
  jand g26725(.dina(n26957), .dinb(n26956), .dout(n26958));
  jand g26726(.dina(n26958), .dinb(n26955), .dout(n26959));
  jand g26727(.dina(n26959), .dinb(n26954), .dout(n26960));
  jxor g26728(.dina(n26960), .dinb(\a[20] ), .dout(n26961));
  jnot g26729(.din(n26961), .dout(n26962));
  jnot g26730(.din(n26844), .dout(n26963));
  jnot g26731(.din(n26850), .dout(n26964));
  jand g26732(.dina(n26964), .dinb(n26963), .dout(n26965));
  jnot g26733(.din(n26965), .dout(n26966));
  jand g26734(.dina(n26850), .dinb(n26844), .dout(n26967));
  jor  g26735(.dina(n26860), .dinb(n26967), .dout(n26968));
  jand g26736(.dina(n26968), .dinb(n26966), .dout(n26969));
  jxor g26737(.dina(n26969), .dinb(n26962), .dout(n26970));
  jxor g26738(.dina(n26970), .dinb(n26953), .dout(n26971));
  jnot g26739(.din(n26761), .dout(n26972));
  jand g26740(.dina(n26767), .dinb(n26972), .dout(n26973));
  jnot g26741(.din(n26973), .dout(n26974));
  jand g26742(.dina(n26768), .dinb(n26761), .dout(n26975));
  jor  g26743(.dina(n26861), .dinb(n26975), .dout(n26976));
  jand g26744(.dina(n26976), .dinb(n26974), .dout(n26977));
  jxor g26745(.dina(n26977), .dinb(n26971), .dout(n26978));
  jxor g26746(.dina(n26978), .dinb(n26878), .dout(n26979));
  jxor g26747(.dina(n26979), .dinb(n26875), .dout(\result[22] ));
  jand g26748(.dina(n26979), .dinb(n26875), .dout(n26981));
  jand g26749(.dina(n26977), .dinb(n26971), .dout(n26982));
  jand g26750(.dina(n26978), .dinb(n26878), .dout(n26983));
  jor  g26751(.dina(n26983), .dinb(n26982), .dout(n26984));
  jand g26752(.dina(n26969), .dinb(n26962), .dout(n26985));
  jand g26753(.dina(n26970), .dinb(n26953), .dout(n26986));
  jor  g26754(.dina(n26986), .dinb(n26985), .dout(n26987));
  jand g26755(.dina(n26944), .dinb(n26887), .dout(n26988));
  jand g26756(.dina(n26952), .dinb(n26945), .dout(n26989));
  jor  g26757(.dina(n26989), .dinb(n26988), .dout(n26990));
  jor  g26758(.dina(n23708), .dinb(n5366), .dout(n26991));
  jor  g26759(.dina(n23710), .dinb(n5499), .dout(n26992));
  jor  g26760(.dina(n23496), .dinb(n5425), .dout(n26993));
  jor  g26761(.dina(n23450), .dinb(n5364), .dout(n26994));
  jand g26762(.dina(n26994), .dinb(n26993), .dout(n26995));
  jand g26763(.dina(n26995), .dinb(n26992), .dout(n26996));
  jand g26764(.dina(n26996), .dinb(n26991), .dout(n26997));
  jxor g26765(.dina(n26997), .dinb(\a[23] ), .dout(n26998));
  jnot g26766(.din(n26998), .dout(n26999));
  jand g26767(.dina(n26900), .dinb(n26896), .dout(n27000));
  jand g26768(.dina(n26943), .dinb(n26901), .dout(n27001));
  jor  g26769(.dina(n27001), .dinb(n27000), .dout(n27002));
  jand g26770(.dina(n26939), .dinb(n26932), .dout(n27003));
  jand g26771(.dina(n26940), .dinb(n26916), .dout(n27004));
  jor  g26772(.dina(n27004), .dinb(n27003), .dout(n27005));
  jor  g26773(.dina(n26930), .dinb(n26801), .dout(n27006));
  jand g26774(.dina(n26931), .dinb(n26918), .dout(n27007));
  jnot g26775(.din(n27007), .dout(n27008));
  jand g26776(.dina(n27008), .dinb(n27006), .dout(n27009));
  jand g26777(.dina(n5003), .dinb(n559), .dout(n27010));
  jand g26778(.dina(n27010), .dinb(n1160), .dout(n27011));
  jand g26779(.dina(n329), .dinb(n82), .dout(n27012));
  jand g26780(.dina(n614), .dinb(n553), .dout(n27013));
  jand g26781(.dina(n27013), .dinb(n27012), .dout(n27014));
  jnot g26782(.din(n1366), .dout(n27015));
  jand g26783(.dina(n1474), .dinb(n27015), .dout(n27016));
  jand g26784(.dina(n27016), .dinb(n27014), .dout(n27017));
  jand g26785(.dina(n12417), .dinb(n3502), .dout(n27018));
  jand g26786(.dina(n27018), .dinb(n27017), .dout(n27019));
  jand g26787(.dina(n27019), .dinb(n27011), .dout(n27020));
  jand g26788(.dina(n3392), .dinb(n1103), .dout(n27021));
  jand g26789(.dina(n27021), .dinb(n27020), .dout(n27022));
  jand g26790(.dina(n27022), .dinb(n25492), .dout(n27023));
  jand g26791(.dina(n27023), .dinb(n7028), .dout(n27024));
  jnot g26792(.din(n27024), .dout(n27025));
  jxor g26793(.dina(n27025), .dinb(n27009), .dout(n27026));
  jand g26794(.dina(n21762), .dinb(n732), .dout(n27027));
  jand g26795(.dina(n19511), .dinb(n3855), .dout(n27028));
  jand g26796(.dina(n19513), .dinb(n3858), .dout(n27029));
  jand g26797(.dina(n19515), .dinb(n3851), .dout(n27030));
  jor  g26798(.dina(n27030), .dinb(n27029), .dout(n27031));
  jor  g26799(.dina(n27031), .dinb(n27028), .dout(n27032));
  jor  g26800(.dina(n27032), .dinb(n27027), .dout(n27033));
  jxor g26801(.dina(n27033), .dinb(n27026), .dout(n27034));
  jxor g26802(.dina(n27034), .dinb(n27005), .dout(n27035));
  jnot g26803(.din(n27035), .dout(n27036));
  jand g26804(.dina(n22250), .dinb(n4449), .dout(n27037));
  jand g26805(.dina(n22248), .dinb(n4453), .dout(n27038));
  jand g26806(.dina(n19758), .dinb(n4457), .dout(n27039));
  jand g26807(.dina(n19510), .dinb(n4461), .dout(n27040));
  jor  g26808(.dina(n27040), .dinb(n27039), .dout(n27041));
  jor  g26809(.dina(n27041), .dinb(n27038), .dout(n27042));
  jor  g26810(.dina(n27042), .dinb(n27037), .dout(n27043));
  jxor g26811(.dina(n27043), .dinb(n88), .dout(n27044));
  jxor g26812(.dina(n27044), .dinb(n27036), .dout(n27045));
  jor  g26813(.dina(n26941), .dinb(n26913), .dout(n27046));
  jand g26814(.dina(n26941), .dinb(n26913), .dout(n27047));
  jor  g26815(.dina(n27047), .dinb(n26910), .dout(n27048));
  jand g26816(.dina(n27048), .dinb(n27046), .dout(n27049));
  jxor g26817(.dina(n27049), .dinb(n27045), .dout(n27050));
  jand g26818(.dina(n22605), .dinb(n75), .dout(n27051));
  jand g26819(.dina(n22603), .dinb(n4933), .dout(n27052));
  jand g26820(.dina(n22539), .dinb(n4918), .dout(n27053));
  jand g26821(.dina(n22540), .dinb(n4745), .dout(n27054));
  jor  g26822(.dina(n27054), .dinb(n27053), .dout(n27055));
  jor  g26823(.dina(n27055), .dinb(n27052), .dout(n27056));
  jor  g26824(.dina(n27056), .dinb(n27051), .dout(n27057));
  jxor g26825(.dina(n27057), .dinb(n68), .dout(n27058));
  jnot g26826(.din(n27058), .dout(n27059));
  jxor g26827(.dina(n27059), .dinb(n27050), .dout(n27060));
  jxor g26828(.dina(n27060), .dinb(n27002), .dout(n27061));
  jxor g26829(.dina(n27061), .dinb(n26999), .dout(n27062));
  jxor g26830(.dina(n27062), .dinb(n26990), .dout(n27063));
  jor  g26831(.dina(n24337), .dinb(n5694), .dout(n27064));
  jor  g26832(.dina(n23921), .dinb(n5692), .dout(n27067));
  jand g26833(.dina(n27067), .dinb(n27064), .dout(n27070));
  jxor g26834(.dina(n27070), .dinb(\a[20] ), .dout(n27071));
  jnot g26835(.din(n27071), .dout(n27072));
  jxor g26836(.dina(n27072), .dinb(n27063), .dout(n27073));
  jxor g26837(.dina(n27073), .dinb(n26987), .dout(n27074));
  jxor g26838(.dina(n27074), .dinb(n26984), .dout(n27075));
  jxor g26839(.dina(n27075), .dinb(n26981), .dout(\result[23] ));
  jand g26840(.dina(n27075), .dinb(n26981), .dout(n27077));
  jnot g26841(.din(n4247), .dout(n27084));
  jor  g26842(.dina(n27060), .dinb(n27002), .dout(n27085));
  jand g26843(.dina(n27060), .dinb(n27002), .dout(n27086));
  jor  g26844(.dina(n27086), .dinb(n26999), .dout(n27087));
  jand g26845(.dina(n27087), .dinb(n27085), .dout(n27088));
  jxor g26846(.dina(n27088), .dinb(n27084), .dout(n27089));
  jand g26847(.dina(n23262), .dinb(n75), .dout(n27090));
  jand g26848(.dina(n23260), .dinb(n4933), .dout(n27091));
  jand g26849(.dina(n22603), .dinb(n4918), .dout(n27092));
  jand g26850(.dina(n22539), .dinb(n4745), .dout(n27093));
  jor  g26851(.dina(n27093), .dinb(n27092), .dout(n27094));
  jor  g26852(.dina(n27094), .dinb(n27091), .dout(n27095));
  jor  g26853(.dina(n27095), .dinb(n27090), .dout(n27096));
  jxor g26854(.dina(n27096), .dinb(n68), .dout(n27097));
  jnot g26855(.din(n27097), .dout(n27098));
  jand g26856(.dina(n12218), .dinb(n1185), .dout(n27099));
  jand g26857(.dina(n27099), .dinb(n1410), .dout(n27100));
  jand g26858(.dina(n853), .dinb(n418), .dout(n27101));
  jand g26859(.dina(n27101), .dinb(n12248), .dout(n27102));
  jand g26860(.dina(n27102), .dinb(n12731), .dout(n27103));
  jand g26861(.dina(n27103), .dinb(n26785), .dout(n27104));
  jand g26862(.dina(n27104), .dinb(n27100), .dout(n27105));
  jand g26863(.dina(n24740), .dinb(n4800), .dout(n27106));
  jand g26864(.dina(n27106), .dinb(n27105), .dout(n27107));
  jand g26865(.dina(n7073), .dinb(n5267), .dout(n27108));
  jand g26866(.dina(n27108), .dinb(n27107), .dout(n27109));
  jand g26867(.dina(n27109), .dinb(n1481), .dout(n27110));
  jxor g26868(.dina(n27110), .dinb(n27025), .dout(n27111));
  jand g26869(.dina(n21750), .dinb(n732), .dout(n27112));
  jand g26870(.dina(n19510), .dinb(n3855), .dout(n27113));
  jand g26871(.dina(n19511), .dinb(n3858), .dout(n27114));
  jand g26872(.dina(n19513), .dinb(n3851), .dout(n27115));
  jor  g26873(.dina(n27115), .dinb(n27114), .dout(n27116));
  jor  g26874(.dina(n27116), .dinb(n27113), .dout(n27117));
  jor  g26875(.dina(n27117), .dinb(n27112), .dout(n27118));
  jxor g26876(.dina(n27118), .dinb(n27111), .dout(n27119));
  jand g26877(.dina(n27025), .dinb(n27009), .dout(n27120));
  jnot g26878(.din(n27120), .dout(n27121));
  jnot g26879(.din(n27009), .dout(n27122));
  jand g26880(.dina(n27024), .dinb(n27122), .dout(n27123));
  jor  g26881(.dina(n27033), .dinb(n27123), .dout(n27124));
  jand g26882(.dina(n27124), .dinb(n27121), .dout(n27125));
  jxor g26883(.dina(n27125), .dinb(n27119), .dout(n27126));
  jnot g26884(.din(n27126), .dout(n27127));
  jand g26885(.dina(n27034), .dinb(n27005), .dout(n27128));
  jnot g26886(.din(n27128), .dout(n27129));
  jor  g26887(.dina(n27044), .dinb(n27036), .dout(n27130));
  jand g26888(.dina(n27130), .dinb(n27129), .dout(n27131));
  jxor g26889(.dina(n27131), .dinb(n27127), .dout(n27132));
  jnot g26890(.din(n27132), .dout(n27133));
  jand g26891(.dina(n22627), .dinb(n4449), .dout(n27134));
  jand g26892(.dina(n22540), .dinb(n4453), .dout(n27135));
  jand g26893(.dina(n22248), .dinb(n4457), .dout(n27136));
  jand g26894(.dina(n19758), .dinb(n4461), .dout(n27137));
  jor  g26895(.dina(n27137), .dinb(n27136), .dout(n27138));
  jor  g26896(.dina(n27138), .dinb(n27135), .dout(n27139));
  jor  g26897(.dina(n27139), .dinb(n27134), .dout(n27140));
  jxor g26898(.dina(n27140), .dinb(n88), .dout(n27141));
  jxor g26899(.dina(n27141), .dinb(n27133), .dout(n27142));
  jxor g26900(.dina(n27142), .dinb(n27098), .dout(n27143));
  jor  g26901(.dina(n27049), .dinb(n27045), .dout(n27144));
  jand g26902(.dina(n27049), .dinb(n27045), .dout(n27145));
  jor  g26903(.dina(n27059), .dinb(n27145), .dout(n27146));
  jand g26904(.dina(n27146), .dinb(n27144), .dout(n27147));
  jxor g26905(.dina(n27147), .dinb(n27143), .dout(n27148));
  jor  g26906(.dina(n23919), .dinb(n5366), .dout(n27149));
  jor  g26907(.dina(n23921), .dinb(n5499), .dout(n27150));
  jor  g26908(.dina(n23710), .dinb(n5425), .dout(n27151));
  jor  g26909(.dina(n23496), .dinb(n5364), .dout(n27152));
  jand g26910(.dina(n27152), .dinb(n27151), .dout(n27153));
  jand g26911(.dina(n27153), .dinb(n27150), .dout(n27154));
  jand g26912(.dina(n27154), .dinb(n27149), .dout(n27155));
  jxor g26913(.dina(n27155), .dinb(\a[23] ), .dout(n27156));
  jnot g26914(.din(n27156), .dout(n27157));
  jxor g26915(.dina(n27157), .dinb(n27148), .dout(n27158));
  jxor g26916(.dina(n27158), .dinb(n27089), .dout(n27159));
  jnot g26917(.din(n26990), .dout(n27160));
  jnot g26918(.din(n27062), .dout(n27161));
  jand g26919(.dina(n27161), .dinb(n27160), .dout(n27162));
  jnot g26920(.din(n27162), .dout(n27163));
  jand g26921(.dina(n27062), .dinb(n26990), .dout(n27164));
  jor  g26922(.dina(n27072), .dinb(n27164), .dout(n27165));
  jand g26923(.dina(n27165), .dinb(n27163), .dout(n27166));
  jxor g26924(.dina(n27166), .dinb(n27159), .dout(n27167));
  jand g26925(.dina(n27073), .dinb(n26987), .dout(n27168));
  jand g26926(.dina(n27074), .dinb(n26984), .dout(n27169));
  jor  g26927(.dina(n27169), .dinb(n27168), .dout(n27170));
  jxor g26928(.dina(n27170), .dinb(n27167), .dout(n27171));
  jxor g26929(.dina(n27171), .dinb(n27077), .dout(\result[24] ));
  jand g26930(.dina(n27171), .dinb(n27077), .dout(n27173));
  jand g26931(.dina(n27166), .dinb(n27159), .dout(n27174));
  jand g26932(.dina(n27170), .dinb(n27167), .dout(n27175));
  jor  g26933(.dina(n27175), .dinb(n27174), .dout(n27176));
  jor  g26934(.dina(n27141), .dinb(n27133), .dout(n27177));
  jand g26935(.dina(n27142), .dinb(n27098), .dout(n27178));
  jnot g26936(.din(n27178), .dout(n27179));
  jand g26937(.dina(n27179), .dinb(n27177), .dout(n27180));
  jnot g26938(.din(n27180), .dout(n27181));
  jor  g26939(.dina(n23494), .dinb(n4747), .dout(n27182));
  jor  g26940(.dina(n23496), .dinb(n4959), .dout(n27183));
  jor  g26941(.dina(n23450), .dinb(n4919), .dout(n27184));
  jor  g26942(.dina(n23449), .dinb(n4746), .dout(n27185));
  jand g26943(.dina(n27185), .dinb(n27184), .dout(n27186));
  jand g26944(.dina(n27186), .dinb(n27183), .dout(n27187));
  jand g26945(.dina(n27187), .dinb(n27182), .dout(n27188));
  jxor g26946(.dina(n27188), .dinb(\a[26] ), .dout(n27189));
  jnot g26947(.din(n27189), .dout(n27190));
  jand g26948(.dina(n27125), .dinb(n27119), .dout(n27191));
  jnot g26949(.din(n27191), .dout(n27192));
  jor  g26950(.dina(n27131), .dinb(n27127), .dout(n27193));
  jand g26951(.dina(n27193), .dinb(n27192), .dout(n27194));
  jnot g26952(.din(n27194), .dout(n27195));
  jor  g26953(.dina(n27110), .dinb(n27025), .dout(n27196));
  jand g26954(.dina(n27118), .dinb(n27111), .dout(n27197));
  jnot g26955(.din(n27197), .dout(n27198));
  jand g26956(.dina(n27198), .dinb(n27196), .dout(n27199));
  jnot g26957(.din(n27199), .dout(n27200));
  jand g26958(.dina(n24593), .dinb(n12959), .dout(n27201));
  jxor g26959(.dina(n27201), .dinb(n4247), .dout(n27202));
  jand g26960(.dina(n4667), .dinb(n1145), .dout(n27203));
  jand g26961(.dina(n27203), .dinb(n1009), .dout(n27204));
  jand g26962(.dina(n689), .dinb(n340), .dout(n27205));
  jand g26963(.dina(n619), .dinb(n476), .dout(n27206));
  jand g26964(.dina(n27206), .dinb(n27205), .dout(n27207));
  jand g26965(.dina(n1975), .dinb(n1205), .dout(n27208));
  jand g26966(.dina(n27208), .dinb(n27207), .dout(n27209));
  jand g26967(.dina(n27209), .dinb(n27204), .dout(n27210));
  jand g26968(.dina(n13626), .dinb(n3299), .dout(n27211));
  jand g26969(.dina(n27211), .dinb(n27210), .dout(n27212));
  jand g26970(.dina(n1488), .dinb(n903), .dout(n27213));
  jand g26971(.dina(n27213), .dinb(n3566), .dout(n27214));
  jand g26972(.dina(n27214), .dinb(n14415), .dout(n27215));
  jand g26973(.dina(n27215), .dinb(n27212), .dout(n27216));
  jand g26974(.dina(n27216), .dinb(n1894), .dout(n27217));
  jand g26975(.dina(n27217), .dinb(n5164), .dout(n27218));
  jxor g26976(.dina(n27218), .dinb(n27024), .dout(n27219));
  jxor g26977(.dina(n27219), .dinb(n27202), .dout(n27220));
  jxor g26978(.dina(n27220), .dinb(n27200), .dout(n27221));
  jand g26979(.dina(n19760), .dinb(n732), .dout(n27222));
  jand g26980(.dina(n19758), .dinb(n3855), .dout(n27223));
  jand g26981(.dina(n19510), .dinb(n3858), .dout(n27224));
  jand g26982(.dina(n19511), .dinb(n3851), .dout(n27225));
  jor  g26983(.dina(n27225), .dinb(n27224), .dout(n27226));
  jor  g26984(.dina(n27226), .dinb(n27223), .dout(n27227));
  jor  g26985(.dina(n27227), .dinb(n27222), .dout(n27228));
  jxor g26986(.dina(n27228), .dinb(n27221), .dout(n27229));
  jxor g26987(.dina(n27229), .dinb(n27195), .dout(n27230));
  jand g26988(.dina(n22617), .dinb(n4449), .dout(n27231));
  jand g26989(.dina(n22539), .dinb(n4453), .dout(n27232));
  jand g26990(.dina(n22540), .dinb(n4457), .dout(n27233));
  jand g26991(.dina(n22248), .dinb(n4461), .dout(n27234));
  jor  g26992(.dina(n27234), .dinb(n27233), .dout(n27235));
  jor  g26993(.dina(n27235), .dinb(n27232), .dout(n27236));
  jor  g26994(.dina(n27236), .dinb(n27231), .dout(n27237));
  jxor g26995(.dina(n27237), .dinb(n88), .dout(n27238));
  jnot g26996(.din(n27238), .dout(n27239));
  jxor g26997(.dina(n27239), .dinb(n27230), .dout(n27240));
  jxor g26998(.dina(n27240), .dinb(n27190), .dout(n27241));
  jxor g26999(.dina(n27241), .dinb(n27181), .dout(n27242));
  jor  g27000(.dina(n24140), .dinb(n5366), .dout(n27243));
  jor  g27001(.dina(n23921), .dinb(n5425), .dout(n27245));
  jor  g27002(.dina(n23710), .dinb(n5364), .dout(n27246));
  jand g27003(.dina(n27246), .dinb(n27245), .dout(n27247));
  jand g27004(.dina(n27247), .dinb(n27243), .dout(n27249));
  jxor g27005(.dina(n27249), .dinb(\a[23] ), .dout(n27250));
  jnot g27006(.din(n27250), .dout(n27251));
  jnot g27007(.din(n27143), .dout(n27252));
  jnot g27008(.din(n27147), .dout(n27253));
  jand g27009(.dina(n27253), .dinb(n27252), .dout(n27254));
  jnot g27010(.din(n27254), .dout(n27255));
  jand g27011(.dina(n27147), .dinb(n27143), .dout(n27256));
  jor  g27012(.dina(n27157), .dinb(n27256), .dout(n27257));
  jand g27013(.dina(n27257), .dinb(n27255), .dout(n27258));
  jxor g27014(.dina(n27258), .dinb(n27251), .dout(n27259));
  jxor g27015(.dina(n27259), .dinb(n27242), .dout(n27260));
  jor  g27016(.dina(n27088), .dinb(n27084), .dout(n27261));
  jand g27017(.dina(n27088), .dinb(n27084), .dout(n27262));
  jor  g27018(.dina(n27158), .dinb(n27262), .dout(n27263));
  jand g27019(.dina(n27263), .dinb(n27261), .dout(n27264));
  jxor g27020(.dina(n27264), .dinb(n27260), .dout(n27265));
  jxor g27021(.dina(n27265), .dinb(n27176), .dout(n27266));
  jxor g27022(.dina(n27266), .dinb(n27173), .dout(\result[25] ));
  jand g27023(.dina(n27266), .dinb(n27173), .dout(n27268));
  jand g27024(.dina(n27264), .dinb(n27260), .dout(n27269));
  jand g27025(.dina(n27265), .dinb(n27176), .dout(n27270));
  jor  g27026(.dina(n27270), .dinb(n27269), .dout(n27271));
  jand g27027(.dina(n27258), .dinb(n27251), .dout(n27272));
  jand g27028(.dina(n27259), .dinb(n27242), .dout(n27273));
  jor  g27029(.dina(n27273), .dinb(n27272), .dout(n27274));
  jand g27030(.dina(n27240), .dinb(n27190), .dout(n27275));
  jand g27031(.dina(n27241), .dinb(n27181), .dout(n27276));
  jor  g27032(.dina(n27276), .dinb(n27275), .dout(n27277));
  jor  g27033(.dina(n27218), .dinb(n27024), .dout(n27278));
  jand g27034(.dina(n27219), .dinb(n27202), .dout(n27279));
  jnot g27035(.din(n27279), .dout(n27280));
  jand g27036(.dina(n27280), .dinb(n27278), .dout(n27281));
  jand g27037(.dina(n424), .dinb(n217), .dout(n27282));
  jand g27038(.dina(n893), .dinb(n249), .dout(n27283));
  jand g27039(.dina(n27283), .dinb(n27282), .dout(n27284));
  jand g27040(.dina(n27284), .dinb(n1183), .dout(n27285));
  jand g27041(.dina(n27285), .dinb(n4183), .dout(n27286));
  jand g27042(.dina(n5549), .dinb(n2413), .dout(n27287));
  jand g27043(.dina(n27287), .dinb(n2547), .dout(n27288));
  jand g27044(.dina(n27288), .dinb(n2472), .dout(n27289));
  jand g27045(.dina(n27289), .dinb(n27286), .dout(n27290));
  jand g27046(.dina(n14473), .dinb(n4075), .dout(n27291));
  jand g27047(.dina(n27291), .dinb(n27290), .dout(n27292));
  jand g27048(.dina(n13217), .dinb(n2511), .dout(n27293));
  jand g27049(.dina(n27293), .dinb(n27292), .dout(n27294));
  jand g27050(.dina(n27294), .dinb(n4807), .dout(n27295));
  jnot g27051(.din(n27295), .dout(n27296));
  jxor g27052(.dina(n27296), .dinb(n27281), .dout(n27297));
  jand g27053(.dina(n22250), .dinb(n732), .dout(n27298));
  jand g27054(.dina(n22248), .dinb(n3855), .dout(n27299));
  jand g27055(.dina(n19758), .dinb(n3858), .dout(n27300));
  jand g27056(.dina(n19510), .dinb(n3851), .dout(n27301));
  jor  g27057(.dina(n27301), .dinb(n27300), .dout(n27302));
  jor  g27058(.dina(n27302), .dinb(n27299), .dout(n27303));
  jor  g27059(.dina(n27303), .dinb(n27298), .dout(n27304));
  jxor g27060(.dina(n27304), .dinb(n27297), .dout(n27305));
  jor  g27061(.dina(n27220), .dinb(n27200), .dout(n27306));
  jand g27062(.dina(n27220), .dinb(n27200), .dout(n27307));
  jor  g27063(.dina(n27228), .dinb(n27307), .dout(n27308));
  jand g27064(.dina(n27308), .dinb(n27306), .dout(n27309));
  jxor g27065(.dina(n27309), .dinb(n27305), .dout(n27310));
  jnot g27066(.din(n27310), .dout(n27311));
  jand g27067(.dina(n22605), .dinb(n4449), .dout(n27312));
  jand g27068(.dina(n22603), .dinb(n4453), .dout(n27313));
  jand g27069(.dina(n22539), .dinb(n4457), .dout(n27314));
  jand g27070(.dina(n22540), .dinb(n4461), .dout(n27315));
  jor  g27071(.dina(n27315), .dinb(n27314), .dout(n27316));
  jor  g27072(.dina(n27316), .dinb(n27313), .dout(n27317));
  jor  g27073(.dina(n27317), .dinb(n27312), .dout(n27318));
  jxor g27074(.dina(n27318), .dinb(n88), .dout(n27319));
  jxor g27075(.dina(n27319), .dinb(n27311), .dout(n27320));
  jor  g27076(.dina(n27229), .dinb(n27195), .dout(n27321));
  jand g27077(.dina(n27229), .dinb(n27195), .dout(n27322));
  jor  g27078(.dina(n27239), .dinb(n27322), .dout(n27323));
  jand g27079(.dina(n27323), .dinb(n27321), .dout(n27324));
  jxor g27080(.dina(n27324), .dinb(n27320), .dout(n27325));
  jor  g27081(.dina(n23708), .dinb(n4747), .dout(n27326));
  jor  g27082(.dina(n23710), .dinb(n4959), .dout(n27327));
  jor  g27083(.dina(n23496), .dinb(n4919), .dout(n27328));
  jor  g27084(.dina(n23450), .dinb(n4746), .dout(n27329));
  jand g27085(.dina(n27329), .dinb(n27328), .dout(n27330));
  jand g27086(.dina(n27330), .dinb(n27327), .dout(n27331));
  jand g27087(.dina(n27331), .dinb(n27326), .dout(n27332));
  jxor g27088(.dina(n27332), .dinb(\a[26] ), .dout(n27333));
  jnot g27089(.din(n27333), .dout(n27334));
  jxor g27090(.dina(n27334), .dinb(n27325), .dout(n27335));
  jxor g27091(.dina(n27335), .dinb(n27277), .dout(n27336));
  jor  g27092(.dina(n24337), .dinb(n5366), .dout(n27337));
  jor  g27093(.dina(n23921), .dinb(n5364), .dout(n27340));
  jand g27094(.dina(n27340), .dinb(n27337), .dout(n27343));
  jxor g27095(.dina(n27343), .dinb(\a[23] ), .dout(n27344));
  jnot g27096(.din(n27344), .dout(n27345));
  jxor g27097(.dina(n27345), .dinb(n27336), .dout(n27346));
  jxor g27098(.dina(n27346), .dinb(n27274), .dout(n27347));
  jxor g27099(.dina(n27347), .dinb(n27271), .dout(n27348));
  jxor g27100(.dina(n27348), .dinb(n27268), .dout(\result[26] ));
  jand g27101(.dina(n27348), .dinb(n27268), .dout(n27350));
  jnot g27102(.din(n72), .dout(n27357));
  jor  g27103(.dina(n27324), .dinb(n27320), .dout(n27358));
  jand g27104(.dina(n27324), .dinb(n27320), .dout(n27359));
  jor  g27105(.dina(n27334), .dinb(n27359), .dout(n27360));
  jand g27106(.dina(n27360), .dinb(n27358), .dout(n27361));
  jxor g27107(.dina(n27361), .dinb(n27357), .dout(n27362));
  jor  g27108(.dina(n23919), .dinb(n4747), .dout(n27363));
  jor  g27109(.dina(n23921), .dinb(n4959), .dout(n27364));
  jor  g27110(.dina(n23710), .dinb(n4919), .dout(n27365));
  jor  g27111(.dina(n23496), .dinb(n4746), .dout(n27366));
  jand g27112(.dina(n27366), .dinb(n27365), .dout(n27367));
  jand g27113(.dina(n27367), .dinb(n27364), .dout(n27368));
  jand g27114(.dina(n27368), .dinb(n27363), .dout(n27369));
  jxor g27115(.dina(n27369), .dinb(\a[26] ), .dout(n27370));
  jnot g27116(.din(n27370), .dout(n27371));
  jand g27117(.dina(n27309), .dinb(n27305), .dout(n27372));
  jnot g27118(.din(n27372), .dout(n27373));
  jor  g27119(.dina(n27319), .dinb(n27311), .dout(n27374));
  jand g27120(.dina(n27374), .dinb(n27373), .dout(n27375));
  jnot g27121(.din(n27375), .dout(n27376));
  jand g27122(.dina(n1185), .dinb(n802), .dout(n27377));
  jand g27123(.dina(n2022), .dinb(n1192), .dout(n27378));
  jand g27124(.dina(n27378), .dinb(n27377), .dout(n27379));
  jand g27125(.dina(n655), .dinb(n441), .dout(n27380));
  jand g27126(.dina(n701), .dinb(n461), .dout(n27381));
  jand g27127(.dina(n27381), .dinb(n27380), .dout(n27382));
  jand g27128(.dina(n2130), .dinb(n1424), .dout(n27383));
  jand g27129(.dina(n27383), .dinb(n27382), .dout(n27384));
  jand g27130(.dina(n14341), .dinb(n12419), .dout(n27385));
  jand g27131(.dina(n27385), .dinb(n27384), .dout(n27386));
  jand g27132(.dina(n27386), .dinb(n27379), .dout(n27387));
  jand g27133(.dina(n25499), .dinb(n22432), .dout(n27388));
  jand g27134(.dina(n27388), .dinb(n27387), .dout(n27389));
  jand g27135(.dina(n27389), .dinb(n20737), .dout(n27390));
  jand g27136(.dina(n27390), .dinb(n4676), .dout(n27391));
  jxor g27137(.dina(n27391), .dinb(n27296), .dout(n27392));
  jand g27138(.dina(n27296), .dinb(n27281), .dout(n27393));
  jnot g27139(.din(n27393), .dout(n27394));
  jnot g27140(.din(n27281), .dout(n27395));
  jand g27141(.dina(n27295), .dinb(n27395), .dout(n27396));
  jor  g27142(.dina(n27304), .dinb(n27396), .dout(n27397));
  jand g27143(.dina(n27397), .dinb(n27394), .dout(n27398));
  jxor g27144(.dina(n27398), .dinb(n27392), .dout(n27399));
  jand g27145(.dina(n22627), .dinb(n732), .dout(n27400));
  jand g27146(.dina(n22540), .dinb(n3855), .dout(n27401));
  jand g27147(.dina(n22248), .dinb(n3858), .dout(n27402));
  jand g27148(.dina(n19758), .dinb(n3851), .dout(n27403));
  jor  g27149(.dina(n27403), .dinb(n27402), .dout(n27404));
  jor  g27150(.dina(n27404), .dinb(n27401), .dout(n27405));
  jor  g27151(.dina(n27405), .dinb(n27400), .dout(n27406));
  jxor g27152(.dina(n27406), .dinb(n27399), .dout(n27407));
  jxor g27153(.dina(n27407), .dinb(n27376), .dout(n27408));
  jnot g27154(.din(n27408), .dout(n27409));
  jand g27155(.dina(n23262), .dinb(n4449), .dout(n27410));
  jand g27156(.dina(n23260), .dinb(n4453), .dout(n27411));
  jand g27157(.dina(n22603), .dinb(n4457), .dout(n27412));
  jand g27158(.dina(n22539), .dinb(n4461), .dout(n27413));
  jor  g27159(.dina(n27413), .dinb(n27412), .dout(n27414));
  jor  g27160(.dina(n27414), .dinb(n27411), .dout(n27415));
  jor  g27161(.dina(n27415), .dinb(n27410), .dout(n27416));
  jxor g27162(.dina(n27416), .dinb(n88), .dout(n27417));
  jxor g27163(.dina(n27417), .dinb(n27409), .dout(n27418));
  jxor g27164(.dina(n27418), .dinb(n27371), .dout(n27419));
  jxor g27165(.dina(n27419), .dinb(n27362), .dout(n27420));
  jor  g27166(.dina(n27335), .dinb(n27277), .dout(n27421));
  jand g27167(.dina(n27335), .dinb(n27277), .dout(n27422));
  jor  g27168(.dina(n27345), .dinb(n27422), .dout(n27423));
  jand g27169(.dina(n27423), .dinb(n27421), .dout(n27424));
  jxor g27170(.dina(n27424), .dinb(n27420), .dout(n27425));
  jand g27171(.dina(n27346), .dinb(n27274), .dout(n27426));
  jand g27172(.dina(n27347), .dinb(n27271), .dout(n27427));
  jor  g27173(.dina(n27427), .dinb(n27426), .dout(n27428));
  jxor g27174(.dina(n27428), .dinb(n27425), .dout(n27429));
  jxor g27175(.dina(n27429), .dinb(n27350), .dout(\result[27] ));
  jand g27176(.dina(n27429), .dinb(n27350), .dout(n27431));
  jand g27177(.dina(n27424), .dinb(n27420), .dout(n27432));
  jand g27178(.dina(n27428), .dinb(n27425), .dout(n27433));
  jor  g27179(.dina(n27433), .dinb(n27432), .dout(n27434));
  jor  g27180(.dina(n27417), .dinb(n27409), .dout(n27435));
  jand g27181(.dina(n27418), .dinb(n27371), .dout(n27436));
  jnot g27182(.din(n27436), .dout(n27437));
  jand g27183(.dina(n27437), .dinb(n27435), .dout(n27438));
  jor  g27184(.dina(n24140), .dinb(n4747), .dout(n27439));
  jor  g27185(.dina(n23921), .dinb(n4919), .dout(n27441));
  jor  g27186(.dina(n23710), .dinb(n4746), .dout(n27442));
  jand g27187(.dina(n27442), .dinb(n27441), .dout(n27443));
  jand g27188(.dina(n27443), .dinb(n27439), .dout(n27445));
  jxor g27189(.dina(n27445), .dinb(\a[26] ), .dout(n27446));
  jxor g27190(.dina(n27446), .dinb(n27438), .dout(n27447));
  jand g27191(.dina(n27406), .dinb(n27399), .dout(n27448));
  jand g27192(.dina(n27407), .dinb(n27376), .dout(n27449));
  jor  g27193(.dina(n27449), .dinb(n27448), .dout(n27450));
  jand g27194(.dina(n27391), .dinb(n27296), .dout(n27451));
  jand g27195(.dina(n27398), .dinb(n27392), .dout(n27452));
  jor  g27196(.dina(n27452), .dinb(n27451), .dout(n27453));
  jand g27197(.dina(n716), .dinb(n371), .dout(n27456));
  jand g27198(.dina(n27456), .dinb(n1285), .dout(n27457));
  jand g27199(.dina(n1997), .dinb(n1057), .dout(n27458));
  jand g27200(.dina(n27458), .dinb(n27457), .dout(n27459));
  jand g27201(.dina(n27459), .dinb(n2366), .dout(n27460));
  jand g27202(.dina(n5748), .dinb(n4366), .dout(n27461));
  jand g27203(.dina(n27461), .dinb(n771), .dout(n27462));
  jand g27204(.dina(n27462), .dinb(n5570), .dout(n27463));
  jand g27205(.dina(n27463), .dinb(n27460), .dout(n27464));
  jand g27206(.dina(n27464), .dinb(n4392), .dout(n27465));
  jand g27207(.dina(n27465), .dinb(n4574), .dout(n27466));
  jand g27208(.dina(n27466), .dinb(n12329), .dout(n27467));
  jxor g27209(.dina(n27467), .dinb(n27391), .dout(n27468));
  jxor g27210(.dina(n27468), .dinb(n72), .dout(n27469));
  jxor g27211(.dina(n27469), .dinb(n27453), .dout(n27470));
  jand g27212(.dina(n22617), .dinb(n732), .dout(n27471));
  jand g27213(.dina(n22539), .dinb(n3855), .dout(n27472));
  jand g27214(.dina(n22540), .dinb(n3858), .dout(n27473));
  jand g27215(.dina(n22248), .dinb(n3851), .dout(n27474));
  jor  g27216(.dina(n27474), .dinb(n27473), .dout(n27475));
  jor  g27217(.dina(n27475), .dinb(n27472), .dout(n27476));
  jor  g27218(.dina(n27476), .dinb(n27471), .dout(n27477));
  jxor g27219(.dina(n27477), .dinb(n27470), .dout(n27478));
  jxor g27220(.dina(n27478), .dinb(n27450), .dout(n27479));
  jor  g27221(.dina(n23494), .dinb(n4724), .dout(n27480));
  jor  g27222(.dina(n23496), .dinb(n4905), .dout(n27481));
  jor  g27223(.dina(n23450), .dinb(n4735), .dout(n27482));
  jor  g27224(.dina(n23449), .dinb(n4733), .dout(n27483));
  jand g27225(.dina(n27483), .dinb(n27482), .dout(n27484));
  jand g27226(.dina(n27484), .dinb(n27481), .dout(n27485));
  jand g27227(.dina(n27485), .dinb(n27480), .dout(n27486));
  jxor g27228(.dina(n27486), .dinb(\a[29] ), .dout(n27487));
  jnot g27229(.din(n27487), .dout(n27488));
  jxor g27230(.dina(n27488), .dinb(n27479), .dout(n27489));
  jxor g27231(.dina(n27489), .dinb(n27447), .dout(n27490));
  jor  g27232(.dina(n27361), .dinb(n27357), .dout(n27491));
  jand g27233(.dina(n27361), .dinb(n27357), .dout(n27492));
  jor  g27234(.dina(n27419), .dinb(n27492), .dout(n27493));
  jand g27235(.dina(n27493), .dinb(n27491), .dout(n27494));
  jxor g27236(.dina(n27494), .dinb(n27490), .dout(n27495));
  jxor g27237(.dina(n27495), .dinb(n27434), .dout(n27496));
  jxor g27238(.dina(n27496), .dinb(n27431), .dout(\result[28] ));
  jand g27239(.dina(n27496), .dinb(n27431), .dout(n27498));
  jand g27240(.dina(n27494), .dinb(n27490), .dout(n27499));
  jand g27241(.dina(n27495), .dinb(n27434), .dout(n27500));
  jor  g27242(.dina(n27500), .dinb(n27499), .dout(n27501));
  jnot g27243(.din(n27438), .dout(n27502));
  jnot g27244(.din(n27446), .dout(n27503));
  jand g27245(.dina(n27503), .dinb(n27502), .dout(n27504));
  jand g27246(.dina(n27489), .dinb(n27447), .dout(n27505));
  jor  g27247(.dina(n27505), .dinb(n27504), .dout(n27506));
  jor  g27248(.dina(n27467), .dinb(n27391), .dout(n27507));
  jand g27249(.dina(n27468), .dinb(n72), .dout(n27508));
  jnot g27250(.din(n27508), .dout(n27509));
  jand g27251(.dina(n27509), .dinb(n27507), .dout(n27510));
  jand g27252(.dina(n2565), .dinb(n277), .dout(n27511));
  jand g27253(.dina(n2301), .dinb(n883), .dout(n27512));
  jand g27254(.dina(n27512), .dinb(n27511), .dout(n27513));
  jand g27255(.dina(n486), .dinb(n476), .dout(n27514));
  jand g27256(.dina(n801), .dinb(n249), .dout(n27515));
  jand g27257(.dina(n27515), .dinb(n27514), .dout(n27516));
  jand g27258(.dina(n27516), .dinb(n13600), .dout(n27517));
  jand g27259(.dina(n27517), .dinb(n27513), .dout(n27518));
  jand g27260(.dina(n2769), .dinb(n355), .dout(n27519));
  jand g27261(.dina(n27519), .dinb(n2663), .dout(n27520));
  jand g27262(.dina(n27520), .dinb(n7117), .dout(n27521));
  jand g27263(.dina(n27521), .dinb(n27518), .dout(n27522));
  jand g27264(.dina(n27522), .dinb(n4381), .dout(n27523));
  jand g27265(.dina(n27523), .dinb(n4340), .dout(n27524));
  jand g27266(.dina(n27524), .dinb(n14323), .dout(n27525));
  jand g27267(.dina(n27525), .dinb(n22578), .dout(n27526));
  jnot g27268(.din(n27526), .dout(n27527));
  jxor g27269(.dina(n27527), .dinb(n27510), .dout(n27528));
  jand g27270(.dina(n22605), .dinb(n732), .dout(n27529));
  jand g27271(.dina(n22603), .dinb(n3855), .dout(n27530));
  jand g27272(.dina(n22539), .dinb(n3858), .dout(n27531));
  jand g27273(.dina(n22540), .dinb(n3851), .dout(n27532));
  jor  g27274(.dina(n27532), .dinb(n27531), .dout(n27533));
  jor  g27275(.dina(n27533), .dinb(n27530), .dout(n27534));
  jor  g27276(.dina(n27534), .dinb(n27529), .dout(n27535));
  jxor g27277(.dina(n27535), .dinb(n27528), .dout(n27536));
  jor  g27278(.dina(n27469), .dinb(n27453), .dout(n27537));
  jand g27279(.dina(n27469), .dinb(n27453), .dout(n27538));
  jor  g27280(.dina(n27477), .dinb(n27538), .dout(n27539));
  jand g27281(.dina(n27539), .dinb(n27537), .dout(n27540));
  jxor g27282(.dina(n27540), .dinb(n27536), .dout(n27541));
  jnot g27283(.din(n27541), .dout(n27542));
  jor  g27284(.dina(n23708), .dinb(n4724), .dout(n27543));
  jor  g27285(.dina(n23710), .dinb(n4905), .dout(n27544));
  jor  g27286(.dina(n23496), .dinb(n4735), .dout(n27545));
  jor  g27287(.dina(n23450), .dinb(n4733), .dout(n27546));
  jand g27288(.dina(n27546), .dinb(n27545), .dout(n27547));
  jand g27289(.dina(n27547), .dinb(n27544), .dout(n27548));
  jand g27290(.dina(n27548), .dinb(n27543), .dout(n27549));
  jxor g27291(.dina(n27549), .dinb(\a[29] ), .dout(n27550));
  jxor g27292(.dina(n27550), .dinb(n27542), .dout(n27551));
  jor  g27293(.dina(n27478), .dinb(n27450), .dout(n27552));
  jand g27294(.dina(n27478), .dinb(n27450), .dout(n27553));
  jor  g27295(.dina(n27488), .dinb(n27553), .dout(n27554));
  jand g27296(.dina(n27554), .dinb(n27552), .dout(n27555));
  jxor g27297(.dina(n27555), .dinb(n27551), .dout(n27556));
  jor  g27298(.dina(n24337), .dinb(n4747), .dout(n27557));
  jor  g27299(.dina(n23921), .dinb(n4746), .dout(n27560));
  jand g27300(.dina(n27560), .dinb(n27557), .dout(n27563));
  jxor g27301(.dina(n27563), .dinb(\a[26] ), .dout(n27564));
  jnot g27302(.din(n27564), .dout(n27565));
  jxor g27303(.dina(n27565), .dinb(n27556), .dout(n27566));
  jxor g27304(.dina(n27566), .dinb(n27506), .dout(n27567));
  jxor g27305(.dina(n27567), .dinb(n27501), .dout(n27568));
  jxor g27306(.dina(n27568), .dinb(n27498), .dout(\result[29] ));
  jand g27307(.dina(n27568), .dinb(n27498), .dout(n27570));
  jand g27308(.dina(n27566), .dinb(n27506), .dout(n27571));
  jand g27309(.dina(n27567), .dinb(n27501), .dout(n27572));
  jor  g27310(.dina(n27572), .dinb(n27571), .dout(n27573));
  jand g27311(.dina(n27540), .dinb(n27536), .dout(n27574));
  jnot g27312(.din(n27574), .dout(n27575));
  jor  g27313(.dina(n27550), .dinb(n27542), .dout(n27576));
  jand g27314(.dina(n27576), .dinb(n27575), .dout(n27577));
  jnot g27315(.din(n27577), .dout(n27578));
  jand g27316(.dina(n12316), .dinb(n4563), .dout(n27579));
  jand g27317(.dina(n27579), .dinb(n3038), .dout(n27580));
  jand g27318(.dina(n4413), .dinb(n4398), .dout(n27581));
  jand g27319(.dina(n27581), .dinb(n4594), .dout(n27582));
  jand g27320(.dina(n27582), .dinb(n27580), .dout(n27583));
  jand g27321(.dina(n27583), .dinb(n22578), .dout(n27584));
  jxor g27322(.dina(n27584), .dinb(n27527), .dout(n27585));
  jand g27323(.dina(n27527), .dinb(n27510), .dout(n27586));
  jnot g27324(.din(n27586), .dout(n27587));
  jnot g27325(.din(n27510), .dout(n27588));
  jand g27326(.dina(n27526), .dinb(n27588), .dout(n27589));
  jor  g27327(.dina(n27535), .dinb(n27589), .dout(n27590));
  jand g27328(.dina(n27590), .dinb(n27587), .dout(n27591));
  jxor g27329(.dina(n27591), .dinb(n27585), .dout(n27592));
  jand g27330(.dina(n23262), .dinb(n732), .dout(n27593));
  jand g27331(.dina(n23260), .dinb(n3855), .dout(n27594));
  jand g27332(.dina(n22603), .dinb(n3858), .dout(n27595));
  jand g27333(.dina(n22539), .dinb(n3851), .dout(n27596));
  jor  g27334(.dina(n27596), .dinb(n27595), .dout(n27597));
  jor  g27335(.dina(n27597), .dinb(n27594), .dout(n27598));
  jor  g27336(.dina(n27598), .dinb(n27593), .dout(n27599));
  jxor g27337(.dina(n27599), .dinb(n27592), .dout(n27600));
  jxor g27338(.dina(n27600), .dinb(n27578), .dout(n27601));
  jor  g27339(.dina(n23919), .dinb(n4724), .dout(n27608));
  jor  g27340(.dina(n23921), .dinb(n4905), .dout(n27609));
  jor  g27341(.dina(n23710), .dinb(n4735), .dout(n27610));
  jor  g27342(.dina(n23496), .dinb(n4733), .dout(n27611));
  jand g27343(.dina(n27611), .dinb(n27610), .dout(n27612));
  jand g27344(.dina(n27612), .dinb(n27609), .dout(n27613));
  jand g27345(.dina(n27613), .dinb(n27608), .dout(n27614));
  jxor g27346(.dina(n27614), .dinb(\a[29] ), .dout(n27615));
  jxor g27347(.dina(n27615), .dinb(n68), .dout(n27616));
  jxor g27348(.dina(n27616), .dinb(n27601), .dout(n27617));
  jor  g27349(.dina(n27555), .dinb(n27551), .dout(n27618));
  jand g27350(.dina(n27555), .dinb(n27551), .dout(n27619));
  jor  g27351(.dina(n27565), .dinb(n27619), .dout(n27620));
  jand g27352(.dina(n27620), .dinb(n27618), .dout(n27621));
  jxor g27353(.dina(n27621), .dinb(n27617), .dout(n27622));
  jxor g27354(.dina(n27622), .dinb(n27573), .dout(n27623));
  jxor g27355(.dina(n27623), .dinb(n27570), .dout(\result[30] ));
  jand g27356(.dina(n27623), .dinb(n27570), .dout(n27625));
  jand g27357(.dina(n24593), .dinb(n22575), .dout(n27626));
  jxor g27358(.dina(n27626), .dinb(n27625), .dout(n27627));
  jand g27359(.dina(n27621), .dinb(n27617), .dout(n27628));
  jand g27360(.dina(n27622), .dinb(n27573), .dout(n27629));
  jor  g27361(.dina(n27629), .dinb(n27628), .dout(n27630));
  jor  g27362(.dina(n27615), .dinb(n68), .dout(n27631));
  jnot g27363(.din(n27601), .dout(n27632));
  jnot g27364(.din(n27616), .dout(n27633));
  jor  g27365(.dina(n27633), .dinb(n27632), .dout(n27634));
  jand g27366(.dina(n27634), .dinb(n27631), .dout(n27635));
  jxor g27367(.dina(n27635), .dinb(n27630), .dout(n27636));
  jxor g27368(.dina(n27636), .dinb(n27527), .dout(n27637));
  jand g27369(.dina(n4628), .dinb(n4583), .dout(n27638));
  jxor g27370(.dina(n27638), .dinb(\a[26] ), .dout(n27639));
  jand g27371(.dina(n27599), .dinb(n27592), .dout(n27640));
  jand g27372(.dina(n27600), .dinb(n27578), .dout(n27641));
  jor  g27373(.dina(n27641), .dinb(n27640), .dout(n27642));
  jor  g27374(.dina(n27584), .dinb(n27527), .dout(n27643));
  jnot g27375(.din(n27585), .dout(n27644));
  jnot g27376(.din(n27591), .dout(n27645));
  jor  g27377(.dina(n27645), .dinb(n27644), .dout(n27646));
  jand g27378(.dina(n27646), .dinb(n27643), .dout(n27647));
  jxor g27379(.dina(n27647), .dinb(n27642), .dout(n27648));
  jor  g27380(.dina(n24140), .dinb(n4724), .dout(n27649));
  jor  g27381(.dina(n24142), .dinb(n4905), .dout(n27650));
  jor  g27382(.dina(n23921), .dinb(n4735), .dout(n27651));
  jor  g27383(.dina(n23710), .dinb(n4733), .dout(n27652));
  jand g27384(.dina(n27652), .dinb(n27651), .dout(n27653));
  jand g27385(.dina(n27653), .dinb(n27650), .dout(n27654));
  jand g27386(.dina(n27654), .dinb(n27649), .dout(n27655));
  jxor g27387(.dina(n27655), .dinb(\a[29] ), .dout(n27656));
  jor  g27388(.dina(n23494), .dinb(n6463), .dout(n27657));
  jor  g27389(.dina(n23496), .dinb(n3854), .dout(n27658));
  jor  g27390(.dina(n23450), .dinb(n24120), .dout(n27659));
  jnot g27391(.din(n3851), .dout(n27660));
  jor  g27392(.dina(n23449), .dinb(n27660), .dout(n27661));
  jand g27393(.dina(n27661), .dinb(n27659), .dout(n27662));
  jand g27394(.dina(n27662), .dinb(n27658), .dout(n27663));
  jand g27395(.dina(n27663), .dinb(n27657), .dout(n27664));
  jxor g27396(.dina(n27664), .dinb(n27656), .dout(n27665));
  jxor g27397(.dina(n27665), .dinb(n27648), .dout(n27666));
  jxor g27398(.dina(n27666), .dinb(n27639), .dout(n27667));
  jxor g27399(.dina(n27667), .dinb(n27637), .dout(n27668));
  jxor g27400(.dina(n27668), .dinb(n27627), .dout(\result[31] ));
endmodule


