// Benchmark "c5315" written by ABC on Wed May 27 22:05:51 2020

module gf_c5315 ( 
    G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
    G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
    G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
    G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140,
    G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173,
    G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209,
    G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251,
    G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293,
    G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338,
    G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389,
    G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523,
    G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691,
    G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717,
    G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34,
    G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76,
    G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103,
    G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
    G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137,
    G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170,
    G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206,
    G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248,
    G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292,
    G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335,
    G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386,
    G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514,
    G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690,
    G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552,
    G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire n314, n316, n318, n320, n321, n325, n326, n327, n328, n329, n330,
    n332, n333, n334, n335, n336, n338, n340, n341, n342, n343, n345, n346,
    n347, n348, n350, n351, n352, n353, n355, n356, n357, n358, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n611, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n663, n664, n665,
    n666, n667, n668, n669, n670, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n776, n777, n778, n779,
    n780, n781, n782, n783, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n810, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n831, n833, n834, n835, n836, n837, n838, n839, n840, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n877, n878, n879, n880, n881, n882, n883,
    n884, n886, n887, n888, n889, n890, n891, n892, n893, n894, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
    n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1215, n1216, n1217, n1218, n1219, n1220, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1238, n1239, n1240, n1241, n1242, n1243, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1253, n1254, n1255, n1256,
    n1257, n1258, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1308, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1360, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1389, n1390, n1391,
    n1392, n1393, n1394, n1395, n1396, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
    n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717;
  jnot g0000(.din(G545), .dout(G594));
  jnot g0001(.din(G348), .dout(G599));
  jnot g0002(.din(G366), .dout(G600));
  jand g0003(.dina(G562), .dinb(G552), .dout(G601));
  jnot g0004(.din(G549), .dout(G602));
  jnot g0005(.din(G338), .dout(G611));
  jnot g0006(.din(G358), .dout(G612));
  jand g0007(.dina(G145), .dinb(G141), .dout(G810));
  jnot g0008(.din(G245), .dout(G848));
  jnot g0009(.din(G552), .dout(G849));
  jnot g0010(.din(G562), .dout(G850));
  jnot g0011(.din(G559), .dout(G851));
  jand g0012(.dina(G373), .dinb(G1), .dout(G634));
  jnot g0013(.din(G3173), .dout(n314));
  jand g0014(.dina(n314), .dinb(G136), .dout(G815));
  jnot g0015(.din(G27), .dout(n316));
  jor  g0016(.dina(G2824), .dinb(n316), .dout(G845));
  jand g0017(.dina(G556), .dinb(G386), .dout(n318));
  jnot g0018(.din(n318), .dout(G847));
  jnot g0019(.din(G140), .dout(n320));
  jnot g0020(.din(G31), .dout(n321));
  jor  g0021(.dina(n321), .dinb(n316), .dout(G809));
  jor  g0022(.dina(G809), .dinb(n320), .dout(G656));
  jnot g0023(.din(G299), .dout(G593));
  jnot g0024(.din(G86), .dout(n325));
  jnot g0025(.din(G2358), .dout(n326));
  jand g0026(.dina(n326), .dinb(n325), .dout(n327));
  jnot g0027(.din(G87), .dout(n328));
  jand g0028(.dina(G2358), .dinb(n328), .dout(n329));
  jor  g0029(.dina(n329), .dinb(G809), .dout(n330));
  jor  g0030(.dina(n330), .dinb(n327), .dout(G636));
  jnot g0031(.din(G88), .dout(n332));
  jand g0032(.dina(n326), .dinb(n332), .dout(n333));
  jnot g0033(.din(G34), .dout(n334));
  jand g0034(.dina(G2358), .dinb(n334), .dout(n335));
  jor  g0035(.dina(n335), .dinb(G809), .dout(n336));
  jor  g0036(.dina(n336), .dinb(n333), .dout(G704));
  jnot g0037(.din(G83), .dout(n338));
  jor  g0038(.dina(G809), .dinb(n338), .dout(G820));
  jand g0039(.dina(n326), .dinb(G24), .dout(n340));
  jand g0040(.dina(G2358), .dinb(G25), .dout(n341));
  jor  g0041(.dina(n341), .dinb(G809), .dout(n342));
  jor  g0042(.dina(n342), .dinb(n340), .dout(n343));
  jand g0043(.dina(n343), .dinb(G141), .dout(G639));
  jand g0044(.dina(n326), .dinb(G26), .dout(n345));
  jand g0045(.dina(G2358), .dinb(G81), .dout(n346));
  jor  g0046(.dina(n346), .dinb(G809), .dout(n347));
  jor  g0047(.dina(n347), .dinb(n345), .dout(n348));
  jand g0048(.dina(n348), .dinb(G141), .dout(G673));
  jand g0049(.dina(n326), .dinb(G79), .dout(n350));
  jand g0050(.dina(G2358), .dinb(G23), .dout(n351));
  jor  g0051(.dina(n351), .dinb(G809), .dout(n352));
  jor  g0052(.dina(n352), .dinb(n350), .dout(n353));
  jand g0053(.dina(n353), .dinb(G141), .dout(G707));
  jand g0054(.dina(G2358), .dinb(G80), .dout(n355));
  jand g0055(.dina(n326), .dinb(G82), .dout(n356));
  jor  g0056(.dina(n356), .dinb(G809), .dout(n357));
  jor  g0057(.dina(n357), .dinb(n355), .dout(n358));
  jand g0058(.dina(n358), .dinb(G141), .dout(G715));
  jand g0059(.dina(G3552), .dinb(G514), .dout(n360));
  jnot g0060(.din(G514), .dout(n361));
  jnot g0061(.din(G3546), .dout(n362));
  jand g0062(.dina(n362), .dinb(n361), .dout(n363));
  jor  g0063(.dina(n363), .dinb(n360), .dout(n364));
  jnot g0064(.din(n364), .dout(n365));
  jnot g0065(.din(G251), .dout(n366));
  jnot g0066(.din(G361), .dout(n367));
  jand g0067(.dina(n367), .dinb(n366), .dout(n368));
  jnot g0068(.din(G248), .dout(n369));
  jand g0069(.dina(G361), .dinb(n369), .dout(n370));
  jor  g0070(.dina(n370), .dinb(n368), .dout(n371));
  jnot g0071(.din(n371), .dout(n372));
  jand g0072(.dina(n372), .dinb(n365), .dout(n373));
  jnot g0073(.din(G351), .dout(n374));
  jnot g0074(.din(G3550), .dout(n375));
  jand g0075(.dina(n375), .dinb(n374), .dout(n376));
  jnot g0076(.din(G534), .dout(n377));
  jnot g0077(.din(G3552), .dout(n378));
  jand g0078(.dina(n378), .dinb(G351), .dout(n379));
  jor  g0079(.dina(n379), .dinb(n377), .dout(n380));
  jor  g0080(.dina(n380), .dinb(n376), .dout(n381));
  jand g0081(.dina(G3546), .dinb(G351), .dout(n382));
  jand g0082(.dina(G3548), .dinb(n374), .dout(n383));
  jor  g0083(.dina(n383), .dinb(n382), .dout(n384));
  jor  g0084(.dina(n384), .dinb(G534), .dout(n385));
  jand g0085(.dina(n385), .dinb(n381), .dout(n386));
  jnot g0086(.din(G341), .dout(n387));
  jand g0087(.dina(n375), .dinb(n387), .dout(n388));
  jnot g0088(.din(G523), .dout(n389));
  jand g0089(.dina(n378), .dinb(G341), .dout(n390));
  jor  g0090(.dina(n390), .dinb(n389), .dout(n391));
  jor  g0091(.dina(n391), .dinb(n388), .dout(n392));
  jand g0092(.dina(G3546), .dinb(G341), .dout(n393));
  jand g0093(.dina(G3548), .dinb(n387), .dout(n394));
  jor  g0094(.dina(n394), .dinb(n393), .dout(n395));
  jor  g0095(.dina(n395), .dinb(G523), .dout(n396));
  jand g0096(.dina(n396), .dinb(n392), .dout(n397));
  jand g0097(.dina(n397), .dinb(n386), .dout(n398));
  jand g0098(.dina(n398), .dinb(n373), .dout(n399));
  jand g0099(.dina(G316), .dinb(G248), .dout(n400));
  jnot g0100(.din(G490), .dout(n401));
  jnot g0101(.din(G316), .dout(n402));
  jand g0102(.dina(n402), .dinb(G251), .dout(n403));
  jor  g0103(.dina(n403), .dinb(n401), .dout(n404));
  jor  g0104(.dina(n404), .dinb(n400), .dout(n405));
  jnot g0105(.din(G254), .dout(n406));
  jand g0106(.dina(n402), .dinb(n406), .dout(n407));
  jnot g0107(.din(G242), .dout(n408));
  jand g0108(.dina(G316), .dinb(n408), .dout(n409));
  jor  g0109(.dina(n409), .dinb(n407), .dout(n410));
  jor  g0110(.dina(n410), .dinb(G490), .dout(n411));
  jand g0111(.dina(n411), .dinb(n405), .dout(n412));
  jand g0112(.dina(G308), .dinb(G248), .dout(n413));
  jnot g0113(.din(G479), .dout(n414));
  jnot g0114(.din(G308), .dout(n415));
  jand g0115(.dina(n415), .dinb(G251), .dout(n416));
  jor  g0116(.dina(n416), .dinb(n414), .dout(n417));
  jor  g0117(.dina(n417), .dinb(n413), .dout(n418));
  jand g0118(.dina(n415), .dinb(n406), .dout(n419));
  jand g0119(.dina(G308), .dinb(n408), .dout(n420));
  jor  g0120(.dina(n420), .dinb(n419), .dout(n421));
  jor  g0121(.dina(n421), .dinb(G479), .dout(n422));
  jand g0122(.dina(n422), .dinb(n418), .dout(n423));
  jand g0123(.dina(n423), .dinb(n412), .dout(n424));
  jnot g0124(.din(G293), .dout(n425));
  jand g0125(.dina(n425), .dinb(n406), .dout(n426));
  jand g0126(.dina(G293), .dinb(n408), .dout(n427));
  jor  g0127(.dina(n427), .dinb(n426), .dout(n428));
  jnot g0128(.din(G302), .dout(n429));
  jand g0129(.dina(n429), .dinb(n366), .dout(n430));
  jand g0130(.dina(G302), .dinb(n369), .dout(n431));
  jor  g0131(.dina(n431), .dinb(n430), .dout(n432));
  jnot g0132(.din(n432), .dout(n433));
  jand g0133(.dina(n433), .dinb(n428), .dout(n434));
  jnot g0134(.din(G324), .dout(n435));
  jand g0135(.dina(n375), .dinb(n435), .dout(n436));
  jnot g0136(.din(G503), .dout(n437));
  jand g0137(.dina(n378), .dinb(G324), .dout(n438));
  jor  g0138(.dina(n438), .dinb(n437), .dout(n439));
  jor  g0139(.dina(n439), .dinb(n436), .dout(n440));
  jand g0140(.dina(G3546), .dinb(G324), .dout(n441));
  jand g0141(.dina(G3548), .dinb(n435), .dout(n442));
  jor  g0142(.dina(n442), .dinb(n441), .dout(n443));
  jor  g0143(.dina(n443), .dinb(G503), .dout(n444));
  jand g0144(.dina(n444), .dinb(n440), .dout(n445));
  jand g0145(.dina(n445), .dinb(n434), .dout(n446));
  jand g0146(.dina(n446), .dinb(n424), .dout(n447));
  jand g0147(.dina(n447), .dinb(n399), .dout(G598));
  jnot g0148(.din(G210), .dout(n449));
  jand g0149(.dina(n375), .dinb(n449), .dout(n450));
  jnot g0150(.din(G457), .dout(n451));
  jand g0151(.dina(n378), .dinb(G210), .dout(n452));
  jor  g0152(.dina(n452), .dinb(n451), .dout(n453));
  jor  g0153(.dina(n453), .dinb(n450), .dout(n454));
  jand g0154(.dina(G3546), .dinb(G210), .dout(n455));
  jand g0155(.dina(G3548), .dinb(n449), .dout(n456));
  jor  g0156(.dina(n456), .dinb(n455), .dout(n457));
  jor  g0157(.dina(n457), .dinb(G457), .dout(n458));
  jand g0158(.dina(n458), .dinb(n454), .dout(n459));
  jnot g0159(.din(G234), .dout(n460));
  jand g0160(.dina(n375), .dinb(n460), .dout(n461));
  jnot g0161(.din(G435), .dout(n462));
  jand g0162(.dina(n378), .dinb(G234), .dout(n463));
  jor  g0163(.dina(n463), .dinb(n462), .dout(n464));
  jor  g0164(.dina(n464), .dinb(n461), .dout(n465));
  jand g0165(.dina(G3546), .dinb(G234), .dout(n466));
  jand g0166(.dina(G3548), .dinb(n460), .dout(n467));
  jor  g0167(.dina(n467), .dinb(n466), .dout(n468));
  jor  g0168(.dina(n468), .dinb(G435), .dout(n469));
  jand g0169(.dina(n469), .dinb(n465), .dout(n470));
  jnot g0170(.din(G273), .dout(n471));
  jand g0171(.dina(n375), .dinb(n471), .dout(n472));
  jnot g0172(.din(G411), .dout(n473));
  jand g0173(.dina(n378), .dinb(G273), .dout(n474));
  jor  g0174(.dina(n474), .dinb(n473), .dout(n475));
  jor  g0175(.dina(n475), .dinb(n472), .dout(n476));
  jand g0176(.dina(G3546), .dinb(G273), .dout(n477));
  jand g0177(.dina(G3548), .dinb(n471), .dout(n478));
  jor  g0178(.dina(n478), .dinb(n477), .dout(n479));
  jor  g0179(.dina(n479), .dinb(G411), .dout(n480));
  jand g0180(.dina(n480), .dinb(n476), .dout(n481));
  jand g0181(.dina(n481), .dinb(n470), .dout(n482));
  jnot g0182(.din(G265), .dout(n483));
  jand g0183(.dina(n375), .dinb(n483), .dout(n484));
  jnot g0184(.din(G400), .dout(n485));
  jand g0185(.dina(n378), .dinb(G265), .dout(n486));
  jor  g0186(.dina(n486), .dinb(n485), .dout(n487));
  jor  g0187(.dina(n487), .dinb(n484), .dout(n488));
  jand g0188(.dina(G3546), .dinb(G265), .dout(n489));
  jand g0189(.dina(G3548), .dinb(n483), .dout(n490));
  jor  g0190(.dina(n490), .dinb(n489), .dout(n491));
  jor  g0191(.dina(n491), .dinb(G400), .dout(n492));
  jand g0192(.dina(n492), .dinb(n488), .dout(n493));
  jnot g0193(.din(G226), .dout(n494));
  jand g0194(.dina(n375), .dinb(n494), .dout(n495));
  jnot g0195(.din(G422), .dout(n496));
  jand g0196(.dina(n378), .dinb(G226), .dout(n497));
  jor  g0197(.dina(n497), .dinb(n496), .dout(n498));
  jor  g0198(.dina(n498), .dinb(n495), .dout(n499));
  jand g0199(.dina(G3546), .dinb(G226), .dout(n500));
  jand g0200(.dina(G3548), .dinb(n494), .dout(n501));
  jor  g0201(.dina(n501), .dinb(n500), .dout(n502));
  jor  g0202(.dina(n502), .dinb(G422), .dout(n503));
  jand g0203(.dina(n503), .dinb(n499), .dout(n504));
  jand g0204(.dina(n504), .dinb(n493), .dout(n505));
  jand g0205(.dina(n505), .dinb(n482), .dout(n506));
  jnot g0206(.din(G218), .dout(n507));
  jand g0207(.dina(n375), .dinb(n507), .dout(n508));
  jnot g0208(.din(G468), .dout(n509));
  jand g0209(.dina(n378), .dinb(G218), .dout(n510));
  jor  g0210(.dina(n510), .dinb(n509), .dout(n511));
  jor  g0211(.dina(n511), .dinb(n508), .dout(n512));
  jand g0212(.dina(G3546), .dinb(G218), .dout(n513));
  jand g0213(.dina(G3548), .dinb(n507), .dout(n514));
  jor  g0214(.dina(n514), .dinb(n513), .dout(n515));
  jor  g0215(.dina(n515), .dinb(G468), .dout(n516));
  jand g0216(.dina(n516), .dinb(n512), .dout(n517));
  jnot g0217(.din(G257), .dout(n518));
  jand g0218(.dina(n375), .dinb(n518), .dout(n519));
  jnot g0219(.din(G389), .dout(n520));
  jand g0220(.dina(n378), .dinb(G257), .dout(n521));
  jor  g0221(.dina(n521), .dinb(n520), .dout(n522));
  jor  g0222(.dina(n522), .dinb(n519), .dout(n523));
  jand g0223(.dina(G3546), .dinb(G257), .dout(n524));
  jand g0224(.dina(G3548), .dinb(n518), .dout(n525));
  jor  g0225(.dina(n525), .dinb(n524), .dout(n526));
  jor  g0226(.dina(n526), .dinb(G389), .dout(n527));
  jand g0227(.dina(n527), .dinb(n523), .dout(n528));
  jand g0228(.dina(n528), .dinb(n517), .dout(n529));
  jnot g0229(.din(G281), .dout(n530));
  jand g0230(.dina(n375), .dinb(n530), .dout(n531));
  jnot g0231(.din(G374), .dout(n532));
  jand g0232(.dina(n378), .dinb(G281), .dout(n533));
  jor  g0233(.dina(n533), .dinb(n532), .dout(n534));
  jor  g0234(.dina(n534), .dinb(n531), .dout(n535));
  jand g0235(.dina(G3546), .dinb(G281), .dout(n536));
  jand g0236(.dina(G3548), .dinb(n530), .dout(n537));
  jor  g0237(.dina(n537), .dinb(n536), .dout(n538));
  jor  g0238(.dina(n538), .dinb(G374), .dout(n539));
  jand g0239(.dina(n539), .dinb(n535), .dout(n540));
  jand g0240(.dina(G248), .dinb(G206), .dout(n541));
  jnot g0241(.din(G446), .dout(n542));
  jnot g0242(.din(G206), .dout(n543));
  jand g0243(.dina(G251), .dinb(n543), .dout(n544));
  jor  g0244(.dina(n544), .dinb(n542), .dout(n545));
  jor  g0245(.dina(n545), .dinb(n541), .dout(n546));
  jand g0246(.dina(n406), .dinb(n543), .dout(n547));
  jand g0247(.dina(n408), .dinb(G206), .dout(n548));
  jor  g0248(.dina(n548), .dinb(n547), .dout(n549));
  jor  g0249(.dina(n549), .dinb(G446), .dout(n550));
  jand g0250(.dina(n550), .dinb(n546), .dout(n551));
  jand g0251(.dina(n551), .dinb(n540), .dout(n552));
  jand g0252(.dina(n552), .dinb(n529), .dout(n553));
  jand g0253(.dina(n553), .dinb(n506), .dout(n554));
  jand g0254(.dina(n554), .dinb(n459), .dout(G610));
  jnot g0255(.din(G335), .dout(n556));
  jand g0256(.dina(n556), .dinb(n530), .dout(n557));
  jnot g0257(.din(n557), .dout(n558));
  jor  g0258(.dina(n556), .dinb(G288), .dout(n559));
  jand g0259(.dina(n559), .dinb(n558), .dout(n560));
  jxor g0260(.dina(n560), .dinb(G374), .dout(n561));
  jand g0261(.dina(n556), .dinb(n471), .dout(n562));
  jnot g0262(.din(n562), .dout(n563));
  jor  g0263(.dina(n556), .dinb(G280), .dout(n564));
  jand g0264(.dina(n564), .dinb(n563), .dout(n565));
  jxor g0265(.dina(n565), .dinb(G411), .dout(n566));
  jand g0266(.dina(n566), .dinb(n561), .dout(n567));
  jnot g0267(.din(n567), .dout(n568));
  jand g0268(.dina(n556), .dinb(n483), .dout(n569));
  jnot g0269(.din(n569), .dout(n570));
  jor  g0270(.dina(n556), .dinb(G272), .dout(n571));
  jand g0271(.dina(n571), .dinb(n570), .dout(n572));
  jxor g0272(.dina(n572), .dinb(G400), .dout(n573));
  jnot g0273(.din(n573), .dout(n574));
  jand g0274(.dina(n556), .dinb(n518), .dout(n575));
  jnot g0275(.din(n575), .dout(n576));
  jor  g0276(.dina(n556), .dinb(G264), .dout(n577));
  jand g0277(.dina(n577), .dinb(n576), .dout(n578));
  jxor g0278(.dina(n578), .dinb(n520), .dout(n579));
  jor  g0279(.dina(n579), .dinb(n574), .dout(n580));
  jor  g0280(.dina(n580), .dinb(n568), .dout(n581));
  jnot g0281(.din(n581), .dout(n582));
  jand g0282(.dina(n556), .dinb(n460), .dout(n583));
  jnot g0283(.din(n583), .dout(n584));
  jor  g0284(.dina(n556), .dinb(G241), .dout(n585));
  jand g0285(.dina(n585), .dinb(n584), .dout(n586));
  jxor g0286(.dina(n586), .dinb(G435), .dout(n587));
  jand g0287(.dina(n587), .dinb(n582), .dout(n588));
  jor  g0288(.dina(G335), .dinb(G206), .dout(n589));
  jor  g0289(.dina(n556), .dinb(G209), .dout(n590));
  jand g0290(.dina(n590), .dinb(n589), .dout(n591));
  jxor g0291(.dina(n591), .dinb(G446), .dout(n592));
  jand g0292(.dina(n556), .dinb(n494), .dout(n593));
  jnot g0293(.din(n593), .dout(n594));
  jor  g0294(.dina(n556), .dinb(G233), .dout(n595));
  jand g0295(.dina(n595), .dinb(n594), .dout(n596));
  jxor g0296(.dina(n596), .dinb(n496), .dout(n597));
  jand g0297(.dina(n556), .dinb(n507), .dout(n598));
  jnot g0298(.din(n598), .dout(n599));
  jor  g0299(.dina(n556), .dinb(G225), .dout(n600));
  jand g0300(.dina(n600), .dinb(n599), .dout(n601));
  jxor g0301(.dina(n601), .dinb(n509), .dout(n602));
  jor  g0302(.dina(n602), .dinb(n597), .dout(n603));
  jand g0303(.dina(n556), .dinb(n449), .dout(n604));
  jnot g0304(.din(n604), .dout(n605));
  jor  g0305(.dina(n556), .dinb(G217), .dout(n606));
  jand g0306(.dina(n606), .dinb(n605), .dout(n607));
  jxor g0307(.dina(n607), .dinb(n451), .dout(n608));
  jor  g0308(.dina(n608), .dinb(n603), .dout(n609));
  jnot g0309(.din(n609), .dout(n610));
  jand g0310(.dina(n610), .dinb(n592), .dout(n611));
  jand g0311(.dina(n611), .dinb(n588), .dout(G588));
  jnot g0312(.din(G332), .dout(n613));
  jand g0313(.dina(n613), .dinb(n435), .dout(n614));
  jnot g0314(.din(n614), .dout(n615));
  jor  g0315(.dina(n613), .dinb(G331), .dout(n616));
  jand g0316(.dina(n616), .dinb(n615), .dout(n617));
  jxor g0317(.dina(n617), .dinb(G503), .dout(n618));
  jor  g0318(.dina(G338), .dinb(n613), .dout(n619));
  jxor g0319(.dina(n619), .dinb(G514), .dout(n620));
  jor  g0320(.dina(G341), .dinb(G332), .dout(n621));
  jor  g0321(.dina(G348), .dinb(n613), .dout(n622));
  jand g0322(.dina(n622), .dinb(n621), .dout(n623));
  jxor g0323(.dina(n623), .dinb(G523), .dout(n624));
  jor  g0324(.dina(G351), .dinb(G332), .dout(n625));
  jor  g0325(.dina(G358), .dinb(n613), .dout(n626));
  jand g0326(.dina(n626), .dinb(n625), .dout(n627));
  jor  g0327(.dina(n627), .dinb(G534), .dout(n628));
  jnot g0328(.din(n625), .dout(n629));
  jand g0329(.dina(G612), .dinb(G332), .dout(n630));
  jor  g0330(.dina(n630), .dinb(n629), .dout(n631));
  jor  g0331(.dina(n631), .dinb(n377), .dout(n632));
  jor  g0332(.dina(G361), .dinb(G332), .dout(n633));
  jor  g0333(.dina(G366), .dinb(n613), .dout(n634));
  jand g0334(.dina(n634), .dinb(n633), .dout(n635));
  jnot g0335(.din(n635), .dout(n636));
  jand g0336(.dina(n636), .dinb(n632), .dout(n637));
  jand g0337(.dina(n637), .dinb(n628), .dout(n638));
  jand g0338(.dina(n638), .dinb(n624), .dout(n639));
  jand g0339(.dina(n639), .dinb(n620), .dout(n640));
  jand g0340(.dina(n640), .dinb(n618), .dout(n641));
  jand g0341(.dina(n613), .dinb(n425), .dout(n642));
  jand g0342(.dina(G332), .dinb(G593), .dout(n643));
  jor  g0343(.dina(n643), .dinb(n642), .dout(n644));
  jand g0344(.dina(n613), .dinb(n429), .dout(n645));
  jnot g0345(.din(n645), .dout(n646));
  jor  g0346(.dina(n613), .dinb(G307), .dout(n647));
  jand g0347(.dina(n647), .dinb(n646), .dout(n648));
  jnot g0348(.din(n648), .dout(n649));
  jand g0349(.dina(n649), .dinb(n644), .dout(n650));
  jor  g0350(.dina(G332), .dinb(G308), .dout(n651));
  jor  g0351(.dina(n613), .dinb(G315), .dout(n652));
  jand g0352(.dina(n652), .dinb(n651), .dout(n653));
  jxor g0353(.dina(n653), .dinb(G479), .dout(n654));
  jand g0354(.dina(n613), .dinb(n402), .dout(n655));
  jnot g0355(.din(n655), .dout(n656));
  jor  g0356(.dina(n613), .dinb(G323), .dout(n657));
  jand g0357(.dina(n657), .dinb(n656), .dout(n658));
  jxor g0358(.dina(n658), .dinb(G490), .dout(n659));
  jand g0359(.dina(n659), .dinb(n654), .dout(n660));
  jand g0360(.dina(n660), .dinb(n650), .dout(n661));
  jand g0361(.dina(n661), .dinb(n641), .dout(G615));
  jxor g0362(.dina(G316), .dinb(G308), .dout(n663));
  jxor g0363(.dina(G302), .dinb(n425), .dout(n664));
  jxor g0364(.dina(n664), .dinb(n663), .dout(n665));
  jxor g0365(.dina(G369), .dinb(G361), .dout(n666));
  jxor g0366(.dina(n666), .dinb(n435), .dout(n667));
  jxor g0367(.dina(G351), .dinb(G341), .dout(n668));
  jxor g0368(.dina(n668), .dinb(n667), .dout(n669));
  jxor g0369(.dina(n669), .dinb(n665), .dout(n670));
  jnot g0370(.din(n670), .dout(G1002));
  jxor g0371(.dina(G226), .dinb(G218), .dout(n672));
  jxor g0372(.dina(G273), .dinb(n483), .dout(n673));
  jxor g0373(.dina(n673), .dinb(n672), .dout(n674));
  jxor g0374(.dina(G289), .dinb(G281), .dout(n675));
  jxor g0375(.dina(G257), .dinb(G234), .dout(n676));
  jxor g0376(.dina(n676), .dinb(n675), .dout(n677));
  jxor g0377(.dina(G210), .dinb(G206), .dout(n678));
  jxor g0378(.dina(n678), .dinb(n677), .dout(n679));
  jxor g0379(.dina(n679), .dinb(n674), .dout(n680));
  jnot g0380(.din(n680), .dout(G1004));
  jand g0381(.dina(n586), .dinb(G435), .dout(n682));
  jnot g0382(.din(n586), .dout(n683));
  jand g0383(.dina(n683), .dinb(n462), .dout(n684));
  jnot g0384(.din(n684), .dout(n685));
  jand g0385(.dina(n578), .dinb(G389), .dout(n686));
  jor  g0386(.dina(n578), .dinb(G389), .dout(n687));
  jnot g0387(.din(n571), .dout(n688));
  jor  g0388(.dina(n688), .dinb(n569), .dout(n689));
  jand g0389(.dina(n689), .dinb(n485), .dout(n690));
  jnot g0390(.din(n690), .dout(n691));
  jand g0391(.dina(n560), .dinb(G374), .dout(n692));
  jor  g0392(.dina(n565), .dinb(G411), .dout(n693));
  jand g0393(.dina(n693), .dinb(n692), .dout(n694));
  jand g0394(.dina(n565), .dinb(G411), .dout(n695));
  jand g0395(.dina(n572), .dinb(G400), .dout(n696));
  jor  g0396(.dina(n696), .dinb(n695), .dout(n697));
  jor  g0397(.dina(n697), .dinb(n694), .dout(n698));
  jand g0398(.dina(n698), .dinb(n691), .dout(n699));
  jand g0399(.dina(n699), .dinb(n687), .dout(n700));
  jor  g0400(.dina(n700), .dinb(n686), .dout(n701));
  jand g0401(.dina(n701), .dinb(n685), .dout(n702));
  jor  g0402(.dina(n702), .dinb(n682), .dout(n703));
  jand g0403(.dina(n703), .dinb(n611), .dout(n704));
  jand g0404(.dina(n591), .dinb(G446), .dout(n705));
  jor  g0405(.dina(n591), .dinb(G446), .dout(n706));
  jand g0406(.dina(n607), .dinb(G457), .dout(n707));
  jor  g0407(.dina(n607), .dinb(G457), .dout(n708));
  jand g0408(.dina(n601), .dinb(G468), .dout(n709));
  jand g0409(.dina(n596), .dinb(G422), .dout(n710));
  jor  g0410(.dina(n601), .dinb(G468), .dout(n711));
  jand g0411(.dina(n711), .dinb(n710), .dout(n712));
  jor  g0412(.dina(n712), .dinb(n709), .dout(n713));
  jand g0413(.dina(n713), .dinb(n708), .dout(n714));
  jor  g0414(.dina(n714), .dinb(n707), .dout(n715));
  jand g0415(.dina(n715), .dinb(n706), .dout(n716));
  jor  g0416(.dina(n716), .dinb(n705), .dout(n717));
  jor  g0417(.dina(n717), .dinb(n704), .dout(G591));
  jand g0418(.dina(n617), .dinb(G503), .dout(n719));
  jor  g0419(.dina(n617), .dinb(G503), .dout(n720));
  jor  g0420(.dina(n619), .dinb(G514), .dout(n721));
  jand g0421(.dina(n619), .dinb(G514), .dout(n722));
  jnot g0422(.din(n621), .dout(n723));
  jand g0423(.dina(G599), .dinb(G332), .dout(n724));
  jor  g0424(.dina(n724), .dinb(n723), .dout(n725));
  jand g0425(.dina(n725), .dinb(n389), .dout(n726));
  jnot g0426(.din(n726), .dout(n727));
  jand g0427(.dina(n635), .dinb(n628), .dout(n728));
  jand g0428(.dina(n623), .dinb(G523), .dout(n729));
  jand g0429(.dina(n627), .dinb(G534), .dout(n730));
  jor  g0430(.dina(n730), .dinb(n729), .dout(n731));
  jor  g0431(.dina(n731), .dinb(n728), .dout(n732));
  jand g0432(.dina(n732), .dinb(n727), .dout(n733));
  jor  g0433(.dina(n733), .dinb(n722), .dout(n734));
  jand g0434(.dina(n734), .dinb(n721), .dout(n735));
  jand g0435(.dina(n735), .dinb(n720), .dout(n736));
  jor  g0436(.dina(n736), .dinb(n719), .dout(n737));
  jand g0437(.dina(n737), .dinb(n660), .dout(n738));
  jnot g0438(.din(n650), .dout(n739));
  jnot g0439(.din(n653), .dout(n740));
  jor  g0440(.dina(n740), .dinb(n414), .dout(n741));
  jand g0441(.dina(n658), .dinb(G490), .dout(n742));
  jand g0442(.dina(n742), .dinb(n654), .dout(n743));
  jnot g0443(.din(n743), .dout(n744));
  jand g0444(.dina(n744), .dinb(n741), .dout(n745));
  jnot g0445(.din(n745), .dout(n746));
  jor  g0446(.dina(n746), .dinb(n739), .dout(n747));
  jor  g0447(.dina(n747), .dinb(n738), .dout(G618));
  jnot g0448(.din(G4091), .dout(n749));
  jand g0449(.dina(G4092), .dinb(n749), .dout(n750));
  jand g0450(.dina(n750), .dinb(G131), .dout(n751));
  jnot g0451(.din(n751), .dout(n752));
  jnot g0452(.din(G54), .dout(n753));
  jxor g0453(.dina(n635), .dinb(n753), .dout(n754));
  jnot g0454(.din(n754), .dout(n755));
  jand g0455(.dina(n755), .dinb(G4091), .dout(n756));
  jand g0456(.dina(n372), .dinb(n749), .dout(n757));
  jor  g0457(.dina(n757), .dinb(G4092), .dout(n758));
  jor  g0458(.dina(n758), .dinb(n756), .dout(n759));
  jand g0459(.dina(n759), .dinb(n752), .dout(G822));
  jand g0460(.dina(n750), .dinb(G129), .dout(n761));
  jnot g0461(.din(n761), .dout(n762));
  jxor g0462(.dina(n627), .dinb(G534), .dout(n763));
  jnot g0463(.din(n763), .dout(n764));
  jand g0464(.dina(n764), .dinb(n635), .dout(n765));
  jor  g0465(.dina(n765), .dinb(n638), .dout(n766));
  jnot g0466(.din(n766), .dout(n767));
  jand g0467(.dina(n767), .dinb(n753), .dout(n768));
  jand g0468(.dina(n763), .dinb(G54), .dout(n769));
  jor  g0469(.dina(n769), .dinb(n768), .dout(n770));
  jand g0470(.dina(n770), .dinb(G4091), .dout(n771));
  jand g0471(.dina(n386), .dinb(n749), .dout(n772));
  jor  g0472(.dina(n772), .dinb(G4092), .dout(n773));
  jor  g0473(.dina(n773), .dinb(n771), .dout(n774));
  jand g0474(.dina(n774), .dinb(n762), .dout(G838));
  jand g0475(.dina(n750), .dinb(G117), .dout(n776));
  jnot g0476(.din(n776), .dout(n777));
  jxor g0477(.dina(n561), .dinb(G4), .dout(n778));
  jnot g0478(.din(n778), .dout(n779));
  jand g0479(.dina(n779), .dinb(G4091), .dout(n780));
  jand g0480(.dina(n540), .dinb(n749), .dout(n781));
  jor  g0481(.dina(n781), .dinb(G4092), .dout(n782));
  jor  g0482(.dina(n782), .dinb(n780), .dout(n783));
  jand g0483(.dina(n783), .dinb(n777), .dout(G861));
  jand g0484(.dina(n641), .dinb(G54), .dout(n785));
  jor  g0485(.dina(n785), .dinb(n737), .dout(n786));
  jand g0486(.dina(n786), .dinb(n660), .dout(n787));
  jor  g0487(.dina(n787), .dinb(n746), .dout(n788));
  jnot g0488(.din(n788), .dout(n789));
  jnot g0489(.din(n644), .dout(n790));
  jxor g0490(.dina(n648), .dinb(n790), .dout(n791));
  jnot g0491(.din(n791), .dout(n792));
  jand g0492(.dina(n792), .dinb(n789), .dout(n793));
  jand g0493(.dina(n788), .dinb(n790), .dout(n794));
  jor  g0494(.dina(n794), .dinb(n793), .dout(n795));
  jnot g0495(.din(n795), .dout(G623));
  jnot g0496(.din(G4088), .dout(n797));
  jnot g0497(.din(G861), .dout(n798));
  jor  g0498(.dina(n798), .dinb(n797), .dout(n799));
  jnot g0499(.din(G4087), .dout(n800));
  jnot g0500(.din(G822), .dout(n801));
  jor  g0501(.dina(n801), .dinb(G4088), .dout(n802));
  jand g0502(.dina(n802), .dinb(n800), .dout(n803));
  jand g0503(.dina(n803), .dinb(n799), .dout(n804));
  jor  g0504(.dina(n797), .dinb(G61), .dout(n805));
  jor  g0505(.dina(G4088), .dinb(G11), .dout(n806));
  jand g0506(.dina(n806), .dinb(G4087), .dout(n807));
  jand g0507(.dina(n807), .dinb(n805), .dout(n808));
  jor  g0508(.dina(n808), .dinb(n804), .dout(G722));
  jand g0509(.dina(n750), .dinb(G52), .dout(n810));
  jnot g0510(.din(n810), .dout(n811));
  jnot g0511(.din(n721), .dout(n812));
  jnot g0512(.din(n722), .dout(n813));
  jand g0513(.dina(n631), .dinb(n377), .dout(n814));
  jor  g0514(.dina(n636), .dinb(n814), .dout(n815));
  jor  g0515(.dina(n725), .dinb(n389), .dout(n816));
  jand g0516(.dina(n632), .dinb(n816), .dout(n817));
  jand g0517(.dina(n817), .dinb(n815), .dout(n818));
  jor  g0518(.dina(n818), .dinb(n726), .dout(n819));
  jand g0519(.dina(n819), .dinb(n813), .dout(n820));
  jor  g0520(.dina(n820), .dinb(n812), .dout(n821));
  jnot g0521(.din(n620), .dout(n822));
  jnot g0522(.din(n639), .dout(n823));
  jor  g0523(.dina(n823), .dinb(n753), .dout(n824));
  jor  g0524(.dina(n824), .dinb(n822), .dout(n825));
  jand g0525(.dina(n825), .dinb(n821), .dout(n826));
  jxor g0526(.dina(n826), .dinb(n618), .dout(n827));
  jand g0527(.dina(n827), .dinb(G4091), .dout(n828));
  jand g0528(.dina(n445), .dinb(n749), .dout(n829));
  jor  g0529(.dina(n829), .dinb(G4092), .dout(n830));
  jor  g0530(.dina(n830), .dinb(n828), .dout(n831));
  jand g0531(.dina(n831), .dinb(n811), .dout(G832));
  jand g0532(.dina(n750), .dinb(G130), .dout(n833));
  jnot g0533(.din(n833), .dout(n834));
  jand g0534(.dina(n824), .dinb(n819), .dout(n835));
  jxor g0535(.dina(n835), .dinb(n620), .dout(n836));
  jand g0536(.dina(n836), .dinb(G4091), .dout(n837));
  jand g0537(.dina(n365), .dinb(n749), .dout(n838));
  jor  g0538(.dina(n838), .dinb(G4092), .dout(n839));
  jor  g0539(.dina(n839), .dinb(n837), .dout(n840));
  jand g0540(.dina(n840), .dinb(n834), .dout(G834));
  jand g0541(.dina(n750), .dinb(G119), .dout(n842));
  jnot g0542(.din(n842), .dout(n843));
  jand g0543(.dina(n397), .dinb(n749), .dout(n844));
  jand g0544(.dina(n637), .dinb(n753), .dout(n845));
  jor  g0545(.dina(n845), .dinb(n814), .dout(n846));
  jxor g0546(.dina(n846), .dinb(n624), .dout(n847));
  jand g0547(.dina(n847), .dinb(G4091), .dout(n848));
  jor  g0548(.dina(n848), .dinb(G4092), .dout(n849));
  jor  g0549(.dina(n849), .dinb(n844), .dout(n850));
  jand g0550(.dina(n850), .dinb(n843), .dout(G836));
  jnot g0551(.din(G4089), .dout(n852));
  jor  g0552(.dina(n798), .dinb(n852), .dout(n853));
  jnot g0553(.din(G4090), .dout(n854));
  jor  g0554(.dina(n801), .dinb(G4089), .dout(n855));
  jand g0555(.dina(n855), .dinb(n854), .dout(n856));
  jand g0556(.dina(n856), .dinb(n853), .dout(n857));
  jor  g0557(.dina(n852), .dinb(G61), .dout(n858));
  jor  g0558(.dina(G4089), .dinb(G11), .dout(n859));
  jand g0559(.dina(n859), .dinb(G4090), .dout(n860));
  jand g0560(.dina(n860), .dinb(n858), .dout(n861));
  jor  g0561(.dina(n861), .dinb(n857), .dout(G859));
  jand g0562(.dina(n750), .dinb(G122), .dout(n863));
  jnot g0563(.din(n863), .dout(n864));
  jnot g0564(.din(n587), .dout(n865));
  jnot g0565(.din(n579), .dout(n866));
  jand g0566(.dina(n567), .dinb(G4), .dout(n867));
  jand g0567(.dina(n867), .dinb(n573), .dout(n868));
  jand g0568(.dina(n868), .dinb(n866), .dout(n869));
  jor  g0569(.dina(n869), .dinb(n701), .dout(n870));
  jxor g0570(.dina(n870), .dinb(n865), .dout(n871));
  jand g0571(.dina(n871), .dinb(G4091), .dout(n872));
  jand g0572(.dina(n470), .dinb(n749), .dout(n873));
  jor  g0573(.dina(n873), .dinb(G4092), .dout(n874));
  jor  g0574(.dina(n874), .dinb(n872), .dout(n875));
  jand g0575(.dina(n875), .dinb(n864), .dout(G871));
  jand g0576(.dina(n750), .dinb(G128), .dout(n877));
  jnot g0577(.din(n877), .dout(n878));
  jor  g0578(.dina(n868), .dinb(n699), .dout(n879));
  jxor g0579(.dina(n879), .dinb(n579), .dout(n880));
  jand g0580(.dina(n880), .dinb(G4091), .dout(n881));
  jand g0581(.dina(n528), .dinb(n749), .dout(n882));
  jor  g0582(.dina(n882), .dinb(G4092), .dout(n883));
  jor  g0583(.dina(n883), .dinb(n881), .dout(n884));
  jand g0584(.dina(n884), .dinb(n878), .dout(G873));
  jand g0585(.dina(n750), .dinb(G127), .dout(n886));
  jnot g0586(.din(n886), .dout(n887));
  jor  g0587(.dina(n694), .dinb(n695), .dout(n888));
  jor  g0588(.dina(n888), .dinb(n867), .dout(n889));
  jxor g0589(.dina(n889), .dinb(n574), .dout(n890));
  jand g0590(.dina(n890), .dinb(G4091), .dout(n891));
  jand g0591(.dina(n493), .dinb(n749), .dout(n892));
  jor  g0592(.dina(n892), .dinb(G4092), .dout(n893));
  jor  g0593(.dina(n893), .dinb(n891), .dout(n894));
  jand g0594(.dina(n894), .dinb(n887), .dout(G875));
  jand g0595(.dina(n750), .dinb(G126), .dout(n896));
  jnot g0596(.din(n896), .dout(n897));
  jnot g0597(.din(n566), .dout(n898));
  jand g0598(.dina(n561), .dinb(G4), .dout(n899));
  jor  g0599(.dina(n899), .dinb(n692), .dout(n900));
  jxor g0600(.dina(n900), .dinb(n898), .dout(n901));
  jand g0601(.dina(n901), .dinb(G4091), .dout(n902));
  jand g0602(.dina(n481), .dinb(n749), .dout(n903));
  jor  g0603(.dina(n903), .dinb(G4092), .dout(n904));
  jor  g0604(.dina(n904), .dinb(n902), .dout(n905));
  jand g0605(.dina(n905), .dinb(n897), .dout(G877));
  jnot g0606(.din(G331), .dout(n907));
  jnot g0607(.din(n619), .dout(n908));
  jand g0608(.dina(n908), .dinb(n907), .dout(n909));
  jand g0609(.dina(n619), .dinb(n617), .dout(n910));
  jor  g0610(.dina(n910), .dinb(n909), .dout(n911));
  jxor g0611(.dina(n911), .dinb(n792), .dout(n912));
  jor  g0612(.dina(G369), .dinb(G332), .dout(n913));
  jor  g0613(.dina(G372), .dinb(n613), .dout(n914));
  jand g0614(.dina(n914), .dinb(n913), .dout(n915));
  jxor g0615(.dina(n915), .dinb(n636), .dout(n916));
  jxor g0616(.dina(n627), .dinb(n725), .dout(n917));
  jxor g0617(.dina(n658), .dinb(n653), .dout(n918));
  jxor g0618(.dina(n918), .dinb(n917), .dout(n919));
  jxor g0619(.dina(n919), .dinb(n916), .dout(n920));
  jxor g0620(.dina(n920), .dinb(n912), .dout(G998));
  jnot g0621(.din(n564), .dout(n922));
  jor  g0622(.dina(n922), .dinb(n562), .dout(n923));
  jxor g0623(.dina(n578), .dinb(n923), .dout(n924));
  jxor g0624(.dina(n572), .dinb(n560), .dout(n925));
  jxor g0625(.dina(n925), .dinb(n924), .dout(n926));
  jor  g0626(.dina(G335), .dinb(G289), .dout(n927));
  jor  g0627(.dina(n556), .dinb(G292), .dout(n928));
  jand g0628(.dina(n928), .dinb(n927), .dout(n929));
  jxor g0629(.dina(n929), .dinb(n591), .dout(n930));
  jxor g0630(.dina(n596), .dinb(n586), .dout(n931));
  jxor g0631(.dina(n607), .dinb(n601), .dout(n932));
  jxor g0632(.dina(n932), .dinb(n931), .dout(n933));
  jxor g0633(.dina(n933), .dinb(n930), .dout(n934));
  jxor g0634(.dina(n934), .dinb(n926), .dout(n935));
  jnot g0635(.din(n935), .dout(G1000));
  jnot g0636(.din(n592), .dout(n937));
  jnot g0637(.din(n715), .dout(n938));
  jor  g0638(.dina(n870), .dinb(n682), .dout(n939));
  jand g0639(.dina(n939), .dinb(n685), .dout(n940));
  jnot g0640(.din(n940), .dout(n941));
  jor  g0641(.dina(n941), .dinb(n609), .dout(n942));
  jand g0642(.dina(n942), .dinb(n938), .dout(n943));
  jxor g0643(.dina(n943), .dinb(n937), .dout(n944));
  jnot g0644(.din(n944), .dout(n945));
  jnot g0645(.din(n603), .dout(n946));
  jand g0646(.dina(n940), .dinb(n946), .dout(n947));
  jor  g0647(.dina(n947), .dinb(n713), .dout(n948));
  jxor g0648(.dina(n948), .dinb(n608), .dout(n949));
  jand g0649(.dina(n949), .dinb(n945), .dout(n950));
  jnot g0650(.din(n602), .dout(n951));
  jnot g0651(.din(n596), .dout(n952));
  jand g0652(.dina(n952), .dinb(n496), .dout(n953));
  jnot g0653(.din(n953), .dout(n954));
  jor  g0654(.dina(n940), .dinb(n710), .dout(n955));
  jand g0655(.dina(n955), .dinb(n954), .dout(n956));
  jxor g0656(.dina(n956), .dinb(n951), .dout(n957));
  jnot g0657(.din(n957), .dout(n958));
  jand g0658(.dina(n890), .dinb(n779), .dout(n959));
  jand g0659(.dina(n959), .dinb(n901), .dout(n960));
  jand g0660(.dina(n960), .dinb(n871), .dout(n961));
  jnot g0661(.din(n597), .dout(n962));
  jxor g0662(.dina(n940), .dinb(n962), .dout(n963));
  jnot g0663(.din(n963), .dout(n964));
  jand g0664(.dina(n964), .dinb(n880), .dout(n965));
  jand g0665(.dina(n965), .dinb(n961), .dout(n966));
  jand g0666(.dina(n966), .dinb(n958), .dout(n967));
  jand g0667(.dina(n967), .dinb(n950), .dout(G575));
  jxor g0668(.dina(n788), .dinb(n649), .dout(n969));
  jnot g0669(.din(n969), .dout(n970));
  jand g0670(.dina(n970), .dinb(n755), .dout(n971));
  jand g0671(.dina(n836), .dinb(G623), .dout(n972));
  jand g0672(.dina(n972), .dinb(n971), .dout(n973));
  jand g0673(.dina(n827), .dinb(n763), .dout(n974));
  jand g0674(.dina(n974), .dinb(n847), .dout(n975));
  jnot g0675(.din(n658), .dout(n976));
  jand g0676(.dina(n976), .dinb(n401), .dout(n977));
  jand g0677(.dina(n977), .dinb(n654), .dout(n978));
  jor  g0678(.dina(n977), .dinb(n654), .dout(n979));
  jnot g0679(.din(n979), .dout(n980));
  jor  g0680(.dina(n786), .dinb(n742), .dout(n981));
  jand g0681(.dina(n981), .dinb(n980), .dout(n982));
  jnot g0682(.din(n981), .dout(n983));
  jand g0683(.dina(n983), .dinb(n654), .dout(n984));
  jor  g0684(.dina(n984), .dinb(n982), .dout(n985));
  jor  g0685(.dina(n985), .dinb(n978), .dout(n986));
  jnot g0686(.din(n986), .dout(n987));
  jnot g0687(.din(n659), .dout(n988));
  jxor g0688(.dina(n786), .dinb(n988), .dout(n989));
  jand g0689(.dina(n989), .dinb(n987), .dout(n990));
  jand g0690(.dina(n990), .dinb(n975), .dout(n991));
  jand g0691(.dina(n991), .dinb(n973), .dout(G585));
  jnot g0692(.din(G1689), .dout(n993));
  jand g0693(.dina(G1690), .dinb(n993), .dout(n994));
  jand g0694(.dina(n994), .dinb(G182), .dout(n995));
  jand g0695(.dina(G1690), .dinb(G1689), .dout(n996));
  jand g0696(.dina(n996), .dinb(G185), .dout(n997));
  jor  g0697(.dina(n798), .dinb(n993), .dout(n998));
  jnot g0698(.din(G1690), .dout(n999));
  jor  g0699(.dina(n801), .dinb(G1689), .dout(n1000));
  jand g0700(.dina(n1000), .dinb(n999), .dout(n1001));
  jand g0701(.dina(n1001), .dinb(n998), .dout(n1002));
  jor  g0702(.dina(n1002), .dinb(n997), .dout(n1003));
  jor  g0703(.dina(n1003), .dinb(n995), .dout(n1004));
  jand g0704(.dina(n1004), .dinb(G137), .dout(G661));
  jor  g0705(.dina(n801), .dinb(G1691), .dout(n1006));
  jnot g0706(.din(G1694), .dout(n1007));
  jnot g0707(.din(G1691), .dout(n1008));
  jor  g0708(.dina(n798), .dinb(n1008), .dout(n1009));
  jand g0709(.dina(n1009), .dinb(n1007), .dout(n1010));
  jand g0710(.dina(n1010), .dinb(n1006), .dout(n1011));
  jand g0711(.dina(G1694), .dinb(G1691), .dout(n1012));
  jand g0712(.dina(n1012), .dinb(G185), .dout(n1013));
  jand g0713(.dina(G1694), .dinb(n1008), .dout(n1014));
  jand g0714(.dina(n1014), .dinb(G182), .dout(n1015));
  jor  g0715(.dina(n1015), .dinb(n1013), .dout(n1016));
  jor  g0716(.dina(n1016), .dinb(n1011), .dout(n1017));
  jand g0717(.dina(n1017), .dinb(G137), .dout(G693));
  jnot g0718(.din(G871), .dout(n1019));
  jor  g0719(.dina(n1019), .dinb(n797), .dout(n1020));
  jnot g0720(.din(G832), .dout(n1021));
  jor  g0721(.dina(n1021), .dinb(G4088), .dout(n1022));
  jand g0722(.dina(n1022), .dinb(n800), .dout(n1023));
  jand g0723(.dina(n1023), .dinb(n1020), .dout(n1024));
  jor  g0724(.dina(n797), .dinb(G37), .dout(n1025));
  jor  g0725(.dina(G4088), .dinb(G43), .dout(n1026));
  jand g0726(.dina(n1026), .dinb(G4087), .dout(n1027));
  jand g0727(.dina(n1027), .dinb(n1025), .dout(n1028));
  jor  g0728(.dina(n1028), .dinb(n1024), .dout(G747));
  jnot g0729(.din(G873), .dout(n1030));
  jor  g0730(.dina(n1030), .dinb(n797), .dout(n1031));
  jnot g0731(.din(G834), .dout(n1032));
  jor  g0732(.dina(n1032), .dinb(G4088), .dout(n1033));
  jand g0733(.dina(n1033), .dinb(n800), .dout(n1034));
  jand g0734(.dina(n1034), .dinb(n1031), .dout(n1035));
  jor  g0735(.dina(n797), .dinb(G20), .dout(n1036));
  jor  g0736(.dina(G4088), .dinb(G76), .dout(n1037));
  jand g0737(.dina(n1037), .dinb(G4087), .dout(n1038));
  jand g0738(.dina(n1038), .dinb(n1036), .dout(n1039));
  jor  g0739(.dina(n1039), .dinb(n1035), .dout(G752));
  jnot g0740(.din(G836), .dout(n1041));
  jor  g0741(.dina(n1041), .dinb(G4088), .dout(n1042));
  jnot g0742(.din(G875), .dout(n1043));
  jor  g0743(.dina(n1043), .dinb(n797), .dout(n1044));
  jand g0744(.dina(n1044), .dinb(n800), .dout(n1045));
  jand g0745(.dina(n1045), .dinb(n1042), .dout(n1046));
  jor  g0746(.dina(n797), .dinb(G17), .dout(n1047));
  jor  g0747(.dina(G4088), .dinb(G73), .dout(n1048));
  jand g0748(.dina(n1048), .dinb(G4087), .dout(n1049));
  jand g0749(.dina(n1049), .dinb(n1047), .dout(n1050));
  jor  g0750(.dina(n1050), .dinb(n1046), .dout(G757));
  jnot g0751(.din(G877), .dout(n1052));
  jor  g0752(.dina(n1052), .dinb(n797), .dout(n1053));
  jnot g0753(.din(G838), .dout(n1054));
  jor  g0754(.dina(n1054), .dinb(G4088), .dout(n1055));
  jand g0755(.dina(n1055), .dinb(n800), .dout(n1056));
  jand g0756(.dina(n1056), .dinb(n1053), .dout(n1057));
  jor  g0757(.dina(n797), .dinb(G70), .dout(n1058));
  jor  g0758(.dina(G4088), .dinb(G67), .dout(n1059));
  jand g0759(.dina(n1059), .dinb(G4087), .dout(n1060));
  jand g0760(.dina(n1060), .dinb(n1058), .dout(n1061));
  jor  g0761(.dina(n1061), .dinb(n1057), .dout(G762));
  jor  g0762(.dina(G4089), .dinb(G43), .dout(n1063));
  jor  g0763(.dina(n852), .dinb(G37), .dout(n1064));
  jand g0764(.dina(n1064), .dinb(G4090), .dout(n1065));
  jand g0765(.dina(n1065), .dinb(n1063), .dout(n1066));
  jor  g0766(.dina(n1021), .dinb(G4089), .dout(n1067));
  jor  g0767(.dina(n1019), .dinb(n852), .dout(n1068));
  jand g0768(.dina(n1068), .dinb(n1067), .dout(n1069));
  jand g0769(.dina(n1069), .dinb(n854), .dout(n1070));
  jor  g0770(.dina(n1070), .dinb(n1066), .dout(G787));
  jor  g0771(.dina(G4089), .dinb(G76), .dout(n1072));
  jor  g0772(.dina(n852), .dinb(G20), .dout(n1073));
  jand g0773(.dina(n1073), .dinb(G4090), .dout(n1074));
  jand g0774(.dina(n1074), .dinb(n1072), .dout(n1075));
  jor  g0775(.dina(n1032), .dinb(G4089), .dout(n1076));
  jor  g0776(.dina(n1030), .dinb(n852), .dout(n1077));
  jand g0777(.dina(n1077), .dinb(n1076), .dout(n1078));
  jand g0778(.dina(n1078), .dinb(n854), .dout(n1079));
  jor  g0779(.dina(n1079), .dinb(n1075), .dout(G792));
  jor  g0780(.dina(G4089), .dinb(G73), .dout(n1081));
  jor  g0781(.dina(n852), .dinb(G17), .dout(n1082));
  jand g0782(.dina(n1082), .dinb(G4090), .dout(n1083));
  jand g0783(.dina(n1083), .dinb(n1081), .dout(n1084));
  jor  g0784(.dina(n1043), .dinb(n852), .dout(n1085));
  jor  g0785(.dina(n1041), .dinb(G4089), .dout(n1086));
  jand g0786(.dina(n1086), .dinb(n1085), .dout(n1087));
  jand g0787(.dina(n1087), .dinb(n854), .dout(n1088));
  jor  g0788(.dina(n1088), .dinb(n1084), .dout(G797));
  jor  g0789(.dina(n1052), .dinb(n852), .dout(n1090));
  jor  g0790(.dina(n1054), .dinb(G4089), .dout(n1091));
  jand g0791(.dina(n1091), .dinb(n854), .dout(n1092));
  jand g0792(.dina(n1092), .dinb(n1090), .dout(n1093));
  jor  g0793(.dina(n852), .dinb(G70), .dout(n1094));
  jor  g0794(.dina(G4089), .dinb(G67), .dout(n1095));
  jand g0795(.dina(n1095), .dinb(G4090), .dout(n1096));
  jand g0796(.dina(n1096), .dinb(n1094), .dout(n1097));
  jor  g0797(.dina(n1097), .dinb(n1093), .dout(G802));
  jor  g0798(.dina(n1021), .dinb(G1689), .dout(n1099));
  jor  g0799(.dina(n1019), .dinb(n993), .dout(n1100));
  jand g0800(.dina(n1100), .dinb(n999), .dout(n1101));
  jand g0801(.dina(n1101), .dinb(n1099), .dout(n1102));
  jand g0802(.dina(n994), .dinb(G200), .dout(n1103));
  jand g0803(.dina(n996), .dinb(G170), .dout(n1104));
  jor  g0804(.dina(n1104), .dinb(n1103), .dout(n1105));
  jor  g0805(.dina(n1105), .dinb(n1102), .dout(n1106));
  jand g0806(.dina(n1106), .dinb(G137), .dout(G642));
  jor  g0807(.dina(n1054), .dinb(G1689), .dout(n1108));
  jor  g0808(.dina(n1052), .dinb(n993), .dout(n1109));
  jand g0809(.dina(n1109), .dinb(n999), .dout(n1110));
  jand g0810(.dina(n1110), .dinb(n1108), .dout(n1111));
  jand g0811(.dina(n994), .dinb(G188), .dout(n1112));
  jand g0812(.dina(n996), .dinb(G158), .dout(n1113));
  jor  g0813(.dina(n1113), .dinb(n1112), .dout(n1114));
  jor  g0814(.dina(n1114), .dinb(n1111), .dout(n1115));
  jand g0815(.dina(n1115), .dinb(G137), .dout(G664));
  jor  g0816(.dina(n1041), .dinb(G1689), .dout(n1117));
  jor  g0817(.dina(n1043), .dinb(n993), .dout(n1118));
  jand g0818(.dina(n1118), .dinb(n999), .dout(n1119));
  jand g0819(.dina(n1119), .dinb(n1117), .dout(n1120));
  jand g0820(.dina(n994), .dinb(G155), .dout(n1121));
  jand g0821(.dina(n996), .dinb(G152), .dout(n1122));
  jor  g0822(.dina(n1122), .dinb(n1121), .dout(n1123));
  jor  g0823(.dina(n1123), .dinb(n1120), .dout(n1124));
  jand g0824(.dina(n1124), .dinb(G137), .dout(G667));
  jor  g0825(.dina(n1032), .dinb(G1689), .dout(n1126));
  jor  g0826(.dina(n1030), .dinb(n993), .dout(n1127));
  jand g0827(.dina(n1127), .dinb(n999), .dout(n1128));
  jand g0828(.dina(n1128), .dinb(n1126), .dout(n1129));
  jand g0829(.dina(n994), .dinb(G149), .dout(n1130));
  jand g0830(.dina(n996), .dinb(G146), .dout(n1131));
  jor  g0831(.dina(n1131), .dinb(n1130), .dout(n1132));
  jor  g0832(.dina(n1132), .dinb(n1129), .dout(n1133));
  jand g0833(.dina(n1133), .dinb(G137), .dout(G670));
  jand g0834(.dina(n1014), .dinb(G200), .dout(n1135));
  jand g0835(.dina(n1012), .dinb(G170), .dout(n1136));
  jor  g0836(.dina(n1019), .dinb(n1008), .dout(n1137));
  jor  g0837(.dina(n1021), .dinb(G1691), .dout(n1138));
  jand g0838(.dina(n1138), .dinb(n1137), .dout(n1139));
  jand g0839(.dina(n1139), .dinb(n1007), .dout(n1140));
  jor  g0840(.dina(n1140), .dinb(n1136), .dout(n1141));
  jor  g0841(.dina(n1141), .dinb(n1135), .dout(n1142));
  jand g0842(.dina(n1142), .dinb(G137), .dout(G676));
  jor  g0843(.dina(n1054), .dinb(G1691), .dout(n1144));
  jor  g0844(.dina(n1052), .dinb(n1008), .dout(n1145));
  jand g0845(.dina(n1145), .dinb(n1007), .dout(n1146));
  jand g0846(.dina(n1146), .dinb(n1144), .dout(n1147));
  jand g0847(.dina(n1014), .dinb(G188), .dout(n1148));
  jand g0848(.dina(n1012), .dinb(G158), .dout(n1149));
  jor  g0849(.dina(n1149), .dinb(n1148), .dout(n1150));
  jor  g0850(.dina(n1150), .dinb(n1147), .dout(n1151));
  jand g0851(.dina(n1151), .dinb(G137), .dout(G696));
  jor  g0852(.dina(n1041), .dinb(G1691), .dout(n1153));
  jor  g0853(.dina(n1043), .dinb(n1008), .dout(n1154));
  jand g0854(.dina(n1154), .dinb(n1007), .dout(n1155));
  jand g0855(.dina(n1155), .dinb(n1153), .dout(n1156));
  jand g0856(.dina(n1014), .dinb(G155), .dout(n1157));
  jand g0857(.dina(n1012), .dinb(G152), .dout(n1158));
  jor  g0858(.dina(n1158), .dinb(n1157), .dout(n1159));
  jor  g0859(.dina(n1159), .dinb(n1156), .dout(n1160));
  jand g0860(.dina(n1160), .dinb(G137), .dout(G699));
  jor  g0861(.dina(n1032), .dinb(G1691), .dout(n1162));
  jor  g0862(.dina(n1030), .dinb(n1008), .dout(n1163));
  jand g0863(.dina(n1163), .dinb(n1007), .dout(n1164));
  jand g0864(.dina(n1164), .dinb(n1162), .dout(n1165));
  jand g0865(.dina(n1014), .dinb(G149), .dout(n1166));
  jand g0866(.dina(n1012), .dinb(G146), .dout(n1167));
  jor  g0867(.dina(n1167), .dinb(n1166), .dout(n1168));
  jor  g0868(.dina(n1168), .dinb(n1165), .dout(n1169));
  jand g0869(.dina(n1169), .dinb(G137), .dout(G702));
  jnot g0870(.din(G135), .dout(n1171));
  jnot g0871(.din(G4115), .dout(n1172));
  jor  g0872(.dina(n1172), .dinb(n1171), .dout(n1173));
  jnot g0873(.din(n428), .dout(n1174));
  jor  g0874(.dina(n1174), .dinb(G3724), .dout(n1175));
  jnot g0875(.din(G3717), .dout(n1176));
  jnot g0876(.din(G3724), .dout(n1177));
  jxor g0877(.dina(n790), .dinb(G132), .dout(n1178));
  jnot g0878(.din(n1178), .dout(n1179));
  jor  g0879(.dina(n1179), .dinb(n1177), .dout(n1180));
  jand g0880(.dina(n1180), .dinb(n1176), .dout(n1181));
  jand g0881(.dina(n1181), .dinb(n1175), .dout(n1182));
  jor  g0882(.dina(n795), .dinb(n1177), .dout(n1183));
  jor  g0883(.dina(G3724), .dinb(G123), .dout(n1184));
  jand g0884(.dina(n1184), .dinb(G3717), .dout(n1185));
  jand g0885(.dina(n1185), .dinb(n1183), .dout(n1186));
  jor  g0886(.dina(n1186), .dinb(n1182), .dout(n1187));
  jand g0887(.dina(n1187), .dinb(n1173), .dout(G818));
  jxor g0888(.dina(n1179), .dinb(n795), .dout(G813));
  jand g0889(.dina(n750), .dinb(G123), .dout(n1190));
  jor  g0890(.dina(n795), .dinb(n749), .dout(n1191));
  jand g0891(.dina(n428), .dinb(n749), .dout(n1192));
  jor  g0892(.dina(n1192), .dinb(G4092), .dout(n1193));
  jnot g0893(.din(n1193), .dout(n1194));
  jand g0894(.dina(n1194), .dinb(n1191), .dout(n1195));
  jor  g0895(.dina(n1195), .dinb(n1190), .dout(n1196));
  jnot g0896(.din(n1196), .dout(G824));
  jand g0897(.dina(n750), .dinb(G121), .dout(n1198));
  jand g0898(.dina(n433), .dinb(n749), .dout(n1199));
  jnot g0899(.din(n1199), .dout(n1200));
  jnot g0900(.din(G4092), .dout(n1201));
  jor  g0901(.dina(n969), .dinb(n749), .dout(n1202));
  jand g0902(.dina(n1202), .dinb(n1201), .dout(n1203));
  jand g0903(.dina(n1203), .dinb(n1200), .dout(n1204));
  jor  g0904(.dina(n1204), .dinb(n1198), .dout(n1205));
  jnot g0905(.din(n1205), .dout(G826));
  jand g0906(.dina(n750), .dinb(G116), .dout(n1207));
  jor  g0907(.dina(n986), .dinb(n749), .dout(n1208));
  jand g0908(.dina(n423), .dinb(n749), .dout(n1209));
  jor  g0909(.dina(n1209), .dinb(G4092), .dout(n1210));
  jnot g0910(.din(n1210), .dout(n1211));
  jand g0911(.dina(n1211), .dinb(n1208), .dout(n1212));
  jor  g0912(.dina(n1212), .dinb(n1207), .dout(n1213));
  jnot g0913(.din(n1213), .dout(G828));
  jand g0914(.dina(n750), .dinb(G112), .dout(n1215));
  jnot g0915(.din(n1215), .dout(n1216));
  jand g0916(.dina(n989), .dinb(G4091), .dout(n1217));
  jand g0917(.dina(n412), .dinb(n749), .dout(n1218));
  jor  g0918(.dina(n1218), .dinb(G4092), .dout(n1219));
  jor  g0919(.dina(n1219), .dinb(n1217), .dout(n1220));
  jand g0920(.dina(n1220), .dinb(n1216), .dout(G830));
  jand g0921(.dina(n680), .dinb(G245), .dout(n1222));
  jand g0922(.dina(n1222), .dinb(n935), .dout(n1223));
  jnot g0923(.din(G998), .dout(n1224));
  jand g0924(.dina(n318), .dinb(G601), .dout(n1225));
  jand g0925(.dina(n1225), .dinb(G559), .dout(n1226));
  jand g0926(.dina(n1226), .dinb(n670), .dout(n1227));
  jand g0927(.dina(n1227), .dinb(n1224), .dout(n1228));
  jand g0928(.dina(n1228), .dinb(n1223), .dout(G854));
  jand g0929(.dina(n750), .dinb(G115), .dout(n1230));
  jand g0930(.dina(n551), .dinb(n749), .dout(n1231));
  jnot g0931(.din(n1231), .dout(n1232));
  jor  g0932(.dina(n944), .dinb(n749), .dout(n1233));
  jand g0933(.dina(n1233), .dinb(n1201), .dout(n1234));
  jand g0934(.dina(n1234), .dinb(n1232), .dout(n1235));
  jor  g0935(.dina(n1235), .dinb(n1230), .dout(n1236));
  jnot g0936(.din(n1236), .dout(G863));
  jand g0937(.dina(n750), .dinb(G114), .dout(n1238));
  jnot g0938(.din(n1238), .dout(n1239));
  jand g0939(.dina(n949), .dinb(G4091), .dout(n1240));
  jand g0940(.dina(n459), .dinb(n749), .dout(n1241));
  jor  g0941(.dina(n1241), .dinb(G4092), .dout(n1242));
  jor  g0942(.dina(n1242), .dinb(n1240), .dout(n1243));
  jand g0943(.dina(n1243), .dinb(n1239), .dout(G865));
  jand g0944(.dina(n750), .dinb(G53), .dout(n1245));
  jand g0945(.dina(n517), .dinb(n749), .dout(n1246));
  jnot g0946(.din(n1246), .dout(n1247));
  jor  g0947(.dina(n957), .dinb(n749), .dout(n1248));
  jand g0948(.dina(n1248), .dinb(n1201), .dout(n1249));
  jand g0949(.dina(n1249), .dinb(n1247), .dout(n1250));
  jor  g0950(.dina(n1250), .dinb(n1245), .dout(n1251));
  jnot g0951(.din(n1251), .dout(G867));
  jand g0952(.dina(n750), .dinb(G113), .dout(n1253));
  jnot g0953(.din(n1253), .dout(n1254));
  jand g0954(.dina(n964), .dinb(G4091), .dout(n1255));
  jand g0955(.dina(n504), .dinb(n749), .dout(n1256));
  jor  g0956(.dina(n1256), .dinb(G4092), .dout(n1257));
  jor  g0957(.dina(n1257), .dinb(n1255), .dout(n1258));
  jand g0958(.dina(n1258), .dinb(n1254), .dout(G869));
  jor  g0959(.dina(G4089), .dinb(G109), .dout(n1260));
  jor  g0960(.dina(n852), .dinb(G106), .dout(n1261));
  jand g0961(.dina(n1261), .dinb(G4090), .dout(n1262));
  jand g0962(.dina(n1262), .dinb(n1260), .dout(n1263));
  jor  g0963(.dina(n1236), .dinb(n852), .dout(n1264));
  jor  g0964(.dina(n1196), .dinb(G4089), .dout(n1265));
  jand g0965(.dina(n1265), .dinb(n854), .dout(n1266));
  jand g0966(.dina(n1266), .dinb(n1264), .dout(n1267));
  jor  g0967(.dina(n1267), .dinb(n1263), .dout(G712));
  jor  g0968(.dina(n1196), .dinb(G4088), .dout(n1269));
  jor  g0969(.dina(n1236), .dinb(n797), .dout(n1270));
  jand g0970(.dina(n1270), .dinb(n800), .dout(n1271));
  jand g0971(.dina(n1271), .dinb(n1269), .dout(n1272));
  jor  g0972(.dina(n797), .dinb(G106), .dout(n1273));
  jor  g0973(.dina(G4088), .dinb(G109), .dout(n1274));
  jand g0974(.dina(n1274), .dinb(G4087), .dout(n1275));
  jand g0975(.dina(n1275), .dinb(n1273), .dout(n1276));
  jor  g0976(.dina(n1276), .dinb(n1272), .dout(G727));
  jor  g0977(.dina(n1205), .dinb(G4088), .dout(n1278));
  jnot g0978(.din(G865), .dout(n1279));
  jor  g0979(.dina(n1279), .dinb(n797), .dout(n1280));
  jand g0980(.dina(n1280), .dinb(n800), .dout(n1281));
  jand g0981(.dina(n1281), .dinb(n1278), .dout(n1282));
  jor  g0982(.dina(n797), .dinb(G49), .dout(n1283));
  jor  g0983(.dina(G4088), .dinb(G46), .dout(n1284));
  jand g0984(.dina(n1284), .dinb(G4087), .dout(n1285));
  jand g0985(.dina(n1285), .dinb(n1283), .dout(n1286));
  jor  g0986(.dina(n1286), .dinb(n1282), .dout(G732));
  jor  g0987(.dina(n1213), .dinb(G4088), .dout(n1288));
  jor  g0988(.dina(n1251), .dinb(n797), .dout(n1289));
  jand g0989(.dina(n1289), .dinb(n800), .dout(n1290));
  jand g0990(.dina(n1290), .dinb(n1288), .dout(n1291));
  jor  g0991(.dina(n797), .dinb(G103), .dout(n1292));
  jor  g0992(.dina(G4088), .dinb(G100), .dout(n1293));
  jand g0993(.dina(n1293), .dinb(G4087), .dout(n1294));
  jand g0994(.dina(n1294), .dinb(n1292), .dout(n1295));
  jor  g0995(.dina(n1295), .dinb(n1291), .dout(G737));
  jnot g0996(.din(G830), .dout(n1297));
  jor  g0997(.dina(n1297), .dinb(G4088), .dout(n1298));
  jnot g0998(.din(G869), .dout(n1299));
  jor  g0999(.dina(n1299), .dinb(n797), .dout(n1300));
  jand g1000(.dina(n1300), .dinb(n800), .dout(n1301));
  jand g1001(.dina(n1301), .dinb(n1298), .dout(n1302));
  jor  g1002(.dina(n797), .dinb(G40), .dout(n1303));
  jor  g1003(.dina(G4088), .dinb(G91), .dout(n1304));
  jand g1004(.dina(n1304), .dinb(G4087), .dout(n1305));
  jand g1005(.dina(n1305), .dinb(n1303), .dout(n1306));
  jor  g1006(.dina(n1306), .dinb(n1302), .dout(G742));
  jor  g1007(.dina(n1205), .dinb(G4089), .dout(n1308));
  jor  g1008(.dina(n1279), .dinb(n852), .dout(n1309));
  jand g1009(.dina(n1309), .dinb(n854), .dout(n1310));
  jand g1010(.dina(n1310), .dinb(n1308), .dout(n1311));
  jor  g1011(.dina(n852), .dinb(G49), .dout(n1312));
  jor  g1012(.dina(G4089), .dinb(G46), .dout(n1313));
  jand g1013(.dina(n1313), .dinb(G4090), .dout(n1314));
  jand g1014(.dina(n1314), .dinb(n1312), .dout(n1315));
  jor  g1015(.dina(n1315), .dinb(n1311), .dout(G772));
  jor  g1016(.dina(n1213), .dinb(G4089), .dout(n1317));
  jor  g1017(.dina(n1251), .dinb(n852), .dout(n1318));
  jand g1018(.dina(n1318), .dinb(n854), .dout(n1319));
  jand g1019(.dina(n1319), .dinb(n1317), .dout(n1320));
  jor  g1020(.dina(n852), .dinb(G103), .dout(n1321));
  jor  g1021(.dina(G4089), .dinb(G100), .dout(n1322));
  jand g1022(.dina(n1322), .dinb(G4090), .dout(n1323));
  jand g1023(.dina(n1323), .dinb(n1321), .dout(n1324));
  jor  g1024(.dina(n1324), .dinb(n1320), .dout(G777));
  jor  g1025(.dina(n1297), .dinb(G4089), .dout(n1326));
  jor  g1026(.dina(n1299), .dinb(n852), .dout(n1327));
  jand g1027(.dina(n1327), .dinb(n854), .dout(n1328));
  jand g1028(.dina(n1328), .dinb(n1326), .dout(n1329));
  jor  g1029(.dina(n852), .dinb(G40), .dout(n1330));
  jor  g1030(.dina(G4089), .dinb(G91), .dout(n1331));
  jand g1031(.dina(n1331), .dinb(G4090), .dout(n1332));
  jand g1032(.dina(n1332), .dinb(n1330), .dout(n1333));
  jor  g1033(.dina(n1333), .dinb(n1329), .dout(G782));
  jor  g1034(.dina(n1297), .dinb(G1689), .dout(n1335));
  jor  g1035(.dina(n1299), .dinb(n993), .dout(n1336));
  jand g1036(.dina(n1336), .dinb(n999), .dout(n1337));
  jand g1037(.dina(n1337), .dinb(n1335), .dout(n1338));
  jand g1038(.dina(n994), .dinb(G203), .dout(n1339));
  jand g1039(.dina(n996), .dinb(G173), .dout(n1340));
  jor  g1040(.dina(n1340), .dinb(n1339), .dout(n1341));
  jor  g1041(.dina(n1341), .dinb(n1338), .dout(n1342));
  jand g1042(.dina(n1342), .dinb(G137), .dout(G645));
  jor  g1043(.dina(n1251), .dinb(n993), .dout(n1344));
  jor  g1044(.dina(n1213), .dinb(G1689), .dout(n1345));
  jand g1045(.dina(n1345), .dinb(n999), .dout(n1346));
  jand g1046(.dina(n1346), .dinb(n1344), .dout(n1347));
  jand g1047(.dina(n994), .dinb(G197), .dout(n1348));
  jand g1048(.dina(n996), .dinb(G167), .dout(n1349));
  jor  g1049(.dina(n1349), .dinb(n1348), .dout(n1350));
  jor  g1050(.dina(n1350), .dinb(n1347), .dout(n1351));
  jand g1051(.dina(n1351), .dinb(G137), .dout(G648));
  jand g1052(.dina(n994), .dinb(G194), .dout(n1353));
  jand g1053(.dina(n996), .dinb(G164), .dout(n1354));
  jor  g1054(.dina(n1354), .dinb(n1353), .dout(n1355));
  jor  g1055(.dina(n1205), .dinb(G1689), .dout(n1356));
  jor  g1056(.dina(n1279), .dinb(n993), .dout(n1357));
  jand g1057(.dina(n1357), .dinb(n1356), .dout(n1358));
  jand g1058(.dina(n1358), .dinb(n999), .dout(n1359));
  jor  g1059(.dina(n1359), .dinb(n1355), .dout(n1360));
  jand g1060(.dina(n1360), .dinb(G137), .dout(G651));
  jand g1061(.dina(n994), .dinb(G191), .dout(n1362));
  jand g1062(.dina(n996), .dinb(G161), .dout(n1363));
  jor  g1063(.dina(n1363), .dinb(n1362), .dout(n1364));
  jor  g1064(.dina(n1196), .dinb(G1689), .dout(n1365));
  jor  g1065(.dina(n1236), .dinb(n993), .dout(n1366));
  jand g1066(.dina(n1366), .dinb(n1365), .dout(n1367));
  jand g1067(.dina(n1367), .dinb(n999), .dout(n1368));
  jor  g1068(.dina(n1368), .dinb(n1364), .dout(n1369));
  jand g1069(.dina(n1369), .dinb(G137), .dout(G654));
  jor  g1070(.dina(n1297), .dinb(G1691), .dout(n1371));
  jor  g1071(.dina(n1299), .dinb(n1008), .dout(n1372));
  jand g1072(.dina(n1372), .dinb(n1007), .dout(n1373));
  jand g1073(.dina(n1373), .dinb(n1371), .dout(n1374));
  jand g1074(.dina(n1014), .dinb(G203), .dout(n1375));
  jand g1075(.dina(n1012), .dinb(G173), .dout(n1376));
  jor  g1076(.dina(n1376), .dinb(n1375), .dout(n1377));
  jor  g1077(.dina(n1377), .dinb(n1374), .dout(n1378));
  jand g1078(.dina(n1378), .dinb(G137), .dout(G679));
  jand g1079(.dina(n1014), .dinb(G197), .dout(n1380));
  jand g1080(.dina(n1012), .dinb(G167), .dout(n1381));
  jor  g1081(.dina(n1381), .dinb(n1380), .dout(n1382));
  jor  g1082(.dina(n1213), .dinb(G1691), .dout(n1383));
  jor  g1083(.dina(n1251), .dinb(n1008), .dout(n1384));
  jand g1084(.dina(n1384), .dinb(n1383), .dout(n1385));
  jand g1085(.dina(n1385), .dinb(n1007), .dout(n1386));
  jor  g1086(.dina(n1386), .dinb(n1382), .dout(n1387));
  jand g1087(.dina(n1387), .dinb(G137), .dout(G682));
  jor  g1088(.dina(n1205), .dinb(G1691), .dout(n1389));
  jor  g1089(.dina(n1279), .dinb(n1008), .dout(n1390));
  jand g1090(.dina(n1390), .dinb(n1007), .dout(n1391));
  jand g1091(.dina(n1391), .dinb(n1389), .dout(n1392));
  jand g1092(.dina(n1014), .dinb(G194), .dout(n1393));
  jand g1093(.dina(n1012), .dinb(G164), .dout(n1394));
  jor  g1094(.dina(n1394), .dinb(n1393), .dout(n1395));
  jor  g1095(.dina(n1395), .dinb(n1392), .dout(n1396));
  jand g1096(.dina(n1396), .dinb(G137), .dout(G685));
  jor  g1097(.dina(n1236), .dinb(n1008), .dout(n1398));
  jor  g1098(.dina(n1196), .dinb(G1691), .dout(n1399));
  jand g1099(.dina(n1399), .dinb(n1007), .dout(n1400));
  jand g1100(.dina(n1400), .dinb(n1398), .dout(n1401));
  jand g1101(.dina(n1014), .dinb(G191), .dout(n1402));
  jand g1102(.dina(n1012), .dinb(G161), .dout(n1403));
  jor  g1103(.dina(n1403), .dinb(n1402), .dout(n1404));
  jor  g1104(.dina(n1404), .dinb(n1401), .dout(n1405));
  jand g1105(.dina(n1405), .dinb(G137), .dout(G688));
  jand g1106(.dina(n746), .dinb(n648), .dout(n1407));
  jxor g1107(.dina(n977), .dinb(n654), .dout(n1408));
  jxor g1108(.dina(n1408), .dinb(n644), .dout(n1409));
  jxor g1109(.dina(n1409), .dinb(n1407), .dout(n1410));
  jor  g1110(.dina(n1410), .dinb(n737), .dout(n1411));
  jnot g1111(.din(G2174), .dout(n1412));
  jnot g1112(.din(n719), .dout(n1413));
  jnot g1113(.din(n720), .dout(n1414));
  jor  g1114(.dina(n821), .dinb(n1414), .dout(n1415));
  jand g1115(.dina(n1415), .dinb(n1413), .dout(n1416));
  jxor g1116(.dina(n742), .dinb(n654), .dout(n1417));
  jxor g1117(.dina(n1417), .dinb(n792), .dout(n1418));
  jnot g1118(.din(n660), .dout(n1419));
  jand g1119(.dina(n745), .dinb(n648), .dout(n1420));
  jand g1120(.dina(n1420), .dinb(n1419), .dout(n1421));
  jxor g1121(.dina(n1421), .dinb(n1418), .dout(n1422));
  jor  g1122(.dina(n1422), .dinb(n1416), .dout(n1423));
  jand g1123(.dina(n1423), .dinb(n1412), .dout(n1424));
  jand g1124(.dina(n1424), .dinb(n1411), .dout(n1425));
  jnot g1125(.din(n1425), .dout(n1426));
  jnot g1126(.din(n641), .dout(n1427));
  jand g1127(.dina(n1416), .dinb(n1427), .dout(n1428));
  jor  g1128(.dina(n1428), .dinb(n1422), .dout(n1429));
  jnot g1129(.din(n1429), .dout(n1430));
  jnot g1130(.din(n1410), .dout(n1431));
  jand g1131(.dina(n1428), .dinb(n1431), .dout(n1432));
  jor  g1132(.dina(n1432), .dinb(n1412), .dout(n1433));
  jor  g1133(.dina(n1433), .dinb(n1430), .dout(n1434));
  jand g1134(.dina(n1434), .dinb(n1426), .dout(n1435));
  jor  g1135(.dina(n728), .dinb(n637), .dout(n1436));
  jxor g1136(.dina(n1436), .dinb(n733), .dout(n1437));
  jxor g1137(.dina(n1437), .dinb(n735), .dout(n1438));
  jor  g1138(.dina(n1438), .dinb(G2174), .dout(n1439));
  jor  g1139(.dina(n735), .dinb(n640), .dout(n1440));
  jor  g1140(.dina(n819), .dinb(n628), .dout(n1441));
  jor  g1141(.dina(n733), .dinb(n814), .dout(n1442));
  jor  g1142(.dina(n1442), .dinb(n639), .dout(n1443));
  jand g1143(.dina(n1443), .dinb(n1441), .dout(n1444));
  jxor g1144(.dina(n1444), .dinb(n1440), .dout(n1445));
  jor  g1145(.dina(n1445), .dinb(n1412), .dout(n1446));
  jand g1146(.dina(n1446), .dinb(n1439), .dout(n1447));
  jxor g1147(.dina(n620), .dinb(n618), .dout(n1448));
  jxor g1148(.dina(n767), .dinb(n624), .dout(n1449));
  jxor g1149(.dina(n1449), .dinb(n1448), .dout(n1450));
  jxor g1150(.dina(n1450), .dinb(n1447), .dout(n1451));
  jnot g1151(.din(n1451), .dout(n1452));
  jand g1152(.dina(n1452), .dinb(n1435), .dout(n1453));
  jor  g1153(.dina(n737), .dinb(n641), .dout(n1454));
  jor  g1154(.dina(n1454), .dinb(n1410), .dout(n1455));
  jand g1155(.dina(n1455), .dinb(G2174), .dout(n1456));
  jand g1156(.dina(n1456), .dinb(n1429), .dout(n1457));
  jor  g1157(.dina(n1457), .dinb(n1425), .dout(n1458));
  jand g1158(.dina(n1451), .dinb(n1458), .dout(n1459));
  jor  g1159(.dina(n1459), .dinb(n749), .dout(n1460));
  jor  g1160(.dina(n1460), .dinb(n1453), .dout(n1461));
  jand g1161(.dina(G351), .dinb(G248), .dout(n1462));
  jand g1162(.dina(n374), .dinb(G251), .dout(n1463));
  jor  g1163(.dina(n1463), .dinb(n377), .dout(n1464));
  jor  g1164(.dina(n1464), .dinb(n1462), .dout(n1465));
  jand g1165(.dina(n374), .dinb(n406), .dout(n1466));
  jand g1166(.dina(G351), .dinb(n408), .dout(n1467));
  jor  g1167(.dina(n1467), .dinb(n1466), .dout(n1468));
  jor  g1168(.dina(n1468), .dinb(G534), .dout(n1469));
  jand g1169(.dina(n1469), .dinb(n1465), .dout(n1470));
  jand g1170(.dina(G341), .dinb(G248), .dout(n1471));
  jand g1171(.dina(n387), .dinb(G251), .dout(n1472));
  jor  g1172(.dina(n1472), .dinb(n389), .dout(n1473));
  jor  g1173(.dina(n1473), .dinb(n1471), .dout(n1474));
  jand g1174(.dina(n387), .dinb(n406), .dout(n1475));
  jand g1175(.dina(G341), .dinb(n408), .dout(n1476));
  jor  g1176(.dina(n1476), .dinb(n1475), .dout(n1477));
  jor  g1177(.dina(n1477), .dinb(G523), .dout(n1478));
  jand g1178(.dina(n1478), .dinb(n1474), .dout(n1479));
  jxor g1179(.dina(n1479), .dinb(n1470), .dout(n1480));
  jor  g1180(.dina(n435), .dinb(n369), .dout(n1481));
  jor  g1181(.dina(G324), .dinb(n366), .dout(n1482));
  jand g1182(.dina(n1482), .dinb(G503), .dout(n1483));
  jand g1183(.dina(n1483), .dinb(n1481), .dout(n1484));
  jor  g1184(.dina(G324), .dinb(G254), .dout(n1485));
  jor  g1185(.dina(n435), .dinb(G242), .dout(n1486));
  jand g1186(.dina(n1486), .dinb(n1485), .dout(n1487));
  jand g1187(.dina(n1487), .dinb(n437), .dout(n1488));
  jor  g1188(.dina(n1488), .dinb(n1484), .dout(n1489));
  jor  g1189(.dina(G514), .dinb(n408), .dout(n1490));
  jor  g1190(.dina(n361), .dinb(G248), .dout(n1491));
  jand g1191(.dina(n1491), .dinb(n1490), .dout(n1492));
  jxor g1192(.dina(n1492), .dinb(n371), .dout(n1493));
  jxor g1193(.dina(n1493), .dinb(n1489), .dout(n1494));
  jxor g1194(.dina(n1494), .dinb(n1480), .dout(n1495));
  jxor g1195(.dina(n433), .dinb(n428), .dout(n1496));
  jxor g1196(.dina(n423), .dinb(n412), .dout(n1497));
  jxor g1197(.dina(n1497), .dinb(n1496), .dout(n1498));
  jxor g1198(.dina(n1498), .dinb(n1495), .dout(n1499));
  jand g1199(.dina(n1499), .dinb(n749), .dout(n1500));
  jnot g1200(.din(n1500), .dout(n1501));
  jand g1201(.dina(n1501), .dinb(n1461), .dout(n1502));
  jor  g1202(.dina(n1502), .dinb(G4092), .dout(n1503));
  jnot g1203(.din(n750), .dout(n1504));
  jor  g1204(.dina(n1504), .dinb(G120), .dout(n1505));
  jand g1205(.dina(n1505), .dinb(n1503), .dout(G843));
  jand g1206(.dina(G273), .dinb(G248), .dout(n1507));
  jand g1207(.dina(n471), .dinb(G251), .dout(n1508));
  jor  g1208(.dina(n1508), .dinb(n473), .dout(n1509));
  jor  g1209(.dina(n1509), .dinb(n1507), .dout(n1510));
  jand g1210(.dina(n471), .dinb(n406), .dout(n1511));
  jand g1211(.dina(G273), .dinb(n408), .dout(n1512));
  jor  g1212(.dina(n1512), .dinb(n1511), .dout(n1513));
  jor  g1213(.dina(n1513), .dinb(G411), .dout(n1514));
  jand g1214(.dina(n1514), .dinb(n1510), .dout(n1515));
  jand g1215(.dina(G281), .dinb(G248), .dout(n1516));
  jand g1216(.dina(n530), .dinb(G251), .dout(n1517));
  jor  g1217(.dina(n1517), .dinb(n532), .dout(n1518));
  jor  g1218(.dina(n1518), .dinb(n1516), .dout(n1519));
  jand g1219(.dina(n530), .dinb(n406), .dout(n1520));
  jand g1220(.dina(G281), .dinb(n408), .dout(n1521));
  jor  g1221(.dina(n1521), .dinb(n1520), .dout(n1522));
  jor  g1222(.dina(n1522), .dinb(G374), .dout(n1523));
  jand g1223(.dina(n1523), .dinb(n1519), .dout(n1524));
  jxor g1224(.dina(n1524), .dinb(n1515), .dout(n1525));
  jor  g1225(.dina(n483), .dinb(n369), .dout(n1526));
  jor  g1226(.dina(G265), .dinb(n366), .dout(n1527));
  jand g1227(.dina(n1527), .dinb(G400), .dout(n1528));
  jand g1228(.dina(n1528), .dinb(n1526), .dout(n1529));
  jor  g1229(.dina(G265), .dinb(G254), .dout(n1530));
  jor  g1230(.dina(n483), .dinb(G242), .dout(n1531));
  jand g1231(.dina(n1531), .dinb(n1530), .dout(n1532));
  jand g1232(.dina(n1532), .dinb(n485), .dout(n1533));
  jor  g1233(.dina(n1533), .dinb(n1529), .dout(n1534));
  jand g1234(.dina(G257), .dinb(G248), .dout(n1535));
  jand g1235(.dina(n518), .dinb(G251), .dout(n1536));
  jor  g1236(.dina(n1536), .dinb(n520), .dout(n1537));
  jor  g1237(.dina(n1537), .dinb(n1535), .dout(n1538));
  jand g1238(.dina(n518), .dinb(n406), .dout(n1539));
  jand g1239(.dina(G257), .dinb(n408), .dout(n1540));
  jor  g1240(.dina(n1540), .dinb(n1539), .dout(n1541));
  jor  g1241(.dina(n1541), .dinb(G389), .dout(n1542));
  jand g1242(.dina(n1542), .dinb(n1538), .dout(n1543));
  jand g1243(.dina(G248), .dinb(G234), .dout(n1544));
  jand g1244(.dina(G251), .dinb(n460), .dout(n1545));
  jor  g1245(.dina(n1545), .dinb(n462), .dout(n1546));
  jor  g1246(.dina(n1546), .dinb(n1544), .dout(n1547));
  jand g1247(.dina(n406), .dinb(n460), .dout(n1548));
  jand g1248(.dina(n408), .dinb(G234), .dout(n1549));
  jor  g1249(.dina(n1549), .dinb(n1548), .dout(n1550));
  jor  g1250(.dina(n1550), .dinb(G435), .dout(n1551));
  jand g1251(.dina(n1551), .dinb(n1547), .dout(n1552));
  jxor g1252(.dina(n1552), .dinb(n1543), .dout(n1553));
  jxor g1253(.dina(n1553), .dinb(n1534), .dout(n1554));
  jxor g1254(.dina(n1554), .dinb(n1525), .dout(n1555));
  jand g1255(.dina(G248), .dinb(G226), .dout(n1556));
  jand g1256(.dina(G251), .dinb(n494), .dout(n1557));
  jor  g1257(.dina(n1557), .dinb(n496), .dout(n1558));
  jor  g1258(.dina(n1558), .dinb(n1556), .dout(n1559));
  jand g1259(.dina(n406), .dinb(n494), .dout(n1560));
  jand g1260(.dina(n408), .dinb(G226), .dout(n1561));
  jor  g1261(.dina(n1561), .dinb(n1560), .dout(n1562));
  jor  g1262(.dina(n1562), .dinb(G422), .dout(n1563));
  jand g1263(.dina(n1563), .dinb(n1559), .dout(n1564));
  jxor g1264(.dina(n1564), .dinb(n551), .dout(n1565));
  jor  g1265(.dina(n369), .dinb(n507), .dout(n1566));
  jor  g1266(.dina(n366), .dinb(G218), .dout(n1567));
  jand g1267(.dina(n1567), .dinb(G468), .dout(n1568));
  jand g1268(.dina(n1568), .dinb(n1566), .dout(n1569));
  jor  g1269(.dina(G254), .dinb(G218), .dout(n1570));
  jor  g1270(.dina(G242), .dinb(n507), .dout(n1571));
  jand g1271(.dina(n1571), .dinb(n1570), .dout(n1572));
  jand g1272(.dina(n1572), .dinb(n509), .dout(n1573));
  jor  g1273(.dina(n1573), .dinb(n1569), .dout(n1574));
  jand g1274(.dina(G248), .dinb(G210), .dout(n1575));
  jand g1275(.dina(G251), .dinb(n449), .dout(n1576));
  jor  g1276(.dina(n1576), .dinb(n451), .dout(n1577));
  jor  g1277(.dina(n1577), .dinb(n1575), .dout(n1578));
  jand g1278(.dina(n406), .dinb(n449), .dout(n1579));
  jand g1279(.dina(n408), .dinb(G210), .dout(n1580));
  jor  g1280(.dina(n1580), .dinb(n1579), .dout(n1581));
  jor  g1281(.dina(n1581), .dinb(G457), .dout(n1582));
  jand g1282(.dina(n1582), .dinb(n1578), .dout(n1583));
  jxor g1283(.dina(n1583), .dinb(n1574), .dout(n1584));
  jxor g1284(.dina(n1584), .dinb(n1565), .dout(n1585));
  jxor g1285(.dina(n1585), .dinb(n1555), .dout(n1586));
  jand g1286(.dina(n1586), .dinb(n749), .dout(n1587));
  jnot g1287(.din(n1587), .dout(n1588));
  jand g1288(.dina(n573), .dinb(n567), .dout(n1589));
  jor  g1289(.dina(n1589), .dinb(n699), .dout(n1590));
  jnot g1290(.din(n559), .dout(n1591));
  jor  g1291(.dina(n1591), .dinb(n557), .dout(n1592));
  jand g1292(.dina(n1592), .dinb(n532), .dout(n1593));
  jnot g1293(.din(n1593), .dout(n1594));
  jor  g1294(.dina(n695), .dinb(n1594), .dout(n1595));
  jand g1295(.dina(n923), .dinb(n473), .dout(n1596));
  jor  g1296(.dina(n1596), .dinb(n1593), .dout(n1597));
  jand g1297(.dina(n1597), .dinb(n1595), .dout(n1598));
  jxor g1298(.dina(n1598), .dinb(n1590), .dout(n1599));
  jnot g1299(.din(n1599), .dout(n1600));
  jnot g1300(.din(n686), .dout(n1601));
  jnot g1301(.din(n687), .dout(n1602));
  jor  g1302(.dina(n1592), .dinb(n532), .dout(n1603));
  jor  g1303(.dina(n1596), .dinb(n1603), .dout(n1604));
  jor  g1304(.dina(n923), .dinb(n473), .dout(n1605));
  jor  g1305(.dina(n689), .dinb(n485), .dout(n1606));
  jand g1306(.dina(n1606), .dinb(n1605), .dout(n1607));
  jand g1307(.dina(n1607), .dinb(n1604), .dout(n1608));
  jor  g1308(.dina(n1608), .dinb(n690), .dout(n1609));
  jor  g1309(.dina(n1609), .dinb(n1602), .dout(n1610));
  jand g1310(.dina(n1610), .dinb(n1601), .dout(n1611));
  jand g1311(.dina(n1611), .dinb(n581), .dout(n1612));
  jxor g1312(.dina(n566), .dinb(n561), .dout(n1613));
  jxor g1313(.dina(n1613), .dinb(n865), .dout(n1614));
  jxor g1314(.dina(n1614), .dinb(n1612), .dout(n1615));
  jnot g1315(.din(n1615), .dout(n1616));
  jand g1316(.dina(n1616), .dinb(n1600), .dout(n1617));
  jnot g1317(.din(G1497), .dout(n1618));
  jand g1318(.dina(n1615), .dinb(n1599), .dout(n1619));
  jor  g1319(.dina(n1619), .dinb(n1618), .dout(n1620));
  jor  g1320(.dina(n1620), .dinb(n1617), .dout(n1621));
  jand g1321(.dina(n1605), .dinb(n1603), .dout(n1622));
  jor  g1322(.dina(n1622), .dinb(n694), .dout(n1623));
  jxor g1323(.dina(n1613), .dinb(n1609), .dout(n1624));
  jxor g1324(.dina(n1624), .dinb(n1623), .dout(n1625));
  jxor g1325(.dina(n1611), .dinb(n865), .dout(n1626));
  jxor g1326(.dina(n1626), .dinb(n1625), .dout(n1627));
  jor  g1327(.dina(n1627), .dinb(G1497), .dout(n1628));
  jand g1328(.dina(n1628), .dinb(n1621), .dout(n1629));
  jxor g1329(.dina(n579), .dinb(n574), .dout(n1630));
  jxor g1330(.dina(n1630), .dinb(n1629), .dout(n1631));
  jnot g1331(.din(n709), .dout(n1632));
  jand g1332(.dina(n1632), .dinb(n953), .dout(n1633));
  jand g1333(.dina(n711), .dinb(n954), .dout(n1634));
  jor  g1334(.dina(n1634), .dinb(n1633), .dout(n1635));
  jxor g1335(.dina(n608), .dinb(n592), .dout(n1636));
  jxor g1336(.dina(n1636), .dinb(n602), .dout(n1637));
  jxor g1337(.dina(n1637), .dinb(n1635), .dout(n1638));
  jor  g1338(.dina(n938), .dinb(n597), .dout(n1639));
  jand g1339(.dina(n609), .dinb(n962), .dout(n1640));
  jor  g1340(.dina(n1640), .dinb(n715), .dout(n1641));
  jand g1341(.dina(n1641), .dinb(n1639), .dout(n1642));
  jxor g1342(.dina(n1642), .dinb(n1638), .dout(n1643));
  jand g1343(.dina(n1643), .dinb(n703), .dout(n1644));
  jnot g1344(.din(n682), .dout(n1645));
  jor  g1345(.dina(n1611), .dinb(n684), .dout(n1646));
  jand g1346(.dina(n1646), .dinb(n1645), .dout(n1647));
  jand g1347(.dina(n713), .dinb(n954), .dout(n1648));
  jor  g1348(.dina(n1648), .dinb(n1633), .dout(n1649));
  jxor g1349(.dina(n1649), .dinb(n938), .dout(n1650));
  jxor g1350(.dina(n1650), .dinb(n1637), .dout(n1651));
  jand g1351(.dina(n1651), .dinb(n1647), .dout(n1652));
  jor  g1352(.dina(n1652), .dinb(n1644), .dout(n1653));
  jor  g1353(.dina(n1653), .dinb(G1497), .dout(n1654));
  jnot g1354(.din(n588), .dout(n1655));
  jand g1355(.dina(n1652), .dinb(n1655), .dout(n1656));
  jor  g1356(.dina(n703), .dinb(n588), .dout(n1657));
  jand g1357(.dina(n1657), .dinb(n1643), .dout(n1658));
  jor  g1358(.dina(n1658), .dinb(n1656), .dout(n1659));
  jor  g1359(.dina(n1659), .dinb(n1618), .dout(n1660));
  jand g1360(.dina(n1660), .dinb(n1654), .dout(n1661));
  jxor g1361(.dina(n1661), .dinb(n1631), .dout(n1662));
  jor  g1362(.dina(n1662), .dinb(n749), .dout(n1663));
  jand g1363(.dina(n1663), .dinb(n1588), .dout(n1664));
  jor  g1364(.dina(n1664), .dinb(G4092), .dout(n1665));
  jor  g1365(.dina(n1504), .dinb(G118), .dout(n1666));
  jand g1366(.dina(n1666), .dinb(n1665), .dout(G882));
  jor  g1367(.dina(G4088), .dinb(G14), .dout(n1668));
  jor  g1368(.dina(n797), .dinb(G64), .dout(n1669));
  jand g1369(.dina(n1669), .dinb(G4087), .dout(n1670));
  jand g1370(.dina(n1670), .dinb(n1668), .dout(n1671));
  jand g1371(.dina(G4092), .dinb(G97), .dout(n1672));
  jnot g1372(.din(n1672), .dout(n1673));
  jand g1373(.dina(n1673), .dinb(n1665), .dout(n1674));
  jnot g1374(.din(n1674), .dout(n1675));
  jor  g1375(.dina(n1675), .dinb(n797), .dout(n1676));
  jand g1376(.dina(G4092), .dinb(G94), .dout(n1677));
  jnot g1377(.din(n1677), .dout(n1678));
  jand g1378(.dina(n1678), .dinb(n1503), .dout(n1679));
  jnot g1379(.din(n1679), .dout(n1680));
  jor  g1380(.dina(n1680), .dinb(G4088), .dout(n1681));
  jand g1381(.dina(n1681), .dinb(n800), .dout(n1682));
  jand g1382(.dina(n1682), .dinb(n1676), .dout(n1683));
  jor  g1383(.dina(n1683), .dinb(n1671), .dout(G767));
  jor  g1384(.dina(G4089), .dinb(G14), .dout(n1685));
  jor  g1385(.dina(n852), .dinb(G64), .dout(n1686));
  jand g1386(.dina(n1686), .dinb(G4090), .dout(n1687));
  jand g1387(.dina(n1687), .dinb(n1685), .dout(n1688));
  jor  g1388(.dina(n1675), .dinb(n852), .dout(n1689));
  jor  g1389(.dina(n1680), .dinb(G4089), .dout(n1690));
  jand g1390(.dina(n1690), .dinb(n854), .dout(n1691));
  jand g1391(.dina(n1691), .dinb(n1689), .dout(n1692));
  jor  g1392(.dina(n1692), .dinb(n1688), .dout(G807));
  jnot g1393(.din(G137), .dout(n1694));
  jnot g1394(.din(G179), .dout(n1695));
  jnot g1395(.din(n996), .dout(n1696));
  jor  g1396(.dina(n1696), .dinb(n1695), .dout(n1697));
  jnot g1397(.din(G176), .dout(n1698));
  jnot g1398(.din(n994), .dout(n1699));
  jor  g1399(.dina(n1699), .dinb(n1698), .dout(n1700));
  jand g1400(.dina(n1674), .dinb(G1689), .dout(n1701));
  jand g1401(.dina(n1679), .dinb(n993), .dout(n1702));
  jor  g1402(.dina(n1702), .dinb(G1690), .dout(n1703));
  jor  g1403(.dina(n1703), .dinb(n1701), .dout(n1704));
  jand g1404(.dina(n1704), .dinb(n1700), .dout(n1705));
  jand g1405(.dina(n1705), .dinb(n1697), .dout(n1706));
  jor  g1406(.dina(n1706), .dinb(n1694), .dout(G658));
  jnot g1407(.din(n1012), .dout(n1708));
  jor  g1408(.dina(n1708), .dinb(n1695), .dout(n1709));
  jnot g1409(.din(n1014), .dout(n1710));
  jor  g1410(.dina(n1710), .dinb(n1698), .dout(n1711));
  jand g1411(.dina(n1674), .dinb(G1691), .dout(n1712));
  jand g1412(.dina(n1679), .dinb(n1008), .dout(n1713));
  jor  g1413(.dina(n1713), .dinb(G1694), .dout(n1714));
  jor  g1414(.dina(n1714), .dinb(n1712), .dout(n1715));
  jand g1415(.dina(n1715), .dinb(n1711), .dout(n1716));
  jand g1416(.dina(n1716), .dinb(n1709), .dout(n1717));
  jor  g1417(.dina(n1717), .dinb(n1694), .dout(G690));
  jdff  g1418(.din(G141), .dout(G144));
  jdff  g1419(.din(G293), .dout(G298));
  jdff  g1420(.din(G3173), .dout(G973));
  jnot g1421(.din(G545), .dout(G603));
  jnot g1422(.din(G545), .dout(G604));
  jdff  g1423(.din(G137), .dout(G926));
  jdff  g1424(.din(G141), .dout(G923));
  jdff  g1425(.din(G1), .dout(G921));
  jdff  g1426(.din(G549), .dout(G892));
  jdff  g1427(.din(G299), .dout(G887));
  jnot g1428(.din(G549), .dout(G606));
  jdff  g1429(.din(G1), .dout(G993));
  jdff  g1430(.din(G1), .dout(G978));
  jdff  g1431(.din(G1), .dout(G949));
  jdff  g1432(.din(G1), .dout(G939));
  jdff  g1433(.din(G299), .dout(G889));
  jor  g1434(.dina(n336), .dinb(n333), .dout(G717));
  jand g1435(.dina(n661), .dinb(n641), .dout(G626));
  jand g1436(.dina(n611), .dinb(n588), .dout(G632));
  jor  g1437(.dina(n717), .dinb(n704), .dout(G621));
  jor  g1438(.dina(n747), .dinb(n738), .dout(G629));
endmodule


