/*

c3540:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jcb: 374
	jdff: 1453
	jand: 535

Summary:
	jxor: 37
	jspl: 206
	jspl3: 356
	jnot: 173
	jcb: 374
	jdff: 1453
	jand: 535
*/

module c3540(gclk, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402);
	input gclk;
	input G1;
	input G13;
	input G20;
	input G33;
	input G41;
	input G45;
	input G50;
	input G58;
	input G68;
	input G77;
	input G87;
	input G97;
	input G107;
	input G116;
	input G124;
	input G125;
	input G128;
	input G132;
	input G137;
	input G143;
	input G150;
	input G159;
	input G169;
	input G179;
	input G190;
	input G200;
	input G213;
	input G222;
	input G223;
	input G226;
	input G232;
	input G238;
	input G244;
	input G250;
	input G257;
	input G264;
	input G270;
	input G274;
	input G283;
	input G294;
	input G303;
	input G311;
	input G317;
	input G322;
	input G326;
	input G329;
	input G330;
	input G343;
	input G1698;
	input G2897;
	output G353;
	output G355;
	output G361;
	output G358;
	output G351;
	output G372;
	output G369;
	output G399;
	output G364;
	output G396;
	output G384;
	output G367;
	output G387;
	output G393;
	output G390;
	output G378;
	output G375;
	output G381;
	output G407;
	output G409;
	output G405;
	output G402;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [2:0] w_G1_2;
	wire [1:0] w_G1_3;
	wire [2:0] w_G13_0;
	wire [1:0] w_G13_1;
	wire [2:0] w_G20_0;
	wire [2:0] w_G20_1;
	wire [2:0] w_G20_2;
	wire [2:0] w_G20_3;
	wire [2:0] w_G20_4;
	wire [2:0] w_G20_5;
	wire [2:0] w_G20_6;
	wire [1:0] w_G20_7;
	wire [2:0] w_G33_0;
	wire [2:0] w_G33_1;
	wire [2:0] w_G33_2;
	wire [2:0] w_G33_3;
	wire [2:0] w_G33_4;
	wire [2:0] w_G33_5;
	wire [2:0] w_G33_6;
	wire [2:0] w_G33_7;
	wire [2:0] w_G33_8;
	wire [2:0] w_G33_9;
	wire [2:0] w_G33_10;
	wire [2:0] w_G33_11;
	wire [2:0] w_G41_0;
	wire [1:0] w_G41_1;
	wire [2:0] w_G45_0;
	wire [2:0] w_G45_1;
	wire [2:0] w_G50_0;
	wire [2:0] w_G50_1;
	wire [2:0] w_G50_2;
	wire [2:0] w_G50_3;
	wire [2:0] w_G50_4;
	wire [2:0] w_G50_5;
	wire [2:0] w_G58_0;
	wire [2:0] w_G58_1;
	wire [2:0] w_G58_2;
	wire [2:0] w_G58_3;
	wire [2:0] w_G58_4;
	wire [1:0] w_G58_5;
	wire [2:0] w_G68_0;
	wire [2:0] w_G68_1;
	wire [2:0] w_G68_2;
	wire [2:0] w_G68_3;
	wire [2:0] w_G68_4;
	wire [1:0] w_G68_5;
	wire [2:0] w_G77_0;
	wire [2:0] w_G77_1;
	wire [2:0] w_G77_2;
	wire [2:0] w_G77_3;
	wire [2:0] w_G77_4;
	wire [1:0] w_G77_5;
	wire [2:0] w_G87_0;
	wire [2:0] w_G87_1;
	wire [2:0] w_G87_2;
	wire [2:0] w_G87_3;
	wire [2:0] w_G97_0;
	wire [2:0] w_G97_1;
	wire [2:0] w_G97_2;
	wire [2:0] w_G97_3;
	wire [2:0] w_G97_4;
	wire [1:0] w_G97_5;
	wire [2:0] w_G107_0;
	wire [2:0] w_G107_1;
	wire [2:0] w_G107_2;
	wire [2:0] w_G107_3;
	wire [2:0] w_G107_4;
	wire [1:0] w_G107_5;
	wire [2:0] w_G116_0;
	wire [2:0] w_G116_1;
	wire [2:0] w_G116_2;
	wire [2:0] w_G116_3;
	wire [2:0] w_G116_4;
	wire [1:0] w_G125_0;
	wire [2:0] w_G128_0;
	wire [2:0] w_G132_0;
	wire [1:0] w_G132_1;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G143_0;
	wire [2:0] w_G143_1;
	wire [1:0] w_G143_2;
	wire [2:0] w_G150_0;
	wire [2:0] w_G150_1;
	wire [2:0] w_G150_2;
	wire [1:0] w_G150_3;
	wire [2:0] w_G159_0;
	wire [2:0] w_G159_1;
	wire [2:0] w_G159_2;
	wire [2:0] w_G159_3;
	wire [2:0] w_G169_0;
	wire [1:0] w_G169_1;
	wire [2:0] w_G179_0;
	wire [2:0] w_G179_1;
	wire [2:0] w_G179_2;
	wire [2:0] w_G190_0;
	wire [2:0] w_G190_1;
	wire [2:0] w_G190_2;
	wire [2:0] w_G190_3;
	wire [1:0] w_G190_4;
	wire [2:0] w_G200_0;
	wire [2:0] w_G200_1;
	wire [2:0] w_G200_2;
	wire [2:0] w_G200_3;
	wire [2:0] w_G200_4;
	wire [2:0] w_G213_0;
	wire [1:0] w_G223_0;
	wire [2:0] w_G226_0;
	wire [1:0] w_G226_1;
	wire [2:0] w_G232_0;
	wire [2:0] w_G232_1;
	wire [2:0] w_G238_0;
	wire [2:0] w_G238_1;
	wire [2:0] w_G244_0;
	wire [2:0] w_G244_1;
	wire [2:0] w_G250_0;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [2:0] w_G264_0;
	wire [1:0] w_G264_1;
	wire [2:0] w_G270_0;
	wire [2:0] w_G274_0;
	wire [2:0] w_G283_0;
	wire [2:0] w_G283_1;
	wire [2:0] w_G283_2;
	wire [2:0] w_G283_3;
	wire [2:0] w_G294_0;
	wire [2:0] w_G294_1;
	wire [2:0] w_G294_2;
	wire [1:0] w_G294_3;
	wire [2:0] w_G303_0;
	wire [2:0] w_G303_1;
	wire [2:0] w_G303_2;
	wire [2:0] w_G311_0;
	wire [2:0] w_G311_1;
	wire [2:0] w_G317_0;
	wire [1:0] w_G317_1;
	wire [2:0] w_G322_0;
	wire [1:0] w_G326_0;
	wire [1:0] w_G330_0;
	wire [1:0] w_G343_0;
	wire [2:0] w_G1698_0;
	wire w_G355_0;
	wire G355_fa_;
	wire [1:0] w_G396_0;
	wire G396_fa_;
	wire w_G384_0;
	wire G384_fa_;
	wire [1:0] w_G387_0;
	wire G387_fa_;
	wire [2:0] w_n72_0;
	wire [1:0] w_n72_1;
	wire [2:0] w_n73_0;
	wire [2:0] w_n73_1;
	wire [2:0] w_n73_2;
	wire [2:0] w_n74_0;
	wire [1:0] w_n74_1;
	wire [2:0] w_n75_0;
	wire [1:0] w_n75_1;
	wire [1:0] w_n76_0;
	wire [1:0] w_n77_0;
	wire [2:0] w_n79_0;
	wire [2:0] w_n80_0;
	wire [1:0] w_n80_1;
	wire [2:0] w_n81_0;
	wire [2:0] w_n85_0;
	wire [1:0] w_n86_0;
	wire [2:0] w_n88_0;
	wire [1:0] w_n88_1;
	wire [2:0] w_n91_0;
	wire [2:0] w_n91_1;
	wire [1:0] w_n93_0;
	wire [2:0] w_n97_0;
	wire [2:0] w_n97_1;
	wire [1:0] w_n97_2;
	wire [2:0] w_n98_0;
	wire [2:0] w_n98_1;
	wire [1:0] w_n98_2;
	wire [2:0] w_n103_0;
	wire [2:0] w_n105_0;
	wire [2:0] w_n105_1;
	wire [1:0] w_n105_2;
	wire [1:0] w_n106_0;
	wire [2:0] w_n112_0;
	wire [2:0] w_n112_1;
	wire [2:0] w_n112_2;
	wire [2:0] w_n112_3;
	wire [2:0] w_n112_4;
	wire [2:0] w_n112_5;
	wire [2:0] w_n113_0;
	wire [2:0] w_n113_1;
	wire [2:0] w_n113_2;
	wire [1:0] w_n113_3;
	wire [2:0] w_n114_0;
	wire [2:0] w_n114_1;
	wire [2:0] w_n115_0;
	wire [1:0] w_n115_1;
	wire [1:0] w_n116_0;
	wire [2:0] w_n118_0;
	wire [2:0] w_n121_0;
	wire [2:0] w_n122_0;
	wire [1:0] w_n122_1;
	wire [2:0] w_n123_0;
	wire [2:0] w_n123_1;
	wire [1:0] w_n131_0;
	wire [1:0] w_n135_0;
	wire [2:0] w_n137_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n144_0;
	wire [2:0] w_n146_0;
	wire [2:0] w_n146_1;
	wire [2:0] w_n146_2;
	wire [2:0] w_n146_3;
	wire [2:0] w_n147_0;
	wire [2:0] w_n148_0;
	wire [2:0] w_n148_1;
	wire [2:0] w_n148_2;
	wire [2:0] w_n148_3;
	wire [2:0] w_n148_4;
	wire [2:0] w_n148_5;
	wire [2:0] w_n148_6;
	wire [2:0] w_n148_7;
	wire [2:0] w_n148_8;
	wire [2:0] w_n148_9;
	wire [2:0] w_n149_0;
	wire [2:0] w_n149_1;
	wire [1:0] w_n149_2;
	wire [2:0] w_n151_0;
	wire [2:0] w_n151_1;
	wire [2:0] w_n151_2;
	wire [2:0] w_n151_3;
	wire [2:0] w_n151_4;
	wire [2:0] w_n152_0;
	wire [2:0] w_n152_1;
	wire [2:0] w_n152_2;
	wire [1:0] w_n152_3;
	wire [1:0] w_n154_0;
	wire [2:0] w_n155_0;
	wire [2:0] w_n155_1;
	wire [2:0] w_n155_2;
	wire [1:0] w_n155_3;
	wire [2:0] w_n157_0;
	wire [2:0] w_n161_0;
	wire [1:0] w_n161_1;
	wire [2:0] w_n162_0;
	wire [1:0] w_n163_0;
	wire [2:0] w_n166_0;
	wire [2:0] w_n166_1;
	wire [2:0] w_n166_2;
	wire [1:0] w_n166_3;
	wire [2:0] w_n170_0;
	wire [1:0] w_n172_0;
	wire [2:0] w_n179_0;
	wire [2:0] w_n179_1;
	wire [1:0] w_n180_0;
	wire [2:0] w_n185_0;
	wire [2:0] w_n185_1;
	wire [2:0] w_n185_2;
	wire [2:0] w_n185_3;
	wire [2:0] w_n189_0;
	wire [2:0] w_n189_1;
	wire [1:0] w_n189_2;
	wire [2:0] w_n190_0;
	wire [2:0] w_n190_1;
	wire [2:0] w_n191_0;
	wire [1:0] w_n195_0;
	wire [2:0] w_n196_0;
	wire [2:0] w_n196_1;
	wire [2:0] w_n196_2;
	wire [2:0] w_n197_0;
	wire [1:0] w_n197_1;
	wire [2:0] w_n199_0;
	wire [1:0] w_n199_1;
	wire [1:0] w_n201_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n206_0;
	wire [2:0] w_n210_0;
	wire [1:0] w_n213_0;
	wire [1:0] w_n214_0;
	wire [1:0] w_n218_0;
	wire [1:0] w_n219_0;
	wire [2:0] w_n221_0;
	wire [1:0] w_n228_0;
	wire [2:0] w_n229_0;
	wire [1:0] w_n230_0;
	wire [2:0] w_n231_0;
	wire [2:0] w_n234_0;
	wire [1:0] w_n241_0;
	wire [2:0] w_n242_0;
	wire [2:0] w_n243_0;
	wire [2:0] w_n246_0;
	wire [1:0] w_n246_1;
	wire [1:0] w_n249_0;
	wire [1:0] w_n255_0;
	wire [1:0] w_n257_0;
	wire [1:0] w_n259_0;
	wire [1:0] w_n261_0;
	wire [1:0] w_n262_0;
	wire [2:0] w_n269_0;
	wire [2:0] w_n269_1;
	wire [1:0] w_n270_0;
	wire [2:0] w_n271_0;
	wire [2:0] w_n271_1;
	wire [2:0] w_n274_0;
	wire [1:0] w_n278_0;
	wire [1:0] w_n279_0;
	wire [1:0] w_n281_0;
	wire [2:0] w_n288_0;
	wire [1:0] w_n288_1;
	wire [1:0] w_n296_0;
	wire [1:0] w_n298_0;
	wire [1:0] w_n300_0;
	wire [1:0] w_n303_0;
	wire [2:0] w_n312_0;
	wire [1:0] w_n312_1;
	wire [1:0] w_n315_0;
	wire [1:0] w_n320_0;
	wire [1:0] w_n324_0;
	wire [1:0] w_n328_0;
	wire [1:0] w_n334_0;
	wire [1:0] w_n339_0;
	wire [2:0] w_n346_0;
	wire [1:0] w_n346_1;
	wire [2:0] w_n355_0;
	wire [1:0] w_n355_1;
	wire [1:0] w_n362_0;
	wire [2:0] w_n367_0;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n374_0;
	wire [1:0] w_n381_0;
	wire [2:0] w_n382_0;
	wire [1:0] w_n382_1;
	wire [2:0] w_n385_0;
	wire [1:0] w_n385_1;
	wire [2:0] w_n387_0;
	wire [1:0] w_n387_1;
	wire [1:0] w_n390_0;
	wire [2:0] w_n401_0;
	wire [2:0] w_n404_0;
	wire [1:0] w_n405_0;
	wire [2:0] w_n407_0;
	wire [2:0] w_n407_1;
	wire [1:0] w_n407_2;
	wire [1:0] w_n412_0;
	wire [2:0] w_n420_0;
	wire [1:0] w_n420_1;
	wire [2:0] w_n425_0;
	wire [2:0] w_n425_1;
	wire [1:0] w_n426_0;
	wire [1:0] w_n430_0;
	wire [2:0] w_n436_0;
	wire [2:0] w_n439_0;
	wire [1:0] w_n439_1;
	wire [1:0] w_n445_0;
	wire [1:0] w_n446_0;
	wire [2:0] w_n455_0;
	wire [2:0] w_n462_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n474_0;
	wire [1:0] w_n475_0;
	wire [1:0] w_n478_0;
	wire [1:0] w_n479_0;
	wire [1:0] w_n483_0;
	wire [1:0] w_n484_0;
	wire [2:0] w_n492_0;
	wire [1:0] w_n507_0;
	wire [1:0] w_n508_0;
	wire [1:0] w_n511_0;
	wire [1:0] w_n512_0;
	wire [1:0] w_n516_0;
	wire [1:0] w_n517_0;
	wire [2:0] w_n519_0;
	wire [2:0] w_n519_1;
	wire [1:0] w_n523_0;
	wire [1:0] w_n524_0;
	wire [1:0] w_n528_0;
	wire [1:0] w_n532_0;
	wire [1:0] w_n534_0;
	wire [2:0] w_n536_0;
	wire [1:0] w_n539_0;
	wire [1:0] w_n541_0;
	wire [2:0] w_n542_0;
	wire [1:0] w_n543_0;
	wire [2:0] w_n548_0;
	wire [1:0] w_n550_0;
	wire [2:0] w_n552_0;
	wire [1:0] w_n552_1;
	wire [2:0] w_n553_0;
	wire [2:0] w_n553_1;
	wire [2:0] w_n553_2;
	wire [2:0] w_n554_0;
	wire [2:0] w_n554_1;
	wire [2:0] w_n554_2;
	wire [2:0] w_n554_3;
	wire [1:0] w_n556_0;
	wire [1:0] w_n557_0;
	wire [2:0] w_n561_0;
	wire [2:0] w_n563_0;
	wire [1:0] w_n564_0;
	wire [1:0] w_n565_0;
	wire [1:0] w_n567_0;
	wire [2:0] w_n571_0;
	wire [2:0] w_n572_0;
	wire [2:0] w_n573_0;
	wire [2:0] w_n576_0;
	wire [1:0] w_n576_1;
	wire [2:0] w_n588_0;
	wire [1:0] w_n588_1;
	wire [2:0] w_n589_0;
	wire [2:0] w_n589_1;
	wire [2:0] w_n591_0;
	wire [1:0] w_n591_1;
	wire [2:0] w_n592_0;
	wire [2:0] w_n592_1;
	wire [1:0] w_n592_2;
	wire [2:0] w_n593_0;
	wire [1:0] w_n602_0;
	wire [2:0] w_n603_0;
	wire [2:0] w_n603_1;
	wire [1:0] w_n603_2;
	wire [2:0] w_n604_0;
	wire [2:0] w_n604_1;
	wire [1:0] w_n604_2;
	wire [2:0] w_n605_0;
	wire [2:0] w_n605_1;
	wire [2:0] w_n608_0;
	wire [2:0] w_n608_1;
	wire [2:0] w_n612_0;
	wire [2:0] w_n612_1;
	wire [2:0] w_n612_2;
	wire [2:0] w_n612_3;
	wire [1:0] w_n612_4;
	wire [2:0] w_n613_0;
	wire [1:0] w_n613_1;
	wire [1:0] w_n615_0;
	wire [1:0] w_n616_0;
	wire [2:0] w_n617_0;
	wire [2:0] w_n617_1;
	wire [2:0] w_n617_2;
	wire [2:0] w_n617_3;
	wire [2:0] w_n617_4;
	wire [2:0] w_n617_5;
	wire [1:0] w_n617_6;
	wire [1:0] w_n619_0;
	wire [1:0] w_n622_0;
	wire [2:0] w_n623_0;
	wire [2:0] w_n623_1;
	wire [2:0] w_n623_2;
	wire [2:0] w_n623_3;
	wire [2:0] w_n623_4;
	wire [1:0] w_n623_5;
	wire [1:0] w_n626_0;
	wire [2:0] w_n627_0;
	wire [2:0] w_n627_1;
	wire [2:0] w_n627_2;
	wire [2:0] w_n627_3;
	wire [2:0] w_n627_4;
	wire [2:0] w_n627_5;
	wire [2:0] w_n627_6;
	wire [1:0] w_n627_7;
	wire [2:0] w_n631_0;
	wire [2:0] w_n631_1;
	wire [2:0] w_n631_2;
	wire [2:0] w_n631_3;
	wire [2:0] w_n631_4;
	wire [2:0] w_n631_5;
	wire [2:0] w_n631_6;
	wire [1:0] w_n631_7;
	wire [2:0] w_n634_0;
	wire [2:0] w_n634_1;
	wire [2:0] w_n634_2;
	wire [2:0] w_n634_3;
	wire [1:0] w_n634_4;
	wire [2:0] w_n636_0;
	wire [2:0] w_n636_1;
	wire [2:0] w_n636_2;
	wire [2:0] w_n636_3;
	wire [2:0] w_n636_4;
	wire [2:0] w_n636_5;
	wire [2:0] w_n636_6;
	wire [1:0] w_n636_7;
	wire [1:0] w_n639_0;
	wire [2:0] w_n640_0;
	wire [2:0] w_n640_1;
	wire [2:0] w_n640_2;
	wire [2:0] w_n640_3;
	wire [2:0] w_n640_4;
	wire [2:0] w_n640_5;
	wire [2:0] w_n640_6;
	wire [1:0] w_n640_7;
	wire [2:0] w_n642_0;
	wire [2:0] w_n642_1;
	wire [2:0] w_n642_2;
	wire [2:0] w_n642_3;
	wire [2:0] w_n642_4;
	wire [2:0] w_n642_5;
	wire [2:0] w_n642_6;
	wire [1:0] w_n642_7;
	wire [1:0] w_n654_0;
	wire [1:0] w_n657_0;
	wire [1:0] w_n661_0;
	wire [2:0] w_n672_0;
	wire [1:0] w_n672_1;
	wire [2:0] w_n675_0;
	wire [1:0] w_n676_0;
	wire [1:0] w_n680_0;
	wire [1:0] w_n692_0;
	wire [2:0] w_n696_0;
	wire [2:0] w_n696_1;
	wire [1:0] w_n717_0;
	wire [1:0] w_n728_0;
	wire [2:0] w_n743_0;
	wire [1:0] w_n743_1;
	wire [1:0] w_n750_0;
	wire [1:0] w_n754_0;
	wire [2:0] w_n758_0;
	wire [1:0] w_n758_1;
	wire [1:0] w_n759_0;
	wire [1:0] w_n760_0;
	wire [2:0] w_n764_0;
	wire [2:0] w_n764_1;
	wire [1:0] w_n769_0;
	wire [2:0] w_n771_0;
	wire [1:0] w_n779_0;
	wire [1:0] w_n797_0;
	wire [1:0] w_n801_0;
	wire [1:0] w_n816_0;
	wire [1:0] w_n823_0;
	wire [1:0] w_n825_0;
	wire [2:0] w_n853_0;
	wire [2:0] w_n855_0;
	wire [2:0] w_n861_0;
	wire [1:0] w_n861_1;
	wire [1:0] w_n863_0;
	wire [1:0] w_n864_0;
	wire [1:0] w_n899_0;
	wire [1:0] w_n909_0;
	wire [2:0] w_n937_0;
	wire [1:0] w_n940_0;
	wire [1:0] w_n962_0;
	wire [2:0] w_n988_0;
	wire [1:0] w_n990_0;
	wire [2:0] w_n991_0;
	wire [1:0] w_n992_0;
	wire [2:0] w_n994_0;
	wire [2:0] w_n996_0;
	wire [1:0] w_n999_0;
	wire [2:0] w_n1001_0;
	wire [2:0] w_n1002_0;
	wire [1:0] w_n1003_0;
	wire [2:0] w_n1049_0;
	wire [1:0] w_n1052_0;
	wire [1:0] w_n1057_0;
	wire [1:0] w_n1059_0;
	wire [1:0] w_n1088_0;
	wire [2:0] w_n1114_0;
	wire [2:0] w_n1162_0;
	wire [1:0] w_n1164_0;
	wire [1:0] w_n1172_0;
	wire [1:0] w_n1175_0;
	wire [1:0] w_n1183_0;
	wire [1:0] w_n1184_0;
	wire [1:0] w_n1187_0;
	wire w_dff_B_DHAEC3iB8_1;
	wire w_dff_B_b8xM2L0C0_1;
	wire w_dff_B_2uIT0MVQ7_0;
	wire w_dff_B_9UNlZxYu7_0;
	wire w_dff_B_g1FTjHUN6_0;
	wire w_dff_A_DG2xMPmt0_1;
	wire w_dff_A_SxUhH09K8_1;
	wire w_dff_A_coblnMg10_0;
	wire w_dff_B_Do0q7fth3_0;
	wire w_dff_B_SXT2Zkzf9_0;
	wire w_dff_B_CjykkLot3_0;
	wire w_dff_B_Rv7m2esg3_0;
	wire w_dff_B_LfoSC3jf1_0;
	wire w_dff_B_RwFA02SY6_0;
	wire w_dff_B_woz0rSSW2_0;
	wire w_dff_B_am17GXv75_0;
	wire w_dff_B_lGxr1js75_0;
	wire w_dff_B_Zzk3xV260_0;
	wire w_dff_B_5iecDHWU5_0;
	wire w_dff_B_BLQN1P1U3_0;
	wire w_dff_B_8vJb4fPa7_0;
	wire w_dff_B_GyZEmpwB0_0;
	wire w_dff_B_XiO6N5Wh8_0;
	wire w_dff_B_UQtWAT099_0;
	wire w_dff_B_ZgwDnQ3j1_0;
	wire w_dff_B_8xEtBd4k8_0;
	wire w_dff_B_6uvlk9mH3_0;
	wire w_dff_B_8rIhmINw8_0;
	wire w_dff_B_6r4cWHNH7_0;
	wire w_dff_B_xSUxJVYv1_1;
	wire w_dff_B_YHtyzqau1_0;
	wire w_dff_B_ddEVRQ7Q7_0;
	wire w_dff_B_3zoO6mt01_0;
	wire w_dff_B_6WTVwIh96_0;
	wire w_dff_B_yVv8qJii1_0;
	wire w_dff_B_EFp0z5Qb6_0;
	wire w_dff_B_2R0WsyJF7_0;
	wire w_dff_B_IsbI2Fv12_0;
	wire w_dff_B_p139BhB06_0;
	wire w_dff_B_0msDaU7S8_0;
	wire w_dff_B_gmGWpgta5_0;
	wire w_dff_B_viTl6LRz7_0;
	wire w_dff_A_3F4ytKjn2_1;
	wire w_dff_A_7X6XhEQy8_1;
	wire w_dff_B_v3w7Yg228_2;
	wire w_dff_B_275f0nXt2_2;
	wire w_dff_B_7L91uwTL8_1;
	wire w_dff_B_YhXlXGjR9_0;
	wire w_dff_B_qXD20aTC1_0;
	wire w_dff_B_nJR4TUuY1_1;
	wire w_dff_B_OTU63Woc9_1;
	wire w_dff_B_0RTIB2M20_1;
	wire w_dff_B_4JaqEF1c5_1;
	wire w_dff_B_lIiPeFPn9_1;
	wire w_dff_B_vPH0PPW99_1;
	wire w_dff_B_oib0qwZT8_1;
	wire w_dff_B_qAQ9g4tO3_1;
	wire w_dff_B_aMA0gFRn7_1;
	wire w_dff_B_EfcMgCN70_1;
	wire w_dff_B_Xga7WSDe7_1;
	wire w_dff_B_MYBZoQKU8_1;
	wire w_dff_B_4FzlR2na7_1;
	wire w_dff_B_XlJT3dCH2_1;
	wire w_dff_B_VreLHDTh9_1;
	wire w_dff_B_swXRbEuM8_1;
	wire w_dff_B_x6SqzwPE6_1;
	wire w_dff_B_iH2R0TEF9_1;
	wire w_dff_B_qSUeiPR88_1;
	wire w_dff_B_E3buoyro4_1;
	wire w_dff_B_jOlsJFD18_1;
	wire w_dff_B_MSqVh61v9_1;
	wire w_dff_B_zYBwZ9ov3_1;
	wire w_dff_B_7yE3ZTQq0_0;
	wire w_dff_B_qDjqAWub7_0;
	wire w_dff_B_dFQcz4hf7_1;
	wire w_dff_A_axV8nzVZ2_1;
	wire w_dff_A_ZB9CuM7a7_1;
	wire w_dff_B_jlaeAtZl5_0;
	wire w_dff_B_QQ5iB8JH2_1;
	wire w_dff_B_EU3V5uT80_1;
	wire w_dff_B_5XShQJNG7_1;
	wire w_dff_B_ohfCSEmq4_1;
	wire w_dff_B_vJ7uPold1_1;
	wire w_dff_B_7nmmNPuO6_1;
	wire w_dff_B_3wfFTdZH3_1;
	wire w_dff_B_IBcbFj835_1;
	wire w_dff_B_jA950uW67_1;
	wire w_dff_B_neeRJMWu1_1;
	wire w_dff_B_jB6Qb3vE6_1;
	wire w_dff_B_MyC8Sz9c4_1;
	wire w_dff_B_skgu4IkI5_1;
	wire w_dff_B_1dbtavxL3_1;
	wire w_dff_B_wFuoGVLd6_1;
	wire w_dff_B_ge0Jm1SX5_1;
	wire w_dff_B_KSktY4Mr6_1;
	wire w_dff_B_giFrDIQ60_1;
	wire w_dff_B_JpAbbAiP6_1;
	wire w_dff_B_qN8Zq43O3_1;
	wire w_dff_A_i9VBFY5u4_0;
	wire w_dff_A_ScFWRy543_0;
	wire w_dff_A_wN0MeD2T1_0;
	wire w_dff_A_tyCRgCWs0_0;
	wire w_dff_A_fzE37sTl9_0;
	wire w_dff_A_diJK79s32_0;
	wire w_dff_A_ZRBmkMcL9_0;
	wire w_dff_A_Qe1V0Qmd0_0;
	wire w_dff_A_br9i2ZRP9_0;
	wire w_dff_A_ZKZiG02d1_0;
	wire w_dff_A_IETcTTfq4_0;
	wire w_dff_A_c72uh5Dh5_0;
	wire w_dff_A_fpkJl5oY0_0;
	wire w_dff_A_UC608D3n8_0;
	wire w_dff_A_1OGrNmsG1_0;
	wire w_dff_A_sjn0rE7i7_0;
	wire w_dff_A_419wEkZg0_0;
	wire w_dff_A_SNPNU4NY5_0;
	wire w_dff_A_unXJm4cd3_1;
	wire w_dff_A_zPvoXHja7_1;
	wire w_dff_A_AfvXZFmK6_1;
	wire w_dff_A_tg6YtNyX5_1;
	wire w_dff_A_75T7SG8l5_1;
	wire w_dff_A_51XrHNuY4_1;
	wire w_dff_A_XswJi0N46_1;
	wire w_dff_A_vtVyJxbu1_1;
	wire w_dff_A_kzuXZDQ53_1;
	wire w_dff_A_0eHIxcLM5_1;
	wire w_dff_A_dF4gTrH22_1;
	wire w_dff_A_yFkfepWh6_1;
	wire w_dff_A_l2EdIA8Y0_1;
	wire w_dff_A_vI6arzXl0_1;
	wire w_dff_A_Tj62m3oB8_1;
	wire w_dff_A_BYOx4pAQ6_1;
	wire w_dff_A_Kt8qZ9wz2_1;
	wire w_dff_A_ZHLQcGmu8_1;
	wire w_dff_A_FkbKZ3nL0_1;
	wire w_dff_A_QNhc1giV7_0;
	wire w_dff_A_1tqHPfDU0_0;
	wire w_dff_B_WGEwa6yO8_1;
	wire w_dff_B_DKx92Ewv1_0;
	wire w_dff_B_8Xg2FRhN2_0;
	wire w_dff_B_dPVwk9Ay5_0;
	wire w_dff_B_Jdb6f3iR3_0;
	wire w_dff_B_3UuxGaOS6_0;
	wire w_dff_B_I4JpWT8j1_0;
	wire w_dff_B_DGak4m8X4_0;
	wire w_dff_B_LxJvPTEC3_0;
	wire w_dff_B_bYYFb0U43_0;
	wire w_dff_B_tApKYSbX2_0;
	wire w_dff_B_oV0HxQMx7_0;
	wire w_dff_B_nFMmOQw68_0;
	wire w_dff_B_PVquzBYK4_1;
	wire w_dff_B_AVSF0Oxw8_1;
	wire w_dff_B_PTsd3AOl7_1;
	wire w_dff_B_xdVHyrCp1_1;
	wire w_dff_B_ijlws6n16_1;
	wire w_dff_B_B3dkUnZH3_1;
	wire w_dff_B_o4aZeyj90_0;
	wire w_dff_B_QZFZsH7S2_0;
	wire w_dff_B_2wW6iHNC3_0;
	wire w_dff_B_2bFDFdJQ3_0;
	wire w_dff_B_iLJQh0yV3_0;
	wire w_dff_B_pbZN7arC8_0;
	wire w_dff_B_ppXrUYdm2_0;
	wire w_dff_B_4zeUQeoC6_1;
	wire w_dff_B_qZohO1Mp1_0;
	wire w_dff_B_OqWtzlI70_0;
	wire w_dff_B_26Vy7vBT7_0;
	wire w_dff_B_2bfFMkNo0_0;
	wire w_dff_B_7MFYz6Q68_0;
	wire w_dff_B_RXABdTP05_1;
	wire w_dff_B_mjJCM2hf6_0;
	wire w_dff_B_Yh40dTcU2_1;
	wire w_dff_B_yb49y52C9_1;
	wire w_dff_B_jYnSfBdI6_1;
	wire w_dff_B_DJYD2Cpt1_0;
	wire w_dff_B_lo148zU95_1;
	wire w_dff_B_jbbSM2MA9_1;
	wire w_dff_B_rSzU9W9K9_1;
	wire w_dff_B_4JQUvYtX3_1;
	wire w_dff_B_V4onKTSI5_1;
	wire w_dff_B_2BA9YJBT0_0;
	wire w_dff_B_WLizeP4z7_0;
	wire w_dff_B_hQWB1MV24_0;
	wire w_dff_B_B7rMKbCp5_0;
	wire w_dff_B_F73aXzK84_1;
	wire w_dff_B_dmMFLBrb2_1;
	wire w_dff_B_IhGxUNJH0_1;
	wire w_dff_A_CzaUIjUg2_1;
	wire w_dff_A_RBGIcHEi1_1;
	wire w_dff_B_u0fVKxXR3_0;
	wire w_dff_B_gT5iOp9K8_1;
	wire w_dff_B_3LIk1Ekd7_1;
	wire w_dff_B_dtN22ksm2_1;
	wire w_dff_B_1kq4zCQq3_1;
	wire w_dff_B_b5Osdyfb3_1;
	wire w_dff_B_dSbXADPr8_1;
	wire w_dff_A_IdP4ctH51_1;
	wire w_dff_A_sYh46rC06_1;
	wire w_dff_A_2huqbXvQ3_1;
	wire w_dff_B_c3brB32t2_0;
	wire w_dff_B_HRJ2qjEE6_0;
	wire w_dff_B_1MxHLlVx4_0;
	wire w_dff_B_Roa0scio0_0;
	wire w_dff_A_oSt1N62k5_0;
	wire w_dff_A_4T6D0jPq0_1;
	wire w_dff_B_IrkBxSno6_0;
	wire w_dff_B_b0bU9vGe5_0;
	wire w_dff_B_EeVSRKdi1_0;
	wire w_dff_B_Oxd3EAzS3_0;
	wire w_dff_B_legx5ooM3_0;
	wire w_dff_B_l47fYpKe0_1;
	wire w_dff_B_u0QRMWvq1_1;
	wire w_dff_B_Fhq7c8ss2_0;
	wire w_dff_B_RTO9is4E1_0;
	wire w_dff_B_Bj8BiRrI3_1;
	wire w_dff_B_4HVNIoJw8_1;
	wire w_dff_B_bGx2WRnA7_1;
	wire w_dff_B_rJw8V6fi8_0;
	wire w_dff_B_kikptGj60_1;
	wire w_dff_B_T6FbOtID0_1;
	wire w_dff_B_LdT9P7kQ6_1;
	wire w_dff_B_wvhPnYKL8_0;
	wire w_dff_B_NmoD7dCD2_2;
	wire w_dff_B_e0kCTptf6_2;
	wire w_dff_B_3NFxnZsM7_2;
	wire w_dff_A_nMX3tB6p1_1;
	wire w_dff_A_jYgrIUsq7_1;
	wire w_dff_A_fcW30N6G1_1;
	wire w_dff_A_7sA1ggSy2_1;
	wire w_dff_A_LqppROXH2_1;
	wire w_dff_B_crVwk4RA1_0;
	wire w_dff_A_kcaawKiK3_0;
	wire w_dff_B_TCA5IC1A5_0;
	wire w_dff_B_RWqRYJSi4_0;
	wire w_dff_B_eQDmSvRQ5_0;
	wire w_dff_B_SyaITMJG9_0;
	wire w_dff_B_LI2DMJ7g8_0;
	wire w_dff_A_SbYlVY0u7_2;
	wire w_dff_A_M88EWdos2_2;
	wire w_dff_A_pdmCXQak7_2;
	wire w_dff_B_8JH86pGa9_0;
	wire w_dff_B_RDYtqR090_0;
	wire w_dff_B_MtfLmKbi8_1;
	wire w_dff_B_I5WQYAhc1_1;
	wire w_dff_B_6LfJIXbT7_0;
	wire w_dff_B_J4fxFNtS0_1;
	wire w_dff_B_JWLVUhxx3_0;
	wire w_dff_B_0EyZIcUc8_0;
	wire w_dff_B_K3IeCsJk6_0;
	wire w_dff_B_xeCC2MJU7_0;
	wire w_dff_B_et0EBgT21_1;
	wire w_dff_B_EeBQm7hU3_1;
	wire w_dff_B_CsuIWoK75_0;
	wire w_dff_A_7AcN7zvh3_2;
	wire w_dff_B_DU2XGEIQ6_2;
	wire w_dff_B_tZTxkOmW8_1;
	wire w_dff_B_QTK8jM607_1;
	wire w_dff_B_bBjhKhHV1_1;
	wire w_dff_B_t7y68eUg3_0;
	wire w_dff_A_5a2f4HA13_0;
	wire w_dff_A_xcnpLyZY2_1;
	wire w_dff_A_LTTgHIkk4_1;
	wire w_dff_A_h0TQx0tk1_1;
	wire w_dff_A_PdBQPsih0_1;
	wire w_dff_A_PA0pLMAL5_2;
	wire w_dff_A_TuMdgiC28_2;
	wire w_dff_A_swxpps9B3_2;
	wire w_dff_B_yW3zibOM5_0;
	wire w_dff_B_NKahejBj1_1;
	wire w_dff_B_u811M5jM0_1;
	wire w_dff_B_V6mBJiHs9_0;
	wire w_dff_B_OGdqf51U6_0;
	wire w_dff_A_BNcqOQnr9_0;
	wire w_dff_A_37fG59s46_0;
	wire w_dff_A_Cu0d6UVD6_0;
	wire w_dff_A_LJEiiwrx0_0;
	wire w_dff_A_Rmpq5NyL1_1;
	wire w_dff_A_ma6Qyv6a7_1;
	wire w_dff_A_99HJibvw4_1;
	wire w_dff_B_MtzuOHMI5_0;
	wire w_dff_A_HeEO2Nmd3_1;
	wire w_dff_A_y3dUgMXB2_1;
	wire w_dff_B_rv7l7Nhd4_1;
	wire w_dff_B_VmrBYFvk2_1;
	wire w_dff_B_DJ7CFo3m2_0;
	wire w_dff_B_xo4Jgk4M3_0;
	wire w_dff_B_BUE8W33A7_0;
	wire w_dff_B_OPcy1Z589_1;
	wire w_dff_B_FGtXuGGF7_1;
	wire w_dff_B_1J4G0RQ80_1;
	wire w_dff_B_0L24BZH86_1;
	wire w_dff_A_WDPW7eG30_1;
	wire w_dff_A_70LQrWZs1_1;
	wire w_dff_B_q6WBqKV42_0;
	wire w_dff_B_khDDenXF7_0;
	wire w_dff_B_K9CLbvgv0_0;
	wire w_dff_B_XoM5BIMh5_3;
	wire w_dff_B_hFsXgRLs2_1;
	wire w_dff_B_ZwcaPGGG5_1;
	wire w_dff_B_JanaiJrn9_0;
	wire w_dff_B_CipYhRss3_0;
	wire w_dff_B_kbCxJTKh5_0;
	wire w_dff_B_oAeiECGu0_0;
	wire w_dff_B_786NVzyQ2_0;
	wire w_dff_B_2Etd3YNq0_0;
	wire w_dff_B_yS816wcL4_1;
	wire w_dff_B_VKqW2bGp3_0;
	wire w_dff_A_AZhXc43T4_0;
	wire w_dff_B_DhQRgtAm4_1;
	wire w_dff_B_ZUSVDj2j0_1;
	wire w_dff_B_qPT0ujuH2_1;
	wire w_dff_B_DwVnuUP80_1;
	wire w_dff_B_WJZSQhCj2_1;
	wire w_dff_B_k9MMBBPr6_1;
	wire w_dff_B_bs5p4BPX4_0;
	wire w_dff_B_hlJjD9Rg6_0;
	wire w_dff_B_5S32BAId0_1;
	wire w_dff_B_V844WwYT9_1;
	wire w_dff_B_MvjyWkCQ5_1;
	wire w_dff_B_BG6W7Crp7_1;
	wire w_dff_B_krmUV8RO2_1;
	wire w_dff_B_KQKiFyKL2_1;
	wire w_dff_B_xVasj5kJ8_1;
	wire w_dff_B_jy15bCAb1_1;
	wire w_dff_B_epMcabcQ1_0;
	wire w_dff_A_G37cgPAn4_2;
	wire w_dff_B_wqUxesZM3_0;
	wire w_dff_B_9d9RryJv7_0;
	wire w_dff_B_YRi0c8Xj3_0;
	wire w_dff_B_oYg0olwJ0_1;
	wire w_dff_B_pxdSli3m3_1;
	wire w_dff_B_iDRMvkcQ1_1;
	wire w_dff_B_1Cq0U0a39_1;
	wire w_dff_B_c5054Njd6_1;
	wire w_dff_B_8VZ402Ky1_1;
	wire w_dff_B_PrT57hO05_1;
	wire w_dff_B_vHxeNTmt0_1;
	wire w_dff_A_HdEUKy3C7_1;
	wire w_dff_A_Yxo3N9Dl4_1;
	wire w_dff_B_QmBhjrpP1_1;
	wire w_dff_B_5KLB4HMo4_1;
	wire w_dff_B_Ve7dusDi5_1;
	wire w_dff_B_8NAA6ogq4_1;
	wire w_dff_A_GMDgsM5t5_0;
	wire w_dff_A_JhtiTWaw7_1;
	wire w_dff_A_eKFFuyiO9_1;
	wire w_dff_A_skVO2sRG1_1;
	wire w_dff_A_GAnDltAD0_2;
	wire w_dff_A_Cr9tn0ke9_2;
	wire w_dff_A_9GBNWQMK3_2;
	wire w_dff_A_9nNLVVbJ4_2;
	wire w_dff_B_QA35yFD00_0;
	wire w_dff_A_3acfUPkO1_0;
	wire w_dff_A_vVDfAQXi7_0;
	wire w_dff_A_Jrn4DL1P6_2;
	wire w_dff_A_tLivtiAV8_2;
	wire w_dff_B_hU0nysu46_0;
	wire w_dff_B_rQOiTh2F7_0;
	wire w_dff_A_c9wDqvvY5_1;
	wire w_dff_A_j3wkjTyJ9_2;
	wire w_dff_A_weg0WuY85_1;
	wire w_dff_A_D9DjRBCi5_2;
	wire w_dff_B_p66zbhX35_1;
	wire w_dff_B_ViLt7ylH0_0;
	wire w_dff_A_SzkP9lAQ1_0;
	wire w_dff_A_xZZrXenR4_1;
	wire w_dff_B_CU5aFT977_1;
	wire w_dff_B_Yvw3WQHh8_0;
	wire w_dff_A_Tiy1oMGB9_0;
	wire w_dff_A_6g9wIwMo1_0;
	wire w_dff_A_7F7lXBco6_0;
	wire w_dff_A_JO8zr94B0_0;
	wire w_dff_A_kHIp0HDB7_0;
	wire w_dff_A_UEPnqtJ47_0;
	wire w_dff_A_t2jFqypB4_1;
	wire w_dff_A_Ba2yrQhG0_1;
	wire w_dff_B_2PCwmbBR7_0;
	wire w_dff_B_Zx7LqFSw7_0;
	wire w_dff_B_FaljJk7V4_0;
	wire w_dff_B_vHDgTMOi9_2;
	wire w_dff_A_TdTjlMHl0_0;
	wire w_dff_A_8WxTUa831_0;
	wire w_dff_B_THST2BMr9_0;
	wire w_dff_B_GTezD0Qw4_0;
	wire w_dff_B_YDTS5TL70_1;
	wire w_dff_B_nb4eicKF1_1;
	wire w_dff_B_kDfzSqZk9_1;
	wire w_dff_B_Ivzg3xIC2_2;
	wire w_dff_B_qFYVwUnH9_1;
	wire w_dff_B_46XW8r5J1_0;
	wire w_dff_A_YLbAZ4IE3_1;
	wire w_dff_A_RtHqXjHw8_1;
	wire w_dff_A_RTF9YcsN6_2;
	wire w_dff_A_88dtetgu2_2;
	wire w_dff_B_fbIPnkxY0_1;
	wire w_dff_B_HZzZqG3p2_1;
	wire w_dff_B_mvi4auYb9_1;
	wire w_dff_B_zwFczmjs6_1;
	wire w_dff_B_Xa2q3nUo6_1;
	wire w_dff_B_1qY5Qug65_1;
	wire w_dff_B_czY4iSWw4_1;
	wire w_dff_B_ZfTKSLIY4_1;
	wire w_dff_B_JjmVLEll5_0;
	wire w_dff_B_cY4O8HI96_1;
	wire w_dff_B_FpeKF35t2_0;
	wire w_dff_B_3wSKf3w46_1;
	wire w_dff_B_dI0eegyn0_0;
	wire w_dff_B_Ol7dW2sh1_3;
	wire w_dff_B_W5QdNekh4_3;
	wire w_dff_B_fFWHIJFq9_3;
	wire w_dff_B_xE9yzJRL6_2;
	wire w_dff_B_m5lLCWo20_2;
	wire w_dff_B_sAp9YiIm4_2;
	wire w_dff_B_89NlwPhh7_0;
	wire w_dff_B_l8LxeCNm6_1;
	wire w_dff_B_gKYk9sFL5_1;
	wire w_dff_B_kjHWZixp2_1;
	wire w_dff_A_xtKFON032_1;
	wire w_dff_A_5KU2o8vn6_1;
	wire w_dff_A_EI2Ilcku7_1;
	wire w_dff_A_MVA5MfC56_2;
	wire w_dff_B_Nf5ZYQsw4_0;
	wire w_dff_B_I8HULOXn1_3;
	wire w_dff_B_fUDQcBrn4_3;
	wire w_dff_B_ug54TCuZ7_3;
	wire w_dff_A_oNML8KrU4_1;
	wire w_dff_A_fkGtClK13_1;
	wire w_dff_A_7zgZhvPP8_1;
	wire w_dff_A_bZ7ijSYX5_1;
	wire w_dff_A_NOiZkSxo8_1;
	wire w_dff_A_IjIfmfFq0_1;
	wire w_dff_A_vnEzpc403_1;
	wire w_dff_A_IXYedGQu8_0;
	wire w_dff_A_XXccezFo3_0;
	wire w_dff_A_mOWTb5FC6_0;
	wire w_dff_A_TZMEC8n68_0;
	wire w_dff_A_SBZocElh5_0;
	wire w_dff_A_4EQ5NfpF9_0;
	wire w_dff_A_A6BCbUAz9_0;
	wire w_dff_A_XVppy1kU6_0;
	wire w_dff_A_Sdz9dIll5_0;
	wire w_dff_A_kpzSiGhz9_2;
	wire w_dff_A_L6gHmMgr3_2;
	wire w_dff_A_jYOdfjyW0_2;
	wire w_dff_A_A3JHM3JR6_2;
	wire w_dff_A_375oD3Ou8_2;
	wire w_dff_A_rvfB9a4U4_2;
	wire w_dff_A_ohTChJrT1_2;
	wire w_dff_A_TgRKKufT2_1;
	wire w_dff_A_WaUW4dsG2_1;
	wire w_dff_A_2ZcylJBQ1_1;
	wire w_dff_A_WXyYF0iP0_1;
	wire w_dff_A_TeFbGmaE3_1;
	wire w_dff_A_jWwQZyvX9_1;
	wire w_dff_A_dICPL2Kz8_1;
	wire w_dff_A_kZcMbeTU7_2;
	wire w_dff_A_weYYilAH6_2;
	wire w_dff_A_6M9fzjsc1_2;
	wire w_dff_A_5iYGyZjj1_2;
	wire w_dff_A_2S75jRV98_2;
	wire w_dff_A_0PsnEPoP3_2;
	wire w_dff_A_9x6Qr2Io4_2;
	wire w_dff_B_VudIogzL6_0;
	wire w_dff_B_aQjpBnWG0_0;
	wire w_dff_B_elJ768Fw9_0;
	wire w_dff_B_o9wqmrq05_0;
	wire w_dff_B_xVPcu1ND6_2;
	wire w_dff_B_41Caj17Y1_2;
	wire w_dff_B_LjJcccF96_2;
	wire w_dff_B_GzgNPC5e4_2;
	wire w_dff_B_fW9xPb2b1_2;
	wire w_dff_B_s6fuivb63_2;
	wire w_dff_B_EOIIpEcT9_2;
	wire w_dff_B_QnSeoWhd6_2;
	wire w_dff_B_YLlFhacG2_2;
	wire w_dff_B_ZYb40iFp0_0;
	wire w_dff_B_h4RtadRs5_0;
	wire w_dff_B_b1pGu6vw9_0;
	wire w_dff_B_nGgjxvac3_0;
	wire w_dff_B_QsZcq38y8_0;
	wire w_dff_B_K6EzFokF1_0;
	wire w_dff_B_b4TGWIg46_0;
	wire w_dff_B_0KBgtigG8_1;
	wire w_dff_B_SAV4Uvhx7_1;
	wire w_dff_B_7jyzD58J2_0;
	wire w_dff_B_eRCI9hCc9_0;
	wire w_dff_B_0E64AsKd0_1;
	wire w_dff_B_uRqsTUXW5_1;
	wire w_dff_A_kiZ2YnPA2_1;
	wire w_dff_A_o4LQQvKM3_2;
	wire w_dff_A_SNqBWfVJ2_1;
	wire w_dff_A_iJUgBwq71_1;
	wire w_dff_A_7p48mYnV6_1;
	wire w_dff_A_hPLRTLOf3_1;
	wire w_dff_A_WVhOwAHD2_2;
	wire w_dff_A_z6SlBdM10_2;
	wire w_dff_A_OWA3kIlo0_2;
	wire w_dff_A_59ogoqPM0_2;
	wire w_dff_A_b5r1Lzgn7_0;
	wire w_dff_A_UT8H2Vic3_0;
	wire w_dff_A_Wbs76ppA6_0;
	wire w_dff_A_8hHkL1PG3_2;
	wire w_dff_A_CSZbFV0d2_2;
	wire w_dff_A_eoz6teQ20_2;
	wire w_dff_B_DktmHrQx5_0;
	wire w_dff_B_sOcuBiPH3_1;
	wire w_dff_B_Q1qvxK2L3_1;
	wire w_dff_B_IdjcOSiq5_0;
	wire w_dff_A_jy5KOk1X7_1;
	wire w_dff_A_H7I5RNYx4_2;
	wire w_dff_B_AS6caYQk9_3;
	wire w_dff_B_iav8vIDC0_3;
	wire w_dff_B_k4zStVQl6_3;
	wire w_dff_B_bC9jIfkQ7_0;
	wire w_dff_A_RufEhbVX7_0;
	wire w_dff_A_oTtkGiLK7_0;
	wire w_dff_A_Mwr1h53n1_1;
	wire w_dff_A_X7KaqByy2_1;
	wire w_dff_A_8Zb4vVrW1_1;
	wire w_dff_A_QCOAP4Qk2_1;
	wire w_dff_B_gY9f2nnX4_0;
	wire w_dff_A_4Oz5YSYp3_1;
	wire w_dff_A_zob0P3cI5_2;
	wire w_dff_B_gbC0DPc77_1;
	wire w_dff_A_85GgCVqu2_1;
	wire w_dff_A_eAk7lmmX5_1;
	wire w_dff_A_zbujm7Tb4_2;
	wire w_dff_A_IBJkRmJa1_2;
	wire w_dff_A_DPRKpDgj8_2;
	wire w_dff_B_gqoWoSKU3_0;
	wire w_dff_B_0ZIerqGo2_0;
	wire w_dff_B_yJpCBKoX8_0;
	wire w_dff_B_CKoaYjSd0_0;
	wire w_dff_A_MKuYlg0D3_0;
	wire w_dff_A_vvO22FOj2_1;
	wire w_dff_A_sWmskyep9_1;
	wire w_dff_A_daKAvAwE4_1;
	wire w_dff_B_keav1kmT0_0;
	wire w_dff_B_dqgSnqHA1_0;
	wire w_dff_B_3fZRx6RI2_0;
	wire w_dff_B_FImqC54b9_0;
	wire w_dff_B_JCQfpg1X7_0;
	wire w_dff_A_rWWVvxsJ8_0;
	wire w_dff_A_k3JGA4C40_0;
	wire w_dff_A_EeZjSg887_2;
	wire w_dff_A_4NmqG9wv9_2;
	wire w_dff_B_pVqq1Jlu5_1;
	wire w_dff_B_t0VQJmnK4_2;
	wire w_dff_A_VTeMM7ch9_0;
	wire w_dff_B_qU8NM3Dz0_3;
	wire w_dff_B_nrXDqPfL0_3;
	wire w_dff_B_c69DTJYd0_3;
	wire w_dff_A_7AYaMK7Q9_1;
	wire w_dff_A_nYsWf3yJ0_1;
	wire w_dff_A_oAWWLL5M1_1;
	wire w_dff_B_t6Zcu4g47_0;
	wire w_dff_A_1LTuX2rb6_1;
	wire w_dff_B_TtNazLUZ4_2;
	wire w_dff_B_Klqcwm7I2_2;
	wire w_dff_B_E2pzOZt54_1;
	wire w_dff_B_k6F7bK6c4_0;
	wire w_dff_B_5R6QWDEa2_0;
	wire w_dff_A_8yy2zotn6_0;
	wire w_dff_A_Ntvkszga7_0;
	wire w_dff_A_JFkCUEOJ0_0;
	wire w_dff_A_95QQxCPE3_1;
	wire w_dff_B_CB45gDrB0_1;
	wire w_dff_B_EmiIeIdo0_1;
	wire w_dff_B_vYoGX6kR4_0;
	wire w_dff_B_15Lwp3E76_0;
	wire w_dff_B_KhwKB54G4_0;
	wire w_dff_B_FtEUyvTn6_0;
	wire w_dff_B_h0wBLRfa5_1;
	wire w_dff_B_aC3Hupml5_1;
	wire w_dff_B_5hryCipb2_1;
	wire w_dff_B_S3vy7CbM2_1;
	wire w_dff_B_g84FQDWf9_1;
	wire w_dff_B_kcBHfiiB6_1;
	wire w_dff_A_KqevKNcd0_0;
	wire w_dff_A_fGoUnq7h8_1;
	wire w_dff_B_FuPue6fb6_1;
	wire w_dff_B_S22Biev41_1;
	wire w_dff_B_BszKyM8a9_1;
	wire w_dff_B_TgVEMjNG0_0;
	wire w_dff_B_C3Zh2WT72_0;
	wire w_dff_B_9Fy2kyov4_0;
	wire w_dff_B_f1dpro7X6_0;
	wire w_dff_B_eUERuVKn4_0;
	wire w_dff_B_pmKtcmWA5_0;
	wire w_dff_A_0RGvImsv3_1;
	wire w_dff_A_JJ9RWBLE3_1;
	wire w_dff_A_yJJP5N8H3_2;
	wire w_dff_A_4Fk1I7i19_2;
	wire w_dff_A_uQxop5AO8_2;
	wire w_dff_B_PDdmklrm3_1;
	wire w_dff_B_HLS7OORf1_1;
	wire w_dff_A_oye51Lho7_0;
	wire w_dff_B_YFNG28sK1_2;
	wire w_dff_A_zymzxxtQ7_1;
	wire w_dff_A_65LzyoxR2_1;
	wire w_dff_A_ptzGm7K20_1;
	wire w_dff_B_nDVKlNPf1_2;
	wire w_dff_B_El1Kyins8_2;
	wire w_dff_B_EQkryD4M1_1;
	wire w_dff_B_pWjzjc0O5_1;
	wire w_dff_B_Tvnatg297_1;
	wire w_dff_B_DwUkk4SC4_1;
	wire w_dff_B_Nvo7ve6m3_0;
	wire w_dff_A_20GyYu6S9_2;
	wire w_dff_B_RecgrcfT2_1;
	wire w_dff_B_INQMja0C0_1;
	wire w_dff_B_LIelNfwt4_1;
	wire w_dff_B_04N51c2S8_1;
	wire w_dff_B_vha6vETx4_1;
	wire w_dff_A_74Wh4UtW0_1;
	wire w_dff_A_rIxLrDBm1_1;
	wire w_dff_A_t7kP4Kj38_1;
	wire w_dff_A_1XGtQpBl9_2;
	wire w_dff_A_GjChyxxK5_2;
	wire w_dff_A_nj2QBwlE1_2;
	wire w_dff_A_gov1gbCz0_1;
	wire w_dff_A_hqL2N1gy3_1;
	wire w_dff_A_b7CJdTKD3_1;
	wire w_dff_A_nQKuoKeb7_2;
	wire w_dff_A_zQKuk2nr8_2;
	wire w_dff_A_kd5ECbCg6_0;
	wire w_dff_A_LiCi63DK0_0;
	wire w_dff_A_VnmzGIqZ9_2;
	wire w_dff_A_qP0PjycH7_2;
	wire w_dff_A_qcAqNnII1_2;
	wire w_dff_A_R2ndmZqm6_2;
	wire w_dff_A_0BjMtfxy1_1;
	wire w_dff_A_XRyOIwwU7_1;
	wire w_dff_A_zBQyaB0w2_1;
	wire w_dff_A_jW3dfybX5_0;
	wire w_dff_A_ldFcLSv06_0;
	wire w_dff_A_ps1pBBQg0_0;
	wire w_dff_A_NlNqZx0B9_2;
	wire w_dff_A_NpK6idSS1_2;
	wire w_dff_A_cDRNt68D6_2;
	wire w_dff_A_bhT07Qpo8_2;
	wire w_dff_A_6b4CzQnG1_0;
	wire w_dff_A_95tQa7W18_0;
	wire w_dff_A_eed2vNmR3_0;
	wire w_dff_B_PYzOnq4l7_0;
	wire w_dff_B_UFkzWYqI2_0;
	wire w_dff_B_g093PoJh8_0;
	wire w_dff_B_k4AlFgau3_0;
	wire w_dff_B_5JxwEWcx5_0;
	wire w_dff_B_XuRRvTNa2_0;
	wire w_dff_A_1UvET2Be9_2;
	wire w_dff_A_efUUGvLH3_2;
	wire w_dff_A_zYsdWECT7_2;
	wire w_dff_A_XTfzI8En2_0;
	wire w_dff_A_EHw4u9ai4_0;
	wire w_dff_B_VEDtvJyM9_1;
	wire w_dff_B_52MHcjgq9_1;
	wire w_dff_B_h4Y4CTa98_1;
	wire w_dff_B_YUqIbko90_1;
	wire w_dff_B_2tEorJjR7_1;
	wire w_dff_B_qy7Dk0eB1_1;
	wire w_dff_B_3P2caIMQ0_1;
	wire w_dff_B_S29NIsBY5_0;
	wire w_dff_B_nCwovcnt8_1;
	wire w_dff_B_Zrtp0TWN6_0;
	wire w_dff_A_Ec9Kqgjw8_0;
	wire w_dff_A_8kX5hHrJ2_0;
	wire w_dff_A_QW2IITbk9_0;
	wire w_dff_A_Ul9C7h3E4_0;
	wire w_dff_A_nTi7pOJZ7_2;
	wire w_dff_A_aVf2RN5x9_2;
	wire w_dff_A_BIlKLNuA7_2;
	wire w_dff_A_KLAYTlk53_2;
	wire w_dff_B_DQhw4aS97_1;
	wire w_dff_B_5ccDlyQl1_0;
	wire w_dff_B_KDY4NsUX0_3;
	wire w_dff_B_pMMLIfB61_3;
	wire w_dff_B_p5xIi9sp7_3;
	wire w_dff_B_86WmmvN65_1;
	wire w_dff_B_MdgUWO5j9_1;
	wire w_dff_A_13t7fpQR2_1;
	wire w_dff_A_JhIdS5Fe6_1;
	wire w_dff_A_wLrENlk49_1;
	wire w_dff_A_VoSx3bgd5_2;
	wire w_dff_A_i2IVPP7p7_2;
	wire w_dff_B_x6nOYpLm4_3;
	wire w_dff_B_8WysDD1G7_3;
	wire w_dff_B_PhCYIDkf7_3;
	wire w_dff_B_JVT5tKHq1_3;
	wire w_dff_B_4B88tn5x2_3;
	wire w_dff_B_t5fzPJDL5_3;
	wire w_dff_A_Ct00FSky8_0;
	wire w_dff_A_d7nwO7Jr9_1;
	wire w_dff_A_XSqLkxZc8_0;
	wire w_dff_A_Sb91akbp9_0;
	wire w_dff_A_7A7o9IQa1_1;
	wire w_dff_B_1kwtdeLX0_3;
	wire w_dff_B_GuEHFn4Z5_3;
	wire w_dff_A_uKnjDzBp6_1;
	wire w_dff_A_Ey0AHIns3_1;
	wire w_dff_A_fCkOyNJy8_2;
	wire w_dff_A_sNGWQ4tz3_2;
	wire w_dff_A_lSokXZRf2_0;
	wire w_dff_A_1Wr1bQN09_0;
	wire w_dff_A_0BzWVpQx9_0;
	wire w_dff_A_TjKxMyW99_2;
	wire w_dff_A_2MWFxzgl8_2;
	wire w_dff_A_SZ6fREAm2_2;
	wire w_dff_A_sRnO9raa1_2;
	wire w_dff_A_lQFdV4Wy1_1;
	wire w_dff_A_ZRrFFLui7_1;
	wire w_dff_A_7itG0YhZ9_1;
	wire w_dff_A_FduOWoSV4_0;
	wire w_dff_A_RswzhSnl3_0;
	wire w_dff_A_xXtWINz73_0;
	wire w_dff_A_RvgJFnRR0_0;
	wire w_dff_A_914Uzl4u8_1;
	wire w_dff_A_3m2KYaT92_1;
	wire w_dff_A_OFynWe806_1;
	wire w_dff_A_UiCAF1gL4_1;
	wire w_dff_A_HlyjsgJx5_1;
	wire w_dff_B_zPIqeoSO7_1;
	wire w_dff_B_iNLtdpIO2_0;
	wire w_dff_A_lmYTnB6T2_0;
	wire w_dff_A_rvbd5L818_0;
	wire w_dff_A_G446uEg82_0;
	wire w_dff_A_o1fgSDMH9_0;
	wire w_dff_A_arW3GOKm9_0;
	wire w_dff_A_7JjrxqHK3_0;
	wire w_dff_A_NecxCShL5_1;
	wire w_dff_A_qn3EYT6o2_1;
	wire w_dff_A_3O7aE85M4_1;
	wire w_dff_A_odEjqQBT9_0;
	wire w_dff_A_tbzMfHWv2_1;
	wire w_dff_A_Y8KSfdHb2_1;
	wire w_dff_A_DU6dpN675_1;
	wire w_dff_A_LYezivm14_1;
	wire w_dff_A_6fc83rfr5_1;
	wire w_dff_A_DvtEd7gf6_1;
	wire w_dff_A_OZ9A1o2l5_1;
	wire w_dff_A_gPvOOn0B3_2;
	wire w_dff_A_DvFUx4YH1_2;
	wire w_dff_A_pB0AHT919_2;
	wire w_dff_A_fGxofY8k0_2;
	wire w_dff_A_8XGHsvdi4_0;
	wire w_dff_A_bKzLMaed4_1;
	wire w_dff_A_dSGJppjg1_1;
	wire w_dff_B_mc5XNW0i3_3;
	wire w_dff_B_p5r3z6Ka3_3;
	wire w_dff_B_YQvH26gl2_3;
	wire w_dff_A_gRoTD7iz4_0;
	wire w_dff_A_fuzE1ysw1_0;
	wire w_dff_A_3d4Cb9cl2_0;
	wire w_dff_A_5MLe7set8_0;
	wire w_dff_A_hVtkSxNU2_0;
	wire w_dff_A_JWLUa8kc1_0;
	wire w_dff_A_yT7VtqIj3_0;
	wire w_dff_A_XgI3rQ976_0;
	wire w_dff_A_c3PGxlbs7_2;
	wire w_dff_A_XPAo245d2_2;
	wire w_dff_A_RmERhBON2_2;
	wire w_dff_A_UvJVFXnw5_2;
	wire w_dff_A_SM7ZPe7K2_2;
	wire w_dff_A_7pMbHm3V3_2;
	wire w_dff_A_X3wMX2hI4_2;
	wire w_dff_A_tcO6s0D57_2;
	wire w_dff_A_d3EBu8i75_1;
	wire w_dff_A_ceDSiX433_1;
	wire w_dff_A_Wj35XI293_1;
	wire w_dff_A_NQgcz3gX4_1;
	wire w_dff_A_seuHrhMy5_2;
	wire w_dff_A_nuaJKMkK5_1;
	wire w_dff_A_MGRcmzfo9_1;
	wire w_dff_A_lqWvE3r74_1;
	wire w_dff_A_iuagizU15_2;
	wire w_dff_A_UOXfvX1p2_2;
	wire w_dff_A_5HJK33pc5_2;
	wire w_dff_A_B8iF0AOI6_0;
	wire w_dff_A_EXPJgVUo8_0;
	wire w_dff_A_hVTreHXn7_0;
	wire w_dff_A_MosWL2Xc7_0;
	wire w_dff_A_6hzNH7Wq9_0;
	wire w_dff_A_kSHJvLUk9_0;
	wire w_dff_A_XvKL8ZfZ2_0;
	wire w_dff_A_9denz4cd7_0;
	wire w_dff_A_4lLPtiA58_0;
	wire w_dff_A_oB09sLbt1_0;
	wire w_dff_A_RaQ0g0xZ2_1;
	wire w_dff_A_ITfKXpn52_1;
	wire w_dff_A_UOpVM55s0_1;
	wire w_dff_A_gOcQMJAL3_1;
	wire w_dff_A_XEUCRZjE9_1;
	wire w_dff_A_8bgwqSiU6_1;
	wire w_dff_A_tc432UJX6_1;
	wire w_dff_A_9eOwMtlQ2_1;
	wire w_dff_A_tIIMMgaG3_1;
	wire w_dff_A_3Nq7jofV2_1;
	wire w_dff_A_vvGvnuOX4_1;
	wire w_dff_A_ohqUtohD0_1;
	wire w_dff_A_iXigC0zp9_1;
	wire w_dff_A_OYlcoSK01_1;
	wire w_dff_A_gEXTiP6o9_1;
	wire w_dff_A_Tl9ag5Oa2_1;
	wire w_dff_A_dtYZgtNk1_1;
	wire w_dff_A_0wOEUyzd3_1;
	wire w_dff_A_JyqdRTrX8_2;
	wire w_dff_A_DojwvyJK9_2;
	wire w_dff_A_67hGSlyt0_2;
	wire w_dff_A_dEjDbPbD9_2;
	wire w_dff_A_oBRutj0d7_2;
	wire w_dff_A_E18gzmfh6_2;
	wire w_dff_A_nS6ihTCi8_2;
	wire w_dff_A_AQJ35VO30_2;
	wire w_dff_A_YTQDqmI01_2;
	wire w_dff_A_GSDAVnE79_2;
	wire w_dff_A_aaUwg8TN3_2;
	wire w_dff_A_Q4uINlbI6_0;
	wire w_dff_A_LLkLYzzG5_0;
	wire w_dff_A_jULG3NAn2_0;
	wire w_dff_A_gMO5Afgd7_1;
	wire w_dff_A_DMtX3I347_1;
	wire w_dff_B_8Fgn1vPH7_0;
	wire w_dff_B_JiVUAAap8_0;
	wire w_dff_A_ZhSqkV059_0;
	wire w_dff_A_6ULOEFua4_0;
	wire w_dff_A_kLIzZhGG6_2;
	wire w_dff_A_AWmVjZRn3_2;
	wire w_dff_A_Afyz80ea3_2;
	wire w_dff_A_2E3IIK0F1_2;
	wire w_dff_A_KGHKFH5d7_2;
	wire w_dff_A_AY9jNJeF9_2;
	wire w_dff_A_eMkn6guf5_2;
	wire w_dff_A_dLX1RnmY5_0;
	wire w_dff_A_OWnSuGej0_0;
	wire w_dff_A_WWHFDgjM6_0;
	wire w_dff_A_C4dNcQlP8_0;
	wire w_dff_A_y12OfxT53_0;
	wire w_dff_A_FYYhgysf1_0;
	wire w_dff_A_g1RxLjhU4_0;
	wire w_dff_A_KaDu34l84_0;
	wire w_dff_A_psX1F1CX9_0;
	wire w_dff_A_XuQLkVNX5_0;
	wire w_dff_A_RKaGtSos7_0;
	wire w_dff_A_k3fbjoaD1_0;
	wire w_dff_A_xQzqKOOf3_0;
	wire w_dff_A_99KqSkib8_0;
	wire w_dff_A_qQ98sBdi6_2;
	wire w_dff_A_W8fROgog4_2;
	wire w_dff_A_g62GXDFM2_2;
	wire w_dff_A_1QtS2Hu31_2;
	wire w_dff_A_evb7rlOY0_2;
	wire w_dff_A_qjpiyGia4_2;
	wire w_dff_A_fOTowXgS5_2;
	wire w_dff_A_xlz6eex52_2;
	wire w_dff_A_qo6zb8tr9_2;
	wire w_dff_A_fx8vizA06_2;
	wire w_dff_B_ZJlqJ5FK5_3;
	wire w_dff_A_T2KnlB2j0_0;
	wire w_dff_A_oWD7Fbko3_0;
	wire w_dff_A_jJo4eJM59_0;
	wire w_dff_A_8U1wUBmo4_0;
	wire w_dff_A_jOSOqfwz8_0;
	wire w_dff_A_AWYJwKgI1_0;
	wire w_dff_A_TSmGjlnZ7_0;
	wire w_dff_A_yrkL9nfY4_0;
	wire w_dff_A_enbsVRWP4_0;
	wire w_dff_A_ouEGlPzD1_0;
	wire w_dff_A_uP2pN1Iw3_0;
	wire w_dff_A_BbfphW8d0_0;
	wire w_dff_A_mYqX3KMD9_0;
	wire w_dff_A_k48sJ4dU4_0;
	wire w_dff_A_0tAfQwI36_0;
	wire w_dff_A_qAo7eWBD2_0;
	wire w_dff_A_lh9QJT3N1_0;
	wire w_dff_A_2D7mIetl1_0;
	wire w_dff_A_Cb3BKH502_0;
	wire w_dff_A_sWvLeDdt9_0;
	wire w_dff_A_Dx84Df5y9_0;
	wire w_dff_A_gdygnVVT6_0;
	wire w_dff_A_hZGV57du9_2;
	wire w_dff_A_zZlJKFXg8_2;
	wire w_dff_A_JcRZ1cNk5_2;
	wire w_dff_A_7aY8PRMZ7_2;
	wire w_dff_A_T6m0G33s8_2;
	wire w_dff_A_TvD462gv0_2;
	wire w_dff_A_N8DzoCir9_2;
	wire w_dff_A_knLSeDn77_2;
	wire w_dff_A_uxs6nHfu0_2;
	wire w_dff_A_qkiXRVFc3_2;
	wire w_dff_A_3eXUnVcQ9_2;
	wire w_dff_A_kcce7wmu0_2;
	wire w_dff_A_mLrwQRJ09_1;
	wire w_dff_A_n5CXs36m9_1;
	wire w_dff_A_pnnxiLey6_1;
	wire w_dff_A_l1y7ttSN8_1;
	wire w_dff_A_ue9GOMuM9_1;
	wire w_dff_A_BaZBveCO0_1;
	wire w_dff_A_CYmuDsfL2_1;
	wire w_dff_A_egzqFENt9_1;
	wire w_dff_A_VXkfY5sT6_1;
	wire w_dff_A_yHY3JlNx6_1;
	wire w_dff_A_DHUjSQ1X3_1;
	wire w_dff_A_N4EYChmd7_2;
	wire w_dff_A_UrMqEtit8_2;
	wire w_dff_A_DdkSMVhT9_2;
	wire w_dff_A_ufzJQTfW8_2;
	wire w_dff_A_aKrx2RoP6_2;
	wire w_dff_A_hqp1s0XK0_2;
	wire w_dff_A_ThhlVpCb8_2;
	wire w_dff_A_8dOLieCe3_2;
	wire w_dff_A_lVqvmdGJ6_2;
	wire w_dff_A_we57jcH39_2;
	wire w_dff_A_A4hFy3VS9_2;
	wire w_dff_B_lVDmVpR90_1;
	wire w_dff_A_FjTBNcjL8_0;
	wire w_dff_A_9ralKSB82_0;
	wire w_dff_A_JALV2n893_2;
	wire w_dff_A_zYqiFtf66_2;
	wire w_dff_A_G8ZFd4Pm3_1;
	wire w_dff_A_Osu92vvW7_1;
	wire w_dff_B_Vkewf4pA1_0;
	wire w_dff_A_tibR6DAP5_1;
	wire w_dff_B_1kLZs6DX8_2;
	wire w_dff_B_cGtmdP1h3_2;
	wire w_dff_B_eElI0crC8_2;
	wire w_dff_B_qDaUGw3r8_0;
	wire w_dff_B_DYgSAR3B4_0;
	wire w_dff_B_218vRI5f9_0;
	wire w_dff_A_dSJwJBTY2_1;
	wire w_dff_A_qkw04i6F0_1;
	wire w_dff_A_J25dw3vL9_1;
	wire w_dff_A_MCUi8aXw4_2;
	wire w_dff_B_Sph0DQDc9_0;
	wire w_dff_A_cSstGaA84_1;
	wire w_dff_B_i1l3Mp175_0;
	wire w_dff_A_y6gSzsOt4_1;
	wire w_dff_A_7G2esgGD7_1;
	wire w_dff_A_KNB7jK4F8_1;
	wire w_dff_A_PnyFohuo6_2;
	wire w_dff_A_bUhcjxrq5_2;
	wire w_dff_B_D9Bk1MgI6_1;
	wire w_dff_B_vEpVHQhZ6_0;
	wire w_dff_A_kIrJMqOC9_0;
	wire w_dff_A_IlnhALf97_0;
	wire w_dff_A_CgQNpzjX4_1;
	wire w_dff_A_XNG8O2VN2_1;
	wire w_dff_A_oirhwcSF6_0;
	wire w_dff_A_cFfobJ8r5_2;
	wire w_dff_A_kv1ybzLQ2_2;
	wire w_dff_A_CIvU00uO4_2;
	wire w_dff_A_K12y90Dv4_2;
	wire w_dff_A_Jefdi59f3_1;
	wire w_dff_A_q9GcptK94_2;
	wire w_dff_A_vbKRF6U80_2;
	wire w_dff_A_LtOaC5ti7_2;
	wire w_dff_A_KFtuu9GJ7_1;
	wire w_dff_A_JSzHfLnD1_2;
	wire w_dff_A_ExMXZJ148_2;
	wire w_dff_A_ZnOsSdK38_0;
	wire w_dff_B_sTdKnjCs0_2;
	wire w_dff_A_G4hzl8R49_0;
	wire w_dff_A_a2K9M8PJ6_0;
	wire w_dff_A_SxnUIRhj3_0;
	wire w_dff_A_QGVfY15l5_0;
	wire w_dff_A_jbHEXkL91_1;
	wire w_dff_A_jWc4I7cD0_1;
	wire w_dff_A_9oEPz5k67_1;
	wire w_dff_A_udX6hQZn4_1;
	wire w_dff_A_21OGRLrO6_1;
	wire w_dff_A_o5lDOTfG0_1;
	wire w_dff_A_cPCngAaW3_0;
	wire w_dff_A_kSMsUd1o0_0;
	wire w_dff_A_iZGzzApM4_1;
	wire w_dff_A_fUYKTDQV8_1;
	wire w_dff_A_GBs9BNAo1_1;
	wire w_dff_A_mI5bW7u41_1;
	wire w_dff_A_ogkQdYD97_2;
	wire w_dff_A_fVvvUUjm7_2;
	wire w_dff_A_jytAgkMy8_1;
	wire w_dff_B_ZsnwmpzD2_0;
	wire w_dff_B_eFv68KBx7_0;
	wire w_dff_A_ENbhoJix7_2;
	wire w_dff_B_UtzkZXLy9_1;
	wire w_dff_B_UDv9v5b98_2;
	wire w_dff_B_c57VbaU79_0;
	wire w_dff_B_Mc9vSWlq9_0;
	wire w_dff_B_bJzwrDL81_1;
	wire w_dff_B_0Br3Y3Xv2_0;
	wire w_dff_A_8E9uyBLA2_1;
	wire w_dff_B_pK93kYGq3_1;
	wire w_dff_A_ZB48YLv05_2;
	wire w_dff_B_DgFaPa4o1_0;
	wire w_dff_B_zDwXkz7L6_0;
	wire w_dff_B_xJhhQOrv7_0;
	wire w_dff_B_IymNsGxt3_1;
	wire w_dff_A_OouquvDn0_1;
	wire w_dff_A_lNlDI1Rb2_1;
	wire w_dff_A_a28Q80VO5_2;
	wire w_dff_A_HEqpfb7G1_2;
	wire w_dff_A_6qkdxHfH4_2;
	wire w_dff_A_mqvqmVgS5_2;
	wire w_dff_A_yVpbMnEO9_2;
	wire w_dff_A_5Fr6r7e69_2;
	wire w_dff_A_gymKLIgf9_0;
	wire w_dff_A_FMppqw4O3_0;
	wire w_dff_A_loB4VqjS4_2;
	wire w_dff_A_GIbWYEPv0_2;
	wire w_dff_A_Gm6slROH2_0;
	wire w_dff_A_CXN2s6KH5_0;
	wire w_dff_A_bmpJ6iiq1_0;
	wire w_dff_A_YcOfHab10_0;
	wire w_dff_A_zdtf3Fyo1_0;
	wire w_dff_A_KdM2oFPR6_0;
	wire w_dff_A_srhLiocW2_0;
	wire w_dff_A_axAXm0vz6_0;
	wire w_dff_A_4SImS4Oy6_0;
	wire w_dff_A_stwUmo9O5_0;
	wire w_dff_A_HfFi8Oi51_0;
	wire w_dff_A_QKFIK7XV4_0;
	wire w_dff_A_lcp8cHKR3_0;
	wire w_dff_A_k928IC5l2_0;
	wire w_dff_A_avztiM3w5_0;
	wire w_dff_A_W0Tp6BaR2_0;
	wire w_dff_A_NZPioaXJ2_0;
	wire w_dff_A_vPczuf2F2_1;
	wire w_dff_A_qRayeMKr2_0;
	wire w_dff_A_Qmrw5kIL7_2;
	wire w_dff_A_iv2p9UGR7_2;
	wire w_dff_A_YaTQG0RH8_2;
	wire w_dff_A_r3TYdPRz8_1;
	wire w_dff_A_HHT873W73_1;
	wire w_dff_A_TupEKacE0_1;
	wire w_dff_A_7cFzR9Dh8_1;
	wire w_dff_A_tQVBHVvz7_1;
	wire w_dff_A_P3wnx4oD8_1;
	wire w_dff_A_lQLBJZEQ1_2;
	wire w_dff_A_vSxQjJ4X3_2;
	wire w_dff_A_qMrvZvq50_2;
	wire w_dff_A_hX56HpIG0_2;
	wire w_dff_A_UfVmVae33_2;
	wire w_dff_A_ploXWUQo9_0;
	wire w_dff_A_ojWxuxiD0_2;
	wire w_dff_A_zrSwBRGm1_0;
	wire w_dff_A_MANApDwJ0_0;
	wire w_dff_A_cFPEjfVC8_1;
	wire w_dff_A_l7lSQxMl7_1;
	wire w_dff_A_juWXiyw33_1;
	wire w_dff_A_bq9azBta7_1;
	wire w_dff_A_QSNq6Oc96_1;
	wire w_dff_A_pgCw6MNt0_1;
	wire w_dff_A_ogwZrAhS2_1;
	wire w_dff_A_k8fhh1kp1_1;
	wire w_dff_A_0CemE09k5_1;
	wire w_dff_A_QUMlrFU18_1;
	wire w_dff_A_WdJmdwBX6_1;
	wire w_dff_A_f9zbZg4C8_1;
	wire w_dff_A_2wRSdLNF4_1;
	wire w_dff_A_9bWExnt25_1;
	wire w_dff_A_aLEHXo812_1;
	wire w_dff_B_wirumzpe5_0;
	wire w_dff_B_IzQrH9399_2;
	wire w_dff_B_8fOJpo850_1;
	wire w_dff_A_oLRdNPdw6_2;
	wire w_dff_A_nP6h92hb4_1;
	wire w_dff_A_t0iXcEPt3_2;
	wire w_dff_B_qA13Ndc32_0;
	wire w_dff_B_yTEEUpH48_0;
	wire w_dff_B_fc3BiEcZ2_0;
	wire w_dff_B_zYYggNLe3_0;
	wire w_dff_B_nh7xxYWg9_1;
	wire w_dff_B_L6FeC3JP5_1;
	wire w_dff_B_i14Gol6C4_1;
	wire w_dff_A_0NDHMjEF6_0;
	wire w_dff_A_g7sa2qLA6_0;
	wire w_dff_A_9ZQvLSfa8_0;
	wire w_dff_A_hjgbbSVR8_0;
	wire w_dff_A_LKMSibzd4_0;
	wire w_dff_A_uqeqgqm72_0;
	wire w_dff_A_zT5VIxUQ5_0;
	wire w_dff_A_nYiQUxpz5_0;
	wire w_dff_A_OtV27sqM7_0;
	wire w_dff_A_8gxL498K9_1;
	wire w_dff_A_X8ZBCkA41_1;
	wire w_dff_A_As1zAiFl1_1;
	wire w_dff_B_WgAINPb89_1;
	wire w_dff_B_wewM4ZSQ5_1;
	wire w_dff_A_l8rs1oAb6_0;
	wire w_dff_A_ybYp2lXE1_1;
	wire w_dff_B_w4Awezhr4_0;
	wire w_dff_B_BzP9mOHK2_1;
	wire w_dff_A_NaxlSU6n5_1;
	wire w_dff_A_ifeXtB8u5_1;
	wire w_dff_A_2J23iolI4_1;
	wire w_dff_A_izkfXpqB4_1;
	wire w_dff_A_Rda2fYaU8_2;
	wire w_dff_A_ZFm3XZBk4_2;
	wire w_dff_A_HK9oBtJF2_2;
	wire w_dff_A_XEEFmGT81_2;
	wire w_dff_A_y8Uk3cet7_2;
	wire w_dff_A_t5wxuhce7_1;
	wire w_dff_B_jwuRkkXK5_0;
	wire w_dff_B_zO1IRGag5_1;
	wire w_dff_B_eta8Muoc4_1;
	wire w_dff_B_lrDaUowg2_0;
	wire w_dff_A_8G0arO6g1_1;
	wire w_dff_A_pGVeTZBk0_0;
	wire w_dff_A_FDiH7MW27_0;
	wire w_dff_B_FO8Gwv0J1_1;
	wire w_dff_B_K7z4jg7I0_1;
	wire w_dff_B_NBjz2sFV6_0;
	wire w_dff_A_4386Ygz54_1;
	wire w_dff_A_i99ftJfc5_1;
	wire w_dff_A_beC0eKaG7_1;
	wire w_dff_A_ONukrniH5_1;
	wire w_dff_A_AsGZYBOs7_2;
	wire w_dff_A_2FUbW2rT0_2;
	wire w_dff_B_prqkqRTk6_0;
	wire w_dff_B_N3cNAHsT0_0;
	wire w_dff_A_8TdrWGBZ9_1;
	wire w_dff_A_rvC2vt7T8_0;
	wire w_dff_A_9ZunfM6Y5_2;
	wire w_dff_B_lw8HqzXo4_1;
	wire w_dff_B_I8qsIiur3_1;
	wire w_dff_A_GQxHmHkp4_0;
	wire w_dff_A_CCEoeB2a5_2;
	wire w_dff_A_hcTSn3R21_2;
	wire w_dff_A_XqgdXkng9_2;
	wire w_dff_A_FrLgA80Y5_0;
	wire w_dff_A_hxr1AAEs1_1;
	wire w_dff_A_BiQXPWQW1_1;
	wire w_dff_A_BJu1r9gt1_2;
	wire w_dff_A_97bTYVVD3_0;
	wire w_dff_A_0HiOQMRJ8_0;
	wire w_dff_A_O2VcMFTg2_0;
	wire w_dff_A_6QVyZ4HI3_1;
	wire w_dff_A_Kw9nV4ns7_1;
	wire w_dff_A_RZwJTBHH0_1;
	wire w_dff_B_l1NMarM66_0;
	wire w_dff_A_CQRgG1Mw5_0;
	wire w_dff_A_uShzZ3Uv1_0;
	wire w_dff_A_al7IYk3V8_1;
	wire w_dff_A_WnxFzNr57_1;
	wire w_dff_A_PDL6C3nK3_0;
	wire w_dff_A_GmVYZNx38_0;
	wire w_dff_A_6SZHnbiP5_0;
	wire w_dff_A_UQq57QqN0_1;
	wire w_dff_A_GawpsW3m4_1;
	wire w_dff_A_g7WmM91Q2_1;
	wire w_dff_A_n2oDV0SI8_1;
	wire w_dff_A_b9bC12Y00_0;
	wire w_dff_A_UYQbUqrz6_0;
	wire w_dff_A_O00dREir7_0;
	wire w_dff_A_iniuKwvB2_2;
	wire w_dff_A_biPj3nGp6_2;
	wire w_dff_A_nzLoglhV6_2;
	wire w_dff_A_W8LYVIsw3_1;
	wire w_dff_A_YBHsC95D4_1;
	wire w_dff_A_axinjCBL2_2;
	wire w_dff_A_j7dOrHzR6_2;
	wire w_dff_A_TH2JGvDg9_1;
	wire w_dff_B_zBzpHhf81_0;
	wire w_dff_B_OaAB421S6_1;
	wire w_dff_A_TuWqKq408_1;
	wire w_dff_A_OHCadVq27_2;
	wire w_dff_A_cYYAdWbW6_0;
	wire w_dff_A_RovLMnhq5_2;
	wire w_dff_A_b7wLZy7l7_0;
	wire w_dff_B_GHq7vOay5_2;
	wire w_dff_A_cTwrrY2b4_0;
	wire w_dff_A_tIMCN33B9_0;
	wire w_dff_A_JgdntH6e3_0;
	wire w_dff_A_e9A7km2s9_0;
	wire w_dff_A_Fou26Hox4_0;
	wire w_dff_A_tZAQhP2l8_1;
	wire w_dff_B_7U7WpZzl4_1;
	wire w_dff_B_JIOC8EHz8_1;
	wire w_dff_A_mU3DqGOy2_0;
	wire w_dff_A_b6fZpL3E6_0;
	wire w_dff_B_I5nmTvxU4_0;
	wire w_dff_A_JeMaVs6t4_0;
	wire w_dff_A_h9DR7GMP4_2;
	wire w_dff_A_8CzCP1zt1_2;
	wire w_dff_A_rsQJNHKW4_2;
	wire w_dff_A_8sWGGBbl3_2;
	wire w_dff_A_EWkT1AOP3_0;
	wire w_dff_B_PT24TNez2_2;
	wire w_dff_A_rcOOxg1z3_0;
	wire w_dff_A_mbURjbvu7_0;
	wire w_dff_A_ygo3ADFz2_0;
	wire w_dff_A_tIDm05Cz1_0;
	wire w_dff_B_xIKDQVJe5_0;
	wire w_dff_B_crRIzxv97_0;
	wire w_dff_B_HZzECxmh4_2;
	wire w_dff_A_HYmMZDFV0_0;
	wire w_dff_A_PwEDttqh4_0;
	wire w_dff_A_94KTuCpr8_0;
	wire w_dff_A_ydIkuUtG6_0;
	wire w_dff_A_cZljE8hi0_1;
	wire w_dff_A_SgbIM5EI2_1;
	wire w_dff_A_Ny0Ff4VQ5_1;
	wire w_dff_A_1vvZxFoU0_2;
	wire w_dff_A_eo3IM3vo2_2;
	wire w_dff_B_lS3T56Se1_3;
	wire w_dff_A_xhAvvTf95_1;
	wire w_dff_B_cKunexlm0_1;
	wire w_dff_B_9COU33x02_1;
	wire w_dff_B_GhdvqHhs9_0;
	wire w_dff_A_xMCwb3Xo0_0;
	wire w_dff_A_cTRfOIBm7_1;
	wire w_dff_A_ugZr37UL0_1;
	wire w_dff_A_4JO5gZAH2_0;
	wire w_dff_A_k8oJfmuI6_0;
	wire w_dff_A_2JC8ADef4_0;
	wire w_dff_A_8tLQ4KOD3_1;
	wire w_dff_A_jmu46CmJ4_1;
	wire w_dff_A_wiJr0S7S8_1;
	wire w_dff_A_QADLD1h01_1;
	wire w_dff_A_icbPBZjK5_0;
	wire w_dff_A_muro9qR59_0;
	wire w_dff_A_9J0G4DIm3_0;
	wire w_dff_A_jqGbUiad9_1;
	wire w_dff_A_7KaqsGwY4_1;
	wire w_dff_A_HY0WJrlP2_1;
	wire w_dff_A_PO9MuSmM7_2;
	wire w_dff_A_44PSQTCf1_2;
	wire w_dff_A_NdF95UbF0_2;
	wire w_dff_A_2Y721u017_0;
	wire w_dff_B_hFHsXgb73_0;
	wire w_dff_B_GRlG9TWL1_0;
	wire w_dff_B_q0dCNmqv6_0;
	wire w_dff_A_Li4Jjbkf8_0;
	wire w_dff_A_v9EzSQWy9_0;
	wire w_dff_A_sVsvKSQR7_0;
	wire w_dff_A_Cxmm5ts75_0;
	wire w_dff_A_dmI39b8w6_1;
	wire w_dff_A_t54hNTpi6_2;
	wire w_dff_A_pxALCa0e1_2;
	wire w_dff_A_Jyv2PZ9J5_2;
	wire w_dff_A_UviIzfNq3_2;
	wire w_dff_A_DFkFYigY0_0;
	wire w_dff_A_4kDaLvsJ5_0;
	wire w_dff_A_BfNynjZ25_0;
	wire w_dff_A_FpJre54a5_0;
	wire w_dff_A_RUd1jwHC1_0;
	wire w_dff_A_ti81mePK8_1;
	wire w_dff_A_C3y9u9Zz6_1;
	wire w_dff_A_1dXG9ppK9_1;
	wire w_dff_A_4d3ZXjKD6_1;
	wire w_dff_B_xmYl4AbE2_1;
	wire w_dff_B_bFExBmbu0_1;
	wire w_dff_B_1cfpiNrB1_0;
	wire w_dff_B_xzZaUamp2_0;
	wire w_dff_B_EGl2WplV9_2;
	wire w_dff_B_tQ5bBQum0_1;
	wire w_dff_B_PrZaD5Zv0_1;
	wire w_dff_B_5wPozv1I6_1;
	wire w_dff_B_ZoCsYINS5_3;
	wire w_dff_A_y5rIwcE93_2;
	wire w_dff_A_siocPJva6_0;
	wire w_dff_A_UxntVVz47_2;
	wire w_dff_A_N10FqqUo3_0;
	wire w_dff_B_FIeyk8Fz8_3;
	wire w_dff_B_9FwPhw8Q1_3;
	wire w_dff_B_l4X8PHtZ6_3;
	wire w_dff_A_AvaVEbvT4_0;
	wire w_dff_A_hKWWXyq27_0;
	wire w_dff_A_ctNigOQu5_0;
	wire w_dff_A_Fc5aWhdd9_0;
	wire w_dff_A_BJplSB7a7_1;
	wire w_dff_A_o8gycTsf9_1;
	wire w_dff_A_CmiBshCD6_1;
	wire w_dff_A_OimBSSv70_1;
	wire w_dff_A_1AsNcgwk6_0;
	wire w_dff_A_XHYTYbR15_0;
	wire w_dff_A_BROATec47_0;
	wire w_dff_A_53Uc2rbS7_0;
	wire w_dff_B_BM9YOQ0C2_1;
	wire w_dff_B_cL8Xs4078_1;
	wire w_dff_B_aCcUphpJ2_0;
	wire w_dff_B_j2zTilF61_0;
	wire w_dff_B_opaONvPE0_0;
	wire w_dff_A_m6CFZT0t9_1;
	wire w_dff_A_gHqlsMsW1_1;
	wire w_dff_A_uXhuoCTd3_1;
	wire w_dff_A_ss9i5BgQ2_2;
	wire w_dff_A_0p1AtjHg8_0;
	wire w_dff_A_nCQ6NDQn7_0;
	wire w_dff_A_hVNnjKgP6_2;
	wire w_dff_A_RCUi5Vvx2_2;
	wire w_dff_A_mKrXYaZq8_2;
	wire w_dff_A_kzFWYfB52_0;
	wire w_dff_A_86qZ2guA2_1;
	wire w_dff_B_DVVSq78l4_1;
	wire w_dff_A_AiFPZa8C2_1;
	wire w_dff_A_xb1N1XZD3_1;
	wire w_dff_A_nQ70BLCU2_1;
	wire w_dff_A_LXJDY3TB2_2;
	wire w_dff_A_8UVLIIqI1_2;
	wire w_dff_A_e7fhqZWt8_2;
	wire w_dff_A_4Koz7mTc1_2;
	wire w_dff_A_rGidlNBb4_2;
	wire w_dff_A_ucjKX2Ip8_2;
	wire w_dff_A_XOGi0qq44_1;
	wire w_dff_A_7DvbtkSk3_1;
	wire w_dff_A_uVI7mBqD7_1;
	wire w_dff_A_kef2gZQk4_2;
	wire w_dff_A_osY162wu3_2;
	wire w_dff_A_dGUtwM5M9_2;
	wire w_dff_A_e3ybj4k98_0;
	wire w_dff_A_G6UuLri30_0;
	wire w_dff_A_yzUpWH5M6_0;
	wire w_dff_A_4u2Un4vU5_1;
	wire w_dff_A_yqm5Cmbs8_0;
	wire w_dff_A_6pRkK9FN2_0;
	wire w_dff_A_ukR2nlQi9_2;
	wire w_dff_A_tKUtTOmO6_2;
	wire w_dff_A_mWHgdEQc4_2;
	wire w_dff_A_vg2Y6Sze3_0;
	wire w_dff_A_uCTlBNek9_0;
	wire w_dff_A_FvwJAaIG2_0;
	wire w_dff_A_zaqVxPXS5_0;
	wire w_dff_A_yoPHyq905_2;
	wire w_dff_A_0m7SaP7A3_2;
	wire w_dff_A_ayIycAJM7_1;
	wire w_dff_A_Dfp0TMCR9_1;
	wire w_dff_A_234SJcZS8_1;
	wire w_dff_A_3Xzilur23_2;
	wire w_dff_A_5FpVGYKY5_2;
	wire w_dff_A_zmKQObbx5_2;
	wire w_dff_A_afzTHK3A5_2;
	wire w_dff_A_56JqZ5B84_1;
	wire w_dff_A_QT5SPFcM2_0;
	wire w_dff_A_CO2XZcYU0_0;
	wire w_dff_A_O8zT6EuW1_2;
	wire w_dff_A_z8K8SKsH1_2;
	wire w_dff_A_hNy8bXX81_2;
	wire w_dff_A_4WU1ylqH1_2;
	wire w_dff_A_bLHzeMOq5_2;
	wire w_dff_A_ssqYW7xV1_0;
	wire w_dff_A_gWXHEB4g6_2;
	wire w_dff_A_mzOzAUZf7_0;
	wire w_dff_A_ttZt2BHE1_0;
	wire w_dff_B_CJBybfjs7_2;
	wire w_dff_A_HLumzEHt0_0;
	wire w_dff_A_Bni4SiGC5_0;
	wire w_dff_A_dznUlpk64_0;
	wire w_dff_A_tCWyG7hq5_2;
	wire w_dff_A_qHGWqIUO4_2;
	wire w_dff_A_qMdiEpKU1_2;
	wire w_dff_A_criETge50_2;
	wire w_dff_A_5YazrCLb8_1;
	wire w_dff_A_fn6533Kk3_1;
	wire w_dff_A_GPRLNY7X4_1;
	wire w_dff_A_C1VcRIZQ0_2;
	wire w_dff_A_krMXfSYv2_0;
	wire w_dff_A_YsH3D4I38_1;
	wire w_dff_A_UWPcFigi2_0;
	wire w_dff_B_EVEz00gg4_0;
	wire w_dff_A_rZ2wUsBs6_0;
	wire w_dff_A_HiU1UimC1_2;
	wire w_dff_A_U5o5NzoL2_0;
	wire w_dff_A_q5Q5q2co5_0;
	wire w_dff_A_a5XfqDH46_0;
	wire w_dff_A_h2y9xBoJ6_0;
	wire w_dff_A_5b4c8wso7_1;
	wire w_dff_A_j7mMMThK7_1;
	wire w_dff_A_wFga1qG85_0;
	wire w_dff_A_OLPawTs87_2;
	wire w_dff_A_q7dzlngA8_2;
	wire w_dff_A_3cucR8oQ9_2;
	wire w_dff_A_0wn3i1iz8_0;
	wire w_dff_A_TY2VhRBY5_0;
	wire w_dff_A_S7dmdcD61_1;
	wire w_dff_A_2kdKdgmT8_1;
	wire w_dff_A_0bxmfvZ33_1;
	wire w_dff_A_npIB8IR04_1;
	wire w_dff_A_F27IqvPM3_2;
	wire w_dff_A_9sBnGlXU2_2;
	wire w_dff_A_DJiarWZ95_2;
	wire w_dff_A_lJhY60M69_0;
	wire w_dff_A_J0qcyDa95_0;
	wire w_dff_A_cQ5cFH192_1;
	wire w_dff_A_2UtXVpAi1_1;
	wire w_dff_A_LmlS4BSt7_0;
	wire w_dff_A_Xnnkyn8u5_2;
	wire w_dff_A_WEIuYqWf0_2;
	wire w_dff_A_puhH3F2G7_1;
	wire w_dff_A_1XfGqOOE2_1;
	wire w_dff_A_1JXlQGbO6_1;
	wire w_dff_A_L9B71FRG1_2;
	wire w_dff_A_VIHtJ1nh8_2;
	wire w_dff_A_uiWlur9c6_2;
	wire w_dff_A_1YvdgI3Y2_1;
	wire w_dff_A_MjRQy9tV0_1;
	wire w_dff_A_W9EB8iqA1_1;
	wire w_dff_A_RRQhBpxU0_2;
	wire w_dff_A_92PNDuK20_0;
	wire w_dff_A_Yqz3Gn3v8_0;
	wire w_dff_A_fJLa1NaZ1_1;
	wire w_dff_A_G6UpWjIo9_1;
	wire w_dff_A_i6QxGQVe1_1;
	wire w_dff_A_2v78RoHI8_2;
	wire w_dff_A_FsqTWjI07_2;
	wire w_dff_A_InfOy5b73_2;
	wire w_dff_A_PrLHja963_0;
	wire w_dff_A_tC83FC8o7_0;
	wire w_dff_A_qkXshSGn7_1;
	wire w_dff_A_JGhT6wNK3_1;
	wire w_dff_A_SEmmsmwT0_1;
	wire w_dff_A_b5uT6m1p0_2;
	wire w_dff_A_h8ARcq9S8_2;
	wire w_dff_A_Vmigz4lE8_1;
	wire w_dff_A_iqj7eGhw3_2;
	wire w_dff_A_ChjD05Oz7_1;
	wire w_dff_A_klL2CcSO6_2;
	wire w_dff_A_2ThYXdQ06_1;
	wire w_dff_A_tOq02BT72_2;
	wire w_dff_A_Ofo02QnI0_0;
	wire w_dff_A_8EkU4qhP9_1;
	wire w_dff_A_XDkJrU828_2;
	wire w_dff_A_d8SxFKtX6_2;
	wire w_dff_A_glmJoVXE4_2;
	wire w_dff_A_11ZkU7Ow7_2;
	wire w_dff_A_OJmdWQiM5_2;
	wire w_dff_A_dPMt59dE4_0;
	wire w_dff_A_gjlubog67_1;
	wire w_dff_A_2PjEZTO05_1;
	wire w_dff_A_0CVfsRU63_2;
	wire w_dff_A_xLxPARyb1_2;
	wire w_dff_A_1hNsEnv72_0;
	wire w_dff_A_zKO6tXtJ2_2;
	wire w_dff_A_4ccyHmp11_0;
	wire w_dff_A_3DuuZRVa7_1;
	wire w_dff_A_gVRr6fTO5_1;
	wire w_dff_A_8OtG8urN5_1;
	wire w_dff_A_ZUfJKdXR1_1;
	wire w_dff_A_BOalHFFR6_2;
	wire w_dff_A_UsWvRPmX7_2;
	wire w_dff_A_IF5vSjQB9_2;
	wire w_dff_A_08fsOT2c1_0;
	wire w_dff_A_dZf0Wm7P0_0;
	wire w_dff_A_93DlXyxW7_0;
	wire w_dff_A_3oN4b9F83_0;
	wire w_dff_A_6uEwpP187_0;
	wire w_dff_A_mDogEzEr3_1;
	wire w_dff_A_gutowc619_1;
	wire w_dff_A_Grg7VoFW1_1;
	wire w_dff_A_sK7Q5PHe8_1;
	wire w_dff_A_2Q8RLOiD5_2;
	wire w_dff_A_TifJx5L45_2;
	wire w_dff_A_xmxtQFrp3_2;
	wire w_dff_A_kv2bcKv06_2;
	wire w_dff_A_H15fiu2u7_2;
	jnot g0000(.din(w_G77_5[1]),.dout(n72),.clk(gclk));
	jnot g0001(.din(w_G50_5[2]),.dout(n73),.clk(gclk));
	jnot g0002(.din(w_G58_5[1]),.dout(n74),.clk(gclk));
	jnot g0003(.din(w_G68_5[1]),.dout(n75),.clk(gclk));
	jand g0004(.dina(w_n75_1[1]),.dinb(w_n74_1[1]),.dout(n76),.clk(gclk));
	jand g0005(.dina(w_n76_0[1]),.dinb(w_n73_2[2]),.dout(n77),.clk(gclk));
	jand g0006(.dina(w_n77_0[1]),.dinb(w_n72_1[1]),.dout(G353),.clk(gclk));
	jnot g0007(.din(w_G97_5[1]),.dout(n79),.clk(gclk));
	jnot g0008(.din(w_G107_5[1]),.dout(n80),.clk(gclk));
	jand g0009(.dina(w_n80_1[1]),.dinb(w_n79_0[2]),.dout(n81),.clk(gclk));
	jnot g0010(.din(w_n81_0[2]),.dout(n82),.clk(gclk));
	jand g0011(.dina(n82),.dinb(w_G87_3[2]),.dout(n83),.clk(gclk));
	jnot g0012(.din(n83),.dout(G355_fa_),.clk(gclk));
	jand g0013(.dina(w_G20_7[1]),.dinb(w_G1_3[1]),.dout(n85),.clk(gclk));
	jnot g0014(.din(w_G226_1[1]),.dout(n86),.clk(gclk));
	jcb g0015(.dina(w_n86_0[1]),.dinb(w_n73_2[1]),.dout(n87));
	jnot g0016(.din(w_G264_1[1]),.dout(n88),.clk(gclk));
	jcb g0017(.dina(w_n88_1[1]),.dinb(w_n80_1[0]),.dout(n89));
	jand g0018(.dina(n89),.dinb(n87),.dout(n90),.clk(gclk));
	jnot g0019(.din(w_G257_1[2]),.dout(n91),.clk(gclk));
	jcb g0020(.dina(w_n91_1[2]),.dinb(w_n79_0[1]),.dout(n92));
	jnot g0021(.din(w_G238_1[2]),.dout(n93),.clk(gclk));
	jcb g0022(.dina(w_n93_0[1]),.dinb(w_n75_1[0]),.dout(n94));
	jand g0023(.dina(n94),.dinb(n92),.dout(n95),.clk(gclk));
	jand g0024(.dina(n95),.dinb(n90),.dout(n96),.clk(gclk));
	jnot g0025(.din(w_G87_3[1]),.dout(n97),.clk(gclk));
	jnot g0026(.din(w_G250_0[2]),.dout(n98),.clk(gclk));
	jcb g0027(.dina(w_n98_2[1]),.dinb(w_n97_2[1]),.dout(n99));
	jnot g0028(.din(w_G232_1[2]),.dout(n100),.clk(gclk));
	jcb g0029(.dina(n100),.dinb(w_n74_1[0]),.dout(n101));
	jand g0030(.dina(n101),.dinb(n99),.dout(n102),.clk(gclk));
	jnot g0031(.din(w_G244_1[2]),.dout(n103),.clk(gclk));
	jcb g0032(.dina(w_n103_0[2]),.dinb(w_n72_1[0]),.dout(n104));
	jnot g0033(.din(w_G116_4[2]),.dout(n105),.clk(gclk));
	jnot g0034(.din(w_G270_0[2]),.dout(n106),.clk(gclk));
	jcb g0035(.dina(w_n106_0[1]),.dinb(w_n105_2[1]),.dout(n107));
	jand g0036(.dina(n107),.dinb(n104),.dout(n108),.clk(gclk));
	jand g0037(.dina(n108),.dinb(n102),.dout(n109),.clk(gclk));
	jand g0038(.dina(n109),.dinb(n96),.dout(n110),.clk(gclk));
	jcb g0039(.dina(n110),.dinb(w_n85_0[2]),.dout(n111));
	jnot g0040(.din(w_G20_7[0]),.dout(n112),.clk(gclk));
	jnot g0041(.din(w_G1_3[0]),.dout(n113),.clk(gclk));
	jnot g0042(.din(w_G13_1[1]),.dout(n114),.clk(gclk));
	jcb g0043(.dina(w_n114_1[2]),.dinb(w_n113_3[1]),.dout(n115));
	jcb g0044(.dina(w_n115_1[1]),.dinb(w_n112_5[2]),.dout(n116));
	jnot g0045(.din(w_n76_0[0]),.dout(n117),.clk(gclk));
	jand g0046(.dina(n117),.dinb(w_G50_5[1]),.dout(n118),.clk(gclk));
	jnot g0047(.din(w_n118_0[2]),.dout(n119),.clk(gclk));
	jcb g0048(.dina(n119),.dinb(w_n116_0[1]),.dout(n120));
	jand g0049(.dina(w_n114_1[1]),.dinb(w_G1_2[2]),.dout(n121),.clk(gclk));
	jand g0050(.dina(w_n121_0[2]),.dinb(w_G20_6[2]),.dout(n122),.clk(gclk));
	jnot g0051(.din(w_n122_1[1]),.dout(n123),.clk(gclk));
	jand g0052(.dina(w_n88_1[0]),.dinb(w_n91_1[1]),.dout(n124),.clk(gclk));
	jcb g0053(.dina(n124),.dinb(w_n98_2[0]),.dout(n125));
	jcb g0054(.dina(w_dff_B_g1FTjHUN6_0),.dinb(w_n123_1[2]),.dout(n126));
	jand g0055(.dina(w_dff_B_2uIT0MVQ7_0),.dinb(n120),.dout(n127),.clk(gclk));
	jand g0056(.dina(n127),.dinb(w_dff_B_b8xM2L0C0_1),.dout(G361),.clk(gclk));
	jxor g0057(.dina(w_G270_0[1]),.dinb(w_G264_1[0]),.dout(n129),.clk(gclk));
	jxor g0058(.dina(w_G257_1[1]),.dinb(w_n98_1[2]),.dout(n130),.clk(gclk));
	jxor g0059(.dina(n130),.dinb(w_dff_B_DhQRgtAm4_1),.dout(n131),.clk(gclk));
	jnot g0060(.din(w_n131_0[1]),.dout(n132),.clk(gclk));
	jxor g0061(.dina(w_G244_1[1]),.dinb(w_G238_1[1]),.dout(n133),.clk(gclk));
	jxor g0062(.dina(w_G232_1[1]),.dinb(w_n86_0[0]),.dout(n134),.clk(gclk));
	jxor g0063(.dina(n134),.dinb(w_dff_B_QmBhjrpP1_1),.dout(n135),.clk(gclk));
	jxor g0064(.dina(w_n135_0[1]),.dinb(n132),.dout(G358),.clk(gclk));
	jxor g0065(.dina(w_G68_5[0]),.dinb(w_G58_5[0]),.dout(n137),.clk(gclk));
	jnot g0066(.din(w_n137_0[2]),.dout(n138),.clk(gclk));
	jxor g0067(.dina(w_G77_5[0]),.dinb(w_G50_5[0]),.dout(n139),.clk(gclk));
	jxor g0068(.dina(w_dff_B_46XW8r5J1_0),.dinb(n138),.dout(n140),.clk(gclk));
	jnot g0069(.din(w_n140_0[1]),.dout(n141),.clk(gclk));
	jxor g0070(.dina(w_G116_4[1]),.dinb(w_G107_5[0]),.dout(n142),.clk(gclk));
	jxor g0071(.dina(w_G97_5[0]),.dinb(w_n97_2[0]),.dout(n143),.clk(gclk));
	jxor g0072(.dina(n143),.dinb(w_dff_B_tZTxkOmW8_1),.dout(n144),.clk(gclk));
	jxor g0073(.dina(w_n144_0[1]),.dinb(n141),.dout(G351),.clk(gclk));
	jnot g0074(.din(w_G169_1[1]),.dout(n146),.clk(gclk));
	jand g0075(.dina(w_G13_1[0]),.dinb(w_G1_2[1]),.dout(n147),.clk(gclk));
	jnot g0076(.din(w_G33_11[2]),.dout(n148),.clk(gclk));
	jnot g0077(.din(w_G41_1[1]),.dout(n149),.clk(gclk));
	jcb g0078(.dina(w_n149_2[1]),.dinb(w_n148_9[2]),.dout(n150));
	jand g0079(.dina(n150),.dinb(w_n147_0[2]),.dout(n151),.clk(gclk));
	jand g0080(.dina(w_G1698_0[2]),.dinb(w_n148_9[1]),.dout(n152),.clk(gclk));
	jand g0081(.dina(w_n152_3[1]),.dinb(w_G244_1[0]),.dout(n153),.clk(gclk));
	jnot g0082(.din(w_G1698_0[1]),.dout(n154),.clk(gclk));
	jand g0083(.dina(w_n154_0[1]),.dinb(w_n148_9[0]),.dout(n155),.clk(gclk));
	jand g0084(.dina(w_n155_3[1]),.dinb(w_G238_1[0]),.dout(n156),.clk(gclk));
	jand g0085(.dina(w_G116_4[0]),.dinb(w_G33_11[1]),.dout(n157),.clk(gclk));
	jcb g0086(.dina(w_n157_0[2]),.dinb(n156),.dout(n158));
	jcb g0087(.dina(n158),.dinb(n153),.dout(n159));
	jand g0088(.dina(n159),.dinb(w_n151_4[2]),.dout(n160),.clk(gclk));
	jnot g0089(.din(w_G45_1[2]),.dout(n161),.clk(gclk));
	jcb g0090(.dina(w_n161_1[1]),.dinb(w_G1_2[0]),.dout(n162));
	jand g0091(.dina(w_n162_0[2]),.dinb(w_n98_1[1]),.dout(n163),.clk(gclk));
	jnot g0092(.din(w_n163_0[1]),.dout(n164),.clk(gclk));
	jand g0093(.dina(w_G41_1[0]),.dinb(w_G33_11[0]),.dout(n165),.clk(gclk));
	jcb g0094(.dina(n165),.dinb(w_n115_1[0]),.dout(n166));
	jcb g0095(.dina(w_n162_0[1]),.dinb(w_G274_0[2]),.dout(n167));
	jand g0096(.dina(n167),.dinb(w_n166_3[1]),.dout(n168),.clk(gclk));
	jand g0097(.dina(w_dff_B_EVEz00gg4_0),.dinb(n164),.dout(n169),.clk(gclk));
	jcb g0098(.dina(n169),.dinb(n160),.dout(n170));
	jand g0099(.dina(w_n170_0[2]),.dinb(w_n146_3[2]),.dout(n171),.clk(gclk));
	jand g0100(.dina(w_G97_4[2]),.dinb(w_G33_10[2]),.dout(n172),.clk(gclk));
	jand g0101(.dina(w_G68_4[2]),.dinb(w_n148_8[2]),.dout(n173),.clk(gclk));
	jcb g0102(.dina(n173),.dinb(w_G20_6[1]),.dout(n174));
	jcb g0103(.dina(n174),.dinb(w_n172_0[1]),.dout(n175));
	jnot g0104(.din(n175),.dout(n176),.clk(gclk));
	jcb g0105(.dina(w_n112_5[1]),.dinb(w_n113_3[0]),.dout(n177));
	jcb g0106(.dina(n177),.dinb(w_n148_8[1]),.dout(n178));
	jand g0107(.dina(n178),.dinb(w_n115_0[2]),.dout(n179),.clk(gclk));
	jand g0108(.dina(w_n81_0[1]),.dinb(w_n97_1[2]),.dout(n180),.clk(gclk));
	jand g0109(.dina(w_n180_0[1]),.dinb(w_G20_6[0]),.dout(n181),.clk(gclk));
	jcb g0110(.dina(n181),.dinb(w_n179_1[2]),.dout(n182));
	jcb g0111(.dina(n182),.dinb(w_dff_B_DVVSq78l4_1),.dout(n183));
	jand g0112(.dina(w_G20_5[2]),.dinb(w_n113_2[2]),.dout(n184),.clk(gclk));
	jand g0113(.dina(n184),.dinb(w_G13_0[2]),.dout(n185),.clk(gclk));
	jand g0114(.dina(w_n185_3[2]),.dinb(w_n97_1[1]),.dout(n186),.clk(gclk));
	jnot g0115(.din(n186),.dout(n187),.clk(gclk));
	jand g0116(.dina(w_n85_0[1]),.dinb(w_G33_10[1]),.dout(n188),.clk(gclk));
	jcb g0117(.dina(n188),.dinb(w_n147_0[1]),.dout(n189));
	jcb g0118(.dina(w_n185_3[1]),.dinb(w_n189_2[1]),.dout(n190));
	jand g0119(.dina(w_G33_10[0]),.dinb(w_n113_2[1]),.dout(n191),.clk(gclk));
	jcb g0120(.dina(w_n191_0[2]),.dinb(w_n97_1[0]),.dout(n192));
	jcb g0121(.dina(w_dff_B_opaONvPE0_0),.dinb(w_n190_1[2]),.dout(n193));
	jand g0122(.dina(w_dff_B_j2zTilF61_0),.dinb(n187),.dout(n194),.clk(gclk));
	jand g0123(.dina(n194),.dinb(w_dff_B_cL8Xs4078_1),.dout(n195),.clk(gclk));
	jnot g0124(.din(w_G179_2[2]),.dout(n196),.clk(gclk));
	jcb g0125(.dina(w_n154_0[0]),.dinb(w_G33_9[2]),.dout(n197));
	jcb g0126(.dina(w_n197_1[1]),.dinb(w_n103_0[1]),.dout(n198));
	jcb g0127(.dina(w_G1698_0[0]),.dinb(w_G33_9[1]),.dout(n199));
	jcb g0128(.dina(w_n199_1[1]),.dinb(w_n93_0[0]),.dout(n200));
	jnot g0129(.din(w_n157_0[1]),.dout(n201),.clk(gclk));
	jand g0130(.dina(w_n201_0[1]),.dinb(w_dff_B_5wPozv1I6_1),.dout(n202),.clk(gclk));
	jand g0131(.dina(n202),.dinb(w_dff_B_PrZaD5Zv0_1),.dout(n203),.clk(gclk));
	jcb g0132(.dina(n203),.dinb(w_n166_3[0]),.dout(n204));
	jnot g0133(.din(w_G274_0[1]),.dout(n205),.clk(gclk));
	jand g0134(.dina(w_G45_1[1]),.dinb(w_n113_2[0]),.dout(n206),.clk(gclk));
	jand g0135(.dina(w_n206_0[1]),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jcb g0136(.dina(n207),.dinb(w_n151_4[1]),.dout(n208));
	jcb g0137(.dina(n208),.dinb(w_n163_0[0]),.dout(n209));
	jand g0138(.dina(w_dff_B_xzZaUamp2_0),.dinb(n204),.dout(n210),.clk(gclk));
	jand g0139(.dina(w_n210_0[2]),.dinb(w_n196_2[2]),.dout(n211),.clk(gclk));
	jcb g0140(.dina(w_dff_B_1cfpiNrB1_0),.dinb(w_n195_0[1]),.dout(n212));
	jcb g0141(.dina(n212),.dinb(w_dff_B_bFExBmbu0_1),.dout(n213));
	jnot g0142(.din(w_n195_0[0]),.dout(n214),.clk(gclk));
	jand g0143(.dina(w_n210_0[1]),.dinb(w_G190_4[1]),.dout(n215),.clk(gclk));
	jand g0144(.dina(w_n170_0[1]),.dinb(w_G200_4[2]),.dout(n216),.clk(gclk));
	jcb g0145(.dina(w_dff_B_q0dCNmqv6_0),.dinb(n215),.dout(n217));
	jcb g0146(.dina(w_dff_B_GRlG9TWL1_0),.dinb(w_n214_0[1]),.dout(n218));
	jand g0147(.dina(w_n218_0[1]),.dinb(w_n213_0[1]),.dout(n219),.clk(gclk));
	jcb g0148(.dina(w_n197_1[0]),.dinb(w_n98_1[0]),.dout(n220));
	jand g0149(.dina(w_G283_3[2]),.dinb(w_G33_9[0]),.dout(n221),.clk(gclk));
	jnot g0150(.din(w_n221_0[2]),.dout(n222),.clk(gclk));
	jcb g0151(.dina(w_n199_1[0]),.dinb(w_n103_0[0]),.dout(n223));
	jand g0152(.dina(w_dff_B_GhdvqHhs9_0),.dinb(n222),.dout(n224),.clk(gclk));
	jand g0153(.dina(n224),.dinb(w_dff_B_9COU33x02_1),.dout(n225),.clk(gclk));
	jcb g0154(.dina(n225),.dinb(w_n166_2[2]),.dout(n226));
	jcb g0155(.dina(w_n151_4[0]),.dinb(w_n205_0[0]),.dout(n227));
	jcb g0156(.dina(w_n162_0[0]),.dinb(w_G41_0[2]),.dout(n228));
	jcb g0157(.dina(w_n228_0[1]),.dinb(n227),.dout(n229));
	jand g0158(.dina(w_n206_0[0]),.dinb(w_n149_2[0]),.dout(n230),.clk(gclk));
	jcb g0159(.dina(w_n230_0[1]),.dinb(w_n151_3[2]),.dout(n231));
	jcb g0160(.dina(w_n231_0[2]),.dinb(w_n91_1[0]),.dout(n232));
	jand g0161(.dina(n232),.dinb(w_n229_0[2]),.dout(n233),.clk(gclk));
	jand g0162(.dina(n233),.dinb(n226),.dout(n234),.clk(gclk));
	jcb g0163(.dina(w_n234_0[2]),.dinb(w_n146_3[1]),.dout(n235));
	jand g0164(.dina(w_n152_3[0]),.dinb(w_G250_0[1]),.dout(n236),.clk(gclk));
	jand g0165(.dina(w_n155_3[0]),.dinb(w_G244_0[2]),.dout(n237),.clk(gclk));
	jcb g0166(.dina(n237),.dinb(w_n221_0[1]),.dout(n238));
	jcb g0167(.dina(n238),.dinb(n236),.dout(n239));
	jand g0168(.dina(n239),.dinb(w_n151_3[1]),.dout(n240),.clk(gclk));
	jand g0169(.dina(w_n166_2[1]),.dinb(w_G274_0[0]),.dout(n241),.clk(gclk));
	jand g0170(.dina(w_n230_0[0]),.dinb(w_n241_0[1]),.dout(n242),.clk(gclk));
	jand g0171(.dina(w_n228_0[0]),.dinb(w_n166_2[0]),.dout(n243),.clk(gclk));
	jand g0172(.dina(w_n243_0[2]),.dinb(w_G257_1[0]),.dout(n244),.clk(gclk));
	jcb g0173(.dina(w_dff_B_crRIzxv97_0),.dinb(w_n242_0[2]),.dout(n245));
	jcb g0174(.dina(n245),.dinb(n240),.dout(n246));
	jcb g0175(.dina(w_n246_1[1]),.dinb(w_n196_2[1]),.dout(n247));
	jand g0176(.dina(w_dff_B_xIKDQVJe5_0),.dinb(n235),.dout(n248),.clk(gclk));
	jand g0177(.dina(w_G107_4[2]),.dinb(w_G33_8[2]),.dout(n249),.clk(gclk));
	jand g0178(.dina(w_G77_4[2]),.dinb(w_n148_8[0]),.dout(n250),.clk(gclk));
	jcb g0179(.dina(n250),.dinb(w_G20_5[1]),.dout(n251));
	jcb g0180(.dina(n251),.dinb(w_n249_0[1]),.dout(n252));
	jand g0181(.dina(w_G107_4[1]),.dinb(w_G97_4[1]),.dout(n253),.clk(gclk));
	jcb g0182(.dina(n253),.dinb(w_n112_5[0]),.dout(n254));
	jcb g0183(.dina(w_dff_B_I5nmTvxU4_0),.dinb(w_n81_0[0]),.dout(n255));
	jand g0184(.dina(w_n255_0[1]),.dinb(n252),.dout(n256),.clk(gclk));
	jand g0185(.dina(n256),.dinb(w_n189_2[0]),.dout(n257),.clk(gclk));
	jnot g0186(.din(w_n257_0[1]),.dout(n258),.clk(gclk));
	jand g0187(.dina(w_n185_3[0]),.dinb(w_n79_0[0]),.dout(n259),.clk(gclk));
	jnot g0188(.din(w_n259_0[1]),.dout(n260),.clk(gclk));
	jnot g0189(.din(w_n191_0[1]),.dout(n261),.clk(gclk));
	jand g0190(.dina(w_n261_0[1]),.dinb(w_G97_4[0]),.dout(n262),.clk(gclk));
	jnot g0191(.din(w_n262_0[1]),.dout(n263),.clk(gclk));
	jcb g0192(.dina(n263),.dinb(w_n190_1[1]),.dout(n264));
	jand g0193(.dina(n264),.dinb(n260),.dout(n265),.clk(gclk));
	jand g0194(.dina(n265),.dinb(w_dff_B_JIOC8EHz8_1),.dout(n266),.clk(gclk));
	jcb g0195(.dina(n266),.dinb(w_dff_B_7U7WpZzl4_1),.dout(n267));
	jand g0196(.dina(w_n246_1[0]),.dinb(w_G200_4[1]),.dout(n268),.clk(gclk));
	jcb g0197(.dina(w_n112_4[2]),.dinb(w_G1_1[2]),.dout(n269));
	jcb g0198(.dina(w_n269_1[2]),.dinb(w_n114_1[0]),.dout(n270));
	jand g0199(.dina(w_n270_0[1]),.dinb(w_n179_1[1]),.dout(n271),.clk(gclk));
	jand g0200(.dina(w_n262_0[0]),.dinb(w_n271_1[2]),.dout(n272),.clk(gclk));
	jcb g0201(.dina(n272),.dinb(w_n259_0[0]),.dout(n273));
	jcb g0202(.dina(n273),.dinb(w_n257_0[0]),.dout(n274));
	jand g0203(.dina(w_n234_0[1]),.dinb(w_G190_4[0]),.dout(n275),.clk(gclk));
	jcb g0204(.dina(n275),.dinb(w_n274_0[2]),.dout(n276));
	jcb g0205(.dina(n276),.dinb(w_dff_B_OaAB421S6_1),.dout(n277));
	jand g0206(.dina(w_dff_B_zBzpHhf81_0),.dinb(n267),.dout(n278),.clk(gclk));
	jand g0207(.dina(w_n278_0[1]),.dinb(w_n219_0[1]),.dout(n279),.clk(gclk));
	jand g0208(.dina(w_n152_2[2]),.dinb(w_G264_0[2]),.dout(n280),.clk(gclk));
	jand g0209(.dina(w_G303_2[2]),.dinb(w_G33_8[1]),.dout(n281),.clk(gclk));
	jand g0210(.dina(w_n155_2[2]),.dinb(w_G257_0[2]),.dout(n282),.clk(gclk));
	jcb g0211(.dina(n282),.dinb(w_n281_0[1]),.dout(n283));
	jcb g0212(.dina(n283),.dinb(n280),.dout(n284));
	jand g0213(.dina(n284),.dinb(w_n151_3[0]),.dout(n285),.clk(gclk));
	jand g0214(.dina(w_n243_0[1]),.dinb(w_G270_0[0]),.dout(n286),.clk(gclk));
	jcb g0215(.dina(w_dff_B_l1NMarM66_0),.dinb(w_n242_0[1]),.dout(n287));
	jcb g0216(.dina(n287),.dinb(n285),.dout(n288));
	jand g0217(.dina(w_n288_1[1]),.dinb(w_n146_3[0]),.dout(n289),.clk(gclk));
	jand g0218(.dina(w_G97_3[2]),.dinb(w_n148_7[2]),.dout(n290),.clk(gclk));
	jcb g0219(.dina(n290),.dinb(w_G20_5[0]),.dout(n291));
	jcb g0220(.dina(n291),.dinb(w_n221_0[0]),.dout(n292));
	jand g0221(.dina(w_n105_2[0]),.dinb(w_G20_4[2]),.dout(n293),.clk(gclk));
	jnot g0222(.din(n293),.dout(n294),.clk(gclk));
	jand g0223(.dina(n294),.dinb(w_n189_1[2]),.dout(n295),.clk(gclk));
	jand g0224(.dina(n295),.dinb(w_dff_B_I8qsIiur3_1),.dout(n296),.clk(gclk));
	jnot g0225(.din(w_n296_0[1]),.dout(n297),.clk(gclk));
	jand g0226(.dina(w_n185_2[2]),.dinb(w_n105_1[2]),.dout(n298),.clk(gclk));
	jnot g0227(.din(w_n298_0[1]),.dout(n299),.clk(gclk));
	jcb g0228(.dina(w_n191_0[0]),.dinb(w_n105_1[1]),.dout(n300));
	jcb g0229(.dina(w_n300_0[1]),.dinb(w_n190_1[0]),.dout(n301));
	jand g0230(.dina(w_dff_B_N3cNAHsT0_0),.dinb(n299),.dout(n302),.clk(gclk));
	jand g0231(.dina(n302),.dinb(n297),.dout(n303),.clk(gclk));
	jcb g0232(.dina(w_n197_0[2]),.dinb(w_n88_0[2]),.dout(n304));
	jnot g0233(.din(w_n281_0[0]),.dout(n305),.clk(gclk));
	jcb g0234(.dina(w_n199_0[2]),.dinb(w_n91_0[2]),.dout(n306));
	jand g0235(.dina(w_dff_B_NBjz2sFV6_0),.dinb(n305),.dout(n307),.clk(gclk));
	jand g0236(.dina(n307),.dinb(w_dff_B_K7z4jg7I0_1),.dout(n308),.clk(gclk));
	jcb g0237(.dina(n308),.dinb(w_n166_1[2]),.dout(n309));
	jcb g0238(.dina(w_n231_0[1]),.dinb(w_n106_0[0]),.dout(n310));
	jand g0239(.dina(n310),.dinb(w_n229_0[1]),.dout(n311),.clk(gclk));
	jand g0240(.dina(n311),.dinb(n309),.dout(n312),.clk(gclk));
	jand g0241(.dina(w_n312_1[1]),.dinb(w_n196_2[0]),.dout(n313),.clk(gclk));
	jcb g0242(.dina(w_dff_B_lrDaUowg2_0),.dinb(w_n303_0[1]),.dout(n314));
	jcb g0243(.dina(n314),.dinb(w_dff_B_eta8Muoc4_1),.dout(n315));
	jand g0244(.dina(w_n288_1[0]),.dinb(w_G200_4[0]),.dout(n316),.clk(gclk));
	jnot g0245(.din(w_n300_0[0]),.dout(n317),.clk(gclk));
	jand g0246(.dina(n317),.dinb(w_n271_1[1]),.dout(n318),.clk(gclk));
	jcb g0247(.dina(n318),.dinb(w_n298_0[0]),.dout(n319));
	jcb g0248(.dina(w_dff_B_jwuRkkXK5_0),.dinb(w_n296_0[0]),.dout(n320));
	jand g0249(.dina(w_n312_1[0]),.dinb(w_G190_3[2]),.dout(n321),.clk(gclk));
	jcb g0250(.dina(n321),.dinb(w_n320_0[1]),.dout(n322));
	jcb g0251(.dina(n322),.dinb(w_dff_B_BzP9mOHK2_1),.dout(n323));
	jand g0252(.dina(w_dff_B_w4Awezhr4_0),.dinb(w_n315_0[1]),.dout(n324),.clk(gclk));
	jcb g0253(.dina(w_n97_0[2]),.dinb(w_G33_8[0]),.dout(n325));
	jand g0254(.dina(n325),.dinb(w_n112_4[1]),.dout(n326),.clk(gclk));
	jand g0255(.dina(n326),.dinb(w_n201_0[0]),.dout(n327),.clk(gclk));
	jcb g0256(.dina(n327),.dinb(w_n179_1[0]),.dout(n328));
	jcb g0257(.dina(w_n328_0[1]),.dinb(w_G20_4[1]),.dout(n329));
	jand g0258(.dina(n329),.dinb(w_G107_4[0]),.dout(n330),.clk(gclk));
	jand g0259(.dina(w_n328_0[0]),.dinb(w_n270_0[0]),.dout(n331),.clk(gclk));
	jcb g0260(.dina(n331),.dinb(n330),.dout(n332));
	jand g0261(.dina(w_n261_0[0]),.dinb(w_G107_3[2]),.dout(n333),.clk(gclk));
	jand g0262(.dina(n333),.dinb(w_n271_1[0]),.dout(n334),.clk(gclk));
	jnot g0263(.din(w_n334_0[1]),.dout(n335),.clk(gclk));
	jand g0264(.dina(n335),.dinb(w_dff_B_wewM4ZSQ5_1),.dout(n336),.clk(gclk));
	jcb g0265(.dina(w_n197_0[1]),.dinb(w_n91_0[1]),.dout(n337));
	jcb g0266(.dina(w_n199_0[1]),.dinb(w_n98_0[2]),.dout(n338));
	jand g0267(.dina(w_G294_3[1]),.dinb(w_G33_7[2]),.dout(n339),.clk(gclk));
	jnot g0268(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jand g0269(.dina(n340),.dinb(w_dff_B_i14Gol6C4_1),.dout(n341),.clk(gclk));
	jand g0270(.dina(n341),.dinb(w_dff_B_L6FeC3JP5_1),.dout(n342),.clk(gclk));
	jcb g0271(.dina(n342),.dinb(w_n166_1[1]),.dout(n343));
	jcb g0272(.dina(w_n231_0[0]),.dinb(w_n88_0[1]),.dout(n344));
	jand g0273(.dina(n344),.dinb(w_n229_0[0]),.dout(n345),.clk(gclk));
	jand g0274(.dina(n345),.dinb(n343),.dout(n346),.clk(gclk));
	jand g0275(.dina(w_n346_1[1]),.dinb(w_n196_1[2]),.dout(n347),.clk(gclk));
	jand g0276(.dina(w_n152_2[1]),.dinb(w_G257_0[1]),.dout(n348),.clk(gclk));
	jand g0277(.dina(w_n155_2[1]),.dinb(w_G250_0[0]),.dout(n349),.clk(gclk));
	jcb g0278(.dina(w_n339_0[0]),.dinb(n349),.dout(n350));
	jcb g0279(.dina(n350),.dinb(n348),.dout(n351));
	jand g0280(.dina(n351),.dinb(w_n151_2[2]),.dout(n352),.clk(gclk));
	jand g0281(.dina(w_n243_0[0]),.dinb(w_G264_0[1]),.dout(n353),.clk(gclk));
	jcb g0282(.dina(w_dff_B_zYYggNLe3_0),.dinb(w_n242_0[0]),.dout(n354));
	jcb g0283(.dina(n354),.dinb(n352),.dout(n355));
	jand g0284(.dina(w_n355_1[1]),.dinb(w_n146_2[2]),.dout(n356),.clk(gclk));
	jcb g0285(.dina(w_dff_B_fc3BiEcZ2_0),.dinb(n347),.dout(n357));
	jcb g0286(.dina(w_dff_B_yTEEUpH48_0),.dinb(n336),.dout(n358));
	jand g0287(.dina(w_G87_3[0]),.dinb(w_n148_7[1]),.dout(n359),.clk(gclk));
	jcb g0288(.dina(n359),.dinb(w_G20_4[0]),.dout(n360));
	jcb g0289(.dina(n360),.dinb(w_n157_0[0]),.dout(n361));
	jand g0290(.dina(n361),.dinb(w_n189_1[1]),.dout(n362),.clk(gclk));
	jand g0291(.dina(w_n362_0[1]),.dinb(w_n112_4[0]),.dout(n363),.clk(gclk));
	jcb g0292(.dina(n363),.dinb(w_n80_0[2]),.dout(n364));
	jcb g0293(.dina(w_n362_0[0]),.dinb(w_n185_2[1]),.dout(n365));
	jand g0294(.dina(w_dff_B_qA13Ndc32_0),.dinb(n364),.dout(n366),.clk(gclk));
	jcb g0295(.dina(w_n334_0[0]),.dinb(n366),.dout(n367));
	jcb g0296(.dina(w_n355_1[0]),.dinb(w_G190_3[1]),.dout(n368));
	jcb g0297(.dina(w_n346_1[0]),.dinb(w_G200_3[2]),.dout(n369));
	jand g0298(.dina(n369),.dinb(w_dff_B_8fOJpo850_1),.dout(n370),.clk(gclk));
	jcb g0299(.dina(n370),.dinb(w_n367_0[2]),.dout(n371));
	jand g0300(.dina(w_n371_0[1]),.dinb(n358),.dout(n372),.clk(gclk));
	jand g0301(.dina(w_n372_0[1]),.dinb(w_n324_0[1]),.dout(n373),.clk(gclk));
	jand g0302(.dina(w_dff_B_wirumzpe5_0),.dinb(w_n279_0[1]),.dout(n374),.clk(gclk));
	jand g0303(.dina(w_n155_2[0]),.dinb(w_G232_1[0]),.dout(n375),.clk(gclk));
	jand g0304(.dina(w_n152_2[0]),.dinb(w_G238_0[2]),.dout(n376),.clk(gclk));
	jcb g0305(.dina(n376),.dinb(w_n249_0[0]),.dout(n377));
	jcb g0306(.dina(n377),.dinb(n375),.dout(n378));
	jand g0307(.dina(n378),.dinb(w_n151_2[1]),.dout(n379),.clk(gclk));
	jand g0308(.dina(w_n161_1[0]),.dinb(w_n149_1[2]),.dout(n380),.clk(gclk));
	jcb g0309(.dina(n380),.dinb(w_G1_1[1]),.dout(n381));
	jand g0310(.dina(w_n381_0[1]),.dinb(w_n166_1[0]),.dout(n382),.clk(gclk));
	jand g0311(.dina(w_n382_1[1]),.dinb(w_G244_0[1]),.dout(n383),.clk(gclk));
	jnot g0312(.din(w_n381_0[0]),.dout(n384),.clk(gclk));
	jand g0313(.dina(n384),.dinb(w_n241_0[0]),.dout(n385),.clk(gclk));
	jcb g0314(.dina(w_n385_1[1]),.dinb(n383),.dout(n386));
	jcb g0315(.dina(n386),.dinb(n379),.dout(n387));
	jand g0316(.dina(w_n387_1[1]),.dinb(w_n146_2[1]),.dout(n388),.clk(gclk));
	jnot g0317(.din(n388),.dout(n389),.clk(gclk));
	jand g0318(.dina(w_G87_2[2]),.dinb(w_G33_7[1]),.dout(n390),.clk(gclk));
	jand g0319(.dina(w_G58_4[2]),.dinb(w_n148_7[0]),.dout(n391),.clk(gclk));
	jcb g0320(.dina(n391),.dinb(w_G20_3[2]),.dout(n392));
	jcb g0321(.dina(n392),.dinb(w_n390_0[1]),.dout(n393));
	jcb g0322(.dina(w_G77_4[1]),.dinb(w_n112_3[2]),.dout(n394));
	jand g0323(.dina(w_dff_B_vEpVHQhZ6_0),.dinb(w_n189_1[0]),.dout(n395),.clk(gclk));
	jand g0324(.dina(n395),.dinb(w_dff_B_D9Bk1MgI6_1),.dout(n396),.clk(gclk));
	jand g0325(.dina(w_n185_2[0]),.dinb(w_n72_0[2]),.dout(n397),.clk(gclk));
	jand g0326(.dina(w_n269_1[1]),.dinb(w_G77_4[0]),.dout(n398),.clk(gclk));
	jand g0327(.dina(w_dff_B_i1l3Mp175_0),.dinb(w_n271_0[2]),.dout(n399),.clk(gclk));
	jcb g0328(.dina(n399),.dinb(n397),.dout(n400));
	jcb g0329(.dina(n400),.dinb(n396),.dout(n401));
	jcb g0330(.dina(w_n387_1[0]),.dinb(w_G179_2[1]),.dout(n402));
	jand g0331(.dina(n402),.dinb(w_n401_0[2]),.dout(n403),.clk(gclk));
	jand g0332(.dina(w_dff_B_Sph0DQDc9_0),.dinb(n389),.dout(n404),.clk(gclk));
	jnot g0333(.din(w_n404_0[2]),.dout(n405),.clk(gclk));
	jand g0334(.dina(w_n387_0[2]),.dinb(w_G200_3[1]),.dout(n406),.clk(gclk));
	jnot g0335(.din(w_G190_3[0]),.dout(n407),.clk(gclk));
	jcb g0336(.dina(w_n387_0[1]),.dinb(w_n407_2[1]),.dout(n408));
	jnot g0337(.din(n408),.dout(n409),.clk(gclk));
	jcb g0338(.dina(n409),.dinb(w_n401_0[1]),.dout(n410));
	jcb g0339(.dina(n410),.dinb(n406),.dout(n411));
	jand g0340(.dina(w_dff_B_218vRI5f9_0),.dinb(w_n405_0[1]),.dout(n412),.clk(gclk));
	jand g0341(.dina(w_n155_1[2]),.dinb(w_G226_1[0]),.dout(n413),.clk(gclk));
	jand g0342(.dina(w_n152_1[2]),.dinb(w_G232_0[2]),.dout(n414),.clk(gclk));
	jcb g0343(.dina(n414),.dinb(w_n172_0[0]),.dout(n415));
	jcb g0344(.dina(n415),.dinb(n413),.dout(n416));
	jand g0345(.dina(n416),.dinb(w_n151_2[0]),.dout(n417),.clk(gclk));
	jand g0346(.dina(w_n382_1[0]),.dinb(w_G238_0[1]),.dout(n418),.clk(gclk));
	jcb g0347(.dina(n418),.dinb(w_n385_1[0]),.dout(n419));
	jcb g0348(.dina(n419),.dinb(n417),.dout(n420));
	jand g0349(.dina(w_n420_1[1]),.dinb(w_n146_2[0]),.dout(n421),.clk(gclk));
	jnot g0350(.din(n421),.dout(n422),.clk(gclk));
	jand g0351(.dina(w_n269_1[0]),.dinb(w_G68_4[1]),.dout(n423),.clk(gclk));
	jand g0352(.dina(w_dff_B_5R6QWDEa2_0),.dinb(w_n271_0[1]),.dout(n424),.clk(gclk));
	jand g0353(.dina(w_n148_6[2]),.dinb(w_n114_0[2]),.dout(n425),.clk(gclk));
	jnot g0354(.din(w_n425_1[2]),.dout(n426),.clk(gclk));
	jand g0355(.dina(w_n426_0[1]),.dinb(w_n85_0[0]),.dout(n427),.clk(gclk));
	jcb g0356(.dina(n427),.dinb(w_n185_1[2]),.dout(n428));
	jand g0357(.dina(n428),.dinb(w_n75_0[2]),.dout(n429),.clk(gclk));
	jand g0358(.dina(w_G77_3[2]),.dinb(w_G33_7[0]),.dout(n430),.clk(gclk));
	jand g0359(.dina(w_G50_4[2]),.dinb(w_n148_6[1]),.dout(n431),.clk(gclk));
	jcb g0360(.dina(n431),.dinb(w_n430_0[1]),.dout(n432));
	jand g0361(.dina(n432),.dinb(w_n112_3[1]),.dout(n433),.clk(gclk));
	jand g0362(.dina(n433),.dinb(w_n189_0[2]),.dout(n434),.clk(gclk));
	jcb g0363(.dina(w_dff_B_k6F7bK6c4_0),.dinb(n429),.dout(n435));
	jcb g0364(.dina(n435),.dinb(w_dff_B_E2pzOZt54_1),.dout(n436));
	jcb g0365(.dina(w_n420_1[0]),.dinb(w_G179_2[0]),.dout(n437));
	jand g0366(.dina(w_dff_B_t6Zcu4g47_0),.dinb(w_n436_0[2]),.dout(n438),.clk(gclk));
	jand g0367(.dina(n438),.dinb(n422),.dout(n439),.clk(gclk));
	jnot g0368(.din(w_n439_1[1]),.dout(n440),.clk(gclk));
	jand g0369(.dina(w_n420_0[2]),.dinb(w_G200_3[0]),.dout(n441),.clk(gclk));
	jcb g0370(.dina(w_n420_0[1]),.dinb(w_n407_2[0]),.dout(n442));
	jnot g0371(.din(n442),.dout(n443),.clk(gclk));
	jcb g0372(.dina(n443),.dinb(w_n436_0[1]),.dout(n444));
	jcb g0373(.dina(n444),.dinb(n441),.dout(n445));
	jand g0374(.dina(w_n445_0[1]),.dinb(n440),.dout(n446),.clk(gclk));
	jand g0375(.dina(w_n446_0[1]),.dinb(w_n412_0[1]),.dout(n447),.clk(gclk));
	jand g0376(.dina(w_n152_1[1]),.dinb(w_G223_0[1]),.dout(n448),.clk(gclk));
	jand g0377(.dina(w_n155_1[1]),.dinb(w_dff_B_HLS7OORf1_1),.dout(n449),.clk(gclk));
	jcb g0378(.dina(n449),.dinb(w_n430_0[0]),.dout(n450));
	jcb g0379(.dina(n450),.dinb(n448),.dout(n451));
	jand g0380(.dina(n451),.dinb(w_n151_1[2]),.dout(n452),.clk(gclk));
	jand g0381(.dina(w_n382_0[2]),.dinb(w_G226_0[2]),.dout(n453),.clk(gclk));
	jcb g0382(.dina(n453),.dinb(w_n385_0[2]),.dout(n454));
	jcb g0383(.dina(n454),.dinb(n452),.dout(n455));
	jand g0384(.dina(w_n455_0[2]),.dinb(w_n146_1[2]),.dout(n456),.clk(gclk));
	jand g0385(.dina(w_n269_0[2]),.dinb(w_G50_4[1]),.dout(n457),.clk(gclk));
	jnot g0386(.din(n457),.dout(n458),.clk(gclk));
	jcb g0387(.dina(n458),.dinb(w_n190_0[2]),.dout(n459));
	jcb g0388(.dina(w_n77_0[0]),.dinb(w_n112_3[0]),.dout(n460));
	jnot g0389(.din(w_G150_3[1]),.dout(n461),.clk(gclk));
	jand g0390(.dina(w_n148_6[0]),.dinb(w_n112_2[2]),.dout(n462),.clk(gclk));
	jnot g0391(.din(w_n462_0[2]),.dout(n463),.clk(gclk));
	jcb g0392(.dina(n463),.dinb(w_dff_B_vha6vETx4_1),.dout(n464));
	jand g0393(.dina(w_G33_6[2]),.dinb(w_n112_2[1]),.dout(n465),.clk(gclk));
	jand g0394(.dina(w_n465_0[1]),.dinb(w_G58_4[1]),.dout(n466),.clk(gclk));
	jnot g0395(.din(n466),.dout(n467),.clk(gclk));
	jand g0396(.dina(n467),.dinb(w_dff_B_LIelNfwt4_1),.dout(n468),.clk(gclk));
	jand g0397(.dina(n468),.dinb(w_dff_B_INQMja0C0_1),.dout(n469),.clk(gclk));
	jcb g0398(.dina(n469),.dinb(w_n179_0[2]),.dout(n470));
	jand g0399(.dina(w_n185_1[1]),.dinb(w_n73_2[0]),.dout(n471),.clk(gclk));
	jnot g0400(.din(n471),.dout(n472),.clk(gclk));
	jand g0401(.dina(w_dff_B_Nvo7ve6m3_0),.dinb(n470),.dout(n473),.clk(gclk));
	jand g0402(.dina(n473),.dinb(w_dff_B_DwUkk4SC4_1),.dout(n474),.clk(gclk));
	jnot g0403(.din(w_n455_0[1]),.dout(n475),.clk(gclk));
	jand g0404(.dina(w_n475_0[1]),.dinb(w_n196_1[1]),.dout(n476),.clk(gclk));
	jcb g0405(.dina(w_dff_B_C3Zh2WT72_0),.dinb(w_n474_0[1]),.dout(n477));
	jcb g0406(.dina(n477),.dinb(w_dff_B_BszKyM8a9_1),.dout(n478));
	jnot g0407(.din(w_n474_0[0]),.dout(n479),.clk(gclk));
	jand g0408(.dina(w_n475_0[0]),.dinb(w_G190_2[2]),.dout(n480),.clk(gclk));
	jand g0409(.dina(w_n455_0[0]),.dinb(w_G200_2[2]),.dout(n481),.clk(gclk));
	jcb g0410(.dina(w_dff_B_pmKtcmWA5_0),.dinb(n480),.dout(n482));
	jcb g0411(.dina(w_dff_B_eUERuVKn4_0),.dinb(w_n479_0[1]),.dout(n483));
	jand g0412(.dina(w_n483_0[1]),.dinb(w_n478_0[1]),.dout(n484),.clk(gclk));
	jand g0413(.dina(w_n152_1[0]),.dinb(w_G226_0[1]),.dout(n485),.clk(gclk));
	jand g0414(.dina(w_n155_1[0]),.dinb(w_G223_0[0]),.dout(n486),.clk(gclk));
	jcb g0415(.dina(n486),.dinb(w_n390_0[0]),.dout(n487));
	jcb g0416(.dina(n487),.dinb(n485),.dout(n488));
	jand g0417(.dina(n488),.dinb(w_n151_1[1]),.dout(n489),.clk(gclk));
	jand g0418(.dina(w_n382_0[1]),.dinb(w_G232_0[1]),.dout(n490),.clk(gclk));
	jcb g0419(.dina(n490),.dinb(w_n385_0[1]),.dout(n491));
	jcb g0420(.dina(n491),.dinb(n489),.dout(n492));
	jand g0421(.dina(w_n492_0[2]),.dinb(w_n146_1[1]),.dout(n493),.clk(gclk));
	jand g0422(.dina(w_n269_0[1]),.dinb(w_G58_4[0]),.dout(n494),.clk(gclk));
	jnot g0423(.din(n494),.dout(n495),.clk(gclk));
	jcb g0424(.dina(n495),.dinb(w_n190_0[1]),.dout(n496));
	jcb g0425(.dina(w_n137_0[1]),.dinb(w_n112_2[0]),.dout(n497));
	jand g0426(.dina(w_n462_0[1]),.dinb(w_G159_3[2]),.dout(n498),.clk(gclk));
	jand g0427(.dina(w_n465_0[0]),.dinb(w_G68_4[0]),.dout(n499),.clk(gclk));
	jcb g0428(.dina(n499),.dinb(n498),.dout(n500));
	jnot g0429(.din(n500),.dout(n501),.clk(gclk));
	jand g0430(.dina(n501),.dinb(w_dff_B_kcBHfiiB6_1),.dout(n502),.clk(gclk));
	jcb g0431(.dina(n502),.dinb(w_n179_0[1]),.dout(n503));
	jand g0432(.dina(w_n185_1[0]),.dinb(w_n74_0[2]),.dout(n504),.clk(gclk));
	jnot g0433(.din(n504),.dout(n505),.clk(gclk));
	jand g0434(.dina(n505),.dinb(n503),.dout(n506),.clk(gclk));
	jand g0435(.dina(n506),.dinb(w_dff_B_5hryCipb2_1),.dout(n507),.clk(gclk));
	jnot g0436(.din(w_n492_0[1]),.dout(n508),.clk(gclk));
	jand g0437(.dina(w_n508_0[1]),.dinb(w_n196_1[0]),.dout(n509),.clk(gclk));
	jcb g0438(.dina(w_dff_B_vYoGX6kR4_0),.dinb(w_n507_0[1]),.dout(n510));
	jcb g0439(.dina(n510),.dinb(w_dff_B_EmiIeIdo0_1),.dout(n511));
	jnot g0440(.din(w_n507_0[0]),.dout(n512),.clk(gclk));
	jand g0441(.dina(w_n508_0[0]),.dinb(w_G190_2[1]),.dout(n513),.clk(gclk));
	jand g0442(.dina(w_n492_0[0]),.dinb(w_G200_2[1]),.dout(n514),.clk(gclk));
	jcb g0443(.dina(w_dff_B_FtEUyvTn6_0),.dinb(n513),.dout(n515));
	jcb g0444(.dina(w_dff_B_KhwKB54G4_0),.dinb(w_n512_0[1]),.dout(n516));
	jand g0445(.dina(w_n516_0[1]),.dinb(w_n511_0[1]),.dout(n517),.clk(gclk));
	jand g0446(.dina(w_n517_0[1]),.dinb(w_n484_0[1]),.dout(n518),.clk(gclk));
	jand g0447(.dina(n518),.dinb(w_dff_B_pVqq1Jlu5_1),.dout(n519),.clk(gclk));
	jand g0448(.dina(w_n519_1[2]),.dinb(w_n374_0[1]),.dout(G372),.clk(gclk));
	jcb g0449(.dina(w_n355_0[2]),.dinb(w_G179_1[2]),.dout(n521));
	jcb g0450(.dina(w_n346_0[2]),.dinb(w_G169_1[0]),.dout(n522));
	jand g0451(.dina(n522),.dinb(w_dff_B_pK93kYGq3_1),.dout(n523),.clk(gclk));
	jand g0452(.dina(w_n523_0[1]),.dinb(w_n367_0[1]),.dout(n524),.clk(gclk));
	jcb g0453(.dina(w_n312_0[2]),.dinb(w_G169_0[2]),.dout(n525));
	jcb g0454(.dina(w_n288_0[2]),.dinb(w_G179_1[1]),.dout(n526));
	jand g0455(.dina(w_dff_B_0Br3Y3Xv2_0),.dinb(w_n320_0[0]),.dout(n527),.clk(gclk));
	jand g0456(.dina(n527),.dinb(w_dff_B_bJzwrDL81_1),.dout(n528),.clk(gclk));
	jand g0457(.dina(w_n371_0[0]),.dinb(w_n528_0[1]),.dout(n529),.clk(gclk));
	jcb g0458(.dina(n529),.dinb(w_n524_0[1]),.dout(n530));
	jand g0459(.dina(w_dff_B_Mc9vSWlq9_0),.dinb(w_n279_0[0]),.dout(n531),.clk(gclk));
	jnot g0460(.din(w_n213_0[0]),.dout(n532),.clk(gclk));
	jand g0461(.dina(w_n246_0[2]),.dinb(w_G169_0[1]),.dout(n533),.clk(gclk));
	jand g0462(.dina(w_n234_0[0]),.dinb(w_G179_1[0]),.dout(n534),.clk(gclk));
	jcb g0463(.dina(w_n534_0[1]),.dinb(w_dff_B_UtzkZXLy9_1),.dout(n535));
	jand g0464(.dina(w_n274_0[1]),.dinb(n535),.dout(n536),.clk(gclk));
	jand g0465(.dina(w_n536_0[2]),.dinb(w_n218_0[0]),.dout(n537),.clk(gclk));
	jcb g0466(.dina(n537),.dinb(w_n532_0[1]),.dout(n538));
	jcb g0467(.dina(w_dff_B_eFv68KBx7_0),.dinb(n531),.dout(n539));
	jand g0468(.dina(w_n539_0[1]),.dinb(w_n519_1[1]),.dout(n540),.clk(gclk));
	jnot g0469(.din(w_n478_0[0]),.dout(n541),.clk(gclk));
	jnot g0470(.din(w_n511_0[0]),.dout(n542),.clk(gclk));
	jcb g0471(.dina(w_n439_1[0]),.dinb(w_n404_0[1]),.dout(n543));
	jand g0472(.dina(w_n543_0[1]),.dinb(w_n445_0[0]),.dout(n544),.clk(gclk));
	jcb g0473(.dina(n544),.dinb(w_n542_0[2]),.dout(n545));
	jand g0474(.dina(n545),.dinb(w_n516_0[0]),.dout(n546),.clk(gclk));
	jcb g0475(.dina(n546),.dinb(w_n541_0[1]),.dout(n547));
	jand g0476(.dina(n547),.dinb(w_n483_0[0]),.dout(n548),.clk(gclk));
	jcb g0477(.dina(w_n548_0[2]),.dinb(n540),.dout(G369));
	jand g0478(.dina(w_n112_1[2]),.dinb(w_G13_0[1]),.dout(n550),.clk(gclk));
	jand g0479(.dina(w_G213_0[2]),.dinb(w_n113_1[2]),.dout(n551),.clk(gclk));
	jand g0480(.dina(n551),.dinb(w_n550_0[1]),.dout(n552),.clk(gclk));
	jand g0481(.dina(w_n552_1[1]),.dinb(w_G343_0[1]),.dout(n553),.clk(gclk));
	jnot g0482(.din(w_n553_2[2]),.dout(n554),.clk(gclk));
	jand g0483(.dina(w_n554_3[2]),.dinb(w_n524_0[0]),.dout(n555),.clk(gclk));
	jand g0484(.dina(w_n554_3[1]),.dinb(w_n528_0[0]),.dout(n556),.clk(gclk));
	jand g0485(.dina(w_n553_2[1]),.dinb(w_n367_0[0]),.dout(n557),.clk(gclk));
	jnot g0486(.din(w_n557_0[1]),.dout(n558),.clk(gclk));
	jand g0487(.dina(w_dff_B_FaljJk7V4_0),.dinb(w_n372_0[0]),.dout(n559),.clk(gclk));
	jand g0488(.dina(w_n557_0[0]),.dinb(w_n523_0[0]),.dout(n560),.clk(gclk));
	jcb g0489(.dina(w_dff_B_Zx7LqFSw7_0),.dinb(n559),.dout(n561));
	jand g0490(.dina(w_n561_0[2]),.dinb(w_n556_0[1]),.dout(n562),.clk(gclk));
	jcb g0491(.dina(n562),.dinb(w_dff_B_ZwcaPGGG5_1),.dout(n563));
	jnot g0492(.din(w_n561_0[1]),.dout(n564),.clk(gclk));
	jnot g0493(.din(w_G330_0[1]),.dout(n565),.clk(gclk));
	jnot g0494(.din(w_n324_0[0]),.dout(n566),.clk(gclk));
	jcb g0495(.dina(w_n554_3[0]),.dinb(w_n303_0[0]),.dout(n567));
	jnot g0496(.din(w_n567_0[1]),.dout(n568),.clk(gclk));
	jcb g0497(.dina(w_dff_B_o9wqmrq05_0),.dinb(n566),.dout(n569));
	jcb g0498(.dina(w_n567_0[0]),.dinb(w_n315_0[0]),.dout(n570));
	jand g0499(.dina(w_dff_B_elJ768Fw9_0),.dinb(n569),.dout(n571),.clk(gclk));
	jcb g0500(.dina(w_n571_0[2]),.dinb(w_n565_0[1]),.dout(n572));
	jcb g0501(.dina(w_n572_0[2]),.dinb(w_n564_0[1]),.dout(n573));
	jnot g0502(.din(w_n573_0[2]),.dout(n574),.clk(gclk));
	jcb g0503(.dina(n574),.dinb(w_n563_0[2]),.dout(G399));
	jand g0504(.dina(w_n554_2[2]),.dinb(w_n539_0[0]),.dout(n576),.clk(gclk));
	jcb g0505(.dina(w_n553_2[0]),.dinb(w_n374_0[0]),.dout(n577));
	jand g0506(.dina(w_n346_0[1]),.dinb(w_n210_0[0]),.dout(n578),.clk(gclk));
	jand g0507(.dina(n578),.dinb(w_n312_0[1]),.dout(n579),.clk(gclk));
	jand g0508(.dina(n579),.dinb(w_n534_0[0]),.dout(n580),.clk(gclk));
	jand g0509(.dina(w_n288_0[1]),.dinb(w_n196_0[2]),.dout(n581),.clk(gclk));
	jand g0510(.dina(w_n355_0[1]),.dinb(w_n246_0[1]),.dout(n582),.clk(gclk));
	jand g0511(.dina(n582),.dinb(w_n170_0[0]),.dout(n583),.clk(gclk));
	jand g0512(.dina(n583),.dinb(w_dff_B_IymNsGxt3_1),.dout(n584),.clk(gclk));
	jcb g0513(.dina(n584),.dinb(w_n554_2[1]),.dout(n585));
	jcb g0514(.dina(w_dff_B_xJhhQOrv7_0),.dinb(n580),.dout(n586));
	jand g0515(.dina(n586),.dinb(w_G330_0[0]),.dout(n587),.clk(gclk));
	jand g0516(.dina(w_dff_B_zDwXkz7L6_0),.dinb(n577),.dout(n588),.clk(gclk));
	jcb g0517(.dina(w_n588_1[1]),.dinb(w_n576_1[1]),.dout(n589));
	jand g0518(.dina(w_n589_1[2]),.dinb(w_n113_1[1]),.dout(n590),.clk(gclk));
	jand g0519(.dina(w_n122_1[0]),.dinb(w_n149_1[1]),.dout(n591),.clk(gclk));
	jnot g0520(.din(w_n591_1[1]),.dout(n592),.clk(gclk));
	jand g0521(.dina(w_n180_0[0]),.dinb(w_n105_1[0]),.dout(n593),.clk(gclk));
	jand g0522(.dina(w_n593_0[2]),.dinb(w_G1_1[0]),.dout(n594),.clk(gclk));
	jand g0523(.dina(n594),.dinb(w_n592_2[1]),.dout(n595),.clk(gclk));
	jand g0524(.dina(w_n591_1[0]),.dinb(w_n118_0[1]),.dout(n596),.clk(gclk));
	jcb g0525(.dina(w_dff_B_am17GXv75_0),.dinb(n595),.dout(n597));
	jcb g0526(.dina(w_dff_B_woz0rSSW2_0),.dinb(n590),.dout(G364));
	jand g0527(.dina(w_n571_0[1]),.dinb(w_n565_0[0]),.dout(n599),.clk(gclk));
	jnot g0528(.din(n599),.dout(n600),.clk(gclk));
	jand g0529(.dina(w_n550_0[0]),.dinb(w_G45_1[0]),.dout(n601),.clk(gclk));
	jcb g0530(.dina(n601),.dinb(w_n113_1[0]),.dout(n602));
	jnot g0531(.din(w_n602_0[1]),.dout(n603),.clk(gclk));
	jand g0532(.dina(w_n603_2[1]),.dinb(w_n592_2[0]),.dout(n604),.clk(gclk));
	jnot g0533(.din(w_n604_2[1]),.dout(n605),.clk(gclk));
	jand g0534(.dina(w_n605_1[2]),.dinb(w_n572_0[1]),.dout(n606),.clk(gclk));
	jand g0535(.dina(w_dff_B_VudIogzL6_0),.dinb(n600),.dout(n607),.clk(gclk));
	jand g0536(.dina(w_n462_0[0]),.dinb(w_n114_0[1]),.dout(n608),.clk(gclk));
	jand g0537(.dina(w_n608_1[2]),.dinb(w_n571_0[0]),.dout(n609),.clk(gclk));
	jnot g0538(.din(n609),.dout(n610),.clk(gclk));
	jand g0539(.dina(w_n146_1[0]),.dinb(w_G20_3[1]),.dout(n611),.clk(gclk));
	jcb g0540(.dina(n611),.dinb(w_n115_0[1]),.dout(n612));
	jand g0541(.dina(w_G179_0[2]),.dinb(w_G20_3[0]),.dout(n613),.clk(gclk));
	jnot g0542(.din(w_n613_1[1]),.dout(n614),.clk(gclk));
	jand g0543(.dina(w_G200_2[0]),.dinb(w_G20_2[2]),.dout(n615),.clk(gclk));
	jand g0544(.dina(w_n615_0[1]),.dinb(n614),.dout(n616),.clk(gclk));
	jand g0545(.dina(w_n616_0[1]),.dinb(w_G190_2[0]),.dout(n617),.clk(gclk));
	jand g0546(.dina(w_n617_6[1]),.dinb(w_G303_2[1]),.dout(n618),.clk(gclk));
	jand g0547(.dina(w_n407_1[2]),.dinb(w_G20_2[1]),.dout(n619),.clk(gclk));
	jnot g0548(.din(w_n619_0[1]),.dout(n620),.clk(gclk));
	jcb g0549(.dina(w_n615_0[0]),.dinb(w_n613_1[0]),.dout(n621));
	jnot g0550(.din(n621),.dout(n622),.clk(gclk));
	jand g0551(.dina(w_n622_0[1]),.dinb(n620),.dout(n623),.clk(gclk));
	jand g0552(.dina(w_n623_5[1]),.dinb(w_G294_3[0]),.dout(n624),.clk(gclk));
	jnot g0553(.din(w_G200_1[2]),.dout(n625),.clk(gclk));
	jand g0554(.dina(w_n613_0[2]),.dinb(n625),.dout(n626),.clk(gclk));
	jand g0555(.dina(w_n626_0[1]),.dinb(w_G190_1[2]),.dout(n627),.clk(gclk));
	jand g0556(.dina(w_n627_7[1]),.dinb(w_G322_0[2]),.dout(n628),.clk(gclk));
	jcb g0557(.dina(w_dff_B_Nf5ZYQsw4_0),.dinb(n624),.dout(n629));
	jcb g0558(.dina(n629),.dinb(n618),.dout(n630));
	jand g0559(.dina(w_n622_0[0]),.dinb(w_n619_0[0]),.dout(n631),.clk(gclk));
	jand g0560(.dina(w_n631_7[1]),.dinb(w_dff_B_kjHWZixp2_1),.dout(n632),.clk(gclk));
	jcb g0561(.dina(n632),.dinb(w_n148_5[2]),.dout(n633));
	jand g0562(.dina(w_n616_0[0]),.dinb(w_n407_1[1]),.dout(n634),.clk(gclk));
	jand g0563(.dina(w_n634_4[1]),.dinb(w_G283_3[1]),.dout(n635),.clk(gclk));
	jand g0564(.dina(w_n626_0[0]),.dinb(w_n407_1[0]),.dout(n636),.clk(gclk));
	jand g0565(.dina(w_n636_7[1]),.dinb(w_G311_1[2]),.dout(n637),.clk(gclk));
	jcb g0566(.dina(w_dff_B_89NlwPhh7_0),.dinb(n635),.dout(n638));
	jand g0567(.dina(w_n613_0[1]),.dinb(w_G200_1[1]),.dout(n639),.clk(gclk));
	jand g0568(.dina(w_n639_0[1]),.dinb(w_G190_1[1]),.dout(n640),.clk(gclk));
	jand g0569(.dina(w_n640_7[1]),.dinb(w_G326_0[1]),.dout(n641),.clk(gclk));
	jand g0570(.dina(w_n639_0[0]),.dinb(w_n407_0[2]),.dout(n642),.clk(gclk));
	jand g0571(.dina(w_n642_7[1]),.dinb(w_G317_1[1]),.dout(n643),.clk(gclk));
	jcb g0572(.dina(n643),.dinb(n641),.dout(n644));
	jcb g0573(.dina(w_dff_B_dI0eegyn0_0),.dinb(n638),.dout(n645));
	jcb g0574(.dina(n645),.dinb(w_dff_B_3wSKf3w46_1),.dout(n646));
	jcb g0575(.dina(n646),.dinb(n630),.dout(n647));
	jand g0576(.dina(w_n631_7[0]),.dinb(w_G159_3[1]),.dout(n648),.clk(gclk));
	jand g0577(.dina(w_n640_7[0]),.dinb(w_G50_4[0]),.dout(n649),.clk(gclk));
	jand g0578(.dina(w_n642_7[0]),.dinb(w_G68_3[2]),.dout(n650),.clk(gclk));
	jcb g0579(.dina(n650),.dinb(n649),.dout(n651));
	jcb g0580(.dina(n651),.dinb(n648),.dout(n652));
	jnot g0581(.din(n652),.dout(n653),.clk(gclk));
	jand g0582(.dina(w_n617_6[0]),.dinb(w_G87_2[1]),.dout(n654),.clk(gclk));
	jnot g0583(.din(w_n654_0[1]),.dout(n655),.clk(gclk));
	jand g0584(.dina(n655),.dinb(w_n148_5[1]),.dout(n656),.clk(gclk));
	jand g0585(.dina(w_n634_4[0]),.dinb(w_G107_3[1]),.dout(n657),.clk(gclk));
	jand g0586(.dina(w_n636_7[0]),.dinb(w_G77_3[1]),.dout(n658),.clk(gclk));
	jcb g0587(.dina(w_dff_B_FpeKF35t2_0),.dinb(w_n657_0[1]),.dout(n659));
	jand g0588(.dina(w_n627_7[0]),.dinb(w_G58_3[2]),.dout(n660),.clk(gclk));
	jand g0589(.dina(w_n623_5[0]),.dinb(w_G97_3[1]),.dout(n661),.clk(gclk));
	jcb g0590(.dina(w_n661_0[1]),.dinb(w_dff_B_cY4O8HI96_1),.dout(n662));
	jcb g0591(.dina(n662),.dinb(n659),.dout(n663));
	jnot g0592(.din(n663),.dout(n664),.clk(gclk));
	jand g0593(.dina(w_dff_B_JjmVLEll5_0),.dinb(n656),.dout(n665),.clk(gclk));
	jand g0594(.dina(n665),.dinb(w_dff_B_ZfTKSLIY4_1),.dout(n666),.clk(gclk));
	jnot g0595(.din(n666),.dout(n667),.clk(gclk));
	jand g0596(.dina(n667),.dinb(w_dff_B_Xa2q3nUo6_1),.dout(n668),.clk(gclk));
	jcb g0597(.dina(n668),.dinb(w_n612_4[1]),.dout(n669));
	jnot g0598(.din(w_n608_1[1]),.dout(n670),.clk(gclk));
	jand g0599(.dina(w_n612_4[0]),.dinb(n670),.dout(n671),.clk(gclk));
	jnot g0600(.din(n671),.dout(n672),.clk(gclk));
	jand g0601(.dina(w_n140_0[0]),.dinb(w_G45_0[2]),.dout(n673),.clk(gclk));
	jand g0602(.dina(w_n118_0[0]),.dinb(w_n161_0[2]),.dout(n674),.clk(gclk));
	jand g0603(.dina(w_n122_0[2]),.dinb(w_G33_6[1]),.dout(n675),.clk(gclk));
	jnot g0604(.din(w_n675_0[2]),.dout(n676),.clk(gclk));
	jcb g0605(.dina(w_n676_0[1]),.dinb(n674),.dout(n677));
	jcb g0606(.dina(n677),.dinb(w_dff_B_qFYVwUnH9_1),.dout(n678));
	jand g0607(.dina(w_n123_1[1]),.dinb(w_n105_0[2]),.dout(n679),.clk(gclk));
	jand g0608(.dina(w_n122_0[1]),.dinb(w_n148_5[0]),.dout(n680),.clk(gclk));
	jand g0609(.dina(w_n680_0[1]),.dinb(w_G355_0),.dout(n681),.clk(gclk));
	jcb g0610(.dina(n681),.dinb(w_dff_B_kDfzSqZk9_1),.dout(n682));
	jnot g0611(.din(n682),.dout(n683),.clk(gclk));
	jand g0612(.dina(n683),.dinb(w_dff_B_nb4eicKF1_1),.dout(n684),.clk(gclk));
	jcb g0613(.dina(n684),.dinb(w_n672_1[1]),.dout(n685));
	jand g0614(.dina(n685),.dinb(w_n604_2[0]),.dout(n686),.clk(gclk));
	jand g0615(.dina(w_dff_B_GTezD0Qw4_0),.dinb(n669),.dout(n687),.clk(gclk));
	jand g0616(.dina(n687),.dinb(n610),.dout(n688),.clk(gclk));
	jcb g0617(.dina(n688),.dinb(n607),.dout(G396_fa_));
	jnot g0618(.din(w_n588_1[0]),.dout(n690),.clk(gclk));
	jnot g0619(.din(w_n401_0[0]),.dout(n691),.clk(gclk));
	jcb g0620(.dina(w_n554_2[0]),.dinb(n691),.dout(n692));
	jand g0621(.dina(w_n692_0[1]),.dinb(w_n412_0[0]),.dout(n693),.clk(gclk));
	jcb g0622(.dina(w_n692_0[0]),.dinb(w_n405_0[0]),.dout(n694));
	jnot g0623(.din(n694),.dout(n695),.clk(gclk));
	jcb g0624(.dina(w_dff_B_Vkewf4pA1_0),.dinb(n693),.dout(n696));
	jxor g0625(.dina(w_n696_1[2]),.dinb(w_n576_1[0]),.dout(n697),.clk(gclk));
	jnot g0626(.din(n697),.dout(n698),.clk(gclk));
	jand g0627(.dina(n698),.dinb(w_dff_B_lVDmVpR90_1),.dout(n699),.clk(gclk));
	jcb g0628(.dina(w_n991_0[2]),.dinb(w_n604_1[2]),.dout(n701));
	jcb g0629(.dina(w_dff_B_JiVUAAap8_0),.dinb(n699),.dout(n702));
	jnot g0630(.din(w_n696_1[1]),.dout(n703),.clk(gclk));
	jand g0631(.dina(n703),.dinb(w_n425_1[1]),.dout(n704),.clk(gclk));
	jnot g0632(.din(n704),.dout(n705),.clk(gclk));
	jand g0633(.dina(w_n631_6[2]),.dinb(w_G132_1[1]),.dout(n706),.clk(gclk));
	jand g0634(.dina(w_n623_4[2]),.dinb(w_G58_3[1]),.dout(n707),.clk(gclk));
	jand g0635(.dina(w_n642_6[2]),.dinb(w_G150_3[0]),.dout(n708),.clk(gclk));
	jcb g0636(.dina(w_dff_B_iNLtdpIO2_0),.dinb(n707),.dout(n709));
	jcb g0637(.dina(n709),.dinb(w_dff_B_zPIqeoSO7_1),.dout(n710));
	jand g0638(.dina(w_n617_5[2]),.dinb(w_G50_3[2]),.dout(n711),.clk(gclk));
	jcb g0639(.dina(n711),.dinb(w_G33_6[0]),.dout(n712));
	jand g0640(.dina(w_n636_6[2]),.dinb(w_G159_3[0]),.dout(n713),.clk(gclk));
	jand g0641(.dina(w_n627_6[2]),.dinb(w_G143_2[1]),.dout(n714),.clk(gclk));
	jcb g0642(.dina(n714),.dinb(n713),.dout(n715));
	jand g0643(.dina(w_n640_6[2]),.dinb(w_G137_1[2]),.dout(n716),.clk(gclk));
	jand g0644(.dina(w_n634_3[2]),.dinb(w_G68_3[1]),.dout(n717),.clk(gclk));
	jcb g0645(.dina(w_n717_0[1]),.dinb(w_dff_B_MdgUWO5j9_1),.dout(n718));
	jcb g0646(.dina(n718),.dinb(w_dff_B_86WmmvN65_1),.dout(n719));
	jcb g0647(.dina(n719),.dinb(n712),.dout(n720));
	jcb g0648(.dina(n720),.dinb(n710),.dout(n721));
	jand g0649(.dina(w_n631_6[1]),.dinb(w_G311_1[1]),.dout(n722),.clk(gclk));
	jand g0650(.dina(w_n617_5[1]),.dinb(w_G107_3[0]),.dout(n723),.clk(gclk));
	jand g0651(.dina(w_n642_6[1]),.dinb(w_G283_3[0]),.dout(n724),.clk(gclk));
	jcb g0652(.dina(w_dff_B_5ccDlyQl1_0),.dinb(n723),.dout(n725));
	jcb g0653(.dina(n725),.dinb(w_dff_B_DQhw4aS97_1),.dout(n726));
	jnot g0654(.din(n726),.dout(n727),.clk(gclk));
	jand g0655(.dina(w_n634_3[1]),.dinb(w_G87_2[0]),.dout(n728),.clk(gclk));
	jnot g0656(.din(w_n728_0[1]),.dout(n729),.clk(gclk));
	jand g0657(.dina(n729),.dinb(w_G33_5[2]),.dout(n730),.clk(gclk));
	jand g0658(.dina(w_n636_6[1]),.dinb(w_G116_3[2]),.dout(n731),.clk(gclk));
	jand g0659(.dina(w_n627_6[1]),.dinb(w_G294_2[2]),.dout(n732),.clk(gclk));
	jcb g0660(.dina(n732),.dinb(n731),.dout(n733));
	jand g0661(.dina(w_n640_6[1]),.dinb(w_G303_2[0]),.dout(n734),.clk(gclk));
	jcb g0662(.dina(w_dff_B_Zrtp0TWN6_0),.dinb(w_n661_0[0]),.dout(n735));
	jcb g0663(.dina(n735),.dinb(w_dff_B_nCwovcnt8_1),.dout(n736));
	jnot g0664(.din(n736),.dout(n737),.clk(gclk));
	jand g0665(.dina(w_dff_B_S29NIsBY5_0),.dinb(n730),.dout(n738),.clk(gclk));
	jand g0666(.dina(n738),.dinb(w_dff_B_3P2caIMQ0_1),.dout(n739),.clk(gclk));
	jnot g0667(.din(n739),.dout(n740),.clk(gclk));
	jand g0668(.dina(n740),.dinb(w_dff_B_2tEorJjR7_1),.dout(n741),.clk(gclk));
	jcb g0669(.dina(n741),.dinb(w_n612_3[2]),.dout(n742));
	jand g0670(.dina(w_n612_3[1]),.dinb(w_n426_0[0]),.dout(n743),.clk(gclk));
	jand g0671(.dina(w_n743_1[1]),.dinb(w_n72_0[1]),.dout(n744),.clk(gclk));
	jcb g0672(.dina(w_dff_B_XuRRvTNa2_0),.dinb(w_n605_1[1]),.dout(n745));
	jnot g0673(.din(n745),.dout(n746),.clk(gclk));
	jand g0674(.dina(w_dff_B_k4AlFgau3_0),.dinb(n742),.dout(n747),.clk(gclk));
	jand g0675(.dina(w_dff_B_PYzOnq4l7_0),.dinb(n705),.dout(n748),.clk(gclk));
	jnot g0676(.din(n748),.dout(n749),.clk(gclk));
	jand g0677(.dina(n749),.dinb(n702),.dout(n750),.clk(gclk));
	jnot g0678(.din(w_n750_0[1]),.dout(G384_fa_),.clk(gclk));
	jnot g0679(.din(w_n552_1[0]),.dout(n752),.clk(gclk));
	jand g0680(.dina(w_dff_B_Roa0scio0_0),.dinb(w_n542_0[1]),.dout(n753),.clk(gclk));
	jand g0681(.dina(w_n552_0[2]),.dinb(w_n512_0[0]),.dout(n754),.clk(gclk));
	jnot g0682(.din(w_n754_0[1]),.dout(n755),.clk(gclk));
	jand g0683(.dina(n755),.dinb(w_n517_0[0]),.dout(n756),.clk(gclk));
	jand g0684(.dina(w_n754_0[0]),.dinb(w_n542_0[0]),.dout(n757),.clk(gclk));
	jcb g0685(.dina(w_dff_B_crVwk4RA1_0),.dinb(n756),.dout(n758));
	jand g0686(.dina(w_n696_1[0]),.dinb(w_n576_0[2]),.dout(n759),.clk(gclk));
	jand g0687(.dina(w_n553_1[2]),.dinb(w_n436_0[0]),.dout(n760),.clk(gclk));
	jnot g0688(.din(w_n760_0[1]),.dout(n761),.clk(gclk));
	jand g0689(.dina(w_dff_B_CKoaYjSd0_0),.dinb(w_n446_0[0]),.dout(n762),.clk(gclk));
	jand g0690(.dina(w_n760_0[0]),.dinb(w_n439_0[2]),.dout(n763),.clk(gclk));
	jcb g0691(.dina(w_dff_B_0ZIerqGo2_0),.dinb(n762),.dout(n764));
	jand g0692(.dina(w_n764_1[2]),.dinb(w_n759_0[1]),.dout(n765),.clk(gclk));
	jcb g0693(.dina(w_n764_1[1]),.dinb(w_n439_0[1]),.dout(n766));
	jand g0694(.dina(w_n554_1[2]),.dinb(w_n543_0[0]),.dout(n767),.clk(gclk));
	jand g0695(.dina(w_dff_B_LI2DMJ7g8_0),.dinb(n766),.dout(n768),.clk(gclk));
	jcb g0696(.dina(w_dff_B_eQDmSvRQ5_0),.dinb(n765),.dout(n769));
	jand g0697(.dina(w_n769_0[1]),.dinb(w_n758_1[1]),.dout(n770),.clk(gclk));
	jcb g0698(.dina(n770),.dinb(w_dff_B_dSbXADPr8_1),.dout(n771));
	jnot g0699(.din(w_n771_0[2]),.dout(n772),.clk(gclk));
	jand g0700(.dina(w_n576_0[1]),.dinb(w_n519_1[0]),.dout(n773),.clk(gclk));
	jcb g0701(.dina(n773),.dinb(w_n548_0[1]),.dout(n774));
	jand g0702(.dina(w_n764_1[0]),.dinb(w_n696_0[2]),.dout(n775),.clk(gclk));
	jand g0703(.dina(n775),.dinb(w_n758_1[0]),.dout(n776),.clk(gclk));
	jxor g0704(.dina(n776),.dinb(w_n519_0[2]),.dout(n777),.clk(gclk));
	jand g0705(.dina(n777),.dinb(w_n588_0[2]),.dout(n778),.clk(gclk));
	jxor g0706(.dina(n778),.dinb(w_dff_B_7L91uwTL8_1),.dout(n779),.clk(gclk));
	jnot g0707(.din(w_n779_0[1]),.dout(n780),.clk(gclk));
	jcb g0708(.dina(n780),.dinb(n772),.dout(n781));
	jcb g0709(.dina(w_n779_0[0]),.dinb(w_n771_0[1]),.dout(n782));
	jnot g0710(.din(w_n121_0[1]),.dout(n783),.clk(gclk));
	jand g0711(.dina(n783),.dinb(w_n116_0[0]),.dout(n784),.clk(gclk));
	jand g0712(.dina(w_dff_B_viTl6LRz7_0),.dinb(n782),.dout(n785),.clk(gclk));
	jand g0713(.dina(n785),.dinb(n781),.dout(n786),.clk(gclk));
	jand g0714(.dina(w_G77_3[0]),.dinb(w_G50_3[1]),.dout(n787),.clk(gclk));
	jand g0715(.dina(n787),.dinb(w_n137_0[0]),.dout(n788),.clk(gclk));
	jand g0716(.dina(w_G68_3[0]),.dinb(w_n73_1[2]),.dout(n789),.clk(gclk));
	jcb g0717(.dina(n789),.dinb(n788),.dout(n790));
	jand g0718(.dina(n790),.dinb(w_n121_0[0]),.dout(n791),.clk(gclk));
	jnot g0719(.din(w_n255_0[0]),.dout(n792),.clk(gclk));
	jand g0720(.dina(w_n147_0[0]),.dinb(w_G116_3[1]),.dout(n793),.clk(gclk));
	jand g0721(.dina(w_dff_B_YHtyzqau1_0),.dinb(n792),.dout(n794),.clk(gclk));
	jcb g0722(.dina(n794),.dinb(w_dff_B_xSUxJVYv1_1),.dout(n795));
	jcb g0723(.dina(w_dff_B_6r4cWHNH7_0),.dinb(n786),.dout(G367));
	jand g0724(.dina(w_n553_1[1]),.dinb(w_n214_0[0]),.dout(n797),.clk(gclk));
	jnot g0725(.din(w_n797_0[1]),.dout(n798),.clk(gclk));
	jand g0726(.dina(n798),.dinb(w_n219_0[0]),.dout(n799),.clk(gclk));
	jand g0727(.dina(w_n797_0[0]),.dinb(w_n532_0[0]),.dout(n800),.clk(gclk));
	jcb g0728(.dina(w_dff_B_wqUxesZM3_0),.dinb(n799),.dout(n801));
	jnot g0729(.din(w_n801_0[1]),.dout(n802),.clk(gclk));
	jand g0730(.dina(n802),.dinb(w_n608_1[0]),.dout(n803),.clk(gclk));
	jnot g0731(.din(n803),.dout(n804),.clk(gclk));
	jand g0732(.dina(w_n631_6[0]),.dinb(w_G317_1[0]),.dout(n805),.clk(gclk));
	jand g0733(.dina(w_n623_4[1]),.dinb(w_G107_2[2]),.dout(n806),.clk(gclk));
	jand g0734(.dina(w_n642_6[0]),.dinb(w_G294_2[1]),.dout(n807),.clk(gclk));
	jcb g0735(.dina(w_dff_B_epMcabcQ1_0),.dinb(n806),.dout(n808));
	jcb g0736(.dina(n808),.dinb(w_dff_B_jy15bCAb1_1),.dout(n809));
	jand g0737(.dina(w_n617_5[0]),.dinb(w_G116_3[0]),.dout(n810),.clk(gclk));
	jcb g0738(.dina(n810),.dinb(w_n148_4[2]),.dout(n811));
	jand g0739(.dina(w_n636_6[0]),.dinb(w_G283_2[2]),.dout(n812),.clk(gclk));
	jand g0740(.dina(w_n627_6[0]),.dinb(w_G303_1[2]),.dout(n813),.clk(gclk));
	jcb g0741(.dina(n813),.dinb(n812),.dout(n814));
	jand g0742(.dina(w_n640_6[0]),.dinb(w_G311_1[0]),.dout(n815),.clk(gclk));
	jand g0743(.dina(w_n634_3[0]),.dinb(w_G97_3[0]),.dout(n816),.clk(gclk));
	jcb g0744(.dina(w_n816_0[1]),.dinb(w_dff_B_xVasj5kJ8_1),.dout(n817));
	jcb g0745(.dina(n817),.dinb(w_dff_B_KQKiFyKL2_1),.dout(n818));
	jcb g0746(.dina(n818),.dinb(n811),.dout(n819));
	jcb g0747(.dina(n819),.dinb(n809),.dout(n820));
	jand g0748(.dina(w_n631_5[2]),.dinb(w_G137_1[1]),.dout(n821),.clk(gclk));
	jnot g0749(.din(n821),.dout(n822),.clk(gclk));
	jand g0750(.dina(w_n623_4[0]),.dinb(w_G68_2[2]),.dout(n823),.clk(gclk));
	jnot g0751(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jand g0752(.dina(w_n634_2[2]),.dinb(w_G77_2[2]),.dout(n825),.clk(gclk));
	jnot g0753(.din(w_n825_0[1]),.dout(n826),.clk(gclk));
	jand g0754(.dina(n826),.dinb(n824),.dout(n827),.clk(gclk));
	jand g0755(.dina(n827),.dinb(w_dff_B_krmUV8RO2_1),.dout(n828),.clk(gclk));
	jand g0756(.dina(w_n642_5[2]),.dinb(w_G159_2[2]),.dout(n829),.clk(gclk));
	jcb g0757(.dina(n829),.dinb(w_G33_5[1]),.dout(n830));
	jand g0758(.dina(w_n640_5[2]),.dinb(w_G143_2[0]),.dout(n831),.clk(gclk));
	jand g0759(.dina(w_n627_5[2]),.dinb(w_G150_2[2]),.dout(n832),.clk(gclk));
	jcb g0760(.dina(n832),.dinb(n831),.dout(n833));
	jand g0761(.dina(w_n636_5[2]),.dinb(w_G50_3[0]),.dout(n834),.clk(gclk));
	jand g0762(.dina(w_n617_4[2]),.dinb(w_G58_3[0]),.dout(n835),.clk(gclk));
	jcb g0763(.dina(n835),.dinb(w_dff_B_MvjyWkCQ5_1),.dout(n836));
	jcb g0764(.dina(n836),.dinb(w_dff_B_V844WwYT9_1),.dout(n837));
	jcb g0765(.dina(n837),.dinb(w_dff_B_5S32BAId0_1),.dout(n838));
	jnot g0766(.din(n838),.dout(n839),.clk(gclk));
	jand g0767(.dina(w_dff_B_hlJjD9Rg6_0),.dinb(n828),.dout(n840),.clk(gclk));
	jnot g0768(.din(n840),.dout(n841),.clk(gclk));
	jand g0769(.dina(n841),.dinb(w_dff_B_k9MMBBPr6_1),.dout(n842),.clk(gclk));
	jcb g0770(.dina(n842),.dinb(w_n612_3[0]),.dout(n843));
	jand g0771(.dina(w_n675_0[1]),.dinb(w_n131_0[0]),.dout(n844),.clk(gclk));
	jand g0772(.dina(w_n123_1[0]),.dinb(w_G87_1[2]),.dout(n845),.clk(gclk));
	jcb g0773(.dina(w_dff_B_VKqW2bGp3_0),.dinb(w_n672_1[0]),.dout(n846));
	jcb g0774(.dina(n846),.dinb(w_dff_B_yS816wcL4_1),.dout(n847));
	jand g0775(.dina(n847),.dinb(w_n604_1[1]),.dout(n848),.clk(gclk));
	jand g0776(.dina(w_dff_B_2Etd3YNq0_0),.dinb(n843),.dout(n849),.clk(gclk));
	jand g0777(.dina(w_dff_B_CipYhRss3_0),.dinb(n804),.dout(n850),.clk(gclk));
	jnot g0778(.din(w_n589_1[1]),.dout(n851),.clk(gclk));
	jxor g0779(.dina(w_n561_0[0]),.dinb(w_n556_0[0]),.dout(n852),.clk(gclk));
	jxor g0780(.dina(n852),.dinb(w_n572_0[0]),.dout(n853),.clk(gclk));
	jnot g0781(.din(w_n853_0[2]),.dout(n854),.clk(gclk));
	jand g0782(.dina(w_dff_B_Yvw3WQHh8_0),.dinb(n851),.dout(n855),.clk(gclk));
	jnot g0783(.din(w_n278_0[0]),.dout(n856),.clk(gclk));
	jand g0784(.dina(w_n553_1[0]),.dinb(w_n274_0[0]),.dout(n857),.clk(gclk));
	jcb g0785(.dina(w_dff_B_K9CLbvgv0_0),.dinb(n856),.dout(n858));
	jand g0786(.dina(w_n553_0[2]),.dinb(w_n536_0[1]),.dout(n859),.clk(gclk));
	jnot g0787(.din(n859),.dout(n860),.clk(gclk));
	jand g0788(.dina(n860),.dinb(n858),.dout(n861),.clk(gclk));
	jxor g0789(.dina(w_n861_1[1]),.dinb(w_n573_0[1]),.dout(n862),.clk(gclk));
	jxor g0790(.dina(n862),.dinb(w_n563_0[1]),.dout(n863),.clk(gclk));
	jand g0791(.dina(w_n863_0[1]),.dinb(w_n855_0[2]),.dout(n864),.clk(gclk));
	jcb g0792(.dina(w_n864_0[1]),.dinb(w_n589_1[0]),.dout(n865));
	jand g0793(.dina(n865),.dinb(w_n591_0[2]),.dout(n866),.clk(gclk));
	jcb g0794(.dina(n866),.dinb(w_n602_0[0]),.dout(n867));
	jand g0795(.dina(w_n554_1[1]),.dinb(w_n536_0[0]),.dout(n868),.clk(gclk));
	jnot g0796(.din(w_n861_1[0]),.dout(n869),.clk(gclk));
	jand g0797(.dina(n869),.dinb(w_n563_0[0]),.dout(n870),.clk(gclk));
	jcb g0798(.dina(n870),.dinb(w_dff_B_0L24BZH86_1),.dout(n871));
	jcb g0799(.dina(w_n861_0[2]),.dinb(w_n573_0[0]),.dout(n872));
	jxor g0800(.dina(w_dff_B_BUE8W33A7_0),.dinb(w_n801_0[0]),.dout(n873),.clk(gclk));
	jxor g0801(.dina(n873),.dinb(n871),.dout(n874),.clk(gclk));
	jnot g0802(.din(n874),.dout(n875),.clk(gclk));
	jand g0803(.dina(w_dff_B_xo4Jgk4M3_0),.dinb(n867),.dout(n876),.clk(gclk));
	jcb g0804(.dina(n876),.dinb(w_dff_B_VmrBYFvk2_1),.dout(G387_fa_));
	jand g0805(.dina(w_n853_0[1]),.dinb(w_n589_0[2]),.dout(n878),.clk(gclk));
	jcb g0806(.dina(w_n855_0[1]),.dinb(w_n592_1[2]),.dout(n879));
	jcb g0807(.dina(n879),.dinb(w_dff_B_CU5aFT977_1),.dout(n880));
	jcb g0808(.dina(w_n853_0[0]),.dinb(w_n603_2[0]),.dout(n881));
	jand g0809(.dina(w_n608_0[2]),.dinb(w_n564_0[0]),.dout(n882),.clk(gclk));
	jand g0810(.dina(w_n631_5[1]),.dinb(w_G326_0[0]),.dout(n883),.clk(gclk));
	jand g0811(.dina(w_n623_3[2]),.dinb(w_G283_2[1]),.dout(n884),.clk(gclk));
	jand g0812(.dina(w_n627_5[1]),.dinb(w_G317_0[2]),.dout(n885),.clk(gclk));
	jcb g0813(.dina(w_dff_B_ViLt7ylH0_0),.dinb(n884),.dout(n886));
	jcb g0814(.dina(n886),.dinb(w_dff_B_p66zbhX35_1),.dout(n887));
	jand g0815(.dina(w_n617_4[1]),.dinb(w_G294_2[0]),.dout(n888),.clk(gclk));
	jcb g0816(.dina(n888),.dinb(w_n148_4[1]),.dout(n889));
	jand g0817(.dina(w_n634_2[1]),.dinb(w_G116_2[2]),.dout(n890),.clk(gclk));
	jand g0818(.dina(w_n636_5[1]),.dinb(w_G303_1[1]),.dout(n891),.clk(gclk));
	jcb g0819(.dina(w_dff_B_rQOiTh2F7_0),.dinb(n890),.dout(n892));
	jand g0820(.dina(w_n640_5[1]),.dinb(w_G322_0[1]),.dout(n893),.clk(gclk));
	jand g0821(.dina(w_n642_5[1]),.dinb(w_G311_0[2]),.dout(n894),.clk(gclk));
	jcb g0822(.dina(n894),.dinb(n893),.dout(n895));
	jcb g0823(.dina(w_dff_B_hU0nysu46_0),.dinb(n892),.dout(n896));
	jcb g0824(.dina(n896),.dinb(n889),.dout(n897));
	jcb g0825(.dina(n897),.dinb(n887),.dout(n898));
	jand g0826(.dina(w_n623_3[1]),.dinb(w_G87_1[1]),.dout(n899),.clk(gclk));
	jand g0827(.dina(w_n642_5[0]),.dinb(w_G58_2[2]),.dout(n900),.clk(gclk));
	jcb g0828(.dina(w_dff_B_QA35yFD00_0),.dinb(w_n816_0[0]),.dout(n901));
	jcb g0829(.dina(n901),.dinb(w_n899_0[1]),.dout(n902));
	jand g0830(.dina(w_n631_5[0]),.dinb(w_G150_2[1]),.dout(n903),.clk(gclk));
	jcb g0831(.dina(n903),.dinb(w_G33_5[0]),.dout(n904));
	jand g0832(.dina(w_n640_5[0]),.dinb(w_G159_2[1]),.dout(n905),.clk(gclk));
	jand g0833(.dina(w_n636_5[0]),.dinb(w_G68_2[1]),.dout(n906),.clk(gclk));
	jcb g0834(.dina(n906),.dinb(n905),.dout(n907));
	jand g0835(.dina(w_n627_5[0]),.dinb(w_G50_2[2]),.dout(n908),.clk(gclk));
	jand g0836(.dina(w_n617_4[0]),.dinb(w_G77_2[1]),.dout(n909),.clk(gclk));
	jcb g0837(.dina(w_n909_0[1]),.dinb(w_dff_B_8NAA6ogq4_1),.dout(n910));
	jcb g0838(.dina(n910),.dinb(w_dff_B_Ve7dusDi5_1),.dout(n911));
	jcb g0839(.dina(n911),.dinb(w_dff_B_5KLB4HMo4_1),.dout(n912));
	jcb g0840(.dina(n912),.dinb(n902),.dout(n913));
	jand g0841(.dina(n913),.dinb(n898),.dout(n914),.clk(gclk));
	jcb g0842(.dina(n914),.dinb(w_n612_2[2]),.dout(n915));
	jand g0843(.dina(w_n135_0[0]),.dinb(w_G45_0[1]),.dout(n916),.clk(gclk));
	jand g0844(.dina(w_G77_2[0]),.dinb(w_G68_2[0]),.dout(n917),.clk(gclk));
	jnot g0845(.din(n917),.dout(n918),.clk(gclk));
	jand g0846(.dina(w_G58_2[1]),.dinb(w_n161_0[1]),.dout(n919),.clk(gclk));
	jand g0847(.dina(n919),.dinb(w_n73_1[1]),.dout(n920),.clk(gclk));
	jand g0848(.dina(n920),.dinb(w_dff_B_vHxeNTmt0_1),.dout(n921),.clk(gclk));
	jand g0849(.dina(n921),.dinb(w_n593_0[1]),.dout(n922),.clk(gclk));
	jcb g0850(.dina(n922),.dinb(w_n676_0[0]),.dout(n923));
	jcb g0851(.dina(n923),.dinb(w_dff_B_PrT57hO05_1),.dout(n924));
	jand g0852(.dina(w_n123_0[2]),.dinb(w_n80_0[1]),.dout(n925),.clk(gclk));
	jnot g0853(.din(w_n593_0[0]),.dout(n926),.clk(gclk));
	jand g0854(.dina(w_n680_0[0]),.dinb(n926),.dout(n927),.clk(gclk));
	jcb g0855(.dina(n927),.dinb(w_dff_B_8VZ402Ky1_1),.dout(n928));
	jnot g0856(.din(n928),.dout(n929),.clk(gclk));
	jand g0857(.dina(n929),.dinb(w_dff_B_c5054Njd6_1),.dout(n930),.clk(gclk));
	jcb g0858(.dina(n930),.dinb(w_n672_0[2]),.dout(n931));
	jand g0859(.dina(n931),.dinb(w_n604_1[0]),.dout(n932),.clk(gclk));
	jand g0860(.dina(n932),.dinb(w_dff_B_iDRMvkcQ1_1),.dout(n933),.clk(gclk));
	jnot g0861(.din(n933),.dout(n934),.clk(gclk));
	jcb g0862(.dina(n934),.dinb(n882),.dout(n935));
	jand g0863(.dina(n935),.dinb(n881),.dout(n936),.clk(gclk));
	jand g0864(.dina(w_dff_B_YRi0c8Xj3_0),.dinb(n880),.dout(n937),.clk(gclk));
	jnot g0865(.din(w_n937_0[2]),.dout(G393),.clk(gclk));
	jnot g0866(.din(w_n855_0[0]),.dout(n939),.clk(gclk));
	jnot g0867(.din(w_n863_0[0]),.dout(n940),.clk(gclk));
	jand g0868(.dina(w_n940_0[1]),.dinb(n939),.dout(n941),.clk(gclk));
	jcb g0869(.dina(w_n864_0[0]),.dinb(w_n592_1[1]),.dout(n942));
	jcb g0870(.dina(w_dff_B_MtzuOHMI5_0),.dinb(n941),.dout(n943));
	jcb g0871(.dina(w_n940_0[0]),.dinb(w_n603_1[2]),.dout(n944));
	jand g0872(.dina(w_n861_0[1]),.dinb(w_n608_0[1]),.dout(n945),.clk(gclk));
	jnot g0873(.din(n945),.dout(n946),.clk(gclk));
	jand g0874(.dina(w_n623_3[0]),.dinb(w_G116_2[1]),.dout(n947),.clk(gclk));
	jand g0875(.dina(w_n617_3[2]),.dinb(w_G283_2[0]),.dout(n948),.clk(gclk));
	jand g0876(.dina(w_n642_4[2]),.dinb(w_G303_1[0]),.dout(n949),.clk(gclk));
	jcb g0877(.dina(w_dff_B_OGdqf51U6_0),.dinb(n948),.dout(n950));
	jcb g0878(.dina(n950),.dinb(n947),.dout(n951));
	jand g0879(.dina(w_n631_4[2]),.dinb(w_G322_0[0]),.dout(n952),.clk(gclk));
	jcb g0880(.dina(n952),.dinb(w_n148_4[0]),.dout(n953));
	jand g0881(.dina(w_n636_4[2]),.dinb(w_G294_1[2]),.dout(n954),.clk(gclk));
	jand g0882(.dina(w_n627_4[2]),.dinb(w_G311_0[1]),.dout(n955),.clk(gclk));
	jcb g0883(.dina(n955),.dinb(n954),.dout(n956));
	jand g0884(.dina(w_n640_4[2]),.dinb(w_G317_0[1]),.dout(n957),.clk(gclk));
	jcb g0885(.dina(w_dff_B_V6mBJiHs9_0),.dinb(w_n657_0[0]),.dout(n958));
	jcb g0886(.dina(n958),.dinb(w_dff_B_u811M5jM0_1),.dout(n959));
	jcb g0887(.dina(n959),.dinb(w_dff_B_NKahejBj1_1),.dout(n960));
	jcb g0888(.dina(n960),.dinb(n951),.dout(n961));
	jand g0889(.dina(w_n623_2[2]),.dinb(w_G77_1[2]),.dout(n962),.clk(gclk));
	jand g0890(.dina(w_n617_3[1]),.dinb(w_G68_1[2]),.dout(n963),.clk(gclk));
	jand g0891(.dina(w_n642_4[1]),.dinb(w_G50_2[1]),.dout(n964),.clk(gclk));
	jcb g0892(.dina(w_dff_B_yW3zibOM5_0),.dinb(n963),.dout(n965));
	jcb g0893(.dina(n965),.dinb(w_n962_0[1]),.dout(n966));
	jand g0894(.dina(w_n631_4[1]),.dinb(w_G143_1[2]),.dout(n967),.clk(gclk));
	jcb g0895(.dina(n967),.dinb(w_G33_4[2]),.dout(n968));
	jand g0896(.dina(w_n636_4[1]),.dinb(w_G58_2[0]),.dout(n969),.clk(gclk));
	jand g0897(.dina(w_n627_4[1]),.dinb(w_G159_2[0]),.dout(n970),.clk(gclk));
	jcb g0898(.dina(n970),.dinb(n969),.dout(n971));
	jand g0899(.dina(w_n640_4[1]),.dinb(w_G150_2[0]),.dout(n972),.clk(gclk));
	jcb g0900(.dina(w_dff_B_t7y68eUg3_0),.dinb(w_n728_0[0]),.dout(n973));
	jcb g0901(.dina(n973),.dinb(w_dff_B_bBjhKhHV1_1),.dout(n974));
	jcb g0902(.dina(n974),.dinb(w_dff_B_QTK8jM607_1),.dout(n975));
	jcb g0903(.dina(n975),.dinb(n966),.dout(n976));
	jand g0904(.dina(n976),.dinb(n961),.dout(n977),.clk(gclk));
	jcb g0905(.dina(n977),.dinb(w_n612_2[1]),.dout(n978));
	jand g0906(.dina(w_n675_0[0]),.dinb(w_n144_0[0]),.dout(n979),.clk(gclk));
	jand g0907(.dina(w_n123_0[1]),.dinb(w_G97_2[2]),.dout(n980),.clk(gclk));
	jcb g0908(.dina(w_dff_B_CsuIWoK75_0),.dinb(w_n672_0[1]),.dout(n981));
	jcb g0909(.dina(n981),.dinb(w_dff_B_EeBQm7hU3_1),.dout(n982));
	jand g0910(.dina(n982),.dinb(w_n604_0[2]),.dout(n983),.clk(gclk));
	jand g0911(.dina(n983),.dinb(w_dff_B_et0EBgT21_1),.dout(n984),.clk(gclk));
	jand g0912(.dina(w_dff_B_xeCC2MJU7_0),.dinb(n946),.dout(n985),.clk(gclk));
	jnot g0913(.din(n985),.dout(n986),.clk(gclk));
	jand g0914(.dina(n986),.dinb(w_dff_B_J4fxFNtS0_1),.dout(n987),.clk(gclk));
	jand g0915(.dina(w_dff_B_6LfJIXbT7_0),.dinb(n943),.dout(n988),.clk(gclk));
	jnot g0916(.din(w_n988_0[2]),.dout(G390),.clk(gclk));
	jnot g0917(.din(w_n758_0[2]),.dout(n990),.clk(gclk));
	jand g0918(.dina(w_n696_0[1]),.dinb(w_n588_0[1]),.dout(n991),.clk(gclk));
	jand g0919(.dina(w_n991_0[1]),.dinb(w_n764_0[2]),.dout(n992),.clk(gclk));
	jxor g0920(.dina(w_n992_0[1]),.dinb(w_n990_0[1]),.dout(n993),.clk(gclk));
	jxor g0921(.dina(n993),.dinb(w_n769_0[0]),.dout(n994),.clk(gclk));
	jand g0922(.dina(w_n589_0[1]),.dinb(w_n519_0[1]),.dout(n995),.clk(gclk));
	jcb g0923(.dina(n995),.dinb(w_n548_0[0]),.dout(n996));
	jand g0924(.dina(w_n554_1[0]),.dinb(w_n404_0[0]),.dout(n997),.clk(gclk));
	jcb g0925(.dina(w_dff_B_JCQfpg1X7_0),.dinb(w_n759_0[0]),.dout(n998));
	jnot g0926(.din(w_n764_0[1]),.dout(n999),.clk(gclk));
	jxor g0927(.dina(w_n991_0[0]),.dinb(w_n999_0[1]),.dout(n1000),.clk(gclk));
	jxor g0928(.dina(n1000),.dinb(w_dff_B_gbC0DPc77_1),.dout(n1001),.clk(gclk));
	jcb g0929(.dina(w_n1001_0[2]),.dinb(w_n996_0[2]),.dout(n1002));
	jcb g0930(.dina(w_n1002_0[2]),.dinb(w_n994_0[2]),.dout(n1003));
	jnot g0931(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jand g0932(.dina(w_n1002_0[1]),.dinb(w_n994_0[1]),.dout(n1005),.clk(gclk));
	jcb g0933(.dina(n1005),.dinb(w_n592_1[0]),.dout(n1006));
	jcb g0934(.dina(n1006),.dinb(n1004),.dout(n1007));
	jcb g0935(.dina(w_n994_0[0]),.dinb(w_n603_1[1]),.dout(n1008));
	jand g0936(.dina(w_n990_0[0]),.dinb(w_n425_1[0]),.dout(n1009),.clk(gclk));
	jnot g0937(.din(n1009),.dout(n1010),.clk(gclk));
	jand g0938(.dina(w_n631_4[0]),.dinb(w_G125_0[1]),.dout(n1011),.clk(gclk));
	jand g0939(.dina(w_n623_2[1]),.dinb(w_G159_1[2]),.dout(n1012),.clk(gclk));
	jand g0940(.dina(w_n642_4[0]),.dinb(w_G137_1[0]),.dout(n1013),.clk(gclk));
	jcb g0941(.dina(w_dff_B_wvhPnYKL8_0),.dinb(n1012),.dout(n1014));
	jcb g0942(.dina(n1014),.dinb(w_dff_B_LdT9P7kQ6_1),.dout(n1015));
	jand g0943(.dina(w_n617_3[0]),.dinb(w_G150_1[2]),.dout(n1016),.clk(gclk));
	jcb g0944(.dina(n1016),.dinb(w_G33_4[1]),.dout(n1017));
	jand g0945(.dina(w_n636_4[0]),.dinb(w_G143_1[1]),.dout(n1018),.clk(gclk));
	jand g0946(.dina(w_n627_4[0]),.dinb(w_G132_1[0]),.dout(n1019),.clk(gclk));
	jcb g0947(.dina(n1019),.dinb(n1018),.dout(n1020));
	jand g0948(.dina(w_n640_4[0]),.dinb(w_G128_0[2]),.dout(n1021),.clk(gclk));
	jand g0949(.dina(w_n634_2[0]),.dinb(w_G50_2[0]),.dout(n1022),.clk(gclk));
	jcb g0950(.dina(n1022),.dinb(w_dff_B_T6FbOtID0_1),.dout(n1023));
	jcb g0951(.dina(n1023),.dinb(w_dff_B_kikptGj60_1),.dout(n1024));
	jcb g0952(.dina(n1024),.dinb(n1017),.dout(n1025));
	jcb g0953(.dina(n1025),.dinb(n1015),.dout(n1026));
	jand g0954(.dina(w_n631_3[2]),.dinb(w_G294_1[1]),.dout(n1027),.clk(gclk));
	jand g0955(.dina(w_n642_3[2]),.dinb(w_G107_2[1]),.dout(n1028),.clk(gclk));
	jcb g0956(.dina(w_dff_B_rJw8V6fi8_0),.dinb(w_n962_0[0]),.dout(n1029));
	jcb g0957(.dina(n1029),.dinb(w_dff_B_bGx2WRnA7_1),.dout(n1030));
	jand g0958(.dina(w_n640_3[2]),.dinb(w_G283_1[2]),.dout(n1031),.clk(gclk));
	jcb g0959(.dina(n1031),.dinb(w_n148_3[2]),.dout(n1032));
	jand g0960(.dina(w_n636_3[2]),.dinb(w_G97_2[1]),.dout(n1033),.clk(gclk));
	jand g0961(.dina(w_n627_3[2]),.dinb(w_G116_2[0]),.dout(n1034),.clk(gclk));
	jcb g0962(.dina(n1034),.dinb(n1033),.dout(n1035));
	jcb g0963(.dina(w_n717_0[0]),.dinb(w_n654_0[0]),.dout(n1036));
	jcb g0964(.dina(n1036),.dinb(w_dff_B_4HVNIoJw8_1),.dout(n1037));
	jcb g0965(.dina(n1037),.dinb(w_dff_B_Bj8BiRrI3_1),.dout(n1038));
	jcb g0966(.dina(n1038),.dinb(n1030),.dout(n1039));
	jand g0967(.dina(n1039),.dinb(n1026),.dout(n1040),.clk(gclk));
	jcb g0968(.dina(n1040),.dinb(w_n612_2[0]),.dout(n1041));
	jand g0969(.dina(w_n743_1[0]),.dinb(w_n74_0[1]),.dout(n1042),.clk(gclk));
	jcb g0970(.dina(w_dff_B_RTO9is4E1_0),.dinb(w_n605_1[0]),.dout(n1043));
	jnot g0971(.din(n1043),.dout(n1044),.clk(gclk));
	jand g0972(.dina(n1044),.dinb(w_dff_B_u0QRMWvq1_1),.dout(n1045),.clk(gclk));
	jand g0973(.dina(w_dff_B_legx5ooM3_0),.dinb(n1010),.dout(n1046),.clk(gclk));
	jnot g0974(.din(n1046),.dout(n1047),.clk(gclk));
	jand g0975(.dina(n1047),.dinb(n1008),.dout(n1048),.clk(gclk));
	jand g0976(.dina(n1048),.dinb(n1007),.dout(n1049),.clk(gclk));
	jnot g0977(.din(w_n1049_0[2]),.dout(G378),.clk(gclk));
	jand g0978(.dina(w_n992_0[0]),.dinb(w_n758_0[1]),.dout(n1051),.clk(gclk));
	jand g0979(.dina(w_n552_0[1]),.dinb(w_n479_0[0]),.dout(n1052),.clk(gclk));
	jnot g0980(.din(w_n1052_0[1]),.dout(n1053),.clk(gclk));
	jand g0981(.dina(n1053),.dinb(w_n484_0[0]),.dout(n1054),.clk(gclk));
	jand g0982(.dina(w_n1052_0[0]),.dinb(w_n541_0[0]),.dout(n1055),.clk(gclk));
	jcb g0983(.dina(w_dff_B_u0fVKxXR3_0),.dinb(n1054),.dout(n1056));
	jnot g0984(.din(n1056),.dout(n1057),.clk(gclk));
	jxor g0985(.dina(w_n1057_0[1]),.dinb(w_n771_0[0]),.dout(n1058),.clk(gclk));
	jxor g0986(.dina(n1058),.dinb(w_dff_B_IhGxUNJH0_1),.dout(n1059),.clk(gclk));
	jcb g0987(.dina(w_n1059_0[1]),.dinb(w_n603_1[0]),.dout(n1060));
	jnot g0988(.din(w_n996_0[1]),.dout(n1061),.clk(gclk));
	jand g0989(.dina(w_n1003_0[0]),.dinb(w_dff_B_dmMFLBrb2_1),.dout(n1062),.clk(gclk));
	jcb g0990(.dina(n1062),.dinb(w_n592_0[2]),.dout(n1063));
	jcb g0991(.dina(n1063),.dinb(w_n1059_0[0]),.dout(n1064));
	jand g0992(.dina(w_n1057_0[0]),.dinb(w_n425_0[2]),.dout(n1065),.clk(gclk));
	jnot g0993(.din(w_n612_1[2]),.dout(n1066),.clk(gclk));
	jand g0994(.dina(w_n642_3[1]),.dinb(w_G132_0[2]),.dout(n1067),.clk(gclk));
	jand g0995(.dina(w_n627_3[1]),.dinb(w_G128_0[1]),.dout(n1068),.clk(gclk));
	jand g0996(.dina(w_n636_3[1]),.dinb(w_G137_0[2]),.dout(n1069),.clk(gclk));
	jcb g0997(.dina(n1069),.dinb(n1068),.dout(n1070));
	jcb g0998(.dina(n1070),.dinb(n1067),.dout(n1071));
	jnot g0999(.din(n1071),.dout(n1072),.clk(gclk));
	jand g1000(.dina(w_n623_2[0]),.dinb(w_G150_1[1]),.dout(n1073),.clk(gclk));
	jnot g1001(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1002(.dina(w_n149_1[0]),.dinb(w_n148_3[1]),.dout(n1075),.clk(gclk));
	jand g1003(.dina(w_dff_B_B7rMKbCp5_0),.dinb(n1074),.dout(n1076),.clk(gclk));
	jand g1004(.dina(w_n640_3[1]),.dinb(w_G125_0[0]),.dout(n1077),.clk(gclk));
	jand g1005(.dina(w_n617_2[2]),.dinb(w_G143_1[0]),.dout(n1078),.clk(gclk));
	jcb g1006(.dina(n1078),.dinb(w_dff_B_V4onKTSI5_1),.dout(n1079));
	jand g1007(.dina(w_n631_3[1]),.dinb(w_dff_B_4JQUvYtX3_1),.dout(n1080),.clk(gclk));
	jand g1008(.dina(w_n634_1[2]),.dinb(w_G159_1[1]),.dout(n1081),.clk(gclk));
	jcb g1009(.dina(n1081),.dinb(w_dff_B_lo148zU95_1),.dout(n1082));
	jcb g1010(.dina(n1082),.dinb(n1079),.dout(n1083));
	jnot g1011(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1012(.dina(w_dff_B_DJYD2Cpt1_0),.dinb(n1076),.dout(n1085),.clk(gclk));
	jand g1013(.dina(n1085),.dinb(w_dff_B_jYnSfBdI6_1),.dout(n1086),.clk(gclk));
	jand g1014(.dina(w_n627_3[0]),.dinb(w_G107_2[0]),.dout(n1087),.clk(gclk));
	jand g1015(.dina(w_n634_1[1]),.dinb(w_G58_1[2]),.dout(n1088),.clk(gclk));
	jand g1016(.dina(w_n636_3[0]),.dinb(w_G87_1[0]),.dout(n1089),.clk(gclk));
	jcb g1017(.dina(w_dff_B_mjJCM2hf6_0),.dinb(w_n1088_0[1]),.dout(n1090));
	jcb g1018(.dina(n1090),.dinb(w_dff_B_RXABdTP05_1),.dout(n1091));
	jnot g1019(.din(n1091),.dout(n1092),.clk(gclk));
	jand g1020(.dina(w_n642_3[0]),.dinb(w_G97_2[0]),.dout(n1093),.clk(gclk));
	jnot g1021(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1022(.dina(w_n149_0[2]),.dinb(w_G33_4[0]),.dout(n1095),.clk(gclk));
	jand g1023(.dina(w_dff_B_7MFYz6Q68_0),.dinb(n1094),.dout(n1096),.clk(gclk));
	jand g1024(.dina(w_n631_3[0]),.dinb(w_G283_1[1]),.dout(n1097),.clk(gclk));
	jcb g1025(.dina(w_dff_B_OqWtzlI70_0),.dinb(w_n823_0[0]),.dout(n1098));
	jand g1026(.dina(w_n640_3[0]),.dinb(w_G116_1[2]),.dout(n1099),.clk(gclk));
	jcb g1027(.dina(w_dff_B_qZohO1Mp1_0),.dinb(w_n909_0[0]),.dout(n1100));
	jcb g1028(.dina(n1100),.dinb(n1098),.dout(n1101));
	jnot g1029(.din(n1101),.dout(n1102),.clk(gclk));
	jand g1030(.dina(n1102),.dinb(n1096),.dout(n1103),.clk(gclk));
	jand g1031(.dina(n1103),.dinb(w_dff_B_4zeUQeoC6_1),.dout(n1104),.clk(gclk));
	jand g1032(.dina(w_n73_1[0]),.dinb(w_G41_0[1]),.dout(n1105),.clk(gclk));
	jcb g1033(.dina(w_dff_B_ppXrUYdm2_0),.dinb(n1104),.dout(n1106));
	jcb g1034(.dina(w_dff_B_o4aZeyj90_0),.dinb(n1086),.dout(n1107));
	jand g1035(.dina(n1107),.dinb(w_dff_B_B3dkUnZH3_1),.dout(n1108),.clk(gclk));
	jand g1036(.dina(w_n743_0[2]),.dinb(w_n73_0[2]),.dout(n1109),.clk(gclk));
	jcb g1037(.dina(w_dff_B_nFMmOQw68_0),.dinb(w_n605_0[2]),.dout(n1110));
	jcb g1038(.dina(w_dff_B_tApKYSbX2_0),.dinb(n1108),.dout(n1111));
	jcb g1039(.dina(w_dff_B_DGak4m8X4_0),.dinb(n1065),.dout(n1112));
	jand g1040(.dina(w_dff_B_dPVwk9Ay5_0),.dinb(n1064),.dout(n1113),.clk(gclk));
	jand g1041(.dina(n1113),.dinb(w_dff_B_WGEwa6yO8_1),.dout(n1114),.clk(gclk));
	jnot g1042(.din(w_n1114_0[2]),.dout(G375),.clk(gclk));
	jand g1043(.dina(w_n1001_0[1]),.dinb(w_n996_0[0]),.dout(n1116),.clk(gclk));
	jnot g1044(.din(n1116),.dout(n1117),.clk(gclk));
	jand g1045(.dina(w_n1002_0[0]),.dinb(w_n591_0[1]),.dout(n1118),.clk(gclk));
	jand g1046(.dina(w_dff_B_gY9f2nnX4_0),.dinb(n1117),.dout(n1119),.clk(gclk));
	jnot g1047(.din(n1119),.dout(n1120),.clk(gclk));
	jcb g1048(.dina(w_n1001_0[0]),.dinb(w_n603_0[2]),.dout(n1121));
	jand g1049(.dina(w_n999_0[0]),.dinb(w_n425_0[1]),.dout(n1122),.clk(gclk));
	jnot g1050(.din(n1122),.dout(n1123),.clk(gclk));
	jand g1051(.dina(w_n623_1[2]),.dinb(w_G50_1[2]),.dout(n1124),.clk(gclk));
	jand g1052(.dina(w_n617_2[1]),.dinb(w_G159_1[0]),.dout(n1125),.clk(gclk));
	jand g1053(.dina(w_n642_2[2]),.dinb(w_G143_0[2]),.dout(n1126),.clk(gclk));
	jcb g1054(.dina(w_dff_B_bC9jIfkQ7_0),.dinb(n1125),.dout(n1127));
	jcb g1055(.dina(n1127),.dinb(n1124),.dout(n1128));
	jand g1056(.dina(w_n631_2[2]),.dinb(w_G128_0[0]),.dout(n1129),.clk(gclk));
	jcb g1057(.dina(n1129),.dinb(w_G33_3[2]),.dout(n1130));
	jand g1058(.dina(w_n636_2[2]),.dinb(w_G150_1[0]),.dout(n1131),.clk(gclk));
	jand g1059(.dina(w_n627_2[2]),.dinb(w_G137_0[1]),.dout(n1132),.clk(gclk));
	jcb g1060(.dina(n1132),.dinb(n1131),.dout(n1133));
	jand g1061(.dina(w_n640_2[2]),.dinb(w_G132_0[1]),.dout(n1134),.clk(gclk));
	jcb g1062(.dina(w_dff_B_IdjcOSiq5_0),.dinb(w_n1088_0[0]),.dout(n1135));
	jcb g1063(.dina(n1135),.dinb(w_dff_B_Q1qvxK2L3_1),.dout(n1136));
	jcb g1064(.dina(n1136),.dinb(w_dff_B_sOcuBiPH3_1),.dout(n1137));
	jcb g1065(.dina(n1137),.dinb(n1128),.dout(n1138));
	jand g1066(.dina(w_n617_2[0]),.dinb(w_G97_1[2]),.dout(n1139),.clk(gclk));
	jand g1067(.dina(w_n640_2[1]),.dinb(w_G294_1[0]),.dout(n1140),.clk(gclk));
	jand g1068(.dina(w_n642_2[1]),.dinb(w_G116_1[1]),.dout(n1141),.clk(gclk));
	jcb g1069(.dina(n1141),.dinb(n1140),.dout(n1142));
	jcb g1070(.dina(w_dff_B_DktmHrQx5_0),.dinb(n1139),.dout(n1143));
	jand g1071(.dina(w_n631_2[1]),.dinb(w_G303_0[2]),.dout(n1144),.clk(gclk));
	jcb g1072(.dina(n1144),.dinb(w_n148_3[0]),.dout(n1145));
	jand g1073(.dina(w_n636_2[1]),.dinb(w_G107_1[2]),.dout(n1146),.clk(gclk));
	jand g1074(.dina(w_n627_2[1]),.dinb(w_G283_1[0]),.dout(n1147),.clk(gclk));
	jcb g1075(.dina(n1147),.dinb(n1146),.dout(n1148));
	jcb g1076(.dina(w_n899_0[0]),.dinb(w_n825_0[0]),.dout(n1149));
	jcb g1077(.dina(n1149),.dinb(w_dff_B_uRqsTUXW5_1),.dout(n1150));
	jcb g1078(.dina(n1150),.dinb(w_dff_B_0E64AsKd0_1),.dout(n1151));
	jcb g1079(.dina(n1151),.dinb(n1143),.dout(n1152));
	jand g1080(.dina(n1152),.dinb(n1138),.dout(n1153),.clk(gclk));
	jcb g1081(.dina(n1153),.dinb(w_n612_1[1]),.dout(n1154));
	jand g1082(.dina(w_n743_0[1]),.dinb(w_n75_0[1]),.dout(n1155),.clk(gclk));
	jcb g1083(.dina(w_dff_B_eRCI9hCc9_0),.dinb(w_n605_0[1]),.dout(n1156));
	jnot g1084(.din(n1156),.dout(n1157),.clk(gclk));
	jand g1085(.dina(n1157),.dinb(w_dff_B_SAV4Uvhx7_1),.dout(n1158),.clk(gclk));
	jand g1086(.dina(w_dff_B_b4TGWIg46_0),.dinb(n1123),.dout(n1159),.clk(gclk));
	jnot g1087(.din(n1159),.dout(n1160),.clk(gclk));
	jand g1088(.dina(n1160),.dinb(n1121),.dout(n1161),.clk(gclk));
	jand g1089(.dina(w_dff_B_b1pGu6vw9_0),.dinb(n1120),.dout(n1162),.clk(gclk));
	jnot g1090(.din(w_n1162_0[2]),.dout(G381),.clk(gclk));
	jand g1091(.dina(w_n1114_0[1]),.dinb(w_n1049_0[1]),.dout(n1164),.clk(gclk));
	jnot g1092(.din(w_G387_0[1]),.dout(n1165),.clk(gclk));
	jnot g1093(.din(w_G396_0[1]),.dout(n1166),.clk(gclk));
	jand g1094(.dina(w_n937_0[1]),.dinb(w_dff_B_dFQcz4hf7_1),.dout(n1167),.clk(gclk));
	jand g1095(.dina(n1167),.dinb(w_n750_0[0]),.dout(n1168),.clk(gclk));
	jand g1096(.dina(n1168),.dinb(w_n988_0[1]),.dout(n1169),.clk(gclk));
	jand g1097(.dina(w_dff_B_qDjqAWub7_0),.dinb(w_n1162_0[1]),.dout(n1170),.clk(gclk));
	jand g1098(.dina(n1170),.dinb(w_dff_B_zYBwZ9ov3_1),.dout(n1171),.clk(gclk));
	jand g1099(.dina(n1171),.dinb(w_n1164_0[1]),.dout(n1172),.clk(gclk));
	jnot g1100(.din(w_n1172_0[1]),.dout(G407),.clk(gclk));
	jnot g1101(.din(w_G213_0[1]),.dout(n1174),.clk(gclk));
	jnot g1102(.din(w_G343_0[0]),.dout(n1175),.clk(gclk));
	jand g1103(.dina(w_n1164_0[0]),.dinb(w_n1175_0[1]),.dout(n1176),.clk(gclk));
	jcb g1104(.dina(n1176),.dinb(w_dff_B_E3buoyro4_1),.dout(n1177));
	jcb g1105(.dina(w_dff_B_qXD20aTC1_0),.dinb(w_n1172_0[0]),.dout(G409));
	jxor g1106(.dina(w_n1162_0[0]),.dinb(w_G384_0),.dout(n1179),.clk(gclk));
	jxor g1107(.dina(w_n937_0[0]),.dinb(w_G396_0[0]),.dout(n1180),.clk(gclk));
	jxor g1108(.dina(w_n988_0[0]),.dinb(w_G387_0[0]),.dout(n1181),.clk(gclk));
	jxor g1109(.dina(n1181),.dinb(w_dff_B_I5WQYAhc1_1),.dout(n1182),.clk(gclk));
	jxor g1110(.dina(w_dff_B_RDYtqR090_0),.dinb(n1179),.dout(n1183),.clk(gclk));
	jand g1111(.dina(w_n1175_0[0]),.dinb(w_G213_0[0]),.dout(n1184),.clk(gclk));
	jnot g1112(.din(w_n1184_0[1]),.dout(n1185),.clk(gclk));
	jcb g1113(.dina(n1185),.dinb(w_dff_B_qN8Zq43O3_1),.dout(n1186));
	jxor g1114(.dina(w_n1114_0[0]),.dinb(w_n1049_0[0]),.dout(n1187),.clk(gclk));
	jcb g1115(.dina(w_n1187_0[1]),.dinb(w_n1184_0[0]),.dout(n1188));
	jand g1116(.dina(n1188),.dinb(w_dff_B_KSktY4Mr6_1),.dout(n1189),.clk(gclk));
	jxor g1117(.dina(w_dff_B_jlaeAtZl5_0),.dinb(w_n1183_0[1]),.dout(G405),.clk(gclk));
	jxor g1118(.dina(w_n1187_0[0]),.dinb(w_n1183_0[0]),.dout(G402),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_dff_A_4ccyHmp11_0),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_dff_A_Fou26Hox4_0),.doutb(w_dff_A_tZAQhP2l8_1),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G1_2(.douta(w_dff_A_1hNsEnv72_0),.doutb(w_G1_2[1]),.doutc(w_dff_A_zKO6tXtJ2_2),.din(w_G1_0[1]));
	jspl jspl_w_G1_3(.douta(w_G1_3[0]),.doutb(w_G1_3[1]),.din(w_G1_0[2]));
	jspl3 jspl3_w_G13_0(.douta(w_G13_0[0]),.doutb(w_dff_A_2PjEZTO05_1),.doutc(w_dff_A_xLxPARyb1_2),.din(G13));
	jspl jspl_w_G13_1(.douta(w_G13_1[0]),.doutb(w_G13_1[1]),.din(w_G13_0[0]));
	jspl3 jspl3_w_G20_0(.douta(w_dff_A_mzOzAUZf7_0),.doutb(w_G20_0[1]),.doutc(w_G20_0[2]),.din(G20));
	jspl3 jspl3_w_G20_1(.douta(w_G20_1[0]),.doutb(w_G20_1[1]),.doutc(w_dff_A_gWXHEB4g6_2),.din(w_G20_0[0]));
	jspl3 jspl3_w_G20_2(.douta(w_G20_2[0]),.doutb(w_dff_A_56JqZ5B84_1),.doutc(w_G20_2[2]),.din(w_G20_0[1]));
	jspl3 jspl3_w_G20_3(.douta(w_G20_3[0]),.doutb(w_dff_A_KFtuu9GJ7_1),.doutc(w_dff_A_ExMXZJ148_2),.din(w_G20_0[2]));
	jspl3 jspl3_w_G20_4(.douta(w_dff_A_FrLgA80Y5_0),.doutb(w_dff_A_BiQXPWQW1_1),.doutc(w_G20_4[2]),.din(w_G20_1[0]));
	jspl3 jspl3_w_G20_5(.douta(w_dff_A_kzFWYfB52_0),.doutb(w_dff_A_86qZ2guA2_1),.doutc(w_G20_5[2]),.din(w_G20_1[1]));
	jspl3 jspl3_w_G20_6(.douta(w_dff_A_ssqYW7xV1_0),.doutb(w_G20_6[1]),.doutc(w_G20_6[2]),.din(w_G20_1[2]));
	jspl jspl_w_G20_7(.douta(w_G20_7[0]),.doutb(w_G20_7[1]),.din(w_G20_2[0]));
	jspl3 jspl3_w_G33_0(.douta(w_dff_A_dPMt59dE4_0),.doutb(w_G33_0[1]),.doutc(w_G33_0[2]),.din(G33));
	jspl3 jspl3_w_G33_1(.douta(w_G33_1[0]),.doutb(w_dff_A_HlyjsgJx5_1),.doutc(w_G33_1[2]),.din(w_G33_0[0]));
	jspl3 jspl3_w_G33_2(.douta(w_G33_2[0]),.doutb(w_G33_2[1]),.doutc(w_G33_2[2]),.din(w_G33_0[1]));
	jspl3 jspl3_w_G33_3(.douta(w_G33_3[0]),.doutb(w_G33_3[1]),.doutc(w_dff_A_OJmdWQiM5_2),.din(w_G33_0[2]));
	jspl3 jspl3_w_G33_4(.douta(w_G33_4[0]),.doutb(w_dff_A_PdBQPsih0_1),.doutc(w_dff_A_swxpps9B3_2),.din(w_G33_1[0]));
	jspl3 jspl3_w_G33_5(.douta(w_G33_5[0]),.doutb(w_G33_5[1]),.doutc(w_dff_A_KLAYTlk53_2),.din(w_G33_1[1]));
	jspl3 jspl3_w_G33_6(.douta(w_dff_A_RvgJFnRR0_0),.doutb(w_dff_A_3m2KYaT92_1),.doutc(w_G33_6[2]),.din(w_G33_1[2]));
	jspl3 jspl3_w_G33_7(.douta(w_G33_7[0]),.doutb(w_G33_7[1]),.doutc(w_G33_7[2]),.din(w_G33_2[0]));
	jspl3 jspl3_w_G33_8(.douta(w_dff_A_tIDm05Cz1_0),.doutb(w_G33_8[1]),.doutc(w_G33_8[2]),.din(w_G33_2[1]));
	jspl3 jspl3_w_G33_9(.douta(w_G33_9[0]),.doutb(w_G33_9[1]),.doutc(w_dff_A_y5rIwcE93_2),.din(w_G33_2[2]));
	jspl3 jspl3_w_G33_10(.douta(w_dff_A_krMXfSYv2_0),.doutb(w_dff_A_YsH3D4I38_1),.doutc(w_G33_10[2]),.din(w_G33_3[0]));
	jspl3 jspl3_w_G33_11(.douta(w_G33_11[0]),.doutb(w_G33_11[1]),.doutc(w_G33_11[2]),.din(w_G33_3[1]));
	jspl3 jspl3_w_G41_0(.douta(w_G41_0[0]),.doutb(w_dff_A_8EkU4qhP9_1),.doutc(w_dff_A_XDkJrU828_2),.din(G41));
	jspl jspl_w_G41_1(.douta(w_G41_1[0]),.doutb(w_G41_1[1]),.din(w_G41_0[0]));
	jspl3 jspl3_w_G45_0(.douta(w_G45_0[0]),.doutb(w_dff_A_npIB8IR04_1),.doutc(w_dff_A_DJiarWZ95_2),.din(G45));
	jspl3 jspl3_w_G45_1(.douta(w_dff_A_TY2VhRBY5_0),.doutb(w_dff_A_S7dmdcD61_1),.doutc(w_G45_1[2]),.din(w_G45_0[0]));
	jspl3 jspl3_w_G50_0(.douta(w_G50_0[0]),.doutb(w_dff_A_7itG0YhZ9_1),.doutc(w_G50_0[2]),.din(G50));
	jspl3 jspl3_w_G50_1(.douta(w_dff_A_ps1pBBQg0_0),.doutb(w_G50_1[1]),.doutc(w_dff_A_bhT07Qpo8_2),.din(w_G50_0[0]));
	jspl3 jspl3_w_G50_2(.douta(w_dff_A_GMDgsM5t5_0),.doutb(w_G50_2[1]),.doutc(w_G50_2[2]),.din(w_G50_0[1]));
	jspl3 jspl3_w_G50_3(.douta(w_dff_A_0BzWVpQx9_0),.doutb(w_G50_3[1]),.doutc(w_dff_A_sRnO9raa1_2),.din(w_G50_0[2]));
	jspl3 jspl3_w_G50_4(.douta(w_dff_A_ldFcLSv06_0),.doutb(w_G50_4[1]),.doutc(w_G50_4[2]),.din(w_G50_1[0]));
	jspl3 jspl3_w_G50_5(.douta(w_G50_5[0]),.doutb(w_dff_A_zBQyaB0w2_1),.doutc(w_G50_5[2]),.din(w_G50_1[1]));
	jspl3 jspl3_w_G58_0(.douta(w_G58_0[0]),.doutb(w_dff_A_Jefdi59f3_1),.doutc(w_dff_A_LtOaC5ti7_2),.din(G58));
	jspl3 jspl3_w_G58_1(.douta(w_dff_A_oirhwcSF6_0),.doutb(w_G58_1[1]),.doutc(w_dff_A_K12y90Dv4_2),.din(w_G58_0[0]));
	jspl3 jspl3_w_G58_2(.douta(w_dff_A_vVDfAQXi7_0),.doutb(w_G58_2[1]),.doutc(w_dff_A_tLivtiAV8_2),.din(w_G58_0[1]));
	jspl3 jspl3_w_G58_3(.douta(w_dff_A_odEjqQBT9_0),.doutb(w_dff_A_tbzMfHWv2_1),.doutc(w_G58_3[2]),.din(w_G58_0[2]));
	jspl3 jspl3_w_G58_4(.douta(w_G58_4[0]),.doutb(w_dff_A_XNG8O2VN2_1),.doutc(w_G58_4[2]),.din(w_G58_1[0]));
	jspl jspl_w_G58_5(.douta(w_G58_5[0]),.doutb(w_G58_5[1]),.din(w_G58_1[1]));
	jspl3 jspl3_w_G68_0(.douta(w_G68_0[0]),.doutb(w_G68_0[1]),.doutc(w_dff_A_bLHzeMOq5_2),.din(G68));
	jspl3 jspl3_w_G68_1(.douta(w_dff_A_CO2XZcYU0_0),.doutb(w_G68_1[1]),.doutc(w_dff_A_4WU1ylqH1_2),.din(w_G68_0[0]));
	jspl3 jspl3_w_G68_2(.douta(w_G68_2[0]),.doutb(w_dff_A_skVO2sRG1_1),.doutc(w_dff_A_9nNLVVbJ4_2),.din(w_G68_0[1]));
	jspl3 jspl3_w_G68_3(.douta(w_G68_3[0]),.doutb(w_dff_A_wLrENlk49_1),.doutc(w_dff_A_i2IVPP7p7_2),.din(w_G68_0[2]));
	jspl3 jspl3_w_G68_4(.douta(w_dff_A_QT5SPFcM2_0),.doutb(w_G68_4[1]),.doutc(w_G68_4[2]),.din(w_G68_1[0]));
	jspl jspl_w_G68_5(.douta(w_G68_5[0]),.doutb(w_G68_5[1]),.din(w_G68_1[1]));
	jspl3 jspl3_w_G77_0(.douta(w_G77_0[0]),.doutb(w_G77_0[1]),.doutc(w_G77_0[2]),.din(G77));
	jspl3 jspl3_w_G77_1(.douta(w_dff_A_JeMaVs6t4_0),.doutb(w_G77_1[1]),.doutc(w_dff_A_8sWGGBbl3_2),.din(w_G77_0[0]));
	jspl3 jspl3_w_G77_2(.douta(w_G77_2[0]),.doutb(w_dff_A_hPLRTLOf3_1),.doutc(w_dff_A_59ogoqPM0_2),.din(w_G77_0[1]));
	jspl3 jspl3_w_G77_3(.douta(w_G77_3[0]),.doutb(w_dff_A_ptzGm7K20_1),.doutc(w_G77_3[2]),.din(w_G77_0[2]));
	jspl3 jspl3_w_G77_4(.douta(w_G77_4[0]),.doutb(w_G77_4[1]),.doutc(w_G77_4[2]),.din(w_G77_1[0]));
	jspl jspl_w_G77_5(.douta(w_G77_5[0]),.doutb(w_G77_5[1]),.din(w_G77_1[1]));
	jspl3 jspl3_w_G87_0(.douta(w_dff_A_FvwJAaIG2_0),.doutb(w_G87_0[1]),.doutc(w_G87_0[2]),.din(G87));
	jspl3 jspl3_w_G87_1(.douta(w_G87_1[0]),.doutb(w_dff_A_kiZ2YnPA2_1),.doutc(w_dff_A_o4LQQvKM3_2),.din(w_G87_0[0]));
	jspl3 jspl3_w_G87_2(.douta(w_dff_A_QGVfY15l5_0),.doutb(w_dff_A_udX6hQZn4_1),.doutc(w_G87_2[2]),.din(w_G87_0[1]));
	jspl3 jspl3_w_G87_3(.douta(w_dff_A_6pRkK9FN2_0),.doutb(w_G87_3[1]),.doutc(w_dff_A_mWHgdEQc4_2),.din(w_G87_0[2]));
	jspl3 jspl3_w_G97_0(.douta(w_G97_0[0]),.doutb(w_dff_A_GPRLNY7X4_1),.doutc(w_dff_A_C1VcRIZQ0_2),.din(G97));
	jspl3 jspl3_w_G97_1(.douta(w_G97_1[0]),.doutb(w_G97_1[1]),.doutc(w_dff_A_criETge50_2),.din(w_G97_0[0]));
	jspl3 jspl3_w_G97_2(.douta(w_G97_2[0]),.doutb(w_G97_2[1]),.doutc(w_dff_A_7AcN7zvh3_2),.din(w_G97_0[1]));
	jspl3 jspl3_w_G97_3(.douta(w_dff_A_O2VcMFTg2_0),.doutb(w_dff_A_RZwJTBHH0_1),.doutc(w_G97_3[2]),.din(w_G97_0[2]));
	jspl3 jspl3_w_G97_4(.douta(w_dff_A_dznUlpk64_0),.doutb(w_G97_4[1]),.doutc(w_G97_4[2]),.din(w_G97_1[0]));
	jspl jspl_w_G97_5(.douta(w_dff_A_yzUpWH5M6_0),.doutb(w_G97_5[1]),.din(w_G97_1[1]));
	jspl3 jspl3_w_G107_0(.douta(w_G107_0[0]),.doutb(w_dff_A_uVI7mBqD7_1),.doutc(w_dff_A_dGUtwM5M9_2),.din(G107));
	jspl3 jspl3_w_G107_1(.douta(w_G107_1[0]),.doutb(w_G107_1[1]),.doutc(w_dff_A_ucjKX2Ip8_2),.din(w_G107_0[0]));
	jspl3 jspl3_w_G107_2(.douta(w_G107_2[0]),.doutb(w_G107_2[1]),.doutc(w_dff_A_G37cgPAn4_2),.din(w_G107_0[1]));
	jspl3 jspl3_w_G107_3(.douta(w_dff_A_l8rs1oAb6_0),.doutb(w_dff_A_ybYp2lXE1_1),.doutc(w_G107_3[2]),.din(w_G107_0[2]));
	jspl3 jspl3_w_G107_4(.douta(w_dff_A_ygo3ADFz2_0),.doutb(w_G107_4[1]),.doutc(w_G107_4[2]),.din(w_G107_1[0]));
	jspl jspl_w_G107_5(.douta(w_G107_5[0]),.doutb(w_G107_5[1]),.din(w_G107_1[1]));
	jspl3 jspl3_w_G116_0(.douta(w_G116_0[0]),.doutb(w_dff_A_W9EB8iqA1_1),.doutc(w_dff_A_RRQhBpxU0_2),.din(G116));
	jspl3 jspl3_w_G116_1(.douta(w_G116_1[0]),.doutb(w_dff_A_1JXlQGbO6_1),.doutc(w_dff_A_uiWlur9c6_2),.din(w_G116_0[0]));
	jspl3 jspl3_w_G116_2(.douta(w_G116_2[0]),.doutb(w_dff_A_c9wDqvvY5_1),.doutc(w_dff_A_j3wkjTyJ9_2),.din(w_G116_0[1]));
	jspl3 jspl3_w_G116_3(.douta(w_dff_A_Ul9C7h3E4_0),.doutb(w_G116_3[1]),.doutc(w_dff_A_aVf2RN5x9_2),.din(w_G116_0[2]));
	jspl3 jspl3_w_G116_4(.douta(w_G116_4[0]),.doutb(w_G116_4[1]),.doutc(w_G116_4[2]),.din(w_G116_1[0]));
	jspl jspl_w_G125_0(.douta(w_G125_0[0]),.doutb(w_G125_0[1]),.din(w_dff_B_3NFxnZsM7_2));
	jspl3 jspl3_w_G128_0(.douta(w_G128_0[0]),.doutb(w_G128_0[1]),.doutc(w_G128_0[2]),.din(w_dff_B_k4zStVQl6_3));
	jspl3 jspl3_w_G132_0(.douta(w_G132_0[0]),.doutb(w_G132_0[1]),.doutc(w_G132_0[2]),.din(w_dff_B_YQvH26gl2_3));
	jspl jspl_w_G132_1(.douta(w_G132_1[0]),.doutb(w_G132_1[1]),.din(w_G132_0[0]));
	jspl3 jspl3_w_G137_0(.douta(w_G137_0[0]),.doutb(w_G137_0[1]),.doutc(w_G137_0[2]),.din(w_dff_B_PhCYIDkf7_3));
	jspl3 jspl3_w_G137_1(.douta(w_G137_1[0]),.doutb(w_G137_1[1]),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G143_0(.douta(w_G143_0[0]),.doutb(w_G143_0[1]),.doutc(w_G143_0[2]),.din(w_dff_B_t5fzPJDL5_3));
	jspl3 jspl3_w_G143_1(.douta(w_dff_A_5a2f4HA13_0),.doutb(w_G143_1[1]),.doutc(w_G143_1[2]),.din(w_G143_0[0]));
	jspl jspl_w_G143_2(.douta(w_G143_2[0]),.doutb(w_G143_2[1]),.din(w_G143_0[1]));
	jspl3 jspl3_w_G150_0(.douta(w_dff_A_7JjrxqHK3_0),.doutb(w_dff_A_3O7aE85M4_1),.doutc(w_G150_0[2]),.din(G150));
	jspl3 jspl3_w_G150_1(.douta(w_G150_1[0]),.doutb(w_dff_A_jy5KOk1X7_1),.doutc(w_dff_A_H7I5RNYx4_2),.din(w_G150_0[0]));
	jspl3 jspl3_w_G150_2(.douta(w_G150_2[0]),.doutb(w_G150_2[1]),.doutc(w_G150_2[2]),.din(w_G150_0[1]));
	jspl jspl_w_G150_3(.douta(w_dff_A_G446uEg82_0),.doutb(w_G150_3[1]),.din(w_G150_0[2]));
	jspl3 jspl3_w_G159_0(.douta(w_dff_A_Sb91akbp9_0),.doutb(w_dff_A_7A7o9IQa1_1),.doutc(w_G159_0[2]),.din(w_dff_B_GuEHFn4Z5_3));
	jspl3 jspl3_w_G159_1(.douta(w_G159_1[0]),.doutb(w_G159_1[1]),.doutc(w_G159_1[2]),.din(w_G159_0[0]));
	jspl3 jspl3_w_G159_2(.douta(w_G159_2[0]),.doutb(w_G159_2[1]),.doutc(w_G159_2[2]),.din(w_G159_0[1]));
	jspl3 jspl3_w_G159_3(.douta(w_dff_A_Ct00FSky8_0),.doutb(w_dff_A_d7nwO7Jr9_1),.doutc(w_G159_3[2]),.din(w_G159_0[2]));
	jspl3 jspl3_w_G169_0(.douta(w_G169_0[0]),.doutb(w_dff_A_sK7Q5PHe8_1),.doutc(w_dff_A_H15fiu2u7_2),.din(G169));
	jspl jspl_w_G169_1(.douta(w_dff_A_6uEwpP187_0),.doutb(w_G169_1[1]),.din(w_G169_0[0]));
	jspl3 jspl3_w_G179_0(.douta(w_dff_A_53Uc2rbS7_0),.doutb(w_G179_0[1]),.doutc(w_G179_0[2]),.din(G179));
	jspl3 jspl3_w_G179_1(.douta(w_dff_A_CXN2s6KH5_0),.doutb(w_G179_1[1]),.doutc(w_G179_1[2]),.din(w_G179_0[0]));
	jspl3 jspl3_w_G179_2(.douta(w_dff_A_Fc5aWhdd9_0),.doutb(w_dff_A_OimBSSv70_1),.doutc(w_G179_2[2]),.din(w_G179_0[1]));
	jspl3 jspl3_w_G190_0(.douta(w_dff_A_RUd1jwHC1_0),.doutb(w_dff_A_1dXG9ppK9_1),.doutc(w_G190_0[2]),.din(G190));
	jspl3 jspl3_w_G190_1(.douta(w_dff_A_BfNynjZ25_0),.doutb(w_G190_1[1]),.doutc(w_G190_1[2]),.din(w_G190_0[0]));
	jspl3 jspl3_w_G190_2(.douta(w_G190_2[0]),.doutb(w_dff_A_Ey0AHIns3_1),.doutc(w_dff_A_sNGWQ4tz3_2),.din(w_G190_0[1]));
	jspl3 jspl3_w_G190_3(.douta(w_G190_3[0]),.doutb(w_dff_A_izkfXpqB4_1),.doutc(w_dff_A_y8Uk3cet7_2),.din(w_G190_0[2]));
	jspl jspl_w_G190_4(.douta(w_G190_4[0]),.doutb(w_G190_4[1]),.din(w_G190_1[0]));
	jspl3 jspl3_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.doutc(w_dff_A_UviIzfNq3_2),.din(G200));
	jspl3 jspl3_w_G200_1(.douta(w_dff_A_Cxmm5ts75_0),.doutb(w_dff_A_dmI39b8w6_1),.doutc(w_G200_1[2]),.din(w_G200_0[0]));
	jspl3 jspl3_w_G200_2(.douta(w_G200_2[0]),.doutb(w_dff_A_OZ9A1o2l5_1),.doutc(w_dff_A_fGxofY8k0_2),.din(w_G200_0[1]));
	jspl3 jspl3_w_G200_3(.douta(w_G200_3[0]),.doutb(w_G200_3[1]),.doutc(w_dff_A_oLRdNPdw6_2),.din(w_G200_0[2]));
	jspl3 jspl3_w_G200_4(.douta(w_G200_4[0]),.doutb(w_G200_4[1]),.doutc(w_G200_4[2]),.din(w_G200_1[0]));
	jspl3 jspl3_w_G213_0(.douta(w_dff_A_ploXWUQo9_0),.doutb(w_G213_0[1]),.doutc(w_dff_A_ojWxuxiD0_2),.din(G213));
	jspl jspl_w_G223_0(.douta(w_G223_0[0]),.doutb(w_G223_0[1]),.din(w_dff_B_El1Kyins8_2));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_dff_A_JJ9RWBLE3_1),.doutc(w_dff_A_uQxop5AO8_2),.din(G226));
	jspl jspl_w_G226_1(.douta(w_dff_A_Ntvkszga7_0),.doutb(w_G226_1[1]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G232_0(.douta(w_G232_0[0]),.doutb(w_dff_A_mI5bW7u41_1),.doutc(w_dff_A_fVvvUUjm7_2),.din(G232));
	jspl3 jspl3_w_G232_1(.douta(w_dff_A_kSMsUd1o0_0),.doutb(w_dff_A_iZGzzApM4_1),.doutc(w_G232_1[2]),.din(w_G232_0[0]));
	jspl3 jspl3_w_G238_0(.douta(w_G238_0[0]),.doutb(w_dff_A_i6QxGQVe1_1),.doutc(w_dff_A_FsqTWjI07_2),.din(G238));
	jspl3 jspl3_w_G238_1(.douta(w_dff_A_Yqz3Gn3v8_0),.doutb(w_G238_1[1]),.doutc(w_G238_1[2]),.din(w_G238_0[0]));
	jspl3 jspl3_w_G244_0(.douta(w_G244_0[0]),.doutb(w_dff_A_SEmmsmwT0_1),.doutc(w_dff_A_h8ARcq9S8_2),.din(G244));
	jspl3 jspl3_w_G244_1(.douta(w_dff_A_tC83FC8o7_0),.doutb(w_G244_1[1]),.doutc(w_G244_1[2]),.din(w_G244_0[0]));
	jspl3 jspl3_w_G250_0(.douta(w_dff_A_J0qcyDa95_0),.doutb(w_dff_A_2UtXVpAi1_1),.doutc(w_G250_0[2]),.din(G250));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_dff_A_Ny0Ff4VQ5_1),.doutc(w_dff_A_eo3IM3vo2_2),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_ydIkuUtG6_0),.doutb(w_dff_A_cZljE8hi0_1),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G264_0(.douta(w_G264_0[0]),.doutb(w_dff_A_YBHsC95D4_1),.doutc(w_dff_A_j7dOrHzR6_2),.din(G264));
	jspl jspl_w_G264_1(.douta(w_G264_1[0]),.doutb(w_G264_1[1]),.din(w_G264_0[0]));
	jspl3 jspl3_w_G270_0(.douta(w_dff_A_uShzZ3Uv1_0),.doutb(w_G270_0[1]),.doutc(w_G270_0[2]),.din(G270));
	jspl3 jspl3_w_G274_0(.douta(w_dff_A_rZ2wUsBs6_0),.doutb(w_G274_0[1]),.doutc(w_dff_A_HiU1UimC1_2),.din(G274));
	jspl3 jspl3_w_G283_0(.douta(w_dff_A_9J0G4DIm3_0),.doutb(w_dff_A_HY0WJrlP2_1),.doutc(w_G283_0[2]),.din(G283));
	jspl3 jspl3_w_G283_1(.douta(w_G283_1[0]),.doutb(w_G283_1[1]),.doutc(w_G283_1[2]),.din(w_G283_0[0]));
	jspl3 jspl3_w_G283_2(.douta(w_dff_A_SzkP9lAQ1_0),.doutb(w_dff_A_xZZrXenR4_1),.doutc(w_G283_2[2]),.din(w_G283_0[1]));
	jspl3 jspl3_w_G283_3(.douta(w_dff_A_2JC8ADef4_0),.doutb(w_dff_A_QADLD1h01_1),.doutc(w_G283_3[2]),.din(w_G283_0[2]));
	jspl3 jspl3_w_G294_0(.douta(w_dff_A_OtV27sqM7_0),.doutb(w_dff_A_As1zAiFl1_1),.doutc(w_G294_0[2]),.din(G294));
	jspl3 jspl3_w_G294_1(.douta(w_G294_1[0]),.doutb(w_G294_1[1]),.doutc(w_G294_1[2]),.din(w_G294_0[0]));
	jspl3 jspl3_w_G294_2(.douta(w_dff_A_Ec9Kqgjw8_0),.doutb(w_G294_2[1]),.doutc(w_G294_2[2]),.din(w_G294_0[1]));
	jspl jspl_w_G294_3(.douta(w_dff_A_uqeqgqm72_0),.doutb(w_G294_3[1]),.din(w_G294_0[2]));
	jspl3 jspl3_w_G303_0(.douta(w_dff_A_O00dREir7_0),.doutb(w_G303_0[1]),.doutc(w_dff_A_nzLoglhV6_2),.din(G303));
	jspl3 jspl3_w_G303_1(.douta(w_G303_1[0]),.doutb(w_G303_1[1]),.doutc(w_G303_1[2]),.din(w_G303_0[0]));
	jspl3 jspl3_w_G303_2(.douta(w_dff_A_6SZHnbiP5_0),.doutb(w_dff_A_n2oDV0SI8_1),.doutc(w_G303_2[2]),.din(w_G303_0[1]));
	jspl3 jspl3_w_G311_0(.douta(w_G311_0[0]),.doutb(w_G311_0[1]),.doutc(w_G311_0[2]),.din(w_dff_B_p5xIi9sp7_3));
	jspl3 jspl3_w_G311_1(.douta(w_G311_1[0]),.doutb(w_G311_1[1]),.doutc(w_G311_1[2]),.din(w_G311_0[0]));
	jspl3 jspl3_w_G317_0(.douta(w_G317_0[0]),.doutb(w_G317_0[1]),.doutc(w_G317_0[2]),.din(w_dff_B_fFWHIJFq9_3));
	jspl jspl_w_G317_1(.douta(w_G317_1[0]),.doutb(w_G317_1[1]),.din(w_G317_0[0]));
	jspl3 jspl3_w_G322_0(.douta(w_G322_0[0]),.doutb(w_G322_0[1]),.doutc(w_G322_0[2]),.din(w_dff_B_ug54TCuZ7_3));
	jspl jspl_w_G326_0(.douta(w_G326_0[0]),.doutb(w_G326_0[1]),.din(w_dff_B_sAp9YiIm4_2));
	jspl jspl_w_G330_0(.douta(w_dff_A_stwUmo9O5_0),.doutb(w_G330_0[1]),.din(G330));
	jspl jspl_w_G343_0(.douta(w_G343_0[0]),.doutb(w_dff_A_9bWExnt25_1),.din(G343));
	jspl3 jspl3_w_G1698_0(.douta(w_G1698_0[0]),.doutb(w_G1698_0[1]),.doutc(w_dff_A_InfOy5b73_2),.din(G1698));
	jspl jspl_w_G355_0(.douta(w_G355_0),.doutb(G355),.din(G355_fa_));
	jspl3 jspl3_w_G396_0(.douta(w_dff_A_8WxTUa831_0),.doutb(w_G396_0[1]),.doutc(G396),.din(G396_fa_));
	jspl jspl_w_G384_0(.douta(w_dff_A_eed2vNmR3_0),.doutb(G384),.din(G384_fa_));
	jspl3 jspl3_w_G387_0(.douta(w_G387_0[0]),.doutb(w_G387_0[1]),.doutc(G387),.din(G387_fa_));
	jspl3 jspl3_w_n72_0(.douta(w_n72_0[0]),.doutb(w_dff_A_KNB7jK4F8_1),.doutc(w_dff_A_bUhcjxrq5_2),.din(n72));
	jspl jspl_w_n72_1(.douta(w_n72_1[0]),.doutb(w_dff_A_SxUhH09K8_1),.din(w_n72_0[0]));
	jspl3 jspl3_w_n73_0(.douta(w_n73_0[0]),.doutb(w_n73_0[1]),.doutc(w_dff_A_R2ndmZqm6_2),.din(n73));
	jspl3 jspl3_w_n73_1(.douta(w_n73_1[0]),.doutb(w_dff_A_HdEUKy3C7_1),.doutc(w_n73_1[2]),.din(w_n73_0[0]));
	jspl3 jspl3_w_n73_2(.douta(w_dff_A_LiCi63DK0_0),.doutb(w_n73_2[1]),.doutc(w_dff_A_VnmzGIqZ9_2),.din(w_n73_0[1]));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_dff_A_b7CJdTKD3_1),.doutc(w_dff_A_zQKuk2nr8_2),.din(n74));
	jspl jspl_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.din(w_n74_0[0]));
	jspl3 jspl3_w_n75_0(.douta(w_n75_0[0]),.doutb(w_dff_A_t7kP4Kj38_1),.doutc(w_dff_A_nj2QBwlE1_2),.din(n75));
	jspl jspl_w_n75_1(.douta(w_n75_1[0]),.doutb(w_n75_1[1]),.din(w_n75_0[0]));
	jspl jspl_w_n76_0(.douta(w_n76_0[0]),.doutb(w_n76_0[1]),.din(n76));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl3 jspl3_w_n79_0(.douta(w_dff_A_G6UuLri30_0),.doutb(w_n79_0[1]),.doutc(w_n79_0[2]),.din(n79));
	jspl3 jspl3_w_n80_0(.douta(w_n80_0[0]),.doutb(w_dff_A_nQ70BLCU2_1),.doutc(w_dff_A_e7fhqZWt8_2),.din(n80));
	jspl jspl_w_n80_1(.douta(w_n80_1[0]),.doutb(w_n80_1[1]),.din(w_n80_0[0]));
	jspl3 jspl3_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.doutc(w_n81_0[2]),.din(n81));
	jspl3 jspl3_w_n85_0(.douta(w_dff_A_nCQ6NDQn7_0),.doutb(w_n85_0[1]),.doutc(w_dff_A_mKrXYaZq8_2),.din(n85));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl3 jspl3_w_n88_0(.douta(w_n88_0[0]),.doutb(w_dff_A_i99ftJfc5_1),.doutc(w_n88_0[2]),.din(n88));
	jspl jspl_w_n88_1(.douta(w_n88_1[0]),.doutb(w_n88_1[1]),.din(w_n88_0[0]));
	jspl3 jspl3_w_n91_0(.douta(w_n91_0[0]),.doutb(w_n91_0[1]),.doutc(w_n91_0[2]),.din(n91));
	jspl3 jspl3_w_n91_1(.douta(w_dff_A_PwEDttqh4_0),.doutb(w_n91_1[1]),.doutc(w_n91_1[2]),.din(w_n91_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n97_0(.douta(w_dff_A_yqm5Cmbs8_0),.doutb(w_n97_0[1]),.doutc(w_n97_0[2]),.din(n97));
	jspl3 jspl3_w_n97_1(.douta(w_n97_1[0]),.doutb(w_dff_A_4u2Un4vU5_1),.doutc(w_n97_1[2]),.din(w_n97_0[0]));
	jspl jspl_w_n97_2(.douta(w_n97_2[0]),.doutb(w_n97_2[1]),.din(w_n97_0[1]));
	jspl3 jspl3_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.doutc(w_n98_0[2]),.din(n98));
	jspl3 jspl3_w_n98_1(.douta(w_n98_1[0]),.doutb(w_n98_1[1]),.doutc(w_n98_1[2]),.din(w_n98_0[0]));
	jspl jspl_w_n98_2(.douta(w_dff_A_coblnMg10_0),.doutb(w_n98_2[1]),.din(w_n98_0[1]));
	jspl3 jspl3_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.doutc(w_n103_0[2]),.din(n103));
	jspl3 jspl3_w_n105_0(.douta(w_dff_A_GQxHmHkp4_0),.doutb(w_n105_0[1]),.doutc(w_dff_A_XqgdXkng9_2),.din(n105));
	jspl3 jspl3_w_n105_1(.douta(w_dff_A_rvC2vt7T8_0),.doutb(w_n105_1[1]),.doutc(w_dff_A_9ZunfM6Y5_2),.din(w_n105_0[0]));
	jspl jspl_w_n105_2(.douta(w_n105_2[0]),.doutb(w_n105_2[1]),.din(w_n105_0[1]));
	jspl jspl_w_n106_0(.douta(w_dff_A_FDiH7MW27_0),.doutb(w_n106_0[1]),.din(n106));
	jspl3 jspl3_w_n112_0(.douta(w_n112_0[0]),.doutb(w_n112_0[1]),.doutc(w_n112_0[2]),.din(n112));
	jspl3 jspl3_w_n112_1(.douta(w_n112_1[0]),.doutb(w_n112_1[1]),.doutc(w_n112_1[2]),.din(w_n112_0[0]));
	jspl3 jspl3_w_n112_2(.douta(w_n112_2[0]),.doutb(w_n112_2[1]),.doutc(w_n112_2[2]),.din(w_n112_0[1]));
	jspl3 jspl3_w_n112_3(.douta(w_dff_A_IlnhALf97_0),.doutb(w_dff_A_CgQNpzjX4_1),.doutc(w_n112_3[2]),.din(w_n112_0[2]));
	jspl3 jspl3_w_n112_4(.douta(w_dff_A_tIMCN33B9_0),.doutb(w_n112_4[1]),.doutc(w_n112_4[2]),.din(w_n112_1[0]));
	jspl3 jspl3_w_n112_5(.douta(w_n112_5[0]),.doutb(w_n112_5[1]),.doutc(w_n112_5[2]),.din(w_n112_1[1]));
	jspl3 jspl3_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.doutc(w_n113_0[2]),.din(n113));
	jspl3 jspl3_w_n113_1(.douta(w_dff_A_MANApDwJ0_0),.doutb(w_dff_A_WdJmdwBX6_1),.doutc(w_n113_1[2]),.din(w_n113_0[0]));
	jspl3 jspl3_w_n113_2(.douta(w_n113_2[0]),.doutb(w_n113_2[1]),.doutc(w_n113_2[2]),.din(w_n113_0[1]));
	jspl jspl_w_n113_3(.douta(w_n113_3[0]),.doutb(w_n113_3[1]),.din(w_n113_0[2]));
	jspl3 jspl3_w_n114_0(.douta(w_n114_0[0]),.doutb(w_dff_A_j7mMMThK7_1),.doutc(w_n114_0[2]),.din(n114));
	jspl3 jspl3_w_n114_1(.douta(w_n114_1[0]),.doutb(w_n114_1[1]),.doutc(w_n114_1[2]),.din(w_n114_0[0]));
	jspl3 jspl3_w_n115_0(.douta(w_n115_0[0]),.doutb(w_dff_A_5b4c8wso7_1),.doutc(w_n115_0[2]),.din(n115));
	jspl jspl_w_n115_1(.douta(w_n115_1[0]),.doutb(w_n115_1[1]),.din(w_n115_0[0]));
	jspl jspl_w_n116_0(.douta(w_n116_0[0]),.doutb(w_dff_A_7X6XhEQy8_1),.din(w_dff_B_275f0nXt2_2));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl3 jspl3_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.doutc(w_n121_0[2]),.din(n121));
	jspl3 jspl3_w_n122_0(.douta(w_n122_0[0]),.doutb(w_n122_0[1]),.doutc(w_n122_0[2]),.din(n122));
	jspl jspl_w_n122_1(.douta(w_n122_1[0]),.doutb(w_n122_1[1]),.din(w_n122_0[0]));
	jspl3 jspl3_w_n123_0(.douta(w_n123_0[0]),.doutb(w_n123_0[1]),.doutc(w_n123_0[2]),.din(n123));
	jspl3 jspl3_w_n123_1(.douta(w_n123_1[0]),.doutb(w_n123_1[1]),.doutc(w_n123_1[2]),.din(w_n123_0[0]));
	jspl jspl_w_n131_0(.douta(w_dff_A_AZhXc43T4_0),.doutb(w_n131_0[1]),.din(n131));
	jspl jspl_w_n135_0(.douta(w_n135_0[0]),.doutb(w_dff_A_Yxo3N9Dl4_1),.din(n135));
	jspl3 jspl3_w_n137_0(.douta(w_n137_0[0]),.doutb(w_n137_0[1]),.doutc(w_n137_0[2]),.din(n137));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(w_dff_B_DU2XGEIQ6_2));
	jspl3 jspl3_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_ZUfJKdXR1_1),.doutc(w_dff_A_IF5vSjQB9_2),.din(n146));
	jspl3 jspl3_w_n146_1(.douta(w_n146_1[0]),.doutb(w_dff_A_lqWvE3r74_1),.doutc(w_dff_A_5HJK33pc5_2),.din(w_n146_0[0]));
	jspl3 jspl3_w_n146_2(.douta(w_n146_2[0]),.doutb(w_n146_2[1]),.doutc(w_n146_2[2]),.din(w_n146_0[1]));
	jspl3 jspl3_w_n146_3(.douta(w_n146_3[0]),.doutb(w_dff_A_3DuuZRVa7_1),.doutc(w_n146_3[2]),.din(w_n146_0[2]));
	jspl3 jspl3_w_n147_0(.douta(w_n147_0[0]),.doutb(w_dff_A_gjlubog67_1),.doutc(w_n147_0[2]),.din(n147));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_dff_A_jULG3NAn2_0),.doutb(w_dff_A_DMtX3I347_1),.doutc(w_n148_1[2]),.din(w_n148_0[0]));
	jspl3 jspl3_w_n148_2(.douta(w_n148_2[0]),.doutb(w_n148_2[1]),.doutc(w_n148_2[2]),.din(w_n148_0[1]));
	jspl3 jspl3_w_n148_3(.douta(w_dff_A_Wbs76ppA6_0),.doutb(w_n148_3[1]),.doutc(w_dff_A_eoz6teQ20_2),.din(w_n148_0[2]));
	jspl3 jspl3_w_n148_4(.douta(w_n148_4[0]),.doutb(w_dff_A_weg0WuY85_1),.doutc(w_dff_A_D9DjRBCi5_2),.din(w_n148_1[0]));
	jspl3 jspl3_w_n148_5(.douta(w_n148_5[0]),.doutb(w_dff_A_EI2Ilcku7_1),.doutc(w_dff_A_MVA5MfC56_2),.din(w_n148_1[1]));
	jspl3 jspl3_w_n148_6(.douta(w_n148_6[0]),.doutb(w_n148_6[1]),.doutc(w_n148_6[2]),.din(w_n148_1[2]));
	jspl3 jspl3_w_n148_7(.douta(w_n148_7[0]),.doutb(w_n148_7[1]),.doutc(w_n148_7[2]),.din(w_n148_2[0]));
	jspl3 jspl3_w_n148_8(.douta(w_n148_8[0]),.doutb(w_n148_8[1]),.doutc(w_n148_8[2]),.din(w_n148_2[1]));
	jspl3 jspl3_w_n148_9(.douta(w_n148_9[0]),.doutb(w_n148_9[1]),.doutc(w_n148_9[2]),.din(w_n148_2[2]));
	jspl3 jspl3_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.doutc(w_n149_0[2]),.din(n149));
	jspl3 jspl3_w_n149_1(.douta(w_n149_1[0]),.doutb(w_dff_A_o5lDOTfG0_1),.doutc(w_n149_1[2]),.din(w_n149_0[0]));
	jspl jspl_w_n149_2(.douta(w_dff_A_Ofo02QnI0_0),.doutb(w_n149_2[1]),.din(w_n149_0[1]));
	jspl3 jspl3_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_2ThYXdQ06_1),.doutc(w_dff_A_tOq02BT72_2),.din(n151));
	jspl3 jspl3_w_n151_1(.douta(w_n151_1[0]),.doutb(w_dff_A_ChjD05Oz7_1),.doutc(w_dff_A_klL2CcSO6_2),.din(w_n151_0[0]));
	jspl3 jspl3_w_n151_2(.douta(w_n151_2[0]),.doutb(w_n151_2[1]),.doutc(w_n151_2[2]),.din(w_n151_0[1]));
	jspl3 jspl3_w_n151_3(.douta(w_n151_3[0]),.doutb(w_n151_3[1]),.doutc(w_n151_3[2]),.din(w_n151_0[2]));
	jspl3 jspl3_w_n151_4(.douta(w_n151_4[0]),.doutb(w_dff_A_Vmigz4lE8_1),.doutc(w_dff_A_iqj7eGhw3_2),.din(w_n151_1[0]));
	jspl3 jspl3_w_n152_0(.douta(w_n152_0[0]),.doutb(w_n152_0[1]),.doutc(w_n152_0[2]),.din(n152));
	jspl3 jspl3_w_n152_1(.douta(w_n152_1[0]),.doutb(w_n152_1[1]),.doutc(w_n152_1[2]),.din(w_n152_0[0]));
	jspl3 jspl3_w_n152_2(.douta(w_n152_2[0]),.doutb(w_n152_2[1]),.doutc(w_n152_2[2]),.din(w_n152_0[1]));
	jspl jspl_w_n152_3(.douta(w_n152_3[0]),.doutb(w_n152_3[1]),.din(w_n152_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_n154_0[1]),.din(n154));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl3 jspl3_w_n155_1(.douta(w_n155_1[0]),.doutb(w_n155_1[1]),.doutc(w_n155_1[2]),.din(w_n155_0[0]));
	jspl3 jspl3_w_n155_2(.douta(w_n155_2[0]),.doutb(w_n155_2[1]),.doutc(w_n155_2[2]),.din(w_n155_0[1]));
	jspl jspl_w_n155_3(.douta(w_n155_3[0]),.doutb(w_n155_3[1]),.din(w_n155_0[2]));
	jspl3 jspl3_w_n157_0(.douta(w_dff_A_LmlS4BSt7_0),.doutb(w_n157_0[1]),.doutc(w_dff_A_WEIuYqWf0_2),.din(n157));
	jspl3 jspl3_w_n161_0(.douta(w_n161_0[0]),.doutb(w_n161_0[1]),.doutc(w_dff_A_3cucR8oQ9_2),.din(n161));
	jspl jspl_w_n161_1(.douta(w_n161_1[0]),.doutb(w_n161_1[1]),.din(w_n161_0[0]));
	jspl3 jspl3_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.doutc(w_n162_0[2]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_dff_A_wFga1qG85_0),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n166_0(.douta(w_dff_A_h2y9xBoJ6_0),.doutb(w_n166_0[1]),.doutc(w_n166_0[2]),.din(n166));
	jspl3 jspl3_w_n166_1(.douta(w_n166_1[0]),.doutb(w_dff_A_ONukrniH5_1),.doutc(w_dff_A_2FUbW2rT0_2),.din(w_n166_0[0]));
	jspl3 jspl3_w_n166_2(.douta(w_n166_2[0]),.doutb(w_n166_2[1]),.doutc(w_dff_A_NdF95UbF0_2),.din(w_n166_0[1]));
	jspl jspl_w_n166_3(.douta(w_dff_A_a5XfqDH46_0),.doutb(w_n166_3[1]),.din(w_n166_0[2]));
	jspl3 jspl3_w_n170_0(.douta(w_dff_A_UWPcFigi2_0),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_dff_A_ttZt2BHE1_0),.doutb(w_n172_0[1]),.din(w_dff_B_CJBybfjs7_2));
	jspl3 jspl3_w_n179_0(.douta(w_n179_0[0]),.doutb(w_dff_A_234SJcZS8_1),.doutc(w_dff_A_afzTHK3A5_2),.din(n179));
	jspl3 jspl3_w_n179_1(.douta(w_dff_A_zaqVxPXS5_0),.doutb(w_n179_1[1]),.doutc(w_dff_A_0m7SaP7A3_2),.din(w_n179_0[0]));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl3 jspl3_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.doutc(w_n185_0[2]),.din(n185));
	jspl3 jspl3_w_n185_1(.douta(w_n185_1[0]),.doutb(w_n185_1[1]),.doutc(w_dff_A_20GyYu6S9_2),.din(w_n185_0[0]));
	jspl3 jspl3_w_n185_2(.douta(w_n185_2[0]),.doutb(w_n185_2[1]),.doutc(w_n185_2[2]),.din(w_n185_0[1]));
	jspl3 jspl3_w_n185_3(.douta(w_n185_3[0]),.doutb(w_n185_3[1]),.doutc(w_n185_3[2]),.din(w_n185_0[2]));
	jspl3 jspl3_w_n189_0(.douta(w_n189_0[0]),.doutb(w_dff_A_uXhuoCTd3_1),.doutc(w_dff_A_ss9i5BgQ2_2),.din(n189));
	jspl3 jspl3_w_n189_1(.douta(w_n189_1[0]),.doutb(w_n189_1[1]),.doutc(w_dff_A_BJu1r9gt1_2),.din(w_n189_0[0]));
	jspl jspl_w_n189_2(.douta(w_n189_2[0]),.doutb(w_n189_2[1]),.din(w_n189_0[1]));
	jspl3 jspl3_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.doutc(w_n190_0[2]),.din(n190));
	jspl3 jspl3_w_n190_1(.douta(w_n190_1[0]),.doutb(w_dff_A_gHqlsMsW1_1),.doutc(w_n190_1[2]),.din(w_n190_0[0]));
	jspl3 jspl3_w_n191_0(.douta(w_n191_0[0]),.doutb(w_n191_0[1]),.doutc(w_n191_0[2]),.din(n191));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl3 jspl3_w_n196_0(.douta(w_dff_A_N10FqqUo3_0),.doutb(w_n196_0[1]),.doutc(w_n196_0[2]),.din(w_dff_B_l4X8PHtZ6_3));
	jspl3 jspl3_w_n196_1(.douta(w_n196_1[0]),.doutb(w_n196_1[1]),.doutc(w_n196_1[2]),.din(w_n196_0[0]));
	jspl3 jspl3_w_n196_2(.douta(w_dff_A_siocPJva6_0),.doutb(w_n196_2[1]),.doutc(w_dff_A_UxntVVz47_2),.din(w_n196_0[1]));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl jspl_w_n197_1(.douta(w_n197_1[0]),.doutb(w_n197_1[1]),.din(w_n197_0[0]));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.doutc(w_n199_0[2]),.din(w_dff_B_ZoCsYINS5_3));
	jspl jspl_w_n199_1(.douta(w_n199_1[0]),.doutb(w_n199_1[1]),.din(w_n199_0[0]));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(n201));
	jspl jspl_w_n205_0(.douta(w_n205_0[0]),.doutb(w_n205_0[1]),.din(w_dff_B_EGl2WplV9_2));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(n206));
	jspl3 jspl3_w_n210_0(.douta(w_n210_0[0]),.doutb(w_n210_0[1]),.doutc(w_n210_0[2]),.din(n210));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_dff_A_4d3ZXjKD6_1),.din(n213));
	jspl jspl_w_n214_0(.douta(w_n214_0[0]),.doutb(w_n214_0[1]),.din(n214));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl jspl_w_n219_0(.douta(w_dff_A_2Y721u017_0),.doutb(w_n219_0[1]),.din(n219));
	jspl3 jspl3_w_n221_0(.douta(w_dff_A_xMCwb3Xo0_0),.doutb(w_dff_A_ugZr37UL0_1),.doutc(w_n221_0[2]),.din(n221));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_dff_A_xhAvvTf95_1),.din(n228));
	jspl3 jspl3_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.doutc(w_n229_0[2]),.din(w_dff_B_lS3T56Se1_3));
	jspl jspl_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.din(n230));
	jspl3 jspl3_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.doutc(w_n231_0[2]),.din(n231));
	jspl3 jspl3_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.doutc(w_n234_0[2]),.din(n234));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.din(w_dff_B_HZzECxmh4_2));
	jspl3 jspl3_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.doutc(w_n242_0[2]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl jspl_w_n246_1(.douta(w_n246_1[0]),.doutb(w_n246_1[1]),.din(w_n246_0[0]));
	jspl jspl_w_n249_0(.douta(w_dff_A_EWkT1AOP3_0),.doutb(w_n249_0[1]),.din(w_dff_B_PT24TNez2_2));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n257_0(.douta(w_dff_A_b6fZpL3E6_0),.doutb(w_n257_0[1]),.din(n257));
	jspl jspl_w_n259_0(.douta(w_dff_A_mU3DqGOy2_0),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.doutc(w_n269_1[2]),.din(w_n269_0[0]));
	jspl jspl_w_n270_0(.douta(w_dff_A_b7wLZy7l7_0),.doutb(w_n270_0[1]),.din(w_dff_B_GHq7vOay5_2));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_dff_A_cYYAdWbW6_0),.doutb(w_n271_1[1]),.doutc(w_dff_A_RovLMnhq5_2),.din(w_n271_0[0]));
	jspl3 jspl3_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_TuWqKq408_1),.doutc(w_dff_A_OHCadVq27_2),.din(n274));
	jspl jspl_w_n278_0(.douta(w_n278_0[0]),.doutb(w_dff_A_TH2JGvDg9_1),.din(n278));
	jspl jspl_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.din(n279));
	jspl jspl_w_n281_0(.douta(w_n281_0[0]),.doutb(w_dff_A_WnxFzNr57_1),.din(n281));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n288_1(.douta(w_n288_1[0]),.doutb(w_n288_1[1]),.din(w_n288_0[0]));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_dff_A_8TdrWGBZ9_1),.din(n300));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_dff_A_8G0arO6g1_1),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_dff_A_t5wxuhce7_1),.din(n320));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n334_0(.douta(w_n334_0[0]),.doutb(w_n334_0[1]),.din(n334));
	jspl jspl_w_n339_0(.douta(w_dff_A_g7sa2qLA6_0),.doutb(w_n339_0[1]),.din(n339));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl jspl_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.din(w_n355_0[0]));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_dff_A_nP6h92hb4_1),.doutc(w_dff_A_t0iXcEPt3_2),.din(n367));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(w_dff_B_IzQrH9399_2));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.din(n372));
	jspl jspl_w_n374_0(.douta(w_n374_0[0]),.doutb(w_dff_A_aLEHXo812_1),.din(n374));
	jspl jspl_w_n381_0(.douta(w_n381_0[0]),.doutb(w_n381_0[1]),.din(n381));
	jspl3 jspl3_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.doutc(w_n382_0[2]),.din(n382));
	jspl jspl_w_n382_1(.douta(w_n382_1[0]),.doutb(w_n382_1[1]),.din(w_n382_0[0]));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl jspl_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n387_1(.douta(w_n387_1[0]),.doutb(w_n387_1[1]),.din(w_n387_0[0]));
	jspl jspl_w_n390_0(.douta(w_dff_A_ZnOsSdK38_0),.doutb(w_n390_0[1]),.din(w_dff_B_sTdKnjCs0_2));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_dff_A_cSstGaA84_1),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.doutc(w_n404_0[2]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n407_0(.douta(w_n407_0[0]),.doutb(w_dff_A_J25dw3vL9_1),.doutc(w_dff_A_MCUi8aXw4_2),.din(n407));
	jspl3 jspl3_w_n407_1(.douta(w_dff_A_8XGHsvdi4_0),.doutb(w_dff_A_dSGJppjg1_1),.doutc(w_n407_1[2]),.din(w_n407_0[0]));
	jspl jspl_w_n407_2(.douta(w_n407_2[0]),.doutb(w_n407_2[1]),.din(w_n407_0[1]));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(n412));
	jspl3 jspl3_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jspl jspl_w_n420_1(.douta(w_n420_1[0]),.doutb(w_n420_1[1]),.din(w_n420_0[0]));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_dff_A_0wOEUyzd3_1),.doutc(w_dff_A_aaUwg8TN3_2),.din(n425));
	jspl3 jspl3_w_n425_1(.douta(w_dff_A_oB09sLbt1_0),.doutb(w_dff_A_tIIMMgaG3_1),.doutc(w_n425_1[2]),.din(w_n425_0[0]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl jspl_w_n430_0(.douta(w_dff_A_oye51Lho7_0),.doutb(w_n430_0[1]),.din(w_dff_B_YFNG28sK1_2));
	jspl3 jspl3_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.doutc(w_n436_0[2]),.din(n436));
	jspl3 jspl3_w_n439_0(.douta(w_n439_0[0]),.doutb(w_dff_A_oAWWLL5M1_1),.doutc(w_n439_0[2]),.din(n439));
	jspl jspl_w_n439_1(.douta(w_n439_1[0]),.doutb(w_n439_1[1]),.din(w_n439_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_dff_A_1LTuX2rb6_1),.din(w_dff_B_Klqcwm7I2_2));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl3 jspl3_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.doutc(w_n455_0[2]),.din(n455));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(n474));
	jspl jspl_w_n475_0(.douta(w_n475_0[0]),.doutb(w_n475_0[1]),.din(n475));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_dff_A_fGoUnq7h8_1),.din(n478));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(n479));
	jspl jspl_w_n483_0(.douta(w_n483_0[0]),.doutb(w_n483_0[1]),.din(n483));
	jspl jspl_w_n484_0(.douta(w_dff_A_VTeMM7ch9_0),.doutb(w_n484_0[1]),.din(n484));
	jspl3 jspl3_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.doutc(w_n492_0[2]),.din(n492));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_dff_A_95QQxCPE3_1),.din(n511));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n516_0(.douta(w_n516_0[0]),.doutb(w_n516_0[1]),.din(n516));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(w_dff_B_t0VQJmnK4_2));
	jspl3 jspl3_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.doutc(w_n519_0[2]),.din(n519));
	jspl3 jspl3_w_n519_1(.douta(w_n519_1[0]),.doutb(w_n519_1[1]),.doutc(w_n519_1[2]),.din(w_n519_0[0]));
	jspl jspl_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_dff_A_8E9uyBLA2_1),.din(n524));
	jspl jspl_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.din(n528));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(w_dff_B_UDv9v5b98_2));
	jspl jspl_w_n534_0(.douta(w_dff_A_Gm6slROH2_0),.doutb(w_n534_0[1]),.din(n534));
	jspl3 jspl3_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.doutc(w_dff_A_ENbhoJix7_2),.din(n536));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_dff_A_jytAgkMy8_1),.din(n539));
	jspl jspl_w_n541_0(.douta(w_dff_A_KqevKNcd0_0),.doutb(w_n541_0[1]),.din(n541));
	jspl3 jspl3_w_n542_0(.douta(w_dff_A_JFkCUEOJ0_0),.doutb(w_n542_0[1]),.doutc(w_n542_0[2]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl3 jspl3_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.doutc(w_n548_0[2]),.din(w_dff_B_c69DTJYd0_3));
	jspl jspl_w_n550_0(.douta(w_n550_0[0]),.doutb(w_n550_0[1]),.din(n550));
	jspl3 jspl3_w_n552_0(.douta(w_n552_0[0]),.doutb(w_dff_A_P3wnx4oD8_1),.doutc(w_dff_A_UfVmVae33_2),.din(n552));
	jspl jspl_w_n552_1(.douta(w_n552_1[0]),.doutb(w_n552_1[1]),.din(w_n552_0[0]));
	jspl3 jspl3_w_n553_0(.douta(w_dff_A_qRayeMKr2_0),.doutb(w_n553_0[1]),.doutc(w_dff_A_YaTQG0RH8_2),.din(n553));
	jspl3 jspl3_w_n553_1(.douta(w_n553_1[0]),.doutb(w_dff_A_daKAvAwE4_1),.doutc(w_n553_1[2]),.din(w_n553_0[0]));
	jspl3 jspl3_w_n553_2(.douta(w_dff_A_NZPioaXJ2_0),.doutb(w_dff_A_vPczuf2F2_1),.doutc(w_n553_2[2]),.din(w_n553_0[1]));
	jspl3 jspl3_w_n554_0(.douta(w_dff_A_FMppqw4O3_0),.doutb(w_n554_0[1]),.doutc(w_dff_A_GIbWYEPv0_2),.din(n554));
	jspl3 jspl3_w_n554_1(.douta(w_n554_1[0]),.doutb(w_n554_1[1]),.doutc(w_n554_1[2]),.din(w_n554_0[0]));
	jspl3 jspl3_w_n554_2(.douta(w_n554_2[0]),.doutb(w_dff_A_lNlDI1Rb2_1),.doutc(w_dff_A_5Fr6r7e69_2),.din(w_n554_0[1]));
	jspl3 jspl3_w_n554_3(.douta(w_n554_3[0]),.doutb(w_n554_3[1]),.doutc(w_n554_3[2]),.din(w_n554_0[2]));
	jspl jspl_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.din(w_dff_B_vHDgTMOi9_2));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl3 jspl3_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.doutc(w_n563_0[2]),.din(w_dff_B_XoM5BIMh5_3));
	jspl jspl_w_n564_0(.douta(w_n564_0[0]),.doutb(w_n564_0[1]),.din(n564));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(w_dff_B_YLlFhacG2_2));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(n567));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_n571_0[2]),.din(n571));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_n573_0[2]),.din(n573));
	jspl3 jspl3_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.doutc(w_n576_0[2]),.din(n576));
	jspl jspl_w_n576_1(.douta(w_n576_1[0]),.doutb(w_n576_1[1]),.din(w_n576_0[0]));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_dff_A_ZB48YLv05_2),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n589_0(.douta(w_n589_0[0]),.doutb(w_n589_0[1]),.doutc(w_n589_0[2]),.din(n589));
	jspl3 jspl3_w_n589_1(.douta(w_dff_A_7F7lXBco6_0),.doutb(w_n589_1[1]),.doutc(w_n589_1[2]),.din(w_n589_0[0]));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_dff_A_DHUjSQ1X3_1),.doutc(w_dff_A_A4hFy3VS9_2),.din(n591));
	jspl jspl_w_n591_1(.douta(w_n591_1[0]),.doutb(w_n591_1[1]),.din(w_n591_0[0]));
	jspl3 jspl3_w_n592_0(.douta(w_dff_A_gdygnVVT6_0),.doutb(w_n592_0[1]),.doutc(w_dff_A_kcce7wmu0_2),.din(n592));
	jspl3 jspl3_w_n592_1(.douta(w_dff_A_UEPnqtJ47_0),.doutb(w_dff_A_t2jFqypB4_1),.doutc(w_n592_1[2]),.din(w_n592_0[0]));
	jspl jspl_w_n592_2(.douta(w_n592_2[0]),.doutb(w_n592_2[1]),.din(w_n592_0[1]));
	jspl3 jspl3_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.doutc(w_n593_0[2]),.din(n593));
	jspl jspl_w_n602_0(.douta(w_dff_A_mYqX3KMD9_0),.doutb(w_n602_0[1]),.din(n602));
	jspl3 jspl3_w_n603_0(.douta(w_dff_A_99KqSkib8_0),.doutb(w_n603_0[1]),.doutc(w_dff_A_fx8vizA06_2),.din(w_dff_B_ZJlqJ5FK5_3));
	jspl3 jspl3_w_n603_1(.douta(w_dff_A_LJEiiwrx0_0),.doutb(w_dff_A_99HJibvw4_1),.doutc(w_n603_1[2]),.din(w_n603_0[0]));
	jspl jspl_w_n603_2(.douta(w_dff_A_FYYhgysf1_0),.doutb(w_n603_2[1]),.din(w_n603_0[1]));
	jspl3 jspl3_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.doutc(w_n604_0[2]),.din(n604));
	jspl3 jspl3_w_n604_1(.douta(w_dff_A_6ULOEFua4_0),.doutb(w_n604_1[1]),.doutc(w_dff_A_eMkn6guf5_2),.din(w_n604_0[0]));
	jspl jspl_w_n604_2(.douta(w_dff_A_EHw4u9ai4_0),.doutb(w_n604_2[1]),.din(w_n604_0[1]));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_dff_A_zYsdWECT7_2),.din(w_n605_0[0]));
	jspl3 jspl3_w_n608_0(.douta(w_n608_0[0]),.doutb(w_dff_A_dICPL2Kz8_1),.doutc(w_dff_A_9x6Qr2Io4_2),.din(n608));
	jspl3 jspl3_w_n608_1(.douta(w_dff_A_Sdz9dIll5_0),.doutb(w_n608_1[1]),.doutc(w_dff_A_ohTChJrT1_2),.din(w_n608_0[0]));
	jspl3 jspl3_w_n612_0(.douta(w_n612_0[0]),.doutb(w_dff_A_NQgcz3gX4_1),.doutc(w_dff_A_seuHrhMy5_2),.din(n612));
	jspl3 jspl3_w_n612_1(.douta(w_dff_A_oTtkGiLK7_0),.doutb(w_dff_A_QCOAP4Qk2_1),.doutc(w_n612_1[2]),.din(w_n612_0[0]));
	jspl3 jspl3_w_n612_2(.douta(w_n612_2[0]),.doutb(w_n612_2[1]),.doutc(w_n612_2[2]),.din(w_n612_0[1]));
	jspl3 jspl3_w_n612_3(.douta(w_dff_A_XgI3rQ976_0),.doutb(w_n612_3[1]),.doutc(w_dff_A_tcO6s0D57_2),.din(w_n612_0[2]));
	jspl jspl_w_n612_4(.douta(w_n612_4[0]),.doutb(w_dff_A_vnEzpc403_1),.din(w_n612_1[0]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl jspl_w_n613_1(.douta(w_n613_1[0]),.doutb(w_n613_1[1]),.din(w_n613_0[0]));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_dff_A_DU6dpN675_1),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl3 jspl3_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.doutc(w_n617_1[2]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n617_2(.douta(w_n617_2[0]),.doutb(w_n617_2[1]),.doutc(w_n617_2[2]),.din(w_n617_0[1]));
	jspl3 jspl3_w_n617_3(.douta(w_n617_3[0]),.doutb(w_n617_3[1]),.doutc(w_n617_3[2]),.din(w_n617_0[2]));
	jspl3 jspl3_w_n617_4(.douta(w_n617_4[0]),.doutb(w_n617_4[1]),.doutc(w_n617_4[2]),.din(w_n617_1[0]));
	jspl3 jspl3_w_n617_5(.douta(w_n617_5[0]),.doutb(w_n617_5[1]),.doutc(w_n617_5[2]),.din(w_n617_1[1]));
	jspl jspl_w_n617_6(.douta(w_n617_6[0]),.doutb(w_n617_6[1]),.din(w_n617_1[2]));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_dff_A_Y8KSfdHb2_1),.din(n622));
	jspl3 jspl3_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.doutc(w_n623_0[2]),.din(n623));
	jspl3 jspl3_w_n623_1(.douta(w_n623_1[0]),.doutb(w_n623_1[1]),.doutc(w_n623_1[2]),.din(w_n623_0[0]));
	jspl3 jspl3_w_n623_2(.douta(w_n623_2[0]),.doutb(w_n623_2[1]),.doutc(w_n623_2[2]),.din(w_n623_0[1]));
	jspl3 jspl3_w_n623_3(.douta(w_n623_3[0]),.doutb(w_n623_3[1]),.doutc(w_n623_3[2]),.din(w_n623_0[2]));
	jspl3 jspl3_w_n623_4(.douta(w_n623_4[0]),.doutb(w_n623_4[1]),.doutc(w_n623_4[2]),.din(w_n623_1[0]));
	jspl jspl_w_n623_5(.douta(w_n623_5[0]),.doutb(w_n623_5[1]),.din(w_n623_1[1]));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(n626));
	jspl3 jspl3_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.doutc(w_n627_0[2]),.din(n627));
	jspl3 jspl3_w_n627_1(.douta(w_n627_1[0]),.doutb(w_n627_1[1]),.doutc(w_n627_1[2]),.din(w_n627_0[0]));
	jspl3 jspl3_w_n627_2(.douta(w_n627_2[0]),.doutb(w_n627_2[1]),.doutc(w_n627_2[2]),.din(w_n627_0[1]));
	jspl3 jspl3_w_n627_3(.douta(w_n627_3[0]),.doutb(w_n627_3[1]),.doutc(w_n627_3[2]),.din(w_n627_0[2]));
	jspl3 jspl3_w_n627_4(.douta(w_n627_4[0]),.doutb(w_n627_4[1]),.doutc(w_n627_4[2]),.din(w_n627_1[0]));
	jspl3 jspl3_w_n627_5(.douta(w_n627_5[0]),.doutb(w_n627_5[1]),.doutc(w_n627_5[2]),.din(w_n627_1[1]));
	jspl3 jspl3_w_n627_6(.douta(w_n627_6[0]),.doutb(w_n627_6[1]),.doutc(w_n627_6[2]),.din(w_n627_1[2]));
	jspl jspl_w_n627_7(.douta(w_n627_7[0]),.doutb(w_n627_7[1]),.din(w_n627_2[0]));
	jspl3 jspl3_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.doutc(w_n631_0[2]),.din(n631));
	jspl3 jspl3_w_n631_1(.douta(w_n631_1[0]),.doutb(w_n631_1[1]),.doutc(w_n631_1[2]),.din(w_n631_0[0]));
	jspl3 jspl3_w_n631_2(.douta(w_n631_2[0]),.doutb(w_n631_2[1]),.doutc(w_n631_2[2]),.din(w_n631_0[1]));
	jspl3 jspl3_w_n631_3(.douta(w_n631_3[0]),.doutb(w_n631_3[1]),.doutc(w_n631_3[2]),.din(w_n631_0[2]));
	jspl3 jspl3_w_n631_4(.douta(w_n631_4[0]),.doutb(w_n631_4[1]),.doutc(w_n631_4[2]),.din(w_n631_1[0]));
	jspl3 jspl3_w_n631_5(.douta(w_n631_5[0]),.doutb(w_n631_5[1]),.doutc(w_n631_5[2]),.din(w_n631_1[1]));
	jspl3 jspl3_w_n631_6(.douta(w_n631_6[0]),.doutb(w_n631_6[1]),.doutc(w_n631_6[2]),.din(w_n631_1[2]));
	jspl jspl_w_n631_7(.douta(w_n631_7[0]),.doutb(w_n631_7[1]),.din(w_n631_2[0]));
	jspl3 jspl3_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.doutc(w_n634_0[2]),.din(n634));
	jspl3 jspl3_w_n634_1(.douta(w_n634_1[0]),.doutb(w_n634_1[1]),.doutc(w_n634_1[2]),.din(w_n634_0[0]));
	jspl3 jspl3_w_n634_2(.douta(w_n634_2[0]),.doutb(w_n634_2[1]),.doutc(w_n634_2[2]),.din(w_n634_0[1]));
	jspl3 jspl3_w_n634_3(.douta(w_n634_3[0]),.doutb(w_n634_3[1]),.doutc(w_n634_3[2]),.din(w_n634_0[2]));
	jspl jspl_w_n634_4(.douta(w_n634_4[0]),.doutb(w_n634_4[1]),.din(w_n634_1[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl3 jspl3_w_n636_1(.douta(w_n636_1[0]),.doutb(w_n636_1[1]),.doutc(w_n636_1[2]),.din(w_n636_0[0]));
	jspl3 jspl3_w_n636_2(.douta(w_n636_2[0]),.doutb(w_n636_2[1]),.doutc(w_n636_2[2]),.din(w_n636_0[1]));
	jspl3 jspl3_w_n636_3(.douta(w_n636_3[0]),.doutb(w_n636_3[1]),.doutc(w_n636_3[2]),.din(w_n636_0[2]));
	jspl3 jspl3_w_n636_4(.douta(w_n636_4[0]),.doutb(w_n636_4[1]),.doutc(w_n636_4[2]),.din(w_n636_1[0]));
	jspl3 jspl3_w_n636_5(.douta(w_n636_5[0]),.doutb(w_n636_5[1]),.doutc(w_n636_5[2]),.din(w_n636_1[1]));
	jspl3 jspl3_w_n636_6(.douta(w_n636_6[0]),.doutb(w_n636_6[1]),.doutc(w_n636_6[2]),.din(w_n636_1[2]));
	jspl jspl_w_n636_7(.douta(w_n636_7[0]),.doutb(w_n636_7[1]),.din(w_n636_2[0]));
	jspl jspl_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.din(n639));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl3 jspl3_w_n640_2(.douta(w_n640_2[0]),.doutb(w_n640_2[1]),.doutc(w_n640_2[2]),.din(w_n640_0[1]));
	jspl3 jspl3_w_n640_3(.douta(w_n640_3[0]),.doutb(w_n640_3[1]),.doutc(w_n640_3[2]),.din(w_n640_0[2]));
	jspl3 jspl3_w_n640_4(.douta(w_n640_4[0]),.doutb(w_n640_4[1]),.doutc(w_n640_4[2]),.din(w_n640_1[0]));
	jspl3 jspl3_w_n640_5(.douta(w_n640_5[0]),.doutb(w_n640_5[1]),.doutc(w_n640_5[2]),.din(w_n640_1[1]));
	jspl3 jspl3_w_n640_6(.douta(w_n640_6[0]),.doutb(w_n640_6[1]),.doutc(w_n640_6[2]),.din(w_n640_1[2]));
	jspl jspl_w_n640_7(.douta(w_n640_7[0]),.doutb(w_n640_7[1]),.din(w_n640_2[0]));
	jspl3 jspl3_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.doutc(w_n642_0[2]),.din(n642));
	jspl3 jspl3_w_n642_1(.douta(w_n642_1[0]),.doutb(w_n642_1[1]),.doutc(w_n642_1[2]),.din(w_n642_0[0]));
	jspl3 jspl3_w_n642_2(.douta(w_n642_2[0]),.doutb(w_n642_2[1]),.doutc(w_n642_2[2]),.din(w_n642_0[1]));
	jspl3 jspl3_w_n642_3(.douta(w_n642_3[0]),.doutb(w_n642_3[1]),.doutc(w_n642_3[2]),.din(w_n642_0[2]));
	jspl3 jspl3_w_n642_4(.douta(w_n642_4[0]),.doutb(w_n642_4[1]),.doutc(w_n642_4[2]),.din(w_n642_1[0]));
	jspl3 jspl3_w_n642_5(.douta(w_n642_5[0]),.doutb(w_n642_5[1]),.doutc(w_n642_5[2]),.din(w_n642_1[1]));
	jspl3 jspl3_w_n642_6(.douta(w_n642_6[0]),.doutb(w_n642_6[1]),.doutc(w_n642_6[2]),.din(w_n642_1[2]));
	jspl jspl_w_n642_7(.douta(w_n642_7[0]),.doutb(w_n642_7[1]),.din(w_n642_2[0]));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(n654));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl3 jspl3_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.doutc(w_dff_A_88dtetgu2_2),.din(n672));
	jspl jspl_w_n672_1(.douta(w_n672_1[0]),.doutb(w_dff_A_RtHqXjHw8_1),.din(w_n672_0[0]));
	jspl3 jspl3_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.doutc(w_n675_0[2]),.din(n675));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(w_dff_B_Ivzg3xIC2_2));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_dff_A_tibR6DAP5_1),.din(w_dff_B_eElI0crC8_2));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_dff_A_Osu92vvW7_1),.doutc(w_n696_0[2]),.din(n696));
	jspl3 jspl3_w_n696_1(.douta(w_dff_A_9ralKSB82_0),.doutb(w_n696_1[1]),.doutc(w_dff_A_zYqiFtf66_2),.din(w_n696_0[0]));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.doutc(w_n743_0[2]),.din(n743));
	jspl jspl_w_n743_1(.douta(w_n743_1[0]),.doutb(w_n743_1[1]),.din(w_n743_0[0]));
	jspl jspl_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl3 jspl3_w_n758_0(.douta(w_n758_0[0]),.doutb(w_dff_A_LqppROXH2_1),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n758_1(.douta(w_n758_1[0]),.doutb(w_dff_A_2huqbXvQ3_1),.din(w_n758_0[0]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_dff_A_MKuYlg0D3_0),.doutb(w_n760_0[1]),.din(n760));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_dff_A_DPRKpDgj8_2),.din(n764));
	jspl3 jspl3_w_n764_1(.douta(w_n764_1[0]),.doutb(w_n764_1[1]),.doutc(w_dff_A_pdmCXQak7_2),.din(w_n764_0[0]));
	jspl jspl_w_n769_0(.douta(w_dff_A_kcaawKiK3_0),.doutb(w_n769_0[1]),.din(n769));
	jspl3 jspl3_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.doutc(w_n771_0[2]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.din(n779));
	jspl jspl_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.din(n797));
	jspl jspl_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.din(n801));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n825_0(.douta(w_n825_0[0]),.doutb(w_n825_0[1]),.din(n825));
	jspl3 jspl3_w_n853_0(.douta(w_n853_0[0]),.doutb(w_dff_A_Ba2yrQhG0_1),.doutc(w_n853_0[2]),.din(n853));
	jspl3 jspl3_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.doutc(w_n855_0[2]),.din(n855));
	jspl3 jspl3_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.doutc(w_n861_0[2]),.din(n861));
	jspl jspl_w_n861_1(.douta(w_n861_1[0]),.doutb(w_n861_1[1]),.din(w_n861_0[0]));
	jspl jspl_w_n863_0(.douta(w_n863_0[0]),.doutb(w_dff_A_70LQrWZs1_1),.din(n863));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.din(n899));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl3 jspl3_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.doutc(w_n937_0[2]),.din(n937));
	jspl jspl_w_n940_0(.douta(w_n940_0[0]),.doutb(w_dff_A_y3dUgMXB2_1),.din(n940));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.doutc(w_n988_0[2]),.din(n988));
	jspl jspl_w_n990_0(.douta(w_n990_0[0]),.doutb(w_dff_A_jYgrIUsq7_1),.din(n990));
	jspl3 jspl3_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.doutc(w_n991_0[2]),.din(n991));
	jspl jspl_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.din(n992));
	jspl3 jspl3_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.doutc(w_n994_0[2]),.din(n994));
	jspl3 jspl3_w_n996_0(.douta(w_dff_A_k3JGA4C40_0),.doutb(w_n996_0[1]),.doutc(w_dff_A_4NmqG9wv9_2),.din(n996));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_dff_A_eAk7lmmX5_1),.din(n999));
	jspl3 jspl3_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.doutc(w_n1001_0[2]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_dff_A_4Oz5YSYp3_1),.doutc(w_dff_A_zob0P3cI5_2),.din(n1002));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl3 jspl3_w_n1049_0(.douta(w_dff_A_oSt1N62k5_0),.doutb(w_dff_A_4T6D0jPq0_1),.doutc(w_n1049_0[2]),.din(n1049));
	jspl jspl_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_dff_A_RBGIcHEi1_1),.din(n1057));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(n1059));
	jspl jspl_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.din(n1088));
	jspl3 jspl3_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.doutc(w_n1114_0[2]),.din(n1114));
	jspl3 jspl3_w_n1162_0(.douta(w_n1162_0[0]),.doutb(w_n1162_0[1]),.doutc(w_n1162_0[2]),.din(n1162));
	jspl jspl_w_n1164_0(.douta(w_n1164_0[0]),.doutb(w_dff_A_ZB9CuM7a7_1),.din(n1164));
	jspl jspl_w_n1172_0(.douta(w_n1172_0[0]),.doutb(w_n1172_0[1]),.din(n1172));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_dff_A_FkbKZ3nL0_1),.din(n1175));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(n1183));
	jspl jspl_w_n1184_0(.douta(w_dff_A_SNPNU4NY5_0),.doutb(w_n1184_0[1]),.din(n1184));
	jspl jspl_w_n1187_0(.douta(w_dff_A_1tqHPfDU0_0),.doutb(w_n1187_0[1]),.din(n1187));
	jdff dff_B_DHAEC3iB8_1(.din(n111),.dout(w_dff_B_DHAEC3iB8_1),.clk(gclk));
	jdff dff_B_b8xM2L0C0_1(.din(w_dff_B_DHAEC3iB8_1),.dout(w_dff_B_b8xM2L0C0_1),.clk(gclk));
	jdff dff_B_2uIT0MVQ7_0(.din(n126),.dout(w_dff_B_2uIT0MVQ7_0),.clk(gclk));
	jdff dff_B_9UNlZxYu7_0(.din(n125),.dout(w_dff_B_9UNlZxYu7_0),.clk(gclk));
	jdff dff_B_g1FTjHUN6_0(.din(w_dff_B_9UNlZxYu7_0),.dout(w_dff_B_g1FTjHUN6_0),.clk(gclk));
	jdff dff_A_DG2xMPmt0_1(.dout(w_n72_1[1]),.din(w_dff_A_DG2xMPmt0_1),.clk(gclk));
	jdff dff_A_SxUhH09K8_1(.dout(w_dff_A_DG2xMPmt0_1),.din(w_dff_A_SxUhH09K8_1),.clk(gclk));
	jdff dff_A_coblnMg10_0(.dout(w_n98_2[0]),.din(w_dff_A_coblnMg10_0),.clk(gclk));
	jdff dff_B_Do0q7fth3_0(.din(n597),.dout(w_dff_B_Do0q7fth3_0),.clk(gclk));
	jdff dff_B_SXT2Zkzf9_0(.din(w_dff_B_Do0q7fth3_0),.dout(w_dff_B_SXT2Zkzf9_0),.clk(gclk));
	jdff dff_B_CjykkLot3_0(.din(w_dff_B_SXT2Zkzf9_0),.dout(w_dff_B_CjykkLot3_0),.clk(gclk));
	jdff dff_B_Rv7m2esg3_0(.din(w_dff_B_CjykkLot3_0),.dout(w_dff_B_Rv7m2esg3_0),.clk(gclk));
	jdff dff_B_LfoSC3jf1_0(.din(w_dff_B_Rv7m2esg3_0),.dout(w_dff_B_LfoSC3jf1_0),.clk(gclk));
	jdff dff_B_RwFA02SY6_0(.din(w_dff_B_LfoSC3jf1_0),.dout(w_dff_B_RwFA02SY6_0),.clk(gclk));
	jdff dff_B_woz0rSSW2_0(.din(w_dff_B_RwFA02SY6_0),.dout(w_dff_B_woz0rSSW2_0),.clk(gclk));
	jdff dff_B_am17GXv75_0(.din(n596),.dout(w_dff_B_am17GXv75_0),.clk(gclk));
	jdff dff_B_lGxr1js75_0(.din(n795),.dout(w_dff_B_lGxr1js75_0),.clk(gclk));
	jdff dff_B_Zzk3xV260_0(.din(w_dff_B_lGxr1js75_0),.dout(w_dff_B_Zzk3xV260_0),.clk(gclk));
	jdff dff_B_5iecDHWU5_0(.din(w_dff_B_Zzk3xV260_0),.dout(w_dff_B_5iecDHWU5_0),.clk(gclk));
	jdff dff_B_BLQN1P1U3_0(.din(w_dff_B_5iecDHWU5_0),.dout(w_dff_B_BLQN1P1U3_0),.clk(gclk));
	jdff dff_B_8vJb4fPa7_0(.din(w_dff_B_BLQN1P1U3_0),.dout(w_dff_B_8vJb4fPa7_0),.clk(gclk));
	jdff dff_B_GyZEmpwB0_0(.din(w_dff_B_8vJb4fPa7_0),.dout(w_dff_B_GyZEmpwB0_0),.clk(gclk));
	jdff dff_B_XiO6N5Wh8_0(.din(w_dff_B_GyZEmpwB0_0),.dout(w_dff_B_XiO6N5Wh8_0),.clk(gclk));
	jdff dff_B_UQtWAT099_0(.din(w_dff_B_XiO6N5Wh8_0),.dout(w_dff_B_UQtWAT099_0),.clk(gclk));
	jdff dff_B_ZgwDnQ3j1_0(.din(w_dff_B_UQtWAT099_0),.dout(w_dff_B_ZgwDnQ3j1_0),.clk(gclk));
	jdff dff_B_8xEtBd4k8_0(.din(w_dff_B_ZgwDnQ3j1_0),.dout(w_dff_B_8xEtBd4k8_0),.clk(gclk));
	jdff dff_B_6uvlk9mH3_0(.din(w_dff_B_8xEtBd4k8_0),.dout(w_dff_B_6uvlk9mH3_0),.clk(gclk));
	jdff dff_B_8rIhmINw8_0(.din(w_dff_B_6uvlk9mH3_0),.dout(w_dff_B_8rIhmINw8_0),.clk(gclk));
	jdff dff_B_6r4cWHNH7_0(.din(w_dff_B_8rIhmINw8_0),.dout(w_dff_B_6r4cWHNH7_0),.clk(gclk));
	jdff dff_B_xSUxJVYv1_1(.din(n791),.dout(w_dff_B_xSUxJVYv1_1),.clk(gclk));
	jdff dff_B_YHtyzqau1_0(.din(n793),.dout(w_dff_B_YHtyzqau1_0),.clk(gclk));
	jdff dff_B_ddEVRQ7Q7_0(.din(n784),.dout(w_dff_B_ddEVRQ7Q7_0),.clk(gclk));
	jdff dff_B_3zoO6mt01_0(.din(w_dff_B_ddEVRQ7Q7_0),.dout(w_dff_B_3zoO6mt01_0),.clk(gclk));
	jdff dff_B_6WTVwIh96_0(.din(w_dff_B_3zoO6mt01_0),.dout(w_dff_B_6WTVwIh96_0),.clk(gclk));
	jdff dff_B_yVv8qJii1_0(.din(w_dff_B_6WTVwIh96_0),.dout(w_dff_B_yVv8qJii1_0),.clk(gclk));
	jdff dff_B_EFp0z5Qb6_0(.din(w_dff_B_yVv8qJii1_0),.dout(w_dff_B_EFp0z5Qb6_0),.clk(gclk));
	jdff dff_B_2R0WsyJF7_0(.din(w_dff_B_EFp0z5Qb6_0),.dout(w_dff_B_2R0WsyJF7_0),.clk(gclk));
	jdff dff_B_IsbI2Fv12_0(.din(w_dff_B_2R0WsyJF7_0),.dout(w_dff_B_IsbI2Fv12_0),.clk(gclk));
	jdff dff_B_p139BhB06_0(.din(w_dff_B_IsbI2Fv12_0),.dout(w_dff_B_p139BhB06_0),.clk(gclk));
	jdff dff_B_0msDaU7S8_0(.din(w_dff_B_p139BhB06_0),.dout(w_dff_B_0msDaU7S8_0),.clk(gclk));
	jdff dff_B_gmGWpgta5_0(.din(w_dff_B_0msDaU7S8_0),.dout(w_dff_B_gmGWpgta5_0),.clk(gclk));
	jdff dff_B_viTl6LRz7_0(.din(w_dff_B_gmGWpgta5_0),.dout(w_dff_B_viTl6LRz7_0),.clk(gclk));
	jdff dff_A_3F4ytKjn2_1(.dout(w_n116_0[1]),.din(w_dff_A_3F4ytKjn2_1),.clk(gclk));
	jdff dff_A_7X6XhEQy8_1(.dout(w_dff_A_3F4ytKjn2_1),.din(w_dff_A_7X6XhEQy8_1),.clk(gclk));
	jdff dff_B_v3w7Yg228_2(.din(n116),.dout(w_dff_B_v3w7Yg228_2),.clk(gclk));
	jdff dff_B_275f0nXt2_2(.din(w_dff_B_v3w7Yg228_2),.dout(w_dff_B_275f0nXt2_2),.clk(gclk));
	jdff dff_B_7L91uwTL8_1(.din(n774),.dout(w_dff_B_7L91uwTL8_1),.clk(gclk));
	jdff dff_B_YhXlXGjR9_0(.din(n1177),.dout(w_dff_B_YhXlXGjR9_0),.clk(gclk));
	jdff dff_B_qXD20aTC1_0(.din(w_dff_B_YhXlXGjR9_0),.dout(w_dff_B_qXD20aTC1_0),.clk(gclk));
	jdff dff_B_nJR4TUuY1_1(.din(n1174),.dout(w_dff_B_nJR4TUuY1_1),.clk(gclk));
	jdff dff_B_OTU63Woc9_1(.din(w_dff_B_nJR4TUuY1_1),.dout(w_dff_B_OTU63Woc9_1),.clk(gclk));
	jdff dff_B_0RTIB2M20_1(.din(w_dff_B_OTU63Woc9_1),.dout(w_dff_B_0RTIB2M20_1),.clk(gclk));
	jdff dff_B_4JaqEF1c5_1(.din(w_dff_B_0RTIB2M20_1),.dout(w_dff_B_4JaqEF1c5_1),.clk(gclk));
	jdff dff_B_lIiPeFPn9_1(.din(w_dff_B_4JaqEF1c5_1),.dout(w_dff_B_lIiPeFPn9_1),.clk(gclk));
	jdff dff_B_vPH0PPW99_1(.din(w_dff_B_lIiPeFPn9_1),.dout(w_dff_B_vPH0PPW99_1),.clk(gclk));
	jdff dff_B_oib0qwZT8_1(.din(w_dff_B_vPH0PPW99_1),.dout(w_dff_B_oib0qwZT8_1),.clk(gclk));
	jdff dff_B_qAQ9g4tO3_1(.din(w_dff_B_oib0qwZT8_1),.dout(w_dff_B_qAQ9g4tO3_1),.clk(gclk));
	jdff dff_B_aMA0gFRn7_1(.din(w_dff_B_qAQ9g4tO3_1),.dout(w_dff_B_aMA0gFRn7_1),.clk(gclk));
	jdff dff_B_EfcMgCN70_1(.din(w_dff_B_aMA0gFRn7_1),.dout(w_dff_B_EfcMgCN70_1),.clk(gclk));
	jdff dff_B_Xga7WSDe7_1(.din(w_dff_B_EfcMgCN70_1),.dout(w_dff_B_Xga7WSDe7_1),.clk(gclk));
	jdff dff_B_MYBZoQKU8_1(.din(w_dff_B_Xga7WSDe7_1),.dout(w_dff_B_MYBZoQKU8_1),.clk(gclk));
	jdff dff_B_4FzlR2na7_1(.din(w_dff_B_MYBZoQKU8_1),.dout(w_dff_B_4FzlR2na7_1),.clk(gclk));
	jdff dff_B_XlJT3dCH2_1(.din(w_dff_B_4FzlR2na7_1),.dout(w_dff_B_XlJT3dCH2_1),.clk(gclk));
	jdff dff_B_VreLHDTh9_1(.din(w_dff_B_XlJT3dCH2_1),.dout(w_dff_B_VreLHDTh9_1),.clk(gclk));
	jdff dff_B_swXRbEuM8_1(.din(w_dff_B_VreLHDTh9_1),.dout(w_dff_B_swXRbEuM8_1),.clk(gclk));
	jdff dff_B_x6SqzwPE6_1(.din(w_dff_B_swXRbEuM8_1),.dout(w_dff_B_x6SqzwPE6_1),.clk(gclk));
	jdff dff_B_iH2R0TEF9_1(.din(w_dff_B_x6SqzwPE6_1),.dout(w_dff_B_iH2R0TEF9_1),.clk(gclk));
	jdff dff_B_qSUeiPR88_1(.din(w_dff_B_iH2R0TEF9_1),.dout(w_dff_B_qSUeiPR88_1),.clk(gclk));
	jdff dff_B_E3buoyro4_1(.din(w_dff_B_qSUeiPR88_1),.dout(w_dff_B_E3buoyro4_1),.clk(gclk));
	jdff dff_B_jOlsJFD18_1(.din(n1165),.dout(w_dff_B_jOlsJFD18_1),.clk(gclk));
	jdff dff_B_MSqVh61v9_1(.din(w_dff_B_jOlsJFD18_1),.dout(w_dff_B_MSqVh61v9_1),.clk(gclk));
	jdff dff_B_zYBwZ9ov3_1(.din(w_dff_B_MSqVh61v9_1),.dout(w_dff_B_zYBwZ9ov3_1),.clk(gclk));
	jdff dff_B_7yE3ZTQq0_0(.din(n1169),.dout(w_dff_B_7yE3ZTQq0_0),.clk(gclk));
	jdff dff_B_qDjqAWub7_0(.din(w_dff_B_7yE3ZTQq0_0),.dout(w_dff_B_qDjqAWub7_0),.clk(gclk));
	jdff dff_B_dFQcz4hf7_1(.din(n1166),.dout(w_dff_B_dFQcz4hf7_1),.clk(gclk));
	jdff dff_A_axV8nzVZ2_1(.dout(w_n1164_0[1]),.din(w_dff_A_axV8nzVZ2_1),.clk(gclk));
	jdff dff_A_ZB9CuM7a7_1(.dout(w_dff_A_axV8nzVZ2_1),.din(w_dff_A_ZB9CuM7a7_1),.clk(gclk));
	jdff dff_B_jlaeAtZl5_0(.din(n1189),.dout(w_dff_B_jlaeAtZl5_0),.clk(gclk));
	jdff dff_B_QQ5iB8JH2_1(.din(n1186),.dout(w_dff_B_QQ5iB8JH2_1),.clk(gclk));
	jdff dff_B_EU3V5uT80_1(.din(w_dff_B_QQ5iB8JH2_1),.dout(w_dff_B_EU3V5uT80_1),.clk(gclk));
	jdff dff_B_5XShQJNG7_1(.din(w_dff_B_EU3V5uT80_1),.dout(w_dff_B_5XShQJNG7_1),.clk(gclk));
	jdff dff_B_ohfCSEmq4_1(.din(w_dff_B_5XShQJNG7_1),.dout(w_dff_B_ohfCSEmq4_1),.clk(gclk));
	jdff dff_B_vJ7uPold1_1(.din(w_dff_B_ohfCSEmq4_1),.dout(w_dff_B_vJ7uPold1_1),.clk(gclk));
	jdff dff_B_7nmmNPuO6_1(.din(w_dff_B_vJ7uPold1_1),.dout(w_dff_B_7nmmNPuO6_1),.clk(gclk));
	jdff dff_B_3wfFTdZH3_1(.din(w_dff_B_7nmmNPuO6_1),.dout(w_dff_B_3wfFTdZH3_1),.clk(gclk));
	jdff dff_B_IBcbFj835_1(.din(w_dff_B_3wfFTdZH3_1),.dout(w_dff_B_IBcbFj835_1),.clk(gclk));
	jdff dff_B_jA950uW67_1(.din(w_dff_B_IBcbFj835_1),.dout(w_dff_B_jA950uW67_1),.clk(gclk));
	jdff dff_B_neeRJMWu1_1(.din(w_dff_B_jA950uW67_1),.dout(w_dff_B_neeRJMWu1_1),.clk(gclk));
	jdff dff_B_jB6Qb3vE6_1(.din(w_dff_B_neeRJMWu1_1),.dout(w_dff_B_jB6Qb3vE6_1),.clk(gclk));
	jdff dff_B_MyC8Sz9c4_1(.din(w_dff_B_jB6Qb3vE6_1),.dout(w_dff_B_MyC8Sz9c4_1),.clk(gclk));
	jdff dff_B_skgu4IkI5_1(.din(w_dff_B_MyC8Sz9c4_1),.dout(w_dff_B_skgu4IkI5_1),.clk(gclk));
	jdff dff_B_1dbtavxL3_1(.din(w_dff_B_skgu4IkI5_1),.dout(w_dff_B_1dbtavxL3_1),.clk(gclk));
	jdff dff_B_wFuoGVLd6_1(.din(w_dff_B_1dbtavxL3_1),.dout(w_dff_B_wFuoGVLd6_1),.clk(gclk));
	jdff dff_B_ge0Jm1SX5_1(.din(w_dff_B_wFuoGVLd6_1),.dout(w_dff_B_ge0Jm1SX5_1),.clk(gclk));
	jdff dff_B_KSktY4Mr6_1(.din(w_dff_B_ge0Jm1SX5_1),.dout(w_dff_B_KSktY4Mr6_1),.clk(gclk));
	jdff dff_B_giFrDIQ60_1(.din(G2897),.dout(w_dff_B_giFrDIQ60_1),.clk(gclk));
	jdff dff_B_JpAbbAiP6_1(.din(w_dff_B_giFrDIQ60_1),.dout(w_dff_B_JpAbbAiP6_1),.clk(gclk));
	jdff dff_B_qN8Zq43O3_1(.din(w_dff_B_JpAbbAiP6_1),.dout(w_dff_B_qN8Zq43O3_1),.clk(gclk));
	jdff dff_A_i9VBFY5u4_0(.dout(w_n1184_0[0]),.din(w_dff_A_i9VBFY5u4_0),.clk(gclk));
	jdff dff_A_ScFWRy543_0(.dout(w_dff_A_i9VBFY5u4_0),.din(w_dff_A_ScFWRy543_0),.clk(gclk));
	jdff dff_A_wN0MeD2T1_0(.dout(w_dff_A_ScFWRy543_0),.din(w_dff_A_wN0MeD2T1_0),.clk(gclk));
	jdff dff_A_tyCRgCWs0_0(.dout(w_dff_A_wN0MeD2T1_0),.din(w_dff_A_tyCRgCWs0_0),.clk(gclk));
	jdff dff_A_fzE37sTl9_0(.dout(w_dff_A_tyCRgCWs0_0),.din(w_dff_A_fzE37sTl9_0),.clk(gclk));
	jdff dff_A_diJK79s32_0(.dout(w_dff_A_fzE37sTl9_0),.din(w_dff_A_diJK79s32_0),.clk(gclk));
	jdff dff_A_ZRBmkMcL9_0(.dout(w_dff_A_diJK79s32_0),.din(w_dff_A_ZRBmkMcL9_0),.clk(gclk));
	jdff dff_A_Qe1V0Qmd0_0(.dout(w_dff_A_ZRBmkMcL9_0),.din(w_dff_A_Qe1V0Qmd0_0),.clk(gclk));
	jdff dff_A_br9i2ZRP9_0(.dout(w_dff_A_Qe1V0Qmd0_0),.din(w_dff_A_br9i2ZRP9_0),.clk(gclk));
	jdff dff_A_ZKZiG02d1_0(.dout(w_dff_A_br9i2ZRP9_0),.din(w_dff_A_ZKZiG02d1_0),.clk(gclk));
	jdff dff_A_IETcTTfq4_0(.dout(w_dff_A_ZKZiG02d1_0),.din(w_dff_A_IETcTTfq4_0),.clk(gclk));
	jdff dff_A_c72uh5Dh5_0(.dout(w_dff_A_IETcTTfq4_0),.din(w_dff_A_c72uh5Dh5_0),.clk(gclk));
	jdff dff_A_fpkJl5oY0_0(.dout(w_dff_A_c72uh5Dh5_0),.din(w_dff_A_fpkJl5oY0_0),.clk(gclk));
	jdff dff_A_UC608D3n8_0(.dout(w_dff_A_fpkJl5oY0_0),.din(w_dff_A_UC608D3n8_0),.clk(gclk));
	jdff dff_A_1OGrNmsG1_0(.dout(w_dff_A_UC608D3n8_0),.din(w_dff_A_1OGrNmsG1_0),.clk(gclk));
	jdff dff_A_sjn0rE7i7_0(.dout(w_dff_A_1OGrNmsG1_0),.din(w_dff_A_sjn0rE7i7_0),.clk(gclk));
	jdff dff_A_419wEkZg0_0(.dout(w_dff_A_sjn0rE7i7_0),.din(w_dff_A_419wEkZg0_0),.clk(gclk));
	jdff dff_A_SNPNU4NY5_0(.dout(w_dff_A_419wEkZg0_0),.din(w_dff_A_SNPNU4NY5_0),.clk(gclk));
	jdff dff_A_unXJm4cd3_1(.dout(w_n1175_0[1]),.din(w_dff_A_unXJm4cd3_1),.clk(gclk));
	jdff dff_A_zPvoXHja7_1(.dout(w_dff_A_unXJm4cd3_1),.din(w_dff_A_zPvoXHja7_1),.clk(gclk));
	jdff dff_A_AfvXZFmK6_1(.dout(w_dff_A_zPvoXHja7_1),.din(w_dff_A_AfvXZFmK6_1),.clk(gclk));
	jdff dff_A_tg6YtNyX5_1(.dout(w_dff_A_AfvXZFmK6_1),.din(w_dff_A_tg6YtNyX5_1),.clk(gclk));
	jdff dff_A_75T7SG8l5_1(.dout(w_dff_A_tg6YtNyX5_1),.din(w_dff_A_75T7SG8l5_1),.clk(gclk));
	jdff dff_A_51XrHNuY4_1(.dout(w_dff_A_75T7SG8l5_1),.din(w_dff_A_51XrHNuY4_1),.clk(gclk));
	jdff dff_A_XswJi0N46_1(.dout(w_dff_A_51XrHNuY4_1),.din(w_dff_A_XswJi0N46_1),.clk(gclk));
	jdff dff_A_vtVyJxbu1_1(.dout(w_dff_A_XswJi0N46_1),.din(w_dff_A_vtVyJxbu1_1),.clk(gclk));
	jdff dff_A_kzuXZDQ53_1(.dout(w_dff_A_vtVyJxbu1_1),.din(w_dff_A_kzuXZDQ53_1),.clk(gclk));
	jdff dff_A_0eHIxcLM5_1(.dout(w_dff_A_kzuXZDQ53_1),.din(w_dff_A_0eHIxcLM5_1),.clk(gclk));
	jdff dff_A_dF4gTrH22_1(.dout(w_dff_A_0eHIxcLM5_1),.din(w_dff_A_dF4gTrH22_1),.clk(gclk));
	jdff dff_A_yFkfepWh6_1(.dout(w_dff_A_dF4gTrH22_1),.din(w_dff_A_yFkfepWh6_1),.clk(gclk));
	jdff dff_A_l2EdIA8Y0_1(.dout(w_dff_A_yFkfepWh6_1),.din(w_dff_A_l2EdIA8Y0_1),.clk(gclk));
	jdff dff_A_vI6arzXl0_1(.dout(w_dff_A_l2EdIA8Y0_1),.din(w_dff_A_vI6arzXl0_1),.clk(gclk));
	jdff dff_A_Tj62m3oB8_1(.dout(w_dff_A_vI6arzXl0_1),.din(w_dff_A_Tj62m3oB8_1),.clk(gclk));
	jdff dff_A_BYOx4pAQ6_1(.dout(w_dff_A_Tj62m3oB8_1),.din(w_dff_A_BYOx4pAQ6_1),.clk(gclk));
	jdff dff_A_Kt8qZ9wz2_1(.dout(w_dff_A_BYOx4pAQ6_1),.din(w_dff_A_Kt8qZ9wz2_1),.clk(gclk));
	jdff dff_A_ZHLQcGmu8_1(.dout(w_dff_A_Kt8qZ9wz2_1),.din(w_dff_A_ZHLQcGmu8_1),.clk(gclk));
	jdff dff_A_FkbKZ3nL0_1(.dout(w_dff_A_ZHLQcGmu8_1),.din(w_dff_A_FkbKZ3nL0_1),.clk(gclk));
	jdff dff_A_QNhc1giV7_0(.dout(w_n1187_0[0]),.din(w_dff_A_QNhc1giV7_0),.clk(gclk));
	jdff dff_A_1tqHPfDU0_0(.dout(w_dff_A_QNhc1giV7_0),.din(w_dff_A_1tqHPfDU0_0),.clk(gclk));
	jdff dff_B_WGEwa6yO8_1(.din(n1060),.dout(w_dff_B_WGEwa6yO8_1),.clk(gclk));
	jdff dff_B_DKx92Ewv1_0(.din(n1112),.dout(w_dff_B_DKx92Ewv1_0),.clk(gclk));
	jdff dff_B_8Xg2FRhN2_0(.din(w_dff_B_DKx92Ewv1_0),.dout(w_dff_B_8Xg2FRhN2_0),.clk(gclk));
	jdff dff_B_dPVwk9Ay5_0(.din(w_dff_B_8Xg2FRhN2_0),.dout(w_dff_B_dPVwk9Ay5_0),.clk(gclk));
	jdff dff_B_Jdb6f3iR3_0(.din(n1111),.dout(w_dff_B_Jdb6f3iR3_0),.clk(gclk));
	jdff dff_B_3UuxGaOS6_0(.din(w_dff_B_Jdb6f3iR3_0),.dout(w_dff_B_3UuxGaOS6_0),.clk(gclk));
	jdff dff_B_I4JpWT8j1_0(.din(w_dff_B_3UuxGaOS6_0),.dout(w_dff_B_I4JpWT8j1_0),.clk(gclk));
	jdff dff_B_DGak4m8X4_0(.din(w_dff_B_I4JpWT8j1_0),.dout(w_dff_B_DGak4m8X4_0),.clk(gclk));
	jdff dff_B_LxJvPTEC3_0(.din(n1110),.dout(w_dff_B_LxJvPTEC3_0),.clk(gclk));
	jdff dff_B_bYYFb0U43_0(.din(w_dff_B_LxJvPTEC3_0),.dout(w_dff_B_bYYFb0U43_0),.clk(gclk));
	jdff dff_B_tApKYSbX2_0(.din(w_dff_B_bYYFb0U43_0),.dout(w_dff_B_tApKYSbX2_0),.clk(gclk));
	jdff dff_B_oV0HxQMx7_0(.din(n1109),.dout(w_dff_B_oV0HxQMx7_0),.clk(gclk));
	jdff dff_B_nFMmOQw68_0(.din(w_dff_B_oV0HxQMx7_0),.dout(w_dff_B_nFMmOQw68_0),.clk(gclk));
	jdff dff_B_PVquzBYK4_1(.din(n1066),.dout(w_dff_B_PVquzBYK4_1),.clk(gclk));
	jdff dff_B_AVSF0Oxw8_1(.din(w_dff_B_PVquzBYK4_1),.dout(w_dff_B_AVSF0Oxw8_1),.clk(gclk));
	jdff dff_B_PTsd3AOl7_1(.din(w_dff_B_AVSF0Oxw8_1),.dout(w_dff_B_PTsd3AOl7_1),.clk(gclk));
	jdff dff_B_xdVHyrCp1_1(.din(w_dff_B_PTsd3AOl7_1),.dout(w_dff_B_xdVHyrCp1_1),.clk(gclk));
	jdff dff_B_ijlws6n16_1(.din(w_dff_B_xdVHyrCp1_1),.dout(w_dff_B_ijlws6n16_1),.clk(gclk));
	jdff dff_B_B3dkUnZH3_1(.din(w_dff_B_ijlws6n16_1),.dout(w_dff_B_B3dkUnZH3_1),.clk(gclk));
	jdff dff_B_o4aZeyj90_0(.din(n1106),.dout(w_dff_B_o4aZeyj90_0),.clk(gclk));
	jdff dff_B_QZFZsH7S2_0(.din(n1105),.dout(w_dff_B_QZFZsH7S2_0),.clk(gclk));
	jdff dff_B_2wW6iHNC3_0(.din(w_dff_B_QZFZsH7S2_0),.dout(w_dff_B_2wW6iHNC3_0),.clk(gclk));
	jdff dff_B_2bFDFdJQ3_0(.din(w_dff_B_2wW6iHNC3_0),.dout(w_dff_B_2bFDFdJQ3_0),.clk(gclk));
	jdff dff_B_iLJQh0yV3_0(.din(w_dff_B_2bFDFdJQ3_0),.dout(w_dff_B_iLJQh0yV3_0),.clk(gclk));
	jdff dff_B_pbZN7arC8_0(.din(w_dff_B_iLJQh0yV3_0),.dout(w_dff_B_pbZN7arC8_0),.clk(gclk));
	jdff dff_B_ppXrUYdm2_0(.din(w_dff_B_pbZN7arC8_0),.dout(w_dff_B_ppXrUYdm2_0),.clk(gclk));
	jdff dff_B_4zeUQeoC6_1(.din(n1092),.dout(w_dff_B_4zeUQeoC6_1),.clk(gclk));
	jdff dff_B_qZohO1Mp1_0(.din(n1099),.dout(w_dff_B_qZohO1Mp1_0),.clk(gclk));
	jdff dff_B_OqWtzlI70_0(.din(n1097),.dout(w_dff_B_OqWtzlI70_0),.clk(gclk));
	jdff dff_B_26Vy7vBT7_0(.din(n1095),.dout(w_dff_B_26Vy7vBT7_0),.clk(gclk));
	jdff dff_B_2bfFMkNo0_0(.din(w_dff_B_26Vy7vBT7_0),.dout(w_dff_B_2bfFMkNo0_0),.clk(gclk));
	jdff dff_B_7MFYz6Q68_0(.din(w_dff_B_2bfFMkNo0_0),.dout(w_dff_B_7MFYz6Q68_0),.clk(gclk));
	jdff dff_B_RXABdTP05_1(.din(n1087),.dout(w_dff_B_RXABdTP05_1),.clk(gclk));
	jdff dff_B_mjJCM2hf6_0(.din(n1089),.dout(w_dff_B_mjJCM2hf6_0),.clk(gclk));
	jdff dff_B_Yh40dTcU2_1(.din(n1072),.dout(w_dff_B_Yh40dTcU2_1),.clk(gclk));
	jdff dff_B_yb49y52C9_1(.din(w_dff_B_Yh40dTcU2_1),.dout(w_dff_B_yb49y52C9_1),.clk(gclk));
	jdff dff_B_jYnSfBdI6_1(.din(w_dff_B_yb49y52C9_1),.dout(w_dff_B_jYnSfBdI6_1),.clk(gclk));
	jdff dff_B_DJYD2Cpt1_0(.din(n1084),.dout(w_dff_B_DJYD2Cpt1_0),.clk(gclk));
	jdff dff_B_lo148zU95_1(.din(n1080),.dout(w_dff_B_lo148zU95_1),.clk(gclk));
	jdff dff_B_jbbSM2MA9_1(.din(G124),.dout(w_dff_B_jbbSM2MA9_1),.clk(gclk));
	jdff dff_B_rSzU9W9K9_1(.din(w_dff_B_jbbSM2MA9_1),.dout(w_dff_B_rSzU9W9K9_1),.clk(gclk));
	jdff dff_B_4JQUvYtX3_1(.din(w_dff_B_rSzU9W9K9_1),.dout(w_dff_B_4JQUvYtX3_1),.clk(gclk));
	jdff dff_B_V4onKTSI5_1(.din(n1077),.dout(w_dff_B_V4onKTSI5_1),.clk(gclk));
	jdff dff_B_2BA9YJBT0_0(.din(n1075),.dout(w_dff_B_2BA9YJBT0_0),.clk(gclk));
	jdff dff_B_WLizeP4z7_0(.din(w_dff_B_2BA9YJBT0_0),.dout(w_dff_B_WLizeP4z7_0),.clk(gclk));
	jdff dff_B_hQWB1MV24_0(.din(w_dff_B_WLizeP4z7_0),.dout(w_dff_B_hQWB1MV24_0),.clk(gclk));
	jdff dff_B_B7rMKbCp5_0(.din(w_dff_B_hQWB1MV24_0),.dout(w_dff_B_B7rMKbCp5_0),.clk(gclk));
	jdff dff_B_F73aXzK84_1(.din(n1061),.dout(w_dff_B_F73aXzK84_1),.clk(gclk));
	jdff dff_B_dmMFLBrb2_1(.din(w_dff_B_F73aXzK84_1),.dout(w_dff_B_dmMFLBrb2_1),.clk(gclk));
	jdff dff_B_IhGxUNJH0_1(.din(n1051),.dout(w_dff_B_IhGxUNJH0_1),.clk(gclk));
	jdff dff_A_CzaUIjUg2_1(.dout(w_n1057_0[1]),.din(w_dff_A_CzaUIjUg2_1),.clk(gclk));
	jdff dff_A_RBGIcHEi1_1(.dout(w_dff_A_CzaUIjUg2_1),.din(w_dff_A_RBGIcHEi1_1),.clk(gclk));
	jdff dff_B_u0fVKxXR3_0(.din(n1055),.dout(w_dff_B_u0fVKxXR3_0),.clk(gclk));
	jdff dff_B_gT5iOp9K8_1(.din(n753),.dout(w_dff_B_gT5iOp9K8_1),.clk(gclk));
	jdff dff_B_3LIk1Ekd7_1(.din(w_dff_B_gT5iOp9K8_1),.dout(w_dff_B_3LIk1Ekd7_1),.clk(gclk));
	jdff dff_B_dtN22ksm2_1(.din(w_dff_B_3LIk1Ekd7_1),.dout(w_dff_B_dtN22ksm2_1),.clk(gclk));
	jdff dff_B_1kq4zCQq3_1(.din(w_dff_B_dtN22ksm2_1),.dout(w_dff_B_1kq4zCQq3_1),.clk(gclk));
	jdff dff_B_b5Osdyfb3_1(.din(w_dff_B_1kq4zCQq3_1),.dout(w_dff_B_b5Osdyfb3_1),.clk(gclk));
	jdff dff_B_dSbXADPr8_1(.din(w_dff_B_b5Osdyfb3_1),.dout(w_dff_B_dSbXADPr8_1),.clk(gclk));
	jdff dff_A_IdP4ctH51_1(.dout(w_n758_1[1]),.din(w_dff_A_IdP4ctH51_1),.clk(gclk));
	jdff dff_A_sYh46rC06_1(.dout(w_dff_A_IdP4ctH51_1),.din(w_dff_A_sYh46rC06_1),.clk(gclk));
	jdff dff_A_2huqbXvQ3_1(.dout(w_dff_A_sYh46rC06_1),.din(w_dff_A_2huqbXvQ3_1),.clk(gclk));
	jdff dff_B_c3brB32t2_0(.din(n752),.dout(w_dff_B_c3brB32t2_0),.clk(gclk));
	jdff dff_B_HRJ2qjEE6_0(.din(w_dff_B_c3brB32t2_0),.dout(w_dff_B_HRJ2qjEE6_0),.clk(gclk));
	jdff dff_B_1MxHLlVx4_0(.din(w_dff_B_HRJ2qjEE6_0),.dout(w_dff_B_1MxHLlVx4_0),.clk(gclk));
	jdff dff_B_Roa0scio0_0(.din(w_dff_B_1MxHLlVx4_0),.dout(w_dff_B_Roa0scio0_0),.clk(gclk));
	jdff dff_A_oSt1N62k5_0(.dout(w_n1049_0[0]),.din(w_dff_A_oSt1N62k5_0),.clk(gclk));
	jdff dff_A_4T6D0jPq0_1(.dout(w_n1049_0[1]),.din(w_dff_A_4T6D0jPq0_1),.clk(gclk));
	jdff dff_B_IrkBxSno6_0(.din(n1045),.dout(w_dff_B_IrkBxSno6_0),.clk(gclk));
	jdff dff_B_b0bU9vGe5_0(.din(w_dff_B_IrkBxSno6_0),.dout(w_dff_B_b0bU9vGe5_0),.clk(gclk));
	jdff dff_B_EeVSRKdi1_0(.din(w_dff_B_b0bU9vGe5_0),.dout(w_dff_B_EeVSRKdi1_0),.clk(gclk));
	jdff dff_B_Oxd3EAzS3_0(.din(w_dff_B_EeVSRKdi1_0),.dout(w_dff_B_Oxd3EAzS3_0),.clk(gclk));
	jdff dff_B_legx5ooM3_0(.din(w_dff_B_Oxd3EAzS3_0),.dout(w_dff_B_legx5ooM3_0),.clk(gclk));
	jdff dff_B_l47fYpKe0_1(.din(n1041),.dout(w_dff_B_l47fYpKe0_1),.clk(gclk));
	jdff dff_B_u0QRMWvq1_1(.din(w_dff_B_l47fYpKe0_1),.dout(w_dff_B_u0QRMWvq1_1),.clk(gclk));
	jdff dff_B_Fhq7c8ss2_0(.din(n1042),.dout(w_dff_B_Fhq7c8ss2_0),.clk(gclk));
	jdff dff_B_RTO9is4E1_0(.din(w_dff_B_Fhq7c8ss2_0),.dout(w_dff_B_RTO9is4E1_0),.clk(gclk));
	jdff dff_B_Bj8BiRrI3_1(.din(n1032),.dout(w_dff_B_Bj8BiRrI3_1),.clk(gclk));
	jdff dff_B_4HVNIoJw8_1(.din(n1035),.dout(w_dff_B_4HVNIoJw8_1),.clk(gclk));
	jdff dff_B_bGx2WRnA7_1(.din(n1027),.dout(w_dff_B_bGx2WRnA7_1),.clk(gclk));
	jdff dff_B_rJw8V6fi8_0(.din(n1028),.dout(w_dff_B_rJw8V6fi8_0),.clk(gclk));
	jdff dff_B_kikptGj60_1(.din(n1020),.dout(w_dff_B_kikptGj60_1),.clk(gclk));
	jdff dff_B_T6FbOtID0_1(.din(n1021),.dout(w_dff_B_T6FbOtID0_1),.clk(gclk));
	jdff dff_B_LdT9P7kQ6_1(.din(n1011),.dout(w_dff_B_LdT9P7kQ6_1),.clk(gclk));
	jdff dff_B_wvhPnYKL8_0(.din(n1013),.dout(w_dff_B_wvhPnYKL8_0),.clk(gclk));
	jdff dff_B_NmoD7dCD2_2(.din(G125),.dout(w_dff_B_NmoD7dCD2_2),.clk(gclk));
	jdff dff_B_e0kCTptf6_2(.din(w_dff_B_NmoD7dCD2_2),.dout(w_dff_B_e0kCTptf6_2),.clk(gclk));
	jdff dff_B_3NFxnZsM7_2(.din(w_dff_B_e0kCTptf6_2),.dout(w_dff_B_3NFxnZsM7_2),.clk(gclk));
	jdff dff_A_nMX3tB6p1_1(.dout(w_n990_0[1]),.din(w_dff_A_nMX3tB6p1_1),.clk(gclk));
	jdff dff_A_jYgrIUsq7_1(.dout(w_dff_A_nMX3tB6p1_1),.din(w_dff_A_jYgrIUsq7_1),.clk(gclk));
	jdff dff_A_fcW30N6G1_1(.dout(w_n758_0[1]),.din(w_dff_A_fcW30N6G1_1),.clk(gclk));
	jdff dff_A_7sA1ggSy2_1(.dout(w_dff_A_fcW30N6G1_1),.din(w_dff_A_7sA1ggSy2_1),.clk(gclk));
	jdff dff_A_LqppROXH2_1(.dout(w_dff_A_7sA1ggSy2_1),.din(w_dff_A_LqppROXH2_1),.clk(gclk));
	jdff dff_B_crVwk4RA1_0(.din(n757),.dout(w_dff_B_crVwk4RA1_0),.clk(gclk));
	jdff dff_A_kcaawKiK3_0(.dout(w_n769_0[0]),.din(w_dff_A_kcaawKiK3_0),.clk(gclk));
	jdff dff_B_TCA5IC1A5_0(.din(n768),.dout(w_dff_B_TCA5IC1A5_0),.clk(gclk));
	jdff dff_B_RWqRYJSi4_0(.din(w_dff_B_TCA5IC1A5_0),.dout(w_dff_B_RWqRYJSi4_0),.clk(gclk));
	jdff dff_B_eQDmSvRQ5_0(.din(w_dff_B_RWqRYJSi4_0),.dout(w_dff_B_eQDmSvRQ5_0),.clk(gclk));
	jdff dff_B_SyaITMJG9_0(.din(n767),.dout(w_dff_B_SyaITMJG9_0),.clk(gclk));
	jdff dff_B_LI2DMJ7g8_0(.din(w_dff_B_SyaITMJG9_0),.dout(w_dff_B_LI2DMJ7g8_0),.clk(gclk));
	jdff dff_A_SbYlVY0u7_2(.dout(w_n764_1[2]),.din(w_dff_A_SbYlVY0u7_2),.clk(gclk));
	jdff dff_A_M88EWdos2_2(.dout(w_dff_A_SbYlVY0u7_2),.din(w_dff_A_M88EWdos2_2),.clk(gclk));
	jdff dff_A_pdmCXQak7_2(.dout(w_dff_A_M88EWdos2_2),.din(w_dff_A_pdmCXQak7_2),.clk(gclk));
	jdff dff_B_8JH86pGa9_0(.din(n1182),.dout(w_dff_B_8JH86pGa9_0),.clk(gclk));
	jdff dff_B_RDYtqR090_0(.din(w_dff_B_8JH86pGa9_0),.dout(w_dff_B_RDYtqR090_0),.clk(gclk));
	jdff dff_B_MtfLmKbi8_1(.din(n1180),.dout(w_dff_B_MtfLmKbi8_1),.clk(gclk));
	jdff dff_B_I5WQYAhc1_1(.din(w_dff_B_MtfLmKbi8_1),.dout(w_dff_B_I5WQYAhc1_1),.clk(gclk));
	jdff dff_B_6LfJIXbT7_0(.din(n987),.dout(w_dff_B_6LfJIXbT7_0),.clk(gclk));
	jdff dff_B_J4fxFNtS0_1(.din(n944),.dout(w_dff_B_J4fxFNtS0_1),.clk(gclk));
	jdff dff_B_JWLVUhxx3_0(.din(n984),.dout(w_dff_B_JWLVUhxx3_0),.clk(gclk));
	jdff dff_B_0EyZIcUc8_0(.din(w_dff_B_JWLVUhxx3_0),.dout(w_dff_B_0EyZIcUc8_0),.clk(gclk));
	jdff dff_B_K3IeCsJk6_0(.din(w_dff_B_0EyZIcUc8_0),.dout(w_dff_B_K3IeCsJk6_0),.clk(gclk));
	jdff dff_B_xeCC2MJU7_0(.din(w_dff_B_K3IeCsJk6_0),.dout(w_dff_B_xeCC2MJU7_0),.clk(gclk));
	jdff dff_B_et0EBgT21_1(.din(n978),.dout(w_dff_B_et0EBgT21_1),.clk(gclk));
	jdff dff_B_EeBQm7hU3_1(.din(n979),.dout(w_dff_B_EeBQm7hU3_1),.clk(gclk));
	jdff dff_B_CsuIWoK75_0(.din(n980),.dout(w_dff_B_CsuIWoK75_0),.clk(gclk));
	jdff dff_A_7AcN7zvh3_2(.dout(w_G97_2[2]),.din(w_dff_A_7AcN7zvh3_2),.clk(gclk));
	jdff dff_B_DU2XGEIQ6_2(.din(n144),.dout(w_dff_B_DU2XGEIQ6_2),.clk(gclk));
	jdff dff_B_tZTxkOmW8_1(.din(n142),.dout(w_dff_B_tZTxkOmW8_1),.clk(gclk));
	jdff dff_B_QTK8jM607_1(.din(n968),.dout(w_dff_B_QTK8jM607_1),.clk(gclk));
	jdff dff_B_bBjhKhHV1_1(.din(n971),.dout(w_dff_B_bBjhKhHV1_1),.clk(gclk));
	jdff dff_B_t7y68eUg3_0(.din(n972),.dout(w_dff_B_t7y68eUg3_0),.clk(gclk));
	jdff dff_A_5a2f4HA13_0(.dout(w_G143_1[0]),.din(w_dff_A_5a2f4HA13_0),.clk(gclk));
	jdff dff_A_xcnpLyZY2_1(.dout(w_G33_4[1]),.din(w_dff_A_xcnpLyZY2_1),.clk(gclk));
	jdff dff_A_LTTgHIkk4_1(.dout(w_dff_A_xcnpLyZY2_1),.din(w_dff_A_LTTgHIkk4_1),.clk(gclk));
	jdff dff_A_h0TQx0tk1_1(.dout(w_dff_A_LTTgHIkk4_1),.din(w_dff_A_h0TQx0tk1_1),.clk(gclk));
	jdff dff_A_PdBQPsih0_1(.dout(w_dff_A_h0TQx0tk1_1),.din(w_dff_A_PdBQPsih0_1),.clk(gclk));
	jdff dff_A_PA0pLMAL5_2(.dout(w_G33_4[2]),.din(w_dff_A_PA0pLMAL5_2),.clk(gclk));
	jdff dff_A_TuMdgiC28_2(.dout(w_dff_A_PA0pLMAL5_2),.din(w_dff_A_TuMdgiC28_2),.clk(gclk));
	jdff dff_A_swxpps9B3_2(.dout(w_dff_A_TuMdgiC28_2),.din(w_dff_A_swxpps9B3_2),.clk(gclk));
	jdff dff_B_yW3zibOM5_0(.din(n964),.dout(w_dff_B_yW3zibOM5_0),.clk(gclk));
	jdff dff_B_NKahejBj1_1(.din(n953),.dout(w_dff_B_NKahejBj1_1),.clk(gclk));
	jdff dff_B_u811M5jM0_1(.din(n956),.dout(w_dff_B_u811M5jM0_1),.clk(gclk));
	jdff dff_B_V6mBJiHs9_0(.din(n957),.dout(w_dff_B_V6mBJiHs9_0),.clk(gclk));
	jdff dff_B_OGdqf51U6_0(.din(n949),.dout(w_dff_B_OGdqf51U6_0),.clk(gclk));
	jdff dff_A_BNcqOQnr9_0(.dout(w_n603_1[0]),.din(w_dff_A_BNcqOQnr9_0),.clk(gclk));
	jdff dff_A_37fG59s46_0(.dout(w_dff_A_BNcqOQnr9_0),.din(w_dff_A_37fG59s46_0),.clk(gclk));
	jdff dff_A_Cu0d6UVD6_0(.dout(w_dff_A_37fG59s46_0),.din(w_dff_A_Cu0d6UVD6_0),.clk(gclk));
	jdff dff_A_LJEiiwrx0_0(.dout(w_dff_A_Cu0d6UVD6_0),.din(w_dff_A_LJEiiwrx0_0),.clk(gclk));
	jdff dff_A_Rmpq5NyL1_1(.dout(w_n603_1[1]),.din(w_dff_A_Rmpq5NyL1_1),.clk(gclk));
	jdff dff_A_ma6Qyv6a7_1(.dout(w_dff_A_Rmpq5NyL1_1),.din(w_dff_A_ma6Qyv6a7_1),.clk(gclk));
	jdff dff_A_99HJibvw4_1(.dout(w_dff_A_ma6Qyv6a7_1),.din(w_dff_A_99HJibvw4_1),.clk(gclk));
	jdff dff_B_MtzuOHMI5_0(.din(n942),.dout(w_dff_B_MtzuOHMI5_0),.clk(gclk));
	jdff dff_A_HeEO2Nmd3_1(.dout(w_n940_0[1]),.din(w_dff_A_HeEO2Nmd3_1),.clk(gclk));
	jdff dff_A_y3dUgMXB2_1(.dout(w_dff_A_HeEO2Nmd3_1),.din(w_dff_A_y3dUgMXB2_1),.clk(gclk));
	jdff dff_B_rv7l7Nhd4_1(.din(n850),.dout(w_dff_B_rv7l7Nhd4_1),.clk(gclk));
	jdff dff_B_VmrBYFvk2_1(.din(w_dff_B_rv7l7Nhd4_1),.dout(w_dff_B_VmrBYFvk2_1),.clk(gclk));
	jdff dff_B_DJ7CFo3m2_0(.din(n875),.dout(w_dff_B_DJ7CFo3m2_0),.clk(gclk));
	jdff dff_B_xo4Jgk4M3_0(.din(w_dff_B_DJ7CFo3m2_0),.dout(w_dff_B_xo4Jgk4M3_0),.clk(gclk));
	jdff dff_B_BUE8W33A7_0(.din(n872),.dout(w_dff_B_BUE8W33A7_0),.clk(gclk));
	jdff dff_B_OPcy1Z589_1(.din(n868),.dout(w_dff_B_OPcy1Z589_1),.clk(gclk));
	jdff dff_B_FGtXuGGF7_1(.din(w_dff_B_OPcy1Z589_1),.dout(w_dff_B_FGtXuGGF7_1),.clk(gclk));
	jdff dff_B_1J4G0RQ80_1(.din(w_dff_B_FGtXuGGF7_1),.dout(w_dff_B_1J4G0RQ80_1),.clk(gclk));
	jdff dff_B_0L24BZH86_1(.din(w_dff_B_1J4G0RQ80_1),.dout(w_dff_B_0L24BZH86_1),.clk(gclk));
	jdff dff_A_WDPW7eG30_1(.dout(w_n863_0[1]),.din(w_dff_A_WDPW7eG30_1),.clk(gclk));
	jdff dff_A_70LQrWZs1_1(.dout(w_dff_A_WDPW7eG30_1),.din(w_dff_A_70LQrWZs1_1),.clk(gclk));
	jdff dff_B_q6WBqKV42_0(.din(n857),.dout(w_dff_B_q6WBqKV42_0),.clk(gclk));
	jdff dff_B_khDDenXF7_0(.din(w_dff_B_q6WBqKV42_0),.dout(w_dff_B_khDDenXF7_0),.clk(gclk));
	jdff dff_B_K9CLbvgv0_0(.din(w_dff_B_khDDenXF7_0),.dout(w_dff_B_K9CLbvgv0_0),.clk(gclk));
	jdff dff_B_XoM5BIMh5_3(.din(n563),.dout(w_dff_B_XoM5BIMh5_3),.clk(gclk));
	jdff dff_B_hFsXgRLs2_1(.din(n555),.dout(w_dff_B_hFsXgRLs2_1),.clk(gclk));
	jdff dff_B_ZwcaPGGG5_1(.din(w_dff_B_hFsXgRLs2_1),.dout(w_dff_B_ZwcaPGGG5_1),.clk(gclk));
	jdff dff_B_JanaiJrn9_0(.din(n849),.dout(w_dff_B_JanaiJrn9_0),.clk(gclk));
	jdff dff_B_CipYhRss3_0(.din(w_dff_B_JanaiJrn9_0),.dout(w_dff_B_CipYhRss3_0),.clk(gclk));
	jdff dff_B_kbCxJTKh5_0(.din(n848),.dout(w_dff_B_kbCxJTKh5_0),.clk(gclk));
	jdff dff_B_oAeiECGu0_0(.din(w_dff_B_kbCxJTKh5_0),.dout(w_dff_B_oAeiECGu0_0),.clk(gclk));
	jdff dff_B_786NVzyQ2_0(.din(w_dff_B_oAeiECGu0_0),.dout(w_dff_B_786NVzyQ2_0),.clk(gclk));
	jdff dff_B_2Etd3YNq0_0(.din(w_dff_B_786NVzyQ2_0),.dout(w_dff_B_2Etd3YNq0_0),.clk(gclk));
	jdff dff_B_yS816wcL4_1(.din(n844),.dout(w_dff_B_yS816wcL4_1),.clk(gclk));
	jdff dff_B_VKqW2bGp3_0(.din(n845),.dout(w_dff_B_VKqW2bGp3_0),.clk(gclk));
	jdff dff_A_AZhXc43T4_0(.dout(w_n131_0[0]),.din(w_dff_A_AZhXc43T4_0),.clk(gclk));
	jdff dff_B_DhQRgtAm4_1(.din(n129),.dout(w_dff_B_DhQRgtAm4_1),.clk(gclk));
	jdff dff_B_ZUSVDj2j0_1(.din(n820),.dout(w_dff_B_ZUSVDj2j0_1),.clk(gclk));
	jdff dff_B_qPT0ujuH2_1(.din(w_dff_B_ZUSVDj2j0_1),.dout(w_dff_B_qPT0ujuH2_1),.clk(gclk));
	jdff dff_B_DwVnuUP80_1(.din(w_dff_B_qPT0ujuH2_1),.dout(w_dff_B_DwVnuUP80_1),.clk(gclk));
	jdff dff_B_WJZSQhCj2_1(.din(w_dff_B_DwVnuUP80_1),.dout(w_dff_B_WJZSQhCj2_1),.clk(gclk));
	jdff dff_B_k9MMBBPr6_1(.din(w_dff_B_WJZSQhCj2_1),.dout(w_dff_B_k9MMBBPr6_1),.clk(gclk));
	jdff dff_B_bs5p4BPX4_0(.din(n839),.dout(w_dff_B_bs5p4BPX4_0),.clk(gclk));
	jdff dff_B_hlJjD9Rg6_0(.din(w_dff_B_bs5p4BPX4_0),.dout(w_dff_B_hlJjD9Rg6_0),.clk(gclk));
	jdff dff_B_5S32BAId0_1(.din(n830),.dout(w_dff_B_5S32BAId0_1),.clk(gclk));
	jdff dff_B_V844WwYT9_1(.din(n833),.dout(w_dff_B_V844WwYT9_1),.clk(gclk));
	jdff dff_B_MvjyWkCQ5_1(.din(n834),.dout(w_dff_B_MvjyWkCQ5_1),.clk(gclk));
	jdff dff_B_BG6W7Crp7_1(.din(n822),.dout(w_dff_B_BG6W7Crp7_1),.clk(gclk));
	jdff dff_B_krmUV8RO2_1(.din(w_dff_B_BG6W7Crp7_1),.dout(w_dff_B_krmUV8RO2_1),.clk(gclk));
	jdff dff_B_KQKiFyKL2_1(.din(n814),.dout(w_dff_B_KQKiFyKL2_1),.clk(gclk));
	jdff dff_B_xVasj5kJ8_1(.din(n815),.dout(w_dff_B_xVasj5kJ8_1),.clk(gclk));
	jdff dff_B_jy15bCAb1_1(.din(n805),.dout(w_dff_B_jy15bCAb1_1),.clk(gclk));
	jdff dff_B_epMcabcQ1_0(.din(n807),.dout(w_dff_B_epMcabcQ1_0),.clk(gclk));
	jdff dff_A_G37cgPAn4_2(.dout(w_G107_2[2]),.din(w_dff_A_G37cgPAn4_2),.clk(gclk));
	jdff dff_B_wqUxesZM3_0(.din(n800),.dout(w_dff_B_wqUxesZM3_0),.clk(gclk));
	jdff dff_B_9d9RryJv7_0(.din(n936),.dout(w_dff_B_9d9RryJv7_0),.clk(gclk));
	jdff dff_B_YRi0c8Xj3_0(.din(w_dff_B_9d9RryJv7_0),.dout(w_dff_B_YRi0c8Xj3_0),.clk(gclk));
	jdff dff_B_oYg0olwJ0_1(.din(n915),.dout(w_dff_B_oYg0olwJ0_1),.clk(gclk));
	jdff dff_B_pxdSli3m3_1(.din(w_dff_B_oYg0olwJ0_1),.dout(w_dff_B_pxdSli3m3_1),.clk(gclk));
	jdff dff_B_iDRMvkcQ1_1(.din(w_dff_B_pxdSli3m3_1),.dout(w_dff_B_iDRMvkcQ1_1),.clk(gclk));
	jdff dff_B_1Cq0U0a39_1(.din(n924),.dout(w_dff_B_1Cq0U0a39_1),.clk(gclk));
	jdff dff_B_c5054Njd6_1(.din(w_dff_B_1Cq0U0a39_1),.dout(w_dff_B_c5054Njd6_1),.clk(gclk));
	jdff dff_B_8VZ402Ky1_1(.din(n925),.dout(w_dff_B_8VZ402Ky1_1),.clk(gclk));
	jdff dff_B_PrT57hO05_1(.din(n916),.dout(w_dff_B_PrT57hO05_1),.clk(gclk));
	jdff dff_B_vHxeNTmt0_1(.din(n918),.dout(w_dff_B_vHxeNTmt0_1),.clk(gclk));
	jdff dff_A_HdEUKy3C7_1(.dout(w_n73_1[1]),.din(w_dff_A_HdEUKy3C7_1),.clk(gclk));
	jdff dff_A_Yxo3N9Dl4_1(.dout(w_n135_0[1]),.din(w_dff_A_Yxo3N9Dl4_1),.clk(gclk));
	jdff dff_B_QmBhjrpP1_1(.din(n133),.dout(w_dff_B_QmBhjrpP1_1),.clk(gclk));
	jdff dff_B_5KLB4HMo4_1(.din(n904),.dout(w_dff_B_5KLB4HMo4_1),.clk(gclk));
	jdff dff_B_Ve7dusDi5_1(.din(n907),.dout(w_dff_B_Ve7dusDi5_1),.clk(gclk));
	jdff dff_B_8NAA6ogq4_1(.din(n908),.dout(w_dff_B_8NAA6ogq4_1),.clk(gclk));
	jdff dff_A_GMDgsM5t5_0(.dout(w_G50_2[0]),.din(w_dff_A_GMDgsM5t5_0),.clk(gclk));
	jdff dff_A_JhtiTWaw7_1(.dout(w_G68_2[1]),.din(w_dff_A_JhtiTWaw7_1),.clk(gclk));
	jdff dff_A_eKFFuyiO9_1(.dout(w_dff_A_JhtiTWaw7_1),.din(w_dff_A_eKFFuyiO9_1),.clk(gclk));
	jdff dff_A_skVO2sRG1_1(.dout(w_dff_A_eKFFuyiO9_1),.din(w_dff_A_skVO2sRG1_1),.clk(gclk));
	jdff dff_A_GAnDltAD0_2(.dout(w_G68_2[2]),.din(w_dff_A_GAnDltAD0_2),.clk(gclk));
	jdff dff_A_Cr9tn0ke9_2(.dout(w_dff_A_GAnDltAD0_2),.din(w_dff_A_Cr9tn0ke9_2),.clk(gclk));
	jdff dff_A_9GBNWQMK3_2(.dout(w_dff_A_Cr9tn0ke9_2),.din(w_dff_A_9GBNWQMK3_2),.clk(gclk));
	jdff dff_A_9nNLVVbJ4_2(.dout(w_dff_A_9GBNWQMK3_2),.din(w_dff_A_9nNLVVbJ4_2),.clk(gclk));
	jdff dff_B_QA35yFD00_0(.din(n900),.dout(w_dff_B_QA35yFD00_0),.clk(gclk));
	jdff dff_A_3acfUPkO1_0(.dout(w_G58_2[0]),.din(w_dff_A_3acfUPkO1_0),.clk(gclk));
	jdff dff_A_vVDfAQXi7_0(.dout(w_dff_A_3acfUPkO1_0),.din(w_dff_A_vVDfAQXi7_0),.clk(gclk));
	jdff dff_A_Jrn4DL1P6_2(.dout(w_G58_2[2]),.din(w_dff_A_Jrn4DL1P6_2),.clk(gclk));
	jdff dff_A_tLivtiAV8_2(.dout(w_dff_A_Jrn4DL1P6_2),.din(w_dff_A_tLivtiAV8_2),.clk(gclk));
	jdff dff_B_hU0nysu46_0(.din(n895),.dout(w_dff_B_hU0nysu46_0),.clk(gclk));
	jdff dff_B_rQOiTh2F7_0(.din(n891),.dout(w_dff_B_rQOiTh2F7_0),.clk(gclk));
	jdff dff_A_c9wDqvvY5_1(.dout(w_G116_2[1]),.din(w_dff_A_c9wDqvvY5_1),.clk(gclk));
	jdff dff_A_j3wkjTyJ9_2(.dout(w_G116_2[2]),.din(w_dff_A_j3wkjTyJ9_2),.clk(gclk));
	jdff dff_A_weg0WuY85_1(.dout(w_n148_4[1]),.din(w_dff_A_weg0WuY85_1),.clk(gclk));
	jdff dff_A_D9DjRBCi5_2(.dout(w_n148_4[2]),.din(w_dff_A_D9DjRBCi5_2),.clk(gclk));
	jdff dff_B_p66zbhX35_1(.din(n883),.dout(w_dff_B_p66zbhX35_1),.clk(gclk));
	jdff dff_B_ViLt7ylH0_0(.din(n885),.dout(w_dff_B_ViLt7ylH0_0),.clk(gclk));
	jdff dff_A_SzkP9lAQ1_0(.dout(w_G283_2[0]),.din(w_dff_A_SzkP9lAQ1_0),.clk(gclk));
	jdff dff_A_xZZrXenR4_1(.dout(w_G283_2[1]),.din(w_dff_A_xZZrXenR4_1),.clk(gclk));
	jdff dff_B_CU5aFT977_1(.din(n878),.dout(w_dff_B_CU5aFT977_1),.clk(gclk));
	jdff dff_B_Yvw3WQHh8_0(.din(n854),.dout(w_dff_B_Yvw3WQHh8_0),.clk(gclk));
	jdff dff_A_Tiy1oMGB9_0(.dout(w_n589_1[0]),.din(w_dff_A_Tiy1oMGB9_0),.clk(gclk));
	jdff dff_A_6g9wIwMo1_0(.dout(w_dff_A_Tiy1oMGB9_0),.din(w_dff_A_6g9wIwMo1_0),.clk(gclk));
	jdff dff_A_7F7lXBco6_0(.dout(w_dff_A_6g9wIwMo1_0),.din(w_dff_A_7F7lXBco6_0),.clk(gclk));
	jdff dff_A_JO8zr94B0_0(.dout(w_n592_1[0]),.din(w_dff_A_JO8zr94B0_0),.clk(gclk));
	jdff dff_A_kHIp0HDB7_0(.dout(w_dff_A_JO8zr94B0_0),.din(w_dff_A_kHIp0HDB7_0),.clk(gclk));
	jdff dff_A_UEPnqtJ47_0(.dout(w_dff_A_kHIp0HDB7_0),.din(w_dff_A_UEPnqtJ47_0),.clk(gclk));
	jdff dff_A_t2jFqypB4_1(.dout(w_n592_1[1]),.din(w_dff_A_t2jFqypB4_1),.clk(gclk));
	jdff dff_A_Ba2yrQhG0_1(.dout(w_n853_0[1]),.din(w_dff_A_Ba2yrQhG0_1),.clk(gclk));
	jdff dff_B_2PCwmbBR7_0(.din(n560),.dout(w_dff_B_2PCwmbBR7_0),.clk(gclk));
	jdff dff_B_Zx7LqFSw7_0(.din(w_dff_B_2PCwmbBR7_0),.dout(w_dff_B_Zx7LqFSw7_0),.clk(gclk));
	jdff dff_B_FaljJk7V4_0(.din(n558),.dout(w_dff_B_FaljJk7V4_0),.clk(gclk));
	jdff dff_B_vHDgTMOi9_2(.din(n556),.dout(w_dff_B_vHDgTMOi9_2),.clk(gclk));
	jdff dff_A_TdTjlMHl0_0(.dout(w_G396_0[0]),.din(w_dff_A_TdTjlMHl0_0),.clk(gclk));
	jdff dff_A_8WxTUa831_0(.dout(w_dff_A_TdTjlMHl0_0),.din(w_dff_A_8WxTUa831_0),.clk(gclk));
	jdff dff_B_THST2BMr9_0(.din(n686),.dout(w_dff_B_THST2BMr9_0),.clk(gclk));
	jdff dff_B_GTezD0Qw4_0(.din(w_dff_B_THST2BMr9_0),.dout(w_dff_B_GTezD0Qw4_0),.clk(gclk));
	jdff dff_B_YDTS5TL70_1(.din(n678),.dout(w_dff_B_YDTS5TL70_1),.clk(gclk));
	jdff dff_B_nb4eicKF1_1(.din(w_dff_B_YDTS5TL70_1),.dout(w_dff_B_nb4eicKF1_1),.clk(gclk));
	jdff dff_B_kDfzSqZk9_1(.din(n679),.dout(w_dff_B_kDfzSqZk9_1),.clk(gclk));
	jdff dff_B_Ivzg3xIC2_2(.din(n680),.dout(w_dff_B_Ivzg3xIC2_2),.clk(gclk));
	jdff dff_B_qFYVwUnH9_1(.din(n673),.dout(w_dff_B_qFYVwUnH9_1),.clk(gclk));
	jdff dff_B_46XW8r5J1_0(.din(n139),.dout(w_dff_B_46XW8r5J1_0),.clk(gclk));
	jdff dff_A_YLbAZ4IE3_1(.dout(w_n672_1[1]),.din(w_dff_A_YLbAZ4IE3_1),.clk(gclk));
	jdff dff_A_RtHqXjHw8_1(.dout(w_dff_A_YLbAZ4IE3_1),.din(w_dff_A_RtHqXjHw8_1),.clk(gclk));
	jdff dff_A_RTF9YcsN6_2(.dout(w_n672_0[2]),.din(w_dff_A_RTF9YcsN6_2),.clk(gclk));
	jdff dff_A_88dtetgu2_2(.dout(w_dff_A_RTF9YcsN6_2),.din(w_dff_A_88dtetgu2_2),.clk(gclk));
	jdff dff_B_fbIPnkxY0_1(.din(n647),.dout(w_dff_B_fbIPnkxY0_1),.clk(gclk));
	jdff dff_B_HZzZqG3p2_1(.din(w_dff_B_fbIPnkxY0_1),.dout(w_dff_B_HZzZqG3p2_1),.clk(gclk));
	jdff dff_B_mvi4auYb9_1(.din(w_dff_B_HZzZqG3p2_1),.dout(w_dff_B_mvi4auYb9_1),.clk(gclk));
	jdff dff_B_zwFczmjs6_1(.din(w_dff_B_mvi4auYb9_1),.dout(w_dff_B_zwFczmjs6_1),.clk(gclk));
	jdff dff_B_Xa2q3nUo6_1(.din(w_dff_B_zwFczmjs6_1),.dout(w_dff_B_Xa2q3nUo6_1),.clk(gclk));
	jdff dff_B_1qY5Qug65_1(.din(n653),.dout(w_dff_B_1qY5Qug65_1),.clk(gclk));
	jdff dff_B_czY4iSWw4_1(.din(w_dff_B_1qY5Qug65_1),.dout(w_dff_B_czY4iSWw4_1),.clk(gclk));
	jdff dff_B_ZfTKSLIY4_1(.din(w_dff_B_czY4iSWw4_1),.dout(w_dff_B_ZfTKSLIY4_1),.clk(gclk));
	jdff dff_B_JjmVLEll5_0(.din(n664),.dout(w_dff_B_JjmVLEll5_0),.clk(gclk));
	jdff dff_B_cY4O8HI96_1(.din(n660),.dout(w_dff_B_cY4O8HI96_1),.clk(gclk));
	jdff dff_B_FpeKF35t2_0(.din(n658),.dout(w_dff_B_FpeKF35t2_0),.clk(gclk));
	jdff dff_B_3wSKf3w46_1(.din(n633),.dout(w_dff_B_3wSKf3w46_1),.clk(gclk));
	jdff dff_B_dI0eegyn0_0(.din(n644),.dout(w_dff_B_dI0eegyn0_0),.clk(gclk));
	jdff dff_B_Ol7dW2sh1_3(.din(G317),.dout(w_dff_B_Ol7dW2sh1_3),.clk(gclk));
	jdff dff_B_W5QdNekh4_3(.din(w_dff_B_Ol7dW2sh1_3),.dout(w_dff_B_W5QdNekh4_3),.clk(gclk));
	jdff dff_B_fFWHIJFq9_3(.din(w_dff_B_W5QdNekh4_3),.dout(w_dff_B_fFWHIJFq9_3),.clk(gclk));
	jdff dff_B_xE9yzJRL6_2(.din(G326),.dout(w_dff_B_xE9yzJRL6_2),.clk(gclk));
	jdff dff_B_m5lLCWo20_2(.din(w_dff_B_xE9yzJRL6_2),.dout(w_dff_B_m5lLCWo20_2),.clk(gclk));
	jdff dff_B_sAp9YiIm4_2(.din(w_dff_B_m5lLCWo20_2),.dout(w_dff_B_sAp9YiIm4_2),.clk(gclk));
	jdff dff_B_89NlwPhh7_0(.din(n637),.dout(w_dff_B_89NlwPhh7_0),.clk(gclk));
	jdff dff_B_l8LxeCNm6_1(.din(G329),.dout(w_dff_B_l8LxeCNm6_1),.clk(gclk));
	jdff dff_B_gKYk9sFL5_1(.din(w_dff_B_l8LxeCNm6_1),.dout(w_dff_B_gKYk9sFL5_1),.clk(gclk));
	jdff dff_B_kjHWZixp2_1(.din(w_dff_B_gKYk9sFL5_1),.dout(w_dff_B_kjHWZixp2_1),.clk(gclk));
	jdff dff_A_xtKFON032_1(.dout(w_n148_5[1]),.din(w_dff_A_xtKFON032_1),.clk(gclk));
	jdff dff_A_5KU2o8vn6_1(.dout(w_dff_A_xtKFON032_1),.din(w_dff_A_5KU2o8vn6_1),.clk(gclk));
	jdff dff_A_EI2Ilcku7_1(.dout(w_dff_A_5KU2o8vn6_1),.din(w_dff_A_EI2Ilcku7_1),.clk(gclk));
	jdff dff_A_MVA5MfC56_2(.dout(w_n148_5[2]),.din(w_dff_A_MVA5MfC56_2),.clk(gclk));
	jdff dff_B_Nf5ZYQsw4_0(.din(n628),.dout(w_dff_B_Nf5ZYQsw4_0),.clk(gclk));
	jdff dff_B_I8HULOXn1_3(.din(G322),.dout(w_dff_B_I8HULOXn1_3),.clk(gclk));
	jdff dff_B_fUDQcBrn4_3(.din(w_dff_B_I8HULOXn1_3),.dout(w_dff_B_fUDQcBrn4_3),.clk(gclk));
	jdff dff_B_ug54TCuZ7_3(.din(w_dff_B_fUDQcBrn4_3),.dout(w_dff_B_ug54TCuZ7_3),.clk(gclk));
	jdff dff_A_oNML8KrU4_1(.dout(w_n612_4[1]),.din(w_dff_A_oNML8KrU4_1),.clk(gclk));
	jdff dff_A_fkGtClK13_1(.dout(w_dff_A_oNML8KrU4_1),.din(w_dff_A_fkGtClK13_1),.clk(gclk));
	jdff dff_A_7zgZhvPP8_1(.dout(w_dff_A_fkGtClK13_1),.din(w_dff_A_7zgZhvPP8_1),.clk(gclk));
	jdff dff_A_bZ7ijSYX5_1(.dout(w_dff_A_7zgZhvPP8_1),.din(w_dff_A_bZ7ijSYX5_1),.clk(gclk));
	jdff dff_A_NOiZkSxo8_1(.dout(w_dff_A_bZ7ijSYX5_1),.din(w_dff_A_NOiZkSxo8_1),.clk(gclk));
	jdff dff_A_IjIfmfFq0_1(.dout(w_dff_A_NOiZkSxo8_1),.din(w_dff_A_IjIfmfFq0_1),.clk(gclk));
	jdff dff_A_vnEzpc403_1(.dout(w_dff_A_IjIfmfFq0_1),.din(w_dff_A_vnEzpc403_1),.clk(gclk));
	jdff dff_A_IXYedGQu8_0(.dout(w_n608_1[0]),.din(w_dff_A_IXYedGQu8_0),.clk(gclk));
	jdff dff_A_XXccezFo3_0(.dout(w_dff_A_IXYedGQu8_0),.din(w_dff_A_XXccezFo3_0),.clk(gclk));
	jdff dff_A_mOWTb5FC6_0(.dout(w_dff_A_XXccezFo3_0),.din(w_dff_A_mOWTb5FC6_0),.clk(gclk));
	jdff dff_A_TZMEC8n68_0(.dout(w_dff_A_mOWTb5FC6_0),.din(w_dff_A_TZMEC8n68_0),.clk(gclk));
	jdff dff_A_SBZocElh5_0(.dout(w_dff_A_TZMEC8n68_0),.din(w_dff_A_SBZocElh5_0),.clk(gclk));
	jdff dff_A_4EQ5NfpF9_0(.dout(w_dff_A_SBZocElh5_0),.din(w_dff_A_4EQ5NfpF9_0),.clk(gclk));
	jdff dff_A_A6BCbUAz9_0(.dout(w_dff_A_4EQ5NfpF9_0),.din(w_dff_A_A6BCbUAz9_0),.clk(gclk));
	jdff dff_A_XVppy1kU6_0(.dout(w_dff_A_A6BCbUAz9_0),.din(w_dff_A_XVppy1kU6_0),.clk(gclk));
	jdff dff_A_Sdz9dIll5_0(.dout(w_dff_A_XVppy1kU6_0),.din(w_dff_A_Sdz9dIll5_0),.clk(gclk));
	jdff dff_A_kpzSiGhz9_2(.dout(w_n608_1[2]),.din(w_dff_A_kpzSiGhz9_2),.clk(gclk));
	jdff dff_A_L6gHmMgr3_2(.dout(w_dff_A_kpzSiGhz9_2),.din(w_dff_A_L6gHmMgr3_2),.clk(gclk));
	jdff dff_A_jYOdfjyW0_2(.dout(w_dff_A_L6gHmMgr3_2),.din(w_dff_A_jYOdfjyW0_2),.clk(gclk));
	jdff dff_A_A3JHM3JR6_2(.dout(w_dff_A_jYOdfjyW0_2),.din(w_dff_A_A3JHM3JR6_2),.clk(gclk));
	jdff dff_A_375oD3Ou8_2(.dout(w_dff_A_A3JHM3JR6_2),.din(w_dff_A_375oD3Ou8_2),.clk(gclk));
	jdff dff_A_rvfB9a4U4_2(.dout(w_dff_A_375oD3Ou8_2),.din(w_dff_A_rvfB9a4U4_2),.clk(gclk));
	jdff dff_A_ohTChJrT1_2(.dout(w_dff_A_rvfB9a4U4_2),.din(w_dff_A_ohTChJrT1_2),.clk(gclk));
	jdff dff_A_TgRKKufT2_1(.dout(w_n608_0[1]),.din(w_dff_A_TgRKKufT2_1),.clk(gclk));
	jdff dff_A_WaUW4dsG2_1(.dout(w_dff_A_TgRKKufT2_1),.din(w_dff_A_WaUW4dsG2_1),.clk(gclk));
	jdff dff_A_2ZcylJBQ1_1(.dout(w_dff_A_WaUW4dsG2_1),.din(w_dff_A_2ZcylJBQ1_1),.clk(gclk));
	jdff dff_A_WXyYF0iP0_1(.dout(w_dff_A_2ZcylJBQ1_1),.din(w_dff_A_WXyYF0iP0_1),.clk(gclk));
	jdff dff_A_TeFbGmaE3_1(.dout(w_dff_A_WXyYF0iP0_1),.din(w_dff_A_TeFbGmaE3_1),.clk(gclk));
	jdff dff_A_jWwQZyvX9_1(.dout(w_dff_A_TeFbGmaE3_1),.din(w_dff_A_jWwQZyvX9_1),.clk(gclk));
	jdff dff_A_dICPL2Kz8_1(.dout(w_dff_A_jWwQZyvX9_1),.din(w_dff_A_dICPL2Kz8_1),.clk(gclk));
	jdff dff_A_kZcMbeTU7_2(.dout(w_n608_0[2]),.din(w_dff_A_kZcMbeTU7_2),.clk(gclk));
	jdff dff_A_weYYilAH6_2(.dout(w_dff_A_kZcMbeTU7_2),.din(w_dff_A_weYYilAH6_2),.clk(gclk));
	jdff dff_A_6M9fzjsc1_2(.dout(w_dff_A_weYYilAH6_2),.din(w_dff_A_6M9fzjsc1_2),.clk(gclk));
	jdff dff_A_5iYGyZjj1_2(.dout(w_dff_A_6M9fzjsc1_2),.din(w_dff_A_5iYGyZjj1_2),.clk(gclk));
	jdff dff_A_2S75jRV98_2(.dout(w_dff_A_5iYGyZjj1_2),.din(w_dff_A_2S75jRV98_2),.clk(gclk));
	jdff dff_A_0PsnEPoP3_2(.dout(w_dff_A_2S75jRV98_2),.din(w_dff_A_0PsnEPoP3_2),.clk(gclk));
	jdff dff_A_9x6Qr2Io4_2(.dout(w_dff_A_0PsnEPoP3_2),.din(w_dff_A_9x6Qr2Io4_2),.clk(gclk));
	jdff dff_B_VudIogzL6_0(.din(n606),.dout(w_dff_B_VudIogzL6_0),.clk(gclk));
	jdff dff_B_aQjpBnWG0_0(.din(n570),.dout(w_dff_B_aQjpBnWG0_0),.clk(gclk));
	jdff dff_B_elJ768Fw9_0(.din(w_dff_B_aQjpBnWG0_0),.dout(w_dff_B_elJ768Fw9_0),.clk(gclk));
	jdff dff_B_o9wqmrq05_0(.din(n568),.dout(w_dff_B_o9wqmrq05_0),.clk(gclk));
	jdff dff_B_xVPcu1ND6_2(.din(n565),.dout(w_dff_B_xVPcu1ND6_2),.clk(gclk));
	jdff dff_B_41Caj17Y1_2(.din(w_dff_B_xVPcu1ND6_2),.dout(w_dff_B_41Caj17Y1_2),.clk(gclk));
	jdff dff_B_LjJcccF96_2(.din(w_dff_B_41Caj17Y1_2),.dout(w_dff_B_LjJcccF96_2),.clk(gclk));
	jdff dff_B_GzgNPC5e4_2(.din(w_dff_B_LjJcccF96_2),.dout(w_dff_B_GzgNPC5e4_2),.clk(gclk));
	jdff dff_B_fW9xPb2b1_2(.din(w_dff_B_GzgNPC5e4_2),.dout(w_dff_B_fW9xPb2b1_2),.clk(gclk));
	jdff dff_B_s6fuivb63_2(.din(w_dff_B_fW9xPb2b1_2),.dout(w_dff_B_s6fuivb63_2),.clk(gclk));
	jdff dff_B_EOIIpEcT9_2(.din(w_dff_B_s6fuivb63_2),.dout(w_dff_B_EOIIpEcT9_2),.clk(gclk));
	jdff dff_B_QnSeoWhd6_2(.din(w_dff_B_EOIIpEcT9_2),.dout(w_dff_B_QnSeoWhd6_2),.clk(gclk));
	jdff dff_B_YLlFhacG2_2(.din(w_dff_B_QnSeoWhd6_2),.dout(w_dff_B_YLlFhacG2_2),.clk(gclk));
	jdff dff_B_ZYb40iFp0_0(.din(n1161),.dout(w_dff_B_ZYb40iFp0_0),.clk(gclk));
	jdff dff_B_h4RtadRs5_0(.din(w_dff_B_ZYb40iFp0_0),.dout(w_dff_B_h4RtadRs5_0),.clk(gclk));
	jdff dff_B_b1pGu6vw9_0(.din(w_dff_B_h4RtadRs5_0),.dout(w_dff_B_b1pGu6vw9_0),.clk(gclk));
	jdff dff_B_nGgjxvac3_0(.din(n1158),.dout(w_dff_B_nGgjxvac3_0),.clk(gclk));
	jdff dff_B_QsZcq38y8_0(.din(w_dff_B_nGgjxvac3_0),.dout(w_dff_B_QsZcq38y8_0),.clk(gclk));
	jdff dff_B_K6EzFokF1_0(.din(w_dff_B_QsZcq38y8_0),.dout(w_dff_B_K6EzFokF1_0),.clk(gclk));
	jdff dff_B_b4TGWIg46_0(.din(w_dff_B_K6EzFokF1_0),.dout(w_dff_B_b4TGWIg46_0),.clk(gclk));
	jdff dff_B_0KBgtigG8_1(.din(n1154),.dout(w_dff_B_0KBgtigG8_1),.clk(gclk));
	jdff dff_B_SAV4Uvhx7_1(.din(w_dff_B_0KBgtigG8_1),.dout(w_dff_B_SAV4Uvhx7_1),.clk(gclk));
	jdff dff_B_7jyzD58J2_0(.din(n1155),.dout(w_dff_B_7jyzD58J2_0),.clk(gclk));
	jdff dff_B_eRCI9hCc9_0(.din(w_dff_B_7jyzD58J2_0),.dout(w_dff_B_eRCI9hCc9_0),.clk(gclk));
	jdff dff_B_0E64AsKd0_1(.din(n1145),.dout(w_dff_B_0E64AsKd0_1),.clk(gclk));
	jdff dff_B_uRqsTUXW5_1(.din(n1148),.dout(w_dff_B_uRqsTUXW5_1),.clk(gclk));
	jdff dff_A_kiZ2YnPA2_1(.dout(w_G87_1[1]),.din(w_dff_A_kiZ2YnPA2_1),.clk(gclk));
	jdff dff_A_o4LQQvKM3_2(.dout(w_G87_1[2]),.din(w_dff_A_o4LQQvKM3_2),.clk(gclk));
	jdff dff_A_SNqBWfVJ2_1(.dout(w_G77_2[1]),.din(w_dff_A_SNqBWfVJ2_1),.clk(gclk));
	jdff dff_A_iJUgBwq71_1(.dout(w_dff_A_SNqBWfVJ2_1),.din(w_dff_A_iJUgBwq71_1),.clk(gclk));
	jdff dff_A_7p48mYnV6_1(.dout(w_dff_A_iJUgBwq71_1),.din(w_dff_A_7p48mYnV6_1),.clk(gclk));
	jdff dff_A_hPLRTLOf3_1(.dout(w_dff_A_7p48mYnV6_1),.din(w_dff_A_hPLRTLOf3_1),.clk(gclk));
	jdff dff_A_WVhOwAHD2_2(.dout(w_G77_2[2]),.din(w_dff_A_WVhOwAHD2_2),.clk(gclk));
	jdff dff_A_z6SlBdM10_2(.dout(w_dff_A_WVhOwAHD2_2),.din(w_dff_A_z6SlBdM10_2),.clk(gclk));
	jdff dff_A_OWA3kIlo0_2(.dout(w_dff_A_z6SlBdM10_2),.din(w_dff_A_OWA3kIlo0_2),.clk(gclk));
	jdff dff_A_59ogoqPM0_2(.dout(w_dff_A_OWA3kIlo0_2),.din(w_dff_A_59ogoqPM0_2),.clk(gclk));
	jdff dff_A_b5r1Lzgn7_0(.dout(w_n148_3[0]),.din(w_dff_A_b5r1Lzgn7_0),.clk(gclk));
	jdff dff_A_UT8H2Vic3_0(.dout(w_dff_A_b5r1Lzgn7_0),.din(w_dff_A_UT8H2Vic3_0),.clk(gclk));
	jdff dff_A_Wbs76ppA6_0(.dout(w_dff_A_UT8H2Vic3_0),.din(w_dff_A_Wbs76ppA6_0),.clk(gclk));
	jdff dff_A_8hHkL1PG3_2(.dout(w_n148_3[2]),.din(w_dff_A_8hHkL1PG3_2),.clk(gclk));
	jdff dff_A_CSZbFV0d2_2(.dout(w_dff_A_8hHkL1PG3_2),.din(w_dff_A_CSZbFV0d2_2),.clk(gclk));
	jdff dff_A_eoz6teQ20_2(.dout(w_dff_A_CSZbFV0d2_2),.din(w_dff_A_eoz6teQ20_2),.clk(gclk));
	jdff dff_B_DktmHrQx5_0(.din(n1142),.dout(w_dff_B_DktmHrQx5_0),.clk(gclk));
	jdff dff_B_sOcuBiPH3_1(.din(n1130),.dout(w_dff_B_sOcuBiPH3_1),.clk(gclk));
	jdff dff_B_Q1qvxK2L3_1(.din(n1133),.dout(w_dff_B_Q1qvxK2L3_1),.clk(gclk));
	jdff dff_B_IdjcOSiq5_0(.din(n1134),.dout(w_dff_B_IdjcOSiq5_0),.clk(gclk));
	jdff dff_A_jy5KOk1X7_1(.dout(w_G150_1[1]),.din(w_dff_A_jy5KOk1X7_1),.clk(gclk));
	jdff dff_A_H7I5RNYx4_2(.dout(w_G150_1[2]),.din(w_dff_A_H7I5RNYx4_2),.clk(gclk));
	jdff dff_B_AS6caYQk9_3(.din(G128),.dout(w_dff_B_AS6caYQk9_3),.clk(gclk));
	jdff dff_B_iav8vIDC0_3(.din(w_dff_B_AS6caYQk9_3),.dout(w_dff_B_iav8vIDC0_3),.clk(gclk));
	jdff dff_B_k4zStVQl6_3(.din(w_dff_B_iav8vIDC0_3),.dout(w_dff_B_k4zStVQl6_3),.clk(gclk));
	jdff dff_B_bC9jIfkQ7_0(.din(n1126),.dout(w_dff_B_bC9jIfkQ7_0),.clk(gclk));
	jdff dff_A_RufEhbVX7_0(.dout(w_n612_1[0]),.din(w_dff_A_RufEhbVX7_0),.clk(gclk));
	jdff dff_A_oTtkGiLK7_0(.dout(w_dff_A_RufEhbVX7_0),.din(w_dff_A_oTtkGiLK7_0),.clk(gclk));
	jdff dff_A_Mwr1h53n1_1(.dout(w_n612_1[1]),.din(w_dff_A_Mwr1h53n1_1),.clk(gclk));
	jdff dff_A_X7KaqByy2_1(.dout(w_dff_A_Mwr1h53n1_1),.din(w_dff_A_X7KaqByy2_1),.clk(gclk));
	jdff dff_A_8Zb4vVrW1_1(.dout(w_dff_A_X7KaqByy2_1),.din(w_dff_A_8Zb4vVrW1_1),.clk(gclk));
	jdff dff_A_QCOAP4Qk2_1(.dout(w_dff_A_8Zb4vVrW1_1),.din(w_dff_A_QCOAP4Qk2_1),.clk(gclk));
	jdff dff_B_gY9f2nnX4_0(.din(n1118),.dout(w_dff_B_gY9f2nnX4_0),.clk(gclk));
	jdff dff_A_4Oz5YSYp3_1(.dout(w_n1002_0[1]),.din(w_dff_A_4Oz5YSYp3_1),.clk(gclk));
	jdff dff_A_zob0P3cI5_2(.dout(w_n1002_0[2]),.din(w_dff_A_zob0P3cI5_2),.clk(gclk));
	jdff dff_B_gbC0DPc77_1(.din(n998),.dout(w_dff_B_gbC0DPc77_1),.clk(gclk));
	jdff dff_A_85GgCVqu2_1(.dout(w_n999_0[1]),.din(w_dff_A_85GgCVqu2_1),.clk(gclk));
	jdff dff_A_eAk7lmmX5_1(.dout(w_dff_A_85GgCVqu2_1),.din(w_dff_A_eAk7lmmX5_1),.clk(gclk));
	jdff dff_A_zbujm7Tb4_2(.dout(w_n764_0[2]),.din(w_dff_A_zbujm7Tb4_2),.clk(gclk));
	jdff dff_A_IBJkRmJa1_2(.dout(w_dff_A_zbujm7Tb4_2),.din(w_dff_A_IBJkRmJa1_2),.clk(gclk));
	jdff dff_A_DPRKpDgj8_2(.dout(w_dff_A_IBJkRmJa1_2),.din(w_dff_A_DPRKpDgj8_2),.clk(gclk));
	jdff dff_B_gqoWoSKU3_0(.din(n763),.dout(w_dff_B_gqoWoSKU3_0),.clk(gclk));
	jdff dff_B_0ZIerqGo2_0(.din(w_dff_B_gqoWoSKU3_0),.dout(w_dff_B_0ZIerqGo2_0),.clk(gclk));
	jdff dff_B_yJpCBKoX8_0(.din(n761),.dout(w_dff_B_yJpCBKoX8_0),.clk(gclk));
	jdff dff_B_CKoaYjSd0_0(.din(w_dff_B_yJpCBKoX8_0),.dout(w_dff_B_CKoaYjSd0_0),.clk(gclk));
	jdff dff_A_MKuYlg0D3_0(.dout(w_n760_0[0]),.din(w_dff_A_MKuYlg0D3_0),.clk(gclk));
	jdff dff_A_vvO22FOj2_1(.dout(w_n553_1[1]),.din(w_dff_A_vvO22FOj2_1),.clk(gclk));
	jdff dff_A_sWmskyep9_1(.dout(w_dff_A_vvO22FOj2_1),.din(w_dff_A_sWmskyep9_1),.clk(gclk));
	jdff dff_A_daKAvAwE4_1(.dout(w_dff_A_sWmskyep9_1),.din(w_dff_A_daKAvAwE4_1),.clk(gclk));
	jdff dff_B_keav1kmT0_0(.din(n997),.dout(w_dff_B_keav1kmT0_0),.clk(gclk));
	jdff dff_B_dqgSnqHA1_0(.din(w_dff_B_keav1kmT0_0),.dout(w_dff_B_dqgSnqHA1_0),.clk(gclk));
	jdff dff_B_3fZRx6RI2_0(.din(w_dff_B_dqgSnqHA1_0),.dout(w_dff_B_3fZRx6RI2_0),.clk(gclk));
	jdff dff_B_FImqC54b9_0(.din(w_dff_B_3fZRx6RI2_0),.dout(w_dff_B_FImqC54b9_0),.clk(gclk));
	jdff dff_B_JCQfpg1X7_0(.din(w_dff_B_FImqC54b9_0),.dout(w_dff_B_JCQfpg1X7_0),.clk(gclk));
	jdff dff_A_rWWVvxsJ8_0(.dout(w_n996_0[0]),.din(w_dff_A_rWWVvxsJ8_0),.clk(gclk));
	jdff dff_A_k3JGA4C40_0(.dout(w_dff_A_rWWVvxsJ8_0),.din(w_dff_A_k3JGA4C40_0),.clk(gclk));
	jdff dff_A_EeZjSg887_2(.dout(w_n996_0[2]),.din(w_dff_A_EeZjSg887_2),.clk(gclk));
	jdff dff_A_4NmqG9wv9_2(.dout(w_dff_A_EeZjSg887_2),.din(w_dff_A_4NmqG9wv9_2),.clk(gclk));
	jdff dff_B_pVqq1Jlu5_1(.din(n447),.dout(w_dff_B_pVqq1Jlu5_1),.clk(gclk));
	jdff dff_B_t0VQJmnK4_2(.din(n517),.dout(w_dff_B_t0VQJmnK4_2),.clk(gclk));
	jdff dff_A_VTeMM7ch9_0(.dout(w_n484_0[0]),.din(w_dff_A_VTeMM7ch9_0),.clk(gclk));
	jdff dff_B_qU8NM3Dz0_3(.din(n548),.dout(w_dff_B_qU8NM3Dz0_3),.clk(gclk));
	jdff dff_B_nrXDqPfL0_3(.din(w_dff_B_qU8NM3Dz0_3),.dout(w_dff_B_nrXDqPfL0_3),.clk(gclk));
	jdff dff_B_c69DTJYd0_3(.din(w_dff_B_nrXDqPfL0_3),.dout(w_dff_B_c69DTJYd0_3),.clk(gclk));
	jdff dff_A_7AYaMK7Q9_1(.dout(w_n439_0[1]),.din(w_dff_A_7AYaMK7Q9_1),.clk(gclk));
	jdff dff_A_nYsWf3yJ0_1(.dout(w_dff_A_7AYaMK7Q9_1),.din(w_dff_A_nYsWf3yJ0_1),.clk(gclk));
	jdff dff_A_oAWWLL5M1_1(.dout(w_dff_A_nYsWf3yJ0_1),.din(w_dff_A_oAWWLL5M1_1),.clk(gclk));
	jdff dff_B_t6Zcu4g47_0(.din(n437),.dout(w_dff_B_t6Zcu4g47_0),.clk(gclk));
	jdff dff_A_1LTuX2rb6_1(.dout(w_n445_0[1]),.din(w_dff_A_1LTuX2rb6_1),.clk(gclk));
	jdff dff_B_TtNazLUZ4_2(.din(n445),.dout(w_dff_B_TtNazLUZ4_2),.clk(gclk));
	jdff dff_B_Klqcwm7I2_2(.din(w_dff_B_TtNazLUZ4_2),.dout(w_dff_B_Klqcwm7I2_2),.clk(gclk));
	jdff dff_B_E2pzOZt54_1(.din(n424),.dout(w_dff_B_E2pzOZt54_1),.clk(gclk));
	jdff dff_B_k6F7bK6c4_0(.din(n434),.dout(w_dff_B_k6F7bK6c4_0),.clk(gclk));
	jdff dff_B_5R6QWDEa2_0(.din(n423),.dout(w_dff_B_5R6QWDEa2_0),.clk(gclk));
	jdff dff_A_8yy2zotn6_0(.dout(w_G226_1[0]),.din(w_dff_A_8yy2zotn6_0),.clk(gclk));
	jdff dff_A_Ntvkszga7_0(.dout(w_dff_A_8yy2zotn6_0),.din(w_dff_A_Ntvkszga7_0),.clk(gclk));
	jdff dff_A_JFkCUEOJ0_0(.dout(w_n542_0[0]),.din(w_dff_A_JFkCUEOJ0_0),.clk(gclk));
	jdff dff_A_95QQxCPE3_1(.dout(w_n511_0[1]),.din(w_dff_A_95QQxCPE3_1),.clk(gclk));
	jdff dff_B_CB45gDrB0_1(.din(n493),.dout(w_dff_B_CB45gDrB0_1),.clk(gclk));
	jdff dff_B_EmiIeIdo0_1(.din(w_dff_B_CB45gDrB0_1),.dout(w_dff_B_EmiIeIdo0_1),.clk(gclk));
	jdff dff_B_vYoGX6kR4_0(.din(n509),.dout(w_dff_B_vYoGX6kR4_0),.clk(gclk));
	jdff dff_B_15Lwp3E76_0(.din(n515),.dout(w_dff_B_15Lwp3E76_0),.clk(gclk));
	jdff dff_B_KhwKB54G4_0(.din(w_dff_B_15Lwp3E76_0),.dout(w_dff_B_KhwKB54G4_0),.clk(gclk));
	jdff dff_B_FtEUyvTn6_0(.din(n514),.dout(w_dff_B_FtEUyvTn6_0),.clk(gclk));
	jdff dff_B_h0wBLRfa5_1(.din(n496),.dout(w_dff_B_h0wBLRfa5_1),.clk(gclk));
	jdff dff_B_aC3Hupml5_1(.din(w_dff_B_h0wBLRfa5_1),.dout(w_dff_B_aC3Hupml5_1),.clk(gclk));
	jdff dff_B_5hryCipb2_1(.din(w_dff_B_aC3Hupml5_1),.dout(w_dff_B_5hryCipb2_1),.clk(gclk));
	jdff dff_B_S3vy7CbM2_1(.din(n497),.dout(w_dff_B_S3vy7CbM2_1),.clk(gclk));
	jdff dff_B_g84FQDWf9_1(.din(w_dff_B_S3vy7CbM2_1),.dout(w_dff_B_g84FQDWf9_1),.clk(gclk));
	jdff dff_B_kcBHfiiB6_1(.din(w_dff_B_g84FQDWf9_1),.dout(w_dff_B_kcBHfiiB6_1),.clk(gclk));
	jdff dff_A_KqevKNcd0_0(.dout(w_n541_0[0]),.din(w_dff_A_KqevKNcd0_0),.clk(gclk));
	jdff dff_A_fGoUnq7h8_1(.dout(w_n478_0[1]),.din(w_dff_A_fGoUnq7h8_1),.clk(gclk));
	jdff dff_B_FuPue6fb6_1(.din(n456),.dout(w_dff_B_FuPue6fb6_1),.clk(gclk));
	jdff dff_B_S22Biev41_1(.din(w_dff_B_FuPue6fb6_1),.dout(w_dff_B_S22Biev41_1),.clk(gclk));
	jdff dff_B_BszKyM8a9_1(.din(w_dff_B_S22Biev41_1),.dout(w_dff_B_BszKyM8a9_1),.clk(gclk));
	jdff dff_B_TgVEMjNG0_0(.din(n476),.dout(w_dff_B_TgVEMjNG0_0),.clk(gclk));
	jdff dff_B_C3Zh2WT72_0(.din(w_dff_B_TgVEMjNG0_0),.dout(w_dff_B_C3Zh2WT72_0),.clk(gclk));
	jdff dff_B_9Fy2kyov4_0(.din(n482),.dout(w_dff_B_9Fy2kyov4_0),.clk(gclk));
	jdff dff_B_f1dpro7X6_0(.din(w_dff_B_9Fy2kyov4_0),.dout(w_dff_B_f1dpro7X6_0),.clk(gclk));
	jdff dff_B_eUERuVKn4_0(.din(w_dff_B_f1dpro7X6_0),.dout(w_dff_B_eUERuVKn4_0),.clk(gclk));
	jdff dff_B_pmKtcmWA5_0(.din(n481),.dout(w_dff_B_pmKtcmWA5_0),.clk(gclk));
	jdff dff_A_0RGvImsv3_1(.dout(w_G226_0[1]),.din(w_dff_A_0RGvImsv3_1),.clk(gclk));
	jdff dff_A_JJ9RWBLE3_1(.dout(w_dff_A_0RGvImsv3_1),.din(w_dff_A_JJ9RWBLE3_1),.clk(gclk));
	jdff dff_A_yJJP5N8H3_2(.dout(w_G226_0[2]),.din(w_dff_A_yJJP5N8H3_2),.clk(gclk));
	jdff dff_A_4Fk1I7i19_2(.dout(w_dff_A_yJJP5N8H3_2),.din(w_dff_A_4Fk1I7i19_2),.clk(gclk));
	jdff dff_A_uQxop5AO8_2(.dout(w_dff_A_4Fk1I7i19_2),.din(w_dff_A_uQxop5AO8_2),.clk(gclk));
	jdff dff_B_PDdmklrm3_1(.din(G222),.dout(w_dff_B_PDdmklrm3_1),.clk(gclk));
	jdff dff_B_HLS7OORf1_1(.din(w_dff_B_PDdmklrm3_1),.dout(w_dff_B_HLS7OORf1_1),.clk(gclk));
	jdff dff_A_oye51Lho7_0(.dout(w_n430_0[0]),.din(w_dff_A_oye51Lho7_0),.clk(gclk));
	jdff dff_B_YFNG28sK1_2(.din(n430),.dout(w_dff_B_YFNG28sK1_2),.clk(gclk));
	jdff dff_A_zymzxxtQ7_1(.dout(w_G77_3[1]),.din(w_dff_A_zymzxxtQ7_1),.clk(gclk));
	jdff dff_A_65LzyoxR2_1(.dout(w_dff_A_zymzxxtQ7_1),.din(w_dff_A_65LzyoxR2_1),.clk(gclk));
	jdff dff_A_ptzGm7K20_1(.dout(w_dff_A_65LzyoxR2_1),.din(w_dff_A_ptzGm7K20_1),.clk(gclk));
	jdff dff_B_nDVKlNPf1_2(.din(G223),.dout(w_dff_B_nDVKlNPf1_2),.clk(gclk));
	jdff dff_B_El1Kyins8_2(.din(w_dff_B_nDVKlNPf1_2),.dout(w_dff_B_El1Kyins8_2),.clk(gclk));
	jdff dff_B_EQkryD4M1_1(.din(n459),.dout(w_dff_B_EQkryD4M1_1),.clk(gclk));
	jdff dff_B_pWjzjc0O5_1(.din(w_dff_B_EQkryD4M1_1),.dout(w_dff_B_pWjzjc0O5_1),.clk(gclk));
	jdff dff_B_Tvnatg297_1(.din(w_dff_B_pWjzjc0O5_1),.dout(w_dff_B_Tvnatg297_1),.clk(gclk));
	jdff dff_B_DwUkk4SC4_1(.din(w_dff_B_Tvnatg297_1),.dout(w_dff_B_DwUkk4SC4_1),.clk(gclk));
	jdff dff_B_Nvo7ve6m3_0(.din(n472),.dout(w_dff_B_Nvo7ve6m3_0),.clk(gclk));
	jdff dff_A_20GyYu6S9_2(.dout(w_n185_1[2]),.din(w_dff_A_20GyYu6S9_2),.clk(gclk));
	jdff dff_B_RecgrcfT2_1(.din(n460),.dout(w_dff_B_RecgrcfT2_1),.clk(gclk));
	jdff dff_B_INQMja0C0_1(.din(w_dff_B_RecgrcfT2_1),.dout(w_dff_B_INQMja0C0_1),.clk(gclk));
	jdff dff_B_LIelNfwt4_1(.din(n464),.dout(w_dff_B_LIelNfwt4_1),.clk(gclk));
	jdff dff_B_04N51c2S8_1(.din(n461),.dout(w_dff_B_04N51c2S8_1),.clk(gclk));
	jdff dff_B_vha6vETx4_1(.din(w_dff_B_04N51c2S8_1),.dout(w_dff_B_vha6vETx4_1),.clk(gclk));
	jdff dff_A_74Wh4UtW0_1(.dout(w_n75_0[1]),.din(w_dff_A_74Wh4UtW0_1),.clk(gclk));
	jdff dff_A_rIxLrDBm1_1(.dout(w_dff_A_74Wh4UtW0_1),.din(w_dff_A_rIxLrDBm1_1),.clk(gclk));
	jdff dff_A_t7kP4Kj38_1(.dout(w_dff_A_rIxLrDBm1_1),.din(w_dff_A_t7kP4Kj38_1),.clk(gclk));
	jdff dff_A_1XGtQpBl9_2(.dout(w_n75_0[2]),.din(w_dff_A_1XGtQpBl9_2),.clk(gclk));
	jdff dff_A_GjChyxxK5_2(.dout(w_dff_A_1XGtQpBl9_2),.din(w_dff_A_GjChyxxK5_2),.clk(gclk));
	jdff dff_A_nj2QBwlE1_2(.dout(w_dff_A_GjChyxxK5_2),.din(w_dff_A_nj2QBwlE1_2),.clk(gclk));
	jdff dff_A_gov1gbCz0_1(.dout(w_n74_0[1]),.din(w_dff_A_gov1gbCz0_1),.clk(gclk));
	jdff dff_A_hqL2N1gy3_1(.dout(w_dff_A_gov1gbCz0_1),.din(w_dff_A_hqL2N1gy3_1),.clk(gclk));
	jdff dff_A_b7CJdTKD3_1(.dout(w_dff_A_hqL2N1gy3_1),.din(w_dff_A_b7CJdTKD3_1),.clk(gclk));
	jdff dff_A_nQKuoKeb7_2(.dout(w_n74_0[2]),.din(w_dff_A_nQKuoKeb7_2),.clk(gclk));
	jdff dff_A_zQKuk2nr8_2(.dout(w_dff_A_nQKuoKeb7_2),.din(w_dff_A_zQKuk2nr8_2),.clk(gclk));
	jdff dff_A_kd5ECbCg6_0(.dout(w_n73_2[0]),.din(w_dff_A_kd5ECbCg6_0),.clk(gclk));
	jdff dff_A_LiCi63DK0_0(.dout(w_dff_A_kd5ECbCg6_0),.din(w_dff_A_LiCi63DK0_0),.clk(gclk));
	jdff dff_A_VnmzGIqZ9_2(.dout(w_n73_2[2]),.din(w_dff_A_VnmzGIqZ9_2),.clk(gclk));
	jdff dff_A_qP0PjycH7_2(.dout(w_n73_0[2]),.din(w_dff_A_qP0PjycH7_2),.clk(gclk));
	jdff dff_A_qcAqNnII1_2(.dout(w_dff_A_qP0PjycH7_2),.din(w_dff_A_qcAqNnII1_2),.clk(gclk));
	jdff dff_A_R2ndmZqm6_2(.dout(w_dff_A_qcAqNnII1_2),.din(w_dff_A_R2ndmZqm6_2),.clk(gclk));
	jdff dff_A_0BjMtfxy1_1(.dout(w_G50_5[1]),.din(w_dff_A_0BjMtfxy1_1),.clk(gclk));
	jdff dff_A_XRyOIwwU7_1(.dout(w_dff_A_0BjMtfxy1_1),.din(w_dff_A_XRyOIwwU7_1),.clk(gclk));
	jdff dff_A_zBQyaB0w2_1(.dout(w_dff_A_XRyOIwwU7_1),.din(w_dff_A_zBQyaB0w2_1),.clk(gclk));
	jdff dff_A_jW3dfybX5_0(.dout(w_G50_4[0]),.din(w_dff_A_jW3dfybX5_0),.clk(gclk));
	jdff dff_A_ldFcLSv06_0(.dout(w_dff_A_jW3dfybX5_0),.din(w_dff_A_ldFcLSv06_0),.clk(gclk));
	jdff dff_A_ps1pBBQg0_0(.dout(w_G50_1[0]),.din(w_dff_A_ps1pBBQg0_0),.clk(gclk));
	jdff dff_A_NlNqZx0B9_2(.dout(w_G50_1[2]),.din(w_dff_A_NlNqZx0B9_2),.clk(gclk));
	jdff dff_A_NpK6idSS1_2(.dout(w_dff_A_NlNqZx0B9_2),.din(w_dff_A_NpK6idSS1_2),.clk(gclk));
	jdff dff_A_cDRNt68D6_2(.dout(w_dff_A_NpK6idSS1_2),.din(w_dff_A_cDRNt68D6_2),.clk(gclk));
	jdff dff_A_bhT07Qpo8_2(.dout(w_dff_A_cDRNt68D6_2),.din(w_dff_A_bhT07Qpo8_2),.clk(gclk));
	jdff dff_A_6b4CzQnG1_0(.dout(w_G384_0),.din(w_dff_A_6b4CzQnG1_0),.clk(gclk));
	jdff dff_A_95tQa7W18_0(.dout(w_dff_A_6b4CzQnG1_0),.din(w_dff_A_95tQa7W18_0),.clk(gclk));
	jdff dff_A_eed2vNmR3_0(.dout(w_dff_A_95tQa7W18_0),.din(w_dff_A_eed2vNmR3_0),.clk(gclk));
	jdff dff_B_PYzOnq4l7_0(.din(n747),.dout(w_dff_B_PYzOnq4l7_0),.clk(gclk));
	jdff dff_B_UFkzWYqI2_0(.din(n746),.dout(w_dff_B_UFkzWYqI2_0),.clk(gclk));
	jdff dff_B_g093PoJh8_0(.din(w_dff_B_UFkzWYqI2_0),.dout(w_dff_B_g093PoJh8_0),.clk(gclk));
	jdff dff_B_k4AlFgau3_0(.din(w_dff_B_g093PoJh8_0),.dout(w_dff_B_k4AlFgau3_0),.clk(gclk));
	jdff dff_B_5JxwEWcx5_0(.din(n744),.dout(w_dff_B_5JxwEWcx5_0),.clk(gclk));
	jdff dff_B_XuRRvTNa2_0(.din(w_dff_B_5JxwEWcx5_0),.dout(w_dff_B_XuRRvTNa2_0),.clk(gclk));
	jdff dff_A_1UvET2Be9_2(.dout(w_n605_1[2]),.din(w_dff_A_1UvET2Be9_2),.clk(gclk));
	jdff dff_A_efUUGvLH3_2(.dout(w_dff_A_1UvET2Be9_2),.din(w_dff_A_efUUGvLH3_2),.clk(gclk));
	jdff dff_A_zYsdWECT7_2(.dout(w_dff_A_efUUGvLH3_2),.din(w_dff_A_zYsdWECT7_2),.clk(gclk));
	jdff dff_A_XTfzI8En2_0(.dout(w_n604_2[0]),.din(w_dff_A_XTfzI8En2_0),.clk(gclk));
	jdff dff_A_EHw4u9ai4_0(.dout(w_dff_A_XTfzI8En2_0),.din(w_dff_A_EHw4u9ai4_0),.clk(gclk));
	jdff dff_B_VEDtvJyM9_1(.din(n721),.dout(w_dff_B_VEDtvJyM9_1),.clk(gclk));
	jdff dff_B_52MHcjgq9_1(.din(w_dff_B_VEDtvJyM9_1),.dout(w_dff_B_52MHcjgq9_1),.clk(gclk));
	jdff dff_B_h4Y4CTa98_1(.din(w_dff_B_52MHcjgq9_1),.dout(w_dff_B_h4Y4CTa98_1),.clk(gclk));
	jdff dff_B_YUqIbko90_1(.din(w_dff_B_h4Y4CTa98_1),.dout(w_dff_B_YUqIbko90_1),.clk(gclk));
	jdff dff_B_2tEorJjR7_1(.din(w_dff_B_YUqIbko90_1),.dout(w_dff_B_2tEorJjR7_1),.clk(gclk));
	jdff dff_B_qy7Dk0eB1_1(.din(n727),.dout(w_dff_B_qy7Dk0eB1_1),.clk(gclk));
	jdff dff_B_3P2caIMQ0_1(.din(w_dff_B_qy7Dk0eB1_1),.dout(w_dff_B_3P2caIMQ0_1),.clk(gclk));
	jdff dff_B_S29NIsBY5_0(.din(n737),.dout(w_dff_B_S29NIsBY5_0),.clk(gclk));
	jdff dff_B_nCwovcnt8_1(.din(n733),.dout(w_dff_B_nCwovcnt8_1),.clk(gclk));
	jdff dff_B_Zrtp0TWN6_0(.din(n734),.dout(w_dff_B_Zrtp0TWN6_0),.clk(gclk));
	jdff dff_A_Ec9Kqgjw8_0(.dout(w_G294_2[0]),.din(w_dff_A_Ec9Kqgjw8_0),.clk(gclk));
	jdff dff_A_8kX5hHrJ2_0(.dout(w_G116_3[0]),.din(w_dff_A_8kX5hHrJ2_0),.clk(gclk));
	jdff dff_A_QW2IITbk9_0(.dout(w_dff_A_8kX5hHrJ2_0),.din(w_dff_A_QW2IITbk9_0),.clk(gclk));
	jdff dff_A_Ul9C7h3E4_0(.dout(w_dff_A_QW2IITbk9_0),.din(w_dff_A_Ul9C7h3E4_0),.clk(gclk));
	jdff dff_A_nTi7pOJZ7_2(.dout(w_G116_3[2]),.din(w_dff_A_nTi7pOJZ7_2),.clk(gclk));
	jdff dff_A_aVf2RN5x9_2(.dout(w_dff_A_nTi7pOJZ7_2),.din(w_dff_A_aVf2RN5x9_2),.clk(gclk));
	jdff dff_A_BIlKLNuA7_2(.dout(w_G33_5[2]),.din(w_dff_A_BIlKLNuA7_2),.clk(gclk));
	jdff dff_A_KLAYTlk53_2(.dout(w_dff_A_BIlKLNuA7_2),.din(w_dff_A_KLAYTlk53_2),.clk(gclk));
	jdff dff_B_DQhw4aS97_1(.din(n722),.dout(w_dff_B_DQhw4aS97_1),.clk(gclk));
	jdff dff_B_5ccDlyQl1_0(.din(n724),.dout(w_dff_B_5ccDlyQl1_0),.clk(gclk));
	jdff dff_B_KDY4NsUX0_3(.din(G311),.dout(w_dff_B_KDY4NsUX0_3),.clk(gclk));
	jdff dff_B_pMMLIfB61_3(.din(w_dff_B_KDY4NsUX0_3),.dout(w_dff_B_pMMLIfB61_3),.clk(gclk));
	jdff dff_B_p5xIi9sp7_3(.din(w_dff_B_pMMLIfB61_3),.dout(w_dff_B_p5xIi9sp7_3),.clk(gclk));
	jdff dff_B_86WmmvN65_1(.din(n715),.dout(w_dff_B_86WmmvN65_1),.clk(gclk));
	jdff dff_B_MdgUWO5j9_1(.din(n716),.dout(w_dff_B_MdgUWO5j9_1),.clk(gclk));
	jdff dff_A_13t7fpQR2_1(.dout(w_G68_3[1]),.din(w_dff_A_13t7fpQR2_1),.clk(gclk));
	jdff dff_A_JhIdS5Fe6_1(.dout(w_dff_A_13t7fpQR2_1),.din(w_dff_A_JhIdS5Fe6_1),.clk(gclk));
	jdff dff_A_wLrENlk49_1(.dout(w_dff_A_JhIdS5Fe6_1),.din(w_dff_A_wLrENlk49_1),.clk(gclk));
	jdff dff_A_VoSx3bgd5_2(.dout(w_G68_3[2]),.din(w_dff_A_VoSx3bgd5_2),.clk(gclk));
	jdff dff_A_i2IVPP7p7_2(.dout(w_dff_A_VoSx3bgd5_2),.din(w_dff_A_i2IVPP7p7_2),.clk(gclk));
	jdff dff_B_x6nOYpLm4_3(.din(G137),.dout(w_dff_B_x6nOYpLm4_3),.clk(gclk));
	jdff dff_B_8WysDD1G7_3(.din(w_dff_B_x6nOYpLm4_3),.dout(w_dff_B_8WysDD1G7_3),.clk(gclk));
	jdff dff_B_PhCYIDkf7_3(.din(w_dff_B_8WysDD1G7_3),.dout(w_dff_B_PhCYIDkf7_3),.clk(gclk));
	jdff dff_B_JVT5tKHq1_3(.din(G143),.dout(w_dff_B_JVT5tKHq1_3),.clk(gclk));
	jdff dff_B_4B88tn5x2_3(.din(w_dff_B_JVT5tKHq1_3),.dout(w_dff_B_4B88tn5x2_3),.clk(gclk));
	jdff dff_B_t5fzPJDL5_3(.din(w_dff_B_4B88tn5x2_3),.dout(w_dff_B_t5fzPJDL5_3),.clk(gclk));
	jdff dff_A_Ct00FSky8_0(.dout(w_G159_3[0]),.din(w_dff_A_Ct00FSky8_0),.clk(gclk));
	jdff dff_A_d7nwO7Jr9_1(.dout(w_G159_3[1]),.din(w_dff_A_d7nwO7Jr9_1),.clk(gclk));
	jdff dff_A_XSqLkxZc8_0(.dout(w_G159_0[0]),.din(w_dff_A_XSqLkxZc8_0),.clk(gclk));
	jdff dff_A_Sb91akbp9_0(.dout(w_dff_A_XSqLkxZc8_0),.din(w_dff_A_Sb91akbp9_0),.clk(gclk));
	jdff dff_A_7A7o9IQa1_1(.dout(w_G159_0[1]),.din(w_dff_A_7A7o9IQa1_1),.clk(gclk));
	jdff dff_B_1kwtdeLX0_3(.din(G159),.dout(w_dff_B_1kwtdeLX0_3),.clk(gclk));
	jdff dff_B_GuEHFn4Z5_3(.din(w_dff_B_1kwtdeLX0_3),.dout(w_dff_B_GuEHFn4Z5_3),.clk(gclk));
	jdff dff_A_uKnjDzBp6_1(.dout(w_G190_2[1]),.din(w_dff_A_uKnjDzBp6_1),.clk(gclk));
	jdff dff_A_Ey0AHIns3_1(.dout(w_dff_A_uKnjDzBp6_1),.din(w_dff_A_Ey0AHIns3_1),.clk(gclk));
	jdff dff_A_fCkOyNJy8_2(.dout(w_G190_2[2]),.din(w_dff_A_fCkOyNJy8_2),.clk(gclk));
	jdff dff_A_sNGWQ4tz3_2(.dout(w_dff_A_fCkOyNJy8_2),.din(w_dff_A_sNGWQ4tz3_2),.clk(gclk));
	jdff dff_A_lSokXZRf2_0(.dout(w_G50_3[0]),.din(w_dff_A_lSokXZRf2_0),.clk(gclk));
	jdff dff_A_1Wr1bQN09_0(.dout(w_dff_A_lSokXZRf2_0),.din(w_dff_A_1Wr1bQN09_0),.clk(gclk));
	jdff dff_A_0BzWVpQx9_0(.dout(w_dff_A_1Wr1bQN09_0),.din(w_dff_A_0BzWVpQx9_0),.clk(gclk));
	jdff dff_A_TjKxMyW99_2(.dout(w_G50_3[2]),.din(w_dff_A_TjKxMyW99_2),.clk(gclk));
	jdff dff_A_2MWFxzgl8_2(.dout(w_dff_A_TjKxMyW99_2),.din(w_dff_A_2MWFxzgl8_2),.clk(gclk));
	jdff dff_A_SZ6fREAm2_2(.dout(w_dff_A_2MWFxzgl8_2),.din(w_dff_A_SZ6fREAm2_2),.clk(gclk));
	jdff dff_A_sRnO9raa1_2(.dout(w_dff_A_SZ6fREAm2_2),.din(w_dff_A_sRnO9raa1_2),.clk(gclk));
	jdff dff_A_lQFdV4Wy1_1(.dout(w_G50_0[1]),.din(w_dff_A_lQFdV4Wy1_1),.clk(gclk));
	jdff dff_A_ZRrFFLui7_1(.dout(w_dff_A_lQFdV4Wy1_1),.din(w_dff_A_ZRrFFLui7_1),.clk(gclk));
	jdff dff_A_7itG0YhZ9_1(.dout(w_dff_A_ZRrFFLui7_1),.din(w_dff_A_7itG0YhZ9_1),.clk(gclk));
	jdff dff_A_FduOWoSV4_0(.dout(w_G33_6[0]),.din(w_dff_A_FduOWoSV4_0),.clk(gclk));
	jdff dff_A_RswzhSnl3_0(.dout(w_dff_A_FduOWoSV4_0),.din(w_dff_A_RswzhSnl3_0),.clk(gclk));
	jdff dff_A_xXtWINz73_0(.dout(w_dff_A_RswzhSnl3_0),.din(w_dff_A_xXtWINz73_0),.clk(gclk));
	jdff dff_A_RvgJFnRR0_0(.dout(w_dff_A_xXtWINz73_0),.din(w_dff_A_RvgJFnRR0_0),.clk(gclk));
	jdff dff_A_914Uzl4u8_1(.dout(w_G33_6[1]),.din(w_dff_A_914Uzl4u8_1),.clk(gclk));
	jdff dff_A_3m2KYaT92_1(.dout(w_dff_A_914Uzl4u8_1),.din(w_dff_A_3m2KYaT92_1),.clk(gclk));
	jdff dff_A_OFynWe806_1(.dout(w_G33_1[1]),.din(w_dff_A_OFynWe806_1),.clk(gclk));
	jdff dff_A_UiCAF1gL4_1(.dout(w_dff_A_OFynWe806_1),.din(w_dff_A_UiCAF1gL4_1),.clk(gclk));
	jdff dff_A_HlyjsgJx5_1(.dout(w_dff_A_UiCAF1gL4_1),.din(w_dff_A_HlyjsgJx5_1),.clk(gclk));
	jdff dff_B_zPIqeoSO7_1(.din(n706),.dout(w_dff_B_zPIqeoSO7_1),.clk(gclk));
	jdff dff_B_iNLtdpIO2_0(.din(n708),.dout(w_dff_B_iNLtdpIO2_0),.clk(gclk));
	jdff dff_A_lmYTnB6T2_0(.dout(w_G150_3[0]),.din(w_dff_A_lmYTnB6T2_0),.clk(gclk));
	jdff dff_A_rvbd5L818_0(.dout(w_dff_A_lmYTnB6T2_0),.din(w_dff_A_rvbd5L818_0),.clk(gclk));
	jdff dff_A_G446uEg82_0(.dout(w_dff_A_rvbd5L818_0),.din(w_dff_A_G446uEg82_0),.clk(gclk));
	jdff dff_A_o1fgSDMH9_0(.dout(w_G150_0[0]),.din(w_dff_A_o1fgSDMH9_0),.clk(gclk));
	jdff dff_A_arW3GOKm9_0(.dout(w_dff_A_o1fgSDMH9_0),.din(w_dff_A_arW3GOKm9_0),.clk(gclk));
	jdff dff_A_7JjrxqHK3_0(.dout(w_dff_A_arW3GOKm9_0),.din(w_dff_A_7JjrxqHK3_0),.clk(gclk));
	jdff dff_A_NecxCShL5_1(.dout(w_G150_0[1]),.din(w_dff_A_NecxCShL5_1),.clk(gclk));
	jdff dff_A_qn3EYT6o2_1(.dout(w_dff_A_NecxCShL5_1),.din(w_dff_A_qn3EYT6o2_1),.clk(gclk));
	jdff dff_A_3O7aE85M4_1(.dout(w_dff_A_qn3EYT6o2_1),.din(w_dff_A_3O7aE85M4_1),.clk(gclk));
	jdff dff_A_odEjqQBT9_0(.dout(w_G58_3[0]),.din(w_dff_A_odEjqQBT9_0),.clk(gclk));
	jdff dff_A_tbzMfHWv2_1(.dout(w_G58_3[1]),.din(w_dff_A_tbzMfHWv2_1),.clk(gclk));
	jdff dff_A_Y8KSfdHb2_1(.dout(w_n622_0[1]),.din(w_dff_A_Y8KSfdHb2_1),.clk(gclk));
	jdff dff_A_DU6dpN675_1(.dout(w_n615_0[1]),.din(w_dff_A_DU6dpN675_1),.clk(gclk));
	jdff dff_A_LYezivm14_1(.dout(w_G200_2[1]),.din(w_dff_A_LYezivm14_1),.clk(gclk));
	jdff dff_A_6fc83rfr5_1(.dout(w_dff_A_LYezivm14_1),.din(w_dff_A_6fc83rfr5_1),.clk(gclk));
	jdff dff_A_DvtEd7gf6_1(.dout(w_dff_A_6fc83rfr5_1),.din(w_dff_A_DvtEd7gf6_1),.clk(gclk));
	jdff dff_A_OZ9A1o2l5_1(.dout(w_dff_A_DvtEd7gf6_1),.din(w_dff_A_OZ9A1o2l5_1),.clk(gclk));
	jdff dff_A_gPvOOn0B3_2(.dout(w_G200_2[2]),.din(w_dff_A_gPvOOn0B3_2),.clk(gclk));
	jdff dff_A_DvFUx4YH1_2(.dout(w_dff_A_gPvOOn0B3_2),.din(w_dff_A_DvFUx4YH1_2),.clk(gclk));
	jdff dff_A_pB0AHT919_2(.dout(w_dff_A_DvFUx4YH1_2),.din(w_dff_A_pB0AHT919_2),.clk(gclk));
	jdff dff_A_fGxofY8k0_2(.dout(w_dff_A_pB0AHT919_2),.din(w_dff_A_fGxofY8k0_2),.clk(gclk));
	jdff dff_A_8XGHsvdi4_0(.dout(w_n407_1[0]),.din(w_dff_A_8XGHsvdi4_0),.clk(gclk));
	jdff dff_A_bKzLMaed4_1(.dout(w_n407_1[1]),.din(w_dff_A_bKzLMaed4_1),.clk(gclk));
	jdff dff_A_dSGJppjg1_1(.dout(w_dff_A_bKzLMaed4_1),.din(w_dff_A_dSGJppjg1_1),.clk(gclk));
	jdff dff_B_mc5XNW0i3_3(.din(G132),.dout(w_dff_B_mc5XNW0i3_3),.clk(gclk));
	jdff dff_B_p5r3z6Ka3_3(.din(w_dff_B_mc5XNW0i3_3),.dout(w_dff_B_p5r3z6Ka3_3),.clk(gclk));
	jdff dff_B_YQvH26gl2_3(.din(w_dff_B_p5r3z6Ka3_3),.dout(w_dff_B_YQvH26gl2_3),.clk(gclk));
	jdff dff_A_gRoTD7iz4_0(.dout(w_n612_3[0]),.din(w_dff_A_gRoTD7iz4_0),.clk(gclk));
	jdff dff_A_fuzE1ysw1_0(.dout(w_dff_A_gRoTD7iz4_0),.din(w_dff_A_fuzE1ysw1_0),.clk(gclk));
	jdff dff_A_3d4Cb9cl2_0(.dout(w_dff_A_fuzE1ysw1_0),.din(w_dff_A_3d4Cb9cl2_0),.clk(gclk));
	jdff dff_A_5MLe7set8_0(.dout(w_dff_A_3d4Cb9cl2_0),.din(w_dff_A_5MLe7set8_0),.clk(gclk));
	jdff dff_A_hVtkSxNU2_0(.dout(w_dff_A_5MLe7set8_0),.din(w_dff_A_hVtkSxNU2_0),.clk(gclk));
	jdff dff_A_JWLUa8kc1_0(.dout(w_dff_A_hVtkSxNU2_0),.din(w_dff_A_JWLUa8kc1_0),.clk(gclk));
	jdff dff_A_yT7VtqIj3_0(.dout(w_dff_A_JWLUa8kc1_0),.din(w_dff_A_yT7VtqIj3_0),.clk(gclk));
	jdff dff_A_XgI3rQ976_0(.dout(w_dff_A_yT7VtqIj3_0),.din(w_dff_A_XgI3rQ976_0),.clk(gclk));
	jdff dff_A_c3PGxlbs7_2(.dout(w_n612_3[2]),.din(w_dff_A_c3PGxlbs7_2),.clk(gclk));
	jdff dff_A_XPAo245d2_2(.dout(w_dff_A_c3PGxlbs7_2),.din(w_dff_A_XPAo245d2_2),.clk(gclk));
	jdff dff_A_RmERhBON2_2(.dout(w_dff_A_XPAo245d2_2),.din(w_dff_A_RmERhBON2_2),.clk(gclk));
	jdff dff_A_UvJVFXnw5_2(.dout(w_dff_A_RmERhBON2_2),.din(w_dff_A_UvJVFXnw5_2),.clk(gclk));
	jdff dff_A_SM7ZPe7K2_2(.dout(w_dff_A_UvJVFXnw5_2),.din(w_dff_A_SM7ZPe7K2_2),.clk(gclk));
	jdff dff_A_7pMbHm3V3_2(.dout(w_dff_A_SM7ZPe7K2_2),.din(w_dff_A_7pMbHm3V3_2),.clk(gclk));
	jdff dff_A_X3wMX2hI4_2(.dout(w_dff_A_7pMbHm3V3_2),.din(w_dff_A_X3wMX2hI4_2),.clk(gclk));
	jdff dff_A_tcO6s0D57_2(.dout(w_dff_A_X3wMX2hI4_2),.din(w_dff_A_tcO6s0D57_2),.clk(gclk));
	jdff dff_A_d3EBu8i75_1(.dout(w_n612_0[1]),.din(w_dff_A_d3EBu8i75_1),.clk(gclk));
	jdff dff_A_ceDSiX433_1(.dout(w_dff_A_d3EBu8i75_1),.din(w_dff_A_ceDSiX433_1),.clk(gclk));
	jdff dff_A_Wj35XI293_1(.dout(w_dff_A_ceDSiX433_1),.din(w_dff_A_Wj35XI293_1),.clk(gclk));
	jdff dff_A_NQgcz3gX4_1(.dout(w_dff_A_Wj35XI293_1),.din(w_dff_A_NQgcz3gX4_1),.clk(gclk));
	jdff dff_A_seuHrhMy5_2(.dout(w_n612_0[2]),.din(w_dff_A_seuHrhMy5_2),.clk(gclk));
	jdff dff_A_nuaJKMkK5_1(.dout(w_n146_1[1]),.din(w_dff_A_nuaJKMkK5_1),.clk(gclk));
	jdff dff_A_MGRcmzfo9_1(.dout(w_dff_A_nuaJKMkK5_1),.din(w_dff_A_MGRcmzfo9_1),.clk(gclk));
	jdff dff_A_lqWvE3r74_1(.dout(w_dff_A_MGRcmzfo9_1),.din(w_dff_A_lqWvE3r74_1),.clk(gclk));
	jdff dff_A_iuagizU15_2(.dout(w_n146_1[2]),.din(w_dff_A_iuagizU15_2),.clk(gclk));
	jdff dff_A_UOXfvX1p2_2(.dout(w_dff_A_iuagizU15_2),.din(w_dff_A_UOXfvX1p2_2),.clk(gclk));
	jdff dff_A_5HJK33pc5_2(.dout(w_dff_A_UOXfvX1p2_2),.din(w_dff_A_5HJK33pc5_2),.clk(gclk));
	jdff dff_A_B8iF0AOI6_0(.dout(w_n425_1[0]),.din(w_dff_A_B8iF0AOI6_0),.clk(gclk));
	jdff dff_A_EXPJgVUo8_0(.dout(w_dff_A_B8iF0AOI6_0),.din(w_dff_A_EXPJgVUo8_0),.clk(gclk));
	jdff dff_A_hVTreHXn7_0(.dout(w_dff_A_EXPJgVUo8_0),.din(w_dff_A_hVTreHXn7_0),.clk(gclk));
	jdff dff_A_MosWL2Xc7_0(.dout(w_dff_A_hVTreHXn7_0),.din(w_dff_A_MosWL2Xc7_0),.clk(gclk));
	jdff dff_A_6hzNH7Wq9_0(.dout(w_dff_A_MosWL2Xc7_0),.din(w_dff_A_6hzNH7Wq9_0),.clk(gclk));
	jdff dff_A_kSHJvLUk9_0(.dout(w_dff_A_6hzNH7Wq9_0),.din(w_dff_A_kSHJvLUk9_0),.clk(gclk));
	jdff dff_A_XvKL8ZfZ2_0(.dout(w_dff_A_kSHJvLUk9_0),.din(w_dff_A_XvKL8ZfZ2_0),.clk(gclk));
	jdff dff_A_9denz4cd7_0(.dout(w_dff_A_XvKL8ZfZ2_0),.din(w_dff_A_9denz4cd7_0),.clk(gclk));
	jdff dff_A_4lLPtiA58_0(.dout(w_dff_A_9denz4cd7_0),.din(w_dff_A_4lLPtiA58_0),.clk(gclk));
	jdff dff_A_oB09sLbt1_0(.dout(w_dff_A_4lLPtiA58_0),.din(w_dff_A_oB09sLbt1_0),.clk(gclk));
	jdff dff_A_RaQ0g0xZ2_1(.dout(w_n425_1[1]),.din(w_dff_A_RaQ0g0xZ2_1),.clk(gclk));
	jdff dff_A_ITfKXpn52_1(.dout(w_dff_A_RaQ0g0xZ2_1),.din(w_dff_A_ITfKXpn52_1),.clk(gclk));
	jdff dff_A_UOpVM55s0_1(.dout(w_dff_A_ITfKXpn52_1),.din(w_dff_A_UOpVM55s0_1),.clk(gclk));
	jdff dff_A_gOcQMJAL3_1(.dout(w_dff_A_UOpVM55s0_1),.din(w_dff_A_gOcQMJAL3_1),.clk(gclk));
	jdff dff_A_XEUCRZjE9_1(.dout(w_dff_A_gOcQMJAL3_1),.din(w_dff_A_XEUCRZjE9_1),.clk(gclk));
	jdff dff_A_8bgwqSiU6_1(.dout(w_dff_A_XEUCRZjE9_1),.din(w_dff_A_8bgwqSiU6_1),.clk(gclk));
	jdff dff_A_tc432UJX6_1(.dout(w_dff_A_8bgwqSiU6_1),.din(w_dff_A_tc432UJX6_1),.clk(gclk));
	jdff dff_A_9eOwMtlQ2_1(.dout(w_dff_A_tc432UJX6_1),.din(w_dff_A_9eOwMtlQ2_1),.clk(gclk));
	jdff dff_A_tIIMMgaG3_1(.dout(w_dff_A_9eOwMtlQ2_1),.din(w_dff_A_tIIMMgaG3_1),.clk(gclk));
	jdff dff_A_3Nq7jofV2_1(.dout(w_n425_0[1]),.din(w_dff_A_3Nq7jofV2_1),.clk(gclk));
	jdff dff_A_vvGvnuOX4_1(.dout(w_dff_A_3Nq7jofV2_1),.din(w_dff_A_vvGvnuOX4_1),.clk(gclk));
	jdff dff_A_ohqUtohD0_1(.dout(w_dff_A_vvGvnuOX4_1),.din(w_dff_A_ohqUtohD0_1),.clk(gclk));
	jdff dff_A_iXigC0zp9_1(.dout(w_dff_A_ohqUtohD0_1),.din(w_dff_A_iXigC0zp9_1),.clk(gclk));
	jdff dff_A_OYlcoSK01_1(.dout(w_dff_A_iXigC0zp9_1),.din(w_dff_A_OYlcoSK01_1),.clk(gclk));
	jdff dff_A_gEXTiP6o9_1(.dout(w_dff_A_OYlcoSK01_1),.din(w_dff_A_gEXTiP6o9_1),.clk(gclk));
	jdff dff_A_Tl9ag5Oa2_1(.dout(w_dff_A_gEXTiP6o9_1),.din(w_dff_A_Tl9ag5Oa2_1),.clk(gclk));
	jdff dff_A_dtYZgtNk1_1(.dout(w_dff_A_Tl9ag5Oa2_1),.din(w_dff_A_dtYZgtNk1_1),.clk(gclk));
	jdff dff_A_0wOEUyzd3_1(.dout(w_dff_A_dtYZgtNk1_1),.din(w_dff_A_0wOEUyzd3_1),.clk(gclk));
	jdff dff_A_JyqdRTrX8_2(.dout(w_n425_0[2]),.din(w_dff_A_JyqdRTrX8_2),.clk(gclk));
	jdff dff_A_DojwvyJK9_2(.dout(w_dff_A_JyqdRTrX8_2),.din(w_dff_A_DojwvyJK9_2),.clk(gclk));
	jdff dff_A_67hGSlyt0_2(.dout(w_dff_A_DojwvyJK9_2),.din(w_dff_A_67hGSlyt0_2),.clk(gclk));
	jdff dff_A_dEjDbPbD9_2(.dout(w_dff_A_67hGSlyt0_2),.din(w_dff_A_dEjDbPbD9_2),.clk(gclk));
	jdff dff_A_oBRutj0d7_2(.dout(w_dff_A_dEjDbPbD9_2),.din(w_dff_A_oBRutj0d7_2),.clk(gclk));
	jdff dff_A_E18gzmfh6_2(.dout(w_dff_A_oBRutj0d7_2),.din(w_dff_A_E18gzmfh6_2),.clk(gclk));
	jdff dff_A_nS6ihTCi8_2(.dout(w_dff_A_E18gzmfh6_2),.din(w_dff_A_nS6ihTCi8_2),.clk(gclk));
	jdff dff_A_AQJ35VO30_2(.dout(w_dff_A_nS6ihTCi8_2),.din(w_dff_A_AQJ35VO30_2),.clk(gclk));
	jdff dff_A_YTQDqmI01_2(.dout(w_dff_A_AQJ35VO30_2),.din(w_dff_A_YTQDqmI01_2),.clk(gclk));
	jdff dff_A_GSDAVnE79_2(.dout(w_dff_A_YTQDqmI01_2),.din(w_dff_A_GSDAVnE79_2),.clk(gclk));
	jdff dff_A_aaUwg8TN3_2(.dout(w_dff_A_GSDAVnE79_2),.din(w_dff_A_aaUwg8TN3_2),.clk(gclk));
	jdff dff_A_Q4uINlbI6_0(.dout(w_n148_1[0]),.din(w_dff_A_Q4uINlbI6_0),.clk(gclk));
	jdff dff_A_LLkLYzzG5_0(.dout(w_dff_A_Q4uINlbI6_0),.din(w_dff_A_LLkLYzzG5_0),.clk(gclk));
	jdff dff_A_jULG3NAn2_0(.dout(w_dff_A_LLkLYzzG5_0),.din(w_dff_A_jULG3NAn2_0),.clk(gclk));
	jdff dff_A_gMO5Afgd7_1(.dout(w_n148_1[1]),.din(w_dff_A_gMO5Afgd7_1),.clk(gclk));
	jdff dff_A_DMtX3I347_1(.dout(w_dff_A_gMO5Afgd7_1),.din(w_dff_A_DMtX3I347_1),.clk(gclk));
	jdff dff_B_8Fgn1vPH7_0(.din(n701),.dout(w_dff_B_8Fgn1vPH7_0),.clk(gclk));
	jdff dff_B_JiVUAAap8_0(.din(w_dff_B_8Fgn1vPH7_0),.dout(w_dff_B_JiVUAAap8_0),.clk(gclk));
	jdff dff_A_ZhSqkV059_0(.dout(w_n604_1[0]),.din(w_dff_A_ZhSqkV059_0),.clk(gclk));
	jdff dff_A_6ULOEFua4_0(.dout(w_dff_A_ZhSqkV059_0),.din(w_dff_A_6ULOEFua4_0),.clk(gclk));
	jdff dff_A_kLIzZhGG6_2(.dout(w_n604_1[2]),.din(w_dff_A_kLIzZhGG6_2),.clk(gclk));
	jdff dff_A_AWmVjZRn3_2(.dout(w_dff_A_kLIzZhGG6_2),.din(w_dff_A_AWmVjZRn3_2),.clk(gclk));
	jdff dff_A_Afyz80ea3_2(.dout(w_dff_A_AWmVjZRn3_2),.din(w_dff_A_Afyz80ea3_2),.clk(gclk));
	jdff dff_A_2E3IIK0F1_2(.dout(w_dff_A_Afyz80ea3_2),.din(w_dff_A_2E3IIK0F1_2),.clk(gclk));
	jdff dff_A_KGHKFH5d7_2(.dout(w_dff_A_2E3IIK0F1_2),.din(w_dff_A_KGHKFH5d7_2),.clk(gclk));
	jdff dff_A_AY9jNJeF9_2(.dout(w_dff_A_KGHKFH5d7_2),.din(w_dff_A_AY9jNJeF9_2),.clk(gclk));
	jdff dff_A_eMkn6guf5_2(.dout(w_dff_A_AY9jNJeF9_2),.din(w_dff_A_eMkn6guf5_2),.clk(gclk));
	jdff dff_A_dLX1RnmY5_0(.dout(w_n603_2[0]),.din(w_dff_A_dLX1RnmY5_0),.clk(gclk));
	jdff dff_A_OWnSuGej0_0(.dout(w_dff_A_dLX1RnmY5_0),.din(w_dff_A_OWnSuGej0_0),.clk(gclk));
	jdff dff_A_WWHFDgjM6_0(.dout(w_dff_A_OWnSuGej0_0),.din(w_dff_A_WWHFDgjM6_0),.clk(gclk));
	jdff dff_A_C4dNcQlP8_0(.dout(w_dff_A_WWHFDgjM6_0),.din(w_dff_A_C4dNcQlP8_0),.clk(gclk));
	jdff dff_A_y12OfxT53_0(.dout(w_dff_A_C4dNcQlP8_0),.din(w_dff_A_y12OfxT53_0),.clk(gclk));
	jdff dff_A_FYYhgysf1_0(.dout(w_dff_A_y12OfxT53_0),.din(w_dff_A_FYYhgysf1_0),.clk(gclk));
	jdff dff_A_g1RxLjhU4_0(.dout(w_n603_0[0]),.din(w_dff_A_g1RxLjhU4_0),.clk(gclk));
	jdff dff_A_KaDu34l84_0(.dout(w_dff_A_g1RxLjhU4_0),.din(w_dff_A_KaDu34l84_0),.clk(gclk));
	jdff dff_A_psX1F1CX9_0(.dout(w_dff_A_KaDu34l84_0),.din(w_dff_A_psX1F1CX9_0),.clk(gclk));
	jdff dff_A_XuQLkVNX5_0(.dout(w_dff_A_psX1F1CX9_0),.din(w_dff_A_XuQLkVNX5_0),.clk(gclk));
	jdff dff_A_RKaGtSos7_0(.dout(w_dff_A_XuQLkVNX5_0),.din(w_dff_A_RKaGtSos7_0),.clk(gclk));
	jdff dff_A_k3fbjoaD1_0(.dout(w_dff_A_RKaGtSos7_0),.din(w_dff_A_k3fbjoaD1_0),.clk(gclk));
	jdff dff_A_xQzqKOOf3_0(.dout(w_dff_A_k3fbjoaD1_0),.din(w_dff_A_xQzqKOOf3_0),.clk(gclk));
	jdff dff_A_99KqSkib8_0(.dout(w_dff_A_xQzqKOOf3_0),.din(w_dff_A_99KqSkib8_0),.clk(gclk));
	jdff dff_A_qQ98sBdi6_2(.dout(w_n603_0[2]),.din(w_dff_A_qQ98sBdi6_2),.clk(gclk));
	jdff dff_A_W8fROgog4_2(.dout(w_dff_A_qQ98sBdi6_2),.din(w_dff_A_W8fROgog4_2),.clk(gclk));
	jdff dff_A_g62GXDFM2_2(.dout(w_dff_A_W8fROgog4_2),.din(w_dff_A_g62GXDFM2_2),.clk(gclk));
	jdff dff_A_1QtS2Hu31_2(.dout(w_dff_A_g62GXDFM2_2),.din(w_dff_A_1QtS2Hu31_2),.clk(gclk));
	jdff dff_A_evb7rlOY0_2(.dout(w_dff_A_1QtS2Hu31_2),.din(w_dff_A_evb7rlOY0_2),.clk(gclk));
	jdff dff_A_qjpiyGia4_2(.dout(w_dff_A_evb7rlOY0_2),.din(w_dff_A_qjpiyGia4_2),.clk(gclk));
	jdff dff_A_fOTowXgS5_2(.dout(w_dff_A_qjpiyGia4_2),.din(w_dff_A_fOTowXgS5_2),.clk(gclk));
	jdff dff_A_xlz6eex52_2(.dout(w_dff_A_fOTowXgS5_2),.din(w_dff_A_xlz6eex52_2),.clk(gclk));
	jdff dff_A_qo6zb8tr9_2(.dout(w_dff_A_xlz6eex52_2),.din(w_dff_A_qo6zb8tr9_2),.clk(gclk));
	jdff dff_A_fx8vizA06_2(.dout(w_dff_A_qo6zb8tr9_2),.din(w_dff_A_fx8vizA06_2),.clk(gclk));
	jdff dff_B_ZJlqJ5FK5_3(.din(n603),.dout(w_dff_B_ZJlqJ5FK5_3),.clk(gclk));
	jdff dff_A_T2KnlB2j0_0(.dout(w_n602_0[0]),.din(w_dff_A_T2KnlB2j0_0),.clk(gclk));
	jdff dff_A_oWD7Fbko3_0(.dout(w_dff_A_T2KnlB2j0_0),.din(w_dff_A_oWD7Fbko3_0),.clk(gclk));
	jdff dff_A_jJo4eJM59_0(.dout(w_dff_A_oWD7Fbko3_0),.din(w_dff_A_jJo4eJM59_0),.clk(gclk));
	jdff dff_A_8U1wUBmo4_0(.dout(w_dff_A_jJo4eJM59_0),.din(w_dff_A_8U1wUBmo4_0),.clk(gclk));
	jdff dff_A_jOSOqfwz8_0(.dout(w_dff_A_8U1wUBmo4_0),.din(w_dff_A_jOSOqfwz8_0),.clk(gclk));
	jdff dff_A_AWYJwKgI1_0(.dout(w_dff_A_jOSOqfwz8_0),.din(w_dff_A_AWYJwKgI1_0),.clk(gclk));
	jdff dff_A_TSmGjlnZ7_0(.dout(w_dff_A_AWYJwKgI1_0),.din(w_dff_A_TSmGjlnZ7_0),.clk(gclk));
	jdff dff_A_yrkL9nfY4_0(.dout(w_dff_A_TSmGjlnZ7_0),.din(w_dff_A_yrkL9nfY4_0),.clk(gclk));
	jdff dff_A_enbsVRWP4_0(.dout(w_dff_A_yrkL9nfY4_0),.din(w_dff_A_enbsVRWP4_0),.clk(gclk));
	jdff dff_A_ouEGlPzD1_0(.dout(w_dff_A_enbsVRWP4_0),.din(w_dff_A_ouEGlPzD1_0),.clk(gclk));
	jdff dff_A_uP2pN1Iw3_0(.dout(w_dff_A_ouEGlPzD1_0),.din(w_dff_A_uP2pN1Iw3_0),.clk(gclk));
	jdff dff_A_BbfphW8d0_0(.dout(w_dff_A_uP2pN1Iw3_0),.din(w_dff_A_BbfphW8d0_0),.clk(gclk));
	jdff dff_A_mYqX3KMD9_0(.dout(w_dff_A_BbfphW8d0_0),.din(w_dff_A_mYqX3KMD9_0),.clk(gclk));
	jdff dff_A_k48sJ4dU4_0(.dout(w_n592_0[0]),.din(w_dff_A_k48sJ4dU4_0),.clk(gclk));
	jdff dff_A_0tAfQwI36_0(.dout(w_dff_A_k48sJ4dU4_0),.din(w_dff_A_0tAfQwI36_0),.clk(gclk));
	jdff dff_A_qAo7eWBD2_0(.dout(w_dff_A_0tAfQwI36_0),.din(w_dff_A_qAo7eWBD2_0),.clk(gclk));
	jdff dff_A_lh9QJT3N1_0(.dout(w_dff_A_qAo7eWBD2_0),.din(w_dff_A_lh9QJT3N1_0),.clk(gclk));
	jdff dff_A_2D7mIetl1_0(.dout(w_dff_A_lh9QJT3N1_0),.din(w_dff_A_2D7mIetl1_0),.clk(gclk));
	jdff dff_A_Cb3BKH502_0(.dout(w_dff_A_2D7mIetl1_0),.din(w_dff_A_Cb3BKH502_0),.clk(gclk));
	jdff dff_A_sWvLeDdt9_0(.dout(w_dff_A_Cb3BKH502_0),.din(w_dff_A_sWvLeDdt9_0),.clk(gclk));
	jdff dff_A_Dx84Df5y9_0(.dout(w_dff_A_sWvLeDdt9_0),.din(w_dff_A_Dx84Df5y9_0),.clk(gclk));
	jdff dff_A_gdygnVVT6_0(.dout(w_dff_A_Dx84Df5y9_0),.din(w_dff_A_gdygnVVT6_0),.clk(gclk));
	jdff dff_A_hZGV57du9_2(.dout(w_n592_0[2]),.din(w_dff_A_hZGV57du9_2),.clk(gclk));
	jdff dff_A_zZlJKFXg8_2(.dout(w_dff_A_hZGV57du9_2),.din(w_dff_A_zZlJKFXg8_2),.clk(gclk));
	jdff dff_A_JcRZ1cNk5_2(.dout(w_dff_A_zZlJKFXg8_2),.din(w_dff_A_JcRZ1cNk5_2),.clk(gclk));
	jdff dff_A_7aY8PRMZ7_2(.dout(w_dff_A_JcRZ1cNk5_2),.din(w_dff_A_7aY8PRMZ7_2),.clk(gclk));
	jdff dff_A_T6m0G33s8_2(.dout(w_dff_A_7aY8PRMZ7_2),.din(w_dff_A_T6m0G33s8_2),.clk(gclk));
	jdff dff_A_TvD462gv0_2(.dout(w_dff_A_T6m0G33s8_2),.din(w_dff_A_TvD462gv0_2),.clk(gclk));
	jdff dff_A_N8DzoCir9_2(.dout(w_dff_A_TvD462gv0_2),.din(w_dff_A_N8DzoCir9_2),.clk(gclk));
	jdff dff_A_knLSeDn77_2(.dout(w_dff_A_N8DzoCir9_2),.din(w_dff_A_knLSeDn77_2),.clk(gclk));
	jdff dff_A_uxs6nHfu0_2(.dout(w_dff_A_knLSeDn77_2),.din(w_dff_A_uxs6nHfu0_2),.clk(gclk));
	jdff dff_A_qkiXRVFc3_2(.dout(w_dff_A_uxs6nHfu0_2),.din(w_dff_A_qkiXRVFc3_2),.clk(gclk));
	jdff dff_A_3eXUnVcQ9_2(.dout(w_dff_A_qkiXRVFc3_2),.din(w_dff_A_3eXUnVcQ9_2),.clk(gclk));
	jdff dff_A_kcce7wmu0_2(.dout(w_dff_A_3eXUnVcQ9_2),.din(w_dff_A_kcce7wmu0_2),.clk(gclk));
	jdff dff_A_mLrwQRJ09_1(.dout(w_n591_0[1]),.din(w_dff_A_mLrwQRJ09_1),.clk(gclk));
	jdff dff_A_n5CXs36m9_1(.dout(w_dff_A_mLrwQRJ09_1),.din(w_dff_A_n5CXs36m9_1),.clk(gclk));
	jdff dff_A_pnnxiLey6_1(.dout(w_dff_A_n5CXs36m9_1),.din(w_dff_A_pnnxiLey6_1),.clk(gclk));
	jdff dff_A_l1y7ttSN8_1(.dout(w_dff_A_pnnxiLey6_1),.din(w_dff_A_l1y7ttSN8_1),.clk(gclk));
	jdff dff_A_ue9GOMuM9_1(.dout(w_dff_A_l1y7ttSN8_1),.din(w_dff_A_ue9GOMuM9_1),.clk(gclk));
	jdff dff_A_BaZBveCO0_1(.dout(w_dff_A_ue9GOMuM9_1),.din(w_dff_A_BaZBveCO0_1),.clk(gclk));
	jdff dff_A_CYmuDsfL2_1(.dout(w_dff_A_BaZBveCO0_1),.din(w_dff_A_CYmuDsfL2_1),.clk(gclk));
	jdff dff_A_egzqFENt9_1(.dout(w_dff_A_CYmuDsfL2_1),.din(w_dff_A_egzqFENt9_1),.clk(gclk));
	jdff dff_A_VXkfY5sT6_1(.dout(w_dff_A_egzqFENt9_1),.din(w_dff_A_VXkfY5sT6_1),.clk(gclk));
	jdff dff_A_yHY3JlNx6_1(.dout(w_dff_A_VXkfY5sT6_1),.din(w_dff_A_yHY3JlNx6_1),.clk(gclk));
	jdff dff_A_DHUjSQ1X3_1(.dout(w_dff_A_yHY3JlNx6_1),.din(w_dff_A_DHUjSQ1X3_1),.clk(gclk));
	jdff dff_A_N4EYChmd7_2(.dout(w_n591_0[2]),.din(w_dff_A_N4EYChmd7_2),.clk(gclk));
	jdff dff_A_UrMqEtit8_2(.dout(w_dff_A_N4EYChmd7_2),.din(w_dff_A_UrMqEtit8_2),.clk(gclk));
	jdff dff_A_DdkSMVhT9_2(.dout(w_dff_A_UrMqEtit8_2),.din(w_dff_A_DdkSMVhT9_2),.clk(gclk));
	jdff dff_A_ufzJQTfW8_2(.dout(w_dff_A_DdkSMVhT9_2),.din(w_dff_A_ufzJQTfW8_2),.clk(gclk));
	jdff dff_A_aKrx2RoP6_2(.dout(w_dff_A_ufzJQTfW8_2),.din(w_dff_A_aKrx2RoP6_2),.clk(gclk));
	jdff dff_A_hqp1s0XK0_2(.dout(w_dff_A_aKrx2RoP6_2),.din(w_dff_A_hqp1s0XK0_2),.clk(gclk));
	jdff dff_A_ThhlVpCb8_2(.dout(w_dff_A_hqp1s0XK0_2),.din(w_dff_A_ThhlVpCb8_2),.clk(gclk));
	jdff dff_A_8dOLieCe3_2(.dout(w_dff_A_ThhlVpCb8_2),.din(w_dff_A_8dOLieCe3_2),.clk(gclk));
	jdff dff_A_lVqvmdGJ6_2(.dout(w_dff_A_8dOLieCe3_2),.din(w_dff_A_lVqvmdGJ6_2),.clk(gclk));
	jdff dff_A_we57jcH39_2(.dout(w_dff_A_lVqvmdGJ6_2),.din(w_dff_A_we57jcH39_2),.clk(gclk));
	jdff dff_A_A4hFy3VS9_2(.dout(w_dff_A_we57jcH39_2),.din(w_dff_A_A4hFy3VS9_2),.clk(gclk));
	jdff dff_B_lVDmVpR90_1(.din(n690),.dout(w_dff_B_lVDmVpR90_1),.clk(gclk));
	jdff dff_A_FjTBNcjL8_0(.dout(w_n696_1[0]),.din(w_dff_A_FjTBNcjL8_0),.clk(gclk));
	jdff dff_A_9ralKSB82_0(.dout(w_dff_A_FjTBNcjL8_0),.din(w_dff_A_9ralKSB82_0),.clk(gclk));
	jdff dff_A_JALV2n893_2(.dout(w_n696_1[2]),.din(w_dff_A_JALV2n893_2),.clk(gclk));
	jdff dff_A_zYqiFtf66_2(.dout(w_dff_A_JALV2n893_2),.din(w_dff_A_zYqiFtf66_2),.clk(gclk));
	jdff dff_A_G8ZFd4Pm3_1(.dout(w_n696_0[1]),.din(w_dff_A_G8ZFd4Pm3_1),.clk(gclk));
	jdff dff_A_Osu92vvW7_1(.dout(w_dff_A_G8ZFd4Pm3_1),.din(w_dff_A_Osu92vvW7_1),.clk(gclk));
	jdff dff_B_Vkewf4pA1_0(.din(n695),.dout(w_dff_B_Vkewf4pA1_0),.clk(gclk));
	jdff dff_A_tibR6DAP5_1(.dout(w_n692_0[1]),.din(w_dff_A_tibR6DAP5_1),.clk(gclk));
	jdff dff_B_1kLZs6DX8_2(.din(n692),.dout(w_dff_B_1kLZs6DX8_2),.clk(gclk));
	jdff dff_B_cGtmdP1h3_2(.din(w_dff_B_1kLZs6DX8_2),.dout(w_dff_B_cGtmdP1h3_2),.clk(gclk));
	jdff dff_B_eElI0crC8_2(.din(w_dff_B_cGtmdP1h3_2),.dout(w_dff_B_eElI0crC8_2),.clk(gclk));
	jdff dff_B_qDaUGw3r8_0(.din(n411),.dout(w_dff_B_qDaUGw3r8_0),.clk(gclk));
	jdff dff_B_DYgSAR3B4_0(.din(w_dff_B_qDaUGw3r8_0),.dout(w_dff_B_DYgSAR3B4_0),.clk(gclk));
	jdff dff_B_218vRI5f9_0(.din(w_dff_B_DYgSAR3B4_0),.dout(w_dff_B_218vRI5f9_0),.clk(gclk));
	jdff dff_A_dSJwJBTY2_1(.dout(w_n407_0[1]),.din(w_dff_A_dSJwJBTY2_1),.clk(gclk));
	jdff dff_A_qkw04i6F0_1(.dout(w_dff_A_dSJwJBTY2_1),.din(w_dff_A_qkw04i6F0_1),.clk(gclk));
	jdff dff_A_J25dw3vL9_1(.dout(w_dff_A_qkw04i6F0_1),.din(w_dff_A_J25dw3vL9_1),.clk(gclk));
	jdff dff_A_MCUi8aXw4_2(.dout(w_n407_0[2]),.din(w_dff_A_MCUi8aXw4_2),.clk(gclk));
	jdff dff_B_Sph0DQDc9_0(.din(n403),.dout(w_dff_B_Sph0DQDc9_0),.clk(gclk));
	jdff dff_A_cSstGaA84_1(.dout(w_n401_0[1]),.din(w_dff_A_cSstGaA84_1),.clk(gclk));
	jdff dff_B_i1l3Mp175_0(.din(n398),.dout(w_dff_B_i1l3Mp175_0),.clk(gclk));
	jdff dff_A_y6gSzsOt4_1(.dout(w_n72_0[1]),.din(w_dff_A_y6gSzsOt4_1),.clk(gclk));
	jdff dff_A_7G2esgGD7_1(.dout(w_dff_A_y6gSzsOt4_1),.din(w_dff_A_7G2esgGD7_1),.clk(gclk));
	jdff dff_A_KNB7jK4F8_1(.dout(w_dff_A_7G2esgGD7_1),.din(w_dff_A_KNB7jK4F8_1),.clk(gclk));
	jdff dff_A_PnyFohuo6_2(.dout(w_n72_0[2]),.din(w_dff_A_PnyFohuo6_2),.clk(gclk));
	jdff dff_A_bUhcjxrq5_2(.dout(w_dff_A_PnyFohuo6_2),.din(w_dff_A_bUhcjxrq5_2),.clk(gclk));
	jdff dff_B_D9Bk1MgI6_1(.din(n393),.dout(w_dff_B_D9Bk1MgI6_1),.clk(gclk));
	jdff dff_B_vEpVHQhZ6_0(.din(n394),.dout(w_dff_B_vEpVHQhZ6_0),.clk(gclk));
	jdff dff_A_kIrJMqOC9_0(.dout(w_n112_3[0]),.din(w_dff_A_kIrJMqOC9_0),.clk(gclk));
	jdff dff_A_IlnhALf97_0(.dout(w_dff_A_kIrJMqOC9_0),.din(w_dff_A_IlnhALf97_0),.clk(gclk));
	jdff dff_A_CgQNpzjX4_1(.dout(w_n112_3[1]),.din(w_dff_A_CgQNpzjX4_1),.clk(gclk));
	jdff dff_A_XNG8O2VN2_1(.dout(w_G58_4[1]),.din(w_dff_A_XNG8O2VN2_1),.clk(gclk));
	jdff dff_A_oirhwcSF6_0(.dout(w_G58_1[0]),.din(w_dff_A_oirhwcSF6_0),.clk(gclk));
	jdff dff_A_cFfobJ8r5_2(.dout(w_G58_1[2]),.din(w_dff_A_cFfobJ8r5_2),.clk(gclk));
	jdff dff_A_kv1ybzLQ2_2(.dout(w_dff_A_cFfobJ8r5_2),.din(w_dff_A_kv1ybzLQ2_2),.clk(gclk));
	jdff dff_A_CIvU00uO4_2(.dout(w_dff_A_kv1ybzLQ2_2),.din(w_dff_A_CIvU00uO4_2),.clk(gclk));
	jdff dff_A_K12y90Dv4_2(.dout(w_dff_A_CIvU00uO4_2),.din(w_dff_A_K12y90Dv4_2),.clk(gclk));
	jdff dff_A_Jefdi59f3_1(.dout(w_G58_0[1]),.din(w_dff_A_Jefdi59f3_1),.clk(gclk));
	jdff dff_A_q9GcptK94_2(.dout(w_G58_0[2]),.din(w_dff_A_q9GcptK94_2),.clk(gclk));
	jdff dff_A_vbKRF6U80_2(.dout(w_dff_A_q9GcptK94_2),.din(w_dff_A_vbKRF6U80_2),.clk(gclk));
	jdff dff_A_LtOaC5ti7_2(.dout(w_dff_A_vbKRF6U80_2),.din(w_dff_A_LtOaC5ti7_2),.clk(gclk));
	jdff dff_A_KFtuu9GJ7_1(.dout(w_G20_3[1]),.din(w_dff_A_KFtuu9GJ7_1),.clk(gclk));
	jdff dff_A_JSzHfLnD1_2(.dout(w_G20_3[2]),.din(w_dff_A_JSzHfLnD1_2),.clk(gclk));
	jdff dff_A_ExMXZJ148_2(.dout(w_dff_A_JSzHfLnD1_2),.din(w_dff_A_ExMXZJ148_2),.clk(gclk));
	jdff dff_A_ZnOsSdK38_0(.dout(w_n390_0[0]),.din(w_dff_A_ZnOsSdK38_0),.clk(gclk));
	jdff dff_B_sTdKnjCs0_2(.din(n390),.dout(w_dff_B_sTdKnjCs0_2),.clk(gclk));
	jdff dff_A_G4hzl8R49_0(.dout(w_G87_2[0]),.din(w_dff_A_G4hzl8R49_0),.clk(gclk));
	jdff dff_A_a2K9M8PJ6_0(.dout(w_dff_A_G4hzl8R49_0),.din(w_dff_A_a2K9M8PJ6_0),.clk(gclk));
	jdff dff_A_SxnUIRhj3_0(.dout(w_dff_A_a2K9M8PJ6_0),.din(w_dff_A_SxnUIRhj3_0),.clk(gclk));
	jdff dff_A_QGVfY15l5_0(.dout(w_dff_A_SxnUIRhj3_0),.din(w_dff_A_QGVfY15l5_0),.clk(gclk));
	jdff dff_A_jbHEXkL91_1(.dout(w_G87_2[1]),.din(w_dff_A_jbHEXkL91_1),.clk(gclk));
	jdff dff_A_jWc4I7cD0_1(.dout(w_dff_A_jbHEXkL91_1),.din(w_dff_A_jWc4I7cD0_1),.clk(gclk));
	jdff dff_A_9oEPz5k67_1(.dout(w_dff_A_jWc4I7cD0_1),.din(w_dff_A_9oEPz5k67_1),.clk(gclk));
	jdff dff_A_udX6hQZn4_1(.dout(w_dff_A_9oEPz5k67_1),.din(w_dff_A_udX6hQZn4_1),.clk(gclk));
	jdff dff_A_21OGRLrO6_1(.dout(w_n149_1[1]),.din(w_dff_A_21OGRLrO6_1),.clk(gclk));
	jdff dff_A_o5lDOTfG0_1(.dout(w_dff_A_21OGRLrO6_1),.din(w_dff_A_o5lDOTfG0_1),.clk(gclk));
	jdff dff_A_cPCngAaW3_0(.dout(w_G232_1[0]),.din(w_dff_A_cPCngAaW3_0),.clk(gclk));
	jdff dff_A_kSMsUd1o0_0(.dout(w_dff_A_cPCngAaW3_0),.din(w_dff_A_kSMsUd1o0_0),.clk(gclk));
	jdff dff_A_iZGzzApM4_1(.dout(w_G232_1[1]),.din(w_dff_A_iZGzzApM4_1),.clk(gclk));
	jdff dff_A_fUYKTDQV8_1(.dout(w_G232_0[1]),.din(w_dff_A_fUYKTDQV8_1),.clk(gclk));
	jdff dff_A_GBs9BNAo1_1(.dout(w_dff_A_fUYKTDQV8_1),.din(w_dff_A_GBs9BNAo1_1),.clk(gclk));
	jdff dff_A_mI5bW7u41_1(.dout(w_dff_A_GBs9BNAo1_1),.din(w_dff_A_mI5bW7u41_1),.clk(gclk));
	jdff dff_A_ogkQdYD97_2(.dout(w_G232_0[2]),.din(w_dff_A_ogkQdYD97_2),.clk(gclk));
	jdff dff_A_fVvvUUjm7_2(.dout(w_dff_A_ogkQdYD97_2),.din(w_dff_A_fVvvUUjm7_2),.clk(gclk));
	jdff dff_A_jytAgkMy8_1(.dout(w_n539_0[1]),.din(w_dff_A_jytAgkMy8_1),.clk(gclk));
	jdff dff_B_ZsnwmpzD2_0(.din(n538),.dout(w_dff_B_ZsnwmpzD2_0),.clk(gclk));
	jdff dff_B_eFv68KBx7_0(.din(w_dff_B_ZsnwmpzD2_0),.dout(w_dff_B_eFv68KBx7_0),.clk(gclk));
	jdff dff_A_ENbhoJix7_2(.dout(w_n536_0[2]),.din(w_dff_A_ENbhoJix7_2),.clk(gclk));
	jdff dff_B_UtzkZXLy9_1(.din(n533),.dout(w_dff_B_UtzkZXLy9_1),.clk(gclk));
	jdff dff_B_UDv9v5b98_2(.din(n532),.dout(w_dff_B_UDv9v5b98_2),.clk(gclk));
	jdff dff_B_c57VbaU79_0(.din(n530),.dout(w_dff_B_c57VbaU79_0),.clk(gclk));
	jdff dff_B_Mc9vSWlq9_0(.din(w_dff_B_c57VbaU79_0),.dout(w_dff_B_Mc9vSWlq9_0),.clk(gclk));
	jdff dff_B_bJzwrDL81_1(.din(n525),.dout(w_dff_B_bJzwrDL81_1),.clk(gclk));
	jdff dff_B_0Br3Y3Xv2_0(.din(n526),.dout(w_dff_B_0Br3Y3Xv2_0),.clk(gclk));
	jdff dff_A_8E9uyBLA2_1(.dout(w_n524_0[1]),.din(w_dff_A_8E9uyBLA2_1),.clk(gclk));
	jdff dff_B_pK93kYGq3_1(.din(n521),.dout(w_dff_B_pK93kYGq3_1),.clk(gclk));
	jdff dff_A_ZB48YLv05_2(.dout(w_n588_0[2]),.din(w_dff_A_ZB48YLv05_2),.clk(gclk));
	jdff dff_B_DgFaPa4o1_0(.din(n587),.dout(w_dff_B_DgFaPa4o1_0),.clk(gclk));
	jdff dff_B_zDwXkz7L6_0(.din(w_dff_B_DgFaPa4o1_0),.dout(w_dff_B_zDwXkz7L6_0),.clk(gclk));
	jdff dff_B_xJhhQOrv7_0(.din(n585),.dout(w_dff_B_xJhhQOrv7_0),.clk(gclk));
	jdff dff_B_IymNsGxt3_1(.din(n581),.dout(w_dff_B_IymNsGxt3_1),.clk(gclk));
	jdff dff_A_OouquvDn0_1(.dout(w_n554_2[1]),.din(w_dff_A_OouquvDn0_1),.clk(gclk));
	jdff dff_A_lNlDI1Rb2_1(.dout(w_dff_A_OouquvDn0_1),.din(w_dff_A_lNlDI1Rb2_1),.clk(gclk));
	jdff dff_A_a28Q80VO5_2(.dout(w_n554_2[2]),.din(w_dff_A_a28Q80VO5_2),.clk(gclk));
	jdff dff_A_HEqpfb7G1_2(.dout(w_dff_A_a28Q80VO5_2),.din(w_dff_A_HEqpfb7G1_2),.clk(gclk));
	jdff dff_A_6qkdxHfH4_2(.dout(w_dff_A_HEqpfb7G1_2),.din(w_dff_A_6qkdxHfH4_2),.clk(gclk));
	jdff dff_A_mqvqmVgS5_2(.dout(w_dff_A_6qkdxHfH4_2),.din(w_dff_A_mqvqmVgS5_2),.clk(gclk));
	jdff dff_A_yVpbMnEO9_2(.dout(w_dff_A_mqvqmVgS5_2),.din(w_dff_A_yVpbMnEO9_2),.clk(gclk));
	jdff dff_A_5Fr6r7e69_2(.dout(w_dff_A_yVpbMnEO9_2),.din(w_dff_A_5Fr6r7e69_2),.clk(gclk));
	jdff dff_A_gymKLIgf9_0(.dout(w_n554_0[0]),.din(w_dff_A_gymKLIgf9_0),.clk(gclk));
	jdff dff_A_FMppqw4O3_0(.dout(w_dff_A_gymKLIgf9_0),.din(w_dff_A_FMppqw4O3_0),.clk(gclk));
	jdff dff_A_loB4VqjS4_2(.dout(w_n554_0[2]),.din(w_dff_A_loB4VqjS4_2),.clk(gclk));
	jdff dff_A_GIbWYEPv0_2(.dout(w_dff_A_loB4VqjS4_2),.din(w_dff_A_GIbWYEPv0_2),.clk(gclk));
	jdff dff_A_Gm6slROH2_0(.dout(w_n534_0[0]),.din(w_dff_A_Gm6slROH2_0),.clk(gclk));
	jdff dff_A_CXN2s6KH5_0(.dout(w_G179_1[0]),.din(w_dff_A_CXN2s6KH5_0),.clk(gclk));
	jdff dff_A_bmpJ6iiq1_0(.dout(w_G330_0[0]),.din(w_dff_A_bmpJ6iiq1_0),.clk(gclk));
	jdff dff_A_YcOfHab10_0(.dout(w_dff_A_bmpJ6iiq1_0),.din(w_dff_A_YcOfHab10_0),.clk(gclk));
	jdff dff_A_zdtf3Fyo1_0(.dout(w_dff_A_YcOfHab10_0),.din(w_dff_A_zdtf3Fyo1_0),.clk(gclk));
	jdff dff_A_KdM2oFPR6_0(.dout(w_dff_A_zdtf3Fyo1_0),.din(w_dff_A_KdM2oFPR6_0),.clk(gclk));
	jdff dff_A_srhLiocW2_0(.dout(w_dff_A_KdM2oFPR6_0),.din(w_dff_A_srhLiocW2_0),.clk(gclk));
	jdff dff_A_axAXm0vz6_0(.dout(w_dff_A_srhLiocW2_0),.din(w_dff_A_axAXm0vz6_0),.clk(gclk));
	jdff dff_A_4SImS4Oy6_0(.dout(w_dff_A_axAXm0vz6_0),.din(w_dff_A_4SImS4Oy6_0),.clk(gclk));
	jdff dff_A_stwUmo9O5_0(.dout(w_dff_A_4SImS4Oy6_0),.din(w_dff_A_stwUmo9O5_0),.clk(gclk));
	jdff dff_A_HfFi8Oi51_0(.dout(w_n553_2[0]),.din(w_dff_A_HfFi8Oi51_0),.clk(gclk));
	jdff dff_A_QKFIK7XV4_0(.dout(w_dff_A_HfFi8Oi51_0),.din(w_dff_A_QKFIK7XV4_0),.clk(gclk));
	jdff dff_A_lcp8cHKR3_0(.dout(w_dff_A_QKFIK7XV4_0),.din(w_dff_A_lcp8cHKR3_0),.clk(gclk));
	jdff dff_A_k928IC5l2_0(.dout(w_dff_A_lcp8cHKR3_0),.din(w_dff_A_k928IC5l2_0),.clk(gclk));
	jdff dff_A_avztiM3w5_0(.dout(w_dff_A_k928IC5l2_0),.din(w_dff_A_avztiM3w5_0),.clk(gclk));
	jdff dff_A_W0Tp6BaR2_0(.dout(w_dff_A_avztiM3w5_0),.din(w_dff_A_W0Tp6BaR2_0),.clk(gclk));
	jdff dff_A_NZPioaXJ2_0(.dout(w_dff_A_W0Tp6BaR2_0),.din(w_dff_A_NZPioaXJ2_0),.clk(gclk));
	jdff dff_A_vPczuf2F2_1(.dout(w_n553_2[1]),.din(w_dff_A_vPczuf2F2_1),.clk(gclk));
	jdff dff_A_qRayeMKr2_0(.dout(w_n553_0[0]),.din(w_dff_A_qRayeMKr2_0),.clk(gclk));
	jdff dff_A_Qmrw5kIL7_2(.dout(w_n553_0[2]),.din(w_dff_A_Qmrw5kIL7_2),.clk(gclk));
	jdff dff_A_iv2p9UGR7_2(.dout(w_dff_A_Qmrw5kIL7_2),.din(w_dff_A_iv2p9UGR7_2),.clk(gclk));
	jdff dff_A_YaTQG0RH8_2(.dout(w_dff_A_iv2p9UGR7_2),.din(w_dff_A_YaTQG0RH8_2),.clk(gclk));
	jdff dff_A_r3TYdPRz8_1(.dout(w_n552_0[1]),.din(w_dff_A_r3TYdPRz8_1),.clk(gclk));
	jdff dff_A_HHT873W73_1(.dout(w_dff_A_r3TYdPRz8_1),.din(w_dff_A_HHT873W73_1),.clk(gclk));
	jdff dff_A_TupEKacE0_1(.dout(w_dff_A_HHT873W73_1),.din(w_dff_A_TupEKacE0_1),.clk(gclk));
	jdff dff_A_7cFzR9Dh8_1(.dout(w_dff_A_TupEKacE0_1),.din(w_dff_A_7cFzR9Dh8_1),.clk(gclk));
	jdff dff_A_tQVBHVvz7_1(.dout(w_dff_A_7cFzR9Dh8_1),.din(w_dff_A_tQVBHVvz7_1),.clk(gclk));
	jdff dff_A_P3wnx4oD8_1(.dout(w_dff_A_tQVBHVvz7_1),.din(w_dff_A_P3wnx4oD8_1),.clk(gclk));
	jdff dff_A_lQLBJZEQ1_2(.dout(w_n552_0[2]),.din(w_dff_A_lQLBJZEQ1_2),.clk(gclk));
	jdff dff_A_vSxQjJ4X3_2(.dout(w_dff_A_lQLBJZEQ1_2),.din(w_dff_A_vSxQjJ4X3_2),.clk(gclk));
	jdff dff_A_qMrvZvq50_2(.dout(w_dff_A_vSxQjJ4X3_2),.din(w_dff_A_qMrvZvq50_2),.clk(gclk));
	jdff dff_A_hX56HpIG0_2(.dout(w_dff_A_qMrvZvq50_2),.din(w_dff_A_hX56HpIG0_2),.clk(gclk));
	jdff dff_A_UfVmVae33_2(.dout(w_dff_A_hX56HpIG0_2),.din(w_dff_A_UfVmVae33_2),.clk(gclk));
	jdff dff_A_ploXWUQo9_0(.dout(w_G213_0[0]),.din(w_dff_A_ploXWUQo9_0),.clk(gclk));
	jdff dff_A_ojWxuxiD0_2(.dout(w_G213_0[2]),.din(w_dff_A_ojWxuxiD0_2),.clk(gclk));
	jdff dff_A_zrSwBRGm1_0(.dout(w_n113_1[0]),.din(w_dff_A_zrSwBRGm1_0),.clk(gclk));
	jdff dff_A_MANApDwJ0_0(.dout(w_dff_A_zrSwBRGm1_0),.din(w_dff_A_MANApDwJ0_0),.clk(gclk));
	jdff dff_A_cFPEjfVC8_1(.dout(w_n113_1[1]),.din(w_dff_A_cFPEjfVC8_1),.clk(gclk));
	jdff dff_A_l7lSQxMl7_1(.dout(w_dff_A_cFPEjfVC8_1),.din(w_dff_A_l7lSQxMl7_1),.clk(gclk));
	jdff dff_A_juWXiyw33_1(.dout(w_dff_A_l7lSQxMl7_1),.din(w_dff_A_juWXiyw33_1),.clk(gclk));
	jdff dff_A_bq9azBta7_1(.dout(w_dff_A_juWXiyw33_1),.din(w_dff_A_bq9azBta7_1),.clk(gclk));
	jdff dff_A_QSNq6Oc96_1(.dout(w_dff_A_bq9azBta7_1),.din(w_dff_A_QSNq6Oc96_1),.clk(gclk));
	jdff dff_A_pgCw6MNt0_1(.dout(w_dff_A_QSNq6Oc96_1),.din(w_dff_A_pgCw6MNt0_1),.clk(gclk));
	jdff dff_A_ogwZrAhS2_1(.dout(w_dff_A_pgCw6MNt0_1),.din(w_dff_A_ogwZrAhS2_1),.clk(gclk));
	jdff dff_A_k8fhh1kp1_1(.dout(w_dff_A_ogwZrAhS2_1),.din(w_dff_A_k8fhh1kp1_1),.clk(gclk));
	jdff dff_A_0CemE09k5_1(.dout(w_dff_A_k8fhh1kp1_1),.din(w_dff_A_0CemE09k5_1),.clk(gclk));
	jdff dff_A_QUMlrFU18_1(.dout(w_dff_A_0CemE09k5_1),.din(w_dff_A_QUMlrFU18_1),.clk(gclk));
	jdff dff_A_WdJmdwBX6_1(.dout(w_dff_A_QUMlrFU18_1),.din(w_dff_A_WdJmdwBX6_1),.clk(gclk));
	jdff dff_A_f9zbZg4C8_1(.dout(w_G343_0[1]),.din(w_dff_A_f9zbZg4C8_1),.clk(gclk));
	jdff dff_A_2wRSdLNF4_1(.dout(w_dff_A_f9zbZg4C8_1),.din(w_dff_A_2wRSdLNF4_1),.clk(gclk));
	jdff dff_A_9bWExnt25_1(.dout(w_dff_A_2wRSdLNF4_1),.din(w_dff_A_9bWExnt25_1),.clk(gclk));
	jdff dff_A_aLEHXo812_1(.dout(w_n374_0[1]),.din(w_dff_A_aLEHXo812_1),.clk(gclk));
	jdff dff_B_wirumzpe5_0(.din(n373),.dout(w_dff_B_wirumzpe5_0),.clk(gclk));
	jdff dff_B_IzQrH9399_2(.din(n371),.dout(w_dff_B_IzQrH9399_2),.clk(gclk));
	jdff dff_B_8fOJpo850_1(.din(n368),.dout(w_dff_B_8fOJpo850_1),.clk(gclk));
	jdff dff_A_oLRdNPdw6_2(.dout(w_G200_3[2]),.din(w_dff_A_oLRdNPdw6_2),.clk(gclk));
	jdff dff_A_nP6h92hb4_1(.dout(w_n367_0[1]),.din(w_dff_A_nP6h92hb4_1),.clk(gclk));
	jdff dff_A_t0iXcEPt3_2(.dout(w_n367_0[2]),.din(w_dff_A_t0iXcEPt3_2),.clk(gclk));
	jdff dff_B_qA13Ndc32_0(.din(n365),.dout(w_dff_B_qA13Ndc32_0),.clk(gclk));
	jdff dff_B_yTEEUpH48_0(.din(n357),.dout(w_dff_B_yTEEUpH48_0),.clk(gclk));
	jdff dff_B_fc3BiEcZ2_0(.din(n356),.dout(w_dff_B_fc3BiEcZ2_0),.clk(gclk));
	jdff dff_B_zYYggNLe3_0(.din(n353),.dout(w_dff_B_zYYggNLe3_0),.clk(gclk));
	jdff dff_B_nh7xxYWg9_1(.din(n337),.dout(w_dff_B_nh7xxYWg9_1),.clk(gclk));
	jdff dff_B_L6FeC3JP5_1(.din(w_dff_B_nh7xxYWg9_1),.dout(w_dff_B_L6FeC3JP5_1),.clk(gclk));
	jdff dff_B_i14Gol6C4_1(.din(n338),.dout(w_dff_B_i14Gol6C4_1),.clk(gclk));
	jdff dff_A_0NDHMjEF6_0(.dout(w_n339_0[0]),.din(w_dff_A_0NDHMjEF6_0),.clk(gclk));
	jdff dff_A_g7sa2qLA6_0(.dout(w_dff_A_0NDHMjEF6_0),.din(w_dff_A_g7sa2qLA6_0),.clk(gclk));
	jdff dff_A_9ZQvLSfa8_0(.dout(w_G294_3[0]),.din(w_dff_A_9ZQvLSfa8_0),.clk(gclk));
	jdff dff_A_hjgbbSVR8_0(.dout(w_dff_A_9ZQvLSfa8_0),.din(w_dff_A_hjgbbSVR8_0),.clk(gclk));
	jdff dff_A_LKMSibzd4_0(.dout(w_dff_A_hjgbbSVR8_0),.din(w_dff_A_LKMSibzd4_0),.clk(gclk));
	jdff dff_A_uqeqgqm72_0(.dout(w_dff_A_LKMSibzd4_0),.din(w_dff_A_uqeqgqm72_0),.clk(gclk));
	jdff dff_A_zT5VIxUQ5_0(.dout(w_G294_0[0]),.din(w_dff_A_zT5VIxUQ5_0),.clk(gclk));
	jdff dff_A_nYiQUxpz5_0(.dout(w_dff_A_zT5VIxUQ5_0),.din(w_dff_A_nYiQUxpz5_0),.clk(gclk));
	jdff dff_A_OtV27sqM7_0(.dout(w_dff_A_nYiQUxpz5_0),.din(w_dff_A_OtV27sqM7_0),.clk(gclk));
	jdff dff_A_8gxL498K9_1(.dout(w_G294_0[1]),.din(w_dff_A_8gxL498K9_1),.clk(gclk));
	jdff dff_A_X8ZBCkA41_1(.dout(w_dff_A_8gxL498K9_1),.din(w_dff_A_X8ZBCkA41_1),.clk(gclk));
	jdff dff_A_As1zAiFl1_1(.dout(w_dff_A_X8ZBCkA41_1),.din(w_dff_A_As1zAiFl1_1),.clk(gclk));
	jdff dff_B_WgAINPb89_1(.din(n332),.dout(w_dff_B_WgAINPb89_1),.clk(gclk));
	jdff dff_B_wewM4ZSQ5_1(.din(w_dff_B_WgAINPb89_1),.dout(w_dff_B_wewM4ZSQ5_1),.clk(gclk));
	jdff dff_A_l8rs1oAb6_0(.dout(w_G107_3[0]),.din(w_dff_A_l8rs1oAb6_0),.clk(gclk));
	jdff dff_A_ybYp2lXE1_1(.dout(w_G107_3[1]),.din(w_dff_A_ybYp2lXE1_1),.clk(gclk));
	jdff dff_B_w4Awezhr4_0(.din(n323),.dout(w_dff_B_w4Awezhr4_0),.clk(gclk));
	jdff dff_B_BzP9mOHK2_1(.din(n316),.dout(w_dff_B_BzP9mOHK2_1),.clk(gclk));
	jdff dff_A_NaxlSU6n5_1(.dout(w_G190_3[1]),.din(w_dff_A_NaxlSU6n5_1),.clk(gclk));
	jdff dff_A_ifeXtB8u5_1(.dout(w_dff_A_NaxlSU6n5_1),.din(w_dff_A_ifeXtB8u5_1),.clk(gclk));
	jdff dff_A_2J23iolI4_1(.dout(w_dff_A_ifeXtB8u5_1),.din(w_dff_A_2J23iolI4_1),.clk(gclk));
	jdff dff_A_izkfXpqB4_1(.dout(w_dff_A_2J23iolI4_1),.din(w_dff_A_izkfXpqB4_1),.clk(gclk));
	jdff dff_A_Rda2fYaU8_2(.dout(w_G190_3[2]),.din(w_dff_A_Rda2fYaU8_2),.clk(gclk));
	jdff dff_A_ZFm3XZBk4_2(.dout(w_dff_A_Rda2fYaU8_2),.din(w_dff_A_ZFm3XZBk4_2),.clk(gclk));
	jdff dff_A_HK9oBtJF2_2(.dout(w_dff_A_ZFm3XZBk4_2),.din(w_dff_A_HK9oBtJF2_2),.clk(gclk));
	jdff dff_A_XEEFmGT81_2(.dout(w_dff_A_HK9oBtJF2_2),.din(w_dff_A_XEEFmGT81_2),.clk(gclk));
	jdff dff_A_y8Uk3cet7_2(.dout(w_dff_A_XEEFmGT81_2),.din(w_dff_A_y8Uk3cet7_2),.clk(gclk));
	jdff dff_A_t5wxuhce7_1(.dout(w_n320_0[1]),.din(w_dff_A_t5wxuhce7_1),.clk(gclk));
	jdff dff_B_jwuRkkXK5_0(.din(n319),.dout(w_dff_B_jwuRkkXK5_0),.clk(gclk));
	jdff dff_B_zO1IRGag5_1(.din(n289),.dout(w_dff_B_zO1IRGag5_1),.clk(gclk));
	jdff dff_B_eta8Muoc4_1(.din(w_dff_B_zO1IRGag5_1),.dout(w_dff_B_eta8Muoc4_1),.clk(gclk));
	jdff dff_B_lrDaUowg2_0(.din(n313),.dout(w_dff_B_lrDaUowg2_0),.clk(gclk));
	jdff dff_A_8G0arO6g1_1(.dout(w_n312_0[1]),.din(w_dff_A_8G0arO6g1_1),.clk(gclk));
	jdff dff_A_pGVeTZBk0_0(.dout(w_n106_0[0]),.din(w_dff_A_pGVeTZBk0_0),.clk(gclk));
	jdff dff_A_FDiH7MW27_0(.dout(w_dff_A_pGVeTZBk0_0),.din(w_dff_A_FDiH7MW27_0),.clk(gclk));
	jdff dff_B_FO8Gwv0J1_1(.din(n304),.dout(w_dff_B_FO8Gwv0J1_1),.clk(gclk));
	jdff dff_B_K7z4jg7I0_1(.din(w_dff_B_FO8Gwv0J1_1),.dout(w_dff_B_K7z4jg7I0_1),.clk(gclk));
	jdff dff_B_NBjz2sFV6_0(.din(n306),.dout(w_dff_B_NBjz2sFV6_0),.clk(gclk));
	jdff dff_A_4386Ygz54_1(.dout(w_n88_0[1]),.din(w_dff_A_4386Ygz54_1),.clk(gclk));
	jdff dff_A_i99ftJfc5_1(.dout(w_dff_A_4386Ygz54_1),.din(w_dff_A_i99ftJfc5_1),.clk(gclk));
	jdff dff_A_beC0eKaG7_1(.dout(w_n166_1[1]),.din(w_dff_A_beC0eKaG7_1),.clk(gclk));
	jdff dff_A_ONukrniH5_1(.dout(w_dff_A_beC0eKaG7_1),.din(w_dff_A_ONukrniH5_1),.clk(gclk));
	jdff dff_A_AsGZYBOs7_2(.dout(w_n166_1[2]),.din(w_dff_A_AsGZYBOs7_2),.clk(gclk));
	jdff dff_A_2FUbW2rT0_2(.dout(w_dff_A_AsGZYBOs7_2),.din(w_dff_A_2FUbW2rT0_2),.clk(gclk));
	jdff dff_B_prqkqRTk6_0(.din(n301),.dout(w_dff_B_prqkqRTk6_0),.clk(gclk));
	jdff dff_B_N3cNAHsT0_0(.din(w_dff_B_prqkqRTk6_0),.dout(w_dff_B_N3cNAHsT0_0),.clk(gclk));
	jdff dff_A_8TdrWGBZ9_1(.dout(w_n300_0[1]),.din(w_dff_A_8TdrWGBZ9_1),.clk(gclk));
	jdff dff_A_rvC2vt7T8_0(.dout(w_n105_1[0]),.din(w_dff_A_rvC2vt7T8_0),.clk(gclk));
	jdff dff_A_9ZunfM6Y5_2(.dout(w_n105_1[2]),.din(w_dff_A_9ZunfM6Y5_2),.clk(gclk));
	jdff dff_B_lw8HqzXo4_1(.din(n292),.dout(w_dff_B_lw8HqzXo4_1),.clk(gclk));
	jdff dff_B_I8qsIiur3_1(.din(w_dff_B_lw8HqzXo4_1),.dout(w_dff_B_I8qsIiur3_1),.clk(gclk));
	jdff dff_A_GQxHmHkp4_0(.dout(w_n105_0[0]),.din(w_dff_A_GQxHmHkp4_0),.clk(gclk));
	jdff dff_A_CCEoeB2a5_2(.dout(w_n105_0[2]),.din(w_dff_A_CCEoeB2a5_2),.clk(gclk));
	jdff dff_A_hcTSn3R21_2(.dout(w_dff_A_CCEoeB2a5_2),.din(w_dff_A_hcTSn3R21_2),.clk(gclk));
	jdff dff_A_XqgdXkng9_2(.dout(w_dff_A_hcTSn3R21_2),.din(w_dff_A_XqgdXkng9_2),.clk(gclk));
	jdff dff_A_FrLgA80Y5_0(.dout(w_G20_4[0]),.din(w_dff_A_FrLgA80Y5_0),.clk(gclk));
	jdff dff_A_hxr1AAEs1_1(.dout(w_G20_4[1]),.din(w_dff_A_hxr1AAEs1_1),.clk(gclk));
	jdff dff_A_BiQXPWQW1_1(.dout(w_dff_A_hxr1AAEs1_1),.din(w_dff_A_BiQXPWQW1_1),.clk(gclk));
	jdff dff_A_BJu1r9gt1_2(.dout(w_n189_1[2]),.din(w_dff_A_BJu1r9gt1_2),.clk(gclk));
	jdff dff_A_97bTYVVD3_0(.dout(w_G97_3[0]),.din(w_dff_A_97bTYVVD3_0),.clk(gclk));
	jdff dff_A_0HiOQMRJ8_0(.dout(w_dff_A_97bTYVVD3_0),.din(w_dff_A_0HiOQMRJ8_0),.clk(gclk));
	jdff dff_A_O2VcMFTg2_0(.dout(w_dff_A_0HiOQMRJ8_0),.din(w_dff_A_O2VcMFTg2_0),.clk(gclk));
	jdff dff_A_6QVyZ4HI3_1(.dout(w_G97_3[1]),.din(w_dff_A_6QVyZ4HI3_1),.clk(gclk));
	jdff dff_A_Kw9nV4ns7_1(.dout(w_dff_A_6QVyZ4HI3_1),.din(w_dff_A_Kw9nV4ns7_1),.clk(gclk));
	jdff dff_A_RZwJTBHH0_1(.dout(w_dff_A_Kw9nV4ns7_1),.din(w_dff_A_RZwJTBHH0_1),.clk(gclk));
	jdff dff_B_l1NMarM66_0(.din(n286),.dout(w_dff_B_l1NMarM66_0),.clk(gclk));
	jdff dff_A_CQRgG1Mw5_0(.dout(w_G270_0[0]),.din(w_dff_A_CQRgG1Mw5_0),.clk(gclk));
	jdff dff_A_uShzZ3Uv1_0(.dout(w_dff_A_CQRgG1Mw5_0),.din(w_dff_A_uShzZ3Uv1_0),.clk(gclk));
	jdff dff_A_al7IYk3V8_1(.dout(w_n281_0[1]),.din(w_dff_A_al7IYk3V8_1),.clk(gclk));
	jdff dff_A_WnxFzNr57_1(.dout(w_dff_A_al7IYk3V8_1),.din(w_dff_A_WnxFzNr57_1),.clk(gclk));
	jdff dff_A_PDL6C3nK3_0(.dout(w_G303_2[0]),.din(w_dff_A_PDL6C3nK3_0),.clk(gclk));
	jdff dff_A_GmVYZNx38_0(.dout(w_dff_A_PDL6C3nK3_0),.din(w_dff_A_GmVYZNx38_0),.clk(gclk));
	jdff dff_A_6SZHnbiP5_0(.dout(w_dff_A_GmVYZNx38_0),.din(w_dff_A_6SZHnbiP5_0),.clk(gclk));
	jdff dff_A_UQq57QqN0_1(.dout(w_G303_2[1]),.din(w_dff_A_UQq57QqN0_1),.clk(gclk));
	jdff dff_A_GawpsW3m4_1(.dout(w_dff_A_UQq57QqN0_1),.din(w_dff_A_GawpsW3m4_1),.clk(gclk));
	jdff dff_A_g7WmM91Q2_1(.dout(w_dff_A_GawpsW3m4_1),.din(w_dff_A_g7WmM91Q2_1),.clk(gclk));
	jdff dff_A_n2oDV0SI8_1(.dout(w_dff_A_g7WmM91Q2_1),.din(w_dff_A_n2oDV0SI8_1),.clk(gclk));
	jdff dff_A_b9bC12Y00_0(.dout(w_G303_0[0]),.din(w_dff_A_b9bC12Y00_0),.clk(gclk));
	jdff dff_A_UYQbUqrz6_0(.dout(w_dff_A_b9bC12Y00_0),.din(w_dff_A_UYQbUqrz6_0),.clk(gclk));
	jdff dff_A_O00dREir7_0(.dout(w_dff_A_UYQbUqrz6_0),.din(w_dff_A_O00dREir7_0),.clk(gclk));
	jdff dff_A_iniuKwvB2_2(.dout(w_G303_0[2]),.din(w_dff_A_iniuKwvB2_2),.clk(gclk));
	jdff dff_A_biPj3nGp6_2(.dout(w_dff_A_iniuKwvB2_2),.din(w_dff_A_biPj3nGp6_2),.clk(gclk));
	jdff dff_A_nzLoglhV6_2(.dout(w_dff_A_biPj3nGp6_2),.din(w_dff_A_nzLoglhV6_2),.clk(gclk));
	jdff dff_A_W8LYVIsw3_1(.dout(w_G264_0[1]),.din(w_dff_A_W8LYVIsw3_1),.clk(gclk));
	jdff dff_A_YBHsC95D4_1(.dout(w_dff_A_W8LYVIsw3_1),.din(w_dff_A_YBHsC95D4_1),.clk(gclk));
	jdff dff_A_axinjCBL2_2(.dout(w_G264_0[2]),.din(w_dff_A_axinjCBL2_2),.clk(gclk));
	jdff dff_A_j7dOrHzR6_2(.dout(w_dff_A_axinjCBL2_2),.din(w_dff_A_j7dOrHzR6_2),.clk(gclk));
	jdff dff_A_TH2JGvDg9_1(.dout(w_n278_0[1]),.din(w_dff_A_TH2JGvDg9_1),.clk(gclk));
	jdff dff_B_zBzpHhf81_0(.din(n277),.dout(w_dff_B_zBzpHhf81_0),.clk(gclk));
	jdff dff_B_OaAB421S6_1(.din(n268),.dout(w_dff_B_OaAB421S6_1),.clk(gclk));
	jdff dff_A_TuWqKq408_1(.dout(w_n274_0[1]),.din(w_dff_A_TuWqKq408_1),.clk(gclk));
	jdff dff_A_OHCadVq27_2(.dout(w_n274_0[2]),.din(w_dff_A_OHCadVq27_2),.clk(gclk));
	jdff dff_A_cYYAdWbW6_0(.dout(w_n271_1[0]),.din(w_dff_A_cYYAdWbW6_0),.clk(gclk));
	jdff dff_A_RovLMnhq5_2(.dout(w_n271_1[2]),.din(w_dff_A_RovLMnhq5_2),.clk(gclk));
	jdff dff_A_b7wLZy7l7_0(.dout(w_n270_0[0]),.din(w_dff_A_b7wLZy7l7_0),.clk(gclk));
	jdff dff_B_GHq7vOay5_2(.din(n270),.dout(w_dff_B_GHq7vOay5_2),.clk(gclk));
	jdff dff_A_cTwrrY2b4_0(.dout(w_n112_4[0]),.din(w_dff_A_cTwrrY2b4_0),.clk(gclk));
	jdff dff_A_tIMCN33B9_0(.dout(w_dff_A_cTwrrY2b4_0),.din(w_dff_A_tIMCN33B9_0),.clk(gclk));
	jdff dff_A_JgdntH6e3_0(.dout(w_G1_1[0]),.din(w_dff_A_JgdntH6e3_0),.clk(gclk));
	jdff dff_A_e9A7km2s9_0(.dout(w_dff_A_JgdntH6e3_0),.din(w_dff_A_e9A7km2s9_0),.clk(gclk));
	jdff dff_A_Fou26Hox4_0(.dout(w_dff_A_e9A7km2s9_0),.din(w_dff_A_Fou26Hox4_0),.clk(gclk));
	jdff dff_A_tZAQhP2l8_1(.dout(w_G1_1[1]),.din(w_dff_A_tZAQhP2l8_1),.clk(gclk));
	jdff dff_B_7U7WpZzl4_1(.din(n248),.dout(w_dff_B_7U7WpZzl4_1),.clk(gclk));
	jdff dff_B_JIOC8EHz8_1(.din(n258),.dout(w_dff_B_JIOC8EHz8_1),.clk(gclk));
	jdff dff_A_mU3DqGOy2_0(.dout(w_n259_0[0]),.din(w_dff_A_mU3DqGOy2_0),.clk(gclk));
	jdff dff_A_b6fZpL3E6_0(.dout(w_n257_0[0]),.din(w_dff_A_b6fZpL3E6_0),.clk(gclk));
	jdff dff_B_I5nmTvxU4_0(.din(n254),.dout(w_dff_B_I5nmTvxU4_0),.clk(gclk));
	jdff dff_A_JeMaVs6t4_0(.dout(w_G77_1[0]),.din(w_dff_A_JeMaVs6t4_0),.clk(gclk));
	jdff dff_A_h9DR7GMP4_2(.dout(w_G77_1[2]),.din(w_dff_A_h9DR7GMP4_2),.clk(gclk));
	jdff dff_A_8CzCP1zt1_2(.dout(w_dff_A_h9DR7GMP4_2),.din(w_dff_A_8CzCP1zt1_2),.clk(gclk));
	jdff dff_A_rsQJNHKW4_2(.dout(w_dff_A_8CzCP1zt1_2),.din(w_dff_A_rsQJNHKW4_2),.clk(gclk));
	jdff dff_A_8sWGGBbl3_2(.dout(w_dff_A_rsQJNHKW4_2),.din(w_dff_A_8sWGGBbl3_2),.clk(gclk));
	jdff dff_A_EWkT1AOP3_0(.dout(w_n249_0[0]),.din(w_dff_A_EWkT1AOP3_0),.clk(gclk));
	jdff dff_B_PT24TNez2_2(.din(n249),.dout(w_dff_B_PT24TNez2_2),.clk(gclk));
	jdff dff_A_rcOOxg1z3_0(.dout(w_G107_4[0]),.din(w_dff_A_rcOOxg1z3_0),.clk(gclk));
	jdff dff_A_mbURjbvu7_0(.dout(w_dff_A_rcOOxg1z3_0),.din(w_dff_A_mbURjbvu7_0),.clk(gclk));
	jdff dff_A_ygo3ADFz2_0(.dout(w_dff_A_mbURjbvu7_0),.din(w_dff_A_ygo3ADFz2_0),.clk(gclk));
	jdff dff_A_tIDm05Cz1_0(.dout(w_G33_8[0]),.din(w_dff_A_tIDm05Cz1_0),.clk(gclk));
	jdff dff_B_xIKDQVJe5_0(.din(n247),.dout(w_dff_B_xIKDQVJe5_0),.clk(gclk));
	jdff dff_B_crRIzxv97_0(.din(n244),.dout(w_dff_B_crRIzxv97_0),.clk(gclk));
	jdff dff_B_HZzECxmh4_2(.din(n241),.dout(w_dff_B_HZzECxmh4_2),.clk(gclk));
	jdff dff_A_HYmMZDFV0_0(.dout(w_n91_1[0]),.din(w_dff_A_HYmMZDFV0_0),.clk(gclk));
	jdff dff_A_PwEDttqh4_0(.dout(w_dff_A_HYmMZDFV0_0),.din(w_dff_A_PwEDttqh4_0),.clk(gclk));
	jdff dff_A_94KTuCpr8_0(.dout(w_G257_1[0]),.din(w_dff_A_94KTuCpr8_0),.clk(gclk));
	jdff dff_A_ydIkuUtG6_0(.dout(w_dff_A_94KTuCpr8_0),.din(w_dff_A_ydIkuUtG6_0),.clk(gclk));
	jdff dff_A_cZljE8hi0_1(.dout(w_G257_1[1]),.din(w_dff_A_cZljE8hi0_1),.clk(gclk));
	jdff dff_A_SgbIM5EI2_1(.dout(w_G257_0[1]),.din(w_dff_A_SgbIM5EI2_1),.clk(gclk));
	jdff dff_A_Ny0Ff4VQ5_1(.dout(w_dff_A_SgbIM5EI2_1),.din(w_dff_A_Ny0Ff4VQ5_1),.clk(gclk));
	jdff dff_A_1vvZxFoU0_2(.dout(w_G257_0[2]),.din(w_dff_A_1vvZxFoU0_2),.clk(gclk));
	jdff dff_A_eo3IM3vo2_2(.dout(w_dff_A_1vvZxFoU0_2),.din(w_dff_A_eo3IM3vo2_2),.clk(gclk));
	jdff dff_B_lS3T56Se1_3(.din(n229),.dout(w_dff_B_lS3T56Se1_3),.clk(gclk));
	jdff dff_A_xhAvvTf95_1(.dout(w_n228_0[1]),.din(w_dff_A_xhAvvTf95_1),.clk(gclk));
	jdff dff_B_cKunexlm0_1(.din(n220),.dout(w_dff_B_cKunexlm0_1),.clk(gclk));
	jdff dff_B_9COU33x02_1(.din(w_dff_B_cKunexlm0_1),.dout(w_dff_B_9COU33x02_1),.clk(gclk));
	jdff dff_B_GhdvqHhs9_0(.din(n223),.dout(w_dff_B_GhdvqHhs9_0),.clk(gclk));
	jdff dff_A_xMCwb3Xo0_0(.dout(w_n221_0[0]),.din(w_dff_A_xMCwb3Xo0_0),.clk(gclk));
	jdff dff_A_cTRfOIBm7_1(.dout(w_n221_0[1]),.din(w_dff_A_cTRfOIBm7_1),.clk(gclk));
	jdff dff_A_ugZr37UL0_1(.dout(w_dff_A_cTRfOIBm7_1),.din(w_dff_A_ugZr37UL0_1),.clk(gclk));
	jdff dff_A_4JO5gZAH2_0(.dout(w_G283_3[0]),.din(w_dff_A_4JO5gZAH2_0),.clk(gclk));
	jdff dff_A_k8oJfmuI6_0(.dout(w_dff_A_4JO5gZAH2_0),.din(w_dff_A_k8oJfmuI6_0),.clk(gclk));
	jdff dff_A_2JC8ADef4_0(.dout(w_dff_A_k8oJfmuI6_0),.din(w_dff_A_2JC8ADef4_0),.clk(gclk));
	jdff dff_A_8tLQ4KOD3_1(.dout(w_G283_3[1]),.din(w_dff_A_8tLQ4KOD3_1),.clk(gclk));
	jdff dff_A_jmu46CmJ4_1(.dout(w_dff_A_8tLQ4KOD3_1),.din(w_dff_A_jmu46CmJ4_1),.clk(gclk));
	jdff dff_A_wiJr0S7S8_1(.dout(w_dff_A_jmu46CmJ4_1),.din(w_dff_A_wiJr0S7S8_1),.clk(gclk));
	jdff dff_A_QADLD1h01_1(.dout(w_dff_A_wiJr0S7S8_1),.din(w_dff_A_QADLD1h01_1),.clk(gclk));
	jdff dff_A_icbPBZjK5_0(.dout(w_G283_0[0]),.din(w_dff_A_icbPBZjK5_0),.clk(gclk));
	jdff dff_A_muro9qR59_0(.dout(w_dff_A_icbPBZjK5_0),.din(w_dff_A_muro9qR59_0),.clk(gclk));
	jdff dff_A_9J0G4DIm3_0(.dout(w_dff_A_muro9qR59_0),.din(w_dff_A_9J0G4DIm3_0),.clk(gclk));
	jdff dff_A_jqGbUiad9_1(.dout(w_G283_0[1]),.din(w_dff_A_jqGbUiad9_1),.clk(gclk));
	jdff dff_A_7KaqsGwY4_1(.dout(w_dff_A_jqGbUiad9_1),.din(w_dff_A_7KaqsGwY4_1),.clk(gclk));
	jdff dff_A_HY0WJrlP2_1(.dout(w_dff_A_7KaqsGwY4_1),.din(w_dff_A_HY0WJrlP2_1),.clk(gclk));
	jdff dff_A_PO9MuSmM7_2(.dout(w_n166_2[2]),.din(w_dff_A_PO9MuSmM7_2),.clk(gclk));
	jdff dff_A_44PSQTCf1_2(.dout(w_dff_A_PO9MuSmM7_2),.din(w_dff_A_44PSQTCf1_2),.clk(gclk));
	jdff dff_A_NdF95UbF0_2(.dout(w_dff_A_44PSQTCf1_2),.din(w_dff_A_NdF95UbF0_2),.clk(gclk));
	jdff dff_A_2Y721u017_0(.dout(w_n219_0[0]),.din(w_dff_A_2Y721u017_0),.clk(gclk));
	jdff dff_B_hFHsXgb73_0(.din(n217),.dout(w_dff_B_hFHsXgb73_0),.clk(gclk));
	jdff dff_B_GRlG9TWL1_0(.din(w_dff_B_hFHsXgb73_0),.dout(w_dff_B_GRlG9TWL1_0),.clk(gclk));
	jdff dff_B_q0dCNmqv6_0(.din(n216),.dout(w_dff_B_q0dCNmqv6_0),.clk(gclk));
	jdff dff_A_Li4Jjbkf8_0(.dout(w_G200_1[0]),.din(w_dff_A_Li4Jjbkf8_0),.clk(gclk));
	jdff dff_A_v9EzSQWy9_0(.dout(w_dff_A_Li4Jjbkf8_0),.din(w_dff_A_v9EzSQWy9_0),.clk(gclk));
	jdff dff_A_sVsvKSQR7_0(.dout(w_dff_A_v9EzSQWy9_0),.din(w_dff_A_sVsvKSQR7_0),.clk(gclk));
	jdff dff_A_Cxmm5ts75_0(.dout(w_dff_A_sVsvKSQR7_0),.din(w_dff_A_Cxmm5ts75_0),.clk(gclk));
	jdff dff_A_dmI39b8w6_1(.dout(w_G200_1[1]),.din(w_dff_A_dmI39b8w6_1),.clk(gclk));
	jdff dff_A_t54hNTpi6_2(.dout(w_G200_0[2]),.din(w_dff_A_t54hNTpi6_2),.clk(gclk));
	jdff dff_A_pxALCa0e1_2(.dout(w_dff_A_t54hNTpi6_2),.din(w_dff_A_pxALCa0e1_2),.clk(gclk));
	jdff dff_A_Jyv2PZ9J5_2(.dout(w_dff_A_pxALCa0e1_2),.din(w_dff_A_Jyv2PZ9J5_2),.clk(gclk));
	jdff dff_A_UviIzfNq3_2(.dout(w_dff_A_Jyv2PZ9J5_2),.din(w_dff_A_UviIzfNq3_2),.clk(gclk));
	jdff dff_A_DFkFYigY0_0(.dout(w_G190_1[0]),.din(w_dff_A_DFkFYigY0_0),.clk(gclk));
	jdff dff_A_4kDaLvsJ5_0(.dout(w_dff_A_DFkFYigY0_0),.din(w_dff_A_4kDaLvsJ5_0),.clk(gclk));
	jdff dff_A_BfNynjZ25_0(.dout(w_dff_A_4kDaLvsJ5_0),.din(w_dff_A_BfNynjZ25_0),.clk(gclk));
	jdff dff_A_FpJre54a5_0(.dout(w_G190_0[0]),.din(w_dff_A_FpJre54a5_0),.clk(gclk));
	jdff dff_A_RUd1jwHC1_0(.dout(w_dff_A_FpJre54a5_0),.din(w_dff_A_RUd1jwHC1_0),.clk(gclk));
	jdff dff_A_ti81mePK8_1(.dout(w_G190_0[1]),.din(w_dff_A_ti81mePK8_1),.clk(gclk));
	jdff dff_A_C3y9u9Zz6_1(.dout(w_dff_A_ti81mePK8_1),.din(w_dff_A_C3y9u9Zz6_1),.clk(gclk));
	jdff dff_A_1dXG9ppK9_1(.dout(w_dff_A_C3y9u9Zz6_1),.din(w_dff_A_1dXG9ppK9_1),.clk(gclk));
	jdff dff_A_4d3ZXjKD6_1(.dout(w_n213_0[1]),.din(w_dff_A_4d3ZXjKD6_1),.clk(gclk));
	jdff dff_B_xmYl4AbE2_1(.din(n171),.dout(w_dff_B_xmYl4AbE2_1),.clk(gclk));
	jdff dff_B_bFExBmbu0_1(.din(w_dff_B_xmYl4AbE2_1),.dout(w_dff_B_bFExBmbu0_1),.clk(gclk));
	jdff dff_B_1cfpiNrB1_0(.din(n211),.dout(w_dff_B_1cfpiNrB1_0),.clk(gclk));
	jdff dff_B_xzZaUamp2_0(.din(n209),.dout(w_dff_B_xzZaUamp2_0),.clk(gclk));
	jdff dff_B_EGl2WplV9_2(.din(n205),.dout(w_dff_B_EGl2WplV9_2),.clk(gclk));
	jdff dff_B_tQ5bBQum0_1(.din(n198),.dout(w_dff_B_tQ5bBQum0_1),.clk(gclk));
	jdff dff_B_PrZaD5Zv0_1(.din(w_dff_B_tQ5bBQum0_1),.dout(w_dff_B_PrZaD5Zv0_1),.clk(gclk));
	jdff dff_B_5wPozv1I6_1(.din(n200),.dout(w_dff_B_5wPozv1I6_1),.clk(gclk));
	jdff dff_B_ZoCsYINS5_3(.din(n199),.dout(w_dff_B_ZoCsYINS5_3),.clk(gclk));
	jdff dff_A_y5rIwcE93_2(.dout(w_G33_9[2]),.din(w_dff_A_y5rIwcE93_2),.clk(gclk));
	jdff dff_A_siocPJva6_0(.dout(w_n196_2[0]),.din(w_dff_A_siocPJva6_0),.clk(gclk));
	jdff dff_A_UxntVVz47_2(.dout(w_n196_2[2]),.din(w_dff_A_UxntVVz47_2),.clk(gclk));
	jdff dff_A_N10FqqUo3_0(.dout(w_n196_0[0]),.din(w_dff_A_N10FqqUo3_0),.clk(gclk));
	jdff dff_B_FIeyk8Fz8_3(.din(n196),.dout(w_dff_B_FIeyk8Fz8_3),.clk(gclk));
	jdff dff_B_9FwPhw8Q1_3(.din(w_dff_B_FIeyk8Fz8_3),.dout(w_dff_B_9FwPhw8Q1_3),.clk(gclk));
	jdff dff_B_l4X8PHtZ6_3(.din(w_dff_B_9FwPhw8Q1_3),.dout(w_dff_B_l4X8PHtZ6_3),.clk(gclk));
	jdff dff_A_AvaVEbvT4_0(.dout(w_G179_2[0]),.din(w_dff_A_AvaVEbvT4_0),.clk(gclk));
	jdff dff_A_hKWWXyq27_0(.dout(w_dff_A_AvaVEbvT4_0),.din(w_dff_A_hKWWXyq27_0),.clk(gclk));
	jdff dff_A_ctNigOQu5_0(.dout(w_dff_A_hKWWXyq27_0),.din(w_dff_A_ctNigOQu5_0),.clk(gclk));
	jdff dff_A_Fc5aWhdd9_0(.dout(w_dff_A_ctNigOQu5_0),.din(w_dff_A_Fc5aWhdd9_0),.clk(gclk));
	jdff dff_A_BJplSB7a7_1(.dout(w_G179_2[1]),.din(w_dff_A_BJplSB7a7_1),.clk(gclk));
	jdff dff_A_o8gycTsf9_1(.dout(w_dff_A_BJplSB7a7_1),.din(w_dff_A_o8gycTsf9_1),.clk(gclk));
	jdff dff_A_CmiBshCD6_1(.dout(w_dff_A_o8gycTsf9_1),.din(w_dff_A_CmiBshCD6_1),.clk(gclk));
	jdff dff_A_OimBSSv70_1(.dout(w_dff_A_CmiBshCD6_1),.din(w_dff_A_OimBSSv70_1),.clk(gclk));
	jdff dff_A_1AsNcgwk6_0(.dout(w_G179_0[0]),.din(w_dff_A_1AsNcgwk6_0),.clk(gclk));
	jdff dff_A_XHYTYbR15_0(.dout(w_dff_A_1AsNcgwk6_0),.din(w_dff_A_XHYTYbR15_0),.clk(gclk));
	jdff dff_A_BROATec47_0(.dout(w_dff_A_XHYTYbR15_0),.din(w_dff_A_BROATec47_0),.clk(gclk));
	jdff dff_A_53Uc2rbS7_0(.dout(w_dff_A_BROATec47_0),.din(w_dff_A_53Uc2rbS7_0),.clk(gclk));
	jdff dff_B_BM9YOQ0C2_1(.din(n183),.dout(w_dff_B_BM9YOQ0C2_1),.clk(gclk));
	jdff dff_B_cL8Xs4078_1(.din(w_dff_B_BM9YOQ0C2_1),.dout(w_dff_B_cL8Xs4078_1),.clk(gclk));
	jdff dff_B_aCcUphpJ2_0(.din(n193),.dout(w_dff_B_aCcUphpJ2_0),.clk(gclk));
	jdff dff_B_j2zTilF61_0(.din(w_dff_B_aCcUphpJ2_0),.dout(w_dff_B_j2zTilF61_0),.clk(gclk));
	jdff dff_B_opaONvPE0_0(.din(n192),.dout(w_dff_B_opaONvPE0_0),.clk(gclk));
	jdff dff_A_m6CFZT0t9_1(.dout(w_n190_1[1]),.din(w_dff_A_m6CFZT0t9_1),.clk(gclk));
	jdff dff_A_gHqlsMsW1_1(.dout(w_dff_A_m6CFZT0t9_1),.din(w_dff_A_gHqlsMsW1_1),.clk(gclk));
	jdff dff_A_uXhuoCTd3_1(.dout(w_n189_0[1]),.din(w_dff_A_uXhuoCTd3_1),.clk(gclk));
	jdff dff_A_ss9i5BgQ2_2(.dout(w_n189_0[2]),.din(w_dff_A_ss9i5BgQ2_2),.clk(gclk));
	jdff dff_A_0p1AtjHg8_0(.dout(w_n85_0[0]),.din(w_dff_A_0p1AtjHg8_0),.clk(gclk));
	jdff dff_A_nCQ6NDQn7_0(.dout(w_dff_A_0p1AtjHg8_0),.din(w_dff_A_nCQ6NDQn7_0),.clk(gclk));
	jdff dff_A_hVNnjKgP6_2(.dout(w_n85_0[2]),.din(w_dff_A_hVNnjKgP6_2),.clk(gclk));
	jdff dff_A_RCUi5Vvx2_2(.dout(w_dff_A_hVNnjKgP6_2),.din(w_dff_A_RCUi5Vvx2_2),.clk(gclk));
	jdff dff_A_mKrXYaZq8_2(.dout(w_dff_A_RCUi5Vvx2_2),.din(w_dff_A_mKrXYaZq8_2),.clk(gclk));
	jdff dff_A_kzFWYfB52_0(.dout(w_G20_5[0]),.din(w_dff_A_kzFWYfB52_0),.clk(gclk));
	jdff dff_A_86qZ2guA2_1(.dout(w_G20_5[1]),.din(w_dff_A_86qZ2guA2_1),.clk(gclk));
	jdff dff_B_DVVSq78l4_1(.din(n176),.dout(w_dff_B_DVVSq78l4_1),.clk(gclk));
	jdff dff_A_AiFPZa8C2_1(.dout(w_n80_0[1]),.din(w_dff_A_AiFPZa8C2_1),.clk(gclk));
	jdff dff_A_xb1N1XZD3_1(.dout(w_dff_A_AiFPZa8C2_1),.din(w_dff_A_xb1N1XZD3_1),.clk(gclk));
	jdff dff_A_nQ70BLCU2_1(.dout(w_dff_A_xb1N1XZD3_1),.din(w_dff_A_nQ70BLCU2_1),.clk(gclk));
	jdff dff_A_LXJDY3TB2_2(.dout(w_n80_0[2]),.din(w_dff_A_LXJDY3TB2_2),.clk(gclk));
	jdff dff_A_8UVLIIqI1_2(.dout(w_dff_A_LXJDY3TB2_2),.din(w_dff_A_8UVLIIqI1_2),.clk(gclk));
	jdff dff_A_e7fhqZWt8_2(.dout(w_dff_A_8UVLIIqI1_2),.din(w_dff_A_e7fhqZWt8_2),.clk(gclk));
	jdff dff_A_4Koz7mTc1_2(.dout(w_G107_1[2]),.din(w_dff_A_4Koz7mTc1_2),.clk(gclk));
	jdff dff_A_rGidlNBb4_2(.dout(w_dff_A_4Koz7mTc1_2),.din(w_dff_A_rGidlNBb4_2),.clk(gclk));
	jdff dff_A_ucjKX2Ip8_2(.dout(w_dff_A_rGidlNBb4_2),.din(w_dff_A_ucjKX2Ip8_2),.clk(gclk));
	jdff dff_A_XOGi0qq44_1(.dout(w_G107_0[1]),.din(w_dff_A_XOGi0qq44_1),.clk(gclk));
	jdff dff_A_7DvbtkSk3_1(.dout(w_dff_A_XOGi0qq44_1),.din(w_dff_A_7DvbtkSk3_1),.clk(gclk));
	jdff dff_A_uVI7mBqD7_1(.dout(w_dff_A_7DvbtkSk3_1),.din(w_dff_A_uVI7mBqD7_1),.clk(gclk));
	jdff dff_A_kef2gZQk4_2(.dout(w_G107_0[2]),.din(w_dff_A_kef2gZQk4_2),.clk(gclk));
	jdff dff_A_osY162wu3_2(.dout(w_dff_A_kef2gZQk4_2),.din(w_dff_A_osY162wu3_2),.clk(gclk));
	jdff dff_A_dGUtwM5M9_2(.dout(w_dff_A_osY162wu3_2),.din(w_dff_A_dGUtwM5M9_2),.clk(gclk));
	jdff dff_A_e3ybj4k98_0(.dout(w_n79_0[0]),.din(w_dff_A_e3ybj4k98_0),.clk(gclk));
	jdff dff_A_G6UuLri30_0(.dout(w_dff_A_e3ybj4k98_0),.din(w_dff_A_G6UuLri30_0),.clk(gclk));
	jdff dff_A_yzUpWH5M6_0(.dout(w_G97_5[0]),.din(w_dff_A_yzUpWH5M6_0),.clk(gclk));
	jdff dff_A_4u2Un4vU5_1(.dout(w_n97_1[1]),.din(w_dff_A_4u2Un4vU5_1),.clk(gclk));
	jdff dff_A_yqm5Cmbs8_0(.dout(w_n97_0[0]),.din(w_dff_A_yqm5Cmbs8_0),.clk(gclk));
	jdff dff_A_6pRkK9FN2_0(.dout(w_G87_3[0]),.din(w_dff_A_6pRkK9FN2_0),.clk(gclk));
	jdff dff_A_ukR2nlQi9_2(.dout(w_G87_3[2]),.din(w_dff_A_ukR2nlQi9_2),.clk(gclk));
	jdff dff_A_tKUtTOmO6_2(.dout(w_dff_A_ukR2nlQi9_2),.din(w_dff_A_tKUtTOmO6_2),.clk(gclk));
	jdff dff_A_mWHgdEQc4_2(.dout(w_dff_A_tKUtTOmO6_2),.din(w_dff_A_mWHgdEQc4_2),.clk(gclk));
	jdff dff_A_vg2Y6Sze3_0(.dout(w_G87_0[0]),.din(w_dff_A_vg2Y6Sze3_0),.clk(gclk));
	jdff dff_A_uCTlBNek9_0(.dout(w_dff_A_vg2Y6Sze3_0),.din(w_dff_A_uCTlBNek9_0),.clk(gclk));
	jdff dff_A_FvwJAaIG2_0(.dout(w_dff_A_uCTlBNek9_0),.din(w_dff_A_FvwJAaIG2_0),.clk(gclk));
	jdff dff_A_zaqVxPXS5_0(.dout(w_n179_1[0]),.din(w_dff_A_zaqVxPXS5_0),.clk(gclk));
	jdff dff_A_yoPHyq905_2(.dout(w_n179_1[2]),.din(w_dff_A_yoPHyq905_2),.clk(gclk));
	jdff dff_A_0m7SaP7A3_2(.dout(w_dff_A_yoPHyq905_2),.din(w_dff_A_0m7SaP7A3_2),.clk(gclk));
	jdff dff_A_ayIycAJM7_1(.dout(w_n179_0[1]),.din(w_dff_A_ayIycAJM7_1),.clk(gclk));
	jdff dff_A_Dfp0TMCR9_1(.dout(w_dff_A_ayIycAJM7_1),.din(w_dff_A_Dfp0TMCR9_1),.clk(gclk));
	jdff dff_A_234SJcZS8_1(.dout(w_dff_A_Dfp0TMCR9_1),.din(w_dff_A_234SJcZS8_1),.clk(gclk));
	jdff dff_A_3Xzilur23_2(.dout(w_n179_0[2]),.din(w_dff_A_3Xzilur23_2),.clk(gclk));
	jdff dff_A_5FpVGYKY5_2(.dout(w_dff_A_3Xzilur23_2),.din(w_dff_A_5FpVGYKY5_2),.clk(gclk));
	jdff dff_A_zmKQObbx5_2(.dout(w_dff_A_5FpVGYKY5_2),.din(w_dff_A_zmKQObbx5_2),.clk(gclk));
	jdff dff_A_afzTHK3A5_2(.dout(w_dff_A_zmKQObbx5_2),.din(w_dff_A_afzTHK3A5_2),.clk(gclk));
	jdff dff_A_56JqZ5B84_1(.dout(w_G20_2[1]),.din(w_dff_A_56JqZ5B84_1),.clk(gclk));
	jdff dff_A_QT5SPFcM2_0(.dout(w_G68_4[0]),.din(w_dff_A_QT5SPFcM2_0),.clk(gclk));
	jdff dff_A_CO2XZcYU0_0(.dout(w_G68_1[0]),.din(w_dff_A_CO2XZcYU0_0),.clk(gclk));
	jdff dff_A_O8zT6EuW1_2(.dout(w_G68_1[2]),.din(w_dff_A_O8zT6EuW1_2),.clk(gclk));
	jdff dff_A_z8K8SKsH1_2(.dout(w_dff_A_O8zT6EuW1_2),.din(w_dff_A_z8K8SKsH1_2),.clk(gclk));
	jdff dff_A_hNy8bXX81_2(.dout(w_dff_A_z8K8SKsH1_2),.din(w_dff_A_hNy8bXX81_2),.clk(gclk));
	jdff dff_A_4WU1ylqH1_2(.dout(w_dff_A_hNy8bXX81_2),.din(w_dff_A_4WU1ylqH1_2),.clk(gclk));
	jdff dff_A_bLHzeMOq5_2(.dout(w_G68_0[2]),.din(w_dff_A_bLHzeMOq5_2),.clk(gclk));
	jdff dff_A_ssqYW7xV1_0(.dout(w_G20_6[0]),.din(w_dff_A_ssqYW7xV1_0),.clk(gclk));
	jdff dff_A_gWXHEB4g6_2(.dout(w_G20_1[2]),.din(w_dff_A_gWXHEB4g6_2),.clk(gclk));
	jdff dff_A_mzOzAUZf7_0(.dout(w_G20_0[0]),.din(w_dff_A_mzOzAUZf7_0),.clk(gclk));
	jdff dff_A_ttZt2BHE1_0(.dout(w_n172_0[0]),.din(w_dff_A_ttZt2BHE1_0),.clk(gclk));
	jdff dff_B_CJBybfjs7_2(.din(n172),.dout(w_dff_B_CJBybfjs7_2),.clk(gclk));
	jdff dff_A_HLumzEHt0_0(.dout(w_G97_4[0]),.din(w_dff_A_HLumzEHt0_0),.clk(gclk));
	jdff dff_A_Bni4SiGC5_0(.dout(w_dff_A_HLumzEHt0_0),.din(w_dff_A_Bni4SiGC5_0),.clk(gclk));
	jdff dff_A_dznUlpk64_0(.dout(w_dff_A_Bni4SiGC5_0),.din(w_dff_A_dznUlpk64_0),.clk(gclk));
	jdff dff_A_tCWyG7hq5_2(.dout(w_G97_1[2]),.din(w_dff_A_tCWyG7hq5_2),.clk(gclk));
	jdff dff_A_qHGWqIUO4_2(.dout(w_dff_A_tCWyG7hq5_2),.din(w_dff_A_qHGWqIUO4_2),.clk(gclk));
	jdff dff_A_qMdiEpKU1_2(.dout(w_dff_A_qHGWqIUO4_2),.din(w_dff_A_qMdiEpKU1_2),.clk(gclk));
	jdff dff_A_criETge50_2(.dout(w_dff_A_qMdiEpKU1_2),.din(w_dff_A_criETge50_2),.clk(gclk));
	jdff dff_A_5YazrCLb8_1(.dout(w_G97_0[1]),.din(w_dff_A_5YazrCLb8_1),.clk(gclk));
	jdff dff_A_fn6533Kk3_1(.dout(w_dff_A_5YazrCLb8_1),.din(w_dff_A_fn6533Kk3_1),.clk(gclk));
	jdff dff_A_GPRLNY7X4_1(.dout(w_dff_A_fn6533Kk3_1),.din(w_dff_A_GPRLNY7X4_1),.clk(gclk));
	jdff dff_A_C1VcRIZQ0_2(.dout(w_G97_0[2]),.din(w_dff_A_C1VcRIZQ0_2),.clk(gclk));
	jdff dff_A_krMXfSYv2_0(.dout(w_G33_10[0]),.din(w_dff_A_krMXfSYv2_0),.clk(gclk));
	jdff dff_A_YsH3D4I38_1(.dout(w_G33_10[1]),.din(w_dff_A_YsH3D4I38_1),.clk(gclk));
	jdff dff_A_UWPcFigi2_0(.dout(w_n170_0[0]),.din(w_dff_A_UWPcFigi2_0),.clk(gclk));
	jdff dff_B_EVEz00gg4_0(.din(n168),.dout(w_dff_B_EVEz00gg4_0),.clk(gclk));
	jdff dff_A_rZ2wUsBs6_0(.dout(w_G274_0[0]),.din(w_dff_A_rZ2wUsBs6_0),.clk(gclk));
	jdff dff_A_HiU1UimC1_2(.dout(w_G274_0[2]),.din(w_dff_A_HiU1UimC1_2),.clk(gclk));
	jdff dff_A_U5o5NzoL2_0(.dout(w_n166_3[0]),.din(w_dff_A_U5o5NzoL2_0),.clk(gclk));
	jdff dff_A_q5Q5q2co5_0(.dout(w_dff_A_U5o5NzoL2_0),.din(w_dff_A_q5Q5q2co5_0),.clk(gclk));
	jdff dff_A_a5XfqDH46_0(.dout(w_dff_A_q5Q5q2co5_0),.din(w_dff_A_a5XfqDH46_0),.clk(gclk));
	jdff dff_A_h2y9xBoJ6_0(.dout(w_n166_0[0]),.din(w_dff_A_h2y9xBoJ6_0),.clk(gclk));
	jdff dff_A_5b4c8wso7_1(.dout(w_n115_0[1]),.din(w_dff_A_5b4c8wso7_1),.clk(gclk));
	jdff dff_A_j7mMMThK7_1(.dout(w_n114_0[1]),.din(w_dff_A_j7mMMThK7_1),.clk(gclk));
	jdff dff_A_wFga1qG85_0(.dout(w_n163_0[0]),.din(w_dff_A_wFga1qG85_0),.clk(gclk));
	jdff dff_A_OLPawTs87_2(.dout(w_n161_0[2]),.din(w_dff_A_OLPawTs87_2),.clk(gclk));
	jdff dff_A_q7dzlngA8_2(.dout(w_dff_A_OLPawTs87_2),.din(w_dff_A_q7dzlngA8_2),.clk(gclk));
	jdff dff_A_3cucR8oQ9_2(.dout(w_dff_A_q7dzlngA8_2),.din(w_dff_A_3cucR8oQ9_2),.clk(gclk));
	jdff dff_A_0wn3i1iz8_0(.dout(w_G45_1[0]),.din(w_dff_A_0wn3i1iz8_0),.clk(gclk));
	jdff dff_A_TY2VhRBY5_0(.dout(w_dff_A_0wn3i1iz8_0),.din(w_dff_A_TY2VhRBY5_0),.clk(gclk));
	jdff dff_A_S7dmdcD61_1(.dout(w_G45_1[1]),.din(w_dff_A_S7dmdcD61_1),.clk(gclk));
	jdff dff_A_2kdKdgmT8_1(.dout(w_G45_0[1]),.din(w_dff_A_2kdKdgmT8_1),.clk(gclk));
	jdff dff_A_0bxmfvZ33_1(.dout(w_dff_A_2kdKdgmT8_1),.din(w_dff_A_0bxmfvZ33_1),.clk(gclk));
	jdff dff_A_npIB8IR04_1(.dout(w_dff_A_0bxmfvZ33_1),.din(w_dff_A_npIB8IR04_1),.clk(gclk));
	jdff dff_A_F27IqvPM3_2(.dout(w_G45_0[2]),.din(w_dff_A_F27IqvPM3_2),.clk(gclk));
	jdff dff_A_9sBnGlXU2_2(.dout(w_dff_A_F27IqvPM3_2),.din(w_dff_A_9sBnGlXU2_2),.clk(gclk));
	jdff dff_A_DJiarWZ95_2(.dout(w_dff_A_9sBnGlXU2_2),.din(w_dff_A_DJiarWZ95_2),.clk(gclk));
	jdff dff_A_lJhY60M69_0(.dout(w_G250_0[0]),.din(w_dff_A_lJhY60M69_0),.clk(gclk));
	jdff dff_A_J0qcyDa95_0(.dout(w_dff_A_lJhY60M69_0),.din(w_dff_A_J0qcyDa95_0),.clk(gclk));
	jdff dff_A_cQ5cFH192_1(.dout(w_G250_0[1]),.din(w_dff_A_cQ5cFH192_1),.clk(gclk));
	jdff dff_A_2UtXVpAi1_1(.dout(w_dff_A_cQ5cFH192_1),.din(w_dff_A_2UtXVpAi1_1),.clk(gclk));
	jdff dff_A_LmlS4BSt7_0(.dout(w_n157_0[0]),.din(w_dff_A_LmlS4BSt7_0),.clk(gclk));
	jdff dff_A_Xnnkyn8u5_2(.dout(w_n157_0[2]),.din(w_dff_A_Xnnkyn8u5_2),.clk(gclk));
	jdff dff_A_WEIuYqWf0_2(.dout(w_dff_A_Xnnkyn8u5_2),.din(w_dff_A_WEIuYqWf0_2),.clk(gclk));
	jdff dff_A_puhH3F2G7_1(.dout(w_G116_1[1]),.din(w_dff_A_puhH3F2G7_1),.clk(gclk));
	jdff dff_A_1XfGqOOE2_1(.dout(w_dff_A_puhH3F2G7_1),.din(w_dff_A_1XfGqOOE2_1),.clk(gclk));
	jdff dff_A_1JXlQGbO6_1(.dout(w_dff_A_1XfGqOOE2_1),.din(w_dff_A_1JXlQGbO6_1),.clk(gclk));
	jdff dff_A_L9B71FRG1_2(.dout(w_G116_1[2]),.din(w_dff_A_L9B71FRG1_2),.clk(gclk));
	jdff dff_A_VIHtJ1nh8_2(.dout(w_dff_A_L9B71FRG1_2),.din(w_dff_A_VIHtJ1nh8_2),.clk(gclk));
	jdff dff_A_uiWlur9c6_2(.dout(w_dff_A_VIHtJ1nh8_2),.din(w_dff_A_uiWlur9c6_2),.clk(gclk));
	jdff dff_A_1YvdgI3Y2_1(.dout(w_G116_0[1]),.din(w_dff_A_1YvdgI3Y2_1),.clk(gclk));
	jdff dff_A_MjRQy9tV0_1(.dout(w_dff_A_1YvdgI3Y2_1),.din(w_dff_A_MjRQy9tV0_1),.clk(gclk));
	jdff dff_A_W9EB8iqA1_1(.dout(w_dff_A_MjRQy9tV0_1),.din(w_dff_A_W9EB8iqA1_1),.clk(gclk));
	jdff dff_A_RRQhBpxU0_2(.dout(w_G116_0[2]),.din(w_dff_A_RRQhBpxU0_2),.clk(gclk));
	jdff dff_A_92PNDuK20_0(.dout(w_G238_1[0]),.din(w_dff_A_92PNDuK20_0),.clk(gclk));
	jdff dff_A_Yqz3Gn3v8_0(.dout(w_dff_A_92PNDuK20_0),.din(w_dff_A_Yqz3Gn3v8_0),.clk(gclk));
	jdff dff_A_fJLa1NaZ1_1(.dout(w_G238_0[1]),.din(w_dff_A_fJLa1NaZ1_1),.clk(gclk));
	jdff dff_A_G6UpWjIo9_1(.dout(w_dff_A_fJLa1NaZ1_1),.din(w_dff_A_G6UpWjIo9_1),.clk(gclk));
	jdff dff_A_i6QxGQVe1_1(.dout(w_dff_A_G6UpWjIo9_1),.din(w_dff_A_i6QxGQVe1_1),.clk(gclk));
	jdff dff_A_2v78RoHI8_2(.dout(w_G238_0[2]),.din(w_dff_A_2v78RoHI8_2),.clk(gclk));
	jdff dff_A_FsqTWjI07_2(.dout(w_dff_A_2v78RoHI8_2),.din(w_dff_A_FsqTWjI07_2),.clk(gclk));
	jdff dff_A_InfOy5b73_2(.dout(w_G1698_0[2]),.din(w_dff_A_InfOy5b73_2),.clk(gclk));
	jdff dff_A_PrLHja963_0(.dout(w_G244_1[0]),.din(w_dff_A_PrLHja963_0),.clk(gclk));
	jdff dff_A_tC83FC8o7_0(.dout(w_dff_A_PrLHja963_0),.din(w_dff_A_tC83FC8o7_0),.clk(gclk));
	jdff dff_A_qkXshSGn7_1(.dout(w_G244_0[1]),.din(w_dff_A_qkXshSGn7_1),.clk(gclk));
	jdff dff_A_JGhT6wNK3_1(.dout(w_dff_A_qkXshSGn7_1),.din(w_dff_A_JGhT6wNK3_1),.clk(gclk));
	jdff dff_A_SEmmsmwT0_1(.dout(w_dff_A_JGhT6wNK3_1),.din(w_dff_A_SEmmsmwT0_1),.clk(gclk));
	jdff dff_A_b5uT6m1p0_2(.dout(w_G244_0[2]),.din(w_dff_A_b5uT6m1p0_2),.clk(gclk));
	jdff dff_A_h8ARcq9S8_2(.dout(w_dff_A_b5uT6m1p0_2),.din(w_dff_A_h8ARcq9S8_2),.clk(gclk));
	jdff dff_A_Vmigz4lE8_1(.dout(w_n151_4[1]),.din(w_dff_A_Vmigz4lE8_1),.clk(gclk));
	jdff dff_A_iqj7eGhw3_2(.dout(w_n151_4[2]),.din(w_dff_A_iqj7eGhw3_2),.clk(gclk));
	jdff dff_A_ChjD05Oz7_1(.dout(w_n151_1[1]),.din(w_dff_A_ChjD05Oz7_1),.clk(gclk));
	jdff dff_A_klL2CcSO6_2(.dout(w_n151_1[2]),.din(w_dff_A_klL2CcSO6_2),.clk(gclk));
	jdff dff_A_2ThYXdQ06_1(.dout(w_n151_0[1]),.din(w_dff_A_2ThYXdQ06_1),.clk(gclk));
	jdff dff_A_tOq02BT72_2(.dout(w_n151_0[2]),.din(w_dff_A_tOq02BT72_2),.clk(gclk));
	jdff dff_A_Ofo02QnI0_0(.dout(w_n149_2[0]),.din(w_dff_A_Ofo02QnI0_0),.clk(gclk));
	jdff dff_A_8EkU4qhP9_1(.dout(w_G41_0[1]),.din(w_dff_A_8EkU4qhP9_1),.clk(gclk));
	jdff dff_A_XDkJrU828_2(.dout(w_G41_0[2]),.din(w_dff_A_XDkJrU828_2),.clk(gclk));
	jdff dff_A_d8SxFKtX6_2(.dout(w_G33_3[2]),.din(w_dff_A_d8SxFKtX6_2),.clk(gclk));
	jdff dff_A_glmJoVXE4_2(.dout(w_dff_A_d8SxFKtX6_2),.din(w_dff_A_glmJoVXE4_2),.clk(gclk));
	jdff dff_A_11ZkU7Ow7_2(.dout(w_dff_A_glmJoVXE4_2),.din(w_dff_A_11ZkU7Ow7_2),.clk(gclk));
	jdff dff_A_OJmdWQiM5_2(.dout(w_dff_A_11ZkU7Ow7_2),.din(w_dff_A_OJmdWQiM5_2),.clk(gclk));
	jdff dff_A_dPMt59dE4_0(.dout(w_G33_0[0]),.din(w_dff_A_dPMt59dE4_0),.clk(gclk));
	jdff dff_A_gjlubog67_1(.dout(w_n147_0[1]),.din(w_dff_A_gjlubog67_1),.clk(gclk));
	jdff dff_A_2PjEZTO05_1(.dout(w_G13_0[1]),.din(w_dff_A_2PjEZTO05_1),.clk(gclk));
	jdff dff_A_0CVfsRU63_2(.dout(w_G13_0[2]),.din(w_dff_A_0CVfsRU63_2),.clk(gclk));
	jdff dff_A_xLxPARyb1_2(.dout(w_dff_A_0CVfsRU63_2),.din(w_dff_A_xLxPARyb1_2),.clk(gclk));
	jdff dff_A_1hNsEnv72_0(.dout(w_G1_2[0]),.din(w_dff_A_1hNsEnv72_0),.clk(gclk));
	jdff dff_A_zKO6tXtJ2_2(.dout(w_G1_2[2]),.din(w_dff_A_zKO6tXtJ2_2),.clk(gclk));
	jdff dff_A_4ccyHmp11_0(.dout(w_G1_0[0]),.din(w_dff_A_4ccyHmp11_0),.clk(gclk));
	jdff dff_A_3DuuZRVa7_1(.dout(w_n146_3[1]),.din(w_dff_A_3DuuZRVa7_1),.clk(gclk));
	jdff dff_A_gVRr6fTO5_1(.dout(w_n146_0[1]),.din(w_dff_A_gVRr6fTO5_1),.clk(gclk));
	jdff dff_A_8OtG8urN5_1(.dout(w_dff_A_gVRr6fTO5_1),.din(w_dff_A_8OtG8urN5_1),.clk(gclk));
	jdff dff_A_ZUfJKdXR1_1(.dout(w_dff_A_8OtG8urN5_1),.din(w_dff_A_ZUfJKdXR1_1),.clk(gclk));
	jdff dff_A_BOalHFFR6_2(.dout(w_n146_0[2]),.din(w_dff_A_BOalHFFR6_2),.clk(gclk));
	jdff dff_A_UsWvRPmX7_2(.dout(w_dff_A_BOalHFFR6_2),.din(w_dff_A_UsWvRPmX7_2),.clk(gclk));
	jdff dff_A_IF5vSjQB9_2(.dout(w_dff_A_UsWvRPmX7_2),.din(w_dff_A_IF5vSjQB9_2),.clk(gclk));
	jdff dff_A_08fsOT2c1_0(.dout(w_G169_1[0]),.din(w_dff_A_08fsOT2c1_0),.clk(gclk));
	jdff dff_A_dZf0Wm7P0_0(.dout(w_dff_A_08fsOT2c1_0),.din(w_dff_A_dZf0Wm7P0_0),.clk(gclk));
	jdff dff_A_93DlXyxW7_0(.dout(w_dff_A_dZf0Wm7P0_0),.din(w_dff_A_93DlXyxW7_0),.clk(gclk));
	jdff dff_A_3oN4b9F83_0(.dout(w_dff_A_93DlXyxW7_0),.din(w_dff_A_3oN4b9F83_0),.clk(gclk));
	jdff dff_A_6uEwpP187_0(.dout(w_dff_A_3oN4b9F83_0),.din(w_dff_A_6uEwpP187_0),.clk(gclk));
	jdff dff_A_mDogEzEr3_1(.dout(w_G169_0[1]),.din(w_dff_A_mDogEzEr3_1),.clk(gclk));
	jdff dff_A_gutowc619_1(.dout(w_dff_A_mDogEzEr3_1),.din(w_dff_A_gutowc619_1),.clk(gclk));
	jdff dff_A_Grg7VoFW1_1(.dout(w_dff_A_gutowc619_1),.din(w_dff_A_Grg7VoFW1_1),.clk(gclk));
	jdff dff_A_sK7Q5PHe8_1(.dout(w_dff_A_Grg7VoFW1_1),.din(w_dff_A_sK7Q5PHe8_1),.clk(gclk));
	jdff dff_A_2Q8RLOiD5_2(.dout(w_G169_0[2]),.din(w_dff_A_2Q8RLOiD5_2),.clk(gclk));
	jdff dff_A_TifJx5L45_2(.dout(w_dff_A_2Q8RLOiD5_2),.din(w_dff_A_TifJx5L45_2),.clk(gclk));
	jdff dff_A_xmxtQFrp3_2(.dout(w_dff_A_TifJx5L45_2),.din(w_dff_A_xmxtQFrp3_2),.clk(gclk));
	jdff dff_A_kv2bcKv06_2(.dout(w_dff_A_xmxtQFrp3_2),.din(w_dff_A_kv2bcKv06_2),.clk(gclk));
	jdff dff_A_H15fiu2u7_2(.dout(w_dff_A_kv2bcKv06_2),.din(w_dff_A_H15fiu2u7_2),.clk(gclk));
endmodule

