/*

c880:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jdff: 781
	jand: 153
	jor: 119

Summary:
	jxor: 27
	jspl: 81
	jspl3: 92
	jnot: 42
	jdff: 781
	jand: 153
	jor: 119

The maximum logic level gap of any gate:
	c880: 5
*/

module rf_c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n101;
	wire n102;
	wire n103;
	wire n105;
	wire n106;
	wire n107;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n118;
	wire n119;
	wire n121;
	wire n122;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire[2:0] w_G1gat_0;
	wire[1:0] w_G1gat_1;
	wire[1:0] w_G8gat_0;
	wire[1:0] w_G13gat_0;
	wire[2:0] w_G17gat_0;
	wire[2:0] w_G17gat_1;
	wire[2:0] w_G17gat_2;
	wire[1:0] w_G26gat_0;
	wire[2:0] w_G29gat_0;
	wire[1:0] w_G36gat_0;
	wire[2:0] w_G42gat_0;
	wire[2:0] w_G42gat_1;
	wire[1:0] w_G42gat_2;
	wire[2:0] w_G51gat_0;
	wire[1:0] w_G51gat_1;
	wire[2:0] w_G55gat_0;
	wire[2:0] w_G59gat_0;
	wire[1:0] w_G59gat_1;
	wire[1:0] w_G68gat_0;
	wire[1:0] w_G75gat_0;
	wire[2:0] w_G80gat_0;
	wire[2:0] w_G91gat_0;
	wire[2:0] w_G96gat_0;
	wire[2:0] w_G101gat_0;
	wire[2:0] w_G106gat_0;
	wire[2:0] w_G111gat_0;
	wire[2:0] w_G116gat_0;
	wire[2:0] w_G121gat_0;
	wire[1:0] w_G126gat_0;
	wire[1:0] w_G130gat_0;
	wire[2:0] w_G138gat_0;
	wire[1:0] w_G138gat_1;
	wire[1:0] w_G143gat_0;
	wire[1:0] w_G146gat_0;
	wire[1:0] w_G149gat_0;
	wire[2:0] w_G153gat_0;
	wire[1:0] w_G156gat_0;
	wire[2:0] w_G159gat_0;
	wire[2:0] w_G159gat_1;
	wire[1:0] w_G159gat_2;
	wire[2:0] w_G165gat_0;
	wire[2:0] w_G165gat_1;
	wire[1:0] w_G165gat_2;
	wire[2:0] w_G171gat_0;
	wire[2:0] w_G171gat_1;
	wire[1:0] w_G171gat_2;
	wire[2:0] w_G177gat_0;
	wire[2:0] w_G177gat_1;
	wire[1:0] w_G177gat_2;
	wire[2:0] w_G183gat_0;
	wire[2:0] w_G183gat_1;
	wire[1:0] w_G183gat_2;
	wire[2:0] w_G189gat_0;
	wire[2:0] w_G189gat_1;
	wire[1:0] w_G189gat_2;
	wire[2:0] w_G195gat_0;
	wire[2:0] w_G195gat_1;
	wire[1:0] w_G195gat_2;
	wire[2:0] w_G201gat_0;
	wire[2:0] w_G201gat_1;
	wire[2:0] w_G201gat_2;
	wire[2:0] w_G210gat_0;
	wire[2:0] w_G210gat_1;
	wire[2:0] w_G210gat_2;
	wire[1:0] w_G210gat_3;
	wire[2:0] w_G219gat_0;
	wire[2:0] w_G219gat_1;
	wire[2:0] w_G219gat_2;
	wire[1:0] w_G219gat_3;
	wire[2:0] w_G228gat_0;
	wire[2:0] w_G228gat_1;
	wire[2:0] w_G228gat_2;
	wire[1:0] w_G228gat_3;
	wire[2:0] w_G237gat_0;
	wire[2:0] w_G237gat_1;
	wire[2:0] w_G237gat_2;
	wire[1:0] w_G237gat_3;
	wire[2:0] w_G246gat_0;
	wire[2:0] w_G246gat_1;
	wire[2:0] w_G246gat_2;
	wire[1:0] w_G246gat_3;
	wire[2:0] w_G255gat_0;
	wire[2:0] w_G261gat_0;
	wire[1:0] w_G268gat_0;
	wire[1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire[2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire[1:0] w_n86_0;
	wire[1:0] w_n88_0;
	wire[2:0] w_n92_0;
	wire[1:0] w_n93_0;
	wire[1:0] w_n96_0;
	wire[1:0] w_n98_0;
	wire[1:0] w_n99_0;
	wire[1:0] w_n101_0;
	wire[1:0] w_n102_0;
	wire[1:0] w_n106_0;
	wire[1:0] w_n107_0;
	wire[1:0] w_n111_0;
	wire[2:0] w_n118_0;
	wire[1:0] w_n121_0;
	wire[1:0] w_n143_0;
	wire[1:0] w_n149_0;
	wire[2:0] w_n153_0;
	wire[2:0] w_n153_1;
	wire[2:0] w_n153_2;
	wire[1:0] w_n153_3;
	wire[1:0] w_n154_0;
	wire[1:0] w_n157_0;
	wire[2:0] w_n159_0;
	wire[1:0] w_n159_1;
	wire[1:0] w_n162_0;
	wire[1:0] w_n163_0;
	wire[2:0] w_n165_0;
	wire[2:0] w_n165_1;
	wire[2:0] w_n167_0;
	wire[1:0] w_n167_1;
	wire[2:0] w_n168_0;
	wire[2:0] w_n181_0;
	wire[2:0] w_n181_1;
	wire[2:0] w_n181_2;
	wire[1:0] w_n181_3;
	wire[2:0] w_n193_0;
	wire[1:0] w_n193_1;
	wire[2:0] w_n194_0;
	wire[1:0] w_n196_0;
	wire[1:0] w_n213_0;
	wire[2:0] w_n217_0;
	wire[1:0] w_n217_1;
	wire[1:0] w_n218_0;
	wire[2:0] w_n222_0;
	wire[1:0] w_n222_1;
	wire[1:0] w_n223_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n228_0;
	wire[1:0] w_n230_0;
	wire[1:0] w_n232_0;
	wire[2:0] w_n236_0;
	wire[1:0] w_n238_0;
	wire[2:0] w_n252_0;
	wire[1:0] w_n255_0;
	wire[2:0] w_n273_0;
	wire[2:0] w_n292_0;
	wire[1:0] w_n292_1;
	wire[2:0] w_n296_0;
	wire[1:0] w_n296_1;
	wire[2:0] w_n299_0;
	wire[1:0] w_n299_1;
	wire[1:0] w_n302_0;
	wire[1:0] w_n303_0;
	wire[2:0] w_n305_0;
	wire[1:0] w_n305_1;
	wire[2:0] w_n312_0;
	wire[1:0] w_n312_1;
	wire[1:0] w_n315_0;
	wire[2:0] w_n321_0;
	wire[1:0] w_n321_1;
	wire[1:0] w_n322_0;
	wire[2:0] w_n328_0;
	wire[1:0] w_n328_1;
	wire[2:0] w_n329_0;
	wire[2:0] w_n330_0;
	wire[1:0] w_n331_0;
	wire[2:0] w_n335_0;
	wire[2:0] w_n337_0;
	wire[1:0] w_n339_0;
	wire[1:0] w_n340_0;
	wire[2:0] w_n346_0;
	wire[1:0] w_n346_1;
	wire[2:0] w_n347_0;
	wire[2:0] w_n367_0;
	wire[2:0] w_n383_0;
	wire[2:0] w_n405_0;
	wire w_dff_B_rcdGIbcJ4_2;
	wire w_dff_B_tiKX16Px0_1;
	wire w_dff_B_e4pn1wKp5_1;
	wire w_dff_A_VbzBPUP40_1;
	wire w_dff_B_TXvRpIgY2_0;
	wire w_dff_B_IhX0KD3f3_1;
	wire w_dff_B_KRLc3MAG8_0;
	wire w_dff_B_enXRNkZg0_0;
	wire w_dff_B_Owi7afwE7_0;
	wire w_dff_B_OHVPmDnQ5_0;
	wire w_dff_B_Nvw7oXI35_0;
	wire w_dff_B_z3ubSxCI4_0;
	wire w_dff_B_HhNG3CKU3_0;
	wire w_dff_B_USfRZPqj1_0;
	wire w_dff_B_AmGWvrWg3_0;
	wire w_dff_B_6vZlHYDc3_0;
	wire w_dff_B_lVb7JkCh4_0;
	wire w_dff_B_ablkYAcJ7_0;
	wire w_dff_B_2tF9mHCD8_0;
	wire w_dff_B_aF4hJVaf0_0;
	wire w_dff_B_Ts0mu9dQ2_0;
	wire w_dff_B_OBt1jgVH8_0;
	wire w_dff_B_LSU65Vw94_0;
	wire w_dff_B_IfUvKnRA3_0;
	wire w_dff_B_e89rPMCW6_0;
	wire w_dff_B_oXLMxhMh5_0;
	wire w_dff_B_EbYTPf9d3_0;
	wire w_dff_B_YqIEs0iB3_0;
	wire w_dff_B_fZttj8oE1_0;
	wire w_dff_B_b07EYonu0_0;
	wire w_dff_A_w1Bf2Yr52_0;
	wire w_dff_A_NVPALc7q9_0;
	wire w_dff_A_6dCSBIm63_0;
	wire w_dff_A_8KFNZSZn2_0;
	wire w_dff_B_TbHt2NqS5_1;
	wire w_dff_B_NPWf3BlC9_1;
	wire w_dff_B_6ntJpehm7_1;
	wire w_dff_B_BYdBkM1K9_1;
	wire w_dff_A_bfFYFjT90_1;
	wire w_dff_A_va8DJXVj6_1;
	wire w_dff_A_nL852zRF6_1;
	wire w_dff_A_lZsuws234_1;
	wire w_dff_B_I9MtPv5B2_0;
	wire w_dff_B_aRKeSmgl0_0;
	wire w_dff_B_LGC1z6e52_0;
	wire w_dff_B_OqDX1mhE5_0;
	wire w_dff_B_JUgQGpSK3_0;
	wire w_dff_B_3PkoWrj11_0;
	wire w_dff_B_GiAlbKGp3_0;
	wire w_dff_B_rOr14aHw5_0;
	wire w_dff_B_dY8HKWI11_0;
	wire w_dff_B_tnMSyusZ3_0;
	wire w_dff_B_UlJzRGsu9_0;
	wire w_dff_B_uQZJAPKj9_0;
	wire w_dff_B_AeskRH0b2_0;
	wire w_dff_B_Ao5ed7Sc2_0;
	wire w_dff_B_3rQfalH84_1;
	wire w_dff_B_NQ4RqetA0_1;
	wire w_dff_B_hbzpXksv7_1;
	wire w_dff_B_foePtHae1_1;
	wire w_dff_A_J2nYIFC01_1;
	wire w_dff_A_LsLfIUFq4_1;
	wire w_dff_A_aE2wYgBZ6_1;
	wire w_dff_A_9h2QmdbG4_1;
	wire w_dff_B_uQ49Dq5p5_0;
	wire w_dff_B_M1Ue3DhB0_0;
	wire w_dff_B_1zNYJEzd3_0;
	wire w_dff_B_QkcrlfEn9_0;
	wire w_dff_B_Lt1awlyo1_0;
	wire w_dff_B_m1dfGMgx5_0;
	wire w_dff_B_jiMhpmyk4_0;
	wire w_dff_B_MtZimH5r2_0;
	wire w_dff_B_A0BDc1nC7_0;
	wire w_dff_B_g681Yg8Y3_0;
	wire w_dff_B_I9IJunoj5_0;
	wire w_dff_B_ldOh7XXr3_0;
	wire w_dff_B_P392CBsC1_0;
	wire w_dff_B_aXzCb0vT9_0;
	wire w_dff_A_xEbT2sl02_1;
	wire w_dff_A_5y9cMeqJ6_1;
	wire w_dff_B_PSsVC57p9_1;
	wire w_dff_B_wQUoV3cU7_1;
	wire w_dff_B_lylyPlAQ1_1;
	wire w_dff_B_j70V6Zra1_1;
	wire w_dff_B_iXPshyrT5_1;
	wire w_dff_B_pXv7gpGb6_1;
	wire w_dff_B_T1LxtHyp1_1;
	wire w_dff_B_4CsWXpvl2_1;
	wire w_dff_B_9SCzL1PZ3_1;
	wire w_dff_B_fePUdM2d9_1;
	wire w_dff_B_R5eBDsPA3_1;
	wire w_dff_B_Vd93AqSE0_1;
	wire w_dff_B_Q0SXByaK0_1;
	wire w_dff_B_U89kJPZY4_1;
	wire w_dff_B_vj6QkmWj3_1;
	wire w_dff_B_4wOsKy8P0_1;
	wire w_dff_B_ue63feuJ8_1;
	wire w_dff_B_URtzJv2O8_1;
	wire w_dff_B_JqCAedvZ7_1;
	wire w_dff_B_UUujBUAM7_0;
	wire w_dff_B_cGkE6gFN0_0;
	wire w_dff_B_IN4gHvf12_0;
	wire w_dff_B_p39H8VW78_0;
	wire w_dff_B_vqWrTDug0_0;
	wire w_dff_B_PWPeztSQ1_0;
	wire w_dff_B_vhlg5ahJ8_0;
	wire w_dff_B_VGeWtE5A5_0;
	wire w_dff_B_JKAPmDKw7_0;
	wire w_dff_B_F5qxVQDB4_0;
	wire w_dff_B_T5cTBSeb9_0;
	wire w_dff_B_1BZcYoJP2_0;
	wire w_dff_B_CUK6ySF87_0;
	wire w_dff_B_QX469E8X6_0;
	wire w_dff_B_KFCGK5jy3_0;
	wire w_dff_A_luHCqTH56_1;
	wire w_dff_A_2q7bebE30_2;
	wire w_dff_A_VrnR1Axb8_0;
	wire w_dff_A_RBJldML08_0;
	wire w_dff_A_XsGDrWzE2_0;
	wire w_dff_A_CcZfl3DE9_0;
	wire w_dff_A_O4BnKZWH7_2;
	wire w_dff_A_TjZN6dMJ0_2;
	wire w_dff_B_PvelPzH93_0;
	wire w_dff_B_Cmgrk6HO6_0;
	wire w_dff_B_OVo8ApWz2_0;
	wire w_dff_B_NJi8DAPx1_0;
	wire w_dff_B_aMUOQhrM9_0;
	wire w_dff_B_BHvrKp0m4_0;
	wire w_dff_B_xzkYETx73_0;
	wire w_dff_A_3c1Tgmvu1_1;
	wire w_dff_A_1UTP8PLS0_1;
	wire w_dff_A_jncO0Wt77_1;
	wire w_dff_A_jkoQySE98_1;
	wire w_dff_A_Rxk9jG7z0_1;
	wire w_dff_A_o42z7cOD5_1;
	wire w_dff_A_fEwDBsn05_1;
	wire w_dff_B_ejuXkCzL1_0;
	wire w_dff_B_bKiJwjb46_0;
	wire w_dff_B_Q5z9qhIY4_0;
	wire w_dff_B_YNtbvHhX4_0;
	wire w_dff_B_vmSlP96T3_0;
	wire w_dff_B_2lmFNbKq1_0;
	wire w_dff_B_qcIiTrxY9_0;
	wire w_dff_B_XFRitF935_0;
	wire w_dff_B_bg76ZjFb0_0;
	wire w_dff_B_MP1MsEYv0_0;
	wire w_dff_B_svDJdJhT9_0;
	wire w_dff_B_m7emHeOP8_0;
	wire w_dff_B_ojYVdEt22_0;
	wire w_dff_B_eiDEt4M17_0;
	wire w_dff_B_EMEVQT7L2_0;
	wire w_dff_B_UDtgVnD31_0;
	wire w_dff_B_LpRmIxIQ1_0;
	wire w_dff_B_vZN3HOEM1_0;
	wire w_dff_B_2Xlx1w636_0;
	wire w_dff_B_6WjvhTfD9_0;
	wire w_dff_B_fvLSBqNQ5_0;
	wire w_dff_B_7hexCDOk7_0;
	wire w_dff_B_lCNVQeRg1_0;
	wire w_dff_B_4yYzpzQZ0_0;
	wire w_dff_B_yhPNafJe5_0;
	wire w_dff_B_eYxYzzQE9_0;
	wire w_dff_A_GrfYJCiC2_1;
	wire w_dff_A_dLR0ShHf5_1;
	wire w_dff_A_1rqDsFLz1_1;
	wire w_dff_A_oW93ECL87_1;
	wire w_dff_A_T43GN7ZP0_1;
	wire w_dff_A_C6VHNfKB4_1;
	wire w_dff_A_BWmG1Y5r6_1;
	wire w_dff_A_ekYEzkko1_1;
	wire w_dff_A_kL7E0WFL2_1;
	wire w_dff_B_y8wriyGN7_1;
	wire w_dff_B_gfoMCJij6_1;
	wire w_dff_B_9P1KBs8x2_1;
	wire w_dff_B_upwepf7Q2_0;
	wire w_dff_B_eRVd6BN99_0;
	wire w_dff_B_Eme59DSZ0_0;
	wire w_dff_B_Mf8HV2vp2_0;
	wire w_dff_A_hVABhXPc1_1;
	wire w_dff_A_vyIiVjNM8_1;
	wire w_dff_A_solfsl5g8_1;
	wire w_dff_A_ZHpQrXdH1_1;
	wire w_dff_B_uubR0MUS1_1;
	wire w_dff_B_ML0mMVFQ9_1;
	wire w_dff_B_alhlfcJh7_1;
	wire w_dff_B_P7J20owu5_0;
	wire w_dff_B_eQtQQ3Um4_0;
	wire w_dff_B_DRLhDGWM8_0;
	wire w_dff_B_gdY9OzYR7_0;
	wire w_dff_A_qFlBrBPR0_1;
	wire w_dff_A_4VrBza8N0_1;
	wire w_dff_A_xwMSUpzW4_1;
	wire w_dff_A_L4YyDJsW5_1;
	wire w_dff_B_VfiQu5VF8_1;
	wire w_dff_B_vuEUIjCo5_1;
	wire w_dff_B_isoGcj515_1;
	wire w_dff_B_qrL2tGue6_1;
	wire w_dff_B_SwdrMDr66_1;
	wire w_dff_B_UkOoVVom8_1;
	wire w_dff_B_2AmxpU0q8_1;
	wire w_dff_B_hwq3fEWR7_0;
	wire w_dff_B_PHn4Iqm46_0;
	wire w_dff_B_n4kuRFsg9_0;
	wire w_dff_B_kmGwrkYe2_0;
	wire w_dff_B_ccCIEoik0_0;
	wire w_dff_B_mWTTLcnW4_0;
	wire w_dff_B_nVWtyN8D2_0;
	wire w_dff_B_S0Dezss19_0;
	wire w_dff_B_PrfmrOam4_0;
	wire w_dff_B_JZYJZQ1Q8_0;
	wire w_dff_B_yIxaJxKJ8_0;
	wire w_dff_B_3BozDWWg7_0;
	wire w_dff_B_b9FJPlqP8_0;
	wire w_dff_B_YN5GQ3cq7_0;
	wire w_dff_B_mFMOqZYj2_0;
	wire w_dff_B_AJSJfjBV2_0;
	wire w_dff_B_ABwgDkzj8_0;
	wire w_dff_B_Hu4cH0Rk2_1;
	wire w_dff_B_fon8S6i46_1;
	wire w_dff_B_PpU2OFFW9_1;
	wire w_dff_B_e1SyOF1o5_1;
	wire w_dff_B_bNLJoKfB2_1;
	wire w_dff_B_cmLMnqV32_1;
	wire w_dff_B_T59eWlDD7_1;
	wire w_dff_B_fI27sppI3_1;
	wire w_dff_B_gYOXGW2O2_1;
	wire w_dff_B_bSf97WbI8_1;
	wire w_dff_B_r0hEydaL2_1;
	wire w_dff_B_IuBiekTt3_1;
	wire w_dff_B_8NxEq6dq0_1;
	wire w_dff_B_Xed15cmI5_1;
	wire w_dff_B_1pNGs2sO1_1;
	wire w_dff_B_j2CIVh7K0_0;
	wire w_dff_B_2HDtAj3D3_0;
	wire w_dff_B_FREj439S2_0;
	wire w_dff_B_mltqWTru1_0;
	wire w_dff_B_LCW2ZACj5_0;
	wire w_dff_B_2kkwxVAz8_0;
	wire w_dff_A_CJMAzMeI6_0;
	wire w_dff_A_7S7PtQTf3_0;
	wire w_dff_A_VZb0BmbH8_0;
	wire w_dff_A_p6whfGDb1_0;
	wire w_dff_A_zAVijECk6_0;
	wire w_dff_A_fJznWadX8_0;
	wire w_dff_A_Zqdv1tL21_2;
	wire w_dff_A_PX2pQ23d1_0;
	wire w_dff_A_6xDU2RAL3_0;
	wire w_dff_A_mIMn5Ykv7_0;
	wire w_dff_A_i2NJ4g9z3_0;
	wire w_dff_A_4QpLVSIA6_0;
	wire w_dff_A_W2JSlw2h6_0;
	wire w_dff_B_G0UghCva0_1;
	wire w_dff_A_1HZBh8Na0_1;
	wire w_dff_A_6iWupodD4_1;
	wire w_dff_A_yGMIvI1r9_1;
	wire w_dff_A_5KNnb36o7_1;
	wire w_dff_A_tOGmhFl81_1;
	wire w_dff_A_t5U60hl49_1;
	wire w_dff_A_DldUsMtM4_1;
	wire w_dff_A_PBhRjxzY1_1;
	wire w_dff_A_YRxUrohg1_1;
	wire w_dff_B_DK7amLpv3_0;
	wire w_dff_B_WgmeGV823_0;
	wire w_dff_B_G5GWcALe2_0;
	wire w_dff_B_56rvIfWm8_0;
	wire w_dff_B_AuPtzbiz8_0;
	wire w_dff_B_Dzq5giEZ1_0;
	wire w_dff_B_CUU6JaBF5_0;
	wire w_dff_B_WflL3jgp8_0;
	wire w_dff_B_8s6KdjQ07_0;
	wire w_dff_B_VibIDv318_0;
	wire w_dff_B_xS3NSyC90_0;
	wire w_dff_B_FdZQ15pz5_0;
	wire w_dff_B_eLkANbUv5_0;
	wire w_dff_B_UPm6L9Nb8_0;
	wire w_dff_B_YkSpfOp92_0;
	wire w_dff_B_vJbsKFLG4_0;
	wire w_dff_B_vYiQ7NLk9_0;
	wire w_dff_B_V0vRGvgv4_0;
	wire w_dff_B_zOsGNssi7_0;
	wire w_dff_B_YpYObPOD1_0;
	wire w_dff_A_2iPPdsSE7_2;
	wire w_dff_B_zwgj93p76_3;
	wire w_dff_B_PFAMbxko0_3;
	wire w_dff_B_MlU0lAIp0_3;
	wire w_dff_B_GIhP74Wg6_3;
	wire w_dff_B_pRq8GCv18_3;
	wire w_dff_B_UpjKneK80_3;
	wire w_dff_B_UJIi8sLE4_3;
	wire w_dff_B_OJh4kz4m2_3;
	wire w_dff_A_Jr3fhXse1_0;
	wire w_dff_A_Vlh8o8fC9_0;
	wire w_dff_A_Qa9NDiWx3_0;
	wire w_dff_A_WmBEmp6c2_0;
	wire w_dff_A_dF3Xy1lW9_0;
	wire w_dff_A_T72zKEQs2_0;
	wire w_dff_A_1HEjBh4a1_0;
	wire w_dff_A_abCT3wmx7_0;
	wire w_dff_A_X5vUCZ1M2_1;
	wire w_dff_A_PKbnaw7G5_1;
	wire w_dff_B_iQVI2BKV5_3;
	wire w_dff_B_iMK9Mlu16_3;
	wire w_dff_B_kW14EWci6_3;
	wire w_dff_B_8Ndi1Zxq2_3;
	wire w_dff_B_E0elwhjG7_3;
	wire w_dff_B_6UNO9qem1_3;
	wire w_dff_B_tbx6iKZj6_3;
	wire w_dff_B_83iLidIz6_3;
	wire w_dff_B_euJtAYGL1_3;
	wire w_dff_B_crlZpAfE1_3;
	wire w_dff_B_rKiurHBS4_1;
	wire w_dff_B_9RCMHPBu0_1;
	wire w_dff_B_RPZmQoZr1_1;
	wire w_dff_B_GXLj3m6L1_1;
	wire w_dff_B_qqUZXOxh3_1;
	wire w_dff_B_8CjKssne5_1;
	wire w_dff_B_EG4wx0MW6_1;
	wire w_dff_B_9yVDhpBE8_1;
	wire w_dff_B_fAWAZmko4_1;
	wire w_dff_B_vNRUB94I4_1;
	wire w_dff_B_lleVSr7Z3_1;
	wire w_dff_B_PnvaJQoS7_1;
	wire w_dff_B_TkBfJ3cD3_1;
	wire w_dff_B_pK3Xx1Um6_1;
	wire w_dff_B_2mhOtTAv5_1;
	wire w_dff_B_YDpaFihz6_1;
	wire w_dff_B_iwS0WEyB8_1;
	wire w_dff_B_oOj2Bofp5_0;
	wire w_dff_B_bMtc4hSB2_0;
	wire w_dff_B_2Wlz6Qyp1_0;
	wire w_dff_B_FNv6dQcA5_0;
	wire w_dff_B_7ByjNhWa2_0;
	wire w_dff_B_iPAFNaLz0_0;
	wire w_dff_B_H7X158O22_0;
	wire w_dff_A_bIRNQoO69_0;
	wire w_dff_A_lqDPTkFj9_0;
	wire w_dff_A_hym8EBkO5_0;
	wire w_dff_A_wiOTDdMU4_0;
	wire w_dff_A_UAmYFGzt6_0;
	wire w_dff_A_BRY6iDHA5_0;
	wire w_dff_A_0Pnsip6t7_0;
	wire w_dff_B_wDYsnYMr6_1;
	wire w_dff_B_l2eRCyw20_1;
	wire w_dff_B_hTzLZthE4_1;
	wire w_dff_B_mcSFyEiD8_1;
	wire w_dff_B_XPX9zK4e7_1;
	wire w_dff_B_H6xxC1vQ8_1;
	wire w_dff_B_nojOaqla9_1;
	wire w_dff_B_NTnOmrvD6_1;
	wire w_dff_B_e3KOWU6d5_1;
	wire w_dff_B_tOdDF97N7_0;
	wire w_dff_A_c7Ea73oJ2_0;
	wire w_dff_B_h7p1nVAO5_1;
	wire w_dff_A_SiQESX4O6_0;
	wire w_dff_A_UpHqMox65_0;
	wire w_dff_A_mZPGkEJ34_0;
	wire w_dff_B_5bvhS0zr2_0;
	wire w_dff_A_d7IZQ9Sj4_0;
	wire w_dff_A_duOlf6nd3_0;
	wire w_dff_A_kkq4hYOp2_0;
	wire w_dff_B_RbD4gjqX9_1;
	wire w_dff_B_vLsphLcm4_1;
	wire w_dff_A_PLo5IAVx8_1;
	wire w_dff_B_aC6KNLd33_2;
	wire w_dff_B_gRcQL1DW6_2;
	wire w_dff_B_HVnYHxUt3_2;
	wire w_dff_B_w4396kB92_2;
	wire w_dff_B_Wdi97rtg3_1;
	wire w_dff_B_lqDVT3hF7_1;
	wire w_dff_B_vqBT7hkr8_1;
	wire w_dff_B_zNfywTMl3_1;
	wire w_dff_B_kowgTTZz9_1;
	wire w_dff_B_Ol54VBa21_1;
	wire w_dff_B_v8lsR8PJ8_1;
	wire w_dff_B_6bYBhQ8m1_1;
	wire w_dff_B_Cy5q0l5Q0_1;
	wire w_dff_B_00CMSlPU3_1;
	wire w_dff_B_EYIGmiwN3_0;
	wire w_dff_B_JX4ZO1KH1_0;
	wire w_dff_B_F4gDpcuX1_2;
	wire w_dff_B_6DhNYeSz7_2;
	wire w_dff_B_vMrHShPs0_2;
	wire w_dff_B_cEECPJF44_2;
	wire w_dff_B_1VoLqFOE1_2;
	wire w_dff_B_N5SRkjjz3_2;
	wire w_dff_B_eja3Zprr7_2;
	wire w_dff_B_9vwFIlb01_2;
	wire w_dff_B_cvM5anir9_2;
	wire w_dff_A_IqsW8ezY1_0;
	wire w_dff_A_opLtEpGM9_1;
	wire w_dff_A_SFxqKb714_1;
	wire w_dff_A_tG4Nq4tb6_1;
	wire w_dff_A_onlv1ElE5_1;
	wire w_dff_A_4QIIxiCh7_1;
	wire w_dff_A_pIASlKGO9_1;
	wire w_dff_A_EJErUeDG7_1;
	wire w_dff_A_tgJgbBm83_1;
	wire w_dff_A_FagwKQkI8_1;
	wire w_dff_A_DxIJJiKv9_1;
	wire w_dff_B_7LyFN7op3_1;
	wire w_dff_A_ZiT1WcL60_1;
	wire w_dff_A_XmYDxrZe7_1;
	wire w_dff_A_pGAtQyKd6_2;
	wire w_dff_A_AMWZ37Nv6_2;
	wire w_dff_A_sdFNJJ7Q5_1;
	wire w_dff_A_3Sp17NIj4_1;
	wire w_dff_A_kApIzi8Z9_2;
	wire w_dff_A_7kPryKTi9_2;
	wire w_dff_B_mUBMt6NB3_0;
	wire w_dff_A_C2Hev3HG1_1;
	wire w_dff_B_ti8FtAkU0_2;
	wire w_dff_B_mJXsWUe91_2;
	wire w_dff_B_ECMNNrAZ5_2;
	wire w_dff_B_5FCgSxWW5_2;
	wire w_dff_A_610Oumgu4_0;
	wire w_dff_A_Y3OHDiIv6_0;
	wire w_dff_A_tohiyxjx3_0;
	wire w_dff_A_RwO6VadG0_0;
	wire w_dff_A_10I71eYm2_0;
	wire w_dff_A_SkXC7s7y6_0;
	wire w_dff_A_LavkY5SI2_0;
	wire w_dff_A_kpotA8MX8_0;
	wire w_dff_B_qRg2ss9o7_0;
	wire w_dff_B_l32VDpjh5_0;
	wire w_dff_B_DLghQFNe1_0;
	wire w_dff_A_wVds7YOW6_1;
	wire w_dff_A_omLyDlCE5_1;
	wire w_dff_A_Yqer7f1Z9_1;
	wire w_dff_A_2Mmiek4i6_1;
	wire w_dff_A_Yk8tPvBx2_1;
	wire w_dff_A_pmkPh0bg4_1;
	wire w_dff_A_6DpZ3zki6_1;
	wire w_dff_A_Ufn7cS606_1;
	wire w_dff_A_TyLlz1ve1_1;
	wire w_dff_B_eCkkmDWn5_0;
	wire w_dff_B_f3GLSOQR9_0;
	wire w_dff_B_lPbYyXpM1_0;
	wire w_dff_B_y0MrhwVI7_0;
	wire w_dff_A_xfZ43KYV4_1;
	wire w_dff_B_JrSDgxZO4_2;
	wire w_dff_B_tqwvZllI5_2;
	wire w_dff_B_h1lEKOyn7_2;
	wire w_dff_B_HZ81dAzI8_2;
	wire w_dff_B_zoCoK8vb1_0;
	wire w_dff_A_12pK7KFc3_2;
	wire w_dff_A_Nveud2mb4_0;
	wire w_dff_A_xoZZ7Jkz7_0;
	wire w_dff_A_Zg9LcbsT3_0;
	wire w_dff_A_QlZpgouh9_0;
	wire w_dff_A_HNUFoqL81_0;
	wire w_dff_A_rrYcQ1I47_0;
	wire w_dff_A_gKljUF238_0;
	wire w_dff_A_IwEWevRP9_0;
	wire w_dff_A_kVEtRdgL9_0;
	wire w_dff_A_nwyhWHvG0_0;
	wire w_dff_A_7M2Y2uWs8_0;
	wire w_dff_A_iGPJBw3f6_0;
	wire w_dff_A_sgUhCVAf1_0;
	wire w_dff_A_3s5spF6g2_0;
	wire w_dff_A_vQYkxVWn0_0;
	wire w_dff_A_Mz7EY8u92_0;
	wire w_dff_A_XRaOVevl0_0;
	wire w_dff_A_YKEeeP0I3_0;
	wire w_dff_A_FYUoAM6L3_2;
	wire w_dff_A_ogZ22fll2_0;
	wire w_dff_A_7UWG0EaP4_0;
	wire w_dff_A_meZ70Nsa8_0;
	wire w_dff_A_vKDZbclY4_0;
	wire w_dff_A_5K1rvWm95_0;
	wire w_dff_A_3I0AGCyS6_0;
	wire w_dff_A_lAuTnL480_0;
	wire w_dff_A_8POfUgPe4_0;
	wire w_dff_A_xxSUZAv19_0;
	wire w_dff_A_ZOicGVPq3_0;
	wire w_dff_A_UqHiV6yw3_0;
	wire w_dff_A_yBosPtPM2_0;
	wire w_dff_A_4caEvDFc9_0;
	wire w_dff_A_3lIBw1P08_0;
	wire w_dff_A_EiHRece77_0;
	wire w_dff_A_DOr5tNY45_0;
	wire w_dff_A_3s61wg1Z0_0;
	wire w_dff_A_H1Mx3OzL2_0;
	wire w_dff_A_EHSzjLlc3_2;
	wire w_dff_A_CHgW6rD36_0;
	wire w_dff_A_WKZJB1pK8_0;
	wire w_dff_A_zwvz0RKX7_0;
	wire w_dff_A_6emzrazG6_0;
	wire w_dff_A_yMYXFCny4_0;
	wire w_dff_A_luCt5MGJ7_0;
	wire w_dff_A_iWBGAb963_0;
	wire w_dff_A_7K20HTUv0_0;
	wire w_dff_A_DR3qcy2o0_0;
	wire w_dff_A_3wc6nGDp3_0;
	wire w_dff_A_d0oS4S9Y3_0;
	wire w_dff_A_fsMYUN2z0_0;
	wire w_dff_A_RxFQS75U2_0;
	wire w_dff_A_Urzsjl4R9_0;
	wire w_dff_A_yKYK3RC75_0;
	wire w_dff_A_eT5arAwv6_0;
	wire w_dff_A_eGguc1PC8_0;
	wire w_dff_A_QsWLzBPp5_0;
	wire w_dff_A_ZCq0xqL09_2;
	wire w_dff_A_OX7zotRu9_0;
	wire w_dff_A_7B1SBpp09_0;
	wire w_dff_A_8eKlMoEv8_0;
	wire w_dff_A_tucDdLNP2_0;
	wire w_dff_A_MAIFzxIl4_0;
	wire w_dff_A_zkYMUutu2_0;
	wire w_dff_A_BmAIfwi21_0;
	wire w_dff_A_JxEO3Ebr1_0;
	wire w_dff_A_twuc0zMm3_0;
	wire w_dff_A_bAFBj0FT7_0;
	wire w_dff_A_QUul71P98_0;
	wire w_dff_A_PmtXLCV48_0;
	wire w_dff_A_ZSPijMuI7_0;
	wire w_dff_A_vmuLVgYq7_0;
	wire w_dff_A_Jb0My8Pv7_0;
	wire w_dff_A_9RpbWCG31_0;
	wire w_dff_A_mrxqTp7K4_0;
	wire w_dff_A_8ESfrLvh2_0;
	wire w_dff_A_QxF9Ckid9_0;
	wire w_dff_A_sp5SF7qA2_2;
	wire w_dff_A_Up6sy3FS0_0;
	wire w_dff_A_uaI8ct1b1_0;
	wire w_dff_A_oD9tbUIl9_0;
	wire w_dff_A_pITwVpZq7_0;
	wire w_dff_A_9jR9Icnk1_0;
	wire w_dff_A_2ShS7tyM6_0;
	wire w_dff_A_hJcR9PoC8_0;
	wire w_dff_A_r5vxBedS4_0;
	wire w_dff_A_dxIJo9643_0;
	wire w_dff_A_SfiwhXMv5_0;
	wire w_dff_A_ulpUGvSQ9_0;
	wire w_dff_A_dhBdF6Sx1_0;
	wire w_dff_A_xTSljTPF5_0;
	wire w_dff_A_ngUQHmGZ0_0;
	wire w_dff_A_3ZSrSQEb4_0;
	wire w_dff_A_F5dugAzX6_0;
	wire w_dff_A_tclHPkqb7_0;
	wire w_dff_A_3joSsVwd5_0;
	wire w_dff_A_JtEJsWvz5_2;
	wire w_dff_A_RgWFr1om1_0;
	wire w_dff_A_z35lUeDj8_0;
	wire w_dff_A_kxs59J0J1_0;
	wire w_dff_A_T6Z5mPxI4_0;
	wire w_dff_A_BPwf4RUr5_0;
	wire w_dff_A_Yowidf4B2_0;
	wire w_dff_A_y4Lb7yxw8_0;
	wire w_dff_A_En05gtRn1_0;
	wire w_dff_A_Xg0EORiO8_0;
	wire w_dff_A_do6nehmm3_0;
	wire w_dff_A_zcAkv89N2_0;
	wire w_dff_A_GxEeDsfF3_0;
	wire w_dff_A_rYnVwgbd8_0;
	wire w_dff_A_zpGG2Epo0_0;
	wire w_dff_A_T9rnltFe9_0;
	wire w_dff_A_ufgHCMDh0_0;
	wire w_dff_A_VXgXdQO33_2;
	wire w_dff_A_QoAfB4xV7_0;
	wire w_dff_A_qdlT4Qmi0_0;
	wire w_dff_A_wKFO3nBv6_0;
	wire w_dff_A_nVaZOBoR7_0;
	wire w_dff_A_klkChoYf7_0;
	wire w_dff_A_HOS84ROD3_0;
	wire w_dff_A_euiWmpy41_0;
	wire w_dff_A_sv8AxLK32_0;
	wire w_dff_A_VN5JsFDp9_0;
	wire w_dff_A_rIALY9Lu8_0;
	wire w_dff_A_MCdaAqhP8_0;
	wire w_dff_A_e7TUax423_0;
	wire w_dff_A_K9RL7O5H6_0;
	wire w_dff_A_1g012K3M1_0;
	wire w_dff_A_jVwmXysm7_0;
	wire w_dff_A_b4LprVON7_0;
	wire w_dff_A_Vy0iPKTt6_0;
	wire w_dff_A_mvmvstLj6_2;
	wire w_dff_A_roSsMDkw8_0;
	wire w_dff_A_rJnnjq135_0;
	wire w_dff_A_aBdCM3vx1_0;
	wire w_dff_A_lTMycKqF8_0;
	wire w_dff_A_mWSbzQui7_0;
	wire w_dff_A_0kwWmSbM3_0;
	wire w_dff_A_HkcuJTrZ8_0;
	wire w_dff_A_xFaU33vH3_0;
	wire w_dff_A_tJ3L6kF58_0;
	wire w_dff_A_8DZTt0635_0;
	wire w_dff_A_PqyY8gLg0_0;
	wire w_dff_A_YVRePyug4_0;
	wire w_dff_A_K4iCGIuu2_0;
	wire w_dff_A_VLntJJmv0_0;
	wire w_dff_A_poeiRc8d5_0;
	wire w_dff_A_ShEdM7Zq4_0;
	wire w_dff_A_zRXboWsx4_0;
	wire w_dff_A_V0h2bNiz8_2;
	wire w_dff_A_VhYTCX0u0_0;
	wire w_dff_A_OQEG2g6w3_0;
	wire w_dff_A_EiyWRMx56_0;
	wire w_dff_A_75ThU4Se8_0;
	wire w_dff_A_ndBHxp119_0;
	wire w_dff_A_Nq2CmN0x1_0;
	wire w_dff_A_osrRrLa16_0;
	wire w_dff_A_XrIWils97_0;
	wire w_dff_A_oVglMcof2_0;
	wire w_dff_A_NZwfK0w07_0;
	wire w_dff_A_Cz4iHh9w7_0;
	wire w_dff_A_zlFk3Zpt3_0;
	wire w_dff_A_9Nhf94Pr2_0;
	wire w_dff_A_asPOGsDj3_0;
	wire w_dff_A_YtitRDRr3_0;
	wire w_dff_A_zMJfpbpH5_0;
	wire w_dff_A_U2gmkXaP9_0;
	wire w_dff_A_ivAHcPXp4_2;
	wire w_dff_A_V8FK9o7q5_0;
	wire w_dff_A_wCwWlHje0_0;
	wire w_dff_A_AG4ASDGc5_0;
	wire w_dff_A_npQicJ6G0_0;
	wire w_dff_A_BOxdcJ2r3_0;
	wire w_dff_A_q2oTiYMh5_0;
	wire w_dff_A_0MO7Ygaz5_0;
	wire w_dff_A_ptWoyQDO7_0;
	wire w_dff_A_Z7SdAHdf9_0;
	wire w_dff_A_LTpyagcE5_0;
	wire w_dff_A_TdrrNlVC7_0;
	wire w_dff_A_RQN5qq0y7_0;
	wire w_dff_A_cN4MUD593_0;
	wire w_dff_A_2BDZbHvk2_0;
	wire w_dff_A_BqanhjYR4_0;
	wire w_dff_A_XDfK61qz5_0;
	wire w_dff_A_vw1sRUCY3_0;
	wire w_dff_A_LqvkWp1d7_0;
	wire w_dff_A_4az9XDkv0_2;
	wire w_dff_A_DNbR0gOT8_0;
	wire w_dff_A_jI86XLkh7_0;
	wire w_dff_A_96ag7xpi2_0;
	wire w_dff_A_VA3YOs9B7_0;
	wire w_dff_A_EWdfiAOS7_0;
	wire w_dff_A_owjYhts39_0;
	wire w_dff_A_509KKv2Y4_0;
	wire w_dff_A_cyIMQczN9_0;
	wire w_dff_A_e62MMZiP0_0;
	wire w_dff_A_NUQstSp63_0;
	wire w_dff_A_bd3IgbbK2_0;
	wire w_dff_A_Ik5DVA7z7_0;
	wire w_dff_A_6IvIwkv89_0;
	wire w_dff_A_4vQ4Uihz0_0;
	wire w_dff_A_of1NuLC28_0;
	wire w_dff_A_FwjUHzgo8_0;
	wire w_dff_A_WuI0a5an7_1;
	wire w_dff_A_weJI9HQ41_0;
	wire w_dff_A_AKunf6VD6_0;
	wire w_dff_A_diOA7yQC8_0;
	wire w_dff_A_6x0iqUGO1_0;
	wire w_dff_A_0JqbgIkv3_0;
	wire w_dff_A_U3pZZzgv1_0;
	wire w_dff_A_lc6C4k3M5_0;
	wire w_dff_A_AogsuvoC4_0;
	wire w_dff_A_hA0u7aOT5_0;
	wire w_dff_A_GKh59UX61_0;
	wire w_dff_A_TutI7v6w2_0;
	wire w_dff_A_IHwdLI531_0;
	wire w_dff_A_TWSbq6RZ2_0;
	wire w_dff_A_84BhZORN9_0;
	wire w_dff_A_eEijS2vl3_0;
	wire w_dff_A_N6hh6wCw7_0;
	wire w_dff_A_tR0UUYRn2_0;
	wire w_dff_A_sKPHJm6Z0_0;
	wire w_dff_A_jR1N3iZq0_2;
	wire w_dff_A_cKyxqtlf9_0;
	wire w_dff_A_KFJitIqo3_0;
	wire w_dff_A_aAVUwLZq8_0;
	wire w_dff_A_xB2QAPUt3_0;
	wire w_dff_A_PcKBPz9O4_0;
	wire w_dff_A_gpeQwYZV5_0;
	wire w_dff_A_u95OFNOR2_0;
	wire w_dff_A_Rm6YChnj1_0;
	wire w_dff_A_LgKvJU7O5_0;
	wire w_dff_A_eUy7NZfC5_0;
	wire w_dff_A_U3Z5fkzs6_0;
	wire w_dff_A_e75DRMSb7_0;
	wire w_dff_A_RyoJMhlL3_0;
	wire w_dff_A_rVhWEfiY7_0;
	wire w_dff_A_1ScZ9tJJ4_0;
	wire w_dff_A_pdf2ggUj7_0;
	wire w_dff_A_sfPjeD881_0;
	wire w_dff_A_jogfoXaH2_2;
	wire w_dff_A_PYaA5tuj5_0;
	wire w_dff_A_8RcVT56I6_0;
	wire w_dff_A_UxH3WkMn3_0;
	wire w_dff_A_6oV0JVcf2_0;
	wire w_dff_A_1GYLlQJV4_0;
	wire w_dff_A_Ynr23nDp5_0;
	wire w_dff_A_28voCodS5_0;
	wire w_dff_A_3NcJpqE30_0;
	wire w_dff_A_AcuqVTbn3_0;
	wire w_dff_A_HnjujpJY0_0;
	wire w_dff_A_fui5hW7b7_0;
	wire w_dff_A_SltGA6xd8_0;
	wire w_dff_A_UFtlop9h0_0;
	wire w_dff_A_AGZUqGvm6_0;
	wire w_dff_A_1rhL1QCK2_0;
	wire w_dff_A_rcbqH4gR9_0;
	wire w_dff_A_YeEfp5zb8_0;
	wire w_dff_A_6SYhABzE8_2;
	wire w_dff_A_U9l8KWph0_0;
	wire w_dff_A_xTRv7I7J8_0;
	wire w_dff_A_4Lor9QnW8_0;
	wire w_dff_A_9BnkiIt54_0;
	wire w_dff_A_qWsc6p1C4_0;
	wire w_dff_A_SaDm0roK8_0;
	wire w_dff_A_yD6iCniA3_0;
	wire w_dff_A_1hnQitfW9_0;
	wire w_dff_A_ef7ZwlsO4_0;
	wire w_dff_A_U6BkSmyZ6_0;
	wire w_dff_A_zsV6ZeO50_0;
	wire w_dff_A_qSKnGyur4_0;
	wire w_dff_A_MSmYgbIt5_0;
	wire w_dff_A_QUDYou8I0_0;
	wire w_dff_A_nZhjkkeD8_0;
	wire w_dff_A_CwiNN6iy1_0;
	wire w_dff_A_Jg3GDmmY5_0;
	wire w_dff_A_hXxK4DLd5_0;
	wire w_dff_A_HjMSVorL4_2;
	wire w_dff_A_8d8VRant6_0;
	wire w_dff_A_EPf7X4f57_0;
	wire w_dff_A_3QNGAKnf1_0;
	wire w_dff_A_EATE4LbZ5_0;
	wire w_dff_A_pxwTyGmv4_0;
	wire w_dff_A_Jhd9VjBL5_0;
	wire w_dff_A_iagwmn7t7_0;
	wire w_dff_A_SC21QAg04_0;
	wire w_dff_A_5riHEL4U7_0;
	wire w_dff_A_UNBskL4w0_0;
	wire w_dff_A_3KoqT49O3_0;
	wire w_dff_A_1gvU1Uhq7_0;
	wire w_dff_A_F60jt1aF1_0;
	wire w_dff_A_H7c7vsDf8_0;
	wire w_dff_A_0dm0PEOh3_0;
	wire w_dff_A_0hgwa0Rq2_0;
	wire w_dff_A_joxD1bRl8_2;
	wire w_dff_A_J13CEXhl5_0;
	wire w_dff_A_pOIz6fq12_0;
	wire w_dff_A_dovxfJBW0_0;
	wire w_dff_A_0dVxO6IS7_0;
	wire w_dff_A_ZiItk0eJ5_0;
	wire w_dff_A_gDherlCp1_0;
	wire w_dff_A_s5VJe8cS8_0;
	wire w_dff_A_83wDDOFU6_0;
	wire w_dff_A_l8jVQVac7_0;
	wire w_dff_A_y59X553Y8_0;
	wire w_dff_A_QtGCyVVl8_0;
	wire w_dff_A_yqlYxW6i3_0;
	wire w_dff_A_BFFUtggX3_0;
	wire w_dff_A_muWherAh0_0;
	wire w_dff_A_77Yh6PNd4_0;
	wire w_dff_A_aDEixSED6_0;
	wire w_dff_A_Hgt1Xa0m0_2;
	wire w_dff_A_vHjowtHT0_0;
	wire w_dff_A_ncYT3LV94_0;
	wire w_dff_A_YumxXzvL1_0;
	wire w_dff_A_hQfwjWuz3_0;
	wire w_dff_A_mtW0mJYG9_0;
	wire w_dff_A_kAG5UFsj0_0;
	wire w_dff_A_Ik4L36mt5_0;
	wire w_dff_A_6DjvaEd45_2;
	wire w_dff_A_7hJsL7Kz2_0;
	wire w_dff_A_ioXI4HxI9_0;
	wire w_dff_A_jdt7MhOb7_0;
	wire w_dff_A_Yomum5wG5_2;
	wire w_dff_A_CaOgh5Yg7_0;
	wire w_dff_A_pL78jcLq3_0;
	wire w_dff_A_9hyLUzWt7_0;
	wire w_dff_A_WotfRuLH0_2;
	wire w_dff_A_3r6LbCBP9_0;
	wire w_dff_A_fps8k8ed6_0;
	wire w_dff_A_e70X0dyi0_0;
	wire w_dff_A_1VAwtGq65_0;
	wire w_dff_A_ksBZVi5i8_0;
	wire w_dff_A_Fm9M2ftm8_2;
	wire w_dff_A_zB1UnxD10_0;
	wire w_dff_A_Pv2dfkZ83_2;
	wire w_dff_A_sW3hjTUa3_0;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(w_dff_A_12pK7KFc3_2),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(w_dff_A_FYUoAM6L3_2),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(w_dff_A_ZCq0xqL09_2),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_G17gat_2[2]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_n92_0[2]),.dout(w_dff_A_sp5SF7qA2_2),.clk(gclk));
	jnot g009(.din(w_n93_0[0]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G1gat_1[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G26gat_0[1]),.dout(n97),.clk(gclk));
	jor g012(.dina(n97),.dinb(w_n96_0[1]),.dout(n98),.clk(gclk));
	jor g013(.dina(w_n98_0[1]),.dinb(n95),.dout(n99),.clk(gclk));
	jor g014(.dina(w_n99_0[1]),.dinb(w_G390gat_0[1]),.dout(w_dff_A_JtEJsWvz5_2),.clk(gclk));
	jnot g015(.din(w_G80gat_0[1]),.dout(n101),.clk(gclk));
	jand g016(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n102),.clk(gclk));
	jnot g017(.din(w_n102_0[1]),.dout(n103),.clk(gclk));
	jor g018(.dina(n103),.dinb(w_n101_0[1]),.dout(w_dff_A_VXgXdQO33_2),.clk(gclk));
	jnot g019(.din(w_G36gat_0[0]),.dout(n105),.clk(gclk));
	jnot g020(.din(w_G59gat_1[0]),.dout(n106),.clk(gclk));
	jor g021(.dina(w_n106_0[1]),.dinb(n105),.dout(n107),.clk(gclk));
	jor g022(.dina(w_n107_0[1]),.dinb(w_n101_0[0]),.dout(w_dff_A_mvmvstLj6_2),.clk(gclk));
	jnot g023(.din(w_G42gat_1[2]),.dout(n109),.clk(gclk));
	jor g024(.dina(w_n107_0[0]),.dinb(w_dff_B_tiKX16Px0_1),.dout(w_dff_A_V0h2bNiz8_2),.clk(gclk));
	jor g025(.dina(G88gat),.dinb(G87gat),.dout(n111),.clk(gclk));
	jand g026(.dina(w_n111_0[1]),.dinb(w_dff_B_e4pn1wKp5_1),.dout(w_dff_A_ivAHcPXp4_2),.clk(gclk));
	jnot g027(.din(w_G390gat_0[0]),.dout(n113),.clk(gclk));
	jor g028(.dina(w_n99_0[0]),.dinb(n113),.dout(w_dff_A_4az9XDkv0_2),.clk(gclk));
	jand g029(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n115),.clk(gclk));
	jand g030(.dina(n115),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g031(.dina(w_G55gat_0[2]),.dinb(w_G13gat_0[0]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_n92_0[1]),.dout(n118),.clk(gclk));
	jand g033(.dina(w_G68gat_0[1]),.dinb(w_G29gat_0[0]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_dff_B_TXvRpIgY2_0),.dinb(w_n118_0[2]),.dout(w_dff_A_jR1N3iZq0_2),.clk(gclk));
	jand g035(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n121),.clk(gclk));
	jand g036(.dina(w_n121_0[1]),.dinb(G74gat),.dout(n122),.clk(gclk));
	jand g037(.dina(n122),.dinb(w_n118_0[1]),.dout(w_dff_A_jogfoXaH2_2),.clk(gclk));
	jand g038(.dina(w_n111_0[0]),.dinb(w_dff_B_IhX0KD3f3_1),.dout(w_dff_A_6SYhABzE8_2),.clk(gclk));
	jxor g039(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n125),.clk(gclk));
	jxor g040(.dina(n125),.dinb(w_G130gat_0[1]),.dout(n126),.clk(gclk));
	jxor g041(.dina(w_G126gat_0[1]),.dinb(w_G121gat_0[2]),.dout(n127),.clk(gclk));
	jxor g042(.dina(n127),.dinb(n126),.dout(n128),.clk(gclk));
	jxor g043(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n129),.clk(gclk));
	jxor g044(.dina(n129),.dinb(G135gat),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(n131),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n128),.dout(w_dff_A_HjMSVorL4_2),.clk(gclk));
	jxor g048(.dina(w_G165gat_2[1]),.dinb(w_G159gat_2[1]),.dout(n134),.clk(gclk));
	jxor g049(.dina(n134),.dinb(w_G130gat_0[0]),.dout(n135),.clk(gclk));
	jxor g050(.dina(w_G201gat_2[2]),.dinb(w_G195gat_2[1]),.dout(n136),.clk(gclk));
	jxor g051(.dina(n136),.dinb(n135),.dout(n137),.clk(gclk));
	jxor g052(.dina(w_G189gat_2[1]),.dinb(w_G183gat_2[1]),.dout(n138),.clk(gclk));
	jxor g053(.dina(n138),.dinb(G207gat),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G177gat_2[1]),.dinb(w_G171gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n137),.dout(w_dff_A_joxD1bRl8_2),.clk(gclk));
	jnot g057(.din(w_G261gat_0[2]),.dout(n143),.clk(gclk));
	jand g058(.dina(w_n102_0[0]),.dinb(w_G42gat_1[1]),.dout(n144),.clk(gclk));
	jnot g059(.din(n144),.dout(n145),.clk(gclk));
	jand g060(.dina(w_G51gat_1[0]),.dinb(w_G17gat_2[1]),.dout(n146),.clk(gclk));
	jand g061(.dina(n146),.dinb(w_n92_0[0]),.dout(n147),.clk(gclk));
	jand g062(.dina(n147),.dinb(n145),.dout(n148),.clk(gclk));
	jand g063(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n149),.clk(gclk));
	jxor g064(.dina(w_G42gat_1[0]),.dinb(w_G17gat_2[0]),.dout(n150),.clk(gclk));
	jand g065(.dina(n150),.dinb(w_n149_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(n151),.dinb(w_G447gat_1),.dout(n152),.clk(gclk));
	jor g067(.dina(w_dff_B_zoCoK8vb1_0),.dinb(n148),.dout(n153),.clk(gclk));
	jand g068(.dina(w_n153_3[1]),.dinb(w_G126gat_0[0]),.dout(n154),.clk(gclk));
	jnot g069(.din(w_G156gat_0[0]),.dout(n155),.clk(gclk));
	jor g070(.dina(n155),.dinb(w_n106_0[0]),.dout(n156),.clk(gclk));
	jand g071(.dina(n156),.dinb(w_G447gat_0[2]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n157_0[1]),.dinb(w_G17gat_1[2]),.dout(n158),.clk(gclk));
	jor g073(.dina(n158),.dinb(w_n96_0[0]),.dout(n159),.clk(gclk));
	jand g074(.dina(w_n159_1[1]),.dinb(w_G153gat_0[2]),.dout(n160),.clk(gclk));
	jand g075(.dina(w_n86_0[0]),.dinb(w_G80gat_0[0]),.dout(n161),.clk(gclk));
	jand g076(.dina(n161),.dinb(w_G447gat_0[1]),.dout(n162),.clk(gclk));
	jnot g077(.din(w_G268gat_0[1]),.dout(n163),.clk(gclk));
	jand g078(.dina(w_n163_0[1]),.dinb(w_G55gat_0[1]),.dout(n164),.clk(gclk));
	jand g079(.dina(w_dff_B_mUBMt6NB3_0),.dinb(w_n162_0[1]),.dout(n165),.clk(gclk));
	jor g080(.dina(w_n165_1[2]),.dinb(n160),.dout(n166),.clk(gclk));
	jor g081(.dina(n166),.dinb(w_n154_0[1]),.dout(n167),.clk(gclk));
	jxor g082(.dina(w_n167_1[1]),.dinb(w_G201gat_2[1]),.dout(n168),.clk(gclk));
	jnot g083(.din(w_n168_0[2]),.dout(n169),.clk(gclk));
	jor g084(.dina(n169),.dinb(w_n143_0[1]),.dout(n170),.clk(gclk));
	jor g085(.dina(w_n168_0[1]),.dinb(w_G261gat_0[1]),.dout(n171),.clk(gclk));
	jand g086(.dina(n171),.dinb(w_G219gat_3[1]),.dout(n172),.clk(gclk));
	jand g087(.dina(n172),.dinb(n170),.dout(n173),.clk(gclk));
	jand g088(.dina(w_n168_0[0]),.dinb(w_G228gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_G237gat_3[1]),.dinb(w_G201gat_2[0]),.dout(n175),.clk(gclk));
	jor g090(.dina(n175),.dinb(w_G246gat_3[1]),.dout(n176),.clk(gclk));
	jand g091(.dina(w_dff_B_6vZlHYDc3_0),.dinb(w_n167_1[0]),.dout(n177),.clk(gclk));
	jand g092(.dina(G72gat),.dinb(w_G42gat_0[2]),.dout(n178),.clk(gclk));
	jand g093(.dina(n178),.dinb(G73gat),.dout(n179),.clk(gclk));
	jand g094(.dina(n179),.dinb(w_n121_0[0]),.dout(n180),.clk(gclk));
	jand g095(.dina(n180),.dinb(w_n118_0[0]),.dout(n181),.clk(gclk));
	jand g096(.dina(w_n181_3[1]),.dinb(w_G201gat_1[2]),.dout(n182),.clk(gclk));
	jand g097(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n183),.clk(gclk));
	jand g098(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n184),.clk(gclk));
	jor g099(.dina(n184),.dinb(n183),.dout(n185),.clk(gclk));
	jor g100(.dina(n185),.dinb(n182),.dout(n186),.clk(gclk));
	jor g101(.dina(w_dff_B_OHVPmDnQ5_0),.dinb(n177),.dout(n187),.clk(gclk));
	jor g102(.dina(n187),.dinb(n174),.dout(n188),.clk(gclk));
	jor g103(.dina(w_dff_B_KRLc3MAG8_0),.dinb(n173),.dout(w_dff_A_Hgt1Xa0m0_2),.clk(gclk));
	jand g104(.dina(w_n159_1[0]),.dinb(w_G143gat_0[1]),.dout(n190),.clk(gclk));
	jand g105(.dina(w_n153_3[0]),.dinb(w_G111gat_0[1]),.dout(n191),.clk(gclk));
	jor g106(.dina(n191),.dinb(w_n165_1[1]),.dout(n192),.clk(gclk));
	jor g107(.dina(n192),.dinb(w_dff_B_7LyFN7op3_1),.dout(n193),.clk(gclk));
	jxor g108(.dina(w_n193_1[1]),.dinb(w_G183gat_2[0]),.dout(n194),.clk(gclk));
	jnot g109(.din(w_n194_0[2]),.dout(n195),.clk(gclk));
	jand g110(.dina(w_n167_0[2]),.dinb(w_G201gat_1[1]),.dout(n196),.clk(gclk));
	jnot g111(.din(w_n196_0[1]),.dout(n197),.clk(gclk));
	jnot g112(.din(w_G201gat_1[0]),.dout(n198),.clk(gclk));
	jnot g113(.din(w_n154_0[0]),.dout(n199),.clk(gclk));
	jnot g114(.din(w_G153gat_0[1]),.dout(n200),.clk(gclk));
	jnot g115(.din(w_G17gat_1[1]),.dout(n201),.clk(gclk));
	jnot g116(.din(w_G51gat_0[2]),.dout(n202),.clk(gclk));
	jor g117(.dina(w_n98_0[0]),.dinb(n202),.dout(n203),.clk(gclk));
	jor g118(.dina(w_n149_0[0]),.dinb(n203),.dout(n204),.clk(gclk));
	jor g119(.dina(n204),.dinb(n201),.dout(n205),.clk(gclk));
	jand g120(.dina(n205),.dinb(w_G1gat_0[1]),.dout(n206),.clk(gclk));
	jor g121(.dina(n206),.dinb(n200),.dout(n207),.clk(gclk));
	jnot g122(.din(w_n165_1[0]),.dout(n208),.clk(gclk));
	jand g123(.dina(w_dff_B_JX4ZO1KH1_0),.dinb(n207),.dout(n209),.clk(gclk));
	jand g124(.dina(n209),.dinb(w_dff_B_00CMSlPU3_1),.dout(n210),.clk(gclk));
	jand g125(.dina(n210),.dinb(w_dff_B_Cy5q0l5Q0_1),.dout(n211),.clk(gclk));
	jor g126(.dina(n211),.dinb(w_n143_0[0]),.dout(n212),.clk(gclk));
	jand g127(.dina(n212),.dinb(w_dff_B_Wdi97rtg3_1),.dout(n213),.clk(gclk));
	jand g128(.dina(w_n159_0[2]),.dinb(w_G146gat_0[1]),.dout(n214),.clk(gclk));
	jand g129(.dina(w_n153_2[2]),.dinb(w_G116gat_0[1]),.dout(n215),.clk(gclk));
	jor g130(.dina(n215),.dinb(w_n165_0[2]),.dout(n216),.clk(gclk));
	jor g131(.dina(n216),.dinb(w_dff_B_vLsphLcm4_1),.dout(n217),.clk(gclk));
	jor g132(.dina(w_n217_1[1]),.dinb(w_G189gat_2[0]),.dout(n218),.clk(gclk));
	jand g133(.dina(w_n159_0[1]),.dinb(w_G149gat_0[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n153_2[1]),.dinb(w_G121gat_0[0]),.dout(n220),.clk(gclk));
	jor g135(.dina(n220),.dinb(w_n165_0[1]),.dout(n221),.clk(gclk));
	jor g136(.dina(n221),.dinb(w_dff_B_RbD4gjqX9_1),.dout(n222),.clk(gclk));
	jor g137(.dina(w_n222_1[1]),.dinb(w_G195gat_2[0]),.dout(n223),.clk(gclk));
	jand g138(.dina(w_n223_0[1]),.dinb(w_n218_0[1]),.dout(n224),.clk(gclk));
	jnot g139(.din(w_n224_0[1]),.dout(n225),.clk(gclk));
	jor g140(.dina(w_dff_B_5bvhS0zr2_0),.dinb(w_n213_0[1]),.dout(n226),.clk(gclk));
	jand g141(.dina(w_n217_1[0]),.dinb(w_G189gat_1[2]),.dout(n227),.clk(gclk));
	jand g142(.dina(w_n222_1[0]),.dinb(w_G195gat_1[2]),.dout(n228),.clk(gclk));
	jand g143(.dina(w_n228_0[1]),.dinb(w_n218_0[0]),.dout(n229),.clk(gclk));
	jor g144(.dina(n229),.dinb(w_dff_B_h7p1nVAO5_1),.dout(n230),.clk(gclk));
	jnot g145(.din(w_n230_0[1]),.dout(n231),.clk(gclk));
	jand g146(.dina(w_dff_B_tOdDF97N7_0),.dinb(n226),.dout(n232),.clk(gclk));
	jor g147(.dina(w_n232_0[1]),.dinb(w_dff_B_BYdBkM1K9_1),.dout(n233),.clk(gclk));
	jor g148(.dina(w_n167_0[1]),.dinb(w_G201gat_0[2]),.dout(n234),.clk(gclk));
	jand g149(.dina(n234),.dinb(w_G261gat_0[0]),.dout(n235),.clk(gclk));
	jor g150(.dina(n235),.dinb(w_n196_0[0]),.dout(n236),.clk(gclk));
	jand g151(.dina(w_n224_0[0]),.dinb(w_n236_0[2]),.dout(n237),.clk(gclk));
	jor g152(.dina(w_n230_0[0]),.dinb(n237),.dout(n238),.clk(gclk));
	jor g153(.dina(w_n238_0[1]),.dinb(w_n194_0[1]),.dout(n239),.clk(gclk));
	jand g154(.dina(n239),.dinb(w_G219gat_3[0]),.dout(n240),.clk(gclk));
	jand g155(.dina(n240),.dinb(n233),.dout(n241),.clk(gclk));
	jand g156(.dina(w_n194_0[0]),.dinb(w_G228gat_3[0]),.dout(n242),.clk(gclk));
	jand g157(.dina(w_G237gat_3[0]),.dinb(w_G183gat_1[2]),.dout(n243),.clk(gclk));
	jor g158(.dina(n243),.dinb(w_G246gat_3[0]),.dout(n244),.clk(gclk));
	jand g159(.dina(w_dff_B_b07EYonu0_0),.dinb(w_n193_1[0]),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n181_3[0]),.dinb(w_G183gat_1[1]),.dout(n246),.clk(gclk));
	jand g161(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n247),.clk(gclk));
	jor g162(.dina(n247),.dinb(n246),.dout(n248),.clk(gclk));
	jor g163(.dina(w_dff_B_IfUvKnRA3_0),.dinb(n245),.dout(n249),.clk(gclk));
	jor g164(.dina(n249),.dinb(n242),.dout(n250),.clk(gclk));
	jor g165(.dina(w_dff_B_Ts0mu9dQ2_0),.dinb(n241),.dout(w_dff_A_6DjvaEd45_2),.clk(gclk));
	jxor g166(.dina(w_n217_0[2]),.dinb(w_G189gat_1[1]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n252_0[2]),.dout(n253),.clk(gclk));
	jand g168(.dina(w_n223_0[0]),.dinb(w_n236_0[1]),.dout(n254),.clk(gclk));
	jor g169(.dina(n254),.dinb(w_n228_0[0]),.dout(n255),.clk(gclk));
	jnot g170(.din(w_n255_0[1]),.dout(n256),.clk(gclk));
	jor g171(.dina(n256),.dinb(w_dff_B_foePtHae1_1),.dout(n257),.clk(gclk));
	jor g172(.dina(w_n255_0[0]),.dinb(w_n252_0[1]),.dout(n258),.clk(gclk));
	jand g173(.dina(n258),.dinb(w_G219gat_2[2]),.dout(n259),.clk(gclk));
	jand g174(.dina(n259),.dinb(n257),.dout(n260),.clk(gclk));
	jand g175(.dina(w_n252_0[0]),.dinb(w_G228gat_2[2]),.dout(n261),.clk(gclk));
	jand g176(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n262),.clk(gclk));
	jor g177(.dina(n262),.dinb(w_G246gat_2[2]),.dout(n263),.clk(gclk));
	jand g178(.dina(w_dff_B_Ao5ed7Sc2_0),.dinb(w_n217_0[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(w_n181_2[2]),.dinb(w_G189gat_0[2]),.dout(n265),.clk(gclk));
	jand g180(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n266),.clk(gclk));
	jand g181(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n267),.clk(gclk));
	jor g182(.dina(n267),.dinb(n266),.dout(n268),.clk(gclk));
	jor g183(.dina(n268),.dinb(n265),.dout(n269),.clk(gclk));
	jor g184(.dina(w_dff_B_rOr14aHw5_0),.dinb(n264),.dout(n270),.clk(gclk));
	jor g185(.dina(n270),.dinb(n261),.dout(n271),.clk(gclk));
	jor g186(.dina(w_dff_B_JUgQGpSK3_0),.dinb(n260),.dout(w_dff_A_Yomum5wG5_2),.clk(gclk));
	jxor g187(.dina(w_n222_0[2]),.dinb(w_G195gat_1[1]),.dout(n273),.clk(gclk));
	jnot g188(.din(w_n273_0[2]),.dout(n274),.clk(gclk));
	jor g189(.dina(w_dff_B_aXzCb0vT9_0),.dinb(w_n213_0[0]),.dout(n275),.clk(gclk));
	jor g190(.dina(w_n273_0[1]),.dinb(w_n236_0[0]),.dout(n276),.clk(gclk));
	jand g191(.dina(n276),.dinb(w_G219gat_2[1]),.dout(n277),.clk(gclk));
	jand g192(.dina(n277),.dinb(n275),.dout(n278),.clk(gclk));
	jand g193(.dina(w_n273_0[0]),.dinb(w_G228gat_2[1]),.dout(n279),.clk(gclk));
	jand g194(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n280),.clk(gclk));
	jor g195(.dina(n280),.dinb(w_G246gat_2[1]),.dout(n281),.clk(gclk));
	jand g196(.dina(w_dff_B_ldOh7XXr3_0),.dinb(w_n222_0[1]),.dout(n282),.clk(gclk));
	jand g197(.dina(w_n181_2[1]),.dinb(w_G195gat_0[2]),.dout(n283),.clk(gclk));
	jand g198(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n284),.clk(gclk));
	jand g199(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n285),.clk(gclk));
	jor g200(.dina(n285),.dinb(n284),.dout(n286),.clk(gclk));
	jor g201(.dina(n286),.dinb(n283),.dout(n287),.clk(gclk));
	jor g202(.dina(w_dff_B_m1dfGMgx5_0),.dinb(n282),.dout(n288),.clk(gclk));
	jor g203(.dina(n288),.dinb(n279),.dout(n289),.clk(gclk));
	jor g204(.dina(w_dff_B_1zNYJEzd3_0),.dinb(n278),.dout(w_dff_A_WotfRuLH0_2),.clk(gclk));
	jand g205(.dina(w_n153_2[0]),.dinb(w_G91gat_0[1]),.dout(n291),.clk(gclk));
	jand g206(.dina(w_n157_0[0]),.dinb(w_G55gat_0[0]),.dout(n292),.clk(gclk));
	jand g207(.dina(w_n292_1[1]),.dinb(w_G143gat_0[0]),.dout(n293),.clk(gclk));
	jand g208(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n294),.clk(gclk));
	jand g209(.dina(w_n163_0[0]),.dinb(w_G17gat_1[0]),.dout(n295),.clk(gclk));
	jand g210(.dina(w_dff_B_y0MrhwVI7_0),.dinb(w_n162_0[0]),.dout(n296),.clk(gclk));
	jor g211(.dina(w_n296_1[1]),.dinb(w_dff_B_9P1KBs8x2_1),.dout(n297),.clk(gclk));
	jor g212(.dina(n297),.dinb(n293),.dout(n298),.clk(gclk));
	jor g213(.dina(n298),.dinb(n291),.dout(n299),.clk(gclk));
	jand g214(.dina(w_n299_1[1]),.dinb(w_G159gat_2[0]),.dout(n300),.clk(gclk));
	jor g215(.dina(w_n299_1[0]),.dinb(w_G159gat_1[2]),.dout(n301),.clk(gclk));
	jand g216(.dina(w_n193_0[2]),.dinb(w_G183gat_1[0]),.dout(n302),.clk(gclk));
	jor g217(.dina(w_n193_0[1]),.dinb(w_G183gat_0[2]),.dout(n303),.clk(gclk));
	jand g218(.dina(w_n238_0[0]),.dinb(w_n303_0[1]),.dout(n304),.clk(gclk));
	jor g219(.dina(n304),.dinb(w_n302_0[1]),.dout(n305),.clk(gclk));
	jnot g220(.din(w_G165gat_2[0]),.dout(n306),.clk(gclk));
	jand g221(.dina(w_n153_1[2]),.dinb(w_G96gat_0[1]),.dout(n307),.clk(gclk));
	jand g222(.dina(w_n292_1[0]),.dinb(w_G146gat_0[0]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n309),.clk(gclk));
	jor g224(.dina(w_dff_B_G5GWcALe2_0),.dinb(w_n296_1[0]),.dout(n310),.clk(gclk));
	jor g225(.dina(n310),.dinb(n308),.dout(n311),.clk(gclk));
	jor g226(.dina(n311),.dinb(n307),.dout(n312),.clk(gclk));
	jnot g227(.din(w_n312_1[1]),.dout(n313),.clk(gclk));
	jand g228(.dina(n313),.dinb(w_dff_B_2AmxpU0q8_1),.dout(n314),.clk(gclk));
	jnot g229(.din(n314),.dout(n315),.clk(gclk));
	jand g230(.dina(w_n153_1[1]),.dinb(w_G101gat_0[1]),.dout(n316),.clk(gclk));
	jand g231(.dina(w_n292_0[2]),.dinb(w_G149gat_0[0]),.dout(n317),.clk(gclk));
	jand g232(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n318),.clk(gclk));
	jor g233(.dina(w_dff_B_lPbYyXpM1_0),.dinb(w_n296_0[2]),.dout(n319),.clk(gclk));
	jor g234(.dina(n319),.dinb(n317),.dout(n320),.clk(gclk));
	jor g235(.dina(n320),.dinb(n316),.dout(n321),.clk(gclk));
	jor g236(.dina(w_n321_1[1]),.dinb(w_G171gat_2[0]),.dout(n322),.clk(gclk));
	jand g237(.dina(w_n153_1[0]),.dinb(w_G106gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_n292_0[1]),.dinb(w_G153gat_0[0]),.dout(n324),.clk(gclk));
	jand g239(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n325),.clk(gclk));
	jor g240(.dina(w_dff_B_DLghQFNe1_0),.dinb(w_n296_0[1]),.dout(n326),.clk(gclk));
	jor g241(.dina(n326),.dinb(n324),.dout(n327),.clk(gclk));
	jor g242(.dina(n327),.dinb(n323),.dout(n328),.clk(gclk));
	jor g243(.dina(w_n328_1[1]),.dinb(w_G177gat_2[0]),.dout(n329),.clk(gclk));
	jand g244(.dina(w_n329_0[2]),.dinb(w_n322_0[1]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n330_0[2]),.dinb(w_n315_0[1]),.dout(n331),.clk(gclk));
	jand g246(.dina(w_n331_0[1]),.dinb(w_n305_1[1]),.dout(n332),.clk(gclk));
	jand g247(.dina(w_n312_1[0]),.dinb(w_G165gat_1[2]),.dout(n333),.clk(gclk));
	jand g248(.dina(w_n321_1[0]),.dinb(w_G171gat_1[2]),.dout(n334),.clk(gclk));
	jand g249(.dina(w_n328_1[0]),.dinb(w_G177gat_1[2]),.dout(n335),.clk(gclk));
	jand g250(.dina(w_n335_0[2]),.dinb(w_n322_0[0]),.dout(n336),.clk(gclk));
	jor g251(.dina(n336),.dinb(w_dff_B_G0UghCva0_1),.dout(n337),.clk(gclk));
	jand g252(.dina(w_n337_0[2]),.dinb(w_n315_0[0]),.dout(n338),.clk(gclk));
	jor g253(.dina(n338),.dinb(w_dff_B_alhlfcJh7_1),.dout(n339),.clk(gclk));
	jor g254(.dina(w_n339_0[1]),.dinb(n332),.dout(n340),.clk(gclk));
	jand g255(.dina(w_n340_0[1]),.dinb(w_dff_B_JqCAedvZ7_1),.dout(n341),.clk(gclk));
	jor g256(.dina(n341),.dinb(w_dff_B_fePUdM2d9_1),.dout(w_dff_A_Fm9M2ftm8_2),.clk(gclk));
	jnot g257(.din(w_n302_0[0]),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n303_0[0]),.dout(n344),.clk(gclk));
	jor g259(.dina(w_n232_0[0]),.dinb(w_dff_B_e3KOWU6d5_1),.dout(n345),.clk(gclk));
	jand g260(.dina(n345),.dinb(w_dff_B_XPX9zK4e7_1),.dout(n346),.clk(gclk));
	jxor g261(.dina(w_n328_0[2]),.dinb(w_G177gat_1[1]),.dout(n347),.clk(gclk));
	jnot g262(.din(w_n347_0[2]),.dout(n348),.clk(gclk));
	jor g263(.dina(w_dff_B_xzkYETx73_0),.dinb(w_n346_1[1]),.dout(n349),.clk(gclk));
	jor g264(.dina(w_n347_0[1]),.dinb(w_n305_1[0]),.dout(n350),.clk(gclk));
	jand g265(.dina(n350),.dinb(w_G219gat_2[0]),.dout(n351),.clk(gclk));
	jand g266(.dina(n351),.dinb(n349),.dout(n352),.clk(gclk));
	jand g267(.dina(w_n347_0[0]),.dinb(w_G228gat_2[0]),.dout(n353),.clk(gclk));
	jand g268(.dina(w_G237gat_2[0]),.dinb(w_G177gat_1[0]),.dout(n354),.clk(gclk));
	jor g269(.dina(n354),.dinb(w_G246gat_2[0]),.dout(n355),.clk(gclk));
	jand g270(.dina(w_dff_B_KFCGK5jy3_0),.dinb(w_n328_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n181_2[0]),.dinb(w_G177gat_0[2]),.dout(n357),.clk(gclk));
	jand g272(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n358),.clk(gclk));
	jor g273(.dina(n358),.dinb(n357),.dout(n359),.clk(gclk));
	jor g274(.dina(w_dff_B_F5qxVQDB4_0),.dinb(n356),.dout(n360),.clk(gclk));
	jor g275(.dina(n360),.dinb(n353),.dout(n361),.clk(gclk));
	jor g276(.dina(w_dff_B_VGeWtE5A5_0),.dinb(n352),.dout(w_dff_A_Pv2dfkZ83_2),.clk(gclk));
	jnot g277(.din(w_n331_0[0]),.dout(n363),.clk(gclk));
	jor g278(.dina(w_dff_B_gdY9OzYR7_0),.dinb(w_n346_1[0]),.dout(n364),.clk(gclk));
	jnot g279(.din(w_n339_0[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_dff_B_Mf8HV2vp2_0),.dinb(n364),.dout(n366),.clk(gclk));
	jxor g281(.dina(w_n299_0[2]),.dinb(w_G159gat_1[1]),.dout(n367),.clk(gclk));
	jnot g282(.din(w_n367_0[2]),.dout(n368),.clk(gclk));
	jor g283(.dina(w_dff_B_eYxYzzQE9_0),.dinb(n366),.dout(n369),.clk(gclk));
	jor g284(.dina(w_n367_0[1]),.dinb(w_n340_0[0]),.dout(n370),.clk(gclk));
	jand g285(.dina(n370),.dinb(w_G219gat_1[2]),.dout(n371),.clk(gclk));
	jand g286(.dina(n371),.dinb(n369),.dout(n372),.clk(gclk));
	jand g287(.dina(w_n367_0[0]),.dinb(w_G228gat_1[2]),.dout(n373),.clk(gclk));
	jand g288(.dina(w_G237gat_1[2]),.dinb(w_G159gat_1[0]),.dout(n374),.clk(gclk));
	jor g289(.dina(n374),.dinb(w_G246gat_1[2]),.dout(n375),.clk(gclk));
	jand g290(.dina(w_dff_B_LpRmIxIQ1_0),.dinb(w_n299_0[1]),.dout(n376),.clk(gclk));
	jand g291(.dina(w_n181_1[2]),.dinb(w_G159gat_0[2]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n378),.clk(gclk));
	jor g293(.dina(n378),.dinb(n377),.dout(n379),.clk(gclk));
	jor g294(.dina(w_dff_B_m7emHeOP8_0),.dinb(n376),.dout(n380),.clk(gclk));
	jor g295(.dina(n380),.dinb(n373),.dout(n381),.clk(gclk));
	jor g296(.dina(w_dff_B_MP1MsEYv0_0),.dinb(n372),.dout(G878gat),.clk(gclk));
	jxor g297(.dina(w_n312_0[2]),.dinb(w_G165gat_1[1]),.dout(n383),.clk(gclk));
	jnot g298(.din(w_n383_0[2]),.dout(n384),.clk(gclk));
	jnot g299(.din(w_n337_0[1]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n330_0[1]),.dout(n386),.clk(gclk));
	jor g301(.dina(w_dff_B_2kkwxVAz8_0),.dinb(w_n346_0[2]),.dout(n387),.clk(gclk));
	jand g302(.dina(n387),.dinb(w_dff_B_1pNGs2sO1_1),.dout(n388),.clk(gclk));
	jor g303(.dina(n388),.dinb(w_dff_B_gYOXGW2O2_1),.dout(n389),.clk(gclk));
	jand g304(.dina(w_n330_0[0]),.dinb(w_n305_0[2]),.dout(n390),.clk(gclk));
	jor g305(.dina(n390),.dinb(w_n337_0[0]),.dout(n391),.clk(gclk));
	jor g306(.dina(n391),.dinb(w_n383_0[1]),.dout(n392),.clk(gclk));
	jand g307(.dina(n392),.dinb(w_G219gat_1[1]),.dout(n393),.clk(gclk));
	jand g308(.dina(n393),.dinb(n389),.dout(n394),.clk(gclk));
	jand g309(.dina(w_n383_0[0]),.dinb(w_G228gat_1[1]),.dout(n395),.clk(gclk));
	jand g310(.dina(w_G237gat_1[1]),.dinb(w_G165gat_1[0]),.dout(n396),.clk(gclk));
	jor g311(.dina(n396),.dinb(w_G246gat_1[1]),.dout(n397),.clk(gclk));
	jand g312(.dina(w_dff_B_ABwgDkzj8_0),.dinb(w_n312_0[1]),.dout(n398),.clk(gclk));
	jand g313(.dina(w_n181_1[1]),.dinb(w_G165gat_0[2]),.dout(n399),.clk(gclk));
	jand g314(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n400),.clk(gclk));
	jor g315(.dina(n400),.dinb(n399),.dout(n401),.clk(gclk));
	jor g316(.dina(w_dff_B_3BozDWWg7_0),.dinb(n398),.dout(n402),.clk(gclk));
	jor g317(.dina(n402),.dinb(n395),.dout(n403),.clk(gclk));
	jor g318(.dina(w_dff_B_JZYJZQ1Q8_0),.dinb(n394),.dout(G879gat),.clk(gclk));
	jxor g319(.dina(w_n321_0[2]),.dinb(w_G171gat_1[1]),.dout(n405),.clk(gclk));
	jnot g320(.din(w_n405_0[2]),.dout(n406),.clk(gclk));
	jnot g321(.din(w_n335_0[1]),.dout(n407),.clk(gclk));
	jnot g322(.din(w_n329_0[1]),.dout(n408),.clk(gclk));
	jor g323(.dina(w_dff_B_H7X158O22_0),.dinb(w_n346_0[1]),.dout(n409),.clk(gclk));
	jand g324(.dina(n409),.dinb(w_dff_B_iwS0WEyB8_1),.dout(n410),.clk(gclk));
	jor g325(.dina(n410),.dinb(w_dff_B_fAWAZmko4_1),.dout(n411),.clk(gclk));
	jand g326(.dina(w_n329_0[0]),.dinb(w_n305_0[1]),.dout(n412),.clk(gclk));
	jor g327(.dina(n412),.dinb(w_n335_0[0]),.dout(n413),.clk(gclk));
	jor g328(.dina(n413),.dinb(w_n405_0[1]),.dout(n414),.clk(gclk));
	jand g329(.dina(n414),.dinb(w_G219gat_1[0]),.dout(n415),.clk(gclk));
	jand g330(.dina(n415),.dinb(n411),.dout(n416),.clk(gclk));
	jand g331(.dina(w_n405_0[0]),.dinb(w_G228gat_1[0]),.dout(n417),.clk(gclk));
	jand g332(.dina(w_G237gat_1[0]),.dinb(w_G171gat_1[0]),.dout(n418),.clk(gclk));
	jor g333(.dina(n418),.dinb(w_G246gat_1[0]),.dout(n419),.clk(gclk));
	jand g334(.dina(w_dff_B_YpYObPOD1_0),.dinb(w_n321_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n181_1[0]),.dinb(w_G171gat_0[2]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jor g337(.dina(n422),.dinb(n421),.dout(n423),.clk(gclk));
	jor g338(.dina(w_dff_B_YkSpfOp92_0),.dinb(n420),.dout(n424),.clk(gclk));
	jor g339(.dina(n424),.dinb(n417),.dout(n425),.clk(gclk));
	jor g340(.dina(w_dff_B_eLkANbUv5_0),.dinb(n416),.dout(G880gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_G13gat_0[1]),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_G17gat_1[0]),.doutb(w_G17gat_1[1]),.doutc(w_G17gat_1[2]),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_G17gat_2[2]),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_G29gat_0[0]),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_G42gat_0[1]),.doutc(w_G42gat_0[2]),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_G42gat_1[0]),.doutb(w_G42gat_1[1]),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_G51gat_1[1]),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_G55gat_0[0]),.doutb(w_G55gat_0[1]),.doutc(w_G55gat_0[2]),.din(G55gat));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_G68gat_0[1]),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_G80gat_0[0]),.doutb(w_G80gat_0[1]),.doutc(w_G80gat_0[2]),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_G91gat_0[1]),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_G96gat_0[1]),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_G101gat_0[1]),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_G106gat_0[0]),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_G111gat_0[1]),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_G116gat_0[1]),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_G121gat_0[0]),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl jspl_w_G126gat_0(.douta(w_G126gat_0[0]),.doutb(w_G126gat_0[1]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_G130gat_0[1]),.din(G130gat));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_dff_A_C2Hev3HG1_1),.din(w_dff_B_5FCgSxWW5_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_dff_A_PLo5IAVx8_1),.din(w_dff_B_w4396kB92_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_dff_A_xfZ43KYV4_1),.din(w_dff_B_HZ81dAzI8_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_G153gat_0[0]),.doutb(w_G153gat_0[1]),.doutc(w_G153gat_0[2]),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_G159gat_0[1]),.doutc(w_G159gat_0[2]),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_G159gat_1[0]),.doutb(w_G159gat_1[1]),.doutc(w_G159gat_1[2]),.din(w_G159gat_0[0]));
	jspl jspl_w_G159gat_2(.douta(w_G159gat_2[0]),.doutb(w_G159gat_2[1]),.din(w_G159gat_0[1]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_G165gat_0[1]),.doutc(w_G165gat_0[2]),.din(G165gat));
	jspl3 jspl3_w_G165gat_1(.douta(w_G165gat_1[0]),.doutb(w_G165gat_1[1]),.doutc(w_G165gat_1[2]),.din(w_G165gat_0[0]));
	jspl jspl_w_G165gat_2(.douta(w_G165gat_2[0]),.doutb(w_G165gat_2[1]),.din(w_G165gat_0[1]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl jspl_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_G177gat_0[1]),.doutc(w_G177gat_0[2]),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_G177gat_1[1]),.doutc(w_G177gat_1[2]),.din(w_G177gat_0[0]));
	jspl jspl_w_G177gat_2(.douta(w_G177gat_2[0]),.doutb(w_G177gat_2[1]),.din(w_G177gat_0[1]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_G183gat_0[2]),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_G183gat_1[0]),.doutb(w_G183gat_1[1]),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl jspl_w_G183gat_2(.douta(w_G183gat_2[0]),.doutb(w_G183gat_2[1]),.din(w_G183gat_0[1]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_G189gat_0[2]),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_G189gat_1[1]),.doutc(w_G189gat_1[2]),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_G189gat_2[0]),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_G195gat_0[2]),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_G195gat_1[1]),.doutc(w_G195gat_1[2]),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_G195gat_2[0]),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_G201gat_0[1]),.doutc(w_G201gat_0[2]),.din(G201gat));
	jspl3 jspl3_w_G201gat_1(.douta(w_G201gat_1[0]),.doutb(w_G201gat_1[1]),.doutc(w_G201gat_1[2]),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G201gat_2(.douta(w_G201gat_2[0]),.doutb(w_G201gat_2[1]),.doutc(w_G201gat_2[2]),.din(w_G201gat_0[1]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_abCT3wmx7_0),.doutb(w_dff_A_PKbnaw7G5_1),.doutc(w_G219gat_0[2]),.din(w_dff_B_crlZpAfE1_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_G219gat_1[0]),.doutb(w_G219gat_1[1]),.doutc(w_G219gat_1[2]),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_CcZfl3DE9_0),.doutb(w_G219gat_2[1]),.doutc(w_dff_A_TjZN6dMJ0_2),.din(w_G219gat_0[1]));
	jspl jspl_w_G219gat_3(.douta(w_dff_A_8KFNZSZn2_0),.doutb(w_G219gat_3[1]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_G228gat_0[0]),.doutb(w_G228gat_0[1]),.doutc(w_dff_A_2iPPdsSE7_2),.din(w_dff_B_OJh4kz4m2_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_G228gat_2[0]),.doutb(w_dff_A_luHCqTH56_1),.doutc(w_dff_A_2q7bebE30_2),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_G228gat_3[1]),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_G237gat_0[0]),.doutb(w_G237gat_0[1]),.doutc(w_G237gat_0[2]),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_G237gat_2[0]),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_G237gat_3[1]),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_G246gat_0[0]),.doutb(w_G246gat_0[1]),.doutc(w_G246gat_0[2]),.din(G246gat));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_G246gat_2[0]),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_G246gat_3[1]),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_G261gat_0[0]),.doutb(w_G261gat_0[1]),.doutc(w_G261gat_0[2]),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_dff_A_VbzBPUP40_1),.doutc(w_dff_A_EHSzjLlc3_2),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_G447gat_0[2]),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(w_dff_A_WuI0a5an7_1),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_n86_0[0]),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl3 jspl3_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.doutc(w_n92_0[2]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_n98_0[0]),.doutb(w_n98_0[1]),.din(n98));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(w_dff_B_rcdGIbcJ4_2));
	jspl jspl_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.din(n102));
	jspl jspl_w_n106_0(.douta(w_n106_0[0]),.doutb(w_n106_0[1]),.din(n106));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n118_0(.douta(w_n118_0[0]),.doutb(w_n118_0[1]),.doutc(w_n118_0[2]),.din(n118));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(w_dff_B_cvM5anir9_2));
	jspl jspl_w_n149_0(.douta(w_n149_0[0]),.doutb(w_n149_0[1]),.din(n149));
	jspl3 jspl3_w_n153_0(.douta(w_n153_0[0]),.doutb(w_n153_0[1]),.doutc(w_n153_0[2]),.din(n153));
	jspl3 jspl3_w_n153_1(.douta(w_n153_1[0]),.doutb(w_n153_1[1]),.doutc(w_n153_1[2]),.din(w_n153_0[0]));
	jspl3 jspl3_w_n153_2(.douta(w_n153_2[0]),.doutb(w_n153_2[1]),.doutc(w_n153_2[2]),.din(w_n153_0[1]));
	jspl jspl_w_n153_3(.douta(w_n153_3[0]),.doutb(w_n153_3[1]),.din(w_n153_0[2]));
	jspl jspl_w_n154_0(.douta(w_n154_0[0]),.doutb(w_dff_A_opLtEpGM9_1),.din(n154));
	jspl jspl_w_n157_0(.douta(w_n157_0[0]),.doutb(w_n157_0[1]),.din(n157));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_n159_0[1]),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl jspl_w_n162_0(.douta(w_n162_0[0]),.doutb(w_n162_0[1]),.din(n162));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl3 jspl3_w_n165_0(.douta(w_n165_0[0]),.doutb(w_dff_A_3Sp17NIj4_1),.doutc(w_dff_A_7kPryKTi9_2),.din(n165));
	jspl3 jspl3_w_n165_1(.douta(w_n165_1[0]),.doutb(w_dff_A_XmYDxrZe7_1),.doutc(w_dff_A_AMWZ37Nv6_2),.din(w_n165_0[0]));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.doutc(w_n167_0[2]),.din(n167));
	jspl jspl_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.doutc(w_n168_0[2]),.din(n168));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n181_2(.douta(w_n181_2[0]),.doutb(w_n181_2[1]),.doutc(w_n181_2[2]),.din(w_n181_0[1]));
	jspl jspl_w_n181_3(.douta(w_n181_3[0]),.doutb(w_n181_3[1]),.din(w_n181_0[2]));
	jspl3 jspl3_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.doutc(w_n193_0[2]),.din(n193));
	jspl jspl_w_n193_1(.douta(w_n193_1[0]),.doutb(w_n193_1[1]),.din(w_n193_0[0]));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_dff_A_lZsuws234_1),.doutc(w_n194_0[2]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_dff_A_IqsW8ezY1_0),.doutb(w_n196_0[1]),.din(n196));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl3 jspl3_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.doutc(w_n217_0[2]),.din(n217));
	jspl jspl_w_n217_1(.douta(w_n217_1[0]),.doutb(w_n217_1[1]),.din(w_n217_0[0]));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(n218));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_n222_0[1]),.doutc(w_n222_0[2]),.din(n222));
	jspl jspl_w_n222_1(.douta(w_n222_1[0]),.doutb(w_n222_1[1]),.din(w_n222_0[0]));
	jspl jspl_w_n223_0(.douta(w_dff_A_kkq4hYOp2_0),.doutb(w_n223_0[1]),.din(n223));
	jspl jspl_w_n224_0(.douta(w_dff_A_d7IZQ9Sj4_0),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n228_0(.douta(w_dff_A_mZPGkEJ34_0),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n230_0(.douta(w_dff_A_c7Ea73oJ2_0),.doutb(w_n230_0[1]),.din(n230));
	jspl jspl_w_n232_0(.douta(w_n232_0[0]),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.doutc(w_n236_0[2]),.din(n236));
	jspl jspl_w_n238_0(.douta(w_n238_0[0]),.doutb(w_n238_0[1]),.din(n238));
	jspl3 jspl3_w_n252_0(.douta(w_n252_0[0]),.doutb(w_dff_A_9h2QmdbG4_1),.doutc(w_n252_0[2]),.din(n252));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_dff_A_5y9cMeqJ6_1),.doutc(w_n273_0[2]),.din(n273));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl jspl_w_n292_1(.douta(w_n292_1[0]),.doutb(w_n292_1[1]),.din(w_n292_0[0]));
	jspl3 jspl3_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.doutc(w_n296_0[2]),.din(n296));
	jspl jspl_w_n296_1(.douta(w_n296_1[0]),.doutb(w_n296_1[1]),.din(w_n296_0[0]));
	jspl3 jspl3_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.doutc(w_n299_0[2]),.din(n299));
	jspl jspl_w_n299_1(.douta(w_n299_1[0]),.doutb(w_n299_1[1]),.din(w_n299_0[0]));
	jspl jspl_w_n302_0(.douta(w_n302_0[0]),.doutb(w_dff_A_DxIJJiKv9_1),.din(n302));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_dff_A_4QIIxiCh7_1),.din(n303));
	jspl3 jspl3_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.doutc(w_n305_0[2]),.din(n305));
	jspl jspl_w_n305_1(.douta(w_n305_1[0]),.doutb(w_n305_1[1]),.din(w_n305_0[0]));
	jspl3 jspl3_w_n312_0(.douta(w_n312_0[0]),.doutb(w_n312_0[1]),.doutc(w_n312_0[2]),.din(n312));
	jspl jspl_w_n312_1(.douta(w_n312_1[0]),.doutb(w_n312_1[1]),.din(w_n312_0[0]));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl3 jspl3_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.doutc(w_n321_0[2]),.din(n321));
	jspl jspl_w_n321_1(.douta(w_n321_1[0]),.doutb(w_n321_1[1]),.din(w_n321_0[0]));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl3 jspl3_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.doutc(w_n328_0[2]),.din(n328));
	jspl jspl_w_n328_1(.douta(w_n328_1[0]),.doutb(w_n328_1[1]),.din(w_n328_0[0]));
	jspl3 jspl3_w_n329_0(.douta(w_dff_A_0Pnsip6t7_0),.doutb(w_n329_0[1]),.doutc(w_n329_0[2]),.din(n329));
	jspl3 jspl3_w_n330_0(.douta(w_dff_A_fJznWadX8_0),.doutb(w_n330_0[1]),.doutc(w_dff_A_Zqdv1tL21_2),.din(n330));
	jspl jspl_w_n331_0(.douta(w_n331_0[0]),.doutb(w_dff_A_L4YyDJsW5_1),.din(n331));
	jspl3 jspl3_w_n335_0(.douta(w_dff_A_kpotA8MX8_0),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl3 jspl3_w_n337_0(.douta(w_dff_A_W2JSlw2h6_0),.doutb(w_n337_0[1]),.doutc(w_n337_0[2]),.din(n337));
	jspl jspl_w_n339_0(.douta(w_n339_0[0]),.doutb(w_dff_A_ZHpQrXdH1_1),.din(n339));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n346_1(.douta(w_n346_1[0]),.doutb(w_n346_1[1]),.din(w_n346_0[0]));
	jspl3 jspl3_w_n347_0(.douta(w_n347_0[0]),.doutb(w_dff_A_fEwDBsn05_1),.doutc(w_n347_0[2]),.din(n347));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_dff_A_kL7E0WFL2_1),.doutc(w_n367_0[2]),.din(n367));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_dff_A_YRxUrohg1_1),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_dff_A_TyLlz1ve1_1),.doutc(w_n405_0[2]),.din(n405));
	jdff dff_B_rcdGIbcJ4_2(.din(n101),.dout(w_dff_B_rcdGIbcJ4_2),.clk(gclk));
	jdff dff_B_tiKX16Px0_1(.din(n109),.dout(w_dff_B_tiKX16Px0_1),.clk(gclk));
	jdff dff_B_e4pn1wKp5_1(.din(G90gat),.dout(w_dff_B_e4pn1wKp5_1),.clk(gclk));
	jdff dff_A_VbzBPUP40_1(.dout(w_G390gat_0[1]),.din(w_dff_A_VbzBPUP40_1),.clk(gclk));
	jdff dff_B_TXvRpIgY2_0(.din(n119),.dout(w_dff_B_TXvRpIgY2_0),.clk(gclk));
	jdff dff_B_IhX0KD3f3_1(.din(G89gat),.dout(w_dff_B_IhX0KD3f3_1),.clk(gclk));
	jdff dff_B_KRLc3MAG8_0(.din(n188),.dout(w_dff_B_KRLc3MAG8_0),.clk(gclk));
	jdff dff_B_enXRNkZg0_0(.din(n186),.dout(w_dff_B_enXRNkZg0_0),.clk(gclk));
	jdff dff_B_Owi7afwE7_0(.din(w_dff_B_enXRNkZg0_0),.dout(w_dff_B_Owi7afwE7_0),.clk(gclk));
	jdff dff_B_OHVPmDnQ5_0(.din(w_dff_B_Owi7afwE7_0),.dout(w_dff_B_OHVPmDnQ5_0),.clk(gclk));
	jdff dff_B_Nvw7oXI35_0(.din(n176),.dout(w_dff_B_Nvw7oXI35_0),.clk(gclk));
	jdff dff_B_z3ubSxCI4_0(.din(w_dff_B_Nvw7oXI35_0),.dout(w_dff_B_z3ubSxCI4_0),.clk(gclk));
	jdff dff_B_HhNG3CKU3_0(.din(w_dff_B_z3ubSxCI4_0),.dout(w_dff_B_HhNG3CKU3_0),.clk(gclk));
	jdff dff_B_USfRZPqj1_0(.din(w_dff_B_HhNG3CKU3_0),.dout(w_dff_B_USfRZPqj1_0),.clk(gclk));
	jdff dff_B_AmGWvrWg3_0(.din(w_dff_B_USfRZPqj1_0),.dout(w_dff_B_AmGWvrWg3_0),.clk(gclk));
	jdff dff_B_6vZlHYDc3_0(.din(w_dff_B_AmGWvrWg3_0),.dout(w_dff_B_6vZlHYDc3_0),.clk(gclk));
	jdff dff_B_lVb7JkCh4_0(.din(n250),.dout(w_dff_B_lVb7JkCh4_0),.clk(gclk));
	jdff dff_B_ablkYAcJ7_0(.din(w_dff_B_lVb7JkCh4_0),.dout(w_dff_B_ablkYAcJ7_0),.clk(gclk));
	jdff dff_B_2tF9mHCD8_0(.din(w_dff_B_ablkYAcJ7_0),.dout(w_dff_B_2tF9mHCD8_0),.clk(gclk));
	jdff dff_B_aF4hJVaf0_0(.din(w_dff_B_2tF9mHCD8_0),.dout(w_dff_B_aF4hJVaf0_0),.clk(gclk));
	jdff dff_B_Ts0mu9dQ2_0(.din(w_dff_B_aF4hJVaf0_0),.dout(w_dff_B_Ts0mu9dQ2_0),.clk(gclk));
	jdff dff_B_OBt1jgVH8_0(.din(n248),.dout(w_dff_B_OBt1jgVH8_0),.clk(gclk));
	jdff dff_B_LSU65Vw94_0(.din(w_dff_B_OBt1jgVH8_0),.dout(w_dff_B_LSU65Vw94_0),.clk(gclk));
	jdff dff_B_IfUvKnRA3_0(.din(w_dff_B_LSU65Vw94_0),.dout(w_dff_B_IfUvKnRA3_0),.clk(gclk));
	jdff dff_B_e89rPMCW6_0(.din(n244),.dout(w_dff_B_e89rPMCW6_0),.clk(gclk));
	jdff dff_B_oXLMxhMh5_0(.din(w_dff_B_e89rPMCW6_0),.dout(w_dff_B_oXLMxhMh5_0),.clk(gclk));
	jdff dff_B_EbYTPf9d3_0(.din(w_dff_B_oXLMxhMh5_0),.dout(w_dff_B_EbYTPf9d3_0),.clk(gclk));
	jdff dff_B_YqIEs0iB3_0(.din(w_dff_B_EbYTPf9d3_0),.dout(w_dff_B_YqIEs0iB3_0),.clk(gclk));
	jdff dff_B_fZttj8oE1_0(.din(w_dff_B_YqIEs0iB3_0),.dout(w_dff_B_fZttj8oE1_0),.clk(gclk));
	jdff dff_B_b07EYonu0_0(.din(w_dff_B_fZttj8oE1_0),.dout(w_dff_B_b07EYonu0_0),.clk(gclk));
	jdff dff_A_w1Bf2Yr52_0(.dout(w_G219gat_3[0]),.din(w_dff_A_w1Bf2Yr52_0),.clk(gclk));
	jdff dff_A_NVPALc7q9_0(.dout(w_dff_A_w1Bf2Yr52_0),.din(w_dff_A_NVPALc7q9_0),.clk(gclk));
	jdff dff_A_6dCSBIm63_0(.dout(w_dff_A_NVPALc7q9_0),.din(w_dff_A_6dCSBIm63_0),.clk(gclk));
	jdff dff_A_8KFNZSZn2_0(.dout(w_dff_A_6dCSBIm63_0),.din(w_dff_A_8KFNZSZn2_0),.clk(gclk));
	jdff dff_B_TbHt2NqS5_1(.din(n195),.dout(w_dff_B_TbHt2NqS5_1),.clk(gclk));
	jdff dff_B_NPWf3BlC9_1(.din(w_dff_B_TbHt2NqS5_1),.dout(w_dff_B_NPWf3BlC9_1),.clk(gclk));
	jdff dff_B_6ntJpehm7_1(.din(w_dff_B_NPWf3BlC9_1),.dout(w_dff_B_6ntJpehm7_1),.clk(gclk));
	jdff dff_B_BYdBkM1K9_1(.din(w_dff_B_6ntJpehm7_1),.dout(w_dff_B_BYdBkM1K9_1),.clk(gclk));
	jdff dff_A_bfFYFjT90_1(.dout(w_n194_0[1]),.din(w_dff_A_bfFYFjT90_1),.clk(gclk));
	jdff dff_A_va8DJXVj6_1(.dout(w_dff_A_bfFYFjT90_1),.din(w_dff_A_va8DJXVj6_1),.clk(gclk));
	jdff dff_A_nL852zRF6_1(.dout(w_dff_A_va8DJXVj6_1),.din(w_dff_A_nL852zRF6_1),.clk(gclk));
	jdff dff_A_lZsuws234_1(.dout(w_dff_A_nL852zRF6_1),.din(w_dff_A_lZsuws234_1),.clk(gclk));
	jdff dff_B_I9MtPv5B2_0(.din(n271),.dout(w_dff_B_I9MtPv5B2_0),.clk(gclk));
	jdff dff_B_aRKeSmgl0_0(.din(w_dff_B_I9MtPv5B2_0),.dout(w_dff_B_aRKeSmgl0_0),.clk(gclk));
	jdff dff_B_LGC1z6e52_0(.din(w_dff_B_aRKeSmgl0_0),.dout(w_dff_B_LGC1z6e52_0),.clk(gclk));
	jdff dff_B_OqDX1mhE5_0(.din(w_dff_B_LGC1z6e52_0),.dout(w_dff_B_OqDX1mhE5_0),.clk(gclk));
	jdff dff_B_JUgQGpSK3_0(.din(w_dff_B_OqDX1mhE5_0),.dout(w_dff_B_JUgQGpSK3_0),.clk(gclk));
	jdff dff_B_3PkoWrj11_0(.din(n269),.dout(w_dff_B_3PkoWrj11_0),.clk(gclk));
	jdff dff_B_GiAlbKGp3_0(.din(w_dff_B_3PkoWrj11_0),.dout(w_dff_B_GiAlbKGp3_0),.clk(gclk));
	jdff dff_B_rOr14aHw5_0(.din(w_dff_B_GiAlbKGp3_0),.dout(w_dff_B_rOr14aHw5_0),.clk(gclk));
	jdff dff_B_dY8HKWI11_0(.din(n263),.dout(w_dff_B_dY8HKWI11_0),.clk(gclk));
	jdff dff_B_tnMSyusZ3_0(.din(w_dff_B_dY8HKWI11_0),.dout(w_dff_B_tnMSyusZ3_0),.clk(gclk));
	jdff dff_B_UlJzRGsu9_0(.din(w_dff_B_tnMSyusZ3_0),.dout(w_dff_B_UlJzRGsu9_0),.clk(gclk));
	jdff dff_B_uQZJAPKj9_0(.din(w_dff_B_UlJzRGsu9_0),.dout(w_dff_B_uQZJAPKj9_0),.clk(gclk));
	jdff dff_B_AeskRH0b2_0(.din(w_dff_B_uQZJAPKj9_0),.dout(w_dff_B_AeskRH0b2_0),.clk(gclk));
	jdff dff_B_Ao5ed7Sc2_0(.din(w_dff_B_AeskRH0b2_0),.dout(w_dff_B_Ao5ed7Sc2_0),.clk(gclk));
	jdff dff_B_3rQfalH84_1(.din(n253),.dout(w_dff_B_3rQfalH84_1),.clk(gclk));
	jdff dff_B_NQ4RqetA0_1(.din(w_dff_B_3rQfalH84_1),.dout(w_dff_B_NQ4RqetA0_1),.clk(gclk));
	jdff dff_B_hbzpXksv7_1(.din(w_dff_B_NQ4RqetA0_1),.dout(w_dff_B_hbzpXksv7_1),.clk(gclk));
	jdff dff_B_foePtHae1_1(.din(w_dff_B_hbzpXksv7_1),.dout(w_dff_B_foePtHae1_1),.clk(gclk));
	jdff dff_A_J2nYIFC01_1(.dout(w_n252_0[1]),.din(w_dff_A_J2nYIFC01_1),.clk(gclk));
	jdff dff_A_LsLfIUFq4_1(.dout(w_dff_A_J2nYIFC01_1),.din(w_dff_A_LsLfIUFq4_1),.clk(gclk));
	jdff dff_A_aE2wYgBZ6_1(.dout(w_dff_A_LsLfIUFq4_1),.din(w_dff_A_aE2wYgBZ6_1),.clk(gclk));
	jdff dff_A_9h2QmdbG4_1(.dout(w_dff_A_aE2wYgBZ6_1),.din(w_dff_A_9h2QmdbG4_1),.clk(gclk));
	jdff dff_B_uQ49Dq5p5_0(.din(n289),.dout(w_dff_B_uQ49Dq5p5_0),.clk(gclk));
	jdff dff_B_M1Ue3DhB0_0(.din(w_dff_B_uQ49Dq5p5_0),.dout(w_dff_B_M1Ue3DhB0_0),.clk(gclk));
	jdff dff_B_1zNYJEzd3_0(.din(w_dff_B_M1Ue3DhB0_0),.dout(w_dff_B_1zNYJEzd3_0),.clk(gclk));
	jdff dff_B_QkcrlfEn9_0(.din(n287),.dout(w_dff_B_QkcrlfEn9_0),.clk(gclk));
	jdff dff_B_Lt1awlyo1_0(.din(w_dff_B_QkcrlfEn9_0),.dout(w_dff_B_Lt1awlyo1_0),.clk(gclk));
	jdff dff_B_m1dfGMgx5_0(.din(w_dff_B_Lt1awlyo1_0),.dout(w_dff_B_m1dfGMgx5_0),.clk(gclk));
	jdff dff_B_jiMhpmyk4_0(.din(n281),.dout(w_dff_B_jiMhpmyk4_0),.clk(gclk));
	jdff dff_B_MtZimH5r2_0(.din(w_dff_B_jiMhpmyk4_0),.dout(w_dff_B_MtZimH5r2_0),.clk(gclk));
	jdff dff_B_A0BDc1nC7_0(.din(w_dff_B_MtZimH5r2_0),.dout(w_dff_B_A0BDc1nC7_0),.clk(gclk));
	jdff dff_B_g681Yg8Y3_0(.din(w_dff_B_A0BDc1nC7_0),.dout(w_dff_B_g681Yg8Y3_0),.clk(gclk));
	jdff dff_B_I9IJunoj5_0(.din(w_dff_B_g681Yg8Y3_0),.dout(w_dff_B_I9IJunoj5_0),.clk(gclk));
	jdff dff_B_ldOh7XXr3_0(.din(w_dff_B_I9IJunoj5_0),.dout(w_dff_B_ldOh7XXr3_0),.clk(gclk));
	jdff dff_B_P392CBsC1_0(.din(n274),.dout(w_dff_B_P392CBsC1_0),.clk(gclk));
	jdff dff_B_aXzCb0vT9_0(.din(w_dff_B_P392CBsC1_0),.dout(w_dff_B_aXzCb0vT9_0),.clk(gclk));
	jdff dff_A_xEbT2sl02_1(.dout(w_n273_0[1]),.din(w_dff_A_xEbT2sl02_1),.clk(gclk));
	jdff dff_A_5y9cMeqJ6_1(.dout(w_dff_A_xEbT2sl02_1),.din(w_dff_A_5y9cMeqJ6_1),.clk(gclk));
	jdff dff_B_PSsVC57p9_1(.din(n300),.dout(w_dff_B_PSsVC57p9_1),.clk(gclk));
	jdff dff_B_wQUoV3cU7_1(.din(w_dff_B_PSsVC57p9_1),.dout(w_dff_B_wQUoV3cU7_1),.clk(gclk));
	jdff dff_B_lylyPlAQ1_1(.din(w_dff_B_wQUoV3cU7_1),.dout(w_dff_B_lylyPlAQ1_1),.clk(gclk));
	jdff dff_B_j70V6Zra1_1(.din(w_dff_B_lylyPlAQ1_1),.dout(w_dff_B_j70V6Zra1_1),.clk(gclk));
	jdff dff_B_iXPshyrT5_1(.din(w_dff_B_j70V6Zra1_1),.dout(w_dff_B_iXPshyrT5_1),.clk(gclk));
	jdff dff_B_pXv7gpGb6_1(.din(w_dff_B_iXPshyrT5_1),.dout(w_dff_B_pXv7gpGb6_1),.clk(gclk));
	jdff dff_B_T1LxtHyp1_1(.din(w_dff_B_pXv7gpGb6_1),.dout(w_dff_B_T1LxtHyp1_1),.clk(gclk));
	jdff dff_B_4CsWXpvl2_1(.din(w_dff_B_T1LxtHyp1_1),.dout(w_dff_B_4CsWXpvl2_1),.clk(gclk));
	jdff dff_B_9SCzL1PZ3_1(.din(w_dff_B_4CsWXpvl2_1),.dout(w_dff_B_9SCzL1PZ3_1),.clk(gclk));
	jdff dff_B_fePUdM2d9_1(.din(w_dff_B_9SCzL1PZ3_1),.dout(w_dff_B_fePUdM2d9_1),.clk(gclk));
	jdff dff_B_R5eBDsPA3_1(.din(n301),.dout(w_dff_B_R5eBDsPA3_1),.clk(gclk));
	jdff dff_B_Vd93AqSE0_1(.din(w_dff_B_R5eBDsPA3_1),.dout(w_dff_B_Vd93AqSE0_1),.clk(gclk));
	jdff dff_B_Q0SXByaK0_1(.din(w_dff_B_Vd93AqSE0_1),.dout(w_dff_B_Q0SXByaK0_1),.clk(gclk));
	jdff dff_B_U89kJPZY4_1(.din(w_dff_B_Q0SXByaK0_1),.dout(w_dff_B_U89kJPZY4_1),.clk(gclk));
	jdff dff_B_vj6QkmWj3_1(.din(w_dff_B_U89kJPZY4_1),.dout(w_dff_B_vj6QkmWj3_1),.clk(gclk));
	jdff dff_B_4wOsKy8P0_1(.din(w_dff_B_vj6QkmWj3_1),.dout(w_dff_B_4wOsKy8P0_1),.clk(gclk));
	jdff dff_B_ue63feuJ8_1(.din(w_dff_B_4wOsKy8P0_1),.dout(w_dff_B_ue63feuJ8_1),.clk(gclk));
	jdff dff_B_URtzJv2O8_1(.din(w_dff_B_ue63feuJ8_1),.dout(w_dff_B_URtzJv2O8_1),.clk(gclk));
	jdff dff_B_JqCAedvZ7_1(.din(w_dff_B_URtzJv2O8_1),.dout(w_dff_B_JqCAedvZ7_1),.clk(gclk));
	jdff dff_B_UUujBUAM7_0(.din(n361),.dout(w_dff_B_UUujBUAM7_0),.clk(gclk));
	jdff dff_B_cGkE6gFN0_0(.din(w_dff_B_UUujBUAM7_0),.dout(w_dff_B_cGkE6gFN0_0),.clk(gclk));
	jdff dff_B_IN4gHvf12_0(.din(w_dff_B_cGkE6gFN0_0),.dout(w_dff_B_IN4gHvf12_0),.clk(gclk));
	jdff dff_B_p39H8VW78_0(.din(w_dff_B_IN4gHvf12_0),.dout(w_dff_B_p39H8VW78_0),.clk(gclk));
	jdff dff_B_vqWrTDug0_0(.din(w_dff_B_p39H8VW78_0),.dout(w_dff_B_vqWrTDug0_0),.clk(gclk));
	jdff dff_B_PWPeztSQ1_0(.din(w_dff_B_vqWrTDug0_0),.dout(w_dff_B_PWPeztSQ1_0),.clk(gclk));
	jdff dff_B_vhlg5ahJ8_0(.din(w_dff_B_PWPeztSQ1_0),.dout(w_dff_B_vhlg5ahJ8_0),.clk(gclk));
	jdff dff_B_VGeWtE5A5_0(.din(w_dff_B_vhlg5ahJ8_0),.dout(w_dff_B_VGeWtE5A5_0),.clk(gclk));
	jdff dff_B_JKAPmDKw7_0(.din(n359),.dout(w_dff_B_JKAPmDKw7_0),.clk(gclk));
	jdff dff_B_F5qxVQDB4_0(.din(w_dff_B_JKAPmDKw7_0),.dout(w_dff_B_F5qxVQDB4_0),.clk(gclk));
	jdff dff_B_T5cTBSeb9_0(.din(n355),.dout(w_dff_B_T5cTBSeb9_0),.clk(gclk));
	jdff dff_B_1BZcYoJP2_0(.din(w_dff_B_T5cTBSeb9_0),.dout(w_dff_B_1BZcYoJP2_0),.clk(gclk));
	jdff dff_B_CUK6ySF87_0(.din(w_dff_B_1BZcYoJP2_0),.dout(w_dff_B_CUK6ySF87_0),.clk(gclk));
	jdff dff_B_QX469E8X6_0(.din(w_dff_B_CUK6ySF87_0),.dout(w_dff_B_QX469E8X6_0),.clk(gclk));
	jdff dff_B_KFCGK5jy3_0(.din(w_dff_B_QX469E8X6_0),.dout(w_dff_B_KFCGK5jy3_0),.clk(gclk));
	jdff dff_A_luHCqTH56_1(.dout(w_G228gat_2[1]),.din(w_dff_A_luHCqTH56_1),.clk(gclk));
	jdff dff_A_2q7bebE30_2(.dout(w_G228gat_2[2]),.din(w_dff_A_2q7bebE30_2),.clk(gclk));
	jdff dff_A_VrnR1Axb8_0(.dout(w_G219gat_2[0]),.din(w_dff_A_VrnR1Axb8_0),.clk(gclk));
	jdff dff_A_RBJldML08_0(.dout(w_dff_A_VrnR1Axb8_0),.din(w_dff_A_RBJldML08_0),.clk(gclk));
	jdff dff_A_XsGDrWzE2_0(.dout(w_dff_A_RBJldML08_0),.din(w_dff_A_XsGDrWzE2_0),.clk(gclk));
	jdff dff_A_CcZfl3DE9_0(.dout(w_dff_A_XsGDrWzE2_0),.din(w_dff_A_CcZfl3DE9_0),.clk(gclk));
	jdff dff_A_O4BnKZWH7_2(.dout(w_G219gat_2[2]),.din(w_dff_A_O4BnKZWH7_2),.clk(gclk));
	jdff dff_A_TjZN6dMJ0_2(.dout(w_dff_A_O4BnKZWH7_2),.din(w_dff_A_TjZN6dMJ0_2),.clk(gclk));
	jdff dff_B_PvelPzH93_0(.din(n348),.dout(w_dff_B_PvelPzH93_0),.clk(gclk));
	jdff dff_B_Cmgrk6HO6_0(.din(w_dff_B_PvelPzH93_0),.dout(w_dff_B_Cmgrk6HO6_0),.clk(gclk));
	jdff dff_B_OVo8ApWz2_0(.din(w_dff_B_Cmgrk6HO6_0),.dout(w_dff_B_OVo8ApWz2_0),.clk(gclk));
	jdff dff_B_NJi8DAPx1_0(.din(w_dff_B_OVo8ApWz2_0),.dout(w_dff_B_NJi8DAPx1_0),.clk(gclk));
	jdff dff_B_aMUOQhrM9_0(.din(w_dff_B_NJi8DAPx1_0),.dout(w_dff_B_aMUOQhrM9_0),.clk(gclk));
	jdff dff_B_BHvrKp0m4_0(.din(w_dff_B_aMUOQhrM9_0),.dout(w_dff_B_BHvrKp0m4_0),.clk(gclk));
	jdff dff_B_xzkYETx73_0(.din(w_dff_B_BHvrKp0m4_0),.dout(w_dff_B_xzkYETx73_0),.clk(gclk));
	jdff dff_A_3c1Tgmvu1_1(.dout(w_n347_0[1]),.din(w_dff_A_3c1Tgmvu1_1),.clk(gclk));
	jdff dff_A_1UTP8PLS0_1(.dout(w_dff_A_3c1Tgmvu1_1),.din(w_dff_A_1UTP8PLS0_1),.clk(gclk));
	jdff dff_A_jncO0Wt77_1(.dout(w_dff_A_1UTP8PLS0_1),.din(w_dff_A_jncO0Wt77_1),.clk(gclk));
	jdff dff_A_jkoQySE98_1(.dout(w_dff_A_jncO0Wt77_1),.din(w_dff_A_jkoQySE98_1),.clk(gclk));
	jdff dff_A_Rxk9jG7z0_1(.dout(w_dff_A_jkoQySE98_1),.din(w_dff_A_Rxk9jG7z0_1),.clk(gclk));
	jdff dff_A_o42z7cOD5_1(.dout(w_dff_A_Rxk9jG7z0_1),.din(w_dff_A_o42z7cOD5_1),.clk(gclk));
	jdff dff_A_fEwDBsn05_1(.dout(w_dff_A_o42z7cOD5_1),.din(w_dff_A_fEwDBsn05_1),.clk(gclk));
	jdff dff_B_ejuXkCzL1_0(.din(n381),.dout(w_dff_B_ejuXkCzL1_0),.clk(gclk));
	jdff dff_B_bKiJwjb46_0(.din(w_dff_B_ejuXkCzL1_0),.dout(w_dff_B_bKiJwjb46_0),.clk(gclk));
	jdff dff_B_Q5z9qhIY4_0(.din(w_dff_B_bKiJwjb46_0),.dout(w_dff_B_Q5z9qhIY4_0),.clk(gclk));
	jdff dff_B_YNtbvHhX4_0(.din(w_dff_B_Q5z9qhIY4_0),.dout(w_dff_B_YNtbvHhX4_0),.clk(gclk));
	jdff dff_B_vmSlP96T3_0(.din(w_dff_B_YNtbvHhX4_0),.dout(w_dff_B_vmSlP96T3_0),.clk(gclk));
	jdff dff_B_2lmFNbKq1_0(.din(w_dff_B_vmSlP96T3_0),.dout(w_dff_B_2lmFNbKq1_0),.clk(gclk));
	jdff dff_B_qcIiTrxY9_0(.din(w_dff_B_2lmFNbKq1_0),.dout(w_dff_B_qcIiTrxY9_0),.clk(gclk));
	jdff dff_B_XFRitF935_0(.din(w_dff_B_qcIiTrxY9_0),.dout(w_dff_B_XFRitF935_0),.clk(gclk));
	jdff dff_B_bg76ZjFb0_0(.din(w_dff_B_XFRitF935_0),.dout(w_dff_B_bg76ZjFb0_0),.clk(gclk));
	jdff dff_B_MP1MsEYv0_0(.din(w_dff_B_bg76ZjFb0_0),.dout(w_dff_B_MP1MsEYv0_0),.clk(gclk));
	jdff dff_B_svDJdJhT9_0(.din(n379),.dout(w_dff_B_svDJdJhT9_0),.clk(gclk));
	jdff dff_B_m7emHeOP8_0(.din(w_dff_B_svDJdJhT9_0),.dout(w_dff_B_m7emHeOP8_0),.clk(gclk));
	jdff dff_B_ojYVdEt22_0(.din(n375),.dout(w_dff_B_ojYVdEt22_0),.clk(gclk));
	jdff dff_B_eiDEt4M17_0(.din(w_dff_B_ojYVdEt22_0),.dout(w_dff_B_eiDEt4M17_0),.clk(gclk));
	jdff dff_B_EMEVQT7L2_0(.din(w_dff_B_eiDEt4M17_0),.dout(w_dff_B_EMEVQT7L2_0),.clk(gclk));
	jdff dff_B_UDtgVnD31_0(.din(w_dff_B_EMEVQT7L2_0),.dout(w_dff_B_UDtgVnD31_0),.clk(gclk));
	jdff dff_B_LpRmIxIQ1_0(.din(w_dff_B_UDtgVnD31_0),.dout(w_dff_B_LpRmIxIQ1_0),.clk(gclk));
	jdff dff_B_vZN3HOEM1_0(.din(n368),.dout(w_dff_B_vZN3HOEM1_0),.clk(gclk));
	jdff dff_B_2Xlx1w636_0(.din(w_dff_B_vZN3HOEM1_0),.dout(w_dff_B_2Xlx1w636_0),.clk(gclk));
	jdff dff_B_6WjvhTfD9_0(.din(w_dff_B_2Xlx1w636_0),.dout(w_dff_B_6WjvhTfD9_0),.clk(gclk));
	jdff dff_B_fvLSBqNQ5_0(.din(w_dff_B_6WjvhTfD9_0),.dout(w_dff_B_fvLSBqNQ5_0),.clk(gclk));
	jdff dff_B_7hexCDOk7_0(.din(w_dff_B_fvLSBqNQ5_0),.dout(w_dff_B_7hexCDOk7_0),.clk(gclk));
	jdff dff_B_lCNVQeRg1_0(.din(w_dff_B_7hexCDOk7_0),.dout(w_dff_B_lCNVQeRg1_0),.clk(gclk));
	jdff dff_B_4yYzpzQZ0_0(.din(w_dff_B_lCNVQeRg1_0),.dout(w_dff_B_4yYzpzQZ0_0),.clk(gclk));
	jdff dff_B_yhPNafJe5_0(.din(w_dff_B_4yYzpzQZ0_0),.dout(w_dff_B_yhPNafJe5_0),.clk(gclk));
	jdff dff_B_eYxYzzQE9_0(.din(w_dff_B_yhPNafJe5_0),.dout(w_dff_B_eYxYzzQE9_0),.clk(gclk));
	jdff dff_A_GrfYJCiC2_1(.dout(w_n367_0[1]),.din(w_dff_A_GrfYJCiC2_1),.clk(gclk));
	jdff dff_A_dLR0ShHf5_1(.dout(w_dff_A_GrfYJCiC2_1),.din(w_dff_A_dLR0ShHf5_1),.clk(gclk));
	jdff dff_A_1rqDsFLz1_1(.dout(w_dff_A_dLR0ShHf5_1),.din(w_dff_A_1rqDsFLz1_1),.clk(gclk));
	jdff dff_A_oW93ECL87_1(.dout(w_dff_A_1rqDsFLz1_1),.din(w_dff_A_oW93ECL87_1),.clk(gclk));
	jdff dff_A_T43GN7ZP0_1(.dout(w_dff_A_oW93ECL87_1),.din(w_dff_A_T43GN7ZP0_1),.clk(gclk));
	jdff dff_A_C6VHNfKB4_1(.dout(w_dff_A_T43GN7ZP0_1),.din(w_dff_A_C6VHNfKB4_1),.clk(gclk));
	jdff dff_A_BWmG1Y5r6_1(.dout(w_dff_A_C6VHNfKB4_1),.din(w_dff_A_BWmG1Y5r6_1),.clk(gclk));
	jdff dff_A_ekYEzkko1_1(.dout(w_dff_A_BWmG1Y5r6_1),.din(w_dff_A_ekYEzkko1_1),.clk(gclk));
	jdff dff_A_kL7E0WFL2_1(.dout(w_dff_A_ekYEzkko1_1),.din(w_dff_A_kL7E0WFL2_1),.clk(gclk));
	jdff dff_B_y8wriyGN7_1(.din(n294),.dout(w_dff_B_y8wriyGN7_1),.clk(gclk));
	jdff dff_B_gfoMCJij6_1(.din(w_dff_B_y8wriyGN7_1),.dout(w_dff_B_gfoMCJij6_1),.clk(gclk));
	jdff dff_B_9P1KBs8x2_1(.din(w_dff_B_gfoMCJij6_1),.dout(w_dff_B_9P1KBs8x2_1),.clk(gclk));
	jdff dff_B_upwepf7Q2_0(.din(n365),.dout(w_dff_B_upwepf7Q2_0),.clk(gclk));
	jdff dff_B_eRVd6BN99_0(.din(w_dff_B_upwepf7Q2_0),.dout(w_dff_B_eRVd6BN99_0),.clk(gclk));
	jdff dff_B_Eme59DSZ0_0(.din(w_dff_B_eRVd6BN99_0),.dout(w_dff_B_Eme59DSZ0_0),.clk(gclk));
	jdff dff_B_Mf8HV2vp2_0(.din(w_dff_B_Eme59DSZ0_0),.dout(w_dff_B_Mf8HV2vp2_0),.clk(gclk));
	jdff dff_A_hVABhXPc1_1(.dout(w_n339_0[1]),.din(w_dff_A_hVABhXPc1_1),.clk(gclk));
	jdff dff_A_vyIiVjNM8_1(.dout(w_dff_A_hVABhXPc1_1),.din(w_dff_A_vyIiVjNM8_1),.clk(gclk));
	jdff dff_A_solfsl5g8_1(.dout(w_dff_A_vyIiVjNM8_1),.din(w_dff_A_solfsl5g8_1),.clk(gclk));
	jdff dff_A_ZHpQrXdH1_1(.dout(w_dff_A_solfsl5g8_1),.din(w_dff_A_ZHpQrXdH1_1),.clk(gclk));
	jdff dff_B_uubR0MUS1_1(.din(n333),.dout(w_dff_B_uubR0MUS1_1),.clk(gclk));
	jdff dff_B_ML0mMVFQ9_1(.din(w_dff_B_uubR0MUS1_1),.dout(w_dff_B_ML0mMVFQ9_1),.clk(gclk));
	jdff dff_B_alhlfcJh7_1(.din(w_dff_B_ML0mMVFQ9_1),.dout(w_dff_B_alhlfcJh7_1),.clk(gclk));
	jdff dff_B_P7J20owu5_0(.din(n363),.dout(w_dff_B_P7J20owu5_0),.clk(gclk));
	jdff dff_B_eQtQQ3Um4_0(.din(w_dff_B_P7J20owu5_0),.dout(w_dff_B_eQtQQ3Um4_0),.clk(gclk));
	jdff dff_B_DRLhDGWM8_0(.din(w_dff_B_eQtQQ3Um4_0),.dout(w_dff_B_DRLhDGWM8_0),.clk(gclk));
	jdff dff_B_gdY9OzYR7_0(.din(w_dff_B_DRLhDGWM8_0),.dout(w_dff_B_gdY9OzYR7_0),.clk(gclk));
	jdff dff_A_qFlBrBPR0_1(.dout(w_n331_0[1]),.din(w_dff_A_qFlBrBPR0_1),.clk(gclk));
	jdff dff_A_4VrBza8N0_1(.dout(w_dff_A_qFlBrBPR0_1),.din(w_dff_A_4VrBza8N0_1),.clk(gclk));
	jdff dff_A_xwMSUpzW4_1(.dout(w_dff_A_4VrBza8N0_1),.din(w_dff_A_xwMSUpzW4_1),.clk(gclk));
	jdff dff_A_L4YyDJsW5_1(.dout(w_dff_A_xwMSUpzW4_1),.din(w_dff_A_L4YyDJsW5_1),.clk(gclk));
	jdff dff_B_VfiQu5VF8_1(.din(n306),.dout(w_dff_B_VfiQu5VF8_1),.clk(gclk));
	jdff dff_B_vuEUIjCo5_1(.din(w_dff_B_VfiQu5VF8_1),.dout(w_dff_B_vuEUIjCo5_1),.clk(gclk));
	jdff dff_B_isoGcj515_1(.din(w_dff_B_vuEUIjCo5_1),.dout(w_dff_B_isoGcj515_1),.clk(gclk));
	jdff dff_B_qrL2tGue6_1(.din(w_dff_B_isoGcj515_1),.dout(w_dff_B_qrL2tGue6_1),.clk(gclk));
	jdff dff_B_SwdrMDr66_1(.din(w_dff_B_qrL2tGue6_1),.dout(w_dff_B_SwdrMDr66_1),.clk(gclk));
	jdff dff_B_UkOoVVom8_1(.din(w_dff_B_SwdrMDr66_1),.dout(w_dff_B_UkOoVVom8_1),.clk(gclk));
	jdff dff_B_2AmxpU0q8_1(.din(w_dff_B_UkOoVVom8_1),.dout(w_dff_B_2AmxpU0q8_1),.clk(gclk));
	jdff dff_B_hwq3fEWR7_0(.din(n403),.dout(w_dff_B_hwq3fEWR7_0),.clk(gclk));
	jdff dff_B_PHn4Iqm46_0(.din(w_dff_B_hwq3fEWR7_0),.dout(w_dff_B_PHn4Iqm46_0),.clk(gclk));
	jdff dff_B_n4kuRFsg9_0(.din(w_dff_B_PHn4Iqm46_0),.dout(w_dff_B_n4kuRFsg9_0),.clk(gclk));
	jdff dff_B_kmGwrkYe2_0(.din(w_dff_B_n4kuRFsg9_0),.dout(w_dff_B_kmGwrkYe2_0),.clk(gclk));
	jdff dff_B_ccCIEoik0_0(.din(w_dff_B_kmGwrkYe2_0),.dout(w_dff_B_ccCIEoik0_0),.clk(gclk));
	jdff dff_B_mWTTLcnW4_0(.din(w_dff_B_ccCIEoik0_0),.dout(w_dff_B_mWTTLcnW4_0),.clk(gclk));
	jdff dff_B_nVWtyN8D2_0(.din(w_dff_B_mWTTLcnW4_0),.dout(w_dff_B_nVWtyN8D2_0),.clk(gclk));
	jdff dff_B_S0Dezss19_0(.din(w_dff_B_nVWtyN8D2_0),.dout(w_dff_B_S0Dezss19_0),.clk(gclk));
	jdff dff_B_PrfmrOam4_0(.din(w_dff_B_S0Dezss19_0),.dout(w_dff_B_PrfmrOam4_0),.clk(gclk));
	jdff dff_B_JZYJZQ1Q8_0(.din(w_dff_B_PrfmrOam4_0),.dout(w_dff_B_JZYJZQ1Q8_0),.clk(gclk));
	jdff dff_B_yIxaJxKJ8_0(.din(n401),.dout(w_dff_B_yIxaJxKJ8_0),.clk(gclk));
	jdff dff_B_3BozDWWg7_0(.din(w_dff_B_yIxaJxKJ8_0),.dout(w_dff_B_3BozDWWg7_0),.clk(gclk));
	jdff dff_B_b9FJPlqP8_0(.din(n397),.dout(w_dff_B_b9FJPlqP8_0),.clk(gclk));
	jdff dff_B_YN5GQ3cq7_0(.din(w_dff_B_b9FJPlqP8_0),.dout(w_dff_B_YN5GQ3cq7_0),.clk(gclk));
	jdff dff_B_mFMOqZYj2_0(.din(w_dff_B_YN5GQ3cq7_0),.dout(w_dff_B_mFMOqZYj2_0),.clk(gclk));
	jdff dff_B_AJSJfjBV2_0(.din(w_dff_B_mFMOqZYj2_0),.dout(w_dff_B_AJSJfjBV2_0),.clk(gclk));
	jdff dff_B_ABwgDkzj8_0(.din(w_dff_B_AJSJfjBV2_0),.dout(w_dff_B_ABwgDkzj8_0),.clk(gclk));
	jdff dff_B_Hu4cH0Rk2_1(.din(n384),.dout(w_dff_B_Hu4cH0Rk2_1),.clk(gclk));
	jdff dff_B_fon8S6i46_1(.din(w_dff_B_Hu4cH0Rk2_1),.dout(w_dff_B_fon8S6i46_1),.clk(gclk));
	jdff dff_B_PpU2OFFW9_1(.din(w_dff_B_fon8S6i46_1),.dout(w_dff_B_PpU2OFFW9_1),.clk(gclk));
	jdff dff_B_e1SyOF1o5_1(.din(w_dff_B_PpU2OFFW9_1),.dout(w_dff_B_e1SyOF1o5_1),.clk(gclk));
	jdff dff_B_bNLJoKfB2_1(.din(w_dff_B_e1SyOF1o5_1),.dout(w_dff_B_bNLJoKfB2_1),.clk(gclk));
	jdff dff_B_cmLMnqV32_1(.din(w_dff_B_bNLJoKfB2_1),.dout(w_dff_B_cmLMnqV32_1),.clk(gclk));
	jdff dff_B_T59eWlDD7_1(.din(w_dff_B_cmLMnqV32_1),.dout(w_dff_B_T59eWlDD7_1),.clk(gclk));
	jdff dff_B_fI27sppI3_1(.din(w_dff_B_T59eWlDD7_1),.dout(w_dff_B_fI27sppI3_1),.clk(gclk));
	jdff dff_B_gYOXGW2O2_1(.din(w_dff_B_fI27sppI3_1),.dout(w_dff_B_gYOXGW2O2_1),.clk(gclk));
	jdff dff_B_bSf97WbI8_1(.din(n385),.dout(w_dff_B_bSf97WbI8_1),.clk(gclk));
	jdff dff_B_r0hEydaL2_1(.din(w_dff_B_bSf97WbI8_1),.dout(w_dff_B_r0hEydaL2_1),.clk(gclk));
	jdff dff_B_IuBiekTt3_1(.din(w_dff_B_r0hEydaL2_1),.dout(w_dff_B_IuBiekTt3_1),.clk(gclk));
	jdff dff_B_8NxEq6dq0_1(.din(w_dff_B_IuBiekTt3_1),.dout(w_dff_B_8NxEq6dq0_1),.clk(gclk));
	jdff dff_B_Xed15cmI5_1(.din(w_dff_B_8NxEq6dq0_1),.dout(w_dff_B_Xed15cmI5_1),.clk(gclk));
	jdff dff_B_1pNGs2sO1_1(.din(w_dff_B_Xed15cmI5_1),.dout(w_dff_B_1pNGs2sO1_1),.clk(gclk));
	jdff dff_B_j2CIVh7K0_0(.din(n386),.dout(w_dff_B_j2CIVh7K0_0),.clk(gclk));
	jdff dff_B_2HDtAj3D3_0(.din(w_dff_B_j2CIVh7K0_0),.dout(w_dff_B_2HDtAj3D3_0),.clk(gclk));
	jdff dff_B_FREj439S2_0(.din(w_dff_B_2HDtAj3D3_0),.dout(w_dff_B_FREj439S2_0),.clk(gclk));
	jdff dff_B_mltqWTru1_0(.din(w_dff_B_FREj439S2_0),.dout(w_dff_B_mltqWTru1_0),.clk(gclk));
	jdff dff_B_LCW2ZACj5_0(.din(w_dff_B_mltqWTru1_0),.dout(w_dff_B_LCW2ZACj5_0),.clk(gclk));
	jdff dff_B_2kkwxVAz8_0(.din(w_dff_B_LCW2ZACj5_0),.dout(w_dff_B_2kkwxVAz8_0),.clk(gclk));
	jdff dff_A_CJMAzMeI6_0(.dout(w_n330_0[0]),.din(w_dff_A_CJMAzMeI6_0),.clk(gclk));
	jdff dff_A_7S7PtQTf3_0(.dout(w_dff_A_CJMAzMeI6_0),.din(w_dff_A_7S7PtQTf3_0),.clk(gclk));
	jdff dff_A_VZb0BmbH8_0(.dout(w_dff_A_7S7PtQTf3_0),.din(w_dff_A_VZb0BmbH8_0),.clk(gclk));
	jdff dff_A_p6whfGDb1_0(.dout(w_dff_A_VZb0BmbH8_0),.din(w_dff_A_p6whfGDb1_0),.clk(gclk));
	jdff dff_A_zAVijECk6_0(.dout(w_dff_A_p6whfGDb1_0),.din(w_dff_A_zAVijECk6_0),.clk(gclk));
	jdff dff_A_fJznWadX8_0(.dout(w_dff_A_zAVijECk6_0),.din(w_dff_A_fJznWadX8_0),.clk(gclk));
	jdff dff_A_Zqdv1tL21_2(.dout(w_n330_0[2]),.din(w_dff_A_Zqdv1tL21_2),.clk(gclk));
	jdff dff_A_PX2pQ23d1_0(.dout(w_n337_0[0]),.din(w_dff_A_PX2pQ23d1_0),.clk(gclk));
	jdff dff_A_6xDU2RAL3_0(.dout(w_dff_A_PX2pQ23d1_0),.din(w_dff_A_6xDU2RAL3_0),.clk(gclk));
	jdff dff_A_mIMn5Ykv7_0(.dout(w_dff_A_6xDU2RAL3_0),.din(w_dff_A_mIMn5Ykv7_0),.clk(gclk));
	jdff dff_A_i2NJ4g9z3_0(.dout(w_dff_A_mIMn5Ykv7_0),.din(w_dff_A_i2NJ4g9z3_0),.clk(gclk));
	jdff dff_A_4QpLVSIA6_0(.dout(w_dff_A_i2NJ4g9z3_0),.din(w_dff_A_4QpLVSIA6_0),.clk(gclk));
	jdff dff_A_W2JSlw2h6_0(.dout(w_dff_A_4QpLVSIA6_0),.din(w_dff_A_W2JSlw2h6_0),.clk(gclk));
	jdff dff_B_G0UghCva0_1(.din(n334),.dout(w_dff_B_G0UghCva0_1),.clk(gclk));
	jdff dff_A_1HZBh8Na0_1(.dout(w_n383_0[1]),.din(w_dff_A_1HZBh8Na0_1),.clk(gclk));
	jdff dff_A_6iWupodD4_1(.dout(w_dff_A_1HZBh8Na0_1),.din(w_dff_A_6iWupodD4_1),.clk(gclk));
	jdff dff_A_yGMIvI1r9_1(.dout(w_dff_A_6iWupodD4_1),.din(w_dff_A_yGMIvI1r9_1),.clk(gclk));
	jdff dff_A_5KNnb36o7_1(.dout(w_dff_A_yGMIvI1r9_1),.din(w_dff_A_5KNnb36o7_1),.clk(gclk));
	jdff dff_A_tOGmhFl81_1(.dout(w_dff_A_5KNnb36o7_1),.din(w_dff_A_tOGmhFl81_1),.clk(gclk));
	jdff dff_A_t5U60hl49_1(.dout(w_dff_A_tOGmhFl81_1),.din(w_dff_A_t5U60hl49_1),.clk(gclk));
	jdff dff_A_DldUsMtM4_1(.dout(w_dff_A_t5U60hl49_1),.din(w_dff_A_DldUsMtM4_1),.clk(gclk));
	jdff dff_A_PBhRjxzY1_1(.dout(w_dff_A_DldUsMtM4_1),.din(w_dff_A_PBhRjxzY1_1),.clk(gclk));
	jdff dff_A_YRxUrohg1_1(.dout(w_dff_A_PBhRjxzY1_1),.din(w_dff_A_YRxUrohg1_1),.clk(gclk));
	jdff dff_B_DK7amLpv3_0(.din(n309),.dout(w_dff_B_DK7amLpv3_0),.clk(gclk));
	jdff dff_B_WgmeGV823_0(.din(w_dff_B_DK7amLpv3_0),.dout(w_dff_B_WgmeGV823_0),.clk(gclk));
	jdff dff_B_G5GWcALe2_0(.din(w_dff_B_WgmeGV823_0),.dout(w_dff_B_G5GWcALe2_0),.clk(gclk));
	jdff dff_B_56rvIfWm8_0(.din(n425),.dout(w_dff_B_56rvIfWm8_0),.clk(gclk));
	jdff dff_B_AuPtzbiz8_0(.din(w_dff_B_56rvIfWm8_0),.dout(w_dff_B_AuPtzbiz8_0),.clk(gclk));
	jdff dff_B_Dzq5giEZ1_0(.din(w_dff_B_AuPtzbiz8_0),.dout(w_dff_B_Dzq5giEZ1_0),.clk(gclk));
	jdff dff_B_CUU6JaBF5_0(.din(w_dff_B_Dzq5giEZ1_0),.dout(w_dff_B_CUU6JaBF5_0),.clk(gclk));
	jdff dff_B_WflL3jgp8_0(.din(w_dff_B_CUU6JaBF5_0),.dout(w_dff_B_WflL3jgp8_0),.clk(gclk));
	jdff dff_B_8s6KdjQ07_0(.din(w_dff_B_WflL3jgp8_0),.dout(w_dff_B_8s6KdjQ07_0),.clk(gclk));
	jdff dff_B_VibIDv318_0(.din(w_dff_B_8s6KdjQ07_0),.dout(w_dff_B_VibIDv318_0),.clk(gclk));
	jdff dff_B_xS3NSyC90_0(.din(w_dff_B_VibIDv318_0),.dout(w_dff_B_xS3NSyC90_0),.clk(gclk));
	jdff dff_B_FdZQ15pz5_0(.din(w_dff_B_xS3NSyC90_0),.dout(w_dff_B_FdZQ15pz5_0),.clk(gclk));
	jdff dff_B_eLkANbUv5_0(.din(w_dff_B_FdZQ15pz5_0),.dout(w_dff_B_eLkANbUv5_0),.clk(gclk));
	jdff dff_B_UPm6L9Nb8_0(.din(n423),.dout(w_dff_B_UPm6L9Nb8_0),.clk(gclk));
	jdff dff_B_YkSpfOp92_0(.din(w_dff_B_UPm6L9Nb8_0),.dout(w_dff_B_YkSpfOp92_0),.clk(gclk));
	jdff dff_B_vJbsKFLG4_0(.din(n419),.dout(w_dff_B_vJbsKFLG4_0),.clk(gclk));
	jdff dff_B_vYiQ7NLk9_0(.din(w_dff_B_vJbsKFLG4_0),.dout(w_dff_B_vYiQ7NLk9_0),.clk(gclk));
	jdff dff_B_V0vRGvgv4_0(.din(w_dff_B_vYiQ7NLk9_0),.dout(w_dff_B_V0vRGvgv4_0),.clk(gclk));
	jdff dff_B_zOsGNssi7_0(.din(w_dff_B_V0vRGvgv4_0),.dout(w_dff_B_zOsGNssi7_0),.clk(gclk));
	jdff dff_B_YpYObPOD1_0(.din(w_dff_B_zOsGNssi7_0),.dout(w_dff_B_YpYObPOD1_0),.clk(gclk));
	jdff dff_A_2iPPdsSE7_2(.dout(w_G228gat_0[2]),.din(w_dff_A_2iPPdsSE7_2),.clk(gclk));
	jdff dff_B_zwgj93p76_3(.din(G228gat),.dout(w_dff_B_zwgj93p76_3),.clk(gclk));
	jdff dff_B_PFAMbxko0_3(.din(w_dff_B_zwgj93p76_3),.dout(w_dff_B_PFAMbxko0_3),.clk(gclk));
	jdff dff_B_MlU0lAIp0_3(.din(w_dff_B_PFAMbxko0_3),.dout(w_dff_B_MlU0lAIp0_3),.clk(gclk));
	jdff dff_B_GIhP74Wg6_3(.din(w_dff_B_MlU0lAIp0_3),.dout(w_dff_B_GIhP74Wg6_3),.clk(gclk));
	jdff dff_B_pRq8GCv18_3(.din(w_dff_B_GIhP74Wg6_3),.dout(w_dff_B_pRq8GCv18_3),.clk(gclk));
	jdff dff_B_UpjKneK80_3(.din(w_dff_B_pRq8GCv18_3),.dout(w_dff_B_UpjKneK80_3),.clk(gclk));
	jdff dff_B_UJIi8sLE4_3(.din(w_dff_B_UpjKneK80_3),.dout(w_dff_B_UJIi8sLE4_3),.clk(gclk));
	jdff dff_B_OJh4kz4m2_3(.din(w_dff_B_UJIi8sLE4_3),.dout(w_dff_B_OJh4kz4m2_3),.clk(gclk));
	jdff dff_A_Jr3fhXse1_0(.dout(w_G219gat_0[0]),.din(w_dff_A_Jr3fhXse1_0),.clk(gclk));
	jdff dff_A_Vlh8o8fC9_0(.dout(w_dff_A_Jr3fhXse1_0),.din(w_dff_A_Vlh8o8fC9_0),.clk(gclk));
	jdff dff_A_Qa9NDiWx3_0(.dout(w_dff_A_Vlh8o8fC9_0),.din(w_dff_A_Qa9NDiWx3_0),.clk(gclk));
	jdff dff_A_WmBEmp6c2_0(.dout(w_dff_A_Qa9NDiWx3_0),.din(w_dff_A_WmBEmp6c2_0),.clk(gclk));
	jdff dff_A_dF3Xy1lW9_0(.dout(w_dff_A_WmBEmp6c2_0),.din(w_dff_A_dF3Xy1lW9_0),.clk(gclk));
	jdff dff_A_T72zKEQs2_0(.dout(w_dff_A_dF3Xy1lW9_0),.din(w_dff_A_T72zKEQs2_0),.clk(gclk));
	jdff dff_A_1HEjBh4a1_0(.dout(w_dff_A_T72zKEQs2_0),.din(w_dff_A_1HEjBh4a1_0),.clk(gclk));
	jdff dff_A_abCT3wmx7_0(.dout(w_dff_A_1HEjBh4a1_0),.din(w_dff_A_abCT3wmx7_0),.clk(gclk));
	jdff dff_A_X5vUCZ1M2_1(.dout(w_G219gat_0[1]),.din(w_dff_A_X5vUCZ1M2_1),.clk(gclk));
	jdff dff_A_PKbnaw7G5_1(.dout(w_dff_A_X5vUCZ1M2_1),.din(w_dff_A_PKbnaw7G5_1),.clk(gclk));
	jdff dff_B_iQVI2BKV5_3(.din(G219gat),.dout(w_dff_B_iQVI2BKV5_3),.clk(gclk));
	jdff dff_B_iMK9Mlu16_3(.din(w_dff_B_iQVI2BKV5_3),.dout(w_dff_B_iMK9Mlu16_3),.clk(gclk));
	jdff dff_B_kW14EWci6_3(.din(w_dff_B_iMK9Mlu16_3),.dout(w_dff_B_kW14EWci6_3),.clk(gclk));
	jdff dff_B_8Ndi1Zxq2_3(.din(w_dff_B_kW14EWci6_3),.dout(w_dff_B_8Ndi1Zxq2_3),.clk(gclk));
	jdff dff_B_E0elwhjG7_3(.din(w_dff_B_8Ndi1Zxq2_3),.dout(w_dff_B_E0elwhjG7_3),.clk(gclk));
	jdff dff_B_6UNO9qem1_3(.din(w_dff_B_E0elwhjG7_3),.dout(w_dff_B_6UNO9qem1_3),.clk(gclk));
	jdff dff_B_tbx6iKZj6_3(.din(w_dff_B_6UNO9qem1_3),.dout(w_dff_B_tbx6iKZj6_3),.clk(gclk));
	jdff dff_B_83iLidIz6_3(.din(w_dff_B_tbx6iKZj6_3),.dout(w_dff_B_83iLidIz6_3),.clk(gclk));
	jdff dff_B_euJtAYGL1_3(.din(w_dff_B_83iLidIz6_3),.dout(w_dff_B_euJtAYGL1_3),.clk(gclk));
	jdff dff_B_crlZpAfE1_3(.din(w_dff_B_euJtAYGL1_3),.dout(w_dff_B_crlZpAfE1_3),.clk(gclk));
	jdff dff_B_rKiurHBS4_1(.din(n406),.dout(w_dff_B_rKiurHBS4_1),.clk(gclk));
	jdff dff_B_9RCMHPBu0_1(.din(w_dff_B_rKiurHBS4_1),.dout(w_dff_B_9RCMHPBu0_1),.clk(gclk));
	jdff dff_B_RPZmQoZr1_1(.din(w_dff_B_9RCMHPBu0_1),.dout(w_dff_B_RPZmQoZr1_1),.clk(gclk));
	jdff dff_B_GXLj3m6L1_1(.din(w_dff_B_RPZmQoZr1_1),.dout(w_dff_B_GXLj3m6L1_1),.clk(gclk));
	jdff dff_B_qqUZXOxh3_1(.din(w_dff_B_GXLj3m6L1_1),.dout(w_dff_B_qqUZXOxh3_1),.clk(gclk));
	jdff dff_B_8CjKssne5_1(.din(w_dff_B_qqUZXOxh3_1),.dout(w_dff_B_8CjKssne5_1),.clk(gclk));
	jdff dff_B_EG4wx0MW6_1(.din(w_dff_B_8CjKssne5_1),.dout(w_dff_B_EG4wx0MW6_1),.clk(gclk));
	jdff dff_B_9yVDhpBE8_1(.din(w_dff_B_EG4wx0MW6_1),.dout(w_dff_B_9yVDhpBE8_1),.clk(gclk));
	jdff dff_B_fAWAZmko4_1(.din(w_dff_B_9yVDhpBE8_1),.dout(w_dff_B_fAWAZmko4_1),.clk(gclk));
	jdff dff_B_vNRUB94I4_1(.din(n407),.dout(w_dff_B_vNRUB94I4_1),.clk(gclk));
	jdff dff_B_lleVSr7Z3_1(.din(w_dff_B_vNRUB94I4_1),.dout(w_dff_B_lleVSr7Z3_1),.clk(gclk));
	jdff dff_B_PnvaJQoS7_1(.din(w_dff_B_lleVSr7Z3_1),.dout(w_dff_B_PnvaJQoS7_1),.clk(gclk));
	jdff dff_B_TkBfJ3cD3_1(.din(w_dff_B_PnvaJQoS7_1),.dout(w_dff_B_TkBfJ3cD3_1),.clk(gclk));
	jdff dff_B_pK3Xx1Um6_1(.din(w_dff_B_TkBfJ3cD3_1),.dout(w_dff_B_pK3Xx1Um6_1),.clk(gclk));
	jdff dff_B_2mhOtTAv5_1(.din(w_dff_B_pK3Xx1Um6_1),.dout(w_dff_B_2mhOtTAv5_1),.clk(gclk));
	jdff dff_B_YDpaFihz6_1(.din(w_dff_B_2mhOtTAv5_1),.dout(w_dff_B_YDpaFihz6_1),.clk(gclk));
	jdff dff_B_iwS0WEyB8_1(.din(w_dff_B_YDpaFihz6_1),.dout(w_dff_B_iwS0WEyB8_1),.clk(gclk));
	jdff dff_B_oOj2Bofp5_0(.din(n408),.dout(w_dff_B_oOj2Bofp5_0),.clk(gclk));
	jdff dff_B_bMtc4hSB2_0(.din(w_dff_B_oOj2Bofp5_0),.dout(w_dff_B_bMtc4hSB2_0),.clk(gclk));
	jdff dff_B_2Wlz6Qyp1_0(.din(w_dff_B_bMtc4hSB2_0),.dout(w_dff_B_2Wlz6Qyp1_0),.clk(gclk));
	jdff dff_B_FNv6dQcA5_0(.din(w_dff_B_2Wlz6Qyp1_0),.dout(w_dff_B_FNv6dQcA5_0),.clk(gclk));
	jdff dff_B_7ByjNhWa2_0(.din(w_dff_B_FNv6dQcA5_0),.dout(w_dff_B_7ByjNhWa2_0),.clk(gclk));
	jdff dff_B_iPAFNaLz0_0(.din(w_dff_B_7ByjNhWa2_0),.dout(w_dff_B_iPAFNaLz0_0),.clk(gclk));
	jdff dff_B_H7X158O22_0(.din(w_dff_B_iPAFNaLz0_0),.dout(w_dff_B_H7X158O22_0),.clk(gclk));
	jdff dff_A_bIRNQoO69_0(.dout(w_n329_0[0]),.din(w_dff_A_bIRNQoO69_0),.clk(gclk));
	jdff dff_A_lqDPTkFj9_0(.dout(w_dff_A_bIRNQoO69_0),.din(w_dff_A_lqDPTkFj9_0),.clk(gclk));
	jdff dff_A_hym8EBkO5_0(.dout(w_dff_A_lqDPTkFj9_0),.din(w_dff_A_hym8EBkO5_0),.clk(gclk));
	jdff dff_A_wiOTDdMU4_0(.dout(w_dff_A_hym8EBkO5_0),.din(w_dff_A_wiOTDdMU4_0),.clk(gclk));
	jdff dff_A_UAmYFGzt6_0(.dout(w_dff_A_wiOTDdMU4_0),.din(w_dff_A_UAmYFGzt6_0),.clk(gclk));
	jdff dff_A_BRY6iDHA5_0(.dout(w_dff_A_UAmYFGzt6_0),.din(w_dff_A_BRY6iDHA5_0),.clk(gclk));
	jdff dff_A_0Pnsip6t7_0(.dout(w_dff_A_BRY6iDHA5_0),.din(w_dff_A_0Pnsip6t7_0),.clk(gclk));
	jdff dff_B_wDYsnYMr6_1(.din(n343),.dout(w_dff_B_wDYsnYMr6_1),.clk(gclk));
	jdff dff_B_l2eRCyw20_1(.din(w_dff_B_wDYsnYMr6_1),.dout(w_dff_B_l2eRCyw20_1),.clk(gclk));
	jdff dff_B_hTzLZthE4_1(.din(w_dff_B_l2eRCyw20_1),.dout(w_dff_B_hTzLZthE4_1),.clk(gclk));
	jdff dff_B_mcSFyEiD8_1(.din(w_dff_B_hTzLZthE4_1),.dout(w_dff_B_mcSFyEiD8_1),.clk(gclk));
	jdff dff_B_XPX9zK4e7_1(.din(w_dff_B_mcSFyEiD8_1),.dout(w_dff_B_XPX9zK4e7_1),.clk(gclk));
	jdff dff_B_H6xxC1vQ8_1(.din(n344),.dout(w_dff_B_H6xxC1vQ8_1),.clk(gclk));
	jdff dff_B_nojOaqla9_1(.din(w_dff_B_H6xxC1vQ8_1),.dout(w_dff_B_nojOaqla9_1),.clk(gclk));
	jdff dff_B_NTnOmrvD6_1(.din(w_dff_B_nojOaqla9_1),.dout(w_dff_B_NTnOmrvD6_1),.clk(gclk));
	jdff dff_B_e3KOWU6d5_1(.din(w_dff_B_NTnOmrvD6_1),.dout(w_dff_B_e3KOWU6d5_1),.clk(gclk));
	jdff dff_B_tOdDF97N7_0(.din(n231),.dout(w_dff_B_tOdDF97N7_0),.clk(gclk));
	jdff dff_A_c7Ea73oJ2_0(.dout(w_n230_0[0]),.din(w_dff_A_c7Ea73oJ2_0),.clk(gclk));
	jdff dff_B_h7p1nVAO5_1(.din(n227),.dout(w_dff_B_h7p1nVAO5_1),.clk(gclk));
	jdff dff_A_SiQESX4O6_0(.dout(w_n228_0[0]),.din(w_dff_A_SiQESX4O6_0),.clk(gclk));
	jdff dff_A_UpHqMox65_0(.dout(w_dff_A_SiQESX4O6_0),.din(w_dff_A_UpHqMox65_0),.clk(gclk));
	jdff dff_A_mZPGkEJ34_0(.dout(w_dff_A_UpHqMox65_0),.din(w_dff_A_mZPGkEJ34_0),.clk(gclk));
	jdff dff_B_5bvhS0zr2_0(.din(n225),.dout(w_dff_B_5bvhS0zr2_0),.clk(gclk));
	jdff dff_A_d7IZQ9Sj4_0(.dout(w_n224_0[0]),.din(w_dff_A_d7IZQ9Sj4_0),.clk(gclk));
	jdff dff_A_duOlf6nd3_0(.dout(w_n223_0[0]),.din(w_dff_A_duOlf6nd3_0),.clk(gclk));
	jdff dff_A_kkq4hYOp2_0(.dout(w_dff_A_duOlf6nd3_0),.din(w_dff_A_kkq4hYOp2_0),.clk(gclk));
	jdff dff_B_RbD4gjqX9_1(.din(n219),.dout(w_dff_B_RbD4gjqX9_1),.clk(gclk));
	jdff dff_B_vLsphLcm4_1(.din(n214),.dout(w_dff_B_vLsphLcm4_1),.clk(gclk));
	jdff dff_A_PLo5IAVx8_1(.dout(w_G146gat_0[1]),.din(w_dff_A_PLo5IAVx8_1),.clk(gclk));
	jdff dff_B_aC6KNLd33_2(.din(G146gat),.dout(w_dff_B_aC6KNLd33_2),.clk(gclk));
	jdff dff_B_gRcQL1DW6_2(.din(w_dff_B_aC6KNLd33_2),.dout(w_dff_B_gRcQL1DW6_2),.clk(gclk));
	jdff dff_B_HVnYHxUt3_2(.din(w_dff_B_gRcQL1DW6_2),.dout(w_dff_B_HVnYHxUt3_2),.clk(gclk));
	jdff dff_B_w4396kB92_2(.din(w_dff_B_HVnYHxUt3_2),.dout(w_dff_B_w4396kB92_2),.clk(gclk));
	jdff dff_B_Wdi97rtg3_1(.din(n197),.dout(w_dff_B_Wdi97rtg3_1),.clk(gclk));
	jdff dff_B_lqDVT3hF7_1(.din(n198),.dout(w_dff_B_lqDVT3hF7_1),.clk(gclk));
	jdff dff_B_vqBT7hkr8_1(.din(w_dff_B_lqDVT3hF7_1),.dout(w_dff_B_vqBT7hkr8_1),.clk(gclk));
	jdff dff_B_zNfywTMl3_1(.din(w_dff_B_vqBT7hkr8_1),.dout(w_dff_B_zNfywTMl3_1),.clk(gclk));
	jdff dff_B_kowgTTZz9_1(.din(w_dff_B_zNfywTMl3_1),.dout(w_dff_B_kowgTTZz9_1),.clk(gclk));
	jdff dff_B_Ol54VBa21_1(.din(w_dff_B_kowgTTZz9_1),.dout(w_dff_B_Ol54VBa21_1),.clk(gclk));
	jdff dff_B_v8lsR8PJ8_1(.din(w_dff_B_Ol54VBa21_1),.dout(w_dff_B_v8lsR8PJ8_1),.clk(gclk));
	jdff dff_B_6bYBhQ8m1_1(.din(w_dff_B_v8lsR8PJ8_1),.dout(w_dff_B_6bYBhQ8m1_1),.clk(gclk));
	jdff dff_B_Cy5q0l5Q0_1(.din(w_dff_B_6bYBhQ8m1_1),.dout(w_dff_B_Cy5q0l5Q0_1),.clk(gclk));
	jdff dff_B_00CMSlPU3_1(.din(n199),.dout(w_dff_B_00CMSlPU3_1),.clk(gclk));
	jdff dff_B_EYIGmiwN3_0(.din(n208),.dout(w_dff_B_EYIGmiwN3_0),.clk(gclk));
	jdff dff_B_JX4ZO1KH1_0(.din(w_dff_B_EYIGmiwN3_0),.dout(w_dff_B_JX4ZO1KH1_0),.clk(gclk));
	jdff dff_B_F4gDpcuX1_2(.din(n143),.dout(w_dff_B_F4gDpcuX1_2),.clk(gclk));
	jdff dff_B_6DhNYeSz7_2(.din(w_dff_B_F4gDpcuX1_2),.dout(w_dff_B_6DhNYeSz7_2),.clk(gclk));
	jdff dff_B_vMrHShPs0_2(.din(w_dff_B_6DhNYeSz7_2),.dout(w_dff_B_vMrHShPs0_2),.clk(gclk));
	jdff dff_B_cEECPJF44_2(.din(w_dff_B_vMrHShPs0_2),.dout(w_dff_B_cEECPJF44_2),.clk(gclk));
	jdff dff_B_1VoLqFOE1_2(.din(w_dff_B_cEECPJF44_2),.dout(w_dff_B_1VoLqFOE1_2),.clk(gclk));
	jdff dff_B_N5SRkjjz3_2(.din(w_dff_B_1VoLqFOE1_2),.dout(w_dff_B_N5SRkjjz3_2),.clk(gclk));
	jdff dff_B_eja3Zprr7_2(.din(w_dff_B_N5SRkjjz3_2),.dout(w_dff_B_eja3Zprr7_2),.clk(gclk));
	jdff dff_B_9vwFIlb01_2(.din(w_dff_B_eja3Zprr7_2),.dout(w_dff_B_9vwFIlb01_2),.clk(gclk));
	jdff dff_B_cvM5anir9_2(.din(w_dff_B_9vwFIlb01_2),.dout(w_dff_B_cvM5anir9_2),.clk(gclk));
	jdff dff_A_IqsW8ezY1_0(.dout(w_n196_0[0]),.din(w_dff_A_IqsW8ezY1_0),.clk(gclk));
	jdff dff_A_opLtEpGM9_1(.dout(w_n154_0[1]),.din(w_dff_A_opLtEpGM9_1),.clk(gclk));
	jdff dff_A_SFxqKb714_1(.dout(w_n303_0[1]),.din(w_dff_A_SFxqKb714_1),.clk(gclk));
	jdff dff_A_tG4Nq4tb6_1(.dout(w_dff_A_SFxqKb714_1),.din(w_dff_A_tG4Nq4tb6_1),.clk(gclk));
	jdff dff_A_onlv1ElE5_1(.dout(w_dff_A_tG4Nq4tb6_1),.din(w_dff_A_onlv1ElE5_1),.clk(gclk));
	jdff dff_A_4QIIxiCh7_1(.dout(w_dff_A_onlv1ElE5_1),.din(w_dff_A_4QIIxiCh7_1),.clk(gclk));
	jdff dff_A_pIASlKGO9_1(.dout(w_n302_0[1]),.din(w_dff_A_pIASlKGO9_1),.clk(gclk));
	jdff dff_A_EJErUeDG7_1(.dout(w_dff_A_pIASlKGO9_1),.din(w_dff_A_EJErUeDG7_1),.clk(gclk));
	jdff dff_A_tgJgbBm83_1(.dout(w_dff_A_EJErUeDG7_1),.din(w_dff_A_tgJgbBm83_1),.clk(gclk));
	jdff dff_A_FagwKQkI8_1(.dout(w_dff_A_tgJgbBm83_1),.din(w_dff_A_FagwKQkI8_1),.clk(gclk));
	jdff dff_A_DxIJJiKv9_1(.dout(w_dff_A_FagwKQkI8_1),.din(w_dff_A_DxIJJiKv9_1),.clk(gclk));
	jdff dff_B_7LyFN7op3_1(.din(n190),.dout(w_dff_B_7LyFN7op3_1),.clk(gclk));
	jdff dff_A_ZiT1WcL60_1(.dout(w_n165_1[1]),.din(w_dff_A_ZiT1WcL60_1),.clk(gclk));
	jdff dff_A_XmYDxrZe7_1(.dout(w_dff_A_ZiT1WcL60_1),.din(w_dff_A_XmYDxrZe7_1),.clk(gclk));
	jdff dff_A_pGAtQyKd6_2(.dout(w_n165_1[2]),.din(w_dff_A_pGAtQyKd6_2),.clk(gclk));
	jdff dff_A_AMWZ37Nv6_2(.dout(w_dff_A_pGAtQyKd6_2),.din(w_dff_A_AMWZ37Nv6_2),.clk(gclk));
	jdff dff_A_sdFNJJ7Q5_1(.dout(w_n165_0[1]),.din(w_dff_A_sdFNJJ7Q5_1),.clk(gclk));
	jdff dff_A_3Sp17NIj4_1(.dout(w_dff_A_sdFNJJ7Q5_1),.din(w_dff_A_3Sp17NIj4_1),.clk(gclk));
	jdff dff_A_kApIzi8Z9_2(.dout(w_n165_0[2]),.din(w_dff_A_kApIzi8Z9_2),.clk(gclk));
	jdff dff_A_7kPryKTi9_2(.dout(w_dff_A_kApIzi8Z9_2),.din(w_dff_A_7kPryKTi9_2),.clk(gclk));
	jdff dff_B_mUBMt6NB3_0(.din(n164),.dout(w_dff_B_mUBMt6NB3_0),.clk(gclk));
	jdff dff_A_C2Hev3HG1_1(.dout(w_G143gat_0[1]),.din(w_dff_A_C2Hev3HG1_1),.clk(gclk));
	jdff dff_B_ti8FtAkU0_2(.din(G143gat),.dout(w_dff_B_ti8FtAkU0_2),.clk(gclk));
	jdff dff_B_mJXsWUe91_2(.din(w_dff_B_ti8FtAkU0_2),.dout(w_dff_B_mJXsWUe91_2),.clk(gclk));
	jdff dff_B_ECMNNrAZ5_2(.din(w_dff_B_mJXsWUe91_2),.dout(w_dff_B_ECMNNrAZ5_2),.clk(gclk));
	jdff dff_B_5FCgSxWW5_2(.din(w_dff_B_ECMNNrAZ5_2),.dout(w_dff_B_5FCgSxWW5_2),.clk(gclk));
	jdff dff_A_610Oumgu4_0(.dout(w_n335_0[0]),.din(w_dff_A_610Oumgu4_0),.clk(gclk));
	jdff dff_A_Y3OHDiIv6_0(.dout(w_dff_A_610Oumgu4_0),.din(w_dff_A_Y3OHDiIv6_0),.clk(gclk));
	jdff dff_A_tohiyxjx3_0(.dout(w_dff_A_Y3OHDiIv6_0),.din(w_dff_A_tohiyxjx3_0),.clk(gclk));
	jdff dff_A_RwO6VadG0_0(.dout(w_dff_A_tohiyxjx3_0),.din(w_dff_A_RwO6VadG0_0),.clk(gclk));
	jdff dff_A_10I71eYm2_0(.dout(w_dff_A_RwO6VadG0_0),.din(w_dff_A_10I71eYm2_0),.clk(gclk));
	jdff dff_A_SkXC7s7y6_0(.dout(w_dff_A_10I71eYm2_0),.din(w_dff_A_SkXC7s7y6_0),.clk(gclk));
	jdff dff_A_LavkY5SI2_0(.dout(w_dff_A_SkXC7s7y6_0),.din(w_dff_A_LavkY5SI2_0),.clk(gclk));
	jdff dff_A_kpotA8MX8_0(.dout(w_dff_A_LavkY5SI2_0),.din(w_dff_A_kpotA8MX8_0),.clk(gclk));
	jdff dff_B_qRg2ss9o7_0(.din(n325),.dout(w_dff_B_qRg2ss9o7_0),.clk(gclk));
	jdff dff_B_l32VDpjh5_0(.din(w_dff_B_qRg2ss9o7_0),.dout(w_dff_B_l32VDpjh5_0),.clk(gclk));
	jdff dff_B_DLghQFNe1_0(.din(w_dff_B_l32VDpjh5_0),.dout(w_dff_B_DLghQFNe1_0),.clk(gclk));
	jdff dff_A_wVds7YOW6_1(.dout(w_n405_0[1]),.din(w_dff_A_wVds7YOW6_1),.clk(gclk));
	jdff dff_A_omLyDlCE5_1(.dout(w_dff_A_wVds7YOW6_1),.din(w_dff_A_omLyDlCE5_1),.clk(gclk));
	jdff dff_A_Yqer7f1Z9_1(.dout(w_dff_A_omLyDlCE5_1),.din(w_dff_A_Yqer7f1Z9_1),.clk(gclk));
	jdff dff_A_2Mmiek4i6_1(.dout(w_dff_A_Yqer7f1Z9_1),.din(w_dff_A_2Mmiek4i6_1),.clk(gclk));
	jdff dff_A_Yk8tPvBx2_1(.dout(w_dff_A_2Mmiek4i6_1),.din(w_dff_A_Yk8tPvBx2_1),.clk(gclk));
	jdff dff_A_pmkPh0bg4_1(.dout(w_dff_A_Yk8tPvBx2_1),.din(w_dff_A_pmkPh0bg4_1),.clk(gclk));
	jdff dff_A_6DpZ3zki6_1(.dout(w_dff_A_pmkPh0bg4_1),.din(w_dff_A_6DpZ3zki6_1),.clk(gclk));
	jdff dff_A_Ufn7cS606_1(.dout(w_dff_A_6DpZ3zki6_1),.din(w_dff_A_Ufn7cS606_1),.clk(gclk));
	jdff dff_A_TyLlz1ve1_1(.dout(w_dff_A_Ufn7cS606_1),.din(w_dff_A_TyLlz1ve1_1),.clk(gclk));
	jdff dff_B_eCkkmDWn5_0(.din(n318),.dout(w_dff_B_eCkkmDWn5_0),.clk(gclk));
	jdff dff_B_f3GLSOQR9_0(.din(w_dff_B_eCkkmDWn5_0),.dout(w_dff_B_f3GLSOQR9_0),.clk(gclk));
	jdff dff_B_lPbYyXpM1_0(.din(w_dff_B_f3GLSOQR9_0),.dout(w_dff_B_lPbYyXpM1_0),.clk(gclk));
	jdff dff_B_y0MrhwVI7_0(.din(n295),.dout(w_dff_B_y0MrhwVI7_0),.clk(gclk));
	jdff dff_A_xfZ43KYV4_1(.dout(w_G149gat_0[1]),.din(w_dff_A_xfZ43KYV4_1),.clk(gclk));
	jdff dff_B_JrSDgxZO4_2(.din(G149gat),.dout(w_dff_B_JrSDgxZO4_2),.clk(gclk));
	jdff dff_B_tqwvZllI5_2(.din(w_dff_B_JrSDgxZO4_2),.dout(w_dff_B_tqwvZllI5_2),.clk(gclk));
	jdff dff_B_h1lEKOyn7_2(.din(w_dff_B_tqwvZllI5_2),.dout(w_dff_B_h1lEKOyn7_2),.clk(gclk));
	jdff dff_B_HZ81dAzI8_2(.din(w_dff_B_h1lEKOyn7_2),.dout(w_dff_B_HZ81dAzI8_2),.clk(gclk));
	jdff dff_B_zoCoK8vb1_0(.din(n152),.dout(w_dff_B_zoCoK8vb1_0),.clk(gclk));
	jdff dff_A_12pK7KFc3_2(.dout(w_dff_A_Nveud2mb4_0),.din(w_dff_A_12pK7KFc3_2),.clk(gclk));
	jdff dff_A_Nveud2mb4_0(.dout(w_dff_A_xoZZ7Jkz7_0),.din(w_dff_A_Nveud2mb4_0),.clk(gclk));
	jdff dff_A_xoZZ7Jkz7_0(.dout(w_dff_A_Zg9LcbsT3_0),.din(w_dff_A_xoZZ7Jkz7_0),.clk(gclk));
	jdff dff_A_Zg9LcbsT3_0(.dout(w_dff_A_QlZpgouh9_0),.din(w_dff_A_Zg9LcbsT3_0),.clk(gclk));
	jdff dff_A_QlZpgouh9_0(.dout(w_dff_A_HNUFoqL81_0),.din(w_dff_A_QlZpgouh9_0),.clk(gclk));
	jdff dff_A_HNUFoqL81_0(.dout(w_dff_A_rrYcQ1I47_0),.din(w_dff_A_HNUFoqL81_0),.clk(gclk));
	jdff dff_A_rrYcQ1I47_0(.dout(w_dff_A_gKljUF238_0),.din(w_dff_A_rrYcQ1I47_0),.clk(gclk));
	jdff dff_A_gKljUF238_0(.dout(w_dff_A_IwEWevRP9_0),.din(w_dff_A_gKljUF238_0),.clk(gclk));
	jdff dff_A_IwEWevRP9_0(.dout(w_dff_A_kVEtRdgL9_0),.din(w_dff_A_IwEWevRP9_0),.clk(gclk));
	jdff dff_A_kVEtRdgL9_0(.dout(w_dff_A_nwyhWHvG0_0),.din(w_dff_A_kVEtRdgL9_0),.clk(gclk));
	jdff dff_A_nwyhWHvG0_0(.dout(w_dff_A_7M2Y2uWs8_0),.din(w_dff_A_nwyhWHvG0_0),.clk(gclk));
	jdff dff_A_7M2Y2uWs8_0(.dout(w_dff_A_iGPJBw3f6_0),.din(w_dff_A_7M2Y2uWs8_0),.clk(gclk));
	jdff dff_A_iGPJBw3f6_0(.dout(w_dff_A_sgUhCVAf1_0),.din(w_dff_A_iGPJBw3f6_0),.clk(gclk));
	jdff dff_A_sgUhCVAf1_0(.dout(w_dff_A_3s5spF6g2_0),.din(w_dff_A_sgUhCVAf1_0),.clk(gclk));
	jdff dff_A_3s5spF6g2_0(.dout(w_dff_A_vQYkxVWn0_0),.din(w_dff_A_3s5spF6g2_0),.clk(gclk));
	jdff dff_A_vQYkxVWn0_0(.dout(w_dff_A_Mz7EY8u92_0),.din(w_dff_A_vQYkxVWn0_0),.clk(gclk));
	jdff dff_A_Mz7EY8u92_0(.dout(w_dff_A_XRaOVevl0_0),.din(w_dff_A_Mz7EY8u92_0),.clk(gclk));
	jdff dff_A_XRaOVevl0_0(.dout(w_dff_A_YKEeeP0I3_0),.din(w_dff_A_XRaOVevl0_0),.clk(gclk));
	jdff dff_A_YKEeeP0I3_0(.dout(G388gat),.din(w_dff_A_YKEeeP0I3_0),.clk(gclk));
	jdff dff_A_FYUoAM6L3_2(.dout(w_dff_A_ogZ22fll2_0),.din(w_dff_A_FYUoAM6L3_2),.clk(gclk));
	jdff dff_A_ogZ22fll2_0(.dout(w_dff_A_7UWG0EaP4_0),.din(w_dff_A_ogZ22fll2_0),.clk(gclk));
	jdff dff_A_7UWG0EaP4_0(.dout(w_dff_A_meZ70Nsa8_0),.din(w_dff_A_7UWG0EaP4_0),.clk(gclk));
	jdff dff_A_meZ70Nsa8_0(.dout(w_dff_A_vKDZbclY4_0),.din(w_dff_A_meZ70Nsa8_0),.clk(gclk));
	jdff dff_A_vKDZbclY4_0(.dout(w_dff_A_5K1rvWm95_0),.din(w_dff_A_vKDZbclY4_0),.clk(gclk));
	jdff dff_A_5K1rvWm95_0(.dout(w_dff_A_3I0AGCyS6_0),.din(w_dff_A_5K1rvWm95_0),.clk(gclk));
	jdff dff_A_3I0AGCyS6_0(.dout(w_dff_A_lAuTnL480_0),.din(w_dff_A_3I0AGCyS6_0),.clk(gclk));
	jdff dff_A_lAuTnL480_0(.dout(w_dff_A_8POfUgPe4_0),.din(w_dff_A_lAuTnL480_0),.clk(gclk));
	jdff dff_A_8POfUgPe4_0(.dout(w_dff_A_xxSUZAv19_0),.din(w_dff_A_8POfUgPe4_0),.clk(gclk));
	jdff dff_A_xxSUZAv19_0(.dout(w_dff_A_ZOicGVPq3_0),.din(w_dff_A_xxSUZAv19_0),.clk(gclk));
	jdff dff_A_ZOicGVPq3_0(.dout(w_dff_A_UqHiV6yw3_0),.din(w_dff_A_ZOicGVPq3_0),.clk(gclk));
	jdff dff_A_UqHiV6yw3_0(.dout(w_dff_A_yBosPtPM2_0),.din(w_dff_A_UqHiV6yw3_0),.clk(gclk));
	jdff dff_A_yBosPtPM2_0(.dout(w_dff_A_4caEvDFc9_0),.din(w_dff_A_yBosPtPM2_0),.clk(gclk));
	jdff dff_A_4caEvDFc9_0(.dout(w_dff_A_3lIBw1P08_0),.din(w_dff_A_4caEvDFc9_0),.clk(gclk));
	jdff dff_A_3lIBw1P08_0(.dout(w_dff_A_EiHRece77_0),.din(w_dff_A_3lIBw1P08_0),.clk(gclk));
	jdff dff_A_EiHRece77_0(.dout(w_dff_A_DOr5tNY45_0),.din(w_dff_A_EiHRece77_0),.clk(gclk));
	jdff dff_A_DOr5tNY45_0(.dout(w_dff_A_3s61wg1Z0_0),.din(w_dff_A_DOr5tNY45_0),.clk(gclk));
	jdff dff_A_3s61wg1Z0_0(.dout(w_dff_A_H1Mx3OzL2_0),.din(w_dff_A_3s61wg1Z0_0),.clk(gclk));
	jdff dff_A_H1Mx3OzL2_0(.dout(G389gat),.din(w_dff_A_H1Mx3OzL2_0),.clk(gclk));
	jdff dff_A_EHSzjLlc3_2(.dout(w_dff_A_CHgW6rD36_0),.din(w_dff_A_EHSzjLlc3_2),.clk(gclk));
	jdff dff_A_CHgW6rD36_0(.dout(w_dff_A_WKZJB1pK8_0),.din(w_dff_A_CHgW6rD36_0),.clk(gclk));
	jdff dff_A_WKZJB1pK8_0(.dout(w_dff_A_zwvz0RKX7_0),.din(w_dff_A_WKZJB1pK8_0),.clk(gclk));
	jdff dff_A_zwvz0RKX7_0(.dout(w_dff_A_6emzrazG6_0),.din(w_dff_A_zwvz0RKX7_0),.clk(gclk));
	jdff dff_A_6emzrazG6_0(.dout(w_dff_A_yMYXFCny4_0),.din(w_dff_A_6emzrazG6_0),.clk(gclk));
	jdff dff_A_yMYXFCny4_0(.dout(w_dff_A_luCt5MGJ7_0),.din(w_dff_A_yMYXFCny4_0),.clk(gclk));
	jdff dff_A_luCt5MGJ7_0(.dout(w_dff_A_iWBGAb963_0),.din(w_dff_A_luCt5MGJ7_0),.clk(gclk));
	jdff dff_A_iWBGAb963_0(.dout(w_dff_A_7K20HTUv0_0),.din(w_dff_A_iWBGAb963_0),.clk(gclk));
	jdff dff_A_7K20HTUv0_0(.dout(w_dff_A_DR3qcy2o0_0),.din(w_dff_A_7K20HTUv0_0),.clk(gclk));
	jdff dff_A_DR3qcy2o0_0(.dout(w_dff_A_3wc6nGDp3_0),.din(w_dff_A_DR3qcy2o0_0),.clk(gclk));
	jdff dff_A_3wc6nGDp3_0(.dout(w_dff_A_d0oS4S9Y3_0),.din(w_dff_A_3wc6nGDp3_0),.clk(gclk));
	jdff dff_A_d0oS4S9Y3_0(.dout(w_dff_A_fsMYUN2z0_0),.din(w_dff_A_d0oS4S9Y3_0),.clk(gclk));
	jdff dff_A_fsMYUN2z0_0(.dout(w_dff_A_RxFQS75U2_0),.din(w_dff_A_fsMYUN2z0_0),.clk(gclk));
	jdff dff_A_RxFQS75U2_0(.dout(w_dff_A_Urzsjl4R9_0),.din(w_dff_A_RxFQS75U2_0),.clk(gclk));
	jdff dff_A_Urzsjl4R9_0(.dout(w_dff_A_yKYK3RC75_0),.din(w_dff_A_Urzsjl4R9_0),.clk(gclk));
	jdff dff_A_yKYK3RC75_0(.dout(w_dff_A_eT5arAwv6_0),.din(w_dff_A_yKYK3RC75_0),.clk(gclk));
	jdff dff_A_eT5arAwv6_0(.dout(w_dff_A_eGguc1PC8_0),.din(w_dff_A_eT5arAwv6_0),.clk(gclk));
	jdff dff_A_eGguc1PC8_0(.dout(w_dff_A_QsWLzBPp5_0),.din(w_dff_A_eGguc1PC8_0),.clk(gclk));
	jdff dff_A_QsWLzBPp5_0(.dout(G390gat),.din(w_dff_A_QsWLzBPp5_0),.clk(gclk));
	jdff dff_A_ZCq0xqL09_2(.dout(w_dff_A_OX7zotRu9_0),.din(w_dff_A_ZCq0xqL09_2),.clk(gclk));
	jdff dff_A_OX7zotRu9_0(.dout(w_dff_A_7B1SBpp09_0),.din(w_dff_A_OX7zotRu9_0),.clk(gclk));
	jdff dff_A_7B1SBpp09_0(.dout(w_dff_A_8eKlMoEv8_0),.din(w_dff_A_7B1SBpp09_0),.clk(gclk));
	jdff dff_A_8eKlMoEv8_0(.dout(w_dff_A_tucDdLNP2_0),.din(w_dff_A_8eKlMoEv8_0),.clk(gclk));
	jdff dff_A_tucDdLNP2_0(.dout(w_dff_A_MAIFzxIl4_0),.din(w_dff_A_tucDdLNP2_0),.clk(gclk));
	jdff dff_A_MAIFzxIl4_0(.dout(w_dff_A_zkYMUutu2_0),.din(w_dff_A_MAIFzxIl4_0),.clk(gclk));
	jdff dff_A_zkYMUutu2_0(.dout(w_dff_A_BmAIfwi21_0),.din(w_dff_A_zkYMUutu2_0),.clk(gclk));
	jdff dff_A_BmAIfwi21_0(.dout(w_dff_A_JxEO3Ebr1_0),.din(w_dff_A_BmAIfwi21_0),.clk(gclk));
	jdff dff_A_JxEO3Ebr1_0(.dout(w_dff_A_twuc0zMm3_0),.din(w_dff_A_JxEO3Ebr1_0),.clk(gclk));
	jdff dff_A_twuc0zMm3_0(.dout(w_dff_A_bAFBj0FT7_0),.din(w_dff_A_twuc0zMm3_0),.clk(gclk));
	jdff dff_A_bAFBj0FT7_0(.dout(w_dff_A_QUul71P98_0),.din(w_dff_A_bAFBj0FT7_0),.clk(gclk));
	jdff dff_A_QUul71P98_0(.dout(w_dff_A_PmtXLCV48_0),.din(w_dff_A_QUul71P98_0),.clk(gclk));
	jdff dff_A_PmtXLCV48_0(.dout(w_dff_A_ZSPijMuI7_0),.din(w_dff_A_PmtXLCV48_0),.clk(gclk));
	jdff dff_A_ZSPijMuI7_0(.dout(w_dff_A_vmuLVgYq7_0),.din(w_dff_A_ZSPijMuI7_0),.clk(gclk));
	jdff dff_A_vmuLVgYq7_0(.dout(w_dff_A_Jb0My8Pv7_0),.din(w_dff_A_vmuLVgYq7_0),.clk(gclk));
	jdff dff_A_Jb0My8Pv7_0(.dout(w_dff_A_9RpbWCG31_0),.din(w_dff_A_Jb0My8Pv7_0),.clk(gclk));
	jdff dff_A_9RpbWCG31_0(.dout(w_dff_A_mrxqTp7K4_0),.din(w_dff_A_9RpbWCG31_0),.clk(gclk));
	jdff dff_A_mrxqTp7K4_0(.dout(w_dff_A_8ESfrLvh2_0),.din(w_dff_A_mrxqTp7K4_0),.clk(gclk));
	jdff dff_A_8ESfrLvh2_0(.dout(w_dff_A_QxF9Ckid9_0),.din(w_dff_A_8ESfrLvh2_0),.clk(gclk));
	jdff dff_A_QxF9Ckid9_0(.dout(G391gat),.din(w_dff_A_QxF9Ckid9_0),.clk(gclk));
	jdff dff_A_sp5SF7qA2_2(.dout(w_dff_A_Up6sy3FS0_0),.din(w_dff_A_sp5SF7qA2_2),.clk(gclk));
	jdff dff_A_Up6sy3FS0_0(.dout(w_dff_A_uaI8ct1b1_0),.din(w_dff_A_Up6sy3FS0_0),.clk(gclk));
	jdff dff_A_uaI8ct1b1_0(.dout(w_dff_A_oD9tbUIl9_0),.din(w_dff_A_uaI8ct1b1_0),.clk(gclk));
	jdff dff_A_oD9tbUIl9_0(.dout(w_dff_A_pITwVpZq7_0),.din(w_dff_A_oD9tbUIl9_0),.clk(gclk));
	jdff dff_A_pITwVpZq7_0(.dout(w_dff_A_9jR9Icnk1_0),.din(w_dff_A_pITwVpZq7_0),.clk(gclk));
	jdff dff_A_9jR9Icnk1_0(.dout(w_dff_A_2ShS7tyM6_0),.din(w_dff_A_9jR9Icnk1_0),.clk(gclk));
	jdff dff_A_2ShS7tyM6_0(.dout(w_dff_A_hJcR9PoC8_0),.din(w_dff_A_2ShS7tyM6_0),.clk(gclk));
	jdff dff_A_hJcR9PoC8_0(.dout(w_dff_A_r5vxBedS4_0),.din(w_dff_A_hJcR9PoC8_0),.clk(gclk));
	jdff dff_A_r5vxBedS4_0(.dout(w_dff_A_dxIJo9643_0),.din(w_dff_A_r5vxBedS4_0),.clk(gclk));
	jdff dff_A_dxIJo9643_0(.dout(w_dff_A_SfiwhXMv5_0),.din(w_dff_A_dxIJo9643_0),.clk(gclk));
	jdff dff_A_SfiwhXMv5_0(.dout(w_dff_A_ulpUGvSQ9_0),.din(w_dff_A_SfiwhXMv5_0),.clk(gclk));
	jdff dff_A_ulpUGvSQ9_0(.dout(w_dff_A_dhBdF6Sx1_0),.din(w_dff_A_ulpUGvSQ9_0),.clk(gclk));
	jdff dff_A_dhBdF6Sx1_0(.dout(w_dff_A_xTSljTPF5_0),.din(w_dff_A_dhBdF6Sx1_0),.clk(gclk));
	jdff dff_A_xTSljTPF5_0(.dout(w_dff_A_ngUQHmGZ0_0),.din(w_dff_A_xTSljTPF5_0),.clk(gclk));
	jdff dff_A_ngUQHmGZ0_0(.dout(w_dff_A_3ZSrSQEb4_0),.din(w_dff_A_ngUQHmGZ0_0),.clk(gclk));
	jdff dff_A_3ZSrSQEb4_0(.dout(w_dff_A_F5dugAzX6_0),.din(w_dff_A_3ZSrSQEb4_0),.clk(gclk));
	jdff dff_A_F5dugAzX6_0(.dout(w_dff_A_tclHPkqb7_0),.din(w_dff_A_F5dugAzX6_0),.clk(gclk));
	jdff dff_A_tclHPkqb7_0(.dout(w_dff_A_3joSsVwd5_0),.din(w_dff_A_tclHPkqb7_0),.clk(gclk));
	jdff dff_A_3joSsVwd5_0(.dout(G418gat),.din(w_dff_A_3joSsVwd5_0),.clk(gclk));
	jdff dff_A_JtEJsWvz5_2(.dout(w_dff_A_RgWFr1om1_0),.din(w_dff_A_JtEJsWvz5_2),.clk(gclk));
	jdff dff_A_RgWFr1om1_0(.dout(w_dff_A_z35lUeDj8_0),.din(w_dff_A_RgWFr1om1_0),.clk(gclk));
	jdff dff_A_z35lUeDj8_0(.dout(w_dff_A_kxs59J0J1_0),.din(w_dff_A_z35lUeDj8_0),.clk(gclk));
	jdff dff_A_kxs59J0J1_0(.dout(w_dff_A_T6Z5mPxI4_0),.din(w_dff_A_kxs59J0J1_0),.clk(gclk));
	jdff dff_A_T6Z5mPxI4_0(.dout(w_dff_A_BPwf4RUr5_0),.din(w_dff_A_T6Z5mPxI4_0),.clk(gclk));
	jdff dff_A_BPwf4RUr5_0(.dout(w_dff_A_Yowidf4B2_0),.din(w_dff_A_BPwf4RUr5_0),.clk(gclk));
	jdff dff_A_Yowidf4B2_0(.dout(w_dff_A_y4Lb7yxw8_0),.din(w_dff_A_Yowidf4B2_0),.clk(gclk));
	jdff dff_A_y4Lb7yxw8_0(.dout(w_dff_A_En05gtRn1_0),.din(w_dff_A_y4Lb7yxw8_0),.clk(gclk));
	jdff dff_A_En05gtRn1_0(.dout(w_dff_A_Xg0EORiO8_0),.din(w_dff_A_En05gtRn1_0),.clk(gclk));
	jdff dff_A_Xg0EORiO8_0(.dout(w_dff_A_do6nehmm3_0),.din(w_dff_A_Xg0EORiO8_0),.clk(gclk));
	jdff dff_A_do6nehmm3_0(.dout(w_dff_A_zcAkv89N2_0),.din(w_dff_A_do6nehmm3_0),.clk(gclk));
	jdff dff_A_zcAkv89N2_0(.dout(w_dff_A_GxEeDsfF3_0),.din(w_dff_A_zcAkv89N2_0),.clk(gclk));
	jdff dff_A_GxEeDsfF3_0(.dout(w_dff_A_rYnVwgbd8_0),.din(w_dff_A_GxEeDsfF3_0),.clk(gclk));
	jdff dff_A_rYnVwgbd8_0(.dout(w_dff_A_zpGG2Epo0_0),.din(w_dff_A_rYnVwgbd8_0),.clk(gclk));
	jdff dff_A_zpGG2Epo0_0(.dout(w_dff_A_T9rnltFe9_0),.din(w_dff_A_zpGG2Epo0_0),.clk(gclk));
	jdff dff_A_T9rnltFe9_0(.dout(w_dff_A_ufgHCMDh0_0),.din(w_dff_A_T9rnltFe9_0),.clk(gclk));
	jdff dff_A_ufgHCMDh0_0(.dout(G419gat),.din(w_dff_A_ufgHCMDh0_0),.clk(gclk));
	jdff dff_A_VXgXdQO33_2(.dout(w_dff_A_QoAfB4xV7_0),.din(w_dff_A_VXgXdQO33_2),.clk(gclk));
	jdff dff_A_QoAfB4xV7_0(.dout(w_dff_A_qdlT4Qmi0_0),.din(w_dff_A_QoAfB4xV7_0),.clk(gclk));
	jdff dff_A_qdlT4Qmi0_0(.dout(w_dff_A_wKFO3nBv6_0),.din(w_dff_A_qdlT4Qmi0_0),.clk(gclk));
	jdff dff_A_wKFO3nBv6_0(.dout(w_dff_A_nVaZOBoR7_0),.din(w_dff_A_wKFO3nBv6_0),.clk(gclk));
	jdff dff_A_nVaZOBoR7_0(.dout(w_dff_A_klkChoYf7_0),.din(w_dff_A_nVaZOBoR7_0),.clk(gclk));
	jdff dff_A_klkChoYf7_0(.dout(w_dff_A_HOS84ROD3_0),.din(w_dff_A_klkChoYf7_0),.clk(gclk));
	jdff dff_A_HOS84ROD3_0(.dout(w_dff_A_euiWmpy41_0),.din(w_dff_A_HOS84ROD3_0),.clk(gclk));
	jdff dff_A_euiWmpy41_0(.dout(w_dff_A_sv8AxLK32_0),.din(w_dff_A_euiWmpy41_0),.clk(gclk));
	jdff dff_A_sv8AxLK32_0(.dout(w_dff_A_VN5JsFDp9_0),.din(w_dff_A_sv8AxLK32_0),.clk(gclk));
	jdff dff_A_VN5JsFDp9_0(.dout(w_dff_A_rIALY9Lu8_0),.din(w_dff_A_VN5JsFDp9_0),.clk(gclk));
	jdff dff_A_rIALY9Lu8_0(.dout(w_dff_A_MCdaAqhP8_0),.din(w_dff_A_rIALY9Lu8_0),.clk(gclk));
	jdff dff_A_MCdaAqhP8_0(.dout(w_dff_A_e7TUax423_0),.din(w_dff_A_MCdaAqhP8_0),.clk(gclk));
	jdff dff_A_e7TUax423_0(.dout(w_dff_A_K9RL7O5H6_0),.din(w_dff_A_e7TUax423_0),.clk(gclk));
	jdff dff_A_K9RL7O5H6_0(.dout(w_dff_A_1g012K3M1_0),.din(w_dff_A_K9RL7O5H6_0),.clk(gclk));
	jdff dff_A_1g012K3M1_0(.dout(w_dff_A_jVwmXysm7_0),.din(w_dff_A_1g012K3M1_0),.clk(gclk));
	jdff dff_A_jVwmXysm7_0(.dout(w_dff_A_b4LprVON7_0),.din(w_dff_A_jVwmXysm7_0),.clk(gclk));
	jdff dff_A_b4LprVON7_0(.dout(w_dff_A_Vy0iPKTt6_0),.din(w_dff_A_b4LprVON7_0),.clk(gclk));
	jdff dff_A_Vy0iPKTt6_0(.dout(G420gat),.din(w_dff_A_Vy0iPKTt6_0),.clk(gclk));
	jdff dff_A_mvmvstLj6_2(.dout(w_dff_A_roSsMDkw8_0),.din(w_dff_A_mvmvstLj6_2),.clk(gclk));
	jdff dff_A_roSsMDkw8_0(.dout(w_dff_A_rJnnjq135_0),.din(w_dff_A_roSsMDkw8_0),.clk(gclk));
	jdff dff_A_rJnnjq135_0(.dout(w_dff_A_aBdCM3vx1_0),.din(w_dff_A_rJnnjq135_0),.clk(gclk));
	jdff dff_A_aBdCM3vx1_0(.dout(w_dff_A_lTMycKqF8_0),.din(w_dff_A_aBdCM3vx1_0),.clk(gclk));
	jdff dff_A_lTMycKqF8_0(.dout(w_dff_A_mWSbzQui7_0),.din(w_dff_A_lTMycKqF8_0),.clk(gclk));
	jdff dff_A_mWSbzQui7_0(.dout(w_dff_A_0kwWmSbM3_0),.din(w_dff_A_mWSbzQui7_0),.clk(gclk));
	jdff dff_A_0kwWmSbM3_0(.dout(w_dff_A_HkcuJTrZ8_0),.din(w_dff_A_0kwWmSbM3_0),.clk(gclk));
	jdff dff_A_HkcuJTrZ8_0(.dout(w_dff_A_xFaU33vH3_0),.din(w_dff_A_HkcuJTrZ8_0),.clk(gclk));
	jdff dff_A_xFaU33vH3_0(.dout(w_dff_A_tJ3L6kF58_0),.din(w_dff_A_xFaU33vH3_0),.clk(gclk));
	jdff dff_A_tJ3L6kF58_0(.dout(w_dff_A_8DZTt0635_0),.din(w_dff_A_tJ3L6kF58_0),.clk(gclk));
	jdff dff_A_8DZTt0635_0(.dout(w_dff_A_PqyY8gLg0_0),.din(w_dff_A_8DZTt0635_0),.clk(gclk));
	jdff dff_A_PqyY8gLg0_0(.dout(w_dff_A_YVRePyug4_0),.din(w_dff_A_PqyY8gLg0_0),.clk(gclk));
	jdff dff_A_YVRePyug4_0(.dout(w_dff_A_K4iCGIuu2_0),.din(w_dff_A_YVRePyug4_0),.clk(gclk));
	jdff dff_A_K4iCGIuu2_0(.dout(w_dff_A_VLntJJmv0_0),.din(w_dff_A_K4iCGIuu2_0),.clk(gclk));
	jdff dff_A_VLntJJmv0_0(.dout(w_dff_A_poeiRc8d5_0),.din(w_dff_A_VLntJJmv0_0),.clk(gclk));
	jdff dff_A_poeiRc8d5_0(.dout(w_dff_A_ShEdM7Zq4_0),.din(w_dff_A_poeiRc8d5_0),.clk(gclk));
	jdff dff_A_ShEdM7Zq4_0(.dout(w_dff_A_zRXboWsx4_0),.din(w_dff_A_ShEdM7Zq4_0),.clk(gclk));
	jdff dff_A_zRXboWsx4_0(.dout(G421gat),.din(w_dff_A_zRXboWsx4_0),.clk(gclk));
	jdff dff_A_V0h2bNiz8_2(.dout(w_dff_A_VhYTCX0u0_0),.din(w_dff_A_V0h2bNiz8_2),.clk(gclk));
	jdff dff_A_VhYTCX0u0_0(.dout(w_dff_A_OQEG2g6w3_0),.din(w_dff_A_VhYTCX0u0_0),.clk(gclk));
	jdff dff_A_OQEG2g6w3_0(.dout(w_dff_A_EiyWRMx56_0),.din(w_dff_A_OQEG2g6w3_0),.clk(gclk));
	jdff dff_A_EiyWRMx56_0(.dout(w_dff_A_75ThU4Se8_0),.din(w_dff_A_EiyWRMx56_0),.clk(gclk));
	jdff dff_A_75ThU4Se8_0(.dout(w_dff_A_ndBHxp119_0),.din(w_dff_A_75ThU4Se8_0),.clk(gclk));
	jdff dff_A_ndBHxp119_0(.dout(w_dff_A_Nq2CmN0x1_0),.din(w_dff_A_ndBHxp119_0),.clk(gclk));
	jdff dff_A_Nq2CmN0x1_0(.dout(w_dff_A_osrRrLa16_0),.din(w_dff_A_Nq2CmN0x1_0),.clk(gclk));
	jdff dff_A_osrRrLa16_0(.dout(w_dff_A_XrIWils97_0),.din(w_dff_A_osrRrLa16_0),.clk(gclk));
	jdff dff_A_XrIWils97_0(.dout(w_dff_A_oVglMcof2_0),.din(w_dff_A_XrIWils97_0),.clk(gclk));
	jdff dff_A_oVglMcof2_0(.dout(w_dff_A_NZwfK0w07_0),.din(w_dff_A_oVglMcof2_0),.clk(gclk));
	jdff dff_A_NZwfK0w07_0(.dout(w_dff_A_Cz4iHh9w7_0),.din(w_dff_A_NZwfK0w07_0),.clk(gclk));
	jdff dff_A_Cz4iHh9w7_0(.dout(w_dff_A_zlFk3Zpt3_0),.din(w_dff_A_Cz4iHh9w7_0),.clk(gclk));
	jdff dff_A_zlFk3Zpt3_0(.dout(w_dff_A_9Nhf94Pr2_0),.din(w_dff_A_zlFk3Zpt3_0),.clk(gclk));
	jdff dff_A_9Nhf94Pr2_0(.dout(w_dff_A_asPOGsDj3_0),.din(w_dff_A_9Nhf94Pr2_0),.clk(gclk));
	jdff dff_A_asPOGsDj3_0(.dout(w_dff_A_YtitRDRr3_0),.din(w_dff_A_asPOGsDj3_0),.clk(gclk));
	jdff dff_A_YtitRDRr3_0(.dout(w_dff_A_zMJfpbpH5_0),.din(w_dff_A_YtitRDRr3_0),.clk(gclk));
	jdff dff_A_zMJfpbpH5_0(.dout(w_dff_A_U2gmkXaP9_0),.din(w_dff_A_zMJfpbpH5_0),.clk(gclk));
	jdff dff_A_U2gmkXaP9_0(.dout(G422gat),.din(w_dff_A_U2gmkXaP9_0),.clk(gclk));
	jdff dff_A_ivAHcPXp4_2(.dout(w_dff_A_V8FK9o7q5_0),.din(w_dff_A_ivAHcPXp4_2),.clk(gclk));
	jdff dff_A_V8FK9o7q5_0(.dout(w_dff_A_wCwWlHje0_0),.din(w_dff_A_V8FK9o7q5_0),.clk(gclk));
	jdff dff_A_wCwWlHje0_0(.dout(w_dff_A_AG4ASDGc5_0),.din(w_dff_A_wCwWlHje0_0),.clk(gclk));
	jdff dff_A_AG4ASDGc5_0(.dout(w_dff_A_npQicJ6G0_0),.din(w_dff_A_AG4ASDGc5_0),.clk(gclk));
	jdff dff_A_npQicJ6G0_0(.dout(w_dff_A_BOxdcJ2r3_0),.din(w_dff_A_npQicJ6G0_0),.clk(gclk));
	jdff dff_A_BOxdcJ2r3_0(.dout(w_dff_A_q2oTiYMh5_0),.din(w_dff_A_BOxdcJ2r3_0),.clk(gclk));
	jdff dff_A_q2oTiYMh5_0(.dout(w_dff_A_0MO7Ygaz5_0),.din(w_dff_A_q2oTiYMh5_0),.clk(gclk));
	jdff dff_A_0MO7Ygaz5_0(.dout(w_dff_A_ptWoyQDO7_0),.din(w_dff_A_0MO7Ygaz5_0),.clk(gclk));
	jdff dff_A_ptWoyQDO7_0(.dout(w_dff_A_Z7SdAHdf9_0),.din(w_dff_A_ptWoyQDO7_0),.clk(gclk));
	jdff dff_A_Z7SdAHdf9_0(.dout(w_dff_A_LTpyagcE5_0),.din(w_dff_A_Z7SdAHdf9_0),.clk(gclk));
	jdff dff_A_LTpyagcE5_0(.dout(w_dff_A_TdrrNlVC7_0),.din(w_dff_A_LTpyagcE5_0),.clk(gclk));
	jdff dff_A_TdrrNlVC7_0(.dout(w_dff_A_RQN5qq0y7_0),.din(w_dff_A_TdrrNlVC7_0),.clk(gclk));
	jdff dff_A_RQN5qq0y7_0(.dout(w_dff_A_cN4MUD593_0),.din(w_dff_A_RQN5qq0y7_0),.clk(gclk));
	jdff dff_A_cN4MUD593_0(.dout(w_dff_A_2BDZbHvk2_0),.din(w_dff_A_cN4MUD593_0),.clk(gclk));
	jdff dff_A_2BDZbHvk2_0(.dout(w_dff_A_BqanhjYR4_0),.din(w_dff_A_2BDZbHvk2_0),.clk(gclk));
	jdff dff_A_BqanhjYR4_0(.dout(w_dff_A_XDfK61qz5_0),.din(w_dff_A_BqanhjYR4_0),.clk(gclk));
	jdff dff_A_XDfK61qz5_0(.dout(w_dff_A_vw1sRUCY3_0),.din(w_dff_A_XDfK61qz5_0),.clk(gclk));
	jdff dff_A_vw1sRUCY3_0(.dout(w_dff_A_LqvkWp1d7_0),.din(w_dff_A_vw1sRUCY3_0),.clk(gclk));
	jdff dff_A_LqvkWp1d7_0(.dout(G423gat),.din(w_dff_A_LqvkWp1d7_0),.clk(gclk));
	jdff dff_A_4az9XDkv0_2(.dout(w_dff_A_DNbR0gOT8_0),.din(w_dff_A_4az9XDkv0_2),.clk(gclk));
	jdff dff_A_DNbR0gOT8_0(.dout(w_dff_A_jI86XLkh7_0),.din(w_dff_A_DNbR0gOT8_0),.clk(gclk));
	jdff dff_A_jI86XLkh7_0(.dout(w_dff_A_96ag7xpi2_0),.din(w_dff_A_jI86XLkh7_0),.clk(gclk));
	jdff dff_A_96ag7xpi2_0(.dout(w_dff_A_VA3YOs9B7_0),.din(w_dff_A_96ag7xpi2_0),.clk(gclk));
	jdff dff_A_VA3YOs9B7_0(.dout(w_dff_A_EWdfiAOS7_0),.din(w_dff_A_VA3YOs9B7_0),.clk(gclk));
	jdff dff_A_EWdfiAOS7_0(.dout(w_dff_A_owjYhts39_0),.din(w_dff_A_EWdfiAOS7_0),.clk(gclk));
	jdff dff_A_owjYhts39_0(.dout(w_dff_A_509KKv2Y4_0),.din(w_dff_A_owjYhts39_0),.clk(gclk));
	jdff dff_A_509KKv2Y4_0(.dout(w_dff_A_cyIMQczN9_0),.din(w_dff_A_509KKv2Y4_0),.clk(gclk));
	jdff dff_A_cyIMQczN9_0(.dout(w_dff_A_e62MMZiP0_0),.din(w_dff_A_cyIMQczN9_0),.clk(gclk));
	jdff dff_A_e62MMZiP0_0(.dout(w_dff_A_NUQstSp63_0),.din(w_dff_A_e62MMZiP0_0),.clk(gclk));
	jdff dff_A_NUQstSp63_0(.dout(w_dff_A_bd3IgbbK2_0),.din(w_dff_A_NUQstSp63_0),.clk(gclk));
	jdff dff_A_bd3IgbbK2_0(.dout(w_dff_A_Ik5DVA7z7_0),.din(w_dff_A_bd3IgbbK2_0),.clk(gclk));
	jdff dff_A_Ik5DVA7z7_0(.dout(w_dff_A_6IvIwkv89_0),.din(w_dff_A_Ik5DVA7z7_0),.clk(gclk));
	jdff dff_A_6IvIwkv89_0(.dout(w_dff_A_4vQ4Uihz0_0),.din(w_dff_A_6IvIwkv89_0),.clk(gclk));
	jdff dff_A_4vQ4Uihz0_0(.dout(w_dff_A_of1NuLC28_0),.din(w_dff_A_4vQ4Uihz0_0),.clk(gclk));
	jdff dff_A_of1NuLC28_0(.dout(w_dff_A_FwjUHzgo8_0),.din(w_dff_A_of1NuLC28_0),.clk(gclk));
	jdff dff_A_FwjUHzgo8_0(.dout(G446gat),.din(w_dff_A_FwjUHzgo8_0),.clk(gclk));
	jdff dff_A_WuI0a5an7_1(.dout(w_dff_A_weJI9HQ41_0),.din(w_dff_A_WuI0a5an7_1),.clk(gclk));
	jdff dff_A_weJI9HQ41_0(.dout(w_dff_A_AKunf6VD6_0),.din(w_dff_A_weJI9HQ41_0),.clk(gclk));
	jdff dff_A_AKunf6VD6_0(.dout(w_dff_A_diOA7yQC8_0),.din(w_dff_A_AKunf6VD6_0),.clk(gclk));
	jdff dff_A_diOA7yQC8_0(.dout(w_dff_A_6x0iqUGO1_0),.din(w_dff_A_diOA7yQC8_0),.clk(gclk));
	jdff dff_A_6x0iqUGO1_0(.dout(w_dff_A_0JqbgIkv3_0),.din(w_dff_A_6x0iqUGO1_0),.clk(gclk));
	jdff dff_A_0JqbgIkv3_0(.dout(w_dff_A_U3pZZzgv1_0),.din(w_dff_A_0JqbgIkv3_0),.clk(gclk));
	jdff dff_A_U3pZZzgv1_0(.dout(w_dff_A_lc6C4k3M5_0),.din(w_dff_A_U3pZZzgv1_0),.clk(gclk));
	jdff dff_A_lc6C4k3M5_0(.dout(w_dff_A_AogsuvoC4_0),.din(w_dff_A_lc6C4k3M5_0),.clk(gclk));
	jdff dff_A_AogsuvoC4_0(.dout(w_dff_A_hA0u7aOT5_0),.din(w_dff_A_AogsuvoC4_0),.clk(gclk));
	jdff dff_A_hA0u7aOT5_0(.dout(w_dff_A_GKh59UX61_0),.din(w_dff_A_hA0u7aOT5_0),.clk(gclk));
	jdff dff_A_GKh59UX61_0(.dout(w_dff_A_TutI7v6w2_0),.din(w_dff_A_GKh59UX61_0),.clk(gclk));
	jdff dff_A_TutI7v6w2_0(.dout(w_dff_A_IHwdLI531_0),.din(w_dff_A_TutI7v6w2_0),.clk(gclk));
	jdff dff_A_IHwdLI531_0(.dout(w_dff_A_TWSbq6RZ2_0),.din(w_dff_A_IHwdLI531_0),.clk(gclk));
	jdff dff_A_TWSbq6RZ2_0(.dout(w_dff_A_84BhZORN9_0),.din(w_dff_A_TWSbq6RZ2_0),.clk(gclk));
	jdff dff_A_84BhZORN9_0(.dout(w_dff_A_eEijS2vl3_0),.din(w_dff_A_84BhZORN9_0),.clk(gclk));
	jdff dff_A_eEijS2vl3_0(.dout(w_dff_A_N6hh6wCw7_0),.din(w_dff_A_eEijS2vl3_0),.clk(gclk));
	jdff dff_A_N6hh6wCw7_0(.dout(w_dff_A_tR0UUYRn2_0),.din(w_dff_A_N6hh6wCw7_0),.clk(gclk));
	jdff dff_A_tR0UUYRn2_0(.dout(w_dff_A_sKPHJm6Z0_0),.din(w_dff_A_tR0UUYRn2_0),.clk(gclk));
	jdff dff_A_sKPHJm6Z0_0(.dout(G447gat),.din(w_dff_A_sKPHJm6Z0_0),.clk(gclk));
	jdff dff_A_jR1N3iZq0_2(.dout(w_dff_A_cKyxqtlf9_0),.din(w_dff_A_jR1N3iZq0_2),.clk(gclk));
	jdff dff_A_cKyxqtlf9_0(.dout(w_dff_A_KFJitIqo3_0),.din(w_dff_A_cKyxqtlf9_0),.clk(gclk));
	jdff dff_A_KFJitIqo3_0(.dout(w_dff_A_aAVUwLZq8_0),.din(w_dff_A_KFJitIqo3_0),.clk(gclk));
	jdff dff_A_aAVUwLZq8_0(.dout(w_dff_A_xB2QAPUt3_0),.din(w_dff_A_aAVUwLZq8_0),.clk(gclk));
	jdff dff_A_xB2QAPUt3_0(.dout(w_dff_A_PcKBPz9O4_0),.din(w_dff_A_xB2QAPUt3_0),.clk(gclk));
	jdff dff_A_PcKBPz9O4_0(.dout(w_dff_A_gpeQwYZV5_0),.din(w_dff_A_PcKBPz9O4_0),.clk(gclk));
	jdff dff_A_gpeQwYZV5_0(.dout(w_dff_A_u95OFNOR2_0),.din(w_dff_A_gpeQwYZV5_0),.clk(gclk));
	jdff dff_A_u95OFNOR2_0(.dout(w_dff_A_Rm6YChnj1_0),.din(w_dff_A_u95OFNOR2_0),.clk(gclk));
	jdff dff_A_Rm6YChnj1_0(.dout(w_dff_A_LgKvJU7O5_0),.din(w_dff_A_Rm6YChnj1_0),.clk(gclk));
	jdff dff_A_LgKvJU7O5_0(.dout(w_dff_A_eUy7NZfC5_0),.din(w_dff_A_LgKvJU7O5_0),.clk(gclk));
	jdff dff_A_eUy7NZfC5_0(.dout(w_dff_A_U3Z5fkzs6_0),.din(w_dff_A_eUy7NZfC5_0),.clk(gclk));
	jdff dff_A_U3Z5fkzs6_0(.dout(w_dff_A_e75DRMSb7_0),.din(w_dff_A_U3Z5fkzs6_0),.clk(gclk));
	jdff dff_A_e75DRMSb7_0(.dout(w_dff_A_RyoJMhlL3_0),.din(w_dff_A_e75DRMSb7_0),.clk(gclk));
	jdff dff_A_RyoJMhlL3_0(.dout(w_dff_A_rVhWEfiY7_0),.din(w_dff_A_RyoJMhlL3_0),.clk(gclk));
	jdff dff_A_rVhWEfiY7_0(.dout(w_dff_A_1ScZ9tJJ4_0),.din(w_dff_A_rVhWEfiY7_0),.clk(gclk));
	jdff dff_A_1ScZ9tJJ4_0(.dout(w_dff_A_pdf2ggUj7_0),.din(w_dff_A_1ScZ9tJJ4_0),.clk(gclk));
	jdff dff_A_pdf2ggUj7_0(.dout(w_dff_A_sfPjeD881_0),.din(w_dff_A_pdf2ggUj7_0),.clk(gclk));
	jdff dff_A_sfPjeD881_0(.dout(G448gat),.din(w_dff_A_sfPjeD881_0),.clk(gclk));
	jdff dff_A_jogfoXaH2_2(.dout(w_dff_A_PYaA5tuj5_0),.din(w_dff_A_jogfoXaH2_2),.clk(gclk));
	jdff dff_A_PYaA5tuj5_0(.dout(w_dff_A_8RcVT56I6_0),.din(w_dff_A_PYaA5tuj5_0),.clk(gclk));
	jdff dff_A_8RcVT56I6_0(.dout(w_dff_A_UxH3WkMn3_0),.din(w_dff_A_8RcVT56I6_0),.clk(gclk));
	jdff dff_A_UxH3WkMn3_0(.dout(w_dff_A_6oV0JVcf2_0),.din(w_dff_A_UxH3WkMn3_0),.clk(gclk));
	jdff dff_A_6oV0JVcf2_0(.dout(w_dff_A_1GYLlQJV4_0),.din(w_dff_A_6oV0JVcf2_0),.clk(gclk));
	jdff dff_A_1GYLlQJV4_0(.dout(w_dff_A_Ynr23nDp5_0),.din(w_dff_A_1GYLlQJV4_0),.clk(gclk));
	jdff dff_A_Ynr23nDp5_0(.dout(w_dff_A_28voCodS5_0),.din(w_dff_A_Ynr23nDp5_0),.clk(gclk));
	jdff dff_A_28voCodS5_0(.dout(w_dff_A_3NcJpqE30_0),.din(w_dff_A_28voCodS5_0),.clk(gclk));
	jdff dff_A_3NcJpqE30_0(.dout(w_dff_A_AcuqVTbn3_0),.din(w_dff_A_3NcJpqE30_0),.clk(gclk));
	jdff dff_A_AcuqVTbn3_0(.dout(w_dff_A_HnjujpJY0_0),.din(w_dff_A_AcuqVTbn3_0),.clk(gclk));
	jdff dff_A_HnjujpJY0_0(.dout(w_dff_A_fui5hW7b7_0),.din(w_dff_A_HnjujpJY0_0),.clk(gclk));
	jdff dff_A_fui5hW7b7_0(.dout(w_dff_A_SltGA6xd8_0),.din(w_dff_A_fui5hW7b7_0),.clk(gclk));
	jdff dff_A_SltGA6xd8_0(.dout(w_dff_A_UFtlop9h0_0),.din(w_dff_A_SltGA6xd8_0),.clk(gclk));
	jdff dff_A_UFtlop9h0_0(.dout(w_dff_A_AGZUqGvm6_0),.din(w_dff_A_UFtlop9h0_0),.clk(gclk));
	jdff dff_A_AGZUqGvm6_0(.dout(w_dff_A_1rhL1QCK2_0),.din(w_dff_A_AGZUqGvm6_0),.clk(gclk));
	jdff dff_A_1rhL1QCK2_0(.dout(w_dff_A_rcbqH4gR9_0),.din(w_dff_A_1rhL1QCK2_0),.clk(gclk));
	jdff dff_A_rcbqH4gR9_0(.dout(w_dff_A_YeEfp5zb8_0),.din(w_dff_A_rcbqH4gR9_0),.clk(gclk));
	jdff dff_A_YeEfp5zb8_0(.dout(G449gat),.din(w_dff_A_YeEfp5zb8_0),.clk(gclk));
	jdff dff_A_6SYhABzE8_2(.dout(w_dff_A_U9l8KWph0_0),.din(w_dff_A_6SYhABzE8_2),.clk(gclk));
	jdff dff_A_U9l8KWph0_0(.dout(w_dff_A_xTRv7I7J8_0),.din(w_dff_A_U9l8KWph0_0),.clk(gclk));
	jdff dff_A_xTRv7I7J8_0(.dout(w_dff_A_4Lor9QnW8_0),.din(w_dff_A_xTRv7I7J8_0),.clk(gclk));
	jdff dff_A_4Lor9QnW8_0(.dout(w_dff_A_9BnkiIt54_0),.din(w_dff_A_4Lor9QnW8_0),.clk(gclk));
	jdff dff_A_9BnkiIt54_0(.dout(w_dff_A_qWsc6p1C4_0),.din(w_dff_A_9BnkiIt54_0),.clk(gclk));
	jdff dff_A_qWsc6p1C4_0(.dout(w_dff_A_SaDm0roK8_0),.din(w_dff_A_qWsc6p1C4_0),.clk(gclk));
	jdff dff_A_SaDm0roK8_0(.dout(w_dff_A_yD6iCniA3_0),.din(w_dff_A_SaDm0roK8_0),.clk(gclk));
	jdff dff_A_yD6iCniA3_0(.dout(w_dff_A_1hnQitfW9_0),.din(w_dff_A_yD6iCniA3_0),.clk(gclk));
	jdff dff_A_1hnQitfW9_0(.dout(w_dff_A_ef7ZwlsO4_0),.din(w_dff_A_1hnQitfW9_0),.clk(gclk));
	jdff dff_A_ef7ZwlsO4_0(.dout(w_dff_A_U6BkSmyZ6_0),.din(w_dff_A_ef7ZwlsO4_0),.clk(gclk));
	jdff dff_A_U6BkSmyZ6_0(.dout(w_dff_A_zsV6ZeO50_0),.din(w_dff_A_U6BkSmyZ6_0),.clk(gclk));
	jdff dff_A_zsV6ZeO50_0(.dout(w_dff_A_qSKnGyur4_0),.din(w_dff_A_zsV6ZeO50_0),.clk(gclk));
	jdff dff_A_qSKnGyur4_0(.dout(w_dff_A_MSmYgbIt5_0),.din(w_dff_A_qSKnGyur4_0),.clk(gclk));
	jdff dff_A_MSmYgbIt5_0(.dout(w_dff_A_QUDYou8I0_0),.din(w_dff_A_MSmYgbIt5_0),.clk(gclk));
	jdff dff_A_QUDYou8I0_0(.dout(w_dff_A_nZhjkkeD8_0),.din(w_dff_A_QUDYou8I0_0),.clk(gclk));
	jdff dff_A_nZhjkkeD8_0(.dout(w_dff_A_CwiNN6iy1_0),.din(w_dff_A_nZhjkkeD8_0),.clk(gclk));
	jdff dff_A_CwiNN6iy1_0(.dout(w_dff_A_Jg3GDmmY5_0),.din(w_dff_A_CwiNN6iy1_0),.clk(gclk));
	jdff dff_A_Jg3GDmmY5_0(.dout(w_dff_A_hXxK4DLd5_0),.din(w_dff_A_Jg3GDmmY5_0),.clk(gclk));
	jdff dff_A_hXxK4DLd5_0(.dout(G450gat),.din(w_dff_A_hXxK4DLd5_0),.clk(gclk));
	jdff dff_A_HjMSVorL4_2(.dout(w_dff_A_8d8VRant6_0),.din(w_dff_A_HjMSVorL4_2),.clk(gclk));
	jdff dff_A_8d8VRant6_0(.dout(w_dff_A_EPf7X4f57_0),.din(w_dff_A_8d8VRant6_0),.clk(gclk));
	jdff dff_A_EPf7X4f57_0(.dout(w_dff_A_3QNGAKnf1_0),.din(w_dff_A_EPf7X4f57_0),.clk(gclk));
	jdff dff_A_3QNGAKnf1_0(.dout(w_dff_A_EATE4LbZ5_0),.din(w_dff_A_3QNGAKnf1_0),.clk(gclk));
	jdff dff_A_EATE4LbZ5_0(.dout(w_dff_A_pxwTyGmv4_0),.din(w_dff_A_EATE4LbZ5_0),.clk(gclk));
	jdff dff_A_pxwTyGmv4_0(.dout(w_dff_A_Jhd9VjBL5_0),.din(w_dff_A_pxwTyGmv4_0),.clk(gclk));
	jdff dff_A_Jhd9VjBL5_0(.dout(w_dff_A_iagwmn7t7_0),.din(w_dff_A_Jhd9VjBL5_0),.clk(gclk));
	jdff dff_A_iagwmn7t7_0(.dout(w_dff_A_SC21QAg04_0),.din(w_dff_A_iagwmn7t7_0),.clk(gclk));
	jdff dff_A_SC21QAg04_0(.dout(w_dff_A_5riHEL4U7_0),.din(w_dff_A_SC21QAg04_0),.clk(gclk));
	jdff dff_A_5riHEL4U7_0(.dout(w_dff_A_UNBskL4w0_0),.din(w_dff_A_5riHEL4U7_0),.clk(gclk));
	jdff dff_A_UNBskL4w0_0(.dout(w_dff_A_3KoqT49O3_0),.din(w_dff_A_UNBskL4w0_0),.clk(gclk));
	jdff dff_A_3KoqT49O3_0(.dout(w_dff_A_1gvU1Uhq7_0),.din(w_dff_A_3KoqT49O3_0),.clk(gclk));
	jdff dff_A_1gvU1Uhq7_0(.dout(w_dff_A_F60jt1aF1_0),.din(w_dff_A_1gvU1Uhq7_0),.clk(gclk));
	jdff dff_A_F60jt1aF1_0(.dout(w_dff_A_H7c7vsDf8_0),.din(w_dff_A_F60jt1aF1_0),.clk(gclk));
	jdff dff_A_H7c7vsDf8_0(.dout(w_dff_A_0dm0PEOh3_0),.din(w_dff_A_H7c7vsDf8_0),.clk(gclk));
	jdff dff_A_0dm0PEOh3_0(.dout(w_dff_A_0hgwa0Rq2_0),.din(w_dff_A_0dm0PEOh3_0),.clk(gclk));
	jdff dff_A_0hgwa0Rq2_0(.dout(G767gat),.din(w_dff_A_0hgwa0Rq2_0),.clk(gclk));
	jdff dff_A_joxD1bRl8_2(.dout(w_dff_A_J13CEXhl5_0),.din(w_dff_A_joxD1bRl8_2),.clk(gclk));
	jdff dff_A_J13CEXhl5_0(.dout(w_dff_A_pOIz6fq12_0),.din(w_dff_A_J13CEXhl5_0),.clk(gclk));
	jdff dff_A_pOIz6fq12_0(.dout(w_dff_A_dovxfJBW0_0),.din(w_dff_A_pOIz6fq12_0),.clk(gclk));
	jdff dff_A_dovxfJBW0_0(.dout(w_dff_A_0dVxO6IS7_0),.din(w_dff_A_dovxfJBW0_0),.clk(gclk));
	jdff dff_A_0dVxO6IS7_0(.dout(w_dff_A_ZiItk0eJ5_0),.din(w_dff_A_0dVxO6IS7_0),.clk(gclk));
	jdff dff_A_ZiItk0eJ5_0(.dout(w_dff_A_gDherlCp1_0),.din(w_dff_A_ZiItk0eJ5_0),.clk(gclk));
	jdff dff_A_gDherlCp1_0(.dout(w_dff_A_s5VJe8cS8_0),.din(w_dff_A_gDherlCp1_0),.clk(gclk));
	jdff dff_A_s5VJe8cS8_0(.dout(w_dff_A_83wDDOFU6_0),.din(w_dff_A_s5VJe8cS8_0),.clk(gclk));
	jdff dff_A_83wDDOFU6_0(.dout(w_dff_A_l8jVQVac7_0),.din(w_dff_A_83wDDOFU6_0),.clk(gclk));
	jdff dff_A_l8jVQVac7_0(.dout(w_dff_A_y59X553Y8_0),.din(w_dff_A_l8jVQVac7_0),.clk(gclk));
	jdff dff_A_y59X553Y8_0(.dout(w_dff_A_QtGCyVVl8_0),.din(w_dff_A_y59X553Y8_0),.clk(gclk));
	jdff dff_A_QtGCyVVl8_0(.dout(w_dff_A_yqlYxW6i3_0),.din(w_dff_A_QtGCyVVl8_0),.clk(gclk));
	jdff dff_A_yqlYxW6i3_0(.dout(w_dff_A_BFFUtggX3_0),.din(w_dff_A_yqlYxW6i3_0),.clk(gclk));
	jdff dff_A_BFFUtggX3_0(.dout(w_dff_A_muWherAh0_0),.din(w_dff_A_BFFUtggX3_0),.clk(gclk));
	jdff dff_A_muWherAh0_0(.dout(w_dff_A_77Yh6PNd4_0),.din(w_dff_A_muWherAh0_0),.clk(gclk));
	jdff dff_A_77Yh6PNd4_0(.dout(w_dff_A_aDEixSED6_0),.din(w_dff_A_77Yh6PNd4_0),.clk(gclk));
	jdff dff_A_aDEixSED6_0(.dout(G768gat),.din(w_dff_A_aDEixSED6_0),.clk(gclk));
	jdff dff_A_Hgt1Xa0m0_2(.dout(w_dff_A_vHjowtHT0_0),.din(w_dff_A_Hgt1Xa0m0_2),.clk(gclk));
	jdff dff_A_vHjowtHT0_0(.dout(w_dff_A_ncYT3LV94_0),.din(w_dff_A_vHjowtHT0_0),.clk(gclk));
	jdff dff_A_ncYT3LV94_0(.dout(w_dff_A_YumxXzvL1_0),.din(w_dff_A_ncYT3LV94_0),.clk(gclk));
	jdff dff_A_YumxXzvL1_0(.dout(w_dff_A_hQfwjWuz3_0),.din(w_dff_A_YumxXzvL1_0),.clk(gclk));
	jdff dff_A_hQfwjWuz3_0(.dout(w_dff_A_mtW0mJYG9_0),.din(w_dff_A_hQfwjWuz3_0),.clk(gclk));
	jdff dff_A_mtW0mJYG9_0(.dout(w_dff_A_kAG5UFsj0_0),.din(w_dff_A_mtW0mJYG9_0),.clk(gclk));
	jdff dff_A_kAG5UFsj0_0(.dout(w_dff_A_Ik4L36mt5_0),.din(w_dff_A_kAG5UFsj0_0),.clk(gclk));
	jdff dff_A_Ik4L36mt5_0(.dout(G850gat),.din(w_dff_A_Ik4L36mt5_0),.clk(gclk));
	jdff dff_A_6DjvaEd45_2(.dout(w_dff_A_7hJsL7Kz2_0),.din(w_dff_A_6DjvaEd45_2),.clk(gclk));
	jdff dff_A_7hJsL7Kz2_0(.dout(w_dff_A_ioXI4HxI9_0),.din(w_dff_A_7hJsL7Kz2_0),.clk(gclk));
	jdff dff_A_ioXI4HxI9_0(.dout(w_dff_A_jdt7MhOb7_0),.din(w_dff_A_ioXI4HxI9_0),.clk(gclk));
	jdff dff_A_jdt7MhOb7_0(.dout(G863gat),.din(w_dff_A_jdt7MhOb7_0),.clk(gclk));
	jdff dff_A_Yomum5wG5_2(.dout(w_dff_A_CaOgh5Yg7_0),.din(w_dff_A_Yomum5wG5_2),.clk(gclk));
	jdff dff_A_CaOgh5Yg7_0(.dout(w_dff_A_pL78jcLq3_0),.din(w_dff_A_CaOgh5Yg7_0),.clk(gclk));
	jdff dff_A_pL78jcLq3_0(.dout(w_dff_A_9hyLUzWt7_0),.din(w_dff_A_pL78jcLq3_0),.clk(gclk));
	jdff dff_A_9hyLUzWt7_0(.dout(G864gat),.din(w_dff_A_9hyLUzWt7_0),.clk(gclk));
	jdff dff_A_WotfRuLH0_2(.dout(w_dff_A_3r6LbCBP9_0),.din(w_dff_A_WotfRuLH0_2),.clk(gclk));
	jdff dff_A_3r6LbCBP9_0(.dout(w_dff_A_fps8k8ed6_0),.din(w_dff_A_3r6LbCBP9_0),.clk(gclk));
	jdff dff_A_fps8k8ed6_0(.dout(w_dff_A_e70X0dyi0_0),.din(w_dff_A_fps8k8ed6_0),.clk(gclk));
	jdff dff_A_e70X0dyi0_0(.dout(w_dff_A_1VAwtGq65_0),.din(w_dff_A_e70X0dyi0_0),.clk(gclk));
	jdff dff_A_1VAwtGq65_0(.dout(w_dff_A_ksBZVi5i8_0),.din(w_dff_A_1VAwtGq65_0),.clk(gclk));
	jdff dff_A_ksBZVi5i8_0(.dout(G865gat),.din(w_dff_A_ksBZVi5i8_0),.clk(gclk));
	jdff dff_A_Fm9M2ftm8_2(.dout(w_dff_A_zB1UnxD10_0),.din(w_dff_A_Fm9M2ftm8_2),.clk(gclk));
	jdff dff_A_zB1UnxD10_0(.dout(G866gat),.din(w_dff_A_zB1UnxD10_0),.clk(gclk));
	jdff dff_A_Pv2dfkZ83_2(.dout(w_dff_A_sW3hjTUa3_0),.din(w_dff_A_Pv2dfkZ83_2),.clk(gclk));
	jdff dff_A_sW3hjTUa3_0(.dout(G874gat),.din(w_dff_A_sW3hjTUa3_0),.clk(gclk));
endmodule

