/*

top:
	jspl: 724
	jspl3: 1211
	jnot: 7
	jand: 1749
	jor: 1404

Summary:
	jspl: 724
	jspl3: 1211
	jnot: 7
	jand: 1749
	jor: 1404

The maximum logic level gap of any gate:
	top: 11
*/

module rf_bar(gclk, a0, a1, a2, a3, a4, a5, a6, a7, a8, a9, a10, a11, a12, a13, a14, a15, a16, a17, a18, a19, a20, a21, a22, a23, a24, a25, a26, a27, a28, a29, a30, a31, a32, a33, a34, a35, a36, a37, a38, a39, a40, a41, a42, a43, a44, a45, a46, a47, a48, a49, a50, a51, a52, a53, a54, a55, a56, a57, a58, a59, a60, a61, a62, a63, a64, a65, a66, a67, a68, a69, a70, a71, a72, a73, a74, a75, a76, a77, a78, a79, a80, a81, a82, a83, a84, a85, a86, a87, a88, a89, a90, a91, a92, a93, a94, a95, a96, a97, a98, a99, a100, a101, a102, a103, a104, a105, a106, a107, a108, a109, a110, a111, a112, a113, a114, a115, a116, a117, a118, a119, a120, a121, a122, a123, a124, a125, a126, a127, shift0, shift1, shift2, shift3, shift4, shift5, shift6, result0, result1, result2, result3, result4, result5, result6, result7, result8, result9, result10, result11, result12, result13, result14, result15, result16, result17, result18, result19, result20, result21, result22, result23, result24, result25, result26, result27, result28, result29, result30, result31, result32, result33, result34, result35, result36, result37, result38, result39, result40, result41, result42, result43, result44, result45, result46, result47, result48, result49, result50, result51, result52, result53, result54, result55, result56, result57, result58, result59, result60, result61, result62, result63, result64, result65, result66, result67, result68, result69, result70, result71, result72, result73, result74, result75, result76, result77, result78, result79, result80, result81, result82, result83, result84, result85, result86, result87, result88, result89, result90, result91, result92, result93, result94, result95, result96, result97, result98, result99, result100, result101, result102, result103, result104, result105, result106, result107, result108, result109, result110, result111, result112, result113, result114, result115, result116, result117, result118, result119, result120, result121, result122, result123, result124, result125, result126, result127);
	input gclk;
	input a0;
	input a1;
	input a2;
	input a3;
	input a4;
	input a5;
	input a6;
	input a7;
	input a8;
	input a9;
	input a10;
	input a11;
	input a12;
	input a13;
	input a14;
	input a15;
	input a16;
	input a17;
	input a18;
	input a19;
	input a20;
	input a21;
	input a22;
	input a23;
	input a24;
	input a25;
	input a26;
	input a27;
	input a28;
	input a29;
	input a30;
	input a31;
	input a32;
	input a33;
	input a34;
	input a35;
	input a36;
	input a37;
	input a38;
	input a39;
	input a40;
	input a41;
	input a42;
	input a43;
	input a44;
	input a45;
	input a46;
	input a47;
	input a48;
	input a49;
	input a50;
	input a51;
	input a52;
	input a53;
	input a54;
	input a55;
	input a56;
	input a57;
	input a58;
	input a59;
	input a60;
	input a61;
	input a62;
	input a63;
	input a64;
	input a65;
	input a66;
	input a67;
	input a68;
	input a69;
	input a70;
	input a71;
	input a72;
	input a73;
	input a74;
	input a75;
	input a76;
	input a77;
	input a78;
	input a79;
	input a80;
	input a81;
	input a82;
	input a83;
	input a84;
	input a85;
	input a86;
	input a87;
	input a88;
	input a89;
	input a90;
	input a91;
	input a92;
	input a93;
	input a94;
	input a95;
	input a96;
	input a97;
	input a98;
	input a99;
	input a100;
	input a101;
	input a102;
	input a103;
	input a104;
	input a105;
	input a106;
	input a107;
	input a108;
	input a109;
	input a110;
	input a111;
	input a112;
	input a113;
	input a114;
	input a115;
	input a116;
	input a117;
	input a118;
	input a119;
	input a120;
	input a121;
	input a122;
	input a123;
	input a124;
	input a125;
	input a126;
	input a127;
	input shift0;
	input shift1;
	input shift2;
	input shift3;
	input shift4;
	input shift5;
	input shift6;
	output result0;
	output result1;
	output result2;
	output result3;
	output result4;
	output result5;
	output result6;
	output result7;
	output result8;
	output result9;
	output result10;
	output result11;
	output result12;
	output result13;
	output result14;
	output result15;
	output result16;
	output result17;
	output result18;
	output result19;
	output result20;
	output result21;
	output result22;
	output result23;
	output result24;
	output result25;
	output result26;
	output result27;
	output result28;
	output result29;
	output result30;
	output result31;
	output result32;
	output result33;
	output result34;
	output result35;
	output result36;
	output result37;
	output result38;
	output result39;
	output result40;
	output result41;
	output result42;
	output result43;
	output result44;
	output result45;
	output result46;
	output result47;
	output result48;
	output result49;
	output result50;
	output result51;
	output result52;
	output result53;
	output result54;
	output result55;
	output result56;
	output result57;
	output result58;
	output result59;
	output result60;
	output result61;
	output result62;
	output result63;
	output result64;
	output result65;
	output result66;
	output result67;
	output result68;
	output result69;
	output result70;
	output result71;
	output result72;
	output result73;
	output result74;
	output result75;
	output result76;
	output result77;
	output result78;
	output result79;
	output result80;
	output result81;
	output result82;
	output result83;
	output result84;
	output result85;
	output result86;
	output result87;
	output result88;
	output result89;
	output result90;
	output result91;
	output result92;
	output result93;
	output result94;
	output result95;
	output result96;
	output result97;
	output result98;
	output result99;
	output result100;
	output result101;
	output result102;
	output result103;
	output result104;
	output result105;
	output result106;
	output result107;
	output result108;
	output result109;
	output result110;
	output result111;
	output result112;
	output result113;
	output result114;
	output result115;
	output result116;
	output result117;
	output result118;
	output result119;
	output result120;
	output result121;
	output result122;
	output result123;
	output result124;
	output result125;
	output result126;
	output result127;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1837;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire n1852;
	wire n1853;
	wire n1854;
	wire n1855;
	wire n1856;
	wire n1857;
	wire n1858;
	wire n1859;
	wire n1860;
	wire n1861;
	wire n1862;
	wire n1863;
	wire n1864;
	wire n1865;
	wire n1866;
	wire n1867;
	wire n1868;
	wire n1869;
	wire n1870;
	wire n1871;
	wire n1872;
	wire n1873;
	wire n1874;
	wire n1875;
	wire n1876;
	wire n1877;
	wire n1878;
	wire n1879;
	wire n1880;
	wire n1881;
	wire n1882;
	wire n1883;
	wire n1884;
	wire n1885;
	wire n1886;
	wire n1887;
	wire n1888;
	wire n1889;
	wire n1890;
	wire n1891;
	wire n1892;
	wire n1893;
	wire n1894;
	wire n1895;
	wire n1896;
	wire n1897;
	wire n1898;
	wire n1899;
	wire n1900;
	wire n1901;
	wire n1902;
	wire n1904;
	wire n1905;
	wire n1906;
	wire n1907;
	wire n1908;
	wire n1909;
	wire n1910;
	wire n1911;
	wire n1912;
	wire n1913;
	wire n1914;
	wire n1915;
	wire n1916;
	wire n1917;
	wire n1918;
	wire n1919;
	wire n1920;
	wire n1921;
	wire n1922;
	wire n1923;
	wire n1924;
	wire n1925;
	wire n1926;
	wire n1927;
	wire n1928;
	wire n1929;
	wire n1930;
	wire n1931;
	wire n1932;
	wire n1933;
	wire n1934;
	wire n1935;
	wire n1936;
	wire n1937;
	wire n1938;
	wire n1939;
	wire n1940;
	wire n1941;
	wire n1942;
	wire n1943;
	wire n1944;
	wire n1945;
	wire n1946;
	wire n1947;
	wire n1948;
	wire n1949;
	wire n1950;
	wire n1951;
	wire n1952;
	wire n1953;
	wire n1954;
	wire n1955;
	wire n1956;
	wire n1957;
	wire n1958;
	wire n1959;
	wire n1960;
	wire n1961;
	wire n1962;
	wire n1963;
	wire n1964;
	wire n1965;
	wire n1966;
	wire n1967;
	wire n1968;
	wire n1969;
	wire n1970;
	wire n1971;
	wire n1972;
	wire n1973;
	wire n1974;
	wire n1975;
	wire n1977;
	wire n1978;
	wire n1979;
	wire n1980;
	wire n1981;
	wire n1982;
	wire n1983;
	wire n1984;
	wire n1985;
	wire n1986;
	wire n1987;
	wire n1988;
	wire n1989;
	wire n1990;
	wire n1991;
	wire n1992;
	wire n1993;
	wire n1994;
	wire n1995;
	wire n1996;
	wire n1997;
	wire n1998;
	wire n1999;
	wire n2000;
	wire n2001;
	wire n2002;
	wire n2003;
	wire n2004;
	wire n2005;
	wire n2006;
	wire n2007;
	wire n2008;
	wire n2009;
	wire n2010;
	wire n2011;
	wire n2012;
	wire n2013;
	wire n2014;
	wire n2015;
	wire n2016;
	wire n2017;
	wire n2018;
	wire n2019;
	wire n2020;
	wire n2021;
	wire n2022;
	wire n2023;
	wire n2024;
	wire n2025;
	wire n2026;
	wire n2027;
	wire n2028;
	wire n2029;
	wire n2030;
	wire n2031;
	wire n2032;
	wire n2033;
	wire n2034;
	wire n2035;
	wire n2036;
	wire n2037;
	wire n2038;
	wire n2039;
	wire n2040;
	wire n2041;
	wire n2042;
	wire n2043;
	wire n2044;
	wire n2045;
	wire n2046;
	wire n2047;
	wire n2048;
	wire n2050;
	wire n2051;
	wire n2052;
	wire n2053;
	wire n2054;
	wire n2055;
	wire n2056;
	wire n2057;
	wire n2058;
	wire n2059;
	wire n2060;
	wire n2061;
	wire n2062;
	wire n2063;
	wire n2064;
	wire n2065;
	wire n2066;
	wire n2067;
	wire n2068;
	wire n2069;
	wire n2070;
	wire n2071;
	wire n2072;
	wire n2073;
	wire n2074;
	wire n2075;
	wire n2076;
	wire n2077;
	wire n2078;
	wire n2079;
	wire n2080;
	wire n2081;
	wire n2082;
	wire n2083;
	wire n2084;
	wire n2085;
	wire n2086;
	wire n2087;
	wire n2088;
	wire n2089;
	wire n2090;
	wire n2091;
	wire n2092;
	wire n2093;
	wire n2094;
	wire n2095;
	wire n2096;
	wire n2097;
	wire n2098;
	wire n2099;
	wire n2100;
	wire n2101;
	wire n2102;
	wire n2103;
	wire n2104;
	wire n2105;
	wire n2106;
	wire n2107;
	wire n2108;
	wire n2109;
	wire n2110;
	wire n2111;
	wire n2112;
	wire n2113;
	wire n2114;
	wire n2115;
	wire n2116;
	wire n2117;
	wire n2118;
	wire n2119;
	wire n2120;
	wire n2121;
	wire n2123;
	wire n2124;
	wire n2125;
	wire n2126;
	wire n2127;
	wire n2128;
	wire n2129;
	wire n2130;
	wire n2131;
	wire n2132;
	wire n2133;
	wire n2134;
	wire n2135;
	wire n2136;
	wire n2137;
	wire n2138;
	wire n2139;
	wire n2140;
	wire n2141;
	wire n2142;
	wire n2143;
	wire n2144;
	wire n2145;
	wire n2146;
	wire n2147;
	wire n2148;
	wire n2149;
	wire n2150;
	wire n2151;
	wire n2152;
	wire n2153;
	wire n2154;
	wire n2155;
	wire n2156;
	wire n2157;
	wire n2158;
	wire n2159;
	wire n2160;
	wire n2161;
	wire n2162;
	wire n2163;
	wire n2164;
	wire n2165;
	wire n2166;
	wire n2167;
	wire n2168;
	wire n2169;
	wire n2170;
	wire n2171;
	wire n2172;
	wire n2173;
	wire n2174;
	wire n2175;
	wire n2176;
	wire n2177;
	wire n2178;
	wire n2179;
	wire n2180;
	wire n2181;
	wire n2182;
	wire n2183;
	wire n2184;
	wire n2185;
	wire n2186;
	wire n2187;
	wire n2188;
	wire n2189;
	wire n2190;
	wire n2191;
	wire n2192;
	wire n2193;
	wire n2194;
	wire n2196;
	wire n2197;
	wire n2198;
	wire n2199;
	wire n2200;
	wire n2201;
	wire n2202;
	wire n2203;
	wire n2204;
	wire n2205;
	wire n2206;
	wire n2207;
	wire n2208;
	wire n2209;
	wire n2210;
	wire n2211;
	wire n2212;
	wire n2213;
	wire n2214;
	wire n2215;
	wire n2216;
	wire n2217;
	wire n2218;
	wire n2219;
	wire n2220;
	wire n2221;
	wire n2222;
	wire n2223;
	wire n2224;
	wire n2225;
	wire n2226;
	wire n2227;
	wire n2228;
	wire n2229;
	wire n2230;
	wire n2231;
	wire n2232;
	wire n2233;
	wire n2234;
	wire n2235;
	wire n2236;
	wire n2237;
	wire n2238;
	wire n2239;
	wire n2240;
	wire n2241;
	wire n2242;
	wire n2243;
	wire n2244;
	wire n2245;
	wire n2246;
	wire n2247;
	wire n2248;
	wire n2249;
	wire n2250;
	wire n2251;
	wire n2252;
	wire n2253;
	wire n2254;
	wire n2255;
	wire n2256;
	wire n2257;
	wire n2258;
	wire n2259;
	wire n2260;
	wire n2261;
	wire n2262;
	wire n2263;
	wire n2264;
	wire n2265;
	wire n2266;
	wire n2267;
	wire n2269;
	wire n2270;
	wire n2271;
	wire n2272;
	wire n2273;
	wire n2274;
	wire n2275;
	wire n2276;
	wire n2277;
	wire n2278;
	wire n2279;
	wire n2280;
	wire n2281;
	wire n2282;
	wire n2283;
	wire n2284;
	wire n2285;
	wire n2286;
	wire n2287;
	wire n2288;
	wire n2289;
	wire n2290;
	wire n2291;
	wire n2292;
	wire n2293;
	wire n2294;
	wire n2295;
	wire n2296;
	wire n2297;
	wire n2298;
	wire n2299;
	wire n2300;
	wire n2301;
	wire n2302;
	wire n2303;
	wire n2304;
	wire n2305;
	wire n2306;
	wire n2307;
	wire n2308;
	wire n2309;
	wire n2310;
	wire n2311;
	wire n2312;
	wire n2313;
	wire n2314;
	wire n2315;
	wire n2316;
	wire n2317;
	wire n2318;
	wire n2319;
	wire n2320;
	wire n2321;
	wire n2322;
	wire n2323;
	wire n2324;
	wire n2325;
	wire n2326;
	wire n2327;
	wire n2328;
	wire n2329;
	wire n2330;
	wire n2331;
	wire n2332;
	wire n2333;
	wire n2334;
	wire n2335;
	wire n2336;
	wire n2337;
	wire n2338;
	wire n2339;
	wire n2340;
	wire n2342;
	wire n2343;
	wire n2344;
	wire n2345;
	wire n2346;
	wire n2347;
	wire n2348;
	wire n2349;
	wire n2350;
	wire n2351;
	wire n2352;
	wire n2353;
	wire n2354;
	wire n2355;
	wire n2356;
	wire n2357;
	wire n2358;
	wire n2359;
	wire n2360;
	wire n2361;
	wire n2362;
	wire n2363;
	wire n2364;
	wire n2365;
	wire n2366;
	wire n2367;
	wire n2368;
	wire n2369;
	wire n2370;
	wire n2371;
	wire n2372;
	wire n2373;
	wire n2374;
	wire n2375;
	wire n2376;
	wire n2377;
	wire n2378;
	wire n2379;
	wire n2380;
	wire n2381;
	wire n2382;
	wire n2383;
	wire n2384;
	wire n2385;
	wire n2386;
	wire n2387;
	wire n2388;
	wire n2389;
	wire n2390;
	wire n2391;
	wire n2392;
	wire n2393;
	wire n2394;
	wire n2395;
	wire n2396;
	wire n2397;
	wire n2398;
	wire n2399;
	wire n2400;
	wire n2401;
	wire n2402;
	wire n2403;
	wire n2404;
	wire n2405;
	wire n2406;
	wire n2407;
	wire n2408;
	wire n2409;
	wire n2410;
	wire n2411;
	wire n2412;
	wire n2413;
	wire n2415;
	wire n2416;
	wire n2417;
	wire n2418;
	wire n2419;
	wire n2420;
	wire n2421;
	wire n2422;
	wire n2423;
	wire n2424;
	wire n2425;
	wire n2426;
	wire n2427;
	wire n2428;
	wire n2429;
	wire n2430;
	wire n2432;
	wire n2433;
	wire n2434;
	wire n2435;
	wire n2436;
	wire n2437;
	wire n2438;
	wire n2439;
	wire n2440;
	wire n2441;
	wire n2442;
	wire n2443;
	wire n2444;
	wire n2445;
	wire n2446;
	wire n2447;
	wire n2449;
	wire n2450;
	wire n2451;
	wire n2452;
	wire n2453;
	wire n2454;
	wire n2455;
	wire n2456;
	wire n2457;
	wire n2458;
	wire n2459;
	wire n2460;
	wire n2461;
	wire n2462;
	wire n2463;
	wire n2464;
	wire n2466;
	wire n2467;
	wire n2468;
	wire n2469;
	wire n2470;
	wire n2471;
	wire n2472;
	wire n2473;
	wire n2474;
	wire n2475;
	wire n2476;
	wire n2477;
	wire n2478;
	wire n2479;
	wire n2480;
	wire n2481;
	wire n2483;
	wire n2484;
	wire n2485;
	wire n2486;
	wire n2487;
	wire n2488;
	wire n2489;
	wire n2490;
	wire n2491;
	wire n2492;
	wire n2493;
	wire n2494;
	wire n2495;
	wire n2496;
	wire n2497;
	wire n2498;
	wire n2500;
	wire n2501;
	wire n2502;
	wire n2503;
	wire n2504;
	wire n2505;
	wire n2506;
	wire n2507;
	wire n2508;
	wire n2509;
	wire n2510;
	wire n2511;
	wire n2512;
	wire n2513;
	wire n2514;
	wire n2515;
	wire n2517;
	wire n2518;
	wire n2519;
	wire n2520;
	wire n2521;
	wire n2522;
	wire n2523;
	wire n2524;
	wire n2525;
	wire n2526;
	wire n2527;
	wire n2528;
	wire n2529;
	wire n2530;
	wire n2531;
	wire n2532;
	wire n2534;
	wire n2535;
	wire n2536;
	wire n2537;
	wire n2538;
	wire n2539;
	wire n2540;
	wire n2541;
	wire n2542;
	wire n2543;
	wire n2544;
	wire n2545;
	wire n2546;
	wire n2547;
	wire n2548;
	wire n2549;
	wire n2551;
	wire n2552;
	wire n2553;
	wire n2554;
	wire n2555;
	wire n2556;
	wire n2557;
	wire n2558;
	wire n2559;
	wire n2560;
	wire n2561;
	wire n2562;
	wire n2563;
	wire n2564;
	wire n2565;
	wire n2566;
	wire n2568;
	wire n2569;
	wire n2570;
	wire n2571;
	wire n2572;
	wire n2573;
	wire n2574;
	wire n2575;
	wire n2576;
	wire n2577;
	wire n2578;
	wire n2579;
	wire n2580;
	wire n2581;
	wire n2582;
	wire n2583;
	wire n2585;
	wire n2586;
	wire n2587;
	wire n2588;
	wire n2589;
	wire n2590;
	wire n2591;
	wire n2592;
	wire n2593;
	wire n2594;
	wire n2595;
	wire n2596;
	wire n2597;
	wire n2598;
	wire n2599;
	wire n2600;
	wire n2602;
	wire n2603;
	wire n2604;
	wire n2605;
	wire n2606;
	wire n2607;
	wire n2608;
	wire n2609;
	wire n2610;
	wire n2611;
	wire n2612;
	wire n2613;
	wire n2614;
	wire n2615;
	wire n2616;
	wire n2617;
	wire n2619;
	wire n2620;
	wire n2621;
	wire n2622;
	wire n2623;
	wire n2624;
	wire n2625;
	wire n2626;
	wire n2627;
	wire n2628;
	wire n2629;
	wire n2630;
	wire n2631;
	wire n2632;
	wire n2633;
	wire n2634;
	wire n2636;
	wire n2637;
	wire n2638;
	wire n2639;
	wire n2640;
	wire n2641;
	wire n2642;
	wire n2643;
	wire n2644;
	wire n2645;
	wire n2646;
	wire n2647;
	wire n2648;
	wire n2649;
	wire n2650;
	wire n2651;
	wire n2653;
	wire n2654;
	wire n2655;
	wire n2656;
	wire n2657;
	wire n2658;
	wire n2659;
	wire n2660;
	wire n2661;
	wire n2662;
	wire n2663;
	wire n2664;
	wire n2665;
	wire n2666;
	wire n2667;
	wire n2668;
	wire n2670;
	wire n2671;
	wire n2672;
	wire n2673;
	wire n2674;
	wire n2675;
	wire n2676;
	wire n2677;
	wire n2678;
	wire n2679;
	wire n2680;
	wire n2681;
	wire n2682;
	wire n2683;
	wire n2684;
	wire n2685;
	wire n2687;
	wire n2688;
	wire n2689;
	wire n2690;
	wire n2691;
	wire n2692;
	wire n2693;
	wire n2694;
	wire n2695;
	wire n2696;
	wire n2697;
	wire n2698;
	wire n2699;
	wire n2700;
	wire n2701;
	wire n2702;
	wire n2704;
	wire n2705;
	wire n2706;
	wire n2707;
	wire n2708;
	wire n2709;
	wire n2710;
	wire n2711;
	wire n2712;
	wire n2713;
	wire n2714;
	wire n2715;
	wire n2716;
	wire n2717;
	wire n2718;
	wire n2719;
	wire n2721;
	wire n2722;
	wire n2723;
	wire n2724;
	wire n2725;
	wire n2726;
	wire n2727;
	wire n2728;
	wire n2729;
	wire n2730;
	wire n2731;
	wire n2732;
	wire n2733;
	wire n2734;
	wire n2735;
	wire n2736;
	wire n2738;
	wire n2739;
	wire n2740;
	wire n2741;
	wire n2742;
	wire n2743;
	wire n2744;
	wire n2745;
	wire n2746;
	wire n2747;
	wire n2748;
	wire n2749;
	wire n2750;
	wire n2751;
	wire n2752;
	wire n2753;
	wire n2755;
	wire n2756;
	wire n2757;
	wire n2758;
	wire n2759;
	wire n2760;
	wire n2761;
	wire n2762;
	wire n2763;
	wire n2764;
	wire n2765;
	wire n2766;
	wire n2767;
	wire n2768;
	wire n2769;
	wire n2770;
	wire n2772;
	wire n2773;
	wire n2774;
	wire n2775;
	wire n2776;
	wire n2777;
	wire n2778;
	wire n2779;
	wire n2780;
	wire n2781;
	wire n2782;
	wire n2783;
	wire n2784;
	wire n2785;
	wire n2786;
	wire n2787;
	wire n2789;
	wire n2790;
	wire n2791;
	wire n2792;
	wire n2793;
	wire n2794;
	wire n2795;
	wire n2796;
	wire n2797;
	wire n2798;
	wire n2799;
	wire n2800;
	wire n2801;
	wire n2802;
	wire n2803;
	wire n2804;
	wire n2806;
	wire n2807;
	wire n2808;
	wire n2809;
	wire n2810;
	wire n2811;
	wire n2812;
	wire n2813;
	wire n2814;
	wire n2815;
	wire n2816;
	wire n2817;
	wire n2818;
	wire n2819;
	wire n2820;
	wire n2821;
	wire n2823;
	wire n2824;
	wire n2825;
	wire n2826;
	wire n2827;
	wire n2828;
	wire n2829;
	wire n2830;
	wire n2831;
	wire n2832;
	wire n2833;
	wire n2834;
	wire n2835;
	wire n2836;
	wire n2837;
	wire n2838;
	wire n2840;
	wire n2841;
	wire n2842;
	wire n2843;
	wire n2844;
	wire n2845;
	wire n2846;
	wire n2847;
	wire n2848;
	wire n2849;
	wire n2850;
	wire n2851;
	wire n2852;
	wire n2853;
	wire n2854;
	wire n2855;
	wire n2857;
	wire n2858;
	wire n2859;
	wire n2860;
	wire n2861;
	wire n2862;
	wire n2863;
	wire n2864;
	wire n2865;
	wire n2866;
	wire n2867;
	wire n2868;
	wire n2869;
	wire n2870;
	wire n2871;
	wire n2872;
	wire n2874;
	wire n2875;
	wire n2876;
	wire n2877;
	wire n2878;
	wire n2879;
	wire n2880;
	wire n2881;
	wire n2882;
	wire n2883;
	wire n2884;
	wire n2885;
	wire n2886;
	wire n2887;
	wire n2888;
	wire n2889;
	wire n2891;
	wire n2892;
	wire n2893;
	wire n2894;
	wire n2895;
	wire n2896;
	wire n2897;
	wire n2898;
	wire n2899;
	wire n2900;
	wire n2901;
	wire n2902;
	wire n2903;
	wire n2904;
	wire n2905;
	wire n2906;
	wire n2908;
	wire n2909;
	wire n2910;
	wire n2911;
	wire n2912;
	wire n2913;
	wire n2914;
	wire n2915;
	wire n2916;
	wire n2917;
	wire n2918;
	wire n2919;
	wire n2920;
	wire n2921;
	wire n2922;
	wire n2923;
	wire n2925;
	wire n2926;
	wire n2927;
	wire n2928;
	wire n2929;
	wire n2930;
	wire n2931;
	wire n2932;
	wire n2933;
	wire n2934;
	wire n2935;
	wire n2936;
	wire n2937;
	wire n2938;
	wire n2939;
	wire n2940;
	wire n2942;
	wire n2943;
	wire n2944;
	wire n2945;
	wire n2946;
	wire n2947;
	wire n2948;
	wire n2949;
	wire n2950;
	wire n2951;
	wire n2952;
	wire n2953;
	wire n2954;
	wire n2955;
	wire n2956;
	wire n2957;
	wire n2959;
	wire n2960;
	wire n2961;
	wire n2962;
	wire n2963;
	wire n2964;
	wire n2965;
	wire n2966;
	wire n2967;
	wire n2968;
	wire n2969;
	wire n2970;
	wire n2971;
	wire n2972;
	wire n2973;
	wire n2974;
	wire n2976;
	wire n2977;
	wire n2978;
	wire n2979;
	wire n2980;
	wire n2981;
	wire n2982;
	wire n2983;
	wire n2984;
	wire n2985;
	wire n2986;
	wire n2987;
	wire n2988;
	wire n2989;
	wire n2990;
	wire n2991;
	wire n2993;
	wire n2994;
	wire n2995;
	wire n2996;
	wire n2997;
	wire n2998;
	wire n2999;
	wire n3000;
	wire n3001;
	wire n3002;
	wire n3003;
	wire n3004;
	wire n3005;
	wire n3006;
	wire n3007;
	wire n3008;
	wire n3010;
	wire n3011;
	wire n3012;
	wire n3013;
	wire n3014;
	wire n3015;
	wire n3016;
	wire n3017;
	wire n3018;
	wire n3019;
	wire n3020;
	wire n3021;
	wire n3022;
	wire n3023;
	wire n3024;
	wire n3025;
	wire n3027;
	wire n3028;
	wire n3029;
	wire n3030;
	wire n3031;
	wire n3032;
	wire n3033;
	wire n3034;
	wire n3035;
	wire n3036;
	wire n3037;
	wire n3038;
	wire n3039;
	wire n3040;
	wire n3041;
	wire n3042;
	wire n3044;
	wire n3045;
	wire n3046;
	wire n3047;
	wire n3048;
	wire n3049;
	wire n3050;
	wire n3051;
	wire n3052;
	wire n3053;
	wire n3054;
	wire n3055;
	wire n3056;
	wire n3057;
	wire n3058;
	wire n3059;
	wire n3061;
	wire n3062;
	wire n3063;
	wire n3064;
	wire n3065;
	wire n3066;
	wire n3067;
	wire n3068;
	wire n3069;
	wire n3070;
	wire n3071;
	wire n3072;
	wire n3073;
	wire n3074;
	wire n3075;
	wire n3076;
	wire n3078;
	wire n3079;
	wire n3080;
	wire n3081;
	wire n3082;
	wire n3083;
	wire n3084;
	wire n3085;
	wire n3086;
	wire n3087;
	wire n3088;
	wire n3089;
	wire n3090;
	wire n3091;
	wire n3092;
	wire n3093;
	wire n3095;
	wire n3096;
	wire n3097;
	wire n3098;
	wire n3099;
	wire n3100;
	wire n3101;
	wire n3102;
	wire n3103;
	wire n3104;
	wire n3105;
	wire n3106;
	wire n3107;
	wire n3108;
	wire n3109;
	wire n3110;
	wire n3112;
	wire n3113;
	wire n3114;
	wire n3115;
	wire n3116;
	wire n3117;
	wire n3118;
	wire n3119;
	wire n3120;
	wire n3121;
	wire n3122;
	wire n3123;
	wire n3124;
	wire n3125;
	wire n3126;
	wire n3127;
	wire n3129;
	wire n3130;
	wire n3131;
	wire n3132;
	wire n3133;
	wire n3134;
	wire n3135;
	wire n3136;
	wire n3137;
	wire n3138;
	wire n3139;
	wire n3140;
	wire n3141;
	wire n3142;
	wire n3143;
	wire n3144;
	wire n3146;
	wire n3147;
	wire n3148;
	wire n3149;
	wire n3150;
	wire n3151;
	wire n3152;
	wire n3153;
	wire n3154;
	wire n3155;
	wire n3156;
	wire n3157;
	wire n3158;
	wire n3159;
	wire n3160;
	wire n3161;
	wire n3163;
	wire n3164;
	wire n3165;
	wire n3166;
	wire n3167;
	wire n3168;
	wire n3169;
	wire n3170;
	wire n3171;
	wire n3172;
	wire n3173;
	wire n3174;
	wire n3175;
	wire n3176;
	wire n3177;
	wire n3178;
	wire n3180;
	wire n3181;
	wire n3182;
	wire n3183;
	wire n3184;
	wire n3185;
	wire n3186;
	wire n3187;
	wire n3188;
	wire n3189;
	wire n3190;
	wire n3191;
	wire n3192;
	wire n3193;
	wire n3194;
	wire n3195;
	wire n3197;
	wire n3198;
	wire n3199;
	wire n3200;
	wire n3201;
	wire n3202;
	wire n3203;
	wire n3204;
	wire n3205;
	wire n3206;
	wire n3207;
	wire n3208;
	wire n3209;
	wire n3210;
	wire n3211;
	wire n3212;
	wire n3214;
	wire n3215;
	wire n3216;
	wire n3217;
	wire n3218;
	wire n3219;
	wire n3220;
	wire n3221;
	wire n3222;
	wire n3223;
	wire n3224;
	wire n3225;
	wire n3226;
	wire n3227;
	wire n3228;
	wire n3229;
	wire n3231;
	wire n3232;
	wire n3234;
	wire n3235;
	wire n3237;
	wire n3238;
	wire n3240;
	wire n3241;
	wire n3243;
	wire n3244;
	wire n3246;
	wire n3247;
	wire n3249;
	wire n3250;
	wire n3252;
	wire n3253;
	wire n3255;
	wire n3256;
	wire n3258;
	wire n3259;
	wire n3261;
	wire n3262;
	wire n3264;
	wire n3265;
	wire n3267;
	wire n3268;
	wire n3270;
	wire n3271;
	wire n3273;
	wire n3274;
	wire n3276;
	wire n3277;
	wire n3279;
	wire n3280;
	wire n3282;
	wire n3283;
	wire n3285;
	wire n3286;
	wire n3288;
	wire n3289;
	wire n3291;
	wire n3292;
	wire n3294;
	wire n3295;
	wire n3297;
	wire n3298;
	wire n3300;
	wire n3301;
	wire n3303;
	wire n3304;
	wire n3306;
	wire n3307;
	wire n3309;
	wire n3310;
	wire n3312;
	wire n3313;
	wire n3315;
	wire n3316;
	wire n3318;
	wire n3319;
	wire n3321;
	wire n3322;
	wire n3324;
	wire n3325;
	wire n3327;
	wire n3328;
	wire n3330;
	wire n3331;
	wire n3333;
	wire n3334;
	wire n3336;
	wire n3337;
	wire n3339;
	wire n3340;
	wire n3342;
	wire n3343;
	wire n3345;
	wire n3346;
	wire n3348;
	wire n3349;
	wire n3351;
	wire n3352;
	wire n3354;
	wire n3355;
	wire n3357;
	wire n3358;
	wire n3360;
	wire n3361;
	wire n3363;
	wire n3364;
	wire n3366;
	wire n3367;
	wire n3369;
	wire n3370;
	wire n3372;
	wire n3373;
	wire n3375;
	wire n3376;
	wire n3378;
	wire n3379;
	wire n3381;
	wire n3382;
	wire n3384;
	wire n3385;
	wire n3387;
	wire n3388;
	wire n3390;
	wire n3391;
	wire n3393;
	wire n3394;
	wire n3396;
	wire n3397;
	wire n3399;
	wire n3400;
	wire n3402;
	wire n3403;
	wire n3405;
	wire n3406;
	wire n3408;
	wire n3409;
	wire n3411;
	wire n3412;
	wire n3414;
	wire n3415;
	wire n3417;
	wire n3418;
	wire n3420;
	wire n3421;
	wire[1:0] w_a0_0;
	wire[1:0] w_a1_0;
	wire[1:0] w_a2_0;
	wire[1:0] w_a3_0;
	wire[1:0] w_a4_0;
	wire[1:0] w_a5_0;
	wire[1:0] w_a6_0;
	wire[1:0] w_a7_0;
	wire[1:0] w_a8_0;
	wire[1:0] w_a9_0;
	wire[1:0] w_a10_0;
	wire[1:0] w_a11_0;
	wire[1:0] w_a12_0;
	wire[1:0] w_a13_0;
	wire[1:0] w_a14_0;
	wire[1:0] w_a15_0;
	wire[1:0] w_a16_0;
	wire[1:0] w_a17_0;
	wire[1:0] w_a18_0;
	wire[1:0] w_a19_0;
	wire[1:0] w_a20_0;
	wire[1:0] w_a21_0;
	wire[1:0] w_a22_0;
	wire[1:0] w_a23_0;
	wire[1:0] w_a24_0;
	wire[1:0] w_a25_0;
	wire[1:0] w_a26_0;
	wire[1:0] w_a27_0;
	wire[1:0] w_a28_0;
	wire[1:0] w_a29_0;
	wire[1:0] w_a30_0;
	wire[1:0] w_a31_0;
	wire[1:0] w_a32_0;
	wire[1:0] w_a33_0;
	wire[1:0] w_a34_0;
	wire[1:0] w_a35_0;
	wire[1:0] w_a36_0;
	wire[1:0] w_a37_0;
	wire[1:0] w_a38_0;
	wire[1:0] w_a39_0;
	wire[1:0] w_a40_0;
	wire[1:0] w_a41_0;
	wire[1:0] w_a42_0;
	wire[1:0] w_a43_0;
	wire[1:0] w_a44_0;
	wire[1:0] w_a45_0;
	wire[1:0] w_a46_0;
	wire[1:0] w_a47_0;
	wire[1:0] w_a48_0;
	wire[1:0] w_a49_0;
	wire[1:0] w_a50_0;
	wire[1:0] w_a51_0;
	wire[1:0] w_a52_0;
	wire[1:0] w_a53_0;
	wire[1:0] w_a54_0;
	wire[1:0] w_a55_0;
	wire[1:0] w_a56_0;
	wire[1:0] w_a57_0;
	wire[1:0] w_a58_0;
	wire[1:0] w_a59_0;
	wire[1:0] w_a60_0;
	wire[1:0] w_a61_0;
	wire[1:0] w_a62_0;
	wire[1:0] w_a63_0;
	wire[1:0] w_a64_0;
	wire[1:0] w_a65_0;
	wire[1:0] w_a66_0;
	wire[1:0] w_a67_0;
	wire[1:0] w_a68_0;
	wire[1:0] w_a69_0;
	wire[1:0] w_a70_0;
	wire[1:0] w_a71_0;
	wire[1:0] w_a72_0;
	wire[1:0] w_a73_0;
	wire[1:0] w_a74_0;
	wire[1:0] w_a75_0;
	wire[1:0] w_a76_0;
	wire[1:0] w_a77_0;
	wire[1:0] w_a78_0;
	wire[1:0] w_a79_0;
	wire[1:0] w_a80_0;
	wire[1:0] w_a81_0;
	wire[1:0] w_a82_0;
	wire[1:0] w_a83_0;
	wire[1:0] w_a84_0;
	wire[1:0] w_a85_0;
	wire[1:0] w_a86_0;
	wire[1:0] w_a87_0;
	wire[1:0] w_a88_0;
	wire[1:0] w_a89_0;
	wire[1:0] w_a90_0;
	wire[1:0] w_a91_0;
	wire[1:0] w_a92_0;
	wire[1:0] w_a93_0;
	wire[1:0] w_a94_0;
	wire[1:0] w_a95_0;
	wire[1:0] w_a96_0;
	wire[1:0] w_a97_0;
	wire[1:0] w_a98_0;
	wire[1:0] w_a99_0;
	wire[1:0] w_a100_0;
	wire[1:0] w_a101_0;
	wire[1:0] w_a102_0;
	wire[1:0] w_a103_0;
	wire[1:0] w_a104_0;
	wire[1:0] w_a105_0;
	wire[1:0] w_a106_0;
	wire[1:0] w_a107_0;
	wire[1:0] w_a108_0;
	wire[1:0] w_a109_0;
	wire[1:0] w_a110_0;
	wire[1:0] w_a111_0;
	wire[1:0] w_a112_0;
	wire[1:0] w_a113_0;
	wire[1:0] w_a114_0;
	wire[1:0] w_a115_0;
	wire[1:0] w_a116_0;
	wire[1:0] w_a117_0;
	wire[1:0] w_a118_0;
	wire[1:0] w_a119_0;
	wire[1:0] w_a120_0;
	wire[1:0] w_a121_0;
	wire[1:0] w_a122_0;
	wire[1:0] w_a123_0;
	wire[1:0] w_a124_0;
	wire[1:0] w_a125_0;
	wire[1:0] w_a126_0;
	wire[1:0] w_a127_0;
	wire[2:0] w_shift0_0;
	wire[2:0] w_shift0_1;
	wire[2:0] w_shift0_2;
	wire[2:0] w_shift0_3;
	wire[2:0] w_shift0_4;
	wire[2:0] w_shift0_5;
	wire[2:0] w_shift0_6;
	wire[2:0] w_shift0_7;
	wire[2:0] w_shift0_8;
	wire[2:0] w_shift0_9;
	wire[2:0] w_shift0_10;
	wire[2:0] w_shift0_11;
	wire[2:0] w_shift0_12;
	wire[2:0] w_shift0_13;
	wire[2:0] w_shift0_14;
	wire[2:0] w_shift0_15;
	wire[2:0] w_shift0_16;
	wire[2:0] w_shift0_17;
	wire[2:0] w_shift0_18;
	wire[2:0] w_shift0_19;
	wire[2:0] w_shift0_20;
	wire[2:0] w_shift0_21;
	wire[2:0] w_shift0_22;
	wire[2:0] w_shift0_23;
	wire[2:0] w_shift0_24;
	wire[2:0] w_shift0_25;
	wire[2:0] w_shift0_26;
	wire[2:0] w_shift0_27;
	wire[2:0] w_shift0_28;
	wire[2:0] w_shift0_29;
	wire[2:0] w_shift0_30;
	wire[2:0] w_shift0_31;
	wire[2:0] w_shift0_32;
	wire[2:0] w_shift0_33;
	wire[2:0] w_shift0_34;
	wire[2:0] w_shift0_35;
	wire[2:0] w_shift0_36;
	wire[2:0] w_shift0_37;
	wire[2:0] w_shift0_38;
	wire[2:0] w_shift0_39;
	wire[2:0] w_shift0_40;
	wire[2:0] w_shift0_41;
	wire[2:0] w_shift0_42;
	wire[2:0] w_shift0_43;
	wire[2:0] w_shift0_44;
	wire[2:0] w_shift0_45;
	wire[2:0] w_shift0_46;
	wire[2:0] w_shift0_47;
	wire[2:0] w_shift0_48;
	wire[2:0] w_shift0_49;
	wire[2:0] w_shift0_50;
	wire[2:0] w_shift0_51;
	wire[2:0] w_shift0_52;
	wire[2:0] w_shift0_53;
	wire[2:0] w_shift0_54;
	wire[2:0] w_shift0_55;
	wire[2:0] w_shift0_56;
	wire[2:0] w_shift0_57;
	wire[2:0] w_shift0_58;
	wire[2:0] w_shift0_59;
	wire[2:0] w_shift0_60;
	wire[2:0] w_shift0_61;
	wire[2:0] w_shift0_62;
	wire[2:0] w_shift0_63;
	wire[2:0] w_shift1_0;
	wire[2:0] w_shift1_1;
	wire[2:0] w_shift1_2;
	wire[2:0] w_shift1_3;
	wire[2:0] w_shift1_4;
	wire[2:0] w_shift1_5;
	wire[2:0] w_shift1_6;
	wire[2:0] w_shift1_7;
	wire[2:0] w_shift1_8;
	wire[2:0] w_shift1_9;
	wire[2:0] w_shift1_10;
	wire[2:0] w_shift1_11;
	wire[2:0] w_shift1_12;
	wire[2:0] w_shift1_13;
	wire[2:0] w_shift1_14;
	wire[2:0] w_shift1_15;
	wire[2:0] w_shift1_16;
	wire[2:0] w_shift1_17;
	wire[2:0] w_shift1_18;
	wire[2:0] w_shift1_19;
	wire[2:0] w_shift1_20;
	wire[2:0] w_shift1_21;
	wire[2:0] w_shift1_22;
	wire[2:0] w_shift1_23;
	wire[2:0] w_shift1_24;
	wire[2:0] w_shift1_25;
	wire[2:0] w_shift1_26;
	wire[2:0] w_shift1_27;
	wire[2:0] w_shift1_28;
	wire[2:0] w_shift1_29;
	wire[2:0] w_shift1_30;
	wire[2:0] w_shift1_31;
	wire[2:0] w_shift1_32;
	wire[2:0] w_shift1_33;
	wire[2:0] w_shift1_34;
	wire[2:0] w_shift1_35;
	wire[2:0] w_shift1_36;
	wire[2:0] w_shift1_37;
	wire[2:0] w_shift1_38;
	wire[2:0] w_shift1_39;
	wire[2:0] w_shift1_40;
	wire[2:0] w_shift1_41;
	wire[2:0] w_shift1_42;
	wire[2:0] w_shift1_43;
	wire[2:0] w_shift1_44;
	wire[2:0] w_shift1_45;
	wire[2:0] w_shift1_46;
	wire[2:0] w_shift1_47;
	wire[2:0] w_shift1_48;
	wire[2:0] w_shift1_49;
	wire[2:0] w_shift1_50;
	wire[2:0] w_shift1_51;
	wire[2:0] w_shift1_52;
	wire[2:0] w_shift1_53;
	wire[2:0] w_shift1_54;
	wire[2:0] w_shift1_55;
	wire[2:0] w_shift1_56;
	wire[2:0] w_shift1_57;
	wire[2:0] w_shift1_58;
	wire[2:0] w_shift1_59;
	wire[2:0] w_shift1_60;
	wire[2:0] w_shift1_61;
	wire[2:0] w_shift1_62;
	wire[2:0] w_shift1_63;
	wire[2:0] w_shift1_64;
	wire[2:0] w_shift1_65;
	wire[2:0] w_shift1_66;
	wire[2:0] w_shift1_67;
	wire[2:0] w_shift1_68;
	wire[2:0] w_shift1_69;
	wire[2:0] w_shift1_70;
	wire[2:0] w_shift1_71;
	wire[2:0] w_shift1_72;
	wire[2:0] w_shift1_73;
	wire[2:0] w_shift1_74;
	wire[2:0] w_shift1_75;
	wire[2:0] w_shift1_76;
	wire[2:0] w_shift1_77;
	wire[2:0] w_shift1_78;
	wire[2:0] w_shift1_79;
	wire[2:0] w_shift1_80;
	wire[2:0] w_shift1_81;
	wire[2:0] w_shift1_82;
	wire[2:0] w_shift1_83;
	wire[2:0] w_shift1_84;
	wire[2:0] w_shift1_85;
	wire[2:0] w_shift1_86;
	wire[2:0] w_shift1_87;
	wire[2:0] w_shift1_88;
	wire[2:0] w_shift1_89;
	wire[2:0] w_shift1_90;
	wire[2:0] w_shift1_91;
	wire[2:0] w_shift1_92;
	wire[2:0] w_shift1_93;
	wire[2:0] w_shift1_94;
	wire[2:0] w_shift1_95;
	wire[2:0] w_shift1_96;
	wire[2:0] w_shift2_0;
	wire[2:0] w_shift3_0;
	wire[2:0] w_shift4_0;
	wire[2:0] w_shift5_0;
	wire[2:0] w_shift6_0;
	wire[2:0] w_shift6_1;
	wire[2:0] w_shift6_2;
	wire[2:0] w_shift6_3;
	wire[2:0] w_shift6_4;
	wire[2:0] w_shift6_5;
	wire[2:0] w_shift6_6;
	wire[2:0] w_shift6_7;
	wire[2:0] w_shift6_8;
	wire[2:0] w_shift6_9;
	wire[2:0] w_shift6_10;
	wire[2:0] w_shift6_11;
	wire[2:0] w_shift6_12;
	wire[2:0] w_shift6_13;
	wire[2:0] w_shift6_14;
	wire[2:0] w_shift6_15;
	wire[2:0] w_shift6_16;
	wire[2:0] w_shift6_17;
	wire[2:0] w_shift6_18;
	wire[2:0] w_shift6_19;
	wire[2:0] w_shift6_20;
	wire[2:0] w_shift6_21;
	wire[2:0] w_shift6_22;
	wire[2:0] w_shift6_23;
	wire[2:0] w_shift6_24;
	wire[2:0] w_shift6_25;
	wire[2:0] w_shift6_26;
	wire[2:0] w_shift6_27;
	wire[2:0] w_shift6_28;
	wire[2:0] w_shift6_29;
	wire[2:0] w_shift6_30;
	wire[2:0] w_shift6_31;
	wire[2:0] w_shift6_32;
	wire[2:0] w_shift6_33;
	wire[2:0] w_shift6_34;
	wire[2:0] w_shift6_35;
	wire[2:0] w_shift6_36;
	wire[2:0] w_shift6_37;
	wire[2:0] w_shift6_38;
	wire[2:0] w_shift6_39;
	wire[2:0] w_shift6_40;
	wire[2:0] w_shift6_41;
	wire[2:0] w_shift6_42;
	wire[2:0] w_shift6_43;
	wire[2:0] w_shift6_44;
	wire[2:0] w_shift6_45;
	wire[2:0] w_shift6_46;
	wire[2:0] w_shift6_47;
	wire[2:0] w_shift6_48;
	wire[2:0] w_shift6_49;
	wire[2:0] w_shift6_50;
	wire[2:0] w_shift6_51;
	wire[2:0] w_shift6_52;
	wire[2:0] w_shift6_53;
	wire[2:0] w_shift6_54;
	wire[2:0] w_shift6_55;
	wire[2:0] w_shift6_56;
	wire[2:0] w_shift6_57;
	wire[2:0] w_shift6_58;
	wire[2:0] w_shift6_59;
	wire[2:0] w_shift6_60;
	wire[2:0] w_shift6_61;
	wire[2:0] w_shift6_62;
	wire[2:0] w_shift6_63;
	wire[2:0] w_n263_0;
	wire[2:0] w_n263_1;
	wire[2:0] w_n263_2;
	wire[2:0] w_n263_3;
	wire[2:0] w_n263_4;
	wire[2:0] w_n263_5;
	wire[2:0] w_n263_6;
	wire[2:0] w_n263_7;
	wire[2:0] w_n263_8;
	wire[2:0] w_n263_9;
	wire[2:0] w_n263_10;
	wire[2:0] w_n263_11;
	wire[2:0] w_n263_12;
	wire[2:0] w_n263_13;
	wire[2:0] w_n263_14;
	wire[2:0] w_n263_15;
	wire[2:0] w_n263_16;
	wire[2:0] w_n263_17;
	wire[2:0] w_n263_18;
	wire[2:0] w_n263_19;
	wire[2:0] w_n263_20;
	wire[2:0] w_n263_21;
	wire[2:0] w_n263_22;
	wire[2:0] w_n263_23;
	wire[2:0] w_n263_24;
	wire[2:0] w_n263_25;
	wire[2:0] w_n263_26;
	wire[2:0] w_n263_27;
	wire[2:0] w_n263_28;
	wire[2:0] w_n263_29;
	wire[2:0] w_n263_30;
	wire[2:0] w_n263_31;
	wire[2:0] w_n263_32;
	wire[2:0] w_n263_33;
	wire[2:0] w_n263_34;
	wire[2:0] w_n263_35;
	wire[2:0] w_n263_36;
	wire[2:0] w_n263_37;
	wire[2:0] w_n263_38;
	wire[2:0] w_n263_39;
	wire[2:0] w_n263_40;
	wire[2:0] w_n263_41;
	wire[2:0] w_n263_42;
	wire[2:0] w_n263_43;
	wire[2:0] w_n263_44;
	wire[2:0] w_n263_45;
	wire[2:0] w_n263_46;
	wire[2:0] w_n263_47;
	wire[2:0] w_n263_48;
	wire[2:0] w_n263_49;
	wire[2:0] w_n263_50;
	wire[2:0] w_n263_51;
	wire[2:0] w_n263_52;
	wire[2:0] w_n263_53;
	wire[2:0] w_n263_54;
	wire[2:0] w_n263_55;
	wire[2:0] w_n263_56;
	wire[2:0] w_n263_57;
	wire[2:0] w_n263_58;
	wire[2:0] w_n263_59;
	wire[2:0] w_n263_60;
	wire[2:0] w_n263_61;
	wire[2:0] w_n263_62;
	wire[1:0] w_n263_63;
	wire[1:0] w_n264_0;
	wire[1:0] w_n265_0;
	wire[2:0] w_n266_0;
	wire[2:0] w_n266_1;
	wire[2:0] w_n266_2;
	wire[2:0] w_n266_3;
	wire[2:0] w_n266_4;
	wire[2:0] w_n266_5;
	wire[2:0] w_n266_6;
	wire[2:0] w_n266_7;
	wire[2:0] w_n266_8;
	wire[2:0] w_n266_9;
	wire[2:0] w_n266_10;
	wire[2:0] w_n266_11;
	wire[2:0] w_n266_12;
	wire[2:0] w_n266_13;
	wire[2:0] w_n266_14;
	wire[2:0] w_n266_15;
	wire[2:0] w_n266_16;
	wire[2:0] w_n266_17;
	wire[2:0] w_n266_18;
	wire[2:0] w_n266_19;
	wire[2:0] w_n266_20;
	wire[2:0] w_n266_21;
	wire[2:0] w_n266_22;
	wire[2:0] w_n266_23;
	wire[2:0] w_n266_24;
	wire[2:0] w_n266_25;
	wire[2:0] w_n266_26;
	wire[2:0] w_n266_27;
	wire[2:0] w_n266_28;
	wire[2:0] w_n266_29;
	wire[2:0] w_n266_30;
	wire[2:0] w_n266_31;
	wire[2:0] w_n266_32;
	wire[2:0] w_n266_33;
	wire[2:0] w_n266_34;
	wire[2:0] w_n266_35;
	wire[2:0] w_n266_36;
	wire[2:0] w_n266_37;
	wire[2:0] w_n266_38;
	wire[2:0] w_n266_39;
	wire[2:0] w_n266_40;
	wire[2:0] w_n266_41;
	wire[2:0] w_n266_42;
	wire[2:0] w_n266_43;
	wire[2:0] w_n266_44;
	wire[2:0] w_n266_45;
	wire[2:0] w_n266_46;
	wire[2:0] w_n266_47;
	wire[2:0] w_n266_48;
	wire[2:0] w_n266_49;
	wire[2:0] w_n266_50;
	wire[2:0] w_n266_51;
	wire[2:0] w_n266_52;
	wire[2:0] w_n266_53;
	wire[2:0] w_n266_54;
	wire[2:0] w_n266_55;
	wire[2:0] w_n266_56;
	wire[2:0] w_n266_57;
	wire[2:0] w_n266_58;
	wire[2:0] w_n266_59;
	wire[2:0] w_n266_60;
	wire[2:0] w_n266_61;
	wire[2:0] w_n266_62;
	wire[1:0] w_n266_63;
	wire[1:0] w_n267_0;
	wire[2:0] w_n269_0;
	wire[2:0] w_n269_1;
	wire[2:0] w_n269_2;
	wire[2:0] w_n269_3;
	wire[2:0] w_n269_4;
	wire[2:0] w_n269_5;
	wire[2:0] w_n269_6;
	wire[2:0] w_n269_7;
	wire[2:0] w_n269_8;
	wire[2:0] w_n269_9;
	wire[2:0] w_n269_10;
	wire[2:0] w_n269_11;
	wire[2:0] w_n269_12;
	wire[2:0] w_n269_13;
	wire[2:0] w_n269_14;
	wire[2:0] w_n269_15;
	wire[2:0] w_n269_16;
	wire[2:0] w_n269_17;
	wire[2:0] w_n269_18;
	wire[2:0] w_n269_19;
	wire[2:0] w_n269_20;
	wire[2:0] w_n269_21;
	wire[2:0] w_n269_22;
	wire[2:0] w_n269_23;
	wire[2:0] w_n269_24;
	wire[2:0] w_n269_25;
	wire[2:0] w_n269_26;
	wire[2:0] w_n269_27;
	wire[2:0] w_n269_28;
	wire[2:0] w_n269_29;
	wire[2:0] w_n269_30;
	wire[2:0] w_n269_31;
	wire[2:0] w_n269_32;
	wire[2:0] w_n269_33;
	wire[2:0] w_n269_34;
	wire[2:0] w_n269_35;
	wire[2:0] w_n269_36;
	wire[2:0] w_n269_37;
	wire[2:0] w_n269_38;
	wire[2:0] w_n269_39;
	wire[2:0] w_n269_40;
	wire[2:0] w_n269_41;
	wire[2:0] w_n269_42;
	wire[2:0] w_n269_43;
	wire[2:0] w_n269_44;
	wire[2:0] w_n269_45;
	wire[2:0] w_n269_46;
	wire[2:0] w_n269_47;
	wire[2:0] w_n269_48;
	wire[2:0] w_n269_49;
	wire[2:0] w_n269_50;
	wire[2:0] w_n269_51;
	wire[2:0] w_n269_52;
	wire[2:0] w_n269_53;
	wire[2:0] w_n269_54;
	wire[2:0] w_n269_55;
	wire[2:0] w_n269_56;
	wire[2:0] w_n269_57;
	wire[2:0] w_n269_58;
	wire[2:0] w_n269_59;
	wire[2:0] w_n269_60;
	wire[2:0] w_n269_61;
	wire[2:0] w_n269_62;
	wire[2:0] w_n269_63;
	wire[2:0] w_n269_64;
	wire[2:0] w_n269_65;
	wire[2:0] w_n269_66;
	wire[2:0] w_n269_67;
	wire[2:0] w_n269_68;
	wire[2:0] w_n269_69;
	wire[2:0] w_n269_70;
	wire[2:0] w_n269_71;
	wire[2:0] w_n269_72;
	wire[2:0] w_n269_73;
	wire[2:0] w_n269_74;
	wire[2:0] w_n269_75;
	wire[2:0] w_n269_76;
	wire[2:0] w_n269_77;
	wire[2:0] w_n269_78;
	wire[2:0] w_n269_79;
	wire[2:0] w_n269_80;
	wire[2:0] w_n269_81;
	wire[2:0] w_n269_82;
	wire[2:0] w_n269_83;
	wire[2:0] w_n269_84;
	wire[2:0] w_n269_85;
	wire[2:0] w_n269_86;
	wire[2:0] w_n269_87;
	wire[2:0] w_n269_88;
	wire[2:0] w_n269_89;
	wire[2:0] w_n269_90;
	wire[2:0] w_n269_91;
	wire[2:0] w_n269_92;
	wire[2:0] w_n269_93;
	wire[2:0] w_n269_94;
	wire[2:0] w_n269_95;
	wire[1:0] w_n269_96;
	wire[2:0] w_n270_0;
	wire[2:0] w_n270_1;
	wire[2:0] w_n270_2;
	wire[2:0] w_n270_3;
	wire[2:0] w_n270_4;
	wire[2:0] w_n270_5;
	wire[2:0] w_n270_6;
	wire[2:0] w_n270_7;
	wire[2:0] w_n270_8;
	wire[2:0] w_n270_9;
	wire[2:0] w_n270_10;
	wire[2:0] w_n270_11;
	wire[2:0] w_n270_12;
	wire[2:0] w_n270_13;
	wire[2:0] w_n270_14;
	wire[2:0] w_n270_15;
	wire[2:0] w_n270_16;
	wire[2:0] w_n270_17;
	wire[2:0] w_n270_18;
	wire[2:0] w_n270_19;
	wire[2:0] w_n270_20;
	wire[2:0] w_n270_21;
	wire[2:0] w_n270_22;
	wire[2:0] w_n270_23;
	wire[2:0] w_n270_24;
	wire[2:0] w_n270_25;
	wire[2:0] w_n270_26;
	wire[2:0] w_n270_27;
	wire[2:0] w_n270_28;
	wire[2:0] w_n270_29;
	wire[2:0] w_n270_30;
	wire[2:0] w_n270_31;
	wire[2:0] w_n270_32;
	wire[2:0] w_n270_33;
	wire[2:0] w_n270_34;
	wire[2:0] w_n270_35;
	wire[2:0] w_n270_36;
	wire[2:0] w_n270_37;
	wire[2:0] w_n270_38;
	wire[2:0] w_n270_39;
	wire[2:0] w_n270_40;
	wire[2:0] w_n270_41;
	wire[2:0] w_n270_42;
	wire[2:0] w_n270_43;
	wire[2:0] w_n270_44;
	wire[2:0] w_n270_45;
	wire[2:0] w_n270_46;
	wire[2:0] w_n270_47;
	wire[2:0] w_n270_48;
	wire[2:0] w_n270_49;
	wire[2:0] w_n270_50;
	wire[2:0] w_n270_51;
	wire[2:0] w_n270_52;
	wire[2:0] w_n270_53;
	wire[2:0] w_n270_54;
	wire[2:0] w_n270_55;
	wire[2:0] w_n270_56;
	wire[2:0] w_n270_57;
	wire[2:0] w_n270_58;
	wire[2:0] w_n270_59;
	wire[2:0] w_n270_60;
	wire[2:0] w_n270_61;
	wire[2:0] w_n270_62;
	wire[1:0] w_n270_63;
	wire[1:0] w_n271_0;
	wire[1:0] w_n274_0;
	wire[1:0] w_n276_0;
	wire[2:0] w_n279_0;
	wire[1:0] w_n279_1;
	wire[2:0] w_n281_0;
	wire[2:0] w_n281_1;
	wire[2:0] w_n281_2;
	wire[2:0] w_n281_3;
	wire[2:0] w_n281_4;
	wire[2:0] w_n281_5;
	wire[2:0] w_n281_6;
	wire[2:0] w_n281_7;
	wire[2:0] w_n281_8;
	wire[2:0] w_n281_9;
	wire[2:0] w_n281_10;
	wire[2:0] w_n281_11;
	wire[2:0] w_n281_12;
	wire[2:0] w_n281_13;
	wire[2:0] w_n281_14;
	wire[2:0] w_n281_15;
	wire[2:0] w_n281_16;
	wire[2:0] w_n281_17;
	wire[2:0] w_n281_18;
	wire[2:0] w_n281_19;
	wire[2:0] w_n281_20;
	wire[2:0] w_n281_21;
	wire[2:0] w_n281_22;
	wire[2:0] w_n281_23;
	wire[2:0] w_n281_24;
	wire[2:0] w_n281_25;
	wire[2:0] w_n281_26;
	wire[2:0] w_n281_27;
	wire[2:0] w_n281_28;
	wire[2:0] w_n281_29;
	wire[2:0] w_n281_30;
	wire[2:0] w_n281_31;
	wire[2:0] w_n281_32;
	wire[2:0] w_n281_33;
	wire[2:0] w_n281_34;
	wire[2:0] w_n281_35;
	wire[2:0] w_n281_36;
	wire[2:0] w_n281_37;
	wire[2:0] w_n281_38;
	wire[2:0] w_n281_39;
	wire[2:0] w_n281_40;
	wire[2:0] w_n281_41;
	wire[2:0] w_n281_42;
	wire[2:0] w_n281_43;
	wire[2:0] w_n281_44;
	wire[2:0] w_n281_45;
	wire[2:0] w_n281_46;
	wire[2:0] w_n281_47;
	wire[2:0] w_n281_48;
	wire[2:0] w_n281_49;
	wire[2:0] w_n281_50;
	wire[2:0] w_n281_51;
	wire[2:0] w_n281_52;
	wire[2:0] w_n281_53;
	wire[2:0] w_n281_54;
	wire[2:0] w_n281_55;
	wire[2:0] w_n281_56;
	wire[2:0] w_n281_57;
	wire[2:0] w_n281_58;
	wire[2:0] w_n281_59;
	wire[2:0] w_n281_60;
	wire[2:0] w_n281_61;
	wire[2:0] w_n281_62;
	wire[1:0] w_n281_63;
	wire[1:0] w_n282_0;
	wire[1:0] w_n284_0;
	wire[1:0] w_n287_0;
	wire[1:0] w_n289_0;
	wire[2:0] w_n292_0;
	wire[1:0] w_n292_1;
	wire[2:0] w_n295_0;
	wire[2:0] w_n295_1;
	wire[2:0] w_n295_2;
	wire[2:0] w_n295_3;
	wire[2:0] w_n295_4;
	wire[2:0] w_n295_5;
	wire[2:0] w_n295_6;
	wire[2:0] w_n295_7;
	wire[2:0] w_n295_8;
	wire[2:0] w_n295_9;
	wire[2:0] w_n295_10;
	wire[2:0] w_n295_11;
	wire[2:0] w_n295_12;
	wire[2:0] w_n295_13;
	wire[2:0] w_n295_14;
	wire[2:0] w_n295_15;
	wire[2:0] w_n295_16;
	wire[2:0] w_n295_17;
	wire[2:0] w_n295_18;
	wire[2:0] w_n295_19;
	wire[2:0] w_n295_20;
	wire[2:0] w_n295_21;
	wire[2:0] w_n295_22;
	wire[2:0] w_n295_23;
	wire[2:0] w_n295_24;
	wire[2:0] w_n295_25;
	wire[2:0] w_n295_26;
	wire[2:0] w_n295_27;
	wire[2:0] w_n295_28;
	wire[2:0] w_n295_29;
	wire[2:0] w_n295_30;
	wire[2:0] w_n295_31;
	wire[2:0] w_n295_32;
	wire[2:0] w_n295_33;
	wire[2:0] w_n295_34;
	wire[2:0] w_n295_35;
	wire[2:0] w_n295_36;
	wire[2:0] w_n295_37;
	wire[2:0] w_n295_38;
	wire[2:0] w_n295_39;
	wire[2:0] w_n295_40;
	wire[2:0] w_n295_41;
	wire[2:0] w_n295_42;
	wire[2:0] w_n295_43;
	wire[2:0] w_n295_44;
	wire[2:0] w_n295_45;
	wire[2:0] w_n295_46;
	wire[2:0] w_n295_47;
	wire[2:0] w_n295_48;
	wire[2:0] w_n295_49;
	wire[2:0] w_n295_50;
	wire[2:0] w_n295_51;
	wire[2:0] w_n295_52;
	wire[2:0] w_n295_53;
	wire[2:0] w_n295_54;
	wire[2:0] w_n295_55;
	wire[2:0] w_n295_56;
	wire[2:0] w_n295_57;
	wire[2:0] w_n295_58;
	wire[2:0] w_n295_59;
	wire[2:0] w_n295_60;
	wire[2:0] w_n295_61;
	wire[2:0] w_n295_62;
	wire[1:0] w_n295_63;
	wire[1:0] w_n296_0;
	wire[1:0] w_n298_0;
	wire[1:0] w_n301_0;
	wire[1:0] w_n303_0;
	wire[2:0] w_n306_0;
	wire[1:0] w_n306_1;
	wire[2:0] w_n308_0;
	wire[2:0] w_n308_1;
	wire[2:0] w_n308_2;
	wire[2:0] w_n308_3;
	wire[2:0] w_n308_4;
	wire[2:0] w_n308_5;
	wire[2:0] w_n308_6;
	wire[2:0] w_n308_7;
	wire[2:0] w_n308_8;
	wire[2:0] w_n308_9;
	wire[2:0] w_n308_10;
	wire[2:0] w_n308_11;
	wire[2:0] w_n308_12;
	wire[2:0] w_n308_13;
	wire[2:0] w_n308_14;
	wire[2:0] w_n308_15;
	wire[2:0] w_n308_16;
	wire[2:0] w_n308_17;
	wire[2:0] w_n308_18;
	wire[2:0] w_n308_19;
	wire[2:0] w_n308_20;
	wire[2:0] w_n308_21;
	wire[2:0] w_n308_22;
	wire[2:0] w_n308_23;
	wire[2:0] w_n308_24;
	wire[2:0] w_n308_25;
	wire[2:0] w_n308_26;
	wire[2:0] w_n308_27;
	wire[2:0] w_n308_28;
	wire[2:0] w_n308_29;
	wire[2:0] w_n308_30;
	wire[2:0] w_n308_31;
	wire[2:0] w_n308_32;
	wire[2:0] w_n308_33;
	wire[2:0] w_n308_34;
	wire[2:0] w_n308_35;
	wire[2:0] w_n308_36;
	wire[2:0] w_n308_37;
	wire[2:0] w_n308_38;
	wire[2:0] w_n308_39;
	wire[2:0] w_n308_40;
	wire[2:0] w_n308_41;
	wire[2:0] w_n308_42;
	wire[2:0] w_n308_43;
	wire[2:0] w_n308_44;
	wire[2:0] w_n308_45;
	wire[2:0] w_n308_46;
	wire[2:0] w_n308_47;
	wire[2:0] w_n308_48;
	wire[2:0] w_n308_49;
	wire[2:0] w_n308_50;
	wire[2:0] w_n308_51;
	wire[2:0] w_n308_52;
	wire[2:0] w_n308_53;
	wire[2:0] w_n308_54;
	wire[2:0] w_n308_55;
	wire[2:0] w_n308_56;
	wire[2:0] w_n308_57;
	wire[2:0] w_n308_58;
	wire[2:0] w_n308_59;
	wire[2:0] w_n308_60;
	wire[2:0] w_n308_61;
	wire[2:0] w_n308_62;
	wire[1:0] w_n308_63;
	wire[1:0] w_n309_0;
	wire[1:0] w_n311_0;
	wire[1:0] w_n314_0;
	wire[1:0] w_n316_0;
	wire[2:0] w_n319_0;
	wire[1:0] w_n319_1;
	wire[2:0] w_n322_0;
	wire[1:0] w_n322_1;
	wire[2:0] w_n323_0;
	wire[2:0] w_n323_1;
	wire[2:0] w_n323_2;
	wire[2:0] w_n323_3;
	wire[2:0] w_n323_4;
	wire[2:0] w_n323_5;
	wire[2:0] w_n323_6;
	wire[2:0] w_n323_7;
	wire[2:0] w_n323_8;
	wire[2:0] w_n323_9;
	wire[2:0] w_n323_10;
	wire[2:0] w_n323_11;
	wire[2:0] w_n323_12;
	wire[2:0] w_n323_13;
	wire[2:0] w_n323_14;
	wire[2:0] w_n323_15;
	wire[2:0] w_n323_16;
	wire[2:0] w_n323_17;
	wire[2:0] w_n323_18;
	wire[2:0] w_n323_19;
	wire[2:0] w_n323_20;
	wire[2:0] w_n323_21;
	wire[2:0] w_n323_22;
	wire[2:0] w_n323_23;
	wire[2:0] w_n323_24;
	wire[2:0] w_n323_25;
	wire[2:0] w_n323_26;
	wire[2:0] w_n323_27;
	wire[2:0] w_n323_28;
	wire[2:0] w_n323_29;
	wire[2:0] w_n323_30;
	wire[2:0] w_n323_31;
	wire[2:0] w_n323_32;
	wire[2:0] w_n323_33;
	wire[2:0] w_n323_34;
	wire[2:0] w_n323_35;
	wire[2:0] w_n323_36;
	wire[2:0] w_n323_37;
	wire[2:0] w_n323_38;
	wire[2:0] w_n323_39;
	wire[2:0] w_n323_40;
	wire[2:0] w_n323_41;
	wire[2:0] w_n323_42;
	wire[2:0] w_n323_43;
	wire[2:0] w_n323_44;
	wire[2:0] w_n323_45;
	wire[2:0] w_n323_46;
	wire[2:0] w_n323_47;
	wire[2:0] w_n323_48;
	wire[2:0] w_n323_49;
	wire[2:0] w_n323_50;
	wire[2:0] w_n323_51;
	wire[2:0] w_n323_52;
	wire[2:0] w_n323_53;
	wire[2:0] w_n323_54;
	wire[2:0] w_n323_55;
	wire[2:0] w_n323_56;
	wire[2:0] w_n323_57;
	wire[2:0] w_n323_58;
	wire[2:0] w_n323_59;
	wire[2:0] w_n323_60;
	wire[2:0] w_n323_61;
	wire[2:0] w_n323_62;
	wire[1:0] w_n323_63;
	wire[1:0] w_n325_0;
	wire[1:0] w_n327_0;
	wire[1:0] w_n330_0;
	wire[1:0] w_n332_0;
	wire[2:0] w_n335_0;
	wire[1:0] w_n335_1;
	wire[1:0] w_n337_0;
	wire[1:0] w_n339_0;
	wire[1:0] w_n342_0;
	wire[1:0] w_n344_0;
	wire[2:0] w_n347_0;
	wire[1:0] w_n347_1;
	wire[1:0] w_n350_0;
	wire[1:0] w_n352_0;
	wire[1:0] w_n355_0;
	wire[1:0] w_n357_0;
	wire[2:0] w_n360_0;
	wire[1:0] w_n360_1;
	wire[1:0] w_n362_0;
	wire[1:0] w_n364_0;
	wire[1:0] w_n367_0;
	wire[1:0] w_n369_0;
	wire[2:0] w_n372_0;
	wire[1:0] w_n372_1;
	wire[2:0] w_n375_0;
	wire[1:0] w_n375_1;
	wire[1:0] w_n376_0;
	wire[2:0] w_n377_0;
	wire[2:0] w_n377_1;
	wire[2:0] w_n377_2;
	wire[2:0] w_n377_3;
	wire[2:0] w_n377_4;
	wire[2:0] w_n377_5;
	wire[2:0] w_n377_6;
	wire[2:0] w_n377_7;
	wire[2:0] w_n377_8;
	wire[2:0] w_n377_9;
	wire[2:0] w_n377_10;
	wire[2:0] w_n377_11;
	wire[2:0] w_n377_12;
	wire[2:0] w_n377_13;
	wire[2:0] w_n377_14;
	wire[2:0] w_n377_15;
	wire[2:0] w_n377_16;
	wire[2:0] w_n377_17;
	wire[2:0] w_n377_18;
	wire[2:0] w_n377_19;
	wire[2:0] w_n377_20;
	wire[2:0] w_n377_21;
	wire[2:0] w_n377_22;
	wire[2:0] w_n377_23;
	wire[2:0] w_n377_24;
	wire[2:0] w_n377_25;
	wire[2:0] w_n377_26;
	wire[2:0] w_n377_27;
	wire[2:0] w_n377_28;
	wire[2:0] w_n377_29;
	wire[2:0] w_n377_30;
	wire[2:0] w_n377_31;
	wire[2:0] w_n377_32;
	wire[2:0] w_n377_33;
	wire[2:0] w_n377_34;
	wire[2:0] w_n377_35;
	wire[2:0] w_n377_36;
	wire[2:0] w_n377_37;
	wire[2:0] w_n377_38;
	wire[2:0] w_n377_39;
	wire[2:0] w_n377_40;
	wire[2:0] w_n377_41;
	wire[2:0] w_n377_42;
	wire[2:0] w_n377_43;
	wire[2:0] w_n377_44;
	wire[2:0] w_n377_45;
	wire[2:0] w_n377_46;
	wire[2:0] w_n377_47;
	wire[2:0] w_n377_48;
	wire[2:0] w_n377_49;
	wire[2:0] w_n377_50;
	wire[2:0] w_n377_51;
	wire[2:0] w_n377_52;
	wire[2:0] w_n377_53;
	wire[2:0] w_n377_54;
	wire[2:0] w_n377_55;
	wire[2:0] w_n377_56;
	wire[2:0] w_n377_57;
	wire[2:0] w_n377_58;
	wire[2:0] w_n377_59;
	wire[2:0] w_n377_60;
	wire[2:0] w_n377_61;
	wire[2:0] w_n377_62;
	wire[1:0] w_n377_63;
	wire[1:0] w_n380_0;
	wire[1:0] w_n382_0;
	wire[1:0] w_n385_0;
	wire[1:0] w_n387_0;
	wire[2:0] w_n390_0;
	wire[1:0] w_n390_1;
	wire[1:0] w_n392_0;
	wire[1:0] w_n394_0;
	wire[1:0] w_n397_0;
	wire[1:0] w_n399_0;
	wire[2:0] w_n402_0;
	wire[1:0] w_n402_1;
	wire[1:0] w_n405_0;
	wire[1:0] w_n407_0;
	wire[1:0] w_n410_0;
	wire[1:0] w_n412_0;
	wire[2:0] w_n415_0;
	wire[1:0] w_n415_1;
	wire[1:0] w_n417_0;
	wire[1:0] w_n419_0;
	wire[1:0] w_n422_0;
	wire[1:0] w_n424_0;
	wire[2:0] w_n427_0;
	wire[1:0] w_n427_1;
	wire[2:0] w_n430_0;
	wire[1:0] w_n430_1;
	wire[1:0] w_n431_0;
	wire[2:0] w_n432_0;
	wire[2:0] w_n432_1;
	wire[2:0] w_n432_2;
	wire[2:0] w_n432_3;
	wire[2:0] w_n432_4;
	wire[2:0] w_n432_5;
	wire[2:0] w_n432_6;
	wire[2:0] w_n432_7;
	wire[2:0] w_n432_8;
	wire[2:0] w_n432_9;
	wire[2:0] w_n432_10;
	wire[2:0] w_n432_11;
	wire[2:0] w_n432_12;
	wire[2:0] w_n432_13;
	wire[2:0] w_n432_14;
	wire[2:0] w_n432_15;
	wire[2:0] w_n432_16;
	wire[2:0] w_n432_17;
	wire[2:0] w_n432_18;
	wire[2:0] w_n432_19;
	wire[2:0] w_n432_20;
	wire[2:0] w_n432_21;
	wire[2:0] w_n432_22;
	wire[2:0] w_n432_23;
	wire[2:0] w_n432_24;
	wire[2:0] w_n432_25;
	wire[2:0] w_n432_26;
	wire[2:0] w_n432_27;
	wire[2:0] w_n432_28;
	wire[2:0] w_n432_29;
	wire[2:0] w_n432_30;
	wire[2:0] w_n432_31;
	wire[2:0] w_n432_32;
	wire[2:0] w_n432_33;
	wire[2:0] w_n432_34;
	wire[2:0] w_n432_35;
	wire[2:0] w_n432_36;
	wire[2:0] w_n432_37;
	wire[2:0] w_n432_38;
	wire[2:0] w_n432_39;
	wire[2:0] w_n432_40;
	wire[2:0] w_n432_41;
	wire[2:0] w_n432_42;
	wire[2:0] w_n432_43;
	wire[2:0] w_n432_44;
	wire[2:0] w_n432_45;
	wire[2:0] w_n432_46;
	wire[2:0] w_n432_47;
	wire[2:0] w_n432_48;
	wire[2:0] w_n432_49;
	wire[2:0] w_n432_50;
	wire[2:0] w_n432_51;
	wire[2:0] w_n432_52;
	wire[2:0] w_n432_53;
	wire[2:0] w_n432_54;
	wire[2:0] w_n432_55;
	wire[2:0] w_n432_56;
	wire[2:0] w_n432_57;
	wire[2:0] w_n432_58;
	wire[2:0] w_n432_59;
	wire[2:0] w_n432_60;
	wire[2:0] w_n432_61;
	wire[2:0] w_n432_62;
	wire[1:0] w_n432_63;
	wire[1:0] w_n434_0;
	wire[1:0] w_n436_0;
	wire[1:0] w_n439_0;
	wire[1:0] w_n441_0;
	wire[2:0] w_n444_0;
	wire[1:0] w_n444_1;
	wire[1:0] w_n446_0;
	wire[1:0] w_n448_0;
	wire[1:0] w_n451_0;
	wire[1:0] w_n453_0;
	wire[2:0] w_n456_0;
	wire[1:0] w_n456_1;
	wire[1:0] w_n459_0;
	wire[1:0] w_n461_0;
	wire[1:0] w_n464_0;
	wire[1:0] w_n466_0;
	wire[2:0] w_n469_0;
	wire[1:0] w_n469_1;
	wire[1:0] w_n471_0;
	wire[1:0] w_n473_0;
	wire[1:0] w_n476_0;
	wire[1:0] w_n478_0;
	wire[2:0] w_n481_0;
	wire[1:0] w_n481_1;
	wire[2:0] w_n484_0;
	wire[1:0] w_n484_1;
	wire[2:0] w_n485_0;
	wire[2:0] w_n485_1;
	wire[2:0] w_n485_2;
	wire[2:0] w_n485_3;
	wire[2:0] w_n485_4;
	wire[2:0] w_n485_5;
	wire[2:0] w_n485_6;
	wire[2:0] w_n485_7;
	wire[2:0] w_n485_8;
	wire[2:0] w_n485_9;
	wire[2:0] w_n485_10;
	wire[2:0] w_n485_11;
	wire[2:0] w_n485_12;
	wire[2:0] w_n485_13;
	wire[2:0] w_n485_14;
	wire[2:0] w_n485_15;
	wire[2:0] w_n485_16;
	wire[2:0] w_n485_17;
	wire[2:0] w_n485_18;
	wire[2:0] w_n485_19;
	wire[2:0] w_n485_20;
	wire[2:0] w_n485_21;
	wire[2:0] w_n485_22;
	wire[2:0] w_n485_23;
	wire[2:0] w_n485_24;
	wire[2:0] w_n485_25;
	wire[2:0] w_n485_26;
	wire[2:0] w_n485_27;
	wire[2:0] w_n485_28;
	wire[2:0] w_n485_29;
	wire[2:0] w_n485_30;
	wire[2:0] w_n485_31;
	wire[2:0] w_n485_32;
	wire[2:0] w_n485_33;
	wire[2:0] w_n485_34;
	wire[2:0] w_n485_35;
	wire[2:0] w_n485_36;
	wire[2:0] w_n485_37;
	wire[2:0] w_n485_38;
	wire[2:0] w_n485_39;
	wire[2:0] w_n485_40;
	wire[2:0] w_n485_41;
	wire[2:0] w_n485_42;
	wire[2:0] w_n485_43;
	wire[2:0] w_n485_44;
	wire[2:0] w_n485_45;
	wire[2:0] w_n485_46;
	wire[2:0] w_n485_47;
	wire[2:0] w_n485_48;
	wire[2:0] w_n485_49;
	wire[2:0] w_n485_50;
	wire[2:0] w_n485_51;
	wire[2:0] w_n485_52;
	wire[2:0] w_n485_53;
	wire[2:0] w_n485_54;
	wire[2:0] w_n485_55;
	wire[2:0] w_n485_56;
	wire[2:0] w_n485_57;
	wire[2:0] w_n485_58;
	wire[2:0] w_n485_59;
	wire[2:0] w_n485_60;
	wire[2:0] w_n485_61;
	wire[2:0] w_n485_62;
	wire[1:0] w_n485_63;
	wire[1:0] w_n488_0;
	wire[1:0] w_n490_0;
	wire[1:0] w_n492_0;
	wire[1:0] w_n495_0;
	wire[1:0] w_n497_0;
	wire[2:0] w_n500_0;
	wire[1:0] w_n500_1;
	wire[1:0] w_n502_0;
	wire[1:0] w_n504_0;
	wire[1:0] w_n507_0;
	wire[1:0] w_n509_0;
	wire[2:0] w_n512_0;
	wire[1:0] w_n512_1;
	wire[1:0] w_n515_0;
	wire[1:0] w_n517_0;
	wire[1:0] w_n520_0;
	wire[1:0] w_n522_0;
	wire[2:0] w_n525_0;
	wire[1:0] w_n525_1;
	wire[1:0] w_n527_0;
	wire[1:0] w_n529_0;
	wire[1:0] w_n532_0;
	wire[1:0] w_n534_0;
	wire[2:0] w_n537_0;
	wire[1:0] w_n537_1;
	wire[2:0] w_n540_0;
	wire[1:0] w_n540_1;
	wire[1:0] w_n542_0;
	wire[1:0] w_n544_0;
	wire[1:0] w_n547_0;
	wire[1:0] w_n549_0;
	wire[2:0] w_n552_0;
	wire[1:0] w_n552_1;
	wire[1:0] w_n554_0;
	wire[1:0] w_n555_0;
	wire[1:0] w_n558_0;
	wire[1:0] w_n559_0;
	wire[2:0] w_n562_0;
	wire[1:0] w_n562_1;
	wire[1:0] w_n565_0;
	wire[1:0] w_n567_0;
	wire[1:0] w_n570_0;
	wire[1:0] w_n572_0;
	wire[2:0] w_n575_0;
	wire[1:0] w_n575_1;
	wire[1:0] w_n577_0;
	wire[1:0] w_n579_0;
	wire[1:0] w_n582_0;
	wire[1:0] w_n584_0;
	wire[2:0] w_n587_0;
	wire[1:0] w_n587_1;
	wire[2:0] w_n590_0;
	wire[1:0] w_n590_1;
	wire[1:0] w_n593_0;
	wire[1:0] w_n595_0;
	wire[1:0] w_n598_0;
	wire[1:0] w_n600_0;
	wire[2:0] w_n603_0;
	wire[1:0] w_n603_1;
	wire[1:0] w_n605_0;
	wire[1:0] w_n607_0;
	wire[1:0] w_n610_0;
	wire[1:0] w_n612_0;
	wire[2:0] w_n615_0;
	wire[1:0] w_n615_1;
	wire[1:0] w_n618_0;
	wire[1:0] w_n620_0;
	wire[1:0] w_n623_0;
	wire[1:0] w_n625_0;
	wire[2:0] w_n628_0;
	wire[1:0] w_n628_1;
	wire[1:0] w_n630_0;
	wire[1:0] w_n632_0;
	wire[1:0] w_n635_0;
	wire[1:0] w_n637_0;
	wire[2:0] w_n640_0;
	wire[1:0] w_n640_1;
	wire[2:0] w_n643_0;
	wire[1:0] w_n643_1;
	wire[1:0] w_n645_0;
	wire[1:0] w_n647_0;
	wire[1:0] w_n650_0;
	wire[1:0] w_n652_0;
	wire[2:0] w_n655_0;
	wire[1:0] w_n655_1;
	wire[1:0] w_n657_0;
	wire[1:0] w_n659_0;
	wire[1:0] w_n662_0;
	wire[1:0] w_n664_0;
	wire[2:0] w_n667_0;
	wire[1:0] w_n667_1;
	wire[1:0] w_n670_0;
	wire[1:0] w_n672_0;
	wire[1:0] w_n675_0;
	wire[1:0] w_n677_0;
	wire[2:0] w_n680_0;
	wire[1:0] w_n680_1;
	wire[1:0] w_n682_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[2:0] w_n692_0;
	wire[1:0] w_n692_1;
	wire[2:0] w_n695_0;
	wire[1:0] w_n695_1;
	wire[1:0] w_n698_0;
	wire[1:0] w_n703_0;
	wire[1:0] w_n707_0;
	wire[2:0] w_n709_0;
	wire[1:0] w_n709_1;
	wire[1:0] w_n713_0;
	wire[1:0] w_n717_0;
	wire[2:0] w_n719_0;
	wire[1:0] w_n719_1;
	wire[1:0] w_n724_0;
	wire[1:0] w_n728_0;
	wire[2:0] w_n730_0;
	wire[1:0] w_n730_1;
	wire[1:0] w_n734_0;
	wire[1:0] w_n738_0;
	wire[2:0] w_n740_0;
	wire[1:0] w_n740_1;
	wire[2:0] w_n743_0;
	wire[1:0] w_n743_1;
	wire[1:0] w_n747_0;
	wire[1:0] w_n751_0;
	wire[2:0] w_n753_0;
	wire[1:0] w_n753_1;
	wire[1:0] w_n757_0;
	wire[1:0] w_n761_0;
	wire[2:0] w_n763_0;
	wire[1:0] w_n763_1;
	wire[1:0] w_n768_0;
	wire[1:0] w_n772_0;
	wire[2:0] w_n774_0;
	wire[1:0] w_n774_1;
	wire[1:0] w_n778_0;
	wire[1:0] w_n782_0;
	wire[2:0] w_n784_0;
	wire[1:0] w_n784_1;
	wire[2:0] w_n787_0;
	wire[1:0] w_n787_1;
	wire[1:0] w_n792_0;
	wire[1:0] w_n796_0;
	wire[2:0] w_n798_0;
	wire[1:0] w_n798_1;
	wire[1:0] w_n802_0;
	wire[1:0] w_n806_0;
	wire[2:0] w_n808_0;
	wire[1:0] w_n808_1;
	wire[1:0] w_n813_0;
	wire[1:0] w_n817_0;
	wire[2:0] w_n819_0;
	wire[1:0] w_n819_1;
	wire[1:0] w_n823_0;
	wire[1:0] w_n827_0;
	wire[2:0] w_n829_0;
	wire[1:0] w_n829_1;
	wire[2:0] w_n832_0;
	wire[1:0] w_n832_1;
	wire[1:0] w_n836_0;
	wire[1:0] w_n840_0;
	wire[2:0] w_n842_0;
	wire[1:0] w_n842_1;
	wire[1:0] w_n846_0;
	wire[1:0] w_n850_0;
	wire[2:0] w_n852_0;
	wire[1:0] w_n852_1;
	wire[1:0] w_n857_0;
	wire[1:0] w_n861_0;
	wire[2:0] w_n863_0;
	wire[1:0] w_n863_1;
	wire[1:0] w_n867_0;
	wire[1:0] w_n871_0;
	wire[2:0] w_n873_0;
	wire[1:0] w_n873_1;
	wire[2:0] w_n876_0;
	wire[1:0] w_n876_1;
	wire[1:0] w_n879_0;
	wire[1:0] w_n883_0;
	wire[1:0] w_n887_0;
	wire[2:0] w_n889_0;
	wire[1:0] w_n889_1;
	wire[1:0] w_n893_0;
	wire[1:0] w_n897_0;
	wire[2:0] w_n899_0;
	wire[1:0] w_n899_1;
	wire[1:0] w_n904_0;
	wire[1:0] w_n908_0;
	wire[2:0] w_n910_0;
	wire[1:0] w_n910_1;
	wire[1:0] w_n914_0;
	wire[1:0] w_n918_0;
	wire[2:0] w_n920_0;
	wire[1:0] w_n920_1;
	wire[2:0] w_n923_0;
	wire[1:0] w_n923_1;
	wire[1:0] w_n927_0;
	wire[1:0] w_n931_0;
	wire[2:0] w_n933_0;
	wire[1:0] w_n933_1;
	wire[1:0] w_n937_0;
	wire[1:0] w_n941_0;
	wire[2:0] w_n943_0;
	wire[1:0] w_n943_1;
	wire[1:0] w_n948_0;
	wire[1:0] w_n952_0;
	wire[2:0] w_n954_0;
	wire[1:0] w_n954_1;
	wire[1:0] w_n958_0;
	wire[1:0] w_n962_0;
	wire[2:0] w_n964_0;
	wire[1:0] w_n964_1;
	wire[2:0] w_n967_0;
	wire[1:0] w_n967_1;
	wire[1:0] w_n972_0;
	wire[1:0] w_n976_0;
	wire[2:0] w_n978_0;
	wire[1:0] w_n978_1;
	wire[1:0] w_n982_0;
	wire[1:0] w_n986_0;
	wire[2:0] w_n988_0;
	wire[1:0] w_n988_1;
	wire[1:0] w_n993_0;
	wire[1:0] w_n997_0;
	wire[2:0] w_n999_0;
	wire[1:0] w_n999_1;
	wire[1:0] w_n1003_0;
	wire[1:0] w_n1007_0;
	wire[2:0] w_n1009_0;
	wire[1:0] w_n1009_1;
	wire[2:0] w_n1012_0;
	wire[1:0] w_n1012_1;
	wire[1:0] w_n1016_0;
	wire[1:0] w_n1018_0;
	wire[1:0] w_n1019_0;
	wire[2:0] w_n1022_0;
	wire[1:0] w_n1022_1;
	wire[1:0] w_n1024_0;
	wire[1:0] w_n1026_0;
	wire[1:0] w_n1029_0;
	wire[1:0] w_n1031_0;
	wire[2:0] w_n1034_0;
	wire[1:0] w_n1034_1;
	wire[1:0] w_n1037_0;
	wire[1:0] w_n1039_0;
	wire[1:0] w_n1042_0;
	wire[1:0] w_n1044_0;
	wire[2:0] w_n1047_0;
	wire[1:0] w_n1047_1;
	wire[1:0] w_n1051_0;
	wire[1:0] w_n1055_0;
	wire[2:0] w_n1057_0;
	wire[1:0] w_n1057_1;
	wire[2:0] w_n1060_0;
	wire[1:0] w_n1060_1;
	wire[1:0] w_n1063_0;
	wire[2:0] w_n1072_0;
	wire[1:0] w_n1072_1;
	wire[2:0] w_n1080_0;
	wire[1:0] w_n1080_1;
	wire[2:0] w_n1089_0;
	wire[1:0] w_n1089_1;
	wire[2:0] w_n1097_0;
	wire[1:0] w_n1097_1;
	wire[2:0] w_n1100_0;
	wire[1:0] w_n1100_1;
	wire[2:0] w_n1108_0;
	wire[1:0] w_n1108_1;
	wire[2:0] w_n1116_0;
	wire[1:0] w_n1116_1;
	wire[2:0] w_n1125_0;
	wire[1:0] w_n1125_1;
	wire[2:0] w_n1133_0;
	wire[1:0] w_n1133_1;
	wire[2:0] w_n1136_0;
	wire[1:0] w_n1136_1;
	wire[2:0] w_n1145_0;
	wire[1:0] w_n1145_1;
	wire[2:0] w_n1153_0;
	wire[1:0] w_n1153_1;
	wire[2:0] w_n1162_0;
	wire[1:0] w_n1162_1;
	wire[2:0] w_n1170_0;
	wire[1:0] w_n1170_1;
	wire[2:0] w_n1173_0;
	wire[1:0] w_n1173_1;
	wire[2:0] w_n1181_0;
	wire[1:0] w_n1181_1;
	wire[2:0] w_n1189_0;
	wire[1:0] w_n1189_1;
	wire[2:0] w_n1198_0;
	wire[1:0] w_n1198_1;
	wire[2:0] w_n1206_0;
	wire[1:0] w_n1206_1;
	wire[2:0] w_n1209_0;
	wire[1:0] w_n1209_1;
	wire[1:0] w_n1212_0;
	wire[2:0] w_n1220_0;
	wire[1:0] w_n1220_1;
	wire[2:0] w_n1228_0;
	wire[1:0] w_n1228_1;
	wire[2:0] w_n1237_0;
	wire[1:0] w_n1237_1;
	wire[2:0] w_n1245_0;
	wire[1:0] w_n1245_1;
	wire[2:0] w_n1248_0;
	wire[1:0] w_n1248_1;
	wire[2:0] w_n1256_0;
	wire[1:0] w_n1256_1;
	wire[2:0] w_n1264_0;
	wire[1:0] w_n1264_1;
	wire[2:0] w_n1273_0;
	wire[1:0] w_n1273_1;
	wire[2:0] w_n1281_0;
	wire[1:0] w_n1281_1;
	wire[2:0] w_n1284_0;
	wire[1:0] w_n1284_1;
	wire[2:0] w_n1293_0;
	wire[1:0] w_n1293_1;
	wire[2:0] w_n1301_0;
	wire[1:0] w_n1301_1;
	wire[2:0] w_n1310_0;
	wire[1:0] w_n1310_1;
	wire[2:0] w_n1318_0;
	wire[1:0] w_n1318_1;
	wire[2:0] w_n1321_0;
	wire[1:0] w_n1321_1;
	wire[2:0] w_n1329_0;
	wire[1:0] w_n1329_1;
	wire[2:0] w_n1337_0;
	wire[1:0] w_n1337_1;
	wire[2:0] w_n1346_0;
	wire[1:0] w_n1346_1;
	wire[2:0] w_n1354_0;
	wire[1:0] w_n1354_1;
	wire[2:0] w_n1357_0;
	wire[1:0] w_n1357_1;
	wire[1:0] w_n1360_0;
	wire[2:0] w_n1365_0;
	wire[1:0] w_n1365_1;
	wire[2:0] w_n1369_0;
	wire[1:0] w_n1369_1;
	wire[2:0] w_n1374_0;
	wire[1:0] w_n1374_1;
	wire[2:0] w_n1378_0;
	wire[1:0] w_n1378_1;
	wire[2:0] w_n1381_0;
	wire[1:0] w_n1381_1;
	wire[2:0] w_n1385_0;
	wire[1:0] w_n1385_1;
	wire[2:0] w_n1389_0;
	wire[1:0] w_n1389_1;
	wire[2:0] w_n1394_0;
	wire[1:0] w_n1394_1;
	wire[2:0] w_n1398_0;
	wire[1:0] w_n1398_1;
	wire[2:0] w_n1401_0;
	wire[1:0] w_n1401_1;
	wire[2:0] w_n1406_0;
	wire[1:0] w_n1406_1;
	wire[2:0] w_n1410_0;
	wire[1:0] w_n1410_1;
	wire[2:0] w_n1415_0;
	wire[1:0] w_n1415_1;
	wire[2:0] w_n1419_0;
	wire[1:0] w_n1419_1;
	wire[2:0] w_n1422_0;
	wire[1:0] w_n1422_1;
	wire[2:0] w_n1426_0;
	wire[1:0] w_n1426_1;
	wire[2:0] w_n1430_0;
	wire[1:0] w_n1430_1;
	wire[2:0] w_n1435_0;
	wire[1:0] w_n1435_1;
	wire[2:0] w_n1439_0;
	wire[1:0] w_n1439_1;
	wire[2:0] w_n1442_0;
	wire[1:0] w_n1442_1;
	wire[1:0] w_n1445_0;
	wire[2:0] w_n1449_0;
	wire[1:0] w_n1449_1;
	wire[2:0] w_n1453_0;
	wire[1:0] w_n1453_1;
	wire[2:0] w_n1458_0;
	wire[1:0] w_n1458_1;
	wire[2:0] w_n1462_0;
	wire[1:0] w_n1462_1;
	wire[2:0] w_n1465_0;
	wire[1:0] w_n1465_1;
	wire[2:0] w_n1469_0;
	wire[1:0] w_n1469_1;
	wire[2:0] w_n1473_0;
	wire[1:0] w_n1473_1;
	wire[2:0] w_n1478_0;
	wire[1:0] w_n1478_1;
	wire[2:0] w_n1482_0;
	wire[1:0] w_n1482_1;
	wire[2:0] w_n1485_0;
	wire[1:0] w_n1485_1;
	wire[2:0] w_n1490_0;
	wire[1:0] w_n1490_1;
	wire[2:0] w_n1496_0;
	wire[1:0] w_n1496_1;
	wire[2:0] w_n1505_0;
	wire[1:0] w_n1505_1;
	wire[2:0] w_n1510_0;
	wire[1:0] w_n1510_1;
	wire[2:0] w_n1513_0;
	wire[1:0] w_n1513_1;
	wire[2:0] w_n1517_0;
	wire[1:0] w_n1517_1;
	wire[2:0] w_n1521_0;
	wire[1:0] w_n1521_1;
	wire[2:0] w_n1526_0;
	wire[1:0] w_n1526_1;
	wire[2:0] w_n1530_0;
	wire[1:0] w_n1530_1;
	wire[2:0] w_n1533_0;
	wire[1:0] w_n1533_1;
	wire[1:0] w_n1536_0;
	wire[2:0] w_n1545_0;
	wire[1:0] w_n1545_1;
	wire[2:0] w_n1553_0;
	wire[1:0] w_n1553_1;
	wire[2:0] w_n1562_0;
	wire[1:0] w_n1562_1;
	wire[2:0] w_n1570_0;
	wire[1:0] w_n1570_1;
	wire[1:0] w_n1573_0;
	wire[2:0] w_n1581_0;
	wire[1:0] w_n1581_1;
	wire[2:0] w_n1589_0;
	wire[1:0] w_n1589_1;
	wire[2:0] w_n1598_0;
	wire[1:0] w_n1598_1;
	wire[2:0] w_n1606_0;
	wire[1:0] w_n1606_1;
	wire[1:0] w_n1609_0;
	wire[2:0] w_n1618_0;
	wire[1:0] w_n1618_1;
	wire[2:0] w_n1626_0;
	wire[1:0] w_n1626_1;
	wire[2:0] w_n1635_0;
	wire[1:0] w_n1635_1;
	wire[2:0] w_n1643_0;
	wire[1:0] w_n1643_1;
	wire[1:0] w_n1646_0;
	wire[2:0] w_n1654_0;
	wire[1:0] w_n1654_1;
	wire[2:0] w_n1662_0;
	wire[1:0] w_n1662_1;
	wire[2:0] w_n1671_0;
	wire[1:0] w_n1671_1;
	wire[2:0] w_n1679_0;
	wire[1:0] w_n1679_1;
	wire[1:0] w_n1682_0;
	wire[2:0] w_n1691_0;
	wire[1:0] w_n1691_1;
	wire[2:0] w_n1699_0;
	wire[1:0] w_n1699_1;
	wire[2:0] w_n1708_0;
	wire[1:0] w_n1708_1;
	wire[2:0] w_n1716_0;
	wire[1:0] w_n1716_1;
	wire[1:0] w_n1719_0;
	wire[2:0] w_n1727_0;
	wire[1:0] w_n1727_1;
	wire[2:0] w_n1735_0;
	wire[1:0] w_n1735_1;
	wire[2:0] w_n1744_0;
	wire[1:0] w_n1744_1;
	wire[2:0] w_n1752_0;
	wire[1:0] w_n1752_1;
	wire[1:0] w_n1755_0;
	wire[2:0] w_n1764_0;
	wire[1:0] w_n1764_1;
	wire[2:0] w_n1772_0;
	wire[1:0] w_n1772_1;
	wire[2:0] w_n1781_0;
	wire[1:0] w_n1781_1;
	wire[2:0] w_n1789_0;
	wire[1:0] w_n1789_1;
	wire[1:0] w_n1792_0;
	wire[2:0] w_n1800_0;
	wire[1:0] w_n1800_1;
	wire[2:0] w_n1808_0;
	wire[1:0] w_n1808_1;
	wire[2:0] w_n1817_0;
	wire[1:0] w_n1817_1;
	wire[2:0] w_n1825_0;
	wire[1:0] w_n1825_1;
	wire[1:0] w_n1828_0;
	wire[2:0] w_n1837_0;
	wire[1:0] w_n1837_1;
	wire[2:0] w_n1845_0;
	wire[1:0] w_n1845_1;
	wire[2:0] w_n1854_0;
	wire[1:0] w_n1854_1;
	wire[2:0] w_n1862_0;
	wire[1:0] w_n1862_1;
	wire[1:0] w_n1865_0;
	wire[2:0] w_n1873_0;
	wire[1:0] w_n1873_1;
	wire[2:0] w_n1881_0;
	wire[1:0] w_n1881_1;
	wire[2:0] w_n1890_0;
	wire[1:0] w_n1890_1;
	wire[2:0] w_n1898_0;
	wire[1:0] w_n1898_1;
	wire[1:0] w_n1901_0;
	wire[2:0] w_n1910_0;
	wire[1:0] w_n1910_1;
	wire[2:0] w_n1918_0;
	wire[1:0] w_n1918_1;
	wire[2:0] w_n1927_0;
	wire[1:0] w_n1927_1;
	wire[2:0] w_n1935_0;
	wire[1:0] w_n1935_1;
	wire[1:0] w_n1938_0;
	wire[2:0] w_n1946_0;
	wire[1:0] w_n1946_1;
	wire[2:0] w_n1954_0;
	wire[1:0] w_n1954_1;
	wire[2:0] w_n1963_0;
	wire[1:0] w_n1963_1;
	wire[2:0] w_n1971_0;
	wire[1:0] w_n1971_1;
	wire[1:0] w_n1974_0;
	wire[2:0] w_n1983_0;
	wire[1:0] w_n1983_1;
	wire[2:0] w_n1991_0;
	wire[1:0] w_n1991_1;
	wire[2:0] w_n2000_0;
	wire[1:0] w_n2000_1;
	wire[2:0] w_n2008_0;
	wire[1:0] w_n2008_1;
	wire[1:0] w_n2011_0;
	wire[2:0] w_n2019_0;
	wire[1:0] w_n2019_1;
	wire[2:0] w_n2027_0;
	wire[1:0] w_n2027_1;
	wire[2:0] w_n2036_0;
	wire[1:0] w_n2036_1;
	wire[2:0] w_n2044_0;
	wire[1:0] w_n2044_1;
	wire[1:0] w_n2047_0;
	wire[2:0] w_n2056_0;
	wire[1:0] w_n2056_1;
	wire[2:0] w_n2064_0;
	wire[1:0] w_n2064_1;
	wire[2:0] w_n2073_0;
	wire[1:0] w_n2073_1;
	wire[2:0] w_n2081_0;
	wire[1:0] w_n2081_1;
	wire[1:0] w_n2084_0;
	wire[2:0] w_n2092_0;
	wire[1:0] w_n2092_1;
	wire[2:0] w_n2100_0;
	wire[1:0] w_n2100_1;
	wire[2:0] w_n2109_0;
	wire[1:0] w_n2109_1;
	wire[2:0] w_n2117_0;
	wire[1:0] w_n2117_1;
	wire[1:0] w_n2120_0;
	wire[2:0] w_n2129_0;
	wire[1:0] w_n2129_1;
	wire[2:0] w_n2137_0;
	wire[1:0] w_n2137_1;
	wire[2:0] w_n2146_0;
	wire[1:0] w_n2146_1;
	wire[2:0] w_n2154_0;
	wire[1:0] w_n2154_1;
	wire[1:0] w_n2157_0;
	wire[2:0] w_n2165_0;
	wire[1:0] w_n2165_1;
	wire[2:0] w_n2173_0;
	wire[1:0] w_n2173_1;
	wire[2:0] w_n2182_0;
	wire[1:0] w_n2182_1;
	wire[2:0] w_n2190_0;
	wire[1:0] w_n2190_1;
	wire[1:0] w_n2193_0;
	wire[2:0] w_n2202_0;
	wire[1:0] w_n2202_1;
	wire[2:0] w_n2210_0;
	wire[1:0] w_n2210_1;
	wire[2:0] w_n2219_0;
	wire[1:0] w_n2219_1;
	wire[2:0] w_n2227_0;
	wire[1:0] w_n2227_1;
	wire[1:0] w_n2230_0;
	wire[2:0] w_n2238_0;
	wire[1:0] w_n2238_1;
	wire[2:0] w_n2246_0;
	wire[1:0] w_n2246_1;
	wire[2:0] w_n2255_0;
	wire[1:0] w_n2255_1;
	wire[2:0] w_n2263_0;
	wire[1:0] w_n2263_1;
	wire[1:0] w_n2266_0;
	wire[2:0] w_n2275_0;
	wire[1:0] w_n2275_1;
	wire[2:0] w_n2283_0;
	wire[1:0] w_n2283_1;
	wire[2:0] w_n2292_0;
	wire[1:0] w_n2292_1;
	wire[2:0] w_n2300_0;
	wire[1:0] w_n2300_1;
	wire[1:0] w_n2303_0;
	wire[2:0] w_n2311_0;
	wire[1:0] w_n2311_1;
	wire[2:0] w_n2319_0;
	wire[1:0] w_n2319_1;
	wire[2:0] w_n2328_0;
	wire[1:0] w_n2328_1;
	wire[2:0] w_n2336_0;
	wire[1:0] w_n2336_1;
	wire[1:0] w_n2339_0;
	wire[2:0] w_n2348_0;
	wire[1:0] w_n2348_1;
	wire[2:0] w_n2356_0;
	wire[1:0] w_n2356_1;
	wire[2:0] w_n2365_0;
	wire[1:0] w_n2365_1;
	wire[2:0] w_n2373_0;
	wire[1:0] w_n2373_1;
	wire[1:0] w_n2376_0;
	wire[2:0] w_n2384_0;
	wire[1:0] w_n2384_1;
	wire[2:0] w_n2392_0;
	wire[1:0] w_n2392_1;
	wire[2:0] w_n2401_0;
	wire[1:0] w_n2401_1;
	wire[2:0] w_n2409_0;
	wire[1:0] w_n2409_1;
	wire[1:0] w_n2412_0;
	wire[1:0] w_n2421_0;
	wire[1:0] w_n2429_0;
	wire[1:0] w_n2438_0;
	wire[1:0] w_n2446_0;
	wire[1:0] w_n2455_0;
	wire[1:0] w_n2463_0;
	wire[1:0] w_n2472_0;
	wire[1:0] w_n2480_0;
	wire[1:0] w_n2489_0;
	wire[1:0] w_n2497_0;
	wire[1:0] w_n2506_0;
	wire[1:0] w_n2514_0;
	wire[1:0] w_n2523_0;
	wire[1:0] w_n2531_0;
	wire[1:0] w_n2540_0;
	wire[1:0] w_n2548_0;
	wire[1:0] w_n2557_0;
	wire[1:0] w_n2565_0;
	wire[1:0] w_n2574_0;
	wire[1:0] w_n2582_0;
	wire[1:0] w_n2591_0;
	wire[1:0] w_n2599_0;
	wire[1:0] w_n2608_0;
	wire[1:0] w_n2616_0;
	wire[1:0] w_n2625_0;
	wire[1:0] w_n2633_0;
	wire[1:0] w_n2642_0;
	wire[1:0] w_n2650_0;
	wire[1:0] w_n2659_0;
	wire[1:0] w_n2667_0;
	wire[1:0] w_n2676_0;
	wire[1:0] w_n2684_0;
	wire[1:0] w_n2693_0;
	wire[1:0] w_n2701_0;
	wire[1:0] w_n2710_0;
	wire[1:0] w_n2718_0;
	wire[1:0] w_n2727_0;
	wire[1:0] w_n2735_0;
	wire[1:0] w_n2744_0;
	wire[1:0] w_n2752_0;
	wire[1:0] w_n2761_0;
	wire[1:0] w_n2769_0;
	wire[1:0] w_n2778_0;
	wire[1:0] w_n2786_0;
	wire[1:0] w_n2795_0;
	wire[1:0] w_n2803_0;
	wire[1:0] w_n2812_0;
	wire[1:0] w_n2820_0;
	wire[1:0] w_n2829_0;
	wire[1:0] w_n2837_0;
	wire[1:0] w_n2846_0;
	wire[1:0] w_n2854_0;
	wire[1:0] w_n2863_0;
	wire[1:0] w_n2871_0;
	wire[1:0] w_n2880_0;
	wire[1:0] w_n2888_0;
	wire[1:0] w_n2897_0;
	wire[1:0] w_n2905_0;
	wire[1:0] w_n2914_0;
	wire[1:0] w_n2922_0;
	wire[1:0] w_n2931_0;
	wire[1:0] w_n2939_0;
	wire[1:0] w_n2948_0;
	wire[1:0] w_n2956_0;
	wire[1:0] w_n2965_0;
	wire[1:0] w_n2973_0;
	wire[1:0] w_n2982_0;
	wire[1:0] w_n2990_0;
	wire[1:0] w_n2999_0;
	wire[1:0] w_n3007_0;
	wire[1:0] w_n3016_0;
	wire[1:0] w_n3024_0;
	wire[1:0] w_n3033_0;
	wire[1:0] w_n3041_0;
	wire[1:0] w_n3050_0;
	wire[1:0] w_n3058_0;
	wire[1:0] w_n3067_0;
	wire[1:0] w_n3075_0;
	wire[1:0] w_n3084_0;
	wire[1:0] w_n3092_0;
	wire[1:0] w_n3101_0;
	wire[1:0] w_n3109_0;
	wire[1:0] w_n3118_0;
	wire[1:0] w_n3126_0;
	wire[1:0] w_n3135_0;
	wire[1:0] w_n3143_0;
	wire[1:0] w_n3152_0;
	wire[1:0] w_n3160_0;
	wire[1:0] w_n3169_0;
	wire[1:0] w_n3177_0;
	wire[1:0] w_n3186_0;
	wire[1:0] w_n3194_0;
	wire[1:0] w_n3203_0;
	wire[1:0] w_n3211_0;
	wire[1:0] w_n3220_0;
	wire[1:0] w_n3228_0;
	jnot g0000(.din(w_shift6_63[2]),.dout(n263),.clk(gclk));
	jnot g0001(.din(w_shift2_0[2]),.dout(n264),.clk(gclk));
	jnot g0002(.din(w_shift3_0[2]),.dout(n265),.clk(gclk));
	jand g0003(.dina(w_n265_0[1]),.dinb(w_n264_0[1]),.dout(n266),.clk(gclk));
	jand g0004(.dina(w_shift0_63[2]),.dinb(w_a79_0[1]),.dout(n267),.clk(gclk));
	jor g0005(.dina(w_n267_0[1]),.dinb(w_shift1_96[2]),.dout(n268),.clk(gclk));
	jnot g0006(.din(w_shift1_96[1]),.dout(n269),.clk(gclk));
	jnot g0007(.din(w_shift0_63[1]),.dout(n270),.clk(gclk));
	jand g0008(.dina(w_n270_63[1]),.dinb(w_a78_0[1]),.dout(n271),.clk(gclk));
	jor g0009(.dina(w_n271_0[1]),.dinb(w_n269_96[1]),.dout(n272),.clk(gclk));
	jand g0010(.dina(n272),.dinb(n268),.dout(n273),.clk(gclk));
	jand g0011(.dina(w_shift0_63[0]),.dinb(w_a77_0[1]),.dout(n274),.clk(gclk));
	jand g0012(.dina(w_n274_0[1]),.dinb(w_shift1_96[0]),.dout(n275),.clk(gclk));
	jand g0013(.dina(w_n270_63[0]),.dinb(w_a80_0[1]),.dout(n276),.clk(gclk));
	jand g0014(.dina(w_n276_0[1]),.dinb(w_n269_96[0]),.dout(n277),.clk(gclk));
	jor g0015(.dina(n277),.dinb(n275),.dout(n278),.clk(gclk));
	jor g0016(.dina(n278),.dinb(n273),.dout(n279),.clk(gclk));
	jand g0017(.dina(w_n279_1[1]),.dinb(w_n266_63[1]),.dout(n280),.clk(gclk));
	jand g0018(.dina(w_shift3_0[1]),.dinb(w_n264_0[0]),.dout(n281),.clk(gclk));
	jand g0019(.dina(w_shift0_62[2]),.dinb(w_a71_0[1]),.dout(n282),.clk(gclk));
	jor g0020(.dina(w_n282_0[1]),.dinb(w_shift1_95[2]),.dout(n283),.clk(gclk));
	jand g0021(.dina(w_n270_62[2]),.dinb(w_a70_0[1]),.dout(n284),.clk(gclk));
	jor g0022(.dina(w_n284_0[1]),.dinb(w_n269_95[2]),.dout(n285),.clk(gclk));
	jand g0023(.dina(n285),.dinb(n283),.dout(n286),.clk(gclk));
	jand g0024(.dina(w_shift0_62[1]),.dinb(w_a69_0[1]),.dout(n287),.clk(gclk));
	jand g0025(.dina(w_n287_0[1]),.dinb(w_shift1_95[1]),.dout(n288),.clk(gclk));
	jand g0026(.dina(w_n270_62[1]),.dinb(w_a72_0[1]),.dout(n289),.clk(gclk));
	jand g0027(.dina(w_n289_0[1]),.dinb(w_n269_95[1]),.dout(n290),.clk(gclk));
	jor g0028(.dina(n290),.dinb(n288),.dout(n291),.clk(gclk));
	jor g0029(.dina(n291),.dinb(n286),.dout(n292),.clk(gclk));
	jand g0030(.dina(w_n292_1[1]),.dinb(w_n281_63[1]),.dout(n293),.clk(gclk));
	jor g0031(.dina(n293),.dinb(n280),.dout(n294),.clk(gclk));
	jand g0032(.dina(w_n265_0[0]),.dinb(w_shift2_0[1]),.dout(n295),.clk(gclk));
	jand g0033(.dina(w_shift0_62[0]),.dinb(w_a75_0[1]),.dout(n296),.clk(gclk));
	jor g0034(.dina(w_n296_0[1]),.dinb(w_shift1_95[0]),.dout(n297),.clk(gclk));
	jand g0035(.dina(w_n270_62[0]),.dinb(w_a74_0[1]),.dout(n298),.clk(gclk));
	jor g0036(.dina(w_n298_0[1]),.dinb(w_n269_95[0]),.dout(n299),.clk(gclk));
	jand g0037(.dina(n299),.dinb(n297),.dout(n300),.clk(gclk));
	jand g0038(.dina(w_shift0_61[2]),.dinb(w_a73_0[1]),.dout(n301),.clk(gclk));
	jand g0039(.dina(w_n301_0[1]),.dinb(w_shift1_94[2]),.dout(n302),.clk(gclk));
	jand g0040(.dina(w_n270_61[2]),.dinb(w_a76_0[1]),.dout(n303),.clk(gclk));
	jand g0041(.dina(w_n303_0[1]),.dinb(w_n269_94[2]),.dout(n304),.clk(gclk));
	jor g0042(.dina(n304),.dinb(n302),.dout(n305),.clk(gclk));
	jor g0043(.dina(n305),.dinb(n300),.dout(n306),.clk(gclk));
	jand g0044(.dina(w_n306_1[1]),.dinb(w_n295_63[1]),.dout(n307),.clk(gclk));
	jand g0045(.dina(w_shift3_0[0]),.dinb(w_shift2_0[0]),.dout(n308),.clk(gclk));
	jand g0046(.dina(w_shift0_61[1]),.dinb(w_a67_0[1]),.dout(n309),.clk(gclk));
	jor g0047(.dina(w_n309_0[1]),.dinb(w_shift1_94[1]),.dout(n310),.clk(gclk));
	jand g0048(.dina(w_n270_61[1]),.dinb(w_a66_0[1]),.dout(n311),.clk(gclk));
	jor g0049(.dina(w_n311_0[1]),.dinb(w_n269_94[1]),.dout(n312),.clk(gclk));
	jand g0050(.dina(n312),.dinb(n310),.dout(n313),.clk(gclk));
	jand g0051(.dina(w_shift0_61[0]),.dinb(w_a65_0[1]),.dout(n314),.clk(gclk));
	jand g0052(.dina(w_n314_0[1]),.dinb(w_shift1_94[0]),.dout(n315),.clk(gclk));
	jand g0053(.dina(w_n270_61[0]),.dinb(w_a68_0[1]),.dout(n316),.clk(gclk));
	jand g0054(.dina(w_n316_0[1]),.dinb(w_n269_94[0]),.dout(n317),.clk(gclk));
	jor g0055(.dina(n317),.dinb(n315),.dout(n318),.clk(gclk));
	jor g0056(.dina(n318),.dinb(n313),.dout(n319),.clk(gclk));
	jand g0057(.dina(w_n319_1[1]),.dinb(w_n308_63[1]),.dout(n320),.clk(gclk));
	jor g0058(.dina(n320),.dinb(n307),.dout(n321),.clk(gclk));
	jor g0059(.dina(n321),.dinb(n294),.dout(n322),.clk(gclk));
	jand g0060(.dina(w_shift5_0[2]),.dinb(w_shift4_0[2]),.dout(n323),.clk(gclk));
	jand g0061(.dina(w_n323_63[1]),.dinb(w_n322_1[1]),.dout(n324),.clk(gclk));
	jand g0062(.dina(w_shift0_60[2]),.dinb(w_a111_0[1]),.dout(n325),.clk(gclk));
	jor g0063(.dina(w_n325_0[1]),.dinb(w_shift1_93[2]),.dout(n326),.clk(gclk));
	jand g0064(.dina(w_n270_60[2]),.dinb(w_a110_0[1]),.dout(n327),.clk(gclk));
	jor g0065(.dina(w_n327_0[1]),.dinb(w_n269_93[2]),.dout(n328),.clk(gclk));
	jand g0066(.dina(n328),.dinb(n326),.dout(n329),.clk(gclk));
	jand g0067(.dina(w_shift0_60[1]),.dinb(w_a109_0[1]),.dout(n330),.clk(gclk));
	jand g0068(.dina(w_n330_0[1]),.dinb(w_shift1_93[1]),.dout(n331),.clk(gclk));
	jand g0069(.dina(w_n270_60[1]),.dinb(w_a112_0[1]),.dout(n332),.clk(gclk));
	jand g0070(.dina(w_n332_0[1]),.dinb(w_n269_93[1]),.dout(n333),.clk(gclk));
	jor g0071(.dina(n333),.dinb(n331),.dout(n334),.clk(gclk));
	jor g0072(.dina(n334),.dinb(n329),.dout(n335),.clk(gclk));
	jand g0073(.dina(w_n335_1[1]),.dinb(w_n266_63[0]),.dout(n336),.clk(gclk));
	jand g0074(.dina(w_shift0_60[0]),.dinb(w_a103_0[1]),.dout(n337),.clk(gclk));
	jor g0075(.dina(w_n337_0[1]),.dinb(w_shift1_93[0]),.dout(n338),.clk(gclk));
	jand g0076(.dina(w_n270_60[0]),.dinb(w_a102_0[1]),.dout(n339),.clk(gclk));
	jor g0077(.dina(w_n339_0[1]),.dinb(w_n269_93[0]),.dout(n340),.clk(gclk));
	jand g0078(.dina(n340),.dinb(n338),.dout(n341),.clk(gclk));
	jand g0079(.dina(w_shift0_59[2]),.dinb(w_a101_0[1]),.dout(n342),.clk(gclk));
	jand g0080(.dina(w_n342_0[1]),.dinb(w_shift1_92[2]),.dout(n343),.clk(gclk));
	jand g0081(.dina(w_n270_59[2]),.dinb(w_a104_0[1]),.dout(n344),.clk(gclk));
	jand g0082(.dina(w_n344_0[1]),.dinb(w_n269_92[2]),.dout(n345),.clk(gclk));
	jor g0083(.dina(n345),.dinb(n343),.dout(n346),.clk(gclk));
	jor g0084(.dina(n346),.dinb(n341),.dout(n347),.clk(gclk));
	jand g0085(.dina(w_n347_1[1]),.dinb(w_n281_63[0]),.dout(n348),.clk(gclk));
	jor g0086(.dina(n348),.dinb(n336),.dout(n349),.clk(gclk));
	jand g0087(.dina(w_shift0_59[1]),.dinb(w_a107_0[1]),.dout(n350),.clk(gclk));
	jor g0088(.dina(w_n350_0[1]),.dinb(w_shift1_92[1]),.dout(n351),.clk(gclk));
	jand g0089(.dina(w_n270_59[1]),.dinb(w_a106_0[1]),.dout(n352),.clk(gclk));
	jor g0090(.dina(w_n352_0[1]),.dinb(w_n269_92[1]),.dout(n353),.clk(gclk));
	jand g0091(.dina(n353),.dinb(n351),.dout(n354),.clk(gclk));
	jand g0092(.dina(w_shift0_59[0]),.dinb(w_a105_0[1]),.dout(n355),.clk(gclk));
	jand g0093(.dina(w_n355_0[1]),.dinb(w_shift1_92[0]),.dout(n356),.clk(gclk));
	jand g0094(.dina(w_n270_59[0]),.dinb(w_a108_0[1]),.dout(n357),.clk(gclk));
	jand g0095(.dina(w_n357_0[1]),.dinb(w_n269_92[0]),.dout(n358),.clk(gclk));
	jor g0096(.dina(n358),.dinb(n356),.dout(n359),.clk(gclk));
	jor g0097(.dina(n359),.dinb(n354),.dout(n360),.clk(gclk));
	jand g0098(.dina(w_n360_1[1]),.dinb(w_n295_63[0]),.dout(n361),.clk(gclk));
	jand g0099(.dina(w_shift0_58[2]),.dinb(w_a99_0[1]),.dout(n362),.clk(gclk));
	jor g0100(.dina(w_n362_0[1]),.dinb(w_shift1_91[2]),.dout(n363),.clk(gclk));
	jand g0101(.dina(w_n270_58[2]),.dinb(w_a98_0[1]),.dout(n364),.clk(gclk));
	jor g0102(.dina(w_n364_0[1]),.dinb(w_n269_91[2]),.dout(n365),.clk(gclk));
	jand g0103(.dina(n365),.dinb(n363),.dout(n366),.clk(gclk));
	jand g0104(.dina(w_shift0_58[1]),.dinb(w_a97_0[1]),.dout(n367),.clk(gclk));
	jand g0105(.dina(w_n367_0[1]),.dinb(w_shift1_91[1]),.dout(n368),.clk(gclk));
	jand g0106(.dina(w_n270_58[1]),.dinb(w_a100_0[1]),.dout(n369),.clk(gclk));
	jand g0107(.dina(w_n369_0[1]),.dinb(w_n269_91[1]),.dout(n370),.clk(gclk));
	jor g0108(.dina(n370),.dinb(n368),.dout(n371),.clk(gclk));
	jor g0109(.dina(n371),.dinb(n366),.dout(n372),.clk(gclk));
	jand g0110(.dina(w_n372_1[1]),.dinb(w_n308_63[0]),.dout(n373),.clk(gclk));
	jor g0111(.dina(n373),.dinb(n361),.dout(n374),.clk(gclk));
	jor g0112(.dina(n374),.dinb(n349),.dout(n375),.clk(gclk));
	jnot g0113(.din(w_shift5_0[1]),.dout(n376),.clk(gclk));
	jand g0114(.dina(w_n376_0[1]),.dinb(w_shift4_0[1]),.dout(n377),.clk(gclk));
	jand g0115(.dina(w_n377_63[1]),.dinb(w_n375_1[1]),.dout(n378),.clk(gclk));
	jor g0116(.dina(n378),.dinb(n324),.dout(n379),.clk(gclk));
	jand g0117(.dina(w_shift0_58[0]),.dinb(w_a95_0[1]),.dout(n380),.clk(gclk));
	jor g0118(.dina(w_n380_0[1]),.dinb(w_shift1_91[0]),.dout(n381),.clk(gclk));
	jand g0119(.dina(w_n270_58[0]),.dinb(w_a94_0[1]),.dout(n382),.clk(gclk));
	jor g0120(.dina(w_n382_0[1]),.dinb(w_n269_91[0]),.dout(n383),.clk(gclk));
	jand g0121(.dina(n383),.dinb(n381),.dout(n384),.clk(gclk));
	jand g0122(.dina(w_shift0_57[2]),.dinb(w_a93_0[1]),.dout(n385),.clk(gclk));
	jand g0123(.dina(w_n385_0[1]),.dinb(w_shift1_90[2]),.dout(n386),.clk(gclk));
	jand g0124(.dina(w_n270_57[2]),.dinb(w_a96_0[1]),.dout(n387),.clk(gclk));
	jand g0125(.dina(w_n387_0[1]),.dinb(w_n269_90[2]),.dout(n388),.clk(gclk));
	jor g0126(.dina(n388),.dinb(n386),.dout(n389),.clk(gclk));
	jor g0127(.dina(n389),.dinb(n384),.dout(n390),.clk(gclk));
	jand g0128(.dina(w_n390_1[1]),.dinb(w_n266_62[2]),.dout(n391),.clk(gclk));
	jand g0129(.dina(w_shift0_57[1]),.dinb(w_a87_0[1]),.dout(n392),.clk(gclk));
	jor g0130(.dina(w_n392_0[1]),.dinb(w_shift1_90[1]),.dout(n393),.clk(gclk));
	jand g0131(.dina(w_n270_57[1]),.dinb(w_a86_0[1]),.dout(n394),.clk(gclk));
	jor g0132(.dina(w_n394_0[1]),.dinb(w_n269_90[1]),.dout(n395),.clk(gclk));
	jand g0133(.dina(n395),.dinb(n393),.dout(n396),.clk(gclk));
	jand g0134(.dina(w_shift0_57[0]),.dinb(w_a85_0[1]),.dout(n397),.clk(gclk));
	jand g0135(.dina(w_n397_0[1]),.dinb(w_shift1_90[0]),.dout(n398),.clk(gclk));
	jand g0136(.dina(w_n270_57[0]),.dinb(w_a88_0[1]),.dout(n399),.clk(gclk));
	jand g0137(.dina(w_n399_0[1]),.dinb(w_n269_90[0]),.dout(n400),.clk(gclk));
	jor g0138(.dina(n400),.dinb(n398),.dout(n401),.clk(gclk));
	jor g0139(.dina(n401),.dinb(n396),.dout(n402),.clk(gclk));
	jand g0140(.dina(w_n402_1[1]),.dinb(w_n281_62[2]),.dout(n403),.clk(gclk));
	jor g0141(.dina(n403),.dinb(n391),.dout(n404),.clk(gclk));
	jand g0142(.dina(w_shift0_56[2]),.dinb(w_a91_0[1]),.dout(n405),.clk(gclk));
	jor g0143(.dina(w_n405_0[1]),.dinb(w_shift1_89[2]),.dout(n406),.clk(gclk));
	jand g0144(.dina(w_n270_56[2]),.dinb(w_a90_0[1]),.dout(n407),.clk(gclk));
	jor g0145(.dina(w_n407_0[1]),.dinb(w_n269_89[2]),.dout(n408),.clk(gclk));
	jand g0146(.dina(n408),.dinb(n406),.dout(n409),.clk(gclk));
	jand g0147(.dina(w_shift0_56[1]),.dinb(w_a89_0[1]),.dout(n410),.clk(gclk));
	jand g0148(.dina(w_n410_0[1]),.dinb(w_shift1_89[1]),.dout(n411),.clk(gclk));
	jand g0149(.dina(w_n270_56[1]),.dinb(w_a92_0[1]),.dout(n412),.clk(gclk));
	jand g0150(.dina(w_n412_0[1]),.dinb(w_n269_89[1]),.dout(n413),.clk(gclk));
	jor g0151(.dina(n413),.dinb(n411),.dout(n414),.clk(gclk));
	jor g0152(.dina(n414),.dinb(n409),.dout(n415),.clk(gclk));
	jand g0153(.dina(w_n415_1[1]),.dinb(w_n295_62[2]),.dout(n416),.clk(gclk));
	jand g0154(.dina(w_shift0_56[0]),.dinb(w_a83_0[1]),.dout(n417),.clk(gclk));
	jor g0155(.dina(w_n417_0[1]),.dinb(w_shift1_89[0]),.dout(n418),.clk(gclk));
	jand g0156(.dina(w_n270_56[0]),.dinb(w_a82_0[1]),.dout(n419),.clk(gclk));
	jor g0157(.dina(w_n419_0[1]),.dinb(w_n269_89[0]),.dout(n420),.clk(gclk));
	jand g0158(.dina(n420),.dinb(n418),.dout(n421),.clk(gclk));
	jand g0159(.dina(w_shift0_55[2]),.dinb(w_a81_0[1]),.dout(n422),.clk(gclk));
	jand g0160(.dina(w_n422_0[1]),.dinb(w_shift1_88[2]),.dout(n423),.clk(gclk));
	jand g0161(.dina(w_n270_55[2]),.dinb(w_a84_0[1]),.dout(n424),.clk(gclk));
	jand g0162(.dina(w_n424_0[1]),.dinb(w_n269_88[2]),.dout(n425),.clk(gclk));
	jor g0163(.dina(n425),.dinb(n423),.dout(n426),.clk(gclk));
	jor g0164(.dina(n426),.dinb(n421),.dout(n427),.clk(gclk));
	jand g0165(.dina(w_n427_1[1]),.dinb(w_n308_62[2]),.dout(n428),.clk(gclk));
	jor g0166(.dina(n428),.dinb(n416),.dout(n429),.clk(gclk));
	jor g0167(.dina(n429),.dinb(n404),.dout(n430),.clk(gclk));
	jnot g0168(.din(w_shift4_0[0]),.dout(n431),.clk(gclk));
	jand g0169(.dina(w_shift5_0[0]),.dinb(w_n431_0[1]),.dout(n432),.clk(gclk));
	jand g0170(.dina(w_n432_63[1]),.dinb(w_n430_1[1]),.dout(n433),.clk(gclk));
	jand g0171(.dina(w_shift0_55[1]),.dinb(w_a127_0[1]),.dout(n434),.clk(gclk));
	jor g0172(.dina(w_n434_0[1]),.dinb(w_shift1_88[1]),.dout(n435),.clk(gclk));
	jand g0173(.dina(w_n270_55[1]),.dinb(w_a126_0[1]),.dout(n436),.clk(gclk));
	jor g0174(.dina(w_n436_0[1]),.dinb(w_n269_88[1]),.dout(n437),.clk(gclk));
	jand g0175(.dina(n437),.dinb(n435),.dout(n438),.clk(gclk));
	jand g0176(.dina(w_shift0_55[0]),.dinb(w_a125_0[1]),.dout(n439),.clk(gclk));
	jand g0177(.dina(w_n439_0[1]),.dinb(w_shift1_88[0]),.dout(n440),.clk(gclk));
	jand g0178(.dina(w_n270_55[0]),.dinb(w_a0_0[1]),.dout(n441),.clk(gclk));
	jand g0179(.dina(w_n441_0[1]),.dinb(w_n269_88[0]),.dout(n442),.clk(gclk));
	jor g0180(.dina(n442),.dinb(n440),.dout(n443),.clk(gclk));
	jor g0181(.dina(n443),.dinb(n438),.dout(n444),.clk(gclk));
	jand g0182(.dina(w_n444_1[1]),.dinb(w_n266_62[1]),.dout(n445),.clk(gclk));
	jand g0183(.dina(w_shift0_54[2]),.dinb(w_a119_0[1]),.dout(n446),.clk(gclk));
	jor g0184(.dina(w_n446_0[1]),.dinb(w_shift1_87[2]),.dout(n447),.clk(gclk));
	jand g0185(.dina(w_n270_54[2]),.dinb(w_a118_0[1]),.dout(n448),.clk(gclk));
	jor g0186(.dina(w_n448_0[1]),.dinb(w_n269_87[2]),.dout(n449),.clk(gclk));
	jand g0187(.dina(n449),.dinb(n447),.dout(n450),.clk(gclk));
	jand g0188(.dina(w_shift0_54[1]),.dinb(w_a117_0[1]),.dout(n451),.clk(gclk));
	jand g0189(.dina(w_n451_0[1]),.dinb(w_shift1_87[1]),.dout(n452),.clk(gclk));
	jand g0190(.dina(w_n270_54[1]),.dinb(w_a120_0[1]),.dout(n453),.clk(gclk));
	jand g0191(.dina(w_n453_0[1]),.dinb(w_n269_87[1]),.dout(n454),.clk(gclk));
	jor g0192(.dina(n454),.dinb(n452),.dout(n455),.clk(gclk));
	jor g0193(.dina(n455),.dinb(n450),.dout(n456),.clk(gclk));
	jand g0194(.dina(w_n456_1[1]),.dinb(w_n281_62[1]),.dout(n457),.clk(gclk));
	jor g0195(.dina(n457),.dinb(n445),.dout(n458),.clk(gclk));
	jand g0196(.dina(w_shift0_54[0]),.dinb(w_a123_0[1]),.dout(n459),.clk(gclk));
	jor g0197(.dina(w_n459_0[1]),.dinb(w_shift1_87[0]),.dout(n460),.clk(gclk));
	jand g0198(.dina(w_n270_54[0]),.dinb(w_a122_0[1]),.dout(n461),.clk(gclk));
	jor g0199(.dina(w_n461_0[1]),.dinb(w_n269_87[0]),.dout(n462),.clk(gclk));
	jand g0200(.dina(n462),.dinb(n460),.dout(n463),.clk(gclk));
	jand g0201(.dina(w_shift0_53[2]),.dinb(w_a121_0[1]),.dout(n464),.clk(gclk));
	jand g0202(.dina(w_n464_0[1]),.dinb(w_shift1_86[2]),.dout(n465),.clk(gclk));
	jand g0203(.dina(w_n270_53[2]),.dinb(w_a124_0[1]),.dout(n466),.clk(gclk));
	jand g0204(.dina(w_n466_0[1]),.dinb(w_n269_86[2]),.dout(n467),.clk(gclk));
	jor g0205(.dina(n467),.dinb(n465),.dout(n468),.clk(gclk));
	jor g0206(.dina(n468),.dinb(n463),.dout(n469),.clk(gclk));
	jand g0207(.dina(w_n469_1[1]),.dinb(w_n295_62[1]),.dout(n470),.clk(gclk));
	jand g0208(.dina(w_shift0_53[1]),.dinb(w_a115_0[1]),.dout(n471),.clk(gclk));
	jor g0209(.dina(w_n471_0[1]),.dinb(w_shift1_86[1]),.dout(n472),.clk(gclk));
	jand g0210(.dina(w_n270_53[1]),.dinb(w_a114_0[1]),.dout(n473),.clk(gclk));
	jor g0211(.dina(w_n473_0[1]),.dinb(w_n269_86[1]),.dout(n474),.clk(gclk));
	jand g0212(.dina(n474),.dinb(n472),.dout(n475),.clk(gclk));
	jand g0213(.dina(w_shift0_53[0]),.dinb(w_a113_0[1]),.dout(n476),.clk(gclk));
	jand g0214(.dina(w_n476_0[1]),.dinb(w_shift1_86[0]),.dout(n477),.clk(gclk));
	jand g0215(.dina(w_n270_53[0]),.dinb(w_a116_0[1]),.dout(n478),.clk(gclk));
	jand g0216(.dina(w_n478_0[1]),.dinb(w_n269_86[0]),.dout(n479),.clk(gclk));
	jor g0217(.dina(n479),.dinb(n477),.dout(n480),.clk(gclk));
	jor g0218(.dina(n480),.dinb(n475),.dout(n481),.clk(gclk));
	jand g0219(.dina(w_n481_1[1]),.dinb(w_n308_62[1]),.dout(n482),.clk(gclk));
	jor g0220(.dina(n482),.dinb(n470),.dout(n483),.clk(gclk));
	jor g0221(.dina(n483),.dinb(n458),.dout(n484),.clk(gclk));
	jand g0222(.dina(w_n376_0[0]),.dinb(w_n431_0[0]),.dout(n485),.clk(gclk));
	jand g0223(.dina(w_n485_63[1]),.dinb(w_n484_1[1]),.dout(n486),.clk(gclk));
	jor g0224(.dina(n486),.dinb(n433),.dout(n487),.clk(gclk));
	jor g0225(.dina(n487),.dinb(n379),.dout(n488),.clk(gclk));
	jand g0226(.dina(w_n488_0[1]),.dinb(w_n263_63[1]),.dout(n489),.clk(gclk));
	jand g0227(.dina(w_shift0_52[2]),.dinb(w_a15_0[1]),.dout(n490),.clk(gclk));
	jor g0228(.dina(w_n490_0[1]),.dinb(w_shift1_85[2]),.dout(n491),.clk(gclk));
	jand g0229(.dina(w_n270_52[2]),.dinb(w_a14_0[1]),.dout(n492),.clk(gclk));
	jor g0230(.dina(w_n492_0[1]),.dinb(w_n269_85[2]),.dout(n493),.clk(gclk));
	jand g0231(.dina(n493),.dinb(n491),.dout(n494),.clk(gclk));
	jand g0232(.dina(w_shift0_52[1]),.dinb(w_a13_0[1]),.dout(n495),.clk(gclk));
	jand g0233(.dina(w_n495_0[1]),.dinb(w_shift1_85[1]),.dout(n496),.clk(gclk));
	jand g0234(.dina(w_n270_52[1]),.dinb(w_a16_0[1]),.dout(n497),.clk(gclk));
	jand g0235(.dina(w_n497_0[1]),.dinb(w_n269_85[1]),.dout(n498),.clk(gclk));
	jor g0236(.dina(n498),.dinb(n496),.dout(n499),.clk(gclk));
	jor g0237(.dina(n499),.dinb(n494),.dout(n500),.clk(gclk));
	jand g0238(.dina(w_n500_1[1]),.dinb(w_n266_62[0]),.dout(n501),.clk(gclk));
	jand g0239(.dina(w_shift0_52[0]),.dinb(w_a7_0[1]),.dout(n502),.clk(gclk));
	jor g0240(.dina(w_n502_0[1]),.dinb(w_shift1_85[0]),.dout(n503),.clk(gclk));
	jand g0241(.dina(w_n270_52[0]),.dinb(w_a6_0[1]),.dout(n504),.clk(gclk));
	jor g0242(.dina(w_n504_0[1]),.dinb(w_n269_85[0]),.dout(n505),.clk(gclk));
	jand g0243(.dina(n505),.dinb(n503),.dout(n506),.clk(gclk));
	jand g0244(.dina(w_shift0_51[2]),.dinb(w_a5_0[1]),.dout(n507),.clk(gclk));
	jand g0245(.dina(w_n507_0[1]),.dinb(w_shift1_84[2]),.dout(n508),.clk(gclk));
	jand g0246(.dina(w_n270_51[2]),.dinb(w_a8_0[1]),.dout(n509),.clk(gclk));
	jand g0247(.dina(w_n509_0[1]),.dinb(w_n269_84[2]),.dout(n510),.clk(gclk));
	jor g0248(.dina(n510),.dinb(n508),.dout(n511),.clk(gclk));
	jor g0249(.dina(n511),.dinb(n506),.dout(n512),.clk(gclk));
	jand g0250(.dina(w_n512_1[1]),.dinb(w_n281_62[0]),.dout(n513),.clk(gclk));
	jor g0251(.dina(n513),.dinb(n501),.dout(n514),.clk(gclk));
	jand g0252(.dina(w_shift0_51[1]),.dinb(w_a11_0[1]),.dout(n515),.clk(gclk));
	jor g0253(.dina(w_n515_0[1]),.dinb(w_shift1_84[1]),.dout(n516),.clk(gclk));
	jand g0254(.dina(w_n270_51[1]),.dinb(w_a10_0[1]),.dout(n517),.clk(gclk));
	jor g0255(.dina(w_n517_0[1]),.dinb(w_n269_84[1]),.dout(n518),.clk(gclk));
	jand g0256(.dina(n518),.dinb(n516),.dout(n519),.clk(gclk));
	jand g0257(.dina(w_shift0_51[0]),.dinb(w_a9_0[1]),.dout(n520),.clk(gclk));
	jand g0258(.dina(w_n520_0[1]),.dinb(w_shift1_84[0]),.dout(n521),.clk(gclk));
	jand g0259(.dina(w_n270_51[0]),.dinb(w_a12_0[1]),.dout(n522),.clk(gclk));
	jand g0260(.dina(w_n522_0[1]),.dinb(w_n269_84[0]),.dout(n523),.clk(gclk));
	jor g0261(.dina(n523),.dinb(n521),.dout(n524),.clk(gclk));
	jor g0262(.dina(n524),.dinb(n519),.dout(n525),.clk(gclk));
	jand g0263(.dina(w_n525_1[1]),.dinb(w_n295_62[0]),.dout(n526),.clk(gclk));
	jand g0264(.dina(w_shift0_50[2]),.dinb(w_a3_0[1]),.dout(n527),.clk(gclk));
	jor g0265(.dina(w_n527_0[1]),.dinb(w_shift1_83[2]),.dout(n528),.clk(gclk));
	jand g0266(.dina(w_n270_50[2]),.dinb(w_a2_0[1]),.dout(n529),.clk(gclk));
	jor g0267(.dina(w_n529_0[1]),.dinb(w_n269_83[2]),.dout(n530),.clk(gclk));
	jand g0268(.dina(n530),.dinb(n528),.dout(n531),.clk(gclk));
	jand g0269(.dina(w_shift0_50[1]),.dinb(w_a1_0[1]),.dout(n532),.clk(gclk));
	jand g0270(.dina(w_n532_0[1]),.dinb(w_shift1_83[1]),.dout(n533),.clk(gclk));
	jand g0271(.dina(w_n270_50[1]),.dinb(w_a4_0[1]),.dout(n534),.clk(gclk));
	jand g0272(.dina(w_n534_0[1]),.dinb(w_n269_83[1]),.dout(n535),.clk(gclk));
	jor g0273(.dina(n535),.dinb(n533),.dout(n536),.clk(gclk));
	jor g0274(.dina(n536),.dinb(n531),.dout(n537),.clk(gclk));
	jand g0275(.dina(w_n537_1[1]),.dinb(w_n308_62[0]),.dout(n538),.clk(gclk));
	jor g0276(.dina(n538),.dinb(n526),.dout(n539),.clk(gclk));
	jor g0277(.dina(n539),.dinb(n514),.dout(n540),.clk(gclk));
	jand g0278(.dina(w_n540_1[1]),.dinb(w_n323_63[0]),.dout(n541),.clk(gclk));
	jand g0279(.dina(w_shift0_50[0]),.dinb(w_a47_0[1]),.dout(n542),.clk(gclk));
	jor g0280(.dina(w_n542_0[1]),.dinb(w_shift1_83[0]),.dout(n543),.clk(gclk));
	jand g0281(.dina(w_n270_50[0]),.dinb(w_a46_0[1]),.dout(n544),.clk(gclk));
	jor g0282(.dina(w_n544_0[1]),.dinb(w_n269_83[0]),.dout(n545),.clk(gclk));
	jand g0283(.dina(n545),.dinb(n543),.dout(n546),.clk(gclk));
	jand g0284(.dina(w_shift0_49[2]),.dinb(w_a45_0[1]),.dout(n547),.clk(gclk));
	jand g0285(.dina(w_n547_0[1]),.dinb(w_shift1_82[2]),.dout(n548),.clk(gclk));
	jand g0286(.dina(w_n270_49[2]),.dinb(w_a48_0[1]),.dout(n549),.clk(gclk));
	jand g0287(.dina(w_n549_0[1]),.dinb(w_n269_82[2]),.dout(n550),.clk(gclk));
	jor g0288(.dina(n550),.dinb(n548),.dout(n551),.clk(gclk));
	jor g0289(.dina(n551),.dinb(n546),.dout(n552),.clk(gclk));
	jand g0290(.dina(w_n552_1[1]),.dinb(w_n266_61[2]),.dout(n553),.clk(gclk));
	jand g0291(.dina(w_n270_49[1]),.dinb(w_a40_0[1]),.dout(n554),.clk(gclk));
	jand g0292(.dina(w_shift0_49[1]),.dinb(w_a39_0[1]),.dout(n555),.clk(gclk));
	jor g0293(.dina(w_n555_0[1]),.dinb(w_n554_0[1]),.dout(n556),.clk(gclk));
	jand g0294(.dina(n556),.dinb(w_n269_82[1]),.dout(n557),.clk(gclk));
	jand g0295(.dina(w_n270_49[0]),.dinb(w_a38_0[1]),.dout(n558),.clk(gclk));
	jand g0296(.dina(w_shift0_49[0]),.dinb(w_a37_0[1]),.dout(n559),.clk(gclk));
	jor g0297(.dina(w_n559_0[1]),.dinb(w_n558_0[1]),.dout(n560),.clk(gclk));
	jand g0298(.dina(n560),.dinb(w_shift1_82[1]),.dout(n561),.clk(gclk));
	jor g0299(.dina(n561),.dinb(n557),.dout(n562),.clk(gclk));
	jand g0300(.dina(w_n562_1[1]),.dinb(w_n281_61[2]),.dout(n563),.clk(gclk));
	jor g0301(.dina(n563),.dinb(n553),.dout(n564),.clk(gclk));
	jand g0302(.dina(w_shift0_48[2]),.dinb(w_a43_0[1]),.dout(n565),.clk(gclk));
	jor g0303(.dina(w_n565_0[1]),.dinb(w_shift1_82[0]),.dout(n566),.clk(gclk));
	jand g0304(.dina(w_n270_48[2]),.dinb(w_a42_0[1]),.dout(n567),.clk(gclk));
	jor g0305(.dina(w_n567_0[1]),.dinb(w_n269_82[0]),.dout(n568),.clk(gclk));
	jand g0306(.dina(n568),.dinb(n566),.dout(n569),.clk(gclk));
	jand g0307(.dina(w_shift0_48[1]),.dinb(w_a41_0[1]),.dout(n570),.clk(gclk));
	jand g0308(.dina(w_n570_0[1]),.dinb(w_shift1_81[2]),.dout(n571),.clk(gclk));
	jand g0309(.dina(w_n270_48[1]),.dinb(w_a44_0[1]),.dout(n572),.clk(gclk));
	jand g0310(.dina(w_n572_0[1]),.dinb(w_n269_81[2]),.dout(n573),.clk(gclk));
	jor g0311(.dina(n573),.dinb(n571),.dout(n574),.clk(gclk));
	jor g0312(.dina(n574),.dinb(n569),.dout(n575),.clk(gclk));
	jand g0313(.dina(w_n575_1[1]),.dinb(w_n295_61[2]),.dout(n576),.clk(gclk));
	jand g0314(.dina(w_shift0_48[0]),.dinb(w_a35_0[1]),.dout(n577),.clk(gclk));
	jor g0315(.dina(w_n577_0[1]),.dinb(w_shift1_81[1]),.dout(n578),.clk(gclk));
	jand g0316(.dina(w_n270_48[0]),.dinb(w_a34_0[1]),.dout(n579),.clk(gclk));
	jor g0317(.dina(w_n579_0[1]),.dinb(w_n269_81[1]),.dout(n580),.clk(gclk));
	jand g0318(.dina(n580),.dinb(n578),.dout(n581),.clk(gclk));
	jand g0319(.dina(w_shift0_47[2]),.dinb(w_a33_0[1]),.dout(n582),.clk(gclk));
	jand g0320(.dina(w_n582_0[1]),.dinb(w_shift1_81[0]),.dout(n583),.clk(gclk));
	jand g0321(.dina(w_n270_47[2]),.dinb(w_a36_0[1]),.dout(n584),.clk(gclk));
	jand g0322(.dina(w_n584_0[1]),.dinb(w_n269_81[0]),.dout(n585),.clk(gclk));
	jor g0323(.dina(n585),.dinb(n583),.dout(n586),.clk(gclk));
	jor g0324(.dina(n586),.dinb(n581),.dout(n587),.clk(gclk));
	jand g0325(.dina(w_n587_1[1]),.dinb(w_n308_61[2]),.dout(n588),.clk(gclk));
	jor g0326(.dina(n588),.dinb(n576),.dout(n589),.clk(gclk));
	jor g0327(.dina(n589),.dinb(n564),.dout(n590),.clk(gclk));
	jand g0328(.dina(w_n590_1[1]),.dinb(w_n377_63[0]),.dout(n591),.clk(gclk));
	jor g0329(.dina(n591),.dinb(n541),.dout(n592),.clk(gclk));
	jand g0330(.dina(w_shift0_47[1]),.dinb(w_a31_0[1]),.dout(n593),.clk(gclk));
	jor g0331(.dina(w_n593_0[1]),.dinb(w_shift1_80[2]),.dout(n594),.clk(gclk));
	jand g0332(.dina(w_n270_47[1]),.dinb(w_a30_0[1]),.dout(n595),.clk(gclk));
	jor g0333(.dina(w_n595_0[1]),.dinb(w_n269_80[2]),.dout(n596),.clk(gclk));
	jand g0334(.dina(n596),.dinb(n594),.dout(n597),.clk(gclk));
	jand g0335(.dina(w_shift0_47[0]),.dinb(w_a29_0[1]),.dout(n598),.clk(gclk));
	jand g0336(.dina(w_n598_0[1]),.dinb(w_shift1_80[1]),.dout(n599),.clk(gclk));
	jand g0337(.dina(w_n270_47[0]),.dinb(w_a32_0[1]),.dout(n600),.clk(gclk));
	jand g0338(.dina(w_n600_0[1]),.dinb(w_n269_80[1]),.dout(n601),.clk(gclk));
	jor g0339(.dina(n601),.dinb(n599),.dout(n602),.clk(gclk));
	jor g0340(.dina(n602),.dinb(n597),.dout(n603),.clk(gclk));
	jand g0341(.dina(w_n603_1[1]),.dinb(w_n266_61[1]),.dout(n604),.clk(gclk));
	jand g0342(.dina(w_shift0_46[2]),.dinb(w_a23_0[1]),.dout(n605),.clk(gclk));
	jor g0343(.dina(w_n605_0[1]),.dinb(w_shift1_80[0]),.dout(n606),.clk(gclk));
	jand g0344(.dina(w_n270_46[2]),.dinb(w_a22_0[1]),.dout(n607),.clk(gclk));
	jor g0345(.dina(w_n607_0[1]),.dinb(w_n269_80[0]),.dout(n608),.clk(gclk));
	jand g0346(.dina(n608),.dinb(n606),.dout(n609),.clk(gclk));
	jand g0347(.dina(w_shift0_46[1]),.dinb(w_a21_0[1]),.dout(n610),.clk(gclk));
	jand g0348(.dina(w_n610_0[1]),.dinb(w_shift1_79[2]),.dout(n611),.clk(gclk));
	jand g0349(.dina(w_n270_46[1]),.dinb(w_a24_0[1]),.dout(n612),.clk(gclk));
	jand g0350(.dina(w_n612_0[1]),.dinb(w_n269_79[2]),.dout(n613),.clk(gclk));
	jor g0351(.dina(n613),.dinb(n611),.dout(n614),.clk(gclk));
	jor g0352(.dina(n614),.dinb(n609),.dout(n615),.clk(gclk));
	jand g0353(.dina(w_n615_1[1]),.dinb(w_n281_61[1]),.dout(n616),.clk(gclk));
	jor g0354(.dina(n616),.dinb(n604),.dout(n617),.clk(gclk));
	jand g0355(.dina(w_shift0_46[0]),.dinb(w_a27_0[1]),.dout(n618),.clk(gclk));
	jor g0356(.dina(w_n618_0[1]),.dinb(w_shift1_79[1]),.dout(n619),.clk(gclk));
	jand g0357(.dina(w_n270_46[0]),.dinb(w_a26_0[1]),.dout(n620),.clk(gclk));
	jor g0358(.dina(w_n620_0[1]),.dinb(w_n269_79[1]),.dout(n621),.clk(gclk));
	jand g0359(.dina(n621),.dinb(n619),.dout(n622),.clk(gclk));
	jand g0360(.dina(w_shift0_45[2]),.dinb(w_a25_0[1]),.dout(n623),.clk(gclk));
	jand g0361(.dina(w_n623_0[1]),.dinb(w_shift1_79[0]),.dout(n624),.clk(gclk));
	jand g0362(.dina(w_n270_45[2]),.dinb(w_a28_0[1]),.dout(n625),.clk(gclk));
	jand g0363(.dina(w_n625_0[1]),.dinb(w_n269_79[0]),.dout(n626),.clk(gclk));
	jor g0364(.dina(n626),.dinb(n624),.dout(n627),.clk(gclk));
	jor g0365(.dina(n627),.dinb(n622),.dout(n628),.clk(gclk));
	jand g0366(.dina(w_n628_1[1]),.dinb(w_n295_61[1]),.dout(n629),.clk(gclk));
	jand g0367(.dina(w_shift0_45[1]),.dinb(w_a19_0[1]),.dout(n630),.clk(gclk));
	jor g0368(.dina(w_n630_0[1]),.dinb(w_shift1_78[2]),.dout(n631),.clk(gclk));
	jand g0369(.dina(w_n270_45[1]),.dinb(w_a18_0[1]),.dout(n632),.clk(gclk));
	jor g0370(.dina(w_n632_0[1]),.dinb(w_n269_78[2]),.dout(n633),.clk(gclk));
	jand g0371(.dina(n633),.dinb(n631),.dout(n634),.clk(gclk));
	jand g0372(.dina(w_shift0_45[0]),.dinb(w_a17_0[1]),.dout(n635),.clk(gclk));
	jand g0373(.dina(w_n635_0[1]),.dinb(w_shift1_78[1]),.dout(n636),.clk(gclk));
	jand g0374(.dina(w_n270_45[0]),.dinb(w_a20_0[1]),.dout(n637),.clk(gclk));
	jand g0375(.dina(w_n637_0[1]),.dinb(w_n269_78[1]),.dout(n638),.clk(gclk));
	jor g0376(.dina(n638),.dinb(n636),.dout(n639),.clk(gclk));
	jor g0377(.dina(n639),.dinb(n634),.dout(n640),.clk(gclk));
	jand g0378(.dina(w_n640_1[1]),.dinb(w_n308_61[1]),.dout(n641),.clk(gclk));
	jor g0379(.dina(n641),.dinb(n629),.dout(n642),.clk(gclk));
	jor g0380(.dina(n642),.dinb(n617),.dout(n643),.clk(gclk));
	jand g0381(.dina(w_n643_1[1]),.dinb(w_n432_63[0]),.dout(n644),.clk(gclk));
	jand g0382(.dina(w_shift0_44[2]),.dinb(w_a63_0[1]),.dout(n645),.clk(gclk));
	jor g0383(.dina(w_n645_0[1]),.dinb(w_shift1_78[0]),.dout(n646),.clk(gclk));
	jand g0384(.dina(w_n270_44[2]),.dinb(w_a62_0[1]),.dout(n647),.clk(gclk));
	jor g0385(.dina(w_n647_0[1]),.dinb(w_n269_78[0]),.dout(n648),.clk(gclk));
	jand g0386(.dina(n648),.dinb(n646),.dout(n649),.clk(gclk));
	jand g0387(.dina(w_shift0_44[1]),.dinb(w_a61_0[1]),.dout(n650),.clk(gclk));
	jand g0388(.dina(w_n650_0[1]),.dinb(w_shift1_77[2]),.dout(n651),.clk(gclk));
	jand g0389(.dina(w_n270_44[1]),.dinb(w_a64_0[1]),.dout(n652),.clk(gclk));
	jand g0390(.dina(w_n652_0[1]),.dinb(w_n269_77[2]),.dout(n653),.clk(gclk));
	jor g0391(.dina(n653),.dinb(n651),.dout(n654),.clk(gclk));
	jor g0392(.dina(n654),.dinb(n649),.dout(n655),.clk(gclk));
	jand g0393(.dina(w_n655_1[1]),.dinb(w_n266_61[0]),.dout(n656),.clk(gclk));
	jand g0394(.dina(w_shift0_44[0]),.dinb(w_a55_0[1]),.dout(n657),.clk(gclk));
	jor g0395(.dina(w_n657_0[1]),.dinb(w_shift1_77[1]),.dout(n658),.clk(gclk));
	jand g0396(.dina(w_n270_44[0]),.dinb(w_a54_0[1]),.dout(n659),.clk(gclk));
	jor g0397(.dina(w_n659_0[1]),.dinb(w_n269_77[1]),.dout(n660),.clk(gclk));
	jand g0398(.dina(n660),.dinb(n658),.dout(n661),.clk(gclk));
	jand g0399(.dina(w_shift0_43[2]),.dinb(w_a53_0[1]),.dout(n662),.clk(gclk));
	jand g0400(.dina(w_n662_0[1]),.dinb(w_shift1_77[0]),.dout(n663),.clk(gclk));
	jand g0401(.dina(w_n270_43[2]),.dinb(w_a56_0[1]),.dout(n664),.clk(gclk));
	jand g0402(.dina(w_n664_0[1]),.dinb(w_n269_77[0]),.dout(n665),.clk(gclk));
	jor g0403(.dina(n665),.dinb(n663),.dout(n666),.clk(gclk));
	jor g0404(.dina(n666),.dinb(n661),.dout(n667),.clk(gclk));
	jand g0405(.dina(w_n667_1[1]),.dinb(w_n281_61[0]),.dout(n668),.clk(gclk));
	jor g0406(.dina(n668),.dinb(n656),.dout(n669),.clk(gclk));
	jand g0407(.dina(w_shift0_43[1]),.dinb(w_a59_0[1]),.dout(n670),.clk(gclk));
	jor g0408(.dina(w_n670_0[1]),.dinb(w_shift1_76[2]),.dout(n671),.clk(gclk));
	jand g0409(.dina(w_n270_43[1]),.dinb(w_a58_0[1]),.dout(n672),.clk(gclk));
	jor g0410(.dina(w_n672_0[1]),.dinb(w_n269_76[2]),.dout(n673),.clk(gclk));
	jand g0411(.dina(n673),.dinb(n671),.dout(n674),.clk(gclk));
	jand g0412(.dina(w_shift0_43[0]),.dinb(w_a57_0[1]),.dout(n675),.clk(gclk));
	jand g0413(.dina(w_n675_0[1]),.dinb(w_shift1_76[1]),.dout(n676),.clk(gclk));
	jand g0414(.dina(w_n270_43[0]),.dinb(w_a60_0[1]),.dout(n677),.clk(gclk));
	jand g0415(.dina(w_n677_0[1]),.dinb(w_n269_76[1]),.dout(n678),.clk(gclk));
	jor g0416(.dina(n678),.dinb(n676),.dout(n679),.clk(gclk));
	jor g0417(.dina(n679),.dinb(n674),.dout(n680),.clk(gclk));
	jand g0418(.dina(w_n680_1[1]),.dinb(w_n295_61[0]),.dout(n681),.clk(gclk));
	jand g0419(.dina(w_shift0_42[2]),.dinb(w_a51_0[1]),.dout(n682),.clk(gclk));
	jor g0420(.dina(w_n682_0[1]),.dinb(w_shift1_76[0]),.dout(n683),.clk(gclk));
	jand g0421(.dina(w_n270_42[2]),.dinb(w_a50_0[1]),.dout(n684),.clk(gclk));
	jor g0422(.dina(w_n684_0[1]),.dinb(w_n269_76[0]),.dout(n685),.clk(gclk));
	jand g0423(.dina(n685),.dinb(n683),.dout(n686),.clk(gclk));
	jand g0424(.dina(w_shift0_42[1]),.dinb(w_a49_0[1]),.dout(n687),.clk(gclk));
	jand g0425(.dina(w_n687_0[1]),.dinb(w_shift1_75[2]),.dout(n688),.clk(gclk));
	jand g0426(.dina(w_n270_42[1]),.dinb(w_a52_0[1]),.dout(n689),.clk(gclk));
	jand g0427(.dina(w_n689_0[1]),.dinb(w_n269_75[2]),.dout(n690),.clk(gclk));
	jor g0428(.dina(n690),.dinb(n688),.dout(n691),.clk(gclk));
	jor g0429(.dina(n691),.dinb(n686),.dout(n692),.clk(gclk));
	jand g0430(.dina(w_n692_1[1]),.dinb(w_n308_61[0]),.dout(n693),.clk(gclk));
	jor g0431(.dina(n693),.dinb(n681),.dout(n694),.clk(gclk));
	jor g0432(.dina(n694),.dinb(n669),.dout(n695),.clk(gclk));
	jand g0433(.dina(w_n695_1[1]),.dinb(w_n485_63[0]),.dout(n696),.clk(gclk));
	jor g0434(.dina(n696),.dinb(n644),.dout(n697),.clk(gclk));
	jor g0435(.dina(n697),.dinb(n592),.dout(n698),.clk(gclk));
	jand g0436(.dina(w_n698_0[1]),.dinb(w_shift6_63[1]),.dout(n699),.clk(gclk));
	jor g0437(.dina(n699),.dinb(n489),.dout(result0),.clk(gclk));
	jor g0438(.dina(w_n270_42[0]),.dinb(w_a78_0[0]),.dout(n701),.clk(gclk));
	jor g0439(.dina(w_shift0_42[0]),.dinb(w_a79_0[0]),.dout(n702),.clk(gclk));
	jand g0440(.dina(n702),.dinb(n701),.dout(n703),.clk(gclk));
	jor g0441(.dina(w_n703_0[1]),.dinb(w_n269_75[1]),.dout(n704),.clk(gclk));
	jor g0442(.dina(w_n270_41[2]),.dinb(w_a80_0[0]),.dout(n705),.clk(gclk));
	jor g0443(.dina(w_shift0_41[2]),.dinb(w_a81_0[0]),.dout(n706),.clk(gclk));
	jand g0444(.dina(n706),.dinb(n705),.dout(n707),.clk(gclk));
	jor g0445(.dina(w_n707_0[1]),.dinb(w_shift1_75[1]),.dout(n708),.clk(gclk));
	jand g0446(.dina(n708),.dinb(n704),.dout(n709),.clk(gclk));
	jand g0447(.dina(w_n709_1[1]),.dinb(w_n266_60[2]),.dout(n710),.clk(gclk));
	jor g0448(.dina(w_n270_41[1]),.dinb(w_a70_0[0]),.dout(n711),.clk(gclk));
	jor g0449(.dina(w_shift0_41[1]),.dinb(w_a71_0[0]),.dout(n712),.clk(gclk));
	jand g0450(.dina(n712),.dinb(n711),.dout(n713),.clk(gclk));
	jor g0451(.dina(w_n713_0[1]),.dinb(w_n269_75[0]),.dout(n714),.clk(gclk));
	jor g0452(.dina(w_n270_41[0]),.dinb(w_a72_0[0]),.dout(n715),.clk(gclk));
	jor g0453(.dina(w_shift0_41[0]),.dinb(w_a73_0[0]),.dout(n716),.clk(gclk));
	jand g0454(.dina(n716),.dinb(n715),.dout(n717),.clk(gclk));
	jor g0455(.dina(w_n717_0[1]),.dinb(w_shift1_75[0]),.dout(n718),.clk(gclk));
	jand g0456(.dina(n718),.dinb(n714),.dout(n719),.clk(gclk));
	jand g0457(.dina(w_n719_1[1]),.dinb(w_n281_60[2]),.dout(n720),.clk(gclk));
	jor g0458(.dina(n720),.dinb(n710),.dout(n721),.clk(gclk));
	jor g0459(.dina(w_n270_40[2]),.dinb(w_a74_0[0]),.dout(n722),.clk(gclk));
	jor g0460(.dina(w_shift0_40[2]),.dinb(w_a75_0[0]),.dout(n723),.clk(gclk));
	jand g0461(.dina(n723),.dinb(n722),.dout(n724),.clk(gclk));
	jor g0462(.dina(w_n724_0[1]),.dinb(w_n269_74[2]),.dout(n725),.clk(gclk));
	jor g0463(.dina(w_n270_40[1]),.dinb(w_a76_0[0]),.dout(n726),.clk(gclk));
	jor g0464(.dina(w_shift0_40[1]),.dinb(w_a77_0[0]),.dout(n727),.clk(gclk));
	jand g0465(.dina(n727),.dinb(n726),.dout(n728),.clk(gclk));
	jor g0466(.dina(w_n728_0[1]),.dinb(w_shift1_74[2]),.dout(n729),.clk(gclk));
	jand g0467(.dina(n729),.dinb(n725),.dout(n730),.clk(gclk));
	jand g0468(.dina(w_n730_1[1]),.dinb(w_n295_60[2]),.dout(n731),.clk(gclk));
	jor g0469(.dina(w_n270_40[0]),.dinb(w_a66_0[0]),.dout(n732),.clk(gclk));
	jor g0470(.dina(w_shift0_40[0]),.dinb(w_a67_0[0]),.dout(n733),.clk(gclk));
	jand g0471(.dina(n733),.dinb(n732),.dout(n734),.clk(gclk));
	jor g0472(.dina(w_n734_0[1]),.dinb(w_n269_74[1]),.dout(n735),.clk(gclk));
	jor g0473(.dina(w_n270_39[2]),.dinb(w_a68_0[0]),.dout(n736),.clk(gclk));
	jor g0474(.dina(w_shift0_39[2]),.dinb(w_a69_0[0]),.dout(n737),.clk(gclk));
	jand g0475(.dina(n737),.dinb(n736),.dout(n738),.clk(gclk));
	jor g0476(.dina(w_n738_0[1]),.dinb(w_shift1_74[1]),.dout(n739),.clk(gclk));
	jand g0477(.dina(n739),.dinb(n735),.dout(n740),.clk(gclk));
	jand g0478(.dina(w_n740_1[1]),.dinb(w_n308_60[2]),.dout(n741),.clk(gclk));
	jor g0479(.dina(n741),.dinb(n731),.dout(n742),.clk(gclk));
	jor g0480(.dina(n742),.dinb(n721),.dout(n743),.clk(gclk));
	jand g0481(.dina(w_n743_1[1]),.dinb(w_n323_62[2]),.dout(n744),.clk(gclk));
	jor g0482(.dina(w_n270_39[1]),.dinb(w_a110_0[0]),.dout(n745),.clk(gclk));
	jor g0483(.dina(w_shift0_39[1]),.dinb(w_a111_0[0]),.dout(n746),.clk(gclk));
	jand g0484(.dina(n746),.dinb(n745),.dout(n747),.clk(gclk));
	jor g0485(.dina(w_n747_0[1]),.dinb(w_n269_74[0]),.dout(n748),.clk(gclk));
	jor g0486(.dina(w_n270_39[0]),.dinb(w_a112_0[0]),.dout(n749),.clk(gclk));
	jor g0487(.dina(w_shift0_39[0]),.dinb(w_a113_0[0]),.dout(n750),.clk(gclk));
	jand g0488(.dina(n750),.dinb(n749),.dout(n751),.clk(gclk));
	jor g0489(.dina(w_n751_0[1]),.dinb(w_shift1_74[0]),.dout(n752),.clk(gclk));
	jand g0490(.dina(n752),.dinb(n748),.dout(n753),.clk(gclk));
	jand g0491(.dina(w_n753_1[1]),.dinb(w_n266_60[1]),.dout(n754),.clk(gclk));
	jor g0492(.dina(w_n270_38[2]),.dinb(w_a102_0[0]),.dout(n755),.clk(gclk));
	jor g0493(.dina(w_shift0_38[2]),.dinb(w_a103_0[0]),.dout(n756),.clk(gclk));
	jand g0494(.dina(n756),.dinb(n755),.dout(n757),.clk(gclk));
	jor g0495(.dina(w_n757_0[1]),.dinb(w_n269_73[2]),.dout(n758),.clk(gclk));
	jor g0496(.dina(w_n270_38[1]),.dinb(w_a104_0[0]),.dout(n759),.clk(gclk));
	jor g0497(.dina(w_shift0_38[1]),.dinb(w_a105_0[0]),.dout(n760),.clk(gclk));
	jand g0498(.dina(n760),.dinb(n759),.dout(n761),.clk(gclk));
	jor g0499(.dina(w_n761_0[1]),.dinb(w_shift1_73[2]),.dout(n762),.clk(gclk));
	jand g0500(.dina(n762),.dinb(n758),.dout(n763),.clk(gclk));
	jand g0501(.dina(w_n763_1[1]),.dinb(w_n281_60[1]),.dout(n764),.clk(gclk));
	jor g0502(.dina(n764),.dinb(n754),.dout(n765),.clk(gclk));
	jor g0503(.dina(w_n270_38[0]),.dinb(w_a106_0[0]),.dout(n766),.clk(gclk));
	jor g0504(.dina(w_shift0_38[0]),.dinb(w_a107_0[0]),.dout(n767),.clk(gclk));
	jand g0505(.dina(n767),.dinb(n766),.dout(n768),.clk(gclk));
	jor g0506(.dina(w_n768_0[1]),.dinb(w_n269_73[1]),.dout(n769),.clk(gclk));
	jor g0507(.dina(w_n270_37[2]),.dinb(w_a108_0[0]),.dout(n770),.clk(gclk));
	jor g0508(.dina(w_shift0_37[2]),.dinb(w_a109_0[0]),.dout(n771),.clk(gclk));
	jand g0509(.dina(n771),.dinb(n770),.dout(n772),.clk(gclk));
	jor g0510(.dina(w_n772_0[1]),.dinb(w_shift1_73[1]),.dout(n773),.clk(gclk));
	jand g0511(.dina(n773),.dinb(n769),.dout(n774),.clk(gclk));
	jand g0512(.dina(w_n774_1[1]),.dinb(w_n295_60[1]),.dout(n775),.clk(gclk));
	jor g0513(.dina(w_n270_37[1]),.dinb(w_a98_0[0]),.dout(n776),.clk(gclk));
	jor g0514(.dina(w_shift0_37[1]),.dinb(w_a99_0[0]),.dout(n777),.clk(gclk));
	jand g0515(.dina(n777),.dinb(n776),.dout(n778),.clk(gclk));
	jor g0516(.dina(w_n778_0[1]),.dinb(w_n269_73[0]),.dout(n779),.clk(gclk));
	jor g0517(.dina(w_n270_37[0]),.dinb(w_a100_0[0]),.dout(n780),.clk(gclk));
	jor g0518(.dina(w_shift0_37[0]),.dinb(w_a101_0[0]),.dout(n781),.clk(gclk));
	jand g0519(.dina(n781),.dinb(n780),.dout(n782),.clk(gclk));
	jor g0520(.dina(w_n782_0[1]),.dinb(w_shift1_73[0]),.dout(n783),.clk(gclk));
	jand g0521(.dina(n783),.dinb(n779),.dout(n784),.clk(gclk));
	jand g0522(.dina(w_n784_1[1]),.dinb(w_n308_60[1]),.dout(n785),.clk(gclk));
	jor g0523(.dina(n785),.dinb(n775),.dout(n786),.clk(gclk));
	jor g0524(.dina(n786),.dinb(n765),.dout(n787),.clk(gclk));
	jand g0525(.dina(w_n787_1[1]),.dinb(w_n377_62[2]),.dout(n788),.clk(gclk));
	jor g0526(.dina(n788),.dinb(n744),.dout(n789),.clk(gclk));
	jor g0527(.dina(w_n270_36[2]),.dinb(w_a94_0[0]),.dout(n790),.clk(gclk));
	jor g0528(.dina(w_shift0_36[2]),.dinb(w_a95_0[0]),.dout(n791),.clk(gclk));
	jand g0529(.dina(n791),.dinb(n790),.dout(n792),.clk(gclk));
	jor g0530(.dina(w_n792_0[1]),.dinb(w_n269_72[2]),.dout(n793),.clk(gclk));
	jor g0531(.dina(w_n270_36[1]),.dinb(w_a96_0[0]),.dout(n794),.clk(gclk));
	jor g0532(.dina(w_shift0_36[1]),.dinb(w_a97_0[0]),.dout(n795),.clk(gclk));
	jand g0533(.dina(n795),.dinb(n794),.dout(n796),.clk(gclk));
	jor g0534(.dina(w_n796_0[1]),.dinb(w_shift1_72[2]),.dout(n797),.clk(gclk));
	jand g0535(.dina(n797),.dinb(n793),.dout(n798),.clk(gclk));
	jand g0536(.dina(w_n798_1[1]),.dinb(w_n266_60[0]),.dout(n799),.clk(gclk));
	jor g0537(.dina(w_n270_36[0]),.dinb(w_a86_0[0]),.dout(n800),.clk(gclk));
	jor g0538(.dina(w_shift0_36[0]),.dinb(w_a87_0[0]),.dout(n801),.clk(gclk));
	jand g0539(.dina(n801),.dinb(n800),.dout(n802),.clk(gclk));
	jor g0540(.dina(w_n802_0[1]),.dinb(w_n269_72[1]),.dout(n803),.clk(gclk));
	jor g0541(.dina(w_n270_35[2]),.dinb(w_a88_0[0]),.dout(n804),.clk(gclk));
	jor g0542(.dina(w_shift0_35[2]),.dinb(w_a89_0[0]),.dout(n805),.clk(gclk));
	jand g0543(.dina(n805),.dinb(n804),.dout(n806),.clk(gclk));
	jor g0544(.dina(w_n806_0[1]),.dinb(w_shift1_72[1]),.dout(n807),.clk(gclk));
	jand g0545(.dina(n807),.dinb(n803),.dout(n808),.clk(gclk));
	jand g0546(.dina(w_n808_1[1]),.dinb(w_n281_60[0]),.dout(n809),.clk(gclk));
	jor g0547(.dina(n809),.dinb(n799),.dout(n810),.clk(gclk));
	jor g0548(.dina(w_n270_35[1]),.dinb(w_a90_0[0]),.dout(n811),.clk(gclk));
	jor g0549(.dina(w_shift0_35[1]),.dinb(w_a91_0[0]),.dout(n812),.clk(gclk));
	jand g0550(.dina(n812),.dinb(n811),.dout(n813),.clk(gclk));
	jor g0551(.dina(w_n813_0[1]),.dinb(w_n269_72[0]),.dout(n814),.clk(gclk));
	jor g0552(.dina(w_n270_35[0]),.dinb(w_a92_0[0]),.dout(n815),.clk(gclk));
	jor g0553(.dina(w_shift0_35[0]),.dinb(w_a93_0[0]),.dout(n816),.clk(gclk));
	jand g0554(.dina(n816),.dinb(n815),.dout(n817),.clk(gclk));
	jor g0555(.dina(w_n817_0[1]),.dinb(w_shift1_72[0]),.dout(n818),.clk(gclk));
	jand g0556(.dina(n818),.dinb(n814),.dout(n819),.clk(gclk));
	jand g0557(.dina(w_n819_1[1]),.dinb(w_n295_60[0]),.dout(n820),.clk(gclk));
	jor g0558(.dina(w_n270_34[2]),.dinb(w_a82_0[0]),.dout(n821),.clk(gclk));
	jor g0559(.dina(w_shift0_34[2]),.dinb(w_a83_0[0]),.dout(n822),.clk(gclk));
	jand g0560(.dina(n822),.dinb(n821),.dout(n823),.clk(gclk));
	jor g0561(.dina(w_n823_0[1]),.dinb(w_n269_71[2]),.dout(n824),.clk(gclk));
	jor g0562(.dina(w_n270_34[1]),.dinb(w_a84_0[0]),.dout(n825),.clk(gclk));
	jor g0563(.dina(w_shift0_34[1]),.dinb(w_a85_0[0]),.dout(n826),.clk(gclk));
	jand g0564(.dina(n826),.dinb(n825),.dout(n827),.clk(gclk));
	jor g0565(.dina(w_n827_0[1]),.dinb(w_shift1_71[2]),.dout(n828),.clk(gclk));
	jand g0566(.dina(n828),.dinb(n824),.dout(n829),.clk(gclk));
	jand g0567(.dina(w_n829_1[1]),.dinb(w_n308_60[0]),.dout(n830),.clk(gclk));
	jor g0568(.dina(n830),.dinb(n820),.dout(n831),.clk(gclk));
	jor g0569(.dina(n831),.dinb(n810),.dout(n832),.clk(gclk));
	jand g0570(.dina(w_n832_1[1]),.dinb(w_n432_62[2]),.dout(n833),.clk(gclk));
	jor g0571(.dina(w_n270_34[0]),.dinb(w_a126_0[0]),.dout(n834),.clk(gclk));
	jor g0572(.dina(w_shift0_34[0]),.dinb(w_a127_0[0]),.dout(n835),.clk(gclk));
	jand g0573(.dina(n835),.dinb(n834),.dout(n836),.clk(gclk));
	jor g0574(.dina(w_n836_0[1]),.dinb(w_n269_71[1]),.dout(n837),.clk(gclk));
	jor g0575(.dina(w_n270_33[2]),.dinb(w_a0_0[0]),.dout(n838),.clk(gclk));
	jor g0576(.dina(w_shift0_33[2]),.dinb(w_a1_0[0]),.dout(n839),.clk(gclk));
	jand g0577(.dina(n839),.dinb(n838),.dout(n840),.clk(gclk));
	jor g0578(.dina(w_n840_0[1]),.dinb(w_shift1_71[1]),.dout(n841),.clk(gclk));
	jand g0579(.dina(n841),.dinb(n837),.dout(n842),.clk(gclk));
	jand g0580(.dina(w_n842_1[1]),.dinb(w_n266_59[2]),.dout(n843),.clk(gclk));
	jor g0581(.dina(w_n270_33[1]),.dinb(w_a118_0[0]),.dout(n844),.clk(gclk));
	jor g0582(.dina(w_shift0_33[1]),.dinb(w_a119_0[0]),.dout(n845),.clk(gclk));
	jand g0583(.dina(n845),.dinb(n844),.dout(n846),.clk(gclk));
	jor g0584(.dina(w_n846_0[1]),.dinb(w_n269_71[0]),.dout(n847),.clk(gclk));
	jor g0585(.dina(w_n270_33[0]),.dinb(w_a120_0[0]),.dout(n848),.clk(gclk));
	jor g0586(.dina(w_shift0_33[0]),.dinb(w_a121_0[0]),.dout(n849),.clk(gclk));
	jand g0587(.dina(n849),.dinb(n848),.dout(n850),.clk(gclk));
	jor g0588(.dina(w_n850_0[1]),.dinb(w_shift1_71[0]),.dout(n851),.clk(gclk));
	jand g0589(.dina(n851),.dinb(n847),.dout(n852),.clk(gclk));
	jand g0590(.dina(w_n852_1[1]),.dinb(w_n281_59[2]),.dout(n853),.clk(gclk));
	jor g0591(.dina(n853),.dinb(n843),.dout(n854),.clk(gclk));
	jor g0592(.dina(w_n270_32[2]),.dinb(w_a122_0[0]),.dout(n855),.clk(gclk));
	jor g0593(.dina(w_shift0_32[2]),.dinb(w_a123_0[0]),.dout(n856),.clk(gclk));
	jand g0594(.dina(n856),.dinb(n855),.dout(n857),.clk(gclk));
	jor g0595(.dina(w_n857_0[1]),.dinb(w_n269_70[2]),.dout(n858),.clk(gclk));
	jor g0596(.dina(w_n270_32[1]),.dinb(w_a124_0[0]),.dout(n859),.clk(gclk));
	jor g0597(.dina(w_shift0_32[1]),.dinb(w_a125_0[0]),.dout(n860),.clk(gclk));
	jand g0598(.dina(n860),.dinb(n859),.dout(n861),.clk(gclk));
	jor g0599(.dina(w_n861_0[1]),.dinb(w_shift1_70[2]),.dout(n862),.clk(gclk));
	jand g0600(.dina(n862),.dinb(n858),.dout(n863),.clk(gclk));
	jand g0601(.dina(w_n863_1[1]),.dinb(w_n295_59[2]),.dout(n864),.clk(gclk));
	jor g0602(.dina(w_n270_32[0]),.dinb(w_a114_0[0]),.dout(n865),.clk(gclk));
	jor g0603(.dina(w_shift0_32[0]),.dinb(w_a115_0[0]),.dout(n866),.clk(gclk));
	jand g0604(.dina(n866),.dinb(n865),.dout(n867),.clk(gclk));
	jor g0605(.dina(w_n867_0[1]),.dinb(w_n269_70[1]),.dout(n868),.clk(gclk));
	jor g0606(.dina(w_n270_31[2]),.dinb(w_a116_0[0]),.dout(n869),.clk(gclk));
	jor g0607(.dina(w_shift0_31[2]),.dinb(w_a117_0[0]),.dout(n870),.clk(gclk));
	jand g0608(.dina(n870),.dinb(n869),.dout(n871),.clk(gclk));
	jor g0609(.dina(w_n871_0[1]),.dinb(w_shift1_70[1]),.dout(n872),.clk(gclk));
	jand g0610(.dina(n872),.dinb(n868),.dout(n873),.clk(gclk));
	jand g0611(.dina(w_n873_1[1]),.dinb(w_n308_59[2]),.dout(n874),.clk(gclk));
	jor g0612(.dina(n874),.dinb(n864),.dout(n875),.clk(gclk));
	jor g0613(.dina(n875),.dinb(n854),.dout(n876),.clk(gclk));
	jand g0614(.dina(w_n876_1[1]),.dinb(w_n485_62[2]),.dout(n877),.clk(gclk));
	jor g0615(.dina(n877),.dinb(n833),.dout(n878),.clk(gclk));
	jor g0616(.dina(n878),.dinb(n789),.dout(n879),.clk(gclk));
	jand g0617(.dina(w_n879_0[1]),.dinb(w_n263_63[0]),.dout(n880),.clk(gclk));
	jor g0618(.dina(w_n270_31[1]),.dinb(w_a62_0[0]),.dout(n881),.clk(gclk));
	jor g0619(.dina(w_shift0_31[1]),.dinb(w_a63_0[0]),.dout(n882),.clk(gclk));
	jand g0620(.dina(n882),.dinb(n881),.dout(n883),.clk(gclk));
	jor g0621(.dina(w_n883_0[1]),.dinb(w_n269_70[0]),.dout(n884),.clk(gclk));
	jor g0622(.dina(w_n270_31[0]),.dinb(w_a64_0[0]),.dout(n885),.clk(gclk));
	jor g0623(.dina(w_shift0_31[0]),.dinb(w_a65_0[0]),.dout(n886),.clk(gclk));
	jand g0624(.dina(n886),.dinb(n885),.dout(n887),.clk(gclk));
	jor g0625(.dina(w_n887_0[1]),.dinb(w_shift1_70[0]),.dout(n888),.clk(gclk));
	jand g0626(.dina(n888),.dinb(n884),.dout(n889),.clk(gclk));
	jand g0627(.dina(w_n889_1[1]),.dinb(w_n266_59[1]),.dout(n890),.clk(gclk));
	jor g0628(.dina(w_n270_30[2]),.dinb(w_a54_0[0]),.dout(n891),.clk(gclk));
	jor g0629(.dina(w_shift0_30[2]),.dinb(w_a55_0[0]),.dout(n892),.clk(gclk));
	jand g0630(.dina(n892),.dinb(n891),.dout(n893),.clk(gclk));
	jor g0631(.dina(w_n893_0[1]),.dinb(w_n269_69[2]),.dout(n894),.clk(gclk));
	jor g0632(.dina(w_n270_30[1]),.dinb(w_a56_0[0]),.dout(n895),.clk(gclk));
	jor g0633(.dina(w_shift0_30[1]),.dinb(w_a57_0[0]),.dout(n896),.clk(gclk));
	jand g0634(.dina(n896),.dinb(n895),.dout(n897),.clk(gclk));
	jor g0635(.dina(w_n897_0[1]),.dinb(w_shift1_69[2]),.dout(n898),.clk(gclk));
	jand g0636(.dina(n898),.dinb(n894),.dout(n899),.clk(gclk));
	jand g0637(.dina(w_n899_1[1]),.dinb(w_n281_59[1]),.dout(n900),.clk(gclk));
	jor g0638(.dina(n900),.dinb(n890),.dout(n901),.clk(gclk));
	jor g0639(.dina(w_n270_30[0]),.dinb(w_a58_0[0]),.dout(n902),.clk(gclk));
	jor g0640(.dina(w_shift0_30[0]),.dinb(w_a59_0[0]),.dout(n903),.clk(gclk));
	jand g0641(.dina(n903),.dinb(n902),.dout(n904),.clk(gclk));
	jor g0642(.dina(w_n904_0[1]),.dinb(w_n269_69[1]),.dout(n905),.clk(gclk));
	jor g0643(.dina(w_n270_29[2]),.dinb(w_a60_0[0]),.dout(n906),.clk(gclk));
	jor g0644(.dina(w_shift0_29[2]),.dinb(w_a61_0[0]),.dout(n907),.clk(gclk));
	jand g0645(.dina(n907),.dinb(n906),.dout(n908),.clk(gclk));
	jor g0646(.dina(w_n908_0[1]),.dinb(w_shift1_69[1]),.dout(n909),.clk(gclk));
	jand g0647(.dina(n909),.dinb(n905),.dout(n910),.clk(gclk));
	jand g0648(.dina(w_n910_1[1]),.dinb(w_n295_59[1]),.dout(n911),.clk(gclk));
	jor g0649(.dina(w_n270_29[1]),.dinb(w_a50_0[0]),.dout(n912),.clk(gclk));
	jor g0650(.dina(w_shift0_29[1]),.dinb(w_a51_0[0]),.dout(n913),.clk(gclk));
	jand g0651(.dina(n913),.dinb(n912),.dout(n914),.clk(gclk));
	jor g0652(.dina(w_n914_0[1]),.dinb(w_n269_69[0]),.dout(n915),.clk(gclk));
	jor g0653(.dina(w_n270_29[0]),.dinb(w_a52_0[0]),.dout(n916),.clk(gclk));
	jor g0654(.dina(w_shift0_29[0]),.dinb(w_a53_0[0]),.dout(n917),.clk(gclk));
	jand g0655(.dina(n917),.dinb(n916),.dout(n918),.clk(gclk));
	jor g0656(.dina(w_n918_0[1]),.dinb(w_shift1_69[0]),.dout(n919),.clk(gclk));
	jand g0657(.dina(n919),.dinb(n915),.dout(n920),.clk(gclk));
	jand g0658(.dina(w_n920_1[1]),.dinb(w_n308_59[1]),.dout(n921),.clk(gclk));
	jor g0659(.dina(n921),.dinb(n911),.dout(n922),.clk(gclk));
	jor g0660(.dina(n922),.dinb(n901),.dout(n923),.clk(gclk));
	jand g0661(.dina(w_n923_1[1]),.dinb(w_n485_62[1]),.dout(n924),.clk(gclk));
	jor g0662(.dina(w_n270_28[2]),.dinb(w_a30_0[0]),.dout(n925),.clk(gclk));
	jor g0663(.dina(w_shift0_28[2]),.dinb(w_a31_0[0]),.dout(n926),.clk(gclk));
	jand g0664(.dina(n926),.dinb(n925),.dout(n927),.clk(gclk));
	jor g0665(.dina(w_n927_0[1]),.dinb(w_n269_68[2]),.dout(n928),.clk(gclk));
	jor g0666(.dina(w_n270_28[1]),.dinb(w_a32_0[0]),.dout(n929),.clk(gclk));
	jor g0667(.dina(w_shift0_28[1]),.dinb(w_a33_0[0]),.dout(n930),.clk(gclk));
	jand g0668(.dina(n930),.dinb(n929),.dout(n931),.clk(gclk));
	jor g0669(.dina(w_n931_0[1]),.dinb(w_shift1_68[2]),.dout(n932),.clk(gclk));
	jand g0670(.dina(n932),.dinb(n928),.dout(n933),.clk(gclk));
	jand g0671(.dina(w_n933_1[1]),.dinb(w_n266_59[0]),.dout(n934),.clk(gclk));
	jor g0672(.dina(w_n270_28[0]),.dinb(w_a22_0[0]),.dout(n935),.clk(gclk));
	jor g0673(.dina(w_shift0_28[0]),.dinb(w_a23_0[0]),.dout(n936),.clk(gclk));
	jand g0674(.dina(n936),.dinb(n935),.dout(n937),.clk(gclk));
	jor g0675(.dina(w_n937_0[1]),.dinb(w_n269_68[1]),.dout(n938),.clk(gclk));
	jor g0676(.dina(w_n270_27[2]),.dinb(w_a24_0[0]),.dout(n939),.clk(gclk));
	jor g0677(.dina(w_shift0_27[2]),.dinb(w_a25_0[0]),.dout(n940),.clk(gclk));
	jand g0678(.dina(n940),.dinb(n939),.dout(n941),.clk(gclk));
	jor g0679(.dina(w_n941_0[1]),.dinb(w_shift1_68[1]),.dout(n942),.clk(gclk));
	jand g0680(.dina(n942),.dinb(n938),.dout(n943),.clk(gclk));
	jand g0681(.dina(w_n943_1[1]),.dinb(w_n281_59[0]),.dout(n944),.clk(gclk));
	jor g0682(.dina(n944),.dinb(n934),.dout(n945),.clk(gclk));
	jor g0683(.dina(w_n270_27[1]),.dinb(w_a26_0[0]),.dout(n946),.clk(gclk));
	jor g0684(.dina(w_shift0_27[1]),.dinb(w_a27_0[0]),.dout(n947),.clk(gclk));
	jand g0685(.dina(n947),.dinb(n946),.dout(n948),.clk(gclk));
	jor g0686(.dina(w_n948_0[1]),.dinb(w_n269_68[0]),.dout(n949),.clk(gclk));
	jor g0687(.dina(w_n270_27[0]),.dinb(w_a28_0[0]),.dout(n950),.clk(gclk));
	jor g0688(.dina(w_shift0_27[0]),.dinb(w_a29_0[0]),.dout(n951),.clk(gclk));
	jand g0689(.dina(n951),.dinb(n950),.dout(n952),.clk(gclk));
	jor g0690(.dina(w_n952_0[1]),.dinb(w_shift1_68[0]),.dout(n953),.clk(gclk));
	jand g0691(.dina(n953),.dinb(n949),.dout(n954),.clk(gclk));
	jand g0692(.dina(w_n954_1[1]),.dinb(w_n295_59[0]),.dout(n955),.clk(gclk));
	jor g0693(.dina(w_n270_26[2]),.dinb(w_a18_0[0]),.dout(n956),.clk(gclk));
	jor g0694(.dina(w_shift0_26[2]),.dinb(w_a19_0[0]),.dout(n957),.clk(gclk));
	jand g0695(.dina(n957),.dinb(n956),.dout(n958),.clk(gclk));
	jor g0696(.dina(w_n958_0[1]),.dinb(w_n269_67[2]),.dout(n959),.clk(gclk));
	jor g0697(.dina(w_n270_26[1]),.dinb(w_a20_0[0]),.dout(n960),.clk(gclk));
	jor g0698(.dina(w_shift0_26[1]),.dinb(w_a21_0[0]),.dout(n961),.clk(gclk));
	jand g0699(.dina(n961),.dinb(n960),.dout(n962),.clk(gclk));
	jor g0700(.dina(w_n962_0[1]),.dinb(w_shift1_67[2]),.dout(n963),.clk(gclk));
	jand g0701(.dina(n963),.dinb(n959),.dout(n964),.clk(gclk));
	jand g0702(.dina(w_n964_1[1]),.dinb(w_n308_59[0]),.dout(n965),.clk(gclk));
	jor g0703(.dina(n965),.dinb(n955),.dout(n966),.clk(gclk));
	jor g0704(.dina(n966),.dinb(n945),.dout(n967),.clk(gclk));
	jand g0705(.dina(w_n967_1[1]),.dinb(w_n432_62[1]),.dout(n968),.clk(gclk));
	jor g0706(.dina(n968),.dinb(n924),.dout(n969),.clk(gclk));
	jor g0707(.dina(w_n270_26[0]),.dinb(w_a14_0[0]),.dout(n970),.clk(gclk));
	jor g0708(.dina(w_shift0_26[0]),.dinb(w_a15_0[0]),.dout(n971),.clk(gclk));
	jand g0709(.dina(n971),.dinb(n970),.dout(n972),.clk(gclk));
	jor g0710(.dina(w_n972_0[1]),.dinb(w_n269_67[1]),.dout(n973),.clk(gclk));
	jor g0711(.dina(w_n270_25[2]),.dinb(w_a16_0[0]),.dout(n974),.clk(gclk));
	jor g0712(.dina(w_shift0_25[2]),.dinb(w_a17_0[0]),.dout(n975),.clk(gclk));
	jand g0713(.dina(n975),.dinb(n974),.dout(n976),.clk(gclk));
	jor g0714(.dina(w_n976_0[1]),.dinb(w_shift1_67[1]),.dout(n977),.clk(gclk));
	jand g0715(.dina(n977),.dinb(n973),.dout(n978),.clk(gclk));
	jand g0716(.dina(w_n978_1[1]),.dinb(w_n266_58[2]),.dout(n979),.clk(gclk));
	jor g0717(.dina(w_n270_25[1]),.dinb(w_a6_0[0]),.dout(n980),.clk(gclk));
	jor g0718(.dina(w_shift0_25[1]),.dinb(w_a7_0[0]),.dout(n981),.clk(gclk));
	jand g0719(.dina(n981),.dinb(n980),.dout(n982),.clk(gclk));
	jor g0720(.dina(w_n982_0[1]),.dinb(w_n269_67[0]),.dout(n983),.clk(gclk));
	jor g0721(.dina(w_n270_25[0]),.dinb(w_a8_0[0]),.dout(n984),.clk(gclk));
	jor g0722(.dina(w_shift0_25[0]),.dinb(w_a9_0[0]),.dout(n985),.clk(gclk));
	jand g0723(.dina(n985),.dinb(n984),.dout(n986),.clk(gclk));
	jor g0724(.dina(w_n986_0[1]),.dinb(w_shift1_67[0]),.dout(n987),.clk(gclk));
	jand g0725(.dina(n987),.dinb(n983),.dout(n988),.clk(gclk));
	jand g0726(.dina(w_n988_1[1]),.dinb(w_n281_58[2]),.dout(n989),.clk(gclk));
	jor g0727(.dina(n989),.dinb(n979),.dout(n990),.clk(gclk));
	jor g0728(.dina(w_n270_24[2]),.dinb(w_a10_0[0]),.dout(n991),.clk(gclk));
	jor g0729(.dina(w_shift0_24[2]),.dinb(w_a11_0[0]),.dout(n992),.clk(gclk));
	jand g0730(.dina(n992),.dinb(n991),.dout(n993),.clk(gclk));
	jor g0731(.dina(w_n993_0[1]),.dinb(w_n269_66[2]),.dout(n994),.clk(gclk));
	jor g0732(.dina(w_n270_24[1]),.dinb(w_a12_0[0]),.dout(n995),.clk(gclk));
	jor g0733(.dina(w_shift0_24[1]),.dinb(w_a13_0[0]),.dout(n996),.clk(gclk));
	jand g0734(.dina(n996),.dinb(n995),.dout(n997),.clk(gclk));
	jor g0735(.dina(w_n997_0[1]),.dinb(w_shift1_66[2]),.dout(n998),.clk(gclk));
	jand g0736(.dina(n998),.dinb(n994),.dout(n999),.clk(gclk));
	jand g0737(.dina(w_n999_1[1]),.dinb(w_n295_58[2]),.dout(n1000),.clk(gclk));
	jor g0738(.dina(w_n270_24[0]),.dinb(w_a2_0[0]),.dout(n1001),.clk(gclk));
	jor g0739(.dina(w_shift0_24[0]),.dinb(w_a3_0[0]),.dout(n1002),.clk(gclk));
	jand g0740(.dina(n1002),.dinb(n1001),.dout(n1003),.clk(gclk));
	jor g0741(.dina(w_n1003_0[1]),.dinb(w_n269_66[1]),.dout(n1004),.clk(gclk));
	jor g0742(.dina(w_n270_23[2]),.dinb(w_a4_0[0]),.dout(n1005),.clk(gclk));
	jor g0743(.dina(w_shift0_23[2]),.dinb(w_a5_0[0]),.dout(n1006),.clk(gclk));
	jand g0744(.dina(n1006),.dinb(n1005),.dout(n1007),.clk(gclk));
	jor g0745(.dina(w_n1007_0[1]),.dinb(w_shift1_66[1]),.dout(n1008),.clk(gclk));
	jand g0746(.dina(n1008),.dinb(n1004),.dout(n1009),.clk(gclk));
	jand g0747(.dina(w_n1009_1[1]),.dinb(w_n308_58[2]),.dout(n1010),.clk(gclk));
	jor g0748(.dina(n1010),.dinb(n1000),.dout(n1011),.clk(gclk));
	jor g0749(.dina(n1011),.dinb(n990),.dout(n1012),.clk(gclk));
	jand g0750(.dina(w_n1012_1[1]),.dinb(w_n323_62[1]),.dout(n1013),.clk(gclk));
	jor g0751(.dina(w_n270_23[1]),.dinb(w_a48_0[0]),.dout(n1014),.clk(gclk));
	jor g0752(.dina(w_shift0_23[1]),.dinb(w_a49_0[0]),.dout(n1015),.clk(gclk));
	jand g0753(.dina(n1015),.dinb(n1014),.dout(n1016),.clk(gclk));
	jand g0754(.dina(w_n1016_0[1]),.dinb(w_n269_66[0]),.dout(n1017),.clk(gclk));
	jand g0755(.dina(w_n270_23[0]),.dinb(w_a47_0[0]),.dout(n1018),.clk(gclk));
	jand g0756(.dina(w_shift0_23[0]),.dinb(w_a46_0[0]),.dout(n1019),.clk(gclk));
	jor g0757(.dina(w_n1019_0[1]),.dinb(w_n1018_0[1]),.dout(n1020),.clk(gclk));
	jand g0758(.dina(n1020),.dinb(w_shift1_66[0]),.dout(n1021),.clk(gclk));
	jor g0759(.dina(n1021),.dinb(n1017),.dout(n1022),.clk(gclk));
	jand g0760(.dina(w_n1022_1[1]),.dinb(w_n266_58[1]),.dout(n1023),.clk(gclk));
	jand g0761(.dina(w_n270_22[2]),.dinb(w_a39_0[0]),.dout(n1024),.clk(gclk));
	jor g0762(.dina(w_n1024_0[1]),.dinb(w_n269_65[2]),.dout(n1025),.clk(gclk));
	jand g0763(.dina(w_n270_22[1]),.dinb(w_a41_0[0]),.dout(n1026),.clk(gclk));
	jor g0764(.dina(w_n1026_0[1]),.dinb(w_shift1_65[2]),.dout(n1027),.clk(gclk));
	jand g0765(.dina(n1027),.dinb(n1025),.dout(n1028),.clk(gclk));
	jand g0766(.dina(w_shift0_22[2]),.dinb(w_a38_0[0]),.dout(n1029),.clk(gclk));
	jand g0767(.dina(w_n1029_0[1]),.dinb(w_shift1_65[1]),.dout(n1030),.clk(gclk));
	jand g0768(.dina(w_shift0_22[1]),.dinb(w_a40_0[0]),.dout(n1031),.clk(gclk));
	jand g0769(.dina(w_n1031_0[1]),.dinb(w_n269_65[1]),.dout(n1032),.clk(gclk));
	jor g0770(.dina(n1032),.dinb(n1030),.dout(n1033),.clk(gclk));
	jor g0771(.dina(n1033),.dinb(n1028),.dout(n1034),.clk(gclk));
	jand g0772(.dina(w_n1034_1[1]),.dinb(w_n281_58[1]),.dout(n1035),.clk(gclk));
	jor g0773(.dina(n1035),.dinb(n1023),.dout(n1036),.clk(gclk));
	jand g0774(.dina(w_shift0_22[0]),.dinb(w_a44_0[0]),.dout(n1037),.clk(gclk));
	jor g0775(.dina(w_n1037_0[1]),.dinb(w_shift1_65[0]),.dout(n1038),.clk(gclk));
	jand g0776(.dina(w_n270_22[0]),.dinb(w_a43_0[0]),.dout(n1039),.clk(gclk));
	jor g0777(.dina(w_n1039_0[1]),.dinb(w_n269_65[0]),.dout(n1040),.clk(gclk));
	jand g0778(.dina(n1040),.dinb(n1038),.dout(n1041),.clk(gclk));
	jand g0779(.dina(w_shift0_21[2]),.dinb(w_a42_0[0]),.dout(n1042),.clk(gclk));
	jand g0780(.dina(w_n1042_0[1]),.dinb(w_shift1_64[2]),.dout(n1043),.clk(gclk));
	jand g0781(.dina(w_n270_21[2]),.dinb(w_a45_0[0]),.dout(n1044),.clk(gclk));
	jand g0782(.dina(w_n1044_0[1]),.dinb(w_n269_64[2]),.dout(n1045),.clk(gclk));
	jor g0783(.dina(n1045),.dinb(n1043),.dout(n1046),.clk(gclk));
	jor g0784(.dina(n1046),.dinb(n1041),.dout(n1047),.clk(gclk));
	jand g0785(.dina(w_n1047_1[1]),.dinb(w_n295_58[1]),.dout(n1048),.clk(gclk));
	jor g0786(.dina(w_n270_21[1]),.dinb(w_a34_0[0]),.dout(n1049),.clk(gclk));
	jor g0787(.dina(w_shift0_21[1]),.dinb(w_a35_0[0]),.dout(n1050),.clk(gclk));
	jand g0788(.dina(n1050),.dinb(n1049),.dout(n1051),.clk(gclk));
	jor g0789(.dina(w_n1051_0[1]),.dinb(w_n269_64[1]),.dout(n1052),.clk(gclk));
	jor g0790(.dina(w_n270_21[0]),.dinb(w_a36_0[0]),.dout(n1053),.clk(gclk));
	jor g0791(.dina(w_shift0_21[0]),.dinb(w_a37_0[0]),.dout(n1054),.clk(gclk));
	jand g0792(.dina(n1054),.dinb(n1053),.dout(n1055),.clk(gclk));
	jor g0793(.dina(w_n1055_0[1]),.dinb(w_shift1_64[1]),.dout(n1056),.clk(gclk));
	jand g0794(.dina(n1056),.dinb(n1052),.dout(n1057),.clk(gclk));
	jand g0795(.dina(w_n1057_1[1]),.dinb(w_n308_58[1]),.dout(n1058),.clk(gclk));
	jor g0796(.dina(n1058),.dinb(n1048),.dout(n1059),.clk(gclk));
	jor g0797(.dina(n1059),.dinb(n1036),.dout(n1060),.clk(gclk));
	jand g0798(.dina(w_n1060_1[1]),.dinb(w_n377_62[1]),.dout(n1061),.clk(gclk));
	jor g0799(.dina(n1061),.dinb(n1013),.dout(n1062),.clk(gclk));
	jor g0800(.dina(n1062),.dinb(n969),.dout(n1063),.clk(gclk));
	jand g0801(.dina(w_n1063_0[1]),.dinb(w_shift6_63[0]),.dout(n1064),.clk(gclk));
	jor g0802(.dina(n1064),.dinb(n880),.dout(result1),.clk(gclk));
	jor g0803(.dina(w_n419_0[0]),.dinb(w_shift1_64[0]),.dout(n1066),.clk(gclk));
	jor g0804(.dina(w_n267_0[0]),.dinb(w_n269_64[0]),.dout(n1067),.clk(gclk));
	jand g0805(.dina(n1067),.dinb(n1066),.dout(n1068),.clk(gclk));
	jand g0806(.dina(w_n276_0[0]),.dinb(w_shift1_63[2]),.dout(n1069),.clk(gclk));
	jand g0807(.dina(w_n422_0[0]),.dinb(w_n269_63[2]),.dout(n1070),.clk(gclk));
	jor g0808(.dina(n1070),.dinb(n1069),.dout(n1071),.clk(gclk));
	jor g0809(.dina(n1071),.dinb(n1068),.dout(n1072),.clk(gclk));
	jand g0810(.dina(w_n1072_1[1]),.dinb(w_n266_58[0]),.dout(n1073),.clk(gclk));
	jor g0811(.dina(w_n298_0[0]),.dinb(w_shift1_63[1]),.dout(n1074),.clk(gclk));
	jor g0812(.dina(w_n282_0[0]),.dinb(w_n269_63[1]),.dout(n1075),.clk(gclk));
	jand g0813(.dina(n1075),.dinb(n1074),.dout(n1076),.clk(gclk));
	jand g0814(.dina(w_n289_0[0]),.dinb(w_shift1_63[0]),.dout(n1077),.clk(gclk));
	jand g0815(.dina(w_n301_0[0]),.dinb(w_n269_63[0]),.dout(n1078),.clk(gclk));
	jor g0816(.dina(n1078),.dinb(n1077),.dout(n1079),.clk(gclk));
	jor g0817(.dina(n1079),.dinb(n1076),.dout(n1080),.clk(gclk));
	jand g0818(.dina(w_n1080_1[1]),.dinb(w_n281_58[0]),.dout(n1081),.clk(gclk));
	jor g0819(.dina(n1081),.dinb(n1073),.dout(n1082),.clk(gclk));
	jor g0820(.dina(w_n271_0[0]),.dinb(w_shift1_62[2]),.dout(n1083),.clk(gclk));
	jor g0821(.dina(w_n296_0[0]),.dinb(w_n269_62[2]),.dout(n1084),.clk(gclk));
	jand g0822(.dina(n1084),.dinb(n1083),.dout(n1085),.clk(gclk));
	jand g0823(.dina(w_n303_0[0]),.dinb(w_shift1_62[1]),.dout(n1086),.clk(gclk));
	jand g0824(.dina(w_n274_0[0]),.dinb(w_n269_62[1]),.dout(n1087),.clk(gclk));
	jor g0825(.dina(n1087),.dinb(n1086),.dout(n1088),.clk(gclk));
	jor g0826(.dina(n1088),.dinb(n1085),.dout(n1089),.clk(gclk));
	jand g0827(.dina(w_n1089_1[1]),.dinb(w_n295_58[0]),.dout(n1090),.clk(gclk));
	jor g0828(.dina(w_n284_0[0]),.dinb(w_shift1_62[0]),.dout(n1091),.clk(gclk));
	jor g0829(.dina(w_n309_0[0]),.dinb(w_n269_62[0]),.dout(n1092),.clk(gclk));
	jand g0830(.dina(n1092),.dinb(n1091),.dout(n1093),.clk(gclk));
	jand g0831(.dina(w_n316_0[0]),.dinb(w_shift1_61[2]),.dout(n1094),.clk(gclk));
	jand g0832(.dina(w_n287_0[0]),.dinb(w_n269_61[2]),.dout(n1095),.clk(gclk));
	jor g0833(.dina(n1095),.dinb(n1094),.dout(n1096),.clk(gclk));
	jor g0834(.dina(n1096),.dinb(n1093),.dout(n1097),.clk(gclk));
	jand g0835(.dina(w_n1097_1[1]),.dinb(w_n308_58[0]),.dout(n1098),.clk(gclk));
	jor g0836(.dina(n1098),.dinb(n1090),.dout(n1099),.clk(gclk));
	jor g0837(.dina(n1099),.dinb(n1082),.dout(n1100),.clk(gclk));
	jand g0838(.dina(w_n1100_1[1]),.dinb(w_n323_62[0]),.dout(n1101),.clk(gclk));
	jor g0839(.dina(w_n473_0[0]),.dinb(w_shift1_61[1]),.dout(n1102),.clk(gclk));
	jor g0840(.dina(w_n325_0[0]),.dinb(w_n269_61[1]),.dout(n1103),.clk(gclk));
	jand g0841(.dina(n1103),.dinb(n1102),.dout(n1104),.clk(gclk));
	jand g0842(.dina(w_n332_0[0]),.dinb(w_shift1_61[0]),.dout(n1105),.clk(gclk));
	jand g0843(.dina(w_n476_0[0]),.dinb(w_n269_61[0]),.dout(n1106),.clk(gclk));
	jor g0844(.dina(n1106),.dinb(n1105),.dout(n1107),.clk(gclk));
	jor g0845(.dina(n1107),.dinb(n1104),.dout(n1108),.clk(gclk));
	jand g0846(.dina(w_n1108_1[1]),.dinb(w_n266_57[2]),.dout(n1109),.clk(gclk));
	jor g0847(.dina(w_n352_0[0]),.dinb(w_shift1_60[2]),.dout(n1110),.clk(gclk));
	jor g0848(.dina(w_n337_0[0]),.dinb(w_n269_60[2]),.dout(n1111),.clk(gclk));
	jand g0849(.dina(n1111),.dinb(n1110),.dout(n1112),.clk(gclk));
	jand g0850(.dina(w_n344_0[0]),.dinb(w_shift1_60[1]),.dout(n1113),.clk(gclk));
	jand g0851(.dina(w_n355_0[0]),.dinb(w_n269_60[1]),.dout(n1114),.clk(gclk));
	jor g0852(.dina(n1114),.dinb(n1113),.dout(n1115),.clk(gclk));
	jor g0853(.dina(n1115),.dinb(n1112),.dout(n1116),.clk(gclk));
	jand g0854(.dina(w_n1116_1[1]),.dinb(w_n281_57[2]),.dout(n1117),.clk(gclk));
	jor g0855(.dina(n1117),.dinb(n1109),.dout(n1118),.clk(gclk));
	jor g0856(.dina(w_n327_0[0]),.dinb(w_shift1_60[0]),.dout(n1119),.clk(gclk));
	jor g0857(.dina(w_n350_0[0]),.dinb(w_n269_60[0]),.dout(n1120),.clk(gclk));
	jand g0858(.dina(n1120),.dinb(n1119),.dout(n1121),.clk(gclk));
	jand g0859(.dina(w_n357_0[0]),.dinb(w_shift1_59[2]),.dout(n1122),.clk(gclk));
	jand g0860(.dina(w_n330_0[0]),.dinb(w_n269_59[2]),.dout(n1123),.clk(gclk));
	jor g0861(.dina(n1123),.dinb(n1122),.dout(n1124),.clk(gclk));
	jor g0862(.dina(n1124),.dinb(n1121),.dout(n1125),.clk(gclk));
	jand g0863(.dina(w_n1125_1[1]),.dinb(w_n295_57[2]),.dout(n1126),.clk(gclk));
	jor g0864(.dina(w_n339_0[0]),.dinb(w_shift1_59[1]),.dout(n1127),.clk(gclk));
	jor g0865(.dina(w_n362_0[0]),.dinb(w_n269_59[1]),.dout(n1128),.clk(gclk));
	jand g0866(.dina(n1128),.dinb(n1127),.dout(n1129),.clk(gclk));
	jand g0867(.dina(w_n369_0[0]),.dinb(w_shift1_59[0]),.dout(n1130),.clk(gclk));
	jand g0868(.dina(w_n342_0[0]),.dinb(w_n269_59[0]),.dout(n1131),.clk(gclk));
	jor g0869(.dina(n1131),.dinb(n1130),.dout(n1132),.clk(gclk));
	jor g0870(.dina(n1132),.dinb(n1129),.dout(n1133),.clk(gclk));
	jand g0871(.dina(w_n1133_1[1]),.dinb(w_n308_57[2]),.dout(n1134),.clk(gclk));
	jor g0872(.dina(n1134),.dinb(n1126),.dout(n1135),.clk(gclk));
	jor g0873(.dina(n1135),.dinb(n1118),.dout(n1136),.clk(gclk));
	jand g0874(.dina(w_n1136_1[1]),.dinb(w_n377_62[0]),.dout(n1137),.clk(gclk));
	jor g0875(.dina(n1137),.dinb(n1101),.dout(n1138),.clk(gclk));
	jor g0876(.dina(w_n364_0[0]),.dinb(w_shift1_58[2]),.dout(n1139),.clk(gclk));
	jor g0877(.dina(w_n380_0[0]),.dinb(w_n269_58[2]),.dout(n1140),.clk(gclk));
	jand g0878(.dina(n1140),.dinb(n1139),.dout(n1141),.clk(gclk));
	jand g0879(.dina(w_n387_0[0]),.dinb(w_shift1_58[1]),.dout(n1142),.clk(gclk));
	jand g0880(.dina(w_n367_0[0]),.dinb(w_n269_58[1]),.dout(n1143),.clk(gclk));
	jor g0881(.dina(n1143),.dinb(n1142),.dout(n1144),.clk(gclk));
	jor g0882(.dina(n1144),.dinb(n1141),.dout(n1145),.clk(gclk));
	jand g0883(.dina(w_n1145_1[1]),.dinb(w_n266_57[1]),.dout(n1146),.clk(gclk));
	jor g0884(.dina(w_n407_0[0]),.dinb(w_shift1_58[0]),.dout(n1147),.clk(gclk));
	jor g0885(.dina(w_n392_0[0]),.dinb(w_n269_58[0]),.dout(n1148),.clk(gclk));
	jand g0886(.dina(n1148),.dinb(n1147),.dout(n1149),.clk(gclk));
	jand g0887(.dina(w_n399_0[0]),.dinb(w_shift1_57[2]),.dout(n1150),.clk(gclk));
	jand g0888(.dina(w_n410_0[0]),.dinb(w_n269_57[2]),.dout(n1151),.clk(gclk));
	jor g0889(.dina(n1151),.dinb(n1150),.dout(n1152),.clk(gclk));
	jor g0890(.dina(n1152),.dinb(n1149),.dout(n1153),.clk(gclk));
	jand g0891(.dina(w_n1153_1[1]),.dinb(w_n281_57[1]),.dout(n1154),.clk(gclk));
	jor g0892(.dina(n1154),.dinb(n1146),.dout(n1155),.clk(gclk));
	jor g0893(.dina(w_n382_0[0]),.dinb(w_shift1_57[1]),.dout(n1156),.clk(gclk));
	jor g0894(.dina(w_n405_0[0]),.dinb(w_n269_57[1]),.dout(n1157),.clk(gclk));
	jand g0895(.dina(n1157),.dinb(n1156),.dout(n1158),.clk(gclk));
	jand g0896(.dina(w_n412_0[0]),.dinb(w_shift1_57[0]),.dout(n1159),.clk(gclk));
	jand g0897(.dina(w_n385_0[0]),.dinb(w_n269_57[0]),.dout(n1160),.clk(gclk));
	jor g0898(.dina(n1160),.dinb(n1159),.dout(n1161),.clk(gclk));
	jor g0899(.dina(n1161),.dinb(n1158),.dout(n1162),.clk(gclk));
	jand g0900(.dina(w_n1162_1[1]),.dinb(w_n295_57[1]),.dout(n1163),.clk(gclk));
	jor g0901(.dina(w_n394_0[0]),.dinb(w_shift1_56[2]),.dout(n1164),.clk(gclk));
	jor g0902(.dina(w_n417_0[0]),.dinb(w_n269_56[2]),.dout(n1165),.clk(gclk));
	jand g0903(.dina(n1165),.dinb(n1164),.dout(n1166),.clk(gclk));
	jand g0904(.dina(w_n424_0[0]),.dinb(w_shift1_56[1]),.dout(n1167),.clk(gclk));
	jand g0905(.dina(w_n397_0[0]),.dinb(w_n269_56[1]),.dout(n1168),.clk(gclk));
	jor g0906(.dina(n1168),.dinb(n1167),.dout(n1169),.clk(gclk));
	jor g0907(.dina(n1169),.dinb(n1166),.dout(n1170),.clk(gclk));
	jand g0908(.dina(w_n1170_1[1]),.dinb(w_n308_57[1]),.dout(n1171),.clk(gclk));
	jor g0909(.dina(n1171),.dinb(n1163),.dout(n1172),.clk(gclk));
	jor g0910(.dina(n1172),.dinb(n1155),.dout(n1173),.clk(gclk));
	jand g0911(.dina(w_n1173_1[1]),.dinb(w_n432_62[0]),.dout(n1174),.clk(gclk));
	jor g0912(.dina(w_n529_0[0]),.dinb(w_shift1_56[0]),.dout(n1175),.clk(gclk));
	jor g0913(.dina(w_n434_0[0]),.dinb(w_n269_56[0]),.dout(n1176),.clk(gclk));
	jand g0914(.dina(n1176),.dinb(n1175),.dout(n1177),.clk(gclk));
	jand g0915(.dina(w_n441_0[0]),.dinb(w_shift1_55[2]),.dout(n1178),.clk(gclk));
	jand g0916(.dina(w_n532_0[0]),.dinb(w_n269_55[2]),.dout(n1179),.clk(gclk));
	jor g0917(.dina(n1179),.dinb(n1178),.dout(n1180),.clk(gclk));
	jor g0918(.dina(n1180),.dinb(n1177),.dout(n1181),.clk(gclk));
	jand g0919(.dina(w_n1181_1[1]),.dinb(w_n266_57[0]),.dout(n1182),.clk(gclk));
	jor g0920(.dina(w_n461_0[0]),.dinb(w_shift1_55[1]),.dout(n1183),.clk(gclk));
	jor g0921(.dina(w_n446_0[0]),.dinb(w_n269_55[1]),.dout(n1184),.clk(gclk));
	jand g0922(.dina(n1184),.dinb(n1183),.dout(n1185),.clk(gclk));
	jand g0923(.dina(w_n453_0[0]),.dinb(w_shift1_55[0]),.dout(n1186),.clk(gclk));
	jand g0924(.dina(w_n464_0[0]),.dinb(w_n269_55[0]),.dout(n1187),.clk(gclk));
	jor g0925(.dina(n1187),.dinb(n1186),.dout(n1188),.clk(gclk));
	jor g0926(.dina(n1188),.dinb(n1185),.dout(n1189),.clk(gclk));
	jand g0927(.dina(w_n1189_1[1]),.dinb(w_n281_57[0]),.dout(n1190),.clk(gclk));
	jor g0928(.dina(n1190),.dinb(n1182),.dout(n1191),.clk(gclk));
	jor g0929(.dina(w_n436_0[0]),.dinb(w_shift1_54[2]),.dout(n1192),.clk(gclk));
	jor g0930(.dina(w_n459_0[0]),.dinb(w_n269_54[2]),.dout(n1193),.clk(gclk));
	jand g0931(.dina(n1193),.dinb(n1192),.dout(n1194),.clk(gclk));
	jand g0932(.dina(w_n466_0[0]),.dinb(w_shift1_54[1]),.dout(n1195),.clk(gclk));
	jand g0933(.dina(w_n439_0[0]),.dinb(w_n269_54[1]),.dout(n1196),.clk(gclk));
	jor g0934(.dina(n1196),.dinb(n1195),.dout(n1197),.clk(gclk));
	jor g0935(.dina(n1197),.dinb(n1194),.dout(n1198),.clk(gclk));
	jand g0936(.dina(w_n1198_1[1]),.dinb(w_n295_57[0]),.dout(n1199),.clk(gclk));
	jor g0937(.dina(w_n448_0[0]),.dinb(w_shift1_54[0]),.dout(n1200),.clk(gclk));
	jor g0938(.dina(w_n471_0[0]),.dinb(w_n269_54[0]),.dout(n1201),.clk(gclk));
	jand g0939(.dina(n1201),.dinb(n1200),.dout(n1202),.clk(gclk));
	jand g0940(.dina(w_n478_0[0]),.dinb(w_shift1_53[2]),.dout(n1203),.clk(gclk));
	jand g0941(.dina(w_n451_0[0]),.dinb(w_n269_53[2]),.dout(n1204),.clk(gclk));
	jor g0942(.dina(n1204),.dinb(n1203),.dout(n1205),.clk(gclk));
	jor g0943(.dina(n1205),.dinb(n1202),.dout(n1206),.clk(gclk));
	jand g0944(.dina(w_n1206_1[1]),.dinb(w_n308_57[0]),.dout(n1207),.clk(gclk));
	jor g0945(.dina(n1207),.dinb(n1199),.dout(n1208),.clk(gclk));
	jor g0946(.dina(n1208),.dinb(n1191),.dout(n1209),.clk(gclk));
	jand g0947(.dina(w_n1209_1[1]),.dinb(w_n485_62[0]),.dout(n1210),.clk(gclk));
	jor g0948(.dina(n1210),.dinb(n1174),.dout(n1211),.clk(gclk));
	jor g0949(.dina(n1211),.dinb(n1138),.dout(n1212),.clk(gclk));
	jand g0950(.dina(w_n1212_0[1]),.dinb(w_n263_62[2]),.dout(n1213),.clk(gclk));
	jor g0951(.dina(w_n311_0[0]),.dinb(w_shift1_53[1]),.dout(n1214),.clk(gclk));
	jor g0952(.dina(w_n645_0[0]),.dinb(w_n269_53[1]),.dout(n1215),.clk(gclk));
	jand g0953(.dina(n1215),.dinb(n1214),.dout(n1216),.clk(gclk));
	jand g0954(.dina(w_n652_0[0]),.dinb(w_shift1_53[0]),.dout(n1217),.clk(gclk));
	jand g0955(.dina(w_n314_0[0]),.dinb(w_n269_53[0]),.dout(n1218),.clk(gclk));
	jor g0956(.dina(n1218),.dinb(n1217),.dout(n1219),.clk(gclk));
	jor g0957(.dina(n1219),.dinb(n1216),.dout(n1220),.clk(gclk));
	jand g0958(.dina(w_n1220_1[1]),.dinb(w_n266_56[2]),.dout(n1221),.clk(gclk));
	jor g0959(.dina(w_n672_0[0]),.dinb(w_shift1_52[2]),.dout(n1222),.clk(gclk));
	jor g0960(.dina(w_n657_0[0]),.dinb(w_n269_52[2]),.dout(n1223),.clk(gclk));
	jand g0961(.dina(n1223),.dinb(n1222),.dout(n1224),.clk(gclk));
	jand g0962(.dina(w_n664_0[0]),.dinb(w_shift1_52[1]),.dout(n1225),.clk(gclk));
	jand g0963(.dina(w_n675_0[0]),.dinb(w_n269_52[1]),.dout(n1226),.clk(gclk));
	jor g0964(.dina(n1226),.dinb(n1225),.dout(n1227),.clk(gclk));
	jor g0965(.dina(n1227),.dinb(n1224),.dout(n1228),.clk(gclk));
	jand g0966(.dina(w_n1228_1[1]),.dinb(w_n281_56[2]),.dout(n1229),.clk(gclk));
	jor g0967(.dina(n1229),.dinb(n1221),.dout(n1230),.clk(gclk));
	jor g0968(.dina(w_n647_0[0]),.dinb(w_shift1_52[0]),.dout(n1231),.clk(gclk));
	jor g0969(.dina(w_n670_0[0]),.dinb(w_n269_52[0]),.dout(n1232),.clk(gclk));
	jand g0970(.dina(n1232),.dinb(n1231),.dout(n1233),.clk(gclk));
	jand g0971(.dina(w_n677_0[0]),.dinb(w_shift1_51[2]),.dout(n1234),.clk(gclk));
	jand g0972(.dina(w_n650_0[0]),.dinb(w_n269_51[2]),.dout(n1235),.clk(gclk));
	jor g0973(.dina(n1235),.dinb(n1234),.dout(n1236),.clk(gclk));
	jor g0974(.dina(n1236),.dinb(n1233),.dout(n1237),.clk(gclk));
	jand g0975(.dina(w_n1237_1[1]),.dinb(w_n295_56[2]),.dout(n1238),.clk(gclk));
	jor g0976(.dina(w_n659_0[0]),.dinb(w_shift1_51[1]),.dout(n1239),.clk(gclk));
	jor g0977(.dina(w_n682_0[0]),.dinb(w_n269_51[1]),.dout(n1240),.clk(gclk));
	jand g0978(.dina(n1240),.dinb(n1239),.dout(n1241),.clk(gclk));
	jand g0979(.dina(w_n689_0[0]),.dinb(w_shift1_51[0]),.dout(n1242),.clk(gclk));
	jand g0980(.dina(w_n662_0[0]),.dinb(w_n269_51[0]),.dout(n1243),.clk(gclk));
	jor g0981(.dina(n1243),.dinb(n1242),.dout(n1244),.clk(gclk));
	jor g0982(.dina(n1244),.dinb(n1241),.dout(n1245),.clk(gclk));
	jand g0983(.dina(w_n1245_1[1]),.dinb(w_n308_56[2]),.dout(n1246),.clk(gclk));
	jor g0984(.dina(n1246),.dinb(n1238),.dout(n1247),.clk(gclk));
	jor g0985(.dina(n1247),.dinb(n1230),.dout(n1248),.clk(gclk));
	jand g0986(.dina(w_n1248_1[1]),.dinb(w_n485_61[2]),.dout(n1249),.clk(gclk));
	jor g0987(.dina(w_n579_0[0]),.dinb(w_shift1_50[2]),.dout(n1250),.clk(gclk));
	jor g0988(.dina(w_n593_0[0]),.dinb(w_n269_50[2]),.dout(n1251),.clk(gclk));
	jand g0989(.dina(n1251),.dinb(n1250),.dout(n1252),.clk(gclk));
	jand g0990(.dina(w_n600_0[0]),.dinb(w_shift1_50[1]),.dout(n1253),.clk(gclk));
	jand g0991(.dina(w_n582_0[0]),.dinb(w_n269_50[1]),.dout(n1254),.clk(gclk));
	jor g0992(.dina(n1254),.dinb(n1253),.dout(n1255),.clk(gclk));
	jor g0993(.dina(n1255),.dinb(n1252),.dout(n1256),.clk(gclk));
	jand g0994(.dina(w_n1256_1[1]),.dinb(w_n266_56[1]),.dout(n1257),.clk(gclk));
	jor g0995(.dina(w_n620_0[0]),.dinb(w_shift1_50[0]),.dout(n1258),.clk(gclk));
	jor g0996(.dina(w_n605_0[0]),.dinb(w_n269_50[0]),.dout(n1259),.clk(gclk));
	jand g0997(.dina(n1259),.dinb(n1258),.dout(n1260),.clk(gclk));
	jand g0998(.dina(w_n612_0[0]),.dinb(w_shift1_49[2]),.dout(n1261),.clk(gclk));
	jand g0999(.dina(w_n623_0[0]),.dinb(w_n269_49[2]),.dout(n1262),.clk(gclk));
	jor g1000(.dina(n1262),.dinb(n1261),.dout(n1263),.clk(gclk));
	jor g1001(.dina(n1263),.dinb(n1260),.dout(n1264),.clk(gclk));
	jand g1002(.dina(w_n1264_1[1]),.dinb(w_n281_56[1]),.dout(n1265),.clk(gclk));
	jor g1003(.dina(n1265),.dinb(n1257),.dout(n1266),.clk(gclk));
	jor g1004(.dina(w_n595_0[0]),.dinb(w_shift1_49[1]),.dout(n1267),.clk(gclk));
	jor g1005(.dina(w_n618_0[0]),.dinb(w_n269_49[1]),.dout(n1268),.clk(gclk));
	jand g1006(.dina(n1268),.dinb(n1267),.dout(n1269),.clk(gclk));
	jand g1007(.dina(w_n625_0[0]),.dinb(w_shift1_49[0]),.dout(n1270),.clk(gclk));
	jand g1008(.dina(w_n598_0[0]),.dinb(w_n269_49[0]),.dout(n1271),.clk(gclk));
	jor g1009(.dina(n1271),.dinb(n1270),.dout(n1272),.clk(gclk));
	jor g1010(.dina(n1272),.dinb(n1269),.dout(n1273),.clk(gclk));
	jand g1011(.dina(w_n1273_1[1]),.dinb(w_n295_56[1]),.dout(n1274),.clk(gclk));
	jor g1012(.dina(w_n607_0[0]),.dinb(w_shift1_48[2]),.dout(n1275),.clk(gclk));
	jor g1013(.dina(w_n630_0[0]),.dinb(w_n269_48[2]),.dout(n1276),.clk(gclk));
	jand g1014(.dina(n1276),.dinb(n1275),.dout(n1277),.clk(gclk));
	jand g1015(.dina(w_n637_0[0]),.dinb(w_shift1_48[1]),.dout(n1278),.clk(gclk));
	jand g1016(.dina(w_n610_0[0]),.dinb(w_n269_48[1]),.dout(n1279),.clk(gclk));
	jor g1017(.dina(n1279),.dinb(n1278),.dout(n1280),.clk(gclk));
	jor g1018(.dina(n1280),.dinb(n1277),.dout(n1281),.clk(gclk));
	jand g1019(.dina(w_n1281_1[1]),.dinb(w_n308_56[1]),.dout(n1282),.clk(gclk));
	jor g1020(.dina(n1282),.dinb(n1274),.dout(n1283),.clk(gclk));
	jor g1021(.dina(n1283),.dinb(n1266),.dout(n1284),.clk(gclk));
	jand g1022(.dina(w_n1284_1[1]),.dinb(w_n432_61[2]),.dout(n1285),.clk(gclk));
	jor g1023(.dina(n1285),.dinb(n1249),.dout(n1286),.clk(gclk));
	jor g1024(.dina(w_n632_0[0]),.dinb(w_shift1_48[0]),.dout(n1287),.clk(gclk));
	jor g1025(.dina(w_n490_0[0]),.dinb(w_n269_48[0]),.dout(n1288),.clk(gclk));
	jand g1026(.dina(n1288),.dinb(n1287),.dout(n1289),.clk(gclk));
	jand g1027(.dina(w_n497_0[0]),.dinb(w_shift1_47[2]),.dout(n1290),.clk(gclk));
	jand g1028(.dina(w_n635_0[0]),.dinb(w_n269_47[2]),.dout(n1291),.clk(gclk));
	jor g1029(.dina(n1291),.dinb(n1290),.dout(n1292),.clk(gclk));
	jor g1030(.dina(n1292),.dinb(n1289),.dout(n1293),.clk(gclk));
	jand g1031(.dina(w_n1293_1[1]),.dinb(w_n266_56[0]),.dout(n1294),.clk(gclk));
	jor g1032(.dina(w_n517_0[0]),.dinb(w_shift1_47[1]),.dout(n1295),.clk(gclk));
	jor g1033(.dina(w_n502_0[0]),.dinb(w_n269_47[1]),.dout(n1296),.clk(gclk));
	jand g1034(.dina(n1296),.dinb(n1295),.dout(n1297),.clk(gclk));
	jand g1035(.dina(w_n509_0[0]),.dinb(w_shift1_47[0]),.dout(n1298),.clk(gclk));
	jand g1036(.dina(w_n520_0[0]),.dinb(w_n269_47[0]),.dout(n1299),.clk(gclk));
	jor g1037(.dina(n1299),.dinb(n1298),.dout(n1300),.clk(gclk));
	jor g1038(.dina(n1300),.dinb(n1297),.dout(n1301),.clk(gclk));
	jand g1039(.dina(w_n1301_1[1]),.dinb(w_n281_56[0]),.dout(n1302),.clk(gclk));
	jor g1040(.dina(n1302),.dinb(n1294),.dout(n1303),.clk(gclk));
	jor g1041(.dina(w_n492_0[0]),.dinb(w_shift1_46[2]),.dout(n1304),.clk(gclk));
	jor g1042(.dina(w_n515_0[0]),.dinb(w_n269_46[2]),.dout(n1305),.clk(gclk));
	jand g1043(.dina(n1305),.dinb(n1304),.dout(n1306),.clk(gclk));
	jand g1044(.dina(w_n522_0[0]),.dinb(w_shift1_46[1]),.dout(n1307),.clk(gclk));
	jand g1045(.dina(w_n495_0[0]),.dinb(w_n269_46[1]),.dout(n1308),.clk(gclk));
	jor g1046(.dina(n1308),.dinb(n1307),.dout(n1309),.clk(gclk));
	jor g1047(.dina(n1309),.dinb(n1306),.dout(n1310),.clk(gclk));
	jand g1048(.dina(w_n1310_1[1]),.dinb(w_n295_56[0]),.dout(n1311),.clk(gclk));
	jor g1049(.dina(w_n504_0[0]),.dinb(w_shift1_46[0]),.dout(n1312),.clk(gclk));
	jor g1050(.dina(w_n527_0[0]),.dinb(w_n269_46[0]),.dout(n1313),.clk(gclk));
	jand g1051(.dina(n1313),.dinb(n1312),.dout(n1314),.clk(gclk));
	jand g1052(.dina(w_n534_0[0]),.dinb(w_shift1_45[2]),.dout(n1315),.clk(gclk));
	jand g1053(.dina(w_n507_0[0]),.dinb(w_n269_45[2]),.dout(n1316),.clk(gclk));
	jor g1054(.dina(n1316),.dinb(n1315),.dout(n1317),.clk(gclk));
	jor g1055(.dina(n1317),.dinb(n1314),.dout(n1318),.clk(gclk));
	jand g1056(.dina(w_n1318_1[1]),.dinb(w_n308_56[0]),.dout(n1319),.clk(gclk));
	jor g1057(.dina(n1319),.dinb(n1311),.dout(n1320),.clk(gclk));
	jor g1058(.dina(n1320),.dinb(n1303),.dout(n1321),.clk(gclk));
	jand g1059(.dina(w_n1321_1[1]),.dinb(w_n323_61[2]),.dout(n1322),.clk(gclk));
	jor g1060(.dina(w_n684_0[0]),.dinb(w_shift1_45[1]),.dout(n1323),.clk(gclk));
	jor g1061(.dina(w_n542_0[0]),.dinb(w_n269_45[1]),.dout(n1324),.clk(gclk));
	jand g1062(.dina(n1324),.dinb(n1323),.dout(n1325),.clk(gclk));
	jand g1063(.dina(w_n549_0[0]),.dinb(w_shift1_45[0]),.dout(n1326),.clk(gclk));
	jand g1064(.dina(w_n687_0[0]),.dinb(w_n269_45[0]),.dout(n1327),.clk(gclk));
	jor g1065(.dina(n1327),.dinb(n1326),.dout(n1328),.clk(gclk));
	jor g1066(.dina(n1328),.dinb(n1325),.dout(n1329),.clk(gclk));
	jand g1067(.dina(w_n1329_1[1]),.dinb(w_n266_55[2]),.dout(n1330),.clk(gclk));
	jor g1068(.dina(w_n555_0[0]),.dinb(w_n269_44[2]),.dout(n1331),.clk(gclk));
	jor g1069(.dina(w_n570_0[0]),.dinb(w_shift1_44[2]),.dout(n1332),.clk(gclk));
	jand g1070(.dina(n1332),.dinb(n1331),.dout(n1333),.clk(gclk));
	jand g1071(.dina(w_n554_0[0]),.dinb(w_shift1_44[1]),.dout(n1334),.clk(gclk));
	jand g1072(.dina(w_n567_0[0]),.dinb(w_n269_44[1]),.dout(n1335),.clk(gclk));
	jor g1073(.dina(n1335),.dinb(n1334),.dout(n1336),.clk(gclk));
	jor g1074(.dina(n1336),.dinb(n1333),.dout(n1337),.clk(gclk));
	jand g1075(.dina(w_n1337_1[1]),.dinb(w_n281_55[2]),.dout(n1338),.clk(gclk));
	jor g1076(.dina(n1338),.dinb(n1330),.dout(n1339),.clk(gclk));
	jor g1077(.dina(w_n547_0[0]),.dinb(w_shift1_44[0]),.dout(n1340),.clk(gclk));
	jor g1078(.dina(w_n572_0[0]),.dinb(w_n269_44[0]),.dout(n1341),.clk(gclk));
	jand g1079(.dina(n1341),.dinb(n1340),.dout(n1342),.clk(gclk));
	jand g1080(.dina(w_n565_0[0]),.dinb(w_shift1_43[2]),.dout(n1343),.clk(gclk));
	jand g1081(.dina(w_n544_0[0]),.dinb(w_n269_43[2]),.dout(n1344),.clk(gclk));
	jor g1082(.dina(n1344),.dinb(n1343),.dout(n1345),.clk(gclk));
	jor g1083(.dina(n1345),.dinb(n1342),.dout(n1346),.clk(gclk));
	jand g1084(.dina(w_n1346_1[1]),.dinb(w_n295_55[2]),.dout(n1347),.clk(gclk));
	jor g1085(.dina(w_n558_0[0]),.dinb(w_shift1_43[1]),.dout(n1348),.clk(gclk));
	jor g1086(.dina(w_n577_0[0]),.dinb(w_n269_43[1]),.dout(n1349),.clk(gclk));
	jand g1087(.dina(n1349),.dinb(n1348),.dout(n1350),.clk(gclk));
	jand g1088(.dina(w_n584_0[0]),.dinb(w_shift1_43[0]),.dout(n1351),.clk(gclk));
	jand g1089(.dina(w_n559_0[0]),.dinb(w_n269_43[0]),.dout(n1352),.clk(gclk));
	jor g1090(.dina(n1352),.dinb(n1351),.dout(n1353),.clk(gclk));
	jor g1091(.dina(n1353),.dinb(n1350),.dout(n1354),.clk(gclk));
	jand g1092(.dina(w_n1354_1[1]),.dinb(w_n308_55[2]),.dout(n1355),.clk(gclk));
	jor g1093(.dina(n1355),.dinb(n1347),.dout(n1356),.clk(gclk));
	jor g1094(.dina(n1356),.dinb(n1339),.dout(n1357),.clk(gclk));
	jand g1095(.dina(w_n1357_1[1]),.dinb(w_n377_61[2]),.dout(n1358),.clk(gclk));
	jor g1096(.dina(n1358),.dinb(n1322),.dout(n1359),.clk(gclk));
	jor g1097(.dina(n1359),.dinb(n1286),.dout(n1360),.clk(gclk));
	jand g1098(.dina(w_n1360_0[1]),.dinb(w_shift6_62[2]),.dout(n1361),.clk(gclk));
	jor g1099(.dina(n1361),.dinb(n1213),.dout(result2),.clk(gclk));
	jor g1100(.dina(w_n751_0[0]),.dinb(w_n269_42[2]),.dout(n1363),.clk(gclk));
	jor g1101(.dina(w_n867_0[0]),.dinb(w_shift1_42[2]),.dout(n1364),.clk(gclk));
	jand g1102(.dina(n1364),.dinb(n1363),.dout(n1365),.clk(gclk));
	jand g1103(.dina(w_n1365_1[1]),.dinb(w_n266_55[1]),.dout(n1366),.clk(gclk));
	jor g1104(.dina(w_n761_0[0]),.dinb(w_n269_42[1]),.dout(n1367),.clk(gclk));
	jor g1105(.dina(w_n768_0[0]),.dinb(w_shift1_42[1]),.dout(n1368),.clk(gclk));
	jand g1106(.dina(n1368),.dinb(n1367),.dout(n1369),.clk(gclk));
	jand g1107(.dina(w_n1369_1[1]),.dinb(w_n281_55[1]),.dout(n1370),.clk(gclk));
	jor g1108(.dina(n1370),.dinb(n1366),.dout(n1371),.clk(gclk));
	jor g1109(.dina(w_n772_0[0]),.dinb(w_n269_42[0]),.dout(n1372),.clk(gclk));
	jor g1110(.dina(w_n747_0[0]),.dinb(w_shift1_42[0]),.dout(n1373),.clk(gclk));
	jand g1111(.dina(n1373),.dinb(n1372),.dout(n1374),.clk(gclk));
	jand g1112(.dina(w_n1374_1[1]),.dinb(w_n295_55[1]),.dout(n1375),.clk(gclk));
	jor g1113(.dina(w_n782_0[0]),.dinb(w_n269_41[2]),.dout(n1376),.clk(gclk));
	jor g1114(.dina(w_n757_0[0]),.dinb(w_shift1_41[2]),.dout(n1377),.clk(gclk));
	jand g1115(.dina(n1377),.dinb(n1376),.dout(n1378),.clk(gclk));
	jand g1116(.dina(w_n1378_1[1]),.dinb(w_n308_55[1]),.dout(n1379),.clk(gclk));
	jor g1117(.dina(n1379),.dinb(n1375),.dout(n1380),.clk(gclk));
	jor g1118(.dina(n1380),.dinb(n1371),.dout(n1381),.clk(gclk));
	jand g1119(.dina(w_n1381_1[1]),.dinb(w_n377_61[1]),.dout(n1382),.clk(gclk));
	jor g1120(.dina(w_n707_0[0]),.dinb(w_n269_41[1]),.dout(n1383),.clk(gclk));
	jor g1121(.dina(w_n823_0[0]),.dinb(w_shift1_41[1]),.dout(n1384),.clk(gclk));
	jand g1122(.dina(n1384),.dinb(n1383),.dout(n1385),.clk(gclk));
	jand g1123(.dina(w_n1385_1[1]),.dinb(w_n266_55[0]),.dout(n1386),.clk(gclk));
	jor g1124(.dina(w_n717_0[0]),.dinb(w_n269_41[0]),.dout(n1387),.clk(gclk));
	jor g1125(.dina(w_n724_0[0]),.dinb(w_shift1_41[0]),.dout(n1388),.clk(gclk));
	jand g1126(.dina(n1388),.dinb(n1387),.dout(n1389),.clk(gclk));
	jand g1127(.dina(w_n1389_1[1]),.dinb(w_n281_55[0]),.dout(n1390),.clk(gclk));
	jor g1128(.dina(n1390),.dinb(n1386),.dout(n1391),.clk(gclk));
	jor g1129(.dina(w_n728_0[0]),.dinb(w_n269_40[2]),.dout(n1392),.clk(gclk));
	jor g1130(.dina(w_n703_0[0]),.dinb(w_shift1_40[2]),.dout(n1393),.clk(gclk));
	jand g1131(.dina(n1393),.dinb(n1392),.dout(n1394),.clk(gclk));
	jand g1132(.dina(w_n1394_1[1]),.dinb(w_n295_55[0]),.dout(n1395),.clk(gclk));
	jor g1133(.dina(w_n738_0[0]),.dinb(w_n269_40[1]),.dout(n1396),.clk(gclk));
	jor g1134(.dina(w_n713_0[0]),.dinb(w_shift1_40[1]),.dout(n1397),.clk(gclk));
	jand g1135(.dina(n1397),.dinb(n1396),.dout(n1398),.clk(gclk));
	jand g1136(.dina(w_n1398_1[1]),.dinb(w_n308_55[0]),.dout(n1399),.clk(gclk));
	jor g1137(.dina(n1399),.dinb(n1395),.dout(n1400),.clk(gclk));
	jor g1138(.dina(n1400),.dinb(n1391),.dout(n1401),.clk(gclk));
	jand g1139(.dina(w_n1401_1[1]),.dinb(w_n323_61[1]),.dout(n1402),.clk(gclk));
	jor g1140(.dina(n1402),.dinb(n1382),.dout(n1403),.clk(gclk));
	jor g1141(.dina(w_n796_0[0]),.dinb(w_n269_40[0]),.dout(n1404),.clk(gclk));
	jor g1142(.dina(w_n778_0[0]),.dinb(w_shift1_40[0]),.dout(n1405),.clk(gclk));
	jand g1143(.dina(n1405),.dinb(n1404),.dout(n1406),.clk(gclk));
	jand g1144(.dina(w_n1406_1[1]),.dinb(w_n266_54[2]),.dout(n1407),.clk(gclk));
	jor g1145(.dina(w_n806_0[0]),.dinb(w_n269_39[2]),.dout(n1408),.clk(gclk));
	jor g1146(.dina(w_n813_0[0]),.dinb(w_shift1_39[2]),.dout(n1409),.clk(gclk));
	jand g1147(.dina(n1409),.dinb(n1408),.dout(n1410),.clk(gclk));
	jand g1148(.dina(w_n1410_1[1]),.dinb(w_n281_54[2]),.dout(n1411),.clk(gclk));
	jor g1149(.dina(n1411),.dinb(n1407),.dout(n1412),.clk(gclk));
	jor g1150(.dina(w_n817_0[0]),.dinb(w_n269_39[1]),.dout(n1413),.clk(gclk));
	jor g1151(.dina(w_n792_0[0]),.dinb(w_shift1_39[1]),.dout(n1414),.clk(gclk));
	jand g1152(.dina(n1414),.dinb(n1413),.dout(n1415),.clk(gclk));
	jand g1153(.dina(w_n1415_1[1]),.dinb(w_n295_54[2]),.dout(n1416),.clk(gclk));
	jor g1154(.dina(w_n827_0[0]),.dinb(w_n269_39[0]),.dout(n1417),.clk(gclk));
	jor g1155(.dina(w_n802_0[0]),.dinb(w_shift1_39[0]),.dout(n1418),.clk(gclk));
	jand g1156(.dina(n1418),.dinb(n1417),.dout(n1419),.clk(gclk));
	jand g1157(.dina(w_n1419_1[1]),.dinb(w_n308_54[2]),.dout(n1420),.clk(gclk));
	jor g1158(.dina(n1420),.dinb(n1416),.dout(n1421),.clk(gclk));
	jor g1159(.dina(n1421),.dinb(n1412),.dout(n1422),.clk(gclk));
	jand g1160(.dina(w_n1422_1[1]),.dinb(w_n432_61[1]),.dout(n1423),.clk(gclk));
	jor g1161(.dina(w_n840_0[0]),.dinb(w_n269_38[2]),.dout(n1424),.clk(gclk));
	jor g1162(.dina(w_n1003_0[0]),.dinb(w_shift1_38[2]),.dout(n1425),.clk(gclk));
	jand g1163(.dina(n1425),.dinb(n1424),.dout(n1426),.clk(gclk));
	jand g1164(.dina(w_n1426_1[1]),.dinb(w_n266_54[1]),.dout(n1427),.clk(gclk));
	jor g1165(.dina(w_n850_0[0]),.dinb(w_n269_38[1]),.dout(n1428),.clk(gclk));
	jor g1166(.dina(w_n857_0[0]),.dinb(w_shift1_38[1]),.dout(n1429),.clk(gclk));
	jand g1167(.dina(n1429),.dinb(n1428),.dout(n1430),.clk(gclk));
	jand g1168(.dina(w_n1430_1[1]),.dinb(w_n281_54[1]),.dout(n1431),.clk(gclk));
	jor g1169(.dina(n1431),.dinb(n1427),.dout(n1432),.clk(gclk));
	jor g1170(.dina(w_n861_0[0]),.dinb(w_n269_38[0]),.dout(n1433),.clk(gclk));
	jor g1171(.dina(w_n836_0[0]),.dinb(w_shift1_38[0]),.dout(n1434),.clk(gclk));
	jand g1172(.dina(n1434),.dinb(n1433),.dout(n1435),.clk(gclk));
	jand g1173(.dina(w_n1435_1[1]),.dinb(w_n295_54[1]),.dout(n1436),.clk(gclk));
	jor g1174(.dina(w_n871_0[0]),.dinb(w_n269_37[2]),.dout(n1437),.clk(gclk));
	jor g1175(.dina(w_n846_0[0]),.dinb(w_shift1_37[2]),.dout(n1438),.clk(gclk));
	jand g1176(.dina(n1438),.dinb(n1437),.dout(n1439),.clk(gclk));
	jand g1177(.dina(w_n1439_1[1]),.dinb(w_n308_54[1]),.dout(n1440),.clk(gclk));
	jor g1178(.dina(n1440),.dinb(n1436),.dout(n1441),.clk(gclk));
	jor g1179(.dina(n1441),.dinb(n1432),.dout(n1442),.clk(gclk));
	jand g1180(.dina(w_n1442_1[1]),.dinb(w_n485_61[1]),.dout(n1443),.clk(gclk));
	jor g1181(.dina(n1443),.dinb(n1423),.dout(n1444),.clk(gclk));
	jor g1182(.dina(n1444),.dinb(n1403),.dout(n1445),.clk(gclk));
	jand g1183(.dina(w_n1445_0[1]),.dinb(w_n263_62[1]),.dout(n1446),.clk(gclk));
	jor g1184(.dina(w_n887_0[0]),.dinb(w_n269_37[1]),.dout(n1447),.clk(gclk));
	jor g1185(.dina(w_n734_0[0]),.dinb(w_shift1_37[1]),.dout(n1448),.clk(gclk));
	jand g1186(.dina(n1448),.dinb(n1447),.dout(n1449),.clk(gclk));
	jand g1187(.dina(w_n1449_1[1]),.dinb(w_n266_54[0]),.dout(n1450),.clk(gclk));
	jor g1188(.dina(w_n897_0[0]),.dinb(w_n269_37[0]),.dout(n1451),.clk(gclk));
	jor g1189(.dina(w_n904_0[0]),.dinb(w_shift1_37[0]),.dout(n1452),.clk(gclk));
	jand g1190(.dina(n1452),.dinb(n1451),.dout(n1453),.clk(gclk));
	jand g1191(.dina(w_n1453_1[1]),.dinb(w_n281_54[0]),.dout(n1454),.clk(gclk));
	jor g1192(.dina(n1454),.dinb(n1450),.dout(n1455),.clk(gclk));
	jor g1193(.dina(w_n908_0[0]),.dinb(w_n269_36[2]),.dout(n1456),.clk(gclk));
	jor g1194(.dina(w_n883_0[0]),.dinb(w_shift1_36[2]),.dout(n1457),.clk(gclk));
	jand g1195(.dina(n1457),.dinb(n1456),.dout(n1458),.clk(gclk));
	jand g1196(.dina(w_n1458_1[1]),.dinb(w_n295_54[0]),.dout(n1459),.clk(gclk));
	jor g1197(.dina(w_n918_0[0]),.dinb(w_n269_36[1]),.dout(n1460),.clk(gclk));
	jor g1198(.dina(w_n893_0[0]),.dinb(w_shift1_36[1]),.dout(n1461),.clk(gclk));
	jand g1199(.dina(n1461),.dinb(n1460),.dout(n1462),.clk(gclk));
	jand g1200(.dina(w_n1462_1[1]),.dinb(w_n308_54[0]),.dout(n1463),.clk(gclk));
	jor g1201(.dina(n1463),.dinb(n1459),.dout(n1464),.clk(gclk));
	jor g1202(.dina(n1464),.dinb(n1455),.dout(n1465),.clk(gclk));
	jand g1203(.dina(w_n1465_1[1]),.dinb(w_n485_61[0]),.dout(n1466),.clk(gclk));
	jor g1204(.dina(w_n931_0[0]),.dinb(w_n269_36[0]),.dout(n1467),.clk(gclk));
	jor g1205(.dina(w_n1051_0[0]),.dinb(w_shift1_36[0]),.dout(n1468),.clk(gclk));
	jand g1206(.dina(n1468),.dinb(n1467),.dout(n1469),.clk(gclk));
	jand g1207(.dina(w_n1469_1[1]),.dinb(w_n266_53[2]),.dout(n1470),.clk(gclk));
	jor g1208(.dina(w_n941_0[0]),.dinb(w_n269_35[2]),.dout(n1471),.clk(gclk));
	jor g1209(.dina(w_n948_0[0]),.dinb(w_shift1_35[2]),.dout(n1472),.clk(gclk));
	jand g1210(.dina(n1472),.dinb(n1471),.dout(n1473),.clk(gclk));
	jand g1211(.dina(w_n1473_1[1]),.dinb(w_n281_53[2]),.dout(n1474),.clk(gclk));
	jor g1212(.dina(n1474),.dinb(n1470),.dout(n1475),.clk(gclk));
	jor g1213(.dina(w_n952_0[0]),.dinb(w_n269_35[1]),.dout(n1476),.clk(gclk));
	jor g1214(.dina(w_n927_0[0]),.dinb(w_shift1_35[1]),.dout(n1477),.clk(gclk));
	jand g1215(.dina(n1477),.dinb(n1476),.dout(n1478),.clk(gclk));
	jand g1216(.dina(w_n1478_1[1]),.dinb(w_n295_53[2]),.dout(n1479),.clk(gclk));
	jor g1217(.dina(w_n962_0[0]),.dinb(w_n269_35[0]),.dout(n1480),.clk(gclk));
	jor g1218(.dina(w_n937_0[0]),.dinb(w_shift1_35[0]),.dout(n1481),.clk(gclk));
	jand g1219(.dina(n1481),.dinb(n1480),.dout(n1482),.clk(gclk));
	jand g1220(.dina(w_n1482_1[1]),.dinb(w_n308_53[2]),.dout(n1483),.clk(gclk));
	jor g1221(.dina(n1483),.dinb(n1479),.dout(n1484),.clk(gclk));
	jor g1222(.dina(n1484),.dinb(n1475),.dout(n1485),.clk(gclk));
	jand g1223(.dina(w_n1485_1[1]),.dinb(w_n432_61[0]),.dout(n1486),.clk(gclk));
	jor g1224(.dina(n1486),.dinb(n1466),.dout(n1487),.clk(gclk));
	jor g1225(.dina(w_n1016_0[0]),.dinb(w_n269_34[2]),.dout(n1488),.clk(gclk));
	jor g1226(.dina(w_n914_0[0]),.dinb(w_shift1_34[2]),.dout(n1489),.clk(gclk));
	jand g1227(.dina(n1489),.dinb(n1488),.dout(n1490),.clk(gclk));
	jand g1228(.dina(w_n1490_1[1]),.dinb(w_n266_53[1]),.dout(n1491),.clk(gclk));
	jor g1229(.dina(w_n1031_0[0]),.dinb(w_n1026_0[0]),.dout(n1492),.clk(gclk));
	jand g1230(.dina(n1492),.dinb(w_shift1_34[1]),.dout(n1493),.clk(gclk));
	jor g1231(.dina(w_n1042_0[0]),.dinb(w_n1039_0[0]),.dout(n1494),.clk(gclk));
	jand g1232(.dina(n1494),.dinb(w_n269_34[1]),.dout(n1495),.clk(gclk));
	jor g1233(.dina(n1495),.dinb(n1493),.dout(n1496),.clk(gclk));
	jand g1234(.dina(w_n1496_1[1]),.dinb(w_n281_53[1]),.dout(n1497),.clk(gclk));
	jor g1235(.dina(n1497),.dinb(n1491),.dout(n1498),.clk(gclk));
	jor g1236(.dina(w_n1019_0[0]),.dinb(w_shift1_34[0]),.dout(n1499),.clk(gclk));
	jor g1237(.dina(w_n1044_0[0]),.dinb(w_n269_34[0]),.dout(n1500),.clk(gclk));
	jand g1238(.dina(n1500),.dinb(n1499),.dout(n1501),.clk(gclk));
	jand g1239(.dina(w_n1037_0[0]),.dinb(w_shift1_33[2]),.dout(n1502),.clk(gclk));
	jand g1240(.dina(w_n1018_0[0]),.dinb(w_n269_33[2]),.dout(n1503),.clk(gclk));
	jor g1241(.dina(n1503),.dinb(n1502),.dout(n1504),.clk(gclk));
	jor g1242(.dina(n1504),.dinb(n1501),.dout(n1505),.clk(gclk));
	jand g1243(.dina(w_n1505_1[1]),.dinb(w_n295_53[1]),.dout(n1506),.clk(gclk));
	jand g1244(.dina(w_n1055_0[0]),.dinb(w_shift1_33[1]),.dout(n1507),.clk(gclk));
	jor g1245(.dina(w_n1029_0[0]),.dinb(w_n1024_0[0]),.dout(n1508),.clk(gclk));
	jand g1246(.dina(n1508),.dinb(w_n269_33[1]),.dout(n1509),.clk(gclk));
	jor g1247(.dina(n1509),.dinb(n1507),.dout(n1510),.clk(gclk));
	jand g1248(.dina(w_n1510_1[1]),.dinb(w_n308_53[1]),.dout(n1511),.clk(gclk));
	jor g1249(.dina(n1511),.dinb(n1506),.dout(n1512),.clk(gclk));
	jor g1250(.dina(n1512),.dinb(n1498),.dout(n1513),.clk(gclk));
	jand g1251(.dina(w_n1513_1[1]),.dinb(w_n377_61[0]),.dout(n1514),.clk(gclk));
	jor g1252(.dina(w_n976_0[0]),.dinb(w_n269_33[0]),.dout(n1515),.clk(gclk));
	jor g1253(.dina(w_n958_0[0]),.dinb(w_shift1_33[0]),.dout(n1516),.clk(gclk));
	jand g1254(.dina(n1516),.dinb(n1515),.dout(n1517),.clk(gclk));
	jand g1255(.dina(w_n1517_1[1]),.dinb(w_n266_53[0]),.dout(n1518),.clk(gclk));
	jor g1256(.dina(w_n986_0[0]),.dinb(w_n269_32[2]),.dout(n1519),.clk(gclk));
	jor g1257(.dina(w_n993_0[0]),.dinb(w_shift1_32[2]),.dout(n1520),.clk(gclk));
	jand g1258(.dina(n1520),.dinb(n1519),.dout(n1521),.clk(gclk));
	jand g1259(.dina(w_n1521_1[1]),.dinb(w_n281_53[0]),.dout(n1522),.clk(gclk));
	jor g1260(.dina(n1522),.dinb(n1518),.dout(n1523),.clk(gclk));
	jor g1261(.dina(w_n997_0[0]),.dinb(w_n269_32[1]),.dout(n1524),.clk(gclk));
	jor g1262(.dina(w_n972_0[0]),.dinb(w_shift1_32[1]),.dout(n1525),.clk(gclk));
	jand g1263(.dina(n1525),.dinb(n1524),.dout(n1526),.clk(gclk));
	jand g1264(.dina(w_n1526_1[1]),.dinb(w_n295_53[0]),.dout(n1527),.clk(gclk));
	jor g1265(.dina(w_n1007_0[0]),.dinb(w_n269_32[0]),.dout(n1528),.clk(gclk));
	jor g1266(.dina(w_n982_0[0]),.dinb(w_shift1_32[0]),.dout(n1529),.clk(gclk));
	jand g1267(.dina(n1529),.dinb(n1528),.dout(n1530),.clk(gclk));
	jand g1268(.dina(w_n1530_1[1]),.dinb(w_n308_53[0]),.dout(n1531),.clk(gclk));
	jor g1269(.dina(n1531),.dinb(n1527),.dout(n1532),.clk(gclk));
	jor g1270(.dina(n1532),.dinb(n1523),.dout(n1533),.clk(gclk));
	jand g1271(.dina(w_n1533_1[1]),.dinb(w_n323_61[0]),.dout(n1534),.clk(gclk));
	jor g1272(.dina(n1534),.dinb(n1514),.dout(n1535),.clk(gclk));
	jor g1273(.dina(n1535),.dinb(n1487),.dout(n1536),.clk(gclk));
	jand g1274(.dina(w_n1536_0[1]),.dinb(w_shift6_62[1]),.dout(n1537),.clk(gclk));
	jor g1275(.dina(n1537),.dinb(n1446),.dout(result3),.clk(gclk));
	jand g1276(.dina(w_n427_1[0]),.dinb(w_n266_52[2]),.dout(n1539),.clk(gclk));
	jand g1277(.dina(w_n306_1[0]),.dinb(w_n281_52[2]),.dout(n1540),.clk(gclk));
	jor g1278(.dina(n1540),.dinb(n1539),.dout(n1541),.clk(gclk));
	jand g1279(.dina(w_n295_52[2]),.dinb(w_n279_1[0]),.dout(n1542),.clk(gclk));
	jand g1280(.dina(w_n308_52[2]),.dinb(w_n292_1[0]),.dout(n1543),.clk(gclk));
	jor g1281(.dina(n1543),.dinb(n1542),.dout(n1544),.clk(gclk));
	jor g1282(.dina(n1544),.dinb(n1541),.dout(n1545),.clk(gclk));
	jand g1283(.dina(w_n1545_1[1]),.dinb(w_n323_60[2]),.dout(n1546),.clk(gclk));
	jand g1284(.dina(w_n481_1[0]),.dinb(w_n266_52[1]),.dout(n1547),.clk(gclk));
	jand g1285(.dina(w_n360_1[0]),.dinb(w_n281_52[1]),.dout(n1548),.clk(gclk));
	jor g1286(.dina(n1548),.dinb(n1547),.dout(n1549),.clk(gclk));
	jand g1287(.dina(w_n335_1[0]),.dinb(w_n295_52[1]),.dout(n1550),.clk(gclk));
	jand g1288(.dina(w_n347_1[0]),.dinb(w_n308_52[1]),.dout(n1551),.clk(gclk));
	jor g1289(.dina(n1551),.dinb(n1550),.dout(n1552),.clk(gclk));
	jor g1290(.dina(n1552),.dinb(n1549),.dout(n1553),.clk(gclk));
	jand g1291(.dina(w_n1553_1[1]),.dinb(w_n377_60[2]),.dout(n1554),.clk(gclk));
	jor g1292(.dina(n1554),.dinb(n1546),.dout(n1555),.clk(gclk));
	jand g1293(.dina(w_n372_1[0]),.dinb(w_n266_52[0]),.dout(n1556),.clk(gclk));
	jand g1294(.dina(w_n415_1[0]),.dinb(w_n281_52[0]),.dout(n1557),.clk(gclk));
	jor g1295(.dina(n1557),.dinb(n1556),.dout(n1558),.clk(gclk));
	jand g1296(.dina(w_n390_1[0]),.dinb(w_n295_52[0]),.dout(n1559),.clk(gclk));
	jand g1297(.dina(w_n402_1[0]),.dinb(w_n308_52[0]),.dout(n1560),.clk(gclk));
	jor g1298(.dina(n1560),.dinb(n1559),.dout(n1561),.clk(gclk));
	jor g1299(.dina(n1561),.dinb(n1558),.dout(n1562),.clk(gclk));
	jand g1300(.dina(w_n1562_1[1]),.dinb(w_n432_60[2]),.dout(n1563),.clk(gclk));
	jand g1301(.dina(w_n537_1[0]),.dinb(w_n266_51[2]),.dout(n1564),.clk(gclk));
	jand g1302(.dina(w_n469_1[0]),.dinb(w_n281_51[2]),.dout(n1565),.clk(gclk));
	jor g1303(.dina(n1565),.dinb(n1564),.dout(n1566),.clk(gclk));
	jand g1304(.dina(w_n444_1[0]),.dinb(w_n295_51[2]),.dout(n1567),.clk(gclk));
	jand g1305(.dina(w_n456_1[0]),.dinb(w_n308_51[2]),.dout(n1568),.clk(gclk));
	jor g1306(.dina(n1568),.dinb(n1567),.dout(n1569),.clk(gclk));
	jor g1307(.dina(n1569),.dinb(n1566),.dout(n1570),.clk(gclk));
	jand g1308(.dina(w_n1570_1[1]),.dinb(w_n485_60[2]),.dout(n1571),.clk(gclk));
	jor g1309(.dina(n1571),.dinb(n1563),.dout(n1572),.clk(gclk));
	jor g1310(.dina(n1572),.dinb(n1555),.dout(n1573),.clk(gclk));
	jand g1311(.dina(w_n1573_0[1]),.dinb(w_n263_62[0]),.dout(n1574),.clk(gclk));
	jand g1312(.dina(w_n692_1[0]),.dinb(w_n266_51[1]),.dout(n1575),.clk(gclk));
	jand g1313(.dina(w_n575_1[0]),.dinb(w_n281_51[1]),.dout(n1576),.clk(gclk));
	jor g1314(.dina(n1576),.dinb(n1575),.dout(n1577),.clk(gclk));
	jand g1315(.dina(w_n552_1[0]),.dinb(w_n295_51[1]),.dout(n1578),.clk(gclk));
	jand g1316(.dina(w_n562_1[0]),.dinb(w_n308_51[1]),.dout(n1579),.clk(gclk));
	jor g1317(.dina(n1579),.dinb(n1578),.dout(n1580),.clk(gclk));
	jor g1318(.dina(n1580),.dinb(n1577),.dout(n1581),.clk(gclk));
	jand g1319(.dina(w_n1581_1[1]),.dinb(w_n377_60[1]),.dout(n1582),.clk(gclk));
	jand g1320(.dina(w_n640_1[0]),.dinb(w_n266_51[0]),.dout(n1583),.clk(gclk));
	jand g1321(.dina(w_n525_1[0]),.dinb(w_n281_51[0]),.dout(n1584),.clk(gclk));
	jor g1322(.dina(n1584),.dinb(n1583),.dout(n1585),.clk(gclk));
	jand g1323(.dina(w_n500_1[0]),.dinb(w_n295_51[0]),.dout(n1586),.clk(gclk));
	jand g1324(.dina(w_n512_1[0]),.dinb(w_n308_51[0]),.dout(n1587),.clk(gclk));
	jor g1325(.dina(n1587),.dinb(n1586),.dout(n1588),.clk(gclk));
	jor g1326(.dina(n1588),.dinb(n1585),.dout(n1589),.clk(gclk));
	jand g1327(.dina(w_n1589_1[1]),.dinb(w_n323_60[1]),.dout(n1590),.clk(gclk));
	jor g1328(.dina(n1590),.dinb(n1582),.dout(n1591),.clk(gclk));
	jand g1329(.dina(w_n319_1[0]),.dinb(w_n266_50[2]),.dout(n1592),.clk(gclk));
	jand g1330(.dina(w_n680_1[0]),.dinb(w_n281_50[2]),.dout(n1593),.clk(gclk));
	jor g1331(.dina(n1593),.dinb(n1592),.dout(n1594),.clk(gclk));
	jand g1332(.dina(w_n655_1[0]),.dinb(w_n295_50[2]),.dout(n1595),.clk(gclk));
	jand g1333(.dina(w_n667_1[0]),.dinb(w_n308_50[2]),.dout(n1596),.clk(gclk));
	jor g1334(.dina(n1596),.dinb(n1595),.dout(n1597),.clk(gclk));
	jor g1335(.dina(n1597),.dinb(n1594),.dout(n1598),.clk(gclk));
	jand g1336(.dina(w_n1598_1[1]),.dinb(w_n485_60[1]),.dout(n1599),.clk(gclk));
	jand g1337(.dina(w_n587_1[0]),.dinb(w_n266_50[1]),.dout(n1600),.clk(gclk));
	jand g1338(.dina(w_n628_1[0]),.dinb(w_n281_50[1]),.dout(n1601),.clk(gclk));
	jor g1339(.dina(n1601),.dinb(n1600),.dout(n1602),.clk(gclk));
	jand g1340(.dina(w_n603_1[0]),.dinb(w_n295_50[1]),.dout(n1603),.clk(gclk));
	jand g1341(.dina(w_n615_1[0]),.dinb(w_n308_50[1]),.dout(n1604),.clk(gclk));
	jor g1342(.dina(n1604),.dinb(n1603),.dout(n1605),.clk(gclk));
	jor g1343(.dina(n1605),.dinb(n1602),.dout(n1606),.clk(gclk));
	jand g1344(.dina(w_n1606_1[1]),.dinb(w_n432_60[1]),.dout(n1607),.clk(gclk));
	jor g1345(.dina(n1607),.dinb(n1599),.dout(n1608),.clk(gclk));
	jor g1346(.dina(n1608),.dinb(n1591),.dout(n1609),.clk(gclk));
	jand g1347(.dina(w_n1609_0[1]),.dinb(w_shift6_62[0]),.dout(n1610),.clk(gclk));
	jor g1348(.dina(n1610),.dinb(n1574),.dout(result4),.clk(gclk));
	jand g1349(.dina(w_n829_1[0]),.dinb(w_n266_50[0]),.dout(n1612),.clk(gclk));
	jand g1350(.dina(w_n730_1[0]),.dinb(w_n281_50[0]),.dout(n1613),.clk(gclk));
	jor g1351(.dina(n1613),.dinb(n1612),.dout(n1614),.clk(gclk));
	jand g1352(.dina(w_n709_1[0]),.dinb(w_n295_50[0]),.dout(n1615),.clk(gclk));
	jand g1353(.dina(w_n719_1[0]),.dinb(w_n308_50[0]),.dout(n1616),.clk(gclk));
	jor g1354(.dina(n1616),.dinb(n1615),.dout(n1617),.clk(gclk));
	jor g1355(.dina(n1617),.dinb(n1614),.dout(n1618),.clk(gclk));
	jand g1356(.dina(w_n1618_1[1]),.dinb(w_n323_60[0]),.dout(n1619),.clk(gclk));
	jand g1357(.dina(w_n873_1[0]),.dinb(w_n266_49[2]),.dout(n1620),.clk(gclk));
	jand g1358(.dina(w_n774_1[0]),.dinb(w_n281_49[2]),.dout(n1621),.clk(gclk));
	jor g1359(.dina(n1621),.dinb(n1620),.dout(n1622),.clk(gclk));
	jand g1360(.dina(w_n753_1[0]),.dinb(w_n295_49[2]),.dout(n1623),.clk(gclk));
	jand g1361(.dina(w_n763_1[0]),.dinb(w_n308_49[2]),.dout(n1624),.clk(gclk));
	jor g1362(.dina(n1624),.dinb(n1623),.dout(n1625),.clk(gclk));
	jor g1363(.dina(n1625),.dinb(n1622),.dout(n1626),.clk(gclk));
	jand g1364(.dina(w_n1626_1[1]),.dinb(w_n377_60[0]),.dout(n1627),.clk(gclk));
	jor g1365(.dina(n1627),.dinb(n1619),.dout(n1628),.clk(gclk));
	jand g1366(.dina(w_n784_1[0]),.dinb(w_n266_49[1]),.dout(n1629),.clk(gclk));
	jand g1367(.dina(w_n819_1[0]),.dinb(w_n281_49[1]),.dout(n1630),.clk(gclk));
	jor g1368(.dina(n1630),.dinb(n1629),.dout(n1631),.clk(gclk));
	jand g1369(.dina(w_n798_1[0]),.dinb(w_n295_49[1]),.dout(n1632),.clk(gclk));
	jand g1370(.dina(w_n808_1[0]),.dinb(w_n308_49[1]),.dout(n1633),.clk(gclk));
	jor g1371(.dina(n1633),.dinb(n1632),.dout(n1634),.clk(gclk));
	jor g1372(.dina(n1634),.dinb(n1631),.dout(n1635),.clk(gclk));
	jand g1373(.dina(w_n1635_1[1]),.dinb(w_n432_60[0]),.dout(n1636),.clk(gclk));
	jand g1374(.dina(w_n1009_1[0]),.dinb(w_n266_49[0]),.dout(n1637),.clk(gclk));
	jand g1375(.dina(w_n863_1[0]),.dinb(w_n281_49[0]),.dout(n1638),.clk(gclk));
	jor g1376(.dina(n1638),.dinb(n1637),.dout(n1639),.clk(gclk));
	jand g1377(.dina(w_n842_1[0]),.dinb(w_n295_49[0]),.dout(n1640),.clk(gclk));
	jand g1378(.dina(w_n852_1[0]),.dinb(w_n308_49[0]),.dout(n1641),.clk(gclk));
	jor g1379(.dina(n1641),.dinb(n1640),.dout(n1642),.clk(gclk));
	jor g1380(.dina(n1642),.dinb(n1639),.dout(n1643),.clk(gclk));
	jand g1381(.dina(w_n1643_1[1]),.dinb(w_n485_60[0]),.dout(n1644),.clk(gclk));
	jor g1382(.dina(n1644),.dinb(n1636),.dout(n1645),.clk(gclk));
	jor g1383(.dina(n1645),.dinb(n1628),.dout(n1646),.clk(gclk));
	jand g1384(.dina(w_n1646_0[1]),.dinb(w_n263_61[2]),.dout(n1647),.clk(gclk));
	jand g1385(.dina(w_n920_1[0]),.dinb(w_n266_48[2]),.dout(n1648),.clk(gclk));
	jand g1386(.dina(w_n1047_1[0]),.dinb(w_n281_48[2]),.dout(n1649),.clk(gclk));
	jor g1387(.dina(n1649),.dinb(n1648),.dout(n1650),.clk(gclk));
	jand g1388(.dina(w_n1022_1[0]),.dinb(w_n295_48[2]),.dout(n1651),.clk(gclk));
	jand g1389(.dina(w_n1034_1[0]),.dinb(w_n308_48[2]),.dout(n1652),.clk(gclk));
	jor g1390(.dina(n1652),.dinb(n1651),.dout(n1653),.clk(gclk));
	jor g1391(.dina(n1653),.dinb(n1650),.dout(n1654),.clk(gclk));
	jand g1392(.dina(w_n1654_1[1]),.dinb(w_n377_59[2]),.dout(n1655),.clk(gclk));
	jand g1393(.dina(w_n964_1[0]),.dinb(w_n266_48[1]),.dout(n1656),.clk(gclk));
	jand g1394(.dina(w_n999_1[0]),.dinb(w_n281_48[1]),.dout(n1657),.clk(gclk));
	jor g1395(.dina(n1657),.dinb(n1656),.dout(n1658),.clk(gclk));
	jand g1396(.dina(w_n978_1[0]),.dinb(w_n295_48[1]),.dout(n1659),.clk(gclk));
	jand g1397(.dina(w_n988_1[0]),.dinb(w_n308_48[1]),.dout(n1660),.clk(gclk));
	jor g1398(.dina(n1660),.dinb(n1659),.dout(n1661),.clk(gclk));
	jor g1399(.dina(n1661),.dinb(n1658),.dout(n1662),.clk(gclk));
	jand g1400(.dina(w_n1662_1[1]),.dinb(w_n323_59[2]),.dout(n1663),.clk(gclk));
	jor g1401(.dina(n1663),.dinb(n1655),.dout(n1664),.clk(gclk));
	jand g1402(.dina(w_n740_1[0]),.dinb(w_n266_48[0]),.dout(n1665),.clk(gclk));
	jand g1403(.dina(w_n910_1[0]),.dinb(w_n281_48[0]),.dout(n1666),.clk(gclk));
	jor g1404(.dina(n1666),.dinb(n1665),.dout(n1667),.clk(gclk));
	jand g1405(.dina(w_n889_1[0]),.dinb(w_n295_48[0]),.dout(n1668),.clk(gclk));
	jand g1406(.dina(w_n899_1[0]),.dinb(w_n308_48[0]),.dout(n1669),.clk(gclk));
	jor g1407(.dina(n1669),.dinb(n1668),.dout(n1670),.clk(gclk));
	jor g1408(.dina(n1670),.dinb(n1667),.dout(n1671),.clk(gclk));
	jand g1409(.dina(w_n1671_1[1]),.dinb(w_n485_59[2]),.dout(n1672),.clk(gclk));
	jand g1410(.dina(w_n1057_1[0]),.dinb(w_n266_47[2]),.dout(n1673),.clk(gclk));
	jand g1411(.dina(w_n954_1[0]),.dinb(w_n281_47[2]),.dout(n1674),.clk(gclk));
	jor g1412(.dina(n1674),.dinb(n1673),.dout(n1675),.clk(gclk));
	jand g1413(.dina(w_n933_1[0]),.dinb(w_n295_47[2]),.dout(n1676),.clk(gclk));
	jand g1414(.dina(w_n943_1[0]),.dinb(w_n308_47[2]),.dout(n1677),.clk(gclk));
	jor g1415(.dina(n1677),.dinb(n1676),.dout(n1678),.clk(gclk));
	jor g1416(.dina(n1678),.dinb(n1675),.dout(n1679),.clk(gclk));
	jand g1417(.dina(w_n1679_1[1]),.dinb(w_n432_59[2]),.dout(n1680),.clk(gclk));
	jor g1418(.dina(n1680),.dinb(n1672),.dout(n1681),.clk(gclk));
	jor g1419(.dina(n1681),.dinb(n1664),.dout(n1682),.clk(gclk));
	jand g1420(.dina(w_n1682_0[1]),.dinb(w_shift6_61[2]),.dout(n1683),.clk(gclk));
	jor g1421(.dina(n1683),.dinb(n1647),.dout(result5),.clk(gclk));
	jand g1422(.dina(w_n1170_1[0]),.dinb(w_n266_47[1]),.dout(n1685),.clk(gclk));
	jand g1423(.dina(w_n1089_1[0]),.dinb(w_n281_47[1]),.dout(n1686),.clk(gclk));
	jor g1424(.dina(n1686),.dinb(n1685),.dout(n1687),.clk(gclk));
	jand g1425(.dina(w_n1072_1[0]),.dinb(w_n295_47[1]),.dout(n1688),.clk(gclk));
	jand g1426(.dina(w_n1080_1[0]),.dinb(w_n308_47[1]),.dout(n1689),.clk(gclk));
	jor g1427(.dina(n1689),.dinb(n1688),.dout(n1690),.clk(gclk));
	jor g1428(.dina(n1690),.dinb(n1687),.dout(n1691),.clk(gclk));
	jand g1429(.dina(w_n1691_1[1]),.dinb(w_n323_59[1]),.dout(n1692),.clk(gclk));
	jand g1430(.dina(w_n1206_1[0]),.dinb(w_n266_47[0]),.dout(n1693),.clk(gclk));
	jand g1431(.dina(w_n1125_1[0]),.dinb(w_n281_47[0]),.dout(n1694),.clk(gclk));
	jor g1432(.dina(n1694),.dinb(n1693),.dout(n1695),.clk(gclk));
	jand g1433(.dina(w_n1108_1[0]),.dinb(w_n295_47[0]),.dout(n1696),.clk(gclk));
	jand g1434(.dina(w_n1116_1[0]),.dinb(w_n308_47[0]),.dout(n1697),.clk(gclk));
	jor g1435(.dina(n1697),.dinb(n1696),.dout(n1698),.clk(gclk));
	jor g1436(.dina(n1698),.dinb(n1695),.dout(n1699),.clk(gclk));
	jand g1437(.dina(w_n1699_1[1]),.dinb(w_n377_59[1]),.dout(n1700),.clk(gclk));
	jor g1438(.dina(n1700),.dinb(n1692),.dout(n1701),.clk(gclk));
	jand g1439(.dina(w_n1133_1[0]),.dinb(w_n266_46[2]),.dout(n1702),.clk(gclk));
	jand g1440(.dina(w_n1162_1[0]),.dinb(w_n281_46[2]),.dout(n1703),.clk(gclk));
	jor g1441(.dina(n1703),.dinb(n1702),.dout(n1704),.clk(gclk));
	jand g1442(.dina(w_n1145_1[0]),.dinb(w_n295_46[2]),.dout(n1705),.clk(gclk));
	jand g1443(.dina(w_n1153_1[0]),.dinb(w_n308_46[2]),.dout(n1706),.clk(gclk));
	jor g1444(.dina(n1706),.dinb(n1705),.dout(n1707),.clk(gclk));
	jor g1445(.dina(n1707),.dinb(n1704),.dout(n1708),.clk(gclk));
	jand g1446(.dina(w_n1708_1[1]),.dinb(w_n432_59[1]),.dout(n1709),.clk(gclk));
	jand g1447(.dina(w_n1318_1[0]),.dinb(w_n266_46[1]),.dout(n1710),.clk(gclk));
	jand g1448(.dina(w_n1198_1[0]),.dinb(w_n281_46[1]),.dout(n1711),.clk(gclk));
	jor g1449(.dina(n1711),.dinb(n1710),.dout(n1712),.clk(gclk));
	jand g1450(.dina(w_n1181_1[0]),.dinb(w_n295_46[1]),.dout(n1713),.clk(gclk));
	jand g1451(.dina(w_n1189_1[0]),.dinb(w_n308_46[1]),.dout(n1714),.clk(gclk));
	jor g1452(.dina(n1714),.dinb(n1713),.dout(n1715),.clk(gclk));
	jor g1453(.dina(n1715),.dinb(n1712),.dout(n1716),.clk(gclk));
	jand g1454(.dina(w_n1716_1[1]),.dinb(w_n485_59[1]),.dout(n1717),.clk(gclk));
	jor g1455(.dina(n1717),.dinb(n1709),.dout(n1718),.clk(gclk));
	jor g1456(.dina(n1718),.dinb(n1701),.dout(n1719),.clk(gclk));
	jand g1457(.dina(w_n1719_0[1]),.dinb(w_n263_61[1]),.dout(n1720),.clk(gclk));
	jand g1458(.dina(w_n1245_1[0]),.dinb(w_n266_46[0]),.dout(n1721),.clk(gclk));
	jand g1459(.dina(w_n1346_1[0]),.dinb(w_n281_46[0]),.dout(n1722),.clk(gclk));
	jor g1460(.dina(n1722),.dinb(n1721),.dout(n1723),.clk(gclk));
	jand g1461(.dina(w_n1329_1[0]),.dinb(w_n295_46[0]),.dout(n1724),.clk(gclk));
	jand g1462(.dina(w_n1337_1[0]),.dinb(w_n308_46[0]),.dout(n1725),.clk(gclk));
	jor g1463(.dina(n1725),.dinb(n1724),.dout(n1726),.clk(gclk));
	jor g1464(.dina(n1726),.dinb(n1723),.dout(n1727),.clk(gclk));
	jand g1465(.dina(w_n1727_1[1]),.dinb(w_n377_59[0]),.dout(n1728),.clk(gclk));
	jand g1466(.dina(w_n1281_1[0]),.dinb(w_n266_45[2]),.dout(n1729),.clk(gclk));
	jand g1467(.dina(w_n1310_1[0]),.dinb(w_n281_45[2]),.dout(n1730),.clk(gclk));
	jor g1468(.dina(n1730),.dinb(n1729),.dout(n1731),.clk(gclk));
	jand g1469(.dina(w_n1293_1[0]),.dinb(w_n295_45[2]),.dout(n1732),.clk(gclk));
	jand g1470(.dina(w_n1301_1[0]),.dinb(w_n308_45[2]),.dout(n1733),.clk(gclk));
	jor g1471(.dina(n1733),.dinb(n1732),.dout(n1734),.clk(gclk));
	jor g1472(.dina(n1734),.dinb(n1731),.dout(n1735),.clk(gclk));
	jand g1473(.dina(w_n1735_1[1]),.dinb(w_n323_59[0]),.dout(n1736),.clk(gclk));
	jor g1474(.dina(n1736),.dinb(n1728),.dout(n1737),.clk(gclk));
	jand g1475(.dina(w_n1097_1[0]),.dinb(w_n266_45[1]),.dout(n1738),.clk(gclk));
	jand g1476(.dina(w_n1237_1[0]),.dinb(w_n281_45[1]),.dout(n1739),.clk(gclk));
	jor g1477(.dina(n1739),.dinb(n1738),.dout(n1740),.clk(gclk));
	jand g1478(.dina(w_n1220_1[0]),.dinb(w_n295_45[1]),.dout(n1741),.clk(gclk));
	jand g1479(.dina(w_n1228_1[0]),.dinb(w_n308_45[1]),.dout(n1742),.clk(gclk));
	jor g1480(.dina(n1742),.dinb(n1741),.dout(n1743),.clk(gclk));
	jor g1481(.dina(n1743),.dinb(n1740),.dout(n1744),.clk(gclk));
	jand g1482(.dina(w_n1744_1[1]),.dinb(w_n485_59[0]),.dout(n1745),.clk(gclk));
	jand g1483(.dina(w_n1354_1[0]),.dinb(w_n266_45[0]),.dout(n1746),.clk(gclk));
	jand g1484(.dina(w_n1273_1[0]),.dinb(w_n281_45[0]),.dout(n1747),.clk(gclk));
	jor g1485(.dina(n1747),.dinb(n1746),.dout(n1748),.clk(gclk));
	jand g1486(.dina(w_n1256_1[0]),.dinb(w_n295_45[0]),.dout(n1749),.clk(gclk));
	jand g1487(.dina(w_n1264_1[0]),.dinb(w_n308_45[0]),.dout(n1750),.clk(gclk));
	jor g1488(.dina(n1750),.dinb(n1749),.dout(n1751),.clk(gclk));
	jor g1489(.dina(n1751),.dinb(n1748),.dout(n1752),.clk(gclk));
	jand g1490(.dina(w_n1752_1[1]),.dinb(w_n432_59[0]),.dout(n1753),.clk(gclk));
	jor g1491(.dina(n1753),.dinb(n1745),.dout(n1754),.clk(gclk));
	jor g1492(.dina(n1754),.dinb(n1737),.dout(n1755),.clk(gclk));
	jand g1493(.dina(w_n1755_0[1]),.dinb(w_shift6_61[1]),.dout(n1756),.clk(gclk));
	jor g1494(.dina(n1756),.dinb(n1720),.dout(result6),.clk(gclk));
	jand g1495(.dina(w_n1419_1[0]),.dinb(w_n266_44[2]),.dout(n1758),.clk(gclk));
	jand g1496(.dina(w_n1394_1[0]),.dinb(w_n281_44[2]),.dout(n1759),.clk(gclk));
	jor g1497(.dina(n1759),.dinb(n1758),.dout(n1760),.clk(gclk));
	jand g1498(.dina(w_n1385_1[0]),.dinb(w_n295_44[2]),.dout(n1761),.clk(gclk));
	jand g1499(.dina(w_n1389_1[0]),.dinb(w_n308_44[2]),.dout(n1762),.clk(gclk));
	jor g1500(.dina(n1762),.dinb(n1761),.dout(n1763),.clk(gclk));
	jor g1501(.dina(n1763),.dinb(n1760),.dout(n1764),.clk(gclk));
	jand g1502(.dina(w_n1764_1[1]),.dinb(w_n323_58[2]),.dout(n1765),.clk(gclk));
	jand g1503(.dina(w_n1439_1[0]),.dinb(w_n266_44[1]),.dout(n1766),.clk(gclk));
	jand g1504(.dina(w_n1374_1[0]),.dinb(w_n281_44[1]),.dout(n1767),.clk(gclk));
	jor g1505(.dina(n1767),.dinb(n1766),.dout(n1768),.clk(gclk));
	jand g1506(.dina(w_n1365_1[0]),.dinb(w_n295_44[1]),.dout(n1769),.clk(gclk));
	jand g1507(.dina(w_n1369_1[0]),.dinb(w_n308_44[1]),.dout(n1770),.clk(gclk));
	jor g1508(.dina(n1770),.dinb(n1769),.dout(n1771),.clk(gclk));
	jor g1509(.dina(n1771),.dinb(n1768),.dout(n1772),.clk(gclk));
	jand g1510(.dina(w_n1772_1[1]),.dinb(w_n377_58[2]),.dout(n1773),.clk(gclk));
	jor g1511(.dina(n1773),.dinb(n1765),.dout(n1774),.clk(gclk));
	jand g1512(.dina(w_n1378_1[0]),.dinb(w_n266_44[0]),.dout(n1775),.clk(gclk));
	jand g1513(.dina(w_n1415_1[0]),.dinb(w_n281_44[0]),.dout(n1776),.clk(gclk));
	jor g1514(.dina(n1776),.dinb(n1775),.dout(n1777),.clk(gclk));
	jand g1515(.dina(w_n1406_1[0]),.dinb(w_n295_44[0]),.dout(n1778),.clk(gclk));
	jand g1516(.dina(w_n1410_1[0]),.dinb(w_n308_44[0]),.dout(n1779),.clk(gclk));
	jor g1517(.dina(n1779),.dinb(n1778),.dout(n1780),.clk(gclk));
	jor g1518(.dina(n1780),.dinb(n1777),.dout(n1781),.clk(gclk));
	jand g1519(.dina(w_n1781_1[1]),.dinb(w_n432_58[2]),.dout(n1782),.clk(gclk));
	jand g1520(.dina(w_n1530_1[0]),.dinb(w_n266_43[2]),.dout(n1783),.clk(gclk));
	jand g1521(.dina(w_n1435_1[0]),.dinb(w_n281_43[2]),.dout(n1784),.clk(gclk));
	jor g1522(.dina(n1784),.dinb(n1783),.dout(n1785),.clk(gclk));
	jand g1523(.dina(w_n1426_1[0]),.dinb(w_n295_43[2]),.dout(n1786),.clk(gclk));
	jand g1524(.dina(w_n1430_1[0]),.dinb(w_n308_43[2]),.dout(n1787),.clk(gclk));
	jor g1525(.dina(n1787),.dinb(n1786),.dout(n1788),.clk(gclk));
	jor g1526(.dina(n1788),.dinb(n1785),.dout(n1789),.clk(gclk));
	jand g1527(.dina(w_n1789_1[1]),.dinb(w_n485_58[2]),.dout(n1790),.clk(gclk));
	jor g1528(.dina(n1790),.dinb(n1782),.dout(n1791),.clk(gclk));
	jor g1529(.dina(n1791),.dinb(n1774),.dout(n1792),.clk(gclk));
	jand g1530(.dina(w_n1792_0[1]),.dinb(w_n263_61[0]),.dout(n1793),.clk(gclk));
	jand g1531(.dina(w_n1490_1[0]),.dinb(w_n295_43[1]),.dout(n1794),.clk(gclk));
	jand g1532(.dina(w_n1462_1[0]),.dinb(w_n266_43[1]),.dout(n1795),.clk(gclk));
	jor g1533(.dina(n1795),.dinb(n1794),.dout(n1796),.clk(gclk));
	jand g1534(.dina(w_n1505_1[0]),.dinb(w_n281_43[1]),.dout(n1797),.clk(gclk));
	jand g1535(.dina(w_n1496_1[0]),.dinb(w_n308_43[1]),.dout(n1798),.clk(gclk));
	jor g1536(.dina(n1798),.dinb(n1797),.dout(n1799),.clk(gclk));
	jor g1537(.dina(n1799),.dinb(n1796),.dout(n1800),.clk(gclk));
	jand g1538(.dina(w_n1800_1[1]),.dinb(w_n377_58[1]),.dout(n1801),.clk(gclk));
	jand g1539(.dina(w_n1482_1[0]),.dinb(w_n266_43[0]),.dout(n1802),.clk(gclk));
	jand g1540(.dina(w_n1526_1[0]),.dinb(w_n281_43[0]),.dout(n1803),.clk(gclk));
	jor g1541(.dina(n1803),.dinb(n1802),.dout(n1804),.clk(gclk));
	jand g1542(.dina(w_n1517_1[0]),.dinb(w_n295_43[0]),.dout(n1805),.clk(gclk));
	jand g1543(.dina(w_n1521_1[0]),.dinb(w_n308_43[0]),.dout(n1806),.clk(gclk));
	jor g1544(.dina(n1806),.dinb(n1805),.dout(n1807),.clk(gclk));
	jor g1545(.dina(n1807),.dinb(n1804),.dout(n1808),.clk(gclk));
	jand g1546(.dina(w_n1808_1[1]),.dinb(w_n323_58[1]),.dout(n1809),.clk(gclk));
	jor g1547(.dina(n1809),.dinb(n1801),.dout(n1810),.clk(gclk));
	jand g1548(.dina(w_n1398_1[0]),.dinb(w_n266_42[2]),.dout(n1811),.clk(gclk));
	jand g1549(.dina(w_n1458_1[0]),.dinb(w_n281_42[2]),.dout(n1812),.clk(gclk));
	jor g1550(.dina(n1812),.dinb(n1811),.dout(n1813),.clk(gclk));
	jand g1551(.dina(w_n1449_1[0]),.dinb(w_n295_42[2]),.dout(n1814),.clk(gclk));
	jand g1552(.dina(w_n1453_1[0]),.dinb(w_n308_42[2]),.dout(n1815),.clk(gclk));
	jor g1553(.dina(n1815),.dinb(n1814),.dout(n1816),.clk(gclk));
	jor g1554(.dina(n1816),.dinb(n1813),.dout(n1817),.clk(gclk));
	jand g1555(.dina(w_n1817_1[1]),.dinb(w_n485_58[1]),.dout(n1818),.clk(gclk));
	jand g1556(.dina(w_n1510_1[0]),.dinb(w_n266_42[1]),.dout(n1819),.clk(gclk));
	jand g1557(.dina(w_n1478_1[0]),.dinb(w_n281_42[1]),.dout(n1820),.clk(gclk));
	jor g1558(.dina(n1820),.dinb(n1819),.dout(n1821),.clk(gclk));
	jand g1559(.dina(w_n1469_1[0]),.dinb(w_n295_42[1]),.dout(n1822),.clk(gclk));
	jand g1560(.dina(w_n1473_1[0]),.dinb(w_n308_42[1]),.dout(n1823),.clk(gclk));
	jor g1561(.dina(n1823),.dinb(n1822),.dout(n1824),.clk(gclk));
	jor g1562(.dina(n1824),.dinb(n1821),.dout(n1825),.clk(gclk));
	jand g1563(.dina(w_n1825_1[1]),.dinb(w_n432_58[1]),.dout(n1826),.clk(gclk));
	jor g1564(.dina(n1826),.dinb(n1818),.dout(n1827),.clk(gclk));
	jor g1565(.dina(n1827),.dinb(n1810),.dout(n1828),.clk(gclk));
	jand g1566(.dina(w_n1828_0[1]),.dinb(w_shift6_61[0]),.dout(n1829),.clk(gclk));
	jor g1567(.dina(n1829),.dinb(n1793),.dout(result7),.clk(gclk));
	jand g1568(.dina(w_n402_0[2]),.dinb(w_n266_42[0]),.dout(n1831),.clk(gclk));
	jand g1569(.dina(w_n281_42[0]),.dinb(w_n279_0[2]),.dout(n1832),.clk(gclk));
	jor g1570(.dina(n1832),.dinb(n1831),.dout(n1833),.clk(gclk));
	jand g1571(.dina(w_n427_0[2]),.dinb(w_n295_42[0]),.dout(n1834),.clk(gclk));
	jand g1572(.dina(w_n308_42[0]),.dinb(w_n306_0[2]),.dout(n1835),.clk(gclk));
	jor g1573(.dina(n1835),.dinb(n1834),.dout(n1836),.clk(gclk));
	jor g1574(.dina(n1836),.dinb(n1833),.dout(n1837),.clk(gclk));
	jand g1575(.dina(w_n1837_1[1]),.dinb(w_n323_58[0]),.dout(n1838),.clk(gclk));
	jand g1576(.dina(w_n456_0[2]),.dinb(w_n266_41[2]),.dout(n1839),.clk(gclk));
	jand g1577(.dina(w_n335_0[2]),.dinb(w_n281_41[2]),.dout(n1840),.clk(gclk));
	jor g1578(.dina(n1840),.dinb(n1839),.dout(n1841),.clk(gclk));
	jand g1579(.dina(w_n481_0[2]),.dinb(w_n295_41[2]),.dout(n1842),.clk(gclk));
	jand g1580(.dina(w_n360_0[2]),.dinb(w_n308_41[2]),.dout(n1843),.clk(gclk));
	jor g1581(.dina(n1843),.dinb(n1842),.dout(n1844),.clk(gclk));
	jor g1582(.dina(n1844),.dinb(n1841),.dout(n1845),.clk(gclk));
	jand g1583(.dina(w_n1845_1[1]),.dinb(w_n377_58[0]),.dout(n1846),.clk(gclk));
	jor g1584(.dina(n1846),.dinb(n1838),.dout(n1847),.clk(gclk));
	jand g1585(.dina(w_n347_0[2]),.dinb(w_n266_41[1]),.dout(n1848),.clk(gclk));
	jand g1586(.dina(w_n390_0[2]),.dinb(w_n281_41[1]),.dout(n1849),.clk(gclk));
	jor g1587(.dina(n1849),.dinb(n1848),.dout(n1850),.clk(gclk));
	jand g1588(.dina(w_n372_0[2]),.dinb(w_n295_41[1]),.dout(n1851),.clk(gclk));
	jand g1589(.dina(w_n415_0[2]),.dinb(w_n308_41[1]),.dout(n1852),.clk(gclk));
	jor g1590(.dina(n1852),.dinb(n1851),.dout(n1853),.clk(gclk));
	jor g1591(.dina(n1853),.dinb(n1850),.dout(n1854),.clk(gclk));
	jand g1592(.dina(w_n1854_1[1]),.dinb(w_n432_58[0]),.dout(n1855),.clk(gclk));
	jand g1593(.dina(w_n512_0[2]),.dinb(w_n266_41[0]),.dout(n1856),.clk(gclk));
	jand g1594(.dina(w_n444_0[2]),.dinb(w_n281_41[0]),.dout(n1857),.clk(gclk));
	jor g1595(.dina(n1857),.dinb(n1856),.dout(n1858),.clk(gclk));
	jand g1596(.dina(w_n537_0[2]),.dinb(w_n295_41[0]),.dout(n1859),.clk(gclk));
	jand g1597(.dina(w_n469_0[2]),.dinb(w_n308_41[0]),.dout(n1860),.clk(gclk));
	jor g1598(.dina(n1860),.dinb(n1859),.dout(n1861),.clk(gclk));
	jor g1599(.dina(n1861),.dinb(n1858),.dout(n1862),.clk(gclk));
	jand g1600(.dina(w_n1862_1[1]),.dinb(w_n485_58[0]),.dout(n1863),.clk(gclk));
	jor g1601(.dina(n1863),.dinb(n1855),.dout(n1864),.clk(gclk));
	jor g1602(.dina(n1864),.dinb(n1847),.dout(n1865),.clk(gclk));
	jand g1603(.dina(w_n1865_0[1]),.dinb(w_n263_60[2]),.dout(n1866),.clk(gclk));
	jand g1604(.dina(w_n667_0[2]),.dinb(w_n266_40[2]),.dout(n1867),.clk(gclk));
	jand g1605(.dina(w_n552_0[2]),.dinb(w_n281_40[2]),.dout(n1868),.clk(gclk));
	jor g1606(.dina(n1868),.dinb(n1867),.dout(n1869),.clk(gclk));
	jand g1607(.dina(w_n692_0[2]),.dinb(w_n295_40[2]),.dout(n1870),.clk(gclk));
	jand g1608(.dina(w_n575_0[2]),.dinb(w_n308_40[2]),.dout(n1871),.clk(gclk));
	jor g1609(.dina(n1871),.dinb(n1870),.dout(n1872),.clk(gclk));
	jor g1610(.dina(n1872),.dinb(n1869),.dout(n1873),.clk(gclk));
	jand g1611(.dina(w_n1873_1[1]),.dinb(w_n377_57[2]),.dout(n1874),.clk(gclk));
	jand g1612(.dina(w_n615_0[2]),.dinb(w_n266_40[1]),.dout(n1875),.clk(gclk));
	jand g1613(.dina(w_n500_0[2]),.dinb(w_n281_40[1]),.dout(n1876),.clk(gclk));
	jor g1614(.dina(n1876),.dinb(n1875),.dout(n1877),.clk(gclk));
	jand g1615(.dina(w_n640_0[2]),.dinb(w_n295_40[1]),.dout(n1878),.clk(gclk));
	jand g1616(.dina(w_n525_0[2]),.dinb(w_n308_40[1]),.dout(n1879),.clk(gclk));
	jor g1617(.dina(n1879),.dinb(n1878),.dout(n1880),.clk(gclk));
	jor g1618(.dina(n1880),.dinb(n1877),.dout(n1881),.clk(gclk));
	jand g1619(.dina(w_n1881_1[1]),.dinb(w_n323_57[2]),.dout(n1882),.clk(gclk));
	jor g1620(.dina(n1882),.dinb(n1874),.dout(n1883),.clk(gclk));
	jand g1621(.dina(w_n292_0[2]),.dinb(w_n266_40[0]),.dout(n1884),.clk(gclk));
	jand g1622(.dina(w_n655_0[2]),.dinb(w_n281_40[0]),.dout(n1885),.clk(gclk));
	jor g1623(.dina(n1885),.dinb(n1884),.dout(n1886),.clk(gclk));
	jand g1624(.dina(w_n319_0[2]),.dinb(w_n295_40[0]),.dout(n1887),.clk(gclk));
	jand g1625(.dina(w_n680_0[2]),.dinb(w_n308_40[0]),.dout(n1888),.clk(gclk));
	jor g1626(.dina(n1888),.dinb(n1887),.dout(n1889),.clk(gclk));
	jor g1627(.dina(n1889),.dinb(n1886),.dout(n1890),.clk(gclk));
	jand g1628(.dina(w_n1890_1[1]),.dinb(w_n485_57[2]),.dout(n1891),.clk(gclk));
	jand g1629(.dina(w_n562_0[2]),.dinb(w_n266_39[2]),.dout(n1892),.clk(gclk));
	jand g1630(.dina(w_n603_0[2]),.dinb(w_n281_39[2]),.dout(n1893),.clk(gclk));
	jor g1631(.dina(n1893),.dinb(n1892),.dout(n1894),.clk(gclk));
	jand g1632(.dina(w_n587_0[2]),.dinb(w_n295_39[2]),.dout(n1895),.clk(gclk));
	jand g1633(.dina(w_n628_0[2]),.dinb(w_n308_39[2]),.dout(n1896),.clk(gclk));
	jor g1634(.dina(n1896),.dinb(n1895),.dout(n1897),.clk(gclk));
	jor g1635(.dina(n1897),.dinb(n1894),.dout(n1898),.clk(gclk));
	jand g1636(.dina(w_n1898_1[1]),.dinb(w_n432_57[2]),.dout(n1899),.clk(gclk));
	jor g1637(.dina(n1899),.dinb(n1891),.dout(n1900),.clk(gclk));
	jor g1638(.dina(n1900),.dinb(n1883),.dout(n1901),.clk(gclk));
	jand g1639(.dina(w_n1901_0[1]),.dinb(w_shift6_60[2]),.dout(n1902),.clk(gclk));
	jor g1640(.dina(n1902),.dinb(n1866),.dout(result8),.clk(gclk));
	jand g1641(.dina(w_n808_0[2]),.dinb(w_n266_39[1]),.dout(n1904),.clk(gclk));
	jand g1642(.dina(w_n709_0[2]),.dinb(w_n281_39[1]),.dout(n1905),.clk(gclk));
	jor g1643(.dina(n1905),.dinb(n1904),.dout(n1906),.clk(gclk));
	jand g1644(.dina(w_n829_0[2]),.dinb(w_n295_39[1]),.dout(n1907),.clk(gclk));
	jand g1645(.dina(w_n730_0[2]),.dinb(w_n308_39[1]),.dout(n1908),.clk(gclk));
	jor g1646(.dina(n1908),.dinb(n1907),.dout(n1909),.clk(gclk));
	jor g1647(.dina(n1909),.dinb(n1906),.dout(n1910),.clk(gclk));
	jand g1648(.dina(w_n1910_1[1]),.dinb(w_n323_57[1]),.dout(n1911),.clk(gclk));
	jand g1649(.dina(w_n852_0[2]),.dinb(w_n266_39[0]),.dout(n1912),.clk(gclk));
	jand g1650(.dina(w_n753_0[2]),.dinb(w_n281_39[0]),.dout(n1913),.clk(gclk));
	jor g1651(.dina(n1913),.dinb(n1912),.dout(n1914),.clk(gclk));
	jand g1652(.dina(w_n873_0[2]),.dinb(w_n295_39[0]),.dout(n1915),.clk(gclk));
	jand g1653(.dina(w_n774_0[2]),.dinb(w_n308_39[0]),.dout(n1916),.clk(gclk));
	jor g1654(.dina(n1916),.dinb(n1915),.dout(n1917),.clk(gclk));
	jor g1655(.dina(n1917),.dinb(n1914),.dout(n1918),.clk(gclk));
	jand g1656(.dina(w_n1918_1[1]),.dinb(w_n377_57[1]),.dout(n1919),.clk(gclk));
	jor g1657(.dina(n1919),.dinb(n1911),.dout(n1920),.clk(gclk));
	jand g1658(.dina(w_n763_0[2]),.dinb(w_n266_38[2]),.dout(n1921),.clk(gclk));
	jand g1659(.dina(w_n798_0[2]),.dinb(w_n281_38[2]),.dout(n1922),.clk(gclk));
	jor g1660(.dina(n1922),.dinb(n1921),.dout(n1923),.clk(gclk));
	jand g1661(.dina(w_n784_0[2]),.dinb(w_n295_38[2]),.dout(n1924),.clk(gclk));
	jand g1662(.dina(w_n819_0[2]),.dinb(w_n308_38[2]),.dout(n1925),.clk(gclk));
	jor g1663(.dina(n1925),.dinb(n1924),.dout(n1926),.clk(gclk));
	jor g1664(.dina(n1926),.dinb(n1923),.dout(n1927),.clk(gclk));
	jand g1665(.dina(w_n1927_1[1]),.dinb(w_n432_57[1]),.dout(n1928),.clk(gclk));
	jand g1666(.dina(w_n988_0[2]),.dinb(w_n266_38[1]),.dout(n1929),.clk(gclk));
	jand g1667(.dina(w_n842_0[2]),.dinb(w_n281_38[1]),.dout(n1930),.clk(gclk));
	jor g1668(.dina(n1930),.dinb(n1929),.dout(n1931),.clk(gclk));
	jand g1669(.dina(w_n1009_0[2]),.dinb(w_n295_38[1]),.dout(n1932),.clk(gclk));
	jand g1670(.dina(w_n863_0[2]),.dinb(w_n308_38[1]),.dout(n1933),.clk(gclk));
	jor g1671(.dina(n1933),.dinb(n1932),.dout(n1934),.clk(gclk));
	jor g1672(.dina(n1934),.dinb(n1931),.dout(n1935),.clk(gclk));
	jand g1673(.dina(w_n1935_1[1]),.dinb(w_n485_57[1]),.dout(n1936),.clk(gclk));
	jor g1674(.dina(n1936),.dinb(n1928),.dout(n1937),.clk(gclk));
	jor g1675(.dina(n1937),.dinb(n1920),.dout(n1938),.clk(gclk));
	jand g1676(.dina(w_n1938_0[1]),.dinb(w_n263_60[1]),.dout(n1939),.clk(gclk));
	jand g1677(.dina(w_n899_0[2]),.dinb(w_n266_38[0]),.dout(n1940),.clk(gclk));
	jand g1678(.dina(w_n1022_0[2]),.dinb(w_n281_38[0]),.dout(n1941),.clk(gclk));
	jor g1679(.dina(n1941),.dinb(n1940),.dout(n1942),.clk(gclk));
	jand g1680(.dina(w_n920_0[2]),.dinb(w_n295_38[0]),.dout(n1943),.clk(gclk));
	jand g1681(.dina(w_n1047_0[2]),.dinb(w_n308_38[0]),.dout(n1944),.clk(gclk));
	jor g1682(.dina(n1944),.dinb(n1943),.dout(n1945),.clk(gclk));
	jor g1683(.dina(n1945),.dinb(n1942),.dout(n1946),.clk(gclk));
	jand g1684(.dina(w_n1946_1[1]),.dinb(w_n377_57[0]),.dout(n1947),.clk(gclk));
	jand g1685(.dina(w_n943_0[2]),.dinb(w_n266_37[2]),.dout(n1948),.clk(gclk));
	jand g1686(.dina(w_n978_0[2]),.dinb(w_n281_37[2]),.dout(n1949),.clk(gclk));
	jor g1687(.dina(n1949),.dinb(n1948),.dout(n1950),.clk(gclk));
	jand g1688(.dina(w_n964_0[2]),.dinb(w_n295_37[2]),.dout(n1951),.clk(gclk));
	jand g1689(.dina(w_n999_0[2]),.dinb(w_n308_37[2]),.dout(n1952),.clk(gclk));
	jor g1690(.dina(n1952),.dinb(n1951),.dout(n1953),.clk(gclk));
	jor g1691(.dina(n1953),.dinb(n1950),.dout(n1954),.clk(gclk));
	jand g1692(.dina(w_n1954_1[1]),.dinb(w_n323_57[0]),.dout(n1955),.clk(gclk));
	jor g1693(.dina(n1955),.dinb(n1947),.dout(n1956),.clk(gclk));
	jand g1694(.dina(w_n719_0[2]),.dinb(w_n266_37[1]),.dout(n1957),.clk(gclk));
	jand g1695(.dina(w_n889_0[2]),.dinb(w_n281_37[1]),.dout(n1958),.clk(gclk));
	jor g1696(.dina(n1958),.dinb(n1957),.dout(n1959),.clk(gclk));
	jand g1697(.dina(w_n740_0[2]),.dinb(w_n295_37[1]),.dout(n1960),.clk(gclk));
	jand g1698(.dina(w_n910_0[2]),.dinb(w_n308_37[1]),.dout(n1961),.clk(gclk));
	jor g1699(.dina(n1961),.dinb(n1960),.dout(n1962),.clk(gclk));
	jor g1700(.dina(n1962),.dinb(n1959),.dout(n1963),.clk(gclk));
	jand g1701(.dina(w_n1963_1[1]),.dinb(w_n485_57[0]),.dout(n1964),.clk(gclk));
	jand g1702(.dina(w_n1034_0[2]),.dinb(w_n266_37[0]),.dout(n1965),.clk(gclk));
	jand g1703(.dina(w_n933_0[2]),.dinb(w_n281_37[0]),.dout(n1966),.clk(gclk));
	jor g1704(.dina(n1966),.dinb(n1965),.dout(n1967),.clk(gclk));
	jand g1705(.dina(w_n1057_0[2]),.dinb(w_n295_37[0]),.dout(n1968),.clk(gclk));
	jand g1706(.dina(w_n954_0[2]),.dinb(w_n308_37[0]),.dout(n1969),.clk(gclk));
	jor g1707(.dina(n1969),.dinb(n1968),.dout(n1970),.clk(gclk));
	jor g1708(.dina(n1970),.dinb(n1967),.dout(n1971),.clk(gclk));
	jand g1709(.dina(w_n1971_1[1]),.dinb(w_n432_57[0]),.dout(n1972),.clk(gclk));
	jor g1710(.dina(n1972),.dinb(n1964),.dout(n1973),.clk(gclk));
	jor g1711(.dina(n1973),.dinb(n1956),.dout(n1974),.clk(gclk));
	jand g1712(.dina(w_n1974_0[1]),.dinb(w_shift6_60[1]),.dout(n1975),.clk(gclk));
	jor g1713(.dina(n1975),.dinb(n1939),.dout(result9),.clk(gclk));
	jand g1714(.dina(w_n1153_0[2]),.dinb(w_n266_36[2]),.dout(n1977),.clk(gclk));
	jand g1715(.dina(w_n1072_0[2]),.dinb(w_n281_36[2]),.dout(n1978),.clk(gclk));
	jor g1716(.dina(n1978),.dinb(n1977),.dout(n1979),.clk(gclk));
	jand g1717(.dina(w_n1170_0[2]),.dinb(w_n295_36[2]),.dout(n1980),.clk(gclk));
	jand g1718(.dina(w_n1089_0[2]),.dinb(w_n308_36[2]),.dout(n1981),.clk(gclk));
	jor g1719(.dina(n1981),.dinb(n1980),.dout(n1982),.clk(gclk));
	jor g1720(.dina(n1982),.dinb(n1979),.dout(n1983),.clk(gclk));
	jand g1721(.dina(w_n1983_1[1]),.dinb(w_n323_56[2]),.dout(n1984),.clk(gclk));
	jand g1722(.dina(w_n1189_0[2]),.dinb(w_n266_36[1]),.dout(n1985),.clk(gclk));
	jand g1723(.dina(w_n1108_0[2]),.dinb(w_n281_36[1]),.dout(n1986),.clk(gclk));
	jor g1724(.dina(n1986),.dinb(n1985),.dout(n1987),.clk(gclk));
	jand g1725(.dina(w_n1206_0[2]),.dinb(w_n295_36[1]),.dout(n1988),.clk(gclk));
	jand g1726(.dina(w_n1125_0[2]),.dinb(w_n308_36[1]),.dout(n1989),.clk(gclk));
	jor g1727(.dina(n1989),.dinb(n1988),.dout(n1990),.clk(gclk));
	jor g1728(.dina(n1990),.dinb(n1987),.dout(n1991),.clk(gclk));
	jand g1729(.dina(w_n1991_1[1]),.dinb(w_n377_56[2]),.dout(n1992),.clk(gclk));
	jor g1730(.dina(n1992),.dinb(n1984),.dout(n1993),.clk(gclk));
	jand g1731(.dina(w_n1116_0[2]),.dinb(w_n266_36[0]),.dout(n1994),.clk(gclk));
	jand g1732(.dina(w_n1145_0[2]),.dinb(w_n281_36[0]),.dout(n1995),.clk(gclk));
	jor g1733(.dina(n1995),.dinb(n1994),.dout(n1996),.clk(gclk));
	jand g1734(.dina(w_n1133_0[2]),.dinb(w_n295_36[0]),.dout(n1997),.clk(gclk));
	jand g1735(.dina(w_n1162_0[2]),.dinb(w_n308_36[0]),.dout(n1998),.clk(gclk));
	jor g1736(.dina(n1998),.dinb(n1997),.dout(n1999),.clk(gclk));
	jor g1737(.dina(n1999),.dinb(n1996),.dout(n2000),.clk(gclk));
	jand g1738(.dina(w_n2000_1[1]),.dinb(w_n432_56[2]),.dout(n2001),.clk(gclk));
	jand g1739(.dina(w_n1301_0[2]),.dinb(w_n266_35[2]),.dout(n2002),.clk(gclk));
	jand g1740(.dina(w_n1181_0[2]),.dinb(w_n281_35[2]),.dout(n2003),.clk(gclk));
	jor g1741(.dina(n2003),.dinb(n2002),.dout(n2004),.clk(gclk));
	jand g1742(.dina(w_n1318_0[2]),.dinb(w_n295_35[2]),.dout(n2005),.clk(gclk));
	jand g1743(.dina(w_n1198_0[2]),.dinb(w_n308_35[2]),.dout(n2006),.clk(gclk));
	jor g1744(.dina(n2006),.dinb(n2005),.dout(n2007),.clk(gclk));
	jor g1745(.dina(n2007),.dinb(n2004),.dout(n2008),.clk(gclk));
	jand g1746(.dina(w_n2008_1[1]),.dinb(w_n485_56[2]),.dout(n2009),.clk(gclk));
	jor g1747(.dina(n2009),.dinb(n2001),.dout(n2010),.clk(gclk));
	jor g1748(.dina(n2010),.dinb(n1993),.dout(n2011),.clk(gclk));
	jand g1749(.dina(w_n2011_0[1]),.dinb(w_n263_60[0]),.dout(n2012),.clk(gclk));
	jand g1750(.dina(w_n1228_0[2]),.dinb(w_n266_35[1]),.dout(n2013),.clk(gclk));
	jand g1751(.dina(w_n1329_0[2]),.dinb(w_n281_35[1]),.dout(n2014),.clk(gclk));
	jor g1752(.dina(n2014),.dinb(n2013),.dout(n2015),.clk(gclk));
	jand g1753(.dina(w_n1245_0[2]),.dinb(w_n295_35[1]),.dout(n2016),.clk(gclk));
	jand g1754(.dina(w_n1346_0[2]),.dinb(w_n308_35[1]),.dout(n2017),.clk(gclk));
	jor g1755(.dina(n2017),.dinb(n2016),.dout(n2018),.clk(gclk));
	jor g1756(.dina(n2018),.dinb(n2015),.dout(n2019),.clk(gclk));
	jand g1757(.dina(w_n2019_1[1]),.dinb(w_n377_56[1]),.dout(n2020),.clk(gclk));
	jand g1758(.dina(w_n1264_0[2]),.dinb(w_n266_35[0]),.dout(n2021),.clk(gclk));
	jand g1759(.dina(w_n1293_0[2]),.dinb(w_n281_35[0]),.dout(n2022),.clk(gclk));
	jor g1760(.dina(n2022),.dinb(n2021),.dout(n2023),.clk(gclk));
	jand g1761(.dina(w_n1281_0[2]),.dinb(w_n295_35[0]),.dout(n2024),.clk(gclk));
	jand g1762(.dina(w_n1310_0[2]),.dinb(w_n308_35[0]),.dout(n2025),.clk(gclk));
	jor g1763(.dina(n2025),.dinb(n2024),.dout(n2026),.clk(gclk));
	jor g1764(.dina(n2026),.dinb(n2023),.dout(n2027),.clk(gclk));
	jand g1765(.dina(w_n2027_1[1]),.dinb(w_n323_56[1]),.dout(n2028),.clk(gclk));
	jor g1766(.dina(n2028),.dinb(n2020),.dout(n2029),.clk(gclk));
	jand g1767(.dina(w_n1080_0[2]),.dinb(w_n266_34[2]),.dout(n2030),.clk(gclk));
	jand g1768(.dina(w_n1220_0[2]),.dinb(w_n281_34[2]),.dout(n2031),.clk(gclk));
	jor g1769(.dina(n2031),.dinb(n2030),.dout(n2032),.clk(gclk));
	jand g1770(.dina(w_n1097_0[2]),.dinb(w_n295_34[2]),.dout(n2033),.clk(gclk));
	jand g1771(.dina(w_n1237_0[2]),.dinb(w_n308_34[2]),.dout(n2034),.clk(gclk));
	jor g1772(.dina(n2034),.dinb(n2033),.dout(n2035),.clk(gclk));
	jor g1773(.dina(n2035),.dinb(n2032),.dout(n2036),.clk(gclk));
	jand g1774(.dina(w_n2036_1[1]),.dinb(w_n485_56[1]),.dout(n2037),.clk(gclk));
	jand g1775(.dina(w_n1337_0[2]),.dinb(w_n266_34[1]),.dout(n2038),.clk(gclk));
	jand g1776(.dina(w_n1256_0[2]),.dinb(w_n281_34[1]),.dout(n2039),.clk(gclk));
	jor g1777(.dina(n2039),.dinb(n2038),.dout(n2040),.clk(gclk));
	jand g1778(.dina(w_n1354_0[2]),.dinb(w_n295_34[1]),.dout(n2041),.clk(gclk));
	jand g1779(.dina(w_n1273_0[2]),.dinb(w_n308_34[1]),.dout(n2042),.clk(gclk));
	jor g1780(.dina(n2042),.dinb(n2041),.dout(n2043),.clk(gclk));
	jor g1781(.dina(n2043),.dinb(n2040),.dout(n2044),.clk(gclk));
	jand g1782(.dina(w_n2044_1[1]),.dinb(w_n432_56[1]),.dout(n2045),.clk(gclk));
	jor g1783(.dina(n2045),.dinb(n2037),.dout(n2046),.clk(gclk));
	jor g1784(.dina(n2046),.dinb(n2029),.dout(n2047),.clk(gclk));
	jand g1785(.dina(w_n2047_0[1]),.dinb(w_shift6_60[0]),.dout(n2048),.clk(gclk));
	jor g1786(.dina(n2048),.dinb(n2012),.dout(result10),.clk(gclk));
	jand g1787(.dina(w_n1410_0[2]),.dinb(w_n266_34[0]),.dout(n2050),.clk(gclk));
	jand g1788(.dina(w_n1385_0[2]),.dinb(w_n281_34[0]),.dout(n2051),.clk(gclk));
	jor g1789(.dina(n2051),.dinb(n2050),.dout(n2052),.clk(gclk));
	jand g1790(.dina(w_n1419_0[2]),.dinb(w_n295_34[0]),.dout(n2053),.clk(gclk));
	jand g1791(.dina(w_n1394_0[2]),.dinb(w_n308_34[0]),.dout(n2054),.clk(gclk));
	jor g1792(.dina(n2054),.dinb(n2053),.dout(n2055),.clk(gclk));
	jor g1793(.dina(n2055),.dinb(n2052),.dout(n2056),.clk(gclk));
	jand g1794(.dina(w_n2056_1[1]),.dinb(w_n323_56[0]),.dout(n2057),.clk(gclk));
	jand g1795(.dina(w_n1430_0[2]),.dinb(w_n266_33[2]),.dout(n2058),.clk(gclk));
	jand g1796(.dina(w_n1365_0[2]),.dinb(w_n281_33[2]),.dout(n2059),.clk(gclk));
	jor g1797(.dina(n2059),.dinb(n2058),.dout(n2060),.clk(gclk));
	jand g1798(.dina(w_n1439_0[2]),.dinb(w_n295_33[2]),.dout(n2061),.clk(gclk));
	jand g1799(.dina(w_n1374_0[2]),.dinb(w_n308_33[2]),.dout(n2062),.clk(gclk));
	jor g1800(.dina(n2062),.dinb(n2061),.dout(n2063),.clk(gclk));
	jor g1801(.dina(n2063),.dinb(n2060),.dout(n2064),.clk(gclk));
	jand g1802(.dina(w_n2064_1[1]),.dinb(w_n377_56[0]),.dout(n2065),.clk(gclk));
	jor g1803(.dina(n2065),.dinb(n2057),.dout(n2066),.clk(gclk));
	jand g1804(.dina(w_n1369_0[2]),.dinb(w_n266_33[1]),.dout(n2067),.clk(gclk));
	jand g1805(.dina(w_n1406_0[2]),.dinb(w_n281_33[1]),.dout(n2068),.clk(gclk));
	jor g1806(.dina(n2068),.dinb(n2067),.dout(n2069),.clk(gclk));
	jand g1807(.dina(w_n1378_0[2]),.dinb(w_n295_33[1]),.dout(n2070),.clk(gclk));
	jand g1808(.dina(w_n1415_0[2]),.dinb(w_n308_33[1]),.dout(n2071),.clk(gclk));
	jor g1809(.dina(n2071),.dinb(n2070),.dout(n2072),.clk(gclk));
	jor g1810(.dina(n2072),.dinb(n2069),.dout(n2073),.clk(gclk));
	jand g1811(.dina(w_n2073_1[1]),.dinb(w_n432_56[0]),.dout(n2074),.clk(gclk));
	jand g1812(.dina(w_n1521_0[2]),.dinb(w_n266_33[0]),.dout(n2075),.clk(gclk));
	jand g1813(.dina(w_n1426_0[2]),.dinb(w_n281_33[0]),.dout(n2076),.clk(gclk));
	jor g1814(.dina(n2076),.dinb(n2075),.dout(n2077),.clk(gclk));
	jand g1815(.dina(w_n1530_0[2]),.dinb(w_n295_33[0]),.dout(n2078),.clk(gclk));
	jand g1816(.dina(w_n1435_0[2]),.dinb(w_n308_33[0]),.dout(n2079),.clk(gclk));
	jor g1817(.dina(n2079),.dinb(n2078),.dout(n2080),.clk(gclk));
	jor g1818(.dina(n2080),.dinb(n2077),.dout(n2081),.clk(gclk));
	jand g1819(.dina(w_n2081_1[1]),.dinb(w_n485_56[0]),.dout(n2082),.clk(gclk));
	jor g1820(.dina(n2082),.dinb(n2074),.dout(n2083),.clk(gclk));
	jor g1821(.dina(n2083),.dinb(n2066),.dout(n2084),.clk(gclk));
	jand g1822(.dina(w_n2084_0[1]),.dinb(w_n263_59[2]),.dout(n2085),.clk(gclk));
	jand g1823(.dina(w_n1453_0[2]),.dinb(w_n266_32[2]),.dout(n2086),.clk(gclk));
	jand g1824(.dina(w_n1462_0[2]),.dinb(w_n295_32[2]),.dout(n2087),.clk(gclk));
	jor g1825(.dina(n2087),.dinb(n2086),.dout(n2088),.clk(gclk));
	jand g1826(.dina(w_n1490_0[2]),.dinb(w_n281_32[2]),.dout(n2089),.clk(gclk));
	jand g1827(.dina(w_n1505_0[2]),.dinb(w_n308_32[2]),.dout(n2090),.clk(gclk));
	jor g1828(.dina(n2090),.dinb(n2089),.dout(n2091),.clk(gclk));
	jor g1829(.dina(n2091),.dinb(n2088),.dout(n2092),.clk(gclk));
	jand g1830(.dina(w_n2092_1[1]),.dinb(w_n377_55[2]),.dout(n2093),.clk(gclk));
	jand g1831(.dina(w_n1473_0[2]),.dinb(w_n266_32[1]),.dout(n2094),.clk(gclk));
	jand g1832(.dina(w_n1517_0[2]),.dinb(w_n281_32[1]),.dout(n2095),.clk(gclk));
	jor g1833(.dina(n2095),.dinb(n2094),.dout(n2096),.clk(gclk));
	jand g1834(.dina(w_n1482_0[2]),.dinb(w_n295_32[1]),.dout(n2097),.clk(gclk));
	jand g1835(.dina(w_n1526_0[2]),.dinb(w_n308_32[1]),.dout(n2098),.clk(gclk));
	jor g1836(.dina(n2098),.dinb(n2097),.dout(n2099),.clk(gclk));
	jor g1837(.dina(n2099),.dinb(n2096),.dout(n2100),.clk(gclk));
	jand g1838(.dina(w_n2100_1[1]),.dinb(w_n323_55[2]),.dout(n2101),.clk(gclk));
	jor g1839(.dina(n2101),.dinb(n2093),.dout(n2102),.clk(gclk));
	jand g1840(.dina(w_n1389_0[2]),.dinb(w_n266_32[0]),.dout(n2103),.clk(gclk));
	jand g1841(.dina(w_n1449_0[2]),.dinb(w_n281_32[0]),.dout(n2104),.clk(gclk));
	jor g1842(.dina(n2104),.dinb(n2103),.dout(n2105),.clk(gclk));
	jand g1843(.dina(w_n1398_0[2]),.dinb(w_n295_32[0]),.dout(n2106),.clk(gclk));
	jand g1844(.dina(w_n1458_0[2]),.dinb(w_n308_32[0]),.dout(n2107),.clk(gclk));
	jor g1845(.dina(n2107),.dinb(n2106),.dout(n2108),.clk(gclk));
	jor g1846(.dina(n2108),.dinb(n2105),.dout(n2109),.clk(gclk));
	jand g1847(.dina(w_n2109_1[1]),.dinb(w_n485_55[2]),.dout(n2110),.clk(gclk));
	jand g1848(.dina(w_n1496_0[2]),.dinb(w_n266_31[2]),.dout(n2111),.clk(gclk));
	jand g1849(.dina(w_n1469_0[2]),.dinb(w_n281_31[2]),.dout(n2112),.clk(gclk));
	jor g1850(.dina(n2112),.dinb(n2111),.dout(n2113),.clk(gclk));
	jand g1851(.dina(w_n1510_0[2]),.dinb(w_n295_31[2]),.dout(n2114),.clk(gclk));
	jand g1852(.dina(w_n1478_0[2]),.dinb(w_n308_31[2]),.dout(n2115),.clk(gclk));
	jor g1853(.dina(n2115),.dinb(n2114),.dout(n2116),.clk(gclk));
	jor g1854(.dina(n2116),.dinb(n2113),.dout(n2117),.clk(gclk));
	jand g1855(.dina(w_n2117_1[1]),.dinb(w_n432_55[2]),.dout(n2118),.clk(gclk));
	jor g1856(.dina(n2118),.dinb(n2110),.dout(n2119),.clk(gclk));
	jor g1857(.dina(n2119),.dinb(n2102),.dout(n2120),.clk(gclk));
	jand g1858(.dina(w_n2120_0[1]),.dinb(w_shift6_59[2]),.dout(n2121),.clk(gclk));
	jor g1859(.dina(n2121),.dinb(n2085),.dout(result11),.clk(gclk));
	jand g1860(.dina(w_n415_0[1]),.dinb(w_n266_31[1]),.dout(n2123),.clk(gclk));
	jand g1861(.dina(w_n427_0[1]),.dinb(w_n281_31[1]),.dout(n2124),.clk(gclk));
	jor g1862(.dina(n2124),.dinb(n2123),.dout(n2125),.clk(gclk));
	jand g1863(.dina(w_n402_0[1]),.dinb(w_n295_31[1]),.dout(n2126),.clk(gclk));
	jand g1864(.dina(w_n308_31[1]),.dinb(w_n279_0[1]),.dout(n2127),.clk(gclk));
	jor g1865(.dina(n2127),.dinb(n2126),.dout(n2128),.clk(gclk));
	jor g1866(.dina(n2128),.dinb(n2125),.dout(n2129),.clk(gclk));
	jand g1867(.dina(w_n2129_1[1]),.dinb(w_n323_55[1]),.dout(n2130),.clk(gclk));
	jand g1868(.dina(w_n469_0[1]),.dinb(w_n266_31[0]),.dout(n2131),.clk(gclk));
	jand g1869(.dina(w_n481_0[1]),.dinb(w_n281_31[0]),.dout(n2132),.clk(gclk));
	jor g1870(.dina(n2132),.dinb(n2131),.dout(n2133),.clk(gclk));
	jand g1871(.dina(w_n456_0[1]),.dinb(w_n295_31[0]),.dout(n2134),.clk(gclk));
	jand g1872(.dina(w_n335_0[1]),.dinb(w_n308_31[0]),.dout(n2135),.clk(gclk));
	jor g1873(.dina(n2135),.dinb(n2134),.dout(n2136),.clk(gclk));
	jor g1874(.dina(n2136),.dinb(n2133),.dout(n2137),.clk(gclk));
	jand g1875(.dina(w_n2137_1[1]),.dinb(w_n377_55[1]),.dout(n2138),.clk(gclk));
	jor g1876(.dina(n2138),.dinb(n2130),.dout(n2139),.clk(gclk));
	jand g1877(.dina(w_n360_0[1]),.dinb(w_n266_30[2]),.dout(n2140),.clk(gclk));
	jand g1878(.dina(w_n372_0[1]),.dinb(w_n281_30[2]),.dout(n2141),.clk(gclk));
	jor g1879(.dina(n2141),.dinb(n2140),.dout(n2142),.clk(gclk));
	jand g1880(.dina(w_n347_0[1]),.dinb(w_n295_30[2]),.dout(n2143),.clk(gclk));
	jand g1881(.dina(w_n390_0[1]),.dinb(w_n308_30[2]),.dout(n2144),.clk(gclk));
	jor g1882(.dina(n2144),.dinb(n2143),.dout(n2145),.clk(gclk));
	jor g1883(.dina(n2145),.dinb(n2142),.dout(n2146),.clk(gclk));
	jand g1884(.dina(w_n2146_1[1]),.dinb(w_n432_55[1]),.dout(n2147),.clk(gclk));
	jand g1885(.dina(w_n525_0[1]),.dinb(w_n266_30[1]),.dout(n2148),.clk(gclk));
	jand g1886(.dina(w_n537_0[1]),.dinb(w_n281_30[1]),.dout(n2149),.clk(gclk));
	jor g1887(.dina(n2149),.dinb(n2148),.dout(n2150),.clk(gclk));
	jand g1888(.dina(w_n512_0[1]),.dinb(w_n295_30[1]),.dout(n2151),.clk(gclk));
	jand g1889(.dina(w_n444_0[1]),.dinb(w_n308_30[1]),.dout(n2152),.clk(gclk));
	jor g1890(.dina(n2152),.dinb(n2151),.dout(n2153),.clk(gclk));
	jor g1891(.dina(n2153),.dinb(n2150),.dout(n2154),.clk(gclk));
	jand g1892(.dina(w_n2154_1[1]),.dinb(w_n485_55[1]),.dout(n2155),.clk(gclk));
	jor g1893(.dina(n2155),.dinb(n2147),.dout(n2156),.clk(gclk));
	jor g1894(.dina(n2156),.dinb(n2139),.dout(n2157),.clk(gclk));
	jand g1895(.dina(w_n2157_0[1]),.dinb(w_n263_59[1]),.dout(n2158),.clk(gclk));
	jand g1896(.dina(w_n680_0[1]),.dinb(w_n266_30[0]),.dout(n2159),.clk(gclk));
	jand g1897(.dina(w_n692_0[1]),.dinb(w_n281_30[0]),.dout(n2160),.clk(gclk));
	jor g1898(.dina(n2160),.dinb(n2159),.dout(n2161),.clk(gclk));
	jand g1899(.dina(w_n667_0[1]),.dinb(w_n295_30[0]),.dout(n2162),.clk(gclk));
	jand g1900(.dina(w_n552_0[1]),.dinb(w_n308_30[0]),.dout(n2163),.clk(gclk));
	jor g1901(.dina(n2163),.dinb(n2162),.dout(n2164),.clk(gclk));
	jor g1902(.dina(n2164),.dinb(n2161),.dout(n2165),.clk(gclk));
	jand g1903(.dina(w_n2165_1[1]),.dinb(w_n377_55[0]),.dout(n2166),.clk(gclk));
	jand g1904(.dina(w_n628_0[1]),.dinb(w_n266_29[2]),.dout(n2167),.clk(gclk));
	jand g1905(.dina(w_n640_0[1]),.dinb(w_n281_29[2]),.dout(n2168),.clk(gclk));
	jor g1906(.dina(n2168),.dinb(n2167),.dout(n2169),.clk(gclk));
	jand g1907(.dina(w_n615_0[1]),.dinb(w_n295_29[2]),.dout(n2170),.clk(gclk));
	jand g1908(.dina(w_n500_0[1]),.dinb(w_n308_29[2]),.dout(n2171),.clk(gclk));
	jor g1909(.dina(n2171),.dinb(n2170),.dout(n2172),.clk(gclk));
	jor g1910(.dina(n2172),.dinb(n2169),.dout(n2173),.clk(gclk));
	jand g1911(.dina(w_n2173_1[1]),.dinb(w_n323_55[0]),.dout(n2174),.clk(gclk));
	jor g1912(.dina(n2174),.dinb(n2166),.dout(n2175),.clk(gclk));
	jand g1913(.dina(w_n306_0[1]),.dinb(w_n266_29[1]),.dout(n2176),.clk(gclk));
	jand g1914(.dina(w_n319_0[1]),.dinb(w_n281_29[1]),.dout(n2177),.clk(gclk));
	jor g1915(.dina(n2177),.dinb(n2176),.dout(n2178),.clk(gclk));
	jand g1916(.dina(w_n295_29[1]),.dinb(w_n292_0[1]),.dout(n2179),.clk(gclk));
	jand g1917(.dina(w_n655_0[1]),.dinb(w_n308_29[1]),.dout(n2180),.clk(gclk));
	jor g1918(.dina(n2180),.dinb(n2179),.dout(n2181),.clk(gclk));
	jor g1919(.dina(n2181),.dinb(n2178),.dout(n2182),.clk(gclk));
	jand g1920(.dina(w_n2182_1[1]),.dinb(w_n485_55[0]),.dout(n2183),.clk(gclk));
	jand g1921(.dina(w_n575_0[1]),.dinb(w_n266_29[0]),.dout(n2184),.clk(gclk));
	jand g1922(.dina(w_n587_0[1]),.dinb(w_n281_29[0]),.dout(n2185),.clk(gclk));
	jor g1923(.dina(n2185),.dinb(n2184),.dout(n2186),.clk(gclk));
	jand g1924(.dina(w_n562_0[1]),.dinb(w_n295_29[0]),.dout(n2187),.clk(gclk));
	jand g1925(.dina(w_n603_0[1]),.dinb(w_n308_29[0]),.dout(n2188),.clk(gclk));
	jor g1926(.dina(n2188),.dinb(n2187),.dout(n2189),.clk(gclk));
	jor g1927(.dina(n2189),.dinb(n2186),.dout(n2190),.clk(gclk));
	jand g1928(.dina(w_n2190_1[1]),.dinb(w_n432_55[0]),.dout(n2191),.clk(gclk));
	jor g1929(.dina(n2191),.dinb(n2183),.dout(n2192),.clk(gclk));
	jor g1930(.dina(n2192),.dinb(n2175),.dout(n2193),.clk(gclk));
	jand g1931(.dina(w_n2193_0[1]),.dinb(w_shift6_59[1]),.dout(n2194),.clk(gclk));
	jor g1932(.dina(n2194),.dinb(n2158),.dout(result12),.clk(gclk));
	jand g1933(.dina(w_n819_0[1]),.dinb(w_n266_28[2]),.dout(n2196),.clk(gclk));
	jand g1934(.dina(w_n829_0[1]),.dinb(w_n281_28[2]),.dout(n2197),.clk(gclk));
	jor g1935(.dina(n2197),.dinb(n2196),.dout(n2198),.clk(gclk));
	jand g1936(.dina(w_n808_0[1]),.dinb(w_n295_28[2]),.dout(n2199),.clk(gclk));
	jand g1937(.dina(w_n709_0[1]),.dinb(w_n308_28[2]),.dout(n2200),.clk(gclk));
	jor g1938(.dina(n2200),.dinb(n2199),.dout(n2201),.clk(gclk));
	jor g1939(.dina(n2201),.dinb(n2198),.dout(n2202),.clk(gclk));
	jand g1940(.dina(w_n2202_1[1]),.dinb(w_n323_54[2]),.dout(n2203),.clk(gclk));
	jand g1941(.dina(w_n863_0[1]),.dinb(w_n266_28[1]),.dout(n2204),.clk(gclk));
	jand g1942(.dina(w_n873_0[1]),.dinb(w_n281_28[1]),.dout(n2205),.clk(gclk));
	jor g1943(.dina(n2205),.dinb(n2204),.dout(n2206),.clk(gclk));
	jand g1944(.dina(w_n852_0[1]),.dinb(w_n295_28[1]),.dout(n2207),.clk(gclk));
	jand g1945(.dina(w_n753_0[1]),.dinb(w_n308_28[1]),.dout(n2208),.clk(gclk));
	jor g1946(.dina(n2208),.dinb(n2207),.dout(n2209),.clk(gclk));
	jor g1947(.dina(n2209),.dinb(n2206),.dout(n2210),.clk(gclk));
	jand g1948(.dina(w_n2210_1[1]),.dinb(w_n377_54[2]),.dout(n2211),.clk(gclk));
	jor g1949(.dina(n2211),.dinb(n2203),.dout(n2212),.clk(gclk));
	jand g1950(.dina(w_n774_0[1]),.dinb(w_n266_28[0]),.dout(n2213),.clk(gclk));
	jand g1951(.dina(w_n784_0[1]),.dinb(w_n281_28[0]),.dout(n2214),.clk(gclk));
	jor g1952(.dina(n2214),.dinb(n2213),.dout(n2215),.clk(gclk));
	jand g1953(.dina(w_n763_0[1]),.dinb(w_n295_28[0]),.dout(n2216),.clk(gclk));
	jand g1954(.dina(w_n798_0[1]),.dinb(w_n308_28[0]),.dout(n2217),.clk(gclk));
	jor g1955(.dina(n2217),.dinb(n2216),.dout(n2218),.clk(gclk));
	jor g1956(.dina(n2218),.dinb(n2215),.dout(n2219),.clk(gclk));
	jand g1957(.dina(w_n2219_1[1]),.dinb(w_n432_54[2]),.dout(n2220),.clk(gclk));
	jand g1958(.dina(w_n999_0[1]),.dinb(w_n266_27[2]),.dout(n2221),.clk(gclk));
	jand g1959(.dina(w_n1009_0[1]),.dinb(w_n281_27[2]),.dout(n2222),.clk(gclk));
	jor g1960(.dina(n2222),.dinb(n2221),.dout(n2223),.clk(gclk));
	jand g1961(.dina(w_n988_0[1]),.dinb(w_n295_27[2]),.dout(n2224),.clk(gclk));
	jand g1962(.dina(w_n842_0[1]),.dinb(w_n308_27[2]),.dout(n2225),.clk(gclk));
	jor g1963(.dina(n2225),.dinb(n2224),.dout(n2226),.clk(gclk));
	jor g1964(.dina(n2226),.dinb(n2223),.dout(n2227),.clk(gclk));
	jand g1965(.dina(w_n2227_1[1]),.dinb(w_n485_54[2]),.dout(n2228),.clk(gclk));
	jor g1966(.dina(n2228),.dinb(n2220),.dout(n2229),.clk(gclk));
	jor g1967(.dina(n2229),.dinb(n2212),.dout(n2230),.clk(gclk));
	jand g1968(.dina(w_n2230_0[1]),.dinb(w_n263_59[0]),.dout(n2231),.clk(gclk));
	jand g1969(.dina(w_n910_0[1]),.dinb(w_n266_27[1]),.dout(n2232),.clk(gclk));
	jand g1970(.dina(w_n920_0[1]),.dinb(w_n281_27[1]),.dout(n2233),.clk(gclk));
	jor g1971(.dina(n2233),.dinb(n2232),.dout(n2234),.clk(gclk));
	jand g1972(.dina(w_n899_0[1]),.dinb(w_n295_27[1]),.dout(n2235),.clk(gclk));
	jand g1973(.dina(w_n1022_0[1]),.dinb(w_n308_27[1]),.dout(n2236),.clk(gclk));
	jor g1974(.dina(n2236),.dinb(n2235),.dout(n2237),.clk(gclk));
	jor g1975(.dina(n2237),.dinb(n2234),.dout(n2238),.clk(gclk));
	jand g1976(.dina(w_n2238_1[1]),.dinb(w_n377_54[1]),.dout(n2239),.clk(gclk));
	jand g1977(.dina(w_n954_0[1]),.dinb(w_n266_27[0]),.dout(n2240),.clk(gclk));
	jand g1978(.dina(w_n964_0[1]),.dinb(w_n281_27[0]),.dout(n2241),.clk(gclk));
	jor g1979(.dina(n2241),.dinb(n2240),.dout(n2242),.clk(gclk));
	jand g1980(.dina(w_n943_0[1]),.dinb(w_n295_27[0]),.dout(n2243),.clk(gclk));
	jand g1981(.dina(w_n978_0[1]),.dinb(w_n308_27[0]),.dout(n2244),.clk(gclk));
	jor g1982(.dina(n2244),.dinb(n2243),.dout(n2245),.clk(gclk));
	jor g1983(.dina(n2245),.dinb(n2242),.dout(n2246),.clk(gclk));
	jand g1984(.dina(w_n2246_1[1]),.dinb(w_n323_54[1]),.dout(n2247),.clk(gclk));
	jor g1985(.dina(n2247),.dinb(n2239),.dout(n2248),.clk(gclk));
	jand g1986(.dina(w_n730_0[1]),.dinb(w_n266_26[2]),.dout(n2249),.clk(gclk));
	jand g1987(.dina(w_n740_0[1]),.dinb(w_n281_26[2]),.dout(n2250),.clk(gclk));
	jor g1988(.dina(n2250),.dinb(n2249),.dout(n2251),.clk(gclk));
	jand g1989(.dina(w_n719_0[1]),.dinb(w_n295_26[2]),.dout(n2252),.clk(gclk));
	jand g1990(.dina(w_n889_0[1]),.dinb(w_n308_26[2]),.dout(n2253),.clk(gclk));
	jor g1991(.dina(n2253),.dinb(n2252),.dout(n2254),.clk(gclk));
	jor g1992(.dina(n2254),.dinb(n2251),.dout(n2255),.clk(gclk));
	jand g1993(.dina(w_n2255_1[1]),.dinb(w_n485_54[1]),.dout(n2256),.clk(gclk));
	jand g1994(.dina(w_n1047_0[1]),.dinb(w_n266_26[1]),.dout(n2257),.clk(gclk));
	jand g1995(.dina(w_n1057_0[1]),.dinb(w_n281_26[1]),.dout(n2258),.clk(gclk));
	jor g1996(.dina(n2258),.dinb(n2257),.dout(n2259),.clk(gclk));
	jand g1997(.dina(w_n1034_0[1]),.dinb(w_n295_26[1]),.dout(n2260),.clk(gclk));
	jand g1998(.dina(w_n933_0[1]),.dinb(w_n308_26[1]),.dout(n2261),.clk(gclk));
	jor g1999(.dina(n2261),.dinb(n2260),.dout(n2262),.clk(gclk));
	jor g2000(.dina(n2262),.dinb(n2259),.dout(n2263),.clk(gclk));
	jand g2001(.dina(w_n2263_1[1]),.dinb(w_n432_54[1]),.dout(n2264),.clk(gclk));
	jor g2002(.dina(n2264),.dinb(n2256),.dout(n2265),.clk(gclk));
	jor g2003(.dina(n2265),.dinb(n2248),.dout(n2266),.clk(gclk));
	jand g2004(.dina(w_n2266_0[1]),.dinb(w_shift6_59[0]),.dout(n2267),.clk(gclk));
	jor g2005(.dina(n2267),.dinb(n2231),.dout(result13),.clk(gclk));
	jand g2006(.dina(w_n1162_0[1]),.dinb(w_n266_26[0]),.dout(n2269),.clk(gclk));
	jand g2007(.dina(w_n1170_0[1]),.dinb(w_n281_26[0]),.dout(n2270),.clk(gclk));
	jor g2008(.dina(n2270),.dinb(n2269),.dout(n2271),.clk(gclk));
	jand g2009(.dina(w_n1153_0[1]),.dinb(w_n295_26[0]),.dout(n2272),.clk(gclk));
	jand g2010(.dina(w_n1072_0[1]),.dinb(w_n308_26[0]),.dout(n2273),.clk(gclk));
	jor g2011(.dina(n2273),.dinb(n2272),.dout(n2274),.clk(gclk));
	jor g2012(.dina(n2274),.dinb(n2271),.dout(n2275),.clk(gclk));
	jand g2013(.dina(w_n2275_1[1]),.dinb(w_n323_54[0]),.dout(n2276),.clk(gclk));
	jand g2014(.dina(w_n1198_0[1]),.dinb(w_n266_25[2]),.dout(n2277),.clk(gclk));
	jand g2015(.dina(w_n1206_0[1]),.dinb(w_n281_25[2]),.dout(n2278),.clk(gclk));
	jor g2016(.dina(n2278),.dinb(n2277),.dout(n2279),.clk(gclk));
	jand g2017(.dina(w_n1189_0[1]),.dinb(w_n295_25[2]),.dout(n2280),.clk(gclk));
	jand g2018(.dina(w_n1108_0[1]),.dinb(w_n308_25[2]),.dout(n2281),.clk(gclk));
	jor g2019(.dina(n2281),.dinb(n2280),.dout(n2282),.clk(gclk));
	jor g2020(.dina(n2282),.dinb(n2279),.dout(n2283),.clk(gclk));
	jand g2021(.dina(w_n2283_1[1]),.dinb(w_n377_54[0]),.dout(n2284),.clk(gclk));
	jor g2022(.dina(n2284),.dinb(n2276),.dout(n2285),.clk(gclk));
	jand g2023(.dina(w_n1125_0[1]),.dinb(w_n266_25[1]),.dout(n2286),.clk(gclk));
	jand g2024(.dina(w_n1133_0[1]),.dinb(w_n281_25[1]),.dout(n2287),.clk(gclk));
	jor g2025(.dina(n2287),.dinb(n2286),.dout(n2288),.clk(gclk));
	jand g2026(.dina(w_n1116_0[1]),.dinb(w_n295_25[1]),.dout(n2289),.clk(gclk));
	jand g2027(.dina(w_n1145_0[1]),.dinb(w_n308_25[1]),.dout(n2290),.clk(gclk));
	jor g2028(.dina(n2290),.dinb(n2289),.dout(n2291),.clk(gclk));
	jor g2029(.dina(n2291),.dinb(n2288),.dout(n2292),.clk(gclk));
	jand g2030(.dina(w_n2292_1[1]),.dinb(w_n432_54[0]),.dout(n2293),.clk(gclk));
	jand g2031(.dina(w_n1310_0[1]),.dinb(w_n266_25[0]),.dout(n2294),.clk(gclk));
	jand g2032(.dina(w_n1318_0[1]),.dinb(w_n281_25[0]),.dout(n2295),.clk(gclk));
	jor g2033(.dina(n2295),.dinb(n2294),.dout(n2296),.clk(gclk));
	jand g2034(.dina(w_n1301_0[1]),.dinb(w_n295_25[0]),.dout(n2297),.clk(gclk));
	jand g2035(.dina(w_n1181_0[1]),.dinb(w_n308_25[0]),.dout(n2298),.clk(gclk));
	jor g2036(.dina(n2298),.dinb(n2297),.dout(n2299),.clk(gclk));
	jor g2037(.dina(n2299),.dinb(n2296),.dout(n2300),.clk(gclk));
	jand g2038(.dina(w_n2300_1[1]),.dinb(w_n485_54[0]),.dout(n2301),.clk(gclk));
	jor g2039(.dina(n2301),.dinb(n2293),.dout(n2302),.clk(gclk));
	jor g2040(.dina(n2302),.dinb(n2285),.dout(n2303),.clk(gclk));
	jand g2041(.dina(w_n2303_0[1]),.dinb(w_n263_58[2]),.dout(n2304),.clk(gclk));
	jand g2042(.dina(w_n1237_0[1]),.dinb(w_n266_24[2]),.dout(n2305),.clk(gclk));
	jand g2043(.dina(w_n1245_0[1]),.dinb(w_n281_24[2]),.dout(n2306),.clk(gclk));
	jor g2044(.dina(n2306),.dinb(n2305),.dout(n2307),.clk(gclk));
	jand g2045(.dina(w_n1228_0[1]),.dinb(w_n295_24[2]),.dout(n2308),.clk(gclk));
	jand g2046(.dina(w_n1329_0[1]),.dinb(w_n308_24[2]),.dout(n2309),.clk(gclk));
	jor g2047(.dina(n2309),.dinb(n2308),.dout(n2310),.clk(gclk));
	jor g2048(.dina(n2310),.dinb(n2307),.dout(n2311),.clk(gclk));
	jand g2049(.dina(w_n2311_1[1]),.dinb(w_n377_53[2]),.dout(n2312),.clk(gclk));
	jand g2050(.dina(w_n1273_0[1]),.dinb(w_n266_24[1]),.dout(n2313),.clk(gclk));
	jand g2051(.dina(w_n1281_0[1]),.dinb(w_n281_24[1]),.dout(n2314),.clk(gclk));
	jor g2052(.dina(n2314),.dinb(n2313),.dout(n2315),.clk(gclk));
	jand g2053(.dina(w_n1264_0[1]),.dinb(w_n295_24[1]),.dout(n2316),.clk(gclk));
	jand g2054(.dina(w_n1293_0[1]),.dinb(w_n308_24[1]),.dout(n2317),.clk(gclk));
	jor g2055(.dina(n2317),.dinb(n2316),.dout(n2318),.clk(gclk));
	jor g2056(.dina(n2318),.dinb(n2315),.dout(n2319),.clk(gclk));
	jand g2057(.dina(w_n2319_1[1]),.dinb(w_n323_53[2]),.dout(n2320),.clk(gclk));
	jor g2058(.dina(n2320),.dinb(n2312),.dout(n2321),.clk(gclk));
	jand g2059(.dina(w_n1089_0[1]),.dinb(w_n266_24[0]),.dout(n2322),.clk(gclk));
	jand g2060(.dina(w_n1097_0[1]),.dinb(w_n281_24[0]),.dout(n2323),.clk(gclk));
	jor g2061(.dina(n2323),.dinb(n2322),.dout(n2324),.clk(gclk));
	jand g2062(.dina(w_n1080_0[1]),.dinb(w_n295_24[0]),.dout(n2325),.clk(gclk));
	jand g2063(.dina(w_n1220_0[1]),.dinb(w_n308_24[0]),.dout(n2326),.clk(gclk));
	jor g2064(.dina(n2326),.dinb(n2325),.dout(n2327),.clk(gclk));
	jor g2065(.dina(n2327),.dinb(n2324),.dout(n2328),.clk(gclk));
	jand g2066(.dina(w_n2328_1[1]),.dinb(w_n485_53[2]),.dout(n2329),.clk(gclk));
	jand g2067(.dina(w_n1346_0[1]),.dinb(w_n266_23[2]),.dout(n2330),.clk(gclk));
	jand g2068(.dina(w_n1354_0[1]),.dinb(w_n281_23[2]),.dout(n2331),.clk(gclk));
	jor g2069(.dina(n2331),.dinb(n2330),.dout(n2332),.clk(gclk));
	jand g2070(.dina(w_n1337_0[1]),.dinb(w_n295_23[2]),.dout(n2333),.clk(gclk));
	jand g2071(.dina(w_n1256_0[1]),.dinb(w_n308_23[2]),.dout(n2334),.clk(gclk));
	jor g2072(.dina(n2334),.dinb(n2333),.dout(n2335),.clk(gclk));
	jor g2073(.dina(n2335),.dinb(n2332),.dout(n2336),.clk(gclk));
	jand g2074(.dina(w_n2336_1[1]),.dinb(w_n432_53[2]),.dout(n2337),.clk(gclk));
	jor g2075(.dina(n2337),.dinb(n2329),.dout(n2338),.clk(gclk));
	jor g2076(.dina(n2338),.dinb(n2321),.dout(n2339),.clk(gclk));
	jand g2077(.dina(w_n2339_0[1]),.dinb(w_shift6_58[2]),.dout(n2340),.clk(gclk));
	jor g2078(.dina(n2340),.dinb(n2304),.dout(result14),.clk(gclk));
	jand g2079(.dina(w_n1415_0[1]),.dinb(w_n266_23[1]),.dout(n2342),.clk(gclk));
	jand g2080(.dina(w_n1419_0[1]),.dinb(w_n281_23[1]),.dout(n2343),.clk(gclk));
	jor g2081(.dina(n2343),.dinb(n2342),.dout(n2344),.clk(gclk));
	jand g2082(.dina(w_n1410_0[1]),.dinb(w_n295_23[1]),.dout(n2345),.clk(gclk));
	jand g2083(.dina(w_n1385_0[1]),.dinb(w_n308_23[1]),.dout(n2346),.clk(gclk));
	jor g2084(.dina(n2346),.dinb(n2345),.dout(n2347),.clk(gclk));
	jor g2085(.dina(n2347),.dinb(n2344),.dout(n2348),.clk(gclk));
	jand g2086(.dina(w_n2348_1[1]),.dinb(w_n323_53[1]),.dout(n2349),.clk(gclk));
	jand g2087(.dina(w_n1435_0[1]),.dinb(w_n266_23[0]),.dout(n2350),.clk(gclk));
	jand g2088(.dina(w_n1439_0[1]),.dinb(w_n281_23[0]),.dout(n2351),.clk(gclk));
	jor g2089(.dina(n2351),.dinb(n2350),.dout(n2352),.clk(gclk));
	jand g2090(.dina(w_n1430_0[1]),.dinb(w_n295_23[0]),.dout(n2353),.clk(gclk));
	jand g2091(.dina(w_n1365_0[1]),.dinb(w_n308_23[0]),.dout(n2354),.clk(gclk));
	jor g2092(.dina(n2354),.dinb(n2353),.dout(n2355),.clk(gclk));
	jor g2093(.dina(n2355),.dinb(n2352),.dout(n2356),.clk(gclk));
	jand g2094(.dina(w_n2356_1[1]),.dinb(w_n377_53[1]),.dout(n2357),.clk(gclk));
	jor g2095(.dina(n2357),.dinb(n2349),.dout(n2358),.clk(gclk));
	jand g2096(.dina(w_n1374_0[1]),.dinb(w_n266_22[2]),.dout(n2359),.clk(gclk));
	jand g2097(.dina(w_n1378_0[1]),.dinb(w_n281_22[2]),.dout(n2360),.clk(gclk));
	jor g2098(.dina(n2360),.dinb(n2359),.dout(n2361),.clk(gclk));
	jand g2099(.dina(w_n1369_0[1]),.dinb(w_n295_22[2]),.dout(n2362),.clk(gclk));
	jand g2100(.dina(w_n1406_0[1]),.dinb(w_n308_22[2]),.dout(n2363),.clk(gclk));
	jor g2101(.dina(n2363),.dinb(n2362),.dout(n2364),.clk(gclk));
	jor g2102(.dina(n2364),.dinb(n2361),.dout(n2365),.clk(gclk));
	jand g2103(.dina(w_n2365_1[1]),.dinb(w_n432_53[1]),.dout(n2366),.clk(gclk));
	jand g2104(.dina(w_n1526_0[1]),.dinb(w_n266_22[1]),.dout(n2367),.clk(gclk));
	jand g2105(.dina(w_n1530_0[1]),.dinb(w_n281_22[1]),.dout(n2368),.clk(gclk));
	jor g2106(.dina(n2368),.dinb(n2367),.dout(n2369),.clk(gclk));
	jand g2107(.dina(w_n1521_0[1]),.dinb(w_n295_22[1]),.dout(n2370),.clk(gclk));
	jand g2108(.dina(w_n1426_0[1]),.dinb(w_n308_22[1]),.dout(n2371),.clk(gclk));
	jor g2109(.dina(n2371),.dinb(n2370),.dout(n2372),.clk(gclk));
	jor g2110(.dina(n2372),.dinb(n2369),.dout(n2373),.clk(gclk));
	jand g2111(.dina(w_n2373_1[1]),.dinb(w_n485_53[1]),.dout(n2374),.clk(gclk));
	jor g2112(.dina(n2374),.dinb(n2366),.dout(n2375),.clk(gclk));
	jor g2113(.dina(n2375),.dinb(n2358),.dout(n2376),.clk(gclk));
	jand g2114(.dina(w_n2376_0[1]),.dinb(w_n263_58[1]),.dout(n2377),.clk(gclk));
	jand g2115(.dina(w_n1458_0[1]),.dinb(w_n266_22[0]),.dout(n2378),.clk(gclk));
	jand g2116(.dina(w_n1462_0[1]),.dinb(w_n281_22[0]),.dout(n2379),.clk(gclk));
	jor g2117(.dina(n2379),.dinb(n2378),.dout(n2380),.clk(gclk));
	jand g2118(.dina(w_n1453_0[1]),.dinb(w_n295_22[0]),.dout(n2381),.clk(gclk));
	jand g2119(.dina(w_n1490_0[1]),.dinb(w_n308_22[0]),.dout(n2382),.clk(gclk));
	jor g2120(.dina(n2382),.dinb(n2381),.dout(n2383),.clk(gclk));
	jor g2121(.dina(n2383),.dinb(n2380),.dout(n2384),.clk(gclk));
	jand g2122(.dina(w_n2384_1[1]),.dinb(w_n377_53[0]),.dout(n2385),.clk(gclk));
	jand g2123(.dina(w_n1478_0[1]),.dinb(w_n266_21[2]),.dout(n2386),.clk(gclk));
	jand g2124(.dina(w_n1482_0[1]),.dinb(w_n281_21[2]),.dout(n2387),.clk(gclk));
	jor g2125(.dina(n2387),.dinb(n2386),.dout(n2388),.clk(gclk));
	jand g2126(.dina(w_n1473_0[1]),.dinb(w_n295_21[2]),.dout(n2389),.clk(gclk));
	jand g2127(.dina(w_n1517_0[1]),.dinb(w_n308_21[2]),.dout(n2390),.clk(gclk));
	jor g2128(.dina(n2390),.dinb(n2389),.dout(n2391),.clk(gclk));
	jor g2129(.dina(n2391),.dinb(n2388),.dout(n2392),.clk(gclk));
	jand g2130(.dina(w_n2392_1[1]),.dinb(w_n323_53[0]),.dout(n2393),.clk(gclk));
	jor g2131(.dina(n2393),.dinb(n2385),.dout(n2394),.clk(gclk));
	jand g2132(.dina(w_n1394_0[1]),.dinb(w_n266_21[1]),.dout(n2395),.clk(gclk));
	jand g2133(.dina(w_n1398_0[1]),.dinb(w_n281_21[1]),.dout(n2396),.clk(gclk));
	jor g2134(.dina(n2396),.dinb(n2395),.dout(n2397),.clk(gclk));
	jand g2135(.dina(w_n1389_0[1]),.dinb(w_n295_21[1]),.dout(n2398),.clk(gclk));
	jand g2136(.dina(w_n1449_0[1]),.dinb(w_n308_21[1]),.dout(n2399),.clk(gclk));
	jor g2137(.dina(n2399),.dinb(n2398),.dout(n2400),.clk(gclk));
	jor g2138(.dina(n2400),.dinb(n2397),.dout(n2401),.clk(gclk));
	jand g2139(.dina(w_n2401_1[1]),.dinb(w_n485_53[0]),.dout(n2402),.clk(gclk));
	jand g2140(.dina(w_n1505_0[1]),.dinb(w_n266_21[0]),.dout(n2403),.clk(gclk));
	jand g2141(.dina(w_n1510_0[1]),.dinb(w_n281_21[0]),.dout(n2404),.clk(gclk));
	jor g2142(.dina(n2404),.dinb(n2403),.dout(n2405),.clk(gclk));
	jand g2143(.dina(w_n1496_0[1]),.dinb(w_n295_21[0]),.dout(n2406),.clk(gclk));
	jand g2144(.dina(w_n1469_0[1]),.dinb(w_n308_21[0]),.dout(n2407),.clk(gclk));
	jor g2145(.dina(n2407),.dinb(n2406),.dout(n2408),.clk(gclk));
	jor g2146(.dina(n2408),.dinb(n2405),.dout(n2409),.clk(gclk));
	jand g2147(.dina(w_n2409_1[1]),.dinb(w_n432_53[0]),.dout(n2410),.clk(gclk));
	jor g2148(.dina(n2410),.dinb(n2402),.dout(n2411),.clk(gclk));
	jor g2149(.dina(n2411),.dinb(n2394),.dout(n2412),.clk(gclk));
	jand g2150(.dina(w_n2412_0[1]),.dinb(w_shift6_58[1]),.dout(n2413),.clk(gclk));
	jor g2151(.dina(n2413),.dinb(n2377),.dout(result15),.clk(gclk));
	jand g2152(.dina(w_n430_1[0]),.dinb(w_n323_52[2]),.dout(n2415),.clk(gclk));
	jand g2153(.dina(w_n484_1[0]),.dinb(w_n377_52[2]),.dout(n2416),.clk(gclk));
	jor g2154(.dina(n2416),.dinb(n2415),.dout(n2417),.clk(gclk));
	jand g2155(.dina(w_n432_52[2]),.dinb(w_n375_1[0]),.dout(n2418),.clk(gclk));
	jand g2156(.dina(w_n540_1[0]),.dinb(w_n485_52[2]),.dout(n2419),.clk(gclk));
	jor g2157(.dina(n2419),.dinb(n2418),.dout(n2420),.clk(gclk));
	jor g2158(.dina(n2420),.dinb(n2417),.dout(n2421),.clk(gclk));
	jand g2159(.dina(w_n2421_0[1]),.dinb(w_n263_58[0]),.dout(n2422),.clk(gclk));
	jand g2160(.dina(w_n485_52[1]),.dinb(w_n322_1[0]),.dout(n2423),.clk(gclk));
	jand g2161(.dina(w_n590_1[0]),.dinb(w_n432_52[1]),.dout(n2424),.clk(gclk));
	jor g2162(.dina(n2424),.dinb(n2423),.dout(n2425),.clk(gclk));
	jand g2163(.dina(w_n643_1[0]),.dinb(w_n323_52[1]),.dout(n2426),.clk(gclk));
	jand g2164(.dina(w_n695_1[0]),.dinb(w_n377_52[1]),.dout(n2427),.clk(gclk));
	jor g2165(.dina(n2427),.dinb(n2426),.dout(n2428),.clk(gclk));
	jor g2166(.dina(n2428),.dinb(n2425),.dout(n2429),.clk(gclk));
	jand g2167(.dina(w_n2429_0[1]),.dinb(w_shift6_58[0]),.dout(n2430),.clk(gclk));
	jor g2168(.dina(n2430),.dinb(n2422),.dout(result16),.clk(gclk));
	jand g2169(.dina(w_n832_1[0]),.dinb(w_n323_52[0]),.dout(n2432),.clk(gclk));
	jand g2170(.dina(w_n876_1[0]),.dinb(w_n377_52[0]),.dout(n2433),.clk(gclk));
	jor g2171(.dina(n2433),.dinb(n2432),.dout(n2434),.clk(gclk));
	jand g2172(.dina(w_n787_1[0]),.dinb(w_n432_52[0]),.dout(n2435),.clk(gclk));
	jand g2173(.dina(w_n1012_1[0]),.dinb(w_n485_52[0]),.dout(n2436),.clk(gclk));
	jor g2174(.dina(n2436),.dinb(n2435),.dout(n2437),.clk(gclk));
	jor g2175(.dina(n2437),.dinb(n2434),.dout(n2438),.clk(gclk));
	jand g2176(.dina(w_n2438_0[1]),.dinb(w_n263_57[2]),.dout(n2439),.clk(gclk));
	jand g2177(.dina(w_n923_1[0]),.dinb(w_n377_51[2]),.dout(n2440),.clk(gclk));
	jand g2178(.dina(w_n967_1[0]),.dinb(w_n323_51[2]),.dout(n2441),.clk(gclk));
	jor g2179(.dina(n2441),.dinb(n2440),.dout(n2442),.clk(gclk));
	jand g2180(.dina(w_n743_1[0]),.dinb(w_n485_51[2]),.dout(n2443),.clk(gclk));
	jand g2181(.dina(w_n1060_1[0]),.dinb(w_n432_51[2]),.dout(n2444),.clk(gclk));
	jor g2182(.dina(n2444),.dinb(n2443),.dout(n2445),.clk(gclk));
	jor g2183(.dina(n2445),.dinb(n2442),.dout(n2446),.clk(gclk));
	jand g2184(.dina(w_n2446_0[1]),.dinb(w_shift6_57[2]),.dout(n2447),.clk(gclk));
	jor g2185(.dina(n2447),.dinb(n2439),.dout(result17),.clk(gclk));
	jand g2186(.dina(w_n1173_1[0]),.dinb(w_n323_51[1]),.dout(n2449),.clk(gclk));
	jand g2187(.dina(w_n1209_1[0]),.dinb(w_n377_51[1]),.dout(n2450),.clk(gclk));
	jor g2188(.dina(n2450),.dinb(n2449),.dout(n2451),.clk(gclk));
	jand g2189(.dina(w_n1136_1[0]),.dinb(w_n432_51[1]),.dout(n2452),.clk(gclk));
	jand g2190(.dina(w_n1321_1[0]),.dinb(w_n485_51[1]),.dout(n2453),.clk(gclk));
	jor g2191(.dina(n2453),.dinb(n2452),.dout(n2454),.clk(gclk));
	jor g2192(.dina(n2454),.dinb(n2451),.dout(n2455),.clk(gclk));
	jand g2193(.dina(w_n2455_0[1]),.dinb(w_n263_57[1]),.dout(n2456),.clk(gclk));
	jand g2194(.dina(w_n1248_1[0]),.dinb(w_n377_51[0]),.dout(n2457),.clk(gclk));
	jand g2195(.dina(w_n1284_1[0]),.dinb(w_n323_51[0]),.dout(n2458),.clk(gclk));
	jor g2196(.dina(n2458),.dinb(n2457),.dout(n2459),.clk(gclk));
	jand g2197(.dina(w_n1100_1[0]),.dinb(w_n485_51[0]),.dout(n2460),.clk(gclk));
	jand g2198(.dina(w_n1357_1[0]),.dinb(w_n432_51[0]),.dout(n2461),.clk(gclk));
	jor g2199(.dina(n2461),.dinb(n2460),.dout(n2462),.clk(gclk));
	jor g2200(.dina(n2462),.dinb(n2459),.dout(n2463),.clk(gclk));
	jand g2201(.dina(w_n2463_0[1]),.dinb(w_shift6_57[1]),.dout(n2464),.clk(gclk));
	jor g2202(.dina(n2464),.dinb(n2456),.dout(result18),.clk(gclk));
	jand g2203(.dina(w_n1381_1[0]),.dinb(w_n432_50[2]),.dout(n2466),.clk(gclk));
	jand g2204(.dina(w_n1533_1[0]),.dinb(w_n485_50[2]),.dout(n2467),.clk(gclk));
	jor g2205(.dina(n2467),.dinb(n2466),.dout(n2468),.clk(gclk));
	jand g2206(.dina(w_n1422_1[0]),.dinb(w_n323_50[2]),.dout(n2469),.clk(gclk));
	jand g2207(.dina(w_n1442_1[0]),.dinb(w_n377_50[2]),.dout(n2470),.clk(gclk));
	jor g2208(.dina(n2470),.dinb(n2469),.dout(n2471),.clk(gclk));
	jor g2209(.dina(n2471),.dinb(n2468),.dout(n2472),.clk(gclk));
	jand g2210(.dina(w_n2472_0[1]),.dinb(w_n263_57[0]),.dout(n2473),.clk(gclk));
	jand g2211(.dina(w_n1465_1[0]),.dinb(w_n377_50[1]),.dout(n2474),.clk(gclk));
	jand g2212(.dina(w_n1513_1[0]),.dinb(w_n432_50[1]),.dout(n2475),.clk(gclk));
	jor g2213(.dina(n2475),.dinb(n2474),.dout(n2476),.clk(gclk));
	jand g2214(.dina(w_n1401_1[0]),.dinb(w_n485_50[1]),.dout(n2477),.clk(gclk));
	jand g2215(.dina(w_n1485_1[0]),.dinb(w_n323_50[1]),.dout(n2478),.clk(gclk));
	jor g2216(.dina(n2478),.dinb(n2477),.dout(n2479),.clk(gclk));
	jor g2217(.dina(n2479),.dinb(n2476),.dout(n2480),.clk(gclk));
	jand g2218(.dina(w_n2480_0[1]),.dinb(w_shift6_57[0]),.dout(n2481),.clk(gclk));
	jor g2219(.dina(n2481),.dinb(n2473),.dout(result19),.clk(gclk));
	jand g2220(.dina(w_n1562_1[0]),.dinb(w_n323_50[0]),.dout(n2483),.clk(gclk));
	jand g2221(.dina(w_n1570_1[0]),.dinb(w_n377_50[0]),.dout(n2484),.clk(gclk));
	jor g2222(.dina(n2484),.dinb(n2483),.dout(n2485),.clk(gclk));
	jand g2223(.dina(w_n1553_1[0]),.dinb(w_n432_50[0]),.dout(n2486),.clk(gclk));
	jand g2224(.dina(w_n1589_1[0]),.dinb(w_n485_50[0]),.dout(n2487),.clk(gclk));
	jor g2225(.dina(n2487),.dinb(n2486),.dout(n2488),.clk(gclk));
	jor g2226(.dina(n2488),.dinb(n2485),.dout(n2489),.clk(gclk));
	jand g2227(.dina(w_n2489_0[1]),.dinb(w_n263_56[2]),.dout(n2490),.clk(gclk));
	jand g2228(.dina(w_n1545_1[0]),.dinb(w_n485_49[2]),.dout(n2491),.clk(gclk));
	jand g2229(.dina(w_n1598_1[0]),.dinb(w_n377_49[2]),.dout(n2492),.clk(gclk));
	jor g2230(.dina(n2492),.dinb(n2491),.dout(n2493),.clk(gclk));
	jand g2231(.dina(w_n1581_1[0]),.dinb(w_n432_49[2]),.dout(n2494),.clk(gclk));
	jand g2232(.dina(w_n1606_1[0]),.dinb(w_n323_49[2]),.dout(n2495),.clk(gclk));
	jor g2233(.dina(n2495),.dinb(n2494),.dout(n2496),.clk(gclk));
	jor g2234(.dina(n2496),.dinb(n2493),.dout(n2497),.clk(gclk));
	jand g2235(.dina(w_n2497_0[1]),.dinb(w_shift6_56[2]),.dout(n2498),.clk(gclk));
	jor g2236(.dina(n2498),.dinb(n2490),.dout(result20),.clk(gclk));
	jand g2237(.dina(w_n1635_1[0]),.dinb(w_n323_49[1]),.dout(n2500),.clk(gclk));
	jand g2238(.dina(w_n1643_1[0]),.dinb(w_n377_49[1]),.dout(n2501),.clk(gclk));
	jor g2239(.dina(n2501),.dinb(n2500),.dout(n2502),.clk(gclk));
	jand g2240(.dina(w_n1626_1[0]),.dinb(w_n432_49[1]),.dout(n2503),.clk(gclk));
	jand g2241(.dina(w_n1662_1[0]),.dinb(w_n485_49[1]),.dout(n2504),.clk(gclk));
	jor g2242(.dina(n2504),.dinb(n2503),.dout(n2505),.clk(gclk));
	jor g2243(.dina(n2505),.dinb(n2502),.dout(n2506),.clk(gclk));
	jand g2244(.dina(w_n2506_0[1]),.dinb(w_n263_56[1]),.dout(n2507),.clk(gclk));
	jand g2245(.dina(w_n1618_1[0]),.dinb(w_n485_49[0]),.dout(n2508),.clk(gclk));
	jand g2246(.dina(w_n1671_1[0]),.dinb(w_n377_49[0]),.dout(n2509),.clk(gclk));
	jor g2247(.dina(n2509),.dinb(n2508),.dout(n2510),.clk(gclk));
	jand g2248(.dina(w_n1654_1[0]),.dinb(w_n432_49[0]),.dout(n2511),.clk(gclk));
	jand g2249(.dina(w_n1679_1[0]),.dinb(w_n323_49[0]),.dout(n2512),.clk(gclk));
	jor g2250(.dina(n2512),.dinb(n2511),.dout(n2513),.clk(gclk));
	jor g2251(.dina(n2513),.dinb(n2510),.dout(n2514),.clk(gclk));
	jand g2252(.dina(w_n2514_0[1]),.dinb(w_shift6_56[1]),.dout(n2515),.clk(gclk));
	jor g2253(.dina(n2515),.dinb(n2507),.dout(result21),.clk(gclk));
	jand g2254(.dina(w_n1708_1[0]),.dinb(w_n323_48[2]),.dout(n2517),.clk(gclk));
	jand g2255(.dina(w_n1716_1[0]),.dinb(w_n377_48[2]),.dout(n2518),.clk(gclk));
	jor g2256(.dina(n2518),.dinb(n2517),.dout(n2519),.clk(gclk));
	jand g2257(.dina(w_n1699_1[0]),.dinb(w_n432_48[2]),.dout(n2520),.clk(gclk));
	jand g2258(.dina(w_n1735_1[0]),.dinb(w_n485_48[2]),.dout(n2521),.clk(gclk));
	jor g2259(.dina(n2521),.dinb(n2520),.dout(n2522),.clk(gclk));
	jor g2260(.dina(n2522),.dinb(n2519),.dout(n2523),.clk(gclk));
	jand g2261(.dina(w_n2523_0[1]),.dinb(w_n263_56[0]),.dout(n2524),.clk(gclk));
	jand g2262(.dina(w_n1691_1[0]),.dinb(w_n485_48[1]),.dout(n2525),.clk(gclk));
	jand g2263(.dina(w_n1744_1[0]),.dinb(w_n377_48[1]),.dout(n2526),.clk(gclk));
	jor g2264(.dina(n2526),.dinb(n2525),.dout(n2527),.clk(gclk));
	jand g2265(.dina(w_n1727_1[0]),.dinb(w_n432_48[1]),.dout(n2528),.clk(gclk));
	jand g2266(.dina(w_n1752_1[0]),.dinb(w_n323_48[1]),.dout(n2529),.clk(gclk));
	jor g2267(.dina(n2529),.dinb(n2528),.dout(n2530),.clk(gclk));
	jor g2268(.dina(n2530),.dinb(n2527),.dout(n2531),.clk(gclk));
	jand g2269(.dina(w_n2531_0[1]),.dinb(w_shift6_56[0]),.dout(n2532),.clk(gclk));
	jor g2270(.dina(n2532),.dinb(n2524),.dout(result22),.clk(gclk));
	jand g2271(.dina(w_n1781_1[0]),.dinb(w_n323_48[0]),.dout(n2534),.clk(gclk));
	jand g2272(.dina(w_n1772_1[0]),.dinb(w_n432_48[0]),.dout(n2535),.clk(gclk));
	jor g2273(.dina(n2535),.dinb(n2534),.dout(n2536),.clk(gclk));
	jand g2274(.dina(w_n1808_1[0]),.dinb(w_n485_48[0]),.dout(n2537),.clk(gclk));
	jand g2275(.dina(w_n1789_1[0]),.dinb(w_n377_48[0]),.dout(n2538),.clk(gclk));
	jor g2276(.dina(n2538),.dinb(n2537),.dout(n2539),.clk(gclk));
	jor g2277(.dina(n2539),.dinb(n2536),.dout(n2540),.clk(gclk));
	jand g2278(.dina(w_n2540_0[1]),.dinb(w_n263_55[2]),.dout(n2541),.clk(gclk));
	jand g2279(.dina(w_n1800_1[0]),.dinb(w_n432_47[2]),.dout(n2542),.clk(gclk));
	jand g2280(.dina(w_n1764_1[0]),.dinb(w_n485_47[2]),.dout(n2543),.clk(gclk));
	jor g2281(.dina(n2543),.dinb(n2542),.dout(n2544),.clk(gclk));
	jand g2282(.dina(w_n1817_1[0]),.dinb(w_n377_47[2]),.dout(n2545),.clk(gclk));
	jand g2283(.dina(w_n1825_1[0]),.dinb(w_n323_47[2]),.dout(n2546),.clk(gclk));
	jor g2284(.dina(n2546),.dinb(n2545),.dout(n2547),.clk(gclk));
	jor g2285(.dina(n2547),.dinb(n2544),.dout(n2548),.clk(gclk));
	jand g2286(.dina(w_n2548_0[1]),.dinb(w_shift6_55[2]),.dout(n2549),.clk(gclk));
	jor g2287(.dina(n2549),.dinb(n2541),.dout(result23),.clk(gclk));
	jand g2288(.dina(w_n1854_1[0]),.dinb(w_n323_47[1]),.dout(n2551),.clk(gclk));
	jand g2289(.dina(w_n1845_1[0]),.dinb(w_n432_47[1]),.dout(n2552),.clk(gclk));
	jor g2290(.dina(n2552),.dinb(n2551),.dout(n2553),.clk(gclk));
	jand g2291(.dina(w_n1881_1[0]),.dinb(w_n485_47[1]),.dout(n2554),.clk(gclk));
	jand g2292(.dina(w_n1862_1[0]),.dinb(w_n377_47[1]),.dout(n2555),.clk(gclk));
	jor g2293(.dina(n2555),.dinb(n2554),.dout(n2556),.clk(gclk));
	jor g2294(.dina(n2556),.dinb(n2553),.dout(n2557),.clk(gclk));
	jand g2295(.dina(w_n2557_0[1]),.dinb(w_n263_55[1]),.dout(n2558),.clk(gclk));
	jand g2296(.dina(w_n1873_1[0]),.dinb(w_n432_47[0]),.dout(n2559),.clk(gclk));
	jand g2297(.dina(w_n1837_1[0]),.dinb(w_n485_47[0]),.dout(n2560),.clk(gclk));
	jor g2298(.dina(n2560),.dinb(n2559),.dout(n2561),.clk(gclk));
	jand g2299(.dina(w_n1890_1[0]),.dinb(w_n377_47[0]),.dout(n2562),.clk(gclk));
	jand g2300(.dina(w_n1898_1[0]),.dinb(w_n323_47[0]),.dout(n2563),.clk(gclk));
	jor g2301(.dina(n2563),.dinb(n2562),.dout(n2564),.clk(gclk));
	jor g2302(.dina(n2564),.dinb(n2561),.dout(n2565),.clk(gclk));
	jand g2303(.dina(w_n2565_0[1]),.dinb(w_shift6_55[1]),.dout(n2566),.clk(gclk));
	jor g2304(.dina(n2566),.dinb(n2558),.dout(result24),.clk(gclk));
	jand g2305(.dina(w_n1927_1[0]),.dinb(w_n323_46[2]),.dout(n2568),.clk(gclk));
	jand g2306(.dina(w_n1918_1[0]),.dinb(w_n432_46[2]),.dout(n2569),.clk(gclk));
	jor g2307(.dina(n2569),.dinb(n2568),.dout(n2570),.clk(gclk));
	jand g2308(.dina(w_n1954_1[0]),.dinb(w_n485_46[2]),.dout(n2571),.clk(gclk));
	jand g2309(.dina(w_n1935_1[0]),.dinb(w_n377_46[2]),.dout(n2572),.clk(gclk));
	jor g2310(.dina(n2572),.dinb(n2571),.dout(n2573),.clk(gclk));
	jor g2311(.dina(n2573),.dinb(n2570),.dout(n2574),.clk(gclk));
	jand g2312(.dina(w_n2574_0[1]),.dinb(w_n263_55[0]),.dout(n2575),.clk(gclk));
	jand g2313(.dina(w_n1946_1[0]),.dinb(w_n432_46[1]),.dout(n2576),.clk(gclk));
	jand g2314(.dina(w_n1910_1[0]),.dinb(w_n485_46[1]),.dout(n2577),.clk(gclk));
	jor g2315(.dina(n2577),.dinb(n2576),.dout(n2578),.clk(gclk));
	jand g2316(.dina(w_n1963_1[0]),.dinb(w_n377_46[1]),.dout(n2579),.clk(gclk));
	jand g2317(.dina(w_n1971_1[0]),.dinb(w_n323_46[1]),.dout(n2580),.clk(gclk));
	jor g2318(.dina(n2580),.dinb(n2579),.dout(n2581),.clk(gclk));
	jor g2319(.dina(n2581),.dinb(n2578),.dout(n2582),.clk(gclk));
	jand g2320(.dina(w_n2582_0[1]),.dinb(w_shift6_55[0]),.dout(n2583),.clk(gclk));
	jor g2321(.dina(n2583),.dinb(n2575),.dout(result25),.clk(gclk));
	jand g2322(.dina(w_n2000_1[0]),.dinb(w_n323_46[0]),.dout(n2585),.clk(gclk));
	jand g2323(.dina(w_n2008_1[0]),.dinb(w_n377_46[0]),.dout(n2586),.clk(gclk));
	jor g2324(.dina(n2586),.dinb(n2585),.dout(n2587),.clk(gclk));
	jand g2325(.dina(w_n1991_1[0]),.dinb(w_n432_46[0]),.dout(n2588),.clk(gclk));
	jand g2326(.dina(w_n2027_1[0]),.dinb(w_n485_46[0]),.dout(n2589),.clk(gclk));
	jor g2327(.dina(n2589),.dinb(n2588),.dout(n2590),.clk(gclk));
	jor g2328(.dina(n2590),.dinb(n2587),.dout(n2591),.clk(gclk));
	jand g2329(.dina(w_n2591_0[1]),.dinb(w_n263_54[2]),.dout(n2592),.clk(gclk));
	jand g2330(.dina(w_n2019_1[0]),.dinb(w_n432_45[2]),.dout(n2593),.clk(gclk));
	jand g2331(.dina(w_n1983_1[0]),.dinb(w_n485_45[2]),.dout(n2594),.clk(gclk));
	jor g2332(.dina(n2594),.dinb(n2593),.dout(n2595),.clk(gclk));
	jand g2333(.dina(w_n2036_1[0]),.dinb(w_n377_45[2]),.dout(n2596),.clk(gclk));
	jand g2334(.dina(w_n2044_1[0]),.dinb(w_n323_45[2]),.dout(n2597),.clk(gclk));
	jor g2335(.dina(n2597),.dinb(n2596),.dout(n2598),.clk(gclk));
	jor g2336(.dina(n2598),.dinb(n2595),.dout(n2599),.clk(gclk));
	jand g2337(.dina(w_n2599_0[1]),.dinb(w_shift6_54[2]),.dout(n2600),.clk(gclk));
	jor g2338(.dina(n2600),.dinb(n2592),.dout(result26),.clk(gclk));
	jand g2339(.dina(w_n2073_1[0]),.dinb(w_n323_45[1]),.dout(n2602),.clk(gclk));
	jand g2340(.dina(w_n2081_1[0]),.dinb(w_n377_45[1]),.dout(n2603),.clk(gclk));
	jor g2341(.dina(n2603),.dinb(n2602),.dout(n2604),.clk(gclk));
	jand g2342(.dina(w_n2064_1[0]),.dinb(w_n432_45[1]),.dout(n2605),.clk(gclk));
	jand g2343(.dina(w_n2100_1[0]),.dinb(w_n485_45[1]),.dout(n2606),.clk(gclk));
	jor g2344(.dina(n2606),.dinb(n2605),.dout(n2607),.clk(gclk));
	jor g2345(.dina(n2607),.dinb(n2604),.dout(n2608),.clk(gclk));
	jand g2346(.dina(w_n2608_0[1]),.dinb(w_n263_54[1]),.dout(n2609),.clk(gclk));
	jand g2347(.dina(w_n2092_1[0]),.dinb(w_n432_45[0]),.dout(n2610),.clk(gclk));
	jand g2348(.dina(w_n2056_1[0]),.dinb(w_n485_45[0]),.dout(n2611),.clk(gclk));
	jor g2349(.dina(n2611),.dinb(n2610),.dout(n2612),.clk(gclk));
	jand g2350(.dina(w_n2109_1[0]),.dinb(w_n377_45[0]),.dout(n2613),.clk(gclk));
	jand g2351(.dina(w_n2117_1[0]),.dinb(w_n323_45[0]),.dout(n2614),.clk(gclk));
	jor g2352(.dina(n2614),.dinb(n2613),.dout(n2615),.clk(gclk));
	jor g2353(.dina(n2615),.dinb(n2612),.dout(n2616),.clk(gclk));
	jand g2354(.dina(w_n2616_0[1]),.dinb(w_shift6_54[1]),.dout(n2617),.clk(gclk));
	jor g2355(.dina(n2617),.dinb(n2609),.dout(result27),.clk(gclk));
	jand g2356(.dina(w_n2146_1[0]),.dinb(w_n323_44[2]),.dout(n2619),.clk(gclk));
	jand g2357(.dina(w_n2154_1[0]),.dinb(w_n377_44[2]),.dout(n2620),.clk(gclk));
	jor g2358(.dina(n2620),.dinb(n2619),.dout(n2621),.clk(gclk));
	jand g2359(.dina(w_n2137_1[0]),.dinb(w_n432_44[2]),.dout(n2622),.clk(gclk));
	jand g2360(.dina(w_n2173_1[0]),.dinb(w_n485_44[2]),.dout(n2623),.clk(gclk));
	jor g2361(.dina(n2623),.dinb(n2622),.dout(n2624),.clk(gclk));
	jor g2362(.dina(n2624),.dinb(n2621),.dout(n2625),.clk(gclk));
	jand g2363(.dina(w_n2625_0[1]),.dinb(w_n263_54[0]),.dout(n2626),.clk(gclk));
	jand g2364(.dina(w_n2165_1[0]),.dinb(w_n432_44[1]),.dout(n2627),.clk(gclk));
	jand g2365(.dina(w_n2129_1[0]),.dinb(w_n485_44[1]),.dout(n2628),.clk(gclk));
	jor g2366(.dina(n2628),.dinb(n2627),.dout(n2629),.clk(gclk));
	jand g2367(.dina(w_n2182_1[0]),.dinb(w_n377_44[1]),.dout(n2630),.clk(gclk));
	jand g2368(.dina(w_n2190_1[0]),.dinb(w_n323_44[1]),.dout(n2631),.clk(gclk));
	jor g2369(.dina(n2631),.dinb(n2630),.dout(n2632),.clk(gclk));
	jor g2370(.dina(n2632),.dinb(n2629),.dout(n2633),.clk(gclk));
	jand g2371(.dina(w_n2633_0[1]),.dinb(w_shift6_54[0]),.dout(n2634),.clk(gclk));
	jor g2372(.dina(n2634),.dinb(n2626),.dout(result28),.clk(gclk));
	jand g2373(.dina(w_n2219_1[0]),.dinb(w_n323_44[0]),.dout(n2636),.clk(gclk));
	jand g2374(.dina(w_n2227_1[0]),.dinb(w_n377_44[0]),.dout(n2637),.clk(gclk));
	jor g2375(.dina(n2637),.dinb(n2636),.dout(n2638),.clk(gclk));
	jand g2376(.dina(w_n2210_1[0]),.dinb(w_n432_44[0]),.dout(n2639),.clk(gclk));
	jand g2377(.dina(w_n2246_1[0]),.dinb(w_n485_44[0]),.dout(n2640),.clk(gclk));
	jor g2378(.dina(n2640),.dinb(n2639),.dout(n2641),.clk(gclk));
	jor g2379(.dina(n2641),.dinb(n2638),.dout(n2642),.clk(gclk));
	jand g2380(.dina(w_n2642_0[1]),.dinb(w_n263_53[2]),.dout(n2643),.clk(gclk));
	jand g2381(.dina(w_n2238_1[0]),.dinb(w_n432_43[2]),.dout(n2644),.clk(gclk));
	jand g2382(.dina(w_n2202_1[0]),.dinb(w_n485_43[2]),.dout(n2645),.clk(gclk));
	jor g2383(.dina(n2645),.dinb(n2644),.dout(n2646),.clk(gclk));
	jand g2384(.dina(w_n2255_1[0]),.dinb(w_n377_43[2]),.dout(n2647),.clk(gclk));
	jand g2385(.dina(w_n2263_1[0]),.dinb(w_n323_43[2]),.dout(n2648),.clk(gclk));
	jor g2386(.dina(n2648),.dinb(n2647),.dout(n2649),.clk(gclk));
	jor g2387(.dina(n2649),.dinb(n2646),.dout(n2650),.clk(gclk));
	jand g2388(.dina(w_n2650_0[1]),.dinb(w_shift6_53[2]),.dout(n2651),.clk(gclk));
	jor g2389(.dina(n2651),.dinb(n2643),.dout(result29),.clk(gclk));
	jand g2390(.dina(w_n2292_1[0]),.dinb(w_n323_43[1]),.dout(n2653),.clk(gclk));
	jand g2391(.dina(w_n2300_1[0]),.dinb(w_n377_43[1]),.dout(n2654),.clk(gclk));
	jor g2392(.dina(n2654),.dinb(n2653),.dout(n2655),.clk(gclk));
	jand g2393(.dina(w_n2283_1[0]),.dinb(w_n432_43[1]),.dout(n2656),.clk(gclk));
	jand g2394(.dina(w_n2319_1[0]),.dinb(w_n485_43[1]),.dout(n2657),.clk(gclk));
	jor g2395(.dina(n2657),.dinb(n2656),.dout(n2658),.clk(gclk));
	jor g2396(.dina(n2658),.dinb(n2655),.dout(n2659),.clk(gclk));
	jand g2397(.dina(w_n2659_0[1]),.dinb(w_n263_53[1]),.dout(n2660),.clk(gclk));
	jand g2398(.dina(w_n2311_1[0]),.dinb(w_n432_43[0]),.dout(n2661),.clk(gclk));
	jand g2399(.dina(w_n2275_1[0]),.dinb(w_n485_43[0]),.dout(n2662),.clk(gclk));
	jor g2400(.dina(n2662),.dinb(n2661),.dout(n2663),.clk(gclk));
	jand g2401(.dina(w_n2328_1[0]),.dinb(w_n377_43[0]),.dout(n2664),.clk(gclk));
	jand g2402(.dina(w_n2336_1[0]),.dinb(w_n323_43[0]),.dout(n2665),.clk(gclk));
	jor g2403(.dina(n2665),.dinb(n2664),.dout(n2666),.clk(gclk));
	jor g2404(.dina(n2666),.dinb(n2663),.dout(n2667),.clk(gclk));
	jand g2405(.dina(w_n2667_0[1]),.dinb(w_shift6_53[1]),.dout(n2668),.clk(gclk));
	jor g2406(.dina(n2668),.dinb(n2660),.dout(result30),.clk(gclk));
	jand g2407(.dina(w_n2365_1[0]),.dinb(w_n323_42[2]),.dout(n2670),.clk(gclk));
	jand g2408(.dina(w_n2373_1[0]),.dinb(w_n377_42[2]),.dout(n2671),.clk(gclk));
	jor g2409(.dina(n2671),.dinb(n2670),.dout(n2672),.clk(gclk));
	jand g2410(.dina(w_n2356_1[0]),.dinb(w_n432_42[2]),.dout(n2673),.clk(gclk));
	jand g2411(.dina(w_n2392_1[0]),.dinb(w_n485_42[2]),.dout(n2674),.clk(gclk));
	jor g2412(.dina(n2674),.dinb(n2673),.dout(n2675),.clk(gclk));
	jor g2413(.dina(n2675),.dinb(n2672),.dout(n2676),.clk(gclk));
	jand g2414(.dina(w_n2676_0[1]),.dinb(w_n263_53[0]),.dout(n2677),.clk(gclk));
	jand g2415(.dina(w_n2384_1[0]),.dinb(w_n432_42[1]),.dout(n2678),.clk(gclk));
	jand g2416(.dina(w_n2348_1[0]),.dinb(w_n485_42[1]),.dout(n2679),.clk(gclk));
	jor g2417(.dina(n2679),.dinb(n2678),.dout(n2680),.clk(gclk));
	jand g2418(.dina(w_n2401_1[0]),.dinb(w_n377_42[1]),.dout(n2681),.clk(gclk));
	jand g2419(.dina(w_n2409_1[0]),.dinb(w_n323_42[1]),.dout(n2682),.clk(gclk));
	jor g2420(.dina(n2682),.dinb(n2681),.dout(n2683),.clk(gclk));
	jor g2421(.dina(n2683),.dinb(n2680),.dout(n2684),.clk(gclk));
	jand g2422(.dina(w_n2684_0[1]),.dinb(w_shift6_53[0]),.dout(n2685),.clk(gclk));
	jor g2423(.dina(n2685),.dinb(n2677),.dout(result31),.clk(gclk));
	jand g2424(.dina(w_n375_0[2]),.dinb(w_n323_42[0]),.dout(n2687),.clk(gclk));
	jand g2425(.dina(w_n540_0[2]),.dinb(w_n377_42[0]),.dout(n2688),.clk(gclk));
	jor g2426(.dina(n2688),.dinb(n2687),.dout(n2689),.clk(gclk));
	jand g2427(.dina(w_n484_0[2]),.dinb(w_n432_42[0]),.dout(n2690),.clk(gclk));
	jand g2428(.dina(w_n643_0[2]),.dinb(w_n485_42[0]),.dout(n2691),.clk(gclk));
	jor g2429(.dina(n2691),.dinb(n2690),.dout(n2692),.clk(gclk));
	jor g2430(.dina(n2692),.dinb(n2689),.dout(n2693),.clk(gclk));
	jand g2431(.dina(w_n2693_0[1]),.dinb(w_n263_52[2]),.dout(n2694),.clk(gclk));
	jand g2432(.dina(w_n377_41[2]),.dinb(w_n322_0[2]),.dout(n2695),.clk(gclk));
	jand g2433(.dina(w_n590_0[2]),.dinb(w_n323_41[2]),.dout(n2696),.clk(gclk));
	jor g2434(.dina(n2696),.dinb(n2695),.dout(n2697),.clk(gclk));
	jand g2435(.dina(w_n485_41[2]),.dinb(w_n430_0[2]),.dout(n2698),.clk(gclk));
	jand g2436(.dina(w_n695_0[2]),.dinb(w_n432_41[2]),.dout(n2699),.clk(gclk));
	jor g2437(.dina(n2699),.dinb(n2698),.dout(n2700),.clk(gclk));
	jor g2438(.dina(n2700),.dinb(n2697),.dout(n2701),.clk(gclk));
	jand g2439(.dina(w_n2701_0[1]),.dinb(w_shift6_52[2]),.dout(n2702),.clk(gclk));
	jor g2440(.dina(n2702),.dinb(n2694),.dout(result32),.clk(gclk));
	jand g2441(.dina(w_n787_0[2]),.dinb(w_n323_41[1]),.dout(n2704),.clk(gclk));
	jand g2442(.dina(w_n1012_0[2]),.dinb(w_n377_41[1]),.dout(n2705),.clk(gclk));
	jor g2443(.dina(n2705),.dinb(n2704),.dout(n2706),.clk(gclk));
	jand g2444(.dina(w_n876_0[2]),.dinb(w_n432_41[1]),.dout(n2707),.clk(gclk));
	jand g2445(.dina(w_n967_0[2]),.dinb(w_n485_41[1]),.dout(n2708),.clk(gclk));
	jor g2446(.dina(n2708),.dinb(n2707),.dout(n2709),.clk(gclk));
	jor g2447(.dina(n2709),.dinb(n2706),.dout(n2710),.clk(gclk));
	jand g2448(.dina(w_n2710_0[1]),.dinb(w_n263_52[1]),.dout(n2711),.clk(gclk));
	jand g2449(.dina(w_n923_0[2]),.dinb(w_n432_41[0]),.dout(n2712),.clk(gclk));
	jand g2450(.dina(w_n832_0[2]),.dinb(w_n485_41[0]),.dout(n2713),.clk(gclk));
	jor g2451(.dina(n2713),.dinb(n2712),.dout(n2714),.clk(gclk));
	jand g2452(.dina(w_n743_0[2]),.dinb(w_n377_41[0]),.dout(n2715),.clk(gclk));
	jand g2453(.dina(w_n1060_0[2]),.dinb(w_n323_41[0]),.dout(n2716),.clk(gclk));
	jor g2454(.dina(n2716),.dinb(n2715),.dout(n2717),.clk(gclk));
	jor g2455(.dina(n2717),.dinb(n2714),.dout(n2718),.clk(gclk));
	jand g2456(.dina(w_n2718_0[1]),.dinb(w_shift6_52[1]),.dout(n2719),.clk(gclk));
	jor g2457(.dina(n2719),.dinb(n2711),.dout(result33),.clk(gclk));
	jand g2458(.dina(w_n1136_0[2]),.dinb(w_n323_40[2]),.dout(n2721),.clk(gclk));
	jand g2459(.dina(w_n1321_0[2]),.dinb(w_n377_40[2]),.dout(n2722),.clk(gclk));
	jor g2460(.dina(n2722),.dinb(n2721),.dout(n2723),.clk(gclk));
	jand g2461(.dina(w_n1209_0[2]),.dinb(w_n432_40[2]),.dout(n2724),.clk(gclk));
	jand g2462(.dina(w_n1284_0[2]),.dinb(w_n485_40[2]),.dout(n2725),.clk(gclk));
	jor g2463(.dina(n2725),.dinb(n2724),.dout(n2726),.clk(gclk));
	jor g2464(.dina(n2726),.dinb(n2723),.dout(n2727),.clk(gclk));
	jand g2465(.dina(w_n2727_0[1]),.dinb(w_n263_52[0]),.dout(n2728),.clk(gclk));
	jand g2466(.dina(w_n1248_0[2]),.dinb(w_n432_40[1]),.dout(n2729),.clk(gclk));
	jand g2467(.dina(w_n1173_0[2]),.dinb(w_n485_40[1]),.dout(n2730),.clk(gclk));
	jor g2468(.dina(n2730),.dinb(n2729),.dout(n2731),.clk(gclk));
	jand g2469(.dina(w_n1100_0[2]),.dinb(w_n377_40[1]),.dout(n2732),.clk(gclk));
	jand g2470(.dina(w_n1357_0[2]),.dinb(w_n323_40[1]),.dout(n2733),.clk(gclk));
	jor g2471(.dina(n2733),.dinb(n2732),.dout(n2734),.clk(gclk));
	jor g2472(.dina(n2734),.dinb(n2731),.dout(n2735),.clk(gclk));
	jand g2473(.dina(w_n2735_0[1]),.dinb(w_shift6_52[0]),.dout(n2736),.clk(gclk));
	jor g2474(.dina(n2736),.dinb(n2728),.dout(result34),.clk(gclk));
	jand g2475(.dina(w_n1381_0[2]),.dinb(w_n323_40[0]),.dout(n2738),.clk(gclk));
	jand g2476(.dina(w_n1533_0[2]),.dinb(w_n377_40[0]),.dout(n2739),.clk(gclk));
	jor g2477(.dina(n2739),.dinb(n2738),.dout(n2740),.clk(gclk));
	jand g2478(.dina(w_n1485_0[2]),.dinb(w_n485_40[0]),.dout(n2741),.clk(gclk));
	jand g2479(.dina(w_n1442_0[2]),.dinb(w_n432_40[0]),.dout(n2742),.clk(gclk));
	jor g2480(.dina(n2742),.dinb(n2741),.dout(n2743),.clk(gclk));
	jor g2481(.dina(n2743),.dinb(n2740),.dout(n2744),.clk(gclk));
	jand g2482(.dina(w_n2744_0[1]),.dinb(w_n263_51[2]),.dout(n2745),.clk(gclk));
	jand g2483(.dina(w_n1465_0[2]),.dinb(w_n432_39[2]),.dout(n2746),.clk(gclk));
	jand g2484(.dina(w_n1401_0[2]),.dinb(w_n377_39[2]),.dout(n2747),.clk(gclk));
	jor g2485(.dina(n2747),.dinb(n2746),.dout(n2748),.clk(gclk));
	jand g2486(.dina(w_n1422_0[2]),.dinb(w_n485_39[2]),.dout(n2749),.clk(gclk));
	jand g2487(.dina(w_n1513_0[2]),.dinb(w_n323_39[2]),.dout(n2750),.clk(gclk));
	jor g2488(.dina(n2750),.dinb(n2749),.dout(n2751),.clk(gclk));
	jor g2489(.dina(n2751),.dinb(n2748),.dout(n2752),.clk(gclk));
	jand g2490(.dina(w_n2752_0[1]),.dinb(w_shift6_51[2]),.dout(n2753),.clk(gclk));
	jor g2491(.dina(n2753),.dinb(n2745),.dout(result35),.clk(gclk));
	jand g2492(.dina(w_n1553_0[2]),.dinb(w_n323_39[1]),.dout(n2755),.clk(gclk));
	jand g2493(.dina(w_n1589_0[2]),.dinb(w_n377_39[1]),.dout(n2756),.clk(gclk));
	jor g2494(.dina(n2756),.dinb(n2755),.dout(n2757),.clk(gclk));
	jand g2495(.dina(w_n1570_0[2]),.dinb(w_n432_39[1]),.dout(n2758),.clk(gclk));
	jand g2496(.dina(w_n1606_0[2]),.dinb(w_n485_39[1]),.dout(n2759),.clk(gclk));
	jor g2497(.dina(n2759),.dinb(n2758),.dout(n2760),.clk(gclk));
	jor g2498(.dina(n2760),.dinb(n2757),.dout(n2761),.clk(gclk));
	jand g2499(.dina(w_n2761_0[1]),.dinb(w_n263_51[1]),.dout(n2762),.clk(gclk));
	jand g2500(.dina(w_n1545_0[2]),.dinb(w_n377_39[0]),.dout(n2763),.clk(gclk));
	jand g2501(.dina(w_n1581_0[2]),.dinb(w_n323_39[0]),.dout(n2764),.clk(gclk));
	jor g2502(.dina(n2764),.dinb(n2763),.dout(n2765),.clk(gclk));
	jand g2503(.dina(w_n1562_0[2]),.dinb(w_n485_39[0]),.dout(n2766),.clk(gclk));
	jand g2504(.dina(w_n1598_0[2]),.dinb(w_n432_39[0]),.dout(n2767),.clk(gclk));
	jor g2505(.dina(n2767),.dinb(n2766),.dout(n2768),.clk(gclk));
	jor g2506(.dina(n2768),.dinb(n2765),.dout(n2769),.clk(gclk));
	jand g2507(.dina(w_n2769_0[1]),.dinb(w_shift6_51[1]),.dout(n2770),.clk(gclk));
	jor g2508(.dina(n2770),.dinb(n2762),.dout(result36),.clk(gclk));
	jand g2509(.dina(w_n1626_0[2]),.dinb(w_n323_38[2]),.dout(n2772),.clk(gclk));
	jand g2510(.dina(w_n1662_0[2]),.dinb(w_n377_38[2]),.dout(n2773),.clk(gclk));
	jor g2511(.dina(n2773),.dinb(n2772),.dout(n2774),.clk(gclk));
	jand g2512(.dina(w_n1643_0[2]),.dinb(w_n432_38[2]),.dout(n2775),.clk(gclk));
	jand g2513(.dina(w_n1679_0[2]),.dinb(w_n485_38[2]),.dout(n2776),.clk(gclk));
	jor g2514(.dina(n2776),.dinb(n2775),.dout(n2777),.clk(gclk));
	jor g2515(.dina(n2777),.dinb(n2774),.dout(n2778),.clk(gclk));
	jand g2516(.dina(w_n2778_0[1]),.dinb(w_n263_51[0]),.dout(n2779),.clk(gclk));
	jand g2517(.dina(w_n1618_0[2]),.dinb(w_n377_38[1]),.dout(n2780),.clk(gclk));
	jand g2518(.dina(w_n1654_0[2]),.dinb(w_n323_38[1]),.dout(n2781),.clk(gclk));
	jor g2519(.dina(n2781),.dinb(n2780),.dout(n2782),.clk(gclk));
	jand g2520(.dina(w_n1635_0[2]),.dinb(w_n485_38[1]),.dout(n2783),.clk(gclk));
	jand g2521(.dina(w_n1671_0[2]),.dinb(w_n432_38[1]),.dout(n2784),.clk(gclk));
	jor g2522(.dina(n2784),.dinb(n2783),.dout(n2785),.clk(gclk));
	jor g2523(.dina(n2785),.dinb(n2782),.dout(n2786),.clk(gclk));
	jand g2524(.dina(w_n2786_0[1]),.dinb(w_shift6_51[0]),.dout(n2787),.clk(gclk));
	jor g2525(.dina(n2787),.dinb(n2779),.dout(result37),.clk(gclk));
	jand g2526(.dina(w_n1699_0[2]),.dinb(w_n323_38[0]),.dout(n2789),.clk(gclk));
	jand g2527(.dina(w_n1735_0[2]),.dinb(w_n377_38[0]),.dout(n2790),.clk(gclk));
	jor g2528(.dina(n2790),.dinb(n2789),.dout(n2791),.clk(gclk));
	jand g2529(.dina(w_n1716_0[2]),.dinb(w_n432_38[0]),.dout(n2792),.clk(gclk));
	jand g2530(.dina(w_n1752_0[2]),.dinb(w_n485_38[0]),.dout(n2793),.clk(gclk));
	jor g2531(.dina(n2793),.dinb(n2792),.dout(n2794),.clk(gclk));
	jor g2532(.dina(n2794),.dinb(n2791),.dout(n2795),.clk(gclk));
	jand g2533(.dina(w_n2795_0[1]),.dinb(w_n263_50[2]),.dout(n2796),.clk(gclk));
	jand g2534(.dina(w_n1691_0[2]),.dinb(w_n377_37[2]),.dout(n2797),.clk(gclk));
	jand g2535(.dina(w_n1727_0[2]),.dinb(w_n323_37[2]),.dout(n2798),.clk(gclk));
	jor g2536(.dina(n2798),.dinb(n2797),.dout(n2799),.clk(gclk));
	jand g2537(.dina(w_n1708_0[2]),.dinb(w_n485_37[2]),.dout(n2800),.clk(gclk));
	jand g2538(.dina(w_n1744_0[2]),.dinb(w_n432_37[2]),.dout(n2801),.clk(gclk));
	jor g2539(.dina(n2801),.dinb(n2800),.dout(n2802),.clk(gclk));
	jor g2540(.dina(n2802),.dinb(n2799),.dout(n2803),.clk(gclk));
	jand g2541(.dina(w_n2803_0[1]),.dinb(w_shift6_50[2]),.dout(n2804),.clk(gclk));
	jor g2542(.dina(n2804),.dinb(n2796),.dout(result38),.clk(gclk));
	jand g2543(.dina(w_n1808_0[2]),.dinb(w_n377_37[1]),.dout(n2806),.clk(gclk));
	jand g2544(.dina(w_n1772_0[2]),.dinb(w_n323_37[1]),.dout(n2807),.clk(gclk));
	jor g2545(.dina(n2807),.dinb(n2806),.dout(n2808),.clk(gclk));
	jand g2546(.dina(w_n1825_0[2]),.dinb(w_n485_37[1]),.dout(n2809),.clk(gclk));
	jand g2547(.dina(w_n1789_0[2]),.dinb(w_n432_37[1]),.dout(n2810),.clk(gclk));
	jor g2548(.dina(n2810),.dinb(n2809),.dout(n2811),.clk(gclk));
	jor g2549(.dina(n2811),.dinb(n2808),.dout(n2812),.clk(gclk));
	jand g2550(.dina(w_n2812_0[1]),.dinb(w_n263_50[1]),.dout(n2813),.clk(gclk));
	jand g2551(.dina(w_n1800_0[2]),.dinb(w_n323_37[0]),.dout(n2814),.clk(gclk));
	jand g2552(.dina(w_n1764_0[2]),.dinb(w_n377_37[0]),.dout(n2815),.clk(gclk));
	jor g2553(.dina(n2815),.dinb(n2814),.dout(n2816),.clk(gclk));
	jand g2554(.dina(w_n1817_0[2]),.dinb(w_n432_37[0]),.dout(n2817),.clk(gclk));
	jand g2555(.dina(w_n1781_0[2]),.dinb(w_n485_37[0]),.dout(n2818),.clk(gclk));
	jor g2556(.dina(n2818),.dinb(n2817),.dout(n2819),.clk(gclk));
	jor g2557(.dina(n2819),.dinb(n2816),.dout(n2820),.clk(gclk));
	jand g2558(.dina(w_n2820_0[1]),.dinb(w_shift6_50[1]),.dout(n2821),.clk(gclk));
	jor g2559(.dina(n2821),.dinb(n2813),.dout(result39),.clk(gclk));
	jand g2560(.dina(w_n1881_0[2]),.dinb(w_n377_36[2]),.dout(n2823),.clk(gclk));
	jand g2561(.dina(w_n1845_0[2]),.dinb(w_n323_36[2]),.dout(n2824),.clk(gclk));
	jor g2562(.dina(n2824),.dinb(n2823),.dout(n2825),.clk(gclk));
	jand g2563(.dina(w_n1898_0[2]),.dinb(w_n485_36[2]),.dout(n2826),.clk(gclk));
	jand g2564(.dina(w_n1862_0[2]),.dinb(w_n432_36[2]),.dout(n2827),.clk(gclk));
	jor g2565(.dina(n2827),.dinb(n2826),.dout(n2828),.clk(gclk));
	jor g2566(.dina(n2828),.dinb(n2825),.dout(n2829),.clk(gclk));
	jand g2567(.dina(w_n2829_0[1]),.dinb(w_n263_50[0]),.dout(n2830),.clk(gclk));
	jand g2568(.dina(w_n1873_0[2]),.dinb(w_n323_36[1]),.dout(n2831),.clk(gclk));
	jand g2569(.dina(w_n1837_0[2]),.dinb(w_n377_36[1]),.dout(n2832),.clk(gclk));
	jor g2570(.dina(n2832),.dinb(n2831),.dout(n2833),.clk(gclk));
	jand g2571(.dina(w_n1890_0[2]),.dinb(w_n432_36[1]),.dout(n2834),.clk(gclk));
	jand g2572(.dina(w_n1854_0[2]),.dinb(w_n485_36[1]),.dout(n2835),.clk(gclk));
	jor g2573(.dina(n2835),.dinb(n2834),.dout(n2836),.clk(gclk));
	jor g2574(.dina(n2836),.dinb(n2833),.dout(n2837),.clk(gclk));
	jand g2575(.dina(w_n2837_0[1]),.dinb(w_shift6_50[0]),.dout(n2838),.clk(gclk));
	jor g2576(.dina(n2838),.dinb(n2830),.dout(result40),.clk(gclk));
	jand g2577(.dina(w_n1954_0[2]),.dinb(w_n377_36[0]),.dout(n2840),.clk(gclk));
	jand g2578(.dina(w_n1918_0[2]),.dinb(w_n323_36[0]),.dout(n2841),.clk(gclk));
	jor g2579(.dina(n2841),.dinb(n2840),.dout(n2842),.clk(gclk));
	jand g2580(.dina(w_n1971_0[2]),.dinb(w_n485_36[0]),.dout(n2843),.clk(gclk));
	jand g2581(.dina(w_n1935_0[2]),.dinb(w_n432_36[0]),.dout(n2844),.clk(gclk));
	jor g2582(.dina(n2844),.dinb(n2843),.dout(n2845),.clk(gclk));
	jor g2583(.dina(n2845),.dinb(n2842),.dout(n2846),.clk(gclk));
	jand g2584(.dina(w_n2846_0[1]),.dinb(w_n263_49[2]),.dout(n2847),.clk(gclk));
	jand g2585(.dina(w_n1946_0[2]),.dinb(w_n323_35[2]),.dout(n2848),.clk(gclk));
	jand g2586(.dina(w_n1910_0[2]),.dinb(w_n377_35[2]),.dout(n2849),.clk(gclk));
	jor g2587(.dina(n2849),.dinb(n2848),.dout(n2850),.clk(gclk));
	jand g2588(.dina(w_n1963_0[2]),.dinb(w_n432_35[2]),.dout(n2851),.clk(gclk));
	jand g2589(.dina(w_n1927_0[2]),.dinb(w_n485_35[2]),.dout(n2852),.clk(gclk));
	jor g2590(.dina(n2852),.dinb(n2851),.dout(n2853),.clk(gclk));
	jor g2591(.dina(n2853),.dinb(n2850),.dout(n2854),.clk(gclk));
	jand g2592(.dina(w_n2854_0[1]),.dinb(w_shift6_49[2]),.dout(n2855),.clk(gclk));
	jor g2593(.dina(n2855),.dinb(n2847),.dout(result41),.clk(gclk));
	jand g2594(.dina(w_n1991_0[2]),.dinb(w_n323_35[1]),.dout(n2857),.clk(gclk));
	jand g2595(.dina(w_n2027_0[2]),.dinb(w_n377_35[1]),.dout(n2858),.clk(gclk));
	jor g2596(.dina(n2858),.dinb(n2857),.dout(n2859),.clk(gclk));
	jand g2597(.dina(w_n2008_0[2]),.dinb(w_n432_35[1]),.dout(n2860),.clk(gclk));
	jand g2598(.dina(w_n2044_0[2]),.dinb(w_n485_35[1]),.dout(n2861),.clk(gclk));
	jor g2599(.dina(n2861),.dinb(n2860),.dout(n2862),.clk(gclk));
	jor g2600(.dina(n2862),.dinb(n2859),.dout(n2863),.clk(gclk));
	jand g2601(.dina(w_n2863_0[1]),.dinb(w_n263_49[1]),.dout(n2864),.clk(gclk));
	jand g2602(.dina(w_n2019_0[2]),.dinb(w_n323_35[0]),.dout(n2865),.clk(gclk));
	jand g2603(.dina(w_n1983_0[2]),.dinb(w_n377_35[0]),.dout(n2866),.clk(gclk));
	jor g2604(.dina(n2866),.dinb(n2865),.dout(n2867),.clk(gclk));
	jand g2605(.dina(w_n2036_0[2]),.dinb(w_n432_35[0]),.dout(n2868),.clk(gclk));
	jand g2606(.dina(w_n2000_0[2]),.dinb(w_n485_35[0]),.dout(n2869),.clk(gclk));
	jor g2607(.dina(n2869),.dinb(n2868),.dout(n2870),.clk(gclk));
	jor g2608(.dina(n2870),.dinb(n2867),.dout(n2871),.clk(gclk));
	jand g2609(.dina(w_n2871_0[1]),.dinb(w_shift6_49[1]),.dout(n2872),.clk(gclk));
	jor g2610(.dina(n2872),.dinb(n2864),.dout(result42),.clk(gclk));
	jand g2611(.dina(w_n2064_0[2]),.dinb(w_n323_34[2]),.dout(n2874),.clk(gclk));
	jand g2612(.dina(w_n2100_0[2]),.dinb(w_n377_34[2]),.dout(n2875),.clk(gclk));
	jor g2613(.dina(n2875),.dinb(n2874),.dout(n2876),.clk(gclk));
	jand g2614(.dina(w_n2081_0[2]),.dinb(w_n432_34[2]),.dout(n2877),.clk(gclk));
	jand g2615(.dina(w_n2117_0[2]),.dinb(w_n485_34[2]),.dout(n2878),.clk(gclk));
	jor g2616(.dina(n2878),.dinb(n2877),.dout(n2879),.clk(gclk));
	jor g2617(.dina(n2879),.dinb(n2876),.dout(n2880),.clk(gclk));
	jand g2618(.dina(w_n2880_0[1]),.dinb(w_n263_49[0]),.dout(n2881),.clk(gclk));
	jand g2619(.dina(w_n2092_0[2]),.dinb(w_n323_34[1]),.dout(n2882),.clk(gclk));
	jand g2620(.dina(w_n2056_0[2]),.dinb(w_n377_34[1]),.dout(n2883),.clk(gclk));
	jor g2621(.dina(n2883),.dinb(n2882),.dout(n2884),.clk(gclk));
	jand g2622(.dina(w_n2109_0[2]),.dinb(w_n432_34[1]),.dout(n2885),.clk(gclk));
	jand g2623(.dina(w_n2073_0[2]),.dinb(w_n485_34[1]),.dout(n2886),.clk(gclk));
	jor g2624(.dina(n2886),.dinb(n2885),.dout(n2887),.clk(gclk));
	jor g2625(.dina(n2887),.dinb(n2884),.dout(n2888),.clk(gclk));
	jand g2626(.dina(w_n2888_0[1]),.dinb(w_shift6_49[0]),.dout(n2889),.clk(gclk));
	jor g2627(.dina(n2889),.dinb(n2881),.dout(result43),.clk(gclk));
	jand g2628(.dina(w_n2137_0[2]),.dinb(w_n323_34[0]),.dout(n2891),.clk(gclk));
	jand g2629(.dina(w_n2173_0[2]),.dinb(w_n377_34[0]),.dout(n2892),.clk(gclk));
	jor g2630(.dina(n2892),.dinb(n2891),.dout(n2893),.clk(gclk));
	jand g2631(.dina(w_n2154_0[2]),.dinb(w_n432_34[0]),.dout(n2894),.clk(gclk));
	jand g2632(.dina(w_n2190_0[2]),.dinb(w_n485_34[0]),.dout(n2895),.clk(gclk));
	jor g2633(.dina(n2895),.dinb(n2894),.dout(n2896),.clk(gclk));
	jor g2634(.dina(n2896),.dinb(n2893),.dout(n2897),.clk(gclk));
	jand g2635(.dina(w_n2897_0[1]),.dinb(w_n263_48[2]),.dout(n2898),.clk(gclk));
	jand g2636(.dina(w_n2165_0[2]),.dinb(w_n323_33[2]),.dout(n2899),.clk(gclk));
	jand g2637(.dina(w_n2129_0[2]),.dinb(w_n377_33[2]),.dout(n2900),.clk(gclk));
	jor g2638(.dina(n2900),.dinb(n2899),.dout(n2901),.clk(gclk));
	jand g2639(.dina(w_n2182_0[2]),.dinb(w_n432_33[2]),.dout(n2902),.clk(gclk));
	jand g2640(.dina(w_n2146_0[2]),.dinb(w_n485_33[2]),.dout(n2903),.clk(gclk));
	jor g2641(.dina(n2903),.dinb(n2902),.dout(n2904),.clk(gclk));
	jor g2642(.dina(n2904),.dinb(n2901),.dout(n2905),.clk(gclk));
	jand g2643(.dina(w_n2905_0[1]),.dinb(w_shift6_48[2]),.dout(n2906),.clk(gclk));
	jor g2644(.dina(n2906),.dinb(n2898),.dout(result44),.clk(gclk));
	jand g2645(.dina(w_n2210_0[2]),.dinb(w_n323_33[1]),.dout(n2908),.clk(gclk));
	jand g2646(.dina(w_n2246_0[2]),.dinb(w_n377_33[1]),.dout(n2909),.clk(gclk));
	jor g2647(.dina(n2909),.dinb(n2908),.dout(n2910),.clk(gclk));
	jand g2648(.dina(w_n2227_0[2]),.dinb(w_n432_33[1]),.dout(n2911),.clk(gclk));
	jand g2649(.dina(w_n2263_0[2]),.dinb(w_n485_33[1]),.dout(n2912),.clk(gclk));
	jor g2650(.dina(n2912),.dinb(n2911),.dout(n2913),.clk(gclk));
	jor g2651(.dina(n2913),.dinb(n2910),.dout(n2914),.clk(gclk));
	jand g2652(.dina(w_n2914_0[1]),.dinb(w_n263_48[1]),.dout(n2915),.clk(gclk));
	jand g2653(.dina(w_n2238_0[2]),.dinb(w_n323_33[0]),.dout(n2916),.clk(gclk));
	jand g2654(.dina(w_n2202_0[2]),.dinb(w_n377_33[0]),.dout(n2917),.clk(gclk));
	jor g2655(.dina(n2917),.dinb(n2916),.dout(n2918),.clk(gclk));
	jand g2656(.dina(w_n2255_0[2]),.dinb(w_n432_33[0]),.dout(n2919),.clk(gclk));
	jand g2657(.dina(w_n2219_0[2]),.dinb(w_n485_33[0]),.dout(n2920),.clk(gclk));
	jor g2658(.dina(n2920),.dinb(n2919),.dout(n2921),.clk(gclk));
	jor g2659(.dina(n2921),.dinb(n2918),.dout(n2922),.clk(gclk));
	jand g2660(.dina(w_n2922_0[1]),.dinb(w_shift6_48[1]),.dout(n2923),.clk(gclk));
	jor g2661(.dina(n2923),.dinb(n2915),.dout(result45),.clk(gclk));
	jand g2662(.dina(w_n2283_0[2]),.dinb(w_n323_32[2]),.dout(n2925),.clk(gclk));
	jand g2663(.dina(w_n2319_0[2]),.dinb(w_n377_32[2]),.dout(n2926),.clk(gclk));
	jor g2664(.dina(n2926),.dinb(n2925),.dout(n2927),.clk(gclk));
	jand g2665(.dina(w_n2300_0[2]),.dinb(w_n432_32[2]),.dout(n2928),.clk(gclk));
	jand g2666(.dina(w_n2336_0[2]),.dinb(w_n485_32[2]),.dout(n2929),.clk(gclk));
	jor g2667(.dina(n2929),.dinb(n2928),.dout(n2930),.clk(gclk));
	jor g2668(.dina(n2930),.dinb(n2927),.dout(n2931),.clk(gclk));
	jand g2669(.dina(w_n2931_0[1]),.dinb(w_n263_48[0]),.dout(n2932),.clk(gclk));
	jand g2670(.dina(w_n2311_0[2]),.dinb(w_n323_32[1]),.dout(n2933),.clk(gclk));
	jand g2671(.dina(w_n2275_0[2]),.dinb(w_n377_32[1]),.dout(n2934),.clk(gclk));
	jor g2672(.dina(n2934),.dinb(n2933),.dout(n2935),.clk(gclk));
	jand g2673(.dina(w_n2328_0[2]),.dinb(w_n432_32[1]),.dout(n2936),.clk(gclk));
	jand g2674(.dina(w_n2292_0[2]),.dinb(w_n485_32[1]),.dout(n2937),.clk(gclk));
	jor g2675(.dina(n2937),.dinb(n2936),.dout(n2938),.clk(gclk));
	jor g2676(.dina(n2938),.dinb(n2935),.dout(n2939),.clk(gclk));
	jand g2677(.dina(w_n2939_0[1]),.dinb(w_shift6_48[0]),.dout(n2940),.clk(gclk));
	jor g2678(.dina(n2940),.dinb(n2932),.dout(result46),.clk(gclk));
	jand g2679(.dina(w_n2356_0[2]),.dinb(w_n323_32[0]),.dout(n2942),.clk(gclk));
	jand g2680(.dina(w_n2392_0[2]),.dinb(w_n377_32[0]),.dout(n2943),.clk(gclk));
	jor g2681(.dina(n2943),.dinb(n2942),.dout(n2944),.clk(gclk));
	jand g2682(.dina(w_n2373_0[2]),.dinb(w_n432_32[0]),.dout(n2945),.clk(gclk));
	jand g2683(.dina(w_n2409_0[2]),.dinb(w_n485_32[0]),.dout(n2946),.clk(gclk));
	jor g2684(.dina(n2946),.dinb(n2945),.dout(n2947),.clk(gclk));
	jor g2685(.dina(n2947),.dinb(n2944),.dout(n2948),.clk(gclk));
	jand g2686(.dina(w_n2948_0[1]),.dinb(w_n263_47[2]),.dout(n2949),.clk(gclk));
	jand g2687(.dina(w_n2384_0[2]),.dinb(w_n323_31[2]),.dout(n2950),.clk(gclk));
	jand g2688(.dina(w_n2348_0[2]),.dinb(w_n377_31[2]),.dout(n2951),.clk(gclk));
	jor g2689(.dina(n2951),.dinb(n2950),.dout(n2952),.clk(gclk));
	jand g2690(.dina(w_n2401_0[2]),.dinb(w_n432_31[2]),.dout(n2953),.clk(gclk));
	jand g2691(.dina(w_n2365_0[2]),.dinb(w_n485_31[2]),.dout(n2954),.clk(gclk));
	jor g2692(.dina(n2954),.dinb(n2953),.dout(n2955),.clk(gclk));
	jor g2693(.dina(n2955),.dinb(n2952),.dout(n2956),.clk(gclk));
	jand g2694(.dina(w_n2956_0[1]),.dinb(w_shift6_47[2]),.dout(n2957),.clk(gclk));
	jor g2695(.dina(n2957),.dinb(n2949),.dout(result47),.clk(gclk));
	jand g2696(.dina(w_n484_0[1]),.dinb(w_n323_31[1]),.dout(n2959),.clk(gclk));
	jand g2697(.dina(w_n643_0[1]),.dinb(w_n377_31[1]),.dout(n2960),.clk(gclk));
	jor g2698(.dina(n2960),.dinb(n2959),.dout(n2961),.clk(gclk));
	jand g2699(.dina(w_n540_0[1]),.dinb(w_n432_31[1]),.dout(n2962),.clk(gclk));
	jand g2700(.dina(w_n590_0[1]),.dinb(w_n485_31[1]),.dout(n2963),.clk(gclk));
	jor g2701(.dina(n2963),.dinb(n2962),.dout(n2964),.clk(gclk));
	jor g2702(.dina(n2964),.dinb(n2961),.dout(n2965),.clk(gclk));
	jand g2703(.dina(w_n2965_0[1]),.dinb(w_n263_47[1]),.dout(n2966),.clk(gclk));
	jand g2704(.dina(w_n432_31[0]),.dinb(w_n322_0[1]),.dout(n2967),.clk(gclk));
	jand g2705(.dina(w_n485_31[0]),.dinb(w_n375_0[1]),.dout(n2968),.clk(gclk));
	jor g2706(.dina(n2968),.dinb(n2967),.dout(n2969),.clk(gclk));
	jand g2707(.dina(w_n430_0[1]),.dinb(w_n377_31[0]),.dout(n2970),.clk(gclk));
	jand g2708(.dina(w_n695_0[1]),.dinb(w_n323_31[0]),.dout(n2971),.clk(gclk));
	jor g2709(.dina(n2971),.dinb(n2970),.dout(n2972),.clk(gclk));
	jor g2710(.dina(n2972),.dinb(n2969),.dout(n2973),.clk(gclk));
	jand g2711(.dina(w_n2973_0[1]),.dinb(w_shift6_47[1]),.dout(n2974),.clk(gclk));
	jor g2712(.dina(n2974),.dinb(n2966),.dout(result48),.clk(gclk));
	jand g2713(.dina(w_n876_0[1]),.dinb(w_n323_30[2]),.dout(n2976),.clk(gclk));
	jand g2714(.dina(w_n967_0[1]),.dinb(w_n377_30[2]),.dout(n2977),.clk(gclk));
	jor g2715(.dina(n2977),.dinb(n2976),.dout(n2978),.clk(gclk));
	jand g2716(.dina(w_n1012_0[1]),.dinb(w_n432_30[2]),.dout(n2979),.clk(gclk));
	jand g2717(.dina(w_n1060_0[1]),.dinb(w_n485_30[2]),.dout(n2980),.clk(gclk));
	jor g2718(.dina(n2980),.dinb(n2979),.dout(n2981),.clk(gclk));
	jor g2719(.dina(n2981),.dinb(n2978),.dout(n2982),.clk(gclk));
	jand g2720(.dina(w_n2982_0[1]),.dinb(w_n263_47[0]),.dout(n2983),.clk(gclk));
	jand g2721(.dina(w_n923_0[1]),.dinb(w_n323_30[1]),.dout(n2984),.clk(gclk));
	jand g2722(.dina(w_n832_0[1]),.dinb(w_n377_30[1]),.dout(n2985),.clk(gclk));
	jor g2723(.dina(n2985),.dinb(n2984),.dout(n2986),.clk(gclk));
	jand g2724(.dina(w_n743_0[1]),.dinb(w_n432_30[1]),.dout(n2987),.clk(gclk));
	jand g2725(.dina(w_n787_0[1]),.dinb(w_n485_30[1]),.dout(n2988),.clk(gclk));
	jor g2726(.dina(n2988),.dinb(n2987),.dout(n2989),.clk(gclk));
	jor g2727(.dina(n2989),.dinb(n2986),.dout(n2990),.clk(gclk));
	jand g2728(.dina(w_n2990_0[1]),.dinb(w_shift6_47[0]),.dout(n2991),.clk(gclk));
	jor g2729(.dina(n2991),.dinb(n2983),.dout(result49),.clk(gclk));
	jand g2730(.dina(w_n1209_0[1]),.dinb(w_n323_30[0]),.dout(n2993),.clk(gclk));
	jand g2731(.dina(w_n1284_0[1]),.dinb(w_n377_30[0]),.dout(n2994),.clk(gclk));
	jor g2732(.dina(n2994),.dinb(n2993),.dout(n2995),.clk(gclk));
	jand g2733(.dina(w_n1321_0[1]),.dinb(w_n432_30[0]),.dout(n2996),.clk(gclk));
	jand g2734(.dina(w_n1357_0[1]),.dinb(w_n485_30[0]),.dout(n2997),.clk(gclk));
	jor g2735(.dina(n2997),.dinb(n2996),.dout(n2998),.clk(gclk));
	jor g2736(.dina(n2998),.dinb(n2995),.dout(n2999),.clk(gclk));
	jand g2737(.dina(w_n2999_0[1]),.dinb(w_n263_46[2]),.dout(n3000),.clk(gclk));
	jand g2738(.dina(w_n1248_0[1]),.dinb(w_n323_29[2]),.dout(n3001),.clk(gclk));
	jand g2739(.dina(w_n1173_0[1]),.dinb(w_n377_29[2]),.dout(n3002),.clk(gclk));
	jor g2740(.dina(n3002),.dinb(n3001),.dout(n3003),.clk(gclk));
	jand g2741(.dina(w_n1100_0[1]),.dinb(w_n432_29[2]),.dout(n3004),.clk(gclk));
	jand g2742(.dina(w_n1136_0[1]),.dinb(w_n485_29[2]),.dout(n3005),.clk(gclk));
	jor g2743(.dina(n3005),.dinb(n3004),.dout(n3006),.clk(gclk));
	jor g2744(.dina(n3006),.dinb(n3003),.dout(n3007),.clk(gclk));
	jand g2745(.dina(w_n3007_0[1]),.dinb(w_shift6_46[2]),.dout(n3008),.clk(gclk));
	jor g2746(.dina(n3008),.dinb(n3000),.dout(result50),.clk(gclk));
	jand g2747(.dina(w_n1513_0[1]),.dinb(w_n485_29[1]),.dout(n3010),.clk(gclk));
	jand g2748(.dina(w_n1533_0[1]),.dinb(w_n432_29[1]),.dout(n3011),.clk(gclk));
	jor g2749(.dina(n3011),.dinb(n3010),.dout(n3012),.clk(gclk));
	jand g2750(.dina(w_n1485_0[1]),.dinb(w_n377_29[1]),.dout(n3013),.clk(gclk));
	jand g2751(.dina(w_n1442_0[1]),.dinb(w_n323_29[1]),.dout(n3014),.clk(gclk));
	jor g2752(.dina(n3014),.dinb(n3013),.dout(n3015),.clk(gclk));
	jor g2753(.dina(n3015),.dinb(n3012),.dout(n3016),.clk(gclk));
	jand g2754(.dina(w_n3016_0[1]),.dinb(w_n263_46[1]),.dout(n3017),.clk(gclk));
	jand g2755(.dina(w_n1465_0[1]),.dinb(w_n323_29[0]),.dout(n3018),.clk(gclk));
	jand g2756(.dina(w_n1422_0[1]),.dinb(w_n377_29[0]),.dout(n3019),.clk(gclk));
	jor g2757(.dina(n3019),.dinb(n3018),.dout(n3020),.clk(gclk));
	jand g2758(.dina(w_n1381_0[1]),.dinb(w_n485_29[0]),.dout(n3021),.clk(gclk));
	jand g2759(.dina(w_n1401_0[1]),.dinb(w_n432_29[0]),.dout(n3022),.clk(gclk));
	jor g2760(.dina(n3022),.dinb(n3021),.dout(n3023),.clk(gclk));
	jor g2761(.dina(n3023),.dinb(n3020),.dout(n3024),.clk(gclk));
	jand g2762(.dina(w_n3024_0[1]),.dinb(w_shift6_46[1]),.dout(n3025),.clk(gclk));
	jor g2763(.dina(n3025),.dinb(n3017),.dout(result51),.clk(gclk));
	jand g2764(.dina(w_n1581_0[1]),.dinb(w_n485_28[2]),.dout(n3027),.clk(gclk));
	jand g2765(.dina(w_n1589_0[1]),.dinb(w_n432_28[2]),.dout(n3028),.clk(gclk));
	jor g2766(.dina(n3028),.dinb(n3027),.dout(n3029),.clk(gclk));
	jand g2767(.dina(w_n1570_0[1]),.dinb(w_n323_28[2]),.dout(n3030),.clk(gclk));
	jand g2768(.dina(w_n1606_0[1]),.dinb(w_n377_28[2]),.dout(n3031),.clk(gclk));
	jor g2769(.dina(n3031),.dinb(n3030),.dout(n3032),.clk(gclk));
	jor g2770(.dina(n3032),.dinb(n3029),.dout(n3033),.clk(gclk));
	jand g2771(.dina(w_n3033_0[1]),.dinb(w_n263_46[0]),.dout(n3034),.clk(gclk));
	jand g2772(.dina(w_n1545_0[1]),.dinb(w_n432_28[1]),.dout(n3035),.clk(gclk));
	jand g2773(.dina(w_n1598_0[1]),.dinb(w_n323_28[1]),.dout(n3036),.clk(gclk));
	jor g2774(.dina(n3036),.dinb(n3035),.dout(n3037),.clk(gclk));
	jand g2775(.dina(w_n1562_0[1]),.dinb(w_n377_28[1]),.dout(n3038),.clk(gclk));
	jand g2776(.dina(w_n1553_0[1]),.dinb(w_n485_28[1]),.dout(n3039),.clk(gclk));
	jor g2777(.dina(n3039),.dinb(n3038),.dout(n3040),.clk(gclk));
	jor g2778(.dina(n3040),.dinb(n3037),.dout(n3041),.clk(gclk));
	jand g2779(.dina(w_n3041_0[1]),.dinb(w_shift6_46[0]),.dout(n3042),.clk(gclk));
	jor g2780(.dina(n3042),.dinb(n3034),.dout(result52),.clk(gclk));
	jand g2781(.dina(w_n1654_0[1]),.dinb(w_n485_28[0]),.dout(n3044),.clk(gclk));
	jand g2782(.dina(w_n1662_0[1]),.dinb(w_n432_28[0]),.dout(n3045),.clk(gclk));
	jor g2783(.dina(n3045),.dinb(n3044),.dout(n3046),.clk(gclk));
	jand g2784(.dina(w_n1643_0[1]),.dinb(w_n323_28[0]),.dout(n3047),.clk(gclk));
	jand g2785(.dina(w_n1679_0[1]),.dinb(w_n377_28[0]),.dout(n3048),.clk(gclk));
	jor g2786(.dina(n3048),.dinb(n3047),.dout(n3049),.clk(gclk));
	jor g2787(.dina(n3049),.dinb(n3046),.dout(n3050),.clk(gclk));
	jand g2788(.dina(w_n3050_0[1]),.dinb(w_n263_45[2]),.dout(n3051),.clk(gclk));
	jand g2789(.dina(w_n1618_0[1]),.dinb(w_n432_27[2]),.dout(n3052),.clk(gclk));
	jand g2790(.dina(w_n1671_0[1]),.dinb(w_n323_27[2]),.dout(n3053),.clk(gclk));
	jor g2791(.dina(n3053),.dinb(n3052),.dout(n3054),.clk(gclk));
	jand g2792(.dina(w_n1635_0[1]),.dinb(w_n377_27[2]),.dout(n3055),.clk(gclk));
	jand g2793(.dina(w_n1626_0[1]),.dinb(w_n485_27[2]),.dout(n3056),.clk(gclk));
	jor g2794(.dina(n3056),.dinb(n3055),.dout(n3057),.clk(gclk));
	jor g2795(.dina(n3057),.dinb(n3054),.dout(n3058),.clk(gclk));
	jand g2796(.dina(w_n3058_0[1]),.dinb(w_shift6_45[2]),.dout(n3059),.clk(gclk));
	jor g2797(.dina(n3059),.dinb(n3051),.dout(result53),.clk(gclk));
	jand g2798(.dina(w_n1727_0[1]),.dinb(w_n485_27[1]),.dout(n3061),.clk(gclk));
	jand g2799(.dina(w_n1735_0[1]),.dinb(w_n432_27[1]),.dout(n3062),.clk(gclk));
	jor g2800(.dina(n3062),.dinb(n3061),.dout(n3063),.clk(gclk));
	jand g2801(.dina(w_n1716_0[1]),.dinb(w_n323_27[1]),.dout(n3064),.clk(gclk));
	jand g2802(.dina(w_n1752_0[1]),.dinb(w_n377_27[1]),.dout(n3065),.clk(gclk));
	jor g2803(.dina(n3065),.dinb(n3064),.dout(n3066),.clk(gclk));
	jor g2804(.dina(n3066),.dinb(n3063),.dout(n3067),.clk(gclk));
	jand g2805(.dina(w_n3067_0[1]),.dinb(w_n263_45[1]),.dout(n3068),.clk(gclk));
	jand g2806(.dina(w_n1691_0[1]),.dinb(w_n432_27[0]),.dout(n3069),.clk(gclk));
	jand g2807(.dina(w_n1744_0[1]),.dinb(w_n323_27[0]),.dout(n3070),.clk(gclk));
	jor g2808(.dina(n3070),.dinb(n3069),.dout(n3071),.clk(gclk));
	jand g2809(.dina(w_n1708_0[1]),.dinb(w_n377_27[0]),.dout(n3072),.clk(gclk));
	jand g2810(.dina(w_n1699_0[1]),.dinb(w_n485_27[0]),.dout(n3073),.clk(gclk));
	jor g2811(.dina(n3073),.dinb(n3072),.dout(n3074),.clk(gclk));
	jor g2812(.dina(n3074),.dinb(n3071),.dout(n3075),.clk(gclk));
	jand g2813(.dina(w_n3075_0[1]),.dinb(w_shift6_45[1]),.dout(n3076),.clk(gclk));
	jor g2814(.dina(n3076),.dinb(n3068),.dout(result54),.clk(gclk));
	jand g2815(.dina(w_n1800_0[1]),.dinb(w_n485_26[2]),.dout(n3078),.clk(gclk));
	jand g2816(.dina(w_n1825_0[1]),.dinb(w_n377_26[2]),.dout(n3079),.clk(gclk));
	jor g2817(.dina(n3079),.dinb(n3078),.dout(n3080),.clk(gclk));
	jand g2818(.dina(w_n1808_0[1]),.dinb(w_n432_26[2]),.dout(n3081),.clk(gclk));
	jand g2819(.dina(w_n1789_0[1]),.dinb(w_n323_26[2]),.dout(n3082),.clk(gclk));
	jor g2820(.dina(n3082),.dinb(n3081),.dout(n3083),.clk(gclk));
	jor g2821(.dina(n3083),.dinb(n3080),.dout(n3084),.clk(gclk));
	jand g2822(.dina(w_n3084_0[1]),.dinb(w_n263_45[0]),.dout(n3085),.clk(gclk));
	jand g2823(.dina(w_n1817_0[1]),.dinb(w_n323_26[1]),.dout(n3086),.clk(gclk));
	jand g2824(.dina(w_n1781_0[1]),.dinb(w_n377_26[1]),.dout(n3087),.clk(gclk));
	jor g2825(.dina(n3087),.dinb(n3086),.dout(n3088),.clk(gclk));
	jand g2826(.dina(w_n1764_0[1]),.dinb(w_n432_26[1]),.dout(n3089),.clk(gclk));
	jand g2827(.dina(w_n1772_0[1]),.dinb(w_n485_26[1]),.dout(n3090),.clk(gclk));
	jor g2828(.dina(n3090),.dinb(n3089),.dout(n3091),.clk(gclk));
	jor g2829(.dina(n3091),.dinb(n3088),.dout(n3092),.clk(gclk));
	jand g2830(.dina(w_n3092_0[1]),.dinb(w_shift6_45[0]),.dout(n3093),.clk(gclk));
	jor g2831(.dina(n3093),.dinb(n3085),.dout(result55),.clk(gclk));
	jand g2832(.dina(w_n1873_0[1]),.dinb(w_n485_26[0]),.dout(n3095),.clk(gclk));
	jand g2833(.dina(w_n1898_0[1]),.dinb(w_n377_26[0]),.dout(n3096),.clk(gclk));
	jor g2834(.dina(n3096),.dinb(n3095),.dout(n3097),.clk(gclk));
	jand g2835(.dina(w_n1881_0[1]),.dinb(w_n432_26[0]),.dout(n3098),.clk(gclk));
	jand g2836(.dina(w_n1862_0[1]),.dinb(w_n323_26[0]),.dout(n3099),.clk(gclk));
	jor g2837(.dina(n3099),.dinb(n3098),.dout(n3100),.clk(gclk));
	jor g2838(.dina(n3100),.dinb(n3097),.dout(n3101),.clk(gclk));
	jand g2839(.dina(w_n3101_0[1]),.dinb(w_n263_44[2]),.dout(n3102),.clk(gclk));
	jand g2840(.dina(w_n1890_0[1]),.dinb(w_n323_25[2]),.dout(n3103),.clk(gclk));
	jand g2841(.dina(w_n1854_0[1]),.dinb(w_n377_25[2]),.dout(n3104),.clk(gclk));
	jor g2842(.dina(n3104),.dinb(n3103),.dout(n3105),.clk(gclk));
	jand g2843(.dina(w_n1837_0[1]),.dinb(w_n432_25[2]),.dout(n3106),.clk(gclk));
	jand g2844(.dina(w_n1845_0[1]),.dinb(w_n485_25[2]),.dout(n3107),.clk(gclk));
	jor g2845(.dina(n3107),.dinb(n3106),.dout(n3108),.clk(gclk));
	jor g2846(.dina(n3108),.dinb(n3105),.dout(n3109),.clk(gclk));
	jand g2847(.dina(w_n3109_0[1]),.dinb(w_shift6_44[2]),.dout(n3110),.clk(gclk));
	jor g2848(.dina(n3110),.dinb(n3102),.dout(result56),.clk(gclk));
	jand g2849(.dina(w_n1946_0[1]),.dinb(w_n485_25[1]),.dout(n3112),.clk(gclk));
	jand g2850(.dina(w_n1971_0[1]),.dinb(w_n377_25[1]),.dout(n3113),.clk(gclk));
	jor g2851(.dina(n3113),.dinb(n3112),.dout(n3114),.clk(gclk));
	jand g2852(.dina(w_n1954_0[1]),.dinb(w_n432_25[1]),.dout(n3115),.clk(gclk));
	jand g2853(.dina(w_n1935_0[1]),.dinb(w_n323_25[1]),.dout(n3116),.clk(gclk));
	jor g2854(.dina(n3116),.dinb(n3115),.dout(n3117),.clk(gclk));
	jor g2855(.dina(n3117),.dinb(n3114),.dout(n3118),.clk(gclk));
	jand g2856(.dina(w_n3118_0[1]),.dinb(w_n263_44[1]),.dout(n3119),.clk(gclk));
	jand g2857(.dina(w_n1963_0[1]),.dinb(w_n323_25[0]),.dout(n3120),.clk(gclk));
	jand g2858(.dina(w_n1927_0[1]),.dinb(w_n377_25[0]),.dout(n3121),.clk(gclk));
	jor g2859(.dina(n3121),.dinb(n3120),.dout(n3122),.clk(gclk));
	jand g2860(.dina(w_n1910_0[1]),.dinb(w_n432_25[0]),.dout(n3123),.clk(gclk));
	jand g2861(.dina(w_n1918_0[1]),.dinb(w_n485_25[0]),.dout(n3124),.clk(gclk));
	jor g2862(.dina(n3124),.dinb(n3123),.dout(n3125),.clk(gclk));
	jor g2863(.dina(n3125),.dinb(n3122),.dout(n3126),.clk(gclk));
	jand g2864(.dina(w_n3126_0[1]),.dinb(w_shift6_44[1]),.dout(n3127),.clk(gclk));
	jor g2865(.dina(n3127),.dinb(n3119),.dout(result57),.clk(gclk));
	jand g2866(.dina(w_n2019_0[1]),.dinb(w_n485_24[2]),.dout(n3129),.clk(gclk));
	jand g2867(.dina(w_n2027_0[1]),.dinb(w_n432_24[2]),.dout(n3130),.clk(gclk));
	jor g2868(.dina(n3130),.dinb(n3129),.dout(n3131),.clk(gclk));
	jand g2869(.dina(w_n2008_0[1]),.dinb(w_n323_24[2]),.dout(n3132),.clk(gclk));
	jand g2870(.dina(w_n2044_0[1]),.dinb(w_n377_24[2]),.dout(n3133),.clk(gclk));
	jor g2871(.dina(n3133),.dinb(n3132),.dout(n3134),.clk(gclk));
	jor g2872(.dina(n3134),.dinb(n3131),.dout(n3135),.clk(gclk));
	jand g2873(.dina(w_n3135_0[1]),.dinb(w_n263_44[0]),.dout(n3136),.clk(gclk));
	jand g2874(.dina(w_n2036_0[1]),.dinb(w_n323_24[1]),.dout(n3137),.clk(gclk));
	jand g2875(.dina(w_n2000_0[1]),.dinb(w_n377_24[1]),.dout(n3138),.clk(gclk));
	jor g2876(.dina(n3138),.dinb(n3137),.dout(n3139),.clk(gclk));
	jand g2877(.dina(w_n1983_0[1]),.dinb(w_n432_24[1]),.dout(n3140),.clk(gclk));
	jand g2878(.dina(w_n1991_0[1]),.dinb(w_n485_24[1]),.dout(n3141),.clk(gclk));
	jor g2879(.dina(n3141),.dinb(n3140),.dout(n3142),.clk(gclk));
	jor g2880(.dina(n3142),.dinb(n3139),.dout(n3143),.clk(gclk));
	jand g2881(.dina(w_n3143_0[1]),.dinb(w_shift6_44[0]),.dout(n3144),.clk(gclk));
	jor g2882(.dina(n3144),.dinb(n3136),.dout(result58),.clk(gclk));
	jand g2883(.dina(w_n2092_0[1]),.dinb(w_n485_24[0]),.dout(n3146),.clk(gclk));
	jand g2884(.dina(w_n2100_0[1]),.dinb(w_n432_24[0]),.dout(n3147),.clk(gclk));
	jor g2885(.dina(n3147),.dinb(n3146),.dout(n3148),.clk(gclk));
	jand g2886(.dina(w_n2081_0[1]),.dinb(w_n323_24[0]),.dout(n3149),.clk(gclk));
	jand g2887(.dina(w_n2117_0[1]),.dinb(w_n377_24[0]),.dout(n3150),.clk(gclk));
	jor g2888(.dina(n3150),.dinb(n3149),.dout(n3151),.clk(gclk));
	jor g2889(.dina(n3151),.dinb(n3148),.dout(n3152),.clk(gclk));
	jand g2890(.dina(w_n3152_0[1]),.dinb(w_n263_43[2]),.dout(n3153),.clk(gclk));
	jand g2891(.dina(w_n2109_0[1]),.dinb(w_n323_23[2]),.dout(n3154),.clk(gclk));
	jand g2892(.dina(w_n2073_0[1]),.dinb(w_n377_23[2]),.dout(n3155),.clk(gclk));
	jor g2893(.dina(n3155),.dinb(n3154),.dout(n3156),.clk(gclk));
	jand g2894(.dina(w_n2056_0[1]),.dinb(w_n432_23[2]),.dout(n3157),.clk(gclk));
	jand g2895(.dina(w_n2064_0[1]),.dinb(w_n485_23[2]),.dout(n3158),.clk(gclk));
	jor g2896(.dina(n3158),.dinb(n3157),.dout(n3159),.clk(gclk));
	jor g2897(.dina(n3159),.dinb(n3156),.dout(n3160),.clk(gclk));
	jand g2898(.dina(w_n3160_0[1]),.dinb(w_shift6_43[2]),.dout(n3161),.clk(gclk));
	jor g2899(.dina(n3161),.dinb(n3153),.dout(result59),.clk(gclk));
	jand g2900(.dina(w_n2165_0[1]),.dinb(w_n485_23[1]),.dout(n3163),.clk(gclk));
	jand g2901(.dina(w_n2173_0[1]),.dinb(w_n432_23[1]),.dout(n3164),.clk(gclk));
	jor g2902(.dina(n3164),.dinb(n3163),.dout(n3165),.clk(gclk));
	jand g2903(.dina(w_n2154_0[1]),.dinb(w_n323_23[1]),.dout(n3166),.clk(gclk));
	jand g2904(.dina(w_n2190_0[1]),.dinb(w_n377_23[1]),.dout(n3167),.clk(gclk));
	jor g2905(.dina(n3167),.dinb(n3166),.dout(n3168),.clk(gclk));
	jor g2906(.dina(n3168),.dinb(n3165),.dout(n3169),.clk(gclk));
	jand g2907(.dina(w_n3169_0[1]),.dinb(w_n263_43[1]),.dout(n3170),.clk(gclk));
	jand g2908(.dina(w_n2182_0[1]),.dinb(w_n323_23[0]),.dout(n3171),.clk(gclk));
	jand g2909(.dina(w_n2146_0[1]),.dinb(w_n377_23[0]),.dout(n3172),.clk(gclk));
	jor g2910(.dina(n3172),.dinb(n3171),.dout(n3173),.clk(gclk));
	jand g2911(.dina(w_n2129_0[1]),.dinb(w_n432_23[0]),.dout(n3174),.clk(gclk));
	jand g2912(.dina(w_n2137_0[1]),.dinb(w_n485_23[0]),.dout(n3175),.clk(gclk));
	jor g2913(.dina(n3175),.dinb(n3174),.dout(n3176),.clk(gclk));
	jor g2914(.dina(n3176),.dinb(n3173),.dout(n3177),.clk(gclk));
	jand g2915(.dina(w_n3177_0[1]),.dinb(w_shift6_43[1]),.dout(n3178),.clk(gclk));
	jor g2916(.dina(n3178),.dinb(n3170),.dout(result60),.clk(gclk));
	jand g2917(.dina(w_n2238_0[1]),.dinb(w_n485_22[2]),.dout(n3180),.clk(gclk));
	jand g2918(.dina(w_n2246_0[1]),.dinb(w_n432_22[2]),.dout(n3181),.clk(gclk));
	jor g2919(.dina(n3181),.dinb(n3180),.dout(n3182),.clk(gclk));
	jand g2920(.dina(w_n2227_0[1]),.dinb(w_n323_22[2]),.dout(n3183),.clk(gclk));
	jand g2921(.dina(w_n2263_0[1]),.dinb(w_n377_22[2]),.dout(n3184),.clk(gclk));
	jor g2922(.dina(n3184),.dinb(n3183),.dout(n3185),.clk(gclk));
	jor g2923(.dina(n3185),.dinb(n3182),.dout(n3186),.clk(gclk));
	jand g2924(.dina(w_n3186_0[1]),.dinb(w_n263_43[0]),.dout(n3187),.clk(gclk));
	jand g2925(.dina(w_n2255_0[1]),.dinb(w_n323_22[1]),.dout(n3188),.clk(gclk));
	jand g2926(.dina(w_n2219_0[1]),.dinb(w_n377_22[1]),.dout(n3189),.clk(gclk));
	jor g2927(.dina(n3189),.dinb(n3188),.dout(n3190),.clk(gclk));
	jand g2928(.dina(w_n2202_0[1]),.dinb(w_n432_22[1]),.dout(n3191),.clk(gclk));
	jand g2929(.dina(w_n2210_0[1]),.dinb(w_n485_22[1]),.dout(n3192),.clk(gclk));
	jor g2930(.dina(n3192),.dinb(n3191),.dout(n3193),.clk(gclk));
	jor g2931(.dina(n3193),.dinb(n3190),.dout(n3194),.clk(gclk));
	jand g2932(.dina(w_n3194_0[1]),.dinb(w_shift6_43[0]),.dout(n3195),.clk(gclk));
	jor g2933(.dina(n3195),.dinb(n3187),.dout(result61),.clk(gclk));
	jand g2934(.dina(w_n2311_0[1]),.dinb(w_n485_22[0]),.dout(n3197),.clk(gclk));
	jand g2935(.dina(w_n2319_0[1]),.dinb(w_n432_22[0]),.dout(n3198),.clk(gclk));
	jor g2936(.dina(n3198),.dinb(n3197),.dout(n3199),.clk(gclk));
	jand g2937(.dina(w_n2300_0[1]),.dinb(w_n323_22[0]),.dout(n3200),.clk(gclk));
	jand g2938(.dina(w_n2336_0[1]),.dinb(w_n377_22[0]),.dout(n3201),.clk(gclk));
	jor g2939(.dina(n3201),.dinb(n3200),.dout(n3202),.clk(gclk));
	jor g2940(.dina(n3202),.dinb(n3199),.dout(n3203),.clk(gclk));
	jand g2941(.dina(w_n3203_0[1]),.dinb(w_n263_42[2]),.dout(n3204),.clk(gclk));
	jand g2942(.dina(w_n2328_0[1]),.dinb(w_n323_21[2]),.dout(n3205),.clk(gclk));
	jand g2943(.dina(w_n2292_0[1]),.dinb(w_n377_21[2]),.dout(n3206),.clk(gclk));
	jor g2944(.dina(n3206),.dinb(n3205),.dout(n3207),.clk(gclk));
	jand g2945(.dina(w_n2275_0[1]),.dinb(w_n432_21[2]),.dout(n3208),.clk(gclk));
	jand g2946(.dina(w_n2283_0[1]),.dinb(w_n485_21[2]),.dout(n3209),.clk(gclk));
	jor g2947(.dina(n3209),.dinb(n3208),.dout(n3210),.clk(gclk));
	jor g2948(.dina(n3210),.dinb(n3207),.dout(n3211),.clk(gclk));
	jand g2949(.dina(w_n3211_0[1]),.dinb(w_shift6_42[2]),.dout(n3212),.clk(gclk));
	jor g2950(.dina(n3212),.dinb(n3204),.dout(result62),.clk(gclk));
	jand g2951(.dina(w_n2384_0[1]),.dinb(w_n485_21[1]),.dout(n3214),.clk(gclk));
	jand g2952(.dina(w_n2392_0[1]),.dinb(w_n432_21[1]),.dout(n3215),.clk(gclk));
	jor g2953(.dina(n3215),.dinb(n3214),.dout(n3216),.clk(gclk));
	jand g2954(.dina(w_n2373_0[1]),.dinb(w_n323_21[1]),.dout(n3217),.clk(gclk));
	jand g2955(.dina(w_n2409_0[1]),.dinb(w_n377_21[1]),.dout(n3218),.clk(gclk));
	jor g2956(.dina(n3218),.dinb(n3217),.dout(n3219),.clk(gclk));
	jor g2957(.dina(n3219),.dinb(n3216),.dout(n3220),.clk(gclk));
	jand g2958(.dina(w_n3220_0[1]),.dinb(w_n263_42[1]),.dout(n3221),.clk(gclk));
	jand g2959(.dina(w_n2401_0[1]),.dinb(w_n323_21[0]),.dout(n3222),.clk(gclk));
	jand g2960(.dina(w_n2365_0[1]),.dinb(w_n377_21[0]),.dout(n3223),.clk(gclk));
	jor g2961(.dina(n3223),.dinb(n3222),.dout(n3224),.clk(gclk));
	jand g2962(.dina(w_n2348_0[1]),.dinb(w_n432_21[0]),.dout(n3225),.clk(gclk));
	jand g2963(.dina(w_n2356_0[1]),.dinb(w_n485_21[0]),.dout(n3226),.clk(gclk));
	jor g2964(.dina(n3226),.dinb(n3225),.dout(n3227),.clk(gclk));
	jor g2965(.dina(n3227),.dinb(n3224),.dout(n3228),.clk(gclk));
	jand g2966(.dina(w_n3228_0[1]),.dinb(w_shift6_42[1]),.dout(n3229),.clk(gclk));
	jor g2967(.dina(n3229),.dinb(n3221),.dout(result63),.clk(gclk));
	jand g2968(.dina(w_n698_0[0]),.dinb(w_n263_42[0]),.dout(n3231),.clk(gclk));
	jand g2969(.dina(w_n488_0[0]),.dinb(w_shift6_42[0]),.dout(n3232),.clk(gclk));
	jor g2970(.dina(n3232),.dinb(n3231),.dout(result64),.clk(gclk));
	jand g2971(.dina(w_n1063_0[0]),.dinb(w_n263_41[2]),.dout(n3234),.clk(gclk));
	jand g2972(.dina(w_n879_0[0]),.dinb(w_shift6_41[2]),.dout(n3235),.clk(gclk));
	jor g2973(.dina(n3235),.dinb(n3234),.dout(result65),.clk(gclk));
	jand g2974(.dina(w_n1360_0[0]),.dinb(w_n263_41[1]),.dout(n3237),.clk(gclk));
	jand g2975(.dina(w_n1212_0[0]),.dinb(w_shift6_41[1]),.dout(n3238),.clk(gclk));
	jor g2976(.dina(n3238),.dinb(n3237),.dout(result66),.clk(gclk));
	jand g2977(.dina(w_n1536_0[0]),.dinb(w_n263_41[0]),.dout(n3240),.clk(gclk));
	jand g2978(.dina(w_n1445_0[0]),.dinb(w_shift6_41[0]),.dout(n3241),.clk(gclk));
	jor g2979(.dina(n3241),.dinb(n3240),.dout(result67),.clk(gclk));
	jand g2980(.dina(w_n1609_0[0]),.dinb(w_n263_40[2]),.dout(n3243),.clk(gclk));
	jand g2981(.dina(w_n1573_0[0]),.dinb(w_shift6_40[2]),.dout(n3244),.clk(gclk));
	jor g2982(.dina(n3244),.dinb(n3243),.dout(result68),.clk(gclk));
	jand g2983(.dina(w_n1682_0[0]),.dinb(w_n263_40[1]),.dout(n3246),.clk(gclk));
	jand g2984(.dina(w_n1646_0[0]),.dinb(w_shift6_40[1]),.dout(n3247),.clk(gclk));
	jor g2985(.dina(n3247),.dinb(n3246),.dout(result69),.clk(gclk));
	jand g2986(.dina(w_n1755_0[0]),.dinb(w_n263_40[0]),.dout(n3249),.clk(gclk));
	jand g2987(.dina(w_n1719_0[0]),.dinb(w_shift6_40[0]),.dout(n3250),.clk(gclk));
	jor g2988(.dina(n3250),.dinb(n3249),.dout(result70),.clk(gclk));
	jand g2989(.dina(w_n1828_0[0]),.dinb(w_n263_39[2]),.dout(n3252),.clk(gclk));
	jand g2990(.dina(w_n1792_0[0]),.dinb(w_shift6_39[2]),.dout(n3253),.clk(gclk));
	jor g2991(.dina(n3253),.dinb(n3252),.dout(result71),.clk(gclk));
	jand g2992(.dina(w_n1901_0[0]),.dinb(w_n263_39[1]),.dout(n3255),.clk(gclk));
	jand g2993(.dina(w_n1865_0[0]),.dinb(w_shift6_39[1]),.dout(n3256),.clk(gclk));
	jor g2994(.dina(n3256),.dinb(n3255),.dout(result72),.clk(gclk));
	jand g2995(.dina(w_n1974_0[0]),.dinb(w_n263_39[0]),.dout(n3258),.clk(gclk));
	jand g2996(.dina(w_n1938_0[0]),.dinb(w_shift6_39[0]),.dout(n3259),.clk(gclk));
	jor g2997(.dina(n3259),.dinb(n3258),.dout(result73),.clk(gclk));
	jand g2998(.dina(w_n2047_0[0]),.dinb(w_n263_38[2]),.dout(n3261),.clk(gclk));
	jand g2999(.dina(w_n2011_0[0]),.dinb(w_shift6_38[2]),.dout(n3262),.clk(gclk));
	jor g3000(.dina(n3262),.dinb(n3261),.dout(result74),.clk(gclk));
	jand g3001(.dina(w_n2120_0[0]),.dinb(w_n263_38[1]),.dout(n3264),.clk(gclk));
	jand g3002(.dina(w_n2084_0[0]),.dinb(w_shift6_38[1]),.dout(n3265),.clk(gclk));
	jor g3003(.dina(n3265),.dinb(n3264),.dout(result75),.clk(gclk));
	jand g3004(.dina(w_n2193_0[0]),.dinb(w_n263_38[0]),.dout(n3267),.clk(gclk));
	jand g3005(.dina(w_n2157_0[0]),.dinb(w_shift6_38[0]),.dout(n3268),.clk(gclk));
	jor g3006(.dina(n3268),.dinb(n3267),.dout(result76),.clk(gclk));
	jand g3007(.dina(w_n2266_0[0]),.dinb(w_n263_37[2]),.dout(n3270),.clk(gclk));
	jand g3008(.dina(w_n2230_0[0]),.dinb(w_shift6_37[2]),.dout(n3271),.clk(gclk));
	jor g3009(.dina(n3271),.dinb(n3270),.dout(result77),.clk(gclk));
	jand g3010(.dina(w_n2339_0[0]),.dinb(w_n263_37[1]),.dout(n3273),.clk(gclk));
	jand g3011(.dina(w_n2303_0[0]),.dinb(w_shift6_37[1]),.dout(n3274),.clk(gclk));
	jor g3012(.dina(n3274),.dinb(n3273),.dout(result78),.clk(gclk));
	jand g3013(.dina(w_n2412_0[0]),.dinb(w_n263_37[0]),.dout(n3276),.clk(gclk));
	jand g3014(.dina(w_n2376_0[0]),.dinb(w_shift6_37[0]),.dout(n3277),.clk(gclk));
	jor g3015(.dina(n3277),.dinb(n3276),.dout(result79),.clk(gclk));
	jand g3016(.dina(w_n2429_0[0]),.dinb(w_n263_36[2]),.dout(n3279),.clk(gclk));
	jand g3017(.dina(w_n2421_0[0]),.dinb(w_shift6_36[2]),.dout(n3280),.clk(gclk));
	jor g3018(.dina(n3280),.dinb(n3279),.dout(result80),.clk(gclk));
	jand g3019(.dina(w_n2446_0[0]),.dinb(w_n263_36[1]),.dout(n3282),.clk(gclk));
	jand g3020(.dina(w_n2438_0[0]),.dinb(w_shift6_36[1]),.dout(n3283),.clk(gclk));
	jor g3021(.dina(n3283),.dinb(n3282),.dout(result81),.clk(gclk));
	jand g3022(.dina(w_n2463_0[0]),.dinb(w_n263_36[0]),.dout(n3285),.clk(gclk));
	jand g3023(.dina(w_n2455_0[0]),.dinb(w_shift6_36[0]),.dout(n3286),.clk(gclk));
	jor g3024(.dina(n3286),.dinb(n3285),.dout(result82),.clk(gclk));
	jand g3025(.dina(w_n2480_0[0]),.dinb(w_n263_35[2]),.dout(n3288),.clk(gclk));
	jand g3026(.dina(w_n2472_0[0]),.dinb(w_shift6_35[2]),.dout(n3289),.clk(gclk));
	jor g3027(.dina(n3289),.dinb(n3288),.dout(result83),.clk(gclk));
	jand g3028(.dina(w_n2497_0[0]),.dinb(w_n263_35[1]),.dout(n3291),.clk(gclk));
	jand g3029(.dina(w_n2489_0[0]),.dinb(w_shift6_35[1]),.dout(n3292),.clk(gclk));
	jor g3030(.dina(n3292),.dinb(n3291),.dout(result84),.clk(gclk));
	jand g3031(.dina(w_n2514_0[0]),.dinb(w_n263_35[0]),.dout(n3294),.clk(gclk));
	jand g3032(.dina(w_n2506_0[0]),.dinb(w_shift6_35[0]),.dout(n3295),.clk(gclk));
	jor g3033(.dina(n3295),.dinb(n3294),.dout(result85),.clk(gclk));
	jand g3034(.dina(w_n2531_0[0]),.dinb(w_n263_34[2]),.dout(n3297),.clk(gclk));
	jand g3035(.dina(w_n2523_0[0]),.dinb(w_shift6_34[2]),.dout(n3298),.clk(gclk));
	jor g3036(.dina(n3298),.dinb(n3297),.dout(result86),.clk(gclk));
	jand g3037(.dina(w_n2548_0[0]),.dinb(w_n263_34[1]),.dout(n3300),.clk(gclk));
	jand g3038(.dina(w_n2540_0[0]),.dinb(w_shift6_34[1]),.dout(n3301),.clk(gclk));
	jor g3039(.dina(n3301),.dinb(n3300),.dout(result87),.clk(gclk));
	jand g3040(.dina(w_n2565_0[0]),.dinb(w_n263_34[0]),.dout(n3303),.clk(gclk));
	jand g3041(.dina(w_n2557_0[0]),.dinb(w_shift6_34[0]),.dout(n3304),.clk(gclk));
	jor g3042(.dina(n3304),.dinb(n3303),.dout(result88),.clk(gclk));
	jand g3043(.dina(w_n2582_0[0]),.dinb(w_n263_33[2]),.dout(n3306),.clk(gclk));
	jand g3044(.dina(w_n2574_0[0]),.dinb(w_shift6_33[2]),.dout(n3307),.clk(gclk));
	jor g3045(.dina(n3307),.dinb(n3306),.dout(result89),.clk(gclk));
	jand g3046(.dina(w_n2599_0[0]),.dinb(w_n263_33[1]),.dout(n3309),.clk(gclk));
	jand g3047(.dina(w_n2591_0[0]),.dinb(w_shift6_33[1]),.dout(n3310),.clk(gclk));
	jor g3048(.dina(n3310),.dinb(n3309),.dout(result90),.clk(gclk));
	jand g3049(.dina(w_n2616_0[0]),.dinb(w_n263_33[0]),.dout(n3312),.clk(gclk));
	jand g3050(.dina(w_n2608_0[0]),.dinb(w_shift6_33[0]),.dout(n3313),.clk(gclk));
	jor g3051(.dina(n3313),.dinb(n3312),.dout(result91),.clk(gclk));
	jand g3052(.dina(w_n2633_0[0]),.dinb(w_n263_32[2]),.dout(n3315),.clk(gclk));
	jand g3053(.dina(w_n2625_0[0]),.dinb(w_shift6_32[2]),.dout(n3316),.clk(gclk));
	jor g3054(.dina(n3316),.dinb(n3315),.dout(result92),.clk(gclk));
	jand g3055(.dina(w_n2650_0[0]),.dinb(w_n263_32[1]),.dout(n3318),.clk(gclk));
	jand g3056(.dina(w_n2642_0[0]),.dinb(w_shift6_32[1]),.dout(n3319),.clk(gclk));
	jor g3057(.dina(n3319),.dinb(n3318),.dout(result93),.clk(gclk));
	jand g3058(.dina(w_n2667_0[0]),.dinb(w_n263_32[0]),.dout(n3321),.clk(gclk));
	jand g3059(.dina(w_n2659_0[0]),.dinb(w_shift6_32[0]),.dout(n3322),.clk(gclk));
	jor g3060(.dina(n3322),.dinb(n3321),.dout(result94),.clk(gclk));
	jand g3061(.dina(w_n2684_0[0]),.dinb(w_n263_31[2]),.dout(n3324),.clk(gclk));
	jand g3062(.dina(w_n2676_0[0]),.dinb(w_shift6_31[2]),.dout(n3325),.clk(gclk));
	jor g3063(.dina(n3325),.dinb(n3324),.dout(result95),.clk(gclk));
	jand g3064(.dina(w_n2701_0[0]),.dinb(w_n263_31[1]),.dout(n3327),.clk(gclk));
	jand g3065(.dina(w_n2693_0[0]),.dinb(w_shift6_31[1]),.dout(n3328),.clk(gclk));
	jor g3066(.dina(n3328),.dinb(n3327),.dout(result96),.clk(gclk));
	jand g3067(.dina(w_n2718_0[0]),.dinb(w_n263_31[0]),.dout(n3330),.clk(gclk));
	jand g3068(.dina(w_n2710_0[0]),.dinb(w_shift6_31[0]),.dout(n3331),.clk(gclk));
	jor g3069(.dina(n3331),.dinb(n3330),.dout(result97),.clk(gclk));
	jand g3070(.dina(w_n2735_0[0]),.dinb(w_n263_30[2]),.dout(n3333),.clk(gclk));
	jand g3071(.dina(w_n2727_0[0]),.dinb(w_shift6_30[2]),.dout(n3334),.clk(gclk));
	jor g3072(.dina(n3334),.dinb(n3333),.dout(result98),.clk(gclk));
	jand g3073(.dina(w_n2752_0[0]),.dinb(w_n263_30[1]),.dout(n3336),.clk(gclk));
	jand g3074(.dina(w_n2744_0[0]),.dinb(w_shift6_30[1]),.dout(n3337),.clk(gclk));
	jor g3075(.dina(n3337),.dinb(n3336),.dout(result99),.clk(gclk));
	jand g3076(.dina(w_n2769_0[0]),.dinb(w_n263_30[0]),.dout(n3339),.clk(gclk));
	jand g3077(.dina(w_n2761_0[0]),.dinb(w_shift6_30[0]),.dout(n3340),.clk(gclk));
	jor g3078(.dina(n3340),.dinb(n3339),.dout(result100),.clk(gclk));
	jand g3079(.dina(w_n2786_0[0]),.dinb(w_n263_29[2]),.dout(n3342),.clk(gclk));
	jand g3080(.dina(w_n2778_0[0]),.dinb(w_shift6_29[2]),.dout(n3343),.clk(gclk));
	jor g3081(.dina(n3343),.dinb(n3342),.dout(result101),.clk(gclk));
	jand g3082(.dina(w_n2803_0[0]),.dinb(w_n263_29[1]),.dout(n3345),.clk(gclk));
	jand g3083(.dina(w_n2795_0[0]),.dinb(w_shift6_29[1]),.dout(n3346),.clk(gclk));
	jor g3084(.dina(n3346),.dinb(n3345),.dout(result102),.clk(gclk));
	jand g3085(.dina(w_n2820_0[0]),.dinb(w_n263_29[0]),.dout(n3348),.clk(gclk));
	jand g3086(.dina(w_n2812_0[0]),.dinb(w_shift6_29[0]),.dout(n3349),.clk(gclk));
	jor g3087(.dina(n3349),.dinb(n3348),.dout(result103),.clk(gclk));
	jand g3088(.dina(w_n2837_0[0]),.dinb(w_n263_28[2]),.dout(n3351),.clk(gclk));
	jand g3089(.dina(w_n2829_0[0]),.dinb(w_shift6_28[2]),.dout(n3352),.clk(gclk));
	jor g3090(.dina(n3352),.dinb(n3351),.dout(result104),.clk(gclk));
	jand g3091(.dina(w_n2854_0[0]),.dinb(w_n263_28[1]),.dout(n3354),.clk(gclk));
	jand g3092(.dina(w_n2846_0[0]),.dinb(w_shift6_28[1]),.dout(n3355),.clk(gclk));
	jor g3093(.dina(n3355),.dinb(n3354),.dout(result105),.clk(gclk));
	jand g3094(.dina(w_n2871_0[0]),.dinb(w_n263_28[0]),.dout(n3357),.clk(gclk));
	jand g3095(.dina(w_n2863_0[0]),.dinb(w_shift6_28[0]),.dout(n3358),.clk(gclk));
	jor g3096(.dina(n3358),.dinb(n3357),.dout(result106),.clk(gclk));
	jand g3097(.dina(w_n2888_0[0]),.dinb(w_n263_27[2]),.dout(n3360),.clk(gclk));
	jand g3098(.dina(w_n2880_0[0]),.dinb(w_shift6_27[2]),.dout(n3361),.clk(gclk));
	jor g3099(.dina(n3361),.dinb(n3360),.dout(result107),.clk(gclk));
	jand g3100(.dina(w_n2905_0[0]),.dinb(w_n263_27[1]),.dout(n3363),.clk(gclk));
	jand g3101(.dina(w_n2897_0[0]),.dinb(w_shift6_27[1]),.dout(n3364),.clk(gclk));
	jor g3102(.dina(n3364),.dinb(n3363),.dout(result108),.clk(gclk));
	jand g3103(.dina(w_n2922_0[0]),.dinb(w_n263_27[0]),.dout(n3366),.clk(gclk));
	jand g3104(.dina(w_n2914_0[0]),.dinb(w_shift6_27[0]),.dout(n3367),.clk(gclk));
	jor g3105(.dina(n3367),.dinb(n3366),.dout(result109),.clk(gclk));
	jand g3106(.dina(w_n2939_0[0]),.dinb(w_n263_26[2]),.dout(n3369),.clk(gclk));
	jand g3107(.dina(w_n2931_0[0]),.dinb(w_shift6_26[2]),.dout(n3370),.clk(gclk));
	jor g3108(.dina(n3370),.dinb(n3369),.dout(result110),.clk(gclk));
	jand g3109(.dina(w_n2956_0[0]),.dinb(w_n263_26[1]),.dout(n3372),.clk(gclk));
	jand g3110(.dina(w_n2948_0[0]),.dinb(w_shift6_26[1]),.dout(n3373),.clk(gclk));
	jor g3111(.dina(n3373),.dinb(n3372),.dout(result111),.clk(gclk));
	jand g3112(.dina(w_n2973_0[0]),.dinb(w_n263_26[0]),.dout(n3375),.clk(gclk));
	jand g3113(.dina(w_n2965_0[0]),.dinb(w_shift6_26[0]),.dout(n3376),.clk(gclk));
	jor g3114(.dina(n3376),.dinb(n3375),.dout(result112),.clk(gclk));
	jand g3115(.dina(w_n2990_0[0]),.dinb(w_n263_25[2]),.dout(n3378),.clk(gclk));
	jand g3116(.dina(w_n2982_0[0]),.dinb(w_shift6_25[2]),.dout(n3379),.clk(gclk));
	jor g3117(.dina(n3379),.dinb(n3378),.dout(result113),.clk(gclk));
	jand g3118(.dina(w_n3007_0[0]),.dinb(w_n263_25[1]),.dout(n3381),.clk(gclk));
	jand g3119(.dina(w_n2999_0[0]),.dinb(w_shift6_25[1]),.dout(n3382),.clk(gclk));
	jor g3120(.dina(n3382),.dinb(n3381),.dout(result114),.clk(gclk));
	jand g3121(.dina(w_n3024_0[0]),.dinb(w_n263_25[0]),.dout(n3384),.clk(gclk));
	jand g3122(.dina(w_n3016_0[0]),.dinb(w_shift6_25[0]),.dout(n3385),.clk(gclk));
	jor g3123(.dina(n3385),.dinb(n3384),.dout(result115),.clk(gclk));
	jand g3124(.dina(w_n3041_0[0]),.dinb(w_n263_24[2]),.dout(n3387),.clk(gclk));
	jand g3125(.dina(w_n3033_0[0]),.dinb(w_shift6_24[2]),.dout(n3388),.clk(gclk));
	jor g3126(.dina(n3388),.dinb(n3387),.dout(result116),.clk(gclk));
	jand g3127(.dina(w_n3058_0[0]),.dinb(w_n263_24[1]),.dout(n3390),.clk(gclk));
	jand g3128(.dina(w_n3050_0[0]),.dinb(w_shift6_24[1]),.dout(n3391),.clk(gclk));
	jor g3129(.dina(n3391),.dinb(n3390),.dout(result117),.clk(gclk));
	jand g3130(.dina(w_n3075_0[0]),.dinb(w_n263_24[0]),.dout(n3393),.clk(gclk));
	jand g3131(.dina(w_n3067_0[0]),.dinb(w_shift6_24[0]),.dout(n3394),.clk(gclk));
	jor g3132(.dina(n3394),.dinb(n3393),.dout(result118),.clk(gclk));
	jand g3133(.dina(w_n3092_0[0]),.dinb(w_n263_23[2]),.dout(n3396),.clk(gclk));
	jand g3134(.dina(w_n3084_0[0]),.dinb(w_shift6_23[2]),.dout(n3397),.clk(gclk));
	jor g3135(.dina(n3397),.dinb(n3396),.dout(result119),.clk(gclk));
	jand g3136(.dina(w_n3109_0[0]),.dinb(w_n263_23[1]),.dout(n3399),.clk(gclk));
	jand g3137(.dina(w_n3101_0[0]),.dinb(w_shift6_23[1]),.dout(n3400),.clk(gclk));
	jor g3138(.dina(n3400),.dinb(n3399),.dout(result120),.clk(gclk));
	jand g3139(.dina(w_n3126_0[0]),.dinb(w_n263_23[0]),.dout(n3402),.clk(gclk));
	jand g3140(.dina(w_n3118_0[0]),.dinb(w_shift6_23[0]),.dout(n3403),.clk(gclk));
	jor g3141(.dina(n3403),.dinb(n3402),.dout(result121),.clk(gclk));
	jand g3142(.dina(w_n3143_0[0]),.dinb(w_n263_22[2]),.dout(n3405),.clk(gclk));
	jand g3143(.dina(w_n3135_0[0]),.dinb(w_shift6_22[2]),.dout(n3406),.clk(gclk));
	jor g3144(.dina(n3406),.dinb(n3405),.dout(result122),.clk(gclk));
	jand g3145(.dina(w_n3160_0[0]),.dinb(w_n263_22[1]),.dout(n3408),.clk(gclk));
	jand g3146(.dina(w_n3152_0[0]),.dinb(w_shift6_22[1]),.dout(n3409),.clk(gclk));
	jor g3147(.dina(n3409),.dinb(n3408),.dout(result123),.clk(gclk));
	jand g3148(.dina(w_n3177_0[0]),.dinb(w_n263_22[0]),.dout(n3411),.clk(gclk));
	jand g3149(.dina(w_n3169_0[0]),.dinb(w_shift6_22[0]),.dout(n3412),.clk(gclk));
	jor g3150(.dina(n3412),.dinb(n3411),.dout(result124),.clk(gclk));
	jand g3151(.dina(w_n3194_0[0]),.dinb(w_n263_21[2]),.dout(n3414),.clk(gclk));
	jand g3152(.dina(w_n3186_0[0]),.dinb(w_shift6_21[2]),.dout(n3415),.clk(gclk));
	jor g3153(.dina(n3415),.dinb(n3414),.dout(result125),.clk(gclk));
	jand g3154(.dina(w_n3211_0[0]),.dinb(w_n263_21[1]),.dout(n3417),.clk(gclk));
	jand g3155(.dina(w_n3203_0[0]),.dinb(w_shift6_21[1]),.dout(n3418),.clk(gclk));
	jor g3156(.dina(n3418),.dinb(n3417),.dout(result126),.clk(gclk));
	jand g3157(.dina(w_n3228_0[0]),.dinb(w_n263_21[0]),.dout(n3420),.clk(gclk));
	jand g3158(.dina(w_n3220_0[0]),.dinb(w_shift6_21[0]),.dout(n3421),.clk(gclk));
	jor g3159(.dina(n3421),.dinb(n3420),.dout(result127),.clk(gclk));
	jspl jspl_w_a0_0(.douta(w_a0_0[0]),.doutb(w_a0_0[1]),.din(a0));
	jspl jspl_w_a1_0(.douta(w_a1_0[0]),.doutb(w_a1_0[1]),.din(a1));
	jspl jspl_w_a2_0(.douta(w_a2_0[0]),.doutb(w_a2_0[1]),.din(a2));
	jspl jspl_w_a3_0(.douta(w_a3_0[0]),.doutb(w_a3_0[1]),.din(a3));
	jspl jspl_w_a4_0(.douta(w_a4_0[0]),.doutb(w_a4_0[1]),.din(a4));
	jspl jspl_w_a5_0(.douta(w_a5_0[0]),.doutb(w_a5_0[1]),.din(a5));
	jspl jspl_w_a6_0(.douta(w_a6_0[0]),.doutb(w_a6_0[1]),.din(a6));
	jspl jspl_w_a7_0(.douta(w_a7_0[0]),.doutb(w_a7_0[1]),.din(a7));
	jspl jspl_w_a8_0(.douta(w_a8_0[0]),.doutb(w_a8_0[1]),.din(a8));
	jspl jspl_w_a9_0(.douta(w_a9_0[0]),.doutb(w_a9_0[1]),.din(a9));
	jspl jspl_w_a10_0(.douta(w_a10_0[0]),.doutb(w_a10_0[1]),.din(a10));
	jspl jspl_w_a11_0(.douta(w_a11_0[0]),.doutb(w_a11_0[1]),.din(a11));
	jspl jspl_w_a12_0(.douta(w_a12_0[0]),.doutb(w_a12_0[1]),.din(a12));
	jspl jspl_w_a13_0(.douta(w_a13_0[0]),.doutb(w_a13_0[1]),.din(a13));
	jspl jspl_w_a14_0(.douta(w_a14_0[0]),.doutb(w_a14_0[1]),.din(a14));
	jspl jspl_w_a15_0(.douta(w_a15_0[0]),.doutb(w_a15_0[1]),.din(a15));
	jspl jspl_w_a16_0(.douta(w_a16_0[0]),.doutb(w_a16_0[1]),.din(a16));
	jspl jspl_w_a17_0(.douta(w_a17_0[0]),.doutb(w_a17_0[1]),.din(a17));
	jspl jspl_w_a18_0(.douta(w_a18_0[0]),.doutb(w_a18_0[1]),.din(a18));
	jspl jspl_w_a19_0(.douta(w_a19_0[0]),.doutb(w_a19_0[1]),.din(a19));
	jspl jspl_w_a20_0(.douta(w_a20_0[0]),.doutb(w_a20_0[1]),.din(a20));
	jspl jspl_w_a21_0(.douta(w_a21_0[0]),.doutb(w_a21_0[1]),.din(a21));
	jspl jspl_w_a22_0(.douta(w_a22_0[0]),.doutb(w_a22_0[1]),.din(a22));
	jspl jspl_w_a23_0(.douta(w_a23_0[0]),.doutb(w_a23_0[1]),.din(a23));
	jspl jspl_w_a24_0(.douta(w_a24_0[0]),.doutb(w_a24_0[1]),.din(a24));
	jspl jspl_w_a25_0(.douta(w_a25_0[0]),.doutb(w_a25_0[1]),.din(a25));
	jspl jspl_w_a26_0(.douta(w_a26_0[0]),.doutb(w_a26_0[1]),.din(a26));
	jspl jspl_w_a27_0(.douta(w_a27_0[0]),.doutb(w_a27_0[1]),.din(a27));
	jspl jspl_w_a28_0(.douta(w_a28_0[0]),.doutb(w_a28_0[1]),.din(a28));
	jspl jspl_w_a29_0(.douta(w_a29_0[0]),.doutb(w_a29_0[1]),.din(a29));
	jspl jspl_w_a30_0(.douta(w_a30_0[0]),.doutb(w_a30_0[1]),.din(a30));
	jspl jspl_w_a31_0(.douta(w_a31_0[0]),.doutb(w_a31_0[1]),.din(a31));
	jspl jspl_w_a32_0(.douta(w_a32_0[0]),.doutb(w_a32_0[1]),.din(a32));
	jspl jspl_w_a33_0(.douta(w_a33_0[0]),.doutb(w_a33_0[1]),.din(a33));
	jspl jspl_w_a34_0(.douta(w_a34_0[0]),.doutb(w_a34_0[1]),.din(a34));
	jspl jspl_w_a35_0(.douta(w_a35_0[0]),.doutb(w_a35_0[1]),.din(a35));
	jspl jspl_w_a36_0(.douta(w_a36_0[0]),.doutb(w_a36_0[1]),.din(a36));
	jspl jspl_w_a37_0(.douta(w_a37_0[0]),.doutb(w_a37_0[1]),.din(a37));
	jspl jspl_w_a38_0(.douta(w_a38_0[0]),.doutb(w_a38_0[1]),.din(a38));
	jspl jspl_w_a39_0(.douta(w_a39_0[0]),.doutb(w_a39_0[1]),.din(a39));
	jspl jspl_w_a40_0(.douta(w_a40_0[0]),.doutb(w_a40_0[1]),.din(a40));
	jspl jspl_w_a41_0(.douta(w_a41_0[0]),.doutb(w_a41_0[1]),.din(a41));
	jspl jspl_w_a42_0(.douta(w_a42_0[0]),.doutb(w_a42_0[1]),.din(a42));
	jspl jspl_w_a43_0(.douta(w_a43_0[0]),.doutb(w_a43_0[1]),.din(a43));
	jspl jspl_w_a44_0(.douta(w_a44_0[0]),.doutb(w_a44_0[1]),.din(a44));
	jspl jspl_w_a45_0(.douta(w_a45_0[0]),.doutb(w_a45_0[1]),.din(a45));
	jspl jspl_w_a46_0(.douta(w_a46_0[0]),.doutb(w_a46_0[1]),.din(a46));
	jspl jspl_w_a47_0(.douta(w_a47_0[0]),.doutb(w_a47_0[1]),.din(a47));
	jspl jspl_w_a48_0(.douta(w_a48_0[0]),.doutb(w_a48_0[1]),.din(a48));
	jspl jspl_w_a49_0(.douta(w_a49_0[0]),.doutb(w_a49_0[1]),.din(a49));
	jspl jspl_w_a50_0(.douta(w_a50_0[0]),.doutb(w_a50_0[1]),.din(a50));
	jspl jspl_w_a51_0(.douta(w_a51_0[0]),.doutb(w_a51_0[1]),.din(a51));
	jspl jspl_w_a52_0(.douta(w_a52_0[0]),.doutb(w_a52_0[1]),.din(a52));
	jspl jspl_w_a53_0(.douta(w_a53_0[0]),.doutb(w_a53_0[1]),.din(a53));
	jspl jspl_w_a54_0(.douta(w_a54_0[0]),.doutb(w_a54_0[1]),.din(a54));
	jspl jspl_w_a55_0(.douta(w_a55_0[0]),.doutb(w_a55_0[1]),.din(a55));
	jspl jspl_w_a56_0(.douta(w_a56_0[0]),.doutb(w_a56_0[1]),.din(a56));
	jspl jspl_w_a57_0(.douta(w_a57_0[0]),.doutb(w_a57_0[1]),.din(a57));
	jspl jspl_w_a58_0(.douta(w_a58_0[0]),.doutb(w_a58_0[1]),.din(a58));
	jspl jspl_w_a59_0(.douta(w_a59_0[0]),.doutb(w_a59_0[1]),.din(a59));
	jspl jspl_w_a60_0(.douta(w_a60_0[0]),.doutb(w_a60_0[1]),.din(a60));
	jspl jspl_w_a61_0(.douta(w_a61_0[0]),.doutb(w_a61_0[1]),.din(a61));
	jspl jspl_w_a62_0(.douta(w_a62_0[0]),.doutb(w_a62_0[1]),.din(a62));
	jspl jspl_w_a63_0(.douta(w_a63_0[0]),.doutb(w_a63_0[1]),.din(a63));
	jspl jspl_w_a64_0(.douta(w_a64_0[0]),.doutb(w_a64_0[1]),.din(a64));
	jspl jspl_w_a65_0(.douta(w_a65_0[0]),.doutb(w_a65_0[1]),.din(a65));
	jspl jspl_w_a66_0(.douta(w_a66_0[0]),.doutb(w_a66_0[1]),.din(a66));
	jspl jspl_w_a67_0(.douta(w_a67_0[0]),.doutb(w_a67_0[1]),.din(a67));
	jspl jspl_w_a68_0(.douta(w_a68_0[0]),.doutb(w_a68_0[1]),.din(a68));
	jspl jspl_w_a69_0(.douta(w_a69_0[0]),.doutb(w_a69_0[1]),.din(a69));
	jspl jspl_w_a70_0(.douta(w_a70_0[0]),.doutb(w_a70_0[1]),.din(a70));
	jspl jspl_w_a71_0(.douta(w_a71_0[0]),.doutb(w_a71_0[1]),.din(a71));
	jspl jspl_w_a72_0(.douta(w_a72_0[0]),.doutb(w_a72_0[1]),.din(a72));
	jspl jspl_w_a73_0(.douta(w_a73_0[0]),.doutb(w_a73_0[1]),.din(a73));
	jspl jspl_w_a74_0(.douta(w_a74_0[0]),.doutb(w_a74_0[1]),.din(a74));
	jspl jspl_w_a75_0(.douta(w_a75_0[0]),.doutb(w_a75_0[1]),.din(a75));
	jspl jspl_w_a76_0(.douta(w_a76_0[0]),.doutb(w_a76_0[1]),.din(a76));
	jspl jspl_w_a77_0(.douta(w_a77_0[0]),.doutb(w_a77_0[1]),.din(a77));
	jspl jspl_w_a78_0(.douta(w_a78_0[0]),.doutb(w_a78_0[1]),.din(a78));
	jspl jspl_w_a79_0(.douta(w_a79_0[0]),.doutb(w_a79_0[1]),.din(a79));
	jspl jspl_w_a80_0(.douta(w_a80_0[0]),.doutb(w_a80_0[1]),.din(a80));
	jspl jspl_w_a81_0(.douta(w_a81_0[0]),.doutb(w_a81_0[1]),.din(a81));
	jspl jspl_w_a82_0(.douta(w_a82_0[0]),.doutb(w_a82_0[1]),.din(a82));
	jspl jspl_w_a83_0(.douta(w_a83_0[0]),.doutb(w_a83_0[1]),.din(a83));
	jspl jspl_w_a84_0(.douta(w_a84_0[0]),.doutb(w_a84_0[1]),.din(a84));
	jspl jspl_w_a85_0(.douta(w_a85_0[0]),.doutb(w_a85_0[1]),.din(a85));
	jspl jspl_w_a86_0(.douta(w_a86_0[0]),.doutb(w_a86_0[1]),.din(a86));
	jspl jspl_w_a87_0(.douta(w_a87_0[0]),.doutb(w_a87_0[1]),.din(a87));
	jspl jspl_w_a88_0(.douta(w_a88_0[0]),.doutb(w_a88_0[1]),.din(a88));
	jspl jspl_w_a89_0(.douta(w_a89_0[0]),.doutb(w_a89_0[1]),.din(a89));
	jspl jspl_w_a90_0(.douta(w_a90_0[0]),.doutb(w_a90_0[1]),.din(a90));
	jspl jspl_w_a91_0(.douta(w_a91_0[0]),.doutb(w_a91_0[1]),.din(a91));
	jspl jspl_w_a92_0(.douta(w_a92_0[0]),.doutb(w_a92_0[1]),.din(a92));
	jspl jspl_w_a93_0(.douta(w_a93_0[0]),.doutb(w_a93_0[1]),.din(a93));
	jspl jspl_w_a94_0(.douta(w_a94_0[0]),.doutb(w_a94_0[1]),.din(a94));
	jspl jspl_w_a95_0(.douta(w_a95_0[0]),.doutb(w_a95_0[1]),.din(a95));
	jspl jspl_w_a96_0(.douta(w_a96_0[0]),.doutb(w_a96_0[1]),.din(a96));
	jspl jspl_w_a97_0(.douta(w_a97_0[0]),.doutb(w_a97_0[1]),.din(a97));
	jspl jspl_w_a98_0(.douta(w_a98_0[0]),.doutb(w_a98_0[1]),.din(a98));
	jspl jspl_w_a99_0(.douta(w_a99_0[0]),.doutb(w_a99_0[1]),.din(a99));
	jspl jspl_w_a100_0(.douta(w_a100_0[0]),.doutb(w_a100_0[1]),.din(a100));
	jspl jspl_w_a101_0(.douta(w_a101_0[0]),.doutb(w_a101_0[1]),.din(a101));
	jspl jspl_w_a102_0(.douta(w_a102_0[0]),.doutb(w_a102_0[1]),.din(a102));
	jspl jspl_w_a103_0(.douta(w_a103_0[0]),.doutb(w_a103_0[1]),.din(a103));
	jspl jspl_w_a104_0(.douta(w_a104_0[0]),.doutb(w_a104_0[1]),.din(a104));
	jspl jspl_w_a105_0(.douta(w_a105_0[0]),.doutb(w_a105_0[1]),.din(a105));
	jspl jspl_w_a106_0(.douta(w_a106_0[0]),.doutb(w_a106_0[1]),.din(a106));
	jspl jspl_w_a107_0(.douta(w_a107_0[0]),.doutb(w_a107_0[1]),.din(a107));
	jspl jspl_w_a108_0(.douta(w_a108_0[0]),.doutb(w_a108_0[1]),.din(a108));
	jspl jspl_w_a109_0(.douta(w_a109_0[0]),.doutb(w_a109_0[1]),.din(a109));
	jspl jspl_w_a110_0(.douta(w_a110_0[0]),.doutb(w_a110_0[1]),.din(a110));
	jspl jspl_w_a111_0(.douta(w_a111_0[0]),.doutb(w_a111_0[1]),.din(a111));
	jspl jspl_w_a112_0(.douta(w_a112_0[0]),.doutb(w_a112_0[1]),.din(a112));
	jspl jspl_w_a113_0(.douta(w_a113_0[0]),.doutb(w_a113_0[1]),.din(a113));
	jspl jspl_w_a114_0(.douta(w_a114_0[0]),.doutb(w_a114_0[1]),.din(a114));
	jspl jspl_w_a115_0(.douta(w_a115_0[0]),.doutb(w_a115_0[1]),.din(a115));
	jspl jspl_w_a116_0(.douta(w_a116_0[0]),.doutb(w_a116_0[1]),.din(a116));
	jspl jspl_w_a117_0(.douta(w_a117_0[0]),.doutb(w_a117_0[1]),.din(a117));
	jspl jspl_w_a118_0(.douta(w_a118_0[0]),.doutb(w_a118_0[1]),.din(a118));
	jspl jspl_w_a119_0(.douta(w_a119_0[0]),.doutb(w_a119_0[1]),.din(a119));
	jspl jspl_w_a120_0(.douta(w_a120_0[0]),.doutb(w_a120_0[1]),.din(a120));
	jspl jspl_w_a121_0(.douta(w_a121_0[0]),.doutb(w_a121_0[1]),.din(a121));
	jspl jspl_w_a122_0(.douta(w_a122_0[0]),.doutb(w_a122_0[1]),.din(a122));
	jspl jspl_w_a123_0(.douta(w_a123_0[0]),.doutb(w_a123_0[1]),.din(a123));
	jspl jspl_w_a124_0(.douta(w_a124_0[0]),.doutb(w_a124_0[1]),.din(a124));
	jspl jspl_w_a125_0(.douta(w_a125_0[0]),.doutb(w_a125_0[1]),.din(a125));
	jspl jspl_w_a126_0(.douta(w_a126_0[0]),.doutb(w_a126_0[1]),.din(a126));
	jspl jspl_w_a127_0(.douta(w_a127_0[0]),.doutb(w_a127_0[1]),.din(a127));
	jspl3 jspl3_w_shift0_0(.douta(w_shift0_0[0]),.doutb(w_shift0_0[1]),.doutc(w_shift0_0[2]),.din(shift0));
	jspl3 jspl3_w_shift0_1(.douta(w_shift0_1[0]),.doutb(w_shift0_1[1]),.doutc(w_shift0_1[2]),.din(w_shift0_0[0]));
	jspl3 jspl3_w_shift0_2(.douta(w_shift0_2[0]),.doutb(w_shift0_2[1]),.doutc(w_shift0_2[2]),.din(w_shift0_0[1]));
	jspl3 jspl3_w_shift0_3(.douta(w_shift0_3[0]),.doutb(w_shift0_3[1]),.doutc(w_shift0_3[2]),.din(w_shift0_0[2]));
	jspl3 jspl3_w_shift0_4(.douta(w_shift0_4[0]),.doutb(w_shift0_4[1]),.doutc(w_shift0_4[2]),.din(w_shift0_1[0]));
	jspl3 jspl3_w_shift0_5(.douta(w_shift0_5[0]),.doutb(w_shift0_5[1]),.doutc(w_shift0_5[2]),.din(w_shift0_1[1]));
	jspl3 jspl3_w_shift0_6(.douta(w_shift0_6[0]),.doutb(w_shift0_6[1]),.doutc(w_shift0_6[2]),.din(w_shift0_1[2]));
	jspl3 jspl3_w_shift0_7(.douta(w_shift0_7[0]),.doutb(w_shift0_7[1]),.doutc(w_shift0_7[2]),.din(w_shift0_2[0]));
	jspl3 jspl3_w_shift0_8(.douta(w_shift0_8[0]),.doutb(w_shift0_8[1]),.doutc(w_shift0_8[2]),.din(w_shift0_2[1]));
	jspl3 jspl3_w_shift0_9(.douta(w_shift0_9[0]),.doutb(w_shift0_9[1]),.doutc(w_shift0_9[2]),.din(w_shift0_2[2]));
	jspl3 jspl3_w_shift0_10(.douta(w_shift0_10[0]),.doutb(w_shift0_10[1]),.doutc(w_shift0_10[2]),.din(w_shift0_3[0]));
	jspl3 jspl3_w_shift0_11(.douta(w_shift0_11[0]),.doutb(w_shift0_11[1]),.doutc(w_shift0_11[2]),.din(w_shift0_3[1]));
	jspl3 jspl3_w_shift0_12(.douta(w_shift0_12[0]),.doutb(w_shift0_12[1]),.doutc(w_shift0_12[2]),.din(w_shift0_3[2]));
	jspl3 jspl3_w_shift0_13(.douta(w_shift0_13[0]),.doutb(w_shift0_13[1]),.doutc(w_shift0_13[2]),.din(w_shift0_4[0]));
	jspl3 jspl3_w_shift0_14(.douta(w_shift0_14[0]),.doutb(w_shift0_14[1]),.doutc(w_shift0_14[2]),.din(w_shift0_4[1]));
	jspl3 jspl3_w_shift0_15(.douta(w_shift0_15[0]),.doutb(w_shift0_15[1]),.doutc(w_shift0_15[2]),.din(w_shift0_4[2]));
	jspl3 jspl3_w_shift0_16(.douta(w_shift0_16[0]),.doutb(w_shift0_16[1]),.doutc(w_shift0_16[2]),.din(w_shift0_5[0]));
	jspl3 jspl3_w_shift0_17(.douta(w_shift0_17[0]),.doutb(w_shift0_17[1]),.doutc(w_shift0_17[2]),.din(w_shift0_5[1]));
	jspl3 jspl3_w_shift0_18(.douta(w_shift0_18[0]),.doutb(w_shift0_18[1]),.doutc(w_shift0_18[2]),.din(w_shift0_5[2]));
	jspl3 jspl3_w_shift0_19(.douta(w_shift0_19[0]),.doutb(w_shift0_19[1]),.doutc(w_shift0_19[2]),.din(w_shift0_6[0]));
	jspl3 jspl3_w_shift0_20(.douta(w_shift0_20[0]),.doutb(w_shift0_20[1]),.doutc(w_shift0_20[2]),.din(w_shift0_6[1]));
	jspl3 jspl3_w_shift0_21(.douta(w_shift0_21[0]),.doutb(w_shift0_21[1]),.doutc(w_shift0_21[2]),.din(w_shift0_6[2]));
	jspl3 jspl3_w_shift0_22(.douta(w_shift0_22[0]),.doutb(w_shift0_22[1]),.doutc(w_shift0_22[2]),.din(w_shift0_7[0]));
	jspl3 jspl3_w_shift0_23(.douta(w_shift0_23[0]),.doutb(w_shift0_23[1]),.doutc(w_shift0_23[2]),.din(w_shift0_7[1]));
	jspl3 jspl3_w_shift0_24(.douta(w_shift0_24[0]),.doutb(w_shift0_24[1]),.doutc(w_shift0_24[2]),.din(w_shift0_7[2]));
	jspl3 jspl3_w_shift0_25(.douta(w_shift0_25[0]),.doutb(w_shift0_25[1]),.doutc(w_shift0_25[2]),.din(w_shift0_8[0]));
	jspl3 jspl3_w_shift0_26(.douta(w_shift0_26[0]),.doutb(w_shift0_26[1]),.doutc(w_shift0_26[2]),.din(w_shift0_8[1]));
	jspl3 jspl3_w_shift0_27(.douta(w_shift0_27[0]),.doutb(w_shift0_27[1]),.doutc(w_shift0_27[2]),.din(w_shift0_8[2]));
	jspl3 jspl3_w_shift0_28(.douta(w_shift0_28[0]),.doutb(w_shift0_28[1]),.doutc(w_shift0_28[2]),.din(w_shift0_9[0]));
	jspl3 jspl3_w_shift0_29(.douta(w_shift0_29[0]),.doutb(w_shift0_29[1]),.doutc(w_shift0_29[2]),.din(w_shift0_9[1]));
	jspl3 jspl3_w_shift0_30(.douta(w_shift0_30[0]),.doutb(w_shift0_30[1]),.doutc(w_shift0_30[2]),.din(w_shift0_9[2]));
	jspl3 jspl3_w_shift0_31(.douta(w_shift0_31[0]),.doutb(w_shift0_31[1]),.doutc(w_shift0_31[2]),.din(w_shift0_10[0]));
	jspl3 jspl3_w_shift0_32(.douta(w_shift0_32[0]),.doutb(w_shift0_32[1]),.doutc(w_shift0_32[2]),.din(w_shift0_10[1]));
	jspl3 jspl3_w_shift0_33(.douta(w_shift0_33[0]),.doutb(w_shift0_33[1]),.doutc(w_shift0_33[2]),.din(w_shift0_10[2]));
	jspl3 jspl3_w_shift0_34(.douta(w_shift0_34[0]),.doutb(w_shift0_34[1]),.doutc(w_shift0_34[2]),.din(w_shift0_11[0]));
	jspl3 jspl3_w_shift0_35(.douta(w_shift0_35[0]),.doutb(w_shift0_35[1]),.doutc(w_shift0_35[2]),.din(w_shift0_11[1]));
	jspl3 jspl3_w_shift0_36(.douta(w_shift0_36[0]),.doutb(w_shift0_36[1]),.doutc(w_shift0_36[2]),.din(w_shift0_11[2]));
	jspl3 jspl3_w_shift0_37(.douta(w_shift0_37[0]),.doutb(w_shift0_37[1]),.doutc(w_shift0_37[2]),.din(w_shift0_12[0]));
	jspl3 jspl3_w_shift0_38(.douta(w_shift0_38[0]),.doutb(w_shift0_38[1]),.doutc(w_shift0_38[2]),.din(w_shift0_12[1]));
	jspl3 jspl3_w_shift0_39(.douta(w_shift0_39[0]),.doutb(w_shift0_39[1]),.doutc(w_shift0_39[2]),.din(w_shift0_12[2]));
	jspl3 jspl3_w_shift0_40(.douta(w_shift0_40[0]),.doutb(w_shift0_40[1]),.doutc(w_shift0_40[2]),.din(w_shift0_13[0]));
	jspl3 jspl3_w_shift0_41(.douta(w_shift0_41[0]),.doutb(w_shift0_41[1]),.doutc(w_shift0_41[2]),.din(w_shift0_13[1]));
	jspl3 jspl3_w_shift0_42(.douta(w_shift0_42[0]),.doutb(w_shift0_42[1]),.doutc(w_shift0_42[2]),.din(w_shift0_13[2]));
	jspl3 jspl3_w_shift0_43(.douta(w_shift0_43[0]),.doutb(w_shift0_43[1]),.doutc(w_shift0_43[2]),.din(w_shift0_14[0]));
	jspl3 jspl3_w_shift0_44(.douta(w_shift0_44[0]),.doutb(w_shift0_44[1]),.doutc(w_shift0_44[2]),.din(w_shift0_14[1]));
	jspl3 jspl3_w_shift0_45(.douta(w_shift0_45[0]),.doutb(w_shift0_45[1]),.doutc(w_shift0_45[2]),.din(w_shift0_14[2]));
	jspl3 jspl3_w_shift0_46(.douta(w_shift0_46[0]),.doutb(w_shift0_46[1]),.doutc(w_shift0_46[2]),.din(w_shift0_15[0]));
	jspl3 jspl3_w_shift0_47(.douta(w_shift0_47[0]),.doutb(w_shift0_47[1]),.doutc(w_shift0_47[2]),.din(w_shift0_15[1]));
	jspl3 jspl3_w_shift0_48(.douta(w_shift0_48[0]),.doutb(w_shift0_48[1]),.doutc(w_shift0_48[2]),.din(w_shift0_15[2]));
	jspl3 jspl3_w_shift0_49(.douta(w_shift0_49[0]),.doutb(w_shift0_49[1]),.doutc(w_shift0_49[2]),.din(w_shift0_16[0]));
	jspl3 jspl3_w_shift0_50(.douta(w_shift0_50[0]),.doutb(w_shift0_50[1]),.doutc(w_shift0_50[2]),.din(w_shift0_16[1]));
	jspl3 jspl3_w_shift0_51(.douta(w_shift0_51[0]),.doutb(w_shift0_51[1]),.doutc(w_shift0_51[2]),.din(w_shift0_16[2]));
	jspl3 jspl3_w_shift0_52(.douta(w_shift0_52[0]),.doutb(w_shift0_52[1]),.doutc(w_shift0_52[2]),.din(w_shift0_17[0]));
	jspl3 jspl3_w_shift0_53(.douta(w_shift0_53[0]),.doutb(w_shift0_53[1]),.doutc(w_shift0_53[2]),.din(w_shift0_17[1]));
	jspl3 jspl3_w_shift0_54(.douta(w_shift0_54[0]),.doutb(w_shift0_54[1]),.doutc(w_shift0_54[2]),.din(w_shift0_17[2]));
	jspl3 jspl3_w_shift0_55(.douta(w_shift0_55[0]),.doutb(w_shift0_55[1]),.doutc(w_shift0_55[2]),.din(w_shift0_18[0]));
	jspl3 jspl3_w_shift0_56(.douta(w_shift0_56[0]),.doutb(w_shift0_56[1]),.doutc(w_shift0_56[2]),.din(w_shift0_18[1]));
	jspl3 jspl3_w_shift0_57(.douta(w_shift0_57[0]),.doutb(w_shift0_57[1]),.doutc(w_shift0_57[2]),.din(w_shift0_18[2]));
	jspl3 jspl3_w_shift0_58(.douta(w_shift0_58[0]),.doutb(w_shift0_58[1]),.doutc(w_shift0_58[2]),.din(w_shift0_19[0]));
	jspl3 jspl3_w_shift0_59(.douta(w_shift0_59[0]),.doutb(w_shift0_59[1]),.doutc(w_shift0_59[2]),.din(w_shift0_19[1]));
	jspl3 jspl3_w_shift0_60(.douta(w_shift0_60[0]),.doutb(w_shift0_60[1]),.doutc(w_shift0_60[2]),.din(w_shift0_19[2]));
	jspl3 jspl3_w_shift0_61(.douta(w_shift0_61[0]),.doutb(w_shift0_61[1]),.doutc(w_shift0_61[2]),.din(w_shift0_20[0]));
	jspl3 jspl3_w_shift0_62(.douta(w_shift0_62[0]),.doutb(w_shift0_62[1]),.doutc(w_shift0_62[2]),.din(w_shift0_20[1]));
	jspl3 jspl3_w_shift0_63(.douta(w_shift0_63[0]),.doutb(w_shift0_63[1]),.doutc(w_shift0_63[2]),.din(w_shift0_20[2]));
	jspl3 jspl3_w_shift1_0(.douta(w_shift1_0[0]),.doutb(w_shift1_0[1]),.doutc(w_shift1_0[2]),.din(shift1));
	jspl3 jspl3_w_shift1_1(.douta(w_shift1_1[0]),.doutb(w_shift1_1[1]),.doutc(w_shift1_1[2]),.din(w_shift1_0[0]));
	jspl3 jspl3_w_shift1_2(.douta(w_shift1_2[0]),.doutb(w_shift1_2[1]),.doutc(w_shift1_2[2]),.din(w_shift1_0[1]));
	jspl3 jspl3_w_shift1_3(.douta(w_shift1_3[0]),.doutb(w_shift1_3[1]),.doutc(w_shift1_3[2]),.din(w_shift1_0[2]));
	jspl3 jspl3_w_shift1_4(.douta(w_shift1_4[0]),.doutb(w_shift1_4[1]),.doutc(w_shift1_4[2]),.din(w_shift1_1[0]));
	jspl3 jspl3_w_shift1_5(.douta(w_shift1_5[0]),.doutb(w_shift1_5[1]),.doutc(w_shift1_5[2]),.din(w_shift1_1[1]));
	jspl3 jspl3_w_shift1_6(.douta(w_shift1_6[0]),.doutb(w_shift1_6[1]),.doutc(w_shift1_6[2]),.din(w_shift1_1[2]));
	jspl3 jspl3_w_shift1_7(.douta(w_shift1_7[0]),.doutb(w_shift1_7[1]),.doutc(w_shift1_7[2]),.din(w_shift1_2[0]));
	jspl3 jspl3_w_shift1_8(.douta(w_shift1_8[0]),.doutb(w_shift1_8[1]),.doutc(w_shift1_8[2]),.din(w_shift1_2[1]));
	jspl3 jspl3_w_shift1_9(.douta(w_shift1_9[0]),.doutb(w_shift1_9[1]),.doutc(w_shift1_9[2]),.din(w_shift1_2[2]));
	jspl3 jspl3_w_shift1_10(.douta(w_shift1_10[0]),.doutb(w_shift1_10[1]),.doutc(w_shift1_10[2]),.din(w_shift1_3[0]));
	jspl3 jspl3_w_shift1_11(.douta(w_shift1_11[0]),.doutb(w_shift1_11[1]),.doutc(w_shift1_11[2]),.din(w_shift1_3[1]));
	jspl3 jspl3_w_shift1_12(.douta(w_shift1_12[0]),.doutb(w_shift1_12[1]),.doutc(w_shift1_12[2]),.din(w_shift1_3[2]));
	jspl3 jspl3_w_shift1_13(.douta(w_shift1_13[0]),.doutb(w_shift1_13[1]),.doutc(w_shift1_13[2]),.din(w_shift1_4[0]));
	jspl3 jspl3_w_shift1_14(.douta(w_shift1_14[0]),.doutb(w_shift1_14[1]),.doutc(w_shift1_14[2]),.din(w_shift1_4[1]));
	jspl3 jspl3_w_shift1_15(.douta(w_shift1_15[0]),.doutb(w_shift1_15[1]),.doutc(w_shift1_15[2]),.din(w_shift1_4[2]));
	jspl3 jspl3_w_shift1_16(.douta(w_shift1_16[0]),.doutb(w_shift1_16[1]),.doutc(w_shift1_16[2]),.din(w_shift1_5[0]));
	jspl3 jspl3_w_shift1_17(.douta(w_shift1_17[0]),.doutb(w_shift1_17[1]),.doutc(w_shift1_17[2]),.din(w_shift1_5[1]));
	jspl3 jspl3_w_shift1_18(.douta(w_shift1_18[0]),.doutb(w_shift1_18[1]),.doutc(w_shift1_18[2]),.din(w_shift1_5[2]));
	jspl3 jspl3_w_shift1_19(.douta(w_shift1_19[0]),.doutb(w_shift1_19[1]),.doutc(w_shift1_19[2]),.din(w_shift1_6[0]));
	jspl3 jspl3_w_shift1_20(.douta(w_shift1_20[0]),.doutb(w_shift1_20[1]),.doutc(w_shift1_20[2]),.din(w_shift1_6[1]));
	jspl3 jspl3_w_shift1_21(.douta(w_shift1_21[0]),.doutb(w_shift1_21[1]),.doutc(w_shift1_21[2]),.din(w_shift1_6[2]));
	jspl3 jspl3_w_shift1_22(.douta(w_shift1_22[0]),.doutb(w_shift1_22[1]),.doutc(w_shift1_22[2]),.din(w_shift1_7[0]));
	jspl3 jspl3_w_shift1_23(.douta(w_shift1_23[0]),.doutb(w_shift1_23[1]),.doutc(w_shift1_23[2]),.din(w_shift1_7[1]));
	jspl3 jspl3_w_shift1_24(.douta(w_shift1_24[0]),.doutb(w_shift1_24[1]),.doutc(w_shift1_24[2]),.din(w_shift1_7[2]));
	jspl3 jspl3_w_shift1_25(.douta(w_shift1_25[0]),.doutb(w_shift1_25[1]),.doutc(w_shift1_25[2]),.din(w_shift1_8[0]));
	jspl3 jspl3_w_shift1_26(.douta(w_shift1_26[0]),.doutb(w_shift1_26[1]),.doutc(w_shift1_26[2]),.din(w_shift1_8[1]));
	jspl3 jspl3_w_shift1_27(.douta(w_shift1_27[0]),.doutb(w_shift1_27[1]),.doutc(w_shift1_27[2]),.din(w_shift1_8[2]));
	jspl3 jspl3_w_shift1_28(.douta(w_shift1_28[0]),.doutb(w_shift1_28[1]),.doutc(w_shift1_28[2]),.din(w_shift1_9[0]));
	jspl3 jspl3_w_shift1_29(.douta(w_shift1_29[0]),.doutb(w_shift1_29[1]),.doutc(w_shift1_29[2]),.din(w_shift1_9[1]));
	jspl3 jspl3_w_shift1_30(.douta(w_shift1_30[0]),.doutb(w_shift1_30[1]),.doutc(w_shift1_30[2]),.din(w_shift1_9[2]));
	jspl3 jspl3_w_shift1_31(.douta(w_shift1_31[0]),.doutb(w_shift1_31[1]),.doutc(w_shift1_31[2]),.din(w_shift1_10[0]));
	jspl3 jspl3_w_shift1_32(.douta(w_shift1_32[0]),.doutb(w_shift1_32[1]),.doutc(w_shift1_32[2]),.din(w_shift1_10[1]));
	jspl3 jspl3_w_shift1_33(.douta(w_shift1_33[0]),.doutb(w_shift1_33[1]),.doutc(w_shift1_33[2]),.din(w_shift1_10[2]));
	jspl3 jspl3_w_shift1_34(.douta(w_shift1_34[0]),.doutb(w_shift1_34[1]),.doutc(w_shift1_34[2]),.din(w_shift1_11[0]));
	jspl3 jspl3_w_shift1_35(.douta(w_shift1_35[0]),.doutb(w_shift1_35[1]),.doutc(w_shift1_35[2]),.din(w_shift1_11[1]));
	jspl3 jspl3_w_shift1_36(.douta(w_shift1_36[0]),.doutb(w_shift1_36[1]),.doutc(w_shift1_36[2]),.din(w_shift1_11[2]));
	jspl3 jspl3_w_shift1_37(.douta(w_shift1_37[0]),.doutb(w_shift1_37[1]),.doutc(w_shift1_37[2]),.din(w_shift1_12[0]));
	jspl3 jspl3_w_shift1_38(.douta(w_shift1_38[0]),.doutb(w_shift1_38[1]),.doutc(w_shift1_38[2]),.din(w_shift1_12[1]));
	jspl3 jspl3_w_shift1_39(.douta(w_shift1_39[0]),.doutb(w_shift1_39[1]),.doutc(w_shift1_39[2]),.din(w_shift1_12[2]));
	jspl3 jspl3_w_shift1_40(.douta(w_shift1_40[0]),.doutb(w_shift1_40[1]),.doutc(w_shift1_40[2]),.din(w_shift1_13[0]));
	jspl3 jspl3_w_shift1_41(.douta(w_shift1_41[0]),.doutb(w_shift1_41[1]),.doutc(w_shift1_41[2]),.din(w_shift1_13[1]));
	jspl3 jspl3_w_shift1_42(.douta(w_shift1_42[0]),.doutb(w_shift1_42[1]),.doutc(w_shift1_42[2]),.din(w_shift1_13[2]));
	jspl3 jspl3_w_shift1_43(.douta(w_shift1_43[0]),.doutb(w_shift1_43[1]),.doutc(w_shift1_43[2]),.din(w_shift1_14[0]));
	jspl3 jspl3_w_shift1_44(.douta(w_shift1_44[0]),.doutb(w_shift1_44[1]),.doutc(w_shift1_44[2]),.din(w_shift1_14[1]));
	jspl3 jspl3_w_shift1_45(.douta(w_shift1_45[0]),.doutb(w_shift1_45[1]),.doutc(w_shift1_45[2]),.din(w_shift1_14[2]));
	jspl3 jspl3_w_shift1_46(.douta(w_shift1_46[0]),.doutb(w_shift1_46[1]),.doutc(w_shift1_46[2]),.din(w_shift1_15[0]));
	jspl3 jspl3_w_shift1_47(.douta(w_shift1_47[0]),.doutb(w_shift1_47[1]),.doutc(w_shift1_47[2]),.din(w_shift1_15[1]));
	jspl3 jspl3_w_shift1_48(.douta(w_shift1_48[0]),.doutb(w_shift1_48[1]),.doutc(w_shift1_48[2]),.din(w_shift1_15[2]));
	jspl3 jspl3_w_shift1_49(.douta(w_shift1_49[0]),.doutb(w_shift1_49[1]),.doutc(w_shift1_49[2]),.din(w_shift1_16[0]));
	jspl3 jspl3_w_shift1_50(.douta(w_shift1_50[0]),.doutb(w_shift1_50[1]),.doutc(w_shift1_50[2]),.din(w_shift1_16[1]));
	jspl3 jspl3_w_shift1_51(.douta(w_shift1_51[0]),.doutb(w_shift1_51[1]),.doutc(w_shift1_51[2]),.din(w_shift1_16[2]));
	jspl3 jspl3_w_shift1_52(.douta(w_shift1_52[0]),.doutb(w_shift1_52[1]),.doutc(w_shift1_52[2]),.din(w_shift1_17[0]));
	jspl3 jspl3_w_shift1_53(.douta(w_shift1_53[0]),.doutb(w_shift1_53[1]),.doutc(w_shift1_53[2]),.din(w_shift1_17[1]));
	jspl3 jspl3_w_shift1_54(.douta(w_shift1_54[0]),.doutb(w_shift1_54[1]),.doutc(w_shift1_54[2]),.din(w_shift1_17[2]));
	jspl3 jspl3_w_shift1_55(.douta(w_shift1_55[0]),.doutb(w_shift1_55[1]),.doutc(w_shift1_55[2]),.din(w_shift1_18[0]));
	jspl3 jspl3_w_shift1_56(.douta(w_shift1_56[0]),.doutb(w_shift1_56[1]),.doutc(w_shift1_56[2]),.din(w_shift1_18[1]));
	jspl3 jspl3_w_shift1_57(.douta(w_shift1_57[0]),.doutb(w_shift1_57[1]),.doutc(w_shift1_57[2]),.din(w_shift1_18[2]));
	jspl3 jspl3_w_shift1_58(.douta(w_shift1_58[0]),.doutb(w_shift1_58[1]),.doutc(w_shift1_58[2]),.din(w_shift1_19[0]));
	jspl3 jspl3_w_shift1_59(.douta(w_shift1_59[0]),.doutb(w_shift1_59[1]),.doutc(w_shift1_59[2]),.din(w_shift1_19[1]));
	jspl3 jspl3_w_shift1_60(.douta(w_shift1_60[0]),.doutb(w_shift1_60[1]),.doutc(w_shift1_60[2]),.din(w_shift1_19[2]));
	jspl3 jspl3_w_shift1_61(.douta(w_shift1_61[0]),.doutb(w_shift1_61[1]),.doutc(w_shift1_61[2]),.din(w_shift1_20[0]));
	jspl3 jspl3_w_shift1_62(.douta(w_shift1_62[0]),.doutb(w_shift1_62[1]),.doutc(w_shift1_62[2]),.din(w_shift1_20[1]));
	jspl3 jspl3_w_shift1_63(.douta(w_shift1_63[0]),.doutb(w_shift1_63[1]),.doutc(w_shift1_63[2]),.din(w_shift1_20[2]));
	jspl3 jspl3_w_shift1_64(.douta(w_shift1_64[0]),.doutb(w_shift1_64[1]),.doutc(w_shift1_64[2]),.din(w_shift1_21[0]));
	jspl3 jspl3_w_shift1_65(.douta(w_shift1_65[0]),.doutb(w_shift1_65[1]),.doutc(w_shift1_65[2]),.din(w_shift1_21[1]));
	jspl3 jspl3_w_shift1_66(.douta(w_shift1_66[0]),.doutb(w_shift1_66[1]),.doutc(w_shift1_66[2]),.din(w_shift1_21[2]));
	jspl3 jspl3_w_shift1_67(.douta(w_shift1_67[0]),.doutb(w_shift1_67[1]),.doutc(w_shift1_67[2]),.din(w_shift1_22[0]));
	jspl3 jspl3_w_shift1_68(.douta(w_shift1_68[0]),.doutb(w_shift1_68[1]),.doutc(w_shift1_68[2]),.din(w_shift1_22[1]));
	jspl3 jspl3_w_shift1_69(.douta(w_shift1_69[0]),.doutb(w_shift1_69[1]),.doutc(w_shift1_69[2]),.din(w_shift1_22[2]));
	jspl3 jspl3_w_shift1_70(.douta(w_shift1_70[0]),.doutb(w_shift1_70[1]),.doutc(w_shift1_70[2]),.din(w_shift1_23[0]));
	jspl3 jspl3_w_shift1_71(.douta(w_shift1_71[0]),.doutb(w_shift1_71[1]),.doutc(w_shift1_71[2]),.din(w_shift1_23[1]));
	jspl3 jspl3_w_shift1_72(.douta(w_shift1_72[0]),.doutb(w_shift1_72[1]),.doutc(w_shift1_72[2]),.din(w_shift1_23[2]));
	jspl3 jspl3_w_shift1_73(.douta(w_shift1_73[0]),.doutb(w_shift1_73[1]),.doutc(w_shift1_73[2]),.din(w_shift1_24[0]));
	jspl3 jspl3_w_shift1_74(.douta(w_shift1_74[0]),.doutb(w_shift1_74[1]),.doutc(w_shift1_74[2]),.din(w_shift1_24[1]));
	jspl3 jspl3_w_shift1_75(.douta(w_shift1_75[0]),.doutb(w_shift1_75[1]),.doutc(w_shift1_75[2]),.din(w_shift1_24[2]));
	jspl3 jspl3_w_shift1_76(.douta(w_shift1_76[0]),.doutb(w_shift1_76[1]),.doutc(w_shift1_76[2]),.din(w_shift1_25[0]));
	jspl3 jspl3_w_shift1_77(.douta(w_shift1_77[0]),.doutb(w_shift1_77[1]),.doutc(w_shift1_77[2]),.din(w_shift1_25[1]));
	jspl3 jspl3_w_shift1_78(.douta(w_shift1_78[0]),.doutb(w_shift1_78[1]),.doutc(w_shift1_78[2]),.din(w_shift1_25[2]));
	jspl3 jspl3_w_shift1_79(.douta(w_shift1_79[0]),.doutb(w_shift1_79[1]),.doutc(w_shift1_79[2]),.din(w_shift1_26[0]));
	jspl3 jspl3_w_shift1_80(.douta(w_shift1_80[0]),.doutb(w_shift1_80[1]),.doutc(w_shift1_80[2]),.din(w_shift1_26[1]));
	jspl3 jspl3_w_shift1_81(.douta(w_shift1_81[0]),.doutb(w_shift1_81[1]),.doutc(w_shift1_81[2]),.din(w_shift1_26[2]));
	jspl3 jspl3_w_shift1_82(.douta(w_shift1_82[0]),.doutb(w_shift1_82[1]),.doutc(w_shift1_82[2]),.din(w_shift1_27[0]));
	jspl3 jspl3_w_shift1_83(.douta(w_shift1_83[0]),.doutb(w_shift1_83[1]),.doutc(w_shift1_83[2]),.din(w_shift1_27[1]));
	jspl3 jspl3_w_shift1_84(.douta(w_shift1_84[0]),.doutb(w_shift1_84[1]),.doutc(w_shift1_84[2]),.din(w_shift1_27[2]));
	jspl3 jspl3_w_shift1_85(.douta(w_shift1_85[0]),.doutb(w_shift1_85[1]),.doutc(w_shift1_85[2]),.din(w_shift1_28[0]));
	jspl3 jspl3_w_shift1_86(.douta(w_shift1_86[0]),.doutb(w_shift1_86[1]),.doutc(w_shift1_86[2]),.din(w_shift1_28[1]));
	jspl3 jspl3_w_shift1_87(.douta(w_shift1_87[0]),.doutb(w_shift1_87[1]),.doutc(w_shift1_87[2]),.din(w_shift1_28[2]));
	jspl3 jspl3_w_shift1_88(.douta(w_shift1_88[0]),.doutb(w_shift1_88[1]),.doutc(w_shift1_88[2]),.din(w_shift1_29[0]));
	jspl3 jspl3_w_shift1_89(.douta(w_shift1_89[0]),.doutb(w_shift1_89[1]),.doutc(w_shift1_89[2]),.din(w_shift1_29[1]));
	jspl3 jspl3_w_shift1_90(.douta(w_shift1_90[0]),.doutb(w_shift1_90[1]),.doutc(w_shift1_90[2]),.din(w_shift1_29[2]));
	jspl3 jspl3_w_shift1_91(.douta(w_shift1_91[0]),.doutb(w_shift1_91[1]),.doutc(w_shift1_91[2]),.din(w_shift1_30[0]));
	jspl3 jspl3_w_shift1_92(.douta(w_shift1_92[0]),.doutb(w_shift1_92[1]),.doutc(w_shift1_92[2]),.din(w_shift1_30[1]));
	jspl3 jspl3_w_shift1_93(.douta(w_shift1_93[0]),.doutb(w_shift1_93[1]),.doutc(w_shift1_93[2]),.din(w_shift1_30[2]));
	jspl3 jspl3_w_shift1_94(.douta(w_shift1_94[0]),.doutb(w_shift1_94[1]),.doutc(w_shift1_94[2]),.din(w_shift1_31[0]));
	jspl3 jspl3_w_shift1_95(.douta(w_shift1_95[0]),.doutb(w_shift1_95[1]),.doutc(w_shift1_95[2]),.din(w_shift1_31[1]));
	jspl3 jspl3_w_shift1_96(.douta(w_shift1_96[0]),.doutb(w_shift1_96[1]),.doutc(w_shift1_96[2]),.din(w_shift1_31[2]));
	jspl3 jspl3_w_shift2_0(.douta(w_shift2_0[0]),.doutb(w_shift2_0[1]),.doutc(w_shift2_0[2]),.din(shift2));
	jspl3 jspl3_w_shift3_0(.douta(w_shift3_0[0]),.doutb(w_shift3_0[1]),.doutc(w_shift3_0[2]),.din(shift3));
	jspl3 jspl3_w_shift4_0(.douta(w_shift4_0[0]),.doutb(w_shift4_0[1]),.doutc(w_shift4_0[2]),.din(shift4));
	jspl3 jspl3_w_shift5_0(.douta(w_shift5_0[0]),.doutb(w_shift5_0[1]),.doutc(w_shift5_0[2]),.din(shift5));
	jspl3 jspl3_w_shift6_0(.douta(w_shift6_0[0]),.doutb(w_shift6_0[1]),.doutc(w_shift6_0[2]),.din(shift6));
	jspl3 jspl3_w_shift6_1(.douta(w_shift6_1[0]),.doutb(w_shift6_1[1]),.doutc(w_shift6_1[2]),.din(w_shift6_0[0]));
	jspl3 jspl3_w_shift6_2(.douta(w_shift6_2[0]),.doutb(w_shift6_2[1]),.doutc(w_shift6_2[2]),.din(w_shift6_0[1]));
	jspl3 jspl3_w_shift6_3(.douta(w_shift6_3[0]),.doutb(w_shift6_3[1]),.doutc(w_shift6_3[2]),.din(w_shift6_0[2]));
	jspl3 jspl3_w_shift6_4(.douta(w_shift6_4[0]),.doutb(w_shift6_4[1]),.doutc(w_shift6_4[2]),.din(w_shift6_1[0]));
	jspl3 jspl3_w_shift6_5(.douta(w_shift6_5[0]),.doutb(w_shift6_5[1]),.doutc(w_shift6_5[2]),.din(w_shift6_1[1]));
	jspl3 jspl3_w_shift6_6(.douta(w_shift6_6[0]),.doutb(w_shift6_6[1]),.doutc(w_shift6_6[2]),.din(w_shift6_1[2]));
	jspl3 jspl3_w_shift6_7(.douta(w_shift6_7[0]),.doutb(w_shift6_7[1]),.doutc(w_shift6_7[2]),.din(w_shift6_2[0]));
	jspl3 jspl3_w_shift6_8(.douta(w_shift6_8[0]),.doutb(w_shift6_8[1]),.doutc(w_shift6_8[2]),.din(w_shift6_2[1]));
	jspl3 jspl3_w_shift6_9(.douta(w_shift6_9[0]),.doutb(w_shift6_9[1]),.doutc(w_shift6_9[2]),.din(w_shift6_2[2]));
	jspl3 jspl3_w_shift6_10(.douta(w_shift6_10[0]),.doutb(w_shift6_10[1]),.doutc(w_shift6_10[2]),.din(w_shift6_3[0]));
	jspl3 jspl3_w_shift6_11(.douta(w_shift6_11[0]),.doutb(w_shift6_11[1]),.doutc(w_shift6_11[2]),.din(w_shift6_3[1]));
	jspl3 jspl3_w_shift6_12(.douta(w_shift6_12[0]),.doutb(w_shift6_12[1]),.doutc(w_shift6_12[2]),.din(w_shift6_3[2]));
	jspl3 jspl3_w_shift6_13(.douta(w_shift6_13[0]),.doutb(w_shift6_13[1]),.doutc(w_shift6_13[2]),.din(w_shift6_4[0]));
	jspl3 jspl3_w_shift6_14(.douta(w_shift6_14[0]),.doutb(w_shift6_14[1]),.doutc(w_shift6_14[2]),.din(w_shift6_4[1]));
	jspl3 jspl3_w_shift6_15(.douta(w_shift6_15[0]),.doutb(w_shift6_15[1]),.doutc(w_shift6_15[2]),.din(w_shift6_4[2]));
	jspl3 jspl3_w_shift6_16(.douta(w_shift6_16[0]),.doutb(w_shift6_16[1]),.doutc(w_shift6_16[2]),.din(w_shift6_5[0]));
	jspl3 jspl3_w_shift6_17(.douta(w_shift6_17[0]),.doutb(w_shift6_17[1]),.doutc(w_shift6_17[2]),.din(w_shift6_5[1]));
	jspl3 jspl3_w_shift6_18(.douta(w_shift6_18[0]),.doutb(w_shift6_18[1]),.doutc(w_shift6_18[2]),.din(w_shift6_5[2]));
	jspl3 jspl3_w_shift6_19(.douta(w_shift6_19[0]),.doutb(w_shift6_19[1]),.doutc(w_shift6_19[2]),.din(w_shift6_6[0]));
	jspl3 jspl3_w_shift6_20(.douta(w_shift6_20[0]),.doutb(w_shift6_20[1]),.doutc(w_shift6_20[2]),.din(w_shift6_6[1]));
	jspl3 jspl3_w_shift6_21(.douta(w_shift6_21[0]),.doutb(w_shift6_21[1]),.doutc(w_shift6_21[2]),.din(w_shift6_6[2]));
	jspl3 jspl3_w_shift6_22(.douta(w_shift6_22[0]),.doutb(w_shift6_22[1]),.doutc(w_shift6_22[2]),.din(w_shift6_7[0]));
	jspl3 jspl3_w_shift6_23(.douta(w_shift6_23[0]),.doutb(w_shift6_23[1]),.doutc(w_shift6_23[2]),.din(w_shift6_7[1]));
	jspl3 jspl3_w_shift6_24(.douta(w_shift6_24[0]),.doutb(w_shift6_24[1]),.doutc(w_shift6_24[2]),.din(w_shift6_7[2]));
	jspl3 jspl3_w_shift6_25(.douta(w_shift6_25[0]),.doutb(w_shift6_25[1]),.doutc(w_shift6_25[2]),.din(w_shift6_8[0]));
	jspl3 jspl3_w_shift6_26(.douta(w_shift6_26[0]),.doutb(w_shift6_26[1]),.doutc(w_shift6_26[2]),.din(w_shift6_8[1]));
	jspl3 jspl3_w_shift6_27(.douta(w_shift6_27[0]),.doutb(w_shift6_27[1]),.doutc(w_shift6_27[2]),.din(w_shift6_8[2]));
	jspl3 jspl3_w_shift6_28(.douta(w_shift6_28[0]),.doutb(w_shift6_28[1]),.doutc(w_shift6_28[2]),.din(w_shift6_9[0]));
	jspl3 jspl3_w_shift6_29(.douta(w_shift6_29[0]),.doutb(w_shift6_29[1]),.doutc(w_shift6_29[2]),.din(w_shift6_9[1]));
	jspl3 jspl3_w_shift6_30(.douta(w_shift6_30[0]),.doutb(w_shift6_30[1]),.doutc(w_shift6_30[2]),.din(w_shift6_9[2]));
	jspl3 jspl3_w_shift6_31(.douta(w_shift6_31[0]),.doutb(w_shift6_31[1]),.doutc(w_shift6_31[2]),.din(w_shift6_10[0]));
	jspl3 jspl3_w_shift6_32(.douta(w_shift6_32[0]),.doutb(w_shift6_32[1]),.doutc(w_shift6_32[2]),.din(w_shift6_10[1]));
	jspl3 jspl3_w_shift6_33(.douta(w_shift6_33[0]),.doutb(w_shift6_33[1]),.doutc(w_shift6_33[2]),.din(w_shift6_10[2]));
	jspl3 jspl3_w_shift6_34(.douta(w_shift6_34[0]),.doutb(w_shift6_34[1]),.doutc(w_shift6_34[2]),.din(w_shift6_11[0]));
	jspl3 jspl3_w_shift6_35(.douta(w_shift6_35[0]),.doutb(w_shift6_35[1]),.doutc(w_shift6_35[2]),.din(w_shift6_11[1]));
	jspl3 jspl3_w_shift6_36(.douta(w_shift6_36[0]),.doutb(w_shift6_36[1]),.doutc(w_shift6_36[2]),.din(w_shift6_11[2]));
	jspl3 jspl3_w_shift6_37(.douta(w_shift6_37[0]),.doutb(w_shift6_37[1]),.doutc(w_shift6_37[2]),.din(w_shift6_12[0]));
	jspl3 jspl3_w_shift6_38(.douta(w_shift6_38[0]),.doutb(w_shift6_38[1]),.doutc(w_shift6_38[2]),.din(w_shift6_12[1]));
	jspl3 jspl3_w_shift6_39(.douta(w_shift6_39[0]),.doutb(w_shift6_39[1]),.doutc(w_shift6_39[2]),.din(w_shift6_12[2]));
	jspl3 jspl3_w_shift6_40(.douta(w_shift6_40[0]),.doutb(w_shift6_40[1]),.doutc(w_shift6_40[2]),.din(w_shift6_13[0]));
	jspl3 jspl3_w_shift6_41(.douta(w_shift6_41[0]),.doutb(w_shift6_41[1]),.doutc(w_shift6_41[2]),.din(w_shift6_13[1]));
	jspl3 jspl3_w_shift6_42(.douta(w_shift6_42[0]),.doutb(w_shift6_42[1]),.doutc(w_shift6_42[2]),.din(w_shift6_13[2]));
	jspl3 jspl3_w_shift6_43(.douta(w_shift6_43[0]),.doutb(w_shift6_43[1]),.doutc(w_shift6_43[2]),.din(w_shift6_14[0]));
	jspl3 jspl3_w_shift6_44(.douta(w_shift6_44[0]),.doutb(w_shift6_44[1]),.doutc(w_shift6_44[2]),.din(w_shift6_14[1]));
	jspl3 jspl3_w_shift6_45(.douta(w_shift6_45[0]),.doutb(w_shift6_45[1]),.doutc(w_shift6_45[2]),.din(w_shift6_14[2]));
	jspl3 jspl3_w_shift6_46(.douta(w_shift6_46[0]),.doutb(w_shift6_46[1]),.doutc(w_shift6_46[2]),.din(w_shift6_15[0]));
	jspl3 jspl3_w_shift6_47(.douta(w_shift6_47[0]),.doutb(w_shift6_47[1]),.doutc(w_shift6_47[2]),.din(w_shift6_15[1]));
	jspl3 jspl3_w_shift6_48(.douta(w_shift6_48[0]),.doutb(w_shift6_48[1]),.doutc(w_shift6_48[2]),.din(w_shift6_15[2]));
	jspl3 jspl3_w_shift6_49(.douta(w_shift6_49[0]),.doutb(w_shift6_49[1]),.doutc(w_shift6_49[2]),.din(w_shift6_16[0]));
	jspl3 jspl3_w_shift6_50(.douta(w_shift6_50[0]),.doutb(w_shift6_50[1]),.doutc(w_shift6_50[2]),.din(w_shift6_16[1]));
	jspl3 jspl3_w_shift6_51(.douta(w_shift6_51[0]),.doutb(w_shift6_51[1]),.doutc(w_shift6_51[2]),.din(w_shift6_16[2]));
	jspl3 jspl3_w_shift6_52(.douta(w_shift6_52[0]),.doutb(w_shift6_52[1]),.doutc(w_shift6_52[2]),.din(w_shift6_17[0]));
	jspl3 jspl3_w_shift6_53(.douta(w_shift6_53[0]),.doutb(w_shift6_53[1]),.doutc(w_shift6_53[2]),.din(w_shift6_17[1]));
	jspl3 jspl3_w_shift6_54(.douta(w_shift6_54[0]),.doutb(w_shift6_54[1]),.doutc(w_shift6_54[2]),.din(w_shift6_17[2]));
	jspl3 jspl3_w_shift6_55(.douta(w_shift6_55[0]),.doutb(w_shift6_55[1]),.doutc(w_shift6_55[2]),.din(w_shift6_18[0]));
	jspl3 jspl3_w_shift6_56(.douta(w_shift6_56[0]),.doutb(w_shift6_56[1]),.doutc(w_shift6_56[2]),.din(w_shift6_18[1]));
	jspl3 jspl3_w_shift6_57(.douta(w_shift6_57[0]),.doutb(w_shift6_57[1]),.doutc(w_shift6_57[2]),.din(w_shift6_18[2]));
	jspl3 jspl3_w_shift6_58(.douta(w_shift6_58[0]),.doutb(w_shift6_58[1]),.doutc(w_shift6_58[2]),.din(w_shift6_19[0]));
	jspl3 jspl3_w_shift6_59(.douta(w_shift6_59[0]),.doutb(w_shift6_59[1]),.doutc(w_shift6_59[2]),.din(w_shift6_19[1]));
	jspl3 jspl3_w_shift6_60(.douta(w_shift6_60[0]),.doutb(w_shift6_60[1]),.doutc(w_shift6_60[2]),.din(w_shift6_19[2]));
	jspl3 jspl3_w_shift6_61(.douta(w_shift6_61[0]),.doutb(w_shift6_61[1]),.doutc(w_shift6_61[2]),.din(w_shift6_20[0]));
	jspl3 jspl3_w_shift6_62(.douta(w_shift6_62[0]),.doutb(w_shift6_62[1]),.doutc(w_shift6_62[2]),.din(w_shift6_20[1]));
	jspl3 jspl3_w_shift6_63(.douta(w_shift6_63[0]),.doutb(w_shift6_63[1]),.doutc(w_shift6_63[2]),.din(w_shift6_20[2]));
	jspl3 jspl3_w_n263_0(.douta(w_n263_0[0]),.doutb(w_n263_0[1]),.doutc(w_n263_0[2]),.din(n263));
	jspl3 jspl3_w_n263_1(.douta(w_n263_1[0]),.doutb(w_n263_1[1]),.doutc(w_n263_1[2]),.din(w_n263_0[0]));
	jspl3 jspl3_w_n263_2(.douta(w_n263_2[0]),.doutb(w_n263_2[1]),.doutc(w_n263_2[2]),.din(w_n263_0[1]));
	jspl3 jspl3_w_n263_3(.douta(w_n263_3[0]),.doutb(w_n263_3[1]),.doutc(w_n263_3[2]),.din(w_n263_0[2]));
	jspl3 jspl3_w_n263_4(.douta(w_n263_4[0]),.doutb(w_n263_4[1]),.doutc(w_n263_4[2]),.din(w_n263_1[0]));
	jspl3 jspl3_w_n263_5(.douta(w_n263_5[0]),.doutb(w_n263_5[1]),.doutc(w_n263_5[2]),.din(w_n263_1[1]));
	jspl3 jspl3_w_n263_6(.douta(w_n263_6[0]),.doutb(w_n263_6[1]),.doutc(w_n263_6[2]),.din(w_n263_1[2]));
	jspl3 jspl3_w_n263_7(.douta(w_n263_7[0]),.doutb(w_n263_7[1]),.doutc(w_n263_7[2]),.din(w_n263_2[0]));
	jspl3 jspl3_w_n263_8(.douta(w_n263_8[0]),.doutb(w_n263_8[1]),.doutc(w_n263_8[2]),.din(w_n263_2[1]));
	jspl3 jspl3_w_n263_9(.douta(w_n263_9[0]),.doutb(w_n263_9[1]),.doutc(w_n263_9[2]),.din(w_n263_2[2]));
	jspl3 jspl3_w_n263_10(.douta(w_n263_10[0]),.doutb(w_n263_10[1]),.doutc(w_n263_10[2]),.din(w_n263_3[0]));
	jspl3 jspl3_w_n263_11(.douta(w_n263_11[0]),.doutb(w_n263_11[1]),.doutc(w_n263_11[2]),.din(w_n263_3[1]));
	jspl3 jspl3_w_n263_12(.douta(w_n263_12[0]),.doutb(w_n263_12[1]),.doutc(w_n263_12[2]),.din(w_n263_3[2]));
	jspl3 jspl3_w_n263_13(.douta(w_n263_13[0]),.doutb(w_n263_13[1]),.doutc(w_n263_13[2]),.din(w_n263_4[0]));
	jspl3 jspl3_w_n263_14(.douta(w_n263_14[0]),.doutb(w_n263_14[1]),.doutc(w_n263_14[2]),.din(w_n263_4[1]));
	jspl3 jspl3_w_n263_15(.douta(w_n263_15[0]),.doutb(w_n263_15[1]),.doutc(w_n263_15[2]),.din(w_n263_4[2]));
	jspl3 jspl3_w_n263_16(.douta(w_n263_16[0]),.doutb(w_n263_16[1]),.doutc(w_n263_16[2]),.din(w_n263_5[0]));
	jspl3 jspl3_w_n263_17(.douta(w_n263_17[0]),.doutb(w_n263_17[1]),.doutc(w_n263_17[2]),.din(w_n263_5[1]));
	jspl3 jspl3_w_n263_18(.douta(w_n263_18[0]),.doutb(w_n263_18[1]),.doutc(w_n263_18[2]),.din(w_n263_5[2]));
	jspl3 jspl3_w_n263_19(.douta(w_n263_19[0]),.doutb(w_n263_19[1]),.doutc(w_n263_19[2]),.din(w_n263_6[0]));
	jspl3 jspl3_w_n263_20(.douta(w_n263_20[0]),.doutb(w_n263_20[1]),.doutc(w_n263_20[2]),.din(w_n263_6[1]));
	jspl3 jspl3_w_n263_21(.douta(w_n263_21[0]),.doutb(w_n263_21[1]),.doutc(w_n263_21[2]),.din(w_n263_6[2]));
	jspl3 jspl3_w_n263_22(.douta(w_n263_22[0]),.doutb(w_n263_22[1]),.doutc(w_n263_22[2]),.din(w_n263_7[0]));
	jspl3 jspl3_w_n263_23(.douta(w_n263_23[0]),.doutb(w_n263_23[1]),.doutc(w_n263_23[2]),.din(w_n263_7[1]));
	jspl3 jspl3_w_n263_24(.douta(w_n263_24[0]),.doutb(w_n263_24[1]),.doutc(w_n263_24[2]),.din(w_n263_7[2]));
	jspl3 jspl3_w_n263_25(.douta(w_n263_25[0]),.doutb(w_n263_25[1]),.doutc(w_n263_25[2]),.din(w_n263_8[0]));
	jspl3 jspl3_w_n263_26(.douta(w_n263_26[0]),.doutb(w_n263_26[1]),.doutc(w_n263_26[2]),.din(w_n263_8[1]));
	jspl3 jspl3_w_n263_27(.douta(w_n263_27[0]),.doutb(w_n263_27[1]),.doutc(w_n263_27[2]),.din(w_n263_8[2]));
	jspl3 jspl3_w_n263_28(.douta(w_n263_28[0]),.doutb(w_n263_28[1]),.doutc(w_n263_28[2]),.din(w_n263_9[0]));
	jspl3 jspl3_w_n263_29(.douta(w_n263_29[0]),.doutb(w_n263_29[1]),.doutc(w_n263_29[2]),.din(w_n263_9[1]));
	jspl3 jspl3_w_n263_30(.douta(w_n263_30[0]),.doutb(w_n263_30[1]),.doutc(w_n263_30[2]),.din(w_n263_9[2]));
	jspl3 jspl3_w_n263_31(.douta(w_n263_31[0]),.doutb(w_n263_31[1]),.doutc(w_n263_31[2]),.din(w_n263_10[0]));
	jspl3 jspl3_w_n263_32(.douta(w_n263_32[0]),.doutb(w_n263_32[1]),.doutc(w_n263_32[2]),.din(w_n263_10[1]));
	jspl3 jspl3_w_n263_33(.douta(w_n263_33[0]),.doutb(w_n263_33[1]),.doutc(w_n263_33[2]),.din(w_n263_10[2]));
	jspl3 jspl3_w_n263_34(.douta(w_n263_34[0]),.doutb(w_n263_34[1]),.doutc(w_n263_34[2]),.din(w_n263_11[0]));
	jspl3 jspl3_w_n263_35(.douta(w_n263_35[0]),.doutb(w_n263_35[1]),.doutc(w_n263_35[2]),.din(w_n263_11[1]));
	jspl3 jspl3_w_n263_36(.douta(w_n263_36[0]),.doutb(w_n263_36[1]),.doutc(w_n263_36[2]),.din(w_n263_11[2]));
	jspl3 jspl3_w_n263_37(.douta(w_n263_37[0]),.doutb(w_n263_37[1]),.doutc(w_n263_37[2]),.din(w_n263_12[0]));
	jspl3 jspl3_w_n263_38(.douta(w_n263_38[0]),.doutb(w_n263_38[1]),.doutc(w_n263_38[2]),.din(w_n263_12[1]));
	jspl3 jspl3_w_n263_39(.douta(w_n263_39[0]),.doutb(w_n263_39[1]),.doutc(w_n263_39[2]),.din(w_n263_12[2]));
	jspl3 jspl3_w_n263_40(.douta(w_n263_40[0]),.doutb(w_n263_40[1]),.doutc(w_n263_40[2]),.din(w_n263_13[0]));
	jspl3 jspl3_w_n263_41(.douta(w_n263_41[0]),.doutb(w_n263_41[1]),.doutc(w_n263_41[2]),.din(w_n263_13[1]));
	jspl3 jspl3_w_n263_42(.douta(w_n263_42[0]),.doutb(w_n263_42[1]),.doutc(w_n263_42[2]),.din(w_n263_13[2]));
	jspl3 jspl3_w_n263_43(.douta(w_n263_43[0]),.doutb(w_n263_43[1]),.doutc(w_n263_43[2]),.din(w_n263_14[0]));
	jspl3 jspl3_w_n263_44(.douta(w_n263_44[0]),.doutb(w_n263_44[1]),.doutc(w_n263_44[2]),.din(w_n263_14[1]));
	jspl3 jspl3_w_n263_45(.douta(w_n263_45[0]),.doutb(w_n263_45[1]),.doutc(w_n263_45[2]),.din(w_n263_14[2]));
	jspl3 jspl3_w_n263_46(.douta(w_n263_46[0]),.doutb(w_n263_46[1]),.doutc(w_n263_46[2]),.din(w_n263_15[0]));
	jspl3 jspl3_w_n263_47(.douta(w_n263_47[0]),.doutb(w_n263_47[1]),.doutc(w_n263_47[2]),.din(w_n263_15[1]));
	jspl3 jspl3_w_n263_48(.douta(w_n263_48[0]),.doutb(w_n263_48[1]),.doutc(w_n263_48[2]),.din(w_n263_15[2]));
	jspl3 jspl3_w_n263_49(.douta(w_n263_49[0]),.doutb(w_n263_49[1]),.doutc(w_n263_49[2]),.din(w_n263_16[0]));
	jspl3 jspl3_w_n263_50(.douta(w_n263_50[0]),.doutb(w_n263_50[1]),.doutc(w_n263_50[2]),.din(w_n263_16[1]));
	jspl3 jspl3_w_n263_51(.douta(w_n263_51[0]),.doutb(w_n263_51[1]),.doutc(w_n263_51[2]),.din(w_n263_16[2]));
	jspl3 jspl3_w_n263_52(.douta(w_n263_52[0]),.doutb(w_n263_52[1]),.doutc(w_n263_52[2]),.din(w_n263_17[0]));
	jspl3 jspl3_w_n263_53(.douta(w_n263_53[0]),.doutb(w_n263_53[1]),.doutc(w_n263_53[2]),.din(w_n263_17[1]));
	jspl3 jspl3_w_n263_54(.douta(w_n263_54[0]),.doutb(w_n263_54[1]),.doutc(w_n263_54[2]),.din(w_n263_17[2]));
	jspl3 jspl3_w_n263_55(.douta(w_n263_55[0]),.doutb(w_n263_55[1]),.doutc(w_n263_55[2]),.din(w_n263_18[0]));
	jspl3 jspl3_w_n263_56(.douta(w_n263_56[0]),.doutb(w_n263_56[1]),.doutc(w_n263_56[2]),.din(w_n263_18[1]));
	jspl3 jspl3_w_n263_57(.douta(w_n263_57[0]),.doutb(w_n263_57[1]),.doutc(w_n263_57[2]),.din(w_n263_18[2]));
	jspl3 jspl3_w_n263_58(.douta(w_n263_58[0]),.doutb(w_n263_58[1]),.doutc(w_n263_58[2]),.din(w_n263_19[0]));
	jspl3 jspl3_w_n263_59(.douta(w_n263_59[0]),.doutb(w_n263_59[1]),.doutc(w_n263_59[2]),.din(w_n263_19[1]));
	jspl3 jspl3_w_n263_60(.douta(w_n263_60[0]),.doutb(w_n263_60[1]),.doutc(w_n263_60[2]),.din(w_n263_19[2]));
	jspl3 jspl3_w_n263_61(.douta(w_n263_61[0]),.doutb(w_n263_61[1]),.doutc(w_n263_61[2]),.din(w_n263_20[0]));
	jspl3 jspl3_w_n263_62(.douta(w_n263_62[0]),.doutb(w_n263_62[1]),.doutc(w_n263_62[2]),.din(w_n263_20[1]));
	jspl jspl_w_n263_63(.douta(w_n263_63[0]),.doutb(w_n263_63[1]),.din(w_n263_20[2]));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(n265));
	jspl3 jspl3_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.doutc(w_n266_0[2]),.din(n266));
	jspl3 jspl3_w_n266_1(.douta(w_n266_1[0]),.doutb(w_n266_1[1]),.doutc(w_n266_1[2]),.din(w_n266_0[0]));
	jspl3 jspl3_w_n266_2(.douta(w_n266_2[0]),.doutb(w_n266_2[1]),.doutc(w_n266_2[2]),.din(w_n266_0[1]));
	jspl3 jspl3_w_n266_3(.douta(w_n266_3[0]),.doutb(w_n266_3[1]),.doutc(w_n266_3[2]),.din(w_n266_0[2]));
	jspl3 jspl3_w_n266_4(.douta(w_n266_4[0]),.doutb(w_n266_4[1]),.doutc(w_n266_4[2]),.din(w_n266_1[0]));
	jspl3 jspl3_w_n266_5(.douta(w_n266_5[0]),.doutb(w_n266_5[1]),.doutc(w_n266_5[2]),.din(w_n266_1[1]));
	jspl3 jspl3_w_n266_6(.douta(w_n266_6[0]),.doutb(w_n266_6[1]),.doutc(w_n266_6[2]),.din(w_n266_1[2]));
	jspl3 jspl3_w_n266_7(.douta(w_n266_7[0]),.doutb(w_n266_7[1]),.doutc(w_n266_7[2]),.din(w_n266_2[0]));
	jspl3 jspl3_w_n266_8(.douta(w_n266_8[0]),.doutb(w_n266_8[1]),.doutc(w_n266_8[2]),.din(w_n266_2[1]));
	jspl3 jspl3_w_n266_9(.douta(w_n266_9[0]),.doutb(w_n266_9[1]),.doutc(w_n266_9[2]),.din(w_n266_2[2]));
	jspl3 jspl3_w_n266_10(.douta(w_n266_10[0]),.doutb(w_n266_10[1]),.doutc(w_n266_10[2]),.din(w_n266_3[0]));
	jspl3 jspl3_w_n266_11(.douta(w_n266_11[0]),.doutb(w_n266_11[1]),.doutc(w_n266_11[2]),.din(w_n266_3[1]));
	jspl3 jspl3_w_n266_12(.douta(w_n266_12[0]),.doutb(w_n266_12[1]),.doutc(w_n266_12[2]),.din(w_n266_3[2]));
	jspl3 jspl3_w_n266_13(.douta(w_n266_13[0]),.doutb(w_n266_13[1]),.doutc(w_n266_13[2]),.din(w_n266_4[0]));
	jspl3 jspl3_w_n266_14(.douta(w_n266_14[0]),.doutb(w_n266_14[1]),.doutc(w_n266_14[2]),.din(w_n266_4[1]));
	jspl3 jspl3_w_n266_15(.douta(w_n266_15[0]),.doutb(w_n266_15[1]),.doutc(w_n266_15[2]),.din(w_n266_4[2]));
	jspl3 jspl3_w_n266_16(.douta(w_n266_16[0]),.doutb(w_n266_16[1]),.doutc(w_n266_16[2]),.din(w_n266_5[0]));
	jspl3 jspl3_w_n266_17(.douta(w_n266_17[0]),.doutb(w_n266_17[1]),.doutc(w_n266_17[2]),.din(w_n266_5[1]));
	jspl3 jspl3_w_n266_18(.douta(w_n266_18[0]),.doutb(w_n266_18[1]),.doutc(w_n266_18[2]),.din(w_n266_5[2]));
	jspl3 jspl3_w_n266_19(.douta(w_n266_19[0]),.doutb(w_n266_19[1]),.doutc(w_n266_19[2]),.din(w_n266_6[0]));
	jspl3 jspl3_w_n266_20(.douta(w_n266_20[0]),.doutb(w_n266_20[1]),.doutc(w_n266_20[2]),.din(w_n266_6[1]));
	jspl3 jspl3_w_n266_21(.douta(w_n266_21[0]),.doutb(w_n266_21[1]),.doutc(w_n266_21[2]),.din(w_n266_6[2]));
	jspl3 jspl3_w_n266_22(.douta(w_n266_22[0]),.doutb(w_n266_22[1]),.doutc(w_n266_22[2]),.din(w_n266_7[0]));
	jspl3 jspl3_w_n266_23(.douta(w_n266_23[0]),.doutb(w_n266_23[1]),.doutc(w_n266_23[2]),.din(w_n266_7[1]));
	jspl3 jspl3_w_n266_24(.douta(w_n266_24[0]),.doutb(w_n266_24[1]),.doutc(w_n266_24[2]),.din(w_n266_7[2]));
	jspl3 jspl3_w_n266_25(.douta(w_n266_25[0]),.doutb(w_n266_25[1]),.doutc(w_n266_25[2]),.din(w_n266_8[0]));
	jspl3 jspl3_w_n266_26(.douta(w_n266_26[0]),.doutb(w_n266_26[1]),.doutc(w_n266_26[2]),.din(w_n266_8[1]));
	jspl3 jspl3_w_n266_27(.douta(w_n266_27[0]),.doutb(w_n266_27[1]),.doutc(w_n266_27[2]),.din(w_n266_8[2]));
	jspl3 jspl3_w_n266_28(.douta(w_n266_28[0]),.doutb(w_n266_28[1]),.doutc(w_n266_28[2]),.din(w_n266_9[0]));
	jspl3 jspl3_w_n266_29(.douta(w_n266_29[0]),.doutb(w_n266_29[1]),.doutc(w_n266_29[2]),.din(w_n266_9[1]));
	jspl3 jspl3_w_n266_30(.douta(w_n266_30[0]),.doutb(w_n266_30[1]),.doutc(w_n266_30[2]),.din(w_n266_9[2]));
	jspl3 jspl3_w_n266_31(.douta(w_n266_31[0]),.doutb(w_n266_31[1]),.doutc(w_n266_31[2]),.din(w_n266_10[0]));
	jspl3 jspl3_w_n266_32(.douta(w_n266_32[0]),.doutb(w_n266_32[1]),.doutc(w_n266_32[2]),.din(w_n266_10[1]));
	jspl3 jspl3_w_n266_33(.douta(w_n266_33[0]),.doutb(w_n266_33[1]),.doutc(w_n266_33[2]),.din(w_n266_10[2]));
	jspl3 jspl3_w_n266_34(.douta(w_n266_34[0]),.doutb(w_n266_34[1]),.doutc(w_n266_34[2]),.din(w_n266_11[0]));
	jspl3 jspl3_w_n266_35(.douta(w_n266_35[0]),.doutb(w_n266_35[1]),.doutc(w_n266_35[2]),.din(w_n266_11[1]));
	jspl3 jspl3_w_n266_36(.douta(w_n266_36[0]),.doutb(w_n266_36[1]),.doutc(w_n266_36[2]),.din(w_n266_11[2]));
	jspl3 jspl3_w_n266_37(.douta(w_n266_37[0]),.doutb(w_n266_37[1]),.doutc(w_n266_37[2]),.din(w_n266_12[0]));
	jspl3 jspl3_w_n266_38(.douta(w_n266_38[0]),.doutb(w_n266_38[1]),.doutc(w_n266_38[2]),.din(w_n266_12[1]));
	jspl3 jspl3_w_n266_39(.douta(w_n266_39[0]),.doutb(w_n266_39[1]),.doutc(w_n266_39[2]),.din(w_n266_12[2]));
	jspl3 jspl3_w_n266_40(.douta(w_n266_40[0]),.doutb(w_n266_40[1]),.doutc(w_n266_40[2]),.din(w_n266_13[0]));
	jspl3 jspl3_w_n266_41(.douta(w_n266_41[0]),.doutb(w_n266_41[1]),.doutc(w_n266_41[2]),.din(w_n266_13[1]));
	jspl3 jspl3_w_n266_42(.douta(w_n266_42[0]),.doutb(w_n266_42[1]),.doutc(w_n266_42[2]),.din(w_n266_13[2]));
	jspl3 jspl3_w_n266_43(.douta(w_n266_43[0]),.doutb(w_n266_43[1]),.doutc(w_n266_43[2]),.din(w_n266_14[0]));
	jspl3 jspl3_w_n266_44(.douta(w_n266_44[0]),.doutb(w_n266_44[1]),.doutc(w_n266_44[2]),.din(w_n266_14[1]));
	jspl3 jspl3_w_n266_45(.douta(w_n266_45[0]),.doutb(w_n266_45[1]),.doutc(w_n266_45[2]),.din(w_n266_14[2]));
	jspl3 jspl3_w_n266_46(.douta(w_n266_46[0]),.doutb(w_n266_46[1]),.doutc(w_n266_46[2]),.din(w_n266_15[0]));
	jspl3 jspl3_w_n266_47(.douta(w_n266_47[0]),.doutb(w_n266_47[1]),.doutc(w_n266_47[2]),.din(w_n266_15[1]));
	jspl3 jspl3_w_n266_48(.douta(w_n266_48[0]),.doutb(w_n266_48[1]),.doutc(w_n266_48[2]),.din(w_n266_15[2]));
	jspl3 jspl3_w_n266_49(.douta(w_n266_49[0]),.doutb(w_n266_49[1]),.doutc(w_n266_49[2]),.din(w_n266_16[0]));
	jspl3 jspl3_w_n266_50(.douta(w_n266_50[0]),.doutb(w_n266_50[1]),.doutc(w_n266_50[2]),.din(w_n266_16[1]));
	jspl3 jspl3_w_n266_51(.douta(w_n266_51[0]),.doutb(w_n266_51[1]),.doutc(w_n266_51[2]),.din(w_n266_16[2]));
	jspl3 jspl3_w_n266_52(.douta(w_n266_52[0]),.doutb(w_n266_52[1]),.doutc(w_n266_52[2]),.din(w_n266_17[0]));
	jspl3 jspl3_w_n266_53(.douta(w_n266_53[0]),.doutb(w_n266_53[1]),.doutc(w_n266_53[2]),.din(w_n266_17[1]));
	jspl3 jspl3_w_n266_54(.douta(w_n266_54[0]),.doutb(w_n266_54[1]),.doutc(w_n266_54[2]),.din(w_n266_17[2]));
	jspl3 jspl3_w_n266_55(.douta(w_n266_55[0]),.doutb(w_n266_55[1]),.doutc(w_n266_55[2]),.din(w_n266_18[0]));
	jspl3 jspl3_w_n266_56(.douta(w_n266_56[0]),.doutb(w_n266_56[1]),.doutc(w_n266_56[2]),.din(w_n266_18[1]));
	jspl3 jspl3_w_n266_57(.douta(w_n266_57[0]),.doutb(w_n266_57[1]),.doutc(w_n266_57[2]),.din(w_n266_18[2]));
	jspl3 jspl3_w_n266_58(.douta(w_n266_58[0]),.doutb(w_n266_58[1]),.doutc(w_n266_58[2]),.din(w_n266_19[0]));
	jspl3 jspl3_w_n266_59(.douta(w_n266_59[0]),.doutb(w_n266_59[1]),.doutc(w_n266_59[2]),.din(w_n266_19[1]));
	jspl3 jspl3_w_n266_60(.douta(w_n266_60[0]),.doutb(w_n266_60[1]),.doutc(w_n266_60[2]),.din(w_n266_19[2]));
	jspl3 jspl3_w_n266_61(.douta(w_n266_61[0]),.doutb(w_n266_61[1]),.doutc(w_n266_61[2]),.din(w_n266_20[0]));
	jspl3 jspl3_w_n266_62(.douta(w_n266_62[0]),.doutb(w_n266_62[1]),.doutc(w_n266_62[2]),.din(w_n266_20[1]));
	jspl jspl_w_n266_63(.douta(w_n266_63[0]),.doutb(w_n266_63[1]),.din(w_n266_20[2]));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(n267));
	jspl3 jspl3_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.doutc(w_n269_0[2]),.din(n269));
	jspl3 jspl3_w_n269_1(.douta(w_n269_1[0]),.doutb(w_n269_1[1]),.doutc(w_n269_1[2]),.din(w_n269_0[0]));
	jspl3 jspl3_w_n269_2(.douta(w_n269_2[0]),.doutb(w_n269_2[1]),.doutc(w_n269_2[2]),.din(w_n269_0[1]));
	jspl3 jspl3_w_n269_3(.douta(w_n269_3[0]),.doutb(w_n269_3[1]),.doutc(w_n269_3[2]),.din(w_n269_0[2]));
	jspl3 jspl3_w_n269_4(.douta(w_n269_4[0]),.doutb(w_n269_4[1]),.doutc(w_n269_4[2]),.din(w_n269_1[0]));
	jspl3 jspl3_w_n269_5(.douta(w_n269_5[0]),.doutb(w_n269_5[1]),.doutc(w_n269_5[2]),.din(w_n269_1[1]));
	jspl3 jspl3_w_n269_6(.douta(w_n269_6[0]),.doutb(w_n269_6[1]),.doutc(w_n269_6[2]),.din(w_n269_1[2]));
	jspl3 jspl3_w_n269_7(.douta(w_n269_7[0]),.doutb(w_n269_7[1]),.doutc(w_n269_7[2]),.din(w_n269_2[0]));
	jspl3 jspl3_w_n269_8(.douta(w_n269_8[0]),.doutb(w_n269_8[1]),.doutc(w_n269_8[2]),.din(w_n269_2[1]));
	jspl3 jspl3_w_n269_9(.douta(w_n269_9[0]),.doutb(w_n269_9[1]),.doutc(w_n269_9[2]),.din(w_n269_2[2]));
	jspl3 jspl3_w_n269_10(.douta(w_n269_10[0]),.doutb(w_n269_10[1]),.doutc(w_n269_10[2]),.din(w_n269_3[0]));
	jspl3 jspl3_w_n269_11(.douta(w_n269_11[0]),.doutb(w_n269_11[1]),.doutc(w_n269_11[2]),.din(w_n269_3[1]));
	jspl3 jspl3_w_n269_12(.douta(w_n269_12[0]),.doutb(w_n269_12[1]),.doutc(w_n269_12[2]),.din(w_n269_3[2]));
	jspl3 jspl3_w_n269_13(.douta(w_n269_13[0]),.doutb(w_n269_13[1]),.doutc(w_n269_13[2]),.din(w_n269_4[0]));
	jspl3 jspl3_w_n269_14(.douta(w_n269_14[0]),.doutb(w_n269_14[1]),.doutc(w_n269_14[2]),.din(w_n269_4[1]));
	jspl3 jspl3_w_n269_15(.douta(w_n269_15[0]),.doutb(w_n269_15[1]),.doutc(w_n269_15[2]),.din(w_n269_4[2]));
	jspl3 jspl3_w_n269_16(.douta(w_n269_16[0]),.doutb(w_n269_16[1]),.doutc(w_n269_16[2]),.din(w_n269_5[0]));
	jspl3 jspl3_w_n269_17(.douta(w_n269_17[0]),.doutb(w_n269_17[1]),.doutc(w_n269_17[2]),.din(w_n269_5[1]));
	jspl3 jspl3_w_n269_18(.douta(w_n269_18[0]),.doutb(w_n269_18[1]),.doutc(w_n269_18[2]),.din(w_n269_5[2]));
	jspl3 jspl3_w_n269_19(.douta(w_n269_19[0]),.doutb(w_n269_19[1]),.doutc(w_n269_19[2]),.din(w_n269_6[0]));
	jspl3 jspl3_w_n269_20(.douta(w_n269_20[0]),.doutb(w_n269_20[1]),.doutc(w_n269_20[2]),.din(w_n269_6[1]));
	jspl3 jspl3_w_n269_21(.douta(w_n269_21[0]),.doutb(w_n269_21[1]),.doutc(w_n269_21[2]),.din(w_n269_6[2]));
	jspl3 jspl3_w_n269_22(.douta(w_n269_22[0]),.doutb(w_n269_22[1]),.doutc(w_n269_22[2]),.din(w_n269_7[0]));
	jspl3 jspl3_w_n269_23(.douta(w_n269_23[0]),.doutb(w_n269_23[1]),.doutc(w_n269_23[2]),.din(w_n269_7[1]));
	jspl3 jspl3_w_n269_24(.douta(w_n269_24[0]),.doutb(w_n269_24[1]),.doutc(w_n269_24[2]),.din(w_n269_7[2]));
	jspl3 jspl3_w_n269_25(.douta(w_n269_25[0]),.doutb(w_n269_25[1]),.doutc(w_n269_25[2]),.din(w_n269_8[0]));
	jspl3 jspl3_w_n269_26(.douta(w_n269_26[0]),.doutb(w_n269_26[1]),.doutc(w_n269_26[2]),.din(w_n269_8[1]));
	jspl3 jspl3_w_n269_27(.douta(w_n269_27[0]),.doutb(w_n269_27[1]),.doutc(w_n269_27[2]),.din(w_n269_8[2]));
	jspl3 jspl3_w_n269_28(.douta(w_n269_28[0]),.doutb(w_n269_28[1]),.doutc(w_n269_28[2]),.din(w_n269_9[0]));
	jspl3 jspl3_w_n269_29(.douta(w_n269_29[0]),.doutb(w_n269_29[1]),.doutc(w_n269_29[2]),.din(w_n269_9[1]));
	jspl3 jspl3_w_n269_30(.douta(w_n269_30[0]),.doutb(w_n269_30[1]),.doutc(w_n269_30[2]),.din(w_n269_9[2]));
	jspl3 jspl3_w_n269_31(.douta(w_n269_31[0]),.doutb(w_n269_31[1]),.doutc(w_n269_31[2]),.din(w_n269_10[0]));
	jspl3 jspl3_w_n269_32(.douta(w_n269_32[0]),.doutb(w_n269_32[1]),.doutc(w_n269_32[2]),.din(w_n269_10[1]));
	jspl3 jspl3_w_n269_33(.douta(w_n269_33[0]),.doutb(w_n269_33[1]),.doutc(w_n269_33[2]),.din(w_n269_10[2]));
	jspl3 jspl3_w_n269_34(.douta(w_n269_34[0]),.doutb(w_n269_34[1]),.doutc(w_n269_34[2]),.din(w_n269_11[0]));
	jspl3 jspl3_w_n269_35(.douta(w_n269_35[0]),.doutb(w_n269_35[1]),.doutc(w_n269_35[2]),.din(w_n269_11[1]));
	jspl3 jspl3_w_n269_36(.douta(w_n269_36[0]),.doutb(w_n269_36[1]),.doutc(w_n269_36[2]),.din(w_n269_11[2]));
	jspl3 jspl3_w_n269_37(.douta(w_n269_37[0]),.doutb(w_n269_37[1]),.doutc(w_n269_37[2]),.din(w_n269_12[0]));
	jspl3 jspl3_w_n269_38(.douta(w_n269_38[0]),.doutb(w_n269_38[1]),.doutc(w_n269_38[2]),.din(w_n269_12[1]));
	jspl3 jspl3_w_n269_39(.douta(w_n269_39[0]),.doutb(w_n269_39[1]),.doutc(w_n269_39[2]),.din(w_n269_12[2]));
	jspl3 jspl3_w_n269_40(.douta(w_n269_40[0]),.doutb(w_n269_40[1]),.doutc(w_n269_40[2]),.din(w_n269_13[0]));
	jspl3 jspl3_w_n269_41(.douta(w_n269_41[0]),.doutb(w_n269_41[1]),.doutc(w_n269_41[2]),.din(w_n269_13[1]));
	jspl3 jspl3_w_n269_42(.douta(w_n269_42[0]),.doutb(w_n269_42[1]),.doutc(w_n269_42[2]),.din(w_n269_13[2]));
	jspl3 jspl3_w_n269_43(.douta(w_n269_43[0]),.doutb(w_n269_43[1]),.doutc(w_n269_43[2]),.din(w_n269_14[0]));
	jspl3 jspl3_w_n269_44(.douta(w_n269_44[0]),.doutb(w_n269_44[1]),.doutc(w_n269_44[2]),.din(w_n269_14[1]));
	jspl3 jspl3_w_n269_45(.douta(w_n269_45[0]),.doutb(w_n269_45[1]),.doutc(w_n269_45[2]),.din(w_n269_14[2]));
	jspl3 jspl3_w_n269_46(.douta(w_n269_46[0]),.doutb(w_n269_46[1]),.doutc(w_n269_46[2]),.din(w_n269_15[0]));
	jspl3 jspl3_w_n269_47(.douta(w_n269_47[0]),.doutb(w_n269_47[1]),.doutc(w_n269_47[2]),.din(w_n269_15[1]));
	jspl3 jspl3_w_n269_48(.douta(w_n269_48[0]),.doutb(w_n269_48[1]),.doutc(w_n269_48[2]),.din(w_n269_15[2]));
	jspl3 jspl3_w_n269_49(.douta(w_n269_49[0]),.doutb(w_n269_49[1]),.doutc(w_n269_49[2]),.din(w_n269_16[0]));
	jspl3 jspl3_w_n269_50(.douta(w_n269_50[0]),.doutb(w_n269_50[1]),.doutc(w_n269_50[2]),.din(w_n269_16[1]));
	jspl3 jspl3_w_n269_51(.douta(w_n269_51[0]),.doutb(w_n269_51[1]),.doutc(w_n269_51[2]),.din(w_n269_16[2]));
	jspl3 jspl3_w_n269_52(.douta(w_n269_52[0]),.doutb(w_n269_52[1]),.doutc(w_n269_52[2]),.din(w_n269_17[0]));
	jspl3 jspl3_w_n269_53(.douta(w_n269_53[0]),.doutb(w_n269_53[1]),.doutc(w_n269_53[2]),.din(w_n269_17[1]));
	jspl3 jspl3_w_n269_54(.douta(w_n269_54[0]),.doutb(w_n269_54[1]),.doutc(w_n269_54[2]),.din(w_n269_17[2]));
	jspl3 jspl3_w_n269_55(.douta(w_n269_55[0]),.doutb(w_n269_55[1]),.doutc(w_n269_55[2]),.din(w_n269_18[0]));
	jspl3 jspl3_w_n269_56(.douta(w_n269_56[0]),.doutb(w_n269_56[1]),.doutc(w_n269_56[2]),.din(w_n269_18[1]));
	jspl3 jspl3_w_n269_57(.douta(w_n269_57[0]),.doutb(w_n269_57[1]),.doutc(w_n269_57[2]),.din(w_n269_18[2]));
	jspl3 jspl3_w_n269_58(.douta(w_n269_58[0]),.doutb(w_n269_58[1]),.doutc(w_n269_58[2]),.din(w_n269_19[0]));
	jspl3 jspl3_w_n269_59(.douta(w_n269_59[0]),.doutb(w_n269_59[1]),.doutc(w_n269_59[2]),.din(w_n269_19[1]));
	jspl3 jspl3_w_n269_60(.douta(w_n269_60[0]),.doutb(w_n269_60[1]),.doutc(w_n269_60[2]),.din(w_n269_19[2]));
	jspl3 jspl3_w_n269_61(.douta(w_n269_61[0]),.doutb(w_n269_61[1]),.doutc(w_n269_61[2]),.din(w_n269_20[0]));
	jspl3 jspl3_w_n269_62(.douta(w_n269_62[0]),.doutb(w_n269_62[1]),.doutc(w_n269_62[2]),.din(w_n269_20[1]));
	jspl3 jspl3_w_n269_63(.douta(w_n269_63[0]),.doutb(w_n269_63[1]),.doutc(w_n269_63[2]),.din(w_n269_20[2]));
	jspl3 jspl3_w_n269_64(.douta(w_n269_64[0]),.doutb(w_n269_64[1]),.doutc(w_n269_64[2]),.din(w_n269_21[0]));
	jspl3 jspl3_w_n269_65(.douta(w_n269_65[0]),.doutb(w_n269_65[1]),.doutc(w_n269_65[2]),.din(w_n269_21[1]));
	jspl3 jspl3_w_n269_66(.douta(w_n269_66[0]),.doutb(w_n269_66[1]),.doutc(w_n269_66[2]),.din(w_n269_21[2]));
	jspl3 jspl3_w_n269_67(.douta(w_n269_67[0]),.doutb(w_n269_67[1]),.doutc(w_n269_67[2]),.din(w_n269_22[0]));
	jspl3 jspl3_w_n269_68(.douta(w_n269_68[0]),.doutb(w_n269_68[1]),.doutc(w_n269_68[2]),.din(w_n269_22[1]));
	jspl3 jspl3_w_n269_69(.douta(w_n269_69[0]),.doutb(w_n269_69[1]),.doutc(w_n269_69[2]),.din(w_n269_22[2]));
	jspl3 jspl3_w_n269_70(.douta(w_n269_70[0]),.doutb(w_n269_70[1]),.doutc(w_n269_70[2]),.din(w_n269_23[0]));
	jspl3 jspl3_w_n269_71(.douta(w_n269_71[0]),.doutb(w_n269_71[1]),.doutc(w_n269_71[2]),.din(w_n269_23[1]));
	jspl3 jspl3_w_n269_72(.douta(w_n269_72[0]),.doutb(w_n269_72[1]),.doutc(w_n269_72[2]),.din(w_n269_23[2]));
	jspl3 jspl3_w_n269_73(.douta(w_n269_73[0]),.doutb(w_n269_73[1]),.doutc(w_n269_73[2]),.din(w_n269_24[0]));
	jspl3 jspl3_w_n269_74(.douta(w_n269_74[0]),.doutb(w_n269_74[1]),.doutc(w_n269_74[2]),.din(w_n269_24[1]));
	jspl3 jspl3_w_n269_75(.douta(w_n269_75[0]),.doutb(w_n269_75[1]),.doutc(w_n269_75[2]),.din(w_n269_24[2]));
	jspl3 jspl3_w_n269_76(.douta(w_n269_76[0]),.doutb(w_n269_76[1]),.doutc(w_n269_76[2]),.din(w_n269_25[0]));
	jspl3 jspl3_w_n269_77(.douta(w_n269_77[0]),.doutb(w_n269_77[1]),.doutc(w_n269_77[2]),.din(w_n269_25[1]));
	jspl3 jspl3_w_n269_78(.douta(w_n269_78[0]),.doutb(w_n269_78[1]),.doutc(w_n269_78[2]),.din(w_n269_25[2]));
	jspl3 jspl3_w_n269_79(.douta(w_n269_79[0]),.doutb(w_n269_79[1]),.doutc(w_n269_79[2]),.din(w_n269_26[0]));
	jspl3 jspl3_w_n269_80(.douta(w_n269_80[0]),.doutb(w_n269_80[1]),.doutc(w_n269_80[2]),.din(w_n269_26[1]));
	jspl3 jspl3_w_n269_81(.douta(w_n269_81[0]),.doutb(w_n269_81[1]),.doutc(w_n269_81[2]),.din(w_n269_26[2]));
	jspl3 jspl3_w_n269_82(.douta(w_n269_82[0]),.doutb(w_n269_82[1]),.doutc(w_n269_82[2]),.din(w_n269_27[0]));
	jspl3 jspl3_w_n269_83(.douta(w_n269_83[0]),.doutb(w_n269_83[1]),.doutc(w_n269_83[2]),.din(w_n269_27[1]));
	jspl3 jspl3_w_n269_84(.douta(w_n269_84[0]),.doutb(w_n269_84[1]),.doutc(w_n269_84[2]),.din(w_n269_27[2]));
	jspl3 jspl3_w_n269_85(.douta(w_n269_85[0]),.doutb(w_n269_85[1]),.doutc(w_n269_85[2]),.din(w_n269_28[0]));
	jspl3 jspl3_w_n269_86(.douta(w_n269_86[0]),.doutb(w_n269_86[1]),.doutc(w_n269_86[2]),.din(w_n269_28[1]));
	jspl3 jspl3_w_n269_87(.douta(w_n269_87[0]),.doutb(w_n269_87[1]),.doutc(w_n269_87[2]),.din(w_n269_28[2]));
	jspl3 jspl3_w_n269_88(.douta(w_n269_88[0]),.doutb(w_n269_88[1]),.doutc(w_n269_88[2]),.din(w_n269_29[0]));
	jspl3 jspl3_w_n269_89(.douta(w_n269_89[0]),.doutb(w_n269_89[1]),.doutc(w_n269_89[2]),.din(w_n269_29[1]));
	jspl3 jspl3_w_n269_90(.douta(w_n269_90[0]),.doutb(w_n269_90[1]),.doutc(w_n269_90[2]),.din(w_n269_29[2]));
	jspl3 jspl3_w_n269_91(.douta(w_n269_91[0]),.doutb(w_n269_91[1]),.doutc(w_n269_91[2]),.din(w_n269_30[0]));
	jspl3 jspl3_w_n269_92(.douta(w_n269_92[0]),.doutb(w_n269_92[1]),.doutc(w_n269_92[2]),.din(w_n269_30[1]));
	jspl3 jspl3_w_n269_93(.douta(w_n269_93[0]),.doutb(w_n269_93[1]),.doutc(w_n269_93[2]),.din(w_n269_30[2]));
	jspl3 jspl3_w_n269_94(.douta(w_n269_94[0]),.doutb(w_n269_94[1]),.doutc(w_n269_94[2]),.din(w_n269_31[0]));
	jspl3 jspl3_w_n269_95(.douta(w_n269_95[0]),.doutb(w_n269_95[1]),.doutc(w_n269_95[2]),.din(w_n269_31[1]));
	jspl jspl_w_n269_96(.douta(w_n269_96[0]),.doutb(w_n269_96[1]),.din(w_n269_31[2]));
	jspl3 jspl3_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.doutc(w_n270_0[2]),.din(n270));
	jspl3 jspl3_w_n270_1(.douta(w_n270_1[0]),.doutb(w_n270_1[1]),.doutc(w_n270_1[2]),.din(w_n270_0[0]));
	jspl3 jspl3_w_n270_2(.douta(w_n270_2[0]),.doutb(w_n270_2[1]),.doutc(w_n270_2[2]),.din(w_n270_0[1]));
	jspl3 jspl3_w_n270_3(.douta(w_n270_3[0]),.doutb(w_n270_3[1]),.doutc(w_n270_3[2]),.din(w_n270_0[2]));
	jspl3 jspl3_w_n270_4(.douta(w_n270_4[0]),.doutb(w_n270_4[1]),.doutc(w_n270_4[2]),.din(w_n270_1[0]));
	jspl3 jspl3_w_n270_5(.douta(w_n270_5[0]),.doutb(w_n270_5[1]),.doutc(w_n270_5[2]),.din(w_n270_1[1]));
	jspl3 jspl3_w_n270_6(.douta(w_n270_6[0]),.doutb(w_n270_6[1]),.doutc(w_n270_6[2]),.din(w_n270_1[2]));
	jspl3 jspl3_w_n270_7(.douta(w_n270_7[0]),.doutb(w_n270_7[1]),.doutc(w_n270_7[2]),.din(w_n270_2[0]));
	jspl3 jspl3_w_n270_8(.douta(w_n270_8[0]),.doutb(w_n270_8[1]),.doutc(w_n270_8[2]),.din(w_n270_2[1]));
	jspl3 jspl3_w_n270_9(.douta(w_n270_9[0]),.doutb(w_n270_9[1]),.doutc(w_n270_9[2]),.din(w_n270_2[2]));
	jspl3 jspl3_w_n270_10(.douta(w_n270_10[0]),.doutb(w_n270_10[1]),.doutc(w_n270_10[2]),.din(w_n270_3[0]));
	jspl3 jspl3_w_n270_11(.douta(w_n270_11[0]),.doutb(w_n270_11[1]),.doutc(w_n270_11[2]),.din(w_n270_3[1]));
	jspl3 jspl3_w_n270_12(.douta(w_n270_12[0]),.doutb(w_n270_12[1]),.doutc(w_n270_12[2]),.din(w_n270_3[2]));
	jspl3 jspl3_w_n270_13(.douta(w_n270_13[0]),.doutb(w_n270_13[1]),.doutc(w_n270_13[2]),.din(w_n270_4[0]));
	jspl3 jspl3_w_n270_14(.douta(w_n270_14[0]),.doutb(w_n270_14[1]),.doutc(w_n270_14[2]),.din(w_n270_4[1]));
	jspl3 jspl3_w_n270_15(.douta(w_n270_15[0]),.doutb(w_n270_15[1]),.doutc(w_n270_15[2]),.din(w_n270_4[2]));
	jspl3 jspl3_w_n270_16(.douta(w_n270_16[0]),.doutb(w_n270_16[1]),.doutc(w_n270_16[2]),.din(w_n270_5[0]));
	jspl3 jspl3_w_n270_17(.douta(w_n270_17[0]),.doutb(w_n270_17[1]),.doutc(w_n270_17[2]),.din(w_n270_5[1]));
	jspl3 jspl3_w_n270_18(.douta(w_n270_18[0]),.doutb(w_n270_18[1]),.doutc(w_n270_18[2]),.din(w_n270_5[2]));
	jspl3 jspl3_w_n270_19(.douta(w_n270_19[0]),.doutb(w_n270_19[1]),.doutc(w_n270_19[2]),.din(w_n270_6[0]));
	jspl3 jspl3_w_n270_20(.douta(w_n270_20[0]),.doutb(w_n270_20[1]),.doutc(w_n270_20[2]),.din(w_n270_6[1]));
	jspl3 jspl3_w_n270_21(.douta(w_n270_21[0]),.doutb(w_n270_21[1]),.doutc(w_n270_21[2]),.din(w_n270_6[2]));
	jspl3 jspl3_w_n270_22(.douta(w_n270_22[0]),.doutb(w_n270_22[1]),.doutc(w_n270_22[2]),.din(w_n270_7[0]));
	jspl3 jspl3_w_n270_23(.douta(w_n270_23[0]),.doutb(w_n270_23[1]),.doutc(w_n270_23[2]),.din(w_n270_7[1]));
	jspl3 jspl3_w_n270_24(.douta(w_n270_24[0]),.doutb(w_n270_24[1]),.doutc(w_n270_24[2]),.din(w_n270_7[2]));
	jspl3 jspl3_w_n270_25(.douta(w_n270_25[0]),.doutb(w_n270_25[1]),.doutc(w_n270_25[2]),.din(w_n270_8[0]));
	jspl3 jspl3_w_n270_26(.douta(w_n270_26[0]),.doutb(w_n270_26[1]),.doutc(w_n270_26[2]),.din(w_n270_8[1]));
	jspl3 jspl3_w_n270_27(.douta(w_n270_27[0]),.doutb(w_n270_27[1]),.doutc(w_n270_27[2]),.din(w_n270_8[2]));
	jspl3 jspl3_w_n270_28(.douta(w_n270_28[0]),.doutb(w_n270_28[1]),.doutc(w_n270_28[2]),.din(w_n270_9[0]));
	jspl3 jspl3_w_n270_29(.douta(w_n270_29[0]),.doutb(w_n270_29[1]),.doutc(w_n270_29[2]),.din(w_n270_9[1]));
	jspl3 jspl3_w_n270_30(.douta(w_n270_30[0]),.doutb(w_n270_30[1]),.doutc(w_n270_30[2]),.din(w_n270_9[2]));
	jspl3 jspl3_w_n270_31(.douta(w_n270_31[0]),.doutb(w_n270_31[1]),.doutc(w_n270_31[2]),.din(w_n270_10[0]));
	jspl3 jspl3_w_n270_32(.douta(w_n270_32[0]),.doutb(w_n270_32[1]),.doutc(w_n270_32[2]),.din(w_n270_10[1]));
	jspl3 jspl3_w_n270_33(.douta(w_n270_33[0]),.doutb(w_n270_33[1]),.doutc(w_n270_33[2]),.din(w_n270_10[2]));
	jspl3 jspl3_w_n270_34(.douta(w_n270_34[0]),.doutb(w_n270_34[1]),.doutc(w_n270_34[2]),.din(w_n270_11[0]));
	jspl3 jspl3_w_n270_35(.douta(w_n270_35[0]),.doutb(w_n270_35[1]),.doutc(w_n270_35[2]),.din(w_n270_11[1]));
	jspl3 jspl3_w_n270_36(.douta(w_n270_36[0]),.doutb(w_n270_36[1]),.doutc(w_n270_36[2]),.din(w_n270_11[2]));
	jspl3 jspl3_w_n270_37(.douta(w_n270_37[0]),.doutb(w_n270_37[1]),.doutc(w_n270_37[2]),.din(w_n270_12[0]));
	jspl3 jspl3_w_n270_38(.douta(w_n270_38[0]),.doutb(w_n270_38[1]),.doutc(w_n270_38[2]),.din(w_n270_12[1]));
	jspl3 jspl3_w_n270_39(.douta(w_n270_39[0]),.doutb(w_n270_39[1]),.doutc(w_n270_39[2]),.din(w_n270_12[2]));
	jspl3 jspl3_w_n270_40(.douta(w_n270_40[0]),.doutb(w_n270_40[1]),.doutc(w_n270_40[2]),.din(w_n270_13[0]));
	jspl3 jspl3_w_n270_41(.douta(w_n270_41[0]),.doutb(w_n270_41[1]),.doutc(w_n270_41[2]),.din(w_n270_13[1]));
	jspl3 jspl3_w_n270_42(.douta(w_n270_42[0]),.doutb(w_n270_42[1]),.doutc(w_n270_42[2]),.din(w_n270_13[2]));
	jspl3 jspl3_w_n270_43(.douta(w_n270_43[0]),.doutb(w_n270_43[1]),.doutc(w_n270_43[2]),.din(w_n270_14[0]));
	jspl3 jspl3_w_n270_44(.douta(w_n270_44[0]),.doutb(w_n270_44[1]),.doutc(w_n270_44[2]),.din(w_n270_14[1]));
	jspl3 jspl3_w_n270_45(.douta(w_n270_45[0]),.doutb(w_n270_45[1]),.doutc(w_n270_45[2]),.din(w_n270_14[2]));
	jspl3 jspl3_w_n270_46(.douta(w_n270_46[0]),.doutb(w_n270_46[1]),.doutc(w_n270_46[2]),.din(w_n270_15[0]));
	jspl3 jspl3_w_n270_47(.douta(w_n270_47[0]),.doutb(w_n270_47[1]),.doutc(w_n270_47[2]),.din(w_n270_15[1]));
	jspl3 jspl3_w_n270_48(.douta(w_n270_48[0]),.doutb(w_n270_48[1]),.doutc(w_n270_48[2]),.din(w_n270_15[2]));
	jspl3 jspl3_w_n270_49(.douta(w_n270_49[0]),.doutb(w_n270_49[1]),.doutc(w_n270_49[2]),.din(w_n270_16[0]));
	jspl3 jspl3_w_n270_50(.douta(w_n270_50[0]),.doutb(w_n270_50[1]),.doutc(w_n270_50[2]),.din(w_n270_16[1]));
	jspl3 jspl3_w_n270_51(.douta(w_n270_51[0]),.doutb(w_n270_51[1]),.doutc(w_n270_51[2]),.din(w_n270_16[2]));
	jspl3 jspl3_w_n270_52(.douta(w_n270_52[0]),.doutb(w_n270_52[1]),.doutc(w_n270_52[2]),.din(w_n270_17[0]));
	jspl3 jspl3_w_n270_53(.douta(w_n270_53[0]),.doutb(w_n270_53[1]),.doutc(w_n270_53[2]),.din(w_n270_17[1]));
	jspl3 jspl3_w_n270_54(.douta(w_n270_54[0]),.doutb(w_n270_54[1]),.doutc(w_n270_54[2]),.din(w_n270_17[2]));
	jspl3 jspl3_w_n270_55(.douta(w_n270_55[0]),.doutb(w_n270_55[1]),.doutc(w_n270_55[2]),.din(w_n270_18[0]));
	jspl3 jspl3_w_n270_56(.douta(w_n270_56[0]),.doutb(w_n270_56[1]),.doutc(w_n270_56[2]),.din(w_n270_18[1]));
	jspl3 jspl3_w_n270_57(.douta(w_n270_57[0]),.doutb(w_n270_57[1]),.doutc(w_n270_57[2]),.din(w_n270_18[2]));
	jspl3 jspl3_w_n270_58(.douta(w_n270_58[0]),.doutb(w_n270_58[1]),.doutc(w_n270_58[2]),.din(w_n270_19[0]));
	jspl3 jspl3_w_n270_59(.douta(w_n270_59[0]),.doutb(w_n270_59[1]),.doutc(w_n270_59[2]),.din(w_n270_19[1]));
	jspl3 jspl3_w_n270_60(.douta(w_n270_60[0]),.doutb(w_n270_60[1]),.doutc(w_n270_60[2]),.din(w_n270_19[2]));
	jspl3 jspl3_w_n270_61(.douta(w_n270_61[0]),.doutb(w_n270_61[1]),.doutc(w_n270_61[2]),.din(w_n270_20[0]));
	jspl3 jspl3_w_n270_62(.douta(w_n270_62[0]),.doutb(w_n270_62[1]),.doutc(w_n270_62[2]),.din(w_n270_20[1]));
	jspl jspl_w_n270_63(.douta(w_n270_63[0]),.doutb(w_n270_63[1]),.din(w_n270_20[2]));
	jspl jspl_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n276_0(.douta(w_n276_0[0]),.doutb(w_n276_0[1]),.din(n276));
	jspl3 jspl3_w_n279_0(.douta(w_n279_0[0]),.doutb(w_n279_0[1]),.doutc(w_n279_0[2]),.din(n279));
	jspl jspl_w_n279_1(.douta(w_n279_1[0]),.doutb(w_n279_1[1]),.din(w_n279_0[0]));
	jspl3 jspl3_w_n281_0(.douta(w_n281_0[0]),.doutb(w_n281_0[1]),.doutc(w_n281_0[2]),.din(n281));
	jspl3 jspl3_w_n281_1(.douta(w_n281_1[0]),.doutb(w_n281_1[1]),.doutc(w_n281_1[2]),.din(w_n281_0[0]));
	jspl3 jspl3_w_n281_2(.douta(w_n281_2[0]),.doutb(w_n281_2[1]),.doutc(w_n281_2[2]),.din(w_n281_0[1]));
	jspl3 jspl3_w_n281_3(.douta(w_n281_3[0]),.doutb(w_n281_3[1]),.doutc(w_n281_3[2]),.din(w_n281_0[2]));
	jspl3 jspl3_w_n281_4(.douta(w_n281_4[0]),.doutb(w_n281_4[1]),.doutc(w_n281_4[2]),.din(w_n281_1[0]));
	jspl3 jspl3_w_n281_5(.douta(w_n281_5[0]),.doutb(w_n281_5[1]),.doutc(w_n281_5[2]),.din(w_n281_1[1]));
	jspl3 jspl3_w_n281_6(.douta(w_n281_6[0]),.doutb(w_n281_6[1]),.doutc(w_n281_6[2]),.din(w_n281_1[2]));
	jspl3 jspl3_w_n281_7(.douta(w_n281_7[0]),.doutb(w_n281_7[1]),.doutc(w_n281_7[2]),.din(w_n281_2[0]));
	jspl3 jspl3_w_n281_8(.douta(w_n281_8[0]),.doutb(w_n281_8[1]),.doutc(w_n281_8[2]),.din(w_n281_2[1]));
	jspl3 jspl3_w_n281_9(.douta(w_n281_9[0]),.doutb(w_n281_9[1]),.doutc(w_n281_9[2]),.din(w_n281_2[2]));
	jspl3 jspl3_w_n281_10(.douta(w_n281_10[0]),.doutb(w_n281_10[1]),.doutc(w_n281_10[2]),.din(w_n281_3[0]));
	jspl3 jspl3_w_n281_11(.douta(w_n281_11[0]),.doutb(w_n281_11[1]),.doutc(w_n281_11[2]),.din(w_n281_3[1]));
	jspl3 jspl3_w_n281_12(.douta(w_n281_12[0]),.doutb(w_n281_12[1]),.doutc(w_n281_12[2]),.din(w_n281_3[2]));
	jspl3 jspl3_w_n281_13(.douta(w_n281_13[0]),.doutb(w_n281_13[1]),.doutc(w_n281_13[2]),.din(w_n281_4[0]));
	jspl3 jspl3_w_n281_14(.douta(w_n281_14[0]),.doutb(w_n281_14[1]),.doutc(w_n281_14[2]),.din(w_n281_4[1]));
	jspl3 jspl3_w_n281_15(.douta(w_n281_15[0]),.doutb(w_n281_15[1]),.doutc(w_n281_15[2]),.din(w_n281_4[2]));
	jspl3 jspl3_w_n281_16(.douta(w_n281_16[0]),.doutb(w_n281_16[1]),.doutc(w_n281_16[2]),.din(w_n281_5[0]));
	jspl3 jspl3_w_n281_17(.douta(w_n281_17[0]),.doutb(w_n281_17[1]),.doutc(w_n281_17[2]),.din(w_n281_5[1]));
	jspl3 jspl3_w_n281_18(.douta(w_n281_18[0]),.doutb(w_n281_18[1]),.doutc(w_n281_18[2]),.din(w_n281_5[2]));
	jspl3 jspl3_w_n281_19(.douta(w_n281_19[0]),.doutb(w_n281_19[1]),.doutc(w_n281_19[2]),.din(w_n281_6[0]));
	jspl3 jspl3_w_n281_20(.douta(w_n281_20[0]),.doutb(w_n281_20[1]),.doutc(w_n281_20[2]),.din(w_n281_6[1]));
	jspl3 jspl3_w_n281_21(.douta(w_n281_21[0]),.doutb(w_n281_21[1]),.doutc(w_n281_21[2]),.din(w_n281_6[2]));
	jspl3 jspl3_w_n281_22(.douta(w_n281_22[0]),.doutb(w_n281_22[1]),.doutc(w_n281_22[2]),.din(w_n281_7[0]));
	jspl3 jspl3_w_n281_23(.douta(w_n281_23[0]),.doutb(w_n281_23[1]),.doutc(w_n281_23[2]),.din(w_n281_7[1]));
	jspl3 jspl3_w_n281_24(.douta(w_n281_24[0]),.doutb(w_n281_24[1]),.doutc(w_n281_24[2]),.din(w_n281_7[2]));
	jspl3 jspl3_w_n281_25(.douta(w_n281_25[0]),.doutb(w_n281_25[1]),.doutc(w_n281_25[2]),.din(w_n281_8[0]));
	jspl3 jspl3_w_n281_26(.douta(w_n281_26[0]),.doutb(w_n281_26[1]),.doutc(w_n281_26[2]),.din(w_n281_8[1]));
	jspl3 jspl3_w_n281_27(.douta(w_n281_27[0]),.doutb(w_n281_27[1]),.doutc(w_n281_27[2]),.din(w_n281_8[2]));
	jspl3 jspl3_w_n281_28(.douta(w_n281_28[0]),.doutb(w_n281_28[1]),.doutc(w_n281_28[2]),.din(w_n281_9[0]));
	jspl3 jspl3_w_n281_29(.douta(w_n281_29[0]),.doutb(w_n281_29[1]),.doutc(w_n281_29[2]),.din(w_n281_9[1]));
	jspl3 jspl3_w_n281_30(.douta(w_n281_30[0]),.doutb(w_n281_30[1]),.doutc(w_n281_30[2]),.din(w_n281_9[2]));
	jspl3 jspl3_w_n281_31(.douta(w_n281_31[0]),.doutb(w_n281_31[1]),.doutc(w_n281_31[2]),.din(w_n281_10[0]));
	jspl3 jspl3_w_n281_32(.douta(w_n281_32[0]),.doutb(w_n281_32[1]),.doutc(w_n281_32[2]),.din(w_n281_10[1]));
	jspl3 jspl3_w_n281_33(.douta(w_n281_33[0]),.doutb(w_n281_33[1]),.doutc(w_n281_33[2]),.din(w_n281_10[2]));
	jspl3 jspl3_w_n281_34(.douta(w_n281_34[0]),.doutb(w_n281_34[1]),.doutc(w_n281_34[2]),.din(w_n281_11[0]));
	jspl3 jspl3_w_n281_35(.douta(w_n281_35[0]),.doutb(w_n281_35[1]),.doutc(w_n281_35[2]),.din(w_n281_11[1]));
	jspl3 jspl3_w_n281_36(.douta(w_n281_36[0]),.doutb(w_n281_36[1]),.doutc(w_n281_36[2]),.din(w_n281_11[2]));
	jspl3 jspl3_w_n281_37(.douta(w_n281_37[0]),.doutb(w_n281_37[1]),.doutc(w_n281_37[2]),.din(w_n281_12[0]));
	jspl3 jspl3_w_n281_38(.douta(w_n281_38[0]),.doutb(w_n281_38[1]),.doutc(w_n281_38[2]),.din(w_n281_12[1]));
	jspl3 jspl3_w_n281_39(.douta(w_n281_39[0]),.doutb(w_n281_39[1]),.doutc(w_n281_39[2]),.din(w_n281_12[2]));
	jspl3 jspl3_w_n281_40(.douta(w_n281_40[0]),.doutb(w_n281_40[1]),.doutc(w_n281_40[2]),.din(w_n281_13[0]));
	jspl3 jspl3_w_n281_41(.douta(w_n281_41[0]),.doutb(w_n281_41[1]),.doutc(w_n281_41[2]),.din(w_n281_13[1]));
	jspl3 jspl3_w_n281_42(.douta(w_n281_42[0]),.doutb(w_n281_42[1]),.doutc(w_n281_42[2]),.din(w_n281_13[2]));
	jspl3 jspl3_w_n281_43(.douta(w_n281_43[0]),.doutb(w_n281_43[1]),.doutc(w_n281_43[2]),.din(w_n281_14[0]));
	jspl3 jspl3_w_n281_44(.douta(w_n281_44[0]),.doutb(w_n281_44[1]),.doutc(w_n281_44[2]),.din(w_n281_14[1]));
	jspl3 jspl3_w_n281_45(.douta(w_n281_45[0]),.doutb(w_n281_45[1]),.doutc(w_n281_45[2]),.din(w_n281_14[2]));
	jspl3 jspl3_w_n281_46(.douta(w_n281_46[0]),.doutb(w_n281_46[1]),.doutc(w_n281_46[2]),.din(w_n281_15[0]));
	jspl3 jspl3_w_n281_47(.douta(w_n281_47[0]),.doutb(w_n281_47[1]),.doutc(w_n281_47[2]),.din(w_n281_15[1]));
	jspl3 jspl3_w_n281_48(.douta(w_n281_48[0]),.doutb(w_n281_48[1]),.doutc(w_n281_48[2]),.din(w_n281_15[2]));
	jspl3 jspl3_w_n281_49(.douta(w_n281_49[0]),.doutb(w_n281_49[1]),.doutc(w_n281_49[2]),.din(w_n281_16[0]));
	jspl3 jspl3_w_n281_50(.douta(w_n281_50[0]),.doutb(w_n281_50[1]),.doutc(w_n281_50[2]),.din(w_n281_16[1]));
	jspl3 jspl3_w_n281_51(.douta(w_n281_51[0]),.doutb(w_n281_51[1]),.doutc(w_n281_51[2]),.din(w_n281_16[2]));
	jspl3 jspl3_w_n281_52(.douta(w_n281_52[0]),.doutb(w_n281_52[1]),.doutc(w_n281_52[2]),.din(w_n281_17[0]));
	jspl3 jspl3_w_n281_53(.douta(w_n281_53[0]),.doutb(w_n281_53[1]),.doutc(w_n281_53[2]),.din(w_n281_17[1]));
	jspl3 jspl3_w_n281_54(.douta(w_n281_54[0]),.doutb(w_n281_54[1]),.doutc(w_n281_54[2]),.din(w_n281_17[2]));
	jspl3 jspl3_w_n281_55(.douta(w_n281_55[0]),.doutb(w_n281_55[1]),.doutc(w_n281_55[2]),.din(w_n281_18[0]));
	jspl3 jspl3_w_n281_56(.douta(w_n281_56[0]),.doutb(w_n281_56[1]),.doutc(w_n281_56[2]),.din(w_n281_18[1]));
	jspl3 jspl3_w_n281_57(.douta(w_n281_57[0]),.doutb(w_n281_57[1]),.doutc(w_n281_57[2]),.din(w_n281_18[2]));
	jspl3 jspl3_w_n281_58(.douta(w_n281_58[0]),.doutb(w_n281_58[1]),.doutc(w_n281_58[2]),.din(w_n281_19[0]));
	jspl3 jspl3_w_n281_59(.douta(w_n281_59[0]),.doutb(w_n281_59[1]),.doutc(w_n281_59[2]),.din(w_n281_19[1]));
	jspl3 jspl3_w_n281_60(.douta(w_n281_60[0]),.doutb(w_n281_60[1]),.doutc(w_n281_60[2]),.din(w_n281_19[2]));
	jspl3 jspl3_w_n281_61(.douta(w_n281_61[0]),.doutb(w_n281_61[1]),.doutc(w_n281_61[2]),.din(w_n281_20[0]));
	jspl3 jspl3_w_n281_62(.douta(w_n281_62[0]),.doutb(w_n281_62[1]),.doutc(w_n281_62[2]),.din(w_n281_20[1]));
	jspl jspl_w_n281_63(.douta(w_n281_63[0]),.doutb(w_n281_63[1]),.din(w_n281_20[2]));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n284_0(.douta(w_n284_0[0]),.doutb(w_n284_0[1]),.din(n284));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl jspl_w_n289_0(.douta(w_n289_0[0]),.doutb(w_n289_0[1]),.din(n289));
	jspl3 jspl3_w_n292_0(.douta(w_n292_0[0]),.doutb(w_n292_0[1]),.doutc(w_n292_0[2]),.din(n292));
	jspl jspl_w_n292_1(.douta(w_n292_1[0]),.doutb(w_n292_1[1]),.din(w_n292_0[0]));
	jspl3 jspl3_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.doutc(w_n295_0[2]),.din(n295));
	jspl3 jspl3_w_n295_1(.douta(w_n295_1[0]),.doutb(w_n295_1[1]),.doutc(w_n295_1[2]),.din(w_n295_0[0]));
	jspl3 jspl3_w_n295_2(.douta(w_n295_2[0]),.doutb(w_n295_2[1]),.doutc(w_n295_2[2]),.din(w_n295_0[1]));
	jspl3 jspl3_w_n295_3(.douta(w_n295_3[0]),.doutb(w_n295_3[1]),.doutc(w_n295_3[2]),.din(w_n295_0[2]));
	jspl3 jspl3_w_n295_4(.douta(w_n295_4[0]),.doutb(w_n295_4[1]),.doutc(w_n295_4[2]),.din(w_n295_1[0]));
	jspl3 jspl3_w_n295_5(.douta(w_n295_5[0]),.doutb(w_n295_5[1]),.doutc(w_n295_5[2]),.din(w_n295_1[1]));
	jspl3 jspl3_w_n295_6(.douta(w_n295_6[0]),.doutb(w_n295_6[1]),.doutc(w_n295_6[2]),.din(w_n295_1[2]));
	jspl3 jspl3_w_n295_7(.douta(w_n295_7[0]),.doutb(w_n295_7[1]),.doutc(w_n295_7[2]),.din(w_n295_2[0]));
	jspl3 jspl3_w_n295_8(.douta(w_n295_8[0]),.doutb(w_n295_8[1]),.doutc(w_n295_8[2]),.din(w_n295_2[1]));
	jspl3 jspl3_w_n295_9(.douta(w_n295_9[0]),.doutb(w_n295_9[1]),.doutc(w_n295_9[2]),.din(w_n295_2[2]));
	jspl3 jspl3_w_n295_10(.douta(w_n295_10[0]),.doutb(w_n295_10[1]),.doutc(w_n295_10[2]),.din(w_n295_3[0]));
	jspl3 jspl3_w_n295_11(.douta(w_n295_11[0]),.doutb(w_n295_11[1]),.doutc(w_n295_11[2]),.din(w_n295_3[1]));
	jspl3 jspl3_w_n295_12(.douta(w_n295_12[0]),.doutb(w_n295_12[1]),.doutc(w_n295_12[2]),.din(w_n295_3[2]));
	jspl3 jspl3_w_n295_13(.douta(w_n295_13[0]),.doutb(w_n295_13[1]),.doutc(w_n295_13[2]),.din(w_n295_4[0]));
	jspl3 jspl3_w_n295_14(.douta(w_n295_14[0]),.doutb(w_n295_14[1]),.doutc(w_n295_14[2]),.din(w_n295_4[1]));
	jspl3 jspl3_w_n295_15(.douta(w_n295_15[0]),.doutb(w_n295_15[1]),.doutc(w_n295_15[2]),.din(w_n295_4[2]));
	jspl3 jspl3_w_n295_16(.douta(w_n295_16[0]),.doutb(w_n295_16[1]),.doutc(w_n295_16[2]),.din(w_n295_5[0]));
	jspl3 jspl3_w_n295_17(.douta(w_n295_17[0]),.doutb(w_n295_17[1]),.doutc(w_n295_17[2]),.din(w_n295_5[1]));
	jspl3 jspl3_w_n295_18(.douta(w_n295_18[0]),.doutb(w_n295_18[1]),.doutc(w_n295_18[2]),.din(w_n295_5[2]));
	jspl3 jspl3_w_n295_19(.douta(w_n295_19[0]),.doutb(w_n295_19[1]),.doutc(w_n295_19[2]),.din(w_n295_6[0]));
	jspl3 jspl3_w_n295_20(.douta(w_n295_20[0]),.doutb(w_n295_20[1]),.doutc(w_n295_20[2]),.din(w_n295_6[1]));
	jspl3 jspl3_w_n295_21(.douta(w_n295_21[0]),.doutb(w_n295_21[1]),.doutc(w_n295_21[2]),.din(w_n295_6[2]));
	jspl3 jspl3_w_n295_22(.douta(w_n295_22[0]),.doutb(w_n295_22[1]),.doutc(w_n295_22[2]),.din(w_n295_7[0]));
	jspl3 jspl3_w_n295_23(.douta(w_n295_23[0]),.doutb(w_n295_23[1]),.doutc(w_n295_23[2]),.din(w_n295_7[1]));
	jspl3 jspl3_w_n295_24(.douta(w_n295_24[0]),.doutb(w_n295_24[1]),.doutc(w_n295_24[2]),.din(w_n295_7[2]));
	jspl3 jspl3_w_n295_25(.douta(w_n295_25[0]),.doutb(w_n295_25[1]),.doutc(w_n295_25[2]),.din(w_n295_8[0]));
	jspl3 jspl3_w_n295_26(.douta(w_n295_26[0]),.doutb(w_n295_26[1]),.doutc(w_n295_26[2]),.din(w_n295_8[1]));
	jspl3 jspl3_w_n295_27(.douta(w_n295_27[0]),.doutb(w_n295_27[1]),.doutc(w_n295_27[2]),.din(w_n295_8[2]));
	jspl3 jspl3_w_n295_28(.douta(w_n295_28[0]),.doutb(w_n295_28[1]),.doutc(w_n295_28[2]),.din(w_n295_9[0]));
	jspl3 jspl3_w_n295_29(.douta(w_n295_29[0]),.doutb(w_n295_29[1]),.doutc(w_n295_29[2]),.din(w_n295_9[1]));
	jspl3 jspl3_w_n295_30(.douta(w_n295_30[0]),.doutb(w_n295_30[1]),.doutc(w_n295_30[2]),.din(w_n295_9[2]));
	jspl3 jspl3_w_n295_31(.douta(w_n295_31[0]),.doutb(w_n295_31[1]),.doutc(w_n295_31[2]),.din(w_n295_10[0]));
	jspl3 jspl3_w_n295_32(.douta(w_n295_32[0]),.doutb(w_n295_32[1]),.doutc(w_n295_32[2]),.din(w_n295_10[1]));
	jspl3 jspl3_w_n295_33(.douta(w_n295_33[0]),.doutb(w_n295_33[1]),.doutc(w_n295_33[2]),.din(w_n295_10[2]));
	jspl3 jspl3_w_n295_34(.douta(w_n295_34[0]),.doutb(w_n295_34[1]),.doutc(w_n295_34[2]),.din(w_n295_11[0]));
	jspl3 jspl3_w_n295_35(.douta(w_n295_35[0]),.doutb(w_n295_35[1]),.doutc(w_n295_35[2]),.din(w_n295_11[1]));
	jspl3 jspl3_w_n295_36(.douta(w_n295_36[0]),.doutb(w_n295_36[1]),.doutc(w_n295_36[2]),.din(w_n295_11[2]));
	jspl3 jspl3_w_n295_37(.douta(w_n295_37[0]),.doutb(w_n295_37[1]),.doutc(w_n295_37[2]),.din(w_n295_12[0]));
	jspl3 jspl3_w_n295_38(.douta(w_n295_38[0]),.doutb(w_n295_38[1]),.doutc(w_n295_38[2]),.din(w_n295_12[1]));
	jspl3 jspl3_w_n295_39(.douta(w_n295_39[0]),.doutb(w_n295_39[1]),.doutc(w_n295_39[2]),.din(w_n295_12[2]));
	jspl3 jspl3_w_n295_40(.douta(w_n295_40[0]),.doutb(w_n295_40[1]),.doutc(w_n295_40[2]),.din(w_n295_13[0]));
	jspl3 jspl3_w_n295_41(.douta(w_n295_41[0]),.doutb(w_n295_41[1]),.doutc(w_n295_41[2]),.din(w_n295_13[1]));
	jspl3 jspl3_w_n295_42(.douta(w_n295_42[0]),.doutb(w_n295_42[1]),.doutc(w_n295_42[2]),.din(w_n295_13[2]));
	jspl3 jspl3_w_n295_43(.douta(w_n295_43[0]),.doutb(w_n295_43[1]),.doutc(w_n295_43[2]),.din(w_n295_14[0]));
	jspl3 jspl3_w_n295_44(.douta(w_n295_44[0]),.doutb(w_n295_44[1]),.doutc(w_n295_44[2]),.din(w_n295_14[1]));
	jspl3 jspl3_w_n295_45(.douta(w_n295_45[0]),.doutb(w_n295_45[1]),.doutc(w_n295_45[2]),.din(w_n295_14[2]));
	jspl3 jspl3_w_n295_46(.douta(w_n295_46[0]),.doutb(w_n295_46[1]),.doutc(w_n295_46[2]),.din(w_n295_15[0]));
	jspl3 jspl3_w_n295_47(.douta(w_n295_47[0]),.doutb(w_n295_47[1]),.doutc(w_n295_47[2]),.din(w_n295_15[1]));
	jspl3 jspl3_w_n295_48(.douta(w_n295_48[0]),.doutb(w_n295_48[1]),.doutc(w_n295_48[2]),.din(w_n295_15[2]));
	jspl3 jspl3_w_n295_49(.douta(w_n295_49[0]),.doutb(w_n295_49[1]),.doutc(w_n295_49[2]),.din(w_n295_16[0]));
	jspl3 jspl3_w_n295_50(.douta(w_n295_50[0]),.doutb(w_n295_50[1]),.doutc(w_n295_50[2]),.din(w_n295_16[1]));
	jspl3 jspl3_w_n295_51(.douta(w_n295_51[0]),.doutb(w_n295_51[1]),.doutc(w_n295_51[2]),.din(w_n295_16[2]));
	jspl3 jspl3_w_n295_52(.douta(w_n295_52[0]),.doutb(w_n295_52[1]),.doutc(w_n295_52[2]),.din(w_n295_17[0]));
	jspl3 jspl3_w_n295_53(.douta(w_n295_53[0]),.doutb(w_n295_53[1]),.doutc(w_n295_53[2]),.din(w_n295_17[1]));
	jspl3 jspl3_w_n295_54(.douta(w_n295_54[0]),.doutb(w_n295_54[1]),.doutc(w_n295_54[2]),.din(w_n295_17[2]));
	jspl3 jspl3_w_n295_55(.douta(w_n295_55[0]),.doutb(w_n295_55[1]),.doutc(w_n295_55[2]),.din(w_n295_18[0]));
	jspl3 jspl3_w_n295_56(.douta(w_n295_56[0]),.doutb(w_n295_56[1]),.doutc(w_n295_56[2]),.din(w_n295_18[1]));
	jspl3 jspl3_w_n295_57(.douta(w_n295_57[0]),.doutb(w_n295_57[1]),.doutc(w_n295_57[2]),.din(w_n295_18[2]));
	jspl3 jspl3_w_n295_58(.douta(w_n295_58[0]),.doutb(w_n295_58[1]),.doutc(w_n295_58[2]),.din(w_n295_19[0]));
	jspl3 jspl3_w_n295_59(.douta(w_n295_59[0]),.doutb(w_n295_59[1]),.doutc(w_n295_59[2]),.din(w_n295_19[1]));
	jspl3 jspl3_w_n295_60(.douta(w_n295_60[0]),.doutb(w_n295_60[1]),.doutc(w_n295_60[2]),.din(w_n295_19[2]));
	jspl3 jspl3_w_n295_61(.douta(w_n295_61[0]),.doutb(w_n295_61[1]),.doutc(w_n295_61[2]),.din(w_n295_20[0]));
	jspl3 jspl3_w_n295_62(.douta(w_n295_62[0]),.doutb(w_n295_62[1]),.doutc(w_n295_62[2]),.din(w_n295_20[1]));
	jspl jspl_w_n295_63(.douta(w_n295_63[0]),.doutb(w_n295_63[1]),.din(w_n295_20[2]));
	jspl jspl_w_n296_0(.douta(w_n296_0[0]),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n301_0(.douta(w_n301_0[0]),.doutb(w_n301_0[1]),.din(n301));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl3 jspl3_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.doutc(w_n306_0[2]),.din(n306));
	jspl jspl_w_n306_1(.douta(w_n306_1[0]),.doutb(w_n306_1[1]),.din(w_n306_0[0]));
	jspl3 jspl3_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.doutc(w_n308_0[2]),.din(n308));
	jspl3 jspl3_w_n308_1(.douta(w_n308_1[0]),.doutb(w_n308_1[1]),.doutc(w_n308_1[2]),.din(w_n308_0[0]));
	jspl3 jspl3_w_n308_2(.douta(w_n308_2[0]),.doutb(w_n308_2[1]),.doutc(w_n308_2[2]),.din(w_n308_0[1]));
	jspl3 jspl3_w_n308_3(.douta(w_n308_3[0]),.doutb(w_n308_3[1]),.doutc(w_n308_3[2]),.din(w_n308_0[2]));
	jspl3 jspl3_w_n308_4(.douta(w_n308_4[0]),.doutb(w_n308_4[1]),.doutc(w_n308_4[2]),.din(w_n308_1[0]));
	jspl3 jspl3_w_n308_5(.douta(w_n308_5[0]),.doutb(w_n308_5[1]),.doutc(w_n308_5[2]),.din(w_n308_1[1]));
	jspl3 jspl3_w_n308_6(.douta(w_n308_6[0]),.doutb(w_n308_6[1]),.doutc(w_n308_6[2]),.din(w_n308_1[2]));
	jspl3 jspl3_w_n308_7(.douta(w_n308_7[0]),.doutb(w_n308_7[1]),.doutc(w_n308_7[2]),.din(w_n308_2[0]));
	jspl3 jspl3_w_n308_8(.douta(w_n308_8[0]),.doutb(w_n308_8[1]),.doutc(w_n308_8[2]),.din(w_n308_2[1]));
	jspl3 jspl3_w_n308_9(.douta(w_n308_9[0]),.doutb(w_n308_9[1]),.doutc(w_n308_9[2]),.din(w_n308_2[2]));
	jspl3 jspl3_w_n308_10(.douta(w_n308_10[0]),.doutb(w_n308_10[1]),.doutc(w_n308_10[2]),.din(w_n308_3[0]));
	jspl3 jspl3_w_n308_11(.douta(w_n308_11[0]),.doutb(w_n308_11[1]),.doutc(w_n308_11[2]),.din(w_n308_3[1]));
	jspl3 jspl3_w_n308_12(.douta(w_n308_12[0]),.doutb(w_n308_12[1]),.doutc(w_n308_12[2]),.din(w_n308_3[2]));
	jspl3 jspl3_w_n308_13(.douta(w_n308_13[0]),.doutb(w_n308_13[1]),.doutc(w_n308_13[2]),.din(w_n308_4[0]));
	jspl3 jspl3_w_n308_14(.douta(w_n308_14[0]),.doutb(w_n308_14[1]),.doutc(w_n308_14[2]),.din(w_n308_4[1]));
	jspl3 jspl3_w_n308_15(.douta(w_n308_15[0]),.doutb(w_n308_15[1]),.doutc(w_n308_15[2]),.din(w_n308_4[2]));
	jspl3 jspl3_w_n308_16(.douta(w_n308_16[0]),.doutb(w_n308_16[1]),.doutc(w_n308_16[2]),.din(w_n308_5[0]));
	jspl3 jspl3_w_n308_17(.douta(w_n308_17[0]),.doutb(w_n308_17[1]),.doutc(w_n308_17[2]),.din(w_n308_5[1]));
	jspl3 jspl3_w_n308_18(.douta(w_n308_18[0]),.doutb(w_n308_18[1]),.doutc(w_n308_18[2]),.din(w_n308_5[2]));
	jspl3 jspl3_w_n308_19(.douta(w_n308_19[0]),.doutb(w_n308_19[1]),.doutc(w_n308_19[2]),.din(w_n308_6[0]));
	jspl3 jspl3_w_n308_20(.douta(w_n308_20[0]),.doutb(w_n308_20[1]),.doutc(w_n308_20[2]),.din(w_n308_6[1]));
	jspl3 jspl3_w_n308_21(.douta(w_n308_21[0]),.doutb(w_n308_21[1]),.doutc(w_n308_21[2]),.din(w_n308_6[2]));
	jspl3 jspl3_w_n308_22(.douta(w_n308_22[0]),.doutb(w_n308_22[1]),.doutc(w_n308_22[2]),.din(w_n308_7[0]));
	jspl3 jspl3_w_n308_23(.douta(w_n308_23[0]),.doutb(w_n308_23[1]),.doutc(w_n308_23[2]),.din(w_n308_7[1]));
	jspl3 jspl3_w_n308_24(.douta(w_n308_24[0]),.doutb(w_n308_24[1]),.doutc(w_n308_24[2]),.din(w_n308_7[2]));
	jspl3 jspl3_w_n308_25(.douta(w_n308_25[0]),.doutb(w_n308_25[1]),.doutc(w_n308_25[2]),.din(w_n308_8[0]));
	jspl3 jspl3_w_n308_26(.douta(w_n308_26[0]),.doutb(w_n308_26[1]),.doutc(w_n308_26[2]),.din(w_n308_8[1]));
	jspl3 jspl3_w_n308_27(.douta(w_n308_27[0]),.doutb(w_n308_27[1]),.doutc(w_n308_27[2]),.din(w_n308_8[2]));
	jspl3 jspl3_w_n308_28(.douta(w_n308_28[0]),.doutb(w_n308_28[1]),.doutc(w_n308_28[2]),.din(w_n308_9[0]));
	jspl3 jspl3_w_n308_29(.douta(w_n308_29[0]),.doutb(w_n308_29[1]),.doutc(w_n308_29[2]),.din(w_n308_9[1]));
	jspl3 jspl3_w_n308_30(.douta(w_n308_30[0]),.doutb(w_n308_30[1]),.doutc(w_n308_30[2]),.din(w_n308_9[2]));
	jspl3 jspl3_w_n308_31(.douta(w_n308_31[0]),.doutb(w_n308_31[1]),.doutc(w_n308_31[2]),.din(w_n308_10[0]));
	jspl3 jspl3_w_n308_32(.douta(w_n308_32[0]),.doutb(w_n308_32[1]),.doutc(w_n308_32[2]),.din(w_n308_10[1]));
	jspl3 jspl3_w_n308_33(.douta(w_n308_33[0]),.doutb(w_n308_33[1]),.doutc(w_n308_33[2]),.din(w_n308_10[2]));
	jspl3 jspl3_w_n308_34(.douta(w_n308_34[0]),.doutb(w_n308_34[1]),.doutc(w_n308_34[2]),.din(w_n308_11[0]));
	jspl3 jspl3_w_n308_35(.douta(w_n308_35[0]),.doutb(w_n308_35[1]),.doutc(w_n308_35[2]),.din(w_n308_11[1]));
	jspl3 jspl3_w_n308_36(.douta(w_n308_36[0]),.doutb(w_n308_36[1]),.doutc(w_n308_36[2]),.din(w_n308_11[2]));
	jspl3 jspl3_w_n308_37(.douta(w_n308_37[0]),.doutb(w_n308_37[1]),.doutc(w_n308_37[2]),.din(w_n308_12[0]));
	jspl3 jspl3_w_n308_38(.douta(w_n308_38[0]),.doutb(w_n308_38[1]),.doutc(w_n308_38[2]),.din(w_n308_12[1]));
	jspl3 jspl3_w_n308_39(.douta(w_n308_39[0]),.doutb(w_n308_39[1]),.doutc(w_n308_39[2]),.din(w_n308_12[2]));
	jspl3 jspl3_w_n308_40(.douta(w_n308_40[0]),.doutb(w_n308_40[1]),.doutc(w_n308_40[2]),.din(w_n308_13[0]));
	jspl3 jspl3_w_n308_41(.douta(w_n308_41[0]),.doutb(w_n308_41[1]),.doutc(w_n308_41[2]),.din(w_n308_13[1]));
	jspl3 jspl3_w_n308_42(.douta(w_n308_42[0]),.doutb(w_n308_42[1]),.doutc(w_n308_42[2]),.din(w_n308_13[2]));
	jspl3 jspl3_w_n308_43(.douta(w_n308_43[0]),.doutb(w_n308_43[1]),.doutc(w_n308_43[2]),.din(w_n308_14[0]));
	jspl3 jspl3_w_n308_44(.douta(w_n308_44[0]),.doutb(w_n308_44[1]),.doutc(w_n308_44[2]),.din(w_n308_14[1]));
	jspl3 jspl3_w_n308_45(.douta(w_n308_45[0]),.doutb(w_n308_45[1]),.doutc(w_n308_45[2]),.din(w_n308_14[2]));
	jspl3 jspl3_w_n308_46(.douta(w_n308_46[0]),.doutb(w_n308_46[1]),.doutc(w_n308_46[2]),.din(w_n308_15[0]));
	jspl3 jspl3_w_n308_47(.douta(w_n308_47[0]),.doutb(w_n308_47[1]),.doutc(w_n308_47[2]),.din(w_n308_15[1]));
	jspl3 jspl3_w_n308_48(.douta(w_n308_48[0]),.doutb(w_n308_48[1]),.doutc(w_n308_48[2]),.din(w_n308_15[2]));
	jspl3 jspl3_w_n308_49(.douta(w_n308_49[0]),.doutb(w_n308_49[1]),.doutc(w_n308_49[2]),.din(w_n308_16[0]));
	jspl3 jspl3_w_n308_50(.douta(w_n308_50[0]),.doutb(w_n308_50[1]),.doutc(w_n308_50[2]),.din(w_n308_16[1]));
	jspl3 jspl3_w_n308_51(.douta(w_n308_51[0]),.doutb(w_n308_51[1]),.doutc(w_n308_51[2]),.din(w_n308_16[2]));
	jspl3 jspl3_w_n308_52(.douta(w_n308_52[0]),.doutb(w_n308_52[1]),.doutc(w_n308_52[2]),.din(w_n308_17[0]));
	jspl3 jspl3_w_n308_53(.douta(w_n308_53[0]),.doutb(w_n308_53[1]),.doutc(w_n308_53[2]),.din(w_n308_17[1]));
	jspl3 jspl3_w_n308_54(.douta(w_n308_54[0]),.doutb(w_n308_54[1]),.doutc(w_n308_54[2]),.din(w_n308_17[2]));
	jspl3 jspl3_w_n308_55(.douta(w_n308_55[0]),.doutb(w_n308_55[1]),.doutc(w_n308_55[2]),.din(w_n308_18[0]));
	jspl3 jspl3_w_n308_56(.douta(w_n308_56[0]),.doutb(w_n308_56[1]),.doutc(w_n308_56[2]),.din(w_n308_18[1]));
	jspl3 jspl3_w_n308_57(.douta(w_n308_57[0]),.doutb(w_n308_57[1]),.doutc(w_n308_57[2]),.din(w_n308_18[2]));
	jspl3 jspl3_w_n308_58(.douta(w_n308_58[0]),.doutb(w_n308_58[1]),.doutc(w_n308_58[2]),.din(w_n308_19[0]));
	jspl3 jspl3_w_n308_59(.douta(w_n308_59[0]),.doutb(w_n308_59[1]),.doutc(w_n308_59[2]),.din(w_n308_19[1]));
	jspl3 jspl3_w_n308_60(.douta(w_n308_60[0]),.doutb(w_n308_60[1]),.doutc(w_n308_60[2]),.din(w_n308_19[2]));
	jspl3 jspl3_w_n308_61(.douta(w_n308_61[0]),.doutb(w_n308_61[1]),.doutc(w_n308_61[2]),.din(w_n308_20[0]));
	jspl3 jspl3_w_n308_62(.douta(w_n308_62[0]),.doutb(w_n308_62[1]),.doutc(w_n308_62[2]),.din(w_n308_20[1]));
	jspl jspl_w_n308_63(.douta(w_n308_63[0]),.doutb(w_n308_63[1]),.din(w_n308_20[2]));
	jspl jspl_w_n309_0(.douta(w_n309_0[0]),.doutb(w_n309_0[1]),.din(n309));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.din(n314));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl3 jspl3_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.doutc(w_n319_0[2]),.din(n319));
	jspl jspl_w_n319_1(.douta(w_n319_1[0]),.doutb(w_n319_1[1]),.din(w_n319_0[0]));
	jspl3 jspl3_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.doutc(w_n322_0[2]),.din(n322));
	jspl jspl_w_n322_1(.douta(w_n322_1[0]),.doutb(w_n322_1[1]),.din(w_n322_0[0]));
	jspl3 jspl3_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.doutc(w_n323_0[2]),.din(n323));
	jspl3 jspl3_w_n323_1(.douta(w_n323_1[0]),.doutb(w_n323_1[1]),.doutc(w_n323_1[2]),.din(w_n323_0[0]));
	jspl3 jspl3_w_n323_2(.douta(w_n323_2[0]),.doutb(w_n323_2[1]),.doutc(w_n323_2[2]),.din(w_n323_0[1]));
	jspl3 jspl3_w_n323_3(.douta(w_n323_3[0]),.doutb(w_n323_3[1]),.doutc(w_n323_3[2]),.din(w_n323_0[2]));
	jspl3 jspl3_w_n323_4(.douta(w_n323_4[0]),.doutb(w_n323_4[1]),.doutc(w_n323_4[2]),.din(w_n323_1[0]));
	jspl3 jspl3_w_n323_5(.douta(w_n323_5[0]),.doutb(w_n323_5[1]),.doutc(w_n323_5[2]),.din(w_n323_1[1]));
	jspl3 jspl3_w_n323_6(.douta(w_n323_6[0]),.doutb(w_n323_6[1]),.doutc(w_n323_6[2]),.din(w_n323_1[2]));
	jspl3 jspl3_w_n323_7(.douta(w_n323_7[0]),.doutb(w_n323_7[1]),.doutc(w_n323_7[2]),.din(w_n323_2[0]));
	jspl3 jspl3_w_n323_8(.douta(w_n323_8[0]),.doutb(w_n323_8[1]),.doutc(w_n323_8[2]),.din(w_n323_2[1]));
	jspl3 jspl3_w_n323_9(.douta(w_n323_9[0]),.doutb(w_n323_9[1]),.doutc(w_n323_9[2]),.din(w_n323_2[2]));
	jspl3 jspl3_w_n323_10(.douta(w_n323_10[0]),.doutb(w_n323_10[1]),.doutc(w_n323_10[2]),.din(w_n323_3[0]));
	jspl3 jspl3_w_n323_11(.douta(w_n323_11[0]),.doutb(w_n323_11[1]),.doutc(w_n323_11[2]),.din(w_n323_3[1]));
	jspl3 jspl3_w_n323_12(.douta(w_n323_12[0]),.doutb(w_n323_12[1]),.doutc(w_n323_12[2]),.din(w_n323_3[2]));
	jspl3 jspl3_w_n323_13(.douta(w_n323_13[0]),.doutb(w_n323_13[1]),.doutc(w_n323_13[2]),.din(w_n323_4[0]));
	jspl3 jspl3_w_n323_14(.douta(w_n323_14[0]),.doutb(w_n323_14[1]),.doutc(w_n323_14[2]),.din(w_n323_4[1]));
	jspl3 jspl3_w_n323_15(.douta(w_n323_15[0]),.doutb(w_n323_15[1]),.doutc(w_n323_15[2]),.din(w_n323_4[2]));
	jspl3 jspl3_w_n323_16(.douta(w_n323_16[0]),.doutb(w_n323_16[1]),.doutc(w_n323_16[2]),.din(w_n323_5[0]));
	jspl3 jspl3_w_n323_17(.douta(w_n323_17[0]),.doutb(w_n323_17[1]),.doutc(w_n323_17[2]),.din(w_n323_5[1]));
	jspl3 jspl3_w_n323_18(.douta(w_n323_18[0]),.doutb(w_n323_18[1]),.doutc(w_n323_18[2]),.din(w_n323_5[2]));
	jspl3 jspl3_w_n323_19(.douta(w_n323_19[0]),.doutb(w_n323_19[1]),.doutc(w_n323_19[2]),.din(w_n323_6[0]));
	jspl3 jspl3_w_n323_20(.douta(w_n323_20[0]),.doutb(w_n323_20[1]),.doutc(w_n323_20[2]),.din(w_n323_6[1]));
	jspl3 jspl3_w_n323_21(.douta(w_n323_21[0]),.doutb(w_n323_21[1]),.doutc(w_n323_21[2]),.din(w_n323_6[2]));
	jspl3 jspl3_w_n323_22(.douta(w_n323_22[0]),.doutb(w_n323_22[1]),.doutc(w_n323_22[2]),.din(w_n323_7[0]));
	jspl3 jspl3_w_n323_23(.douta(w_n323_23[0]),.doutb(w_n323_23[1]),.doutc(w_n323_23[2]),.din(w_n323_7[1]));
	jspl3 jspl3_w_n323_24(.douta(w_n323_24[0]),.doutb(w_n323_24[1]),.doutc(w_n323_24[2]),.din(w_n323_7[2]));
	jspl3 jspl3_w_n323_25(.douta(w_n323_25[0]),.doutb(w_n323_25[1]),.doutc(w_n323_25[2]),.din(w_n323_8[0]));
	jspl3 jspl3_w_n323_26(.douta(w_n323_26[0]),.doutb(w_n323_26[1]),.doutc(w_n323_26[2]),.din(w_n323_8[1]));
	jspl3 jspl3_w_n323_27(.douta(w_n323_27[0]),.doutb(w_n323_27[1]),.doutc(w_n323_27[2]),.din(w_n323_8[2]));
	jspl3 jspl3_w_n323_28(.douta(w_n323_28[0]),.doutb(w_n323_28[1]),.doutc(w_n323_28[2]),.din(w_n323_9[0]));
	jspl3 jspl3_w_n323_29(.douta(w_n323_29[0]),.doutb(w_n323_29[1]),.doutc(w_n323_29[2]),.din(w_n323_9[1]));
	jspl3 jspl3_w_n323_30(.douta(w_n323_30[0]),.doutb(w_n323_30[1]),.doutc(w_n323_30[2]),.din(w_n323_9[2]));
	jspl3 jspl3_w_n323_31(.douta(w_n323_31[0]),.doutb(w_n323_31[1]),.doutc(w_n323_31[2]),.din(w_n323_10[0]));
	jspl3 jspl3_w_n323_32(.douta(w_n323_32[0]),.doutb(w_n323_32[1]),.doutc(w_n323_32[2]),.din(w_n323_10[1]));
	jspl3 jspl3_w_n323_33(.douta(w_n323_33[0]),.doutb(w_n323_33[1]),.doutc(w_n323_33[2]),.din(w_n323_10[2]));
	jspl3 jspl3_w_n323_34(.douta(w_n323_34[0]),.doutb(w_n323_34[1]),.doutc(w_n323_34[2]),.din(w_n323_11[0]));
	jspl3 jspl3_w_n323_35(.douta(w_n323_35[0]),.doutb(w_n323_35[1]),.doutc(w_n323_35[2]),.din(w_n323_11[1]));
	jspl3 jspl3_w_n323_36(.douta(w_n323_36[0]),.doutb(w_n323_36[1]),.doutc(w_n323_36[2]),.din(w_n323_11[2]));
	jspl3 jspl3_w_n323_37(.douta(w_n323_37[0]),.doutb(w_n323_37[1]),.doutc(w_n323_37[2]),.din(w_n323_12[0]));
	jspl3 jspl3_w_n323_38(.douta(w_n323_38[0]),.doutb(w_n323_38[1]),.doutc(w_n323_38[2]),.din(w_n323_12[1]));
	jspl3 jspl3_w_n323_39(.douta(w_n323_39[0]),.doutb(w_n323_39[1]),.doutc(w_n323_39[2]),.din(w_n323_12[2]));
	jspl3 jspl3_w_n323_40(.douta(w_n323_40[0]),.doutb(w_n323_40[1]),.doutc(w_n323_40[2]),.din(w_n323_13[0]));
	jspl3 jspl3_w_n323_41(.douta(w_n323_41[0]),.doutb(w_n323_41[1]),.doutc(w_n323_41[2]),.din(w_n323_13[1]));
	jspl3 jspl3_w_n323_42(.douta(w_n323_42[0]),.doutb(w_n323_42[1]),.doutc(w_n323_42[2]),.din(w_n323_13[2]));
	jspl3 jspl3_w_n323_43(.douta(w_n323_43[0]),.doutb(w_n323_43[1]),.doutc(w_n323_43[2]),.din(w_n323_14[0]));
	jspl3 jspl3_w_n323_44(.douta(w_n323_44[0]),.doutb(w_n323_44[1]),.doutc(w_n323_44[2]),.din(w_n323_14[1]));
	jspl3 jspl3_w_n323_45(.douta(w_n323_45[0]),.doutb(w_n323_45[1]),.doutc(w_n323_45[2]),.din(w_n323_14[2]));
	jspl3 jspl3_w_n323_46(.douta(w_n323_46[0]),.doutb(w_n323_46[1]),.doutc(w_n323_46[2]),.din(w_n323_15[0]));
	jspl3 jspl3_w_n323_47(.douta(w_n323_47[0]),.doutb(w_n323_47[1]),.doutc(w_n323_47[2]),.din(w_n323_15[1]));
	jspl3 jspl3_w_n323_48(.douta(w_n323_48[0]),.doutb(w_n323_48[1]),.doutc(w_n323_48[2]),.din(w_n323_15[2]));
	jspl3 jspl3_w_n323_49(.douta(w_n323_49[0]),.doutb(w_n323_49[1]),.doutc(w_n323_49[2]),.din(w_n323_16[0]));
	jspl3 jspl3_w_n323_50(.douta(w_n323_50[0]),.doutb(w_n323_50[1]),.doutc(w_n323_50[2]),.din(w_n323_16[1]));
	jspl3 jspl3_w_n323_51(.douta(w_n323_51[0]),.doutb(w_n323_51[1]),.doutc(w_n323_51[2]),.din(w_n323_16[2]));
	jspl3 jspl3_w_n323_52(.douta(w_n323_52[0]),.doutb(w_n323_52[1]),.doutc(w_n323_52[2]),.din(w_n323_17[0]));
	jspl3 jspl3_w_n323_53(.douta(w_n323_53[0]),.doutb(w_n323_53[1]),.doutc(w_n323_53[2]),.din(w_n323_17[1]));
	jspl3 jspl3_w_n323_54(.douta(w_n323_54[0]),.doutb(w_n323_54[1]),.doutc(w_n323_54[2]),.din(w_n323_17[2]));
	jspl3 jspl3_w_n323_55(.douta(w_n323_55[0]),.doutb(w_n323_55[1]),.doutc(w_n323_55[2]),.din(w_n323_18[0]));
	jspl3 jspl3_w_n323_56(.douta(w_n323_56[0]),.doutb(w_n323_56[1]),.doutc(w_n323_56[2]),.din(w_n323_18[1]));
	jspl3 jspl3_w_n323_57(.douta(w_n323_57[0]),.doutb(w_n323_57[1]),.doutc(w_n323_57[2]),.din(w_n323_18[2]));
	jspl3 jspl3_w_n323_58(.douta(w_n323_58[0]),.doutb(w_n323_58[1]),.doutc(w_n323_58[2]),.din(w_n323_19[0]));
	jspl3 jspl3_w_n323_59(.douta(w_n323_59[0]),.doutb(w_n323_59[1]),.doutc(w_n323_59[2]),.din(w_n323_19[1]));
	jspl3 jspl3_w_n323_60(.douta(w_n323_60[0]),.doutb(w_n323_60[1]),.doutc(w_n323_60[2]),.din(w_n323_19[2]));
	jspl3 jspl3_w_n323_61(.douta(w_n323_61[0]),.doutb(w_n323_61[1]),.doutc(w_n323_61[2]),.din(w_n323_20[0]));
	jspl3 jspl3_w_n323_62(.douta(w_n323_62[0]),.doutb(w_n323_62[1]),.doutc(w_n323_62[2]),.din(w_n323_20[1]));
	jspl jspl_w_n323_63(.douta(w_n323_63[0]),.doutb(w_n323_63[1]),.din(w_n323_20[2]));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(n327));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(n330));
	jspl jspl_w_n332_0(.douta(w_n332_0[0]),.doutb(w_n332_0[1]),.din(n332));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl jspl_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.din(w_n335_0[0]));
	jspl jspl_w_n337_0(.douta(w_n337_0[0]),.doutb(w_n337_0[1]),.din(n337));
	jspl jspl_w_n339_0(.douta(w_n339_0[0]),.doutb(w_n339_0[1]),.din(n339));
	jspl jspl_w_n342_0(.douta(w_n342_0[0]),.doutb(w_n342_0[1]),.din(n342));
	jspl jspl_w_n344_0(.douta(w_n344_0[0]),.doutb(w_n344_0[1]),.din(n344));
	jspl3 jspl3_w_n347_0(.douta(w_n347_0[0]),.doutb(w_n347_0[1]),.doutc(w_n347_0[2]),.din(n347));
	jspl jspl_w_n347_1(.douta(w_n347_1[0]),.doutb(w_n347_1[1]),.din(w_n347_0[0]));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n352_0(.douta(w_n352_0[0]),.doutb(w_n352_0[1]),.din(n352));
	jspl jspl_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl3 jspl3_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.doutc(w_n360_0[2]),.din(n360));
	jspl jspl_w_n360_1(.douta(w_n360_1[0]),.doutb(w_n360_1[1]),.din(w_n360_0[0]));
	jspl jspl_w_n362_0(.douta(w_n362_0[0]),.doutb(w_n362_0[1]),.din(n362));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.din(n367));
	jspl jspl_w_n369_0(.douta(w_n369_0[0]),.doutb(w_n369_0[1]),.din(n369));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.doutc(w_n372_0[2]),.din(n372));
	jspl jspl_w_n372_1(.douta(w_n372_1[0]),.doutb(w_n372_1[1]),.din(w_n372_0[0]));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl jspl_w_n375_1(.douta(w_n375_1[0]),.doutb(w_n375_1[1]),.din(w_n375_0[0]));
	jspl jspl_w_n376_0(.douta(w_n376_0[0]),.doutb(w_n376_0[1]),.din(n376));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_n377_0[2]),.din(n377));
	jspl3 jspl3_w_n377_1(.douta(w_n377_1[0]),.doutb(w_n377_1[1]),.doutc(w_n377_1[2]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n377_2(.douta(w_n377_2[0]),.doutb(w_n377_2[1]),.doutc(w_n377_2[2]),.din(w_n377_0[1]));
	jspl3 jspl3_w_n377_3(.douta(w_n377_3[0]),.doutb(w_n377_3[1]),.doutc(w_n377_3[2]),.din(w_n377_0[2]));
	jspl3 jspl3_w_n377_4(.douta(w_n377_4[0]),.doutb(w_n377_4[1]),.doutc(w_n377_4[2]),.din(w_n377_1[0]));
	jspl3 jspl3_w_n377_5(.douta(w_n377_5[0]),.doutb(w_n377_5[1]),.doutc(w_n377_5[2]),.din(w_n377_1[1]));
	jspl3 jspl3_w_n377_6(.douta(w_n377_6[0]),.doutb(w_n377_6[1]),.doutc(w_n377_6[2]),.din(w_n377_1[2]));
	jspl3 jspl3_w_n377_7(.douta(w_n377_7[0]),.doutb(w_n377_7[1]),.doutc(w_n377_7[2]),.din(w_n377_2[0]));
	jspl3 jspl3_w_n377_8(.douta(w_n377_8[0]),.doutb(w_n377_8[1]),.doutc(w_n377_8[2]),.din(w_n377_2[1]));
	jspl3 jspl3_w_n377_9(.douta(w_n377_9[0]),.doutb(w_n377_9[1]),.doutc(w_n377_9[2]),.din(w_n377_2[2]));
	jspl3 jspl3_w_n377_10(.douta(w_n377_10[0]),.doutb(w_n377_10[1]),.doutc(w_n377_10[2]),.din(w_n377_3[0]));
	jspl3 jspl3_w_n377_11(.douta(w_n377_11[0]),.doutb(w_n377_11[1]),.doutc(w_n377_11[2]),.din(w_n377_3[1]));
	jspl3 jspl3_w_n377_12(.douta(w_n377_12[0]),.doutb(w_n377_12[1]),.doutc(w_n377_12[2]),.din(w_n377_3[2]));
	jspl3 jspl3_w_n377_13(.douta(w_n377_13[0]),.doutb(w_n377_13[1]),.doutc(w_n377_13[2]),.din(w_n377_4[0]));
	jspl3 jspl3_w_n377_14(.douta(w_n377_14[0]),.doutb(w_n377_14[1]),.doutc(w_n377_14[2]),.din(w_n377_4[1]));
	jspl3 jspl3_w_n377_15(.douta(w_n377_15[0]),.doutb(w_n377_15[1]),.doutc(w_n377_15[2]),.din(w_n377_4[2]));
	jspl3 jspl3_w_n377_16(.douta(w_n377_16[0]),.doutb(w_n377_16[1]),.doutc(w_n377_16[2]),.din(w_n377_5[0]));
	jspl3 jspl3_w_n377_17(.douta(w_n377_17[0]),.doutb(w_n377_17[1]),.doutc(w_n377_17[2]),.din(w_n377_5[1]));
	jspl3 jspl3_w_n377_18(.douta(w_n377_18[0]),.doutb(w_n377_18[1]),.doutc(w_n377_18[2]),.din(w_n377_5[2]));
	jspl3 jspl3_w_n377_19(.douta(w_n377_19[0]),.doutb(w_n377_19[1]),.doutc(w_n377_19[2]),.din(w_n377_6[0]));
	jspl3 jspl3_w_n377_20(.douta(w_n377_20[0]),.doutb(w_n377_20[1]),.doutc(w_n377_20[2]),.din(w_n377_6[1]));
	jspl3 jspl3_w_n377_21(.douta(w_n377_21[0]),.doutb(w_n377_21[1]),.doutc(w_n377_21[2]),.din(w_n377_6[2]));
	jspl3 jspl3_w_n377_22(.douta(w_n377_22[0]),.doutb(w_n377_22[1]),.doutc(w_n377_22[2]),.din(w_n377_7[0]));
	jspl3 jspl3_w_n377_23(.douta(w_n377_23[0]),.doutb(w_n377_23[1]),.doutc(w_n377_23[2]),.din(w_n377_7[1]));
	jspl3 jspl3_w_n377_24(.douta(w_n377_24[0]),.doutb(w_n377_24[1]),.doutc(w_n377_24[2]),.din(w_n377_7[2]));
	jspl3 jspl3_w_n377_25(.douta(w_n377_25[0]),.doutb(w_n377_25[1]),.doutc(w_n377_25[2]),.din(w_n377_8[0]));
	jspl3 jspl3_w_n377_26(.douta(w_n377_26[0]),.doutb(w_n377_26[1]),.doutc(w_n377_26[2]),.din(w_n377_8[1]));
	jspl3 jspl3_w_n377_27(.douta(w_n377_27[0]),.doutb(w_n377_27[1]),.doutc(w_n377_27[2]),.din(w_n377_8[2]));
	jspl3 jspl3_w_n377_28(.douta(w_n377_28[0]),.doutb(w_n377_28[1]),.doutc(w_n377_28[2]),.din(w_n377_9[0]));
	jspl3 jspl3_w_n377_29(.douta(w_n377_29[0]),.doutb(w_n377_29[1]),.doutc(w_n377_29[2]),.din(w_n377_9[1]));
	jspl3 jspl3_w_n377_30(.douta(w_n377_30[0]),.doutb(w_n377_30[1]),.doutc(w_n377_30[2]),.din(w_n377_9[2]));
	jspl3 jspl3_w_n377_31(.douta(w_n377_31[0]),.doutb(w_n377_31[1]),.doutc(w_n377_31[2]),.din(w_n377_10[0]));
	jspl3 jspl3_w_n377_32(.douta(w_n377_32[0]),.doutb(w_n377_32[1]),.doutc(w_n377_32[2]),.din(w_n377_10[1]));
	jspl3 jspl3_w_n377_33(.douta(w_n377_33[0]),.doutb(w_n377_33[1]),.doutc(w_n377_33[2]),.din(w_n377_10[2]));
	jspl3 jspl3_w_n377_34(.douta(w_n377_34[0]),.doutb(w_n377_34[1]),.doutc(w_n377_34[2]),.din(w_n377_11[0]));
	jspl3 jspl3_w_n377_35(.douta(w_n377_35[0]),.doutb(w_n377_35[1]),.doutc(w_n377_35[2]),.din(w_n377_11[1]));
	jspl3 jspl3_w_n377_36(.douta(w_n377_36[0]),.doutb(w_n377_36[1]),.doutc(w_n377_36[2]),.din(w_n377_11[2]));
	jspl3 jspl3_w_n377_37(.douta(w_n377_37[0]),.doutb(w_n377_37[1]),.doutc(w_n377_37[2]),.din(w_n377_12[0]));
	jspl3 jspl3_w_n377_38(.douta(w_n377_38[0]),.doutb(w_n377_38[1]),.doutc(w_n377_38[2]),.din(w_n377_12[1]));
	jspl3 jspl3_w_n377_39(.douta(w_n377_39[0]),.doutb(w_n377_39[1]),.doutc(w_n377_39[2]),.din(w_n377_12[2]));
	jspl3 jspl3_w_n377_40(.douta(w_n377_40[0]),.doutb(w_n377_40[1]),.doutc(w_n377_40[2]),.din(w_n377_13[0]));
	jspl3 jspl3_w_n377_41(.douta(w_n377_41[0]),.doutb(w_n377_41[1]),.doutc(w_n377_41[2]),.din(w_n377_13[1]));
	jspl3 jspl3_w_n377_42(.douta(w_n377_42[0]),.doutb(w_n377_42[1]),.doutc(w_n377_42[2]),.din(w_n377_13[2]));
	jspl3 jspl3_w_n377_43(.douta(w_n377_43[0]),.doutb(w_n377_43[1]),.doutc(w_n377_43[2]),.din(w_n377_14[0]));
	jspl3 jspl3_w_n377_44(.douta(w_n377_44[0]),.doutb(w_n377_44[1]),.doutc(w_n377_44[2]),.din(w_n377_14[1]));
	jspl3 jspl3_w_n377_45(.douta(w_n377_45[0]),.doutb(w_n377_45[1]),.doutc(w_n377_45[2]),.din(w_n377_14[2]));
	jspl3 jspl3_w_n377_46(.douta(w_n377_46[0]),.doutb(w_n377_46[1]),.doutc(w_n377_46[2]),.din(w_n377_15[0]));
	jspl3 jspl3_w_n377_47(.douta(w_n377_47[0]),.doutb(w_n377_47[1]),.doutc(w_n377_47[2]),.din(w_n377_15[1]));
	jspl3 jspl3_w_n377_48(.douta(w_n377_48[0]),.doutb(w_n377_48[1]),.doutc(w_n377_48[2]),.din(w_n377_15[2]));
	jspl3 jspl3_w_n377_49(.douta(w_n377_49[0]),.doutb(w_n377_49[1]),.doutc(w_n377_49[2]),.din(w_n377_16[0]));
	jspl3 jspl3_w_n377_50(.douta(w_n377_50[0]),.doutb(w_n377_50[1]),.doutc(w_n377_50[2]),.din(w_n377_16[1]));
	jspl3 jspl3_w_n377_51(.douta(w_n377_51[0]),.doutb(w_n377_51[1]),.doutc(w_n377_51[2]),.din(w_n377_16[2]));
	jspl3 jspl3_w_n377_52(.douta(w_n377_52[0]),.doutb(w_n377_52[1]),.doutc(w_n377_52[2]),.din(w_n377_17[0]));
	jspl3 jspl3_w_n377_53(.douta(w_n377_53[0]),.doutb(w_n377_53[1]),.doutc(w_n377_53[2]),.din(w_n377_17[1]));
	jspl3 jspl3_w_n377_54(.douta(w_n377_54[0]),.doutb(w_n377_54[1]),.doutc(w_n377_54[2]),.din(w_n377_17[2]));
	jspl3 jspl3_w_n377_55(.douta(w_n377_55[0]),.doutb(w_n377_55[1]),.doutc(w_n377_55[2]),.din(w_n377_18[0]));
	jspl3 jspl3_w_n377_56(.douta(w_n377_56[0]),.doutb(w_n377_56[1]),.doutc(w_n377_56[2]),.din(w_n377_18[1]));
	jspl3 jspl3_w_n377_57(.douta(w_n377_57[0]),.doutb(w_n377_57[1]),.doutc(w_n377_57[2]),.din(w_n377_18[2]));
	jspl3 jspl3_w_n377_58(.douta(w_n377_58[0]),.doutb(w_n377_58[1]),.doutc(w_n377_58[2]),.din(w_n377_19[0]));
	jspl3 jspl3_w_n377_59(.douta(w_n377_59[0]),.doutb(w_n377_59[1]),.doutc(w_n377_59[2]),.din(w_n377_19[1]));
	jspl3 jspl3_w_n377_60(.douta(w_n377_60[0]),.doutb(w_n377_60[1]),.doutc(w_n377_60[2]),.din(w_n377_19[2]));
	jspl3 jspl3_w_n377_61(.douta(w_n377_61[0]),.doutb(w_n377_61[1]),.doutc(w_n377_61[2]),.din(w_n377_20[0]));
	jspl3 jspl3_w_n377_62(.douta(w_n377_62[0]),.doutb(w_n377_62[1]),.doutc(w_n377_62[2]),.din(w_n377_20[1]));
	jspl jspl_w_n377_63(.douta(w_n377_63[0]),.doutb(w_n377_63[1]),.din(w_n377_20[2]));
	jspl jspl_w_n380_0(.douta(w_n380_0[0]),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.din(n382));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl jspl_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.din(n387));
	jspl3 jspl3_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.doutc(w_n390_0[2]),.din(n390));
	jspl jspl_w_n390_1(.douta(w_n390_1[0]),.doutb(w_n390_1[1]),.din(w_n390_0[0]));
	jspl jspl_w_n392_0(.douta(w_n392_0[0]),.doutb(w_n392_0[1]),.din(n392));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n399_0(.douta(w_n399_0[0]),.doutb(w_n399_0[1]),.din(n399));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl jspl_w_n402_1(.douta(w_n402_1[0]),.doutb(w_n402_1[1]),.din(w_n402_0[0]));
	jspl jspl_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.din(n405));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl jspl_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.din(n410));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(n412));
	jspl3 jspl3_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.doutc(w_n415_0[2]),.din(n415));
	jspl jspl_w_n415_1(.douta(w_n415_1[0]),.doutb(w_n415_1[1]),.din(w_n415_0[0]));
	jspl jspl_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.din(n417));
	jspl jspl_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.din(n419));
	jspl jspl_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.din(n422));
	jspl jspl_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.din(n424));
	jspl3 jspl3_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.doutc(w_n427_0[2]),.din(n427));
	jspl jspl_w_n427_1(.douta(w_n427_1[0]),.doutb(w_n427_1[1]),.din(w_n427_0[0]));
	jspl3 jspl3_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.doutc(w_n430_0[2]),.din(n430));
	jspl jspl_w_n430_1(.douta(w_n430_1[0]),.doutb(w_n430_1[1]),.din(w_n430_0[0]));
	jspl jspl_w_n431_0(.douta(w_n431_0[0]),.doutb(w_n431_0[1]),.din(n431));
	jspl3 jspl3_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.doutc(w_n432_0[2]),.din(n432));
	jspl3 jspl3_w_n432_1(.douta(w_n432_1[0]),.doutb(w_n432_1[1]),.doutc(w_n432_1[2]),.din(w_n432_0[0]));
	jspl3 jspl3_w_n432_2(.douta(w_n432_2[0]),.doutb(w_n432_2[1]),.doutc(w_n432_2[2]),.din(w_n432_0[1]));
	jspl3 jspl3_w_n432_3(.douta(w_n432_3[0]),.doutb(w_n432_3[1]),.doutc(w_n432_3[2]),.din(w_n432_0[2]));
	jspl3 jspl3_w_n432_4(.douta(w_n432_4[0]),.doutb(w_n432_4[1]),.doutc(w_n432_4[2]),.din(w_n432_1[0]));
	jspl3 jspl3_w_n432_5(.douta(w_n432_5[0]),.doutb(w_n432_5[1]),.doutc(w_n432_5[2]),.din(w_n432_1[1]));
	jspl3 jspl3_w_n432_6(.douta(w_n432_6[0]),.doutb(w_n432_6[1]),.doutc(w_n432_6[2]),.din(w_n432_1[2]));
	jspl3 jspl3_w_n432_7(.douta(w_n432_7[0]),.doutb(w_n432_7[1]),.doutc(w_n432_7[2]),.din(w_n432_2[0]));
	jspl3 jspl3_w_n432_8(.douta(w_n432_8[0]),.doutb(w_n432_8[1]),.doutc(w_n432_8[2]),.din(w_n432_2[1]));
	jspl3 jspl3_w_n432_9(.douta(w_n432_9[0]),.doutb(w_n432_9[1]),.doutc(w_n432_9[2]),.din(w_n432_2[2]));
	jspl3 jspl3_w_n432_10(.douta(w_n432_10[0]),.doutb(w_n432_10[1]),.doutc(w_n432_10[2]),.din(w_n432_3[0]));
	jspl3 jspl3_w_n432_11(.douta(w_n432_11[0]),.doutb(w_n432_11[1]),.doutc(w_n432_11[2]),.din(w_n432_3[1]));
	jspl3 jspl3_w_n432_12(.douta(w_n432_12[0]),.doutb(w_n432_12[1]),.doutc(w_n432_12[2]),.din(w_n432_3[2]));
	jspl3 jspl3_w_n432_13(.douta(w_n432_13[0]),.doutb(w_n432_13[1]),.doutc(w_n432_13[2]),.din(w_n432_4[0]));
	jspl3 jspl3_w_n432_14(.douta(w_n432_14[0]),.doutb(w_n432_14[1]),.doutc(w_n432_14[2]),.din(w_n432_4[1]));
	jspl3 jspl3_w_n432_15(.douta(w_n432_15[0]),.doutb(w_n432_15[1]),.doutc(w_n432_15[2]),.din(w_n432_4[2]));
	jspl3 jspl3_w_n432_16(.douta(w_n432_16[0]),.doutb(w_n432_16[1]),.doutc(w_n432_16[2]),.din(w_n432_5[0]));
	jspl3 jspl3_w_n432_17(.douta(w_n432_17[0]),.doutb(w_n432_17[1]),.doutc(w_n432_17[2]),.din(w_n432_5[1]));
	jspl3 jspl3_w_n432_18(.douta(w_n432_18[0]),.doutb(w_n432_18[1]),.doutc(w_n432_18[2]),.din(w_n432_5[2]));
	jspl3 jspl3_w_n432_19(.douta(w_n432_19[0]),.doutb(w_n432_19[1]),.doutc(w_n432_19[2]),.din(w_n432_6[0]));
	jspl3 jspl3_w_n432_20(.douta(w_n432_20[0]),.doutb(w_n432_20[1]),.doutc(w_n432_20[2]),.din(w_n432_6[1]));
	jspl3 jspl3_w_n432_21(.douta(w_n432_21[0]),.doutb(w_n432_21[1]),.doutc(w_n432_21[2]),.din(w_n432_6[2]));
	jspl3 jspl3_w_n432_22(.douta(w_n432_22[0]),.doutb(w_n432_22[1]),.doutc(w_n432_22[2]),.din(w_n432_7[0]));
	jspl3 jspl3_w_n432_23(.douta(w_n432_23[0]),.doutb(w_n432_23[1]),.doutc(w_n432_23[2]),.din(w_n432_7[1]));
	jspl3 jspl3_w_n432_24(.douta(w_n432_24[0]),.doutb(w_n432_24[1]),.doutc(w_n432_24[2]),.din(w_n432_7[2]));
	jspl3 jspl3_w_n432_25(.douta(w_n432_25[0]),.doutb(w_n432_25[1]),.doutc(w_n432_25[2]),.din(w_n432_8[0]));
	jspl3 jspl3_w_n432_26(.douta(w_n432_26[0]),.doutb(w_n432_26[1]),.doutc(w_n432_26[2]),.din(w_n432_8[1]));
	jspl3 jspl3_w_n432_27(.douta(w_n432_27[0]),.doutb(w_n432_27[1]),.doutc(w_n432_27[2]),.din(w_n432_8[2]));
	jspl3 jspl3_w_n432_28(.douta(w_n432_28[0]),.doutb(w_n432_28[1]),.doutc(w_n432_28[2]),.din(w_n432_9[0]));
	jspl3 jspl3_w_n432_29(.douta(w_n432_29[0]),.doutb(w_n432_29[1]),.doutc(w_n432_29[2]),.din(w_n432_9[1]));
	jspl3 jspl3_w_n432_30(.douta(w_n432_30[0]),.doutb(w_n432_30[1]),.doutc(w_n432_30[2]),.din(w_n432_9[2]));
	jspl3 jspl3_w_n432_31(.douta(w_n432_31[0]),.doutb(w_n432_31[1]),.doutc(w_n432_31[2]),.din(w_n432_10[0]));
	jspl3 jspl3_w_n432_32(.douta(w_n432_32[0]),.doutb(w_n432_32[1]),.doutc(w_n432_32[2]),.din(w_n432_10[1]));
	jspl3 jspl3_w_n432_33(.douta(w_n432_33[0]),.doutb(w_n432_33[1]),.doutc(w_n432_33[2]),.din(w_n432_10[2]));
	jspl3 jspl3_w_n432_34(.douta(w_n432_34[0]),.doutb(w_n432_34[1]),.doutc(w_n432_34[2]),.din(w_n432_11[0]));
	jspl3 jspl3_w_n432_35(.douta(w_n432_35[0]),.doutb(w_n432_35[1]),.doutc(w_n432_35[2]),.din(w_n432_11[1]));
	jspl3 jspl3_w_n432_36(.douta(w_n432_36[0]),.doutb(w_n432_36[1]),.doutc(w_n432_36[2]),.din(w_n432_11[2]));
	jspl3 jspl3_w_n432_37(.douta(w_n432_37[0]),.doutb(w_n432_37[1]),.doutc(w_n432_37[2]),.din(w_n432_12[0]));
	jspl3 jspl3_w_n432_38(.douta(w_n432_38[0]),.doutb(w_n432_38[1]),.doutc(w_n432_38[2]),.din(w_n432_12[1]));
	jspl3 jspl3_w_n432_39(.douta(w_n432_39[0]),.doutb(w_n432_39[1]),.doutc(w_n432_39[2]),.din(w_n432_12[2]));
	jspl3 jspl3_w_n432_40(.douta(w_n432_40[0]),.doutb(w_n432_40[1]),.doutc(w_n432_40[2]),.din(w_n432_13[0]));
	jspl3 jspl3_w_n432_41(.douta(w_n432_41[0]),.doutb(w_n432_41[1]),.doutc(w_n432_41[2]),.din(w_n432_13[1]));
	jspl3 jspl3_w_n432_42(.douta(w_n432_42[0]),.doutb(w_n432_42[1]),.doutc(w_n432_42[2]),.din(w_n432_13[2]));
	jspl3 jspl3_w_n432_43(.douta(w_n432_43[0]),.doutb(w_n432_43[1]),.doutc(w_n432_43[2]),.din(w_n432_14[0]));
	jspl3 jspl3_w_n432_44(.douta(w_n432_44[0]),.doutb(w_n432_44[1]),.doutc(w_n432_44[2]),.din(w_n432_14[1]));
	jspl3 jspl3_w_n432_45(.douta(w_n432_45[0]),.doutb(w_n432_45[1]),.doutc(w_n432_45[2]),.din(w_n432_14[2]));
	jspl3 jspl3_w_n432_46(.douta(w_n432_46[0]),.doutb(w_n432_46[1]),.doutc(w_n432_46[2]),.din(w_n432_15[0]));
	jspl3 jspl3_w_n432_47(.douta(w_n432_47[0]),.doutb(w_n432_47[1]),.doutc(w_n432_47[2]),.din(w_n432_15[1]));
	jspl3 jspl3_w_n432_48(.douta(w_n432_48[0]),.doutb(w_n432_48[1]),.doutc(w_n432_48[2]),.din(w_n432_15[2]));
	jspl3 jspl3_w_n432_49(.douta(w_n432_49[0]),.doutb(w_n432_49[1]),.doutc(w_n432_49[2]),.din(w_n432_16[0]));
	jspl3 jspl3_w_n432_50(.douta(w_n432_50[0]),.doutb(w_n432_50[1]),.doutc(w_n432_50[2]),.din(w_n432_16[1]));
	jspl3 jspl3_w_n432_51(.douta(w_n432_51[0]),.doutb(w_n432_51[1]),.doutc(w_n432_51[2]),.din(w_n432_16[2]));
	jspl3 jspl3_w_n432_52(.douta(w_n432_52[0]),.doutb(w_n432_52[1]),.doutc(w_n432_52[2]),.din(w_n432_17[0]));
	jspl3 jspl3_w_n432_53(.douta(w_n432_53[0]),.doutb(w_n432_53[1]),.doutc(w_n432_53[2]),.din(w_n432_17[1]));
	jspl3 jspl3_w_n432_54(.douta(w_n432_54[0]),.doutb(w_n432_54[1]),.doutc(w_n432_54[2]),.din(w_n432_17[2]));
	jspl3 jspl3_w_n432_55(.douta(w_n432_55[0]),.doutb(w_n432_55[1]),.doutc(w_n432_55[2]),.din(w_n432_18[0]));
	jspl3 jspl3_w_n432_56(.douta(w_n432_56[0]),.doutb(w_n432_56[1]),.doutc(w_n432_56[2]),.din(w_n432_18[1]));
	jspl3 jspl3_w_n432_57(.douta(w_n432_57[0]),.doutb(w_n432_57[1]),.doutc(w_n432_57[2]),.din(w_n432_18[2]));
	jspl3 jspl3_w_n432_58(.douta(w_n432_58[0]),.doutb(w_n432_58[1]),.doutc(w_n432_58[2]),.din(w_n432_19[0]));
	jspl3 jspl3_w_n432_59(.douta(w_n432_59[0]),.doutb(w_n432_59[1]),.doutc(w_n432_59[2]),.din(w_n432_19[1]));
	jspl3 jspl3_w_n432_60(.douta(w_n432_60[0]),.doutb(w_n432_60[1]),.doutc(w_n432_60[2]),.din(w_n432_19[2]));
	jspl3 jspl3_w_n432_61(.douta(w_n432_61[0]),.doutb(w_n432_61[1]),.doutc(w_n432_61[2]),.din(w_n432_20[0]));
	jspl3 jspl3_w_n432_62(.douta(w_n432_62[0]),.doutb(w_n432_62[1]),.doutc(w_n432_62[2]),.din(w_n432_20[1]));
	jspl jspl_w_n432_63(.douta(w_n432_63[0]),.doutb(w_n432_63[1]),.din(w_n432_20[2]));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl jspl_w_n436_0(.douta(w_n436_0[0]),.doutb(w_n436_0[1]),.din(n436));
	jspl jspl_w_n439_0(.douta(w_n439_0[0]),.doutb(w_n439_0[1]),.din(n439));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl3 jspl3_w_n444_0(.douta(w_n444_0[0]),.doutb(w_n444_0[1]),.doutc(w_n444_0[2]),.din(n444));
	jspl jspl_w_n444_1(.douta(w_n444_1[0]),.doutb(w_n444_1[1]),.din(w_n444_0[0]));
	jspl jspl_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.din(n446));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.din(n448));
	jspl jspl_w_n451_0(.douta(w_n451_0[0]),.doutb(w_n451_0[1]),.din(n451));
	jspl jspl_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.din(n453));
	jspl3 jspl3_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.doutc(w_n456_0[2]),.din(n456));
	jspl jspl_w_n456_1(.douta(w_n456_1[0]),.doutb(w_n456_1[1]),.din(w_n456_0[0]));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(n459));
	jspl jspl_w_n461_0(.douta(w_n461_0[0]),.doutb(w_n461_0[1]),.din(n461));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(n464));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(n466));
	jspl3 jspl3_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.doutc(w_n469_0[2]),.din(n469));
	jspl jspl_w_n469_1(.douta(w_n469_1[0]),.doutb(w_n469_1[1]),.din(w_n469_0[0]));
	jspl jspl_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.din(n471));
	jspl jspl_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.din(n473));
	jspl jspl_w_n476_0(.douta(w_n476_0[0]),.doutb(w_n476_0[1]),.din(n476));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl3 jspl3_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.doutc(w_n481_0[2]),.din(n481));
	jspl jspl_w_n481_1(.douta(w_n481_1[0]),.doutb(w_n481_1[1]),.din(w_n481_0[0]));
	jspl3 jspl3_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.doutc(w_n484_0[2]),.din(n484));
	jspl jspl_w_n484_1(.douta(w_n484_1[0]),.doutb(w_n484_1[1]),.din(w_n484_0[0]));
	jspl3 jspl3_w_n485_0(.douta(w_n485_0[0]),.doutb(w_n485_0[1]),.doutc(w_n485_0[2]),.din(n485));
	jspl3 jspl3_w_n485_1(.douta(w_n485_1[0]),.doutb(w_n485_1[1]),.doutc(w_n485_1[2]),.din(w_n485_0[0]));
	jspl3 jspl3_w_n485_2(.douta(w_n485_2[0]),.doutb(w_n485_2[1]),.doutc(w_n485_2[2]),.din(w_n485_0[1]));
	jspl3 jspl3_w_n485_3(.douta(w_n485_3[0]),.doutb(w_n485_3[1]),.doutc(w_n485_3[2]),.din(w_n485_0[2]));
	jspl3 jspl3_w_n485_4(.douta(w_n485_4[0]),.doutb(w_n485_4[1]),.doutc(w_n485_4[2]),.din(w_n485_1[0]));
	jspl3 jspl3_w_n485_5(.douta(w_n485_5[0]),.doutb(w_n485_5[1]),.doutc(w_n485_5[2]),.din(w_n485_1[1]));
	jspl3 jspl3_w_n485_6(.douta(w_n485_6[0]),.doutb(w_n485_6[1]),.doutc(w_n485_6[2]),.din(w_n485_1[2]));
	jspl3 jspl3_w_n485_7(.douta(w_n485_7[0]),.doutb(w_n485_7[1]),.doutc(w_n485_7[2]),.din(w_n485_2[0]));
	jspl3 jspl3_w_n485_8(.douta(w_n485_8[0]),.doutb(w_n485_8[1]),.doutc(w_n485_8[2]),.din(w_n485_2[1]));
	jspl3 jspl3_w_n485_9(.douta(w_n485_9[0]),.doutb(w_n485_9[1]),.doutc(w_n485_9[2]),.din(w_n485_2[2]));
	jspl3 jspl3_w_n485_10(.douta(w_n485_10[0]),.doutb(w_n485_10[1]),.doutc(w_n485_10[2]),.din(w_n485_3[0]));
	jspl3 jspl3_w_n485_11(.douta(w_n485_11[0]),.doutb(w_n485_11[1]),.doutc(w_n485_11[2]),.din(w_n485_3[1]));
	jspl3 jspl3_w_n485_12(.douta(w_n485_12[0]),.doutb(w_n485_12[1]),.doutc(w_n485_12[2]),.din(w_n485_3[2]));
	jspl3 jspl3_w_n485_13(.douta(w_n485_13[0]),.doutb(w_n485_13[1]),.doutc(w_n485_13[2]),.din(w_n485_4[0]));
	jspl3 jspl3_w_n485_14(.douta(w_n485_14[0]),.doutb(w_n485_14[1]),.doutc(w_n485_14[2]),.din(w_n485_4[1]));
	jspl3 jspl3_w_n485_15(.douta(w_n485_15[0]),.doutb(w_n485_15[1]),.doutc(w_n485_15[2]),.din(w_n485_4[2]));
	jspl3 jspl3_w_n485_16(.douta(w_n485_16[0]),.doutb(w_n485_16[1]),.doutc(w_n485_16[2]),.din(w_n485_5[0]));
	jspl3 jspl3_w_n485_17(.douta(w_n485_17[0]),.doutb(w_n485_17[1]),.doutc(w_n485_17[2]),.din(w_n485_5[1]));
	jspl3 jspl3_w_n485_18(.douta(w_n485_18[0]),.doutb(w_n485_18[1]),.doutc(w_n485_18[2]),.din(w_n485_5[2]));
	jspl3 jspl3_w_n485_19(.douta(w_n485_19[0]),.doutb(w_n485_19[1]),.doutc(w_n485_19[2]),.din(w_n485_6[0]));
	jspl3 jspl3_w_n485_20(.douta(w_n485_20[0]),.doutb(w_n485_20[1]),.doutc(w_n485_20[2]),.din(w_n485_6[1]));
	jspl3 jspl3_w_n485_21(.douta(w_n485_21[0]),.doutb(w_n485_21[1]),.doutc(w_n485_21[2]),.din(w_n485_6[2]));
	jspl3 jspl3_w_n485_22(.douta(w_n485_22[0]),.doutb(w_n485_22[1]),.doutc(w_n485_22[2]),.din(w_n485_7[0]));
	jspl3 jspl3_w_n485_23(.douta(w_n485_23[0]),.doutb(w_n485_23[1]),.doutc(w_n485_23[2]),.din(w_n485_7[1]));
	jspl3 jspl3_w_n485_24(.douta(w_n485_24[0]),.doutb(w_n485_24[1]),.doutc(w_n485_24[2]),.din(w_n485_7[2]));
	jspl3 jspl3_w_n485_25(.douta(w_n485_25[0]),.doutb(w_n485_25[1]),.doutc(w_n485_25[2]),.din(w_n485_8[0]));
	jspl3 jspl3_w_n485_26(.douta(w_n485_26[0]),.doutb(w_n485_26[1]),.doutc(w_n485_26[2]),.din(w_n485_8[1]));
	jspl3 jspl3_w_n485_27(.douta(w_n485_27[0]),.doutb(w_n485_27[1]),.doutc(w_n485_27[2]),.din(w_n485_8[2]));
	jspl3 jspl3_w_n485_28(.douta(w_n485_28[0]),.doutb(w_n485_28[1]),.doutc(w_n485_28[2]),.din(w_n485_9[0]));
	jspl3 jspl3_w_n485_29(.douta(w_n485_29[0]),.doutb(w_n485_29[1]),.doutc(w_n485_29[2]),.din(w_n485_9[1]));
	jspl3 jspl3_w_n485_30(.douta(w_n485_30[0]),.doutb(w_n485_30[1]),.doutc(w_n485_30[2]),.din(w_n485_9[2]));
	jspl3 jspl3_w_n485_31(.douta(w_n485_31[0]),.doutb(w_n485_31[1]),.doutc(w_n485_31[2]),.din(w_n485_10[0]));
	jspl3 jspl3_w_n485_32(.douta(w_n485_32[0]),.doutb(w_n485_32[1]),.doutc(w_n485_32[2]),.din(w_n485_10[1]));
	jspl3 jspl3_w_n485_33(.douta(w_n485_33[0]),.doutb(w_n485_33[1]),.doutc(w_n485_33[2]),.din(w_n485_10[2]));
	jspl3 jspl3_w_n485_34(.douta(w_n485_34[0]),.doutb(w_n485_34[1]),.doutc(w_n485_34[2]),.din(w_n485_11[0]));
	jspl3 jspl3_w_n485_35(.douta(w_n485_35[0]),.doutb(w_n485_35[1]),.doutc(w_n485_35[2]),.din(w_n485_11[1]));
	jspl3 jspl3_w_n485_36(.douta(w_n485_36[0]),.doutb(w_n485_36[1]),.doutc(w_n485_36[2]),.din(w_n485_11[2]));
	jspl3 jspl3_w_n485_37(.douta(w_n485_37[0]),.doutb(w_n485_37[1]),.doutc(w_n485_37[2]),.din(w_n485_12[0]));
	jspl3 jspl3_w_n485_38(.douta(w_n485_38[0]),.doutb(w_n485_38[1]),.doutc(w_n485_38[2]),.din(w_n485_12[1]));
	jspl3 jspl3_w_n485_39(.douta(w_n485_39[0]),.doutb(w_n485_39[1]),.doutc(w_n485_39[2]),.din(w_n485_12[2]));
	jspl3 jspl3_w_n485_40(.douta(w_n485_40[0]),.doutb(w_n485_40[1]),.doutc(w_n485_40[2]),.din(w_n485_13[0]));
	jspl3 jspl3_w_n485_41(.douta(w_n485_41[0]),.doutb(w_n485_41[1]),.doutc(w_n485_41[2]),.din(w_n485_13[1]));
	jspl3 jspl3_w_n485_42(.douta(w_n485_42[0]),.doutb(w_n485_42[1]),.doutc(w_n485_42[2]),.din(w_n485_13[2]));
	jspl3 jspl3_w_n485_43(.douta(w_n485_43[0]),.doutb(w_n485_43[1]),.doutc(w_n485_43[2]),.din(w_n485_14[0]));
	jspl3 jspl3_w_n485_44(.douta(w_n485_44[0]),.doutb(w_n485_44[1]),.doutc(w_n485_44[2]),.din(w_n485_14[1]));
	jspl3 jspl3_w_n485_45(.douta(w_n485_45[0]),.doutb(w_n485_45[1]),.doutc(w_n485_45[2]),.din(w_n485_14[2]));
	jspl3 jspl3_w_n485_46(.douta(w_n485_46[0]),.doutb(w_n485_46[1]),.doutc(w_n485_46[2]),.din(w_n485_15[0]));
	jspl3 jspl3_w_n485_47(.douta(w_n485_47[0]),.doutb(w_n485_47[1]),.doutc(w_n485_47[2]),.din(w_n485_15[1]));
	jspl3 jspl3_w_n485_48(.douta(w_n485_48[0]),.doutb(w_n485_48[1]),.doutc(w_n485_48[2]),.din(w_n485_15[2]));
	jspl3 jspl3_w_n485_49(.douta(w_n485_49[0]),.doutb(w_n485_49[1]),.doutc(w_n485_49[2]),.din(w_n485_16[0]));
	jspl3 jspl3_w_n485_50(.douta(w_n485_50[0]),.doutb(w_n485_50[1]),.doutc(w_n485_50[2]),.din(w_n485_16[1]));
	jspl3 jspl3_w_n485_51(.douta(w_n485_51[0]),.doutb(w_n485_51[1]),.doutc(w_n485_51[2]),.din(w_n485_16[2]));
	jspl3 jspl3_w_n485_52(.douta(w_n485_52[0]),.doutb(w_n485_52[1]),.doutc(w_n485_52[2]),.din(w_n485_17[0]));
	jspl3 jspl3_w_n485_53(.douta(w_n485_53[0]),.doutb(w_n485_53[1]),.doutc(w_n485_53[2]),.din(w_n485_17[1]));
	jspl3 jspl3_w_n485_54(.douta(w_n485_54[0]),.doutb(w_n485_54[1]),.doutc(w_n485_54[2]),.din(w_n485_17[2]));
	jspl3 jspl3_w_n485_55(.douta(w_n485_55[0]),.doutb(w_n485_55[1]),.doutc(w_n485_55[2]),.din(w_n485_18[0]));
	jspl3 jspl3_w_n485_56(.douta(w_n485_56[0]),.doutb(w_n485_56[1]),.doutc(w_n485_56[2]),.din(w_n485_18[1]));
	jspl3 jspl3_w_n485_57(.douta(w_n485_57[0]),.doutb(w_n485_57[1]),.doutc(w_n485_57[2]),.din(w_n485_18[2]));
	jspl3 jspl3_w_n485_58(.douta(w_n485_58[0]),.doutb(w_n485_58[1]),.doutc(w_n485_58[2]),.din(w_n485_19[0]));
	jspl3 jspl3_w_n485_59(.douta(w_n485_59[0]),.doutb(w_n485_59[1]),.doutc(w_n485_59[2]),.din(w_n485_19[1]));
	jspl3 jspl3_w_n485_60(.douta(w_n485_60[0]),.doutb(w_n485_60[1]),.doutc(w_n485_60[2]),.din(w_n485_19[2]));
	jspl3 jspl3_w_n485_61(.douta(w_n485_61[0]),.doutb(w_n485_61[1]),.doutc(w_n485_61[2]),.din(w_n485_20[0]));
	jspl3 jspl3_w_n485_62(.douta(w_n485_62[0]),.doutb(w_n485_62[1]),.doutc(w_n485_62[2]),.din(w_n485_20[1]));
	jspl jspl_w_n485_63(.douta(w_n485_63[0]),.doutb(w_n485_63[1]),.din(w_n485_20[2]));
	jspl jspl_w_n488_0(.douta(w_n488_0[0]),.doutb(w_n488_0[1]),.din(n488));
	jspl jspl_w_n490_0(.douta(w_n490_0[0]),.doutb(w_n490_0[1]),.din(n490));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.din(n495));
	jspl jspl_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.din(n497));
	jspl3 jspl3_w_n500_0(.douta(w_n500_0[0]),.doutb(w_n500_0[1]),.doutc(w_n500_0[2]),.din(n500));
	jspl jspl_w_n500_1(.douta(w_n500_1[0]),.doutb(w_n500_1[1]),.din(w_n500_0[0]));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(n509));
	jspl3 jspl3_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.doutc(w_n512_0[2]),.din(n512));
	jspl jspl_w_n512_1(.douta(w_n512_1[0]),.doutb(w_n512_1[1]),.din(w_n512_0[0]));
	jspl jspl_w_n515_0(.douta(w_n515_0[0]),.doutb(w_n515_0[1]),.din(n515));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n525_0(.douta(w_n525_0[0]),.doutb(w_n525_0[1]),.doutc(w_n525_0[2]),.din(n525));
	jspl jspl_w_n525_1(.douta(w_n525_1[0]),.doutb(w_n525_1[1]),.din(w_n525_0[0]));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_n529_0[0]),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(n532));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl3 jspl3_w_n537_0(.douta(w_n537_0[0]),.doutb(w_n537_0[1]),.doutc(w_n537_0[2]),.din(n537));
	jspl jspl_w_n537_1(.douta(w_n537_1[0]),.doutb(w_n537_1[1]),.din(w_n537_0[0]));
	jspl3 jspl3_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.doutc(w_n540_0[2]),.din(n540));
	jspl jspl_w_n540_1(.douta(w_n540_1[0]),.doutb(w_n540_1[1]),.din(w_n540_0[0]));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(n547));
	jspl jspl_w_n549_0(.douta(w_n549_0[0]),.doutb(w_n549_0[1]),.din(n549));
	jspl3 jspl3_w_n552_0(.douta(w_n552_0[0]),.doutb(w_n552_0[1]),.doutc(w_n552_0[2]),.din(n552));
	jspl jspl_w_n552_1(.douta(w_n552_1[0]),.doutb(w_n552_1[1]),.din(w_n552_0[0]));
	jspl jspl_w_n554_0(.douta(w_n554_0[0]),.doutb(w_n554_0[1]),.din(n554));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n558_0(.douta(w_n558_0[0]),.doutb(w_n558_0[1]),.din(n558));
	jspl jspl_w_n559_0(.douta(w_n559_0[0]),.doutb(w_n559_0[1]),.din(n559));
	jspl3 jspl3_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.doutc(w_n562_0[2]),.din(n562));
	jspl jspl_w_n562_1(.douta(w_n562_1[0]),.doutb(w_n562_1[1]),.din(w_n562_0[0]));
	jspl jspl_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.din(n565));
	jspl jspl_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.din(n567));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl jspl_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.din(n572));
	jspl3 jspl3_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.doutc(w_n575_0[2]),.din(n575));
	jspl jspl_w_n575_1(.douta(w_n575_1[0]),.doutb(w_n575_1[1]),.din(w_n575_0[0]));
	jspl jspl_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.din(n577));
	jspl jspl_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.din(n579));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl jspl_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.din(n584));
	jspl3 jspl3_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.doutc(w_n587_0[2]),.din(n587));
	jspl jspl_w_n587_1(.douta(w_n587_1[0]),.doutb(w_n587_1[1]),.din(w_n587_0[0]));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.doutc(w_n590_0[2]),.din(n590));
	jspl jspl_w_n590_1(.douta(w_n590_1[0]),.doutb(w_n590_1[1]),.din(w_n590_0[0]));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(n593));
	jspl jspl_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.din(n595));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(n598));
	jspl jspl_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.din(n600));
	jspl3 jspl3_w_n603_0(.douta(w_n603_0[0]),.doutb(w_n603_0[1]),.doutc(w_n603_0[2]),.din(n603));
	jspl jspl_w_n603_1(.douta(w_n603_1[0]),.doutb(w_n603_1[1]),.din(w_n603_0[0]));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl jspl_w_n610_0(.douta(w_n610_0[0]),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl3 jspl3_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.doutc(w_n615_0[2]),.din(n615));
	jspl jspl_w_n615_1(.douta(w_n615_1[0]),.doutb(w_n615_1[1]),.din(w_n615_0[0]));
	jspl jspl_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.din(n618));
	jspl jspl_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.din(n620));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.din(n625));
	jspl3 jspl3_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.doutc(w_n628_0[2]),.din(n628));
	jspl jspl_w_n628_1(.douta(w_n628_1[0]),.doutb(w_n628_1[1]),.din(w_n628_0[0]));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(n632));
	jspl jspl_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.din(n635));
	jspl jspl_w_n637_0(.douta(w_n637_0[0]),.doutb(w_n637_0[1]),.din(n637));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_n640_0[2]),.din(n640));
	jspl jspl_w_n640_1(.douta(w_n640_1[0]),.doutb(w_n640_1[1]),.din(w_n640_0[0]));
	jspl3 jspl3_w_n643_0(.douta(w_n643_0[0]),.doutb(w_n643_0[1]),.doutc(w_n643_0[2]),.din(n643));
	jspl jspl_w_n643_1(.douta(w_n643_1[0]),.doutb(w_n643_1[1]),.din(w_n643_0[0]));
	jspl jspl_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(n647));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl3 jspl3_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.doutc(w_n655_0[2]),.din(n655));
	jspl jspl_w_n655_1(.douta(w_n655_1[0]),.doutb(w_n655_1[1]),.din(w_n655_0[0]));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(n662));
	jspl jspl_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.din(n664));
	jspl3 jspl3_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.doutc(w_n667_0[2]),.din(n667));
	jspl jspl_w_n667_1(.douta(w_n667_1[0]),.doutb(w_n667_1[1]),.din(w_n667_0[0]));
	jspl jspl_w_n670_0(.douta(w_n670_0[0]),.doutb(w_n670_0[1]),.din(n670));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.din(n675));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl3 jspl3_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.doutc(w_n680_0[2]),.din(n680));
	jspl jspl_w_n680_1(.douta(w_n680_1[0]),.doutb(w_n680_1[1]),.din(w_n680_0[0]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(n684));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl3 jspl3_w_n692_0(.douta(w_n692_0[0]),.doutb(w_n692_0[1]),.doutc(w_n692_0[2]),.din(n692));
	jspl jspl_w_n692_1(.douta(w_n692_1[0]),.doutb(w_n692_1[1]),.din(w_n692_0[0]));
	jspl3 jspl3_w_n695_0(.douta(w_n695_0[0]),.doutb(w_n695_0[1]),.doutc(w_n695_0[2]),.din(n695));
	jspl jspl_w_n695_1(.douta(w_n695_1[0]),.doutb(w_n695_1[1]),.din(w_n695_0[0]));
	jspl jspl_w_n698_0(.douta(w_n698_0[0]),.doutb(w_n698_0[1]),.din(n698));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.din(n703));
	jspl jspl_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.din(n707));
	jspl3 jspl3_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.doutc(w_n709_0[2]),.din(n709));
	jspl jspl_w_n709_1(.douta(w_n709_1[0]),.doutb(w_n709_1[1]),.din(w_n709_0[0]));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl3 jspl3_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.doutc(w_n719_0[2]),.din(n719));
	jspl jspl_w_n719_1(.douta(w_n719_1[0]),.doutb(w_n719_1[1]),.din(w_n719_0[0]));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(n724));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n730_0(.douta(w_n730_0[0]),.doutb(w_n730_0[1]),.doutc(w_n730_0[2]),.din(n730));
	jspl jspl_w_n730_1(.douta(w_n730_1[0]),.doutb(w_n730_1[1]),.din(w_n730_0[0]));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(n734));
	jspl jspl_w_n738_0(.douta(w_n738_0[0]),.doutb(w_n738_0[1]),.din(n738));
	jspl3 jspl3_w_n740_0(.douta(w_n740_0[0]),.doutb(w_n740_0[1]),.doutc(w_n740_0[2]),.din(n740));
	jspl jspl_w_n740_1(.douta(w_n740_1[0]),.doutb(w_n740_1[1]),.din(w_n740_0[0]));
	jspl3 jspl3_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.doutc(w_n743_0[2]),.din(n743));
	jspl jspl_w_n743_1(.douta(w_n743_1[0]),.doutb(w_n743_1[1]),.din(w_n743_0[0]));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(n747));
	jspl jspl_w_n751_0(.douta(w_n751_0[0]),.doutb(w_n751_0[1]),.din(n751));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.doutc(w_n753_0[2]),.din(n753));
	jspl jspl_w_n753_1(.douta(w_n753_1[0]),.doutb(w_n753_1[1]),.din(w_n753_0[0]));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.din(n761));
	jspl3 jspl3_w_n763_0(.douta(w_n763_0[0]),.doutb(w_n763_0[1]),.doutc(w_n763_0[2]),.din(n763));
	jspl jspl_w_n763_1(.douta(w_n763_1[0]),.doutb(w_n763_1[1]),.din(w_n763_0[0]));
	jspl jspl_w_n768_0(.douta(w_n768_0[0]),.doutb(w_n768_0[1]),.din(n768));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(n772));
	jspl3 jspl3_w_n774_0(.douta(w_n774_0[0]),.doutb(w_n774_0[1]),.doutc(w_n774_0[2]),.din(n774));
	jspl jspl_w_n774_1(.douta(w_n774_1[0]),.doutb(w_n774_1[1]),.din(w_n774_0[0]));
	jspl jspl_w_n778_0(.douta(w_n778_0[0]),.doutb(w_n778_0[1]),.din(n778));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(n782));
	jspl3 jspl3_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.doutc(w_n784_0[2]),.din(n784));
	jspl jspl_w_n784_1(.douta(w_n784_1[0]),.doutb(w_n784_1[1]),.din(w_n784_0[0]));
	jspl3 jspl3_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.doutc(w_n787_0[2]),.din(n787));
	jspl jspl_w_n787_1(.douta(w_n787_1[0]),.doutb(w_n787_1[1]),.din(w_n787_0[0]));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl3 jspl3_w_n798_0(.douta(w_n798_0[0]),.doutb(w_n798_0[1]),.doutc(w_n798_0[2]),.din(n798));
	jspl jspl_w_n798_1(.douta(w_n798_1[0]),.doutb(w_n798_1[1]),.din(w_n798_0[0]));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.din(n806));
	jspl3 jspl3_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.doutc(w_n808_0[2]),.din(n808));
	jspl jspl_w_n808_1(.douta(w_n808_1[0]),.doutb(w_n808_1[1]),.din(w_n808_0[0]));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(n817));
	jspl3 jspl3_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.doutc(w_n819_0[2]),.din(n819));
	jspl jspl_w_n819_1(.douta(w_n819_1[0]),.doutb(w_n819_1[1]),.din(w_n819_0[0]));
	jspl jspl_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl3 jspl3_w_n829_0(.douta(w_n829_0[0]),.doutb(w_n829_0[1]),.doutc(w_n829_0[2]),.din(n829));
	jspl jspl_w_n829_1(.douta(w_n829_1[0]),.doutb(w_n829_1[1]),.din(w_n829_0[0]));
	jspl3 jspl3_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.doutc(w_n832_0[2]),.din(n832));
	jspl jspl_w_n832_1(.douta(w_n832_1[0]),.doutb(w_n832_1[1]),.din(w_n832_0[0]));
	jspl jspl_w_n836_0(.douta(w_n836_0[0]),.doutb(w_n836_0[1]),.din(n836));
	jspl jspl_w_n840_0(.douta(w_n840_0[0]),.doutb(w_n840_0[1]),.din(n840));
	jspl3 jspl3_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.doutc(w_n842_0[2]),.din(n842));
	jspl jspl_w_n842_1(.douta(w_n842_1[0]),.doutb(w_n842_1[1]),.din(w_n842_0[0]));
	jspl jspl_w_n846_0(.douta(w_n846_0[0]),.doutb(w_n846_0[1]),.din(n846));
	jspl jspl_w_n850_0(.douta(w_n850_0[0]),.doutb(w_n850_0[1]),.din(n850));
	jspl3 jspl3_w_n852_0(.douta(w_n852_0[0]),.doutb(w_n852_0[1]),.doutc(w_n852_0[2]),.din(n852));
	jspl jspl_w_n852_1(.douta(w_n852_1[0]),.doutb(w_n852_1[1]),.din(w_n852_0[0]));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(n857));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(n861));
	jspl3 jspl3_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.doutc(w_n863_0[2]),.din(n863));
	jspl jspl_w_n863_1(.douta(w_n863_1[0]),.doutb(w_n863_1[1]),.din(w_n863_0[0]));
	jspl jspl_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.din(n867));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl3 jspl3_w_n873_0(.douta(w_n873_0[0]),.doutb(w_n873_0[1]),.doutc(w_n873_0[2]),.din(n873));
	jspl jspl_w_n873_1(.douta(w_n873_1[0]),.doutb(w_n873_1[1]),.din(w_n873_0[0]));
	jspl3 jspl3_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.doutc(w_n876_0[2]),.din(n876));
	jspl jspl_w_n876_1(.douta(w_n876_1[0]),.doutb(w_n876_1[1]),.din(w_n876_0[0]));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n883_0(.douta(w_n883_0[0]),.doutb(w_n883_0[1]),.din(n883));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_n887_0[1]),.din(n887));
	jspl3 jspl3_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.doutc(w_n889_0[2]),.din(n889));
	jspl jspl_w_n889_1(.douta(w_n889_1[0]),.doutb(w_n889_1[1]),.din(w_n889_0[0]));
	jspl jspl_w_n893_0(.douta(w_n893_0[0]),.doutb(w_n893_0[1]),.din(n893));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl3 jspl3_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.doutc(w_n899_0[2]),.din(n899));
	jspl jspl_w_n899_1(.douta(w_n899_1[0]),.doutb(w_n899_1[1]),.din(w_n899_0[0]));
	jspl jspl_w_n904_0(.douta(w_n904_0[0]),.doutb(w_n904_0[1]),.din(n904));
	jspl jspl_w_n908_0(.douta(w_n908_0[0]),.doutb(w_n908_0[1]),.din(n908));
	jspl3 jspl3_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.doutc(w_n910_0[2]),.din(n910));
	jspl jspl_w_n910_1(.douta(w_n910_1[0]),.doutb(w_n910_1[1]),.din(w_n910_0[0]));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.din(n918));
	jspl3 jspl3_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.doutc(w_n920_0[2]),.din(n920));
	jspl jspl_w_n920_1(.douta(w_n920_1[0]),.doutb(w_n920_1[1]),.din(w_n920_0[0]));
	jspl3 jspl3_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.doutc(w_n923_0[2]),.din(n923));
	jspl jspl_w_n923_1(.douta(w_n923_1[0]),.doutb(w_n923_1[1]),.din(w_n923_0[0]));
	jspl jspl_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.din(n927));
	jspl jspl_w_n931_0(.douta(w_n931_0[0]),.doutb(w_n931_0[1]),.din(n931));
	jspl3 jspl3_w_n933_0(.douta(w_n933_0[0]),.doutb(w_n933_0[1]),.doutc(w_n933_0[2]),.din(n933));
	jspl jspl_w_n933_1(.douta(w_n933_1[0]),.doutb(w_n933_1[1]),.din(w_n933_0[0]));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n941_0(.douta(w_n941_0[0]),.doutb(w_n941_0[1]),.din(n941));
	jspl3 jspl3_w_n943_0(.douta(w_n943_0[0]),.doutb(w_n943_0[1]),.doutc(w_n943_0[2]),.din(n943));
	jspl jspl_w_n943_1(.douta(w_n943_1[0]),.doutb(w_n943_1[1]),.din(w_n943_0[0]));
	jspl jspl_w_n948_0(.douta(w_n948_0[0]),.doutb(w_n948_0[1]),.din(n948));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl3 jspl3_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.doutc(w_n954_0[2]),.din(n954));
	jspl jspl_w_n954_1(.douta(w_n954_1[0]),.doutb(w_n954_1[1]),.din(w_n954_0[0]));
	jspl jspl_w_n958_0(.douta(w_n958_0[0]),.doutb(w_n958_0[1]),.din(n958));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl3 jspl3_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.doutc(w_n964_0[2]),.din(n964));
	jspl jspl_w_n964_1(.douta(w_n964_1[0]),.doutb(w_n964_1[1]),.din(w_n964_0[0]));
	jspl3 jspl3_w_n967_0(.douta(w_n967_0[0]),.doutb(w_n967_0[1]),.doutc(w_n967_0[2]),.din(n967));
	jspl jspl_w_n967_1(.douta(w_n967_1[0]),.doutb(w_n967_1[1]),.din(w_n967_0[0]));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n976_0(.douta(w_n976_0[0]),.doutb(w_n976_0[1]),.din(n976));
	jspl3 jspl3_w_n978_0(.douta(w_n978_0[0]),.doutb(w_n978_0[1]),.doutc(w_n978_0[2]),.din(n978));
	jspl jspl_w_n978_1(.douta(w_n978_1[0]),.doutb(w_n978_1[1]),.din(w_n978_0[0]));
	jspl jspl_w_n982_0(.douta(w_n982_0[0]),.doutb(w_n982_0[1]),.din(n982));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(n986));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.doutc(w_n988_0[2]),.din(n988));
	jspl jspl_w_n988_1(.douta(w_n988_1[0]),.doutb(w_n988_1[1]),.din(w_n988_0[0]));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_n993_0[1]),.din(n993));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.doutc(w_n999_0[2]),.din(n999));
	jspl jspl_w_n999_1(.douta(w_n999_1[0]),.doutb(w_n999_1[1]),.din(w_n999_0[0]));
	jspl jspl_w_n1003_0(.douta(w_n1003_0[0]),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl3 jspl3_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.doutc(w_n1009_0[2]),.din(n1009));
	jspl jspl_w_n1009_1(.douta(w_n1009_1[0]),.doutb(w_n1009_1[1]),.din(w_n1009_0[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl jspl_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.din(w_n1012_0[0]));
	jspl jspl_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.din(n1016));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(n1018));
	jspl jspl_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.din(n1019));
	jspl3 jspl3_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.doutc(w_n1022_0[2]),.din(n1022));
	jspl jspl_w_n1022_1(.douta(w_n1022_1[0]),.doutb(w_n1022_1[1]),.din(w_n1022_0[0]));
	jspl jspl_w_n1024_0(.douta(w_n1024_0[0]),.doutb(w_n1024_0[1]),.din(n1024));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.din(n1029));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl3 jspl3_w_n1034_0(.douta(w_n1034_0[0]),.doutb(w_n1034_0[1]),.doutc(w_n1034_0[2]),.din(n1034));
	jspl jspl_w_n1034_1(.douta(w_n1034_1[0]),.doutb(w_n1034_1[1]),.din(w_n1034_0[0]));
	jspl jspl_w_n1037_0(.douta(w_n1037_0[0]),.doutb(w_n1037_0[1]),.din(n1037));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.din(n1039));
	jspl jspl_w_n1042_0(.douta(w_n1042_0[0]),.doutb(w_n1042_0[1]),.din(n1042));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(n1044));
	jspl3 jspl3_w_n1047_0(.douta(w_n1047_0[0]),.doutb(w_n1047_0[1]),.doutc(w_n1047_0[2]),.din(n1047));
	jspl jspl_w_n1047_1(.douta(w_n1047_1[0]),.doutb(w_n1047_1[1]),.din(w_n1047_0[0]));
	jspl jspl_w_n1051_0(.douta(w_n1051_0[0]),.doutb(w_n1051_0[1]),.din(n1051));
	jspl jspl_w_n1055_0(.douta(w_n1055_0[0]),.doutb(w_n1055_0[1]),.din(n1055));
	jspl3 jspl3_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.doutc(w_n1057_0[2]),.din(n1057));
	jspl jspl_w_n1057_1(.douta(w_n1057_1[0]),.doutb(w_n1057_1[1]),.din(w_n1057_0[0]));
	jspl3 jspl3_w_n1060_0(.douta(w_n1060_0[0]),.doutb(w_n1060_0[1]),.doutc(w_n1060_0[2]),.din(n1060));
	jspl jspl_w_n1060_1(.douta(w_n1060_1[0]),.doutb(w_n1060_1[1]),.din(w_n1060_0[0]));
	jspl jspl_w_n1063_0(.douta(w_n1063_0[0]),.doutb(w_n1063_0[1]),.din(n1063));
	jspl3 jspl3_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.doutc(w_n1072_0[2]),.din(n1072));
	jspl jspl_w_n1072_1(.douta(w_n1072_1[0]),.doutb(w_n1072_1[1]),.din(w_n1072_0[0]));
	jspl3 jspl3_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.doutc(w_n1080_0[2]),.din(n1080));
	jspl jspl_w_n1080_1(.douta(w_n1080_1[0]),.doutb(w_n1080_1[1]),.din(w_n1080_0[0]));
	jspl3 jspl3_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.doutc(w_n1089_0[2]),.din(n1089));
	jspl jspl_w_n1089_1(.douta(w_n1089_1[0]),.doutb(w_n1089_1[1]),.din(w_n1089_0[0]));
	jspl3 jspl3_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.doutc(w_n1097_0[2]),.din(n1097));
	jspl jspl_w_n1097_1(.douta(w_n1097_1[0]),.doutb(w_n1097_1[1]),.din(w_n1097_0[0]));
	jspl3 jspl3_w_n1100_0(.douta(w_n1100_0[0]),.doutb(w_n1100_0[1]),.doutc(w_n1100_0[2]),.din(n1100));
	jspl jspl_w_n1100_1(.douta(w_n1100_1[0]),.doutb(w_n1100_1[1]),.din(w_n1100_0[0]));
	jspl3 jspl3_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_n1108_0[1]),.doutc(w_n1108_0[2]),.din(n1108));
	jspl jspl_w_n1108_1(.douta(w_n1108_1[0]),.doutb(w_n1108_1[1]),.din(w_n1108_0[0]));
	jspl3 jspl3_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.doutc(w_n1116_0[2]),.din(n1116));
	jspl jspl_w_n1116_1(.douta(w_n1116_1[0]),.doutb(w_n1116_1[1]),.din(w_n1116_0[0]));
	jspl3 jspl3_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.doutc(w_n1125_0[2]),.din(n1125));
	jspl jspl_w_n1125_1(.douta(w_n1125_1[0]),.doutb(w_n1125_1[1]),.din(w_n1125_0[0]));
	jspl3 jspl3_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.doutc(w_n1133_0[2]),.din(n1133));
	jspl jspl_w_n1133_1(.douta(w_n1133_1[0]),.doutb(w_n1133_1[1]),.din(w_n1133_0[0]));
	jspl3 jspl3_w_n1136_0(.douta(w_n1136_0[0]),.doutb(w_n1136_0[1]),.doutc(w_n1136_0[2]),.din(n1136));
	jspl jspl_w_n1136_1(.douta(w_n1136_1[0]),.doutb(w_n1136_1[1]),.din(w_n1136_0[0]));
	jspl3 jspl3_w_n1145_0(.douta(w_n1145_0[0]),.doutb(w_n1145_0[1]),.doutc(w_n1145_0[2]),.din(n1145));
	jspl jspl_w_n1145_1(.douta(w_n1145_1[0]),.doutb(w_n1145_1[1]),.din(w_n1145_0[0]));
	jspl3 jspl3_w_n1153_0(.douta(w_n1153_0[0]),.doutb(w_n1153_0[1]),.doutc(w_n1153_0[2]),.din(n1153));
	jspl jspl_w_n1153_1(.douta(w_n1153_1[0]),.doutb(w_n1153_1[1]),.din(w_n1153_0[0]));
	jspl3 jspl3_w_n1162_0(.douta(w_n1162_0[0]),.doutb(w_n1162_0[1]),.doutc(w_n1162_0[2]),.din(n1162));
	jspl jspl_w_n1162_1(.douta(w_n1162_1[0]),.doutb(w_n1162_1[1]),.din(w_n1162_0[0]));
	jspl3 jspl3_w_n1170_0(.douta(w_n1170_0[0]),.doutb(w_n1170_0[1]),.doutc(w_n1170_0[2]),.din(n1170));
	jspl jspl_w_n1170_1(.douta(w_n1170_1[0]),.doutb(w_n1170_1[1]),.din(w_n1170_0[0]));
	jspl3 jspl3_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.doutc(w_n1173_0[2]),.din(n1173));
	jspl jspl_w_n1173_1(.douta(w_n1173_1[0]),.doutb(w_n1173_1[1]),.din(w_n1173_0[0]));
	jspl3 jspl3_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.doutc(w_n1181_0[2]),.din(n1181));
	jspl jspl_w_n1181_1(.douta(w_n1181_1[0]),.doutb(w_n1181_1[1]),.din(w_n1181_0[0]));
	jspl3 jspl3_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.doutc(w_n1189_0[2]),.din(n1189));
	jspl jspl_w_n1189_1(.douta(w_n1189_1[0]),.doutb(w_n1189_1[1]),.din(w_n1189_0[0]));
	jspl3 jspl3_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.doutc(w_n1198_0[2]),.din(n1198));
	jspl jspl_w_n1198_1(.douta(w_n1198_1[0]),.doutb(w_n1198_1[1]),.din(w_n1198_0[0]));
	jspl3 jspl3_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.doutc(w_n1206_0[2]),.din(n1206));
	jspl jspl_w_n1206_1(.douta(w_n1206_1[0]),.doutb(w_n1206_1[1]),.din(w_n1206_0[0]));
	jspl3 jspl3_w_n1209_0(.douta(w_n1209_0[0]),.doutb(w_n1209_0[1]),.doutc(w_n1209_0[2]),.din(n1209));
	jspl jspl_w_n1209_1(.douta(w_n1209_1[0]),.doutb(w_n1209_1[1]),.din(w_n1209_0[0]));
	jspl jspl_w_n1212_0(.douta(w_n1212_0[0]),.doutb(w_n1212_0[1]),.din(n1212));
	jspl3 jspl3_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.doutc(w_n1220_0[2]),.din(n1220));
	jspl jspl_w_n1220_1(.douta(w_n1220_1[0]),.doutb(w_n1220_1[1]),.din(w_n1220_0[0]));
	jspl3 jspl3_w_n1228_0(.douta(w_n1228_0[0]),.doutb(w_n1228_0[1]),.doutc(w_n1228_0[2]),.din(n1228));
	jspl jspl_w_n1228_1(.douta(w_n1228_1[0]),.doutb(w_n1228_1[1]),.din(w_n1228_0[0]));
	jspl3 jspl3_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.doutc(w_n1237_0[2]),.din(n1237));
	jspl jspl_w_n1237_1(.douta(w_n1237_1[0]),.doutb(w_n1237_1[1]),.din(w_n1237_0[0]));
	jspl3 jspl3_w_n1245_0(.douta(w_n1245_0[0]),.doutb(w_n1245_0[1]),.doutc(w_n1245_0[2]),.din(n1245));
	jspl jspl_w_n1245_1(.douta(w_n1245_1[0]),.doutb(w_n1245_1[1]),.din(w_n1245_0[0]));
	jspl3 jspl3_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.doutc(w_n1248_0[2]),.din(n1248));
	jspl jspl_w_n1248_1(.douta(w_n1248_1[0]),.doutb(w_n1248_1[1]),.din(w_n1248_0[0]));
	jspl3 jspl3_w_n1256_0(.douta(w_n1256_0[0]),.doutb(w_n1256_0[1]),.doutc(w_n1256_0[2]),.din(n1256));
	jspl jspl_w_n1256_1(.douta(w_n1256_1[0]),.doutb(w_n1256_1[1]),.din(w_n1256_0[0]));
	jspl3 jspl3_w_n1264_0(.douta(w_n1264_0[0]),.doutb(w_n1264_0[1]),.doutc(w_n1264_0[2]),.din(n1264));
	jspl jspl_w_n1264_1(.douta(w_n1264_1[0]),.doutb(w_n1264_1[1]),.din(w_n1264_0[0]));
	jspl3 jspl3_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.doutc(w_n1273_0[2]),.din(n1273));
	jspl jspl_w_n1273_1(.douta(w_n1273_1[0]),.doutb(w_n1273_1[1]),.din(w_n1273_0[0]));
	jspl3 jspl3_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.doutc(w_n1281_0[2]),.din(n1281));
	jspl jspl_w_n1281_1(.douta(w_n1281_1[0]),.doutb(w_n1281_1[1]),.din(w_n1281_0[0]));
	jspl3 jspl3_w_n1284_0(.douta(w_n1284_0[0]),.doutb(w_n1284_0[1]),.doutc(w_n1284_0[2]),.din(n1284));
	jspl jspl_w_n1284_1(.douta(w_n1284_1[0]),.doutb(w_n1284_1[1]),.din(w_n1284_0[0]));
	jspl3 jspl3_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.doutc(w_n1293_0[2]),.din(n1293));
	jspl jspl_w_n1293_1(.douta(w_n1293_1[0]),.doutb(w_n1293_1[1]),.din(w_n1293_0[0]));
	jspl3 jspl3_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.doutc(w_n1301_0[2]),.din(n1301));
	jspl jspl_w_n1301_1(.douta(w_n1301_1[0]),.doutb(w_n1301_1[1]),.din(w_n1301_0[0]));
	jspl3 jspl3_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.doutc(w_n1310_0[2]),.din(n1310));
	jspl jspl_w_n1310_1(.douta(w_n1310_1[0]),.doutb(w_n1310_1[1]),.din(w_n1310_0[0]));
	jspl3 jspl3_w_n1318_0(.douta(w_n1318_0[0]),.doutb(w_n1318_0[1]),.doutc(w_n1318_0[2]),.din(n1318));
	jspl jspl_w_n1318_1(.douta(w_n1318_1[0]),.doutb(w_n1318_1[1]),.din(w_n1318_0[0]));
	jspl3 jspl3_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.doutc(w_n1321_0[2]),.din(n1321));
	jspl jspl_w_n1321_1(.douta(w_n1321_1[0]),.doutb(w_n1321_1[1]),.din(w_n1321_0[0]));
	jspl3 jspl3_w_n1329_0(.douta(w_n1329_0[0]),.doutb(w_n1329_0[1]),.doutc(w_n1329_0[2]),.din(n1329));
	jspl jspl_w_n1329_1(.douta(w_n1329_1[0]),.doutb(w_n1329_1[1]),.din(w_n1329_0[0]));
	jspl3 jspl3_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.doutc(w_n1337_0[2]),.din(n1337));
	jspl jspl_w_n1337_1(.douta(w_n1337_1[0]),.doutb(w_n1337_1[1]),.din(w_n1337_0[0]));
	jspl3 jspl3_w_n1346_0(.douta(w_n1346_0[0]),.doutb(w_n1346_0[1]),.doutc(w_n1346_0[2]),.din(n1346));
	jspl jspl_w_n1346_1(.douta(w_n1346_1[0]),.doutb(w_n1346_1[1]),.din(w_n1346_0[0]));
	jspl3 jspl3_w_n1354_0(.douta(w_n1354_0[0]),.doutb(w_n1354_0[1]),.doutc(w_n1354_0[2]),.din(n1354));
	jspl jspl_w_n1354_1(.douta(w_n1354_1[0]),.doutb(w_n1354_1[1]),.din(w_n1354_0[0]));
	jspl3 jspl3_w_n1357_0(.douta(w_n1357_0[0]),.doutb(w_n1357_0[1]),.doutc(w_n1357_0[2]),.din(n1357));
	jspl jspl_w_n1357_1(.douta(w_n1357_1[0]),.doutb(w_n1357_1[1]),.din(w_n1357_0[0]));
	jspl jspl_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.din(n1360));
	jspl3 jspl3_w_n1365_0(.douta(w_n1365_0[0]),.doutb(w_n1365_0[1]),.doutc(w_n1365_0[2]),.din(n1365));
	jspl jspl_w_n1365_1(.douta(w_n1365_1[0]),.doutb(w_n1365_1[1]),.din(w_n1365_0[0]));
	jspl3 jspl3_w_n1369_0(.douta(w_n1369_0[0]),.doutb(w_n1369_0[1]),.doutc(w_n1369_0[2]),.din(n1369));
	jspl jspl_w_n1369_1(.douta(w_n1369_1[0]),.doutb(w_n1369_1[1]),.din(w_n1369_0[0]));
	jspl3 jspl3_w_n1374_0(.douta(w_n1374_0[0]),.doutb(w_n1374_0[1]),.doutc(w_n1374_0[2]),.din(n1374));
	jspl jspl_w_n1374_1(.douta(w_n1374_1[0]),.doutb(w_n1374_1[1]),.din(w_n1374_0[0]));
	jspl3 jspl3_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.doutc(w_n1378_0[2]),.din(n1378));
	jspl jspl_w_n1378_1(.douta(w_n1378_1[0]),.doutb(w_n1378_1[1]),.din(w_n1378_0[0]));
	jspl3 jspl3_w_n1381_0(.douta(w_n1381_0[0]),.doutb(w_n1381_0[1]),.doutc(w_n1381_0[2]),.din(n1381));
	jspl jspl_w_n1381_1(.douta(w_n1381_1[0]),.doutb(w_n1381_1[1]),.din(w_n1381_0[0]));
	jspl3 jspl3_w_n1385_0(.douta(w_n1385_0[0]),.doutb(w_n1385_0[1]),.doutc(w_n1385_0[2]),.din(n1385));
	jspl jspl_w_n1385_1(.douta(w_n1385_1[0]),.doutb(w_n1385_1[1]),.din(w_n1385_0[0]));
	jspl3 jspl3_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.doutc(w_n1389_0[2]),.din(n1389));
	jspl jspl_w_n1389_1(.douta(w_n1389_1[0]),.doutb(w_n1389_1[1]),.din(w_n1389_0[0]));
	jspl3 jspl3_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.doutc(w_n1394_0[2]),.din(n1394));
	jspl jspl_w_n1394_1(.douta(w_n1394_1[0]),.doutb(w_n1394_1[1]),.din(w_n1394_0[0]));
	jspl3 jspl3_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.doutc(w_n1398_0[2]),.din(n1398));
	jspl jspl_w_n1398_1(.douta(w_n1398_1[0]),.doutb(w_n1398_1[1]),.din(w_n1398_0[0]));
	jspl3 jspl3_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_n1401_0[1]),.doutc(w_n1401_0[2]),.din(n1401));
	jspl jspl_w_n1401_1(.douta(w_n1401_1[0]),.doutb(w_n1401_1[1]),.din(w_n1401_0[0]));
	jspl3 jspl3_w_n1406_0(.douta(w_n1406_0[0]),.doutb(w_n1406_0[1]),.doutc(w_n1406_0[2]),.din(n1406));
	jspl jspl_w_n1406_1(.douta(w_n1406_1[0]),.doutb(w_n1406_1[1]),.din(w_n1406_0[0]));
	jspl3 jspl3_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.doutc(w_n1410_0[2]),.din(n1410));
	jspl jspl_w_n1410_1(.douta(w_n1410_1[0]),.doutb(w_n1410_1[1]),.din(w_n1410_0[0]));
	jspl3 jspl3_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.doutc(w_n1415_0[2]),.din(n1415));
	jspl jspl_w_n1415_1(.douta(w_n1415_1[0]),.doutb(w_n1415_1[1]),.din(w_n1415_0[0]));
	jspl3 jspl3_w_n1419_0(.douta(w_n1419_0[0]),.doutb(w_n1419_0[1]),.doutc(w_n1419_0[2]),.din(n1419));
	jspl jspl_w_n1419_1(.douta(w_n1419_1[0]),.doutb(w_n1419_1[1]),.din(w_n1419_0[0]));
	jspl3 jspl3_w_n1422_0(.douta(w_n1422_0[0]),.doutb(w_n1422_0[1]),.doutc(w_n1422_0[2]),.din(n1422));
	jspl jspl_w_n1422_1(.douta(w_n1422_1[0]),.doutb(w_n1422_1[1]),.din(w_n1422_0[0]));
	jspl3 jspl3_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.doutc(w_n1426_0[2]),.din(n1426));
	jspl jspl_w_n1426_1(.douta(w_n1426_1[0]),.doutb(w_n1426_1[1]),.din(w_n1426_0[0]));
	jspl3 jspl3_w_n1430_0(.douta(w_n1430_0[0]),.doutb(w_n1430_0[1]),.doutc(w_n1430_0[2]),.din(n1430));
	jspl jspl_w_n1430_1(.douta(w_n1430_1[0]),.doutb(w_n1430_1[1]),.din(w_n1430_0[0]));
	jspl3 jspl3_w_n1435_0(.douta(w_n1435_0[0]),.doutb(w_n1435_0[1]),.doutc(w_n1435_0[2]),.din(n1435));
	jspl jspl_w_n1435_1(.douta(w_n1435_1[0]),.doutb(w_n1435_1[1]),.din(w_n1435_0[0]));
	jspl3 jspl3_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.doutc(w_n1439_0[2]),.din(n1439));
	jspl jspl_w_n1439_1(.douta(w_n1439_1[0]),.doutb(w_n1439_1[1]),.din(w_n1439_0[0]));
	jspl3 jspl3_w_n1442_0(.douta(w_n1442_0[0]),.doutb(w_n1442_0[1]),.doutc(w_n1442_0[2]),.din(n1442));
	jspl jspl_w_n1442_1(.douta(w_n1442_1[0]),.doutb(w_n1442_1[1]),.din(w_n1442_0[0]));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl3 jspl3_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.doutc(w_n1449_0[2]),.din(n1449));
	jspl jspl_w_n1449_1(.douta(w_n1449_1[0]),.doutb(w_n1449_1[1]),.din(w_n1449_0[0]));
	jspl3 jspl3_w_n1453_0(.douta(w_n1453_0[0]),.doutb(w_n1453_0[1]),.doutc(w_n1453_0[2]),.din(n1453));
	jspl jspl_w_n1453_1(.douta(w_n1453_1[0]),.doutb(w_n1453_1[1]),.din(w_n1453_0[0]));
	jspl3 jspl3_w_n1458_0(.douta(w_n1458_0[0]),.doutb(w_n1458_0[1]),.doutc(w_n1458_0[2]),.din(n1458));
	jspl jspl_w_n1458_1(.douta(w_n1458_1[0]),.doutb(w_n1458_1[1]),.din(w_n1458_0[0]));
	jspl3 jspl3_w_n1462_0(.douta(w_n1462_0[0]),.doutb(w_n1462_0[1]),.doutc(w_n1462_0[2]),.din(n1462));
	jspl jspl_w_n1462_1(.douta(w_n1462_1[0]),.doutb(w_n1462_1[1]),.din(w_n1462_0[0]));
	jspl3 jspl3_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.doutc(w_n1465_0[2]),.din(n1465));
	jspl jspl_w_n1465_1(.douta(w_n1465_1[0]),.doutb(w_n1465_1[1]),.din(w_n1465_0[0]));
	jspl3 jspl3_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.doutc(w_n1469_0[2]),.din(n1469));
	jspl jspl_w_n1469_1(.douta(w_n1469_1[0]),.doutb(w_n1469_1[1]),.din(w_n1469_0[0]));
	jspl3 jspl3_w_n1473_0(.douta(w_n1473_0[0]),.doutb(w_n1473_0[1]),.doutc(w_n1473_0[2]),.din(n1473));
	jspl jspl_w_n1473_1(.douta(w_n1473_1[0]),.doutb(w_n1473_1[1]),.din(w_n1473_0[0]));
	jspl3 jspl3_w_n1478_0(.douta(w_n1478_0[0]),.doutb(w_n1478_0[1]),.doutc(w_n1478_0[2]),.din(n1478));
	jspl jspl_w_n1478_1(.douta(w_n1478_1[0]),.doutb(w_n1478_1[1]),.din(w_n1478_0[0]));
	jspl3 jspl3_w_n1482_0(.douta(w_n1482_0[0]),.doutb(w_n1482_0[1]),.doutc(w_n1482_0[2]),.din(n1482));
	jspl jspl_w_n1482_1(.douta(w_n1482_1[0]),.doutb(w_n1482_1[1]),.din(w_n1482_0[0]));
	jspl3 jspl3_w_n1485_0(.douta(w_n1485_0[0]),.doutb(w_n1485_0[1]),.doutc(w_n1485_0[2]),.din(n1485));
	jspl jspl_w_n1485_1(.douta(w_n1485_1[0]),.doutb(w_n1485_1[1]),.din(w_n1485_0[0]));
	jspl3 jspl3_w_n1490_0(.douta(w_n1490_0[0]),.doutb(w_n1490_0[1]),.doutc(w_n1490_0[2]),.din(n1490));
	jspl jspl_w_n1490_1(.douta(w_n1490_1[0]),.doutb(w_n1490_1[1]),.din(w_n1490_0[0]));
	jspl3 jspl3_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.doutc(w_n1496_0[2]),.din(n1496));
	jspl jspl_w_n1496_1(.douta(w_n1496_1[0]),.doutb(w_n1496_1[1]),.din(w_n1496_0[0]));
	jspl3 jspl3_w_n1505_0(.douta(w_n1505_0[0]),.doutb(w_n1505_0[1]),.doutc(w_n1505_0[2]),.din(n1505));
	jspl jspl_w_n1505_1(.douta(w_n1505_1[0]),.doutb(w_n1505_1[1]),.din(w_n1505_0[0]));
	jspl3 jspl3_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.doutc(w_n1510_0[2]),.din(n1510));
	jspl jspl_w_n1510_1(.douta(w_n1510_1[0]),.doutb(w_n1510_1[1]),.din(w_n1510_0[0]));
	jspl3 jspl3_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.doutc(w_n1513_0[2]),.din(n1513));
	jspl jspl_w_n1513_1(.douta(w_n1513_1[0]),.doutb(w_n1513_1[1]),.din(w_n1513_0[0]));
	jspl3 jspl3_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.doutc(w_n1517_0[2]),.din(n1517));
	jspl jspl_w_n1517_1(.douta(w_n1517_1[0]),.doutb(w_n1517_1[1]),.din(w_n1517_0[0]));
	jspl3 jspl3_w_n1521_0(.douta(w_n1521_0[0]),.doutb(w_n1521_0[1]),.doutc(w_n1521_0[2]),.din(n1521));
	jspl jspl_w_n1521_1(.douta(w_n1521_1[0]),.doutb(w_n1521_1[1]),.din(w_n1521_0[0]));
	jspl3 jspl3_w_n1526_0(.douta(w_n1526_0[0]),.doutb(w_n1526_0[1]),.doutc(w_n1526_0[2]),.din(n1526));
	jspl jspl_w_n1526_1(.douta(w_n1526_1[0]),.doutb(w_n1526_1[1]),.din(w_n1526_0[0]));
	jspl3 jspl3_w_n1530_0(.douta(w_n1530_0[0]),.doutb(w_n1530_0[1]),.doutc(w_n1530_0[2]),.din(n1530));
	jspl jspl_w_n1530_1(.douta(w_n1530_1[0]),.doutb(w_n1530_1[1]),.din(w_n1530_0[0]));
	jspl3 jspl3_w_n1533_0(.douta(w_n1533_0[0]),.doutb(w_n1533_0[1]),.doutc(w_n1533_0[2]),.din(n1533));
	jspl jspl_w_n1533_1(.douta(w_n1533_1[0]),.doutb(w_n1533_1[1]),.din(w_n1533_0[0]));
	jspl jspl_w_n1536_0(.douta(w_n1536_0[0]),.doutb(w_n1536_0[1]),.din(n1536));
	jspl3 jspl3_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.doutc(w_n1545_0[2]),.din(n1545));
	jspl jspl_w_n1545_1(.douta(w_n1545_1[0]),.doutb(w_n1545_1[1]),.din(w_n1545_0[0]));
	jspl3 jspl3_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.doutc(w_n1553_0[2]),.din(n1553));
	jspl jspl_w_n1553_1(.douta(w_n1553_1[0]),.doutb(w_n1553_1[1]),.din(w_n1553_0[0]));
	jspl3 jspl3_w_n1562_0(.douta(w_n1562_0[0]),.doutb(w_n1562_0[1]),.doutc(w_n1562_0[2]),.din(n1562));
	jspl jspl_w_n1562_1(.douta(w_n1562_1[0]),.doutb(w_n1562_1[1]),.din(w_n1562_0[0]));
	jspl3 jspl3_w_n1570_0(.douta(w_n1570_0[0]),.doutb(w_n1570_0[1]),.doutc(w_n1570_0[2]),.din(n1570));
	jspl jspl_w_n1570_1(.douta(w_n1570_1[0]),.doutb(w_n1570_1[1]),.din(w_n1570_0[0]));
	jspl jspl_w_n1573_0(.douta(w_n1573_0[0]),.doutb(w_n1573_0[1]),.din(n1573));
	jspl3 jspl3_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_n1581_0[1]),.doutc(w_n1581_0[2]),.din(n1581));
	jspl jspl_w_n1581_1(.douta(w_n1581_1[0]),.doutb(w_n1581_1[1]),.din(w_n1581_0[0]));
	jspl3 jspl3_w_n1589_0(.douta(w_n1589_0[0]),.doutb(w_n1589_0[1]),.doutc(w_n1589_0[2]),.din(n1589));
	jspl jspl_w_n1589_1(.douta(w_n1589_1[0]),.doutb(w_n1589_1[1]),.din(w_n1589_0[0]));
	jspl3 jspl3_w_n1598_0(.douta(w_n1598_0[0]),.doutb(w_n1598_0[1]),.doutc(w_n1598_0[2]),.din(n1598));
	jspl jspl_w_n1598_1(.douta(w_n1598_1[0]),.doutb(w_n1598_1[1]),.din(w_n1598_0[0]));
	jspl3 jspl3_w_n1606_0(.douta(w_n1606_0[0]),.doutb(w_n1606_0[1]),.doutc(w_n1606_0[2]),.din(n1606));
	jspl jspl_w_n1606_1(.douta(w_n1606_1[0]),.doutb(w_n1606_1[1]),.din(w_n1606_0[0]));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl3 jspl3_w_n1618_0(.douta(w_n1618_0[0]),.doutb(w_n1618_0[1]),.doutc(w_n1618_0[2]),.din(n1618));
	jspl jspl_w_n1618_1(.douta(w_n1618_1[0]),.doutb(w_n1618_1[1]),.din(w_n1618_0[0]));
	jspl3 jspl3_w_n1626_0(.douta(w_n1626_0[0]),.doutb(w_n1626_0[1]),.doutc(w_n1626_0[2]),.din(n1626));
	jspl jspl_w_n1626_1(.douta(w_n1626_1[0]),.doutb(w_n1626_1[1]),.din(w_n1626_0[0]));
	jspl3 jspl3_w_n1635_0(.douta(w_n1635_0[0]),.doutb(w_n1635_0[1]),.doutc(w_n1635_0[2]),.din(n1635));
	jspl jspl_w_n1635_1(.douta(w_n1635_1[0]),.doutb(w_n1635_1[1]),.din(w_n1635_0[0]));
	jspl3 jspl3_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.doutc(w_n1643_0[2]),.din(n1643));
	jspl jspl_w_n1643_1(.douta(w_n1643_1[0]),.doutb(w_n1643_1[1]),.din(w_n1643_0[0]));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(n1646));
	jspl3 jspl3_w_n1654_0(.douta(w_n1654_0[0]),.doutb(w_n1654_0[1]),.doutc(w_n1654_0[2]),.din(n1654));
	jspl jspl_w_n1654_1(.douta(w_n1654_1[0]),.doutb(w_n1654_1[1]),.din(w_n1654_0[0]));
	jspl3 jspl3_w_n1662_0(.douta(w_n1662_0[0]),.doutb(w_n1662_0[1]),.doutc(w_n1662_0[2]),.din(n1662));
	jspl jspl_w_n1662_1(.douta(w_n1662_1[0]),.doutb(w_n1662_1[1]),.din(w_n1662_0[0]));
	jspl3 jspl3_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.doutc(w_n1671_0[2]),.din(n1671));
	jspl jspl_w_n1671_1(.douta(w_n1671_1[0]),.doutb(w_n1671_1[1]),.din(w_n1671_0[0]));
	jspl3 jspl3_w_n1679_0(.douta(w_n1679_0[0]),.doutb(w_n1679_0[1]),.doutc(w_n1679_0[2]),.din(n1679));
	jspl jspl_w_n1679_1(.douta(w_n1679_1[0]),.doutb(w_n1679_1[1]),.din(w_n1679_0[0]));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(n1682));
	jspl3 jspl3_w_n1691_0(.douta(w_n1691_0[0]),.doutb(w_n1691_0[1]),.doutc(w_n1691_0[2]),.din(n1691));
	jspl jspl_w_n1691_1(.douta(w_n1691_1[0]),.doutb(w_n1691_1[1]),.din(w_n1691_0[0]));
	jspl3 jspl3_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.doutc(w_n1699_0[2]),.din(n1699));
	jspl jspl_w_n1699_1(.douta(w_n1699_1[0]),.doutb(w_n1699_1[1]),.din(w_n1699_0[0]));
	jspl3 jspl3_w_n1708_0(.douta(w_n1708_0[0]),.doutb(w_n1708_0[1]),.doutc(w_n1708_0[2]),.din(n1708));
	jspl jspl_w_n1708_1(.douta(w_n1708_1[0]),.doutb(w_n1708_1[1]),.din(w_n1708_0[0]));
	jspl3 jspl3_w_n1716_0(.douta(w_n1716_0[0]),.doutb(w_n1716_0[1]),.doutc(w_n1716_0[2]),.din(n1716));
	jspl jspl_w_n1716_1(.douta(w_n1716_1[0]),.doutb(w_n1716_1[1]),.din(w_n1716_0[0]));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl3 jspl3_w_n1727_0(.douta(w_n1727_0[0]),.doutb(w_n1727_0[1]),.doutc(w_n1727_0[2]),.din(n1727));
	jspl jspl_w_n1727_1(.douta(w_n1727_1[0]),.doutb(w_n1727_1[1]),.din(w_n1727_0[0]));
	jspl3 jspl3_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.doutc(w_n1735_0[2]),.din(n1735));
	jspl jspl_w_n1735_1(.douta(w_n1735_1[0]),.doutb(w_n1735_1[1]),.din(w_n1735_0[0]));
	jspl3 jspl3_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.doutc(w_n1744_0[2]),.din(n1744));
	jspl jspl_w_n1744_1(.douta(w_n1744_1[0]),.doutb(w_n1744_1[1]),.din(w_n1744_0[0]));
	jspl3 jspl3_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.doutc(w_n1752_0[2]),.din(n1752));
	jspl jspl_w_n1752_1(.douta(w_n1752_1[0]),.doutb(w_n1752_1[1]),.din(w_n1752_0[0]));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl3 jspl3_w_n1764_0(.douta(w_n1764_0[0]),.doutb(w_n1764_0[1]),.doutc(w_n1764_0[2]),.din(n1764));
	jspl jspl_w_n1764_1(.douta(w_n1764_1[0]),.doutb(w_n1764_1[1]),.din(w_n1764_0[0]));
	jspl3 jspl3_w_n1772_0(.douta(w_n1772_0[0]),.doutb(w_n1772_0[1]),.doutc(w_n1772_0[2]),.din(n1772));
	jspl jspl_w_n1772_1(.douta(w_n1772_1[0]),.doutb(w_n1772_1[1]),.din(w_n1772_0[0]));
	jspl3 jspl3_w_n1781_0(.douta(w_n1781_0[0]),.doutb(w_n1781_0[1]),.doutc(w_n1781_0[2]),.din(n1781));
	jspl jspl_w_n1781_1(.douta(w_n1781_1[0]),.doutb(w_n1781_1[1]),.din(w_n1781_0[0]));
	jspl3 jspl3_w_n1789_0(.douta(w_n1789_0[0]),.doutb(w_n1789_0[1]),.doutc(w_n1789_0[2]),.din(n1789));
	jspl jspl_w_n1789_1(.douta(w_n1789_1[0]),.doutb(w_n1789_1[1]),.din(w_n1789_0[0]));
	jspl jspl_w_n1792_0(.douta(w_n1792_0[0]),.doutb(w_n1792_0[1]),.din(n1792));
	jspl3 jspl3_w_n1800_0(.douta(w_n1800_0[0]),.doutb(w_n1800_0[1]),.doutc(w_n1800_0[2]),.din(n1800));
	jspl jspl_w_n1800_1(.douta(w_n1800_1[0]),.doutb(w_n1800_1[1]),.din(w_n1800_0[0]));
	jspl3 jspl3_w_n1808_0(.douta(w_n1808_0[0]),.doutb(w_n1808_0[1]),.doutc(w_n1808_0[2]),.din(n1808));
	jspl jspl_w_n1808_1(.douta(w_n1808_1[0]),.doutb(w_n1808_1[1]),.din(w_n1808_0[0]));
	jspl3 jspl3_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_n1817_0[1]),.doutc(w_n1817_0[2]),.din(n1817));
	jspl jspl_w_n1817_1(.douta(w_n1817_1[0]),.doutb(w_n1817_1[1]),.din(w_n1817_0[0]));
	jspl3 jspl3_w_n1825_0(.douta(w_n1825_0[0]),.doutb(w_n1825_0[1]),.doutc(w_n1825_0[2]),.din(n1825));
	jspl jspl_w_n1825_1(.douta(w_n1825_1[0]),.doutb(w_n1825_1[1]),.din(w_n1825_0[0]));
	jspl jspl_w_n1828_0(.douta(w_n1828_0[0]),.doutb(w_n1828_0[1]),.din(n1828));
	jspl3 jspl3_w_n1837_0(.douta(w_n1837_0[0]),.doutb(w_n1837_0[1]),.doutc(w_n1837_0[2]),.din(n1837));
	jspl jspl_w_n1837_1(.douta(w_n1837_1[0]),.doutb(w_n1837_1[1]),.din(w_n1837_0[0]));
	jspl3 jspl3_w_n1845_0(.douta(w_n1845_0[0]),.doutb(w_n1845_0[1]),.doutc(w_n1845_0[2]),.din(n1845));
	jspl jspl_w_n1845_1(.douta(w_n1845_1[0]),.doutb(w_n1845_1[1]),.din(w_n1845_0[0]));
	jspl3 jspl3_w_n1854_0(.douta(w_n1854_0[0]),.doutb(w_n1854_0[1]),.doutc(w_n1854_0[2]),.din(n1854));
	jspl jspl_w_n1854_1(.douta(w_n1854_1[0]),.doutb(w_n1854_1[1]),.din(w_n1854_0[0]));
	jspl3 jspl3_w_n1862_0(.douta(w_n1862_0[0]),.doutb(w_n1862_0[1]),.doutc(w_n1862_0[2]),.din(n1862));
	jspl jspl_w_n1862_1(.douta(w_n1862_1[0]),.doutb(w_n1862_1[1]),.din(w_n1862_0[0]));
	jspl jspl_w_n1865_0(.douta(w_n1865_0[0]),.doutb(w_n1865_0[1]),.din(n1865));
	jspl3 jspl3_w_n1873_0(.douta(w_n1873_0[0]),.doutb(w_n1873_0[1]),.doutc(w_n1873_0[2]),.din(n1873));
	jspl jspl_w_n1873_1(.douta(w_n1873_1[0]),.doutb(w_n1873_1[1]),.din(w_n1873_0[0]));
	jspl3 jspl3_w_n1881_0(.douta(w_n1881_0[0]),.doutb(w_n1881_0[1]),.doutc(w_n1881_0[2]),.din(n1881));
	jspl jspl_w_n1881_1(.douta(w_n1881_1[0]),.doutb(w_n1881_1[1]),.din(w_n1881_0[0]));
	jspl3 jspl3_w_n1890_0(.douta(w_n1890_0[0]),.doutb(w_n1890_0[1]),.doutc(w_n1890_0[2]),.din(n1890));
	jspl jspl_w_n1890_1(.douta(w_n1890_1[0]),.doutb(w_n1890_1[1]),.din(w_n1890_0[0]));
	jspl3 jspl3_w_n1898_0(.douta(w_n1898_0[0]),.doutb(w_n1898_0[1]),.doutc(w_n1898_0[2]),.din(n1898));
	jspl jspl_w_n1898_1(.douta(w_n1898_1[0]),.doutb(w_n1898_1[1]),.din(w_n1898_0[0]));
	jspl jspl_w_n1901_0(.douta(w_n1901_0[0]),.doutb(w_n1901_0[1]),.din(n1901));
	jspl3 jspl3_w_n1910_0(.douta(w_n1910_0[0]),.doutb(w_n1910_0[1]),.doutc(w_n1910_0[2]),.din(n1910));
	jspl jspl_w_n1910_1(.douta(w_n1910_1[0]),.doutb(w_n1910_1[1]),.din(w_n1910_0[0]));
	jspl3 jspl3_w_n1918_0(.douta(w_n1918_0[0]),.doutb(w_n1918_0[1]),.doutc(w_n1918_0[2]),.din(n1918));
	jspl jspl_w_n1918_1(.douta(w_n1918_1[0]),.doutb(w_n1918_1[1]),.din(w_n1918_0[0]));
	jspl3 jspl3_w_n1927_0(.douta(w_n1927_0[0]),.doutb(w_n1927_0[1]),.doutc(w_n1927_0[2]),.din(n1927));
	jspl jspl_w_n1927_1(.douta(w_n1927_1[0]),.doutb(w_n1927_1[1]),.din(w_n1927_0[0]));
	jspl3 jspl3_w_n1935_0(.douta(w_n1935_0[0]),.doutb(w_n1935_0[1]),.doutc(w_n1935_0[2]),.din(n1935));
	jspl jspl_w_n1935_1(.douta(w_n1935_1[0]),.doutb(w_n1935_1[1]),.din(w_n1935_0[0]));
	jspl jspl_w_n1938_0(.douta(w_n1938_0[0]),.doutb(w_n1938_0[1]),.din(n1938));
	jspl3 jspl3_w_n1946_0(.douta(w_n1946_0[0]),.doutb(w_n1946_0[1]),.doutc(w_n1946_0[2]),.din(n1946));
	jspl jspl_w_n1946_1(.douta(w_n1946_1[0]),.doutb(w_n1946_1[1]),.din(w_n1946_0[0]));
	jspl3 jspl3_w_n1954_0(.douta(w_n1954_0[0]),.doutb(w_n1954_0[1]),.doutc(w_n1954_0[2]),.din(n1954));
	jspl jspl_w_n1954_1(.douta(w_n1954_1[0]),.doutb(w_n1954_1[1]),.din(w_n1954_0[0]));
	jspl3 jspl3_w_n1963_0(.douta(w_n1963_0[0]),.doutb(w_n1963_0[1]),.doutc(w_n1963_0[2]),.din(n1963));
	jspl jspl_w_n1963_1(.douta(w_n1963_1[0]),.doutb(w_n1963_1[1]),.din(w_n1963_0[0]));
	jspl3 jspl3_w_n1971_0(.douta(w_n1971_0[0]),.doutb(w_n1971_0[1]),.doutc(w_n1971_0[2]),.din(n1971));
	jspl jspl_w_n1971_1(.douta(w_n1971_1[0]),.doutb(w_n1971_1[1]),.din(w_n1971_0[0]));
	jspl jspl_w_n1974_0(.douta(w_n1974_0[0]),.doutb(w_n1974_0[1]),.din(n1974));
	jspl3 jspl3_w_n1983_0(.douta(w_n1983_0[0]),.doutb(w_n1983_0[1]),.doutc(w_n1983_0[2]),.din(n1983));
	jspl jspl_w_n1983_1(.douta(w_n1983_1[0]),.doutb(w_n1983_1[1]),.din(w_n1983_0[0]));
	jspl3 jspl3_w_n1991_0(.douta(w_n1991_0[0]),.doutb(w_n1991_0[1]),.doutc(w_n1991_0[2]),.din(n1991));
	jspl jspl_w_n1991_1(.douta(w_n1991_1[0]),.doutb(w_n1991_1[1]),.din(w_n1991_0[0]));
	jspl3 jspl3_w_n2000_0(.douta(w_n2000_0[0]),.doutb(w_n2000_0[1]),.doutc(w_n2000_0[2]),.din(n2000));
	jspl jspl_w_n2000_1(.douta(w_n2000_1[0]),.doutb(w_n2000_1[1]),.din(w_n2000_0[0]));
	jspl3 jspl3_w_n2008_0(.douta(w_n2008_0[0]),.doutb(w_n2008_0[1]),.doutc(w_n2008_0[2]),.din(n2008));
	jspl jspl_w_n2008_1(.douta(w_n2008_1[0]),.doutb(w_n2008_1[1]),.din(w_n2008_0[0]));
	jspl jspl_w_n2011_0(.douta(w_n2011_0[0]),.doutb(w_n2011_0[1]),.din(n2011));
	jspl3 jspl3_w_n2019_0(.douta(w_n2019_0[0]),.doutb(w_n2019_0[1]),.doutc(w_n2019_0[2]),.din(n2019));
	jspl jspl_w_n2019_1(.douta(w_n2019_1[0]),.doutb(w_n2019_1[1]),.din(w_n2019_0[0]));
	jspl3 jspl3_w_n2027_0(.douta(w_n2027_0[0]),.doutb(w_n2027_0[1]),.doutc(w_n2027_0[2]),.din(n2027));
	jspl jspl_w_n2027_1(.douta(w_n2027_1[0]),.doutb(w_n2027_1[1]),.din(w_n2027_0[0]));
	jspl3 jspl3_w_n2036_0(.douta(w_n2036_0[0]),.doutb(w_n2036_0[1]),.doutc(w_n2036_0[2]),.din(n2036));
	jspl jspl_w_n2036_1(.douta(w_n2036_1[0]),.doutb(w_n2036_1[1]),.din(w_n2036_0[0]));
	jspl3 jspl3_w_n2044_0(.douta(w_n2044_0[0]),.doutb(w_n2044_0[1]),.doutc(w_n2044_0[2]),.din(n2044));
	jspl jspl_w_n2044_1(.douta(w_n2044_1[0]),.doutb(w_n2044_1[1]),.din(w_n2044_0[0]));
	jspl jspl_w_n2047_0(.douta(w_n2047_0[0]),.doutb(w_n2047_0[1]),.din(n2047));
	jspl3 jspl3_w_n2056_0(.douta(w_n2056_0[0]),.doutb(w_n2056_0[1]),.doutc(w_n2056_0[2]),.din(n2056));
	jspl jspl_w_n2056_1(.douta(w_n2056_1[0]),.doutb(w_n2056_1[1]),.din(w_n2056_0[0]));
	jspl3 jspl3_w_n2064_0(.douta(w_n2064_0[0]),.doutb(w_n2064_0[1]),.doutc(w_n2064_0[2]),.din(n2064));
	jspl jspl_w_n2064_1(.douta(w_n2064_1[0]),.doutb(w_n2064_1[1]),.din(w_n2064_0[0]));
	jspl3 jspl3_w_n2073_0(.douta(w_n2073_0[0]),.doutb(w_n2073_0[1]),.doutc(w_n2073_0[2]),.din(n2073));
	jspl jspl_w_n2073_1(.douta(w_n2073_1[0]),.doutb(w_n2073_1[1]),.din(w_n2073_0[0]));
	jspl3 jspl3_w_n2081_0(.douta(w_n2081_0[0]),.doutb(w_n2081_0[1]),.doutc(w_n2081_0[2]),.din(n2081));
	jspl jspl_w_n2081_1(.douta(w_n2081_1[0]),.doutb(w_n2081_1[1]),.din(w_n2081_0[0]));
	jspl jspl_w_n2084_0(.douta(w_n2084_0[0]),.doutb(w_n2084_0[1]),.din(n2084));
	jspl3 jspl3_w_n2092_0(.douta(w_n2092_0[0]),.doutb(w_n2092_0[1]),.doutc(w_n2092_0[2]),.din(n2092));
	jspl jspl_w_n2092_1(.douta(w_n2092_1[0]),.doutb(w_n2092_1[1]),.din(w_n2092_0[0]));
	jspl3 jspl3_w_n2100_0(.douta(w_n2100_0[0]),.doutb(w_n2100_0[1]),.doutc(w_n2100_0[2]),.din(n2100));
	jspl jspl_w_n2100_1(.douta(w_n2100_1[0]),.doutb(w_n2100_1[1]),.din(w_n2100_0[0]));
	jspl3 jspl3_w_n2109_0(.douta(w_n2109_0[0]),.doutb(w_n2109_0[1]),.doutc(w_n2109_0[2]),.din(n2109));
	jspl jspl_w_n2109_1(.douta(w_n2109_1[0]),.doutb(w_n2109_1[1]),.din(w_n2109_0[0]));
	jspl3 jspl3_w_n2117_0(.douta(w_n2117_0[0]),.doutb(w_n2117_0[1]),.doutc(w_n2117_0[2]),.din(n2117));
	jspl jspl_w_n2117_1(.douta(w_n2117_1[0]),.doutb(w_n2117_1[1]),.din(w_n2117_0[0]));
	jspl jspl_w_n2120_0(.douta(w_n2120_0[0]),.doutb(w_n2120_0[1]),.din(n2120));
	jspl3 jspl3_w_n2129_0(.douta(w_n2129_0[0]),.doutb(w_n2129_0[1]),.doutc(w_n2129_0[2]),.din(n2129));
	jspl jspl_w_n2129_1(.douta(w_n2129_1[0]),.doutb(w_n2129_1[1]),.din(w_n2129_0[0]));
	jspl3 jspl3_w_n2137_0(.douta(w_n2137_0[0]),.doutb(w_n2137_0[1]),.doutc(w_n2137_0[2]),.din(n2137));
	jspl jspl_w_n2137_1(.douta(w_n2137_1[0]),.doutb(w_n2137_1[1]),.din(w_n2137_0[0]));
	jspl3 jspl3_w_n2146_0(.douta(w_n2146_0[0]),.doutb(w_n2146_0[1]),.doutc(w_n2146_0[2]),.din(n2146));
	jspl jspl_w_n2146_1(.douta(w_n2146_1[0]),.doutb(w_n2146_1[1]),.din(w_n2146_0[0]));
	jspl3 jspl3_w_n2154_0(.douta(w_n2154_0[0]),.doutb(w_n2154_0[1]),.doutc(w_n2154_0[2]),.din(n2154));
	jspl jspl_w_n2154_1(.douta(w_n2154_1[0]),.doutb(w_n2154_1[1]),.din(w_n2154_0[0]));
	jspl jspl_w_n2157_0(.douta(w_n2157_0[0]),.doutb(w_n2157_0[1]),.din(n2157));
	jspl3 jspl3_w_n2165_0(.douta(w_n2165_0[0]),.doutb(w_n2165_0[1]),.doutc(w_n2165_0[2]),.din(n2165));
	jspl jspl_w_n2165_1(.douta(w_n2165_1[0]),.doutb(w_n2165_1[1]),.din(w_n2165_0[0]));
	jspl3 jspl3_w_n2173_0(.douta(w_n2173_0[0]),.doutb(w_n2173_0[1]),.doutc(w_n2173_0[2]),.din(n2173));
	jspl jspl_w_n2173_1(.douta(w_n2173_1[0]),.doutb(w_n2173_1[1]),.din(w_n2173_0[0]));
	jspl3 jspl3_w_n2182_0(.douta(w_n2182_0[0]),.doutb(w_n2182_0[1]),.doutc(w_n2182_0[2]),.din(n2182));
	jspl jspl_w_n2182_1(.douta(w_n2182_1[0]),.doutb(w_n2182_1[1]),.din(w_n2182_0[0]));
	jspl3 jspl3_w_n2190_0(.douta(w_n2190_0[0]),.doutb(w_n2190_0[1]),.doutc(w_n2190_0[2]),.din(n2190));
	jspl jspl_w_n2190_1(.douta(w_n2190_1[0]),.doutb(w_n2190_1[1]),.din(w_n2190_0[0]));
	jspl jspl_w_n2193_0(.douta(w_n2193_0[0]),.doutb(w_n2193_0[1]),.din(n2193));
	jspl3 jspl3_w_n2202_0(.douta(w_n2202_0[0]),.doutb(w_n2202_0[1]),.doutc(w_n2202_0[2]),.din(n2202));
	jspl jspl_w_n2202_1(.douta(w_n2202_1[0]),.doutb(w_n2202_1[1]),.din(w_n2202_0[0]));
	jspl3 jspl3_w_n2210_0(.douta(w_n2210_0[0]),.doutb(w_n2210_0[1]),.doutc(w_n2210_0[2]),.din(n2210));
	jspl jspl_w_n2210_1(.douta(w_n2210_1[0]),.doutb(w_n2210_1[1]),.din(w_n2210_0[0]));
	jspl3 jspl3_w_n2219_0(.douta(w_n2219_0[0]),.doutb(w_n2219_0[1]),.doutc(w_n2219_0[2]),.din(n2219));
	jspl jspl_w_n2219_1(.douta(w_n2219_1[0]),.doutb(w_n2219_1[1]),.din(w_n2219_0[0]));
	jspl3 jspl3_w_n2227_0(.douta(w_n2227_0[0]),.doutb(w_n2227_0[1]),.doutc(w_n2227_0[2]),.din(n2227));
	jspl jspl_w_n2227_1(.douta(w_n2227_1[0]),.doutb(w_n2227_1[1]),.din(w_n2227_0[0]));
	jspl jspl_w_n2230_0(.douta(w_n2230_0[0]),.doutb(w_n2230_0[1]),.din(n2230));
	jspl3 jspl3_w_n2238_0(.douta(w_n2238_0[0]),.doutb(w_n2238_0[1]),.doutc(w_n2238_0[2]),.din(n2238));
	jspl jspl_w_n2238_1(.douta(w_n2238_1[0]),.doutb(w_n2238_1[1]),.din(w_n2238_0[0]));
	jspl3 jspl3_w_n2246_0(.douta(w_n2246_0[0]),.doutb(w_n2246_0[1]),.doutc(w_n2246_0[2]),.din(n2246));
	jspl jspl_w_n2246_1(.douta(w_n2246_1[0]),.doutb(w_n2246_1[1]),.din(w_n2246_0[0]));
	jspl3 jspl3_w_n2255_0(.douta(w_n2255_0[0]),.doutb(w_n2255_0[1]),.doutc(w_n2255_0[2]),.din(n2255));
	jspl jspl_w_n2255_1(.douta(w_n2255_1[0]),.doutb(w_n2255_1[1]),.din(w_n2255_0[0]));
	jspl3 jspl3_w_n2263_0(.douta(w_n2263_0[0]),.doutb(w_n2263_0[1]),.doutc(w_n2263_0[2]),.din(n2263));
	jspl jspl_w_n2263_1(.douta(w_n2263_1[0]),.doutb(w_n2263_1[1]),.din(w_n2263_0[0]));
	jspl jspl_w_n2266_0(.douta(w_n2266_0[0]),.doutb(w_n2266_0[1]),.din(n2266));
	jspl3 jspl3_w_n2275_0(.douta(w_n2275_0[0]),.doutb(w_n2275_0[1]),.doutc(w_n2275_0[2]),.din(n2275));
	jspl jspl_w_n2275_1(.douta(w_n2275_1[0]),.doutb(w_n2275_1[1]),.din(w_n2275_0[0]));
	jspl3 jspl3_w_n2283_0(.douta(w_n2283_0[0]),.doutb(w_n2283_0[1]),.doutc(w_n2283_0[2]),.din(n2283));
	jspl jspl_w_n2283_1(.douta(w_n2283_1[0]),.doutb(w_n2283_1[1]),.din(w_n2283_0[0]));
	jspl3 jspl3_w_n2292_0(.douta(w_n2292_0[0]),.doutb(w_n2292_0[1]),.doutc(w_n2292_0[2]),.din(n2292));
	jspl jspl_w_n2292_1(.douta(w_n2292_1[0]),.doutb(w_n2292_1[1]),.din(w_n2292_0[0]));
	jspl3 jspl3_w_n2300_0(.douta(w_n2300_0[0]),.doutb(w_n2300_0[1]),.doutc(w_n2300_0[2]),.din(n2300));
	jspl jspl_w_n2300_1(.douta(w_n2300_1[0]),.doutb(w_n2300_1[1]),.din(w_n2300_0[0]));
	jspl jspl_w_n2303_0(.douta(w_n2303_0[0]),.doutb(w_n2303_0[1]),.din(n2303));
	jspl3 jspl3_w_n2311_0(.douta(w_n2311_0[0]),.doutb(w_n2311_0[1]),.doutc(w_n2311_0[2]),.din(n2311));
	jspl jspl_w_n2311_1(.douta(w_n2311_1[0]),.doutb(w_n2311_1[1]),.din(w_n2311_0[0]));
	jspl3 jspl3_w_n2319_0(.douta(w_n2319_0[0]),.doutb(w_n2319_0[1]),.doutc(w_n2319_0[2]),.din(n2319));
	jspl jspl_w_n2319_1(.douta(w_n2319_1[0]),.doutb(w_n2319_1[1]),.din(w_n2319_0[0]));
	jspl3 jspl3_w_n2328_0(.douta(w_n2328_0[0]),.doutb(w_n2328_0[1]),.doutc(w_n2328_0[2]),.din(n2328));
	jspl jspl_w_n2328_1(.douta(w_n2328_1[0]),.doutb(w_n2328_1[1]),.din(w_n2328_0[0]));
	jspl3 jspl3_w_n2336_0(.douta(w_n2336_0[0]),.doutb(w_n2336_0[1]),.doutc(w_n2336_0[2]),.din(n2336));
	jspl jspl_w_n2336_1(.douta(w_n2336_1[0]),.doutb(w_n2336_1[1]),.din(w_n2336_0[0]));
	jspl jspl_w_n2339_0(.douta(w_n2339_0[0]),.doutb(w_n2339_0[1]),.din(n2339));
	jspl3 jspl3_w_n2348_0(.douta(w_n2348_0[0]),.doutb(w_n2348_0[1]),.doutc(w_n2348_0[2]),.din(n2348));
	jspl jspl_w_n2348_1(.douta(w_n2348_1[0]),.doutb(w_n2348_1[1]),.din(w_n2348_0[0]));
	jspl3 jspl3_w_n2356_0(.douta(w_n2356_0[0]),.doutb(w_n2356_0[1]),.doutc(w_n2356_0[2]),.din(n2356));
	jspl jspl_w_n2356_1(.douta(w_n2356_1[0]),.doutb(w_n2356_1[1]),.din(w_n2356_0[0]));
	jspl3 jspl3_w_n2365_0(.douta(w_n2365_0[0]),.doutb(w_n2365_0[1]),.doutc(w_n2365_0[2]),.din(n2365));
	jspl jspl_w_n2365_1(.douta(w_n2365_1[0]),.doutb(w_n2365_1[1]),.din(w_n2365_0[0]));
	jspl3 jspl3_w_n2373_0(.douta(w_n2373_0[0]),.doutb(w_n2373_0[1]),.doutc(w_n2373_0[2]),.din(n2373));
	jspl jspl_w_n2373_1(.douta(w_n2373_1[0]),.doutb(w_n2373_1[1]),.din(w_n2373_0[0]));
	jspl jspl_w_n2376_0(.douta(w_n2376_0[0]),.doutb(w_n2376_0[1]),.din(n2376));
	jspl3 jspl3_w_n2384_0(.douta(w_n2384_0[0]),.doutb(w_n2384_0[1]),.doutc(w_n2384_0[2]),.din(n2384));
	jspl jspl_w_n2384_1(.douta(w_n2384_1[0]),.doutb(w_n2384_1[1]),.din(w_n2384_0[0]));
	jspl3 jspl3_w_n2392_0(.douta(w_n2392_0[0]),.doutb(w_n2392_0[1]),.doutc(w_n2392_0[2]),.din(n2392));
	jspl jspl_w_n2392_1(.douta(w_n2392_1[0]),.doutb(w_n2392_1[1]),.din(w_n2392_0[0]));
	jspl3 jspl3_w_n2401_0(.douta(w_n2401_0[0]),.doutb(w_n2401_0[1]),.doutc(w_n2401_0[2]),.din(n2401));
	jspl jspl_w_n2401_1(.douta(w_n2401_1[0]),.doutb(w_n2401_1[1]),.din(w_n2401_0[0]));
	jspl3 jspl3_w_n2409_0(.douta(w_n2409_0[0]),.doutb(w_n2409_0[1]),.doutc(w_n2409_0[2]),.din(n2409));
	jspl jspl_w_n2409_1(.douta(w_n2409_1[0]),.doutb(w_n2409_1[1]),.din(w_n2409_0[0]));
	jspl jspl_w_n2412_0(.douta(w_n2412_0[0]),.doutb(w_n2412_0[1]),.din(n2412));
	jspl jspl_w_n2421_0(.douta(w_n2421_0[0]),.doutb(w_n2421_0[1]),.din(n2421));
	jspl jspl_w_n2429_0(.douta(w_n2429_0[0]),.doutb(w_n2429_0[1]),.din(n2429));
	jspl jspl_w_n2438_0(.douta(w_n2438_0[0]),.doutb(w_n2438_0[1]),.din(n2438));
	jspl jspl_w_n2446_0(.douta(w_n2446_0[0]),.doutb(w_n2446_0[1]),.din(n2446));
	jspl jspl_w_n2455_0(.douta(w_n2455_0[0]),.doutb(w_n2455_0[1]),.din(n2455));
	jspl jspl_w_n2463_0(.douta(w_n2463_0[0]),.doutb(w_n2463_0[1]),.din(n2463));
	jspl jspl_w_n2472_0(.douta(w_n2472_0[0]),.doutb(w_n2472_0[1]),.din(n2472));
	jspl jspl_w_n2480_0(.douta(w_n2480_0[0]),.doutb(w_n2480_0[1]),.din(n2480));
	jspl jspl_w_n2489_0(.douta(w_n2489_0[0]),.doutb(w_n2489_0[1]),.din(n2489));
	jspl jspl_w_n2497_0(.douta(w_n2497_0[0]),.doutb(w_n2497_0[1]),.din(n2497));
	jspl jspl_w_n2506_0(.douta(w_n2506_0[0]),.doutb(w_n2506_0[1]),.din(n2506));
	jspl jspl_w_n2514_0(.douta(w_n2514_0[0]),.doutb(w_n2514_0[1]),.din(n2514));
	jspl jspl_w_n2523_0(.douta(w_n2523_0[0]),.doutb(w_n2523_0[1]),.din(n2523));
	jspl jspl_w_n2531_0(.douta(w_n2531_0[0]),.doutb(w_n2531_0[1]),.din(n2531));
	jspl jspl_w_n2540_0(.douta(w_n2540_0[0]),.doutb(w_n2540_0[1]),.din(n2540));
	jspl jspl_w_n2548_0(.douta(w_n2548_0[0]),.doutb(w_n2548_0[1]),.din(n2548));
	jspl jspl_w_n2557_0(.douta(w_n2557_0[0]),.doutb(w_n2557_0[1]),.din(n2557));
	jspl jspl_w_n2565_0(.douta(w_n2565_0[0]),.doutb(w_n2565_0[1]),.din(n2565));
	jspl jspl_w_n2574_0(.douta(w_n2574_0[0]),.doutb(w_n2574_0[1]),.din(n2574));
	jspl jspl_w_n2582_0(.douta(w_n2582_0[0]),.doutb(w_n2582_0[1]),.din(n2582));
	jspl jspl_w_n2591_0(.douta(w_n2591_0[0]),.doutb(w_n2591_0[1]),.din(n2591));
	jspl jspl_w_n2599_0(.douta(w_n2599_0[0]),.doutb(w_n2599_0[1]),.din(n2599));
	jspl jspl_w_n2608_0(.douta(w_n2608_0[0]),.doutb(w_n2608_0[1]),.din(n2608));
	jspl jspl_w_n2616_0(.douta(w_n2616_0[0]),.doutb(w_n2616_0[1]),.din(n2616));
	jspl jspl_w_n2625_0(.douta(w_n2625_0[0]),.doutb(w_n2625_0[1]),.din(n2625));
	jspl jspl_w_n2633_0(.douta(w_n2633_0[0]),.doutb(w_n2633_0[1]),.din(n2633));
	jspl jspl_w_n2642_0(.douta(w_n2642_0[0]),.doutb(w_n2642_0[1]),.din(n2642));
	jspl jspl_w_n2650_0(.douta(w_n2650_0[0]),.doutb(w_n2650_0[1]),.din(n2650));
	jspl jspl_w_n2659_0(.douta(w_n2659_0[0]),.doutb(w_n2659_0[1]),.din(n2659));
	jspl jspl_w_n2667_0(.douta(w_n2667_0[0]),.doutb(w_n2667_0[1]),.din(n2667));
	jspl jspl_w_n2676_0(.douta(w_n2676_0[0]),.doutb(w_n2676_0[1]),.din(n2676));
	jspl jspl_w_n2684_0(.douta(w_n2684_0[0]),.doutb(w_n2684_0[1]),.din(n2684));
	jspl jspl_w_n2693_0(.douta(w_n2693_0[0]),.doutb(w_n2693_0[1]),.din(n2693));
	jspl jspl_w_n2701_0(.douta(w_n2701_0[0]),.doutb(w_n2701_0[1]),.din(n2701));
	jspl jspl_w_n2710_0(.douta(w_n2710_0[0]),.doutb(w_n2710_0[1]),.din(n2710));
	jspl jspl_w_n2718_0(.douta(w_n2718_0[0]),.doutb(w_n2718_0[1]),.din(n2718));
	jspl jspl_w_n2727_0(.douta(w_n2727_0[0]),.doutb(w_n2727_0[1]),.din(n2727));
	jspl jspl_w_n2735_0(.douta(w_n2735_0[0]),.doutb(w_n2735_0[1]),.din(n2735));
	jspl jspl_w_n2744_0(.douta(w_n2744_0[0]),.doutb(w_n2744_0[1]),.din(n2744));
	jspl jspl_w_n2752_0(.douta(w_n2752_0[0]),.doutb(w_n2752_0[1]),.din(n2752));
	jspl jspl_w_n2761_0(.douta(w_n2761_0[0]),.doutb(w_n2761_0[1]),.din(n2761));
	jspl jspl_w_n2769_0(.douta(w_n2769_0[0]),.doutb(w_n2769_0[1]),.din(n2769));
	jspl jspl_w_n2778_0(.douta(w_n2778_0[0]),.doutb(w_n2778_0[1]),.din(n2778));
	jspl jspl_w_n2786_0(.douta(w_n2786_0[0]),.doutb(w_n2786_0[1]),.din(n2786));
	jspl jspl_w_n2795_0(.douta(w_n2795_0[0]),.doutb(w_n2795_0[1]),.din(n2795));
	jspl jspl_w_n2803_0(.douta(w_n2803_0[0]),.doutb(w_n2803_0[1]),.din(n2803));
	jspl jspl_w_n2812_0(.douta(w_n2812_0[0]),.doutb(w_n2812_0[1]),.din(n2812));
	jspl jspl_w_n2820_0(.douta(w_n2820_0[0]),.doutb(w_n2820_0[1]),.din(n2820));
	jspl jspl_w_n2829_0(.douta(w_n2829_0[0]),.doutb(w_n2829_0[1]),.din(n2829));
	jspl jspl_w_n2837_0(.douta(w_n2837_0[0]),.doutb(w_n2837_0[1]),.din(n2837));
	jspl jspl_w_n2846_0(.douta(w_n2846_0[0]),.doutb(w_n2846_0[1]),.din(n2846));
	jspl jspl_w_n2854_0(.douta(w_n2854_0[0]),.doutb(w_n2854_0[1]),.din(n2854));
	jspl jspl_w_n2863_0(.douta(w_n2863_0[0]),.doutb(w_n2863_0[1]),.din(n2863));
	jspl jspl_w_n2871_0(.douta(w_n2871_0[0]),.doutb(w_n2871_0[1]),.din(n2871));
	jspl jspl_w_n2880_0(.douta(w_n2880_0[0]),.doutb(w_n2880_0[1]),.din(n2880));
	jspl jspl_w_n2888_0(.douta(w_n2888_0[0]),.doutb(w_n2888_0[1]),.din(n2888));
	jspl jspl_w_n2897_0(.douta(w_n2897_0[0]),.doutb(w_n2897_0[1]),.din(n2897));
	jspl jspl_w_n2905_0(.douta(w_n2905_0[0]),.doutb(w_n2905_0[1]),.din(n2905));
	jspl jspl_w_n2914_0(.douta(w_n2914_0[0]),.doutb(w_n2914_0[1]),.din(n2914));
	jspl jspl_w_n2922_0(.douta(w_n2922_0[0]),.doutb(w_n2922_0[1]),.din(n2922));
	jspl jspl_w_n2931_0(.douta(w_n2931_0[0]),.doutb(w_n2931_0[1]),.din(n2931));
	jspl jspl_w_n2939_0(.douta(w_n2939_0[0]),.doutb(w_n2939_0[1]),.din(n2939));
	jspl jspl_w_n2948_0(.douta(w_n2948_0[0]),.doutb(w_n2948_0[1]),.din(n2948));
	jspl jspl_w_n2956_0(.douta(w_n2956_0[0]),.doutb(w_n2956_0[1]),.din(n2956));
	jspl jspl_w_n2965_0(.douta(w_n2965_0[0]),.doutb(w_n2965_0[1]),.din(n2965));
	jspl jspl_w_n2973_0(.douta(w_n2973_0[0]),.doutb(w_n2973_0[1]),.din(n2973));
	jspl jspl_w_n2982_0(.douta(w_n2982_0[0]),.doutb(w_n2982_0[1]),.din(n2982));
	jspl jspl_w_n2990_0(.douta(w_n2990_0[0]),.doutb(w_n2990_0[1]),.din(n2990));
	jspl jspl_w_n2999_0(.douta(w_n2999_0[0]),.doutb(w_n2999_0[1]),.din(n2999));
	jspl jspl_w_n3007_0(.douta(w_n3007_0[0]),.doutb(w_n3007_0[1]),.din(n3007));
	jspl jspl_w_n3016_0(.douta(w_n3016_0[0]),.doutb(w_n3016_0[1]),.din(n3016));
	jspl jspl_w_n3024_0(.douta(w_n3024_0[0]),.doutb(w_n3024_0[1]),.din(n3024));
	jspl jspl_w_n3033_0(.douta(w_n3033_0[0]),.doutb(w_n3033_0[1]),.din(n3033));
	jspl jspl_w_n3041_0(.douta(w_n3041_0[0]),.doutb(w_n3041_0[1]),.din(n3041));
	jspl jspl_w_n3050_0(.douta(w_n3050_0[0]),.doutb(w_n3050_0[1]),.din(n3050));
	jspl jspl_w_n3058_0(.douta(w_n3058_0[0]),.doutb(w_n3058_0[1]),.din(n3058));
	jspl jspl_w_n3067_0(.douta(w_n3067_0[0]),.doutb(w_n3067_0[1]),.din(n3067));
	jspl jspl_w_n3075_0(.douta(w_n3075_0[0]),.doutb(w_n3075_0[1]),.din(n3075));
	jspl jspl_w_n3084_0(.douta(w_n3084_0[0]),.doutb(w_n3084_0[1]),.din(n3084));
	jspl jspl_w_n3092_0(.douta(w_n3092_0[0]),.doutb(w_n3092_0[1]),.din(n3092));
	jspl jspl_w_n3101_0(.douta(w_n3101_0[0]),.doutb(w_n3101_0[1]),.din(n3101));
	jspl jspl_w_n3109_0(.douta(w_n3109_0[0]),.doutb(w_n3109_0[1]),.din(n3109));
	jspl jspl_w_n3118_0(.douta(w_n3118_0[0]),.doutb(w_n3118_0[1]),.din(n3118));
	jspl jspl_w_n3126_0(.douta(w_n3126_0[0]),.doutb(w_n3126_0[1]),.din(n3126));
	jspl jspl_w_n3135_0(.douta(w_n3135_0[0]),.doutb(w_n3135_0[1]),.din(n3135));
	jspl jspl_w_n3143_0(.douta(w_n3143_0[0]),.doutb(w_n3143_0[1]),.din(n3143));
	jspl jspl_w_n3152_0(.douta(w_n3152_0[0]),.doutb(w_n3152_0[1]),.din(n3152));
	jspl jspl_w_n3160_0(.douta(w_n3160_0[0]),.doutb(w_n3160_0[1]),.din(n3160));
	jspl jspl_w_n3169_0(.douta(w_n3169_0[0]),.doutb(w_n3169_0[1]),.din(n3169));
	jspl jspl_w_n3177_0(.douta(w_n3177_0[0]),.doutb(w_n3177_0[1]),.din(n3177));
	jspl jspl_w_n3186_0(.douta(w_n3186_0[0]),.doutb(w_n3186_0[1]),.din(n3186));
	jspl jspl_w_n3194_0(.douta(w_n3194_0[0]),.doutb(w_n3194_0[1]),.din(n3194));
	jspl jspl_w_n3203_0(.douta(w_n3203_0[0]),.doutb(w_n3203_0[1]),.din(n3203));
	jspl jspl_w_n3211_0(.douta(w_n3211_0[0]),.doutb(w_n3211_0[1]),.din(n3211));
	jspl jspl_w_n3220_0(.douta(w_n3220_0[0]),.doutb(w_n3220_0[1]),.din(n3220));
	jspl jspl_w_n3228_0(.douta(w_n3228_0[0]),.doutb(w_n3228_0[1]),.din(n3228));
endmodule

