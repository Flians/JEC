/*

c880:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jdff: 1588
	jand: 151
	jor: 122

Summary:
	jxor: 26
	jspl: 85
	jspl3: 90
	jnot: 48
	jdff: 1588
	jand: 151
	jor: 122
*/

module c880(gclk, G1gat, G8gat, G13gat, G17gat, G26gat, G29gat, G36gat, G42gat, G51gat, G55gat, G59gat, G68gat, G72gat, G73gat, G74gat, G75gat, G80gat, G85gat, G86gat, G87gat, G88gat, G89gat, G90gat, G91gat, G96gat, G101gat, G106gat, G111gat, G116gat, G121gat, G126gat, G130gat, G135gat, G138gat, G143gat, G146gat, G149gat, G152gat, G153gat, G156gat, G159gat, G165gat, G171gat, G177gat, G183gat, G189gat, G195gat, G201gat, G207gat, G210gat, G219gat, G228gat, G237gat, G246gat, G255gat, G259gat, G260gat, G261gat, G267gat, G268gat, G388gat, G389gat, G390gat, G391gat, G418gat, G419gat, G420gat, G421gat, G422gat, G423gat, G446gat, G447gat, G448gat, G449gat, G450gat, G767gat, G768gat, G850gat, G863gat, G864gat, G865gat, G866gat, G874gat, G878gat, G879gat, G880gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G13gat;
	input G17gat;
	input G26gat;
	input G29gat;
	input G36gat;
	input G42gat;
	input G51gat;
	input G55gat;
	input G59gat;
	input G68gat;
	input G72gat;
	input G73gat;
	input G74gat;
	input G75gat;
	input G80gat;
	input G85gat;
	input G86gat;
	input G87gat;
	input G88gat;
	input G89gat;
	input G90gat;
	input G91gat;
	input G96gat;
	input G101gat;
	input G106gat;
	input G111gat;
	input G116gat;
	input G121gat;
	input G126gat;
	input G130gat;
	input G135gat;
	input G138gat;
	input G143gat;
	input G146gat;
	input G149gat;
	input G152gat;
	input G153gat;
	input G156gat;
	input G159gat;
	input G165gat;
	input G171gat;
	input G177gat;
	input G183gat;
	input G189gat;
	input G195gat;
	input G201gat;
	input G207gat;
	input G210gat;
	input G219gat;
	input G228gat;
	input G237gat;
	input G246gat;
	input G255gat;
	input G259gat;
	input G260gat;
	input G261gat;
	input G267gat;
	input G268gat;
	output G388gat;
	output G389gat;
	output G390gat;
	output G391gat;
	output G418gat;
	output G419gat;
	output G420gat;
	output G421gat;
	output G422gat;
	output G423gat;
	output G446gat;
	output G447gat;
	output G448gat;
	output G449gat;
	output G450gat;
	output G767gat;
	output G768gat;
	output G850gat;
	output G863gat;
	output G864gat;
	output G865gat;
	output G866gat;
	output G874gat;
	output G878gat;
	output G879gat;
	output G880gat;
	wire n86;
	wire n88;
	wire n92;
	wire n93;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n103;
	wire n104;
	wire n105;
	wire n107;
	wire n108;
	wire n109;
	wire n111;
	wire n113;
	wire n115;
	wire n117;
	wire n119;
	wire n120;
	wire n122;
	wire n123;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire [2:0] w_G1gat_0;
	wire [1:0] w_G1gat_1;
	wire [1:0] w_G8gat_0;
	wire [1:0] w_G13gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G17gat_1;
	wire [2:0] w_G17gat_2;
	wire [1:0] w_G26gat_0;
	wire [2:0] w_G29gat_0;
	wire [1:0] w_G36gat_0;
	wire [2:0] w_G42gat_0;
	wire [2:0] w_G42gat_1;
	wire [1:0] w_G42gat_2;
	wire [2:0] w_G51gat_0;
	wire [1:0] w_G51gat_1;
	wire [2:0] w_G55gat_0;
	wire [2:0] w_G59gat_0;
	wire [1:0] w_G59gat_1;
	wire [1:0] w_G68gat_0;
	wire [1:0] w_G75gat_0;
	wire [2:0] w_G80gat_0;
	wire [2:0] w_G91gat_0;
	wire [2:0] w_G96gat_0;
	wire [2:0] w_G101gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G111gat_0;
	wire [2:0] w_G116gat_0;
	wire [2:0] w_G121gat_0;
	wire [2:0] w_G126gat_0;
	wire [1:0] w_G130gat_0;
	wire [2:0] w_G138gat_0;
	wire [1:0] w_G138gat_1;
	wire [1:0] w_G143gat_0;
	wire [1:0] w_G146gat_0;
	wire [1:0] w_G149gat_0;
	wire [2:0] w_G153gat_0;
	wire [1:0] w_G156gat_0;
	wire [2:0] w_G159gat_0;
	wire [2:0] w_G159gat_1;
	wire [2:0] w_G165gat_0;
	wire [2:0] w_G165gat_1;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [2:0] w_G177gat_0;
	wire [2:0] w_G177gat_1;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G183gat_1;
	wire [2:0] w_G189gat_0;
	wire [2:0] w_G189gat_1;
	wire [1:0] w_G189gat_2;
	wire [2:0] w_G195gat_0;
	wire [2:0] w_G195gat_1;
	wire [1:0] w_G195gat_2;
	wire [2:0] w_G201gat_0;
	wire [1:0] w_G201gat_1;
	wire [2:0] w_G210gat_0;
	wire [2:0] w_G210gat_1;
	wire [2:0] w_G210gat_2;
	wire [1:0] w_G210gat_3;
	wire [2:0] w_G219gat_0;
	wire [2:0] w_G219gat_1;
	wire [2:0] w_G219gat_2;
	wire [2:0] w_G219gat_3;
	wire [2:0] w_G228gat_0;
	wire [2:0] w_G228gat_1;
	wire [2:0] w_G228gat_2;
	wire [1:0] w_G228gat_3;
	wire [2:0] w_G237gat_0;
	wire [2:0] w_G237gat_1;
	wire [2:0] w_G237gat_2;
	wire [1:0] w_G237gat_3;
	wire [2:0] w_G246gat_0;
	wire [2:0] w_G246gat_1;
	wire [2:0] w_G246gat_2;
	wire [1:0] w_G246gat_3;
	wire [2:0] w_G255gat_0;
	wire [2:0] w_G261gat_0;
	wire [1:0] w_G268gat_0;
	wire [1:0] w_G390gat_0;
	wire G390gat_fa_;
	wire [2:0] w_G447gat_0;
	wire w_G447gat_1;
	wire G447gat_fa_;
	wire [1:0] w_n86_0;
	wire [1:0] w_n88_0;
	wire [1:0] w_n92_0;
	wire [1:0] w_n93_0;
	wire [2:0] w_n95_0;
	wire [1:0] w_n97_0;
	wire [1:0] w_n99_0;
	wire [1:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n109_0;
	wire [1:0] w_n111_0;
	wire [1:0] w_n113_0;
	wire [2:0] w_n119_0;
	wire [1:0] w_n122_0;
	wire [1:0] w_n144_0;
	wire [1:0] w_n146_0;
	wire [2:0] w_n148_0;
	wire [2:0] w_n148_1;
	wire [1:0] w_n149_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n152_0;
	wire [1:0] w_n162_0;
	wire [2:0] w_n164_0;
	wire [2:0] w_n164_1;
	wire [2:0] w_n164_2;
	wire [1:0] w_n164_3;
	wire [1:0] w_n167_0;
	wire [1:0] w_n168_0;
	wire [2:0] w_n170_0;
	wire [1:0] w_n170_1;
	wire [1:0] w_n173_0;
	wire [2:0] w_n178_0;
	wire [2:0] w_n178_1;
	wire [2:0] w_n178_2;
	wire [1:0] w_n178_3;
	wire [2:0] w_n181_0;
	wire [1:0] w_n185_0;
	wire [2:0] w_n197_0;
	wire [2:0] w_n198_0;
	wire [1:0] w_n200_0;
	wire [1:0] w_n209_0;
	wire [2:0] w_n218_0;
	wire [1:0] w_n218_1;
	wire [2:0] w_n219_0;
	wire [2:0] w_n222_0;
	wire [2:0] w_n233_0;
	wire [1:0] w_n233_1;
	wire [1:0] w_n234_0;
	wire [1:0] w_n235_0;
	wire [2:0] w_n239_0;
	wire [1:0] w_n239_1;
	wire [1:0] w_n240_0;
	wire [1:0] w_n241_0;
	wire [1:0] w_n242_0;
	wire [1:0] w_n245_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n258_0;
	wire [1:0] w_n260_0;
	wire [1:0] w_n262_0;
	wire [2:0] w_n267_0;
	wire [2:0] w_n285_0;
	wire [2:0] w_n303_0;
	wire [1:0] w_n303_1;
	wire [2:0] w_n306_0;
	wire [1:0] w_n306_1;
	wire [2:0] w_n311_0;
	wire [2:0] w_n311_1;
	wire [2:0] w_n319_0;
	wire [2:0] w_n319_1;
	wire [1:0] w_n320_0;
	wire [1:0] w_n321_0;
	wire [2:0] w_n327_0;
	wire [2:0] w_n327_1;
	wire [1:0] w_n328_0;
	wire [1:0] w_n329_0;
	wire [2:0] w_n335_0;
	wire [1:0] w_n335_1;
	wire [2:0] w_n336_0;
	wire [1:0] w_n339_0;
	wire [1:0] w_n343_0;
	wire [1:0] w_n346_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n350_0;
	wire [1:0] w_n352_0;
	wire [1:0] w_n355_0;
	wire [1:0] w_n361_0;
	wire [2:0] w_n377_0;
	wire [1:0] w_n391_0;
	wire [1:0] w_n393_0;
	wire [2:0] w_n404_0;
	wire [2:0] w_n420_0;
	wire w_dff_B_7UlRVwTw9_2;
	wire w_dff_B_jm6eXLIy3_1;
	wire w_dff_B_UsegxPG92_1;
	wire w_dff_B_rCIjOu890_1;
	wire w_dff_A_Mp84KvMm0_1;
	wire w_dff_A_qZXECBCX7_1;
	wire w_dff_B_tjY6mTfZ5_1;
	wire w_dff_B_8XYJYpfg6_1;
	wire w_dff_B_WVTmUIe00_1;
	wire w_dff_B_iwGeSgRi3_1;
	wire w_dff_B_Ul7hI5tG2_1;
	wire w_dff_B_rPt4A9FB8_1;
	wire w_dff_B_7qFlguCr1_1;
	wire w_dff_A_t3vhnhtj8_1;
	wire w_dff_B_GCcZzlST4_1;
	wire w_dff_B_FshnuNUN2_1;
	wire w_dff_B_dweSJyXE7_1;
	wire w_dff_B_RY5HtDGj1_1;
	wire w_dff_B_MfuJcyUF1_1;
	wire w_dff_B_8UW0a6hs8_1;
	wire w_dff_B_WoauTbc81_0;
	wire w_dff_B_YLyCys8s2_0;
	wire w_dff_B_NGwO7JMM5_0;
	wire w_dff_B_hC8WYbeE4_0;
	wire w_dff_B_fM8BQZxK7_0;
	wire w_dff_B_u6fiRcjm4_0;
	wire w_dff_B_yqChSveb7_0;
	wire w_dff_B_1GYBylOX6_0;
	wire w_dff_B_FpHV7IlO9_0;
	wire w_dff_B_dQlbsjPQ2_0;
	wire w_dff_B_mV64A36W0_0;
	wire w_dff_B_q2Mmt25B3_0;
	wire w_dff_B_1SdJrmBv2_0;
	wire w_dff_B_49ONw7UW7_0;
	wire w_dff_A_y76Rzs7J3_0;
	wire w_dff_A_ei1QMaBS2_0;
	wire w_dff_A_WILyofej2_0;
	wire w_dff_A_e6G37ysD6_0;
	wire w_dff_B_q7n4idcE4_1;
	wire w_dff_B_N6Tfx1Ar5_1;
	wire w_dff_B_kDcwAYjq9_1;
	wire w_dff_B_NKZFhnVf6_1;
	wire w_dff_B_u0Hj6Ey13_1;
	wire w_dff_B_chD6sUN56_1;
	wire w_dff_B_Zy4hPM1a2_1;
	wire w_dff_B_6PUZVafV9_1;
	wire w_dff_B_FGQFoZA48_1;
	wire w_dff_B_3MF9MMpJ7_1;
	wire w_dff_B_4S9JlBsT8_1;
	wire w_dff_B_937gr0qJ4_1;
	wire w_dff_B_eNvjwhZd4_1;
	wire w_dff_B_Skhb3sQy7_1;
	wire w_dff_B_4sDERiW18_1;
	wire w_dff_B_3SS9q1EH8_1;
	wire w_dff_B_mzVXuXBw2_1;
	wire w_dff_B_KHPx0GP12_1;
	wire w_dff_B_yrA6AFeh2_1;
	wire w_dff_B_zI0EUErO1_1;
	wire w_dff_B_n6JYwdGJ7_1;
	wire w_dff_B_g0kUmBXv6_0;
	wire w_dff_B_LWQkaye88_0;
	wire w_dff_B_N9NDx65W8_0;
	wire w_dff_B_3uoepQeC1_0;
	wire w_dff_B_0FLcXZ3g0_0;
	wire w_dff_B_YQ2SxZa59_0;
	wire w_dff_B_Rqvbevwl8_0;
	wire w_dff_B_fVBiDBSq8_0;
	wire w_dff_A_WxfrdtCB9_1;
	wire w_dff_A_nES0KIdl6_1;
	wire w_dff_A_5hwc9EMo6_1;
	wire w_dff_A_qyfNGqSj3_1;
	wire w_dff_A_xdnUc8VM1_1;
	wire w_dff_A_RJLwdD6t4_1;
	wire w_dff_A_ElR4gAoP2_1;
	wire w_dff_A_d4bHz1mU6_1;
	wire w_dff_A_3wgMOOQ69_1;
	wire w_dff_A_9fCcpP7I3_0;
	wire w_dff_A_T7XbUg8G8_0;
	wire w_dff_A_Xm1iaeH91_0;
	wire w_dff_A_Hx6YmaQx0_0;
	wire w_dff_A_KxpzTuRX8_1;
	wire w_dff_A_3Ua3kYjk4_1;
	wire w_dff_A_v6aPyT290_1;
	wire w_dff_A_Yx7gMPpu3_1;
	wire w_dff_A_lNxowiTO0_1;
	wire w_dff_A_QXDDZelg7_1;
	wire w_dff_A_qfPZP3rV5_1;
	wire w_dff_A_HC7Nf5MP7_1;
	wire w_dff_A_rksPqlv74_1;
	wire w_dff_B_svI9Jd4Y5_1;
	wire w_dff_B_sNDaXlOl5_1;
	wire w_dff_B_9743cxsy9_1;
	wire w_dff_B_qKHZi9Qz3_1;
	wire w_dff_B_M5R1DhEI3_1;
	wire w_dff_B_EEoS2hDm7_1;
	wire w_dff_B_62diWx547_0;
	wire w_dff_B_dEK1uI2L2_0;
	wire w_dff_B_z2k3bJfc6_0;
	wire w_dff_B_cqmCFRno5_0;
	wire w_dff_A_0lrckFhS8_0;
	wire w_dff_A_O1GOhNL70_0;
	wire w_dff_A_bTSBTNYh3_0;
	wire w_dff_A_xj9rrQLS1_1;
	wire w_dff_A_cOAz7LA88_1;
	wire w_dff_A_eJlvrSJz1_1;
	wire w_dff_A_63S5tTKF5_1;
	wire w_dff_A_2NJtDy212_1;
	wire w_dff_B_UnPMVXid7_1;
	wire w_dff_B_PTxwytmR2_0;
	wire w_dff_B_EeKn8Uay2_0;
	wire w_dff_B_piIehyoL8_0;
	wire w_dff_B_rkhPEvKP7_0;
	wire w_dff_B_N5WUdfXS6_1;
	wire w_dff_B_mpGiSs4C5_1;
	wire w_dff_B_GcVIOolo0_1;
	wire w_dff_B_vrb2f6Eq5_1;
	wire w_dff_B_akiqZQJF7_1;
	wire w_dff_B_RyYg89Tg4_1;
	wire w_dff_B_leIemAES2_1;
	wire w_dff_B_LFFLHu1r9_1;
	wire w_dff_B_AF3tlUxG8_1;
	wire w_dff_B_C224M06e0_1;
	wire w_dff_B_Ck0f7Him3_1;
	wire w_dff_B_Pyg5iKqF8_1;
	wire w_dff_B_TCsd3mpf6_0;
	wire w_dff_B_czOdfPvk2_0;
	wire w_dff_B_mY9Sqhs87_0;
	wire w_dff_B_XFJMWFuF9_0;
	wire w_dff_B_jvq62fAN3_0;
	wire w_dff_B_2tEvSQQL6_0;
	wire w_dff_A_eoQKWcvc0_1;
	wire w_dff_A_vHhr7IKu0_1;
	wire w_dff_A_DOrvQ7ON2_1;
	wire w_dff_A_Hqkzsl6L6_1;
	wire w_dff_A_WuhLNmxI1_1;
	wire w_dff_B_RsEIk6Gb6_1;
	wire w_dff_B_T80HOhX68_1;
	wire w_dff_B_hvvMwwgx5_1;
	wire w_dff_B_fF2QgabW1_1;
	wire w_dff_B_BdyNMImr7_0;
	wire w_dff_B_taFFIebQ6_0;
	wire w_dff_B_wEPRavaN2_1;
	wire w_dff_B_xcvs9gbx6_0;
	wire w_dff_B_ovA5gLQj8_0;
	wire w_dff_B_UCoh4UA02_0;
	wire w_dff_B_XB3EYXri9_0;
	wire w_dff_B_8Biy8HoB6_0;
	wire w_dff_B_4yAYi2zR9_0;
	wire w_dff_B_kddekpHh7_0;
	wire w_dff_B_IaTZyc2r2_0;
	wire w_dff_B_etzueml98_1;
	wire w_dff_B_InCJkVUG4_1;
	wire w_dff_B_mOLi3xb05_1;
	wire w_dff_B_P5yEMZo09_1;
	wire w_dff_B_ze1z8i5u7_1;
	wire w_dff_B_SyRsljGN8_1;
	wire w_dff_B_o8kDHWXS4_1;
	wire w_dff_B_8okNkrcH4_1;
	wire w_dff_B_IX2gNa7v7_0;
	wire w_dff_B_2NDYToDA8_0;
	wire w_dff_B_LrOKdEeB7_0;
	wire w_dff_B_oxQqHDfP1_0;
	wire w_dff_B_E03DlSsn5_0;
	wire w_dff_B_fFdRJIrJ7_0;
	wire w_dff_A_iDbQWpUL7_1;
	wire w_dff_A_1rB99uad4_1;
	wire w_dff_A_rusbvijp6_1;
	wire w_dff_B_kSsJKgwg1_1;
	wire w_dff_B_43B09MBs2_1;
	wire w_dff_B_Op1CpqzH5_1;
	wire w_dff_B_0vWjKmTn5_1;
	wire w_dff_B_cu8ntCVH0_1;
	wire w_dff_B_uc8tjbyv6_1;
	wire w_dff_B_uoBxPFug8_1;
	wire w_dff_B_e7sIoZUy2_1;
	wire w_dff_B_qXp7vjer1_1;
	wire w_dff_B_nUQ1juD46_1;
	wire w_dff_B_Fbs1rSb97_1;
	wire w_dff_B_bkOfII9t6_1;
	wire w_dff_B_IaomOtqn8_1;
	wire w_dff_B_UOxabOif8_1;
	wire w_dff_B_739TqVXR9_1;
	wire w_dff_B_y0EVvG4E1_1;
	wire w_dff_B_LpLr2JyZ2_1;
	wire w_dff_B_I5b885YO1_1;
	wire w_dff_B_d0IVv4Ub4_1;
	wire w_dff_B_beWCevmd1_1;
	wire w_dff_B_KEE8T8tc0_1;
	wire w_dff_B_VGdy73zl8_1;
	wire w_dff_B_5YsVXXsZ7_1;
	wire w_dff_B_sUM1eFew4_1;
	wire w_dff_B_FA4LMIaE2_1;
	wire w_dff_B_uTybdJek4_1;
	wire w_dff_B_NOvm9CIC9_1;
	wire w_dff_B_Ltyj8zTE9_1;
	wire w_dff_B_5CGT7VBX5_1;
	wire w_dff_A_sMswmXfh8_0;
	wire w_dff_A_g1wpCx1M3_0;
	wire w_dff_A_pvIYsaCQ1_0;
	wire w_dff_A_cdhk59nc5_0;
	wire w_dff_A_2iBPq9uz9_0;
	wire w_dff_A_hudM42rt9_0;
	wire w_dff_A_UlSE4vDR4_0;
	wire w_dff_A_5bLlU6QD3_0;
	wire w_dff_A_zhBzgukI2_0;
	wire w_dff_A_Sqhp3Ll85_1;
	wire w_dff_A_4gHLy7o37_1;
	wire w_dff_A_ARIYx2xm2_1;
	wire w_dff_A_WJ1a99Eu2_1;
	wire w_dff_A_CF5LVvPB8_1;
	wire w_dff_A_3Gv9hCnB8_1;
	wire w_dff_A_3fl3KfOT1_1;
	wire w_dff_A_xvf3G3pH2_1;
	wire w_dff_A_7uwBozfY0_1;
	wire w_dff_B_7ml3irGR4_1;
	wire w_dff_B_1j2Q1vXK1_1;
	wire w_dff_B_hdSk64Iz4_0;
	wire w_dff_B_mufPi80S3_0;
	wire w_dff_B_jOm5GwFl3_0;
	wire w_dff_B_5eDNN2EO0_0;
	wire w_dff_B_JCJhpumM3_0;
	wire w_dff_B_cr61jGFc1_0;
	wire w_dff_B_l4r2TkkW4_0;
	wire w_dff_B_ve2Urtnk4_0;
	wire w_dff_B_mzrTgbZ98_0;
	wire w_dff_B_xRbMtTXj2_0;
	wire w_dff_B_I7wZJAGP9_0;
	wire w_dff_B_dNpIQaZa4_0;
	wire w_dff_B_mYeIAa6e7_0;
	wire w_dff_B_ZrWmph8z4_1;
	wire w_dff_B_b78AtUI52_1;
	wire w_dff_B_Uzu2GLJV8_1;
	wire w_dff_B_Tf9lao5j4_1;
	wire w_dff_A_8FX0cMhG3_0;
	wire w_dff_A_cJALGAt54_0;
	wire w_dff_A_JqRJhMZx7_0;
	wire w_dff_A_cT7LEdyK6_0;
	wire w_dff_A_Xzygf2yW8_0;
	wire w_dff_A_t3rNkFgf8_0;
	wire w_dff_A_qMjKUJIc7_0;
	wire w_dff_A_4c2qsVTd9_0;
	wire w_dff_A_ZbXT1eMg1_0;
	wire w_dff_A_nUpXirUW7_0;
	wire w_dff_A_W7RQboxT6_0;
	wire w_dff_A_uvat82rS3_0;
	wire w_dff_A_M8hCgQuY4_0;
	wire w_dff_A_W32VJuG51_0;
	wire w_dff_A_V930wQB33_0;
	wire w_dff_A_xQjEh6la9_0;
	wire w_dff_A_kUbHugkv4_0;
	wire w_dff_A_msuOIyv83_0;
	wire w_dff_A_5QjO1zHm3_0;
	wire w_dff_A_bBt8WHv93_0;
	wire w_dff_A_taTrXRn34_0;
	wire w_dff_A_WExNutIZ2_0;
	wire w_dff_A_6PzrO9ha8_0;
	wire w_dff_A_JDXWOT8h5_0;
	wire w_dff_A_EnobATnd6_0;
	wire w_dff_A_SF9bc0cb3_0;
	wire w_dff_A_S4IMaqBt1_0;
	wire w_dff_A_8lffngNi1_0;
	wire w_dff_B_dnFacWZS8_1;
	wire w_dff_B_ChAj5V7s1_1;
	wire w_dff_B_vcGy6fu08_1;
	wire w_dff_B_YZDxEaTx5_1;
	wire w_dff_B_3o8olskU4_1;
	wire w_dff_B_SAMtjTEq0_1;
	wire w_dff_B_ROjGXolF2_1;
	wire w_dff_B_2d5NJLya1_1;
	wire w_dff_A_HwTXhXM91_0;
	wire w_dff_A_SQ9Ieeev8_0;
	wire w_dff_A_fE1fGi9P7_0;
	wire w_dff_A_2h074jhv1_0;
	wire w_dff_A_LbMPQRS23_0;
	wire w_dff_A_6Y535p2A7_1;
	wire w_dff_A_E5e6dLfm8_1;
	wire w_dff_A_0svlEpfE3_1;
	wire w_dff_A_hQC7yUKo5_1;
	wire w_dff_A_aUXG5iXh7_1;
	wire w_dff_A_sEEF8IXs3_0;
	wire w_dff_A_l8Ou2Oup8_0;
	wire w_dff_A_sLMlHiQa3_0;
	wire w_dff_A_IOMLg2xW7_0;
	wire w_dff_A_hS4x2fMT4_0;
	wire w_dff_A_v00IdZma0_0;
	wire w_dff_A_Y9GoIESn6_0;
	wire w_dff_A_Ml7zHJL61_0;
	wire w_dff_A_LucvfUrM8_0;
	wire w_dff_A_ugG0IBNP3_0;
	wire w_dff_B_hetlFEwP1_1;
	wire w_dff_B_bAsJDF3r8_1;
	wire w_dff_B_CuATVhDw1_1;
	wire w_dff_B_KX6B9jr39_1;
	wire w_dff_B_pycnsQ9g2_1;
	wire w_dff_B_DRk5VQ9g3_1;
	wire w_dff_B_Rp3sBDlO8_1;
	wire w_dff_B_SnILTlOj6_1;
	wire w_dff_B_2Owu4vM60_1;
	wire w_dff_B_5TqY3Od33_1;
	wire w_dff_B_mHLYSgYu5_1;
	wire w_dff_B_E3TxnA6D4_1;
	wire w_dff_B_ySyv817e3_1;
	wire w_dff_B_BOuBIw5n9_1;
	wire w_dff_B_EBZndK3K6_0;
	wire w_dff_B_4HyA0wIj7_0;
	wire w_dff_B_7nSN1BmL7_0;
	wire w_dff_B_Mn4qUrrj7_0;
	wire w_dff_B_0htFlQng5_0;
	wire w_dff_B_fpSwq8P94_0;
	wire w_dff_B_UT5tplb66_0;
	wire w_dff_B_1E6aVRxq1_0;
	wire w_dff_B_QJ13foVS7_0;
	wire w_dff_B_gYq8QZHH3_0;
	wire w_dff_B_GoXSQxgj3_0;
	wire w_dff_B_H8v8jYX84_0;
	wire w_dff_B_QEWIw3vD5_0;
	wire w_dff_B_QRPM9spZ3_1;
	wire w_dff_B_kelSn6tj3_1;
	wire w_dff_B_LuaotrBh6_1;
	wire w_dff_B_T95ZiaqZ8_1;
	wire w_dff_B_KBtDMrJr2_1;
	wire w_dff_B_R2vPl1S98_1;
	wire w_dff_B_TlhEKaBq6_1;
	wire w_dff_B_f9IH6ZEw6_1;
	wire w_dff_B_7iMcDOUP1_1;
	wire w_dff_B_hAv3xOsb5_1;
	wire w_dff_B_KZ88IVSD8_1;
	wire w_dff_B_NCXRkPjm8_1;
	wire w_dff_B_iy63Giph4_1;
	wire w_dff_B_0uytZM3i5_1;
	wire w_dff_B_ILAq4wtu3_1;
	wire w_dff_B_KUj9xLIJ2_1;
	wire w_dff_B_jzw0ZPRT0_1;
	wire w_dff_B_11LjaTYV3_1;
	wire w_dff_B_wyAxp38r0_1;
	wire w_dff_B_U71aS9Tm2_1;
	wire w_dff_B_gdwCuFFa6_1;
	wire w_dff_B_HpV3k66f6_1;
	wire w_dff_B_oMivBNZI9_1;
	wire w_dff_A_UOBezrC63_1;
	wire w_dff_A_tj08DVM04_1;
	wire w_dff_A_GlX34DJ62_1;
	wire w_dff_A_Eq1zp2Dw6_1;
	wire w_dff_A_FfZrgR9U5_1;
	wire w_dff_A_4vPJs7jD0_1;
	wire w_dff_A_46M3CdYD9_1;
	wire w_dff_A_CA4pmh520_1;
	wire w_dff_A_PXVCfAFW4_1;
	wire w_dff_A_xACCcJFQ1_1;
	wire w_dff_A_GxpxLcHC6_1;
	wire w_dff_A_5xKtEQe73_1;
	wire w_dff_A_7n9azYfH2_1;
	wire w_dff_A_VQBmQ5rn6_1;
	wire w_dff_A_79Bw3fkS3_1;
	wire w_dff_A_QHEB5vvC2_1;
	wire w_dff_A_QM3FYHyt2_1;
	wire w_dff_A_hSBQleYN1_1;
	wire w_dff_A_8WffbtJj9_1;
	wire w_dff_A_5XZFMBH08_1;
	wire w_dff_A_M4FMebO84_1;
	wire w_dff_A_lbx1p6qA3_1;
	wire w_dff_A_FtpnX7Gw5_1;
	wire w_dff_A_Pv1iwvnC9_1;
	wire w_dff_A_1Gws1uM55_1;
	wire w_dff_A_XJ8O74G11_0;
	wire w_dff_A_2iVKTzZv7_0;
	wire w_dff_A_YYYq4rAK1_0;
	wire w_dff_A_uFtfOXYX4_0;
	wire w_dff_A_GVEcGpgF3_0;
	wire w_dff_A_q4TbT11D1_0;
	wire w_dff_A_XUXWmUkq8_0;
	wire w_dff_A_DpfGHxbG0_0;
	wire w_dff_A_qGQ6gt3I0_1;
	wire w_dff_A_RyUJF3wM7_1;
	wire w_dff_A_BgrZISZv1_1;
	wire w_dff_A_jgFwIr5U7_1;
	wire w_dff_A_Oc9mLevZ3_1;
	wire w_dff_A_1FZQV4Ma1_1;
	wire w_dff_A_w9yjRRAl0_1;
	wire w_dff_A_0OM3pxNM4_1;
	wire w_dff_B_CuOGcm1S0_1;
	wire w_dff_B_Z0YVqnoq3_0;
	wire w_dff_B_CRcWHqIK8_0;
	wire w_dff_B_9OUsEcae6_0;
	wire w_dff_B_td3bFAe70_0;
	wire w_dff_B_KtuRsVeg7_0;
	wire w_dff_B_qKMce3FS2_0;
	wire w_dff_B_0OwU0sfQ2_0;
	wire w_dff_B_21aDwmQi0_0;
	wire w_dff_B_UmnxBDse4_0;
	wire w_dff_B_TxpAa5yk6_0;
	wire w_dff_B_y2ynUSV36_0;
	wire w_dff_B_biX3YSsp4_0;
	wire w_dff_A_59cUwoyC3_1;
	wire w_dff_A_gVympQoA6_1;
	wire w_dff_A_UFWYzOYZ4_1;
	wire w_dff_A_9aXzQHFG3_1;
	wire w_dff_A_H1v2ywFF4_1;
	wire w_dff_A_JX1KFojR5_1;
	wire w_dff_A_ZcDVxExB4_1;
	wire w_dff_A_32pX3Qta9_1;
	wire w_dff_A_aRe9hpuv5_1;
	wire w_dff_A_LXmpmsgf0_1;
	wire w_dff_A_InLg641k6_1;
	wire w_dff_A_rCpwzjQz6_1;
	wire w_dff_A_CP52tFaI4_1;
	wire w_dff_A_bBur5LSG3_1;
	wire w_dff_B_vetATD6j3_1;
	wire w_dff_B_T0wICkI14_0;
	wire w_dff_B_FANpPhwB5_0;
	wire w_dff_B_10ZvEDF80_0;
	wire w_dff_B_pyicbREB9_0;
	wire w_dff_B_UwvsC6jy9_0;
	wire w_dff_B_Bw7zreyl4_0;
	wire w_dff_B_wWgacB2x5_1;
	wire w_dff_A_NrDX6v2g9_1;
	wire w_dff_A_qesOdUex1_1;
	wire w_dff_A_WkeiUzpd4_1;
	wire w_dff_A_Pd4xpJIf5_1;
	wire w_dff_A_DKQFbzJV8_1;
	wire w_dff_A_03RQZdCF5_1;
	wire w_dff_A_VcOZFsjM3_1;
	wire w_dff_A_7H3GdROP4_1;
	wire w_dff_A_AhPRc8qB6_1;
	wire w_dff_A_Dpyy9W5a8_2;
	wire w_dff_A_r5uO8BJM1_2;
	wire w_dff_A_N1DY7i6J2_2;
	wire w_dff_A_rsIkIIhy3_2;
	wire w_dff_A_4GB2XfD99_2;
	wire w_dff_A_BYklxgVr5_2;
	wire w_dff_A_aOsX3niG4_2;
	wire w_dff_A_D5LscFzv6_2;
	wire w_dff_A_m4bfDoaB5_2;
	wire w_dff_A_xH1AbGAZ5_2;
	wire w_dff_A_7PmScMsT7_2;
	wire w_dff_B_vZh3sQ576_1;
	wire w_dff_B_QbP7DQ4V1_1;
	wire w_dff_B_jieyf3aQ0_1;
	wire w_dff_B_bM3Ld3Co3_1;
	wire w_dff_B_g67Qs0BX0_1;
	wire w_dff_B_Bv12QFqb9_1;
	wire w_dff_B_vgCJhJqx7_1;
	wire w_dff_B_l5h5YGp65_1;
	wire w_dff_B_5046kXT62_1;
	wire w_dff_B_QwRYwze47_1;
	wire w_dff_B_UQrHe30V6_1;
	wire w_dff_B_T5248S5W0_1;
	wire w_dff_B_PtM3Dr2W9_0;
	wire w_dff_B_rjY96nYx6_0;
	wire w_dff_B_8UJVHaaO8_0;
	wire w_dff_B_Ko8ulaEL1_0;
	wire w_dff_B_EFte2PZh5_0;
	wire w_dff_B_O1Og2UUj2_0;
	wire w_dff_B_i93QyhJt3_0;
	wire w_dff_B_LufdEjVa5_0;
	wire w_dff_B_JXcNqjgB5_0;
	wire w_dff_B_rfQbAPgC3_0;
	wire w_dff_B_3qyVJZYN9_0;
	wire w_dff_B_7Pit0s874_1;
	wire w_dff_B_UBCQA1KC5_1;
	wire w_dff_B_JzdIy3vP0_1;
	wire w_dff_B_E7FeexCx6_1;
	wire w_dff_B_iOkVEekg7_1;
	wire w_dff_B_xr8kS8ob6_1;
	wire w_dff_B_1InQcKpH7_1;
	wire w_dff_B_yKijsFl48_1;
	wire w_dff_B_XYGPfLPa7_1;
	wire w_dff_B_pKHPn9e06_1;
	wire w_dff_B_1utYZW6O4_1;
	wire w_dff_B_DHFwIxVo5_1;
	wire w_dff_B_SweBN5zZ6_1;
	wire w_dff_B_sDvaAJgS4_1;
	wire w_dff_B_Grw3UOcM2_1;
	wire w_dff_B_Ql2kUoG23_1;
	wire w_dff_B_wPbLM3uh5_1;
	wire w_dff_B_wk5YgdTi4_1;
	wire w_dff_B_OwT51m6A4_1;
	wire w_dff_A_6VJrT6Q04_1;
	wire w_dff_A_Eeqwj9sL2_1;
	wire w_dff_A_9toAGEIR6_1;
	wire w_dff_A_T12HvpLQ2_1;
	wire w_dff_A_b2vtq1xz3_1;
	wire w_dff_A_iccYKbFn6_1;
	wire w_dff_A_8xgd9K394_1;
	wire w_dff_A_WW5FOQ2g6_1;
	wire w_dff_A_wmBO8hgq5_1;
	wire w_dff_A_SA2XWHV18_1;
	wire w_dff_A_tv7AzjQJ7_1;
	wire w_dff_A_udiWCKmO9_1;
	wire w_dff_A_EIkbPqy40_1;
	wire w_dff_A_fqioc4hn6_1;
	wire w_dff_A_xHhtf05p2_1;
	wire w_dff_A_P2v0pyPP4_1;
	wire w_dff_A_VZWadwJ72_1;
	wire w_dff_A_LlGqN3Mo9_1;
	wire w_dff_A_e5X4VvEw4_1;
	wire w_dff_A_HRj135OL9_1;
	wire w_dff_A_uiynUS0O5_1;
	wire w_dff_A_F0gyBVJH0_0;
	wire w_dff_A_nxGnwvvR9_0;
	wire w_dff_A_CJvQSQl91_0;
	wire w_dff_A_EWNHvqtf6_0;
	wire w_dff_A_dc8ThQtv3_0;
	wire w_dff_A_zCAx90Vt7_0;
	wire w_dff_A_Srky7VtO1_0;
	wire w_dff_A_38k4Dps60_0;
	wire w_dff_A_umCUVVI01_0;
	wire w_dff_A_3KgmhgZJ7_1;
	wire w_dff_A_FGqvfwLq0_1;
	wire w_dff_A_jZIaruy44_1;
	wire w_dff_A_6P1esCKU2_1;
	wire w_dff_A_gXH4ucZ47_1;
	wire w_dff_A_TEcjQdqf6_1;
	wire w_dff_A_N8YKFdqL5_1;
	wire w_dff_A_Ea4uFO2l8_1;
	wire w_dff_A_bcwERkRS3_1;
	wire w_dff_B_ykPKv9fg2_1;
	wire w_dff_B_jfrwmKXx8_0;
	wire w_dff_B_aNK4sIva0_0;
	wire w_dff_B_2grKY5GW2_0;
	wire w_dff_B_omz9XJ0y8_0;
	wire w_dff_B_h0RbNmS50_0;
	wire w_dff_B_wK80aSpe8_0;
	wire w_dff_B_dWQMcvUP9_0;
	wire w_dff_B_tPrZ7pkb8_0;
	wire w_dff_B_3eZQpfrg2_0;
	wire w_dff_B_eJUlmpTO5_0;
	wire w_dff_B_bTXwLdX74_0;
	wire w_dff_B_88IJbZFB0_0;
	wire w_dff_A_8Fw7Cyt83_1;
	wire w_dff_A_djKevLiJ2_1;
	wire w_dff_A_RXeM7CTo8_1;
	wire w_dff_A_s7KWYlr42_1;
	wire w_dff_A_hhccyiDD4_1;
	wire w_dff_A_iRg79Aqh2_1;
	wire w_dff_A_DRcLU07w7_1;
	wire w_dff_A_61nbhmew8_1;
	wire w_dff_A_e5ILXfQq6_1;
	wire w_dff_A_Dl3G6LQf0_1;
	wire w_dff_A_dUSFqEcb6_1;
	wire w_dff_A_b6AHIqUo2_1;
	wire w_dff_A_5VvKMCik3_1;
	wire w_dff_A_rNfMDcpZ5_1;
	wire w_dff_A_XLAPQinO1_1;
	wire w_dff_A_7alIDhDI4_1;
	wire w_dff_A_mKDxqvHc9_1;
	wire w_dff_A_uoaCAX433_1;
	wire w_dff_B_IWySEGWJ5_0;
	wire w_dff_B_OX3LEpD00_0;
	wire w_dff_B_8Fc9rkR46_0;
	wire w_dff_B_TTtzqLXh9_0;
	wire w_dff_B_1NlFHSi64_0;
	wire w_dff_A_2MjEC4Z57_0;
	wire w_dff_A_BNV2YFLi3_0;
	wire w_dff_A_QEAajFoc6_1;
	wire w_dff_A_Aror5NMl5_1;
	wire w_dff_A_EhApnEyJ6_1;
	wire w_dff_A_RPlFmqo16_1;
	wire w_dff_A_bT7jQvhl1_1;
	wire w_dff_A_3amFmrMm6_1;
	wire w_dff_A_MlTYgtO17_1;
	wire w_dff_A_1AgLbiWv4_1;
	wire w_dff_A_k6mPRUsv1_2;
	wire w_dff_A_WxKp6Ttt4_2;
	wire w_dff_A_aXYBMq7V4_2;
	wire w_dff_A_UENpWxHM5_2;
	wire w_dff_A_1w0hamCF8_2;
	wire w_dff_A_PB6FsCxF0_2;
	wire w_dff_A_1qF4CLvp5_2;
	wire w_dff_A_298pn4NC8_2;
	wire w_dff_A_LPDgjxLY2_2;
	wire w_dff_A_bJNZScVw7_2;
	wire w_dff_B_JItRWBQW9_3;
	wire w_dff_B_j3mZBrun8_1;
	wire w_dff_B_SWfn3xHP0_1;
	wire w_dff_B_zv0iiJYS0_1;
	wire w_dff_B_9CdR91dx3_1;
	wire w_dff_B_0B2Kby3U8_1;
	wire w_dff_B_quZmBvAP5_1;
	wire w_dff_B_qYqgYkN95_1;
	wire w_dff_B_fpwSqhsz0_1;
	wire w_dff_B_U0G8QVwx8_1;
	wire w_dff_B_zwOOlXSY7_1;
	wire w_dff_B_aVeVvnDx5_1;
	wire w_dff_B_50nYNajY8_1;
	wire w_dff_B_nQ74u1A52_1;
	wire w_dff_B_sDVeZaKg0_1;
	wire w_dff_B_z8dkGq7T6_1;
	wire w_dff_B_pndSr3IK8_1;
	wire w_dff_B_FoaT62Es1_1;
	wire w_dff_B_w2mCSZRx3_1;
	wire w_dff_B_vYmNCp3o7_1;
	wire w_dff_B_3rD6pZGq8_1;
	wire w_dff_B_2AmrlOwa8_1;
	wire w_dff_B_jracUH0O1_0;
	wire w_dff_A_sPkWwMba2_1;
	wire w_dff_A_xUjB7yms6_1;
	wire w_dff_A_B81bi5UN8_2;
	wire w_dff_A_5Snwdjtc3_2;
	wire w_dff_A_foZW5O332_2;
	wire w_dff_A_dbuGOjr01_2;
	wire w_dff_A_BLjNfsyj6_0;
	wire w_dff_A_gzDGlbFK2_0;
	wire w_dff_A_FJcBoJQt8_0;
	wire w_dff_A_faq1I0Ji9_0;
	wire w_dff_A_QbAPkKYA4_0;
	wire w_dff_A_6SQldnJf4_0;
	wire w_dff_A_nbptmbQi5_0;
	wire w_dff_A_UAygJ8aK3_0;
	wire w_dff_A_QDzD2JfG6_0;
	wire w_dff_A_NplqoaS60_1;
	wire w_dff_B_uk05Dcmc8_3;
	wire w_dff_B_sLop7rVf9_3;
	wire w_dff_B_ANpwJDwI1_3;
	wire w_dff_B_JvU5D3g95_3;
	wire w_dff_B_IIDP34hE8_3;
	wire w_dff_B_kERcH4e84_3;
	wire w_dff_B_k00DyxE73_3;
	wire w_dff_B_w5mZq1nO9_3;
	wire w_dff_B_OPtafDMO3_3;
	wire w_dff_B_Vm5QE5b82_3;
	wire w_dff_B_FLjWXDwp4_3;
	wire w_dff_B_0lpOHo1W6_3;
	wire w_dff_B_sNrNHi2Z1_0;
	wire w_dff_B_WQUWdl4E3_0;
	wire w_dff_B_hNCpO3UZ2_0;
	wire w_dff_B_gOkFCPuS6_0;
	wire w_dff_B_2J2GUgQg6_0;
	wire w_dff_B_R6SoFP8o6_0;
	wire w_dff_B_KW8igGK98_0;
	wire w_dff_B_nsnNKdcK2_0;
	wire w_dff_B_8cj5bpxF6_0;
	wire w_dff_B_oqg5uijF4_1;
	wire w_dff_B_5rUUiEGJ8_1;
	wire w_dff_B_mfTyZGju3_1;
	wire w_dff_B_nRbGTyVN2_1;
	wire w_dff_B_Th2SJlN16_1;
	wire w_dff_B_WtXRA1ld5_1;
	wire w_dff_B_rstrKNJd9_1;
	wire w_dff_B_WBbSlcL66_1;
	wire w_dff_B_P8Amf1Ii6_1;
	wire w_dff_B_oqJwv3pa1_1;
	wire w_dff_B_bizyuQ3c8_1;
	wire w_dff_B_vU79NiWV1_1;
	wire w_dff_B_9OqRy8FR4_1;
	wire w_dff_B_OS01naCz7_1;
	wire w_dff_B_FNU1id9n2_1;
	wire w_dff_B_DOzp6tmT5_1;
	wire w_dff_B_eP1m1TJH8_1;
	wire w_dff_B_9xyLXn9B4_1;
	wire w_dff_B_wlKVFxMU3_1;
	wire w_dff_B_dKGR2FA92_1;
	wire w_dff_B_EA1D05Qk2_1;
	wire w_dff_B_CGyvMpLi8_1;
	wire w_dff_B_OxgmYRwT3_1;
	wire w_dff_B_wSLV5KIX0_1;
	wire w_dff_B_a50DAPam4_1;
	wire w_dff_B_F7IlVEb42_1;
	wire w_dff_B_Zzo3shUD6_1;
	wire w_dff_B_rpB8y5Sp7_1;
	wire w_dff_B_LzIDozHE7_1;
	wire w_dff_A_OMBCyLHr2_1;
	wire w_dff_B_bi6WFPIu5_2;
	wire w_dff_B_8IudweDH8_2;
	wire w_dff_B_Sb1PajTg8_2;
	wire w_dff_B_TkSNEB3m5_2;
	wire w_dff_B_mxpB1oQ99_2;
	wire w_dff_B_2wF5YYm92_2;
	wire w_dff_B_gY9tg5BZ1_2;
	wire w_dff_B_MY5bGOmQ9_2;
	wire w_dff_B_m4CVuFCK4_2;
	wire w_dff_A_OSv6XK8A7_0;
	wire w_dff_A_NWo7Y8IW9_0;
	wire w_dff_A_BKBe6dXk9_0;
	wire w_dff_A_lS9CqEuB1_0;
	wire w_dff_A_TLkUr34r9_0;
	wire w_dff_A_QBERo3H81_0;
	wire w_dff_A_uXqbUymm0_0;
	wire w_dff_A_6aJZEYCH1_0;
	wire w_dff_A_ZDsl5Lcn6_0;
	wire w_dff_A_eW8E8Ysa1_0;
	wire w_dff_A_gvvmMb2i6_2;
	wire w_dff_A_nXia7lYJ7_2;
	wire w_dff_A_jr6JBQgN5_2;
	wire w_dff_A_wC8V2YAR2_2;
	wire w_dff_A_5XdvEl584_2;
	wire w_dff_A_9D3OSMVh9_2;
	wire w_dff_A_Ftvykmck4_2;
	wire w_dff_A_mCwaDtVM6_2;
	wire w_dff_A_WXlMYB3o1_2;
	wire w_dff_A_4uGeR0Mo1_2;
	wire w_dff_A_qtE1DAht0_0;
	wire w_dff_B_qXTKOI5C0_1;
	wire w_dff_B_2cxF5EFe8_1;
	wire w_dff_B_2D3NmVGD1_1;
	wire w_dff_B_khQssahd6_1;
	wire w_dff_B_SVHRydft8_1;
	wire w_dff_B_2ZMWjlJC5_1;
	wire w_dff_B_ewqprN978_1;
	wire w_dff_B_Q0Knbh0l8_1;
	wire w_dff_B_88ohiOGL1_1;
	wire w_dff_B_ZzQs6d4t2_1;
	wire w_dff_B_ArAGjGG74_1;
	wire w_dff_B_5qfs6eGb0_1;
	wire w_dff_A_Xle9Dmgz2_1;
	wire w_dff_A_z4XKVlhK2_1;
	wire w_dff_A_jfUGE5tT0_1;
	wire w_dff_A_PFPzP88J5_1;
	wire w_dff_A_MDG70IGx8_1;
	wire w_dff_A_pRUoTZao7_1;
	wire w_dff_B_bPaiuNPW7_3;
	wire w_dff_B_JfWnVgFu5_3;
	wire w_dff_B_Y9XE2ZZg8_3;
	wire w_dff_B_KGvslmRa9_3;
	wire w_dff_B_r3Df2uqj6_3;
	wire w_dff_B_7xvuNP4j7_3;
	wire w_dff_B_5V7Qa8fd0_3;
	wire w_dff_B_OITevaWi2_3;
	wire w_dff_A_zfivgzQD7_1;
	wire w_dff_A_xpW9u7715_1;
	wire w_dff_A_OJsL894y4_1;
	wire w_dff_A_ZvFnALLa1_1;
	wire w_dff_A_uvvfuUbd9_1;
	wire w_dff_A_wuKu8Twq6_1;
	wire w_dff_A_VR0JYUqs3_1;
	wire w_dff_A_zFw44dvQ9_1;
	wire w_dff_A_9fbgEdg66_1;
	wire w_dff_A_z4qfyLAF0_1;
	wire w_dff_A_nEbG1Hc63_1;
	wire w_dff_A_TPrcG7s28_1;
	wire w_dff_A_1m2tPiys5_1;
	wire w_dff_A_QQetPoYP3_1;
	wire w_dff_A_G9UY5Wjl4_1;
	wire w_dff_A_QWdUFinA3_1;
	wire w_dff_A_44uvJDc92_1;
	wire w_dff_A_5nr9JNoN4_1;
	wire w_dff_A_YaQ6DfTj4_1;
	wire w_dff_A_8FFtGJvN1_1;
	wire w_dff_A_1b21DjhC1_2;
	wire w_dff_A_PJg3mHst9_2;
	wire w_dff_A_MuqMFDeA2_2;
	wire w_dff_A_l7hXzU142_2;
	wire w_dff_A_ztQ9x2QQ4_2;
	wire w_dff_A_YoXKZITh4_2;
	wire w_dff_A_UNHbRGcD2_2;
	wire w_dff_A_T6GTcP1f5_2;
	wire w_dff_A_8a8iIFTM4_1;
	wire w_dff_A_FfVdTNP35_1;
	wire w_dff_A_F8EUEhhI8_1;
	wire w_dff_A_KyteEw716_1;
	wire w_dff_A_UKS2OG6w5_0;
	wire w_dff_A_IvZc5PzL8_0;
	wire w_dff_A_uVzCD2xt2_0;
	wire w_dff_A_RHud1xLO8_0;
	wire w_dff_A_pCLLzebd9_0;
	wire w_dff_A_dUBtC1qd6_0;
	wire w_dff_A_4kgXKw3Q4_0;
	wire w_dff_A_8nxSezyE0_0;
	wire w_dff_A_bdxg8klS9_0;
	wire w_dff_A_Dtk9iih96_0;
	wire w_dff_A_xnniHpW95_0;
	wire w_dff_A_3jlUaKb16_0;
	wire w_dff_A_qldccWpz1_0;
	wire w_dff_A_va40lpK76_0;
	wire w_dff_A_paX5FpD35_2;
	wire w_dff_A_83v3Ptnb2_2;
	wire w_dff_A_066jas2T6_2;
	wire w_dff_A_INSPVGEJ9_2;
	wire w_dff_A_hT3JGetU5_1;
	wire w_dff_A_oUvkHlAV4_1;
	wire w_dff_A_GFdWze8v3_1;
	wire w_dff_A_q9ZKECyl4_1;
	wire w_dff_A_vkKBmERZ0_1;
	wire w_dff_A_x0CfwG637_1;
	wire w_dff_A_mGyWlh4m6_1;
	wire w_dff_A_J9YVKSMT2_1;
	wire w_dff_A_TE1LYzJ55_1;
	wire w_dff_A_NROoXcQx5_1;
	wire w_dff_A_8SHpV8Nt2_1;
	wire w_dff_A_Nh81YyjX3_1;
	wire w_dff_A_sUwDPp9l2_1;
	wire w_dff_A_GhiR5F3t9_2;
	wire w_dff_A_MFHuu97o5_2;
	wire w_dff_A_0EOctvqZ9_2;
	wire w_dff_A_306pFsMo8_2;
	wire w_dff_A_Ak6kEMNY0_2;
	wire w_dff_A_I3HcGDLJ5_2;
	wire w_dff_A_0DpHexeU4_2;
	wire w_dff_A_Ht5CjNyr0_2;
	wire w_dff_A_zAfpDSX87_1;
	wire w_dff_A_cOcRJlFR6_1;
	wire w_dff_A_o6lfSWg87_1;
	wire w_dff_A_voUozTFw6_1;
	wire w_dff_A_rsFIe1aH5_1;
	wire w_dff_A_p9nyq2QR8_1;
	wire w_dff_A_itxIFKPu8_1;
	wire w_dff_B_D0vffpct1_2;
	wire w_dff_B_mIIJ43376_2;
	wire w_dff_B_yyJouFsP9_2;
	wire w_dff_B_y1SzNhuL3_2;
	wire w_dff_A_RNBdg8Ms9_1;
	wire w_dff_A_rClJEoJn2_1;
	wire w_dff_A_NgCqrEpS2_1;
	wire w_dff_A_JNhs96JO1_1;
	wire w_dff_A_xn0pxsVC0_1;
	wire w_dff_A_6ylewrAP0_1;
	wire w_dff_A_exW2EZWI8_0;
	wire w_dff_A_L2KCFRc49_0;
	wire w_dff_A_ju2QhJQJ5_0;
	wire w_dff_A_RATGlef17_0;
	wire w_dff_A_sV33Isf88_0;
	wire w_dff_A_wC9MZx0i8_0;
	wire w_dff_A_20GTuGzz7_0;
	wire w_dff_A_bb2z6G8Z2_0;
	wire w_dff_A_P1CXzswa6_2;
	wire w_dff_A_yJ1wKhIb6_2;
	wire w_dff_A_fSYQQfb87_2;
	wire w_dff_A_zjT6Xz1q5_2;
	wire w_dff_A_im0Atm1c4_0;
	wire w_dff_A_XaOxr14T7_0;
	wire w_dff_A_lusLN7lH4_0;
	wire w_dff_A_ljsR9KFd9_0;
	wire w_dff_A_NLs4hC7u2_0;
	wire w_dff_A_n6gYM2im1_0;
	wire w_dff_B_9uarQ1Is4_1;
	wire w_dff_B_3qBlOM3f6_1;
	wire w_dff_B_nU0ZGq4l6_1;
	wire w_dff_B_d9HnqHjg6_1;
	wire w_dff_B_Sea4Laxb4_1;
	wire w_dff_B_HDMLwBiH1_1;
	wire w_dff_B_WSpepJWM5_1;
	wire w_dff_B_7c8zefUi4_1;
	wire w_dff_A_1276Se0U6_1;
	wire w_dff_A_UvhdSvIW7_1;
	wire w_dff_A_A0sc5vW81_1;
	wire w_dff_A_N6wcWuk02_1;
	wire w_dff_A_qOyCYc875_1;
	wire w_dff_A_eN5PGpMF1_1;
	wire w_dff_A_0C0f06Tg1_1;
	wire w_dff_A_dVLCxt2u1_1;
	wire w_dff_A_WTQitkku9_0;
	wire w_dff_A_KZy4AgKK7_0;
	wire w_dff_A_RGUelmQ76_0;
	wire w_dff_A_9XrtnsfL1_1;
	wire w_dff_B_PbmYmigO7_2;
	wire w_dff_B_LN0jDN862_2;
	wire w_dff_B_NQ3Az6R77_2;
	wire w_dff_B_W2ds2gT87_2;
	wire w_dff_A_KX4xrdus9_2;
	wire w_dff_A_cZ6N61VB0_2;
	wire w_dff_A_9klrine08_1;
	wire w_dff_A_BzAvCowr5_1;
	wire w_dff_A_1dS8OmZd0_1;
	wire w_dff_A_7XkwRaaW3_1;
	wire w_dff_A_cTxiTtCl2_1;
	wire w_dff_A_lv8FHbdM0_1;
	wire w_dff_A_OlVTpwZU4_2;
	wire w_dff_A_gDVyWr702_2;
	wire w_dff_A_buhkmTua3_2;
	wire w_dff_A_k9kVHTqQ3_2;
	wire w_dff_A_u7tzo7zk0_2;
	wire w_dff_A_ah55yj4e8_2;
	wire w_dff_A_8bgxasnh3_2;
	wire w_dff_A_siOi6SOO6_2;
	wire w_dff_A_HNYOv0cD4_0;
	wire w_dff_A_Lm7BwhMC1_0;
	wire w_dff_A_6n5evL4g2_0;
	wire w_dff_A_sR5Q5RPH8_0;
	wire w_dff_A_qLueEBvD8_0;
	wire w_dff_A_eAF7bSiM8_0;
	wire w_dff_A_5A1BFLOD0_0;
	wire w_dff_B_lnS2vrXY0_1;
	wire w_dff_B_JrDdZA3y2_1;
	wire w_dff_B_pDCYbpM12_1;
	wire w_dff_B_Dc7TnKSD0_1;
	wire w_dff_B_7aBGlWGu1_1;
	wire w_dff_B_cTxHss4A7_1;
	wire w_dff_B_U7cJsRJT2_1;
	wire w_dff_B_axxf9eNX1_1;
	wire w_dff_B_8sAH4KSb6_1;
	wire w_dff_A_6l4WfGqp4_2;
	wire w_dff_A_oGHeM9ZH6_2;
	wire w_dff_A_lMEn3ARL2_2;
	wire w_dff_A_Sl90eJT38_2;
	wire w_dff_A_sGm1VWF71_2;
	wire w_dff_A_8htcuhXY7_2;
	wire w_dff_A_y9Y7Sc8U7_2;
	wire w_dff_A_tvP2TVC82_2;
	wire w_dff_A_46IsRfaU5_2;
	wire w_dff_B_8lj84eFO9_0;
	wire w_dff_B_RqulqVkV4_0;
	wire w_dff_B_NkXKTgrX3_0;
	wire w_dff_B_BUhoOciU0_0;
	wire w_dff_B_8l7w3nKv2_0;
	wire w_dff_A_HJxgksb40_0;
	wire w_dff_A_OfQHsrTF6_0;
	wire w_dff_A_RHKRwJjA2_0;
	wire w_dff_A_8gyjgMM89_0;
	wire w_dff_A_2EFgIYXW6_2;
	wire w_dff_A_enq2Zzxs7_2;
	wire w_dff_A_9o9dBuND3_2;
	wire w_dff_A_fSnEzeN89_2;
	wire w_dff_A_mxXocBMM9_2;
	wire w_dff_A_L62tc7Dd0_0;
	wire w_dff_A_a4qT7Xu44_0;
	wire w_dff_A_1xzprc0w0_0;
	wire w_dff_A_L6VAPfac5_0;
	wire w_dff_A_klsIOVKv9_0;
	wire w_dff_A_V3oXX5jK6_0;
	wire w_dff_A_8VgGHXUs0_1;
	wire w_dff_A_GbhNhxNH8_1;
	wire w_dff_A_PisMM5Bj4_1;
	wire w_dff_A_TqH7orVF0_1;
	wire w_dff_A_Oz6QmTxr1_1;
	wire w_dff_A_TdVLNlCS0_1;
	wire w_dff_A_rvSm0j1y6_1;
	wire w_dff_A_AkP1uF6n0_1;
	wire w_dff_A_Rxs8MonY8_1;
	wire w_dff_A_Vt5OnxID0_1;
	wire w_dff_A_ILWbdHPl1_1;
	wire w_dff_A_JBxxJOJA1_1;
	wire w_dff_A_da8ugNZc1_1;
	wire w_dff_A_qoIWz5a47_2;
	wire w_dff_A_q3X0KEwW9_2;
	wire w_dff_A_730LaZ7j1_2;
	wire w_dff_A_eY3Mqnvi9_2;
	wire w_dff_A_noMmOXyy1_2;
	wire w_dff_A_QCiMM3Yr2_2;
	wire w_dff_A_xY7Von7i7_2;
	wire w_dff_A_Twmi2ZNt9_2;
	wire w_dff_A_Mc204LWe0_2;
	wire w_dff_B_fPSD0pYd9_1;
	wire w_dff_B_DTU96SJW7_0;
	wire w_dff_B_uepjOYpG2_0;
	wire w_dff_A_ALhd4WmP7_0;
	wire w_dff_A_UZ8gk4Pj5_0;
	wire w_dff_A_MYSTLQrl9_0;
	wire w_dff_A_KImW2BEJ3_0;
	wire w_dff_A_XdXQYG6W9_0;
	wire w_dff_A_ZzO4hFMM8_0;
	wire w_dff_A_aY5nKX752_0;
	wire w_dff_A_fLHp83Dq1_0;
	wire w_dff_A_950OsaRw7_2;
	wire w_dff_A_GC1gLHOV3_2;
	wire w_dff_A_sSuLM3c61_2;
	wire w_dff_A_39Baepz57_2;
	wire w_dff_A_wyp1YpKB4_2;
	wire w_dff_A_BXFiDA3H5_2;
	wire w_dff_A_NRrZTE351_2;
	wire w_dff_B_Fdz3JHdN9_3;
	wire w_dff_B_zw2JVQPw8_0;
	wire w_dff_B_wGz6DyCH2_0;
	wire w_dff_B_4cD81alE6_0;
	wire w_dff_B_QNW1eCAA6_0;
	wire w_dff_B_NUzTcCaO1_0;
	wire w_dff_B_92g3k8ZW4_0;
	wire w_dff_B_YR8dbmug6_0;
	wire w_dff_B_xP34Jod42_0;
	wire w_dff_B_KDbK71tq5_0;
	wire w_dff_B_76toLV5I0_0;
	wire w_dff_A_SriR0mtm0_1;
	wire w_dff_A_9tXpX3St5_1;
	wire w_dff_A_twc62EEK4_1;
	wire w_dff_A_NKLBGq8R1_1;
	wire w_dff_A_GJnujMiz2_1;
	wire w_dff_A_J5WWu8vw3_1;
	wire w_dff_A_XseHY1Bc0_0;
	wire w_dff_A_GV7MT6a02_0;
	wire w_dff_A_V3Qm89lt7_0;
	wire w_dff_A_Nx2WuXS21_0;
	wire w_dff_A_4hjn560R5_0;
	wire w_dff_A_h00G7oYg4_0;
	wire w_dff_A_34xTxBlh3_0;
	wire w_dff_A_m56LLBKI0_0;
	wire w_dff_A_kpnReuMh1_0;
	wire w_dff_A_ZnRoYSm69_0;
	wire w_dff_A_OzA84GwL3_0;
	wire w_dff_B_9l6yyhOS4_3;
	wire w_dff_B_A4JFNNgI4_3;
	wire w_dff_B_PZsI1MeH8_3;
	wire w_dff_B_tWTJ7AHu0_3;
	wire w_dff_B_4mQzefYm8_3;
	wire w_dff_B_MOzoEuXH0_3;
	wire w_dff_B_xKtEAKwg1_3;
	wire w_dff_B_4LaYW1xw5_3;
	wire w_dff_B_KbHsGt928_3;
	wire w_dff_B_9o2qWziS6_0;
	wire w_dff_B_tiTsG5Uz1_0;
	wire w_dff_B_FomnhM4z3_0;
	wire w_dff_B_NpP7XHZp8_0;
	wire w_dff_B_y0VubNw90_0;
	wire w_dff_A_sKjzEtp54_1;
	wire w_dff_B_7XqWas4T8_2;
	wire w_dff_B_5uZwh7n95_2;
	wire w_dff_B_bdNmndIN0_2;
	wire w_dff_B_1vyeyFvv6_2;
	wire w_dff_A_oSWM9JoE8_0;
	wire w_dff_B_v1kqLZzI0_1;
	wire w_dff_B_5rUP3GbJ8_1;
	wire w_dff_A_N45xjSrR7_0;
	wire w_dff_A_wcdBy92T7_0;
	wire w_dff_B_UjZgYGR24_2;
	wire w_dff_A_cpCu6avO1_0;
	wire w_dff_A_NSZkdbwm2_0;
	wire w_dff_A_0oyhkhfG6_1;
	wire w_dff_A_mXyGRX4a1_0;
	wire w_dff_A_9AvQxqe39_0;
	wire w_dff_A_RCCusdtM6_0;
	wire w_dff_A_n4EJj6SZ6_0;
	wire w_dff_A_Tu6IBioy6_2;
	wire w_dff_A_xdF2g7xZ1_2;
	wire w_dff_A_lvPQA1Dz7_2;
	wire w_dff_A_yTbhX3DK6_2;
	wire w_dff_A_CmXasMQG4_1;
	wire w_dff_A_gX0bUCa55_1;
	wire w_dff_A_3gMeFb358_1;
	wire w_dff_A_ktBrAn0o7_1;
	wire w_dff_A_04GdtLtn4_1;
	wire w_dff_A_XWhEy3fA5_1;
	wire w_dff_A_xWOPtsL63_1;
	wire w_dff_A_jwd2PVLX6_1;
	wire w_dff_A_tWGjU2hY2_2;
	wire w_dff_A_drFSEFik4_2;
	wire w_dff_A_WeDFvyBK6_2;
	wire w_dff_A_vtFqyFjw7_1;
	wire w_dff_A_BRHNwvHb2_0;
	wire w_dff_A_OYyvent54_0;
	wire w_dff_A_l1lgeYc16_2;
	wire w_dff_A_96QlWdhU9_0;
	wire w_dff_A_vSZJR51x1_0;
	wire w_dff_A_obUGa6ao4_0;
	wire w_dff_A_34mUYBoW0_0;
	wire w_dff_A_Fbey7Ie68_0;
	wire w_dff_A_dPDWhqCa3_0;
	wire w_dff_A_nOjcjacW6_0;
	wire w_dff_A_3IrxBpCR3_0;
	wire w_dff_A_0P3NhH3m6_0;
	wire w_dff_A_wflFVMgs8_1;
	wire w_dff_A_H3WSC5Cr7_1;
	wire w_dff_A_SzktELqp8_1;
	wire w_dff_B_rIwknfaB5_2;
	wire w_dff_B_RErpIhdZ2_2;
	wire w_dff_B_lmnB0qBT2_2;
	wire w_dff_B_GpVk69285_2;
	wire w_dff_A_r2bFMfYK2_0;
	wire w_dff_A_L1iI4IxQ0_0;
	wire w_dff_A_dT8BkolX6_0;
	wire w_dff_A_GaCu5nFp5_0;
	wire w_dff_A_htwfXtvx6_0;
	wire w_dff_A_lq4FohJn7_0;
	wire w_dff_A_hbdbuWOr4_0;
	wire w_dff_A_7yRMoRsM6_0;
	wire w_dff_A_J5vPYbcI0_0;
	wire w_dff_A_laDFa2zu2_2;
	wire w_dff_A_9OPS5w880_2;
	wire w_dff_A_LLc8bT972_2;
	wire w_dff_A_b1ljgJmY3_2;
	wire w_dff_A_nNpQaDzM0_2;
	wire w_dff_A_dB3LscY20_2;
	wire w_dff_A_xHp1pKxb1_2;
	wire w_dff_A_SjoOAylz5_2;
	wire w_dff_A_PL2qUMNt7_2;
	wire w_dff_A_MfkAFl0a6_0;
	wire w_dff_A_Odny8Msv7_0;
	wire w_dff_A_piYXRAxf0_0;
	wire w_dff_A_XtQmeaet3_0;
	wire w_dff_A_rdNs4Fft0_0;
	wire w_dff_A_lkCyxoMw0_0;
	wire w_dff_B_b8ZWjFh27_0;
	wire w_dff_A_hDQvtrfi8_1;
	wire w_dff_A_quODDAjE7_1;
	wire w_dff_A_QmySZphF4_1;
	wire w_dff_A_LroE6Vnx5_1;
	wire w_dff_A_o9pMM5bp2_1;
	wire w_dff_A_qojV7tH43_1;
	wire w_dff_A_8qlIpxDT9_1;
	wire w_dff_A_NdxYmoco0_1;
	wire w_dff_A_WqJex0pj3_2;
	wire w_dff_A_cO8ebXUQ9_1;
	wire w_dff_A_wIKXo2rm0_1;
	wire w_dff_A_bXzyRzKZ0_1;
	wire w_dff_A_fRIkdtgf0_1;
	wire w_dff_A_zMhrg1dP1_1;
	wire w_dff_A_4UdvMskC3_1;
	wire w_dff_A_xMdlOa8c6_0;
	wire w_dff_A_3GW2ZMyL9_1;
	wire w_dff_A_xlfd0ulf6_1;
	wire w_dff_B_NANhh2Uw2_3;
	wire w_dff_B_Xcmk5ta43_3;
	wire w_dff_A_kPrmW1xA7_1;
	wire w_dff_A_QaRVHLuf2_1;
	wire w_dff_A_WL3akhXN1_1;
	wire w_dff_A_Jw0iRXoy0_1;
	wire w_dff_A_6mUDeEdE6_1;
	wire w_dff_A_FfLDhcoP8_1;
	wire w_dff_A_zuYUgyF44_1;
	wire w_dff_A_wVTUoFv55_1;
	wire w_dff_A_mBVIAkts0_1;
	wire w_dff_A_CYnoMac51_2;
	wire w_dff_A_fTM6ixcC6_2;
	wire w_dff_A_WYgSgO6b6_2;
	wire w_dff_A_pxeYE0363_2;
	wire w_dff_A_VdK6Yi0k4_2;
	wire w_dff_A_6qrrPZvc4_2;
	wire w_dff_A_LrqkyobM3_2;
	wire w_dff_A_yJXLWBp65_2;
	wire w_dff_A_wLEibnnH4_2;
	wire w_dff_A_EUmFp00M3_2;
	wire w_dff_A_5SJuxCkp4_2;
	wire w_dff_A_HSjTpPa27_2;
	wire w_dff_A_idGuKr9w1_0;
	wire w_dff_A_vg55lHw58_0;
	wire w_dff_A_rzYNMmVB3_0;
	wire w_dff_A_PRplB95s9_0;
	wire w_dff_A_7aX1TLdR2_0;
	wire w_dff_A_sK38tr9E7_0;
	wire w_dff_A_WyhyoSTf0_0;
	wire w_dff_A_DwZrHQHc2_0;
	wire w_dff_A_mXbgThea2_0;
	wire w_dff_A_r0TA22Mu1_0;
	wire w_dff_A_NFRYoIXw7_0;
	wire w_dff_A_TbKnCqjP0_0;
	wire w_dff_A_Gol52KhP8_0;
	wire w_dff_A_OzaMz4Ag7_0;
	wire w_dff_A_3EHQgUGu1_0;
	wire w_dff_A_NUZ2tYBl2_0;
	wire w_dff_A_Ce8vzDI03_0;
	wire w_dff_A_tioiS3R20_0;
	wire w_dff_A_86xQDTQk2_0;
	wire w_dff_A_zZ4yhI6G8_0;
	wire w_dff_A_5s27TObq3_0;
	wire w_dff_A_Xp999MZh7_0;
	wire w_dff_A_cH18MPb36_0;
	wire w_dff_A_SGf4mYTT3_0;
	wire w_dff_A_Z0eio7q67_0;
	wire w_dff_A_f9jfGi1f8_2;
	wire w_dff_A_HMwz0DNp8_0;
	wire w_dff_A_HV3zwfae1_0;
	wire w_dff_A_D6Sv39Nd2_0;
	wire w_dff_A_LMREqGFh0_0;
	wire w_dff_A_ca35UtDb1_0;
	wire w_dff_A_fd6Tv5PF4_0;
	wire w_dff_A_HWwoIRTV6_0;
	wire w_dff_A_L1MFaNGw5_0;
	wire w_dff_A_gFWabiwQ6_0;
	wire w_dff_A_cSwBo1S84_0;
	wire w_dff_A_296taM8l5_0;
	wire w_dff_A_jYimi9zI3_0;
	wire w_dff_A_B2ceTytw6_0;
	wire w_dff_A_uzxHMbEa7_0;
	wire w_dff_A_RVlSOjWJ5_0;
	wire w_dff_A_p8j1fZJX5_0;
	wire w_dff_A_p3UBz73t9_0;
	wire w_dff_A_Dq2CU8ir5_0;
	wire w_dff_A_uNVvBkCR0_0;
	wire w_dff_A_q3j452TK6_0;
	wire w_dff_A_FbW9FTP21_0;
	wire w_dff_A_b36pVjRq4_0;
	wire w_dff_A_oECxZpiS8_0;
	wire w_dff_A_6w8racrw7_0;
	wire w_dff_A_4BaqbvN94_0;
	wire w_dff_A_xEjasLss1_2;
	wire w_dff_A_S4BSjuEv6_0;
	wire w_dff_A_u0TSUPbc6_0;
	wire w_dff_A_AE9M0Kb65_0;
	wire w_dff_A_h3Pgjv6l0_0;
	wire w_dff_A_obBNlIvk1_0;
	wire w_dff_A_WbJC8jyf2_0;
	wire w_dff_A_0JLLsif19_0;
	wire w_dff_A_iLzIIg2s4_0;
	wire w_dff_A_HXdi2wXa4_0;
	wire w_dff_A_qud9klAs1_0;
	wire w_dff_A_vryFEqRx4_0;
	wire w_dff_A_Ac9i4vmv3_0;
	wire w_dff_A_60t3tQxw1_0;
	wire w_dff_A_daHJC0Hc7_0;
	wire w_dff_A_3SGc56OH4_0;
	wire w_dff_A_daKrQNTC3_0;
	wire w_dff_A_KnwKOTlc6_0;
	wire w_dff_A_ytdODurQ0_0;
	wire w_dff_A_ivYdgyuy5_0;
	wire w_dff_A_PbTYPrLf1_0;
	wire w_dff_A_u0x9AqAx3_0;
	wire w_dff_A_4lOJXUlQ6_0;
	wire w_dff_A_0gIa4O151_0;
	wire w_dff_A_wNt5qoBd0_0;
	wire w_dff_A_o0SInsMd8_0;
	wire w_dff_A_Cbt2rFAg8_2;
	wire w_dff_A_1MyEp29m8_0;
	wire w_dff_A_XvKS7zT87_0;
	wire w_dff_A_YlJyR9GJ6_0;
	wire w_dff_A_a0weg2kE5_0;
	wire w_dff_A_TQM7qa7r1_0;
	wire w_dff_A_S9G4N98N7_0;
	wire w_dff_A_cqp1KyIn0_0;
	wire w_dff_A_NhjFSoQ59_0;
	wire w_dff_A_1jGBqCSY7_0;
	wire w_dff_A_BCeEtFbI2_0;
	wire w_dff_A_D80TTEYH3_0;
	wire w_dff_A_l9kjwhD18_0;
	wire w_dff_A_r1HOiBy80_0;
	wire w_dff_A_WrP7NWcZ3_0;
	wire w_dff_A_SObQLSJS2_0;
	wire w_dff_A_trccRMOl7_0;
	wire w_dff_A_eFKgkVmo2_0;
	wire w_dff_A_vOK49FMM8_0;
	wire w_dff_A_cByvQm4W0_0;
	wire w_dff_A_zXxNE0wq8_0;
	wire w_dff_A_2CNvd6hu5_0;
	wire w_dff_A_gUL5Fqwn9_0;
	wire w_dff_A_8hs3jjnI3_0;
	wire w_dff_A_aFRDWzMY2_0;
	wire w_dff_A_VTodtSkO6_0;
	wire w_dff_A_h4I0Sdyv3_0;
	wire w_dff_A_JJMPLPol7_2;
	wire w_dff_A_zxJ2Df549_0;
	wire w_dff_A_yBRMDJhx8_0;
	wire w_dff_A_kwigkLOH3_0;
	wire w_dff_A_MCQAO53A7_0;
	wire w_dff_A_iBEuXitr9_0;
	wire w_dff_A_4bafrp5H0_0;
	wire w_dff_A_dcKDPXzk9_0;
	wire w_dff_A_jrUf9jZz0_0;
	wire w_dff_A_ChxVa4a04_0;
	wire w_dff_A_A3bHpQhj3_0;
	wire w_dff_A_XsRhZxzX1_0;
	wire w_dff_A_jB7Si0fg3_0;
	wire w_dff_A_z8h3eS3X4_0;
	wire w_dff_A_BIEDadFO7_0;
	wire w_dff_A_Jv4vFuU77_0;
	wire w_dff_A_VBju6Dg06_0;
	wire w_dff_A_Qb0xrRd38_0;
	wire w_dff_A_N3n2jcgj9_0;
	wire w_dff_A_Z1HAv0Te5_0;
	wire w_dff_A_3cQgvXZ49_0;
	wire w_dff_A_hOUyfhGo9_0;
	wire w_dff_A_s6LtyaQZ9_0;
	wire w_dff_A_vWmPcjBe7_0;
	wire w_dff_A_jV1i1rqS4_0;
	wire w_dff_A_a7ON3QTw2_2;
	wire w_dff_A_DTgA1dQF9_0;
	wire w_dff_A_Xcmqkp3J5_0;
	wire w_dff_A_Cm5WgIml4_0;
	wire w_dff_A_0GzK5Pvj4_0;
	wire w_dff_A_JV9dQzFw4_0;
	wire w_dff_A_U389dqkI3_0;
	wire w_dff_A_dzGRMpLF4_0;
	wire w_dff_A_2xWTgVTf8_0;
	wire w_dff_A_lXs6Jn781_0;
	wire w_dff_A_imRzTusE1_0;
	wire w_dff_A_FulKy1cM0_0;
	wire w_dff_A_1JEw5cSI1_0;
	wire w_dff_A_efmcyHqd5_0;
	wire w_dff_A_A7mAtw7O5_0;
	wire w_dff_A_GEZ9vhTE6_0;
	wire w_dff_A_EYkfTLMA4_0;
	wire w_dff_A_yNFT2uKZ8_0;
	wire w_dff_A_ye6WrywS0_0;
	wire w_dff_A_I60293s53_0;
	wire w_dff_A_fP4q7mAE3_0;
	wire w_dff_A_daZmWlMT8_0;
	wire w_dff_A_TnxqdI4c1_0;
	wire w_dff_A_sGkqRViV5_2;
	wire w_dff_A_7xCTlbl73_0;
	wire w_dff_A_FbKaRzbb5_0;
	wire w_dff_A_Oq84gOft3_0;
	wire w_dff_A_PpDO167k2_0;
	wire w_dff_A_Y455jQ0n4_0;
	wire w_dff_A_TtXrNHfD9_0;
	wire w_dff_A_KvGDVl7u2_0;
	wire w_dff_A_1cXROs9R2_0;
	wire w_dff_A_7q2YFTi09_0;
	wire w_dff_A_tBKDfHWq7_0;
	wire w_dff_A_U5wuA1fv2_0;
	wire w_dff_A_5ND1oFoY5_0;
	wire w_dff_A_LA91jVVJ0_0;
	wire w_dff_A_j5En6ecb7_0;
	wire w_dff_A_JC8OGn1F0_0;
	wire w_dff_A_tPYt13Bd3_0;
	wire w_dff_A_UCbCiM7p0_0;
	wire w_dff_A_3aksizyi0_0;
	wire w_dff_A_Nw4UEA4k9_0;
	wire w_dff_A_18YPC1vo5_0;
	wire w_dff_A_km4XTKFV5_0;
	wire w_dff_A_hQAagMdR9_0;
	wire w_dff_A_pFwlOgAu4_0;
	wire w_dff_A_Yz1levAm9_0;
	wire w_dff_A_BHZ57keO2_2;
	wire w_dff_A_taGKzJPg3_0;
	wire w_dff_A_EbK3gKnN3_0;
	wire w_dff_A_fzw0d7ND8_0;
	wire w_dff_A_Y6kPJhE06_0;
	wire w_dff_A_qxPrS9xV0_0;
	wire w_dff_A_Eaj43ibm4_0;
	wire w_dff_A_JYvudEBN0_0;
	wire w_dff_A_whqszE3R1_0;
	wire w_dff_A_xU6hoIzQ9_0;
	wire w_dff_A_ntLWWh2T0_0;
	wire w_dff_A_k5sL1d9Y5_0;
	wire w_dff_A_Gjl8uLap7_0;
	wire w_dff_A_hGpaFSkD3_0;
	wire w_dff_A_VTGlvQ4I5_0;
	wire w_dff_A_QihP0Aci1_0;
	wire w_dff_A_cX9qwrjL3_0;
	wire w_dff_A_V7dbeJo28_0;
	wire w_dff_A_PDG6DZXt0_0;
	wire w_dff_A_anMJzwjP0_0;
	wire w_dff_A_esdq5fg16_0;
	wire w_dff_A_oc3xFxVt5_0;
	wire w_dff_A_HcZgitik1_0;
	wire w_dff_A_eYRAqSb62_0;
	wire w_dff_A_jTIiErZg3_0;
	wire w_dff_A_NliuMYGZ6_2;
	wire w_dff_A_CFniME9j9_0;
	wire w_dff_A_McNRy9Yo9_0;
	wire w_dff_A_cGZP2Qm32_0;
	wire w_dff_A_FQgyl4FQ6_0;
	wire w_dff_A_Y0mWhTRw7_0;
	wire w_dff_A_jJunn7vf3_0;
	wire w_dff_A_hk2NxoL14_0;
	wire w_dff_A_8soCHyqz9_0;
	wire w_dff_A_zkWQI8Kg0_0;
	wire w_dff_A_v1ffeCSe4_0;
	wire w_dff_A_pFTUNJCc4_0;
	wire w_dff_A_qedkkuD08_0;
	wire w_dff_A_StBpS3jA8_0;
	wire w_dff_A_nptZEgg33_0;
	wire w_dff_A_6i0osKXe2_0;
	wire w_dff_A_PTevI6bL9_0;
	wire w_dff_A_j8esl1S99_0;
	wire w_dff_A_psNGMqjG3_0;
	wire w_dff_A_XewaMgJw4_0;
	wire w_dff_A_ENaEuGdi8_0;
	wire w_dff_A_XcLFnf3w2_0;
	wire w_dff_A_WM3so4VJ7_0;
	wire w_dff_A_4xocwfny9_0;
	wire w_dff_A_85WkFkzR8_0;
	wire w_dff_A_iuAfvJlo7_2;
	wire w_dff_A_7zyp774y3_0;
	wire w_dff_A_o0QDc4Lj0_0;
	wire w_dff_A_Z9xshVnD3_0;
	wire w_dff_A_2U4ebGGE2_0;
	wire w_dff_A_JpcVDTG93_0;
	wire w_dff_A_dED0aKgU3_0;
	wire w_dff_A_fFck0DHD1_0;
	wire w_dff_A_j6hya3RE5_0;
	wire w_dff_A_8uijJj7v2_0;
	wire w_dff_A_cKWoBNME2_0;
	wire w_dff_A_fVRFjDS67_0;
	wire w_dff_A_dfitOVYm9_0;
	wire w_dff_A_FpDDf8581_0;
	wire w_dff_A_xEveGCUn3_0;
	wire w_dff_A_EN62yg8U2_0;
	wire w_dff_A_j90Emxzm1_0;
	wire w_dff_A_9wadJcyZ9_0;
	wire w_dff_A_EemJd0qx1_0;
	wire w_dff_A_wMVKlU2i0_0;
	wire w_dff_A_mG2gUNQ59_0;
	wire w_dff_A_YASmzfXQ1_0;
	wire w_dff_A_V5VILOyP8_0;
	wire w_dff_A_e5W7SCNd9_0;
	wire w_dff_A_IlmZkdRu3_0;
	wire w_dff_A_pJD6yBb64_0;
	wire w_dff_A_L5QySJRo8_2;
	wire w_dff_A_F2qGzpBA7_0;
	wire w_dff_A_TQ2wNTcd7_0;
	wire w_dff_A_nzGkn6xV0_0;
	wire w_dff_A_6xVT5N4Z7_0;
	wire w_dff_A_7vDB6KNm7_0;
	wire w_dff_A_1MQN4qje1_0;
	wire w_dff_A_JYPV7wm15_0;
	wire w_dff_A_2GsegVcI0_0;
	wire w_dff_A_YzrW7Ovp0_0;
	wire w_dff_A_gjnV77zI2_0;
	wire w_dff_A_PNNuSGOK1_0;
	wire w_dff_A_3bqyUTnF6_0;
	wire w_dff_A_9evnXDIv3_0;
	wire w_dff_A_xtU66SQn3_0;
	wire w_dff_A_JFyU1dCK7_0;
	wire w_dff_A_aQADH9PS5_0;
	wire w_dff_A_7seewoh85_0;
	wire w_dff_A_CBENJXHJ6_0;
	wire w_dff_A_HO9PsLxw8_0;
	wire w_dff_A_xFSUe6E94_0;
	wire w_dff_A_lC6Hynj40_0;
	wire w_dff_A_uRT7JYxG0_0;
	wire w_dff_A_gk8fR03i2_1;
	wire w_dff_A_e47X5IZU5_0;
	wire w_dff_A_EfVOVywg4_0;
	wire w_dff_A_qcV3iOse3_0;
	wire w_dff_A_okgCl0jt8_0;
	wire w_dff_A_PK7eK3ZX3_0;
	wire w_dff_A_FCstpzfG0_0;
	wire w_dff_A_zNiaWqLi7_0;
	wire w_dff_A_16Ca2n3i1_0;
	wire w_dff_A_wstXoahf6_0;
	wire w_dff_A_tG95oNRl6_0;
	wire w_dff_A_uI4KyswJ8_0;
	wire w_dff_A_DelgB37r1_0;
	wire w_dff_A_sqY7QrJQ1_0;
	wire w_dff_A_wdhRcQGc3_0;
	wire w_dff_A_skfRXWvu2_0;
	wire w_dff_A_ODTZmUmu6_0;
	wire w_dff_A_JWibhQgc3_0;
	wire w_dff_A_F4Zc1xLN0_0;
	wire w_dff_A_IUnrGZDz2_0;
	wire w_dff_A_uBXI9UD37_0;
	wire w_dff_A_yuZRqyvC1_0;
	wire w_dff_A_g2M7lntS1_0;
	wire w_dff_A_44p5UJvB5_0;
	wire w_dff_A_pdQtL1Zb0_0;
	wire w_dff_A_JPt2ryYJ4_0;
	wire w_dff_A_z8F8E7fH6_2;
	wire w_dff_A_N6tYl2Vm4_0;
	wire w_dff_A_itiq37yH1_0;
	wire w_dff_A_EklhlN0Z8_0;
	wire w_dff_A_yliVfoSD3_0;
	wire w_dff_A_3a6PNsEi4_0;
	wire w_dff_A_tYRR5tEV3_0;
	wire w_dff_A_cDdU84Np2_0;
	wire w_dff_A_iuFlyMMf6_0;
	wire w_dff_A_T3FUjRtb4_0;
	wire w_dff_A_PCnx4Ua85_0;
	wire w_dff_A_PihY6KjF4_0;
	wire w_dff_A_YT5GUfvM0_0;
	wire w_dff_A_qoEQlI4f8_0;
	wire w_dff_A_abDVmSIk8_0;
	wire w_dff_A_FtgM57jl7_0;
	wire w_dff_A_vz1tj4NN9_0;
	wire w_dff_A_G2Bulu845_0;
	wire w_dff_A_1Vq4zG4Y3_0;
	wire w_dff_A_H57ICmdt0_0;
	wire w_dff_A_qWBwVJn27_0;
	wire w_dff_A_ySES4hWu9_0;
	wire w_dff_A_du7yM5w39_0;
	wire w_dff_A_35UzA5Ss9_2;
	wire w_dff_A_0Ptgjekn0_0;
	wire w_dff_A_j8Ii4hMS8_0;
	wire w_dff_A_lM2R0Pch0_0;
	wire w_dff_A_j84R6Ve84_0;
	wire w_dff_A_Mv0tkdQm6_0;
	wire w_dff_A_77Fev5oC7_0;
	wire w_dff_A_1b5cLdGh4_0;
	wire w_dff_A_diSnmqkp3_0;
	wire w_dff_A_q84iModq4_0;
	wire w_dff_A_AwWNJQoM4_0;
	wire w_dff_A_2uFWQlNp4_0;
	wire w_dff_A_ELE8zD7S1_0;
	wire w_dff_A_4BXwUa9W2_0;
	wire w_dff_A_shJNXAUR0_0;
	wire w_dff_A_vK0pB3BG3_0;
	wire w_dff_A_IakdHtb17_0;
	wire w_dff_A_i2CTfwHc6_0;
	wire w_dff_A_8OXctc0o6_0;
	wire w_dff_A_k0UJc8H90_0;
	wire w_dff_A_y1D5oWcT5_0;
	wire w_dff_A_YUq6vmec7_0;
	wire w_dff_A_LXlVsLMV9_0;
	wire w_dff_A_Cm3FyGve2_2;
	wire w_dff_A_31Ad5Iot4_0;
	wire w_dff_A_NfA965aN3_0;
	wire w_dff_A_G58gEOws6_0;
	wire w_dff_A_IU2e1hUv2_0;
	wire w_dff_A_KOZq2ZvW6_0;
	wire w_dff_A_joH00s858_0;
	wire w_dff_A_8lFmZ9hw9_0;
	wire w_dff_A_iRdDOUiF8_0;
	wire w_dff_A_zuCDbIFm5_0;
	wire w_dff_A_7cCx4HiP1_0;
	wire w_dff_A_9OOROhO05_0;
	wire w_dff_A_IcCDwTRV7_0;
	wire w_dff_A_DQ4gr52g4_0;
	wire w_dff_A_XRm1YKov8_0;
	wire w_dff_A_htqpJaBP0_0;
	wire w_dff_A_ZLO8NrNs5_0;
	wire w_dff_A_xE0I3a5k5_0;
	wire w_dff_A_12k9JVQK0_0;
	wire w_dff_A_e9byq4wk7_0;
	wire w_dff_A_1dRJWU1m6_0;
	wire w_dff_A_tmHVEUtT4_0;
	wire w_dff_A_6ZSNF53G6_0;
	wire w_dff_A_JkHaEiYN3_0;
	wire w_dff_A_OrUcK1n14_0;
	wire w_dff_A_yBV16ocd2_0;
	wire w_dff_A_Tfh5LF372_2;
	wire w_dff_A_uPvHRNLG3_0;
	wire w_dff_A_Uy02UmIo8_0;
	wire w_dff_A_m1Vt2YBx6_0;
	wire w_dff_A_dyAkftY82_0;
	wire w_dff_A_D53pIOFt5_0;
	wire w_dff_A_CvzpfV0D9_0;
	wire w_dff_A_ZoPtnveL5_0;
	wire w_dff_A_WPlGyvyq0_0;
	wire w_dff_A_JKOIBxQq9_0;
	wire w_dff_A_u1It9b1q6_0;
	wire w_dff_A_oRS2jfnE2_0;
	wire w_dff_A_niqioGRP2_0;
	wire w_dff_A_NSirViKM5_0;
	wire w_dff_A_YHqalQIW2_0;
	wire w_dff_A_gnDyFYLu4_0;
	wire w_dff_A_dPSSX9k19_0;
	wire w_dff_A_vIuqw2K54_0;
	wire w_dff_A_SoKFsxUJ2_0;
	wire w_dff_A_DrjcHeE33_0;
	wire w_dff_A_hopkUYEs1_0;
	wire w_dff_A_EAjv4duJ1_0;
	wire w_dff_A_zz2fzF9F7_0;
	wire w_dff_A_0wNKKP4D7_0;
	wire w_dff_A_9HXCWLs03_2;
	wire w_dff_A_Zvi0FnSB8_0;
	wire w_dff_A_MTai2li04_0;
	wire w_dff_A_ZxCGqh3S5_0;
	wire w_dff_A_KBHhX25z7_0;
	wire w_dff_A_ygILS7ks5_0;
	wire w_dff_A_mXZT9Yf57_0;
	wire w_dff_A_w9f46bQM2_0;
	wire w_dff_A_aUqLlwpE2_0;
	wire w_dff_A_RXQZh2Bh6_0;
	wire w_dff_A_FKsLlO5G5_0;
	wire w_dff_A_YFaKUnug7_0;
	wire w_dff_A_FKUAsMtU8_0;
	wire w_dff_A_dBQoEy1P7_0;
	wire w_dff_A_mshbxTQ17_0;
	wire w_dff_A_RyOrPpx31_0;
	wire w_dff_A_wGDEOBAO3_0;
	wire w_dff_A_7ZHxunlr6_0;
	wire w_dff_A_EofVAvGa0_0;
	wire w_dff_A_5ccZHtLU6_0;
	wire w_dff_A_IpKG5eOQ7_0;
	wire w_dff_A_MLPK6q7u3_0;
	wire w_dff_A_jKRHPVkF7_0;
	wire w_dff_A_baKIWzB34_0;
	wire w_dff_A_XpWbAcL04_2;
	wire w_dff_A_2Gn6GIy29_0;
	wire w_dff_A_1lALqmkr3_0;
	wire w_dff_A_8swZOnoU1_0;
	wire w_dff_A_QEaCdejI2_0;
	wire w_dff_A_yFJ7F2XZ4_0;
	wire w_dff_A_uY6qbbZk2_0;
	wire w_dff_A_YgoEzABX5_0;
	wire w_dff_A_erC9KmhN4_0;
	wire w_dff_A_zu3e41Xj6_0;
	wire w_dff_A_qz7hHSpY3_0;
	wire w_dff_A_NyZhUtfT3_0;
	wire w_dff_A_qbDNvsOO4_0;
	wire w_dff_A_4HrvKHDq8_2;
	wire w_dff_A_ZTkAA7oB6_0;
	wire w_dff_A_bbsihPsa0_0;
	wire w_dff_A_Ouqn9SIP4_0;
	wire w_dff_A_MDe9hBTy5_0;
	wire w_dff_A_FmKbmgVM8_0;
	wire w_dff_A_a3cHNdpE2_0;
	wire w_dff_A_BvwwH1tn7_0;
	wire w_dff_A_UT8qrq8w4_2;
	wire w_dff_A_Z7zdoE9J2_0;
	wire w_dff_A_GF43g0tL7_0;
	wire w_dff_A_GSg1tmyc9_0;
	wire w_dff_A_jyqkSZWD5_0;
	wire w_dff_A_NO5UTTHf5_0;
	wire w_dff_A_U0i1pmL48_0;
	wire w_dff_A_wpYFfFYg9_0;
	wire w_dff_A_xOVi91633_0;
	wire w_dff_A_xxYGU16b4_0;
	wire w_dff_A_iVhb6Mw44_2;
	wire w_dff_A_SKTtECSv5_0;
	wire w_dff_A_ztrwt2oI9_0;
	wire w_dff_A_gJ1UJKoo7_0;
	wire w_dff_A_zMBmsAcS3_0;
	wire w_dff_A_Ur4qw2Wy9_0;
	wire w_dff_A_ekL7g0Qy7_0;
	wire w_dff_A_s7lnhHck6_0;
	wire w_dff_A_QtxOKwNC8_0;
	wire w_dff_A_fFR7xMcQ5_0;
	wire w_dff_A_Z7sUUe0q7_0;
	wire w_dff_A_mDhjMDqr1_0;
	wire w_dff_A_WiHHet6v3_2;
	wire w_dff_A_XWW50pqM5_0;
	wire w_dff_A_xA640cQm0_2;
	wire w_dff_A_qV1VhWRJ7_0;
	wire w_dff_A_SJQjbrIe3_0;
	wire w_dff_A_AdgVd7bd8_0;
	wire w_dff_A_cXd4Sbxm0_0;
	wire w_dff_A_0JlrbuTL8_2;
	wire w_dff_A_esbwER353_0;
	wire w_dff_A_y8Z8qDZW3_2;
	wire w_dff_A_ZHQ0hDa74_0;
	wire w_dff_A_16jvoNja6_0;
	wire w_dff_A_vchR78ye5_0;
	jand g000(.dina(w_G75gat_0[1]),.dinb(w_G29gat_0[2]),.dout(n86),.clk(gclk));
	jand g001(.dina(w_n86_0[1]),.dinb(w_G42gat_2[1]),.dout(w_dff_A_HSjTpPa27_2),.clk(gclk));
	jand g002(.dina(w_G36gat_0[1]),.dinb(w_G29gat_0[1]),.dout(n88),.clk(gclk));
	jand g003(.dina(w_n88_0[1]),.dinb(w_G80gat_0[2]),.dout(w_dff_A_f9jfGi1f8_2),.clk(gclk));
	jand g004(.dina(w_n88_0[0]),.dinb(w_G42gat_2[0]),.dout(G390gat_fa_),.clk(gclk));
	jand g005(.dina(G86gat),.dinb(G85gat),.dout(w_dff_A_Cbt2rFAg8_2),.clk(gclk));
	jand g006(.dina(w_G8gat_0[1]),.dinb(w_G1gat_1[1]),.dout(n92),.clk(gclk));
	jand g007(.dina(w_n92_0[1]),.dinb(w_G13gat_0[1]),.dout(n93),.clk(gclk));
	jand g008(.dina(w_n93_0[1]),.dinb(w_G17gat_2[2]),.dout(w_dff_A_JJMPLPol7_2),.clk(gclk));
	jnot g009(.din(w_G17gat_2[1]),.dout(n95),.clk(gclk));
	jnot g010(.din(w_G13gat_0[0]),.dout(n96),.clk(gclk));
	jnot g011(.din(w_G1gat_1[0]),.dout(n97),.clk(gclk));
	jnot g012(.din(w_G26gat_0[1]),.dout(n98),.clk(gclk));
	jor g013(.dina(n98),.dinb(w_n97_0[1]),.dout(n99),.clk(gclk));
	jor g014(.dina(w_n99_0[1]),.dinb(w_dff_B_rCIjOu890_1),.dout(n100),.clk(gclk));
	jor g015(.dina(n100),.dinb(w_n95_0[2]),.dout(n101),.clk(gclk));
	jor g016(.dina(w_n101_0[1]),.dinb(w_G390gat_0[1]),.dout(w_dff_A_a7ON3QTw2_2),.clk(gclk));
	jnot g017(.din(w_G80gat_0[1]),.dout(n103),.clk(gclk));
	jand g018(.dina(w_G75gat_0[0]),.dinb(w_G59gat_1[1]),.dout(n104),.clk(gclk));
	jnot g019(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jor g020(.dina(n105),.dinb(w_n103_0[1]),.dout(w_dff_A_sGkqRViV5_2),.clk(gclk));
	jnot g021(.din(w_G36gat_0[0]),.dout(n107),.clk(gclk));
	jnot g022(.din(w_G59gat_1[0]),.dout(n108),.clk(gclk));
	jor g023(.dina(w_n108_0[1]),.dinb(n107),.dout(n109),.clk(gclk));
	jor g024(.dina(w_n109_0[1]),.dinb(w_n103_0[0]),.dout(w_dff_A_BHZ57keO2_2),.clk(gclk));
	jnot g025(.din(w_G42gat_1[2]),.dout(n111),.clk(gclk));
	jor g026(.dina(w_n109_0[0]),.dinb(w_n111_0[1]),.dout(w_dff_A_NliuMYGZ6_2),.clk(gclk));
	jor g027(.dina(G88gat),.dinb(G87gat),.dout(n113),.clk(gclk));
	jand g028(.dina(w_n113_0[1]),.dinb(w_dff_B_jm6eXLIy3_1),.dout(w_dff_A_iuAfvJlo7_2),.clk(gclk));
	jnot g029(.din(w_G390gat_0[0]),.dout(n115),.clk(gclk));
	jor g030(.dina(w_n101_0[0]),.dinb(w_dff_B_UsegxPG92_1),.dout(w_dff_A_L5QySJRo8_2),.clk(gclk));
	jand g031(.dina(w_G26gat_0[0]),.dinb(w_G1gat_0[2]),.dout(n117),.clk(gclk));
	jand g032(.dina(n117),.dinb(w_G51gat_1[1]),.dout(G447gat_fa_),.clk(gclk));
	jand g033(.dina(w_n93_0[0]),.dinb(w_G55gat_0[2]),.dout(n119),.clk(gclk));
	jand g034(.dina(w_n119_0[2]),.dinb(w_G29gat_0[0]),.dout(n120),.clk(gclk));
	jand g035(.dina(n120),.dinb(w_G68gat_0[1]),.dout(w_dff_A_z8F8E7fH6_2),.clk(gclk));
	jand g036(.dina(w_G68gat_0[0]),.dinb(w_G59gat_0[2]),.dout(n122),.clk(gclk));
	jand g037(.dina(w_n119_0[1]),.dinb(w_dff_B_WVTmUIe00_1),.dout(n123),.clk(gclk));
	jand g038(.dina(n123),.dinb(w_n122_0[1]),.dout(w_dff_A_35UzA5Ss9_2),.clk(gclk));
	jand g039(.dina(w_n113_0[0]),.dinb(w_dff_B_iwGeSgRi3_1),.dout(w_dff_A_Cm3FyGve2_2),.clk(gclk));
	jxor g040(.dina(w_G116gat_0[2]),.dinb(w_G111gat_0[2]),.dout(n126),.clk(gclk));
	jxor g041(.dina(n126),.dinb(w_dff_B_rPt4A9FB8_1),.dout(n127),.clk(gclk));
	jxor g042(.dina(w_G96gat_0[2]),.dinb(w_G91gat_0[2]),.dout(n128),.clk(gclk));
	jxor g043(.dina(n128),.dinb(w_G130gat_0[1]),.dout(n129),.clk(gclk));
	jxor g044(.dina(w_G106gat_0[2]),.dinb(w_G101gat_0[2]),.dout(n130),.clk(gclk));
	jxor g045(.dina(w_G126gat_0[2]),.dinb(w_G121gat_0[2]),.dout(n131),.clk(gclk));
	jxor g046(.dina(n131),.dinb(n130),.dout(n132),.clk(gclk));
	jxor g047(.dina(n132),.dinb(n129),.dout(n133),.clk(gclk));
	jxor g048(.dina(n133),.dinb(w_dff_B_Ul7hI5tG2_1),.dout(w_dff_A_Tfh5LF372_2),.clk(gclk));
	jxor g049(.dina(w_G189gat_2[1]),.dinb(w_G183gat_1[2]),.dout(n135),.clk(gclk));
	jxor g050(.dina(n135),.dinb(w_dff_B_GCcZzlST4_1),.dout(n136),.clk(gclk));
	jxor g051(.dina(w_G159gat_1[2]),.dinb(w_G130gat_0[0]),.dout(n137),.clk(gclk));
	jxor g052(.dina(n137),.dinb(w_G165gat_1[2]),.dout(n138),.clk(gclk));
	jxor g053(.dina(w_G177gat_1[2]),.dinb(w_G171gat_1[2]),.dout(n139),.clk(gclk));
	jxor g054(.dina(w_G201gat_1[1]),.dinb(w_G195gat_2[1]),.dout(n140),.clk(gclk));
	jxor g055(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g056(.dina(n141),.dinb(n138),.dout(n142),.clk(gclk));
	jxor g057(.dina(n142),.dinb(w_dff_B_7qFlguCr1_1),.dout(w_dff_A_9HXCWLs03_2),.clk(gclk));
	jnot g058(.din(w_G268gat_0[1]),.dout(n144),.clk(gclk));
	jand g059(.dina(w_G447gat_1),.dinb(w_G80gat_0[0]),.dout(n145),.clk(gclk));
	jand g060(.dina(n145),.dinb(w_n86_0[0]),.dout(n146),.clk(gclk));
	jand g061(.dina(w_n146_0[1]),.dinb(w_G55gat_0[1]),.dout(n147),.clk(gclk));
	jand g062(.dina(n147),.dinb(w_n144_0[1]),.dout(n148),.clk(gclk));
	jand g063(.dina(w_n111_0[0]),.dinb(w_n95_0[1]),.dout(n149),.clk(gclk));
	jnot g064(.din(w_n149_0[1]),.dout(n150),.clk(gclk));
	jand g065(.dina(w_G156gat_0[1]),.dinb(w_G59gat_0[1]),.dout(n151),.clk(gclk));
	jand g066(.dina(w_G42gat_1[1]),.dinb(w_G17gat_2[0]),.dout(n152),.clk(gclk));
	jnot g067(.din(w_n152_0[1]),.dout(n153),.clk(gclk));
	jand g068(.dina(n153),.dinb(w_n151_0[1]),.dout(n154),.clk(gclk));
	jand g069(.dina(n154),.dinb(w_G447gat_0[2]),.dout(n155),.clk(gclk));
	jand g070(.dina(n155),.dinb(w_dff_B_5rUP3GbJ8_1),.dout(n156),.clk(gclk));
	jnot g071(.din(w_n92_0[0]),.dout(n157),.clk(gclk));
	jand g072(.dina(w_n104_0[0]),.dinb(w_G42gat_1[0]),.dout(n158),.clk(gclk));
	jand g073(.dina(w_G51gat_1[0]),.dinb(w_G17gat_1[2]),.dout(n159),.clk(gclk));
	jnot g074(.din(n159),.dout(n160),.clk(gclk));
	jor g075(.dina(n160),.dinb(n158),.dout(n161),.clk(gclk));
	jor g076(.dina(n161),.dinb(w_dff_B_v1kqLZzI0_1),.dout(n162),.clk(gclk));
	jnot g077(.din(w_n162_0[1]),.dout(n163),.clk(gclk));
	jor g078(.dina(n163),.dinb(n156),.dout(n164),.clk(gclk));
	jand g079(.dina(w_n164_3[1]),.dinb(w_G126gat_0[1]),.dout(n165),.clk(gclk));
	jnot g080(.din(w_G156gat_0[0]),.dout(n166),.clk(gclk));
	jor g081(.dina(n166),.dinb(w_n108_0[0]),.dout(n167),.clk(gclk));
	jand g082(.dina(w_n167_0[1]),.dinb(w_G447gat_0[1]),.dout(n168),.clk(gclk));
	jand g083(.dina(w_n168_0[1]),.dinb(w_G17gat_1[1]),.dout(n169),.clk(gclk));
	jor g084(.dina(n169),.dinb(w_n97_0[0]),.dout(n170),.clk(gclk));
	jand g085(.dina(w_n170_1[1]),.dinb(w_G153gat_0[2]),.dout(n171),.clk(gclk));
	jor g086(.dina(w_dff_B_jracUH0O1_0),.dinb(n165),.dout(n172),.clk(gclk));
	jor g087(.dina(n172),.dinb(w_n148_1[2]),.dout(n173),.clk(gclk));
	jand g088(.dina(w_n173_0[1]),.dinb(w_G246gat_3[1]),.dout(n174),.clk(gclk));
	jand g089(.dina(w_n122_0[0]),.dinb(w_G42gat_0[2]),.dout(n175),.clk(gclk));
	jand g090(.dina(G73gat),.dinb(G72gat),.dout(n176),.clk(gclk));
	jand g091(.dina(w_dff_B_b8ZWjFh27_0),.dinb(n175),.dout(n177),.clk(gclk));
	jand g092(.dina(n177),.dinb(w_n119_0[0]),.dout(n178),.clk(gclk));
	jand g093(.dina(w_n178_3[1]),.dinb(w_G201gat_1[0]),.dout(n179),.clk(gclk));
	jor g094(.dina(w_dff_B_49ONw7UW7_0),.dinb(n174),.dout(n180),.clk(gclk));
	jnot g095(.din(w_G201gat_0[2]),.dout(n181),.clk(gclk));
	jnot g096(.din(w_n148_1[1]),.dout(n182),.clk(gclk));
	jnot g097(.din(w_G126gat_0[0]),.dout(n183),.clk(gclk));
	jnot g098(.din(w_G51gat_0[2]),.dout(n184),.clk(gclk));
	jor g099(.dina(w_n99_0[0]),.dinb(w_dff_B_5qfs6eGb0_1),.dout(n185),.clk(gclk));
	jor g100(.dina(w_n152_0[0]),.dinb(w_n167_0[0]),.dout(n186),.clk(gclk));
	jor g101(.dina(n186),.dinb(w_n185_0[1]),.dout(n187),.clk(gclk));
	jor g102(.dina(n187),.dinb(w_n149_0[0]),.dout(n188),.clk(gclk));
	jand g103(.dina(w_n162_0[0]),.dinb(n188),.dout(n189),.clk(gclk));
	jor g104(.dina(n189),.dinb(w_dff_B_ArAGjGG74_1),.dout(n190),.clk(gclk));
	jnot g105(.din(w_G153gat_0[1]),.dout(n191),.clk(gclk));
	jor g106(.dina(w_n151_0[0]),.dinb(w_n185_0[0]),.dout(n192),.clk(gclk));
	jor g107(.dina(n192),.dinb(w_n95_0[0]),.dout(n193),.clk(gclk));
	jand g108(.dina(n193),.dinb(w_G1gat_0[1]),.dout(n194),.clk(gclk));
	jor g109(.dina(n194),.dinb(w_dff_B_2ZMWjlJC5_1),.dout(n195),.clk(gclk));
	jand g110(.dina(n195),.dinb(n190),.dout(n196),.clk(gclk));
	jand g111(.dina(n196),.dinb(w_dff_B_qXTKOI5C0_1),.dout(n197),.clk(gclk));
	jxor g112(.dina(w_n197_0[2]),.dinb(w_n181_0[2]),.dout(n198),.clk(gclk));
	jand g113(.dina(w_n198_0[2]),.dinb(w_G228gat_3[1]),.dout(n199),.clk(gclk));
	jand g114(.dina(w_n173_0[0]),.dinb(w_G201gat_0[1]),.dout(n200),.clk(gclk));
	jand g115(.dina(w_n200_0[1]),.dinb(w_G237gat_3[1]),.dout(n201),.clk(gclk));
	jand g116(.dina(w_G210gat_3[1]),.dinb(w_G121gat_0[1]),.dout(n202),.clk(gclk));
	jand g117(.dina(G267gat),.dinb(w_G255gat_0[2]),.dout(n203),.clk(gclk));
	jor g118(.dina(n203),.dinb(n202),.dout(n204),.clk(gclk));
	jor g119(.dina(w_dff_B_FpHV7IlO9_0),.dinb(n201),.dout(n205),.clk(gclk));
	jor g120(.dina(n205),.dinb(w_dff_B_8UW0a6hs8_1),.dout(n206),.clk(gclk));
	jor g121(.dina(n206),.dinb(w_dff_B_MfuJcyUF1_1),.dout(n207),.clk(gclk));
	jor g122(.dina(w_n198_0[1]),.dinb(w_G261gat_0[2]),.dout(n208),.clk(gclk));
	jnot g123(.din(w_G261gat_0[1]),.dout(n209),.clk(gclk));
	jnot g124(.din(w_n198_0[0]),.dout(n210),.clk(gclk));
	jor g125(.dina(n210),.dinb(w_n209_0[1]),.dout(n211),.clk(gclk));
	jand g126(.dina(n211),.dinb(w_G219gat_3[2]),.dout(n212),.clk(gclk));
	jand g127(.dina(n212),.dinb(w_dff_B_dweSJyXE7_1),.dout(n213),.clk(gclk));
	jor g128(.dina(n213),.dinb(n207),.dout(w_dff_A_XpWbAcL04_2),.clk(gclk));
	jand g129(.dina(w_n164_3[0]),.dinb(w_G111gat_0[1]),.dout(n215),.clk(gclk));
	jand g130(.dina(w_n170_1[0]),.dinb(w_G143gat_0[1]),.dout(n216),.clk(gclk));
	jor g131(.dina(n216),.dinb(w_n148_1[0]),.dout(n217),.clk(gclk));
	jor g132(.dina(n217),.dinb(n215),.dout(n218),.clk(gclk));
	jxor g133(.dina(w_n218_1[1]),.dinb(w_G183gat_1[1]),.dout(n219),.clk(gclk));
	jand g134(.dina(w_n219_0[2]),.dinb(w_G228gat_3[0]),.dout(n220),.clk(gclk));
	jand g135(.dina(w_n178_3[0]),.dinb(w_G183gat_1[0]),.dout(n221),.clk(gclk));
	jand g136(.dina(w_n218_1[0]),.dinb(w_G183gat_0[2]),.dout(n222),.clk(gclk));
	jand g137(.dina(w_n222_0[2]),.dinb(w_G237gat_3[0]),.dout(n223),.clk(gclk));
	jand g138(.dina(w_n218_0[2]),.dinb(w_G246gat_3[0]),.dout(n224),.clk(gclk));
	jand g139(.dina(w_G210gat_3[0]),.dinb(w_G106gat_0[1]),.dout(n225),.clk(gclk));
	jor g140(.dina(w_dff_B_fVBiDBSq8_0),.dinb(n224),.dout(n226),.clk(gclk));
	jor g141(.dina(n226),.dinb(n223),.dout(n227),.clk(gclk));
	jor g142(.dina(n227),.dinb(w_dff_B_n6JYwdGJ7_1),.dout(n228),.clk(gclk));
	jor g143(.dina(n228),.dinb(w_dff_B_4sDERiW18_1),.dout(n229),.clk(gclk));
	jand g144(.dina(w_n164_2[2]),.dinb(w_G116gat_0[1]),.dout(n230),.clk(gclk));
	jand g145(.dina(w_n170_0[2]),.dinb(w_G146gat_0[1]),.dout(n231),.clk(gclk));
	jor g146(.dina(n231),.dinb(w_n148_0[2]),.dout(n232),.clk(gclk));
	jor g147(.dina(n232),.dinb(n230),.dout(n233),.clk(gclk));
	jand g148(.dina(w_n233_1[1]),.dinb(w_G189gat_2[0]),.dout(n234),.clk(gclk));
	jor g149(.dina(w_n233_1[0]),.dinb(w_G189gat_1[2]),.dout(n235),.clk(gclk));
	jand g150(.dina(w_n164_2[1]),.dinb(w_G121gat_0[0]),.dout(n236),.clk(gclk));
	jand g151(.dina(w_n170_0[1]),.dinb(w_G149gat_0[1]),.dout(n237),.clk(gclk));
	jor g152(.dina(n237),.dinb(w_n148_0[1]),.dout(n238),.clk(gclk));
	jor g153(.dina(n238),.dinb(n236),.dout(n239),.clk(gclk));
	jand g154(.dina(w_n239_1[1]),.dinb(w_G195gat_2[0]),.dout(n240),.clk(gclk));
	jor g155(.dina(w_n239_1[0]),.dinb(w_G195gat_1[2]),.dout(n241),.clk(gclk));
	jand g156(.dina(w_n197_0[1]),.dinb(w_n181_0[1]),.dout(n242),.clk(gclk));
	jnot g157(.din(w_n242_0[1]),.dout(n243),.clk(gclk));
	jor g158(.dina(w_n200_0[0]),.dinb(w_G261gat_0[0]),.dout(n244),.clk(gclk));
	jand g159(.dina(n244),.dinb(n243),.dout(n245),.clk(gclk));
	jand g160(.dina(w_n245_0[1]),.dinb(w_n241_0[1]),.dout(n246),.clk(gclk));
	jor g161(.dina(n246),.dinb(w_n240_0[1]),.dout(n247),.clk(gclk));
	jand g162(.dina(w_n247_0[1]),.dinb(w_n235_0[1]),.dout(n248),.clk(gclk));
	jor g163(.dina(n248),.dinb(w_n234_0[1]),.dout(n249),.clk(gclk));
	jor g164(.dina(w_n249_0[1]),.dinb(w_n219_0[1]),.dout(n250),.clk(gclk));
	jnot g165(.din(w_n219_0[0]),.dout(n251),.clk(gclk));
	jnot g166(.din(w_n234_0[0]),.dout(n252),.clk(gclk));
	jnot g167(.din(w_n235_0[0]),.dout(n253),.clk(gclk));
	jnot g168(.din(w_n240_0[0]),.dout(n254),.clk(gclk));
	jnot g169(.din(w_n241_0[0]),.dout(n255),.clk(gclk));
	jor g170(.dina(w_n197_0[0]),.dinb(w_n181_0[0]),.dout(n256),.clk(gclk));
	jand g171(.dina(n256),.dinb(w_n209_0[0]),.dout(n257),.clk(gclk));
	jor g172(.dina(n257),.dinb(w_n242_0[0]),.dout(n258),.clk(gclk));
	jor g173(.dina(w_n258_0[1]),.dinb(w_dff_B_LzIDozHE7_1),.dout(n259),.clk(gclk));
	jand g174(.dina(n259),.dinb(w_dff_B_Zzo3shUD6_1),.dout(n260),.clk(gclk));
	jor g175(.dina(w_n260_0[1]),.dinb(w_dff_B_wSLV5KIX0_1),.dout(n261),.clk(gclk));
	jand g176(.dina(n261),.dinb(w_dff_B_dKGR2FA92_1),.dout(n262),.clk(gclk));
	jor g177(.dina(w_n262_0[1]),.dinb(w_dff_B_eNvjwhZd4_1),.dout(n263),.clk(gclk));
	jand g178(.dina(n263),.dinb(w_G219gat_3[1]),.dout(n264),.clk(gclk));
	jand g179(.dina(n264),.dinb(w_dff_B_Zy4hPM1a2_1),.dout(n265),.clk(gclk));
	jor g180(.dina(n265),.dinb(w_dff_B_chD6sUN56_1),.dout(w_dff_A_4HrvKHDq8_2),.clk(gclk));
	jxor g181(.dina(w_n233_0[2]),.dinb(w_G189gat_1[1]),.dout(n267),.clk(gclk));
	jand g182(.dina(w_n267_0[2]),.dinb(w_G228gat_2[2]),.dout(n268),.clk(gclk));
	jand g183(.dina(w_G210gat_2[2]),.dinb(w_G111gat_0[0]),.dout(n269),.clk(gclk));
	jand g184(.dina(w_G237gat_2[2]),.dinb(w_G189gat_1[0]),.dout(n270),.clk(gclk));
	jor g185(.dina(n270),.dinb(w_G246gat_2[2]),.dout(n271),.clk(gclk));
	jand g186(.dina(w_dff_B_2tEvSQQL6_0),.dinb(w_n233_0[1]),.dout(n272),.clk(gclk));
	jor g187(.dina(n272),.dinb(w_dff_B_Pyg5iKqF8_1),.dout(n273),.clk(gclk));
	jand g188(.dina(G259gat),.dinb(w_G255gat_0[1]),.dout(n274),.clk(gclk));
	jand g189(.dina(w_n178_2[2]),.dinb(w_G189gat_0[2]),.dout(n275),.clk(gclk));
	jor g190(.dina(n275),.dinb(w_dff_B_vrb2f6Eq5_1),.dout(n276),.clk(gclk));
	jor g191(.dina(w_dff_B_rkhPEvKP7_0),.dinb(n273),.dout(n277),.clk(gclk));
	jor g192(.dina(n277),.dinb(w_dff_B_UnPMVXid7_1),.dout(n278),.clk(gclk));
	jor g193(.dina(w_n267_0[1]),.dinb(w_n247_0[0]),.dout(n279),.clk(gclk));
	jnot g194(.din(w_n267_0[0]),.dout(n280),.clk(gclk));
	jor g195(.dina(w_dff_B_cqmCFRno5_0),.dinb(w_n260_0[0]),.dout(n281),.clk(gclk));
	jand g196(.dina(n281),.dinb(w_G219gat_3[0]),.dout(n282),.clk(gclk));
	jand g197(.dina(n282),.dinb(w_dff_B_EEoS2hDm7_1),.dout(n283),.clk(gclk));
	jor g198(.dina(n283),.dinb(w_dff_B_M5R1DhEI3_1),.dout(w_dff_A_UT8qrq8w4_2),.clk(gclk));
	jxor g199(.dina(w_n239_0[2]),.dinb(w_G195gat_1[1]),.dout(n285),.clk(gclk));
	jand g200(.dina(w_n285_0[2]),.dinb(w_G228gat_2[1]),.dout(n286),.clk(gclk));
	jand g201(.dina(w_G210gat_2[1]),.dinb(w_G116gat_0[0]),.dout(n287),.clk(gclk));
	jand g202(.dina(w_G237gat_2[1]),.dinb(w_G195gat_1[0]),.dout(n288),.clk(gclk));
	jor g203(.dina(n288),.dinb(w_G246gat_2[1]),.dout(n289),.clk(gclk));
	jand g204(.dina(w_dff_B_fFdRJIrJ7_0),.dinb(w_n239_0[1]),.dout(n290),.clk(gclk));
	jor g205(.dina(n290),.dinb(w_dff_B_8okNkrcH4_1),.dout(n291),.clk(gclk));
	jand g206(.dina(w_n178_2[1]),.dinb(w_G195gat_0[2]),.dout(n292),.clk(gclk));
	jand g207(.dina(G260gat),.dinb(w_G255gat_0[0]),.dout(n293),.clk(gclk));
	jor g208(.dina(w_dff_B_IaTZyc2r2_0),.dinb(n292),.dout(n294),.clk(gclk));
	jor g209(.dina(w_dff_B_XB3EYXri9_0),.dinb(n291),.dout(n295),.clk(gclk));
	jor g210(.dina(n295),.dinb(w_dff_B_wEPRavaN2_1),.dout(n296),.clk(gclk));
	jor g211(.dina(w_n285_0[1]),.dinb(w_n245_0[0]),.dout(n297),.clk(gclk));
	jnot g212(.din(w_n285_0[0]),.dout(n298),.clk(gclk));
	jor g213(.dina(w_dff_B_taFFIebQ6_0),.dinb(w_n258_0[0]),.dout(n299),.clk(gclk));
	jand g214(.dina(n299),.dinb(w_G219gat_2[2]),.dout(n300),.clk(gclk));
	jand g215(.dina(n300),.dinb(w_dff_B_fF2QgabW1_1),.dout(n301),.clk(gclk));
	jor g216(.dina(n301),.dinb(w_dff_B_hvvMwwgx5_1),.dout(w_dff_A_iVhb6Mw44_2),.clk(gclk));
	jand g217(.dina(w_n168_0[0]),.dinb(w_G55gat_0[0]),.dout(n303),.clk(gclk));
	jand g218(.dina(w_n303_1[1]),.dinb(w_G143gat_0[0]),.dout(n304),.clk(gclk));
	jand g219(.dina(w_n146_0[0]),.dinb(w_G17gat_1[0]),.dout(n305),.clk(gclk));
	jand g220(.dina(n305),.dinb(w_n144_0[0]),.dout(n306),.clk(gclk));
	jor g221(.dina(w_n306_1[1]),.dinb(w_dff_B_wWgacB2x5_1),.dout(n307),.clk(gclk));
	jand g222(.dina(w_n164_2[0]),.dinb(w_G91gat_0[1]),.dout(n308),.clk(gclk));
	jand g223(.dina(w_G138gat_1[1]),.dinb(w_G8gat_0[0]),.dout(n309),.clk(gclk));
	jor g224(.dina(w_dff_B_Bw7zreyl4_0),.dinb(n308),.dout(n310),.clk(gclk));
	jor g225(.dina(n310),.dinb(w_dff_B_vetATD6j3_1),.dout(n311),.clk(gclk));
	jand g226(.dina(w_n311_1[2]),.dinb(w_G159gat_1[1]),.dout(n312),.clk(gclk));
	jor g227(.dina(w_n311_1[1]),.dinb(w_G159gat_1[0]),.dout(n313),.clk(gclk));
	jand g228(.dina(w_n164_1[2]),.dinb(w_G96gat_0[1]),.dout(n314),.clk(gclk));
	jand g229(.dina(w_n303_1[0]),.dinb(w_G146gat_0[0]),.dout(n315),.clk(gclk));
	jand g230(.dina(w_G138gat_1[0]),.dinb(w_G51gat_0[1]),.dout(n316),.clk(gclk));
	jor g231(.dina(w_dff_B_1NlFHSi64_0),.dinb(n315),.dout(n317),.clk(gclk));
	jor g232(.dina(w_dff_B_IWySEGWJ5_0),.dinb(n314),.dout(n318),.clk(gclk));
	jor g233(.dina(n318),.dinb(w_n306_1[0]),.dout(n319),.clk(gclk));
	jand g234(.dina(w_n319_1[2]),.dinb(w_G165gat_1[1]),.dout(n320),.clk(gclk));
	jor g235(.dina(w_n319_1[1]),.dinb(w_G165gat_1[0]),.dout(n321),.clk(gclk));
	jand g236(.dina(w_n164_1[1]),.dinb(w_G101gat_0[1]),.dout(n322),.clk(gclk));
	jand g237(.dina(w_n303_0[2]),.dinb(w_G149gat_0[0]),.dout(n323),.clk(gclk));
	jand g238(.dina(w_G138gat_0[2]),.dinb(w_G17gat_0[2]),.dout(n324),.clk(gclk));
	jor g239(.dina(w_dff_B_y0VubNw90_0),.dinb(n323),.dout(n325),.clk(gclk));
	jor g240(.dina(w_dff_B_9o2qWziS6_0),.dinb(n322),.dout(n326),.clk(gclk));
	jor g241(.dina(n326),.dinb(w_n306_0[2]),.dout(n327),.clk(gclk));
	jand g242(.dina(w_n327_1[2]),.dinb(w_G171gat_1[1]),.dout(n328),.clk(gclk));
	jor g243(.dina(w_n327_1[1]),.dinb(w_G171gat_1[0]),.dout(n329),.clk(gclk));
	jand g244(.dina(w_n164_1[0]),.dinb(w_G106gat_0[0]),.dout(n330),.clk(gclk));
	jand g245(.dina(w_n303_0[1]),.dinb(w_G153gat_0[0]),.dout(n331),.clk(gclk));
	jand g246(.dina(G152gat),.dinb(w_G138gat_0[1]),.dout(n332),.clk(gclk));
	jor g247(.dina(w_dff_B_8l7w3nKv2_0),.dinb(n331),.dout(n333),.clk(gclk));
	jor g248(.dina(w_dff_B_8lj84eFO9_0),.dinb(n330),.dout(n334),.clk(gclk));
	jor g249(.dina(n334),.dinb(w_n306_0[1]),.dout(n335),.clk(gclk));
	jand g250(.dina(w_n335_1[1]),.dinb(w_G177gat_1[1]),.dout(n336),.clk(gclk));
	jnot g251(.din(w_G177gat_1[0]),.dout(n337),.clk(gclk));
	jnot g252(.din(w_n335_1[0]),.dout(n338),.clk(gclk));
	jand g253(.dina(n338),.dinb(w_dff_B_8sAH4KSb6_1),.dout(n339),.clk(gclk));
	jnot g254(.din(w_n339_0[1]),.dout(n340),.clk(gclk));
	jnot g255(.din(w_G183gat_0[1]),.dout(n341),.clk(gclk));
	jnot g256(.din(w_n218_0[1]),.dout(n342),.clk(gclk));
	jand g257(.dina(n342),.dinb(w_dff_B_7c8zefUi4_1),.dout(n343),.clk(gclk));
	jnot g258(.din(w_n343_0[1]),.dout(n344),.clk(gclk));
	jand g259(.dina(w_n249_0[0]),.dinb(w_dff_B_2AmrlOwa8_1),.dout(n345),.clk(gclk));
	jor g260(.dina(n345),.dinb(w_n222_0[1]),.dout(n346),.clk(gclk));
	jand g261(.dina(w_n346_0[1]),.dinb(w_dff_B_pndSr3IK8_1),.dout(n347),.clk(gclk));
	jor g262(.dina(n347),.dinb(w_n336_0[2]),.dout(n348),.clk(gclk));
	jand g263(.dina(w_n348_0[1]),.dinb(w_n329_0[1]),.dout(n349),.clk(gclk));
	jor g264(.dina(n349),.dinb(w_n328_0[1]),.dout(n350),.clk(gclk));
	jand g265(.dina(w_n350_0[1]),.dinb(w_n321_0[1]),.dout(n351),.clk(gclk));
	jor g266(.dina(n351),.dinb(w_n320_0[1]),.dout(n352),.clk(gclk));
	jand g267(.dina(w_n352_0[1]),.dinb(w_dff_B_5CGT7VBX5_1),.dout(n353),.clk(gclk));
	jor g268(.dina(n353),.dinb(w_dff_B_739TqVXR9_1),.dout(w_dff_A_WiHHet6v3_2),.clk(gclk));
	jxor g269(.dina(w_n335_0[2]),.dinb(w_G177gat_0[2]),.dout(n355),.clk(gclk));
	jnot g270(.din(w_n355_0[1]),.dout(n356),.clk(gclk));
	jand g271(.dina(w_n346_0[0]),.dinb(w_G219gat_2[1]),.dout(n357),.clk(gclk));
	jand g272(.dina(n357),.dinb(w_dff_B_2d5NJLya1_1),.dout(n358),.clk(gclk));
	jnot g273(.din(w_n222_0[0]),.dout(n359),.clk(gclk));
	jor g274(.dina(w_n262_0[0]),.dinb(w_n343_0[0]),.dout(n360),.clk(gclk));
	jand g275(.dina(n360),.dinb(w_dff_B_FNU1id9n2_1),.dout(n361),.clk(gclk));
	jand g276(.dina(w_n361_0[1]),.dinb(w_G219gat_2[0]),.dout(n362),.clk(gclk));
	jor g277(.dina(n362),.dinb(w_G228gat_2[0]),.dout(n363),.clk(gclk));
	jand g278(.dina(n363),.dinb(w_n355_0[0]),.dout(n364),.clk(gclk));
	jand g279(.dina(w_n336_0[1]),.dinb(w_G237gat_2[0]),.dout(n365),.clk(gclk));
	jand g280(.dina(w_n335_0[1]),.dinb(w_G246gat_2[0]),.dout(n366),.clk(gclk));
	jand g281(.dina(w_G210gat_2[0]),.dinb(w_G101gat_0[0]),.dout(n367),.clk(gclk));
	jand g282(.dina(w_n178_2[0]),.dinb(w_G177gat_0[1]),.dout(n368),.clk(gclk));
	jor g283(.dina(n368),.dinb(w_dff_B_Tf9lao5j4_1),.dout(n369),.clk(gclk));
	jor g284(.dina(w_dff_B_mYeIAa6e7_0),.dinb(n366),.dout(n370),.clk(gclk));
	jor g285(.dina(n370),.dinb(n365),.dout(n371),.clk(gclk));
	jor g286(.dina(w_dff_B_mzrTgbZ98_0),.dinb(n364),.dout(n372),.clk(gclk));
	jor g287(.dina(n372),.dinb(w_dff_B_1j2Q1vXK1_1),.dout(w_dff_A_xA640cQm0_2),.clk(gclk));
	jand g288(.dina(w_n311_1[0]),.dinb(w_G237gat_1[2]),.dout(n374),.clk(gclk));
	jor g289(.dina(n374),.dinb(w_n178_1[2]),.dout(n375),.clk(gclk));
	jand g290(.dina(n375),.dinb(w_G159gat_0[2]),.dout(n376),.clk(gclk));
	jxor g291(.dina(w_n311_0[2]),.dinb(w_G159gat_0[1]),.dout(n377),.clk(gclk));
	jand g292(.dina(w_n377_0[2]),.dinb(w_G228gat_1[2]),.dout(n378),.clk(gclk));
	jand g293(.dina(w_G268gat_0[0]),.dinb(w_G210gat_1[2]),.dout(n379),.clk(gclk));
	jor g294(.dina(w_dff_B_biX3YSsp4_0),.dinb(n378),.dout(n380),.clk(gclk));
	jand g295(.dina(w_n311_0[1]),.dinb(w_G246gat_1[2]),.dout(n381),.clk(gclk));
	jor g296(.dina(w_dff_B_CRcWHqIK8_0),.dinb(n380),.dout(n382),.clk(gclk));
	jor g297(.dina(n382),.dinb(w_dff_B_CuOGcm1S0_1),.dout(n383),.clk(gclk));
	jor g298(.dina(w_n377_0[1]),.dinb(w_n352_0[0]),.dout(n384),.clk(gclk));
	jnot g299(.din(w_n320_0[0]),.dout(n385),.clk(gclk));
	jnot g300(.din(w_n321_0[0]),.dout(n386),.clk(gclk));
	jnot g301(.din(w_n328_0[0]),.dout(n387),.clk(gclk));
	jnot g302(.din(w_n329_0[0]),.dout(n388),.clk(gclk));
	jnot g303(.din(w_n336_0[0]),.dout(n389),.clk(gclk));
	jor g304(.dina(w_n361_0[0]),.dinb(w_n339_0[0]),.dout(n390),.clk(gclk));
	jand g305(.dina(n390),.dinb(w_dff_B_WBbSlcL66_1),.dout(n391),.clk(gclk));
	jor g306(.dina(w_n391_0[1]),.dinb(w_dff_B_OwT51m6A4_1),.dout(n392),.clk(gclk));
	jand g307(.dina(n392),.dinb(w_dff_B_pKHPn9e06_1),.dout(n393),.clk(gclk));
	jor g308(.dina(w_n393_0[1]),.dinb(w_dff_B_oMivBNZI9_1),.dout(n394),.clk(gclk));
	jand g309(.dina(n394),.dinb(w_dff_B_NCXRkPjm8_1),.dout(n395),.clk(gclk));
	jnot g310(.din(w_n377_0[0]),.dout(n396),.clk(gclk));
	jor g311(.dina(w_dff_B_QEWIw3vD5_0),.dinb(n395),.dout(n397),.clk(gclk));
	jand g312(.dina(n397),.dinb(w_G219gat_1[2]),.dout(n398),.clk(gclk));
	jand g313(.dina(n398),.dinb(w_dff_B_BOuBIw5n9_1),.dout(n399),.clk(gclk));
	jor g314(.dina(n399),.dinb(w_dff_B_ySyv817e3_1),.dout(G878gat),.clk(gclk));
	jand g315(.dina(w_n319_1[0]),.dinb(w_G237gat_1[1]),.dout(n401),.clk(gclk));
	jor g316(.dina(n401),.dinb(w_n178_1[1]),.dout(n402),.clk(gclk));
	jand g317(.dina(n402),.dinb(w_G165gat_0[2]),.dout(n403),.clk(gclk));
	jxor g318(.dina(w_n319_0[2]),.dinb(w_G165gat_0[1]),.dout(n404),.clk(gclk));
	jand g319(.dina(w_n404_0[2]),.dinb(w_G228gat_1[1]),.dout(n405),.clk(gclk));
	jand g320(.dina(w_G210gat_1[1]),.dinb(w_G91gat_0[0]),.dout(n406),.clk(gclk));
	jor g321(.dina(w_dff_B_88IJbZFB0_0),.dinb(n405),.dout(n407),.clk(gclk));
	jand g322(.dina(w_n319_0[1]),.dinb(w_G246gat_1[1]),.dout(n408),.clk(gclk));
	jor g323(.dina(w_dff_B_aNK4sIva0_0),.dinb(n407),.dout(n409),.clk(gclk));
	jor g324(.dina(n409),.dinb(w_dff_B_ykPKv9fg2_1),.dout(n410),.clk(gclk));
	jor g325(.dina(w_n404_0[1]),.dinb(w_n350_0[0]),.dout(n411),.clk(gclk));
	jnot g326(.din(w_n404_0[0]),.dout(n412),.clk(gclk));
	jor g327(.dina(w_dff_B_3qyVJZYN9_0),.dinb(w_n393_0[0]),.dout(n413),.clk(gclk));
	jand g328(.dina(n413),.dinb(w_G219gat_1[1]),.dout(n414),.clk(gclk));
	jand g329(.dina(n414),.dinb(w_dff_B_T5248S5W0_1),.dout(n415),.clk(gclk));
	jor g330(.dina(n415),.dinb(w_dff_B_UQrHe30V6_1),.dout(w_dff_A_0JlrbuTL8_2),.clk(gclk));
	jand g331(.dina(w_n327_1[0]),.dinb(w_G237gat_1[0]),.dout(n417),.clk(gclk));
	jor g332(.dina(n417),.dinb(w_n178_1[0]),.dout(n418),.clk(gclk));
	jand g333(.dina(n418),.dinb(w_G171gat_0[2]),.dout(n419),.clk(gclk));
	jxor g334(.dina(w_n327_0[2]),.dinb(w_G171gat_0[1]),.dout(n420),.clk(gclk));
	jand g335(.dina(w_n420_0[2]),.dinb(w_G228gat_1[0]),.dout(n421),.clk(gclk));
	jand g336(.dina(w_G210gat_1[0]),.dinb(w_G96gat_0[0]),.dout(n422),.clk(gclk));
	jor g337(.dina(w_dff_B_76toLV5I0_0),.dinb(n421),.dout(n423),.clk(gclk));
	jand g338(.dina(w_n327_0[1]),.dinb(w_G246gat_1[0]),.dout(n424),.clk(gclk));
	jor g339(.dina(w_dff_B_uepjOYpG2_0),.dinb(n423),.dout(n425),.clk(gclk));
	jor g340(.dina(n425),.dinb(w_dff_B_fPSD0pYd9_1),.dout(n426),.clk(gclk));
	jnot g341(.din(w_n420_0[1]),.dout(n427),.clk(gclk));
	jor g342(.dina(w_dff_B_8cj5bpxF6_0),.dinb(w_n391_0[0]),.dout(n428),.clk(gclk));
	jor g343(.dina(w_n420_0[0]),.dinb(w_n348_0[0]),.dout(n429),.clk(gclk));
	jand g344(.dina(n429),.dinb(w_G219gat_1[0]),.dout(n430),.clk(gclk));
	jand g345(.dina(n430),.dinb(w_dff_B_zwOOlXSY7_1),.dout(n431),.clk(gclk));
	jor g346(.dina(n431),.dinb(w_dff_B_U0G8QVwx8_1),.dout(w_dff_A_y8Z8qDZW3_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_dff_A_zMhrg1dP1_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl jspl_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.din(w_G1gat_0[0]));
	jspl jspl_w_G8gat_0(.douta(w_G8gat_0[0]),.doutb(w_G8gat_0[1]),.din(G8gat));
	jspl jspl_w_G13gat_0(.douta(w_G13gat_0[0]),.doutb(w_dff_A_4UdvMskC3_1),.din(G13gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_G17gat_0[0]),.doutb(w_G17gat_0[1]),.doutc(w_G17gat_0[2]),.din(G17gat));
	jspl3 jspl3_w_G17gat_1(.douta(w_dff_A_0P3NhH3m6_0),.doutb(w_dff_A_SzktELqp8_1),.doutc(w_G17gat_1[2]),.din(w_G17gat_0[0]));
	jspl3 jspl3_w_G17gat_2(.douta(w_G17gat_2[0]),.doutb(w_G17gat_2[1]),.doutc(w_dff_A_yTbhX3DK6_2),.din(w_G17gat_0[1]));
	jspl jspl_w_G26gat_0(.douta(w_G26gat_0[0]),.doutb(w_G26gat_0[1]),.din(G26gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_dff_A_Fbey7Ie68_0),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl jspl_w_G36gat_0(.douta(w_G36gat_0[0]),.doutb(w_G36gat_0[1]),.din(G36gat));
	jspl3 jspl3_w_G42gat_0(.douta(w_G42gat_0[0]),.doutb(w_dff_A_NdxYmoco0_1),.doutc(w_dff_A_WqJex0pj3_2),.din(G42gat));
	jspl3 jspl3_w_G42gat_1(.douta(w_dff_A_mXyGRX4a1_0),.doutb(w_G42gat_1[1]),.doutc(w_G42gat_1[2]),.din(w_G42gat_0[0]));
	jspl jspl_w_G42gat_2(.douta(w_G42gat_2[0]),.doutb(w_G42gat_2[1]),.din(w_G42gat_0[1]));
	jspl3 jspl3_w_G51gat_0(.douta(w_G51gat_0[0]),.doutb(w_G51gat_0[1]),.doutc(w_G51gat_0[2]),.din(G51gat));
	jspl jspl_w_G51gat_1(.douta(w_G51gat_1[0]),.doutb(w_dff_A_vtFqyFjw7_1),.din(w_G51gat_0[0]));
	jspl3 jspl3_w_G55gat_0(.douta(w_dff_A_xMdlOa8c6_0),.doutb(w_dff_A_xlfd0ulf6_1),.doutc(w_G55gat_0[2]),.din(w_dff_B_Xcmk5ta43_3));
	jspl3 jspl3_w_G59gat_0(.douta(w_G59gat_0[0]),.doutb(w_G59gat_0[1]),.doutc(w_G59gat_0[2]),.din(G59gat));
	jspl jspl_w_G59gat_1(.douta(w_G59gat_1[0]),.doutb(w_G59gat_1[1]),.din(w_G59gat_0[0]));
	jspl jspl_w_G68gat_0(.douta(w_G68gat_0[0]),.doutb(w_dff_A_8qlIpxDT9_1),.din(G68gat));
	jspl jspl_w_G75gat_0(.douta(w_G75gat_0[0]),.doutb(w_G75gat_0[1]),.din(G75gat));
	jspl3 jspl3_w_G80gat_0(.douta(w_dff_A_OYyvent54_0),.doutb(w_G80gat_0[1]),.doutc(w_dff_A_l1lgeYc16_2),.din(G80gat));
	jspl3 jspl3_w_G91gat_0(.douta(w_G91gat_0[0]),.doutb(w_dff_A_iRg79Aqh2_1),.doutc(w_G91gat_0[2]),.din(G91gat));
	jspl3 jspl3_w_G96gat_0(.douta(w_G96gat_0[0]),.doutb(w_dff_A_J5WWu8vw3_1),.doutc(w_G96gat_0[2]),.din(G96gat));
	jspl3 jspl3_w_G101gat_0(.douta(w_G101gat_0[0]),.doutb(w_dff_A_XWhEy3fA5_1),.doutc(w_G101gat_0[2]),.din(G101gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_V3oXX5jK6_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G111gat_0(.douta(w_G111gat_0[0]),.doutb(w_dff_A_lv8FHbdM0_1),.doutc(w_G111gat_0[2]),.din(G111gat));
	jspl3 jspl3_w_G116gat_0(.douta(w_G116gat_0[0]),.doutb(w_dff_A_6ylewrAP0_1),.doutc(w_G116gat_0[2]),.din(G116gat));
	jspl3 jspl3_w_G121gat_0(.douta(w_dff_A_dUBtC1qd6_0),.doutb(w_G121gat_0[1]),.doutc(w_G121gat_0[2]),.din(G121gat));
	jspl3 jspl3_w_G126gat_0(.douta(w_G126gat_0[0]),.doutb(w_dff_A_pRUoTZao7_1),.doutc(w_G126gat_0[2]),.din(G126gat));
	jspl jspl_w_G130gat_0(.douta(w_G130gat_0[0]),.doutb(w_dff_A_t3vhnhtj8_1),.din(G130gat));
	jspl3 jspl3_w_G138gat_0(.douta(w_G138gat_0[0]),.doutb(w_G138gat_0[1]),.doutc(w_G138gat_0[2]),.din(G138gat));
	jspl jspl_w_G138gat_1(.douta(w_G138gat_1[0]),.doutb(w_G138gat_1[1]),.din(w_G138gat_0[0]));
	jspl jspl_w_G143gat_0(.douta(w_G143gat_0[0]),.doutb(w_dff_A_9XrtnsfL1_1),.din(w_dff_B_W2ds2gT87_2));
	jspl jspl_w_G146gat_0(.douta(w_G146gat_0[0]),.doutb(w_dff_A_itxIFKPu8_1),.din(w_dff_B_y1SzNhuL3_2));
	jspl jspl_w_G149gat_0(.douta(w_G149gat_0[0]),.doutb(w_dff_A_sKjzEtp54_1),.din(w_dff_B_1vyeyFvv6_2));
	jspl3 jspl3_w_G153gat_0(.douta(w_dff_A_8gyjgMM89_0),.doutb(w_G153gat_0[1]),.doutc(w_dff_A_mxXocBMM9_2),.din(G153gat));
	jspl jspl_w_G156gat_0(.douta(w_G156gat_0[0]),.doutb(w_G156gat_0[1]),.din(G156gat));
	jspl3 jspl3_w_G159gat_0(.douta(w_G159gat_0[0]),.doutb(w_dff_A_AhPRc8qB6_1),.doutc(w_dff_A_7PmScMsT7_2),.din(G159gat));
	jspl3 jspl3_w_G159gat_1(.douta(w_dff_A_zhBzgukI2_0),.doutb(w_dff_A_7uwBozfY0_1),.doutc(w_G159gat_1[2]),.din(w_G159gat_0[0]));
	jspl3 jspl3_w_G165gat_0(.douta(w_G165gat_0[0]),.doutb(w_dff_A_1AgLbiWv4_1),.doutc(w_dff_A_bJNZScVw7_2),.din(w_dff_B_JItRWBQW9_3));
	jspl3 jspl3_w_G165gat_1(.douta(w_dff_A_DpfGHxbG0_0),.doutb(w_dff_A_0OM3pxNM4_1),.doutc(w_G165gat_1[2]),.din(w_G165gat_0[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_dff_A_mBVIAkts0_1),.doutc(w_dff_A_5SJuxCkp4_2),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_dff_A_umCUVVI01_0),.doutb(w_dff_A_bcwERkRS3_1),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G177gat_0(.douta(w_G177gat_0[0]),.doutb(w_dff_A_da8ugNZc1_1),.doutc(w_dff_A_Mc204LWe0_2),.din(G177gat));
	jspl3 jspl3_w_G177gat_1(.douta(w_G177gat_1[0]),.doutb(w_dff_A_Rxs8MonY8_1),.doutc(w_G177gat_1[2]),.din(w_G177gat_0[0]));
	jspl3 jspl3_w_G183gat_0(.douta(w_G183gat_0[0]),.doutb(w_G183gat_0[1]),.doutc(w_dff_A_siOi6SOO6_2),.din(G183gat));
	jspl3 jspl3_w_G183gat_1(.douta(w_dff_A_Hx6YmaQx0_0),.doutb(w_dff_A_HC7Nf5MP7_1),.doutc(w_G183gat_1[2]),.din(w_G183gat_0[0]));
	jspl3 jspl3_w_G189gat_0(.douta(w_G189gat_0[0]),.doutb(w_G189gat_0[1]),.doutc(w_dff_A_zjT6Xz1q5_2),.din(G189gat));
	jspl3 jspl3_w_G189gat_1(.douta(w_G189gat_1[0]),.doutb(w_dff_A_sUwDPp9l2_1),.doutc(w_dff_A_Ht5CjNyr0_2),.din(w_G189gat_0[0]));
	jspl jspl_w_G189gat_2(.douta(w_dff_A_bb2z6G8Z2_0),.doutb(w_G189gat_2[1]),.din(w_G189gat_0[1]));
	jspl3 jspl3_w_G195gat_0(.douta(w_G195gat_0[0]),.doutb(w_G195gat_0[1]),.doutc(w_dff_A_INSPVGEJ9_2),.din(G195gat));
	jspl3 jspl3_w_G195gat_1(.douta(w_G195gat_1[0]),.doutb(w_dff_A_8FFtGJvN1_1),.doutc(w_dff_A_T6GTcP1f5_2),.din(w_G195gat_0[0]));
	jspl jspl_w_G195gat_2(.douta(w_dff_A_va40lpK76_0),.doutb(w_G195gat_2[1]),.din(w_G195gat_0[1]));
	jspl3 jspl3_w_G201gat_0(.douta(w_G201gat_0[0]),.doutb(w_dff_A_9fbgEdg66_1),.doutc(w_G201gat_0[2]),.din(G201gat));
	jspl jspl_w_G201gat_1(.douta(w_dff_A_e6G37ysD6_0),.doutb(w_G201gat_1[1]),.din(w_G201gat_0[0]));
	jspl3 jspl3_w_G210gat_0(.douta(w_G210gat_0[0]),.doutb(w_G210gat_0[1]),.doutc(w_G210gat_0[2]),.din(G210gat));
	jspl3 jspl3_w_G210gat_1(.douta(w_G210gat_1[0]),.doutb(w_G210gat_1[1]),.doutc(w_G210gat_1[2]),.din(w_G210gat_0[0]));
	jspl3 jspl3_w_G210gat_2(.douta(w_G210gat_2[0]),.doutb(w_G210gat_2[1]),.doutc(w_G210gat_2[2]),.din(w_G210gat_0[1]));
	jspl jspl_w_G210gat_3(.douta(w_G210gat_3[0]),.doutb(w_G210gat_3[1]),.din(w_G210gat_0[2]));
	jspl3 jspl3_w_G219gat_0(.douta(w_dff_A_QDzD2JfG6_0),.doutb(w_dff_A_NplqoaS60_1),.doutc(w_G219gat_0[2]),.din(w_dff_B_0lpOHo1W6_3));
	jspl3 jspl3_w_G219gat_1(.douta(w_G219gat_1[0]),.doutb(w_dff_A_xUjB7yms6_1),.doutc(w_dff_A_dbuGOjr01_2),.din(w_G219gat_0[0]));
	jspl3 jspl3_w_G219gat_2(.douta(w_dff_A_LbMPQRS23_0),.doutb(w_dff_A_aUXG5iXh7_1),.doutc(w_G219gat_2[2]),.din(w_G219gat_0[1]));
	jspl3 jspl3_w_G219gat_3(.douta(w_dff_A_bTSBTNYh3_0),.doutb(w_dff_A_2NJtDy212_1),.doutc(w_G219gat_3[2]),.din(w_G219gat_0[2]));
	jspl3 jspl3_w_G228gat_0(.douta(w_dff_A_OzA84GwL3_0),.doutb(w_G228gat_0[1]),.doutc(w_G228gat_0[2]),.din(w_dff_B_KbHsGt928_3));
	jspl3 jspl3_w_G228gat_1(.douta(w_G228gat_1[0]),.doutb(w_G228gat_1[1]),.doutc(w_G228gat_1[2]),.din(w_G228gat_0[0]));
	jspl3 jspl3_w_G228gat_2(.douta(w_dff_A_8lffngNi1_0),.doutb(w_G228gat_2[1]),.doutc(w_G228gat_2[2]),.din(w_G228gat_0[1]));
	jspl jspl_w_G228gat_3(.douta(w_G228gat_3[0]),.doutb(w_dff_A_rksPqlv74_1),.din(w_G228gat_0[2]));
	jspl3 jspl3_w_G237gat_0(.douta(w_dff_A_J5vPYbcI0_0),.doutb(w_G237gat_0[1]),.doutc(w_dff_A_PL2qUMNt7_2),.din(G237gat));
	jspl3 jspl3_w_G237gat_1(.douta(w_G237gat_1[0]),.doutb(w_G237gat_1[1]),.doutc(w_G237gat_1[2]),.din(w_G237gat_0[0]));
	jspl3 jspl3_w_G237gat_2(.douta(w_dff_A_msuOIyv83_0),.doutb(w_G237gat_2[1]),.doutc(w_G237gat_2[2]),.din(w_G237gat_0[1]));
	jspl jspl_w_G237gat_3(.douta(w_G237gat_3[0]),.doutb(w_dff_A_nES0KIdl6_1),.din(w_G237gat_0[2]));
	jspl3 jspl3_w_G246gat_0(.douta(w_dff_A_fLHp83Dq1_0),.doutb(w_G246gat_0[1]),.doutc(w_dff_A_NRrZTE351_2),.din(w_dff_B_Fdz3JHdN9_3));
	jspl3 jspl3_w_G246gat_1(.douta(w_G246gat_1[0]),.doutb(w_G246gat_1[1]),.doutc(w_G246gat_1[2]),.din(w_G246gat_0[0]));
	jspl3 jspl3_w_G246gat_2(.douta(w_dff_A_4c2qsVTd9_0),.doutb(w_G246gat_2[1]),.doutc(w_G246gat_2[2]),.din(w_G246gat_0[1]));
	jspl jspl_w_G246gat_3(.douta(w_G246gat_3[0]),.doutb(w_dff_A_WxfrdtCB9_1),.din(w_G246gat_0[2]));
	jspl3 jspl3_w_G255gat_0(.douta(w_G255gat_0[0]),.doutb(w_G255gat_0[1]),.doutc(w_G255gat_0[2]),.din(G255gat));
	jspl3 jspl3_w_G261gat_0(.douta(w_dff_A_eW8E8Ysa1_0),.doutb(w_G261gat_0[1]),.doutc(w_dff_A_4uGeR0Mo1_2),.din(G261gat));
	jspl jspl_w_G268gat_0(.douta(w_G268gat_0[0]),.doutb(w_G268gat_0[1]),.din(G268gat));
	jspl3 jspl3_w_G390gat_0(.douta(w_G390gat_0[0]),.doutb(w_dff_A_qZXECBCX7_1),.doutc(w_dff_A_xEjasLss1_2),.din(G390gat_fa_));
	jspl3 jspl3_w_G447gat_0(.douta(w_G447gat_0[0]),.doutb(w_G447gat_0[1]),.doutc(w_dff_A_WeDFvyBK6_2),.din(G447gat_fa_));
	jspl jspl_w_G447gat_1(.douta(w_G447gat_1),.doutb(w_dff_A_gk8fR03i2_1),.din(w_G447gat_0[0]));
	jspl jspl_w_n86_0(.douta(w_dff_A_vSZJR51x1_0),.doutb(w_n86_0[1]),.din(n86));
	jspl jspl_w_n88_0(.douta(w_n88_0[0]),.doutb(w_n88_0[1]),.din(n88));
	jspl jspl_w_n92_0(.douta(w_n92_0[0]),.doutb(w_n92_0[1]),.din(n92));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n95_0(.douta(w_dff_A_n4EJj6SZ6_0),.doutb(w_n95_0[1]),.doutc(w_dff_A_xdF2g7xZ1_2),.din(n95));
	jspl jspl_w_n97_0(.douta(w_dff_A_RGUelmQ76_0),.doutb(w_n97_0[1]),.din(n97));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl jspl_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_n103_0[1]),.din(w_dff_B_7UlRVwTw9_2));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n109_0(.douta(w_n109_0[0]),.doutb(w_n109_0[1]),.din(n109));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_dff_A_0oyhkhfG6_1),.din(n111));
	jspl jspl_w_n113_0(.douta(w_n113_0[0]),.doutb(w_n113_0[1]),.din(n113));
	jspl3 jspl3_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.doutc(w_n119_0[2]),.din(n119));
	jspl jspl_w_n122_0(.douta(w_n122_0[0]),.doutb(w_dff_A_QmySZphF4_1),.din(n122));
	jspl jspl_w_n144_0(.douta(w_n144_0[0]),.doutb(w_n144_0[1]),.din(w_dff_B_GpVk69285_2));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_n146_0[1]),.din(n146));
	jspl3 jspl3_w_n148_0(.douta(w_n148_0[0]),.doutb(w_n148_0[1]),.doutc(w_n148_0[2]),.din(n148));
	jspl3 jspl3_w_n148_1(.douta(w_n148_1[0]),.doutb(w_n148_1[1]),.doutc(w_dff_A_cZ6N61VB0_2),.din(w_n148_0[0]));
	jspl jspl_w_n149_0(.douta(w_dff_A_NSZkdbwm2_0),.doutb(w_n149_0[1]),.din(n149));
	jspl jspl_w_n151_0(.douta(w_dff_A_wcdBy92T7_0),.doutb(w_n151_0[1]),.din(w_dff_B_UjZgYGR24_2));
	jspl jspl_w_n152_0(.douta(w_dff_A_N45xjSrR7_0),.doutb(w_n152_0[1]),.din(n152));
	jspl jspl_w_n162_0(.douta(w_dff_A_oSWM9JoE8_0),.doutb(w_n162_0[1]),.din(n162));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_n164_0[1]),.doutc(w_n164_0[2]),.din(n164));
	jspl3 jspl3_w_n164_1(.douta(w_n164_1[0]),.doutb(w_n164_1[1]),.doutc(w_n164_1[2]),.din(w_n164_0[0]));
	jspl3 jspl3_w_n164_2(.douta(w_n164_2[0]),.doutb(w_n164_2[1]),.doutc(w_n164_2[2]),.din(w_n164_0[1]));
	jspl jspl_w_n164_3(.douta(w_n164_3[0]),.doutb(w_n164_3[1]),.din(w_n164_0[2]));
	jspl jspl_w_n167_0(.douta(w_n167_0[0]),.doutb(w_n167_0[1]),.din(n167));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.doutc(w_n170_0[2]),.din(n170));
	jspl jspl_w_n170_1(.douta(w_n170_1[0]),.doutb(w_n170_1[1]),.din(w_n170_0[0]));
	jspl jspl_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.din(n173));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_lkCyxoMw0_0),.doutb(w_n178_0[1]),.doutc(w_n178_0[2]),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_n178_1[1]),.doutc(w_n178_1[2]),.din(w_n178_0[0]));
	jspl3 jspl3_w_n178_2(.douta(w_n178_2[0]),.doutb(w_n178_2[1]),.doutc(w_n178_2[2]),.din(w_n178_0[1]));
	jspl jspl_w_n178_3(.douta(w_n178_3[0]),.doutb(w_n178_3[1]),.din(w_n178_0[2]));
	jspl3 jspl3_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.doutc(w_n181_0[2]),.din(w_dff_B_OITevaWi2_3));
	jspl jspl_w_n185_0(.douta(w_n185_0[0]),.doutb(w_n185_0[1]),.din(n185));
	jspl3 jspl3_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.doutc(w_n197_0[2]),.din(n197));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_n198_0[2]),.din(n198));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(n200));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_dff_A_OMBCyLHr2_1),.din(w_dff_B_m4CVuFCK4_2));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_n218_0[2]),.din(n218));
	jspl jspl_w_n218_1(.douta(w_n218_1[0]),.doutb(w_n218_1[1]),.din(w_n218_0[0]));
	jspl3 jspl3_w_n219_0(.douta(w_n219_0[0]),.doutb(w_dff_A_3wgMOOQ69_1),.doutc(w_n219_0[2]),.din(n219));
	jspl3 jspl3_w_n222_0(.douta(w_n222_0[0]),.doutb(w_dff_A_dVLCxt2u1_1),.doutc(w_n222_0[2]),.din(n222));
	jspl3 jspl3_w_n233_0(.douta(w_n233_0[0]),.doutb(w_n233_0[1]),.doutc(w_n233_0[2]),.din(n233));
	jspl jspl_w_n233_1(.douta(w_n233_1[0]),.doutb(w_n233_1[1]),.din(w_n233_0[0]));
	jspl jspl_w_n234_0(.douta(w_n234_0[0]),.doutb(w_dff_A_p9nyq2QR8_1),.din(n234));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_dff_A_vkKBmERZ0_1),.din(n235));
	jspl3 jspl3_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.doutc(w_n239_0[2]),.din(n239));
	jspl jspl_w_n239_1(.douta(w_n239_1[0]),.doutb(w_n239_1[1]),.din(w_n239_0[0]));
	jspl jspl_w_n240_0(.douta(w_n240_0[0]),.doutb(w_dff_A_KyteEw716_1),.din(n240));
	jspl jspl_w_n241_0(.douta(w_n241_0[0]),.doutb(w_dff_A_TPrcG7s28_1),.din(n241));
	jspl jspl_w_n242_0(.douta(w_dff_A_qtE1DAht0_0),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n245_0(.douta(w_n245_0[0]),.doutb(w_n245_0[1]),.din(n245));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n258_0(.douta(w_n258_0[0]),.doutb(w_n258_0[1]),.din(n258));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl jspl_w_n262_0(.douta(w_n262_0[0]),.doutb(w_n262_0[1]),.din(n262));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_dff_A_WuhLNmxI1_1),.doutc(w_n267_0[2]),.din(n267));
	jspl3 jspl3_w_n285_0(.douta(w_n285_0[0]),.doutb(w_dff_A_rusbvijp6_1),.doutc(w_n285_0[2]),.din(n285));
	jspl3 jspl3_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.doutc(w_n303_0[2]),.din(n303));
	jspl jspl_w_n303_1(.douta(w_n303_1[0]),.doutb(w_n303_1[1]),.din(w_n303_0[0]));
	jspl3 jspl3_w_n306_0(.douta(w_n306_0[0]),.doutb(w_dff_A_jwd2PVLX6_1),.doutc(w_dff_A_drFSEFik4_2),.din(n306));
	jspl jspl_w_n306_1(.douta(w_dff_A_BNV2YFLi3_0),.doutb(w_n306_1[1]),.din(w_n306_0[0]));
	jspl3 jspl3_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.doutc(w_n311_0[2]),.din(n311));
	jspl3 jspl3_w_n311_1(.douta(w_n311_1[0]),.doutb(w_n311_1[1]),.doutc(w_n311_1[2]),.din(w_n311_0[0]));
	jspl3 jspl3_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.doutc(w_n319_0[2]),.din(n319));
	jspl3 jspl3_w_n319_1(.douta(w_n319_1[0]),.doutb(w_n319_1[1]),.doutc(w_n319_1[2]),.din(w_n319_0[0]));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_dff_A_1Gws1uM55_1),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_dff_A_5xKtEQe73_1),.din(n321));
	jspl3 jspl3_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.doutc(w_n327_0[2]),.din(n327));
	jspl3 jspl3_w_n327_1(.douta(w_n327_1[0]),.doutb(w_n327_1[1]),.doutc(w_n327_1[2]),.din(w_n327_0[0]));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_dff_A_uiynUS0O5_1),.din(n328));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_dff_A_SA2XWHV18_1),.din(n329));
	jspl3 jspl3_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.doutc(w_n335_0[2]),.din(n335));
	jspl jspl_w_n335_1(.douta(w_n335_1[0]),.doutb(w_n335_1[1]),.din(w_n335_0[0]));
	jspl3 jspl3_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.doutc(w_dff_A_46IsRfaU5_2),.din(n336));
	jspl jspl_w_n339_0(.douta(w_dff_A_5A1BFLOD0_0),.doutb(w_n339_0[1]),.din(n339));
	jspl jspl_w_n343_0(.douta(w_dff_A_n6gYM2im1_0),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(n348));
	jspl jspl_w_n350_0(.douta(w_n350_0[0]),.doutb(w_n350_0[1]),.din(n350));
	jspl jspl_w_n352_0(.douta(w_n352_0[0]),.doutb(w_n352_0[1]),.din(n352));
	jspl jspl_w_n355_0(.douta(w_dff_A_ugG0IBNP3_0),.doutb(w_n355_0[1]),.din(n355));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_dff_A_bBur5LSG3_1),.doutc(w_n377_0[2]),.din(n377));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(n391));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl3 jspl3_w_n404_0(.douta(w_n404_0[0]),.doutb(w_dff_A_uoaCAX433_1),.doutc(w_n404_0[2]),.din(n404));
	jspl3 jspl3_w_n420_0(.douta(w_dff_A_ZnRoYSm69_0),.doutb(w_n420_0[1]),.doutc(w_n420_0[2]),.din(n420));
	jdff dff_B_7UlRVwTw9_2(.din(n103),.dout(w_dff_B_7UlRVwTw9_2),.clk(gclk));
	jdff dff_B_jm6eXLIy3_1(.din(G90gat),.dout(w_dff_B_jm6eXLIy3_1),.clk(gclk));
	jdff dff_B_UsegxPG92_1(.din(n115),.dout(w_dff_B_UsegxPG92_1),.clk(gclk));
	jdff dff_B_rCIjOu890_1(.din(n96),.dout(w_dff_B_rCIjOu890_1),.clk(gclk));
	jdff dff_A_Mp84KvMm0_1(.dout(w_G390gat_0[1]),.din(w_dff_A_Mp84KvMm0_1),.clk(gclk));
	jdff dff_A_qZXECBCX7_1(.dout(w_dff_A_Mp84KvMm0_1),.din(w_dff_A_qZXECBCX7_1),.clk(gclk));
	jdff dff_B_tjY6mTfZ5_1(.din(G74gat),.dout(w_dff_B_tjY6mTfZ5_1),.clk(gclk));
	jdff dff_B_8XYJYpfg6_1(.din(w_dff_B_tjY6mTfZ5_1),.dout(w_dff_B_8XYJYpfg6_1),.clk(gclk));
	jdff dff_B_WVTmUIe00_1(.din(w_dff_B_8XYJYpfg6_1),.dout(w_dff_B_WVTmUIe00_1),.clk(gclk));
	jdff dff_B_iwGeSgRi3_1(.din(G89gat),.dout(w_dff_B_iwGeSgRi3_1),.clk(gclk));
	jdff dff_B_Ul7hI5tG2_1(.din(n127),.dout(w_dff_B_Ul7hI5tG2_1),.clk(gclk));
	jdff dff_B_rPt4A9FB8_1(.din(G135gat),.dout(w_dff_B_rPt4A9FB8_1),.clk(gclk));
	jdff dff_B_7qFlguCr1_1(.din(n136),.dout(w_dff_B_7qFlguCr1_1),.clk(gclk));
	jdff dff_A_t3vhnhtj8_1(.dout(w_G130gat_0[1]),.din(w_dff_A_t3vhnhtj8_1),.clk(gclk));
	jdff dff_B_GCcZzlST4_1(.din(G207gat),.dout(w_dff_B_GCcZzlST4_1),.clk(gclk));
	jdff dff_B_FshnuNUN2_1(.din(n208),.dout(w_dff_B_FshnuNUN2_1),.clk(gclk));
	jdff dff_B_dweSJyXE7_1(.din(w_dff_B_FshnuNUN2_1),.dout(w_dff_B_dweSJyXE7_1),.clk(gclk));
	jdff dff_B_RY5HtDGj1_1(.din(n180),.dout(w_dff_B_RY5HtDGj1_1),.clk(gclk));
	jdff dff_B_MfuJcyUF1_1(.din(w_dff_B_RY5HtDGj1_1),.dout(w_dff_B_MfuJcyUF1_1),.clk(gclk));
	jdff dff_B_8UW0a6hs8_1(.din(n199),.dout(w_dff_B_8UW0a6hs8_1),.clk(gclk));
	jdff dff_B_WoauTbc81_0(.din(n204),.dout(w_dff_B_WoauTbc81_0),.clk(gclk));
	jdff dff_B_YLyCys8s2_0(.din(w_dff_B_WoauTbc81_0),.dout(w_dff_B_YLyCys8s2_0),.clk(gclk));
	jdff dff_B_NGwO7JMM5_0(.din(w_dff_B_YLyCys8s2_0),.dout(w_dff_B_NGwO7JMM5_0),.clk(gclk));
	jdff dff_B_hC8WYbeE4_0(.din(w_dff_B_NGwO7JMM5_0),.dout(w_dff_B_hC8WYbeE4_0),.clk(gclk));
	jdff dff_B_fM8BQZxK7_0(.din(w_dff_B_hC8WYbeE4_0),.dout(w_dff_B_fM8BQZxK7_0),.clk(gclk));
	jdff dff_B_u6fiRcjm4_0(.din(w_dff_B_fM8BQZxK7_0),.dout(w_dff_B_u6fiRcjm4_0),.clk(gclk));
	jdff dff_B_yqChSveb7_0(.din(w_dff_B_u6fiRcjm4_0),.dout(w_dff_B_yqChSveb7_0),.clk(gclk));
	jdff dff_B_1GYBylOX6_0(.din(w_dff_B_yqChSveb7_0),.dout(w_dff_B_1GYBylOX6_0),.clk(gclk));
	jdff dff_B_FpHV7IlO9_0(.din(w_dff_B_1GYBylOX6_0),.dout(w_dff_B_FpHV7IlO9_0),.clk(gclk));
	jdff dff_B_dQlbsjPQ2_0(.din(n179),.dout(w_dff_B_dQlbsjPQ2_0),.clk(gclk));
	jdff dff_B_mV64A36W0_0(.din(w_dff_B_dQlbsjPQ2_0),.dout(w_dff_B_mV64A36W0_0),.clk(gclk));
	jdff dff_B_q2Mmt25B3_0(.din(w_dff_B_mV64A36W0_0),.dout(w_dff_B_q2Mmt25B3_0),.clk(gclk));
	jdff dff_B_1SdJrmBv2_0(.din(w_dff_B_q2Mmt25B3_0),.dout(w_dff_B_1SdJrmBv2_0),.clk(gclk));
	jdff dff_B_49ONw7UW7_0(.din(w_dff_B_1SdJrmBv2_0),.dout(w_dff_B_49ONw7UW7_0),.clk(gclk));
	jdff dff_A_y76Rzs7J3_0(.dout(w_G201gat_1[0]),.din(w_dff_A_y76Rzs7J3_0),.clk(gclk));
	jdff dff_A_ei1QMaBS2_0(.dout(w_dff_A_y76Rzs7J3_0),.din(w_dff_A_ei1QMaBS2_0),.clk(gclk));
	jdff dff_A_WILyofej2_0(.dout(w_dff_A_ei1QMaBS2_0),.din(w_dff_A_WILyofej2_0),.clk(gclk));
	jdff dff_A_e6G37ysD6_0(.dout(w_dff_A_WILyofej2_0),.din(w_dff_A_e6G37ysD6_0),.clk(gclk));
	jdff dff_B_q7n4idcE4_1(.din(n229),.dout(w_dff_B_q7n4idcE4_1),.clk(gclk));
	jdff dff_B_N6Tfx1Ar5_1(.din(w_dff_B_q7n4idcE4_1),.dout(w_dff_B_N6Tfx1Ar5_1),.clk(gclk));
	jdff dff_B_kDcwAYjq9_1(.din(w_dff_B_N6Tfx1Ar5_1),.dout(w_dff_B_kDcwAYjq9_1),.clk(gclk));
	jdff dff_B_NKZFhnVf6_1(.din(w_dff_B_kDcwAYjq9_1),.dout(w_dff_B_NKZFhnVf6_1),.clk(gclk));
	jdff dff_B_u0Hj6Ey13_1(.din(w_dff_B_NKZFhnVf6_1),.dout(w_dff_B_u0Hj6Ey13_1),.clk(gclk));
	jdff dff_B_chD6sUN56_1(.din(w_dff_B_u0Hj6Ey13_1),.dout(w_dff_B_chD6sUN56_1),.clk(gclk));
	jdff dff_B_Zy4hPM1a2_1(.din(n250),.dout(w_dff_B_Zy4hPM1a2_1),.clk(gclk));
	jdff dff_B_6PUZVafV9_1(.din(n251),.dout(w_dff_B_6PUZVafV9_1),.clk(gclk));
	jdff dff_B_FGQFoZA48_1(.din(w_dff_B_6PUZVafV9_1),.dout(w_dff_B_FGQFoZA48_1),.clk(gclk));
	jdff dff_B_3MF9MMpJ7_1(.din(w_dff_B_FGQFoZA48_1),.dout(w_dff_B_3MF9MMpJ7_1),.clk(gclk));
	jdff dff_B_4S9JlBsT8_1(.din(w_dff_B_3MF9MMpJ7_1),.dout(w_dff_B_4S9JlBsT8_1),.clk(gclk));
	jdff dff_B_937gr0qJ4_1(.din(w_dff_B_4S9JlBsT8_1),.dout(w_dff_B_937gr0qJ4_1),.clk(gclk));
	jdff dff_B_eNvjwhZd4_1(.din(w_dff_B_937gr0qJ4_1),.dout(w_dff_B_eNvjwhZd4_1),.clk(gclk));
	jdff dff_B_Skhb3sQy7_1(.din(n220),.dout(w_dff_B_Skhb3sQy7_1),.clk(gclk));
	jdff dff_B_4sDERiW18_1(.din(w_dff_B_Skhb3sQy7_1),.dout(w_dff_B_4sDERiW18_1),.clk(gclk));
	jdff dff_B_3SS9q1EH8_1(.din(n221),.dout(w_dff_B_3SS9q1EH8_1),.clk(gclk));
	jdff dff_B_mzVXuXBw2_1(.din(w_dff_B_3SS9q1EH8_1),.dout(w_dff_B_mzVXuXBw2_1),.clk(gclk));
	jdff dff_B_KHPx0GP12_1(.din(w_dff_B_mzVXuXBw2_1),.dout(w_dff_B_KHPx0GP12_1),.clk(gclk));
	jdff dff_B_yrA6AFeh2_1(.din(w_dff_B_KHPx0GP12_1),.dout(w_dff_B_yrA6AFeh2_1),.clk(gclk));
	jdff dff_B_zI0EUErO1_1(.din(w_dff_B_yrA6AFeh2_1),.dout(w_dff_B_zI0EUErO1_1),.clk(gclk));
	jdff dff_B_n6JYwdGJ7_1(.din(w_dff_B_zI0EUErO1_1),.dout(w_dff_B_n6JYwdGJ7_1),.clk(gclk));
	jdff dff_B_g0kUmBXv6_0(.din(n225),.dout(w_dff_B_g0kUmBXv6_0),.clk(gclk));
	jdff dff_B_LWQkaye88_0(.din(w_dff_B_g0kUmBXv6_0),.dout(w_dff_B_LWQkaye88_0),.clk(gclk));
	jdff dff_B_N9NDx65W8_0(.din(w_dff_B_LWQkaye88_0),.dout(w_dff_B_N9NDx65W8_0),.clk(gclk));
	jdff dff_B_3uoepQeC1_0(.din(w_dff_B_N9NDx65W8_0),.dout(w_dff_B_3uoepQeC1_0),.clk(gclk));
	jdff dff_B_0FLcXZ3g0_0(.din(w_dff_B_3uoepQeC1_0),.dout(w_dff_B_0FLcXZ3g0_0),.clk(gclk));
	jdff dff_B_YQ2SxZa59_0(.din(w_dff_B_0FLcXZ3g0_0),.dout(w_dff_B_YQ2SxZa59_0),.clk(gclk));
	jdff dff_B_Rqvbevwl8_0(.din(w_dff_B_YQ2SxZa59_0),.dout(w_dff_B_Rqvbevwl8_0),.clk(gclk));
	jdff dff_B_fVBiDBSq8_0(.din(w_dff_B_Rqvbevwl8_0),.dout(w_dff_B_fVBiDBSq8_0),.clk(gclk));
	jdff dff_A_WxfrdtCB9_1(.dout(w_G246gat_3[1]),.din(w_dff_A_WxfrdtCB9_1),.clk(gclk));
	jdff dff_A_nES0KIdl6_1(.dout(w_G237gat_3[1]),.din(w_dff_A_nES0KIdl6_1),.clk(gclk));
	jdff dff_A_5hwc9EMo6_1(.dout(w_n219_0[1]),.din(w_dff_A_5hwc9EMo6_1),.clk(gclk));
	jdff dff_A_qyfNGqSj3_1(.dout(w_dff_A_5hwc9EMo6_1),.din(w_dff_A_qyfNGqSj3_1),.clk(gclk));
	jdff dff_A_xdnUc8VM1_1(.dout(w_dff_A_qyfNGqSj3_1),.din(w_dff_A_xdnUc8VM1_1),.clk(gclk));
	jdff dff_A_RJLwdD6t4_1(.dout(w_dff_A_xdnUc8VM1_1),.din(w_dff_A_RJLwdD6t4_1),.clk(gclk));
	jdff dff_A_ElR4gAoP2_1(.dout(w_dff_A_RJLwdD6t4_1),.din(w_dff_A_ElR4gAoP2_1),.clk(gclk));
	jdff dff_A_d4bHz1mU6_1(.dout(w_dff_A_ElR4gAoP2_1),.din(w_dff_A_d4bHz1mU6_1),.clk(gclk));
	jdff dff_A_3wgMOOQ69_1(.dout(w_dff_A_d4bHz1mU6_1),.din(w_dff_A_3wgMOOQ69_1),.clk(gclk));
	jdff dff_A_9fCcpP7I3_0(.dout(w_G183gat_1[0]),.din(w_dff_A_9fCcpP7I3_0),.clk(gclk));
	jdff dff_A_T7XbUg8G8_0(.dout(w_dff_A_9fCcpP7I3_0),.din(w_dff_A_T7XbUg8G8_0),.clk(gclk));
	jdff dff_A_Xm1iaeH91_0(.dout(w_dff_A_T7XbUg8G8_0),.din(w_dff_A_Xm1iaeH91_0),.clk(gclk));
	jdff dff_A_Hx6YmaQx0_0(.dout(w_dff_A_Xm1iaeH91_0),.din(w_dff_A_Hx6YmaQx0_0),.clk(gclk));
	jdff dff_A_KxpzTuRX8_1(.dout(w_G183gat_1[1]),.din(w_dff_A_KxpzTuRX8_1),.clk(gclk));
	jdff dff_A_3Ua3kYjk4_1(.dout(w_dff_A_KxpzTuRX8_1),.din(w_dff_A_3Ua3kYjk4_1),.clk(gclk));
	jdff dff_A_v6aPyT290_1(.dout(w_dff_A_3Ua3kYjk4_1),.din(w_dff_A_v6aPyT290_1),.clk(gclk));
	jdff dff_A_Yx7gMPpu3_1(.dout(w_dff_A_v6aPyT290_1),.din(w_dff_A_Yx7gMPpu3_1),.clk(gclk));
	jdff dff_A_lNxowiTO0_1(.dout(w_dff_A_Yx7gMPpu3_1),.din(w_dff_A_lNxowiTO0_1),.clk(gclk));
	jdff dff_A_QXDDZelg7_1(.dout(w_dff_A_lNxowiTO0_1),.din(w_dff_A_QXDDZelg7_1),.clk(gclk));
	jdff dff_A_qfPZP3rV5_1(.dout(w_dff_A_QXDDZelg7_1),.din(w_dff_A_qfPZP3rV5_1),.clk(gclk));
	jdff dff_A_HC7Nf5MP7_1(.dout(w_dff_A_qfPZP3rV5_1),.din(w_dff_A_HC7Nf5MP7_1),.clk(gclk));
	jdff dff_A_rksPqlv74_1(.dout(w_G228gat_3[1]),.din(w_dff_A_rksPqlv74_1),.clk(gclk));
	jdff dff_B_svI9Jd4Y5_1(.din(n278),.dout(w_dff_B_svI9Jd4Y5_1),.clk(gclk));
	jdff dff_B_sNDaXlOl5_1(.din(w_dff_B_svI9Jd4Y5_1),.dout(w_dff_B_sNDaXlOl5_1),.clk(gclk));
	jdff dff_B_9743cxsy9_1(.din(w_dff_B_sNDaXlOl5_1),.dout(w_dff_B_9743cxsy9_1),.clk(gclk));
	jdff dff_B_qKHZi9Qz3_1(.din(w_dff_B_9743cxsy9_1),.dout(w_dff_B_qKHZi9Qz3_1),.clk(gclk));
	jdff dff_B_M5R1DhEI3_1(.din(w_dff_B_qKHZi9Qz3_1),.dout(w_dff_B_M5R1DhEI3_1),.clk(gclk));
	jdff dff_B_EEoS2hDm7_1(.din(n279),.dout(w_dff_B_EEoS2hDm7_1),.clk(gclk));
	jdff dff_B_62diWx547_0(.din(n280),.dout(w_dff_B_62diWx547_0),.clk(gclk));
	jdff dff_B_dEK1uI2L2_0(.din(w_dff_B_62diWx547_0),.dout(w_dff_B_dEK1uI2L2_0),.clk(gclk));
	jdff dff_B_z2k3bJfc6_0(.din(w_dff_B_dEK1uI2L2_0),.dout(w_dff_B_z2k3bJfc6_0),.clk(gclk));
	jdff dff_B_cqmCFRno5_0(.din(w_dff_B_z2k3bJfc6_0),.dout(w_dff_B_cqmCFRno5_0),.clk(gclk));
	jdff dff_A_0lrckFhS8_0(.dout(w_G219gat_3[0]),.din(w_dff_A_0lrckFhS8_0),.clk(gclk));
	jdff dff_A_O1GOhNL70_0(.dout(w_dff_A_0lrckFhS8_0),.din(w_dff_A_O1GOhNL70_0),.clk(gclk));
	jdff dff_A_bTSBTNYh3_0(.dout(w_dff_A_O1GOhNL70_0),.din(w_dff_A_bTSBTNYh3_0),.clk(gclk));
	jdff dff_A_xj9rrQLS1_1(.dout(w_G219gat_3[1]),.din(w_dff_A_xj9rrQLS1_1),.clk(gclk));
	jdff dff_A_cOAz7LA88_1(.dout(w_dff_A_xj9rrQLS1_1),.din(w_dff_A_cOAz7LA88_1),.clk(gclk));
	jdff dff_A_eJlvrSJz1_1(.dout(w_dff_A_cOAz7LA88_1),.din(w_dff_A_eJlvrSJz1_1),.clk(gclk));
	jdff dff_A_63S5tTKF5_1(.dout(w_dff_A_eJlvrSJz1_1),.din(w_dff_A_63S5tTKF5_1),.clk(gclk));
	jdff dff_A_2NJtDy212_1(.dout(w_dff_A_63S5tTKF5_1),.din(w_dff_A_2NJtDy212_1),.clk(gclk));
	jdff dff_B_UnPMVXid7_1(.din(n268),.dout(w_dff_B_UnPMVXid7_1),.clk(gclk));
	jdff dff_B_PTxwytmR2_0(.din(n276),.dout(w_dff_B_PTxwytmR2_0),.clk(gclk));
	jdff dff_B_EeKn8Uay2_0(.din(w_dff_B_PTxwytmR2_0),.dout(w_dff_B_EeKn8Uay2_0),.clk(gclk));
	jdff dff_B_piIehyoL8_0(.din(w_dff_B_EeKn8Uay2_0),.dout(w_dff_B_piIehyoL8_0),.clk(gclk));
	jdff dff_B_rkhPEvKP7_0(.din(w_dff_B_piIehyoL8_0),.dout(w_dff_B_rkhPEvKP7_0),.clk(gclk));
	jdff dff_B_N5WUdfXS6_1(.din(n274),.dout(w_dff_B_N5WUdfXS6_1),.clk(gclk));
	jdff dff_B_mpGiSs4C5_1(.din(w_dff_B_N5WUdfXS6_1),.dout(w_dff_B_mpGiSs4C5_1),.clk(gclk));
	jdff dff_B_GcVIOolo0_1(.din(w_dff_B_mpGiSs4C5_1),.dout(w_dff_B_GcVIOolo0_1),.clk(gclk));
	jdff dff_B_vrb2f6Eq5_1(.din(w_dff_B_GcVIOolo0_1),.dout(w_dff_B_vrb2f6Eq5_1),.clk(gclk));
	jdff dff_B_akiqZQJF7_1(.din(n269),.dout(w_dff_B_akiqZQJF7_1),.clk(gclk));
	jdff dff_B_RyYg89Tg4_1(.din(w_dff_B_akiqZQJF7_1),.dout(w_dff_B_RyYg89Tg4_1),.clk(gclk));
	jdff dff_B_leIemAES2_1(.din(w_dff_B_RyYg89Tg4_1),.dout(w_dff_B_leIemAES2_1),.clk(gclk));
	jdff dff_B_LFFLHu1r9_1(.din(w_dff_B_leIemAES2_1),.dout(w_dff_B_LFFLHu1r9_1),.clk(gclk));
	jdff dff_B_AF3tlUxG8_1(.din(w_dff_B_LFFLHu1r9_1),.dout(w_dff_B_AF3tlUxG8_1),.clk(gclk));
	jdff dff_B_C224M06e0_1(.din(w_dff_B_AF3tlUxG8_1),.dout(w_dff_B_C224M06e0_1),.clk(gclk));
	jdff dff_B_Ck0f7Him3_1(.din(w_dff_B_C224M06e0_1),.dout(w_dff_B_Ck0f7Him3_1),.clk(gclk));
	jdff dff_B_Pyg5iKqF8_1(.din(w_dff_B_Ck0f7Him3_1),.dout(w_dff_B_Pyg5iKqF8_1),.clk(gclk));
	jdff dff_B_TCsd3mpf6_0(.din(n271),.dout(w_dff_B_TCsd3mpf6_0),.clk(gclk));
	jdff dff_B_czOdfPvk2_0(.din(w_dff_B_TCsd3mpf6_0),.dout(w_dff_B_czOdfPvk2_0),.clk(gclk));
	jdff dff_B_mY9Sqhs87_0(.din(w_dff_B_czOdfPvk2_0),.dout(w_dff_B_mY9Sqhs87_0),.clk(gclk));
	jdff dff_B_XFJMWFuF9_0(.din(w_dff_B_mY9Sqhs87_0),.dout(w_dff_B_XFJMWFuF9_0),.clk(gclk));
	jdff dff_B_jvq62fAN3_0(.din(w_dff_B_XFJMWFuF9_0),.dout(w_dff_B_jvq62fAN3_0),.clk(gclk));
	jdff dff_B_2tEvSQQL6_0(.din(w_dff_B_jvq62fAN3_0),.dout(w_dff_B_2tEvSQQL6_0),.clk(gclk));
	jdff dff_A_eoQKWcvc0_1(.dout(w_n267_0[1]),.din(w_dff_A_eoQKWcvc0_1),.clk(gclk));
	jdff dff_A_vHhr7IKu0_1(.dout(w_dff_A_eoQKWcvc0_1),.din(w_dff_A_vHhr7IKu0_1),.clk(gclk));
	jdff dff_A_DOrvQ7ON2_1(.dout(w_dff_A_vHhr7IKu0_1),.din(w_dff_A_DOrvQ7ON2_1),.clk(gclk));
	jdff dff_A_Hqkzsl6L6_1(.dout(w_dff_A_DOrvQ7ON2_1),.din(w_dff_A_Hqkzsl6L6_1),.clk(gclk));
	jdff dff_A_WuhLNmxI1_1(.dout(w_dff_A_Hqkzsl6L6_1),.din(w_dff_A_WuhLNmxI1_1),.clk(gclk));
	jdff dff_B_RsEIk6Gb6_1(.din(n296),.dout(w_dff_B_RsEIk6Gb6_1),.clk(gclk));
	jdff dff_B_T80HOhX68_1(.din(w_dff_B_RsEIk6Gb6_1),.dout(w_dff_B_T80HOhX68_1),.clk(gclk));
	jdff dff_B_hvvMwwgx5_1(.din(w_dff_B_T80HOhX68_1),.dout(w_dff_B_hvvMwwgx5_1),.clk(gclk));
	jdff dff_B_fF2QgabW1_1(.din(n297),.dout(w_dff_B_fF2QgabW1_1),.clk(gclk));
	jdff dff_B_BdyNMImr7_0(.din(n298),.dout(w_dff_B_BdyNMImr7_0),.clk(gclk));
	jdff dff_B_taFFIebQ6_0(.din(w_dff_B_BdyNMImr7_0),.dout(w_dff_B_taFFIebQ6_0),.clk(gclk));
	jdff dff_B_wEPRavaN2_1(.din(n286),.dout(w_dff_B_wEPRavaN2_1),.clk(gclk));
	jdff dff_B_xcvs9gbx6_0(.din(n294),.dout(w_dff_B_xcvs9gbx6_0),.clk(gclk));
	jdff dff_B_ovA5gLQj8_0(.din(w_dff_B_xcvs9gbx6_0),.dout(w_dff_B_ovA5gLQj8_0),.clk(gclk));
	jdff dff_B_UCoh4UA02_0(.din(w_dff_B_ovA5gLQj8_0),.dout(w_dff_B_UCoh4UA02_0),.clk(gclk));
	jdff dff_B_XB3EYXri9_0(.din(w_dff_B_UCoh4UA02_0),.dout(w_dff_B_XB3EYXri9_0),.clk(gclk));
	jdff dff_B_8Biy8HoB6_0(.din(n293),.dout(w_dff_B_8Biy8HoB6_0),.clk(gclk));
	jdff dff_B_4yAYi2zR9_0(.din(w_dff_B_8Biy8HoB6_0),.dout(w_dff_B_4yAYi2zR9_0),.clk(gclk));
	jdff dff_B_kddekpHh7_0(.din(w_dff_B_4yAYi2zR9_0),.dout(w_dff_B_kddekpHh7_0),.clk(gclk));
	jdff dff_B_IaTZyc2r2_0(.din(w_dff_B_kddekpHh7_0),.dout(w_dff_B_IaTZyc2r2_0),.clk(gclk));
	jdff dff_B_etzueml98_1(.din(n287),.dout(w_dff_B_etzueml98_1),.clk(gclk));
	jdff dff_B_InCJkVUG4_1(.din(w_dff_B_etzueml98_1),.dout(w_dff_B_InCJkVUG4_1),.clk(gclk));
	jdff dff_B_mOLi3xb05_1(.din(w_dff_B_InCJkVUG4_1),.dout(w_dff_B_mOLi3xb05_1),.clk(gclk));
	jdff dff_B_P5yEMZo09_1(.din(w_dff_B_mOLi3xb05_1),.dout(w_dff_B_P5yEMZo09_1),.clk(gclk));
	jdff dff_B_ze1z8i5u7_1(.din(w_dff_B_P5yEMZo09_1),.dout(w_dff_B_ze1z8i5u7_1),.clk(gclk));
	jdff dff_B_SyRsljGN8_1(.din(w_dff_B_ze1z8i5u7_1),.dout(w_dff_B_SyRsljGN8_1),.clk(gclk));
	jdff dff_B_o8kDHWXS4_1(.din(w_dff_B_SyRsljGN8_1),.dout(w_dff_B_o8kDHWXS4_1),.clk(gclk));
	jdff dff_B_8okNkrcH4_1(.din(w_dff_B_o8kDHWXS4_1),.dout(w_dff_B_8okNkrcH4_1),.clk(gclk));
	jdff dff_B_IX2gNa7v7_0(.din(n289),.dout(w_dff_B_IX2gNa7v7_0),.clk(gclk));
	jdff dff_B_2NDYToDA8_0(.din(w_dff_B_IX2gNa7v7_0),.dout(w_dff_B_2NDYToDA8_0),.clk(gclk));
	jdff dff_B_LrOKdEeB7_0(.din(w_dff_B_2NDYToDA8_0),.dout(w_dff_B_LrOKdEeB7_0),.clk(gclk));
	jdff dff_B_oxQqHDfP1_0(.din(w_dff_B_LrOKdEeB7_0),.dout(w_dff_B_oxQqHDfP1_0),.clk(gclk));
	jdff dff_B_E03DlSsn5_0(.din(w_dff_B_oxQqHDfP1_0),.dout(w_dff_B_E03DlSsn5_0),.clk(gclk));
	jdff dff_B_fFdRJIrJ7_0(.din(w_dff_B_E03DlSsn5_0),.dout(w_dff_B_fFdRJIrJ7_0),.clk(gclk));
	jdff dff_A_iDbQWpUL7_1(.dout(w_n285_0[1]),.din(w_dff_A_iDbQWpUL7_1),.clk(gclk));
	jdff dff_A_1rB99uad4_1(.dout(w_dff_A_iDbQWpUL7_1),.din(w_dff_A_1rB99uad4_1),.clk(gclk));
	jdff dff_A_rusbvijp6_1(.dout(w_dff_A_1rB99uad4_1),.din(w_dff_A_rusbvijp6_1),.clk(gclk));
	jdff dff_B_kSsJKgwg1_1(.din(n312),.dout(w_dff_B_kSsJKgwg1_1),.clk(gclk));
	jdff dff_B_43B09MBs2_1(.din(w_dff_B_kSsJKgwg1_1),.dout(w_dff_B_43B09MBs2_1),.clk(gclk));
	jdff dff_B_Op1CpqzH5_1(.din(w_dff_B_43B09MBs2_1),.dout(w_dff_B_Op1CpqzH5_1),.clk(gclk));
	jdff dff_B_0vWjKmTn5_1(.din(w_dff_B_Op1CpqzH5_1),.dout(w_dff_B_0vWjKmTn5_1),.clk(gclk));
	jdff dff_B_cu8ntCVH0_1(.din(w_dff_B_0vWjKmTn5_1),.dout(w_dff_B_cu8ntCVH0_1),.clk(gclk));
	jdff dff_B_uc8tjbyv6_1(.din(w_dff_B_cu8ntCVH0_1),.dout(w_dff_B_uc8tjbyv6_1),.clk(gclk));
	jdff dff_B_uoBxPFug8_1(.din(w_dff_B_uc8tjbyv6_1),.dout(w_dff_B_uoBxPFug8_1),.clk(gclk));
	jdff dff_B_e7sIoZUy2_1(.din(w_dff_B_uoBxPFug8_1),.dout(w_dff_B_e7sIoZUy2_1),.clk(gclk));
	jdff dff_B_qXp7vjer1_1(.din(w_dff_B_e7sIoZUy2_1),.dout(w_dff_B_qXp7vjer1_1),.clk(gclk));
	jdff dff_B_nUQ1juD46_1(.din(w_dff_B_qXp7vjer1_1),.dout(w_dff_B_nUQ1juD46_1),.clk(gclk));
	jdff dff_B_Fbs1rSb97_1(.din(w_dff_B_nUQ1juD46_1),.dout(w_dff_B_Fbs1rSb97_1),.clk(gclk));
	jdff dff_B_bkOfII9t6_1(.din(w_dff_B_Fbs1rSb97_1),.dout(w_dff_B_bkOfII9t6_1),.clk(gclk));
	jdff dff_B_IaomOtqn8_1(.din(w_dff_B_bkOfII9t6_1),.dout(w_dff_B_IaomOtqn8_1),.clk(gclk));
	jdff dff_B_UOxabOif8_1(.din(w_dff_B_IaomOtqn8_1),.dout(w_dff_B_UOxabOif8_1),.clk(gclk));
	jdff dff_B_739TqVXR9_1(.din(w_dff_B_UOxabOif8_1),.dout(w_dff_B_739TqVXR9_1),.clk(gclk));
	jdff dff_B_y0EVvG4E1_1(.din(n313),.dout(w_dff_B_y0EVvG4E1_1),.clk(gclk));
	jdff dff_B_LpLr2JyZ2_1(.din(w_dff_B_y0EVvG4E1_1),.dout(w_dff_B_LpLr2JyZ2_1),.clk(gclk));
	jdff dff_B_I5b885YO1_1(.din(w_dff_B_LpLr2JyZ2_1),.dout(w_dff_B_I5b885YO1_1),.clk(gclk));
	jdff dff_B_d0IVv4Ub4_1(.din(w_dff_B_I5b885YO1_1),.dout(w_dff_B_d0IVv4Ub4_1),.clk(gclk));
	jdff dff_B_beWCevmd1_1(.din(w_dff_B_d0IVv4Ub4_1),.dout(w_dff_B_beWCevmd1_1),.clk(gclk));
	jdff dff_B_KEE8T8tc0_1(.din(w_dff_B_beWCevmd1_1),.dout(w_dff_B_KEE8T8tc0_1),.clk(gclk));
	jdff dff_B_VGdy73zl8_1(.din(w_dff_B_KEE8T8tc0_1),.dout(w_dff_B_VGdy73zl8_1),.clk(gclk));
	jdff dff_B_5YsVXXsZ7_1(.din(w_dff_B_VGdy73zl8_1),.dout(w_dff_B_5YsVXXsZ7_1),.clk(gclk));
	jdff dff_B_sUM1eFew4_1(.din(w_dff_B_5YsVXXsZ7_1),.dout(w_dff_B_sUM1eFew4_1),.clk(gclk));
	jdff dff_B_FA4LMIaE2_1(.din(w_dff_B_sUM1eFew4_1),.dout(w_dff_B_FA4LMIaE2_1),.clk(gclk));
	jdff dff_B_uTybdJek4_1(.din(w_dff_B_FA4LMIaE2_1),.dout(w_dff_B_uTybdJek4_1),.clk(gclk));
	jdff dff_B_NOvm9CIC9_1(.din(w_dff_B_uTybdJek4_1),.dout(w_dff_B_NOvm9CIC9_1),.clk(gclk));
	jdff dff_B_Ltyj8zTE9_1(.din(w_dff_B_NOvm9CIC9_1),.dout(w_dff_B_Ltyj8zTE9_1),.clk(gclk));
	jdff dff_B_5CGT7VBX5_1(.din(w_dff_B_Ltyj8zTE9_1),.dout(w_dff_B_5CGT7VBX5_1),.clk(gclk));
	jdff dff_A_sMswmXfh8_0(.dout(w_G159gat_1[0]),.din(w_dff_A_sMswmXfh8_0),.clk(gclk));
	jdff dff_A_g1wpCx1M3_0(.dout(w_dff_A_sMswmXfh8_0),.din(w_dff_A_g1wpCx1M3_0),.clk(gclk));
	jdff dff_A_pvIYsaCQ1_0(.dout(w_dff_A_g1wpCx1M3_0),.din(w_dff_A_pvIYsaCQ1_0),.clk(gclk));
	jdff dff_A_cdhk59nc5_0(.dout(w_dff_A_pvIYsaCQ1_0),.din(w_dff_A_cdhk59nc5_0),.clk(gclk));
	jdff dff_A_2iBPq9uz9_0(.dout(w_dff_A_cdhk59nc5_0),.din(w_dff_A_2iBPq9uz9_0),.clk(gclk));
	jdff dff_A_hudM42rt9_0(.dout(w_dff_A_2iBPq9uz9_0),.din(w_dff_A_hudM42rt9_0),.clk(gclk));
	jdff dff_A_UlSE4vDR4_0(.dout(w_dff_A_hudM42rt9_0),.din(w_dff_A_UlSE4vDR4_0),.clk(gclk));
	jdff dff_A_5bLlU6QD3_0(.dout(w_dff_A_UlSE4vDR4_0),.din(w_dff_A_5bLlU6QD3_0),.clk(gclk));
	jdff dff_A_zhBzgukI2_0(.dout(w_dff_A_5bLlU6QD3_0),.din(w_dff_A_zhBzgukI2_0),.clk(gclk));
	jdff dff_A_Sqhp3Ll85_1(.dout(w_G159gat_1[1]),.din(w_dff_A_Sqhp3Ll85_1),.clk(gclk));
	jdff dff_A_4gHLy7o37_1(.dout(w_dff_A_Sqhp3Ll85_1),.din(w_dff_A_4gHLy7o37_1),.clk(gclk));
	jdff dff_A_ARIYx2xm2_1(.dout(w_dff_A_4gHLy7o37_1),.din(w_dff_A_ARIYx2xm2_1),.clk(gclk));
	jdff dff_A_WJ1a99Eu2_1(.dout(w_dff_A_ARIYx2xm2_1),.din(w_dff_A_WJ1a99Eu2_1),.clk(gclk));
	jdff dff_A_CF5LVvPB8_1(.dout(w_dff_A_WJ1a99Eu2_1),.din(w_dff_A_CF5LVvPB8_1),.clk(gclk));
	jdff dff_A_3Gv9hCnB8_1(.dout(w_dff_A_CF5LVvPB8_1),.din(w_dff_A_3Gv9hCnB8_1),.clk(gclk));
	jdff dff_A_3fl3KfOT1_1(.dout(w_dff_A_3Gv9hCnB8_1),.din(w_dff_A_3fl3KfOT1_1),.clk(gclk));
	jdff dff_A_xvf3G3pH2_1(.dout(w_dff_A_3fl3KfOT1_1),.din(w_dff_A_xvf3G3pH2_1),.clk(gclk));
	jdff dff_A_7uwBozfY0_1(.dout(w_dff_A_xvf3G3pH2_1),.din(w_dff_A_7uwBozfY0_1),.clk(gclk));
	jdff dff_B_7ml3irGR4_1(.din(n358),.dout(w_dff_B_7ml3irGR4_1),.clk(gclk));
	jdff dff_B_1j2Q1vXK1_1(.din(w_dff_B_7ml3irGR4_1),.dout(w_dff_B_1j2Q1vXK1_1),.clk(gclk));
	jdff dff_B_hdSk64Iz4_0(.din(n371),.dout(w_dff_B_hdSk64Iz4_0),.clk(gclk));
	jdff dff_B_mufPi80S3_0(.din(w_dff_B_hdSk64Iz4_0),.dout(w_dff_B_mufPi80S3_0),.clk(gclk));
	jdff dff_B_jOm5GwFl3_0(.din(w_dff_B_mufPi80S3_0),.dout(w_dff_B_jOm5GwFl3_0),.clk(gclk));
	jdff dff_B_5eDNN2EO0_0(.din(w_dff_B_jOm5GwFl3_0),.dout(w_dff_B_5eDNN2EO0_0),.clk(gclk));
	jdff dff_B_JCJhpumM3_0(.din(w_dff_B_5eDNN2EO0_0),.dout(w_dff_B_JCJhpumM3_0),.clk(gclk));
	jdff dff_B_cr61jGFc1_0(.din(w_dff_B_JCJhpumM3_0),.dout(w_dff_B_cr61jGFc1_0),.clk(gclk));
	jdff dff_B_l4r2TkkW4_0(.din(w_dff_B_cr61jGFc1_0),.dout(w_dff_B_l4r2TkkW4_0),.clk(gclk));
	jdff dff_B_ve2Urtnk4_0(.din(w_dff_B_l4r2TkkW4_0),.dout(w_dff_B_ve2Urtnk4_0),.clk(gclk));
	jdff dff_B_mzrTgbZ98_0(.din(w_dff_B_ve2Urtnk4_0),.dout(w_dff_B_mzrTgbZ98_0),.clk(gclk));
	jdff dff_B_xRbMtTXj2_0(.din(n369),.dout(w_dff_B_xRbMtTXj2_0),.clk(gclk));
	jdff dff_B_I7wZJAGP9_0(.din(w_dff_B_xRbMtTXj2_0),.dout(w_dff_B_I7wZJAGP9_0),.clk(gclk));
	jdff dff_B_dNpIQaZa4_0(.din(w_dff_B_I7wZJAGP9_0),.dout(w_dff_B_dNpIQaZa4_0),.clk(gclk));
	jdff dff_B_mYeIAa6e7_0(.din(w_dff_B_dNpIQaZa4_0),.dout(w_dff_B_mYeIAa6e7_0),.clk(gclk));
	jdff dff_B_ZrWmph8z4_1(.din(n367),.dout(w_dff_B_ZrWmph8z4_1),.clk(gclk));
	jdff dff_B_b78AtUI52_1(.din(w_dff_B_ZrWmph8z4_1),.dout(w_dff_B_b78AtUI52_1),.clk(gclk));
	jdff dff_B_Uzu2GLJV8_1(.din(w_dff_B_b78AtUI52_1),.dout(w_dff_B_Uzu2GLJV8_1),.clk(gclk));
	jdff dff_B_Tf9lao5j4_1(.din(w_dff_B_Uzu2GLJV8_1),.dout(w_dff_B_Tf9lao5j4_1),.clk(gclk));
	jdff dff_A_8FX0cMhG3_0(.dout(w_G246gat_2[0]),.din(w_dff_A_8FX0cMhG3_0),.clk(gclk));
	jdff dff_A_cJALGAt54_0(.dout(w_dff_A_8FX0cMhG3_0),.din(w_dff_A_cJALGAt54_0),.clk(gclk));
	jdff dff_A_JqRJhMZx7_0(.dout(w_dff_A_cJALGAt54_0),.din(w_dff_A_JqRJhMZx7_0),.clk(gclk));
	jdff dff_A_cT7LEdyK6_0(.dout(w_dff_A_JqRJhMZx7_0),.din(w_dff_A_cT7LEdyK6_0),.clk(gclk));
	jdff dff_A_Xzygf2yW8_0(.dout(w_dff_A_cT7LEdyK6_0),.din(w_dff_A_Xzygf2yW8_0),.clk(gclk));
	jdff dff_A_t3rNkFgf8_0(.dout(w_dff_A_Xzygf2yW8_0),.din(w_dff_A_t3rNkFgf8_0),.clk(gclk));
	jdff dff_A_qMjKUJIc7_0(.dout(w_dff_A_t3rNkFgf8_0),.din(w_dff_A_qMjKUJIc7_0),.clk(gclk));
	jdff dff_A_4c2qsVTd9_0(.dout(w_dff_A_qMjKUJIc7_0),.din(w_dff_A_4c2qsVTd9_0),.clk(gclk));
	jdff dff_A_ZbXT1eMg1_0(.dout(w_G237gat_2[0]),.din(w_dff_A_ZbXT1eMg1_0),.clk(gclk));
	jdff dff_A_nUpXirUW7_0(.dout(w_dff_A_ZbXT1eMg1_0),.din(w_dff_A_nUpXirUW7_0),.clk(gclk));
	jdff dff_A_W7RQboxT6_0(.dout(w_dff_A_nUpXirUW7_0),.din(w_dff_A_W7RQboxT6_0),.clk(gclk));
	jdff dff_A_uvat82rS3_0(.dout(w_dff_A_W7RQboxT6_0),.din(w_dff_A_uvat82rS3_0),.clk(gclk));
	jdff dff_A_M8hCgQuY4_0(.dout(w_dff_A_uvat82rS3_0),.din(w_dff_A_M8hCgQuY4_0),.clk(gclk));
	jdff dff_A_W32VJuG51_0(.dout(w_dff_A_M8hCgQuY4_0),.din(w_dff_A_W32VJuG51_0),.clk(gclk));
	jdff dff_A_V930wQB33_0(.dout(w_dff_A_W32VJuG51_0),.din(w_dff_A_V930wQB33_0),.clk(gclk));
	jdff dff_A_xQjEh6la9_0(.dout(w_dff_A_V930wQB33_0),.din(w_dff_A_xQjEh6la9_0),.clk(gclk));
	jdff dff_A_kUbHugkv4_0(.dout(w_dff_A_xQjEh6la9_0),.din(w_dff_A_kUbHugkv4_0),.clk(gclk));
	jdff dff_A_msuOIyv83_0(.dout(w_dff_A_kUbHugkv4_0),.din(w_dff_A_msuOIyv83_0),.clk(gclk));
	jdff dff_A_5QjO1zHm3_0(.dout(w_G228gat_2[0]),.din(w_dff_A_5QjO1zHm3_0),.clk(gclk));
	jdff dff_A_bBt8WHv93_0(.dout(w_dff_A_5QjO1zHm3_0),.din(w_dff_A_bBt8WHv93_0),.clk(gclk));
	jdff dff_A_taTrXRn34_0(.dout(w_dff_A_bBt8WHv93_0),.din(w_dff_A_taTrXRn34_0),.clk(gclk));
	jdff dff_A_WExNutIZ2_0(.dout(w_dff_A_taTrXRn34_0),.din(w_dff_A_WExNutIZ2_0),.clk(gclk));
	jdff dff_A_6PzrO9ha8_0(.dout(w_dff_A_WExNutIZ2_0),.din(w_dff_A_6PzrO9ha8_0),.clk(gclk));
	jdff dff_A_JDXWOT8h5_0(.dout(w_dff_A_6PzrO9ha8_0),.din(w_dff_A_JDXWOT8h5_0),.clk(gclk));
	jdff dff_A_EnobATnd6_0(.dout(w_dff_A_JDXWOT8h5_0),.din(w_dff_A_EnobATnd6_0),.clk(gclk));
	jdff dff_A_SF9bc0cb3_0(.dout(w_dff_A_EnobATnd6_0),.din(w_dff_A_SF9bc0cb3_0),.clk(gclk));
	jdff dff_A_S4IMaqBt1_0(.dout(w_dff_A_SF9bc0cb3_0),.din(w_dff_A_S4IMaqBt1_0),.clk(gclk));
	jdff dff_A_8lffngNi1_0(.dout(w_dff_A_S4IMaqBt1_0),.din(w_dff_A_8lffngNi1_0),.clk(gclk));
	jdff dff_B_dnFacWZS8_1(.din(n356),.dout(w_dff_B_dnFacWZS8_1),.clk(gclk));
	jdff dff_B_ChAj5V7s1_1(.din(w_dff_B_dnFacWZS8_1),.dout(w_dff_B_ChAj5V7s1_1),.clk(gclk));
	jdff dff_B_vcGy6fu08_1(.din(w_dff_B_ChAj5V7s1_1),.dout(w_dff_B_vcGy6fu08_1),.clk(gclk));
	jdff dff_B_YZDxEaTx5_1(.din(w_dff_B_vcGy6fu08_1),.dout(w_dff_B_YZDxEaTx5_1),.clk(gclk));
	jdff dff_B_3o8olskU4_1(.din(w_dff_B_YZDxEaTx5_1),.dout(w_dff_B_3o8olskU4_1),.clk(gclk));
	jdff dff_B_SAMtjTEq0_1(.din(w_dff_B_3o8olskU4_1),.dout(w_dff_B_SAMtjTEq0_1),.clk(gclk));
	jdff dff_B_ROjGXolF2_1(.din(w_dff_B_SAMtjTEq0_1),.dout(w_dff_B_ROjGXolF2_1),.clk(gclk));
	jdff dff_B_2d5NJLya1_1(.din(w_dff_B_ROjGXolF2_1),.dout(w_dff_B_2d5NJLya1_1),.clk(gclk));
	jdff dff_A_HwTXhXM91_0(.dout(w_G219gat_2[0]),.din(w_dff_A_HwTXhXM91_0),.clk(gclk));
	jdff dff_A_SQ9Ieeev8_0(.dout(w_dff_A_HwTXhXM91_0),.din(w_dff_A_SQ9Ieeev8_0),.clk(gclk));
	jdff dff_A_fE1fGi9P7_0(.dout(w_dff_A_SQ9Ieeev8_0),.din(w_dff_A_fE1fGi9P7_0),.clk(gclk));
	jdff dff_A_2h074jhv1_0(.dout(w_dff_A_fE1fGi9P7_0),.din(w_dff_A_2h074jhv1_0),.clk(gclk));
	jdff dff_A_LbMPQRS23_0(.dout(w_dff_A_2h074jhv1_0),.din(w_dff_A_LbMPQRS23_0),.clk(gclk));
	jdff dff_A_6Y535p2A7_1(.dout(w_G219gat_2[1]),.din(w_dff_A_6Y535p2A7_1),.clk(gclk));
	jdff dff_A_E5e6dLfm8_1(.dout(w_dff_A_6Y535p2A7_1),.din(w_dff_A_E5e6dLfm8_1),.clk(gclk));
	jdff dff_A_0svlEpfE3_1(.dout(w_dff_A_E5e6dLfm8_1),.din(w_dff_A_0svlEpfE3_1),.clk(gclk));
	jdff dff_A_hQC7yUKo5_1(.dout(w_dff_A_0svlEpfE3_1),.din(w_dff_A_hQC7yUKo5_1),.clk(gclk));
	jdff dff_A_aUXG5iXh7_1(.dout(w_dff_A_hQC7yUKo5_1),.din(w_dff_A_aUXG5iXh7_1),.clk(gclk));
	jdff dff_A_sEEF8IXs3_0(.dout(w_n355_0[0]),.din(w_dff_A_sEEF8IXs3_0),.clk(gclk));
	jdff dff_A_l8Ou2Oup8_0(.dout(w_dff_A_sEEF8IXs3_0),.din(w_dff_A_l8Ou2Oup8_0),.clk(gclk));
	jdff dff_A_sLMlHiQa3_0(.dout(w_dff_A_l8Ou2Oup8_0),.din(w_dff_A_sLMlHiQa3_0),.clk(gclk));
	jdff dff_A_IOMLg2xW7_0(.dout(w_dff_A_sLMlHiQa3_0),.din(w_dff_A_IOMLg2xW7_0),.clk(gclk));
	jdff dff_A_hS4x2fMT4_0(.dout(w_dff_A_IOMLg2xW7_0),.din(w_dff_A_hS4x2fMT4_0),.clk(gclk));
	jdff dff_A_v00IdZma0_0(.dout(w_dff_A_hS4x2fMT4_0),.din(w_dff_A_v00IdZma0_0),.clk(gclk));
	jdff dff_A_Y9GoIESn6_0(.dout(w_dff_A_v00IdZma0_0),.din(w_dff_A_Y9GoIESn6_0),.clk(gclk));
	jdff dff_A_Ml7zHJL61_0(.dout(w_dff_A_Y9GoIESn6_0),.din(w_dff_A_Ml7zHJL61_0),.clk(gclk));
	jdff dff_A_LucvfUrM8_0(.dout(w_dff_A_Ml7zHJL61_0),.din(w_dff_A_LucvfUrM8_0),.clk(gclk));
	jdff dff_A_ugG0IBNP3_0(.dout(w_dff_A_LucvfUrM8_0),.din(w_dff_A_ugG0IBNP3_0),.clk(gclk));
	jdff dff_B_hetlFEwP1_1(.din(n383),.dout(w_dff_B_hetlFEwP1_1),.clk(gclk));
	jdff dff_B_bAsJDF3r8_1(.din(w_dff_B_hetlFEwP1_1),.dout(w_dff_B_bAsJDF3r8_1),.clk(gclk));
	jdff dff_B_CuATVhDw1_1(.din(w_dff_B_bAsJDF3r8_1),.dout(w_dff_B_CuATVhDw1_1),.clk(gclk));
	jdff dff_B_KX6B9jr39_1(.din(w_dff_B_CuATVhDw1_1),.dout(w_dff_B_KX6B9jr39_1),.clk(gclk));
	jdff dff_B_pycnsQ9g2_1(.din(w_dff_B_KX6B9jr39_1),.dout(w_dff_B_pycnsQ9g2_1),.clk(gclk));
	jdff dff_B_DRk5VQ9g3_1(.din(w_dff_B_pycnsQ9g2_1),.dout(w_dff_B_DRk5VQ9g3_1),.clk(gclk));
	jdff dff_B_Rp3sBDlO8_1(.din(w_dff_B_DRk5VQ9g3_1),.dout(w_dff_B_Rp3sBDlO8_1),.clk(gclk));
	jdff dff_B_SnILTlOj6_1(.din(w_dff_B_Rp3sBDlO8_1),.dout(w_dff_B_SnILTlOj6_1),.clk(gclk));
	jdff dff_B_2Owu4vM60_1(.din(w_dff_B_SnILTlOj6_1),.dout(w_dff_B_2Owu4vM60_1),.clk(gclk));
	jdff dff_B_5TqY3Od33_1(.din(w_dff_B_2Owu4vM60_1),.dout(w_dff_B_5TqY3Od33_1),.clk(gclk));
	jdff dff_B_mHLYSgYu5_1(.din(w_dff_B_5TqY3Od33_1),.dout(w_dff_B_mHLYSgYu5_1),.clk(gclk));
	jdff dff_B_E3TxnA6D4_1(.din(w_dff_B_mHLYSgYu5_1),.dout(w_dff_B_E3TxnA6D4_1),.clk(gclk));
	jdff dff_B_ySyv817e3_1(.din(w_dff_B_E3TxnA6D4_1),.dout(w_dff_B_ySyv817e3_1),.clk(gclk));
	jdff dff_B_BOuBIw5n9_1(.din(n384),.dout(w_dff_B_BOuBIw5n9_1),.clk(gclk));
	jdff dff_B_EBZndK3K6_0(.din(n396),.dout(w_dff_B_EBZndK3K6_0),.clk(gclk));
	jdff dff_B_4HyA0wIj7_0(.din(w_dff_B_EBZndK3K6_0),.dout(w_dff_B_4HyA0wIj7_0),.clk(gclk));
	jdff dff_B_7nSN1BmL7_0(.din(w_dff_B_4HyA0wIj7_0),.dout(w_dff_B_7nSN1BmL7_0),.clk(gclk));
	jdff dff_B_Mn4qUrrj7_0(.din(w_dff_B_7nSN1BmL7_0),.dout(w_dff_B_Mn4qUrrj7_0),.clk(gclk));
	jdff dff_B_0htFlQng5_0(.din(w_dff_B_Mn4qUrrj7_0),.dout(w_dff_B_0htFlQng5_0),.clk(gclk));
	jdff dff_B_fpSwq8P94_0(.din(w_dff_B_0htFlQng5_0),.dout(w_dff_B_fpSwq8P94_0),.clk(gclk));
	jdff dff_B_UT5tplb66_0(.din(w_dff_B_fpSwq8P94_0),.dout(w_dff_B_UT5tplb66_0),.clk(gclk));
	jdff dff_B_1E6aVRxq1_0(.din(w_dff_B_UT5tplb66_0),.dout(w_dff_B_1E6aVRxq1_0),.clk(gclk));
	jdff dff_B_QJ13foVS7_0(.din(w_dff_B_1E6aVRxq1_0),.dout(w_dff_B_QJ13foVS7_0),.clk(gclk));
	jdff dff_B_gYq8QZHH3_0(.din(w_dff_B_QJ13foVS7_0),.dout(w_dff_B_gYq8QZHH3_0),.clk(gclk));
	jdff dff_B_GoXSQxgj3_0(.din(w_dff_B_gYq8QZHH3_0),.dout(w_dff_B_GoXSQxgj3_0),.clk(gclk));
	jdff dff_B_H8v8jYX84_0(.din(w_dff_B_GoXSQxgj3_0),.dout(w_dff_B_H8v8jYX84_0),.clk(gclk));
	jdff dff_B_QEWIw3vD5_0(.din(w_dff_B_H8v8jYX84_0),.dout(w_dff_B_QEWIw3vD5_0),.clk(gclk));
	jdff dff_B_QRPM9spZ3_1(.din(n385),.dout(w_dff_B_QRPM9spZ3_1),.clk(gclk));
	jdff dff_B_kelSn6tj3_1(.din(w_dff_B_QRPM9spZ3_1),.dout(w_dff_B_kelSn6tj3_1),.clk(gclk));
	jdff dff_B_LuaotrBh6_1(.din(w_dff_B_kelSn6tj3_1),.dout(w_dff_B_LuaotrBh6_1),.clk(gclk));
	jdff dff_B_T95ZiaqZ8_1(.din(w_dff_B_LuaotrBh6_1),.dout(w_dff_B_T95ZiaqZ8_1),.clk(gclk));
	jdff dff_B_KBtDMrJr2_1(.din(w_dff_B_T95ZiaqZ8_1),.dout(w_dff_B_KBtDMrJr2_1),.clk(gclk));
	jdff dff_B_R2vPl1S98_1(.din(w_dff_B_KBtDMrJr2_1),.dout(w_dff_B_R2vPl1S98_1),.clk(gclk));
	jdff dff_B_TlhEKaBq6_1(.din(w_dff_B_R2vPl1S98_1),.dout(w_dff_B_TlhEKaBq6_1),.clk(gclk));
	jdff dff_B_f9IH6ZEw6_1(.din(w_dff_B_TlhEKaBq6_1),.dout(w_dff_B_f9IH6ZEw6_1),.clk(gclk));
	jdff dff_B_7iMcDOUP1_1(.din(w_dff_B_f9IH6ZEw6_1),.dout(w_dff_B_7iMcDOUP1_1),.clk(gclk));
	jdff dff_B_hAv3xOsb5_1(.din(w_dff_B_7iMcDOUP1_1),.dout(w_dff_B_hAv3xOsb5_1),.clk(gclk));
	jdff dff_B_KZ88IVSD8_1(.din(w_dff_B_hAv3xOsb5_1),.dout(w_dff_B_KZ88IVSD8_1),.clk(gclk));
	jdff dff_B_NCXRkPjm8_1(.din(w_dff_B_KZ88IVSD8_1),.dout(w_dff_B_NCXRkPjm8_1),.clk(gclk));
	jdff dff_B_iy63Giph4_1(.din(n386),.dout(w_dff_B_iy63Giph4_1),.clk(gclk));
	jdff dff_B_0uytZM3i5_1(.din(w_dff_B_iy63Giph4_1),.dout(w_dff_B_0uytZM3i5_1),.clk(gclk));
	jdff dff_B_ILAq4wtu3_1(.din(w_dff_B_0uytZM3i5_1),.dout(w_dff_B_ILAq4wtu3_1),.clk(gclk));
	jdff dff_B_KUj9xLIJ2_1(.din(w_dff_B_ILAq4wtu3_1),.dout(w_dff_B_KUj9xLIJ2_1),.clk(gclk));
	jdff dff_B_jzw0ZPRT0_1(.din(w_dff_B_KUj9xLIJ2_1),.dout(w_dff_B_jzw0ZPRT0_1),.clk(gclk));
	jdff dff_B_11LjaTYV3_1(.din(w_dff_B_jzw0ZPRT0_1),.dout(w_dff_B_11LjaTYV3_1),.clk(gclk));
	jdff dff_B_wyAxp38r0_1(.din(w_dff_B_11LjaTYV3_1),.dout(w_dff_B_wyAxp38r0_1),.clk(gclk));
	jdff dff_B_U71aS9Tm2_1(.din(w_dff_B_wyAxp38r0_1),.dout(w_dff_B_U71aS9Tm2_1),.clk(gclk));
	jdff dff_B_gdwCuFFa6_1(.din(w_dff_B_U71aS9Tm2_1),.dout(w_dff_B_gdwCuFFa6_1),.clk(gclk));
	jdff dff_B_HpV3k66f6_1(.din(w_dff_B_gdwCuFFa6_1),.dout(w_dff_B_HpV3k66f6_1),.clk(gclk));
	jdff dff_B_oMivBNZI9_1(.din(w_dff_B_HpV3k66f6_1),.dout(w_dff_B_oMivBNZI9_1),.clk(gclk));
	jdff dff_A_UOBezrC63_1(.dout(w_n321_0[1]),.din(w_dff_A_UOBezrC63_1),.clk(gclk));
	jdff dff_A_tj08DVM04_1(.dout(w_dff_A_UOBezrC63_1),.din(w_dff_A_tj08DVM04_1),.clk(gclk));
	jdff dff_A_GlX34DJ62_1(.dout(w_dff_A_tj08DVM04_1),.din(w_dff_A_GlX34DJ62_1),.clk(gclk));
	jdff dff_A_Eq1zp2Dw6_1(.dout(w_dff_A_GlX34DJ62_1),.din(w_dff_A_Eq1zp2Dw6_1),.clk(gclk));
	jdff dff_A_FfZrgR9U5_1(.dout(w_dff_A_Eq1zp2Dw6_1),.din(w_dff_A_FfZrgR9U5_1),.clk(gclk));
	jdff dff_A_4vPJs7jD0_1(.dout(w_dff_A_FfZrgR9U5_1),.din(w_dff_A_4vPJs7jD0_1),.clk(gclk));
	jdff dff_A_46M3CdYD9_1(.dout(w_dff_A_4vPJs7jD0_1),.din(w_dff_A_46M3CdYD9_1),.clk(gclk));
	jdff dff_A_CA4pmh520_1(.dout(w_dff_A_46M3CdYD9_1),.din(w_dff_A_CA4pmh520_1),.clk(gclk));
	jdff dff_A_PXVCfAFW4_1(.dout(w_dff_A_CA4pmh520_1),.din(w_dff_A_PXVCfAFW4_1),.clk(gclk));
	jdff dff_A_xACCcJFQ1_1(.dout(w_dff_A_PXVCfAFW4_1),.din(w_dff_A_xACCcJFQ1_1),.clk(gclk));
	jdff dff_A_GxpxLcHC6_1(.dout(w_dff_A_xACCcJFQ1_1),.din(w_dff_A_GxpxLcHC6_1),.clk(gclk));
	jdff dff_A_5xKtEQe73_1(.dout(w_dff_A_GxpxLcHC6_1),.din(w_dff_A_5xKtEQe73_1),.clk(gclk));
	jdff dff_A_7n9azYfH2_1(.dout(w_n320_0[1]),.din(w_dff_A_7n9azYfH2_1),.clk(gclk));
	jdff dff_A_VQBmQ5rn6_1(.dout(w_dff_A_7n9azYfH2_1),.din(w_dff_A_VQBmQ5rn6_1),.clk(gclk));
	jdff dff_A_79Bw3fkS3_1(.dout(w_dff_A_VQBmQ5rn6_1),.din(w_dff_A_79Bw3fkS3_1),.clk(gclk));
	jdff dff_A_QHEB5vvC2_1(.dout(w_dff_A_79Bw3fkS3_1),.din(w_dff_A_QHEB5vvC2_1),.clk(gclk));
	jdff dff_A_QM3FYHyt2_1(.dout(w_dff_A_QHEB5vvC2_1),.din(w_dff_A_QM3FYHyt2_1),.clk(gclk));
	jdff dff_A_hSBQleYN1_1(.dout(w_dff_A_QM3FYHyt2_1),.din(w_dff_A_hSBQleYN1_1),.clk(gclk));
	jdff dff_A_8WffbtJj9_1(.dout(w_dff_A_hSBQleYN1_1),.din(w_dff_A_8WffbtJj9_1),.clk(gclk));
	jdff dff_A_5XZFMBH08_1(.dout(w_dff_A_8WffbtJj9_1),.din(w_dff_A_5XZFMBH08_1),.clk(gclk));
	jdff dff_A_M4FMebO84_1(.dout(w_dff_A_5XZFMBH08_1),.din(w_dff_A_M4FMebO84_1),.clk(gclk));
	jdff dff_A_lbx1p6qA3_1(.dout(w_dff_A_M4FMebO84_1),.din(w_dff_A_lbx1p6qA3_1),.clk(gclk));
	jdff dff_A_FtpnX7Gw5_1(.dout(w_dff_A_lbx1p6qA3_1),.din(w_dff_A_FtpnX7Gw5_1),.clk(gclk));
	jdff dff_A_Pv1iwvnC9_1(.dout(w_dff_A_FtpnX7Gw5_1),.din(w_dff_A_Pv1iwvnC9_1),.clk(gclk));
	jdff dff_A_1Gws1uM55_1(.dout(w_dff_A_Pv1iwvnC9_1),.din(w_dff_A_1Gws1uM55_1),.clk(gclk));
	jdff dff_A_XJ8O74G11_0(.dout(w_G165gat_1[0]),.din(w_dff_A_XJ8O74G11_0),.clk(gclk));
	jdff dff_A_2iVKTzZv7_0(.dout(w_dff_A_XJ8O74G11_0),.din(w_dff_A_2iVKTzZv7_0),.clk(gclk));
	jdff dff_A_YYYq4rAK1_0(.dout(w_dff_A_2iVKTzZv7_0),.din(w_dff_A_YYYq4rAK1_0),.clk(gclk));
	jdff dff_A_uFtfOXYX4_0(.dout(w_dff_A_YYYq4rAK1_0),.din(w_dff_A_uFtfOXYX4_0),.clk(gclk));
	jdff dff_A_GVEcGpgF3_0(.dout(w_dff_A_uFtfOXYX4_0),.din(w_dff_A_GVEcGpgF3_0),.clk(gclk));
	jdff dff_A_q4TbT11D1_0(.dout(w_dff_A_GVEcGpgF3_0),.din(w_dff_A_q4TbT11D1_0),.clk(gclk));
	jdff dff_A_XUXWmUkq8_0(.dout(w_dff_A_q4TbT11D1_0),.din(w_dff_A_XUXWmUkq8_0),.clk(gclk));
	jdff dff_A_DpfGHxbG0_0(.dout(w_dff_A_XUXWmUkq8_0),.din(w_dff_A_DpfGHxbG0_0),.clk(gclk));
	jdff dff_A_qGQ6gt3I0_1(.dout(w_G165gat_1[1]),.din(w_dff_A_qGQ6gt3I0_1),.clk(gclk));
	jdff dff_A_RyUJF3wM7_1(.dout(w_dff_A_qGQ6gt3I0_1),.din(w_dff_A_RyUJF3wM7_1),.clk(gclk));
	jdff dff_A_BgrZISZv1_1(.dout(w_dff_A_RyUJF3wM7_1),.din(w_dff_A_BgrZISZv1_1),.clk(gclk));
	jdff dff_A_jgFwIr5U7_1(.dout(w_dff_A_BgrZISZv1_1),.din(w_dff_A_jgFwIr5U7_1),.clk(gclk));
	jdff dff_A_Oc9mLevZ3_1(.dout(w_dff_A_jgFwIr5U7_1),.din(w_dff_A_Oc9mLevZ3_1),.clk(gclk));
	jdff dff_A_1FZQV4Ma1_1(.dout(w_dff_A_Oc9mLevZ3_1),.din(w_dff_A_1FZQV4Ma1_1),.clk(gclk));
	jdff dff_A_w9yjRRAl0_1(.dout(w_dff_A_1FZQV4Ma1_1),.din(w_dff_A_w9yjRRAl0_1),.clk(gclk));
	jdff dff_A_0OM3pxNM4_1(.dout(w_dff_A_w9yjRRAl0_1),.din(w_dff_A_0OM3pxNM4_1),.clk(gclk));
	jdff dff_B_CuOGcm1S0_1(.din(n376),.dout(w_dff_B_CuOGcm1S0_1),.clk(gclk));
	jdff dff_B_Z0YVqnoq3_0(.din(n381),.dout(w_dff_B_Z0YVqnoq3_0),.clk(gclk));
	jdff dff_B_CRcWHqIK8_0(.din(w_dff_B_Z0YVqnoq3_0),.dout(w_dff_B_CRcWHqIK8_0),.clk(gclk));
	jdff dff_B_9OUsEcae6_0(.din(n379),.dout(w_dff_B_9OUsEcae6_0),.clk(gclk));
	jdff dff_B_td3bFAe70_0(.din(w_dff_B_9OUsEcae6_0),.dout(w_dff_B_td3bFAe70_0),.clk(gclk));
	jdff dff_B_KtuRsVeg7_0(.din(w_dff_B_td3bFAe70_0),.dout(w_dff_B_KtuRsVeg7_0),.clk(gclk));
	jdff dff_B_qKMce3FS2_0(.din(w_dff_B_KtuRsVeg7_0),.dout(w_dff_B_qKMce3FS2_0),.clk(gclk));
	jdff dff_B_0OwU0sfQ2_0(.din(w_dff_B_qKMce3FS2_0),.dout(w_dff_B_0OwU0sfQ2_0),.clk(gclk));
	jdff dff_B_21aDwmQi0_0(.din(w_dff_B_0OwU0sfQ2_0),.dout(w_dff_B_21aDwmQi0_0),.clk(gclk));
	jdff dff_B_UmnxBDse4_0(.din(w_dff_B_21aDwmQi0_0),.dout(w_dff_B_UmnxBDse4_0),.clk(gclk));
	jdff dff_B_TxpAa5yk6_0(.din(w_dff_B_UmnxBDse4_0),.dout(w_dff_B_TxpAa5yk6_0),.clk(gclk));
	jdff dff_B_y2ynUSV36_0(.din(w_dff_B_TxpAa5yk6_0),.dout(w_dff_B_y2ynUSV36_0),.clk(gclk));
	jdff dff_B_biX3YSsp4_0(.din(w_dff_B_y2ynUSV36_0),.dout(w_dff_B_biX3YSsp4_0),.clk(gclk));
	jdff dff_A_59cUwoyC3_1(.dout(w_n377_0[1]),.din(w_dff_A_59cUwoyC3_1),.clk(gclk));
	jdff dff_A_gVympQoA6_1(.dout(w_dff_A_59cUwoyC3_1),.din(w_dff_A_gVympQoA6_1),.clk(gclk));
	jdff dff_A_UFWYzOYZ4_1(.dout(w_dff_A_gVympQoA6_1),.din(w_dff_A_UFWYzOYZ4_1),.clk(gclk));
	jdff dff_A_9aXzQHFG3_1(.dout(w_dff_A_UFWYzOYZ4_1),.din(w_dff_A_9aXzQHFG3_1),.clk(gclk));
	jdff dff_A_H1v2ywFF4_1(.dout(w_dff_A_9aXzQHFG3_1),.din(w_dff_A_H1v2ywFF4_1),.clk(gclk));
	jdff dff_A_JX1KFojR5_1(.dout(w_dff_A_H1v2ywFF4_1),.din(w_dff_A_JX1KFojR5_1),.clk(gclk));
	jdff dff_A_ZcDVxExB4_1(.dout(w_dff_A_JX1KFojR5_1),.din(w_dff_A_ZcDVxExB4_1),.clk(gclk));
	jdff dff_A_32pX3Qta9_1(.dout(w_dff_A_ZcDVxExB4_1),.din(w_dff_A_32pX3Qta9_1),.clk(gclk));
	jdff dff_A_aRe9hpuv5_1(.dout(w_dff_A_32pX3Qta9_1),.din(w_dff_A_aRe9hpuv5_1),.clk(gclk));
	jdff dff_A_LXmpmsgf0_1(.dout(w_dff_A_aRe9hpuv5_1),.din(w_dff_A_LXmpmsgf0_1),.clk(gclk));
	jdff dff_A_InLg641k6_1(.dout(w_dff_A_LXmpmsgf0_1),.din(w_dff_A_InLg641k6_1),.clk(gclk));
	jdff dff_A_rCpwzjQz6_1(.dout(w_dff_A_InLg641k6_1),.din(w_dff_A_rCpwzjQz6_1),.clk(gclk));
	jdff dff_A_CP52tFaI4_1(.dout(w_dff_A_rCpwzjQz6_1),.din(w_dff_A_CP52tFaI4_1),.clk(gclk));
	jdff dff_A_bBur5LSG3_1(.dout(w_dff_A_CP52tFaI4_1),.din(w_dff_A_bBur5LSG3_1),.clk(gclk));
	jdff dff_B_vetATD6j3_1(.din(n307),.dout(w_dff_B_vetATD6j3_1),.clk(gclk));
	jdff dff_B_T0wICkI14_0(.din(n309),.dout(w_dff_B_T0wICkI14_0),.clk(gclk));
	jdff dff_B_FANpPhwB5_0(.din(w_dff_B_T0wICkI14_0),.dout(w_dff_B_FANpPhwB5_0),.clk(gclk));
	jdff dff_B_10ZvEDF80_0(.din(w_dff_B_FANpPhwB5_0),.dout(w_dff_B_10ZvEDF80_0),.clk(gclk));
	jdff dff_B_pyicbREB9_0(.din(w_dff_B_10ZvEDF80_0),.dout(w_dff_B_pyicbREB9_0),.clk(gclk));
	jdff dff_B_UwvsC6jy9_0(.din(w_dff_B_pyicbREB9_0),.dout(w_dff_B_UwvsC6jy9_0),.clk(gclk));
	jdff dff_B_Bw7zreyl4_0(.din(w_dff_B_UwvsC6jy9_0),.dout(w_dff_B_Bw7zreyl4_0),.clk(gclk));
	jdff dff_B_wWgacB2x5_1(.din(n304),.dout(w_dff_B_wWgacB2x5_1),.clk(gclk));
	jdff dff_A_NrDX6v2g9_1(.dout(w_G159gat_0[1]),.din(w_dff_A_NrDX6v2g9_1),.clk(gclk));
	jdff dff_A_qesOdUex1_1(.dout(w_dff_A_NrDX6v2g9_1),.din(w_dff_A_qesOdUex1_1),.clk(gclk));
	jdff dff_A_WkeiUzpd4_1(.dout(w_dff_A_qesOdUex1_1),.din(w_dff_A_WkeiUzpd4_1),.clk(gclk));
	jdff dff_A_Pd4xpJIf5_1(.dout(w_dff_A_WkeiUzpd4_1),.din(w_dff_A_Pd4xpJIf5_1),.clk(gclk));
	jdff dff_A_DKQFbzJV8_1(.dout(w_dff_A_Pd4xpJIf5_1),.din(w_dff_A_DKQFbzJV8_1),.clk(gclk));
	jdff dff_A_03RQZdCF5_1(.dout(w_dff_A_DKQFbzJV8_1),.din(w_dff_A_03RQZdCF5_1),.clk(gclk));
	jdff dff_A_VcOZFsjM3_1(.dout(w_dff_A_03RQZdCF5_1),.din(w_dff_A_VcOZFsjM3_1),.clk(gclk));
	jdff dff_A_7H3GdROP4_1(.dout(w_dff_A_VcOZFsjM3_1),.din(w_dff_A_7H3GdROP4_1),.clk(gclk));
	jdff dff_A_AhPRc8qB6_1(.dout(w_dff_A_7H3GdROP4_1),.din(w_dff_A_AhPRc8qB6_1),.clk(gclk));
	jdff dff_A_Dpyy9W5a8_2(.dout(w_G159gat_0[2]),.din(w_dff_A_Dpyy9W5a8_2),.clk(gclk));
	jdff dff_A_r5uO8BJM1_2(.dout(w_dff_A_Dpyy9W5a8_2),.din(w_dff_A_r5uO8BJM1_2),.clk(gclk));
	jdff dff_A_N1DY7i6J2_2(.dout(w_dff_A_r5uO8BJM1_2),.din(w_dff_A_N1DY7i6J2_2),.clk(gclk));
	jdff dff_A_rsIkIIhy3_2(.dout(w_dff_A_N1DY7i6J2_2),.din(w_dff_A_rsIkIIhy3_2),.clk(gclk));
	jdff dff_A_4GB2XfD99_2(.dout(w_dff_A_rsIkIIhy3_2),.din(w_dff_A_4GB2XfD99_2),.clk(gclk));
	jdff dff_A_BYklxgVr5_2(.dout(w_dff_A_4GB2XfD99_2),.din(w_dff_A_BYklxgVr5_2),.clk(gclk));
	jdff dff_A_aOsX3niG4_2(.dout(w_dff_A_BYklxgVr5_2),.din(w_dff_A_aOsX3niG4_2),.clk(gclk));
	jdff dff_A_D5LscFzv6_2(.dout(w_dff_A_aOsX3niG4_2),.din(w_dff_A_D5LscFzv6_2),.clk(gclk));
	jdff dff_A_m4bfDoaB5_2(.dout(w_dff_A_D5LscFzv6_2),.din(w_dff_A_m4bfDoaB5_2),.clk(gclk));
	jdff dff_A_xH1AbGAZ5_2(.dout(w_dff_A_m4bfDoaB5_2),.din(w_dff_A_xH1AbGAZ5_2),.clk(gclk));
	jdff dff_A_7PmScMsT7_2(.dout(w_dff_A_xH1AbGAZ5_2),.din(w_dff_A_7PmScMsT7_2),.clk(gclk));
	jdff dff_B_vZh3sQ576_1(.din(n410),.dout(w_dff_B_vZh3sQ576_1),.clk(gclk));
	jdff dff_B_QbP7DQ4V1_1(.din(w_dff_B_vZh3sQ576_1),.dout(w_dff_B_QbP7DQ4V1_1),.clk(gclk));
	jdff dff_B_jieyf3aQ0_1(.din(w_dff_B_QbP7DQ4V1_1),.dout(w_dff_B_jieyf3aQ0_1),.clk(gclk));
	jdff dff_B_bM3Ld3Co3_1(.din(w_dff_B_jieyf3aQ0_1),.dout(w_dff_B_bM3Ld3Co3_1),.clk(gclk));
	jdff dff_B_g67Qs0BX0_1(.din(w_dff_B_bM3Ld3Co3_1),.dout(w_dff_B_g67Qs0BX0_1),.clk(gclk));
	jdff dff_B_Bv12QFqb9_1(.din(w_dff_B_g67Qs0BX0_1),.dout(w_dff_B_Bv12QFqb9_1),.clk(gclk));
	jdff dff_B_vgCJhJqx7_1(.din(w_dff_B_Bv12QFqb9_1),.dout(w_dff_B_vgCJhJqx7_1),.clk(gclk));
	jdff dff_B_l5h5YGp65_1(.din(w_dff_B_vgCJhJqx7_1),.dout(w_dff_B_l5h5YGp65_1),.clk(gclk));
	jdff dff_B_5046kXT62_1(.din(w_dff_B_l5h5YGp65_1),.dout(w_dff_B_5046kXT62_1),.clk(gclk));
	jdff dff_B_QwRYwze47_1(.din(w_dff_B_5046kXT62_1),.dout(w_dff_B_QwRYwze47_1),.clk(gclk));
	jdff dff_B_UQrHe30V6_1(.din(w_dff_B_QwRYwze47_1),.dout(w_dff_B_UQrHe30V6_1),.clk(gclk));
	jdff dff_B_T5248S5W0_1(.din(n411),.dout(w_dff_B_T5248S5W0_1),.clk(gclk));
	jdff dff_B_PtM3Dr2W9_0(.din(n412),.dout(w_dff_B_PtM3Dr2W9_0),.clk(gclk));
	jdff dff_B_rjY96nYx6_0(.din(w_dff_B_PtM3Dr2W9_0),.dout(w_dff_B_rjY96nYx6_0),.clk(gclk));
	jdff dff_B_8UJVHaaO8_0(.din(w_dff_B_rjY96nYx6_0),.dout(w_dff_B_8UJVHaaO8_0),.clk(gclk));
	jdff dff_B_Ko8ulaEL1_0(.din(w_dff_B_8UJVHaaO8_0),.dout(w_dff_B_Ko8ulaEL1_0),.clk(gclk));
	jdff dff_B_EFte2PZh5_0(.din(w_dff_B_Ko8ulaEL1_0),.dout(w_dff_B_EFte2PZh5_0),.clk(gclk));
	jdff dff_B_O1Og2UUj2_0(.din(w_dff_B_EFte2PZh5_0),.dout(w_dff_B_O1Og2UUj2_0),.clk(gclk));
	jdff dff_B_i93QyhJt3_0(.din(w_dff_B_O1Og2UUj2_0),.dout(w_dff_B_i93QyhJt3_0),.clk(gclk));
	jdff dff_B_LufdEjVa5_0(.din(w_dff_B_i93QyhJt3_0),.dout(w_dff_B_LufdEjVa5_0),.clk(gclk));
	jdff dff_B_JXcNqjgB5_0(.din(w_dff_B_LufdEjVa5_0),.dout(w_dff_B_JXcNqjgB5_0),.clk(gclk));
	jdff dff_B_rfQbAPgC3_0(.din(w_dff_B_JXcNqjgB5_0),.dout(w_dff_B_rfQbAPgC3_0),.clk(gclk));
	jdff dff_B_3qyVJZYN9_0(.din(w_dff_B_rfQbAPgC3_0),.dout(w_dff_B_3qyVJZYN9_0),.clk(gclk));
	jdff dff_B_7Pit0s874_1(.din(n387),.dout(w_dff_B_7Pit0s874_1),.clk(gclk));
	jdff dff_B_UBCQA1KC5_1(.din(w_dff_B_7Pit0s874_1),.dout(w_dff_B_UBCQA1KC5_1),.clk(gclk));
	jdff dff_B_JzdIy3vP0_1(.din(w_dff_B_UBCQA1KC5_1),.dout(w_dff_B_JzdIy3vP0_1),.clk(gclk));
	jdff dff_B_E7FeexCx6_1(.din(w_dff_B_JzdIy3vP0_1),.dout(w_dff_B_E7FeexCx6_1),.clk(gclk));
	jdff dff_B_iOkVEekg7_1(.din(w_dff_B_E7FeexCx6_1),.dout(w_dff_B_iOkVEekg7_1),.clk(gclk));
	jdff dff_B_xr8kS8ob6_1(.din(w_dff_B_iOkVEekg7_1),.dout(w_dff_B_xr8kS8ob6_1),.clk(gclk));
	jdff dff_B_1InQcKpH7_1(.din(w_dff_B_xr8kS8ob6_1),.dout(w_dff_B_1InQcKpH7_1),.clk(gclk));
	jdff dff_B_yKijsFl48_1(.din(w_dff_B_1InQcKpH7_1),.dout(w_dff_B_yKijsFl48_1),.clk(gclk));
	jdff dff_B_XYGPfLPa7_1(.din(w_dff_B_yKijsFl48_1),.dout(w_dff_B_XYGPfLPa7_1),.clk(gclk));
	jdff dff_B_pKHPn9e06_1(.din(w_dff_B_XYGPfLPa7_1),.dout(w_dff_B_pKHPn9e06_1),.clk(gclk));
	jdff dff_B_1utYZW6O4_1(.din(n388),.dout(w_dff_B_1utYZW6O4_1),.clk(gclk));
	jdff dff_B_DHFwIxVo5_1(.din(w_dff_B_1utYZW6O4_1),.dout(w_dff_B_DHFwIxVo5_1),.clk(gclk));
	jdff dff_B_SweBN5zZ6_1(.din(w_dff_B_DHFwIxVo5_1),.dout(w_dff_B_SweBN5zZ6_1),.clk(gclk));
	jdff dff_B_sDvaAJgS4_1(.din(w_dff_B_SweBN5zZ6_1),.dout(w_dff_B_sDvaAJgS4_1),.clk(gclk));
	jdff dff_B_Grw3UOcM2_1(.din(w_dff_B_sDvaAJgS4_1),.dout(w_dff_B_Grw3UOcM2_1),.clk(gclk));
	jdff dff_B_Ql2kUoG23_1(.din(w_dff_B_Grw3UOcM2_1),.dout(w_dff_B_Ql2kUoG23_1),.clk(gclk));
	jdff dff_B_wPbLM3uh5_1(.din(w_dff_B_Ql2kUoG23_1),.dout(w_dff_B_wPbLM3uh5_1),.clk(gclk));
	jdff dff_B_wk5YgdTi4_1(.din(w_dff_B_wPbLM3uh5_1),.dout(w_dff_B_wk5YgdTi4_1),.clk(gclk));
	jdff dff_B_OwT51m6A4_1(.din(w_dff_B_wk5YgdTi4_1),.dout(w_dff_B_OwT51m6A4_1),.clk(gclk));
	jdff dff_A_6VJrT6Q04_1(.dout(w_n329_0[1]),.din(w_dff_A_6VJrT6Q04_1),.clk(gclk));
	jdff dff_A_Eeqwj9sL2_1(.dout(w_dff_A_6VJrT6Q04_1),.din(w_dff_A_Eeqwj9sL2_1),.clk(gclk));
	jdff dff_A_9toAGEIR6_1(.dout(w_dff_A_Eeqwj9sL2_1),.din(w_dff_A_9toAGEIR6_1),.clk(gclk));
	jdff dff_A_T12HvpLQ2_1(.dout(w_dff_A_9toAGEIR6_1),.din(w_dff_A_T12HvpLQ2_1),.clk(gclk));
	jdff dff_A_b2vtq1xz3_1(.dout(w_dff_A_T12HvpLQ2_1),.din(w_dff_A_b2vtq1xz3_1),.clk(gclk));
	jdff dff_A_iccYKbFn6_1(.dout(w_dff_A_b2vtq1xz3_1),.din(w_dff_A_iccYKbFn6_1),.clk(gclk));
	jdff dff_A_8xgd9K394_1(.dout(w_dff_A_iccYKbFn6_1),.din(w_dff_A_8xgd9K394_1),.clk(gclk));
	jdff dff_A_WW5FOQ2g6_1(.dout(w_dff_A_8xgd9K394_1),.din(w_dff_A_WW5FOQ2g6_1),.clk(gclk));
	jdff dff_A_wmBO8hgq5_1(.dout(w_dff_A_WW5FOQ2g6_1),.din(w_dff_A_wmBO8hgq5_1),.clk(gclk));
	jdff dff_A_SA2XWHV18_1(.dout(w_dff_A_wmBO8hgq5_1),.din(w_dff_A_SA2XWHV18_1),.clk(gclk));
	jdff dff_A_tv7AzjQJ7_1(.dout(w_n328_0[1]),.din(w_dff_A_tv7AzjQJ7_1),.clk(gclk));
	jdff dff_A_udiWCKmO9_1(.dout(w_dff_A_tv7AzjQJ7_1),.din(w_dff_A_udiWCKmO9_1),.clk(gclk));
	jdff dff_A_EIkbPqy40_1(.dout(w_dff_A_udiWCKmO9_1),.din(w_dff_A_EIkbPqy40_1),.clk(gclk));
	jdff dff_A_fqioc4hn6_1(.dout(w_dff_A_EIkbPqy40_1),.din(w_dff_A_fqioc4hn6_1),.clk(gclk));
	jdff dff_A_xHhtf05p2_1(.dout(w_dff_A_fqioc4hn6_1),.din(w_dff_A_xHhtf05p2_1),.clk(gclk));
	jdff dff_A_P2v0pyPP4_1(.dout(w_dff_A_xHhtf05p2_1),.din(w_dff_A_P2v0pyPP4_1),.clk(gclk));
	jdff dff_A_VZWadwJ72_1(.dout(w_dff_A_P2v0pyPP4_1),.din(w_dff_A_VZWadwJ72_1),.clk(gclk));
	jdff dff_A_LlGqN3Mo9_1(.dout(w_dff_A_VZWadwJ72_1),.din(w_dff_A_LlGqN3Mo9_1),.clk(gclk));
	jdff dff_A_e5X4VvEw4_1(.dout(w_dff_A_LlGqN3Mo9_1),.din(w_dff_A_e5X4VvEw4_1),.clk(gclk));
	jdff dff_A_HRj135OL9_1(.dout(w_dff_A_e5X4VvEw4_1),.din(w_dff_A_HRj135OL9_1),.clk(gclk));
	jdff dff_A_uiynUS0O5_1(.dout(w_dff_A_HRj135OL9_1),.din(w_dff_A_uiynUS0O5_1),.clk(gclk));
	jdff dff_A_F0gyBVJH0_0(.dout(w_G171gat_1[0]),.din(w_dff_A_F0gyBVJH0_0),.clk(gclk));
	jdff dff_A_nxGnwvvR9_0(.dout(w_dff_A_F0gyBVJH0_0),.din(w_dff_A_nxGnwvvR9_0),.clk(gclk));
	jdff dff_A_CJvQSQl91_0(.dout(w_dff_A_nxGnwvvR9_0),.din(w_dff_A_CJvQSQl91_0),.clk(gclk));
	jdff dff_A_EWNHvqtf6_0(.dout(w_dff_A_CJvQSQl91_0),.din(w_dff_A_EWNHvqtf6_0),.clk(gclk));
	jdff dff_A_dc8ThQtv3_0(.dout(w_dff_A_EWNHvqtf6_0),.din(w_dff_A_dc8ThQtv3_0),.clk(gclk));
	jdff dff_A_zCAx90Vt7_0(.dout(w_dff_A_dc8ThQtv3_0),.din(w_dff_A_zCAx90Vt7_0),.clk(gclk));
	jdff dff_A_Srky7VtO1_0(.dout(w_dff_A_zCAx90Vt7_0),.din(w_dff_A_Srky7VtO1_0),.clk(gclk));
	jdff dff_A_38k4Dps60_0(.dout(w_dff_A_Srky7VtO1_0),.din(w_dff_A_38k4Dps60_0),.clk(gclk));
	jdff dff_A_umCUVVI01_0(.dout(w_dff_A_38k4Dps60_0),.din(w_dff_A_umCUVVI01_0),.clk(gclk));
	jdff dff_A_3KgmhgZJ7_1(.dout(w_G171gat_1[1]),.din(w_dff_A_3KgmhgZJ7_1),.clk(gclk));
	jdff dff_A_FGqvfwLq0_1(.dout(w_dff_A_3KgmhgZJ7_1),.din(w_dff_A_FGqvfwLq0_1),.clk(gclk));
	jdff dff_A_jZIaruy44_1(.dout(w_dff_A_FGqvfwLq0_1),.din(w_dff_A_jZIaruy44_1),.clk(gclk));
	jdff dff_A_6P1esCKU2_1(.dout(w_dff_A_jZIaruy44_1),.din(w_dff_A_6P1esCKU2_1),.clk(gclk));
	jdff dff_A_gXH4ucZ47_1(.dout(w_dff_A_6P1esCKU2_1),.din(w_dff_A_gXH4ucZ47_1),.clk(gclk));
	jdff dff_A_TEcjQdqf6_1(.dout(w_dff_A_gXH4ucZ47_1),.din(w_dff_A_TEcjQdqf6_1),.clk(gclk));
	jdff dff_A_N8YKFdqL5_1(.dout(w_dff_A_TEcjQdqf6_1),.din(w_dff_A_N8YKFdqL5_1),.clk(gclk));
	jdff dff_A_Ea4uFO2l8_1(.dout(w_dff_A_N8YKFdqL5_1),.din(w_dff_A_Ea4uFO2l8_1),.clk(gclk));
	jdff dff_A_bcwERkRS3_1(.dout(w_dff_A_Ea4uFO2l8_1),.din(w_dff_A_bcwERkRS3_1),.clk(gclk));
	jdff dff_B_ykPKv9fg2_1(.din(n403),.dout(w_dff_B_ykPKv9fg2_1),.clk(gclk));
	jdff dff_B_jfrwmKXx8_0(.din(n408),.dout(w_dff_B_jfrwmKXx8_0),.clk(gclk));
	jdff dff_B_aNK4sIva0_0(.din(w_dff_B_jfrwmKXx8_0),.dout(w_dff_B_aNK4sIva0_0),.clk(gclk));
	jdff dff_B_2grKY5GW2_0(.din(n406),.dout(w_dff_B_2grKY5GW2_0),.clk(gclk));
	jdff dff_B_omz9XJ0y8_0(.din(w_dff_B_2grKY5GW2_0),.dout(w_dff_B_omz9XJ0y8_0),.clk(gclk));
	jdff dff_B_h0RbNmS50_0(.din(w_dff_B_omz9XJ0y8_0),.dout(w_dff_B_h0RbNmS50_0),.clk(gclk));
	jdff dff_B_wK80aSpe8_0(.din(w_dff_B_h0RbNmS50_0),.dout(w_dff_B_wK80aSpe8_0),.clk(gclk));
	jdff dff_B_dWQMcvUP9_0(.din(w_dff_B_wK80aSpe8_0),.dout(w_dff_B_dWQMcvUP9_0),.clk(gclk));
	jdff dff_B_tPrZ7pkb8_0(.din(w_dff_B_dWQMcvUP9_0),.dout(w_dff_B_tPrZ7pkb8_0),.clk(gclk));
	jdff dff_B_3eZQpfrg2_0(.din(w_dff_B_tPrZ7pkb8_0),.dout(w_dff_B_3eZQpfrg2_0),.clk(gclk));
	jdff dff_B_eJUlmpTO5_0(.din(w_dff_B_3eZQpfrg2_0),.dout(w_dff_B_eJUlmpTO5_0),.clk(gclk));
	jdff dff_B_bTXwLdX74_0(.din(w_dff_B_eJUlmpTO5_0),.dout(w_dff_B_bTXwLdX74_0),.clk(gclk));
	jdff dff_B_88IJbZFB0_0(.din(w_dff_B_bTXwLdX74_0),.dout(w_dff_B_88IJbZFB0_0),.clk(gclk));
	jdff dff_A_8Fw7Cyt83_1(.dout(w_G91gat_0[1]),.din(w_dff_A_8Fw7Cyt83_1),.clk(gclk));
	jdff dff_A_djKevLiJ2_1(.dout(w_dff_A_8Fw7Cyt83_1),.din(w_dff_A_djKevLiJ2_1),.clk(gclk));
	jdff dff_A_RXeM7CTo8_1(.dout(w_dff_A_djKevLiJ2_1),.din(w_dff_A_RXeM7CTo8_1),.clk(gclk));
	jdff dff_A_s7KWYlr42_1(.dout(w_dff_A_RXeM7CTo8_1),.din(w_dff_A_s7KWYlr42_1),.clk(gclk));
	jdff dff_A_hhccyiDD4_1(.dout(w_dff_A_s7KWYlr42_1),.din(w_dff_A_hhccyiDD4_1),.clk(gclk));
	jdff dff_A_iRg79Aqh2_1(.dout(w_dff_A_hhccyiDD4_1),.din(w_dff_A_iRg79Aqh2_1),.clk(gclk));
	jdff dff_A_DRcLU07w7_1(.dout(w_n404_0[1]),.din(w_dff_A_DRcLU07w7_1),.clk(gclk));
	jdff dff_A_61nbhmew8_1(.dout(w_dff_A_DRcLU07w7_1),.din(w_dff_A_61nbhmew8_1),.clk(gclk));
	jdff dff_A_e5ILXfQq6_1(.dout(w_dff_A_61nbhmew8_1),.din(w_dff_A_e5ILXfQq6_1),.clk(gclk));
	jdff dff_A_Dl3G6LQf0_1(.dout(w_dff_A_e5ILXfQq6_1),.din(w_dff_A_Dl3G6LQf0_1),.clk(gclk));
	jdff dff_A_dUSFqEcb6_1(.dout(w_dff_A_Dl3G6LQf0_1),.din(w_dff_A_dUSFqEcb6_1),.clk(gclk));
	jdff dff_A_b6AHIqUo2_1(.dout(w_dff_A_dUSFqEcb6_1),.din(w_dff_A_b6AHIqUo2_1),.clk(gclk));
	jdff dff_A_5VvKMCik3_1(.dout(w_dff_A_b6AHIqUo2_1),.din(w_dff_A_5VvKMCik3_1),.clk(gclk));
	jdff dff_A_rNfMDcpZ5_1(.dout(w_dff_A_5VvKMCik3_1),.din(w_dff_A_rNfMDcpZ5_1),.clk(gclk));
	jdff dff_A_XLAPQinO1_1(.dout(w_dff_A_rNfMDcpZ5_1),.din(w_dff_A_XLAPQinO1_1),.clk(gclk));
	jdff dff_A_7alIDhDI4_1(.dout(w_dff_A_XLAPQinO1_1),.din(w_dff_A_7alIDhDI4_1),.clk(gclk));
	jdff dff_A_mKDxqvHc9_1(.dout(w_dff_A_7alIDhDI4_1),.din(w_dff_A_mKDxqvHc9_1),.clk(gclk));
	jdff dff_A_uoaCAX433_1(.dout(w_dff_A_mKDxqvHc9_1),.din(w_dff_A_uoaCAX433_1),.clk(gclk));
	jdff dff_B_IWySEGWJ5_0(.din(n317),.dout(w_dff_B_IWySEGWJ5_0),.clk(gclk));
	jdff dff_B_OX3LEpD00_0(.din(n316),.dout(w_dff_B_OX3LEpD00_0),.clk(gclk));
	jdff dff_B_8Fc9rkR46_0(.din(w_dff_B_OX3LEpD00_0),.dout(w_dff_B_8Fc9rkR46_0),.clk(gclk));
	jdff dff_B_TTtzqLXh9_0(.din(w_dff_B_8Fc9rkR46_0),.dout(w_dff_B_TTtzqLXh9_0),.clk(gclk));
	jdff dff_B_1NlFHSi64_0(.din(w_dff_B_TTtzqLXh9_0),.dout(w_dff_B_1NlFHSi64_0),.clk(gclk));
	jdff dff_A_2MjEC4Z57_0(.dout(w_n306_1[0]),.din(w_dff_A_2MjEC4Z57_0),.clk(gclk));
	jdff dff_A_BNV2YFLi3_0(.dout(w_dff_A_2MjEC4Z57_0),.din(w_dff_A_BNV2YFLi3_0),.clk(gclk));
	jdff dff_A_QEAajFoc6_1(.dout(w_G165gat_0[1]),.din(w_dff_A_QEAajFoc6_1),.clk(gclk));
	jdff dff_A_Aror5NMl5_1(.dout(w_dff_A_QEAajFoc6_1),.din(w_dff_A_Aror5NMl5_1),.clk(gclk));
	jdff dff_A_EhApnEyJ6_1(.dout(w_dff_A_Aror5NMl5_1),.din(w_dff_A_EhApnEyJ6_1),.clk(gclk));
	jdff dff_A_RPlFmqo16_1(.dout(w_dff_A_EhApnEyJ6_1),.din(w_dff_A_RPlFmqo16_1),.clk(gclk));
	jdff dff_A_bT7jQvhl1_1(.dout(w_dff_A_RPlFmqo16_1),.din(w_dff_A_bT7jQvhl1_1),.clk(gclk));
	jdff dff_A_3amFmrMm6_1(.dout(w_dff_A_bT7jQvhl1_1),.din(w_dff_A_3amFmrMm6_1),.clk(gclk));
	jdff dff_A_MlTYgtO17_1(.dout(w_dff_A_3amFmrMm6_1),.din(w_dff_A_MlTYgtO17_1),.clk(gclk));
	jdff dff_A_1AgLbiWv4_1(.dout(w_dff_A_MlTYgtO17_1),.din(w_dff_A_1AgLbiWv4_1),.clk(gclk));
	jdff dff_A_k6mPRUsv1_2(.dout(w_G165gat_0[2]),.din(w_dff_A_k6mPRUsv1_2),.clk(gclk));
	jdff dff_A_WxKp6Ttt4_2(.dout(w_dff_A_k6mPRUsv1_2),.din(w_dff_A_WxKp6Ttt4_2),.clk(gclk));
	jdff dff_A_aXYBMq7V4_2(.dout(w_dff_A_WxKp6Ttt4_2),.din(w_dff_A_aXYBMq7V4_2),.clk(gclk));
	jdff dff_A_UENpWxHM5_2(.dout(w_dff_A_aXYBMq7V4_2),.din(w_dff_A_UENpWxHM5_2),.clk(gclk));
	jdff dff_A_1w0hamCF8_2(.dout(w_dff_A_UENpWxHM5_2),.din(w_dff_A_1w0hamCF8_2),.clk(gclk));
	jdff dff_A_PB6FsCxF0_2(.dout(w_dff_A_1w0hamCF8_2),.din(w_dff_A_PB6FsCxF0_2),.clk(gclk));
	jdff dff_A_1qF4CLvp5_2(.dout(w_dff_A_PB6FsCxF0_2),.din(w_dff_A_1qF4CLvp5_2),.clk(gclk));
	jdff dff_A_298pn4NC8_2(.dout(w_dff_A_1qF4CLvp5_2),.din(w_dff_A_298pn4NC8_2),.clk(gclk));
	jdff dff_A_LPDgjxLY2_2(.dout(w_dff_A_298pn4NC8_2),.din(w_dff_A_LPDgjxLY2_2),.clk(gclk));
	jdff dff_A_bJNZScVw7_2(.dout(w_dff_A_LPDgjxLY2_2),.din(w_dff_A_bJNZScVw7_2),.clk(gclk));
	jdff dff_B_JItRWBQW9_3(.din(G165gat),.dout(w_dff_B_JItRWBQW9_3),.clk(gclk));
	jdff dff_B_j3mZBrun8_1(.din(n426),.dout(w_dff_B_j3mZBrun8_1),.clk(gclk));
	jdff dff_B_SWfn3xHP0_1(.din(w_dff_B_j3mZBrun8_1),.dout(w_dff_B_SWfn3xHP0_1),.clk(gclk));
	jdff dff_B_zv0iiJYS0_1(.din(w_dff_B_SWfn3xHP0_1),.dout(w_dff_B_zv0iiJYS0_1),.clk(gclk));
	jdff dff_B_9CdR91dx3_1(.din(w_dff_B_zv0iiJYS0_1),.dout(w_dff_B_9CdR91dx3_1),.clk(gclk));
	jdff dff_B_0B2Kby3U8_1(.din(w_dff_B_9CdR91dx3_1),.dout(w_dff_B_0B2Kby3U8_1),.clk(gclk));
	jdff dff_B_quZmBvAP5_1(.din(w_dff_B_0B2Kby3U8_1),.dout(w_dff_B_quZmBvAP5_1),.clk(gclk));
	jdff dff_B_qYqgYkN95_1(.din(w_dff_B_quZmBvAP5_1),.dout(w_dff_B_qYqgYkN95_1),.clk(gclk));
	jdff dff_B_fpwSqhsz0_1(.din(w_dff_B_qYqgYkN95_1),.dout(w_dff_B_fpwSqhsz0_1),.clk(gclk));
	jdff dff_B_U0G8QVwx8_1(.din(w_dff_B_fpwSqhsz0_1),.dout(w_dff_B_U0G8QVwx8_1),.clk(gclk));
	jdff dff_B_zwOOlXSY7_1(.din(n428),.dout(w_dff_B_zwOOlXSY7_1),.clk(gclk));
	jdff dff_B_aVeVvnDx5_1(.din(n340),.dout(w_dff_B_aVeVvnDx5_1),.clk(gclk));
	jdff dff_B_50nYNajY8_1(.din(w_dff_B_aVeVvnDx5_1),.dout(w_dff_B_50nYNajY8_1),.clk(gclk));
	jdff dff_B_nQ74u1A52_1(.din(w_dff_B_50nYNajY8_1),.dout(w_dff_B_nQ74u1A52_1),.clk(gclk));
	jdff dff_B_sDVeZaKg0_1(.din(w_dff_B_nQ74u1A52_1),.dout(w_dff_B_sDVeZaKg0_1),.clk(gclk));
	jdff dff_B_z8dkGq7T6_1(.din(w_dff_B_sDVeZaKg0_1),.dout(w_dff_B_z8dkGq7T6_1),.clk(gclk));
	jdff dff_B_pndSr3IK8_1(.din(w_dff_B_z8dkGq7T6_1),.dout(w_dff_B_pndSr3IK8_1),.clk(gclk));
	jdff dff_B_FoaT62Es1_1(.din(n344),.dout(w_dff_B_FoaT62Es1_1),.clk(gclk));
	jdff dff_B_w2mCSZRx3_1(.din(w_dff_B_FoaT62Es1_1),.dout(w_dff_B_w2mCSZRx3_1),.clk(gclk));
	jdff dff_B_vYmNCp3o7_1(.din(w_dff_B_w2mCSZRx3_1),.dout(w_dff_B_vYmNCp3o7_1),.clk(gclk));
	jdff dff_B_3rD6pZGq8_1(.din(w_dff_B_vYmNCp3o7_1),.dout(w_dff_B_3rD6pZGq8_1),.clk(gclk));
	jdff dff_B_2AmrlOwa8_1(.din(w_dff_B_3rD6pZGq8_1),.dout(w_dff_B_2AmrlOwa8_1),.clk(gclk));
	jdff dff_B_jracUH0O1_0(.din(n171),.dout(w_dff_B_jracUH0O1_0),.clk(gclk));
	jdff dff_A_sPkWwMba2_1(.dout(w_G219gat_1[1]),.din(w_dff_A_sPkWwMba2_1),.clk(gclk));
	jdff dff_A_xUjB7yms6_1(.dout(w_dff_A_sPkWwMba2_1),.din(w_dff_A_xUjB7yms6_1),.clk(gclk));
	jdff dff_A_B81bi5UN8_2(.dout(w_G219gat_1[2]),.din(w_dff_A_B81bi5UN8_2),.clk(gclk));
	jdff dff_A_5Snwdjtc3_2(.dout(w_dff_A_B81bi5UN8_2),.din(w_dff_A_5Snwdjtc3_2),.clk(gclk));
	jdff dff_A_foZW5O332_2(.dout(w_dff_A_5Snwdjtc3_2),.din(w_dff_A_foZW5O332_2),.clk(gclk));
	jdff dff_A_dbuGOjr01_2(.dout(w_dff_A_foZW5O332_2),.din(w_dff_A_dbuGOjr01_2),.clk(gclk));
	jdff dff_A_BLjNfsyj6_0(.dout(w_G219gat_0[0]),.din(w_dff_A_BLjNfsyj6_0),.clk(gclk));
	jdff dff_A_gzDGlbFK2_0(.dout(w_dff_A_BLjNfsyj6_0),.din(w_dff_A_gzDGlbFK2_0),.clk(gclk));
	jdff dff_A_FJcBoJQt8_0(.dout(w_dff_A_gzDGlbFK2_0),.din(w_dff_A_FJcBoJQt8_0),.clk(gclk));
	jdff dff_A_faq1I0Ji9_0(.dout(w_dff_A_FJcBoJQt8_0),.din(w_dff_A_faq1I0Ji9_0),.clk(gclk));
	jdff dff_A_QbAPkKYA4_0(.dout(w_dff_A_faq1I0Ji9_0),.din(w_dff_A_QbAPkKYA4_0),.clk(gclk));
	jdff dff_A_6SQldnJf4_0(.dout(w_dff_A_QbAPkKYA4_0),.din(w_dff_A_6SQldnJf4_0),.clk(gclk));
	jdff dff_A_nbptmbQi5_0(.dout(w_dff_A_6SQldnJf4_0),.din(w_dff_A_nbptmbQi5_0),.clk(gclk));
	jdff dff_A_UAygJ8aK3_0(.dout(w_dff_A_nbptmbQi5_0),.din(w_dff_A_UAygJ8aK3_0),.clk(gclk));
	jdff dff_A_QDzD2JfG6_0(.dout(w_dff_A_UAygJ8aK3_0),.din(w_dff_A_QDzD2JfG6_0),.clk(gclk));
	jdff dff_A_NplqoaS60_1(.dout(w_G219gat_0[1]),.din(w_dff_A_NplqoaS60_1),.clk(gclk));
	jdff dff_B_uk05Dcmc8_3(.din(G219gat),.dout(w_dff_B_uk05Dcmc8_3),.clk(gclk));
	jdff dff_B_sLop7rVf9_3(.din(w_dff_B_uk05Dcmc8_3),.dout(w_dff_B_sLop7rVf9_3),.clk(gclk));
	jdff dff_B_ANpwJDwI1_3(.din(w_dff_B_sLop7rVf9_3),.dout(w_dff_B_ANpwJDwI1_3),.clk(gclk));
	jdff dff_B_JvU5D3g95_3(.din(w_dff_B_ANpwJDwI1_3),.dout(w_dff_B_JvU5D3g95_3),.clk(gclk));
	jdff dff_B_IIDP34hE8_3(.din(w_dff_B_JvU5D3g95_3),.dout(w_dff_B_IIDP34hE8_3),.clk(gclk));
	jdff dff_B_kERcH4e84_3(.din(w_dff_B_IIDP34hE8_3),.dout(w_dff_B_kERcH4e84_3),.clk(gclk));
	jdff dff_B_k00DyxE73_3(.din(w_dff_B_kERcH4e84_3),.dout(w_dff_B_k00DyxE73_3),.clk(gclk));
	jdff dff_B_w5mZq1nO9_3(.din(w_dff_B_k00DyxE73_3),.dout(w_dff_B_w5mZq1nO9_3),.clk(gclk));
	jdff dff_B_OPtafDMO3_3(.din(w_dff_B_w5mZq1nO9_3),.dout(w_dff_B_OPtafDMO3_3),.clk(gclk));
	jdff dff_B_Vm5QE5b82_3(.din(w_dff_B_OPtafDMO3_3),.dout(w_dff_B_Vm5QE5b82_3),.clk(gclk));
	jdff dff_B_FLjWXDwp4_3(.din(w_dff_B_Vm5QE5b82_3),.dout(w_dff_B_FLjWXDwp4_3),.clk(gclk));
	jdff dff_B_0lpOHo1W6_3(.din(w_dff_B_FLjWXDwp4_3),.dout(w_dff_B_0lpOHo1W6_3),.clk(gclk));
	jdff dff_B_sNrNHi2Z1_0(.din(n427),.dout(w_dff_B_sNrNHi2Z1_0),.clk(gclk));
	jdff dff_B_WQUWdl4E3_0(.din(w_dff_B_sNrNHi2Z1_0),.dout(w_dff_B_WQUWdl4E3_0),.clk(gclk));
	jdff dff_B_hNCpO3UZ2_0(.din(w_dff_B_WQUWdl4E3_0),.dout(w_dff_B_hNCpO3UZ2_0),.clk(gclk));
	jdff dff_B_gOkFCPuS6_0(.din(w_dff_B_hNCpO3UZ2_0),.dout(w_dff_B_gOkFCPuS6_0),.clk(gclk));
	jdff dff_B_2J2GUgQg6_0(.din(w_dff_B_gOkFCPuS6_0),.dout(w_dff_B_2J2GUgQg6_0),.clk(gclk));
	jdff dff_B_R6SoFP8o6_0(.din(w_dff_B_2J2GUgQg6_0),.dout(w_dff_B_R6SoFP8o6_0),.clk(gclk));
	jdff dff_B_KW8igGK98_0(.din(w_dff_B_R6SoFP8o6_0),.dout(w_dff_B_KW8igGK98_0),.clk(gclk));
	jdff dff_B_nsnNKdcK2_0(.din(w_dff_B_KW8igGK98_0),.dout(w_dff_B_nsnNKdcK2_0),.clk(gclk));
	jdff dff_B_8cj5bpxF6_0(.din(w_dff_B_nsnNKdcK2_0),.dout(w_dff_B_8cj5bpxF6_0),.clk(gclk));
	jdff dff_B_oqg5uijF4_1(.din(n389),.dout(w_dff_B_oqg5uijF4_1),.clk(gclk));
	jdff dff_B_5rUUiEGJ8_1(.din(w_dff_B_oqg5uijF4_1),.dout(w_dff_B_5rUUiEGJ8_1),.clk(gclk));
	jdff dff_B_mfTyZGju3_1(.din(w_dff_B_5rUUiEGJ8_1),.dout(w_dff_B_mfTyZGju3_1),.clk(gclk));
	jdff dff_B_nRbGTyVN2_1(.din(w_dff_B_mfTyZGju3_1),.dout(w_dff_B_nRbGTyVN2_1),.clk(gclk));
	jdff dff_B_Th2SJlN16_1(.din(w_dff_B_nRbGTyVN2_1),.dout(w_dff_B_Th2SJlN16_1),.clk(gclk));
	jdff dff_B_WtXRA1ld5_1(.din(w_dff_B_Th2SJlN16_1),.dout(w_dff_B_WtXRA1ld5_1),.clk(gclk));
	jdff dff_B_rstrKNJd9_1(.din(w_dff_B_WtXRA1ld5_1),.dout(w_dff_B_rstrKNJd9_1),.clk(gclk));
	jdff dff_B_WBbSlcL66_1(.din(w_dff_B_rstrKNJd9_1),.dout(w_dff_B_WBbSlcL66_1),.clk(gclk));
	jdff dff_B_P8Amf1Ii6_1(.din(n359),.dout(w_dff_B_P8Amf1Ii6_1),.clk(gclk));
	jdff dff_B_oqJwv3pa1_1(.din(w_dff_B_P8Amf1Ii6_1),.dout(w_dff_B_oqJwv3pa1_1),.clk(gclk));
	jdff dff_B_bizyuQ3c8_1(.din(w_dff_B_oqJwv3pa1_1),.dout(w_dff_B_bizyuQ3c8_1),.clk(gclk));
	jdff dff_B_vU79NiWV1_1(.din(w_dff_B_bizyuQ3c8_1),.dout(w_dff_B_vU79NiWV1_1),.clk(gclk));
	jdff dff_B_9OqRy8FR4_1(.din(w_dff_B_vU79NiWV1_1),.dout(w_dff_B_9OqRy8FR4_1),.clk(gclk));
	jdff dff_B_OS01naCz7_1(.din(w_dff_B_9OqRy8FR4_1),.dout(w_dff_B_OS01naCz7_1),.clk(gclk));
	jdff dff_B_FNU1id9n2_1(.din(w_dff_B_OS01naCz7_1),.dout(w_dff_B_FNU1id9n2_1),.clk(gclk));
	jdff dff_B_DOzp6tmT5_1(.din(n252),.dout(w_dff_B_DOzp6tmT5_1),.clk(gclk));
	jdff dff_B_eP1m1TJH8_1(.din(w_dff_B_DOzp6tmT5_1),.dout(w_dff_B_eP1m1TJH8_1),.clk(gclk));
	jdff dff_B_9xyLXn9B4_1(.din(w_dff_B_eP1m1TJH8_1),.dout(w_dff_B_9xyLXn9B4_1),.clk(gclk));
	jdff dff_B_wlKVFxMU3_1(.din(w_dff_B_9xyLXn9B4_1),.dout(w_dff_B_wlKVFxMU3_1),.clk(gclk));
	jdff dff_B_dKGR2FA92_1(.din(w_dff_B_wlKVFxMU3_1),.dout(w_dff_B_dKGR2FA92_1),.clk(gclk));
	jdff dff_B_EA1D05Qk2_1(.din(n253),.dout(w_dff_B_EA1D05Qk2_1),.clk(gclk));
	jdff dff_B_CGyvMpLi8_1(.din(w_dff_B_EA1D05Qk2_1),.dout(w_dff_B_CGyvMpLi8_1),.clk(gclk));
	jdff dff_B_OxgmYRwT3_1(.din(w_dff_B_CGyvMpLi8_1),.dout(w_dff_B_OxgmYRwT3_1),.clk(gclk));
	jdff dff_B_wSLV5KIX0_1(.din(w_dff_B_OxgmYRwT3_1),.dout(w_dff_B_wSLV5KIX0_1),.clk(gclk));
	jdff dff_B_a50DAPam4_1(.din(n254),.dout(w_dff_B_a50DAPam4_1),.clk(gclk));
	jdff dff_B_F7IlVEb42_1(.din(w_dff_B_a50DAPam4_1),.dout(w_dff_B_F7IlVEb42_1),.clk(gclk));
	jdff dff_B_Zzo3shUD6_1(.din(w_dff_B_F7IlVEb42_1),.dout(w_dff_B_Zzo3shUD6_1),.clk(gclk));
	jdff dff_B_rpB8y5Sp7_1(.din(n255),.dout(w_dff_B_rpB8y5Sp7_1),.clk(gclk));
	jdff dff_B_LzIDozHE7_1(.din(w_dff_B_rpB8y5Sp7_1),.dout(w_dff_B_LzIDozHE7_1),.clk(gclk));
	jdff dff_A_OMBCyLHr2_1(.dout(w_n209_0[1]),.din(w_dff_A_OMBCyLHr2_1),.clk(gclk));
	jdff dff_B_bi6WFPIu5_2(.din(n209),.dout(w_dff_B_bi6WFPIu5_2),.clk(gclk));
	jdff dff_B_8IudweDH8_2(.din(w_dff_B_bi6WFPIu5_2),.dout(w_dff_B_8IudweDH8_2),.clk(gclk));
	jdff dff_B_Sb1PajTg8_2(.din(w_dff_B_8IudweDH8_2),.dout(w_dff_B_Sb1PajTg8_2),.clk(gclk));
	jdff dff_B_TkSNEB3m5_2(.din(w_dff_B_Sb1PajTg8_2),.dout(w_dff_B_TkSNEB3m5_2),.clk(gclk));
	jdff dff_B_mxpB1oQ99_2(.din(w_dff_B_TkSNEB3m5_2),.dout(w_dff_B_mxpB1oQ99_2),.clk(gclk));
	jdff dff_B_2wF5YYm92_2(.din(w_dff_B_mxpB1oQ99_2),.dout(w_dff_B_2wF5YYm92_2),.clk(gclk));
	jdff dff_B_gY9tg5BZ1_2(.din(w_dff_B_2wF5YYm92_2),.dout(w_dff_B_gY9tg5BZ1_2),.clk(gclk));
	jdff dff_B_MY5bGOmQ9_2(.din(w_dff_B_gY9tg5BZ1_2),.dout(w_dff_B_MY5bGOmQ9_2),.clk(gclk));
	jdff dff_B_m4CVuFCK4_2(.din(w_dff_B_MY5bGOmQ9_2),.dout(w_dff_B_m4CVuFCK4_2),.clk(gclk));
	jdff dff_A_OSv6XK8A7_0(.dout(w_G261gat_0[0]),.din(w_dff_A_OSv6XK8A7_0),.clk(gclk));
	jdff dff_A_NWo7Y8IW9_0(.dout(w_dff_A_OSv6XK8A7_0),.din(w_dff_A_NWo7Y8IW9_0),.clk(gclk));
	jdff dff_A_BKBe6dXk9_0(.dout(w_dff_A_NWo7Y8IW9_0),.din(w_dff_A_BKBe6dXk9_0),.clk(gclk));
	jdff dff_A_lS9CqEuB1_0(.dout(w_dff_A_BKBe6dXk9_0),.din(w_dff_A_lS9CqEuB1_0),.clk(gclk));
	jdff dff_A_TLkUr34r9_0(.dout(w_dff_A_lS9CqEuB1_0),.din(w_dff_A_TLkUr34r9_0),.clk(gclk));
	jdff dff_A_QBERo3H81_0(.dout(w_dff_A_TLkUr34r9_0),.din(w_dff_A_QBERo3H81_0),.clk(gclk));
	jdff dff_A_uXqbUymm0_0(.dout(w_dff_A_QBERo3H81_0),.din(w_dff_A_uXqbUymm0_0),.clk(gclk));
	jdff dff_A_6aJZEYCH1_0(.dout(w_dff_A_uXqbUymm0_0),.din(w_dff_A_6aJZEYCH1_0),.clk(gclk));
	jdff dff_A_ZDsl5Lcn6_0(.dout(w_dff_A_6aJZEYCH1_0),.din(w_dff_A_ZDsl5Lcn6_0),.clk(gclk));
	jdff dff_A_eW8E8Ysa1_0(.dout(w_dff_A_ZDsl5Lcn6_0),.din(w_dff_A_eW8E8Ysa1_0),.clk(gclk));
	jdff dff_A_gvvmMb2i6_2(.dout(w_G261gat_0[2]),.din(w_dff_A_gvvmMb2i6_2),.clk(gclk));
	jdff dff_A_nXia7lYJ7_2(.dout(w_dff_A_gvvmMb2i6_2),.din(w_dff_A_nXia7lYJ7_2),.clk(gclk));
	jdff dff_A_jr6JBQgN5_2(.dout(w_dff_A_nXia7lYJ7_2),.din(w_dff_A_jr6JBQgN5_2),.clk(gclk));
	jdff dff_A_wC8V2YAR2_2(.dout(w_dff_A_jr6JBQgN5_2),.din(w_dff_A_wC8V2YAR2_2),.clk(gclk));
	jdff dff_A_5XdvEl584_2(.dout(w_dff_A_wC8V2YAR2_2),.din(w_dff_A_5XdvEl584_2),.clk(gclk));
	jdff dff_A_9D3OSMVh9_2(.dout(w_dff_A_5XdvEl584_2),.din(w_dff_A_9D3OSMVh9_2),.clk(gclk));
	jdff dff_A_Ftvykmck4_2(.dout(w_dff_A_9D3OSMVh9_2),.din(w_dff_A_Ftvykmck4_2),.clk(gclk));
	jdff dff_A_mCwaDtVM6_2(.dout(w_dff_A_Ftvykmck4_2),.din(w_dff_A_mCwaDtVM6_2),.clk(gclk));
	jdff dff_A_WXlMYB3o1_2(.dout(w_dff_A_mCwaDtVM6_2),.din(w_dff_A_WXlMYB3o1_2),.clk(gclk));
	jdff dff_A_4uGeR0Mo1_2(.dout(w_dff_A_WXlMYB3o1_2),.din(w_dff_A_4uGeR0Mo1_2),.clk(gclk));
	jdff dff_A_qtE1DAht0_0(.dout(w_n242_0[0]),.din(w_dff_A_qtE1DAht0_0),.clk(gclk));
	jdff dff_B_qXTKOI5C0_1(.din(n182),.dout(w_dff_B_qXTKOI5C0_1),.clk(gclk));
	jdff dff_B_2cxF5EFe8_1(.din(n191),.dout(w_dff_B_2cxF5EFe8_1),.clk(gclk));
	jdff dff_B_2D3NmVGD1_1(.din(w_dff_B_2cxF5EFe8_1),.dout(w_dff_B_2D3NmVGD1_1),.clk(gclk));
	jdff dff_B_khQssahd6_1(.din(w_dff_B_2D3NmVGD1_1),.dout(w_dff_B_khQssahd6_1),.clk(gclk));
	jdff dff_B_SVHRydft8_1(.din(w_dff_B_khQssahd6_1),.dout(w_dff_B_SVHRydft8_1),.clk(gclk));
	jdff dff_B_2ZMWjlJC5_1(.din(w_dff_B_SVHRydft8_1),.dout(w_dff_B_2ZMWjlJC5_1),.clk(gclk));
	jdff dff_B_ewqprN978_1(.din(n183),.dout(w_dff_B_ewqprN978_1),.clk(gclk));
	jdff dff_B_Q0Knbh0l8_1(.din(w_dff_B_ewqprN978_1),.dout(w_dff_B_Q0Knbh0l8_1),.clk(gclk));
	jdff dff_B_88ohiOGL1_1(.din(w_dff_B_Q0Knbh0l8_1),.dout(w_dff_B_88ohiOGL1_1),.clk(gclk));
	jdff dff_B_ZzQs6d4t2_1(.din(w_dff_B_88ohiOGL1_1),.dout(w_dff_B_ZzQs6d4t2_1),.clk(gclk));
	jdff dff_B_ArAGjGG74_1(.din(w_dff_B_ZzQs6d4t2_1),.dout(w_dff_B_ArAGjGG74_1),.clk(gclk));
	jdff dff_B_5qfs6eGb0_1(.din(n184),.dout(w_dff_B_5qfs6eGb0_1),.clk(gclk));
	jdff dff_A_Xle9Dmgz2_1(.dout(w_G126gat_0[1]),.din(w_dff_A_Xle9Dmgz2_1),.clk(gclk));
	jdff dff_A_z4XKVlhK2_1(.dout(w_dff_A_Xle9Dmgz2_1),.din(w_dff_A_z4XKVlhK2_1),.clk(gclk));
	jdff dff_A_jfUGE5tT0_1(.dout(w_dff_A_z4XKVlhK2_1),.din(w_dff_A_jfUGE5tT0_1),.clk(gclk));
	jdff dff_A_PFPzP88J5_1(.dout(w_dff_A_jfUGE5tT0_1),.din(w_dff_A_PFPzP88J5_1),.clk(gclk));
	jdff dff_A_MDG70IGx8_1(.dout(w_dff_A_PFPzP88J5_1),.din(w_dff_A_MDG70IGx8_1),.clk(gclk));
	jdff dff_A_pRUoTZao7_1(.dout(w_dff_A_MDG70IGx8_1),.din(w_dff_A_pRUoTZao7_1),.clk(gclk));
	jdff dff_B_bPaiuNPW7_3(.din(n181),.dout(w_dff_B_bPaiuNPW7_3),.clk(gclk));
	jdff dff_B_JfWnVgFu5_3(.din(w_dff_B_bPaiuNPW7_3),.dout(w_dff_B_JfWnVgFu5_3),.clk(gclk));
	jdff dff_B_Y9XE2ZZg8_3(.din(w_dff_B_JfWnVgFu5_3),.dout(w_dff_B_Y9XE2ZZg8_3),.clk(gclk));
	jdff dff_B_KGvslmRa9_3(.din(w_dff_B_Y9XE2ZZg8_3),.dout(w_dff_B_KGvslmRa9_3),.clk(gclk));
	jdff dff_B_r3Df2uqj6_3(.din(w_dff_B_KGvslmRa9_3),.dout(w_dff_B_r3Df2uqj6_3),.clk(gclk));
	jdff dff_B_7xvuNP4j7_3(.din(w_dff_B_r3Df2uqj6_3),.dout(w_dff_B_7xvuNP4j7_3),.clk(gclk));
	jdff dff_B_5V7Qa8fd0_3(.din(w_dff_B_7xvuNP4j7_3),.dout(w_dff_B_5V7Qa8fd0_3),.clk(gclk));
	jdff dff_B_OITevaWi2_3(.din(w_dff_B_5V7Qa8fd0_3),.dout(w_dff_B_OITevaWi2_3),.clk(gclk));
	jdff dff_A_zfivgzQD7_1(.dout(w_G201gat_0[1]),.din(w_dff_A_zfivgzQD7_1),.clk(gclk));
	jdff dff_A_xpW9u7715_1(.dout(w_dff_A_zfivgzQD7_1),.din(w_dff_A_xpW9u7715_1),.clk(gclk));
	jdff dff_A_OJsL894y4_1(.dout(w_dff_A_xpW9u7715_1),.din(w_dff_A_OJsL894y4_1),.clk(gclk));
	jdff dff_A_ZvFnALLa1_1(.dout(w_dff_A_OJsL894y4_1),.din(w_dff_A_ZvFnALLa1_1),.clk(gclk));
	jdff dff_A_uvvfuUbd9_1(.dout(w_dff_A_ZvFnALLa1_1),.din(w_dff_A_uvvfuUbd9_1),.clk(gclk));
	jdff dff_A_wuKu8Twq6_1(.dout(w_dff_A_uvvfuUbd9_1),.din(w_dff_A_wuKu8Twq6_1),.clk(gclk));
	jdff dff_A_VR0JYUqs3_1(.dout(w_dff_A_wuKu8Twq6_1),.din(w_dff_A_VR0JYUqs3_1),.clk(gclk));
	jdff dff_A_zFw44dvQ9_1(.dout(w_dff_A_VR0JYUqs3_1),.din(w_dff_A_zFw44dvQ9_1),.clk(gclk));
	jdff dff_A_9fbgEdg66_1(.dout(w_dff_A_zFw44dvQ9_1),.din(w_dff_A_9fbgEdg66_1),.clk(gclk));
	jdff dff_A_z4qfyLAF0_1(.dout(w_n241_0[1]),.din(w_dff_A_z4qfyLAF0_1),.clk(gclk));
	jdff dff_A_nEbG1Hc63_1(.dout(w_dff_A_z4qfyLAF0_1),.din(w_dff_A_nEbG1Hc63_1),.clk(gclk));
	jdff dff_A_TPrcG7s28_1(.dout(w_dff_A_nEbG1Hc63_1),.din(w_dff_A_TPrcG7s28_1),.clk(gclk));
	jdff dff_A_1m2tPiys5_1(.dout(w_G195gat_1[1]),.din(w_dff_A_1m2tPiys5_1),.clk(gclk));
	jdff dff_A_QQetPoYP3_1(.dout(w_dff_A_1m2tPiys5_1),.din(w_dff_A_QQetPoYP3_1),.clk(gclk));
	jdff dff_A_G9UY5Wjl4_1(.dout(w_dff_A_QQetPoYP3_1),.din(w_dff_A_G9UY5Wjl4_1),.clk(gclk));
	jdff dff_A_QWdUFinA3_1(.dout(w_dff_A_G9UY5Wjl4_1),.din(w_dff_A_QWdUFinA3_1),.clk(gclk));
	jdff dff_A_44uvJDc92_1(.dout(w_dff_A_QWdUFinA3_1),.din(w_dff_A_44uvJDc92_1),.clk(gclk));
	jdff dff_A_5nr9JNoN4_1(.dout(w_dff_A_44uvJDc92_1),.din(w_dff_A_5nr9JNoN4_1),.clk(gclk));
	jdff dff_A_YaQ6DfTj4_1(.dout(w_dff_A_5nr9JNoN4_1),.din(w_dff_A_YaQ6DfTj4_1),.clk(gclk));
	jdff dff_A_8FFtGJvN1_1(.dout(w_dff_A_YaQ6DfTj4_1),.din(w_dff_A_8FFtGJvN1_1),.clk(gclk));
	jdff dff_A_1b21DjhC1_2(.dout(w_G195gat_1[2]),.din(w_dff_A_1b21DjhC1_2),.clk(gclk));
	jdff dff_A_PJg3mHst9_2(.dout(w_dff_A_1b21DjhC1_2),.din(w_dff_A_PJg3mHst9_2),.clk(gclk));
	jdff dff_A_MuqMFDeA2_2(.dout(w_dff_A_PJg3mHst9_2),.din(w_dff_A_MuqMFDeA2_2),.clk(gclk));
	jdff dff_A_l7hXzU142_2(.dout(w_dff_A_MuqMFDeA2_2),.din(w_dff_A_l7hXzU142_2),.clk(gclk));
	jdff dff_A_ztQ9x2QQ4_2(.dout(w_dff_A_l7hXzU142_2),.din(w_dff_A_ztQ9x2QQ4_2),.clk(gclk));
	jdff dff_A_YoXKZITh4_2(.dout(w_dff_A_ztQ9x2QQ4_2),.din(w_dff_A_YoXKZITh4_2),.clk(gclk));
	jdff dff_A_UNHbRGcD2_2(.dout(w_dff_A_YoXKZITh4_2),.din(w_dff_A_UNHbRGcD2_2),.clk(gclk));
	jdff dff_A_T6GTcP1f5_2(.dout(w_dff_A_UNHbRGcD2_2),.din(w_dff_A_T6GTcP1f5_2),.clk(gclk));
	jdff dff_A_8a8iIFTM4_1(.dout(w_n240_0[1]),.din(w_dff_A_8a8iIFTM4_1),.clk(gclk));
	jdff dff_A_FfVdTNP35_1(.dout(w_dff_A_8a8iIFTM4_1),.din(w_dff_A_FfVdTNP35_1),.clk(gclk));
	jdff dff_A_F8EUEhhI8_1(.dout(w_dff_A_FfVdTNP35_1),.din(w_dff_A_F8EUEhhI8_1),.clk(gclk));
	jdff dff_A_KyteEw716_1(.dout(w_dff_A_F8EUEhhI8_1),.din(w_dff_A_KyteEw716_1),.clk(gclk));
	jdff dff_A_UKS2OG6w5_0(.dout(w_G121gat_0[0]),.din(w_dff_A_UKS2OG6w5_0),.clk(gclk));
	jdff dff_A_IvZc5PzL8_0(.dout(w_dff_A_UKS2OG6w5_0),.din(w_dff_A_IvZc5PzL8_0),.clk(gclk));
	jdff dff_A_uVzCD2xt2_0(.dout(w_dff_A_IvZc5PzL8_0),.din(w_dff_A_uVzCD2xt2_0),.clk(gclk));
	jdff dff_A_RHud1xLO8_0(.dout(w_dff_A_uVzCD2xt2_0),.din(w_dff_A_RHud1xLO8_0),.clk(gclk));
	jdff dff_A_pCLLzebd9_0(.dout(w_dff_A_RHud1xLO8_0),.din(w_dff_A_pCLLzebd9_0),.clk(gclk));
	jdff dff_A_dUBtC1qd6_0(.dout(w_dff_A_pCLLzebd9_0),.din(w_dff_A_dUBtC1qd6_0),.clk(gclk));
	jdff dff_A_4kgXKw3Q4_0(.dout(w_G195gat_2[0]),.din(w_dff_A_4kgXKw3Q4_0),.clk(gclk));
	jdff dff_A_8nxSezyE0_0(.dout(w_dff_A_4kgXKw3Q4_0),.din(w_dff_A_8nxSezyE0_0),.clk(gclk));
	jdff dff_A_bdxg8klS9_0(.dout(w_dff_A_8nxSezyE0_0),.din(w_dff_A_bdxg8klS9_0),.clk(gclk));
	jdff dff_A_Dtk9iih96_0(.dout(w_dff_A_bdxg8klS9_0),.din(w_dff_A_Dtk9iih96_0),.clk(gclk));
	jdff dff_A_xnniHpW95_0(.dout(w_dff_A_Dtk9iih96_0),.din(w_dff_A_xnniHpW95_0),.clk(gclk));
	jdff dff_A_3jlUaKb16_0(.dout(w_dff_A_xnniHpW95_0),.din(w_dff_A_3jlUaKb16_0),.clk(gclk));
	jdff dff_A_qldccWpz1_0(.dout(w_dff_A_3jlUaKb16_0),.din(w_dff_A_qldccWpz1_0),.clk(gclk));
	jdff dff_A_va40lpK76_0(.dout(w_dff_A_qldccWpz1_0),.din(w_dff_A_va40lpK76_0),.clk(gclk));
	jdff dff_A_paX5FpD35_2(.dout(w_G195gat_0[2]),.din(w_dff_A_paX5FpD35_2),.clk(gclk));
	jdff dff_A_83v3Ptnb2_2(.dout(w_dff_A_paX5FpD35_2),.din(w_dff_A_83v3Ptnb2_2),.clk(gclk));
	jdff dff_A_066jas2T6_2(.dout(w_dff_A_83v3Ptnb2_2),.din(w_dff_A_066jas2T6_2),.clk(gclk));
	jdff dff_A_INSPVGEJ9_2(.dout(w_dff_A_066jas2T6_2),.din(w_dff_A_INSPVGEJ9_2),.clk(gclk));
	jdff dff_A_hT3JGetU5_1(.dout(w_n235_0[1]),.din(w_dff_A_hT3JGetU5_1),.clk(gclk));
	jdff dff_A_oUvkHlAV4_1(.dout(w_dff_A_hT3JGetU5_1),.din(w_dff_A_oUvkHlAV4_1),.clk(gclk));
	jdff dff_A_GFdWze8v3_1(.dout(w_dff_A_oUvkHlAV4_1),.din(w_dff_A_GFdWze8v3_1),.clk(gclk));
	jdff dff_A_q9ZKECyl4_1(.dout(w_dff_A_GFdWze8v3_1),.din(w_dff_A_q9ZKECyl4_1),.clk(gclk));
	jdff dff_A_vkKBmERZ0_1(.dout(w_dff_A_q9ZKECyl4_1),.din(w_dff_A_vkKBmERZ0_1),.clk(gclk));
	jdff dff_A_x0CfwG637_1(.dout(w_G189gat_1[1]),.din(w_dff_A_x0CfwG637_1),.clk(gclk));
	jdff dff_A_mGyWlh4m6_1(.dout(w_dff_A_x0CfwG637_1),.din(w_dff_A_mGyWlh4m6_1),.clk(gclk));
	jdff dff_A_J9YVKSMT2_1(.dout(w_dff_A_mGyWlh4m6_1),.din(w_dff_A_J9YVKSMT2_1),.clk(gclk));
	jdff dff_A_TE1LYzJ55_1(.dout(w_dff_A_J9YVKSMT2_1),.din(w_dff_A_TE1LYzJ55_1),.clk(gclk));
	jdff dff_A_NROoXcQx5_1(.dout(w_dff_A_TE1LYzJ55_1),.din(w_dff_A_NROoXcQx5_1),.clk(gclk));
	jdff dff_A_8SHpV8Nt2_1(.dout(w_dff_A_NROoXcQx5_1),.din(w_dff_A_8SHpV8Nt2_1),.clk(gclk));
	jdff dff_A_Nh81YyjX3_1(.dout(w_dff_A_8SHpV8Nt2_1),.din(w_dff_A_Nh81YyjX3_1),.clk(gclk));
	jdff dff_A_sUwDPp9l2_1(.dout(w_dff_A_Nh81YyjX3_1),.din(w_dff_A_sUwDPp9l2_1),.clk(gclk));
	jdff dff_A_GhiR5F3t9_2(.dout(w_G189gat_1[2]),.din(w_dff_A_GhiR5F3t9_2),.clk(gclk));
	jdff dff_A_MFHuu97o5_2(.dout(w_dff_A_GhiR5F3t9_2),.din(w_dff_A_MFHuu97o5_2),.clk(gclk));
	jdff dff_A_0EOctvqZ9_2(.dout(w_dff_A_MFHuu97o5_2),.din(w_dff_A_0EOctvqZ9_2),.clk(gclk));
	jdff dff_A_306pFsMo8_2(.dout(w_dff_A_0EOctvqZ9_2),.din(w_dff_A_306pFsMo8_2),.clk(gclk));
	jdff dff_A_Ak6kEMNY0_2(.dout(w_dff_A_306pFsMo8_2),.din(w_dff_A_Ak6kEMNY0_2),.clk(gclk));
	jdff dff_A_I3HcGDLJ5_2(.dout(w_dff_A_Ak6kEMNY0_2),.din(w_dff_A_I3HcGDLJ5_2),.clk(gclk));
	jdff dff_A_0DpHexeU4_2(.dout(w_dff_A_I3HcGDLJ5_2),.din(w_dff_A_0DpHexeU4_2),.clk(gclk));
	jdff dff_A_Ht5CjNyr0_2(.dout(w_dff_A_0DpHexeU4_2),.din(w_dff_A_Ht5CjNyr0_2),.clk(gclk));
	jdff dff_A_zAfpDSX87_1(.dout(w_n234_0[1]),.din(w_dff_A_zAfpDSX87_1),.clk(gclk));
	jdff dff_A_cOcRJlFR6_1(.dout(w_dff_A_zAfpDSX87_1),.din(w_dff_A_cOcRJlFR6_1),.clk(gclk));
	jdff dff_A_o6lfSWg87_1(.dout(w_dff_A_cOcRJlFR6_1),.din(w_dff_A_o6lfSWg87_1),.clk(gclk));
	jdff dff_A_voUozTFw6_1(.dout(w_dff_A_o6lfSWg87_1),.din(w_dff_A_voUozTFw6_1),.clk(gclk));
	jdff dff_A_rsFIe1aH5_1(.dout(w_dff_A_voUozTFw6_1),.din(w_dff_A_rsFIe1aH5_1),.clk(gclk));
	jdff dff_A_p9nyq2QR8_1(.dout(w_dff_A_rsFIe1aH5_1),.din(w_dff_A_p9nyq2QR8_1),.clk(gclk));
	jdff dff_A_itxIFKPu8_1(.dout(w_G146gat_0[1]),.din(w_dff_A_itxIFKPu8_1),.clk(gclk));
	jdff dff_B_D0vffpct1_2(.din(G146gat),.dout(w_dff_B_D0vffpct1_2),.clk(gclk));
	jdff dff_B_mIIJ43376_2(.din(w_dff_B_D0vffpct1_2),.dout(w_dff_B_mIIJ43376_2),.clk(gclk));
	jdff dff_B_yyJouFsP9_2(.din(w_dff_B_mIIJ43376_2),.dout(w_dff_B_yyJouFsP9_2),.clk(gclk));
	jdff dff_B_y1SzNhuL3_2(.din(w_dff_B_yyJouFsP9_2),.dout(w_dff_B_y1SzNhuL3_2),.clk(gclk));
	jdff dff_A_RNBdg8Ms9_1(.dout(w_G116gat_0[1]),.din(w_dff_A_RNBdg8Ms9_1),.clk(gclk));
	jdff dff_A_rClJEoJn2_1(.dout(w_dff_A_RNBdg8Ms9_1),.din(w_dff_A_rClJEoJn2_1),.clk(gclk));
	jdff dff_A_NgCqrEpS2_1(.dout(w_dff_A_rClJEoJn2_1),.din(w_dff_A_NgCqrEpS2_1),.clk(gclk));
	jdff dff_A_JNhs96JO1_1(.dout(w_dff_A_NgCqrEpS2_1),.din(w_dff_A_JNhs96JO1_1),.clk(gclk));
	jdff dff_A_xn0pxsVC0_1(.dout(w_dff_A_JNhs96JO1_1),.din(w_dff_A_xn0pxsVC0_1),.clk(gclk));
	jdff dff_A_6ylewrAP0_1(.dout(w_dff_A_xn0pxsVC0_1),.din(w_dff_A_6ylewrAP0_1),.clk(gclk));
	jdff dff_A_exW2EZWI8_0(.dout(w_G189gat_2[0]),.din(w_dff_A_exW2EZWI8_0),.clk(gclk));
	jdff dff_A_L2KCFRc49_0(.dout(w_dff_A_exW2EZWI8_0),.din(w_dff_A_L2KCFRc49_0),.clk(gclk));
	jdff dff_A_ju2QhJQJ5_0(.dout(w_dff_A_L2KCFRc49_0),.din(w_dff_A_ju2QhJQJ5_0),.clk(gclk));
	jdff dff_A_RATGlef17_0(.dout(w_dff_A_ju2QhJQJ5_0),.din(w_dff_A_RATGlef17_0),.clk(gclk));
	jdff dff_A_sV33Isf88_0(.dout(w_dff_A_RATGlef17_0),.din(w_dff_A_sV33Isf88_0),.clk(gclk));
	jdff dff_A_wC9MZx0i8_0(.dout(w_dff_A_sV33Isf88_0),.din(w_dff_A_wC9MZx0i8_0),.clk(gclk));
	jdff dff_A_20GTuGzz7_0(.dout(w_dff_A_wC9MZx0i8_0),.din(w_dff_A_20GTuGzz7_0),.clk(gclk));
	jdff dff_A_bb2z6G8Z2_0(.dout(w_dff_A_20GTuGzz7_0),.din(w_dff_A_bb2z6G8Z2_0),.clk(gclk));
	jdff dff_A_P1CXzswa6_2(.dout(w_G189gat_0[2]),.din(w_dff_A_P1CXzswa6_2),.clk(gclk));
	jdff dff_A_yJ1wKhIb6_2(.dout(w_dff_A_P1CXzswa6_2),.din(w_dff_A_yJ1wKhIb6_2),.clk(gclk));
	jdff dff_A_fSYQQfb87_2(.dout(w_dff_A_yJ1wKhIb6_2),.din(w_dff_A_fSYQQfb87_2),.clk(gclk));
	jdff dff_A_zjT6Xz1q5_2(.dout(w_dff_A_fSYQQfb87_2),.din(w_dff_A_zjT6Xz1q5_2),.clk(gclk));
	jdff dff_A_im0Atm1c4_0(.dout(w_n343_0[0]),.din(w_dff_A_im0Atm1c4_0),.clk(gclk));
	jdff dff_A_XaOxr14T7_0(.dout(w_dff_A_im0Atm1c4_0),.din(w_dff_A_XaOxr14T7_0),.clk(gclk));
	jdff dff_A_lusLN7lH4_0(.dout(w_dff_A_XaOxr14T7_0),.din(w_dff_A_lusLN7lH4_0),.clk(gclk));
	jdff dff_A_ljsR9KFd9_0(.dout(w_dff_A_lusLN7lH4_0),.din(w_dff_A_ljsR9KFd9_0),.clk(gclk));
	jdff dff_A_NLs4hC7u2_0(.dout(w_dff_A_ljsR9KFd9_0),.din(w_dff_A_NLs4hC7u2_0),.clk(gclk));
	jdff dff_A_n6gYM2im1_0(.dout(w_dff_A_NLs4hC7u2_0),.din(w_dff_A_n6gYM2im1_0),.clk(gclk));
	jdff dff_B_9uarQ1Is4_1(.din(n341),.dout(w_dff_B_9uarQ1Is4_1),.clk(gclk));
	jdff dff_B_3qBlOM3f6_1(.din(w_dff_B_9uarQ1Is4_1),.dout(w_dff_B_3qBlOM3f6_1),.clk(gclk));
	jdff dff_B_nU0ZGq4l6_1(.din(w_dff_B_3qBlOM3f6_1),.dout(w_dff_B_nU0ZGq4l6_1),.clk(gclk));
	jdff dff_B_d9HnqHjg6_1(.din(w_dff_B_nU0ZGq4l6_1),.dout(w_dff_B_d9HnqHjg6_1),.clk(gclk));
	jdff dff_B_Sea4Laxb4_1(.din(w_dff_B_d9HnqHjg6_1),.dout(w_dff_B_Sea4Laxb4_1),.clk(gclk));
	jdff dff_B_HDMLwBiH1_1(.din(w_dff_B_Sea4Laxb4_1),.dout(w_dff_B_HDMLwBiH1_1),.clk(gclk));
	jdff dff_B_WSpepJWM5_1(.din(w_dff_B_HDMLwBiH1_1),.dout(w_dff_B_WSpepJWM5_1),.clk(gclk));
	jdff dff_B_7c8zefUi4_1(.din(w_dff_B_WSpepJWM5_1),.dout(w_dff_B_7c8zefUi4_1),.clk(gclk));
	jdff dff_A_1276Se0U6_1(.dout(w_n222_0[1]),.din(w_dff_A_1276Se0U6_1),.clk(gclk));
	jdff dff_A_UvhdSvIW7_1(.dout(w_dff_A_1276Se0U6_1),.din(w_dff_A_UvhdSvIW7_1),.clk(gclk));
	jdff dff_A_A0sc5vW81_1(.dout(w_dff_A_UvhdSvIW7_1),.din(w_dff_A_A0sc5vW81_1),.clk(gclk));
	jdff dff_A_N6wcWuk02_1(.dout(w_dff_A_A0sc5vW81_1),.din(w_dff_A_N6wcWuk02_1),.clk(gclk));
	jdff dff_A_qOyCYc875_1(.dout(w_dff_A_N6wcWuk02_1),.din(w_dff_A_qOyCYc875_1),.clk(gclk));
	jdff dff_A_eN5PGpMF1_1(.dout(w_dff_A_qOyCYc875_1),.din(w_dff_A_eN5PGpMF1_1),.clk(gclk));
	jdff dff_A_0C0f06Tg1_1(.dout(w_dff_A_eN5PGpMF1_1),.din(w_dff_A_0C0f06Tg1_1),.clk(gclk));
	jdff dff_A_dVLCxt2u1_1(.dout(w_dff_A_0C0f06Tg1_1),.din(w_dff_A_dVLCxt2u1_1),.clk(gclk));
	jdff dff_A_WTQitkku9_0(.dout(w_n97_0[0]),.din(w_dff_A_WTQitkku9_0),.clk(gclk));
	jdff dff_A_KZy4AgKK7_0(.dout(w_dff_A_WTQitkku9_0),.din(w_dff_A_KZy4AgKK7_0),.clk(gclk));
	jdff dff_A_RGUelmQ76_0(.dout(w_dff_A_KZy4AgKK7_0),.din(w_dff_A_RGUelmQ76_0),.clk(gclk));
	jdff dff_A_9XrtnsfL1_1(.dout(w_G143gat_0[1]),.din(w_dff_A_9XrtnsfL1_1),.clk(gclk));
	jdff dff_B_PbmYmigO7_2(.din(G143gat),.dout(w_dff_B_PbmYmigO7_2),.clk(gclk));
	jdff dff_B_LN0jDN862_2(.din(w_dff_B_PbmYmigO7_2),.dout(w_dff_B_LN0jDN862_2),.clk(gclk));
	jdff dff_B_NQ3Az6R77_2(.din(w_dff_B_LN0jDN862_2),.dout(w_dff_B_NQ3Az6R77_2),.clk(gclk));
	jdff dff_B_W2ds2gT87_2(.din(w_dff_B_NQ3Az6R77_2),.dout(w_dff_B_W2ds2gT87_2),.clk(gclk));
	jdff dff_A_KX4xrdus9_2(.dout(w_n148_1[2]),.din(w_dff_A_KX4xrdus9_2),.clk(gclk));
	jdff dff_A_cZ6N61VB0_2(.dout(w_dff_A_KX4xrdus9_2),.din(w_dff_A_cZ6N61VB0_2),.clk(gclk));
	jdff dff_A_9klrine08_1(.dout(w_G111gat_0[1]),.din(w_dff_A_9klrine08_1),.clk(gclk));
	jdff dff_A_BzAvCowr5_1(.dout(w_dff_A_9klrine08_1),.din(w_dff_A_BzAvCowr5_1),.clk(gclk));
	jdff dff_A_1dS8OmZd0_1(.dout(w_dff_A_BzAvCowr5_1),.din(w_dff_A_1dS8OmZd0_1),.clk(gclk));
	jdff dff_A_7XkwRaaW3_1(.dout(w_dff_A_1dS8OmZd0_1),.din(w_dff_A_7XkwRaaW3_1),.clk(gclk));
	jdff dff_A_cTxiTtCl2_1(.dout(w_dff_A_7XkwRaaW3_1),.din(w_dff_A_cTxiTtCl2_1),.clk(gclk));
	jdff dff_A_lv8FHbdM0_1(.dout(w_dff_A_cTxiTtCl2_1),.din(w_dff_A_lv8FHbdM0_1),.clk(gclk));
	jdff dff_A_OlVTpwZU4_2(.dout(w_G183gat_0[2]),.din(w_dff_A_OlVTpwZU4_2),.clk(gclk));
	jdff dff_A_gDVyWr702_2(.dout(w_dff_A_OlVTpwZU4_2),.din(w_dff_A_gDVyWr702_2),.clk(gclk));
	jdff dff_A_buhkmTua3_2(.dout(w_dff_A_gDVyWr702_2),.din(w_dff_A_buhkmTua3_2),.clk(gclk));
	jdff dff_A_k9kVHTqQ3_2(.dout(w_dff_A_buhkmTua3_2),.din(w_dff_A_k9kVHTqQ3_2),.clk(gclk));
	jdff dff_A_u7tzo7zk0_2(.dout(w_dff_A_k9kVHTqQ3_2),.din(w_dff_A_u7tzo7zk0_2),.clk(gclk));
	jdff dff_A_ah55yj4e8_2(.dout(w_dff_A_u7tzo7zk0_2),.din(w_dff_A_ah55yj4e8_2),.clk(gclk));
	jdff dff_A_8bgxasnh3_2(.dout(w_dff_A_ah55yj4e8_2),.din(w_dff_A_8bgxasnh3_2),.clk(gclk));
	jdff dff_A_siOi6SOO6_2(.dout(w_dff_A_8bgxasnh3_2),.din(w_dff_A_siOi6SOO6_2),.clk(gclk));
	jdff dff_A_HNYOv0cD4_0(.dout(w_n339_0[0]),.din(w_dff_A_HNYOv0cD4_0),.clk(gclk));
	jdff dff_A_Lm7BwhMC1_0(.dout(w_dff_A_HNYOv0cD4_0),.din(w_dff_A_Lm7BwhMC1_0),.clk(gclk));
	jdff dff_A_6n5evL4g2_0(.dout(w_dff_A_Lm7BwhMC1_0),.din(w_dff_A_6n5evL4g2_0),.clk(gclk));
	jdff dff_A_sR5Q5RPH8_0(.dout(w_dff_A_6n5evL4g2_0),.din(w_dff_A_sR5Q5RPH8_0),.clk(gclk));
	jdff dff_A_qLueEBvD8_0(.dout(w_dff_A_sR5Q5RPH8_0),.din(w_dff_A_qLueEBvD8_0),.clk(gclk));
	jdff dff_A_eAF7bSiM8_0(.dout(w_dff_A_qLueEBvD8_0),.din(w_dff_A_eAF7bSiM8_0),.clk(gclk));
	jdff dff_A_5A1BFLOD0_0(.dout(w_dff_A_eAF7bSiM8_0),.din(w_dff_A_5A1BFLOD0_0),.clk(gclk));
	jdff dff_B_lnS2vrXY0_1(.din(n337),.dout(w_dff_B_lnS2vrXY0_1),.clk(gclk));
	jdff dff_B_JrDdZA3y2_1(.din(w_dff_B_lnS2vrXY0_1),.dout(w_dff_B_JrDdZA3y2_1),.clk(gclk));
	jdff dff_B_pDCYbpM12_1(.din(w_dff_B_JrDdZA3y2_1),.dout(w_dff_B_pDCYbpM12_1),.clk(gclk));
	jdff dff_B_Dc7TnKSD0_1(.din(w_dff_B_pDCYbpM12_1),.dout(w_dff_B_Dc7TnKSD0_1),.clk(gclk));
	jdff dff_B_7aBGlWGu1_1(.din(w_dff_B_Dc7TnKSD0_1),.dout(w_dff_B_7aBGlWGu1_1),.clk(gclk));
	jdff dff_B_cTxHss4A7_1(.din(w_dff_B_7aBGlWGu1_1),.dout(w_dff_B_cTxHss4A7_1),.clk(gclk));
	jdff dff_B_U7cJsRJT2_1(.din(w_dff_B_cTxHss4A7_1),.dout(w_dff_B_U7cJsRJT2_1),.clk(gclk));
	jdff dff_B_axxf9eNX1_1(.din(w_dff_B_U7cJsRJT2_1),.dout(w_dff_B_axxf9eNX1_1),.clk(gclk));
	jdff dff_B_8sAH4KSb6_1(.din(w_dff_B_axxf9eNX1_1),.dout(w_dff_B_8sAH4KSb6_1),.clk(gclk));
	jdff dff_A_6l4WfGqp4_2(.dout(w_n336_0[2]),.din(w_dff_A_6l4WfGqp4_2),.clk(gclk));
	jdff dff_A_oGHeM9ZH6_2(.dout(w_dff_A_6l4WfGqp4_2),.din(w_dff_A_oGHeM9ZH6_2),.clk(gclk));
	jdff dff_A_lMEn3ARL2_2(.dout(w_dff_A_oGHeM9ZH6_2),.din(w_dff_A_lMEn3ARL2_2),.clk(gclk));
	jdff dff_A_Sl90eJT38_2(.dout(w_dff_A_lMEn3ARL2_2),.din(w_dff_A_Sl90eJT38_2),.clk(gclk));
	jdff dff_A_sGm1VWF71_2(.dout(w_dff_A_Sl90eJT38_2),.din(w_dff_A_sGm1VWF71_2),.clk(gclk));
	jdff dff_A_8htcuhXY7_2(.dout(w_dff_A_sGm1VWF71_2),.din(w_dff_A_8htcuhXY7_2),.clk(gclk));
	jdff dff_A_y9Y7Sc8U7_2(.dout(w_dff_A_8htcuhXY7_2),.din(w_dff_A_y9Y7Sc8U7_2),.clk(gclk));
	jdff dff_A_tvP2TVC82_2(.dout(w_dff_A_y9Y7Sc8U7_2),.din(w_dff_A_tvP2TVC82_2),.clk(gclk));
	jdff dff_A_46IsRfaU5_2(.dout(w_dff_A_tvP2TVC82_2),.din(w_dff_A_46IsRfaU5_2),.clk(gclk));
	jdff dff_B_8lj84eFO9_0(.din(n333),.dout(w_dff_B_8lj84eFO9_0),.clk(gclk));
	jdff dff_B_RqulqVkV4_0(.din(n332),.dout(w_dff_B_RqulqVkV4_0),.clk(gclk));
	jdff dff_B_NkXKTgrX3_0(.din(w_dff_B_RqulqVkV4_0),.dout(w_dff_B_NkXKTgrX3_0),.clk(gclk));
	jdff dff_B_BUhoOciU0_0(.din(w_dff_B_NkXKTgrX3_0),.dout(w_dff_B_BUhoOciU0_0),.clk(gclk));
	jdff dff_B_8l7w3nKv2_0(.din(w_dff_B_BUhoOciU0_0),.dout(w_dff_B_8l7w3nKv2_0),.clk(gclk));
	jdff dff_A_HJxgksb40_0(.dout(w_G153gat_0[0]),.din(w_dff_A_HJxgksb40_0),.clk(gclk));
	jdff dff_A_OfQHsrTF6_0(.dout(w_dff_A_HJxgksb40_0),.din(w_dff_A_OfQHsrTF6_0),.clk(gclk));
	jdff dff_A_RHKRwJjA2_0(.dout(w_dff_A_OfQHsrTF6_0),.din(w_dff_A_RHKRwJjA2_0),.clk(gclk));
	jdff dff_A_8gyjgMM89_0(.dout(w_dff_A_RHKRwJjA2_0),.din(w_dff_A_8gyjgMM89_0),.clk(gclk));
	jdff dff_A_2EFgIYXW6_2(.dout(w_G153gat_0[2]),.din(w_dff_A_2EFgIYXW6_2),.clk(gclk));
	jdff dff_A_enq2Zzxs7_2(.dout(w_dff_A_2EFgIYXW6_2),.din(w_dff_A_enq2Zzxs7_2),.clk(gclk));
	jdff dff_A_9o9dBuND3_2(.dout(w_dff_A_enq2Zzxs7_2),.din(w_dff_A_9o9dBuND3_2),.clk(gclk));
	jdff dff_A_fSnEzeN89_2(.dout(w_dff_A_9o9dBuND3_2),.din(w_dff_A_fSnEzeN89_2),.clk(gclk));
	jdff dff_A_mxXocBMM9_2(.dout(w_dff_A_fSnEzeN89_2),.din(w_dff_A_mxXocBMM9_2),.clk(gclk));
	jdff dff_A_L62tc7Dd0_0(.dout(w_G106gat_0[0]),.din(w_dff_A_L62tc7Dd0_0),.clk(gclk));
	jdff dff_A_a4qT7Xu44_0(.dout(w_dff_A_L62tc7Dd0_0),.din(w_dff_A_a4qT7Xu44_0),.clk(gclk));
	jdff dff_A_1xzprc0w0_0(.dout(w_dff_A_a4qT7Xu44_0),.din(w_dff_A_1xzprc0w0_0),.clk(gclk));
	jdff dff_A_L6VAPfac5_0(.dout(w_dff_A_1xzprc0w0_0),.din(w_dff_A_L6VAPfac5_0),.clk(gclk));
	jdff dff_A_klsIOVKv9_0(.dout(w_dff_A_L6VAPfac5_0),.din(w_dff_A_klsIOVKv9_0),.clk(gclk));
	jdff dff_A_V3oXX5jK6_0(.dout(w_dff_A_klsIOVKv9_0),.din(w_dff_A_V3oXX5jK6_0),.clk(gclk));
	jdff dff_A_8VgGHXUs0_1(.dout(w_G177gat_1[1]),.din(w_dff_A_8VgGHXUs0_1),.clk(gclk));
	jdff dff_A_GbhNhxNH8_1(.dout(w_dff_A_8VgGHXUs0_1),.din(w_dff_A_GbhNhxNH8_1),.clk(gclk));
	jdff dff_A_PisMM5Bj4_1(.dout(w_dff_A_GbhNhxNH8_1),.din(w_dff_A_PisMM5Bj4_1),.clk(gclk));
	jdff dff_A_TqH7orVF0_1(.dout(w_dff_A_PisMM5Bj4_1),.din(w_dff_A_TqH7orVF0_1),.clk(gclk));
	jdff dff_A_Oz6QmTxr1_1(.dout(w_dff_A_TqH7orVF0_1),.din(w_dff_A_Oz6QmTxr1_1),.clk(gclk));
	jdff dff_A_TdVLNlCS0_1(.dout(w_dff_A_Oz6QmTxr1_1),.din(w_dff_A_TdVLNlCS0_1),.clk(gclk));
	jdff dff_A_rvSm0j1y6_1(.dout(w_dff_A_TdVLNlCS0_1),.din(w_dff_A_rvSm0j1y6_1),.clk(gclk));
	jdff dff_A_AkP1uF6n0_1(.dout(w_dff_A_rvSm0j1y6_1),.din(w_dff_A_AkP1uF6n0_1),.clk(gclk));
	jdff dff_A_Rxs8MonY8_1(.dout(w_dff_A_AkP1uF6n0_1),.din(w_dff_A_Rxs8MonY8_1),.clk(gclk));
	jdff dff_A_Vt5OnxID0_1(.dout(w_G177gat_0[1]),.din(w_dff_A_Vt5OnxID0_1),.clk(gclk));
	jdff dff_A_ILWbdHPl1_1(.dout(w_dff_A_Vt5OnxID0_1),.din(w_dff_A_ILWbdHPl1_1),.clk(gclk));
	jdff dff_A_JBxxJOJA1_1(.dout(w_dff_A_ILWbdHPl1_1),.din(w_dff_A_JBxxJOJA1_1),.clk(gclk));
	jdff dff_A_da8ugNZc1_1(.dout(w_dff_A_JBxxJOJA1_1),.din(w_dff_A_da8ugNZc1_1),.clk(gclk));
	jdff dff_A_qoIWz5a47_2(.dout(w_G177gat_0[2]),.din(w_dff_A_qoIWz5a47_2),.clk(gclk));
	jdff dff_A_q3X0KEwW9_2(.dout(w_dff_A_qoIWz5a47_2),.din(w_dff_A_q3X0KEwW9_2),.clk(gclk));
	jdff dff_A_730LaZ7j1_2(.dout(w_dff_A_q3X0KEwW9_2),.din(w_dff_A_730LaZ7j1_2),.clk(gclk));
	jdff dff_A_eY3Mqnvi9_2(.dout(w_dff_A_730LaZ7j1_2),.din(w_dff_A_eY3Mqnvi9_2),.clk(gclk));
	jdff dff_A_noMmOXyy1_2(.dout(w_dff_A_eY3Mqnvi9_2),.din(w_dff_A_noMmOXyy1_2),.clk(gclk));
	jdff dff_A_QCiMM3Yr2_2(.dout(w_dff_A_noMmOXyy1_2),.din(w_dff_A_QCiMM3Yr2_2),.clk(gclk));
	jdff dff_A_xY7Von7i7_2(.dout(w_dff_A_QCiMM3Yr2_2),.din(w_dff_A_xY7Von7i7_2),.clk(gclk));
	jdff dff_A_Twmi2ZNt9_2(.dout(w_dff_A_xY7Von7i7_2),.din(w_dff_A_Twmi2ZNt9_2),.clk(gclk));
	jdff dff_A_Mc204LWe0_2(.dout(w_dff_A_Twmi2ZNt9_2),.din(w_dff_A_Mc204LWe0_2),.clk(gclk));
	jdff dff_B_fPSD0pYd9_1(.din(n419),.dout(w_dff_B_fPSD0pYd9_1),.clk(gclk));
	jdff dff_B_DTU96SJW7_0(.din(n424),.dout(w_dff_B_DTU96SJW7_0),.clk(gclk));
	jdff dff_B_uepjOYpG2_0(.din(w_dff_B_DTU96SJW7_0),.dout(w_dff_B_uepjOYpG2_0),.clk(gclk));
	jdff dff_A_ALhd4WmP7_0(.dout(w_G246gat_0[0]),.din(w_dff_A_ALhd4WmP7_0),.clk(gclk));
	jdff dff_A_UZ8gk4Pj5_0(.dout(w_dff_A_ALhd4WmP7_0),.din(w_dff_A_UZ8gk4Pj5_0),.clk(gclk));
	jdff dff_A_MYSTLQrl9_0(.dout(w_dff_A_UZ8gk4Pj5_0),.din(w_dff_A_MYSTLQrl9_0),.clk(gclk));
	jdff dff_A_KImW2BEJ3_0(.dout(w_dff_A_MYSTLQrl9_0),.din(w_dff_A_KImW2BEJ3_0),.clk(gclk));
	jdff dff_A_XdXQYG6W9_0(.dout(w_dff_A_KImW2BEJ3_0),.din(w_dff_A_XdXQYG6W9_0),.clk(gclk));
	jdff dff_A_ZzO4hFMM8_0(.dout(w_dff_A_XdXQYG6W9_0),.din(w_dff_A_ZzO4hFMM8_0),.clk(gclk));
	jdff dff_A_aY5nKX752_0(.dout(w_dff_A_ZzO4hFMM8_0),.din(w_dff_A_aY5nKX752_0),.clk(gclk));
	jdff dff_A_fLHp83Dq1_0(.dout(w_dff_A_aY5nKX752_0),.din(w_dff_A_fLHp83Dq1_0),.clk(gclk));
	jdff dff_A_950OsaRw7_2(.dout(w_G246gat_0[2]),.din(w_dff_A_950OsaRw7_2),.clk(gclk));
	jdff dff_A_GC1gLHOV3_2(.dout(w_dff_A_950OsaRw7_2),.din(w_dff_A_GC1gLHOV3_2),.clk(gclk));
	jdff dff_A_sSuLM3c61_2(.dout(w_dff_A_GC1gLHOV3_2),.din(w_dff_A_sSuLM3c61_2),.clk(gclk));
	jdff dff_A_39Baepz57_2(.dout(w_dff_A_sSuLM3c61_2),.din(w_dff_A_39Baepz57_2),.clk(gclk));
	jdff dff_A_wyp1YpKB4_2(.dout(w_dff_A_39Baepz57_2),.din(w_dff_A_wyp1YpKB4_2),.clk(gclk));
	jdff dff_A_BXFiDA3H5_2(.dout(w_dff_A_wyp1YpKB4_2),.din(w_dff_A_BXFiDA3H5_2),.clk(gclk));
	jdff dff_A_NRrZTE351_2(.dout(w_dff_A_BXFiDA3H5_2),.din(w_dff_A_NRrZTE351_2),.clk(gclk));
	jdff dff_B_Fdz3JHdN9_3(.din(G246gat),.dout(w_dff_B_Fdz3JHdN9_3),.clk(gclk));
	jdff dff_B_zw2JVQPw8_0(.din(n422),.dout(w_dff_B_zw2JVQPw8_0),.clk(gclk));
	jdff dff_B_wGz6DyCH2_0(.din(w_dff_B_zw2JVQPw8_0),.dout(w_dff_B_wGz6DyCH2_0),.clk(gclk));
	jdff dff_B_4cD81alE6_0(.din(w_dff_B_wGz6DyCH2_0),.dout(w_dff_B_4cD81alE6_0),.clk(gclk));
	jdff dff_B_QNW1eCAA6_0(.din(w_dff_B_4cD81alE6_0),.dout(w_dff_B_QNW1eCAA6_0),.clk(gclk));
	jdff dff_B_NUzTcCaO1_0(.din(w_dff_B_QNW1eCAA6_0),.dout(w_dff_B_NUzTcCaO1_0),.clk(gclk));
	jdff dff_B_92g3k8ZW4_0(.din(w_dff_B_NUzTcCaO1_0),.dout(w_dff_B_92g3k8ZW4_0),.clk(gclk));
	jdff dff_B_YR8dbmug6_0(.din(w_dff_B_92g3k8ZW4_0),.dout(w_dff_B_YR8dbmug6_0),.clk(gclk));
	jdff dff_B_xP34Jod42_0(.din(w_dff_B_YR8dbmug6_0),.dout(w_dff_B_xP34Jod42_0),.clk(gclk));
	jdff dff_B_KDbK71tq5_0(.din(w_dff_B_xP34Jod42_0),.dout(w_dff_B_KDbK71tq5_0),.clk(gclk));
	jdff dff_B_76toLV5I0_0(.din(w_dff_B_KDbK71tq5_0),.dout(w_dff_B_76toLV5I0_0),.clk(gclk));
	jdff dff_A_SriR0mtm0_1(.dout(w_G96gat_0[1]),.din(w_dff_A_SriR0mtm0_1),.clk(gclk));
	jdff dff_A_9tXpX3St5_1(.dout(w_dff_A_SriR0mtm0_1),.din(w_dff_A_9tXpX3St5_1),.clk(gclk));
	jdff dff_A_twc62EEK4_1(.dout(w_dff_A_9tXpX3St5_1),.din(w_dff_A_twc62EEK4_1),.clk(gclk));
	jdff dff_A_NKLBGq8R1_1(.dout(w_dff_A_twc62EEK4_1),.din(w_dff_A_NKLBGq8R1_1),.clk(gclk));
	jdff dff_A_GJnujMiz2_1(.dout(w_dff_A_NKLBGq8R1_1),.din(w_dff_A_GJnujMiz2_1),.clk(gclk));
	jdff dff_A_J5WWu8vw3_1(.dout(w_dff_A_GJnujMiz2_1),.din(w_dff_A_J5WWu8vw3_1),.clk(gclk));
	jdff dff_A_XseHY1Bc0_0(.dout(w_n420_0[0]),.din(w_dff_A_XseHY1Bc0_0),.clk(gclk));
	jdff dff_A_GV7MT6a02_0(.dout(w_dff_A_XseHY1Bc0_0),.din(w_dff_A_GV7MT6a02_0),.clk(gclk));
	jdff dff_A_V3Qm89lt7_0(.dout(w_dff_A_GV7MT6a02_0),.din(w_dff_A_V3Qm89lt7_0),.clk(gclk));
	jdff dff_A_Nx2WuXS21_0(.dout(w_dff_A_V3Qm89lt7_0),.din(w_dff_A_Nx2WuXS21_0),.clk(gclk));
	jdff dff_A_4hjn560R5_0(.dout(w_dff_A_Nx2WuXS21_0),.din(w_dff_A_4hjn560R5_0),.clk(gclk));
	jdff dff_A_h00G7oYg4_0(.dout(w_dff_A_4hjn560R5_0),.din(w_dff_A_h00G7oYg4_0),.clk(gclk));
	jdff dff_A_34xTxBlh3_0(.dout(w_dff_A_h00G7oYg4_0),.din(w_dff_A_34xTxBlh3_0),.clk(gclk));
	jdff dff_A_m56LLBKI0_0(.dout(w_dff_A_34xTxBlh3_0),.din(w_dff_A_m56LLBKI0_0),.clk(gclk));
	jdff dff_A_kpnReuMh1_0(.dout(w_dff_A_m56LLBKI0_0),.din(w_dff_A_kpnReuMh1_0),.clk(gclk));
	jdff dff_A_ZnRoYSm69_0(.dout(w_dff_A_kpnReuMh1_0),.din(w_dff_A_ZnRoYSm69_0),.clk(gclk));
	jdff dff_A_OzA84GwL3_0(.dout(w_G228gat_0[0]),.din(w_dff_A_OzA84GwL3_0),.clk(gclk));
	jdff dff_B_9l6yyhOS4_3(.din(G228gat),.dout(w_dff_B_9l6yyhOS4_3),.clk(gclk));
	jdff dff_B_A4JFNNgI4_3(.din(w_dff_B_9l6yyhOS4_3),.dout(w_dff_B_A4JFNNgI4_3),.clk(gclk));
	jdff dff_B_PZsI1MeH8_3(.din(w_dff_B_A4JFNNgI4_3),.dout(w_dff_B_PZsI1MeH8_3),.clk(gclk));
	jdff dff_B_tWTJ7AHu0_3(.din(w_dff_B_PZsI1MeH8_3),.dout(w_dff_B_tWTJ7AHu0_3),.clk(gclk));
	jdff dff_B_4mQzefYm8_3(.din(w_dff_B_tWTJ7AHu0_3),.dout(w_dff_B_4mQzefYm8_3),.clk(gclk));
	jdff dff_B_MOzoEuXH0_3(.din(w_dff_B_4mQzefYm8_3),.dout(w_dff_B_MOzoEuXH0_3),.clk(gclk));
	jdff dff_B_xKtEAKwg1_3(.din(w_dff_B_MOzoEuXH0_3),.dout(w_dff_B_xKtEAKwg1_3),.clk(gclk));
	jdff dff_B_4LaYW1xw5_3(.din(w_dff_B_xKtEAKwg1_3),.dout(w_dff_B_4LaYW1xw5_3),.clk(gclk));
	jdff dff_B_KbHsGt928_3(.din(w_dff_B_4LaYW1xw5_3),.dout(w_dff_B_KbHsGt928_3),.clk(gclk));
	jdff dff_B_9o2qWziS6_0(.din(n325),.dout(w_dff_B_9o2qWziS6_0),.clk(gclk));
	jdff dff_B_tiTsG5Uz1_0(.din(n324),.dout(w_dff_B_tiTsG5Uz1_0),.clk(gclk));
	jdff dff_B_FomnhM4z3_0(.din(w_dff_B_tiTsG5Uz1_0),.dout(w_dff_B_FomnhM4z3_0),.clk(gclk));
	jdff dff_B_NpP7XHZp8_0(.din(w_dff_B_FomnhM4z3_0),.dout(w_dff_B_NpP7XHZp8_0),.clk(gclk));
	jdff dff_B_y0VubNw90_0(.din(w_dff_B_NpP7XHZp8_0),.dout(w_dff_B_y0VubNw90_0),.clk(gclk));
	jdff dff_A_sKjzEtp54_1(.dout(w_G149gat_0[1]),.din(w_dff_A_sKjzEtp54_1),.clk(gclk));
	jdff dff_B_7XqWas4T8_2(.din(G149gat),.dout(w_dff_B_7XqWas4T8_2),.clk(gclk));
	jdff dff_B_5uZwh7n95_2(.din(w_dff_B_7XqWas4T8_2),.dout(w_dff_B_5uZwh7n95_2),.clk(gclk));
	jdff dff_B_bdNmndIN0_2(.din(w_dff_B_5uZwh7n95_2),.dout(w_dff_B_bdNmndIN0_2),.clk(gclk));
	jdff dff_B_1vyeyFvv6_2(.din(w_dff_B_bdNmndIN0_2),.dout(w_dff_B_1vyeyFvv6_2),.clk(gclk));
	jdff dff_A_oSWM9JoE8_0(.dout(w_n162_0[0]),.din(w_dff_A_oSWM9JoE8_0),.clk(gclk));
	jdff dff_B_v1kqLZzI0_1(.din(n157),.dout(w_dff_B_v1kqLZzI0_1),.clk(gclk));
	jdff dff_B_5rUP3GbJ8_1(.din(n150),.dout(w_dff_B_5rUP3GbJ8_1),.clk(gclk));
	jdff dff_A_N45xjSrR7_0(.dout(w_n152_0[0]),.din(w_dff_A_N45xjSrR7_0),.clk(gclk));
	jdff dff_A_wcdBy92T7_0(.dout(w_n151_0[0]),.din(w_dff_A_wcdBy92T7_0),.clk(gclk));
	jdff dff_B_UjZgYGR24_2(.din(n151),.dout(w_dff_B_UjZgYGR24_2),.clk(gclk));
	jdff dff_A_cpCu6avO1_0(.dout(w_n149_0[0]),.din(w_dff_A_cpCu6avO1_0),.clk(gclk));
	jdff dff_A_NSZkdbwm2_0(.dout(w_dff_A_cpCu6avO1_0),.din(w_dff_A_NSZkdbwm2_0),.clk(gclk));
	jdff dff_A_0oyhkhfG6_1(.dout(w_n111_0[1]),.din(w_dff_A_0oyhkhfG6_1),.clk(gclk));
	jdff dff_A_mXyGRX4a1_0(.dout(w_G42gat_1[0]),.din(w_dff_A_mXyGRX4a1_0),.clk(gclk));
	jdff dff_A_9AvQxqe39_0(.dout(w_n95_0[0]),.din(w_dff_A_9AvQxqe39_0),.clk(gclk));
	jdff dff_A_RCCusdtM6_0(.dout(w_dff_A_9AvQxqe39_0),.din(w_dff_A_RCCusdtM6_0),.clk(gclk));
	jdff dff_A_n4EJj6SZ6_0(.dout(w_dff_A_RCCusdtM6_0),.din(w_dff_A_n4EJj6SZ6_0),.clk(gclk));
	jdff dff_A_Tu6IBioy6_2(.dout(w_n95_0[2]),.din(w_dff_A_Tu6IBioy6_2),.clk(gclk));
	jdff dff_A_xdF2g7xZ1_2(.dout(w_dff_A_Tu6IBioy6_2),.din(w_dff_A_xdF2g7xZ1_2),.clk(gclk));
	jdff dff_A_lvPQA1Dz7_2(.dout(w_G17gat_2[2]),.din(w_dff_A_lvPQA1Dz7_2),.clk(gclk));
	jdff dff_A_yTbhX3DK6_2(.dout(w_dff_A_lvPQA1Dz7_2),.din(w_dff_A_yTbhX3DK6_2),.clk(gclk));
	jdff dff_A_CmXasMQG4_1(.dout(w_G101gat_0[1]),.din(w_dff_A_CmXasMQG4_1),.clk(gclk));
	jdff dff_A_gX0bUCa55_1(.dout(w_dff_A_CmXasMQG4_1),.din(w_dff_A_gX0bUCa55_1),.clk(gclk));
	jdff dff_A_3gMeFb358_1(.dout(w_dff_A_gX0bUCa55_1),.din(w_dff_A_3gMeFb358_1),.clk(gclk));
	jdff dff_A_ktBrAn0o7_1(.dout(w_dff_A_3gMeFb358_1),.din(w_dff_A_ktBrAn0o7_1),.clk(gclk));
	jdff dff_A_04GdtLtn4_1(.dout(w_dff_A_ktBrAn0o7_1),.din(w_dff_A_04GdtLtn4_1),.clk(gclk));
	jdff dff_A_XWhEy3fA5_1(.dout(w_dff_A_04GdtLtn4_1),.din(w_dff_A_XWhEy3fA5_1),.clk(gclk));
	jdff dff_A_xWOPtsL63_1(.dout(w_n306_0[1]),.din(w_dff_A_xWOPtsL63_1),.clk(gclk));
	jdff dff_A_jwd2PVLX6_1(.dout(w_dff_A_xWOPtsL63_1),.din(w_dff_A_jwd2PVLX6_1),.clk(gclk));
	jdff dff_A_tWGjU2hY2_2(.dout(w_n306_0[2]),.din(w_dff_A_tWGjU2hY2_2),.clk(gclk));
	jdff dff_A_drFSEFik4_2(.dout(w_dff_A_tWGjU2hY2_2),.din(w_dff_A_drFSEFik4_2),.clk(gclk));
	jdff dff_A_WeDFvyBK6_2(.dout(w_G447gat_0[2]),.din(w_dff_A_WeDFvyBK6_2),.clk(gclk));
	jdff dff_A_vtFqyFjw7_1(.dout(w_G51gat_1[1]),.din(w_dff_A_vtFqyFjw7_1),.clk(gclk));
	jdff dff_A_BRHNwvHb2_0(.dout(w_G80gat_0[0]),.din(w_dff_A_BRHNwvHb2_0),.clk(gclk));
	jdff dff_A_OYyvent54_0(.dout(w_dff_A_BRHNwvHb2_0),.din(w_dff_A_OYyvent54_0),.clk(gclk));
	jdff dff_A_l1lgeYc16_2(.dout(w_G80gat_0[2]),.din(w_dff_A_l1lgeYc16_2),.clk(gclk));
	jdff dff_A_96QlWdhU9_0(.dout(w_n86_0[0]),.din(w_dff_A_96QlWdhU9_0),.clk(gclk));
	jdff dff_A_vSZJR51x1_0(.dout(w_dff_A_96QlWdhU9_0),.din(w_dff_A_vSZJR51x1_0),.clk(gclk));
	jdff dff_A_obUGa6ao4_0(.dout(w_G29gat_0[0]),.din(w_dff_A_obUGa6ao4_0),.clk(gclk));
	jdff dff_A_34mUYBoW0_0(.dout(w_dff_A_obUGa6ao4_0),.din(w_dff_A_34mUYBoW0_0),.clk(gclk));
	jdff dff_A_Fbey7Ie68_0(.dout(w_dff_A_34mUYBoW0_0),.din(w_dff_A_Fbey7Ie68_0),.clk(gclk));
	jdff dff_A_dPDWhqCa3_0(.dout(w_G17gat_1[0]),.din(w_dff_A_dPDWhqCa3_0),.clk(gclk));
	jdff dff_A_nOjcjacW6_0(.dout(w_dff_A_dPDWhqCa3_0),.din(w_dff_A_nOjcjacW6_0),.clk(gclk));
	jdff dff_A_3IrxBpCR3_0(.dout(w_dff_A_nOjcjacW6_0),.din(w_dff_A_3IrxBpCR3_0),.clk(gclk));
	jdff dff_A_0P3NhH3m6_0(.dout(w_dff_A_3IrxBpCR3_0),.din(w_dff_A_0P3NhH3m6_0),.clk(gclk));
	jdff dff_A_wflFVMgs8_1(.dout(w_G17gat_1[1]),.din(w_dff_A_wflFVMgs8_1),.clk(gclk));
	jdff dff_A_H3WSC5Cr7_1(.dout(w_dff_A_wflFVMgs8_1),.din(w_dff_A_H3WSC5Cr7_1),.clk(gclk));
	jdff dff_A_SzktELqp8_1(.dout(w_dff_A_H3WSC5Cr7_1),.din(w_dff_A_SzktELqp8_1),.clk(gclk));
	jdff dff_B_rIwknfaB5_2(.din(n144),.dout(w_dff_B_rIwknfaB5_2),.clk(gclk));
	jdff dff_B_RErpIhdZ2_2(.din(w_dff_B_rIwknfaB5_2),.dout(w_dff_B_RErpIhdZ2_2),.clk(gclk));
	jdff dff_B_lmnB0qBT2_2(.din(w_dff_B_RErpIhdZ2_2),.dout(w_dff_B_lmnB0qBT2_2),.clk(gclk));
	jdff dff_B_GpVk69285_2(.din(w_dff_B_lmnB0qBT2_2),.dout(w_dff_B_GpVk69285_2),.clk(gclk));
	jdff dff_A_r2bFMfYK2_0(.dout(w_G237gat_0[0]),.din(w_dff_A_r2bFMfYK2_0),.clk(gclk));
	jdff dff_A_L1iI4IxQ0_0(.dout(w_dff_A_r2bFMfYK2_0),.din(w_dff_A_L1iI4IxQ0_0),.clk(gclk));
	jdff dff_A_dT8BkolX6_0(.dout(w_dff_A_L1iI4IxQ0_0),.din(w_dff_A_dT8BkolX6_0),.clk(gclk));
	jdff dff_A_GaCu5nFp5_0(.dout(w_dff_A_dT8BkolX6_0),.din(w_dff_A_GaCu5nFp5_0),.clk(gclk));
	jdff dff_A_htwfXtvx6_0(.dout(w_dff_A_GaCu5nFp5_0),.din(w_dff_A_htwfXtvx6_0),.clk(gclk));
	jdff dff_A_lq4FohJn7_0(.dout(w_dff_A_htwfXtvx6_0),.din(w_dff_A_lq4FohJn7_0),.clk(gclk));
	jdff dff_A_hbdbuWOr4_0(.dout(w_dff_A_lq4FohJn7_0),.din(w_dff_A_hbdbuWOr4_0),.clk(gclk));
	jdff dff_A_7yRMoRsM6_0(.dout(w_dff_A_hbdbuWOr4_0),.din(w_dff_A_7yRMoRsM6_0),.clk(gclk));
	jdff dff_A_J5vPYbcI0_0(.dout(w_dff_A_7yRMoRsM6_0),.din(w_dff_A_J5vPYbcI0_0),.clk(gclk));
	jdff dff_A_laDFa2zu2_2(.dout(w_G237gat_0[2]),.din(w_dff_A_laDFa2zu2_2),.clk(gclk));
	jdff dff_A_9OPS5w880_2(.dout(w_dff_A_laDFa2zu2_2),.din(w_dff_A_9OPS5w880_2),.clk(gclk));
	jdff dff_A_LLc8bT972_2(.dout(w_dff_A_9OPS5w880_2),.din(w_dff_A_LLc8bT972_2),.clk(gclk));
	jdff dff_A_b1ljgJmY3_2(.dout(w_dff_A_LLc8bT972_2),.din(w_dff_A_b1ljgJmY3_2),.clk(gclk));
	jdff dff_A_nNpQaDzM0_2(.dout(w_dff_A_b1ljgJmY3_2),.din(w_dff_A_nNpQaDzM0_2),.clk(gclk));
	jdff dff_A_dB3LscY20_2(.dout(w_dff_A_nNpQaDzM0_2),.din(w_dff_A_dB3LscY20_2),.clk(gclk));
	jdff dff_A_xHp1pKxb1_2(.dout(w_dff_A_dB3LscY20_2),.din(w_dff_A_xHp1pKxb1_2),.clk(gclk));
	jdff dff_A_SjoOAylz5_2(.dout(w_dff_A_xHp1pKxb1_2),.din(w_dff_A_SjoOAylz5_2),.clk(gclk));
	jdff dff_A_PL2qUMNt7_2(.dout(w_dff_A_SjoOAylz5_2),.din(w_dff_A_PL2qUMNt7_2),.clk(gclk));
	jdff dff_A_MfkAFl0a6_0(.dout(w_n178_0[0]),.din(w_dff_A_MfkAFl0a6_0),.clk(gclk));
	jdff dff_A_Odny8Msv7_0(.dout(w_dff_A_MfkAFl0a6_0),.din(w_dff_A_Odny8Msv7_0),.clk(gclk));
	jdff dff_A_piYXRAxf0_0(.dout(w_dff_A_Odny8Msv7_0),.din(w_dff_A_piYXRAxf0_0),.clk(gclk));
	jdff dff_A_XtQmeaet3_0(.dout(w_dff_A_piYXRAxf0_0),.din(w_dff_A_XtQmeaet3_0),.clk(gclk));
	jdff dff_A_rdNs4Fft0_0(.dout(w_dff_A_XtQmeaet3_0),.din(w_dff_A_rdNs4Fft0_0),.clk(gclk));
	jdff dff_A_lkCyxoMw0_0(.dout(w_dff_A_rdNs4Fft0_0),.din(w_dff_A_lkCyxoMw0_0),.clk(gclk));
	jdff dff_B_b8ZWjFh27_0(.din(n176),.dout(w_dff_B_b8ZWjFh27_0),.clk(gclk));
	jdff dff_A_hDQvtrfi8_1(.dout(w_n122_0[1]),.din(w_dff_A_hDQvtrfi8_1),.clk(gclk));
	jdff dff_A_quODDAjE7_1(.dout(w_dff_A_hDQvtrfi8_1),.din(w_dff_A_quODDAjE7_1),.clk(gclk));
	jdff dff_A_QmySZphF4_1(.dout(w_dff_A_quODDAjE7_1),.din(w_dff_A_QmySZphF4_1),.clk(gclk));
	jdff dff_A_LroE6Vnx5_1(.dout(w_G68gat_0[1]),.din(w_dff_A_LroE6Vnx5_1),.clk(gclk));
	jdff dff_A_o9pMM5bp2_1(.dout(w_dff_A_LroE6Vnx5_1),.din(w_dff_A_o9pMM5bp2_1),.clk(gclk));
	jdff dff_A_qojV7tH43_1(.dout(w_dff_A_o9pMM5bp2_1),.din(w_dff_A_qojV7tH43_1),.clk(gclk));
	jdff dff_A_8qlIpxDT9_1(.dout(w_dff_A_qojV7tH43_1),.din(w_dff_A_8qlIpxDT9_1),.clk(gclk));
	jdff dff_A_NdxYmoco0_1(.dout(w_G42gat_0[1]),.din(w_dff_A_NdxYmoco0_1),.clk(gclk));
	jdff dff_A_WqJex0pj3_2(.dout(w_G42gat_0[2]),.din(w_dff_A_WqJex0pj3_2),.clk(gclk));
	jdff dff_A_cO8ebXUQ9_1(.dout(w_G1gat_0[1]),.din(w_dff_A_cO8ebXUQ9_1),.clk(gclk));
	jdff dff_A_wIKXo2rm0_1(.dout(w_dff_A_cO8ebXUQ9_1),.din(w_dff_A_wIKXo2rm0_1),.clk(gclk));
	jdff dff_A_bXzyRzKZ0_1(.dout(w_dff_A_wIKXo2rm0_1),.din(w_dff_A_bXzyRzKZ0_1),.clk(gclk));
	jdff dff_A_fRIkdtgf0_1(.dout(w_dff_A_bXzyRzKZ0_1),.din(w_dff_A_fRIkdtgf0_1),.clk(gclk));
	jdff dff_A_zMhrg1dP1_1(.dout(w_dff_A_fRIkdtgf0_1),.din(w_dff_A_zMhrg1dP1_1),.clk(gclk));
	jdff dff_A_4UdvMskC3_1(.dout(w_G13gat_0[1]),.din(w_dff_A_4UdvMskC3_1),.clk(gclk));
	jdff dff_A_xMdlOa8c6_0(.dout(w_G55gat_0[0]),.din(w_dff_A_xMdlOa8c6_0),.clk(gclk));
	jdff dff_A_3GW2ZMyL9_1(.dout(w_G55gat_0[1]),.din(w_dff_A_3GW2ZMyL9_1),.clk(gclk));
	jdff dff_A_xlfd0ulf6_1(.dout(w_dff_A_3GW2ZMyL9_1),.din(w_dff_A_xlfd0ulf6_1),.clk(gclk));
	jdff dff_B_NANhh2Uw2_3(.din(G55gat),.dout(w_dff_B_NANhh2Uw2_3),.clk(gclk));
	jdff dff_B_Xcmk5ta43_3(.din(w_dff_B_NANhh2Uw2_3),.dout(w_dff_B_Xcmk5ta43_3),.clk(gclk));
	jdff dff_A_kPrmW1xA7_1(.dout(w_G171gat_0[1]),.din(w_dff_A_kPrmW1xA7_1),.clk(gclk));
	jdff dff_A_QaRVHLuf2_1(.dout(w_dff_A_kPrmW1xA7_1),.din(w_dff_A_QaRVHLuf2_1),.clk(gclk));
	jdff dff_A_WL3akhXN1_1(.dout(w_dff_A_QaRVHLuf2_1),.din(w_dff_A_WL3akhXN1_1),.clk(gclk));
	jdff dff_A_Jw0iRXoy0_1(.dout(w_dff_A_WL3akhXN1_1),.din(w_dff_A_Jw0iRXoy0_1),.clk(gclk));
	jdff dff_A_6mUDeEdE6_1(.dout(w_dff_A_Jw0iRXoy0_1),.din(w_dff_A_6mUDeEdE6_1),.clk(gclk));
	jdff dff_A_FfLDhcoP8_1(.dout(w_dff_A_6mUDeEdE6_1),.din(w_dff_A_FfLDhcoP8_1),.clk(gclk));
	jdff dff_A_zuYUgyF44_1(.dout(w_dff_A_FfLDhcoP8_1),.din(w_dff_A_zuYUgyF44_1),.clk(gclk));
	jdff dff_A_wVTUoFv55_1(.dout(w_dff_A_zuYUgyF44_1),.din(w_dff_A_wVTUoFv55_1),.clk(gclk));
	jdff dff_A_mBVIAkts0_1(.dout(w_dff_A_wVTUoFv55_1),.din(w_dff_A_mBVIAkts0_1),.clk(gclk));
	jdff dff_A_CYnoMac51_2(.dout(w_G171gat_0[2]),.din(w_dff_A_CYnoMac51_2),.clk(gclk));
	jdff dff_A_fTM6ixcC6_2(.dout(w_dff_A_CYnoMac51_2),.din(w_dff_A_fTM6ixcC6_2),.clk(gclk));
	jdff dff_A_WYgSgO6b6_2(.dout(w_dff_A_fTM6ixcC6_2),.din(w_dff_A_WYgSgO6b6_2),.clk(gclk));
	jdff dff_A_pxeYE0363_2(.dout(w_dff_A_WYgSgO6b6_2),.din(w_dff_A_pxeYE0363_2),.clk(gclk));
	jdff dff_A_VdK6Yi0k4_2(.dout(w_dff_A_pxeYE0363_2),.din(w_dff_A_VdK6Yi0k4_2),.clk(gclk));
	jdff dff_A_6qrrPZvc4_2(.dout(w_dff_A_VdK6Yi0k4_2),.din(w_dff_A_6qrrPZvc4_2),.clk(gclk));
	jdff dff_A_LrqkyobM3_2(.dout(w_dff_A_6qrrPZvc4_2),.din(w_dff_A_LrqkyobM3_2),.clk(gclk));
	jdff dff_A_yJXLWBp65_2(.dout(w_dff_A_LrqkyobM3_2),.din(w_dff_A_yJXLWBp65_2),.clk(gclk));
	jdff dff_A_wLEibnnH4_2(.dout(w_dff_A_yJXLWBp65_2),.din(w_dff_A_wLEibnnH4_2),.clk(gclk));
	jdff dff_A_EUmFp00M3_2(.dout(w_dff_A_wLEibnnH4_2),.din(w_dff_A_EUmFp00M3_2),.clk(gclk));
	jdff dff_A_5SJuxCkp4_2(.dout(w_dff_A_EUmFp00M3_2),.din(w_dff_A_5SJuxCkp4_2),.clk(gclk));
	jdff dff_A_HSjTpPa27_2(.dout(w_dff_A_idGuKr9w1_0),.din(w_dff_A_HSjTpPa27_2),.clk(gclk));
	jdff dff_A_idGuKr9w1_0(.dout(w_dff_A_vg55lHw58_0),.din(w_dff_A_idGuKr9w1_0),.clk(gclk));
	jdff dff_A_vg55lHw58_0(.dout(w_dff_A_rzYNMmVB3_0),.din(w_dff_A_vg55lHw58_0),.clk(gclk));
	jdff dff_A_rzYNMmVB3_0(.dout(w_dff_A_PRplB95s9_0),.din(w_dff_A_rzYNMmVB3_0),.clk(gclk));
	jdff dff_A_PRplB95s9_0(.dout(w_dff_A_7aX1TLdR2_0),.din(w_dff_A_PRplB95s9_0),.clk(gclk));
	jdff dff_A_7aX1TLdR2_0(.dout(w_dff_A_sK38tr9E7_0),.din(w_dff_A_7aX1TLdR2_0),.clk(gclk));
	jdff dff_A_sK38tr9E7_0(.dout(w_dff_A_WyhyoSTf0_0),.din(w_dff_A_sK38tr9E7_0),.clk(gclk));
	jdff dff_A_WyhyoSTf0_0(.dout(w_dff_A_DwZrHQHc2_0),.din(w_dff_A_WyhyoSTf0_0),.clk(gclk));
	jdff dff_A_DwZrHQHc2_0(.dout(w_dff_A_mXbgThea2_0),.din(w_dff_A_DwZrHQHc2_0),.clk(gclk));
	jdff dff_A_mXbgThea2_0(.dout(w_dff_A_r0TA22Mu1_0),.din(w_dff_A_mXbgThea2_0),.clk(gclk));
	jdff dff_A_r0TA22Mu1_0(.dout(w_dff_A_NFRYoIXw7_0),.din(w_dff_A_r0TA22Mu1_0),.clk(gclk));
	jdff dff_A_NFRYoIXw7_0(.dout(w_dff_A_TbKnCqjP0_0),.din(w_dff_A_NFRYoIXw7_0),.clk(gclk));
	jdff dff_A_TbKnCqjP0_0(.dout(w_dff_A_Gol52KhP8_0),.din(w_dff_A_TbKnCqjP0_0),.clk(gclk));
	jdff dff_A_Gol52KhP8_0(.dout(w_dff_A_OzaMz4Ag7_0),.din(w_dff_A_Gol52KhP8_0),.clk(gclk));
	jdff dff_A_OzaMz4Ag7_0(.dout(w_dff_A_3EHQgUGu1_0),.din(w_dff_A_OzaMz4Ag7_0),.clk(gclk));
	jdff dff_A_3EHQgUGu1_0(.dout(w_dff_A_NUZ2tYBl2_0),.din(w_dff_A_3EHQgUGu1_0),.clk(gclk));
	jdff dff_A_NUZ2tYBl2_0(.dout(w_dff_A_Ce8vzDI03_0),.din(w_dff_A_NUZ2tYBl2_0),.clk(gclk));
	jdff dff_A_Ce8vzDI03_0(.dout(w_dff_A_tioiS3R20_0),.din(w_dff_A_Ce8vzDI03_0),.clk(gclk));
	jdff dff_A_tioiS3R20_0(.dout(w_dff_A_86xQDTQk2_0),.din(w_dff_A_tioiS3R20_0),.clk(gclk));
	jdff dff_A_86xQDTQk2_0(.dout(w_dff_A_zZ4yhI6G8_0),.din(w_dff_A_86xQDTQk2_0),.clk(gclk));
	jdff dff_A_zZ4yhI6G8_0(.dout(w_dff_A_5s27TObq3_0),.din(w_dff_A_zZ4yhI6G8_0),.clk(gclk));
	jdff dff_A_5s27TObq3_0(.dout(w_dff_A_Xp999MZh7_0),.din(w_dff_A_5s27TObq3_0),.clk(gclk));
	jdff dff_A_Xp999MZh7_0(.dout(w_dff_A_cH18MPb36_0),.din(w_dff_A_Xp999MZh7_0),.clk(gclk));
	jdff dff_A_cH18MPb36_0(.dout(w_dff_A_SGf4mYTT3_0),.din(w_dff_A_cH18MPb36_0),.clk(gclk));
	jdff dff_A_SGf4mYTT3_0(.dout(w_dff_A_Z0eio7q67_0),.din(w_dff_A_SGf4mYTT3_0),.clk(gclk));
	jdff dff_A_Z0eio7q67_0(.dout(G388gat),.din(w_dff_A_Z0eio7q67_0),.clk(gclk));
	jdff dff_A_f9jfGi1f8_2(.dout(w_dff_A_HMwz0DNp8_0),.din(w_dff_A_f9jfGi1f8_2),.clk(gclk));
	jdff dff_A_HMwz0DNp8_0(.dout(w_dff_A_HV3zwfae1_0),.din(w_dff_A_HMwz0DNp8_0),.clk(gclk));
	jdff dff_A_HV3zwfae1_0(.dout(w_dff_A_D6Sv39Nd2_0),.din(w_dff_A_HV3zwfae1_0),.clk(gclk));
	jdff dff_A_D6Sv39Nd2_0(.dout(w_dff_A_LMREqGFh0_0),.din(w_dff_A_D6Sv39Nd2_0),.clk(gclk));
	jdff dff_A_LMREqGFh0_0(.dout(w_dff_A_ca35UtDb1_0),.din(w_dff_A_LMREqGFh0_0),.clk(gclk));
	jdff dff_A_ca35UtDb1_0(.dout(w_dff_A_fd6Tv5PF4_0),.din(w_dff_A_ca35UtDb1_0),.clk(gclk));
	jdff dff_A_fd6Tv5PF4_0(.dout(w_dff_A_HWwoIRTV6_0),.din(w_dff_A_fd6Tv5PF4_0),.clk(gclk));
	jdff dff_A_HWwoIRTV6_0(.dout(w_dff_A_L1MFaNGw5_0),.din(w_dff_A_HWwoIRTV6_0),.clk(gclk));
	jdff dff_A_L1MFaNGw5_0(.dout(w_dff_A_gFWabiwQ6_0),.din(w_dff_A_L1MFaNGw5_0),.clk(gclk));
	jdff dff_A_gFWabiwQ6_0(.dout(w_dff_A_cSwBo1S84_0),.din(w_dff_A_gFWabiwQ6_0),.clk(gclk));
	jdff dff_A_cSwBo1S84_0(.dout(w_dff_A_296taM8l5_0),.din(w_dff_A_cSwBo1S84_0),.clk(gclk));
	jdff dff_A_296taM8l5_0(.dout(w_dff_A_jYimi9zI3_0),.din(w_dff_A_296taM8l5_0),.clk(gclk));
	jdff dff_A_jYimi9zI3_0(.dout(w_dff_A_B2ceTytw6_0),.din(w_dff_A_jYimi9zI3_0),.clk(gclk));
	jdff dff_A_B2ceTytw6_0(.dout(w_dff_A_uzxHMbEa7_0),.din(w_dff_A_B2ceTytw6_0),.clk(gclk));
	jdff dff_A_uzxHMbEa7_0(.dout(w_dff_A_RVlSOjWJ5_0),.din(w_dff_A_uzxHMbEa7_0),.clk(gclk));
	jdff dff_A_RVlSOjWJ5_0(.dout(w_dff_A_p8j1fZJX5_0),.din(w_dff_A_RVlSOjWJ5_0),.clk(gclk));
	jdff dff_A_p8j1fZJX5_0(.dout(w_dff_A_p3UBz73t9_0),.din(w_dff_A_p8j1fZJX5_0),.clk(gclk));
	jdff dff_A_p3UBz73t9_0(.dout(w_dff_A_Dq2CU8ir5_0),.din(w_dff_A_p3UBz73t9_0),.clk(gclk));
	jdff dff_A_Dq2CU8ir5_0(.dout(w_dff_A_uNVvBkCR0_0),.din(w_dff_A_Dq2CU8ir5_0),.clk(gclk));
	jdff dff_A_uNVvBkCR0_0(.dout(w_dff_A_q3j452TK6_0),.din(w_dff_A_uNVvBkCR0_0),.clk(gclk));
	jdff dff_A_q3j452TK6_0(.dout(w_dff_A_FbW9FTP21_0),.din(w_dff_A_q3j452TK6_0),.clk(gclk));
	jdff dff_A_FbW9FTP21_0(.dout(w_dff_A_b36pVjRq4_0),.din(w_dff_A_FbW9FTP21_0),.clk(gclk));
	jdff dff_A_b36pVjRq4_0(.dout(w_dff_A_oECxZpiS8_0),.din(w_dff_A_b36pVjRq4_0),.clk(gclk));
	jdff dff_A_oECxZpiS8_0(.dout(w_dff_A_6w8racrw7_0),.din(w_dff_A_oECxZpiS8_0),.clk(gclk));
	jdff dff_A_6w8racrw7_0(.dout(w_dff_A_4BaqbvN94_0),.din(w_dff_A_6w8racrw7_0),.clk(gclk));
	jdff dff_A_4BaqbvN94_0(.dout(G389gat),.din(w_dff_A_4BaqbvN94_0),.clk(gclk));
	jdff dff_A_xEjasLss1_2(.dout(w_dff_A_S4BSjuEv6_0),.din(w_dff_A_xEjasLss1_2),.clk(gclk));
	jdff dff_A_S4BSjuEv6_0(.dout(w_dff_A_u0TSUPbc6_0),.din(w_dff_A_S4BSjuEv6_0),.clk(gclk));
	jdff dff_A_u0TSUPbc6_0(.dout(w_dff_A_AE9M0Kb65_0),.din(w_dff_A_u0TSUPbc6_0),.clk(gclk));
	jdff dff_A_AE9M0Kb65_0(.dout(w_dff_A_h3Pgjv6l0_0),.din(w_dff_A_AE9M0Kb65_0),.clk(gclk));
	jdff dff_A_h3Pgjv6l0_0(.dout(w_dff_A_obBNlIvk1_0),.din(w_dff_A_h3Pgjv6l0_0),.clk(gclk));
	jdff dff_A_obBNlIvk1_0(.dout(w_dff_A_WbJC8jyf2_0),.din(w_dff_A_obBNlIvk1_0),.clk(gclk));
	jdff dff_A_WbJC8jyf2_0(.dout(w_dff_A_0JLLsif19_0),.din(w_dff_A_WbJC8jyf2_0),.clk(gclk));
	jdff dff_A_0JLLsif19_0(.dout(w_dff_A_iLzIIg2s4_0),.din(w_dff_A_0JLLsif19_0),.clk(gclk));
	jdff dff_A_iLzIIg2s4_0(.dout(w_dff_A_HXdi2wXa4_0),.din(w_dff_A_iLzIIg2s4_0),.clk(gclk));
	jdff dff_A_HXdi2wXa4_0(.dout(w_dff_A_qud9klAs1_0),.din(w_dff_A_HXdi2wXa4_0),.clk(gclk));
	jdff dff_A_qud9klAs1_0(.dout(w_dff_A_vryFEqRx4_0),.din(w_dff_A_qud9klAs1_0),.clk(gclk));
	jdff dff_A_vryFEqRx4_0(.dout(w_dff_A_Ac9i4vmv3_0),.din(w_dff_A_vryFEqRx4_0),.clk(gclk));
	jdff dff_A_Ac9i4vmv3_0(.dout(w_dff_A_60t3tQxw1_0),.din(w_dff_A_Ac9i4vmv3_0),.clk(gclk));
	jdff dff_A_60t3tQxw1_0(.dout(w_dff_A_daHJC0Hc7_0),.din(w_dff_A_60t3tQxw1_0),.clk(gclk));
	jdff dff_A_daHJC0Hc7_0(.dout(w_dff_A_3SGc56OH4_0),.din(w_dff_A_daHJC0Hc7_0),.clk(gclk));
	jdff dff_A_3SGc56OH4_0(.dout(w_dff_A_daKrQNTC3_0),.din(w_dff_A_3SGc56OH4_0),.clk(gclk));
	jdff dff_A_daKrQNTC3_0(.dout(w_dff_A_KnwKOTlc6_0),.din(w_dff_A_daKrQNTC3_0),.clk(gclk));
	jdff dff_A_KnwKOTlc6_0(.dout(w_dff_A_ytdODurQ0_0),.din(w_dff_A_KnwKOTlc6_0),.clk(gclk));
	jdff dff_A_ytdODurQ0_0(.dout(w_dff_A_ivYdgyuy5_0),.din(w_dff_A_ytdODurQ0_0),.clk(gclk));
	jdff dff_A_ivYdgyuy5_0(.dout(w_dff_A_PbTYPrLf1_0),.din(w_dff_A_ivYdgyuy5_0),.clk(gclk));
	jdff dff_A_PbTYPrLf1_0(.dout(w_dff_A_u0x9AqAx3_0),.din(w_dff_A_PbTYPrLf1_0),.clk(gclk));
	jdff dff_A_u0x9AqAx3_0(.dout(w_dff_A_4lOJXUlQ6_0),.din(w_dff_A_u0x9AqAx3_0),.clk(gclk));
	jdff dff_A_4lOJXUlQ6_0(.dout(w_dff_A_0gIa4O151_0),.din(w_dff_A_4lOJXUlQ6_0),.clk(gclk));
	jdff dff_A_0gIa4O151_0(.dout(w_dff_A_wNt5qoBd0_0),.din(w_dff_A_0gIa4O151_0),.clk(gclk));
	jdff dff_A_wNt5qoBd0_0(.dout(w_dff_A_o0SInsMd8_0),.din(w_dff_A_wNt5qoBd0_0),.clk(gclk));
	jdff dff_A_o0SInsMd8_0(.dout(G390gat),.din(w_dff_A_o0SInsMd8_0),.clk(gclk));
	jdff dff_A_Cbt2rFAg8_2(.dout(w_dff_A_1MyEp29m8_0),.din(w_dff_A_Cbt2rFAg8_2),.clk(gclk));
	jdff dff_A_1MyEp29m8_0(.dout(w_dff_A_XvKS7zT87_0),.din(w_dff_A_1MyEp29m8_0),.clk(gclk));
	jdff dff_A_XvKS7zT87_0(.dout(w_dff_A_YlJyR9GJ6_0),.din(w_dff_A_XvKS7zT87_0),.clk(gclk));
	jdff dff_A_YlJyR9GJ6_0(.dout(w_dff_A_a0weg2kE5_0),.din(w_dff_A_YlJyR9GJ6_0),.clk(gclk));
	jdff dff_A_a0weg2kE5_0(.dout(w_dff_A_TQM7qa7r1_0),.din(w_dff_A_a0weg2kE5_0),.clk(gclk));
	jdff dff_A_TQM7qa7r1_0(.dout(w_dff_A_S9G4N98N7_0),.din(w_dff_A_TQM7qa7r1_0),.clk(gclk));
	jdff dff_A_S9G4N98N7_0(.dout(w_dff_A_cqp1KyIn0_0),.din(w_dff_A_S9G4N98N7_0),.clk(gclk));
	jdff dff_A_cqp1KyIn0_0(.dout(w_dff_A_NhjFSoQ59_0),.din(w_dff_A_cqp1KyIn0_0),.clk(gclk));
	jdff dff_A_NhjFSoQ59_0(.dout(w_dff_A_1jGBqCSY7_0),.din(w_dff_A_NhjFSoQ59_0),.clk(gclk));
	jdff dff_A_1jGBqCSY7_0(.dout(w_dff_A_BCeEtFbI2_0),.din(w_dff_A_1jGBqCSY7_0),.clk(gclk));
	jdff dff_A_BCeEtFbI2_0(.dout(w_dff_A_D80TTEYH3_0),.din(w_dff_A_BCeEtFbI2_0),.clk(gclk));
	jdff dff_A_D80TTEYH3_0(.dout(w_dff_A_l9kjwhD18_0),.din(w_dff_A_D80TTEYH3_0),.clk(gclk));
	jdff dff_A_l9kjwhD18_0(.dout(w_dff_A_r1HOiBy80_0),.din(w_dff_A_l9kjwhD18_0),.clk(gclk));
	jdff dff_A_r1HOiBy80_0(.dout(w_dff_A_WrP7NWcZ3_0),.din(w_dff_A_r1HOiBy80_0),.clk(gclk));
	jdff dff_A_WrP7NWcZ3_0(.dout(w_dff_A_SObQLSJS2_0),.din(w_dff_A_WrP7NWcZ3_0),.clk(gclk));
	jdff dff_A_SObQLSJS2_0(.dout(w_dff_A_trccRMOl7_0),.din(w_dff_A_SObQLSJS2_0),.clk(gclk));
	jdff dff_A_trccRMOl7_0(.dout(w_dff_A_eFKgkVmo2_0),.din(w_dff_A_trccRMOl7_0),.clk(gclk));
	jdff dff_A_eFKgkVmo2_0(.dout(w_dff_A_vOK49FMM8_0),.din(w_dff_A_eFKgkVmo2_0),.clk(gclk));
	jdff dff_A_vOK49FMM8_0(.dout(w_dff_A_cByvQm4W0_0),.din(w_dff_A_vOK49FMM8_0),.clk(gclk));
	jdff dff_A_cByvQm4W0_0(.dout(w_dff_A_zXxNE0wq8_0),.din(w_dff_A_cByvQm4W0_0),.clk(gclk));
	jdff dff_A_zXxNE0wq8_0(.dout(w_dff_A_2CNvd6hu5_0),.din(w_dff_A_zXxNE0wq8_0),.clk(gclk));
	jdff dff_A_2CNvd6hu5_0(.dout(w_dff_A_gUL5Fqwn9_0),.din(w_dff_A_2CNvd6hu5_0),.clk(gclk));
	jdff dff_A_gUL5Fqwn9_0(.dout(w_dff_A_8hs3jjnI3_0),.din(w_dff_A_gUL5Fqwn9_0),.clk(gclk));
	jdff dff_A_8hs3jjnI3_0(.dout(w_dff_A_aFRDWzMY2_0),.din(w_dff_A_8hs3jjnI3_0),.clk(gclk));
	jdff dff_A_aFRDWzMY2_0(.dout(w_dff_A_VTodtSkO6_0),.din(w_dff_A_aFRDWzMY2_0),.clk(gclk));
	jdff dff_A_VTodtSkO6_0(.dout(w_dff_A_h4I0Sdyv3_0),.din(w_dff_A_VTodtSkO6_0),.clk(gclk));
	jdff dff_A_h4I0Sdyv3_0(.dout(G391gat),.din(w_dff_A_h4I0Sdyv3_0),.clk(gclk));
	jdff dff_A_JJMPLPol7_2(.dout(w_dff_A_zxJ2Df549_0),.din(w_dff_A_JJMPLPol7_2),.clk(gclk));
	jdff dff_A_zxJ2Df549_0(.dout(w_dff_A_yBRMDJhx8_0),.din(w_dff_A_zxJ2Df549_0),.clk(gclk));
	jdff dff_A_yBRMDJhx8_0(.dout(w_dff_A_kwigkLOH3_0),.din(w_dff_A_yBRMDJhx8_0),.clk(gclk));
	jdff dff_A_kwigkLOH3_0(.dout(w_dff_A_MCQAO53A7_0),.din(w_dff_A_kwigkLOH3_0),.clk(gclk));
	jdff dff_A_MCQAO53A7_0(.dout(w_dff_A_iBEuXitr9_0),.din(w_dff_A_MCQAO53A7_0),.clk(gclk));
	jdff dff_A_iBEuXitr9_0(.dout(w_dff_A_4bafrp5H0_0),.din(w_dff_A_iBEuXitr9_0),.clk(gclk));
	jdff dff_A_4bafrp5H0_0(.dout(w_dff_A_dcKDPXzk9_0),.din(w_dff_A_4bafrp5H0_0),.clk(gclk));
	jdff dff_A_dcKDPXzk9_0(.dout(w_dff_A_jrUf9jZz0_0),.din(w_dff_A_dcKDPXzk9_0),.clk(gclk));
	jdff dff_A_jrUf9jZz0_0(.dout(w_dff_A_ChxVa4a04_0),.din(w_dff_A_jrUf9jZz0_0),.clk(gclk));
	jdff dff_A_ChxVa4a04_0(.dout(w_dff_A_A3bHpQhj3_0),.din(w_dff_A_ChxVa4a04_0),.clk(gclk));
	jdff dff_A_A3bHpQhj3_0(.dout(w_dff_A_XsRhZxzX1_0),.din(w_dff_A_A3bHpQhj3_0),.clk(gclk));
	jdff dff_A_XsRhZxzX1_0(.dout(w_dff_A_jB7Si0fg3_0),.din(w_dff_A_XsRhZxzX1_0),.clk(gclk));
	jdff dff_A_jB7Si0fg3_0(.dout(w_dff_A_z8h3eS3X4_0),.din(w_dff_A_jB7Si0fg3_0),.clk(gclk));
	jdff dff_A_z8h3eS3X4_0(.dout(w_dff_A_BIEDadFO7_0),.din(w_dff_A_z8h3eS3X4_0),.clk(gclk));
	jdff dff_A_BIEDadFO7_0(.dout(w_dff_A_Jv4vFuU77_0),.din(w_dff_A_BIEDadFO7_0),.clk(gclk));
	jdff dff_A_Jv4vFuU77_0(.dout(w_dff_A_VBju6Dg06_0),.din(w_dff_A_Jv4vFuU77_0),.clk(gclk));
	jdff dff_A_VBju6Dg06_0(.dout(w_dff_A_Qb0xrRd38_0),.din(w_dff_A_VBju6Dg06_0),.clk(gclk));
	jdff dff_A_Qb0xrRd38_0(.dout(w_dff_A_N3n2jcgj9_0),.din(w_dff_A_Qb0xrRd38_0),.clk(gclk));
	jdff dff_A_N3n2jcgj9_0(.dout(w_dff_A_Z1HAv0Te5_0),.din(w_dff_A_N3n2jcgj9_0),.clk(gclk));
	jdff dff_A_Z1HAv0Te5_0(.dout(w_dff_A_3cQgvXZ49_0),.din(w_dff_A_Z1HAv0Te5_0),.clk(gclk));
	jdff dff_A_3cQgvXZ49_0(.dout(w_dff_A_hOUyfhGo9_0),.din(w_dff_A_3cQgvXZ49_0),.clk(gclk));
	jdff dff_A_hOUyfhGo9_0(.dout(w_dff_A_s6LtyaQZ9_0),.din(w_dff_A_hOUyfhGo9_0),.clk(gclk));
	jdff dff_A_s6LtyaQZ9_0(.dout(w_dff_A_vWmPcjBe7_0),.din(w_dff_A_s6LtyaQZ9_0),.clk(gclk));
	jdff dff_A_vWmPcjBe7_0(.dout(w_dff_A_jV1i1rqS4_0),.din(w_dff_A_vWmPcjBe7_0),.clk(gclk));
	jdff dff_A_jV1i1rqS4_0(.dout(G418gat),.din(w_dff_A_jV1i1rqS4_0),.clk(gclk));
	jdff dff_A_a7ON3QTw2_2(.dout(w_dff_A_DTgA1dQF9_0),.din(w_dff_A_a7ON3QTw2_2),.clk(gclk));
	jdff dff_A_DTgA1dQF9_0(.dout(w_dff_A_Xcmqkp3J5_0),.din(w_dff_A_DTgA1dQF9_0),.clk(gclk));
	jdff dff_A_Xcmqkp3J5_0(.dout(w_dff_A_Cm5WgIml4_0),.din(w_dff_A_Xcmqkp3J5_0),.clk(gclk));
	jdff dff_A_Cm5WgIml4_0(.dout(w_dff_A_0GzK5Pvj4_0),.din(w_dff_A_Cm5WgIml4_0),.clk(gclk));
	jdff dff_A_0GzK5Pvj4_0(.dout(w_dff_A_JV9dQzFw4_0),.din(w_dff_A_0GzK5Pvj4_0),.clk(gclk));
	jdff dff_A_JV9dQzFw4_0(.dout(w_dff_A_U389dqkI3_0),.din(w_dff_A_JV9dQzFw4_0),.clk(gclk));
	jdff dff_A_U389dqkI3_0(.dout(w_dff_A_dzGRMpLF4_0),.din(w_dff_A_U389dqkI3_0),.clk(gclk));
	jdff dff_A_dzGRMpLF4_0(.dout(w_dff_A_2xWTgVTf8_0),.din(w_dff_A_dzGRMpLF4_0),.clk(gclk));
	jdff dff_A_2xWTgVTf8_0(.dout(w_dff_A_lXs6Jn781_0),.din(w_dff_A_2xWTgVTf8_0),.clk(gclk));
	jdff dff_A_lXs6Jn781_0(.dout(w_dff_A_imRzTusE1_0),.din(w_dff_A_lXs6Jn781_0),.clk(gclk));
	jdff dff_A_imRzTusE1_0(.dout(w_dff_A_FulKy1cM0_0),.din(w_dff_A_imRzTusE1_0),.clk(gclk));
	jdff dff_A_FulKy1cM0_0(.dout(w_dff_A_1JEw5cSI1_0),.din(w_dff_A_FulKy1cM0_0),.clk(gclk));
	jdff dff_A_1JEw5cSI1_0(.dout(w_dff_A_efmcyHqd5_0),.din(w_dff_A_1JEw5cSI1_0),.clk(gclk));
	jdff dff_A_efmcyHqd5_0(.dout(w_dff_A_A7mAtw7O5_0),.din(w_dff_A_efmcyHqd5_0),.clk(gclk));
	jdff dff_A_A7mAtw7O5_0(.dout(w_dff_A_GEZ9vhTE6_0),.din(w_dff_A_A7mAtw7O5_0),.clk(gclk));
	jdff dff_A_GEZ9vhTE6_0(.dout(w_dff_A_EYkfTLMA4_0),.din(w_dff_A_GEZ9vhTE6_0),.clk(gclk));
	jdff dff_A_EYkfTLMA4_0(.dout(w_dff_A_yNFT2uKZ8_0),.din(w_dff_A_EYkfTLMA4_0),.clk(gclk));
	jdff dff_A_yNFT2uKZ8_0(.dout(w_dff_A_ye6WrywS0_0),.din(w_dff_A_yNFT2uKZ8_0),.clk(gclk));
	jdff dff_A_ye6WrywS0_0(.dout(w_dff_A_I60293s53_0),.din(w_dff_A_ye6WrywS0_0),.clk(gclk));
	jdff dff_A_I60293s53_0(.dout(w_dff_A_fP4q7mAE3_0),.din(w_dff_A_I60293s53_0),.clk(gclk));
	jdff dff_A_fP4q7mAE3_0(.dout(w_dff_A_daZmWlMT8_0),.din(w_dff_A_fP4q7mAE3_0),.clk(gclk));
	jdff dff_A_daZmWlMT8_0(.dout(w_dff_A_TnxqdI4c1_0),.din(w_dff_A_daZmWlMT8_0),.clk(gclk));
	jdff dff_A_TnxqdI4c1_0(.dout(G419gat),.din(w_dff_A_TnxqdI4c1_0),.clk(gclk));
	jdff dff_A_sGkqRViV5_2(.dout(w_dff_A_7xCTlbl73_0),.din(w_dff_A_sGkqRViV5_2),.clk(gclk));
	jdff dff_A_7xCTlbl73_0(.dout(w_dff_A_FbKaRzbb5_0),.din(w_dff_A_7xCTlbl73_0),.clk(gclk));
	jdff dff_A_FbKaRzbb5_0(.dout(w_dff_A_Oq84gOft3_0),.din(w_dff_A_FbKaRzbb5_0),.clk(gclk));
	jdff dff_A_Oq84gOft3_0(.dout(w_dff_A_PpDO167k2_0),.din(w_dff_A_Oq84gOft3_0),.clk(gclk));
	jdff dff_A_PpDO167k2_0(.dout(w_dff_A_Y455jQ0n4_0),.din(w_dff_A_PpDO167k2_0),.clk(gclk));
	jdff dff_A_Y455jQ0n4_0(.dout(w_dff_A_TtXrNHfD9_0),.din(w_dff_A_Y455jQ0n4_0),.clk(gclk));
	jdff dff_A_TtXrNHfD9_0(.dout(w_dff_A_KvGDVl7u2_0),.din(w_dff_A_TtXrNHfD9_0),.clk(gclk));
	jdff dff_A_KvGDVl7u2_0(.dout(w_dff_A_1cXROs9R2_0),.din(w_dff_A_KvGDVl7u2_0),.clk(gclk));
	jdff dff_A_1cXROs9R2_0(.dout(w_dff_A_7q2YFTi09_0),.din(w_dff_A_1cXROs9R2_0),.clk(gclk));
	jdff dff_A_7q2YFTi09_0(.dout(w_dff_A_tBKDfHWq7_0),.din(w_dff_A_7q2YFTi09_0),.clk(gclk));
	jdff dff_A_tBKDfHWq7_0(.dout(w_dff_A_U5wuA1fv2_0),.din(w_dff_A_tBKDfHWq7_0),.clk(gclk));
	jdff dff_A_U5wuA1fv2_0(.dout(w_dff_A_5ND1oFoY5_0),.din(w_dff_A_U5wuA1fv2_0),.clk(gclk));
	jdff dff_A_5ND1oFoY5_0(.dout(w_dff_A_LA91jVVJ0_0),.din(w_dff_A_5ND1oFoY5_0),.clk(gclk));
	jdff dff_A_LA91jVVJ0_0(.dout(w_dff_A_j5En6ecb7_0),.din(w_dff_A_LA91jVVJ0_0),.clk(gclk));
	jdff dff_A_j5En6ecb7_0(.dout(w_dff_A_JC8OGn1F0_0),.din(w_dff_A_j5En6ecb7_0),.clk(gclk));
	jdff dff_A_JC8OGn1F0_0(.dout(w_dff_A_tPYt13Bd3_0),.din(w_dff_A_JC8OGn1F0_0),.clk(gclk));
	jdff dff_A_tPYt13Bd3_0(.dout(w_dff_A_UCbCiM7p0_0),.din(w_dff_A_tPYt13Bd3_0),.clk(gclk));
	jdff dff_A_UCbCiM7p0_0(.dout(w_dff_A_3aksizyi0_0),.din(w_dff_A_UCbCiM7p0_0),.clk(gclk));
	jdff dff_A_3aksizyi0_0(.dout(w_dff_A_Nw4UEA4k9_0),.din(w_dff_A_3aksizyi0_0),.clk(gclk));
	jdff dff_A_Nw4UEA4k9_0(.dout(w_dff_A_18YPC1vo5_0),.din(w_dff_A_Nw4UEA4k9_0),.clk(gclk));
	jdff dff_A_18YPC1vo5_0(.dout(w_dff_A_km4XTKFV5_0),.din(w_dff_A_18YPC1vo5_0),.clk(gclk));
	jdff dff_A_km4XTKFV5_0(.dout(w_dff_A_hQAagMdR9_0),.din(w_dff_A_km4XTKFV5_0),.clk(gclk));
	jdff dff_A_hQAagMdR9_0(.dout(w_dff_A_pFwlOgAu4_0),.din(w_dff_A_hQAagMdR9_0),.clk(gclk));
	jdff dff_A_pFwlOgAu4_0(.dout(w_dff_A_Yz1levAm9_0),.din(w_dff_A_pFwlOgAu4_0),.clk(gclk));
	jdff dff_A_Yz1levAm9_0(.dout(G420gat),.din(w_dff_A_Yz1levAm9_0),.clk(gclk));
	jdff dff_A_BHZ57keO2_2(.dout(w_dff_A_taGKzJPg3_0),.din(w_dff_A_BHZ57keO2_2),.clk(gclk));
	jdff dff_A_taGKzJPg3_0(.dout(w_dff_A_EbK3gKnN3_0),.din(w_dff_A_taGKzJPg3_0),.clk(gclk));
	jdff dff_A_EbK3gKnN3_0(.dout(w_dff_A_fzw0d7ND8_0),.din(w_dff_A_EbK3gKnN3_0),.clk(gclk));
	jdff dff_A_fzw0d7ND8_0(.dout(w_dff_A_Y6kPJhE06_0),.din(w_dff_A_fzw0d7ND8_0),.clk(gclk));
	jdff dff_A_Y6kPJhE06_0(.dout(w_dff_A_qxPrS9xV0_0),.din(w_dff_A_Y6kPJhE06_0),.clk(gclk));
	jdff dff_A_qxPrS9xV0_0(.dout(w_dff_A_Eaj43ibm4_0),.din(w_dff_A_qxPrS9xV0_0),.clk(gclk));
	jdff dff_A_Eaj43ibm4_0(.dout(w_dff_A_JYvudEBN0_0),.din(w_dff_A_Eaj43ibm4_0),.clk(gclk));
	jdff dff_A_JYvudEBN0_0(.dout(w_dff_A_whqszE3R1_0),.din(w_dff_A_JYvudEBN0_0),.clk(gclk));
	jdff dff_A_whqszE3R1_0(.dout(w_dff_A_xU6hoIzQ9_0),.din(w_dff_A_whqszE3R1_0),.clk(gclk));
	jdff dff_A_xU6hoIzQ9_0(.dout(w_dff_A_ntLWWh2T0_0),.din(w_dff_A_xU6hoIzQ9_0),.clk(gclk));
	jdff dff_A_ntLWWh2T0_0(.dout(w_dff_A_k5sL1d9Y5_0),.din(w_dff_A_ntLWWh2T0_0),.clk(gclk));
	jdff dff_A_k5sL1d9Y5_0(.dout(w_dff_A_Gjl8uLap7_0),.din(w_dff_A_k5sL1d9Y5_0),.clk(gclk));
	jdff dff_A_Gjl8uLap7_0(.dout(w_dff_A_hGpaFSkD3_0),.din(w_dff_A_Gjl8uLap7_0),.clk(gclk));
	jdff dff_A_hGpaFSkD3_0(.dout(w_dff_A_VTGlvQ4I5_0),.din(w_dff_A_hGpaFSkD3_0),.clk(gclk));
	jdff dff_A_VTGlvQ4I5_0(.dout(w_dff_A_QihP0Aci1_0),.din(w_dff_A_VTGlvQ4I5_0),.clk(gclk));
	jdff dff_A_QihP0Aci1_0(.dout(w_dff_A_cX9qwrjL3_0),.din(w_dff_A_QihP0Aci1_0),.clk(gclk));
	jdff dff_A_cX9qwrjL3_0(.dout(w_dff_A_V7dbeJo28_0),.din(w_dff_A_cX9qwrjL3_0),.clk(gclk));
	jdff dff_A_V7dbeJo28_0(.dout(w_dff_A_PDG6DZXt0_0),.din(w_dff_A_V7dbeJo28_0),.clk(gclk));
	jdff dff_A_PDG6DZXt0_0(.dout(w_dff_A_anMJzwjP0_0),.din(w_dff_A_PDG6DZXt0_0),.clk(gclk));
	jdff dff_A_anMJzwjP0_0(.dout(w_dff_A_esdq5fg16_0),.din(w_dff_A_anMJzwjP0_0),.clk(gclk));
	jdff dff_A_esdq5fg16_0(.dout(w_dff_A_oc3xFxVt5_0),.din(w_dff_A_esdq5fg16_0),.clk(gclk));
	jdff dff_A_oc3xFxVt5_0(.dout(w_dff_A_HcZgitik1_0),.din(w_dff_A_oc3xFxVt5_0),.clk(gclk));
	jdff dff_A_HcZgitik1_0(.dout(w_dff_A_eYRAqSb62_0),.din(w_dff_A_HcZgitik1_0),.clk(gclk));
	jdff dff_A_eYRAqSb62_0(.dout(w_dff_A_jTIiErZg3_0),.din(w_dff_A_eYRAqSb62_0),.clk(gclk));
	jdff dff_A_jTIiErZg3_0(.dout(G421gat),.din(w_dff_A_jTIiErZg3_0),.clk(gclk));
	jdff dff_A_NliuMYGZ6_2(.dout(w_dff_A_CFniME9j9_0),.din(w_dff_A_NliuMYGZ6_2),.clk(gclk));
	jdff dff_A_CFniME9j9_0(.dout(w_dff_A_McNRy9Yo9_0),.din(w_dff_A_CFniME9j9_0),.clk(gclk));
	jdff dff_A_McNRy9Yo9_0(.dout(w_dff_A_cGZP2Qm32_0),.din(w_dff_A_McNRy9Yo9_0),.clk(gclk));
	jdff dff_A_cGZP2Qm32_0(.dout(w_dff_A_FQgyl4FQ6_0),.din(w_dff_A_cGZP2Qm32_0),.clk(gclk));
	jdff dff_A_FQgyl4FQ6_0(.dout(w_dff_A_Y0mWhTRw7_0),.din(w_dff_A_FQgyl4FQ6_0),.clk(gclk));
	jdff dff_A_Y0mWhTRw7_0(.dout(w_dff_A_jJunn7vf3_0),.din(w_dff_A_Y0mWhTRw7_0),.clk(gclk));
	jdff dff_A_jJunn7vf3_0(.dout(w_dff_A_hk2NxoL14_0),.din(w_dff_A_jJunn7vf3_0),.clk(gclk));
	jdff dff_A_hk2NxoL14_0(.dout(w_dff_A_8soCHyqz9_0),.din(w_dff_A_hk2NxoL14_0),.clk(gclk));
	jdff dff_A_8soCHyqz9_0(.dout(w_dff_A_zkWQI8Kg0_0),.din(w_dff_A_8soCHyqz9_0),.clk(gclk));
	jdff dff_A_zkWQI8Kg0_0(.dout(w_dff_A_v1ffeCSe4_0),.din(w_dff_A_zkWQI8Kg0_0),.clk(gclk));
	jdff dff_A_v1ffeCSe4_0(.dout(w_dff_A_pFTUNJCc4_0),.din(w_dff_A_v1ffeCSe4_0),.clk(gclk));
	jdff dff_A_pFTUNJCc4_0(.dout(w_dff_A_qedkkuD08_0),.din(w_dff_A_pFTUNJCc4_0),.clk(gclk));
	jdff dff_A_qedkkuD08_0(.dout(w_dff_A_StBpS3jA8_0),.din(w_dff_A_qedkkuD08_0),.clk(gclk));
	jdff dff_A_StBpS3jA8_0(.dout(w_dff_A_nptZEgg33_0),.din(w_dff_A_StBpS3jA8_0),.clk(gclk));
	jdff dff_A_nptZEgg33_0(.dout(w_dff_A_6i0osKXe2_0),.din(w_dff_A_nptZEgg33_0),.clk(gclk));
	jdff dff_A_6i0osKXe2_0(.dout(w_dff_A_PTevI6bL9_0),.din(w_dff_A_6i0osKXe2_0),.clk(gclk));
	jdff dff_A_PTevI6bL9_0(.dout(w_dff_A_j8esl1S99_0),.din(w_dff_A_PTevI6bL9_0),.clk(gclk));
	jdff dff_A_j8esl1S99_0(.dout(w_dff_A_psNGMqjG3_0),.din(w_dff_A_j8esl1S99_0),.clk(gclk));
	jdff dff_A_psNGMqjG3_0(.dout(w_dff_A_XewaMgJw4_0),.din(w_dff_A_psNGMqjG3_0),.clk(gclk));
	jdff dff_A_XewaMgJw4_0(.dout(w_dff_A_ENaEuGdi8_0),.din(w_dff_A_XewaMgJw4_0),.clk(gclk));
	jdff dff_A_ENaEuGdi8_0(.dout(w_dff_A_XcLFnf3w2_0),.din(w_dff_A_ENaEuGdi8_0),.clk(gclk));
	jdff dff_A_XcLFnf3w2_0(.dout(w_dff_A_WM3so4VJ7_0),.din(w_dff_A_XcLFnf3w2_0),.clk(gclk));
	jdff dff_A_WM3so4VJ7_0(.dout(w_dff_A_4xocwfny9_0),.din(w_dff_A_WM3so4VJ7_0),.clk(gclk));
	jdff dff_A_4xocwfny9_0(.dout(w_dff_A_85WkFkzR8_0),.din(w_dff_A_4xocwfny9_0),.clk(gclk));
	jdff dff_A_85WkFkzR8_0(.dout(G422gat),.din(w_dff_A_85WkFkzR8_0),.clk(gclk));
	jdff dff_A_iuAfvJlo7_2(.dout(w_dff_A_7zyp774y3_0),.din(w_dff_A_iuAfvJlo7_2),.clk(gclk));
	jdff dff_A_7zyp774y3_0(.dout(w_dff_A_o0QDc4Lj0_0),.din(w_dff_A_7zyp774y3_0),.clk(gclk));
	jdff dff_A_o0QDc4Lj0_0(.dout(w_dff_A_Z9xshVnD3_0),.din(w_dff_A_o0QDc4Lj0_0),.clk(gclk));
	jdff dff_A_Z9xshVnD3_0(.dout(w_dff_A_2U4ebGGE2_0),.din(w_dff_A_Z9xshVnD3_0),.clk(gclk));
	jdff dff_A_2U4ebGGE2_0(.dout(w_dff_A_JpcVDTG93_0),.din(w_dff_A_2U4ebGGE2_0),.clk(gclk));
	jdff dff_A_JpcVDTG93_0(.dout(w_dff_A_dED0aKgU3_0),.din(w_dff_A_JpcVDTG93_0),.clk(gclk));
	jdff dff_A_dED0aKgU3_0(.dout(w_dff_A_fFck0DHD1_0),.din(w_dff_A_dED0aKgU3_0),.clk(gclk));
	jdff dff_A_fFck0DHD1_0(.dout(w_dff_A_j6hya3RE5_0),.din(w_dff_A_fFck0DHD1_0),.clk(gclk));
	jdff dff_A_j6hya3RE5_0(.dout(w_dff_A_8uijJj7v2_0),.din(w_dff_A_j6hya3RE5_0),.clk(gclk));
	jdff dff_A_8uijJj7v2_0(.dout(w_dff_A_cKWoBNME2_0),.din(w_dff_A_8uijJj7v2_0),.clk(gclk));
	jdff dff_A_cKWoBNME2_0(.dout(w_dff_A_fVRFjDS67_0),.din(w_dff_A_cKWoBNME2_0),.clk(gclk));
	jdff dff_A_fVRFjDS67_0(.dout(w_dff_A_dfitOVYm9_0),.din(w_dff_A_fVRFjDS67_0),.clk(gclk));
	jdff dff_A_dfitOVYm9_0(.dout(w_dff_A_FpDDf8581_0),.din(w_dff_A_dfitOVYm9_0),.clk(gclk));
	jdff dff_A_FpDDf8581_0(.dout(w_dff_A_xEveGCUn3_0),.din(w_dff_A_FpDDf8581_0),.clk(gclk));
	jdff dff_A_xEveGCUn3_0(.dout(w_dff_A_EN62yg8U2_0),.din(w_dff_A_xEveGCUn3_0),.clk(gclk));
	jdff dff_A_EN62yg8U2_0(.dout(w_dff_A_j90Emxzm1_0),.din(w_dff_A_EN62yg8U2_0),.clk(gclk));
	jdff dff_A_j90Emxzm1_0(.dout(w_dff_A_9wadJcyZ9_0),.din(w_dff_A_j90Emxzm1_0),.clk(gclk));
	jdff dff_A_9wadJcyZ9_0(.dout(w_dff_A_EemJd0qx1_0),.din(w_dff_A_9wadJcyZ9_0),.clk(gclk));
	jdff dff_A_EemJd0qx1_0(.dout(w_dff_A_wMVKlU2i0_0),.din(w_dff_A_EemJd0qx1_0),.clk(gclk));
	jdff dff_A_wMVKlU2i0_0(.dout(w_dff_A_mG2gUNQ59_0),.din(w_dff_A_wMVKlU2i0_0),.clk(gclk));
	jdff dff_A_mG2gUNQ59_0(.dout(w_dff_A_YASmzfXQ1_0),.din(w_dff_A_mG2gUNQ59_0),.clk(gclk));
	jdff dff_A_YASmzfXQ1_0(.dout(w_dff_A_V5VILOyP8_0),.din(w_dff_A_YASmzfXQ1_0),.clk(gclk));
	jdff dff_A_V5VILOyP8_0(.dout(w_dff_A_e5W7SCNd9_0),.din(w_dff_A_V5VILOyP8_0),.clk(gclk));
	jdff dff_A_e5W7SCNd9_0(.dout(w_dff_A_IlmZkdRu3_0),.din(w_dff_A_e5W7SCNd9_0),.clk(gclk));
	jdff dff_A_IlmZkdRu3_0(.dout(w_dff_A_pJD6yBb64_0),.din(w_dff_A_IlmZkdRu3_0),.clk(gclk));
	jdff dff_A_pJD6yBb64_0(.dout(G423gat),.din(w_dff_A_pJD6yBb64_0),.clk(gclk));
	jdff dff_A_L5QySJRo8_2(.dout(w_dff_A_F2qGzpBA7_0),.din(w_dff_A_L5QySJRo8_2),.clk(gclk));
	jdff dff_A_F2qGzpBA7_0(.dout(w_dff_A_TQ2wNTcd7_0),.din(w_dff_A_F2qGzpBA7_0),.clk(gclk));
	jdff dff_A_TQ2wNTcd7_0(.dout(w_dff_A_nzGkn6xV0_0),.din(w_dff_A_TQ2wNTcd7_0),.clk(gclk));
	jdff dff_A_nzGkn6xV0_0(.dout(w_dff_A_6xVT5N4Z7_0),.din(w_dff_A_nzGkn6xV0_0),.clk(gclk));
	jdff dff_A_6xVT5N4Z7_0(.dout(w_dff_A_7vDB6KNm7_0),.din(w_dff_A_6xVT5N4Z7_0),.clk(gclk));
	jdff dff_A_7vDB6KNm7_0(.dout(w_dff_A_1MQN4qje1_0),.din(w_dff_A_7vDB6KNm7_0),.clk(gclk));
	jdff dff_A_1MQN4qje1_0(.dout(w_dff_A_JYPV7wm15_0),.din(w_dff_A_1MQN4qje1_0),.clk(gclk));
	jdff dff_A_JYPV7wm15_0(.dout(w_dff_A_2GsegVcI0_0),.din(w_dff_A_JYPV7wm15_0),.clk(gclk));
	jdff dff_A_2GsegVcI0_0(.dout(w_dff_A_YzrW7Ovp0_0),.din(w_dff_A_2GsegVcI0_0),.clk(gclk));
	jdff dff_A_YzrW7Ovp0_0(.dout(w_dff_A_gjnV77zI2_0),.din(w_dff_A_YzrW7Ovp0_0),.clk(gclk));
	jdff dff_A_gjnV77zI2_0(.dout(w_dff_A_PNNuSGOK1_0),.din(w_dff_A_gjnV77zI2_0),.clk(gclk));
	jdff dff_A_PNNuSGOK1_0(.dout(w_dff_A_3bqyUTnF6_0),.din(w_dff_A_PNNuSGOK1_0),.clk(gclk));
	jdff dff_A_3bqyUTnF6_0(.dout(w_dff_A_9evnXDIv3_0),.din(w_dff_A_3bqyUTnF6_0),.clk(gclk));
	jdff dff_A_9evnXDIv3_0(.dout(w_dff_A_xtU66SQn3_0),.din(w_dff_A_9evnXDIv3_0),.clk(gclk));
	jdff dff_A_xtU66SQn3_0(.dout(w_dff_A_JFyU1dCK7_0),.din(w_dff_A_xtU66SQn3_0),.clk(gclk));
	jdff dff_A_JFyU1dCK7_0(.dout(w_dff_A_aQADH9PS5_0),.din(w_dff_A_JFyU1dCK7_0),.clk(gclk));
	jdff dff_A_aQADH9PS5_0(.dout(w_dff_A_7seewoh85_0),.din(w_dff_A_aQADH9PS5_0),.clk(gclk));
	jdff dff_A_7seewoh85_0(.dout(w_dff_A_CBENJXHJ6_0),.din(w_dff_A_7seewoh85_0),.clk(gclk));
	jdff dff_A_CBENJXHJ6_0(.dout(w_dff_A_HO9PsLxw8_0),.din(w_dff_A_CBENJXHJ6_0),.clk(gclk));
	jdff dff_A_HO9PsLxw8_0(.dout(w_dff_A_xFSUe6E94_0),.din(w_dff_A_HO9PsLxw8_0),.clk(gclk));
	jdff dff_A_xFSUe6E94_0(.dout(w_dff_A_lC6Hynj40_0),.din(w_dff_A_xFSUe6E94_0),.clk(gclk));
	jdff dff_A_lC6Hynj40_0(.dout(w_dff_A_uRT7JYxG0_0),.din(w_dff_A_lC6Hynj40_0),.clk(gclk));
	jdff dff_A_uRT7JYxG0_0(.dout(G446gat),.din(w_dff_A_uRT7JYxG0_0),.clk(gclk));
	jdff dff_A_gk8fR03i2_1(.dout(w_dff_A_e47X5IZU5_0),.din(w_dff_A_gk8fR03i2_1),.clk(gclk));
	jdff dff_A_e47X5IZU5_0(.dout(w_dff_A_EfVOVywg4_0),.din(w_dff_A_e47X5IZU5_0),.clk(gclk));
	jdff dff_A_EfVOVywg4_0(.dout(w_dff_A_qcV3iOse3_0),.din(w_dff_A_EfVOVywg4_0),.clk(gclk));
	jdff dff_A_qcV3iOse3_0(.dout(w_dff_A_okgCl0jt8_0),.din(w_dff_A_qcV3iOse3_0),.clk(gclk));
	jdff dff_A_okgCl0jt8_0(.dout(w_dff_A_PK7eK3ZX3_0),.din(w_dff_A_okgCl0jt8_0),.clk(gclk));
	jdff dff_A_PK7eK3ZX3_0(.dout(w_dff_A_FCstpzfG0_0),.din(w_dff_A_PK7eK3ZX3_0),.clk(gclk));
	jdff dff_A_FCstpzfG0_0(.dout(w_dff_A_zNiaWqLi7_0),.din(w_dff_A_FCstpzfG0_0),.clk(gclk));
	jdff dff_A_zNiaWqLi7_0(.dout(w_dff_A_16Ca2n3i1_0),.din(w_dff_A_zNiaWqLi7_0),.clk(gclk));
	jdff dff_A_16Ca2n3i1_0(.dout(w_dff_A_wstXoahf6_0),.din(w_dff_A_16Ca2n3i1_0),.clk(gclk));
	jdff dff_A_wstXoahf6_0(.dout(w_dff_A_tG95oNRl6_0),.din(w_dff_A_wstXoahf6_0),.clk(gclk));
	jdff dff_A_tG95oNRl6_0(.dout(w_dff_A_uI4KyswJ8_0),.din(w_dff_A_tG95oNRl6_0),.clk(gclk));
	jdff dff_A_uI4KyswJ8_0(.dout(w_dff_A_DelgB37r1_0),.din(w_dff_A_uI4KyswJ8_0),.clk(gclk));
	jdff dff_A_DelgB37r1_0(.dout(w_dff_A_sqY7QrJQ1_0),.din(w_dff_A_DelgB37r1_0),.clk(gclk));
	jdff dff_A_sqY7QrJQ1_0(.dout(w_dff_A_wdhRcQGc3_0),.din(w_dff_A_sqY7QrJQ1_0),.clk(gclk));
	jdff dff_A_wdhRcQGc3_0(.dout(w_dff_A_skfRXWvu2_0),.din(w_dff_A_wdhRcQGc3_0),.clk(gclk));
	jdff dff_A_skfRXWvu2_0(.dout(w_dff_A_ODTZmUmu6_0),.din(w_dff_A_skfRXWvu2_0),.clk(gclk));
	jdff dff_A_ODTZmUmu6_0(.dout(w_dff_A_JWibhQgc3_0),.din(w_dff_A_ODTZmUmu6_0),.clk(gclk));
	jdff dff_A_JWibhQgc3_0(.dout(w_dff_A_F4Zc1xLN0_0),.din(w_dff_A_JWibhQgc3_0),.clk(gclk));
	jdff dff_A_F4Zc1xLN0_0(.dout(w_dff_A_IUnrGZDz2_0),.din(w_dff_A_F4Zc1xLN0_0),.clk(gclk));
	jdff dff_A_IUnrGZDz2_0(.dout(w_dff_A_uBXI9UD37_0),.din(w_dff_A_IUnrGZDz2_0),.clk(gclk));
	jdff dff_A_uBXI9UD37_0(.dout(w_dff_A_yuZRqyvC1_0),.din(w_dff_A_uBXI9UD37_0),.clk(gclk));
	jdff dff_A_yuZRqyvC1_0(.dout(w_dff_A_g2M7lntS1_0),.din(w_dff_A_yuZRqyvC1_0),.clk(gclk));
	jdff dff_A_g2M7lntS1_0(.dout(w_dff_A_44p5UJvB5_0),.din(w_dff_A_g2M7lntS1_0),.clk(gclk));
	jdff dff_A_44p5UJvB5_0(.dout(w_dff_A_pdQtL1Zb0_0),.din(w_dff_A_44p5UJvB5_0),.clk(gclk));
	jdff dff_A_pdQtL1Zb0_0(.dout(w_dff_A_JPt2ryYJ4_0),.din(w_dff_A_pdQtL1Zb0_0),.clk(gclk));
	jdff dff_A_JPt2ryYJ4_0(.dout(G447gat),.din(w_dff_A_JPt2ryYJ4_0),.clk(gclk));
	jdff dff_A_z8F8E7fH6_2(.dout(w_dff_A_N6tYl2Vm4_0),.din(w_dff_A_z8F8E7fH6_2),.clk(gclk));
	jdff dff_A_N6tYl2Vm4_0(.dout(w_dff_A_itiq37yH1_0),.din(w_dff_A_N6tYl2Vm4_0),.clk(gclk));
	jdff dff_A_itiq37yH1_0(.dout(w_dff_A_EklhlN0Z8_0),.din(w_dff_A_itiq37yH1_0),.clk(gclk));
	jdff dff_A_EklhlN0Z8_0(.dout(w_dff_A_yliVfoSD3_0),.din(w_dff_A_EklhlN0Z8_0),.clk(gclk));
	jdff dff_A_yliVfoSD3_0(.dout(w_dff_A_3a6PNsEi4_0),.din(w_dff_A_yliVfoSD3_0),.clk(gclk));
	jdff dff_A_3a6PNsEi4_0(.dout(w_dff_A_tYRR5tEV3_0),.din(w_dff_A_3a6PNsEi4_0),.clk(gclk));
	jdff dff_A_tYRR5tEV3_0(.dout(w_dff_A_cDdU84Np2_0),.din(w_dff_A_tYRR5tEV3_0),.clk(gclk));
	jdff dff_A_cDdU84Np2_0(.dout(w_dff_A_iuFlyMMf6_0),.din(w_dff_A_cDdU84Np2_0),.clk(gclk));
	jdff dff_A_iuFlyMMf6_0(.dout(w_dff_A_T3FUjRtb4_0),.din(w_dff_A_iuFlyMMf6_0),.clk(gclk));
	jdff dff_A_T3FUjRtb4_0(.dout(w_dff_A_PCnx4Ua85_0),.din(w_dff_A_T3FUjRtb4_0),.clk(gclk));
	jdff dff_A_PCnx4Ua85_0(.dout(w_dff_A_PihY6KjF4_0),.din(w_dff_A_PCnx4Ua85_0),.clk(gclk));
	jdff dff_A_PihY6KjF4_0(.dout(w_dff_A_YT5GUfvM0_0),.din(w_dff_A_PihY6KjF4_0),.clk(gclk));
	jdff dff_A_YT5GUfvM0_0(.dout(w_dff_A_qoEQlI4f8_0),.din(w_dff_A_YT5GUfvM0_0),.clk(gclk));
	jdff dff_A_qoEQlI4f8_0(.dout(w_dff_A_abDVmSIk8_0),.din(w_dff_A_qoEQlI4f8_0),.clk(gclk));
	jdff dff_A_abDVmSIk8_0(.dout(w_dff_A_FtgM57jl7_0),.din(w_dff_A_abDVmSIk8_0),.clk(gclk));
	jdff dff_A_FtgM57jl7_0(.dout(w_dff_A_vz1tj4NN9_0),.din(w_dff_A_FtgM57jl7_0),.clk(gclk));
	jdff dff_A_vz1tj4NN9_0(.dout(w_dff_A_G2Bulu845_0),.din(w_dff_A_vz1tj4NN9_0),.clk(gclk));
	jdff dff_A_G2Bulu845_0(.dout(w_dff_A_1Vq4zG4Y3_0),.din(w_dff_A_G2Bulu845_0),.clk(gclk));
	jdff dff_A_1Vq4zG4Y3_0(.dout(w_dff_A_H57ICmdt0_0),.din(w_dff_A_1Vq4zG4Y3_0),.clk(gclk));
	jdff dff_A_H57ICmdt0_0(.dout(w_dff_A_qWBwVJn27_0),.din(w_dff_A_H57ICmdt0_0),.clk(gclk));
	jdff dff_A_qWBwVJn27_0(.dout(w_dff_A_ySES4hWu9_0),.din(w_dff_A_qWBwVJn27_0),.clk(gclk));
	jdff dff_A_ySES4hWu9_0(.dout(w_dff_A_du7yM5w39_0),.din(w_dff_A_ySES4hWu9_0),.clk(gclk));
	jdff dff_A_du7yM5w39_0(.dout(G448gat),.din(w_dff_A_du7yM5w39_0),.clk(gclk));
	jdff dff_A_35UzA5Ss9_2(.dout(w_dff_A_0Ptgjekn0_0),.din(w_dff_A_35UzA5Ss9_2),.clk(gclk));
	jdff dff_A_0Ptgjekn0_0(.dout(w_dff_A_j8Ii4hMS8_0),.din(w_dff_A_0Ptgjekn0_0),.clk(gclk));
	jdff dff_A_j8Ii4hMS8_0(.dout(w_dff_A_lM2R0Pch0_0),.din(w_dff_A_j8Ii4hMS8_0),.clk(gclk));
	jdff dff_A_lM2R0Pch0_0(.dout(w_dff_A_j84R6Ve84_0),.din(w_dff_A_lM2R0Pch0_0),.clk(gclk));
	jdff dff_A_j84R6Ve84_0(.dout(w_dff_A_Mv0tkdQm6_0),.din(w_dff_A_j84R6Ve84_0),.clk(gclk));
	jdff dff_A_Mv0tkdQm6_0(.dout(w_dff_A_77Fev5oC7_0),.din(w_dff_A_Mv0tkdQm6_0),.clk(gclk));
	jdff dff_A_77Fev5oC7_0(.dout(w_dff_A_1b5cLdGh4_0),.din(w_dff_A_77Fev5oC7_0),.clk(gclk));
	jdff dff_A_1b5cLdGh4_0(.dout(w_dff_A_diSnmqkp3_0),.din(w_dff_A_1b5cLdGh4_0),.clk(gclk));
	jdff dff_A_diSnmqkp3_0(.dout(w_dff_A_q84iModq4_0),.din(w_dff_A_diSnmqkp3_0),.clk(gclk));
	jdff dff_A_q84iModq4_0(.dout(w_dff_A_AwWNJQoM4_0),.din(w_dff_A_q84iModq4_0),.clk(gclk));
	jdff dff_A_AwWNJQoM4_0(.dout(w_dff_A_2uFWQlNp4_0),.din(w_dff_A_AwWNJQoM4_0),.clk(gclk));
	jdff dff_A_2uFWQlNp4_0(.dout(w_dff_A_ELE8zD7S1_0),.din(w_dff_A_2uFWQlNp4_0),.clk(gclk));
	jdff dff_A_ELE8zD7S1_0(.dout(w_dff_A_4BXwUa9W2_0),.din(w_dff_A_ELE8zD7S1_0),.clk(gclk));
	jdff dff_A_4BXwUa9W2_0(.dout(w_dff_A_shJNXAUR0_0),.din(w_dff_A_4BXwUa9W2_0),.clk(gclk));
	jdff dff_A_shJNXAUR0_0(.dout(w_dff_A_vK0pB3BG3_0),.din(w_dff_A_shJNXAUR0_0),.clk(gclk));
	jdff dff_A_vK0pB3BG3_0(.dout(w_dff_A_IakdHtb17_0),.din(w_dff_A_vK0pB3BG3_0),.clk(gclk));
	jdff dff_A_IakdHtb17_0(.dout(w_dff_A_i2CTfwHc6_0),.din(w_dff_A_IakdHtb17_0),.clk(gclk));
	jdff dff_A_i2CTfwHc6_0(.dout(w_dff_A_8OXctc0o6_0),.din(w_dff_A_i2CTfwHc6_0),.clk(gclk));
	jdff dff_A_8OXctc0o6_0(.dout(w_dff_A_k0UJc8H90_0),.din(w_dff_A_8OXctc0o6_0),.clk(gclk));
	jdff dff_A_k0UJc8H90_0(.dout(w_dff_A_y1D5oWcT5_0),.din(w_dff_A_k0UJc8H90_0),.clk(gclk));
	jdff dff_A_y1D5oWcT5_0(.dout(w_dff_A_YUq6vmec7_0),.din(w_dff_A_y1D5oWcT5_0),.clk(gclk));
	jdff dff_A_YUq6vmec7_0(.dout(w_dff_A_LXlVsLMV9_0),.din(w_dff_A_YUq6vmec7_0),.clk(gclk));
	jdff dff_A_LXlVsLMV9_0(.dout(G449gat),.din(w_dff_A_LXlVsLMV9_0),.clk(gclk));
	jdff dff_A_Cm3FyGve2_2(.dout(w_dff_A_31Ad5Iot4_0),.din(w_dff_A_Cm3FyGve2_2),.clk(gclk));
	jdff dff_A_31Ad5Iot4_0(.dout(w_dff_A_NfA965aN3_0),.din(w_dff_A_31Ad5Iot4_0),.clk(gclk));
	jdff dff_A_NfA965aN3_0(.dout(w_dff_A_G58gEOws6_0),.din(w_dff_A_NfA965aN3_0),.clk(gclk));
	jdff dff_A_G58gEOws6_0(.dout(w_dff_A_IU2e1hUv2_0),.din(w_dff_A_G58gEOws6_0),.clk(gclk));
	jdff dff_A_IU2e1hUv2_0(.dout(w_dff_A_KOZq2ZvW6_0),.din(w_dff_A_IU2e1hUv2_0),.clk(gclk));
	jdff dff_A_KOZq2ZvW6_0(.dout(w_dff_A_joH00s858_0),.din(w_dff_A_KOZq2ZvW6_0),.clk(gclk));
	jdff dff_A_joH00s858_0(.dout(w_dff_A_8lFmZ9hw9_0),.din(w_dff_A_joH00s858_0),.clk(gclk));
	jdff dff_A_8lFmZ9hw9_0(.dout(w_dff_A_iRdDOUiF8_0),.din(w_dff_A_8lFmZ9hw9_0),.clk(gclk));
	jdff dff_A_iRdDOUiF8_0(.dout(w_dff_A_zuCDbIFm5_0),.din(w_dff_A_iRdDOUiF8_0),.clk(gclk));
	jdff dff_A_zuCDbIFm5_0(.dout(w_dff_A_7cCx4HiP1_0),.din(w_dff_A_zuCDbIFm5_0),.clk(gclk));
	jdff dff_A_7cCx4HiP1_0(.dout(w_dff_A_9OOROhO05_0),.din(w_dff_A_7cCx4HiP1_0),.clk(gclk));
	jdff dff_A_9OOROhO05_0(.dout(w_dff_A_IcCDwTRV7_0),.din(w_dff_A_9OOROhO05_0),.clk(gclk));
	jdff dff_A_IcCDwTRV7_0(.dout(w_dff_A_DQ4gr52g4_0),.din(w_dff_A_IcCDwTRV7_0),.clk(gclk));
	jdff dff_A_DQ4gr52g4_0(.dout(w_dff_A_XRm1YKov8_0),.din(w_dff_A_DQ4gr52g4_0),.clk(gclk));
	jdff dff_A_XRm1YKov8_0(.dout(w_dff_A_htqpJaBP0_0),.din(w_dff_A_XRm1YKov8_0),.clk(gclk));
	jdff dff_A_htqpJaBP0_0(.dout(w_dff_A_ZLO8NrNs5_0),.din(w_dff_A_htqpJaBP0_0),.clk(gclk));
	jdff dff_A_ZLO8NrNs5_0(.dout(w_dff_A_xE0I3a5k5_0),.din(w_dff_A_ZLO8NrNs5_0),.clk(gclk));
	jdff dff_A_xE0I3a5k5_0(.dout(w_dff_A_12k9JVQK0_0),.din(w_dff_A_xE0I3a5k5_0),.clk(gclk));
	jdff dff_A_12k9JVQK0_0(.dout(w_dff_A_e9byq4wk7_0),.din(w_dff_A_12k9JVQK0_0),.clk(gclk));
	jdff dff_A_e9byq4wk7_0(.dout(w_dff_A_1dRJWU1m6_0),.din(w_dff_A_e9byq4wk7_0),.clk(gclk));
	jdff dff_A_1dRJWU1m6_0(.dout(w_dff_A_tmHVEUtT4_0),.din(w_dff_A_1dRJWU1m6_0),.clk(gclk));
	jdff dff_A_tmHVEUtT4_0(.dout(w_dff_A_6ZSNF53G6_0),.din(w_dff_A_tmHVEUtT4_0),.clk(gclk));
	jdff dff_A_6ZSNF53G6_0(.dout(w_dff_A_JkHaEiYN3_0),.din(w_dff_A_6ZSNF53G6_0),.clk(gclk));
	jdff dff_A_JkHaEiYN3_0(.dout(w_dff_A_OrUcK1n14_0),.din(w_dff_A_JkHaEiYN3_0),.clk(gclk));
	jdff dff_A_OrUcK1n14_0(.dout(w_dff_A_yBV16ocd2_0),.din(w_dff_A_OrUcK1n14_0),.clk(gclk));
	jdff dff_A_yBV16ocd2_0(.dout(G450gat),.din(w_dff_A_yBV16ocd2_0),.clk(gclk));
	jdff dff_A_Tfh5LF372_2(.dout(w_dff_A_uPvHRNLG3_0),.din(w_dff_A_Tfh5LF372_2),.clk(gclk));
	jdff dff_A_uPvHRNLG3_0(.dout(w_dff_A_Uy02UmIo8_0),.din(w_dff_A_uPvHRNLG3_0),.clk(gclk));
	jdff dff_A_Uy02UmIo8_0(.dout(w_dff_A_m1Vt2YBx6_0),.din(w_dff_A_Uy02UmIo8_0),.clk(gclk));
	jdff dff_A_m1Vt2YBx6_0(.dout(w_dff_A_dyAkftY82_0),.din(w_dff_A_m1Vt2YBx6_0),.clk(gclk));
	jdff dff_A_dyAkftY82_0(.dout(w_dff_A_D53pIOFt5_0),.din(w_dff_A_dyAkftY82_0),.clk(gclk));
	jdff dff_A_D53pIOFt5_0(.dout(w_dff_A_CvzpfV0D9_0),.din(w_dff_A_D53pIOFt5_0),.clk(gclk));
	jdff dff_A_CvzpfV0D9_0(.dout(w_dff_A_ZoPtnveL5_0),.din(w_dff_A_CvzpfV0D9_0),.clk(gclk));
	jdff dff_A_ZoPtnveL5_0(.dout(w_dff_A_WPlGyvyq0_0),.din(w_dff_A_ZoPtnveL5_0),.clk(gclk));
	jdff dff_A_WPlGyvyq0_0(.dout(w_dff_A_JKOIBxQq9_0),.din(w_dff_A_WPlGyvyq0_0),.clk(gclk));
	jdff dff_A_JKOIBxQq9_0(.dout(w_dff_A_u1It9b1q6_0),.din(w_dff_A_JKOIBxQq9_0),.clk(gclk));
	jdff dff_A_u1It9b1q6_0(.dout(w_dff_A_oRS2jfnE2_0),.din(w_dff_A_u1It9b1q6_0),.clk(gclk));
	jdff dff_A_oRS2jfnE2_0(.dout(w_dff_A_niqioGRP2_0),.din(w_dff_A_oRS2jfnE2_0),.clk(gclk));
	jdff dff_A_niqioGRP2_0(.dout(w_dff_A_NSirViKM5_0),.din(w_dff_A_niqioGRP2_0),.clk(gclk));
	jdff dff_A_NSirViKM5_0(.dout(w_dff_A_YHqalQIW2_0),.din(w_dff_A_NSirViKM5_0),.clk(gclk));
	jdff dff_A_YHqalQIW2_0(.dout(w_dff_A_gnDyFYLu4_0),.din(w_dff_A_YHqalQIW2_0),.clk(gclk));
	jdff dff_A_gnDyFYLu4_0(.dout(w_dff_A_dPSSX9k19_0),.din(w_dff_A_gnDyFYLu4_0),.clk(gclk));
	jdff dff_A_dPSSX9k19_0(.dout(w_dff_A_vIuqw2K54_0),.din(w_dff_A_dPSSX9k19_0),.clk(gclk));
	jdff dff_A_vIuqw2K54_0(.dout(w_dff_A_SoKFsxUJ2_0),.din(w_dff_A_vIuqw2K54_0),.clk(gclk));
	jdff dff_A_SoKFsxUJ2_0(.dout(w_dff_A_DrjcHeE33_0),.din(w_dff_A_SoKFsxUJ2_0),.clk(gclk));
	jdff dff_A_DrjcHeE33_0(.dout(w_dff_A_hopkUYEs1_0),.din(w_dff_A_DrjcHeE33_0),.clk(gclk));
	jdff dff_A_hopkUYEs1_0(.dout(w_dff_A_EAjv4duJ1_0),.din(w_dff_A_hopkUYEs1_0),.clk(gclk));
	jdff dff_A_EAjv4duJ1_0(.dout(w_dff_A_zz2fzF9F7_0),.din(w_dff_A_EAjv4duJ1_0),.clk(gclk));
	jdff dff_A_zz2fzF9F7_0(.dout(w_dff_A_0wNKKP4D7_0),.din(w_dff_A_zz2fzF9F7_0),.clk(gclk));
	jdff dff_A_0wNKKP4D7_0(.dout(G767gat),.din(w_dff_A_0wNKKP4D7_0),.clk(gclk));
	jdff dff_A_9HXCWLs03_2(.dout(w_dff_A_Zvi0FnSB8_0),.din(w_dff_A_9HXCWLs03_2),.clk(gclk));
	jdff dff_A_Zvi0FnSB8_0(.dout(w_dff_A_MTai2li04_0),.din(w_dff_A_Zvi0FnSB8_0),.clk(gclk));
	jdff dff_A_MTai2li04_0(.dout(w_dff_A_ZxCGqh3S5_0),.din(w_dff_A_MTai2li04_0),.clk(gclk));
	jdff dff_A_ZxCGqh3S5_0(.dout(w_dff_A_KBHhX25z7_0),.din(w_dff_A_ZxCGqh3S5_0),.clk(gclk));
	jdff dff_A_KBHhX25z7_0(.dout(w_dff_A_ygILS7ks5_0),.din(w_dff_A_KBHhX25z7_0),.clk(gclk));
	jdff dff_A_ygILS7ks5_0(.dout(w_dff_A_mXZT9Yf57_0),.din(w_dff_A_ygILS7ks5_0),.clk(gclk));
	jdff dff_A_mXZT9Yf57_0(.dout(w_dff_A_w9f46bQM2_0),.din(w_dff_A_mXZT9Yf57_0),.clk(gclk));
	jdff dff_A_w9f46bQM2_0(.dout(w_dff_A_aUqLlwpE2_0),.din(w_dff_A_w9f46bQM2_0),.clk(gclk));
	jdff dff_A_aUqLlwpE2_0(.dout(w_dff_A_RXQZh2Bh6_0),.din(w_dff_A_aUqLlwpE2_0),.clk(gclk));
	jdff dff_A_RXQZh2Bh6_0(.dout(w_dff_A_FKsLlO5G5_0),.din(w_dff_A_RXQZh2Bh6_0),.clk(gclk));
	jdff dff_A_FKsLlO5G5_0(.dout(w_dff_A_YFaKUnug7_0),.din(w_dff_A_FKsLlO5G5_0),.clk(gclk));
	jdff dff_A_YFaKUnug7_0(.dout(w_dff_A_FKUAsMtU8_0),.din(w_dff_A_YFaKUnug7_0),.clk(gclk));
	jdff dff_A_FKUAsMtU8_0(.dout(w_dff_A_dBQoEy1P7_0),.din(w_dff_A_FKUAsMtU8_0),.clk(gclk));
	jdff dff_A_dBQoEy1P7_0(.dout(w_dff_A_mshbxTQ17_0),.din(w_dff_A_dBQoEy1P7_0),.clk(gclk));
	jdff dff_A_mshbxTQ17_0(.dout(w_dff_A_RyOrPpx31_0),.din(w_dff_A_mshbxTQ17_0),.clk(gclk));
	jdff dff_A_RyOrPpx31_0(.dout(w_dff_A_wGDEOBAO3_0),.din(w_dff_A_RyOrPpx31_0),.clk(gclk));
	jdff dff_A_wGDEOBAO3_0(.dout(w_dff_A_7ZHxunlr6_0),.din(w_dff_A_wGDEOBAO3_0),.clk(gclk));
	jdff dff_A_7ZHxunlr6_0(.dout(w_dff_A_EofVAvGa0_0),.din(w_dff_A_7ZHxunlr6_0),.clk(gclk));
	jdff dff_A_EofVAvGa0_0(.dout(w_dff_A_5ccZHtLU6_0),.din(w_dff_A_EofVAvGa0_0),.clk(gclk));
	jdff dff_A_5ccZHtLU6_0(.dout(w_dff_A_IpKG5eOQ7_0),.din(w_dff_A_5ccZHtLU6_0),.clk(gclk));
	jdff dff_A_IpKG5eOQ7_0(.dout(w_dff_A_MLPK6q7u3_0),.din(w_dff_A_IpKG5eOQ7_0),.clk(gclk));
	jdff dff_A_MLPK6q7u3_0(.dout(w_dff_A_jKRHPVkF7_0),.din(w_dff_A_MLPK6q7u3_0),.clk(gclk));
	jdff dff_A_jKRHPVkF7_0(.dout(w_dff_A_baKIWzB34_0),.din(w_dff_A_jKRHPVkF7_0),.clk(gclk));
	jdff dff_A_baKIWzB34_0(.dout(G768gat),.din(w_dff_A_baKIWzB34_0),.clk(gclk));
	jdff dff_A_XpWbAcL04_2(.dout(w_dff_A_2Gn6GIy29_0),.din(w_dff_A_XpWbAcL04_2),.clk(gclk));
	jdff dff_A_2Gn6GIy29_0(.dout(w_dff_A_1lALqmkr3_0),.din(w_dff_A_2Gn6GIy29_0),.clk(gclk));
	jdff dff_A_1lALqmkr3_0(.dout(w_dff_A_8swZOnoU1_0),.din(w_dff_A_1lALqmkr3_0),.clk(gclk));
	jdff dff_A_8swZOnoU1_0(.dout(w_dff_A_QEaCdejI2_0),.din(w_dff_A_8swZOnoU1_0),.clk(gclk));
	jdff dff_A_QEaCdejI2_0(.dout(w_dff_A_yFJ7F2XZ4_0),.din(w_dff_A_QEaCdejI2_0),.clk(gclk));
	jdff dff_A_yFJ7F2XZ4_0(.dout(w_dff_A_uY6qbbZk2_0),.din(w_dff_A_yFJ7F2XZ4_0),.clk(gclk));
	jdff dff_A_uY6qbbZk2_0(.dout(w_dff_A_YgoEzABX5_0),.din(w_dff_A_uY6qbbZk2_0),.clk(gclk));
	jdff dff_A_YgoEzABX5_0(.dout(w_dff_A_erC9KmhN4_0),.din(w_dff_A_YgoEzABX5_0),.clk(gclk));
	jdff dff_A_erC9KmhN4_0(.dout(w_dff_A_zu3e41Xj6_0),.din(w_dff_A_erC9KmhN4_0),.clk(gclk));
	jdff dff_A_zu3e41Xj6_0(.dout(w_dff_A_qz7hHSpY3_0),.din(w_dff_A_zu3e41Xj6_0),.clk(gclk));
	jdff dff_A_qz7hHSpY3_0(.dout(w_dff_A_NyZhUtfT3_0),.din(w_dff_A_qz7hHSpY3_0),.clk(gclk));
	jdff dff_A_NyZhUtfT3_0(.dout(w_dff_A_qbDNvsOO4_0),.din(w_dff_A_NyZhUtfT3_0),.clk(gclk));
	jdff dff_A_qbDNvsOO4_0(.dout(G850gat),.din(w_dff_A_qbDNvsOO4_0),.clk(gclk));
	jdff dff_A_4HrvKHDq8_2(.dout(w_dff_A_ZTkAA7oB6_0),.din(w_dff_A_4HrvKHDq8_2),.clk(gclk));
	jdff dff_A_ZTkAA7oB6_0(.dout(w_dff_A_bbsihPsa0_0),.din(w_dff_A_ZTkAA7oB6_0),.clk(gclk));
	jdff dff_A_bbsihPsa0_0(.dout(w_dff_A_Ouqn9SIP4_0),.din(w_dff_A_bbsihPsa0_0),.clk(gclk));
	jdff dff_A_Ouqn9SIP4_0(.dout(w_dff_A_MDe9hBTy5_0),.din(w_dff_A_Ouqn9SIP4_0),.clk(gclk));
	jdff dff_A_MDe9hBTy5_0(.dout(w_dff_A_FmKbmgVM8_0),.din(w_dff_A_MDe9hBTy5_0),.clk(gclk));
	jdff dff_A_FmKbmgVM8_0(.dout(w_dff_A_a3cHNdpE2_0),.din(w_dff_A_FmKbmgVM8_0),.clk(gclk));
	jdff dff_A_a3cHNdpE2_0(.dout(w_dff_A_BvwwH1tn7_0),.din(w_dff_A_a3cHNdpE2_0),.clk(gclk));
	jdff dff_A_BvwwH1tn7_0(.dout(G863gat),.din(w_dff_A_BvwwH1tn7_0),.clk(gclk));
	jdff dff_A_UT8qrq8w4_2(.dout(w_dff_A_Z7zdoE9J2_0),.din(w_dff_A_UT8qrq8w4_2),.clk(gclk));
	jdff dff_A_Z7zdoE9J2_0(.dout(w_dff_A_GF43g0tL7_0),.din(w_dff_A_Z7zdoE9J2_0),.clk(gclk));
	jdff dff_A_GF43g0tL7_0(.dout(w_dff_A_GSg1tmyc9_0),.din(w_dff_A_GF43g0tL7_0),.clk(gclk));
	jdff dff_A_GSg1tmyc9_0(.dout(w_dff_A_jyqkSZWD5_0),.din(w_dff_A_GSg1tmyc9_0),.clk(gclk));
	jdff dff_A_jyqkSZWD5_0(.dout(w_dff_A_NO5UTTHf5_0),.din(w_dff_A_jyqkSZWD5_0),.clk(gclk));
	jdff dff_A_NO5UTTHf5_0(.dout(w_dff_A_U0i1pmL48_0),.din(w_dff_A_NO5UTTHf5_0),.clk(gclk));
	jdff dff_A_U0i1pmL48_0(.dout(w_dff_A_wpYFfFYg9_0),.din(w_dff_A_U0i1pmL48_0),.clk(gclk));
	jdff dff_A_wpYFfFYg9_0(.dout(w_dff_A_xOVi91633_0),.din(w_dff_A_wpYFfFYg9_0),.clk(gclk));
	jdff dff_A_xOVi91633_0(.dout(w_dff_A_xxYGU16b4_0),.din(w_dff_A_xOVi91633_0),.clk(gclk));
	jdff dff_A_xxYGU16b4_0(.dout(G864gat),.din(w_dff_A_xxYGU16b4_0),.clk(gclk));
	jdff dff_A_iVhb6Mw44_2(.dout(w_dff_A_SKTtECSv5_0),.din(w_dff_A_iVhb6Mw44_2),.clk(gclk));
	jdff dff_A_SKTtECSv5_0(.dout(w_dff_A_ztrwt2oI9_0),.din(w_dff_A_SKTtECSv5_0),.clk(gclk));
	jdff dff_A_ztrwt2oI9_0(.dout(w_dff_A_gJ1UJKoo7_0),.din(w_dff_A_ztrwt2oI9_0),.clk(gclk));
	jdff dff_A_gJ1UJKoo7_0(.dout(w_dff_A_zMBmsAcS3_0),.din(w_dff_A_gJ1UJKoo7_0),.clk(gclk));
	jdff dff_A_zMBmsAcS3_0(.dout(w_dff_A_Ur4qw2Wy9_0),.din(w_dff_A_zMBmsAcS3_0),.clk(gclk));
	jdff dff_A_Ur4qw2Wy9_0(.dout(w_dff_A_ekL7g0Qy7_0),.din(w_dff_A_Ur4qw2Wy9_0),.clk(gclk));
	jdff dff_A_ekL7g0Qy7_0(.dout(w_dff_A_s7lnhHck6_0),.din(w_dff_A_ekL7g0Qy7_0),.clk(gclk));
	jdff dff_A_s7lnhHck6_0(.dout(w_dff_A_QtxOKwNC8_0),.din(w_dff_A_s7lnhHck6_0),.clk(gclk));
	jdff dff_A_QtxOKwNC8_0(.dout(w_dff_A_fFR7xMcQ5_0),.din(w_dff_A_QtxOKwNC8_0),.clk(gclk));
	jdff dff_A_fFR7xMcQ5_0(.dout(w_dff_A_Z7sUUe0q7_0),.din(w_dff_A_fFR7xMcQ5_0),.clk(gclk));
	jdff dff_A_Z7sUUe0q7_0(.dout(w_dff_A_mDhjMDqr1_0),.din(w_dff_A_Z7sUUe0q7_0),.clk(gclk));
	jdff dff_A_mDhjMDqr1_0(.dout(G865gat),.din(w_dff_A_mDhjMDqr1_0),.clk(gclk));
	jdff dff_A_WiHHet6v3_2(.dout(w_dff_A_XWW50pqM5_0),.din(w_dff_A_WiHHet6v3_2),.clk(gclk));
	jdff dff_A_XWW50pqM5_0(.dout(G866gat),.din(w_dff_A_XWW50pqM5_0),.clk(gclk));
	jdff dff_A_xA640cQm0_2(.dout(w_dff_A_qV1VhWRJ7_0),.din(w_dff_A_xA640cQm0_2),.clk(gclk));
	jdff dff_A_qV1VhWRJ7_0(.dout(w_dff_A_SJQjbrIe3_0),.din(w_dff_A_qV1VhWRJ7_0),.clk(gclk));
	jdff dff_A_SJQjbrIe3_0(.dout(w_dff_A_AdgVd7bd8_0),.din(w_dff_A_SJQjbrIe3_0),.clk(gclk));
	jdff dff_A_AdgVd7bd8_0(.dout(w_dff_A_cXd4Sbxm0_0),.din(w_dff_A_AdgVd7bd8_0),.clk(gclk));
	jdff dff_A_cXd4Sbxm0_0(.dout(G874gat),.din(w_dff_A_cXd4Sbxm0_0),.clk(gclk));
	jdff dff_A_0JlrbuTL8_2(.dout(w_dff_A_esbwER353_0),.din(w_dff_A_0JlrbuTL8_2),.clk(gclk));
	jdff dff_A_esbwER353_0(.dout(G879gat),.din(w_dff_A_esbwER353_0),.clk(gclk));
	jdff dff_A_y8Z8qDZW3_2(.dout(w_dff_A_ZHQ0hDa74_0),.din(w_dff_A_y8Z8qDZW3_2),.clk(gclk));
	jdff dff_A_ZHQ0hDa74_0(.dout(w_dff_A_16jvoNja6_0),.din(w_dff_A_ZHQ0hDa74_0),.clk(gclk));
	jdff dff_A_16jvoNja6_0(.dout(w_dff_A_vchR78ye5_0),.din(w_dff_A_16jvoNja6_0),.clk(gclk));
	jdff dff_A_vchR78ye5_0(.dout(G880gat),.din(w_dff_A_vchR78ye5_0),.clk(gclk));
endmodule

