module rf_c880(G268gat, G267gat, G111gat, G87gat, G130gat, G159gat, G261gat, G101gat, G152gat, G86gat, G29gat, G13gat, G106gat, G74gat, G96gat, G91gat, G149gat, G73gat, G80gat, G138gat, G72gat, G90gat, G8gat, G51gat, G143gat, G26gat, G55gat, G36gat, G153gat, G17gat, G246gat, G85gat, G59gat, G116gat, G121gat, G146gat, G126gat, G135gat, G89gat, G219gat, G68gat, G156gat, G165gat, G42gat, G171gat, G177gat, G195gat, G259gat, G183gat, G88gat, G189gat, G210gat, G237gat, G201gat, G75gat, G1gat, G207gat, G228gat, G255gat, G260gat, G879gat, G878gat, G874gat, G865gat, G864gat, G767gat, G450gat, G423gat, G850gat, G389gat, G390gat, G447gat, G880gat, G449gat, G391gat, G418gat, G863gat, G419gat, G768gat, G422gat, G420gat, G421gat, G448gat, G866gat, G388gat, G446gat);
    input G268gat, G267gat, G111gat, G87gat, G130gat, G159gat, G261gat, G101gat, G152gat, G86gat, G29gat, G13gat, G106gat, G74gat, G96gat, G91gat, G149gat, G73gat, G80gat, G138gat, G72gat, G90gat, G8gat, G51gat, G143gat, G26gat, G55gat, G36gat, G153gat, G17gat, G246gat, G85gat, G59gat, G116gat, G121gat, G146gat, G126gat, G135gat, G89gat, G219gat, G68gat, G156gat, G165gat, G42gat, G171gat, G177gat, G195gat, G259gat, G183gat, G88gat, G189gat, G210gat, G237gat, G201gat, G75gat, G1gat, G207gat, G228gat, G255gat, G260gat;
    output G879gat, G878gat, G874gat, G865gat, G864gat, G767gat, G450gat, G423gat, G850gat, G389gat, G390gat, G447gat, G880gat, G449gat, G391gat, G418gat, G863gat, G419gat, G768gat, G422gat, G420gat, G421gat, G448gat, G866gat, G388gat, G446gat;
    wire n89;
    wire n93;
    wire n97;
    wire n101;
    wire n105;
    wire n109;
    wire n113;
    wire n117;
    wire n121;
    wire n124;
    wire n127;
    wire n130;
    wire n134;
    wire n138;
    wire n142;
    wire n145;
    wire n149;
    wire n152;
    wire n156;
    wire n159;
    wire n162;
    wire n166;
    wire n170;
    wire n173;
    wire n177;
    wire n181;
    wire n185;
    wire n188;
    wire n192;
    wire n196;
    wire n200;
    wire n204;
    wire n208;
    wire n212;
    wire n216;
    wire n220;
    wire n224;
    wire n228;
    wire n232;
    wire n236;
    wire n240;
    wire n244;
    wire n248;
    wire n252;
    wire n256;
    wire n260;
    wire n264;
    wire n268;
    wire n272;
    wire n276;
    wire n280;
    wire n284;
    wire n288;
    wire n292;
    wire n296;
    wire n300;
    wire n304;
    wire n307;
    wire n311;
    wire n314;
    wire n318;
    wire n322;
    wire n326;
    wire n330;
    wire n334;
    wire n338;
    wire n342;
    wire n346;
    wire n350;
    wire n353;
    wire n357;
    wire n361;
    wire n365;
    wire n369;
    wire n373;
    wire n377;
    wire n381;
    wire n384;
    wire n388;
    wire n392;
    wire n396;
    wire n400;
    wire n404;
    wire n407;
    wire n411;
    wire n415;
    wire n419;
    wire n423;
    wire n427;
    wire n431;
    wire n435;
    wire n439;
    wire n443;
    wire n447;
    wire n451;
    wire n455;
    wire n459;
    wire n463;
    wire n467;
    wire n471;
    wire n475;
    wire n479;
    wire n483;
    wire n487;
    wire n491;
    wire n495;
    wire n499;
    wire n503;
    wire n507;
    wire n510;
    wire n514;
    wire n517;
    wire n520;
    wire n523;
    wire n526;
    wire n529;
    wire n532;
    wire n536;
    wire n540;
    wire n544;
    wire n548;
    wire n552;
    wire n555;
    wire n559;
    wire n563;
    wire n567;
    wire n571;
    wire n575;
    wire n579;
    wire n583;
    wire n587;
    wire n591;
    wire n595;
    wire n599;
    wire n603;
    wire n607;
    wire n611;
    wire n615;
    wire n619;
    wire n622;
    wire n626;
    wire n630;
    wire n634;
    wire n638;
    wire n642;
    wire n645;
    wire n649;
    wire n653;
    wire n657;
    wire n661;
    wire n665;
    wire n669;
    wire n673;
    wire n677;
    wire n681;
    wire n685;
    wire n689;
    wire n693;
    wire n697;
    wire n701;
    wire n705;
    wire n709;
    wire n713;
    wire n717;
    wire n721;
    wire n725;
    wire n729;
    wire n732;
    wire n736;
    wire n740;
    wire n743;
    wire n747;
    wire n751;
    wire n755;
    wire n759;
    wire n763;
    wire n767;
    wire n771;
    wire n775;
    wire n779;
    wire n783;
    wire n787;
    wire n791;
    wire n795;
    wire n799;
    wire n803;
    wire n807;
    wire n811;
    wire n814;
    wire n818;
    wire n822;
    wire n826;
    wire n830;
    wire n834;
    wire n838;
    wire n842;
    wire n846;
    wire n850;
    wire n854;
    wire n858;
    wire n862;
    wire n866;
    wire n870;
    wire n874;
    wire n878;
    wire n882;
    wire n886;
    wire n890;
    wire n894;
    wire n898;
    wire n902;
    wire n906;
    wire n910;
    wire n914;
    wire n918;
    wire n922;
    wire n926;
    wire n930;
    wire n934;
    wire n938;
    wire n941;
    wire n945;
    wire n949;
    wire n953;
    wire n957;
    wire n961;
    wire n965;
    wire n968;
    wire n972;
    wire n975;
    wire n979;
    wire n983;
    wire n987;
    wire n991;
    wire n995;
    wire n999;
    wire n1003;
    wire n1007;
    wire n1011;
    wire n1015;
    wire n1019;
    wire n1023;
    wire n1027;
    wire n1031;
    wire n1035;
    wire n1039;
    wire n1043;
    wire n1047;
    wire n1051;
    wire n1055;
    wire n1059;
    wire n1063;
    wire n1067;
    wire n1071;
    wire n1075;
    wire n1079;
    wire n1083;
    wire n1086;
    wire n1089;
    wire n1093;
    wire n1097;
    wire n1101;
    wire n1104;
    wire n1108;
    wire n1112;
    wire n1116;
    wire n1120;
    wire n1124;
    wire n1128;
    wire n1132;
    wire n1136;
    wire n1140;
    wire n1144;
    wire n1148;
    wire n1152;
    wire n1156;
    wire n1160;
    wire n1163;
    wire n1167;
    wire n1170;
    wire n1174;
    wire n1178;
    wire n1181;
    wire n1185;
    wire n1189;
    wire n1193;
    wire n1197;
    wire n1201;
    wire n1205;
    wire n1209;
    wire n1213;
    wire n1217;
    wire n1221;
    wire n1225;
    wire n1229;
    wire n1233;
    wire n1241;
    wire n1244;
    wire n1247;
    wire n1250;
    wire n1254;
    wire n1258;
    wire n1262;
    wire n1266;
    wire n1270;
    wire n1274;
    wire n1278;
    wire n1282;
    wire n1286;
    wire n1290;
    wire n1294;
    wire n1298;
    wire n1302;
    wire n1306;
    wire n1310;
    wire n1314;
    wire n1318;
    wire n1326;
    wire n1329;
    wire n1332;
    wire n1335;
    wire n1339;
    wire n1343;
    wire n1347;
    wire n1351;
    wire n1355;
    wire n1359;
    wire n1363;
    wire n1367;
    wire n1371;
    wire n1375;
    wire n1379;
    wire n1383;
    wire n1387;
    wire n1391;
    wire n1395;
    wire n1399;
    wire n1403;
    wire n2021;
    wire n2024;
    wire n2027;
    wire n2029;
    wire n2033;
    wire n2036;
    wire n2039;
    wire n2042;
    wire n2045;
    wire n2048;
    wire n2051;
    wire n2054;
    wire n2057;
    wire n2060;
    wire n2063;
    wire n2066;
    wire n2069;
    wire n2072;
    wire n2075;
    wire n2078;
    wire n2081;
    wire n2084;
    wire n2087;
    wire n2090;
    wire n2093;
    wire n2096;
    wire n2099;
    wire n2101;
    wire n2104;
    wire n2107;
    wire n2110;
    wire n2113;
    wire n2116;
    wire n2119;
    wire n2122;
    wire n2126;
    wire n2129;
    wire n2132;
    wire n2135;
    wire n2138;
    wire n2141;
    wire n2144;
    wire n2147;
    wire n2150;
    wire n2153;
    wire n2156;
    wire n2159;
    wire n2162;
    wire n2165;
    wire n2168;
    wire n2171;
    wire n2174;
    wire n2177;
    wire n2179;
    wire n2182;
    wire n2185;
    wire n2188;
    wire n2192;
    wire n2195;
    wire n2198;
    wire n2201;
    wire n2203;
    wire n2206;
    wire n2209;
    wire n2212;
    wire n2215;
    wire n2218;
    wire n2221;
    wire n2224;
    wire n2227;
    wire n2230;
    wire n2233;
    wire n2236;
    wire n2240;
    wire n2243;
    wire n2246;
    wire n2249;
    wire n2252;
    wire n2255;
    wire n2258;
    wire n2261;
    wire n2264;
    wire n2267;
    wire n2270;
    wire n2273;
    wire n2276;
    wire n2279;
    wire n2282;
    wire n2285;
    wire n2288;
    wire n2291;
    wire n2294;
    wire n2297;
    wire n2300;
    wire n2302;
    wire n2305;
    wire n2308;
    wire n2311;
    wire n2315;
    wire n2318;
    wire n2321;
    wire n2324;
    wire n2327;
    wire n2330;
    wire n2333;
    wire n2336;
    wire n2339;
    wire n2342;
    wire n2345;
    wire n2348;
    wire n2351;
    wire n2354;
    wire n2357;
    wire n2360;
    wire n2363;
    wire n2365;
    wire n2368;
    wire n2372;
    wire n2375;
    wire n2378;
    wire n2381;
    wire n2384;
    wire n2387;
    wire n2390;
    wire n2393;
    wire n2396;
    wire n2399;
    wire n2402;
    wire n2405;
    wire n2408;
    wire n2411;
    wire n2414;
    wire n2417;
    wire n2420;
    wire n2423;
    wire n2426;
    wire n2428;
    wire n2431;
    wire n2434;
    wire n2437;
    wire n2440;
    wire n2443;
    wire n2446;
    wire n2450;
    wire n2453;
    wire n2456;
    wire n2459;
    wire n2462;
    wire n2465;
    wire n2468;
    wire n2471;
    wire n2474;
    wire n2477;
    wire n2480;
    wire n2483;
    wire n2486;
    wire n2489;
    wire n2492;
    wire n2495;
    wire n2498;
    wire n2501;
    wire n2504;
    wire n2506;
    wire n2509;
    wire n2512;
    wire n2515;
    wire n2518;
    wire n2521;
    wire n2524;
    wire n2527;
    wire n2531;
    wire n2534;
    wire n2537;
    wire n2540;
    wire n2543;
    wire n2546;
    wire n2549;
    wire n2551;
    wire n2554;
    wire n2557;
    wire n2560;
    wire n2563;
    wire n2566;
    wire n2569;
    wire n2573;
    wire n2576;
    wire n2579;
    wire n2582;
    wire n2585;
    wire n2588;
    wire n2591;
    wire n2594;
    wire n2597;
    wire n2600;
    wire n2603;
    wire n2606;
    wire n2609;
    wire n2612;
    wire n2615;
    wire n2618;
    wire n2621;
    wire n2624;
    wire n2627;
    wire n2630;
    wire n2633;
    wire n2636;
    wire n2639;
    wire n2642;
    wire n2645;
    wire n2648;
    wire n2651;
    wire n2654;
    wire n2657;
    wire n2660;
    wire n2662;
    wire n2665;
    wire n2668;
    wire n2671;
    wire n2674;
    wire n2677;
    wire n2680;
    wire n2683;
    wire n2686;
    wire n2690;
    wire n2693;
    wire n2696;
    wire n2698;
    wire n2701;
    wire n2704;
    wire n2707;
    wire n2710;
    wire n2713;
    wire n2716;
    wire n2719;
    wire n2722;
    wire n2725;
    wire n2728;
    wire n2731;
    wire n2734;
    wire n2737;
    wire n2740;
    wire n2743;
    wire n2746;
    wire n2749;
    wire n2753;
    wire n2756;
    wire n2759;
    wire n2762;
    wire n2764;
    wire n2767;
    wire n2770;
    wire n2773;
    wire n2777;
    wire n2780;
    wire n2783;
    wire n2786;
    wire n2789;
    wire n2792;
    wire n2795;
    wire n2797;
    wire n2800;
    wire n2803;
    wire n2806;
    wire n2810;
    wire n2813;
    wire n2816;
    wire n2819;
    wire n2822;
    wire n2825;
    wire n2828;
    wire n2831;
    wire n2834;
    wire n2837;
    wire n2840;
    wire n2843;
    wire n2846;
    wire n2849;
    wire n2852;
    wire n2855;
    wire n2858;
    wire n2861;
    wire n2864;
    wire n2867;
    wire n2870;
    wire n2873;
    wire n2876;
    wire n2878;
    wire n2881;
    wire n2884;
    wire n2887;
    wire n2890;
    wire n2894;
    wire n2897;
    wire n2900;
    wire n2903;
    wire n2906;
    wire n2909;
    wire n2912;
    wire n2915;
    wire n2918;
    wire n2921;
    wire n2924;
    wire n2927;
    wire n2930;
    wire n2933;
    wire n2936;
    wire n2939;
    wire n2942;
    wire n2945;
    wire n2948;
    wire n2951;
    wire n2954;
    wire n2957;
    wire n2960;
    wire n2963;
    wire n2966;
    wire n2969;
    wire n2971;
    wire n2974;
    wire n2977;
    wire n2980;
    wire n2983;
    wire n2986;
    wire n2989;
    wire n2992;
    wire n2995;
    wire n2998;
    wire n3001;
    wire n3004;
    wire n3007;
    wire n3011;
    wire n3013;
    wire n3016;
    wire n3019;
    wire n3022;
    wire n3025;
    wire n3028;
    wire n3031;
    wire n3034;
    wire n3037;
    wire n3040;
    wire n3043;
    wire n3046;
    wire n3049;
    wire n3052;
    wire n3055;
    wire n3058;
    wire n3062;
    wire n3065;
    wire n3068;
    wire n3070;
    wire n3073;
    wire n3076;
    wire n3079;
    wire n3082;
    wire n3085;
    wire n3088;
    wire n3091;
    wire n3094;
    wire n3097;
    wire n3100;
    wire n3103;
    wire n3106;
    wire n3109;
    wire n3112;
    wire n3115;
    wire n3118;
    wire n3121;
    wire n3125;
    wire n3128;
    wire n3131;
    wire n3134;
    wire n3137;
    wire n3140;
    wire n3143;
    wire n3146;
    wire n3149;
    wire n3152;
    wire n3155;
    wire n3158;
    wire n3161;
    wire n3164;
    wire n3167;
    wire n3170;
    wire n3172;
    wire n3175;
    wire n3178;
    wire n3181;
    wire n3184;
    wire n3188;
    wire n3190;
    wire n3193;
    wire n3197;
    wire n3200;
    wire n3203;
    wire n3206;
    wire n3209;
    wire n3212;
    wire n3214;
    wire n3218;
    wire n3221;
    wire n3224;
    wire n3227;
    wire n3230;
    wire n3233;
    wire n3236;
    wire n3239;
    wire n3241;
    wire n3244;
    wire n3247;
    wire n3250;
    wire n3253;
    wire n3256;
    wire n3259;
    wire n3262;
    wire n3265;
    wire n3268;
    wire n3272;
    wire n3275;
    wire n3278;
    wire n3281;
    wire n3284;
    wire n3287;
    wire n3290;
    wire n3293;
    wire n3296;
    wire n3299;
    wire n3302;
    wire n3305;
    wire n3308;
    wire n3311;
    wire n3314;
    wire n3317;
    wire n3320;
    wire n3323;
    wire n3326;
    wire n3329;
    wire n3332;
    wire n3335;
    wire n3338;
    wire n3341;
    wire n3344;
    wire n3347;
    wire n3350;
    wire n3353;
    wire n3356;
    wire n3359;
    wire n3362;
    wire n3365;
    wire n3368;
    wire n3371;
    wire n3373;
    wire n3376;
    wire n3379;
    wire n3382;
    wire n3385;
    wire n3388;
    wire n3391;
    wire n3394;
    wire n3397;
    wire n3400;
    wire n3403;
    wire n3406;
    wire n3409;
    wire n3412;
    wire n3416;
    wire n3419;
    wire n3422;
    wire n3425;
    wire n3428;
    wire n3431;
    wire n3434;
    wire n3437;
    wire n3440;
    wire n3443;
    wire n3445;
    wire n3449;
    wire n3451;
    wire n3454;
    wire n3457;
    wire n3460;
    wire n3463;
    wire n3466;
    wire n3469;
    wire n3472;
    wire n3475;
    wire n3478;
    wire n3481;
    wire n3484;
    wire n3487;
    wire n3490;
    wire n3493;
    wire n3496;
    wire n3499;
    wire n3502;
    wire n3505;
    wire n3508;
    wire n3511;
    wire n3514;
    wire n3517;
    wire n3520;
    wire n3523;
    wire n3526;
    wire n3529;
    wire n3532;
    wire n3535;
    wire n3538;
    wire n3541;
    wire n3544;
    wire n3547;
    wire n3550;
    wire n3553;
    wire n3557;
    wire n3559;
    wire n3562;
    wire n3565;
    wire n3569;
    wire n3571;
    wire n3574;
    wire n3577;
    wire n3580;
    wire n3583;
    wire n3586;
    wire n3589;
    wire n3592;
    wire n3595;
    wire n3598;
    wire n3601;
    wire n3604;
    wire n3607;
    wire n3610;
    wire n3613;
    wire n3616;
    wire n3619;
    wire n3623;
    wire n3625;
    wire n3628;
    wire n3631;
    wire n3634;
    wire n3637;
    wire n3640;
    wire n3644;
    wire n3647;
    wire n3650;
    wire n3653;
    wire n3655;
    wire n3658;
    wire n3661;
    wire n3664;
    wire n3667;
    wire n3670;
    wire n3673;
    wire n3676;
    wire n3679;
    wire n3682;
    wire n3685;
    wire n3688;
    wire n3692;
    wire n3695;
    wire n3698;
    wire n3701;
    wire n3704;
    wire n3707;
    wire n3710;
    wire n3713;
    wire n3716;
    wire n3719;
    wire n3722;
    wire n3725;
    wire n3728;
    wire n3731;
    wire n3734;
    wire n3737;
    wire n3740;
    wire n3743;
    wire n3746;
    wire n3749;
    wire n3752;
    wire n3755;
    wire n3758;
    wire n3761;
    wire n3764;
    wire n3767;
    wire n3770;
    wire n3773;
    wire n3776;
    wire n3779;
    wire n3781;
    wire n3784;
    wire n3787;
    wire n3790;
    wire n3793;
    wire n3796;
    wire n3799;
    wire n3802;
    wire n3805;
    wire n3808;
    wire n3811;
    wire n3814;
    wire n3817;
    wire n3820;
    wire n3823;
    wire n3826;
    wire n3829;
    wire n3832;
    wire n3835;
    wire n3838;
    wire n3841;
    wire n3844;
    wire n3847;
    wire n3850;
    wire n3853;
    wire n3856;
    wire n3859;
    wire n3862;
    wire n3865;
    wire n3868;
    wire n3871;
    wire n3874;
    wire n3877;
    wire n3880;
    wire n3883;
    wire n3886;
    wire n3889;
    wire n3892;
    wire n3895;
    wire n3898;
    wire n3901;
    wire n3904;
    wire n3907;
    wire n3910;
    wire n3913;
    wire n3916;
    wire n3919;
    wire n3922;
    wire n3925;
    wire n3928;
    wire n3931;
    wire n3934;
    wire n3937;
    wire n3940;
    wire n3944;
    wire n3946;
    wire n3949;
    wire n3952;
    wire n3955;
    wire n3958;
    wire n3961;
    wire n3964;
    wire n3967;
    wire n3970;
    wire n3973;
    wire n3976;
    wire n3979;
    wire n3982;
    wire n3986;
    wire n3988;
    wire n3991;
    wire n3994;
    wire n3997;
    wire n4001;
    wire n4004;
    wire n4007;
    wire n4010;
    wire n4012;
    wire n4015;
    wire n4018;
    wire n4021;
    wire n4024;
    wire n4027;
    wire n4030;
    wire n4033;
    wire n4036;
    wire n4039;
    wire n4042;
    wire n4045;
    wire n4048;
    wire n4051;
    wire n4054;
    wire n4057;
    wire n4060;
    wire n4063;
    wire n4066;
    wire n4069;
    wire n4072;
    wire n4075;
    wire n4078;
    wire n4081;
    wire n4084;
    wire n4087;
    wire n4090;
    wire n4093;
    wire n4097;
    wire n4100;
    wire n4103;
    wire n4105;
    wire n4108;
    wire n4111;
    wire n4114;
    wire n4117;
    wire n4120;
    wire n4123;
    wire n4126;
    wire n4129;
    wire n4132;
    wire n4135;
    wire n4138;
    wire n4141;
    wire n4144;
    wire n4147;
    wire n4150;
    wire n4153;
    wire n4156;
    wire n4159;
    wire n4162;
    wire n4165;
    wire n4168;
    wire n4171;
    wire n4174;
    wire n4177;
    wire n4180;
    wire n4183;
    wire n4186;
    wire n4189;
    wire n4192;
    wire n4195;
    wire n4198;
    wire n4201;
    wire n4204;
    wire n4207;
    wire n4210;
    wire n4213;
    wire n4216;
    wire n4219;
    wire n4222;
    wire n4225;
    wire n4229;
    wire n4232;
    wire n4235;
    wire n4238;
    wire n4240;
    wire n4243;
    wire n4246;
    wire n4249;
    wire n4252;
    wire n4255;
    wire n4258;
    wire n4261;
    wire n4264;
    wire n4267;
    wire n4270;
    wire n4274;
    wire n4277;
    wire n4280;
    wire n4283;
    wire n4286;
    wire n4288;
    wire n4291;
    wire n4295;
    wire n4297;
    wire n4300;
    wire n4303;
    wire n4306;
    wire n4309;
    wire n4312;
    wire n4315;
    wire n4318;
    wire n4321;
    wire n4324;
    wire n4327;
    wire n4330;
    wire n4333;
    wire n4336;
    wire n4339;
    wire n4342;
    wire n4345;
    wire n4348;
    wire n4351;
    wire n4354;
    wire n4357;
    wire n4360;
    wire n4363;
    wire n4366;
    wire n4369;
    wire n4372;
    wire n4375;
    wire n4378;
    wire n4381;
    wire n4384;
    wire n4387;
    wire n4390;
    wire n4393;
    wire n4396;
    wire n4399;
    wire n4402;
    wire n4405;
    wire n4408;
    wire n4411;
    wire n4414;
    wire n4417;
    wire n4420;
    wire n4423;
    wire n4426;
    wire n4429;
    wire n4432;
    wire n4435;
    wire n4438;
    wire n4441;
    wire n4447;
    wire n4450;
    wire n4453;
    wire n4456;
    wire n4459;
    wire n4462;
    wire n4465;
    wire n4468;
    wire n4471;
    wire n4474;
    wire n4477;
    wire n4480;
    wire n4483;
    wire n4486;
    wire n4489;
    wire n4492;
    wire n4495;
    wire n4498;
    wire n4504;
    wire n4507;
    wire n4510;
    wire n4513;
    wire n4516;
    wire n4519;
    wire n4522;
    wire n4525;
    wire n4528;
    wire n4531;
    wire n4534;
    wire n4537;
    wire n4540;
    wire n4543;
    wire n4546;
    wire n4549;
    wire n4552;
    wire n4555;
    wire n4561;
    wire n4564;
    wire n4567;
    wire n4570;
    wire n4573;
    wire n4576;
    wire n4579;
    wire n4582;
    wire n4585;
    wire n4588;
    wire n4591;
    wire n4594;
    wire n4597;
    wire n4600;
    wire n4603;
    wire n4606;
    wire n4609;
    wire n4612;
    wire n4615;
    wire n4621;
    wire n4624;
    wire n4627;
    wire n4630;
    wire n4633;
    wire n4636;
    wire n4639;
    wire n4642;
    wire n4645;
    wire n4648;
    wire n4651;
    wire n4654;
    wire n4657;
    wire n4660;
    wire n4663;
    wire n4666;
    wire n4669;
    wire n4672;
    wire n4678;
    wire n4681;
    wire n4684;
    wire n4687;
    wire n4690;
    wire n4693;
    wire n4696;
    wire n4699;
    wire n4702;
    wire n4705;
    wire n4708;
    wire n4711;
    wire n4714;
    wire n4717;
    wire n4720;
    wire n4723;
    wire n4729;
    wire n4732;
    wire n4735;
    wire n4738;
    wire n4741;
    wire n4744;
    wire n4747;
    wire n4750;
    wire n4753;
    wire n4756;
    wire n4759;
    wire n4762;
    wire n4765;
    wire n4768;
    wire n4771;
    wire n4774;
    wire n4777;
    wire n4783;
    wire n4786;
    wire n4789;
    wire n4792;
    wire n4795;
    wire n4798;
    wire n4801;
    wire n4804;
    wire n4807;
    wire n4810;
    wire n4813;
    wire n4816;
    wire n4819;
    wire n4822;
    wire n4825;
    wire n4828;
    wire n4831;
    wire n4837;
    wire n4840;
    wire n4843;
    wire n4846;
    wire n4849;
    wire n4852;
    wire n4855;
    wire n4858;
    wire n4861;
    wire n4864;
    wire n4867;
    wire n4870;
    wire n4873;
    wire n4876;
    wire n4879;
    wire n4882;
    wire n4885;
    wire n4891;
    wire n4894;
    wire n4897;
    wire n4900;
    wire n4903;
    wire n4906;
    wire n4909;
    wire n4912;
    wire n4915;
    wire n4918;
    wire n4921;
    wire n4924;
    wire n4927;
    wire n4930;
    wire n4933;
    wire n4936;
    wire n4939;
    wire n4942;
    wire n4948;
    wire n4951;
    wire n4954;
    wire n4957;
    wire n4960;
    wire n4963;
    wire n4966;
    wire n4969;
    wire n4972;
    wire n4975;
    wire n4978;
    wire n4981;
    wire n4984;
    wire n4987;
    wire n4990;
    wire n4993;
    wire n4999;
    wire n5002;
    wire n5005;
    wire n5008;
    wire n5011;
    wire n5014;
    wire n5017;
    wire n5020;
    wire n5023;
    wire n5026;
    wire n5029;
    wire n5032;
    wire n5035;
    wire n5038;
    wire n5041;
    wire n5044;
    wire n5047;
    wire n5050;
    wire n5056;
    wire n5059;
    wire n5062;
    wire n5065;
    wire n5068;
    wire n5071;
    wire n5074;
    wire n5077;
    wire n5080;
    wire n5083;
    wire n5086;
    wire n5089;
    wire n5092;
    wire n5095;
    wire n5098;
    wire n5101;
    wire n5104;
    wire n5110;
    wire n5113;
    wire n5116;
    wire n5119;
    wire n5122;
    wire n5125;
    wire n5128;
    wire n5131;
    wire n5134;
    wire n5137;
    wire n5140;
    wire n5143;
    wire n5146;
    wire n5149;
    wire n5152;
    wire n5155;
    wire n5158;
    wire n5164;
    wire n5167;
    wire n5170;
    wire n5173;
    wire n5176;
    wire n5179;
    wire n5182;
    wire n5185;
    wire n5188;
    wire n5191;
    wire n5194;
    wire n5197;
    wire n5200;
    wire n5203;
    wire n5206;
    wire n5209;
    wire n5212;
    wire n5215;
    wire n5221;
    wire n5224;
    wire n5227;
    wire n5230;
    wire n5233;
    wire n5236;
    wire n5239;
    wire n5242;
    wire n5245;
    wire n5248;
    wire n5251;
    wire n5254;
    wire n5257;
    wire n5260;
    wire n5263;
    wire n5266;
    wire n5272;
    wire n5275;
    wire n5278;
    wire n5281;
    wire n5284;
    wire n5287;
    wire n5290;
    wire n5293;
    wire n5296;
    wire n5299;
    wire n5302;
    wire n5305;
    wire n5308;
    wire n5311;
    wire n5314;
    wire n5317;
    wire n5323;
    wire n5326;
    wire n5329;
    wire n5332;
    wire n5335;
    wire n5338;
    wire n5341;
    wire n5347;
    wire n5350;
    wire n5353;
    wire n5359;
    wire n5362;
    wire n5365;
    wire n5371;
    wire n5374;
    wire n5377;
    wire n5380;
    wire n5383;
    wire n5389;
    wire n5395;
    jand g000(.dinb(G29gat), .dina(G75gat), .dout(n89));
    jand g001(.dinb(n4318), .dina(n89), .dout(n93));
    jand g002(.dinb(G29gat), .dina(G36gat), .dout(n97));
    jand g003(.dinb(n4255), .dina(n97), .dout(n101));
    jand g004(.dinb(n4318), .dina(n97), .dout(n105));
    jand g005(.dinb(G85gat), .dina(G86gat), .dout(n109));
    jand g006(.dinb(G1gat), .dina(G8gat), .dout(n113));
    jand g007(.dinb(G13gat), .dina(G17gat), .dout(n117));
    jand g008(.dinb(n113), .dina(n117), .dout(n121));
    jnot g009(.din(n117), .dout(n124));
    jnot g010(.din(G1gat), .dout(n127));
    jnot g011(.din(G26gat), .dout(n130));
    jor g012(.dinb(n127), .dina(n130), .dout(n134));
    jor g013(.dinb(n124), .dina(n134), .dout(n138));
    jor g014(.dinb(n2029), .dina(n138), .dout(n142));
    jnot g015(.din(G80gat), .dout(n145));
    jand g016(.dinb(G59gat), .dina(G75gat), .dout(n149));
    jnot g017(.din(n149), .dout(n152));
    jor g018(.dinb(n2021), .dina(n152), .dout(n156));
    jnot g019(.din(G36gat), .dout(n159));
    jnot g020(.din(G59gat), .dout(n162));
    jor g021(.dinb(n159), .dina(n162), .dout(n166));
    jor g022(.dinb(n2021), .dina(n166), .dout(n170));
    jnot g023(.din(G42gat), .dout(n173));
    jor g024(.dinb(n2024), .dina(n166), .dout(n177));
    jor g025(.dinb(G87gat), .dina(G88gat), .dout(n181));
    jand g026(.dinb(n2027), .dina(n181), .dout(n185));
    jnot g027(.din(n105), .dout(n188));
    jor g028(.dinb(n188), .dina(n138), .dout(n192));
    jand g029(.dinb(G1gat), .dina(G26gat), .dout(n196));
    jand g030(.dinb(n4297), .dina(n196), .dout(n200));
    jand g031(.dinb(G13gat), .dina(G55gat), .dout(n204));
    jand g032(.dinb(n113), .dina(n204), .dout(n208));
    jand g033(.dinb(G29gat), .dina(G68gat), .dout(n212));
    jand g034(.dinb(n208), .dina(n2033), .dout(n216));
    jand g035(.dinb(G59gat), .dina(G68gat), .dout(n220));
    jand g036(.dinb(n2036), .dina(n220), .dout(n224));
    jand g037(.dinb(n208), .dina(n224), .dout(n228));
    jand g038(.dinb(n2039), .dina(n181), .dout(n232));
    jxor g039(.dinb(G91gat), .dina(G96gat), .dout(n236));
    jxor g040(.dinb(n2060), .dina(n236), .dout(n240));
    jxor g041(.dinb(G121gat), .dina(G126gat), .dout(n244));
    jxor g042(.dinb(n240), .dina(n2048), .dout(n248));
    jxor g043(.dinb(G111gat), .dina(G116gat), .dout(n252));
    jxor g044(.dinb(n2045), .dina(n252), .dout(n256));
    jxor g045(.dinb(G101gat), .dina(G106gat), .dout(n260));
    jxor g046(.dinb(n256), .dina(n2042), .dout(n264));
    jxor g047(.dinb(n248), .dina(n264), .dout(n268));
    jxor g048(.dinb(G159gat), .dina(G165gat), .dout(n272));
    jxor g049(.dinb(n2060), .dina(n272), .dout(n276));
    jxor g050(.dinb(G195gat), .dina(G201gat), .dout(n280));
    jxor g051(.dinb(n276), .dina(n2057), .dout(n284));
    jxor g052(.dinb(G183gat), .dina(G189gat), .dout(n288));
    jxor g053(.dinb(n2054), .dina(n288), .dout(n292));
    jxor g054(.dinb(G171gat), .dina(G177gat), .dout(n296));
    jxor g055(.dinb(n292), .dina(n2051), .dout(n300));
    jxor g056(.dinb(n284), .dina(n300), .dout(n304));
    jnot g057(.din(G261gat), .dout(n307));
    jand g058(.dinb(n4315), .dina(n149), .dout(n311));
    jnot g059(.din(n311), .dout(n314));
    jand g060(.dinb(G17gat), .dina(G51gat), .dout(n318));
    jand g061(.dinb(n113), .dina(n318), .dout(n322));
    jand g062(.dinb(n314), .dina(n4295), .dout(n326));
    jand g063(.dinb(G59gat), .dina(G156gat), .dout(n330));
    jxor g064(.dinb(G17gat), .dina(G42gat), .dout(n334));
    jand g065(.dinb(n330), .dina(n334), .dout(n338));
    jand g066(.dinb(n200), .dina(n338), .dout(n342));
    jor g067(.dinb(n326), .dina(n4286), .dout(n346));
    jand g068(.dinb(n3841), .dina(n346), .dout(n350));
    jnot g069(.din(G156gat), .dout(n353));
    jor g070(.dinb(n162), .dina(n353), .dout(n357));
    jand g071(.dinb(n200), .dina(n357), .dout(n361));
    jand g072(.dinb(n4243), .dina(n361), .dout(n365));
    jor g073(.dinb(n3988), .dina(n365), .dout(n369));
    jand g074(.dinb(n4117), .dina(n369), .dout(n373));
    jand g075(.dinb(n4252), .dina(n89), .dout(n377));
    jand g076(.dinb(n200), .dina(n377), .dout(n381));
    jnot g077(.din(G268gat), .dout(n384));
    jand g078(.dinb(n4267), .dina(n384), .dout(n388));
    jand g079(.dinb(n381), .dina(n3986), .dout(n392));
    jor g080(.dinb(n373), .dina(n3967), .dout(n396));
    jor g081(.dinb(n3838), .dina(n396), .dout(n400));
    jxor g082(.dinb(n2101), .dina(n400), .dout(n404));
    jnot g083(.din(n404), .dout(n407));
    jor g084(.dinb(n3779), .dina(n407), .dout(n411));
    jor g085(.dinb(n3808), .dina(n404), .dout(n415));
    jand g086(.dinb(n3299), .dina(n415), .dout(n419));
    jand g087(.dinb(n411), .dina(n419), .dout(n423));
    jand g088(.dinb(n3214), .dina(n404), .dout(n427));
    jand g089(.dinb(G201gat), .dina(G237gat), .dout(n431));
    jor g090(.dinb(n3212), .dina(n431), .dout(n435));
    jand g091(.dinb(n400), .dina(n2099), .dout(n439));
    jand g092(.dinb(G42gat), .dina(G72gat), .dout(n443));
    jand g093(.dinb(n3188), .dina(n443), .dout(n447));
    jand g094(.dinb(n3190), .dina(n447), .dout(n451));
    jand g095(.dinb(n3193), .dina(n451), .dout(n455));
    jand g096(.dinb(n3880), .dina(n455), .dout(n459));
    jand g097(.dinb(G121gat), .dina(G210gat), .dout(n463));
    jand g098(.dinb(G255gat), .dina(G267gat), .dout(n467));
    jor g099(.dinb(n463), .dina(n467), .dout(n471));
    jor g100(.dinb(n459), .dina(n2081), .dout(n475));
    jor g101(.dinb(n439), .dina(n2072), .dout(n479));
    jor g102(.dinb(n427), .dina(n479), .dout(n483));
    jor g103(.dinb(n423), .dina(n2063), .dout(n487));
    jand g104(.dinb(n3997), .dina(n369), .dout(n491));
    jand g105(.dinb(n3946), .dina(n346), .dout(n495));
    jor g106(.dinb(n3961), .dina(n495), .dout(n499));
    jor g107(.dinb(n3944), .dina(n499), .dout(n503));
    jxor g108(.dinb(n2215), .dina(n503), .dout(n507));
    jnot g109(.din(n507), .dout(n510));
    jand g110(.dinb(n3856), .dina(n400), .dout(n514));
    jnot g111(.din(n514), .dout(n517));
    jnot g112(.din(G201gat), .dout(n520));
    jnot g113(.din(n350), .dout(n523));
    jnot g114(.din(G153gat), .dout(n526));
    jnot g115(.din(G17gat), .dout(n529));
    jnot g116(.din(G51gat), .dout(n532));
    jor g117(.dinb(n3752), .dina(n134), .dout(n536));
    jor g118(.dinb(n536), .dina(n4288), .dout(n540));
    jor g119(.dinb(n3749), .dina(n540), .dout(n544));
    jand g120(.dinb(n4300), .dina(n544), .dout(n548));
    jor g121(.dinb(n3740), .dina(n548), .dout(n552));
    jnot g122(.din(n392), .dout(n555));
    jand g123(.dinb(n552), .dina(n3725), .dout(n559));
    jand g124(.dinb(n3719), .dina(n559), .dout(n563));
    jand g125(.dinb(n3716), .dina(n563), .dout(n567));
    jor g126(.dinb(n3779), .dina(n567), .dout(n571));
    jand g127(.dinb(n3692), .dina(n571), .dout(n575));
    jand g128(.dinb(n3640), .dina(n369), .dout(n579));
    jand g129(.dinb(n3625), .dina(n346), .dout(n583));
    jor g130(.dinb(n3979), .dina(n583), .dout(n587));
    jor g131(.dinb(n3623), .dina(n587), .dout(n591));
    jor g132(.dinb(n3655), .dina(n591), .dout(n595));
    jand g133(.dinb(n4270), .dina(n369), .dout(n599));
    jand g134(.dinb(n3571), .dina(n346), .dout(n603));
    jor g135(.dinb(n3973), .dina(n603), .dout(n607));
    jor g136(.dinb(n3569), .dina(n607), .dout(n611));
    jor g137(.dinb(n3586), .dina(n611), .dout(n615));
    jand g138(.dinb(n595), .dina(n615), .dout(n619));
    jnot g139(.din(n619), .dout(n622));
    jor g140(.dinb(n575), .dina(n3557), .dout(n626));
    jand g141(.dinb(n3532), .dina(n591), .dout(n630));
    jand g142(.dinb(n3484), .dina(n611), .dout(n634));
    jand g143(.dinb(n595), .dina(n634), .dout(n638));
    jor g144(.dinb(n3449), .dina(n638), .dout(n642));
    jnot g145(.din(n642), .dout(n645));
    jand g146(.dinb(n626), .dina(n3443), .dout(n649));
    jor g147(.dinb(n2201), .dina(n649), .dout(n653));
    jor g148(.dinb(n3892), .dina(n400), .dout(n657));
    jand g149(.dinb(n3781), .dina(n657), .dout(n661));
    jor g150(.dinb(n3835), .dina(n661), .dout(n665));
    jand g151(.dinb(n665), .dina(n3559), .dout(n669));
    jor g152(.dinb(n669), .dina(n3445), .dout(n673));
    jor g153(.dinb(n2203), .dina(n673), .dout(n677));
    jand g154(.dinb(n2179), .dina(n677), .dout(n681));
    jand g155(.dinb(n653), .dina(n681), .dout(n685));
    jand g156(.dinb(n3214), .dina(n507), .dout(n689));
    jand g157(.dinb(G183gat), .dina(G237gat), .dout(n693));
    jor g158(.dinb(n3212), .dina(n693), .dout(n697));
    jand g159(.dinb(n503), .dina(n2177), .dout(n701));
    jand g160(.dinb(n4036), .dina(n455), .dout(n705));
    jand g161(.dinb(G106gat), .dina(G210gat), .dout(n709));
    jor g162(.dinb(n705), .dina(n2159), .dout(n713));
    jor g163(.dinb(n701), .dina(n2147), .dout(n717));
    jor g164(.dinb(n689), .dina(n717), .dout(n721));
    jor g165(.dinb(n685), .dina(n2138), .dout(n725));
    jxor g166(.dinb(n3508), .dina(n591), .dout(n729));
    jnot g167(.din(n729), .dout(n732));
    jand g168(.dinb(n665), .dina(n3562), .dout(n736));
    jor g169(.dinb(n3451), .dina(n736), .dout(n740));
    jnot g170(.din(n740), .dout(n743));
    jor g171(.dinb(n2300), .dina(n743), .dout(n747));
    jor g172(.dinb(n2302), .dina(n740), .dout(n751));
    jand g173(.dinb(n2524), .dina(n751), .dout(n755));
    jand g174(.dinb(n747), .dina(n755), .dout(n759));
    jand g175(.dinb(n2509), .dina(n729), .dout(n763));
    jand g176(.dinb(G189gat), .dina(G237gat), .dout(n767));
    jor g177(.dinb(n3212), .dina(n767), .dout(n771));
    jand g178(.dinb(n591), .dina(n2288), .dout(n775));
    jand g179(.dinb(n3679), .dina(n455), .dout(n779));
    jand g180(.dinb(G111gat), .dina(G210gat), .dout(n783));
    jand g181(.dinb(G255gat), .dina(G259gat), .dout(n787));
    jor g182(.dinb(n783), .dina(n787), .dout(n791));
    jor g183(.dinb(n779), .dina(n2270), .dout(n795));
    jor g184(.dinb(n775), .dina(n2261), .dout(n799));
    jor g185(.dinb(n763), .dina(n799), .dout(n803));
    jor g186(.dinb(n759), .dina(n2252), .dout(n807));
    jxor g187(.dinb(n3460), .dina(n611), .dout(n811));
    jnot g188(.din(n811), .dout(n814));
    jor g189(.dinb(n575), .dina(n2363), .dout(n818));
    jor g190(.dinb(n665), .dina(n2365), .dout(n822));
    jand g191(.dinb(n3265), .dina(n822), .dout(n826));
    jand g192(.dinb(n818), .dina(n826), .dout(n830));
    jand g193(.dinb(n2506), .dina(n811), .dout(n834));
    jand g194(.dinb(G195gat), .dina(G237gat), .dout(n838));
    jor g195(.dinb(n3212), .dina(n838), .dout(n842));
    jand g196(.dinb(n611), .dina(n2357), .dout(n846));
    jand g197(.dinb(n3610), .dina(n455), .dout(n850));
    jand g198(.dinb(G116gat), .dina(G210gat), .dout(n854));
    jand g199(.dinb(G255gat), .dina(G260gat), .dout(n858));
    jor g200(.dinb(n854), .dina(n858), .dout(n862));
    jor g201(.dinb(n850), .dina(n2339), .dout(n866));
    jor g202(.dinb(n846), .dina(n2330), .dout(n870));
    jor g203(.dinb(n834), .dina(n870), .dout(n874));
    jor g204(.dinb(n830), .dina(n2321), .dout(n878));
    jand g205(.dinb(n2878), .dina(n346), .dout(n882));
    jand g206(.dinb(n4258), .dina(n361), .dout(n886));
    jand g207(.dinb(n4010), .dina(n886), .dout(n890));
    jand g208(.dinb(G8gat), .dina(G138gat), .dout(n894));
    jand g209(.dinb(n4240), .dina(n384), .dout(n898));
    jand g210(.dinb(n381), .dina(n4238), .dout(n902));
    jor g211(.dinb(n2696), .dina(n902), .dout(n906));
    jor g212(.dinb(n890), .dina(n906), .dout(n910));
    jor g213(.dinb(n882), .dina(n910), .dout(n914));
    jand g214(.dinb(n2428), .dina(n914), .dout(n918));
    jor g215(.dinb(n2719), .dina(n914), .dout(n922));
    jand g216(.dinb(n4012), .dina(n503), .dout(n926));
    jor g217(.dinb(n4048), .dina(n503), .dout(n930));
    jand g218(.dinb(n3916), .dina(n673), .dout(n934));
    jor g219(.dinb(n3928), .dina(n934), .dout(n938));
    jnot g220(.din(G165gat), .dout(n941));
    jand g221(.dinb(n3172), .dina(n346), .dout(n945));
    jand g222(.dinb(n3653), .dina(n886), .dout(n949));
    jand g223(.dinb(G51gat), .dina(G138gat), .dout(n953));
    jor g224(.dinb(n902), .dina(n3068), .dout(n957));
    jor g225(.dinb(n949), .dina(n957), .dout(n961));
    jor g226(.dinb(n945), .dina(n961), .dout(n965));
    jnot g227(.din(n965), .dout(n968));
    jand g228(.dinb(n2828), .dina(n968), .dout(n972));
    jnot g229(.din(n972), .dout(n975));
    jand g230(.dinb(n4321), .dina(n346), .dout(n979));
    jand g231(.dinb(n4283), .dina(n886), .dout(n983));
    jand g232(.dinb(G17gat), .dina(G138gat), .dout(n987));
    jor g233(.dinb(n902), .dina(n4235), .dout(n991));
    jor g234(.dinb(n983), .dina(n991), .dout(n995));
    jor g235(.dinb(n979), .dina(n995), .dout(n999));
    jor g236(.dinb(n3013), .dina(n999), .dout(n1003));
    jand g237(.dinb(n4132), .dina(n346), .dout(n1007));
    jand g238(.dinb(n4105), .dina(n886), .dout(n1011));
    jand g239(.dinb(G138gat), .dina(G152gat), .dout(n1015));
    jor g240(.dinb(n902), .dina(n4103), .dout(n1019));
    jor g241(.dinb(n1011), .dina(n1019), .dout(n1023));
    jor g242(.dinb(n1007), .dina(n1023), .dout(n1027));
    jor g243(.dinb(n3394), .dina(n1027), .dout(n1031));
    jand g244(.dinb(n1003), .dina(n1031), .dout(n1035));
    jand g245(.dinb(n975), .dina(n2989), .dout(n1039));
    jand g246(.dinb(n938), .dina(n2797), .dout(n1043));
    jand g247(.dinb(n3091), .dina(n965), .dout(n1047));
    jand g248(.dinb(n4357), .dina(n999), .dout(n1051));
    jand g249(.dinb(n4168), .dina(n1027), .dout(n1055));
    jand g250(.dinb(n1003), .dina(n1055), .dout(n1059));
    jor g251(.dinb(n3011), .dina(n1059), .dout(n1063));
    jand g252(.dinb(n975), .dina(n1063), .dout(n1067));
    jor g253(.dinb(n2783), .dina(n1067), .dout(n1071));
    jor g254(.dinb(n1043), .dina(n2764), .dout(n1075));
    jand g255(.dinb(n2426), .dina(n1075), .dout(n1079));
    jor g256(.dinb(n2399), .dina(n1079), .dout(n1083));
    jnot g257(.din(n926), .dout(n1086));
    jnot g258(.din(n930), .dout(n1089));
    jor g259(.dinb(n3440), .dina(n649), .dout(n1093));
    jand g260(.dinb(n3428), .dina(n1093), .dout(n1097));
    jxor g261(.dinb(n4147), .dina(n1027), .dout(n1101));
    jnot g262(.din(n1101), .dout(n1104));
    jor g263(.dinb(n1097), .dina(n2549), .dout(n1108));
    jor g264(.dinb(n938), .dina(n2551), .dout(n1112));
    jand g265(.dinb(n2512), .dina(n1112), .dout(n1116));
    jand g266(.dinb(n1108), .dina(n1116), .dout(n1120));
    jand g267(.dinb(n3239), .dina(n1101), .dout(n1124));
    jand g268(.dinb(G177gat), .dina(G237gat), .dout(n1128));
    jor g269(.dinb(n3212), .dina(n1128), .dout(n1132));
    jand g270(.dinb(n1027), .dina(n2504), .dout(n1136));
    jand g271(.dinb(n4189), .dina(n455), .dout(n1140));
    jand g272(.dinb(G101gat), .dina(G210gat), .dout(n1144));
    jor g273(.dinb(n1140), .dina(n2489), .dout(n1148));
    jor g274(.dinb(n1136), .dina(n2477), .dout(n1152));
    jor g275(.dinb(n1124), .dina(n1152), .dout(n1156));
    jor g276(.dinb(n1120), .dina(n2471), .dout(n1160));
    jnot g277(.din(n1039), .dout(n1163));
    jor g278(.dinb(n1097), .dina(n2795), .dout(n1167));
    jnot g279(.din(n1071), .dout(n1170));
    jand g280(.dinb(n1167), .dina(n2762), .dout(n1174));
    jxor g281(.dinb(n2698), .dina(n914), .dout(n1178));
    jnot g282(.din(n1178), .dout(n1181));
    jor g283(.dinb(n1174), .dina(n2660), .dout(n1185));
    jor g284(.dinb(n1075), .dina(n2662), .dout(n1189));
    jand g285(.dinb(n3241), .dina(n1189), .dout(n1193));
    jand g286(.dinb(n1185), .dina(n1193), .dout(n1197));
    jand g287(.dinb(n3239), .dina(n1178), .dout(n1201));
    jand g288(.dinb(G159gat), .dina(G237gat), .dout(n1205));
    jor g289(.dinb(n3212), .dina(n1205), .dout(n1209));
    jand g290(.dinb(n914), .dina(n2633), .dout(n1213));
    jand g291(.dinb(n2740), .dina(n455), .dout(n1217));
    jand g292(.dinb(G210gat), .dina(G268gat), .dout(n1221));
    jor g293(.dinb(n1217), .dina(n2618), .dout(n1225));
    jor g294(.dinb(n1213), .dina(n2606), .dout(n1229));
    jor g295(.dinb(n1201), .dina(n1229), .dout(n1233));
    jor g296(.dinb(n1197), .dina(n2600), .dout(G878gat));
    jxor g297(.dinb(n3070), .dina(n965), .dout(n1241));
    jnot g298(.din(n1241), .dout(n1244));
    jnot g299(.din(n1063), .dout(n1247));
    jnot g300(.din(n1035), .dout(n1250));
    jor g301(.dinb(n1097), .dina(n2969), .dout(n1254));
    jand g302(.dinb(n2951), .dina(n1254), .dout(n1258));
    jor g303(.dinb(n2933), .dina(n1258), .dout(n1262));
    jand g304(.dinb(n938), .dina(n2971), .dout(n1266));
    jor g305(.dinb(n2992), .dina(n1266), .dout(n1270));
    jor g306(.dinb(n3034), .dina(n1270), .dout(n1274));
    jand g307(.dinb(n3241), .dina(n1274), .dout(n1278));
    jand g308(.dinb(n1262), .dina(n1278), .dout(n1282));
    jand g309(.dinb(n3239), .dina(n1241), .dout(n1286));
    jand g310(.dinb(G165gat), .dina(G237gat), .dout(n1290));
    jor g311(.dinb(n3212), .dina(n1290), .dout(n1294));
    jand g312(.dinb(n965), .dina(n2906), .dout(n1298));
    jand g313(.dinb(n3112), .dina(n455), .dout(n1302));
    jand g314(.dinb(G91gat), .dina(G210gat), .dout(n1306));
    jor g315(.dinb(n1302), .dina(n2876), .dout(n1310));
    jor g316(.dinb(n1298), .dina(n2864), .dout(n1314));
    jor g317(.dinb(n1286), .dina(n1314), .dout(n1318));
    jor g318(.dinb(n1282), .dina(n2858), .dout(G879gat));
    jxor g319(.dinb(n4336), .dina(n999), .dout(n1326));
    jnot g320(.din(n1326), .dout(n1329));
    jnot g321(.din(n1055), .dout(n1332));
    jnot g322(.din(n1031), .dout(n1335));
    jor g323(.dinb(n1097), .dina(n3371), .dout(n1339));
    jand g324(.dinb(n3350), .dina(n1339), .dout(n1343));
    jor g325(.dinb(n3326), .dina(n1343), .dout(n1347));
    jand g326(.dinb(n938), .dina(n3373), .dout(n1351));
    jor g327(.dinb(n4072), .dina(n1351), .dout(n1355));
    jor g328(.dinb(n4201), .dina(n1355), .dout(n1359));
    jand g329(.dinb(n3241), .dina(n1359), .dout(n1363));
    jand g330(.dinb(n1347), .dina(n1363), .dout(n1367));
    jand g331(.dinb(n3239), .dina(n1326), .dout(n1371));
    jand g332(.dinb(G171gat), .dina(G237gat), .dout(n1375));
    jor g333(.dinb(n3212), .dina(n1375), .dout(n1379));
    jand g334(.dinb(n999), .dina(n3209), .dout(n1383));
    jand g335(.dinb(n4378), .dina(n455), .dout(n1387));
    jand g336(.dinb(G96gat), .dina(G210gat), .dout(n1391));
    jor g337(.dinb(n1387), .dina(n3170), .dout(n1395));
    jor g338(.dinb(n1383), .dina(n3158), .dout(n1399));
    jor g339(.dinb(n1371), .dina(n1399), .dout(n1403));
    jor g340(.dinb(n1367), .dina(n3152), .dout(G880gat));
    jdff dff_A_bCGK6ity0_0(.din(n5395), .dout(G874gat));
    jdff dff_A_4uviTJyN4_2(.din(n1160), .dout(n5395));
    jdff dff_A_sr7IBH1k9_0(.din(n5389), .dout(G866gat));
    jdff dff_A_k24t8EOj8_2(.din(n1083), .dout(n5389));
    jdff dff_A_NUrM0tWc5_0(.din(n5383), .dout(G865gat));
    jdff dff_A_uqNWdzWx9_0(.din(n5380), .dout(n5383));
    jdff dff_A_z1oCuJhh8_0(.din(n5377), .dout(n5380));
    jdff dff_A_cUuhVVoP3_0(.din(n5374), .dout(n5377));
    jdff dff_A_sworGvl53_0(.din(n5371), .dout(n5374));
    jdff dff_A_yKfR0GGH1_2(.din(n878), .dout(n5371));
    jdff dff_A_j82oyDVy1_0(.din(n5365), .dout(G864gat));
    jdff dff_A_pTdiBhOH3_0(.din(n5362), .dout(n5365));
    jdff dff_A_wq0l5bdW9_0(.din(n5359), .dout(n5362));
    jdff dff_A_VWu5r75i1_2(.din(n807), .dout(n5359));
    jdff dff_A_nO3QnoHq0_0(.din(n5353), .dout(G863gat));
    jdff dff_A_utUMXrRq9_0(.din(n5350), .dout(n5353));
    jdff dff_A_y1E9JOjN1_0(.din(n5347), .dout(n5350));
    jdff dff_A_mgcnRDmm4_2(.din(n725), .dout(n5347));
    jdff dff_A_EGj3SVRD2_0(.din(n5341), .dout(G850gat));
    jdff dff_A_SCKs2Omb9_0(.din(n5338), .dout(n5341));
    jdff dff_A_ht8ABj3t4_0(.din(n5335), .dout(n5338));
    jdff dff_A_YoqysCiO4_0(.din(n5332), .dout(n5335));
    jdff dff_A_J21VZuxz4_0(.din(n5329), .dout(n5332));
    jdff dff_A_aYieiXnk6_0(.din(n5326), .dout(n5329));
    jdff dff_A_gX40HpxM5_0(.din(n5323), .dout(n5326));
    jdff dff_A_7W4PhO7b3_2(.din(n487), .dout(n5323));
    jdff dff_A_ROsCN0oV9_0(.din(n5317), .dout(G768gat));
    jdff dff_A_CUal9O1N1_0(.din(n5314), .dout(n5317));
    jdff dff_A_UEJG2x9F1_0(.din(n5311), .dout(n5314));
    jdff dff_A_SC76EtqL9_0(.din(n5308), .dout(n5311));
    jdff dff_A_qUN49Yui5_0(.din(n5305), .dout(n5308));
    jdff dff_A_Hzkem6hU8_0(.din(n5302), .dout(n5305));
    jdff dff_A_2SuZKbSr9_0(.din(n5299), .dout(n5302));
    jdff dff_A_1QrvILdF1_0(.din(n5296), .dout(n5299));
    jdff dff_A_4MpTUQrL9_0(.din(n5293), .dout(n5296));
    jdff dff_A_L6iLODd12_0(.din(n5290), .dout(n5293));
    jdff dff_A_ZzdwRnFU3_0(.din(n5287), .dout(n5290));
    jdff dff_A_6Pw5vc0f1_0(.din(n5284), .dout(n5287));
    jdff dff_A_DtIC18th4_0(.din(n5281), .dout(n5284));
    jdff dff_A_0eEcsSck5_0(.din(n5278), .dout(n5281));
    jdff dff_A_pWu2FU9w1_0(.din(n5275), .dout(n5278));
    jdff dff_A_2Sfk8hZq5_0(.din(n5272), .dout(n5275));
    jdff dff_A_4vD5BJ2U0_2(.din(n304), .dout(n5272));
    jdff dff_A_0IlwTYZ81_0(.din(n5266), .dout(G767gat));
    jdff dff_A_As6zZmd30_0(.din(n5263), .dout(n5266));
    jdff dff_A_sJmRVQDw9_0(.din(n5260), .dout(n5263));
    jdff dff_A_CugvgRr46_0(.din(n5257), .dout(n5260));
    jdff dff_A_20bCMobo8_0(.din(n5254), .dout(n5257));
    jdff dff_A_hV6sMuhr8_0(.din(n5251), .dout(n5254));
    jdff dff_A_aMpIvDcO3_0(.din(n5248), .dout(n5251));
    jdff dff_A_QVyTf5I20_0(.din(n5245), .dout(n5248));
    jdff dff_A_viuvkxgk6_0(.din(n5242), .dout(n5245));
    jdff dff_A_IlpauXBo3_0(.din(n5239), .dout(n5242));
    jdff dff_A_fbfY82HE3_0(.din(n5236), .dout(n5239));
    jdff dff_A_QflP8YtV6_0(.din(n5233), .dout(n5236));
    jdff dff_A_JPLBFfI53_0(.din(n5230), .dout(n5233));
    jdff dff_A_3G9WnZxV1_0(.din(n5227), .dout(n5230));
    jdff dff_A_Im3bDWIN7_0(.din(n5224), .dout(n5227));
    jdff dff_A_uaor30g26_0(.din(n5221), .dout(n5224));
    jdff dff_A_xsrmNVkq7_2(.din(n268), .dout(n5221));
    jdff dff_A_svC8UNFs8_0(.din(n5215), .dout(G450gat));
    jdff dff_A_32HHgdDc0_0(.din(n5212), .dout(n5215));
    jdff dff_A_nNZP1V5O0_0(.din(n5209), .dout(n5212));
    jdff dff_A_PHgt0RCM2_0(.din(n5206), .dout(n5209));
    jdff dff_A_f5aOjsHf0_0(.din(n5203), .dout(n5206));
    jdff dff_A_08gBmKcK0_0(.din(n5200), .dout(n5203));
    jdff dff_A_oq6czHbW5_0(.din(n5197), .dout(n5200));
    jdff dff_A_nlOkYiMg2_0(.din(n5194), .dout(n5197));
    jdff dff_A_kEVaACIG0_0(.din(n5191), .dout(n5194));
    jdff dff_A_ZOeJBvtb0_0(.din(n5188), .dout(n5191));
    jdff dff_A_1b1w5zwa7_0(.din(n5185), .dout(n5188));
    jdff dff_A_0O1rlOkM9_0(.din(n5182), .dout(n5185));
    jdff dff_A_5HHzlktf9_0(.din(n5179), .dout(n5182));
    jdff dff_A_IsILClwD4_0(.din(n5176), .dout(n5179));
    jdff dff_A_TFxh5nxS0_0(.din(n5173), .dout(n5176));
    jdff dff_A_00R8rm1m6_0(.din(n5170), .dout(n5173));
    jdff dff_A_wp5znw2A7_0(.din(n5167), .dout(n5170));
    jdff dff_A_gQCgLpuQ3_0(.din(n5164), .dout(n5167));
    jdff dff_A_CrUGfiSX7_2(.din(n232), .dout(n5164));
    jdff dff_A_eRsuRZUc0_0(.din(n5158), .dout(G449gat));
    jdff dff_A_2NM1ELsb7_0(.din(n5155), .dout(n5158));
    jdff dff_A_niKJqv7r5_0(.din(n5152), .dout(n5155));
    jdff dff_A_uVEAPLAS1_0(.din(n5149), .dout(n5152));
    jdff dff_A_UtEUmA5r4_0(.din(n5146), .dout(n5149));
    jdff dff_A_5zFJQRLR1_0(.din(n5143), .dout(n5146));
    jdff dff_A_x9c69HAT5_0(.din(n5140), .dout(n5143));
    jdff dff_A_EfRRtaOF5_0(.din(n5137), .dout(n5140));
    jdff dff_A_JeZJ3xhm8_0(.din(n5134), .dout(n5137));
    jdff dff_A_dt74t9FM2_0(.din(n5131), .dout(n5134));
    jdff dff_A_fEYCxMoo8_0(.din(n5128), .dout(n5131));
    jdff dff_A_864MDl3i8_0(.din(n5125), .dout(n5128));
    jdff dff_A_OjXFrgtr1_0(.din(n5122), .dout(n5125));
    jdff dff_A_1kUW6dBg2_0(.din(n5119), .dout(n5122));
    jdff dff_A_iySXuQF41_0(.din(n5116), .dout(n5119));
    jdff dff_A_XPMuzRkf4_0(.din(n5113), .dout(n5116));
    jdff dff_A_mkY1nLu22_0(.din(n5110), .dout(n5113));
    jdff dff_A_csl3aRhX5_2(.din(n228), .dout(n5110));
    jdff dff_A_oaRMwzhY2_0(.din(n5104), .dout(G448gat));
    jdff dff_A_MkRBpyr40_0(.din(n5101), .dout(n5104));
    jdff dff_A_W3dLmgUe1_0(.din(n5098), .dout(n5101));
    jdff dff_A_XweZXmXJ1_0(.din(n5095), .dout(n5098));
    jdff dff_A_rck1oucl5_0(.din(n5092), .dout(n5095));
    jdff dff_A_xgwledVq0_0(.din(n5089), .dout(n5092));
    jdff dff_A_8LJkgOP54_0(.din(n5086), .dout(n5089));
    jdff dff_A_5SSV1iub4_0(.din(n5083), .dout(n5086));
    jdff dff_A_7gVl9CFj9_0(.din(n5080), .dout(n5083));
    jdff dff_A_UiTCakOA9_0(.din(n5077), .dout(n5080));
    jdff dff_A_aafD2M4u7_0(.din(n5074), .dout(n5077));
    jdff dff_A_w33NIjZJ6_0(.din(n5071), .dout(n5074));
    jdff dff_A_xtUb4BHg8_0(.din(n5068), .dout(n5071));
    jdff dff_A_iwvqaTI53_0(.din(n5065), .dout(n5068));
    jdff dff_A_yXgFXQGu6_0(.din(n5062), .dout(n5065));
    jdff dff_A_aHk1J1aU1_0(.din(n5059), .dout(n5062));
    jdff dff_A_IjVS0GVL5_0(.din(n5056), .dout(n5059));
    jdff dff_A_up1EhJML0_2(.din(n216), .dout(n5056));
    jdff dff_A_zmegFpcB2_0(.din(n5050), .dout(G447gat));
    jdff dff_A_HGE1uK6W9_0(.din(n5047), .dout(n5050));
    jdff dff_A_EKKJA5do1_0(.din(n5044), .dout(n5047));
    jdff dff_A_mvOK2W9h7_0(.din(n5041), .dout(n5044));
    jdff dff_A_60hFFASs2_0(.din(n5038), .dout(n5041));
    jdff dff_A_MSP2qFW88_0(.din(n5035), .dout(n5038));
    jdff dff_A_peBbtvtG6_0(.din(n5032), .dout(n5035));
    jdff dff_A_wciQpmws5_0(.din(n5029), .dout(n5032));
    jdff dff_A_Cr7eBnNh4_0(.din(n5026), .dout(n5029));
    jdff dff_A_A9ztUOAT4_0(.din(n5023), .dout(n5026));
    jdff dff_A_4RU2KqSQ4_0(.din(n5020), .dout(n5023));
    jdff dff_A_WgwIgCm09_0(.din(n5017), .dout(n5020));
    jdff dff_A_k2fvyJjP1_0(.din(n5014), .dout(n5017));
    jdff dff_A_WPd6hMJ60_0(.din(n5011), .dout(n5014));
    jdff dff_A_dnb8rUiS2_0(.din(n5008), .dout(n5011));
    jdff dff_A_1T43lxQM8_0(.din(n5005), .dout(n5008));
    jdff dff_A_5ibh62iE0_0(.din(n5002), .dout(n5005));
    jdff dff_A_I9x3h4qN1_0(.din(n4999), .dout(n5002));
    jdff dff_A_4aE1HHNH6_1(.din(n200), .dout(n4999));
    jdff dff_A_XNxCifA49_0(.din(n4993), .dout(G446gat));
    jdff dff_A_RUQd7QgF4_0(.din(n4990), .dout(n4993));
    jdff dff_A_1dCwUPHy5_0(.din(n4987), .dout(n4990));
    jdff dff_A_GET4LZId2_0(.din(n4984), .dout(n4987));
    jdff dff_A_r3vJIeo42_0(.din(n4981), .dout(n4984));
    jdff dff_A_J99FjoF71_0(.din(n4978), .dout(n4981));
    jdff dff_A_SURhRANd5_0(.din(n4975), .dout(n4978));
    jdff dff_A_6ngXizyP7_0(.din(n4972), .dout(n4975));
    jdff dff_A_7modmixP5_0(.din(n4969), .dout(n4972));
    jdff dff_A_9RROfpFx0_0(.din(n4966), .dout(n4969));
    jdff dff_A_VqeBgFVJ2_0(.din(n4963), .dout(n4966));
    jdff dff_A_LDyGWqCN4_0(.din(n4960), .dout(n4963));
    jdff dff_A_F2VvoqcI3_0(.din(n4957), .dout(n4960));
    jdff dff_A_QdI9JvV67_0(.din(n4954), .dout(n4957));
    jdff dff_A_Wo8dyX5s4_0(.din(n4951), .dout(n4954));
    jdff dff_A_OjT0IQyU4_0(.din(n4948), .dout(n4951));
    jdff dff_A_K9PJEWpm2_2(.din(n192), .dout(n4948));
    jdff dff_A_4EjUyHLf3_0(.din(n4942), .dout(G423gat));
    jdff dff_A_3qMyA9P25_0(.din(n4939), .dout(n4942));
    jdff dff_A_KRmvczNF6_0(.din(n4936), .dout(n4939));
    jdff dff_A_SnGkx1gH4_0(.din(n4933), .dout(n4936));
    jdff dff_A_I7IoKrtQ2_0(.din(n4930), .dout(n4933));
    jdff dff_A_zN488CAe4_0(.din(n4927), .dout(n4930));
    jdff dff_A_PJrSBVSY8_0(.din(n4924), .dout(n4927));
    jdff dff_A_ascmzqmL6_0(.din(n4921), .dout(n4924));
    jdff dff_A_nCXLlWfk0_0(.din(n4918), .dout(n4921));
    jdff dff_A_Un5Z3Ob27_0(.din(n4915), .dout(n4918));
    jdff dff_A_Teh4GM4H0_0(.din(n4912), .dout(n4915));
    jdff dff_A_lsF9shlh8_0(.din(n4909), .dout(n4912));
    jdff dff_A_4rqMQxgh1_0(.din(n4906), .dout(n4909));
    jdff dff_A_EioGrX3Z4_0(.din(n4903), .dout(n4906));
    jdff dff_A_IPn94Egd6_0(.din(n4900), .dout(n4903));
    jdff dff_A_iBunZqcK2_0(.din(n4897), .dout(n4900));
    jdff dff_A_2t4rJmJw5_0(.din(n4894), .dout(n4897));
    jdff dff_A_9xtsT3pm2_0(.din(n4891), .dout(n4894));
    jdff dff_A_398D8Blp3_2(.din(n185), .dout(n4891));
    jdff dff_A_aprmP46e1_0(.din(n4885), .dout(G422gat));
    jdff dff_A_lmZZyiBz7_0(.din(n4882), .dout(n4885));
    jdff dff_A_z7J8qGh39_0(.din(n4879), .dout(n4882));
    jdff dff_B_20dLN3zF8_2(.din(n145), .dout(n2021));
    jdff dff_B_imBdP2hB7_1(.din(n173), .dout(n2024));
    jdff dff_B_bSewn0At8_1(.din(G90gat), .dout(n2027));
    jdff dff_A_HGAmaQlw0_1(.din(n105), .dout(n2029));
    jdff dff_B_p1spw8vZ3_0(.din(n212), .dout(n2033));
    jdff dff_B_0SVk7vvA0_1(.din(G74gat), .dout(n2036));
    jdff dff_B_grGLpViM1_1(.din(G89gat), .dout(n2039));
    jdff dff_B_Ph8WKAOg1_0(.din(n260), .dout(n2042));
    jdff dff_B_rhfo69NT1_1(.din(G135gat), .dout(n2045));
    jdff dff_B_B5B76rGU8_0(.din(n244), .dout(n2048));
    jdff dff_B_0Ti6aoJG7_0(.din(n296), .dout(n2051));
    jdff dff_B_qHOAPsD99_1(.din(G207gat), .dout(n2054));
    jdff dff_B_gaEppACI8_0(.din(n280), .dout(n2057));
    jdff dff_B_QgsYS31O1_2(.din(G130gat), .dout(n2060));
    jdff dff_B_YGClbl2b5_0(.din(n483), .dout(n2063));
    jdff dff_B_O4xtUkOQ4_0(.din(n475), .dout(n2066));
    jdff dff_B_ybglk5AV2_0(.din(n2066), .dout(n2069));
    jdff dff_B_AzrEMCtS5_0(.din(n2069), .dout(n2072));
    jdff dff_B_p8U5SauZ6_0(.din(n471), .dout(n2075));
    jdff dff_B_ixm5HORf2_0(.din(n2075), .dout(n2078));
    jdff dff_B_1Ckw5jTi5_0(.din(n2078), .dout(n2081));
    jdff dff_B_9ONUZyXy5_0(.din(n435), .dout(n2084));
    jdff dff_B_5sfbu1df6_0(.din(n2084), .dout(n2087));
    jdff dff_B_gsRf9kRE5_0(.din(n2087), .dout(n2090));
    jdff dff_B_ay7CdLwp0_0(.din(n2090), .dout(n2093));
    jdff dff_B_lCubPa2y6_0(.din(n2093), .dout(n2096));
    jdff dff_B_e4tEbFwq7_0(.din(n2096), .dout(n2099));
    jdff dff_A_uyBtC1KM4_1(.din(n2104), .dout(n2101));
    jdff dff_A_d02kyb4O8_1(.din(n2107), .dout(n2104));
    jdff dff_A_zG0SrBk54_1(.din(n2110), .dout(n2107));
    jdff dff_A_NsjjrEY33_1(.din(n2113), .dout(n2110));
    jdff dff_A_BU2ztQuX6_1(.din(n2116), .dout(n2113));
    jdff dff_A_d5I7JrIA4_1(.din(n2119), .dout(n2116));
    jdff dff_A_y8SpNbTV6_1(.din(n2122), .dout(n2119));
    jdff dff_A_91NrIlWL9_1(.din(G201gat), .dout(n2122));
    jdff dff_B_gLJK9rfG7_0(.din(n721), .dout(n2126));
    jdff dff_B_wqovFkR87_0(.din(n2126), .dout(n2129));
    jdff dff_B_IFrpMZ5N0_0(.din(n2129), .dout(n2132));
    jdff dff_B_buhThgss7_0(.din(n2132), .dout(n2135));
    jdff dff_B_AHzH8W2L4_0(.din(n2135), .dout(n2138));
    jdff dff_B_T8PDaqa59_0(.din(n713), .dout(n2141));
    jdff dff_B_GiovWExW0_0(.din(n2141), .dout(n2144));
    jdff dff_B_gbJbg8IZ7_0(.din(n2144), .dout(n2147));
    jdff dff_B_9pbRBZMr3_0(.din(n709), .dout(n2150));
    jdff dff_B_5yE5FOPw1_0(.din(n2150), .dout(n2153));
    jdff dff_B_eny3aYSx1_0(.din(n2153), .dout(n2156));
    jdff dff_B_TBYpJrwa5_0(.din(n2156), .dout(n2159));
    jdff dff_B_LlKdc5LR6_0(.din(n697), .dout(n2162));
    jdff dff_B_Lq3Kd2KJ5_0(.din(n2162), .dout(n2165));
    jdff dff_B_Rhy7Vwpy6_0(.din(n2165), .dout(n2168));
    jdff dff_B_0X2DTZyU9_0(.din(n2168), .dout(n2171));
    jdff dff_B_2KGvhXHX7_0(.din(n2171), .dout(n2174));
    jdff dff_B_PkuvAbhw4_0(.din(n2174), .dout(n2177));
    jdff dff_A_71SzKjgp3_0(.din(n2182), .dout(n2179));
    jdff dff_A_kMQa9KPt0_0(.din(n2185), .dout(n2182));
    jdff dff_A_r5yEQohJ0_0(.din(n2188), .dout(n2185));
    jdff dff_A_kfV1ScLC4_0(.din(n3299), .dout(n2188));
    jdff dff_B_ARNxSAtR9_1(.din(n510), .dout(n2192));
    jdff dff_B_44Lon0vO1_1(.din(n2192), .dout(n2195));
    jdff dff_B_3aKBqgG15_1(.din(n2195), .dout(n2198));
    jdff dff_B_OnGJBMIS9_1(.din(n2198), .dout(n2201));
    jdff dff_A_dqYIZIoN4_1(.din(n2206), .dout(n2203));
    jdff dff_A_bPr74adn8_1(.din(n2209), .dout(n2206));
    jdff dff_A_2i2VcIGE8_1(.din(n2212), .dout(n2209));
    jdff dff_A_zrKGkpZa4_1(.din(n507), .dout(n2212));
    jdff dff_A_3j60n8el0_0(.din(n2218), .dout(n2215));
    jdff dff_A_KjYrMeKG1_0(.din(n2221), .dout(n2218));
    jdff dff_A_U55PGDX44_0(.din(n2224), .dout(n2221));
    jdff dff_A_p6xXJuug1_0(.din(n2227), .dout(n2224));
    jdff dff_A_hHVkuQgB7_0(.din(n2230), .dout(n2227));
    jdff dff_A_aumyIOC68_0(.din(n2233), .dout(n2230));
    jdff dff_A_zlP5GoH65_0(.din(n2236), .dout(n2233));
    jdff dff_A_8UXupTrs7_0(.din(G183gat), .dout(n2236));
    jdff dff_B_jKblZ1Io3_0(.din(n803), .dout(n2240));
    jdff dff_B_4Oh6NWAF2_0(.din(n2240), .dout(n2243));
    jdff dff_B_K1mWKtft0_0(.din(n2243), .dout(n2246));
    jdff dff_B_AC8deFa16_0(.din(n2246), .dout(n2249));
    jdff dff_B_Azjf68mi8_0(.din(n2249), .dout(n2252));
    jdff dff_B_PwwxRCIU4_0(.din(n795), .dout(n2255));
    jdff dff_B_PKOBX8gL3_0(.din(n2255), .dout(n2258));
    jdff dff_B_Z8JMqWBH9_0(.din(n2258), .dout(n2261));
    jdff dff_B_RGC0gZks6_0(.din(n791), .dout(n2264));
    jdff dff_B_2ewSbTsW5_0(.din(n2264), .dout(n2267));
    jdff dff_B_MniE1BeU3_0(.din(n2267), .dout(n2270));
    jdff dff_B_MPxPuv9U3_0(.din(n771), .dout(n2273));
    jdff dff_B_1B1che8B6_0(.din(n2273), .dout(n2276));
    jdff dff_B_utPzGWY18_0(.din(n2276), .dout(n2279));
    jdff dff_B_hM4RozQr3_0(.din(n2279), .dout(n2282));
    jdff dff_B_UNzA1csy7_0(.din(n2282), .dout(n2285));
    jdff dff_B_AHbSZy1E6_0(.din(n2285), .dout(n2288));
    jdff dff_B_jlP1OLvK8_1(.din(n732), .dout(n2291));
    jdff dff_B_sCrphbuU2_1(.din(n2291), .dout(n2294));
    jdff dff_B_LSni4cBE7_1(.din(n2294), .dout(n2297));
    jdff dff_B_5g2hOEDC3_1(.din(n2297), .dout(n2300));
    jdff dff_A_GrPBqO918_1(.din(n2305), .dout(n2302));
    jdff dff_A_bnscJa248_1(.din(n2308), .dout(n2305));
    jdff dff_A_DxyktazZ8_1(.din(n2311), .dout(n2308));
    jdff dff_A_9rSqPCBT7_1(.din(n729), .dout(n2311));
    jdff dff_B_e5bnfAO46_0(.din(n874), .dout(n2315));
    jdff dff_B_bkPu8vnq1_0(.din(n2315), .dout(n2318));
    jdff dff_B_mXZ9OooB6_0(.din(n2318), .dout(n2321));
    jdff dff_B_Yf4oWFVd6_0(.din(n866), .dout(n2324));
    jdff dff_B_7Nw6Hepr2_0(.din(n2324), .dout(n2327));
    jdff dff_B_mM67qCh82_0(.din(n2327), .dout(n2330));
    jdff dff_B_HOwL5CEw0_0(.din(n862), .dout(n2333));
    jdff dff_B_ovZcmco80_0(.din(n2333), .dout(n2336));
    jdff dff_B_UbIOBVj62_0(.din(n2336), .dout(n2339));
    jdff dff_B_EDmjy9Uf2_0(.din(n842), .dout(n2342));
    jdff dff_B_CKNTQsoL2_0(.din(n2342), .dout(n2345));
    jdff dff_B_BLQanJGl2_0(.din(n2345), .dout(n2348));
    jdff dff_B_XHEiAOyR0_0(.din(n2348), .dout(n2351));
    jdff dff_B_8BqY0Q968_0(.din(n2351), .dout(n2354));
    jdff dff_B_NLR683bv2_0(.din(n2354), .dout(n2357));
    jdff dff_B_4Uma8bE48_0(.din(n814), .dout(n2360));
    jdff dff_B_htQwsgFs6_0(.din(n2360), .dout(n2363));
    jdff dff_A_HLvrnQlk3_1(.din(n2368), .dout(n2365));
    jdff dff_A_XRHeV7YM6_1(.din(n811), .dout(n2368));
    jdff dff_B_9xZT2iRI4_1(.din(n918), .dout(n2372));
    jdff dff_B_pHcCZFPs0_1(.din(n2372), .dout(n2375));
    jdff dff_B_vRnS05bD7_1(.din(n2375), .dout(n2378));
    jdff dff_B_nwHzjng78_1(.din(n2378), .dout(n2381));
    jdff dff_B_Zawc3RUZ2_1(.din(n2381), .dout(n2384));
    jdff dff_B_taifWXKy4_1(.din(n2384), .dout(n2387));
    jdff dff_B_aWax5gil0_1(.din(n2387), .dout(n2390));
    jdff dff_B_ekJRrZl70_1(.din(n2390), .dout(n2393));
    jdff dff_B_FJtONLbG5_1(.din(n2393), .dout(n2396));
    jdff dff_B_Vu62d98T6_1(.din(n2396), .dout(n2399));
    jdff dff_B_x8TNGM6s2_1(.din(n922), .dout(n2402));
    jdff dff_B_bmBLbOZ03_1(.din(n2402), .dout(n2405));
    jdff dff_B_E54BZqYM6_1(.din(n2405), .dout(n2408));
    jdff dff_B_QG6DV6Jm6_1(.din(n2408), .dout(n2411));
    jdff dff_B_ZZklmh1s0_1(.din(n2411), .dout(n2414));
    jdff dff_B_ht8GZpwO0_1(.din(n2414), .dout(n2417));
    jdff dff_B_91k8CrMr2_1(.din(n2417), .dout(n2420));
    jdff dff_B_Gu84OHbr3_1(.din(n2420), .dout(n2423));
    jdff dff_B_bCNiqDY01_1(.din(n2423), .dout(n2426));
    jdff dff_A_zOBPkLcQ4_0(.din(n2431), .dout(n2428));
    jdff dff_A_MWDaFW5U3_0(.din(n2434), .dout(n2431));
    jdff dff_A_EH6Ydh4c5_0(.din(n2437), .dout(n2434));
    jdff dff_A_W3Rzjnlm1_0(.din(n2440), .dout(n2437));
    jdff dff_A_YUbiW5946_0(.din(n2443), .dout(n2440));
    jdff dff_A_QxkZQQRA3_0(.din(n2446), .dout(n2443));
    jdff dff_A_Gk5jogLs6_0(.din(G159gat), .dout(n2446));
    jdff dff_B_8FQ52lYY8_0(.din(n1156), .dout(n2450));
    jdff dff_B_IX1kvsFC3_0(.din(n2450), .dout(n2453));
    jdff dff_B_RcHhDRc17_0(.din(n2453), .dout(n2456));
    jdff dff_B_l8StTNXe4_0(.din(n2456), .dout(n2459));
    jdff dff_B_pXwGRbk69_0(.din(n2459), .dout(n2462));
    jdff dff_B_hZSntnMI9_0(.din(n2462), .dout(n2465));
    jdff dff_B_WFQYmM1L3_0(.din(n2465), .dout(n2468));
    jdff dff_B_TaQMXKwf6_0(.din(n2468), .dout(n2471));
    jdff dff_B_QRwLWZYo2_0(.din(n1148), .dout(n2474));
    jdff dff_B_vwu3chqa7_0(.din(n2474), .dout(n2477));
    jdff dff_B_9JYDDdE36_0(.din(n1144), .dout(n2480));
    jdff dff_B_smpALfaa5_0(.din(n2480), .dout(n2483));
    jdff dff_B_iJ5QzUeg2_0(.din(n2483), .dout(n2486));
    jdff dff_B_XSfu6jy41_0(.din(n2486), .dout(n2489));
    jdff dff_B_iq5ceS9A8_0(.din(n1132), .dout(n2492));
    jdff dff_B_3I4pFtGl9_0(.din(n2492), .dout(n2495));
    jdff dff_B_bjeD6pub3_0(.din(n2495), .dout(n2498));
    jdff dff_B_7KXbOgVN3_0(.din(n2498), .dout(n2501));
    jdff dff_B_939bfeFA6_0(.din(n2501), .dout(n2504));
    jdff dff_A_qpejjR656_1(.din(n3239), .dout(n2506));
    jdff dff_A_ZGrPnzK36_2(.din(n3239), .dout(n2509));
    jdff dff_A_azNFpMhM8_0(.din(n2515), .dout(n2512));
    jdff dff_A_e7CKnUIu7_0(.din(n2518), .dout(n2515));
    jdff dff_A_T9jjpiEI2_0(.din(n2521), .dout(n2518));
    jdff dff_A_2ubPBvQG8_0(.din(n3265), .dout(n2521));
    jdff dff_A_dY5lbPeH2_2(.din(n2527), .dout(n2524));
    jdff dff_A_Y0KSzmJG1_2(.din(n3265), .dout(n2527));
    jdff dff_B_ocmLXuYB1_0(.din(n1104), .dout(n2531));
    jdff dff_B_QSNp8d8W0_0(.din(n2531), .dout(n2534));
    jdff dff_B_x1gLVjkK1_0(.din(n2534), .dout(n2537));
    jdff dff_B_8nRvfffo3_0(.din(n2537), .dout(n2540));
    jdff dff_B_UgI77JXC7_0(.din(n2540), .dout(n2543));
    jdff dff_B_8vVYtivF3_0(.din(n2543), .dout(n2546));
    jdff dff_B_ZATPpVoE5_0(.din(n2546), .dout(n2549));
    jdff dff_A_Hf4R2y4P9_1(.din(n2554), .dout(n2551));
    jdff dff_A_fnZaLzfw6_1(.din(n2557), .dout(n2554));
    jdff dff_A_iAJ93bts7_1(.din(n2560), .dout(n2557));
    jdff dff_A_izT8ZUpC3_1(.din(n2563), .dout(n2560));
    jdff dff_A_wUV9aZlo1_1(.din(n2566), .dout(n2563));
    jdff dff_A_7x4rsCSo3_1(.din(n2569), .dout(n2566));
    jdff dff_A_3Y6MdOJP6_1(.din(n1101), .dout(n2569));
    jdff dff_B_YP1ptw8m1_0(.din(n1233), .dout(n2573));
    jdff dff_B_qyAHTwhB0_0(.din(n2573), .dout(n2576));
    jdff dff_B_34uARqsn6_0(.din(n2576), .dout(n2579));
    jdff dff_B_vQMMS74M7_0(.din(n2579), .dout(n2582));
    jdff dff_B_6429jJEN6_0(.din(n2582), .dout(n2585));
    jdff dff_B_oC0b5SRv8_0(.din(n2585), .dout(n2588));
    jdff dff_B_hZWEU94y7_0(.din(n2588), .dout(n2591));
    jdff dff_B_AfRRtiyr7_0(.din(n2591), .dout(n2594));
    jdff dff_B_Fo1aHILk9_0(.din(n2594), .dout(n2597));
    jdff dff_B_Izf4783V0_0(.din(n2597), .dout(n2600));
    jdff dff_B_ym3pvic20_0(.din(n1225), .dout(n2603));
    jdff dff_B_MIHLAari6_0(.din(n2603), .dout(n2606));
    jdff dff_B_YtlP2FKE4_0(.din(n1221), .dout(n2609));
    jdff dff_B_Tcu6c5IJ4_0(.din(n2609), .dout(n2612));
    jdff dff_B_sgHWmJTp7_0(.din(n2612), .dout(n2615));
    jdff dff_B_jjcIAjEI9_0(.din(n2615), .dout(n2618));
    jdff dff_B_hgt6o9t34_0(.din(n1209), .dout(n2621));
    jdff dff_B_MlJi8swA5_0(.din(n2621), .dout(n2624));
    jdff dff_B_3DYU1nwt0_0(.din(n2624), .dout(n2627));
    jdff dff_B_utkHbiUL4_0(.din(n2627), .dout(n2630));
    jdff dff_B_Wh4Yu1TF4_0(.din(n2630), .dout(n2633));
    jdff dff_B_lQd04rdX2_0(.din(n1181), .dout(n2636));
    jdff dff_B_T9QDIIpq3_0(.din(n2636), .dout(n2639));
    jdff dff_B_sBvHmArP9_0(.din(n2639), .dout(n2642));
    jdff dff_B_1TRPL6zQ8_0(.din(n2642), .dout(n2645));
    jdff dff_B_2dDd7thp5_0(.din(n2645), .dout(n2648));
    jdff dff_B_cN5Fl1bl3_0(.din(n2648), .dout(n2651));
    jdff dff_B_lNQigljw6_0(.din(n2651), .dout(n2654));
    jdff dff_B_9qONROA47_0(.din(n2654), .dout(n2657));
    jdff dff_B_PNoVvop11_0(.din(n2657), .dout(n2660));
    jdff dff_A_GGqPTmaf8_1(.din(n2665), .dout(n2662));
    jdff dff_A_qJlR1Via2_1(.din(n2668), .dout(n2665));
    jdff dff_A_1c6f6JN29_1(.din(n2671), .dout(n2668));
    jdff dff_A_fYQhOLMb1_1(.din(n2674), .dout(n2671));
    jdff dff_A_PuEJQdU62_1(.din(n2677), .dout(n2674));
    jdff dff_A_glE6YjOI9_1(.din(n2680), .dout(n2677));
    jdff dff_A_DD5VzlQI2_1(.din(n2683), .dout(n2680));
    jdff dff_A_yLKQHjhw5_1(.din(n2686), .dout(n2683));
    jdff dff_A_zguWoSTU8_1(.din(n1178), .dout(n2686));
    jdff dff_B_Njars19K6_1(.din(n894), .dout(n2690));
    jdff dff_B_T1w9DNB23_1(.din(n2690), .dout(n2693));
    jdff dff_B_nBOiScYI3_1(.din(n2693), .dout(n2696));
    jdff dff_A_3NFqrWk85_1(.din(n2701), .dout(n2698));
    jdff dff_A_XJ75fKMM1_1(.din(n2704), .dout(n2701));
    jdff dff_A_4sauANMr5_1(.din(n2707), .dout(n2704));
    jdff dff_A_5Rc1NTn82_1(.din(n2710), .dout(n2707));
    jdff dff_A_22EzaNRH2_1(.din(n2713), .dout(n2710));
    jdff dff_A_YFVx8Hve1_1(.din(n2716), .dout(n2713));
    jdff dff_A_3CXBDjGy9_1(.din(G159gat), .dout(n2716));
    jdff dff_A_ONychntC1_2(.din(n2722), .dout(n2719));
    jdff dff_A_4GwYeHZU7_2(.din(n2725), .dout(n2722));
    jdff dff_A_rZWI63BR4_2(.din(n2728), .dout(n2725));
    jdff dff_A_rCHswxiA2_2(.din(n2731), .dout(n2728));
    jdff dff_A_4CYVFgmW9_2(.din(n2734), .dout(n2731));
    jdff dff_A_1b3pr0Eu8_2(.din(n2737), .dout(n2734));
    jdff dff_A_pFZYmTHO8_2(.din(G159gat), .dout(n2737));
    jdff dff_A_7j1cYmm35_2(.din(n2743), .dout(n2740));
    jdff dff_A_7QNwRjLL8_2(.din(n2746), .dout(n2743));
    jdff dff_A_VALLlZDi7_2(.din(n2749), .dout(n2746));
    jdff dff_A_Y7MJgL9w2_2(.din(G159gat), .dout(n2749));
    jdff dff_B_fI6OMezF4_0(.din(n1170), .dout(n2753));
    jdff dff_B_PUoCACqF5_0(.din(n2753), .dout(n2756));
    jdff dff_B_FCcmQtCQ5_0(.din(n2756), .dout(n2759));
    jdff dff_B_WjlhjVFz8_0(.din(n2759), .dout(n2762));
    jdff dff_A_L73bfKqD5_1(.din(n2767), .dout(n2764));
    jdff dff_A_QRSBxjvm0_1(.din(n2770), .dout(n2767));
    jdff dff_A_smHjJcy14_1(.din(n2773), .dout(n2770));
    jdff dff_A_AbClJDsC1_1(.din(n1071), .dout(n2773));
    jdff dff_B_JLFDRsbE1_1(.din(n1047), .dout(n2777));
    jdff dff_B_TI3tV9FD4_1(.din(n2777), .dout(n2780));
    jdff dff_B_6W5xi0fm4_1(.din(n2780), .dout(n2783));
    jdff dff_B_mLJ7Ql8H6_0(.din(n1163), .dout(n2786));
    jdff dff_B_7URkGVGW8_0(.din(n2786), .dout(n2789));
    jdff dff_B_EPuOvwon3_0(.din(n2789), .dout(n2792));
    jdff dff_B_LpuWcMhc0_0(.din(n2792), .dout(n2795));
    jdff dff_A_d5WapaAd8_1(.din(n2800), .dout(n2797));
    jdff dff_A_j39aCgnn3_1(.din(n2803), .dout(n2800));
    jdff dff_A_Aga2VbG81_1(.din(n2806), .dout(n2803));
    jdff dff_A_W22bFRvE6_1(.din(n1039), .dout(n2806));
    jdff dff_B_OJKZr1Pa1_1(.din(n941), .dout(n2810));
    jdff dff_B_VE2PbU0n4_1(.din(n2810), .dout(n2813));
    jdff dff_B_PdEw4Pai8_1(.din(n2813), .dout(n2816));
    jdff dff_B_YbtlO2aU0_1(.din(n2816), .dout(n2819));
    jdff dff_B_U9yoAtHN1_1(.din(n2819), .dout(n2822));
    jdff dff_B_UsVqLjAM8_1(.din(n2822), .dout(n2825));
    jdff dff_B_pRJznE1q4_1(.din(n2825), .dout(n2828));
    jdff dff_B_CO0TEYyV5_0(.din(n1318), .dout(n2831));
    jdff dff_B_RfywZe636_0(.din(n2831), .dout(n2834));
    jdff dff_B_7q6IeY6F4_0(.din(n2834), .dout(n2837));
    jdff dff_B_R2TlDJIS9_0(.din(n2837), .dout(n2840));
    jdff dff_B_V8mtbQ7e9_0(.din(n2840), .dout(n2843));
    jdff dff_B_KiN71b3D9_0(.din(n2843), .dout(n2846));
    jdff dff_B_Feks7tyM3_0(.din(n2846), .dout(n2849));
    jdff dff_B_pD7DtAH65_0(.din(n2849), .dout(n2852));
    jdff dff_B_PxDM8Pdk2_0(.din(n2852), .dout(n2855));
    jdff dff_B_knFNQfaJ1_0(.din(n2855), .dout(n2858));
    jdff dff_B_TkBwFMYm3_0(.din(n1310), .dout(n2861));
    jdff dff_B_2spQn6sk2_0(.din(n2861), .dout(n2864));
    jdff dff_B_mKHVLYLl6_0(.din(n1306), .dout(n2867));
    jdff dff_B_r4tmjpNV0_0(.din(n2867), .dout(n2870));
    jdff dff_B_MBICdgy26_0(.din(n2870), .dout(n2873));
    jdff dff_B_qyXVzmYJ7_0(.din(n2873), .dout(n2876));
    jdff dff_A_hA9yRRx98_1(.din(n2881), .dout(n2878));
    jdff dff_A_EKF1ZGSF3_1(.din(n2884), .dout(n2881));
    jdff dff_A_hBLY9SOv4_1(.din(n2887), .dout(n2884));
    jdff dff_A_pBohs5H37_1(.din(n2890), .dout(n2887));
    jdff dff_A_6LWhfFPr7_1(.din(G91gat), .dout(n2890));
    jdff dff_B_cB1AxH6V7_0(.din(n1294), .dout(n2894));
    jdff dff_B_KKaxXAic3_0(.din(n2894), .dout(n2897));
    jdff dff_B_CH4j4C5Y7_0(.din(n2897), .dout(n2900));
    jdff dff_B_ZAcBpBG22_0(.din(n2900), .dout(n2903));
    jdff dff_B_GJ3Zrlbj5_0(.din(n2903), .dout(n2906));
    jdff dff_B_t4CSkoIp3_1(.din(n1244), .dout(n2909));
    jdff dff_B_ow44jL611_1(.din(n2909), .dout(n2912));
    jdff dff_B_N35O9IcH8_1(.din(n2912), .dout(n2915));
    jdff dff_B_U8Jo871b9_1(.din(n2915), .dout(n2918));
    jdff dff_B_efg2qdYU1_1(.din(n2918), .dout(n2921));
    jdff dff_B_emH93ejM9_1(.din(n2921), .dout(n2924));
    jdff dff_B_mrW5kCZ85_1(.din(n2924), .dout(n2927));
    jdff dff_B_HQAup70o0_1(.din(n2927), .dout(n2930));
    jdff dff_B_OelSTeiU1_1(.din(n2930), .dout(n2933));
    jdff dff_B_mZuN47YQ3_1(.din(n1247), .dout(n2936));
    jdff dff_B_Jr5ZHMyQ0_1(.din(n2936), .dout(n2939));
    jdff dff_B_kn2ms3Rz5_1(.din(n2939), .dout(n2942));
    jdff dff_B_q4xEbWFW2_1(.din(n2942), .dout(n2945));
    jdff dff_B_QNGxCLSY9_1(.din(n2945), .dout(n2948));
    jdff dff_B_fkPCQbba7_1(.din(n2948), .dout(n2951));
    jdff dff_B_AlOKLYwV3_0(.din(n1250), .dout(n2954));
    jdff dff_B_FvY63EkL9_0(.din(n2954), .dout(n2957));
    jdff dff_B_fNYjGCB03_0(.din(n2957), .dout(n2960));
    jdff dff_B_f84puu9g0_0(.din(n2960), .dout(n2963));
    jdff dff_B_4z0SVa6o3_0(.din(n2963), .dout(n2966));
    jdff dff_B_3XQtlWSc7_0(.din(n2966), .dout(n2969));
    jdff dff_A_D5s9Hsp36_0(.din(n2974), .dout(n2971));
    jdff dff_A_3VFNgtBl1_0(.din(n2977), .dout(n2974));
    jdff dff_A_eiCg0iHe0_0(.din(n2980), .dout(n2977));
    jdff dff_A_YwyFruk58_0(.din(n2983), .dout(n2980));
    jdff dff_A_J8mq48JQ0_0(.din(n2986), .dout(n2983));
    jdff dff_A_dfDj8RWL9_0(.din(n1035), .dout(n2986));
    jdff dff_A_KbcVS7sh7_2(.din(n1035), .dout(n2989));
    jdff dff_A_KnGvYnNg0_0(.din(n2995), .dout(n2992));
    jdff dff_A_rIpQowp34_0(.din(n2998), .dout(n2995));
    jdff dff_A_qJKfoSUw4_0(.din(n3001), .dout(n2998));
    jdff dff_A_bPA3mF5m3_0(.din(n3004), .dout(n3001));
    jdff dff_A_90RkIKWw4_0(.din(n3007), .dout(n3004));
    jdff dff_A_wS7nXe1t7_0(.din(n1063), .dout(n3007));
    jdff dff_B_lkdbdiPE2_1(.din(n1051), .dout(n3011));
    jdff dff_A_Ko2xzVei3_0(.din(n3016), .dout(n3013));
    jdff dff_A_wuiXzE2p2_0(.din(n3019), .dout(n3016));
    jdff dff_A_5xkH4MHd4_0(.din(n3022), .dout(n3019));
    jdff dff_A_oLAu9PgN6_0(.din(n3025), .dout(n3022));
    jdff dff_A_DmMZkXHQ6_0(.din(n3028), .dout(n3025));
    jdff dff_A_UoymzHYZ3_0(.din(n3031), .dout(n3028));
    jdff dff_A_KPkjkTHf0_0(.din(G171gat), .dout(n3031));
    jdff dff_A_iKnk4anM6_1(.din(n3037), .dout(n3034));
    jdff dff_A_ddbxkrov7_1(.din(n3040), .dout(n3037));
    jdff dff_A_Y1Bdosnl9_1(.din(n3043), .dout(n3040));
    jdff dff_A_diCDEsHX2_1(.din(n3046), .dout(n3043));
    jdff dff_A_RVw0n8sK9_1(.din(n3049), .dout(n3046));
    jdff dff_A_pndzv8ct0_1(.din(n3052), .dout(n3049));
    jdff dff_A_yMQ6iL6S3_1(.din(n3055), .dout(n3052));
    jdff dff_A_alIZJUzz0_1(.din(n3058), .dout(n3055));
    jdff dff_A_UJ7N9NOf9_1(.din(n1241), .dout(n3058));
    jdff dff_B_5CABIsTw2_0(.din(n953), .dout(n3062));
    jdff dff_B_TjBTKXoi7_0(.din(n3062), .dout(n3065));
    jdff dff_B_i5cAmkLc7_0(.din(n3065), .dout(n3068));
    jdff dff_A_jvc0pF3Z5_1(.din(n3073), .dout(n3070));
    jdff dff_A_eJxtZOeL6_1(.din(n3076), .dout(n3073));
    jdff dff_A_j6aI7Icb3_1(.din(n3079), .dout(n3076));
    jdff dff_A_lTYqFZCO3_1(.din(n3082), .dout(n3079));
    jdff dff_A_TJCZ1xdI6_1(.din(n3085), .dout(n3082));
    jdff dff_A_WnLAxBC29_1(.din(n3088), .dout(n3085));
    jdff dff_A_jc7HTzSh1_1(.din(G165gat), .dout(n3088));
    jdff dff_A_bsCysOS74_2(.din(n3094), .dout(n3091));
    jdff dff_A_vFormJ3P0_2(.din(n3097), .dout(n3094));
    jdff dff_A_jxuKexFD5_2(.din(n3100), .dout(n3097));
    jdff dff_A_pIJI1wR47_2(.din(n3103), .dout(n3100));
    jdff dff_A_sbFtc1u37_2(.din(n3106), .dout(n3103));
    jdff dff_A_VaX0XcJM4_2(.din(n3109), .dout(n3106));
    jdff dff_A_5KNPP9EU7_2(.din(G165gat), .dout(n3109));
    jdff dff_A_eterAJUo3_2(.din(n3115), .dout(n3112));
    jdff dff_A_RYypYTir9_2(.din(n3118), .dout(n3115));
    jdff dff_A_7LdjYk5T4_2(.din(n3121), .dout(n3118));
    jdff dff_A_8XpGyw5C6_2(.din(G165gat), .dout(n3121));
    jdff dff_B_zeyF7S7C6_0(.din(n1403), .dout(n3125));
    jdff dff_B_i6oBulh41_0(.din(n3125), .dout(n3128));
    jdff dff_B_EgtbQ1og3_0(.din(n3128), .dout(n3131));
    jdff dff_B_uGwKqtyq4_0(.din(n3131), .dout(n3134));
    jdff dff_B_ssY13juN7_0(.din(n3134), .dout(n3137));
    jdff dff_B_3ZBUr4P26_0(.din(n3137), .dout(n3140));
    jdff dff_B_pMpnmSFT7_0(.din(n3140), .dout(n3143));
    jdff dff_B_qMGeSdpT8_0(.din(n3143), .dout(n3146));
    jdff dff_B_xXJGaZgs1_0(.din(n3146), .dout(n3149));
    jdff dff_B_bBEt4ZWG5_0(.din(n3149), .dout(n3152));
    jdff dff_B_cYhKNdA75_0(.din(n1395), .dout(n3155));
    jdff dff_B_nBQKbeDD7_0(.din(n3155), .dout(n3158));
    jdff dff_B_LovpfXDU5_0(.din(n1391), .dout(n3161));
    jdff dff_B_ANnB8LUY2_0(.din(n3161), .dout(n3164));
    jdff dff_B_z0Aue9fS2_0(.din(n3164), .dout(n3167));
    jdff dff_B_Pv1yspMa9_0(.din(n3167), .dout(n3170));
    jdff dff_A_it6uYGN15_1(.din(n3175), .dout(n3172));
    jdff dff_A_N6o8wclS5_1(.din(n3178), .dout(n3175));
    jdff dff_A_F2bI8AQq9_1(.din(n3181), .dout(n3178));
    jdff dff_A_iKwxcC1S7_1(.din(n3184), .dout(n3181));
    jdff dff_A_98YQrYo79_1(.din(G96gat), .dout(n3184));
    jdff dff_B_vTI34gNP8_1(.din(G73gat), .dout(n3188));
    jdff dff_A_LxxNHobh5_0(.din(n220), .dout(n3190));
    jdff dff_A_shD5mLGa3_0(.din(n208), .dout(n3193));
    jdff dff_B_CrHvogc18_0(.din(n1379), .dout(n3197));
    jdff dff_B_k7j50dZ35_0(.din(n3197), .dout(n3200));
    jdff dff_B_lzpiCVSF1_0(.din(n3200), .dout(n3203));
    jdff dff_B_RckJwQxV6_0(.din(n3203), .dout(n3206));
    jdff dff_B_Gm0kNzhg3_0(.din(n3206), .dout(n3209));
    jdff dff_B_0gjBhWBg7_3(.din(G246gat), .dout(n3212));
    jdff dff_A_JhAco3gd1_2(.din(n3239), .dout(n3214));
    jdff dff_B_yH1b8k1E3_3(.din(G228gat), .dout(n3218));
    jdff dff_B_ZB59Gv4L7_3(.din(n3218), .dout(n3221));
    jdff dff_B_7sgX5yrC5_3(.din(n3221), .dout(n3224));
    jdff dff_B_OdRa28TU4_3(.din(n3224), .dout(n3227));
    jdff dff_B_Wy3Gey7V3_3(.din(n3227), .dout(n3230));
    jdff dff_B_T8GuwOpR6_3(.din(n3230), .dout(n3233));
    jdff dff_B_MSA3xcpb2_3(.din(n3233), .dout(n3236));
    jdff dff_B_cunaExpD1_3(.din(n3236), .dout(n3239));
    jdff dff_A_FWaJm0wq7_0(.din(n3244), .dout(n3241));
    jdff dff_A_s3hp9UnE5_0(.din(n3247), .dout(n3244));
    jdff dff_A_RcxMbyay4_0(.din(n3250), .dout(n3247));
    jdff dff_A_XopyLnzA5_0(.din(n3253), .dout(n3250));
    jdff dff_A_yvWTABtl4_0(.din(n3256), .dout(n3253));
    jdff dff_A_ViQqoSan2_0(.din(n3259), .dout(n3256));
    jdff dff_A_dL1MpdZe6_0(.din(n3262), .dout(n3259));
    jdff dff_A_2WeA3owF7_0(.din(n3299), .dout(n3262));
    jdff dff_A_WIADCNa01_1(.din(n3268), .dout(n3265));
    jdff dff_A_j2mV2HVv6_1(.din(n3299), .dout(n3268));
    jdff dff_B_LECh1TG46_3(.din(G219gat), .dout(n3272));
    jdff dff_B_k2ACAfl64_3(.din(n3272), .dout(n3275));
    jdff dff_B_QAiyhTQn6_3(.din(n3275), .dout(n3278));
    jdff dff_B_hTK7h19Q7_3(.din(n3278), .dout(n3281));
    jdff dff_B_Wrja4ard4_3(.din(n3281), .dout(n3284));
    jdff dff_B_Zb8Mnr6N1_3(.din(n3284), .dout(n3287));
    jdff dff_B_JABA05kb4_3(.din(n3287), .dout(n3290));
    jdff dff_B_js1SSsc40_3(.din(n3290), .dout(n3293));
    jdff dff_B_iTMyeUSy8_3(.din(n3293), .dout(n3296));
    jdff dff_B_ZL8ZAyZh2_3(.din(n3296), .dout(n3299));
    jdff dff_B_NiV2AKPp7_1(.din(n1329), .dout(n3302));
    jdff dff_B_90CIGYAP8_1(.din(n3302), .dout(n3305));
    jdff dff_B_O7GIOyoc4_1(.din(n3305), .dout(n3308));
    jdff dff_B_MQ5HIeHj0_1(.din(n3308), .dout(n3311));
    jdff dff_B_ligpKIir9_1(.din(n3311), .dout(n3314));
    jdff dff_B_zy5x0kiP4_1(.din(n3314), .dout(n3317));
    jdff dff_B_VpozsdDg7_1(.din(n3317), .dout(n3320));
    jdff dff_B_2esykH8h4_1(.din(n3320), .dout(n3323));
    jdff dff_B_NLszNRtg2_1(.din(n3323), .dout(n3326));
    jdff dff_B_lYounoyC7_1(.din(n1332), .dout(n3329));
    jdff dff_B_fRQc0Ubi5_1(.din(n3329), .dout(n3332));
    jdff dff_B_PWsRhbmR1_1(.din(n3332), .dout(n3335));
    jdff dff_B_HVkZ9dnD0_1(.din(n3335), .dout(n3338));
    jdff dff_B_kHP8xzmV3_1(.din(n3338), .dout(n3341));
    jdff dff_B_0q7Y0Ifp9_1(.din(n3341), .dout(n3344));
    jdff dff_B_dvgKbKCL6_1(.din(n3344), .dout(n3347));
    jdff dff_B_QyXeecTJ0_1(.din(n3347), .dout(n3350));
    jdff dff_B_VLbt0aoS7_0(.din(n1335), .dout(n3353));
    jdff dff_B_tkk7Pp4Y7_0(.din(n3353), .dout(n3356));
    jdff dff_B_Fw2zGQ9u2_0(.din(n3356), .dout(n3359));
    jdff dff_B_u8LhLyL08_0(.din(n3359), .dout(n3362));
    jdff dff_B_3dK4KEEy6_0(.din(n3362), .dout(n3365));
    jdff dff_B_gorGpyFJ5_0(.din(n3365), .dout(n3368));
    jdff dff_B_L0320AkD2_0(.din(n3368), .dout(n3371));
    jdff dff_A_0lyqxPsZ5_0(.din(n3376), .dout(n3373));
    jdff dff_A_WzPbRMYu6_0(.din(n3379), .dout(n3376));
    jdff dff_A_tlvt9k2R0_0(.din(n3382), .dout(n3379));
    jdff dff_A_s3zgy9cj0_0(.din(n3385), .dout(n3382));
    jdff dff_A_OCJEHcr90_0(.din(n3388), .dout(n3385));
    jdff dff_A_burd5mjC4_0(.din(n3391), .dout(n3388));
    jdff dff_A_kScFJcsb4_0(.din(n1031), .dout(n3391));
    jdff dff_A_WK3aLGhH9_0(.din(n3397), .dout(n3394));
    jdff dff_A_jw1L4KQf4_0(.din(n3400), .dout(n3397));
    jdff dff_A_gF8O0kOx7_0(.din(n3403), .dout(n3400));
    jdff dff_A_h3AlJXLC9_0(.din(n3406), .dout(n3403));
    jdff dff_A_pX56OMCk2_0(.din(n3409), .dout(n3406));
    jdff dff_A_ZXyQHwlc3_0(.din(n3412), .dout(n3409));
    jdff dff_A_kPNf8Wh39_0(.din(G177gat), .dout(n3412));
    jdff dff_B_M8u8lpIW6_1(.din(n1086), .dout(n3416));
    jdff dff_B_dfzaaTg61_1(.din(n3416), .dout(n3419));
    jdff dff_B_5JtSqqhk2_1(.din(n3419), .dout(n3422));
    jdff dff_B_XEQnazf80_1(.din(n3422), .dout(n3425));
    jdff dff_B_FxFBpVrk9_1(.din(n3425), .dout(n3428));
    jdff dff_B_wJ5ruUjE4_1(.din(n1089), .dout(n3431));
    jdff dff_B_NzKj01Qv2_1(.din(n3431), .dout(n3434));
    jdff dff_B_maYxTiIJ7_1(.din(n3434), .dout(n3437));
    jdff dff_B_BU8RXXAE6_1(.din(n3437), .dout(n3440));
    jdff dff_B_zCTWHUUc0_0(.din(n645), .dout(n3443));
    jdff dff_A_U8VkxY2G1_0(.din(n642), .dout(n3445));
    jdff dff_B_HJhhk2Za1_1(.din(n630), .dout(n3449));
    jdff dff_A_yAdCop6Z3_0(.din(n3454), .dout(n3451));
    jdff dff_A_xMfnZn0I7_0(.din(n3457), .dout(n3454));
    jdff dff_A_C4oHFx8z8_0(.din(n634), .dout(n3457));
    jdff dff_A_0UYYGZAd7_1(.din(n3463), .dout(n3460));
    jdff dff_A_dKYJ5aZf9_1(.din(n3466), .dout(n3463));
    jdff dff_A_aZn7jFaW6_1(.din(n3469), .dout(n3466));
    jdff dff_A_9LjsbrFf8_1(.din(n3472), .dout(n3469));
    jdff dff_A_pF2s8jJy7_1(.din(n3475), .dout(n3472));
    jdff dff_A_VB2fzTlZ8_1(.din(n3478), .dout(n3475));
    jdff dff_A_h6fWmWR07_1(.din(n3481), .dout(n3478));
    jdff dff_A_DTUD1R403_1(.din(G195gat), .dout(n3481));
    jdff dff_A_JHMj1Keu4_2(.din(n3487), .dout(n3484));
    jdff dff_A_NaguskDQ5_2(.din(n3490), .dout(n3487));
    jdff dff_A_aZxjJvh80_2(.din(n3493), .dout(n3490));
    jdff dff_A_BjECwNAx5_2(.din(n3496), .dout(n3493));
    jdff dff_A_RqT43T9y2_2(.din(n3499), .dout(n3496));
    jdff dff_A_rCeAFLiN1_2(.din(n3502), .dout(n3499));
    jdff dff_A_Qv1SyCfy9_2(.din(n3505), .dout(n3502));
    jdff dff_A_fsxYyJjG3_2(.din(G195gat), .dout(n3505));
    jdff dff_A_t2VKqC012_1(.din(n3511), .dout(n3508));
    jdff dff_A_rKur3qzb4_1(.din(n3514), .dout(n3511));
    jdff dff_A_6FlEJPGT6_1(.din(n3517), .dout(n3514));
    jdff dff_A_8s9P6lSF8_1(.din(n3520), .dout(n3517));
    jdff dff_A_ED5y1Mrd2_1(.din(n3523), .dout(n3520));
    jdff dff_A_rG8SlCZZ8_1(.din(n3526), .dout(n3523));
    jdff dff_A_jN2amZtz9_1(.din(n3529), .dout(n3526));
    jdff dff_A_Bk71gHeV9_1(.din(G189gat), .dout(n3529));
    jdff dff_A_Ml3LPoRN6_2(.din(n3535), .dout(n3532));
    jdff dff_A_Cb2IXG5A8_2(.din(n3538), .dout(n3535));
    jdff dff_A_W7xMu0jm8_2(.din(n3541), .dout(n3538));
    jdff dff_A_U46mvkgj9_2(.din(n3544), .dout(n3541));
    jdff dff_A_KSUlxIVK5_2(.din(n3547), .dout(n3544));
    jdff dff_A_XkLLA4j06_2(.din(n3550), .dout(n3547));
    jdff dff_A_hMy2MXLM0_2(.din(n3553), .dout(n3550));
    jdff dff_A_ihUrwOyU2_2(.din(G189gat), .dout(n3553));
    jdff dff_B_7A8CQ8wf1_0(.din(n622), .dout(n3557));
    jdff dff_A_c2yYKDc01_0(.din(n619), .dout(n3559));
    jdff dff_A_WkSOeeeh6_0(.din(n3565), .dout(n3562));
    jdff dff_A_EEBKWNz20_0(.din(n615), .dout(n3565));
    jdff dff_B_rRvGpYtZ9_1(.din(n599), .dout(n3569));
    jdff dff_A_v5nfyNWc3_0(.din(n3574), .dout(n3571));
    jdff dff_A_Eq6Muw3W5_0(.din(n3577), .dout(n3574));
    jdff dff_A_VQx0RyiS8_0(.din(n3580), .dout(n3577));
    jdff dff_A_OKECXWQi5_0(.din(n3583), .dout(n3580));
    jdff dff_A_fyBPgIOs4_0(.din(G121gat), .dout(n3583));
    jdff dff_A_7WBawzON4_0(.din(n3589), .dout(n3586));
    jdff dff_A_QmSLiku04_0(.din(n3592), .dout(n3589));
    jdff dff_A_xFXitK0D6_0(.din(n3595), .dout(n3592));
    jdff dff_A_ksId0XEv9_0(.din(n3598), .dout(n3595));
    jdff dff_A_3C6fbs1i9_0(.din(n3601), .dout(n3598));
    jdff dff_A_FMfH9g317_0(.din(n3604), .dout(n3601));
    jdff dff_A_9XhzZTb43_0(.din(n3607), .dout(n3604));
    jdff dff_A_IpqDrjdh0_0(.din(G195gat), .dout(n3607));
    jdff dff_A_HZkf69Kn8_2(.din(n3613), .dout(n3610));
    jdff dff_A_jrjUOp1I0_2(.din(n3616), .dout(n3613));
    jdff dff_A_vn9IGqtz7_2(.din(n3619), .dout(n3616));
    jdff dff_A_7tnFYHLD3_2(.din(G195gat), .dout(n3619));
    jdff dff_B_HP1pRa9y2_1(.din(n579), .dout(n3623));
    jdff dff_A_K4JB3bi80_1(.din(n3628), .dout(n3625));
    jdff dff_A_rLOPMm421_1(.din(n3631), .dout(n3628));
    jdff dff_A_O2Gy59Yd5_1(.din(n3634), .dout(n3631));
    jdff dff_A_eNwx5A8U0_1(.din(n3637), .dout(n3634));
    jdff dff_A_4J4xqKLW5_1(.din(G116gat), .dout(n3637));
    jdff dff_A_kvfY68hY2_1(.din(n3653), .dout(n3640));
    jdff dff_B_g8xrYXn64_2(.din(G146gat), .dout(n3644));
    jdff dff_B_ZDNC6rPy5_2(.din(n3644), .dout(n3647));
    jdff dff_B_LrlYXd8T1_2(.din(n3647), .dout(n3650));
    jdff dff_B_piD0i7Xt2_2(.din(n3650), .dout(n3653));
    jdff dff_A_avSQB05u4_0(.din(n3658), .dout(n3655));
    jdff dff_A_ohMpxTvy5_0(.din(n3661), .dout(n3658));
    jdff dff_A_18xIItvs4_0(.din(n3664), .dout(n3661));
    jdff dff_A_ZJEF9ZSQ7_0(.din(n3667), .dout(n3664));
    jdff dff_A_uLTmUqcE9_0(.din(n3670), .dout(n3667));
    jdff dff_A_gAhvSEBA2_0(.din(n3673), .dout(n3670));
    jdff dff_A_5MuUyKNx9_0(.din(n3676), .dout(n3673));
    jdff dff_A_PNmlGw7p8_0(.din(G189gat), .dout(n3676));
    jdff dff_A_WKhiULLH2_2(.din(n3682), .dout(n3679));
    jdff dff_A_3evzTTmu8_2(.din(n3685), .dout(n3682));
    jdff dff_A_oqqOtPtr9_2(.din(n3688), .dout(n3685));
    jdff dff_A_7awGszEe9_2(.din(G189gat), .dout(n3688));
    jdff dff_B_Bj9Xhqiq0_1(.din(n517), .dout(n3692));
    jdff dff_B_YWJF9daW1_1(.din(n520), .dout(n3695));
    jdff dff_B_0aZHIupd6_1(.din(n3695), .dout(n3698));
    jdff dff_B_zp8Q2MNX9_1(.din(n3698), .dout(n3701));
    jdff dff_B_Scid7VSd1_1(.din(n3701), .dout(n3704));
    jdff dff_B_6QO0Oz3U5_1(.din(n3704), .dout(n3707));
    jdff dff_B_kboDXVne9_1(.din(n3707), .dout(n3710));
    jdff dff_B_l3EjJiUZ8_1(.din(n3710), .dout(n3713));
    jdff dff_B_skd7gkZr8_1(.din(n3713), .dout(n3716));
    jdff dff_B_CRE4zai05_1(.din(n523), .dout(n3719));
    jdff dff_B_aaNCrRes6_0(.din(n555), .dout(n3722));
    jdff dff_B_teIs8hoA6_0(.din(n3722), .dout(n3725));
    jdff dff_B_F6Wksyvu4_1(.din(n526), .dout(n3728));
    jdff dff_B_Ji6T9NuC1_1(.din(n3728), .dout(n3731));
    jdff dff_B_1maUqPPy8_1(.din(n3731), .dout(n3734));
    jdff dff_B_aGrgTfJx5_1(.din(n3734), .dout(n3737));
    jdff dff_B_308swCCT8_1(.din(n3737), .dout(n3740));
    jdff dff_B_WHqEB5UA4_1(.din(n529), .dout(n3743));
    jdff dff_B_RgedzBox4_1(.din(n3743), .dout(n3746));
    jdff dff_B_zcWU9T686_1(.din(n3746), .dout(n3749));
    jdff dff_B_CEyhQme00_1(.din(n532), .dout(n3752));
    jdff dff_B_OT2NGZCo5_2(.din(n307), .dout(n3755));
    jdff dff_B_o62SLLAi8_2(.din(n3755), .dout(n3758));
    jdff dff_B_weoeNh1Z2_2(.din(n3758), .dout(n3761));
    jdff dff_B_QLqm9Rjl5_2(.din(n3761), .dout(n3764));
    jdff dff_B_fqdGfhSa0_2(.din(n3764), .dout(n3767));
    jdff dff_B_jlAjge222_2(.din(n3767), .dout(n3770));
    jdff dff_B_PNREf1H55_2(.din(n3770), .dout(n3773));
    jdff dff_B_O7IYYnW93_2(.din(n3773), .dout(n3776));
    jdff dff_B_W8buxaVQ2_2(.din(n3776), .dout(n3779));
    jdff dff_A_eI1hEaNQ3_0(.din(n3784), .dout(n3781));
    jdff dff_A_eEZuc3JX5_0(.din(n3787), .dout(n3784));
    jdff dff_A_gzGnGGAu2_0(.din(n3790), .dout(n3787));
    jdff dff_A_BXzaIjEq7_0(.din(n3793), .dout(n3790));
    jdff dff_A_6N9GaMhU6_0(.din(n3796), .dout(n3793));
    jdff dff_A_PqkO6H438_0(.din(n3799), .dout(n3796));
    jdff dff_A_MDCxWnEX0_0(.din(n3802), .dout(n3799));
    jdff dff_A_SkK6WUdn5_0(.din(n3805), .dout(n3802));
    jdff dff_A_EPD7r3wi6_0(.din(G261gat), .dout(n3805));
    jdff dff_A_Zx2Dsoyo2_1(.din(n3811), .dout(n3808));
    jdff dff_A_xVZx3eOO5_1(.din(n3814), .dout(n3811));
    jdff dff_A_yy4Xcum80_1(.din(n3817), .dout(n3814));
    jdff dff_A_IKIePTK22_1(.din(n3820), .dout(n3817));
    jdff dff_A_xCoL9wn42_1(.din(n3823), .dout(n3820));
    jdff dff_A_ArIkvXv60_1(.din(n3826), .dout(n3823));
    jdff dff_A_xODEzUgS7_1(.din(n3829), .dout(n3826));
    jdff dff_A_gQitHaxw7_1(.din(n3832), .dout(n3829));
    jdff dff_A_fwjkoGRV6_1(.din(G261gat), .dout(n3832));
    jdff dff_A_bSvZyBQD0_0(.din(n514), .dout(n3835));
    jdff dff_A_WmCX4QAd4_1(.din(n350), .dout(n3838));
    jdff dff_A_Ozb6AsFn9_0(.din(n3844), .dout(n3841));
    jdff dff_A_BZzvcps99_0(.din(n3847), .dout(n3844));
    jdff dff_A_NmSiOZAZ2_0(.din(n3850), .dout(n3847));
    jdff dff_A_9Q1Z28lf8_0(.din(n3853), .dout(n3850));
    jdff dff_A_WeingIaf9_0(.din(G126gat), .dout(n3853));
    jdff dff_A_GWKmMSds5_1(.din(n3859), .dout(n3856));
    jdff dff_A_MZNSBQMW6_1(.din(n3862), .dout(n3859));
    jdff dff_A_dHCIQLS56_1(.din(n3865), .dout(n3862));
    jdff dff_A_CqfVyh1X8_1(.din(n3868), .dout(n3865));
    jdff dff_A_ZoFaf9jF1_1(.din(n3871), .dout(n3868));
    jdff dff_A_faiL1H6P0_1(.din(n3874), .dout(n3871));
    jdff dff_A_nbBr9Jmr4_1(.din(n3877), .dout(n3874));
    jdff dff_A_KCKcfahM1_1(.din(G201gat), .dout(n3877));
    jdff dff_A_fqYz0gn91_2(.din(n3883), .dout(n3880));
    jdff dff_A_KkK22m7r8_2(.din(n3886), .dout(n3883));
    jdff dff_A_WyfH7fgS7_2(.din(n3889), .dout(n3886));
    jdff dff_A_bt1n3pah3_2(.din(G201gat), .dout(n3889));
    jdff dff_A_nNciEC3p7_2(.din(n3895), .dout(n3892));
    jdff dff_A_Q4679qAd0_2(.din(n3898), .dout(n3895));
    jdff dff_A_f9bvKH217_2(.din(n3901), .dout(n3898));
    jdff dff_A_I0eyeOdC1_2(.din(n3904), .dout(n3901));
    jdff dff_A_V0DLYVtI8_2(.din(n3907), .dout(n3904));
    jdff dff_A_AWcbRMiQ4_2(.din(n3910), .dout(n3907));
    jdff dff_A_zpr6cEBJ4_2(.din(n3913), .dout(n3910));
    jdff dff_A_QZg04gcl8_2(.din(G201gat), .dout(n3913));
    jdff dff_A_7PhRkVid1_1(.din(n3919), .dout(n3916));
    jdff dff_A_dr9yFtro2_1(.din(n3922), .dout(n3919));
    jdff dff_A_eXq9rgTs1_1(.din(n3925), .dout(n3922));
    jdff dff_A_yqcEP5M88_1(.din(n930), .dout(n3925));
    jdff dff_A_d6UTlw6b8_1(.din(n3931), .dout(n3928));
    jdff dff_A_t1XsacIZ5_1(.din(n3934), .dout(n3931));
    jdff dff_A_VUDk8WcB1_1(.din(n3937), .dout(n3934));
    jdff dff_A_gKAnkFhG8_1(.din(n3940), .dout(n3937));
    jdff dff_A_YWGPJBXF6_1(.din(n926), .dout(n3940));
    jdff dff_B_DGX4PC4T2_1(.din(n491), .dout(n3944));
    jdff dff_A_HVyJZuJi9_1(.din(n3949), .dout(n3946));
    jdff dff_A_iAL4fUL74_1(.din(n3952), .dout(n3949));
    jdff dff_A_VWf8y2e67_1(.din(n3955), .dout(n3952));
    jdff dff_A_7RlY8bLN9_1(.din(n3958), .dout(n3955));
    jdff dff_A_uIjmtxar9_1(.din(G111gat), .dout(n3958));
    jdff dff_A_tfwqjyyU3_1(.din(n3964), .dout(n3961));
    jdff dff_A_EftGHX5V2_1(.din(n392), .dout(n3964));
    jdff dff_A_8oI9TO9J2_2(.din(n3970), .dout(n3967));
    jdff dff_A_vUIuLwci3_2(.din(n392), .dout(n3970));
    jdff dff_A_ddvr60bq8_1(.din(n3976), .dout(n3973));
    jdff dff_A_rKyPGpVz7_1(.din(n392), .dout(n3976));
    jdff dff_A_QlSQTq4C2_2(.din(n3982), .dout(n3979));
    jdff dff_A_w9FWJmsQ3_2(.din(n392), .dout(n3982));
    jdff dff_B_8kWAgWBF9_0(.din(n388), .dout(n3986));
    jdff dff_A_wI6DRQ022_0(.din(n3991), .dout(n3988));
    jdff dff_A_jds7d27L4_0(.din(n3994), .dout(n3991));
    jdff dff_A_Wzfu0KCD4_0(.din(n127), .dout(n3994));
    jdff dff_A_XR9CSE6t7_1(.din(n4010), .dout(n3997));
    jdff dff_B_XOaP6XDE5_2(.din(G143gat), .dout(n4001));
    jdff dff_B_ttmPs0EQ7_2(.din(n4001), .dout(n4004));
    jdff dff_B_zp4lH0lP0_2(.din(n4004), .dout(n4007));
    jdff dff_B_SKyVliyN8_2(.din(n4007), .dout(n4010));
    jdff dff_A_1W0H5qBI4_0(.din(n4015), .dout(n4012));
    jdff dff_A_wSAYqYIq6_0(.din(n4018), .dout(n4015));
    jdff dff_A_KTxNf5Mh6_0(.din(n4021), .dout(n4018));
    jdff dff_A_PomoBPfT4_0(.din(n4024), .dout(n4021));
    jdff dff_A_jMBcLWEX5_0(.din(n4027), .dout(n4024));
    jdff dff_A_ClVOk8HB2_0(.din(n4030), .dout(n4027));
    jdff dff_A_UztsRuXl7_0(.din(n4033), .dout(n4030));
    jdff dff_A_vSNtDbIa9_0(.din(G183gat), .dout(n4033));
    jdff dff_A_jXmvuQg96_1(.din(n4039), .dout(n4036));
    jdff dff_A_pWHCK0eD6_1(.din(n4042), .dout(n4039));
    jdff dff_A_RE7WW2799_1(.din(n4045), .dout(n4042));
    jdff dff_A_M3JOp4nt7_1(.din(G183gat), .dout(n4045));
    jdff dff_A_MAXA9IyN0_2(.din(n4051), .dout(n4048));
    jdff dff_A_bCaJ9rnB5_2(.din(n4054), .dout(n4051));
    jdff dff_A_iyvIJL261_2(.din(n4057), .dout(n4054));
    jdff dff_A_jKmKaN8m1_2(.din(n4060), .dout(n4057));
    jdff dff_A_i0ZiWJD53_2(.din(n4063), .dout(n4060));
    jdff dff_A_wjUNbkYd0_2(.din(n4066), .dout(n4063));
    jdff dff_A_NrRqS20P0_2(.din(n4069), .dout(n4066));
    jdff dff_A_bESZbtfo6_2(.din(G183gat), .dout(n4069));
    jdff dff_A_mO5uSkrM3_0(.din(n4075), .dout(n4072));
    jdff dff_A_ZBKepXBW4_0(.din(n4078), .dout(n4075));
    jdff dff_A_iYAmN6LJ7_0(.din(n4081), .dout(n4078));
    jdff dff_A_yaXvQ9sw2_0(.din(n4084), .dout(n4081));
    jdff dff_A_hM2aoxTy5_0(.din(n4087), .dout(n4084));
    jdff dff_A_K8RBRrLP4_0(.din(n4090), .dout(n4087));
    jdff dff_A_PBBSU47T0_0(.din(n4093), .dout(n4090));
    jdff dff_A_AQyWoWVP1_0(.din(n1055), .dout(n4093));
    jdff dff_B_Ts3otrzS6_0(.din(n1015), .dout(n4097));
    jdff dff_B_6AipjvpJ7_0(.din(n4097), .dout(n4100));
    jdff dff_B_p6SyBldd6_0(.din(n4100), .dout(n4103));
    jdff dff_A_QTP6IFPs4_0(.din(n4108), .dout(n4105));
    jdff dff_A_d8ZqSQZm5_0(.din(n4111), .dout(n4108));
    jdff dff_A_wMZJN35v9_0(.din(n4114), .dout(n4111));
    jdff dff_A_X6eRaYX78_0(.din(G153gat), .dout(n4114));
    jdff dff_A_HEsdDwwn8_2(.din(n4120), .dout(n4117));
    jdff dff_A_Jw8bTo2j2_2(.din(n4123), .dout(n4120));
    jdff dff_A_6pFHfPs42_2(.din(n4126), .dout(n4123));
    jdff dff_A_SVAwRhBm6_2(.din(n4129), .dout(n4126));
    jdff dff_A_qQHNDwii7_2(.din(G153gat), .dout(n4129));
    jdff dff_A_yWMPujIT7_0(.din(n4135), .dout(n4132));
    jdff dff_A_AGG8RYi54_0(.din(n4138), .dout(n4135));
    jdff dff_A_ajWd8BSR1_0(.din(n4141), .dout(n4138));
    jdff dff_A_NUAbXkWe9_0(.din(n4144), .dout(n4141));
    jdff dff_A_7M8ANXzy7_0(.din(G106gat), .dout(n4144));
    jdff dff_A_yD0VGvYK8_1(.din(n4150), .dout(n4147));
    jdff dff_A_FgeEyTeZ8_1(.din(n4153), .dout(n4150));
    jdff dff_A_1tBzBOUQ3_1(.din(n4156), .dout(n4153));
    jdff dff_A_j2xZuIC02_1(.din(n4159), .dout(n4156));
    jdff dff_A_yeHP93kZ5_1(.din(n4162), .dout(n4159));
    jdff dff_A_x3c0XfEU5_1(.din(n4165), .dout(n4162));
    jdff dff_A_m4k7EtwD6_1(.din(G177gat), .dout(n4165));
    jdff dff_A_BdwHBUHD2_2(.din(n4171), .dout(n4168));
    jdff dff_A_KMn96lEg1_2(.din(n4174), .dout(n4171));
    jdff dff_A_CY8P0kfJ7_2(.din(n4177), .dout(n4174));
    jdff dff_A_WSKquXtZ5_2(.din(n4180), .dout(n4177));
    jdff dff_A_nNQ9DpNP8_2(.din(n4183), .dout(n4180));
    jdff dff_A_MTZAPu169_2(.din(n4186), .dout(n4183));
    jdff dff_A_szDrL2Wm8_2(.din(G177gat), .dout(n4186));
    jdff dff_A_Z1jsBvNe5_2(.din(n4192), .dout(n4189));
    jdff dff_A_KmZYAzur6_2(.din(n4195), .dout(n4192));
    jdff dff_A_cHBGzICT0_2(.din(n4198), .dout(n4195));
    jdff dff_A_rP3rK1Vr4_2(.din(G177gat), .dout(n4198));
    jdff dff_A_ECHHZQPu9_1(.din(n4204), .dout(n4201));
    jdff dff_A_XoYtyOy69_1(.din(n4207), .dout(n4204));
    jdff dff_A_a07NDFPc2_1(.din(n4210), .dout(n4207));
    jdff dff_A_FH4QgV1M8_1(.din(n4213), .dout(n4210));
    jdff dff_A_cM7tMsys0_1(.din(n4216), .dout(n4213));
    jdff dff_A_jvyYKYyr3_1(.din(n4219), .dout(n4216));
    jdff dff_A_qjnqF0wv6_1(.din(n4222), .dout(n4219));
    jdff dff_A_XaSQRJzn9_1(.din(n4225), .dout(n4222));
    jdff dff_A_t8uQFiOZ9_1(.din(n1326), .dout(n4225));
    jdff dff_B_zM4IdtOI4_0(.din(n987), .dout(n4229));
    jdff dff_B_vUYxz9TH0_0(.din(n4229), .dout(n4232));
    jdff dff_B_yNPXiZOq1_0(.din(n4232), .dout(n4235));
    jdff dff_B_b3prPnl21_0(.din(n898), .dout(n4238));
    jdff dff_A_LRt7OTZo0_0(.din(G17gat), .dout(n4240));
    jdff dff_A_DFPhiLNs1_2(.din(n4246), .dout(n4243));
    jdff dff_A_yRtBaMq77_2(.din(n4249), .dout(n4246));
    jdff dff_A_v4FSawgS7_2(.din(G17gat), .dout(n4249));
    jdff dff_A_nlkU6uhQ0_0(.din(G80gat), .dout(n4252));
    jdff dff_A_A9E8vdJ38_2(.din(G80gat), .dout(n4255));
    jdff dff_A_RDYRiz6I3_0(.din(n4261), .dout(n4258));
    jdff dff_A_bibeQP7Q3_0(.din(n4264), .dout(n4261));
    jdff dff_A_49kWzJ3N9_0(.din(G55gat), .dout(n4264));
    jdff dff_A_vRztP4pg7_1(.din(G55gat), .dout(n4267));
    jdff dff_A_QhYn5t4m1_1(.din(n4283), .dout(n4270));
    jdff dff_B_zvOTUrU43_2(.din(G149gat), .dout(n4274));
    jdff dff_B_Zt7zWCQB8_2(.din(n4274), .dout(n4277));
    jdff dff_B_pL2mCnru0_2(.din(n4277), .dout(n4280));
    jdff dff_B_ds0xvXlA6_2(.din(n4280), .dout(n4283));
    jdff dff_B_ZRw0s8gv8_0(.din(n342), .dout(n4286));
    jdff dff_A_jbDHMsX74_0(.din(n4291), .dout(n4288));
    jdff dff_A_WXECFDTI9_0(.din(n330), .dout(n4291));
    jdff dff_B_7pT4tBQP9_0(.din(n322), .dout(n4295));
    jdff dff_A_8DmXtU3j6_1(.din(G51gat), .dout(n4297));
    jdff dff_A_iI9RsNaw6_1(.din(n4303), .dout(n4300));
    jdff dff_A_HavkOJJE6_1(.din(n4306), .dout(n4303));
    jdff dff_A_bywnkVAZ2_1(.din(n4309), .dout(n4306));
    jdff dff_A_i8iMz5ip7_1(.din(n4312), .dout(n4309));
    jdff dff_A_3vyI5rie3_1(.din(G1gat), .dout(n4312));
    jdff dff_A_JzK7kycc4_1(.din(G42gat), .dout(n4315));
    jdff dff_A_qtEIuVFu9_1(.din(G42gat), .dout(n4318));
    jdff dff_A_EDqdme8J4_1(.din(n4324), .dout(n4321));
    jdff dff_A_oOBWseRU9_1(.din(n4327), .dout(n4324));
    jdff dff_A_be5oHboV7_1(.din(n4330), .dout(n4327));
    jdff dff_A_YZrrfRrS1_1(.din(n4333), .dout(n4330));
    jdff dff_A_nayQiYXK3_1(.din(G101gat), .dout(n4333));
    jdff dff_A_9tSlHmkX2_1(.din(n4339), .dout(n4336));
    jdff dff_A_0OEzxPyU6_1(.din(n4342), .dout(n4339));
    jdff dff_A_Jr6sG1Ph8_1(.din(n4345), .dout(n4342));
    jdff dff_A_izl34Adi5_1(.din(n4348), .dout(n4345));
    jdff dff_A_RHfp2CIP1_1(.din(n4351), .dout(n4348));
    jdff dff_A_ryF2tkFQ7_1(.din(n4354), .dout(n4351));
    jdff dff_A_qRKbhJJt7_1(.din(G171gat), .dout(n4354));
    jdff dff_A_1E524EgH1_2(.din(n4360), .dout(n4357));
    jdff dff_A_5DUnFiR40_2(.din(n4363), .dout(n4360));
    jdff dff_A_GkJHd3ou9_2(.din(n4366), .dout(n4363));
    jdff dff_A_zIU79f7v9_2(.din(n4369), .dout(n4366));
    jdff dff_A_AwXPWF3r1_2(.din(n4372), .dout(n4369));
    jdff dff_A_moQLh0bi9_2(.din(n4375), .dout(n4372));
    jdff dff_A_zDzKJnBE0_2(.din(G171gat), .dout(n4375));
    jdff dff_A_wkhht0JW4_2(.din(n4381), .dout(n4378));
    jdff dff_A_zjRwJyqb7_2(.din(n4384), .dout(n4381));
    jdff dff_A_jtDD79jW1_2(.din(n4387), .dout(n4384));
    jdff dff_A_sBkbIeom1_2(.din(G171gat), .dout(n4387));
    jdff dff_A_X0kHbAdb7_2(.din(n93), .dout(n4390));
    jdff dff_A_GuAOCVhn2_0(.din(n4390), .dout(n4393));
    jdff dff_A_LKlLEh6J0_0(.din(n4393), .dout(n4396));
    jdff dff_A_QY1HNHBJ4_0(.din(n4396), .dout(n4399));
    jdff dff_A_aW2Db9OB6_0(.din(n4399), .dout(n4402));
    jdff dff_A_ppDEx3IG8_0(.din(n4402), .dout(n4405));
    jdff dff_A_hBXJmn1q4_0(.din(n4405), .dout(n4408));
    jdff dff_A_FcZzibNF5_0(.din(n4408), .dout(n4411));
    jdff dff_A_RjGobxKk6_0(.din(n4411), .dout(n4414));
    jdff dff_A_KLsQ9dIp4_0(.din(n4414), .dout(n4417));
    jdff dff_A_RvwfMsgN3_0(.din(n4417), .dout(n4420));
    jdff dff_A_7tU4sIsA9_0(.din(n4420), .dout(n4423));
    jdff dff_A_aZ6oFDTS2_0(.din(n4423), .dout(n4426));
    jdff dff_A_jrV05aOS6_0(.din(n4426), .dout(n4429));
    jdff dff_A_6q7s0qdu3_0(.din(n4429), .dout(n4432));
    jdff dff_A_nkt1lD8z7_0(.din(n4432), .dout(n4435));
    jdff dff_A_eNFRzgiG5_0(.din(n4435), .dout(n4438));
    jdff dff_A_ITEFn8wP3_0(.din(n4438), .dout(n4441));
    jdff dff_A_7i9jumX77_0(.din(n4441), .dout(G388gat));
    jdff dff_A_Y1nK9cE15_2(.din(n101), .dout(n4447));
    jdff dff_A_pxVP3Bml5_0(.din(n4447), .dout(n4450));
    jdff dff_A_uS7IE3Xd3_0(.din(n4450), .dout(n4453));
    jdff dff_A_xBieCWyF6_0(.din(n4453), .dout(n4456));
    jdff dff_A_vZnXxdw23_0(.din(n4456), .dout(n4459));
    jdff dff_A_DhjSzHIZ5_0(.din(n4459), .dout(n4462));
    jdff dff_A_q8JscRw53_0(.din(n4462), .dout(n4465));
    jdff dff_A_HT3gbkfU4_0(.din(n4465), .dout(n4468));
    jdff dff_A_qXGm286t0_0(.din(n4468), .dout(n4471));
    jdff dff_A_jO4U8LkB2_0(.din(n4471), .dout(n4474));
    jdff dff_A_HIBjT0qA1_0(.din(n4474), .dout(n4477));
    jdff dff_A_BtI0d3MF4_0(.din(n4477), .dout(n4480));
    jdff dff_A_S9KIXEaX7_0(.din(n4480), .dout(n4483));
    jdff dff_A_rlDvStwN0_0(.din(n4483), .dout(n4486));
    jdff dff_A_vUSHjRba9_0(.din(n4486), .dout(n4489));
    jdff dff_A_XySDXnhr5_0(.din(n4489), .dout(n4492));
    jdff dff_A_rchMZ7zR7_0(.din(n4492), .dout(n4495));
    jdff dff_A_52z0K9tC3_0(.din(n4495), .dout(n4498));
    jdff dff_A_8dNA4qOz6_0(.din(n4498), .dout(G389gat));
    jdff dff_A_ZXpPQbxW2_2(.din(n105), .dout(n4504));
    jdff dff_A_OTiqX9dw5_0(.din(n4504), .dout(n4507));
    jdff dff_A_pTDW5cen9_0(.din(n4507), .dout(n4510));
    jdff dff_A_zhlrvFaz9_0(.din(n4510), .dout(n4513));
    jdff dff_A_EKQQIoI42_0(.din(n4513), .dout(n4516));
    jdff dff_A_p3CTsA2X3_0(.din(n4516), .dout(n4519));
    jdff dff_A_0tBTn4xp7_0(.din(n4519), .dout(n4522));
    jdff dff_A_x4uE6wDa7_0(.din(n4522), .dout(n4525));
    jdff dff_A_188jnfxY0_0(.din(n4525), .dout(n4528));
    jdff dff_A_vfiaz7JC2_0(.din(n4528), .dout(n4531));
    jdff dff_A_0QEDlCjd3_0(.din(n4531), .dout(n4534));
    jdff dff_A_2CcnYQGP6_0(.din(n4534), .dout(n4537));
    jdff dff_A_M45ZyP6K8_0(.din(n4537), .dout(n4540));
    jdff dff_A_jy5KxXSS5_0(.din(n4540), .dout(n4543));
    jdff dff_A_AkCJCekU5_0(.din(n4543), .dout(n4546));
    jdff dff_A_vhmXD8te8_0(.din(n4546), .dout(n4549));
    jdff dff_A_5ntqW6Wo7_0(.din(n4549), .dout(n4552));
    jdff dff_A_f6hGMEQq3_0(.din(n4552), .dout(n4555));
    jdff dff_A_cJAURovK3_0(.din(n4555), .dout(G390gat));
    jdff dff_A_SpizB91N3_2(.din(n109), .dout(n4561));
    jdff dff_A_wFiDbO0J6_0(.din(n4561), .dout(n4564));
    jdff dff_A_k1Y13Y8V4_0(.din(n4564), .dout(n4567));
    jdff dff_A_b1VoSuUE0_0(.din(n4567), .dout(n4570));
    jdff dff_A_vWAO6IYk0_0(.din(n4570), .dout(n4573));
    jdff dff_A_1A2nlKG22_0(.din(n4573), .dout(n4576));
    jdff dff_A_IicdvabJ4_0(.din(n4576), .dout(n4579));
    jdff dff_A_I8ekCjS71_0(.din(n4579), .dout(n4582));
    jdff dff_A_peuVB3pl6_0(.din(n4582), .dout(n4585));
    jdff dff_A_UlI71KH61_0(.din(n4585), .dout(n4588));
    jdff dff_A_vauKkLvB3_0(.din(n4588), .dout(n4591));
    jdff dff_A_gZPnn3N70_0(.din(n4591), .dout(n4594));
    jdff dff_A_RmHT7Dty3_0(.din(n4594), .dout(n4597));
    jdff dff_A_zUP43K6b4_0(.din(n4597), .dout(n4600));
    jdff dff_A_7iflffAH3_0(.din(n4600), .dout(n4603));
    jdff dff_A_7qbnZ8U06_0(.din(n4603), .dout(n4606));
    jdff dff_A_8Soj1kAF1_0(.din(n4606), .dout(n4609));
    jdff dff_A_IZgVQmPA7_0(.din(n4609), .dout(n4612));
    jdff dff_A_jAQp9lAk2_0(.din(n4612), .dout(n4615));
    jdff dff_A_DTCDeFvN1_0(.din(n4615), .dout(G391gat));
    jdff dff_A_DaA0Cm0b8_2(.din(n121), .dout(n4621));
    jdff dff_A_kcvgynvC2_0(.din(n4621), .dout(n4624));
    jdff dff_A_pVzYYPWE4_0(.din(n4624), .dout(n4627));
    jdff dff_A_udigj5878_0(.din(n4627), .dout(n4630));
    jdff dff_A_AmwrHkzk7_0(.din(n4630), .dout(n4633));
    jdff dff_A_CpqIqHEB8_0(.din(n4633), .dout(n4636));
    jdff dff_A_gOD43Cmg6_0(.din(n4636), .dout(n4639));
    jdff dff_A_THoY87Un0_0(.din(n4639), .dout(n4642));
    jdff dff_A_kxVaw1Yf9_0(.din(n4642), .dout(n4645));
    jdff dff_A_X58358Id2_0(.din(n4645), .dout(n4648));
    jdff dff_A_321Hbrh97_0(.din(n4648), .dout(n4651));
    jdff dff_A_GVXUdRe55_0(.din(n4651), .dout(n4654));
    jdff dff_A_VCRxQNCe3_0(.din(n4654), .dout(n4657));
    jdff dff_A_Vtr8G3At1_0(.din(n4657), .dout(n4660));
    jdff dff_A_b8SS2enS3_0(.din(n4660), .dout(n4663));
    jdff dff_A_r9khn0Sj8_0(.din(n4663), .dout(n4666));
    jdff dff_A_kK4gBzNY9_0(.din(n4666), .dout(n4669));
    jdff dff_A_gm97eV5i6_0(.din(n4669), .dout(n4672));
    jdff dff_A_076S63OU4_0(.din(n4672), .dout(G418gat));
    jdff dff_A_Q7Y9z1ZK3_2(.din(n142), .dout(n4678));
    jdff dff_A_HzPxqt1Z6_0(.din(n4678), .dout(n4681));
    jdff dff_A_U6M9yE166_0(.din(n4681), .dout(n4684));
    jdff dff_A_YNdaR6bh9_0(.din(n4684), .dout(n4687));
    jdff dff_A_9Cy8yFQN2_0(.din(n4687), .dout(n4690));
    jdff dff_A_dQvVwmBJ9_0(.din(n4690), .dout(n4693));
    jdff dff_A_K9H0oYzO8_0(.din(n4693), .dout(n4696));
    jdff dff_A_XeIn005r7_0(.din(n4696), .dout(n4699));
    jdff dff_A_HRA0lOJY5_0(.din(n4699), .dout(n4702));
    jdff dff_A_ZnsDw7zE3_0(.din(n4702), .dout(n4705));
    jdff dff_A_HVRVC1VK8_0(.din(n4705), .dout(n4708));
    jdff dff_A_geW4UDfo4_0(.din(n4708), .dout(n4711));
    jdff dff_A_BKRIBCOx6_0(.din(n4711), .dout(n4714));
    jdff dff_A_7Tn18E0L6_0(.din(n4714), .dout(n4717));
    jdff dff_A_kHreSdkd2_0(.din(n4717), .dout(n4720));
    jdff dff_A_lkLcpaEg1_0(.din(n4720), .dout(n4723));
    jdff dff_A_uwCUJgbf2_0(.din(n4723), .dout(G419gat));
    jdff dff_A_PC6qmYf30_2(.din(n156), .dout(n4729));
    jdff dff_A_0FdV3wTW3_0(.din(n4729), .dout(n4732));
    jdff dff_A_Z8nbjcKD3_0(.din(n4732), .dout(n4735));
    jdff dff_A_z6pwVCWP5_0(.din(n4735), .dout(n4738));
    jdff dff_A_2ZC5W0XD0_0(.din(n4738), .dout(n4741));
    jdff dff_A_pDR1iKwO0_0(.din(n4741), .dout(n4744));
    jdff dff_A_uxUs2PCY8_0(.din(n4744), .dout(n4747));
    jdff dff_A_8I4fbpua4_0(.din(n4747), .dout(n4750));
    jdff dff_A_aTCXI97f2_0(.din(n4750), .dout(n4753));
    jdff dff_A_CR55BGBM5_0(.din(n4753), .dout(n4756));
    jdff dff_A_jSRamrSx0_0(.din(n4756), .dout(n4759));
    jdff dff_A_9hCgF8fD4_0(.din(n4759), .dout(n4762));
    jdff dff_A_qML2Jkjc9_0(.din(n4762), .dout(n4765));
    jdff dff_A_TCjHZf5d7_0(.din(n4765), .dout(n4768));
    jdff dff_A_kanGzhW38_0(.din(n4768), .dout(n4771));
    jdff dff_A_GEWHvxaL8_0(.din(n4771), .dout(n4774));
    jdff dff_A_52Fa1Yns7_0(.din(n4774), .dout(n4777));
    jdff dff_A_rLmSjeJg4_0(.din(n4777), .dout(G420gat));
    jdff dff_A_KVpRZNKx4_2(.din(n170), .dout(n4783));
    jdff dff_A_Rhynn9945_0(.din(n4783), .dout(n4786));
    jdff dff_A_wigCtVz05_0(.din(n4786), .dout(n4789));
    jdff dff_A_YKYRJEAY4_0(.din(n4789), .dout(n4792));
    jdff dff_A_RYjya74O8_0(.din(n4792), .dout(n4795));
    jdff dff_A_1caixoAE3_0(.din(n4795), .dout(n4798));
    jdff dff_A_gDP94gmv7_0(.din(n4798), .dout(n4801));
    jdff dff_A_rgVVfYiv7_0(.din(n4801), .dout(n4804));
    jdff dff_A_d2BtERMW8_0(.din(n4804), .dout(n4807));
    jdff dff_A_l7NK7DFj6_0(.din(n4807), .dout(n4810));
    jdff dff_A_iMxUOqYy0_0(.din(n4810), .dout(n4813));
    jdff dff_A_Ocz9z1wh1_0(.din(n4813), .dout(n4816));
    jdff dff_A_zj7HAygN9_0(.din(n4816), .dout(n4819));
    jdff dff_A_JBKPhhKh7_0(.din(n4819), .dout(n4822));
    jdff dff_A_jEc1bim20_0(.din(n4822), .dout(n4825));
    jdff dff_A_BFp5owVO5_0(.din(n4825), .dout(n4828));
    jdff dff_A_QNVKxMMM6_0(.din(n4828), .dout(n4831));
    jdff dff_A_yg0VlKrA6_0(.din(n4831), .dout(G421gat));
    jdff dff_A_e8sPWf7F8_2(.din(n177), .dout(n4837));
    jdff dff_A_SI057U6r4_0(.din(n4837), .dout(n4840));
    jdff dff_A_nA3S8Bqt0_0(.din(n4840), .dout(n4843));
    jdff dff_A_qdFba6oH0_0(.din(n4843), .dout(n4846));
    jdff dff_A_0kFxVnYG9_0(.din(n4846), .dout(n4849));
    jdff dff_A_dePyAu5j6_0(.din(n4849), .dout(n4852));
    jdff dff_A_0jL7wY0t2_0(.din(n4852), .dout(n4855));
    jdff dff_A_WDyrjHUh8_0(.din(n4855), .dout(n4858));
    jdff dff_A_HQy7LTtE8_0(.din(n4858), .dout(n4861));
    jdff dff_A_drtiOR7H3_0(.din(n4861), .dout(n4864));
    jdff dff_A_okes5AJ46_0(.din(n4864), .dout(n4867));
    jdff dff_A_OLSXyivU0_0(.din(n4867), .dout(n4870));
    jdff dff_A_zBpAOFK81_0(.din(n4870), .dout(n4873));
    jdff dff_A_xHrPpOCF5_0(.din(n4873), .dout(n4876));
    jdff dff_A_mPN3NODv5_0(.din(n4876), .dout(n4879));
endmodule

