/*

c432:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jdff: 1153
	jand: 111
	jor: 110

Summary:
	jxor: 3
	jspl: 93
	jspl3: 51
	jnot: 50
	jdff: 1153
	jand: 111
	jor: 110
*/

module c432(gclk, G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat);
	input gclk;
	input G1gat;
	input G4gat;
	input G8gat;
	input G11gat;
	input G14gat;
	input G17gat;
	input G21gat;
	input G24gat;
	input G27gat;
	input G30gat;
	input G34gat;
	input G37gat;
	input G40gat;
	input G43gat;
	input G47gat;
	input G50gat;
	input G53gat;
	input G56gat;
	input G60gat;
	input G63gat;
	input G66gat;
	input G69gat;
	input G73gat;
	input G76gat;
	input G79gat;
	input G82gat;
	input G86gat;
	input G89gat;
	input G92gat;
	input G95gat;
	input G99gat;
	input G102gat;
	input G105gat;
	input G108gat;
	input G112gat;
	input G115gat;
	output G223gat;
	output G329gat;
	output G370gat;
	output G421gat;
	output G430gat;
	output G431gat;
	output G432gat;
	wire n43;
	wire n44;
	wire n45;
	wire n46;
	wire n47;
	wire n48;
	wire n49;
	wire n50;
	wire n51;
	wire n52;
	wire n53;
	wire n54;
	wire n55;
	wire n56;
	wire n57;
	wire n58;
	wire n59;
	wire n60;
	wire n61;
	wire n62;
	wire n63;
	wire n64;
	wire n65;
	wire n66;
	wire n67;
	wire n69;
	wire n70;
	wire n71;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n150;
	wire n151;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n182;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n191;
	wire n192;
	wire n193;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n217;
	wire n218;
	wire n219;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n235;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n244;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n262;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G4gat_0;
	wire [2:0] w_G8gat_0;
	wire [2:0] w_G11gat_0;
	wire [2:0] w_G14gat_0;
	wire [2:0] w_G17gat_0;
	wire [2:0] w_G21gat_0;
	wire [1:0] w_G21gat_1;
	wire [1:0] w_G24gat_0;
	wire [1:0] w_G27gat_0;
	wire [1:0] w_G30gat_0;
	wire [2:0] w_G34gat_0;
	wire [2:0] w_G37gat_0;
	wire [1:0] w_G40gat_0;
	wire [2:0] w_G43gat_0;
	wire [1:0] w_G43gat_1;
	wire [1:0] w_G47gat_0;
	wire [2:0] w_G50gat_0;
	wire [1:0] w_G53gat_0;
	wire [2:0] w_G56gat_0;
	wire [2:0] w_G60gat_0;
	wire [2:0] w_G63gat_0;
	wire [1:0] w_G66gat_0;
	wire [2:0] w_G69gat_0;
	wire [2:0] w_G73gat_0;
	wire [1:0] w_G76gat_0;
	wire [1:0] w_G79gat_0;
	wire [2:0] w_G82gat_0;
	wire [2:0] w_G86gat_0;
	wire [1:0] w_G86gat_1;
	wire [2:0] w_G89gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G95gat_0;
	wire [2:0] w_G99gat_0;
	wire [2:0] w_G102gat_0;
	wire [1:0] w_G105gat_0;
	wire [2:0] w_G108gat_0;
	wire [2:0] w_G112gat_0;
	wire [1:0] w_G115gat_0;
	wire [2:0] w_G223gat_0;
	wire [2:0] w_G223gat_1;
	wire [2:0] w_G223gat_2;
	wire [1:0] w_G223gat_3;
	wire G223gat_fa_;
	wire [2:0] w_G329gat_0;
	wire [2:0] w_G329gat_1;
	wire [2:0] w_G329gat_2;
	wire [2:0] w_G329gat_3;
	wire [2:0] w_G329gat_4;
	wire [2:0] w_G329gat_5;
	wire w_G329gat_6;
	wire G329gat_fa_;
	wire [2:0] w_G370gat_0;
	wire [2:0] w_G370gat_1;
	wire w_G370gat_2;
	wire G370gat_fa_;
	wire w_G430gat_0;
	wire G430gat_fa_;
	wire [1:0] w_n43_0;
	wire [1:0] w_n44_0;
	wire [1:0] w_n47_0;
	wire [1:0] w_n52_0;
	wire [1:0] w_n53_0;
	wire [1:0] w_n56_0;
	wire [1:0] w_n58_0;
	wire [1:0] w_n61_0;
	wire [1:0] w_n63_0;
	wire [1:0] w_n69_0;
	wire [1:0] w_n71_0;
	wire [1:0] w_n72_0;
	wire [1:0] w_n73_0;
	wire [1:0] w_n77_0;
	wire [1:0] w_n78_0;
	wire [1:0] w_n79_0;
	wire [1:0] w_n82_0;
	wire [1:0] w_n84_0;
	wire [1:0] w_n87_0;
	wire [1:0] w_n89_0;
	wire [2:0] w_n94_0;
	wire [2:0] w_n94_1;
	wire [2:0] w_n94_2;
	wire [2:0] w_n94_3;
	wire [1:0] w_n94_4;
	wire [1:0] w_n96_0;
	wire [1:0] w_n98_0;
	wire [1:0] w_n100_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n109_0;
	wire [2:0] w_n114_0;
	wire [1:0] w_n115_0;
	wire [1:0] w_n119_0;
	wire [1:0] w_n121_0;
	wire [1:0] w_n123_0;
	wire [2:0] w_n126_0;
	wire [1:0] w_n128_0;
	wire [2:0] w_n130_0;
	wire [1:0] w_n132_0;
	wire [1:0] w_n139_0;
	wire [1:0] w_n141_0;
	wire [1:0] w_n142_0;
	wire [1:0] w_n145_0;
	wire [1:0] w_n146_0;
	wire [1:0] w_n147_0;
	wire [1:0] w_n150_0;
	wire [1:0] w_n151_0;
	wire [1:0] w_n154_0;
	wire [1:0] w_n156_0;
	wire [1:0] w_n159_0;
	wire [1:0] w_n164_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n174_0;
	wire [1:0] w_n177_0;
	wire [2:0] w_n182_0;
	wire [2:0] w_n182_1;
	wire [2:0] w_n182_2;
	wire [1:0] w_n182_3;
	wire [1:0] w_n184_0;
	wire [1:0] w_n188_0;
	wire [1:0] w_n191_0;
	wire [1:0] w_n193_0;
	wire [1:0] w_n197_0;
	wire [1:0] w_n198_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n205_0;
	wire [1:0] w_n217_0;
	wire [1:0] w_n219_0;
	wire [1:0] w_n222_0;
	wire [1:0] w_n224_0;
	wire [1:0] w_n231_0;
	wire [1:0] w_n254_0;
	wire [1:0] w_n260_0;
	wire [2:0] w_n271_0;
	wire [2:0] w_n271_1;
	wire [2:0] w_n271_2;
	wire [1:0] w_n271_3;
	wire [1:0] w_n274_0;
	wire [1:0] w_n281_0;
	wire [1:0] w_n283_0;
	wire [1:0] w_n286_0;
	wire [1:0] w_n290_0;
	wire [1:0] w_n293_0;
	wire [1:0] w_n296_0;
	wire [1:0] w_n303_0;
	wire [1:0] w_n305_0;
	wire [1:0] w_n313_0;
	wire [1:0] w_n314_0;
	wire [2:0] w_n317_0;
	wire [1:0] w_n319_0;
	wire w_dff_B_GSnDh2kE5_1;
	wire w_dff_B_hIduJqmc9_1;
	wire w_dff_B_VIrjoWqg4_1;
	wire w_dff_B_czkWL5uQ7_0;
	wire w_dff_B_jDyP1OjQ3_0;
	wire w_dff_B_ariQ0ZvI5_0;
	wire w_dff_B_CyL4EsOq2_0;
	wire w_dff_B_9zOLbmIy1_0;
	wire w_dff_B_ZYoFFb5A6_1;
	wire w_dff_A_X7vp4PL19_0;
	wire w_dff_B_xLjl8rKw0_0;
	wire w_dff_B_Tx7d7DJC6_0;
	wire w_dff_B_CSQEN4uL9_0;
	wire w_dff_B_O8kTvuKD0_0;
	wire w_dff_B_dVyWw4fQ3_0;
	wire w_dff_A_pLfHtfeN2_0;
	wire w_dff_B_KXmdAilH7_1;
	wire w_dff_B_zDDe9ktI8_0;
	wire w_dff_B_M7M6Hzdg9_0;
	wire w_dff_B_hKUYCX0D1_0;
	wire w_dff_B_KCxFHtaV2_0;
	wire w_dff_B_qxgHqkJt9_0;
	wire w_dff_A_laMmicQ84_0;
	wire w_dff_A_HY9rZFi71_0;
	wire w_dff_A_WFT3tQ0g0_0;
	wire w_dff_A_FmfjjktR9_0;
	wire w_dff_A_y0kxChaU5_0;
	wire w_dff_A_ygXpwAxh3_0;
	wire w_dff_A_WmmXD38Y6_0;
	wire w_dff_B_xHxGJ5Ny8_1;
	wire w_dff_B_oeQS6wIZ6_1;
	wire w_dff_B_NnICCbs74_1;
	wire w_dff_B_7mLxy2vQ7_1;
	wire w_dff_B_kXbpKEBk3_1;
	wire w_dff_B_OAL6iOP00_1;
	wire w_dff_B_WVRZKLQ06_1;
	wire w_dff_B_4lf6p1SM7_1;
	wire w_dff_B_vb4owMNK2_1;
	wire w_dff_B_2gInBCgu9_1;
	wire w_dff_B_CGrQXk1L9_1;
	wire w_dff_B_8vYHROXb7_1;
	wire w_dff_B_D8sSyh4c1_1;
	wire w_dff_B_7xphdRD70_1;
	wire w_dff_B_R88nFhvk8_1;
	wire w_dff_B_F7c70FBE9_1;
	wire w_dff_B_CG7TzqnV4_1;
	wire w_dff_B_TRhcUU752_1;
	wire w_dff_B_BHWgLUzc9_1;
	wire w_dff_B_qAxORBmV6_1;
	wire w_dff_B_bl2fhLvS6_1;
	wire w_dff_B_5D7c1szW3_1;
	wire w_dff_B_6KNdW3L09_1;
	wire w_dff_B_3EXKWv7H2_1;
	wire w_dff_B_BTec5vnc7_1;
	wire w_dff_B_hWCdCurf8_1;
	wire w_dff_B_TihVYKXx0_1;
	wire w_dff_B_lVg0OwBZ2_0;
	wire w_dff_B_mkjwvadh6_0;
	wire w_dff_B_fU6PONy31_0;
	wire w_dff_A_WvE99bJX6_1;
	wire w_dff_A_6186ux1M5_1;
	wire w_dff_A_WFd7z3iY9_1;
	wire w_dff_A_Y6qPYb1y9_1;
	wire w_dff_A_eahucu861_1;
	wire w_dff_A_Dx6iqY3E7_1;
	wire w_dff_B_V16kZFy51_1;
	wire w_dff_B_LPZI1See8_0;
	wire w_dff_B_hcxHYc191_0;
	wire w_dff_B_6eoxg8OF6_0;
	wire w_dff_B_0TbexHT18_0;
	wire w_dff_B_FbCoXbMV1_0;
	wire w_dff_B_LVxx1fIm2_1;
	wire w_dff_B_22sCyIcv4_0;
	wire w_dff_B_ARh6LNE23_0;
	wire w_dff_B_PmwhMaNd7_0;
	wire w_dff_B_4WmcnZt15_0;
	wire w_dff_A_iG3ii5kw4_0;
	wire w_dff_A_LVk07qnr8_0;
	wire w_dff_A_fqjjwXgZ7_0;
	wire w_dff_A_SaJ3X7Bv2_0;
	wire w_dff_A_Hacp7Wwv0_0;
	wire w_dff_A_25w1lPMr9_0;
	wire w_dff_A_VcVnZbwv6_0;
	wire w_dff_A_OAWoaVVb9_0;
	wire w_dff_A_XiFcFEo62_0;
	wire w_dff_A_8TQkw6lt7_0;
	wire w_dff_A_HGwRYJUM1_0;
	wire w_dff_A_OzVYxTJp1_0;
	wire w_dff_A_fnqeUtC94_0;
	wire w_dff_A_F02wDE6p8_0;
	wire w_dff_A_DWFINrfc8_0;
	wire w_dff_A_3xb3bOl61_0;
	wire w_dff_A_tUq7FhWe6_0;
	wire w_dff_A_woeQ6xX11_0;
	wire w_dff_B_VMJWkdGw0_0;
	wire w_dff_B_xwAI8yyP8_0;
	wire w_dff_B_GIKci5Mb3_0;
	wire w_dff_B_feggU7DD0_0;
	wire w_dff_B_YH9V6D4u8_0;
	wire w_dff_B_qkWew6ny7_0;
	wire w_dff_B_ELQB5Iqi7_1;
	wire w_dff_B_GNSqXq4E6_1;
	wire w_dff_B_kIK7VG9F5_1;
	wire w_dff_A_8kvUfK8O1_0;
	wire w_dff_A_3MYg9Swm8_0;
	wire w_dff_A_4dlXNgHr5_0;
	wire w_dff_A_9KT6QPQ52_0;
	wire w_dff_A_UH48UZ7X9_0;
	wire w_dff_A_nnUpAHli6_0;
	wire w_dff_A_yBpJdM7k4_0;
	wire w_dff_A_5bTae3JN6_0;
	wire w_dff_A_5P8rL2ZA6_0;
	wire w_dff_A_O1jOcvJz0_0;
	wire w_dff_A_bbCfdq1r1_0;
	wire w_dff_B_YdMERaM50_2;
	wire w_dff_B_hyyEkbhs8_2;
	wire w_dff_B_IbWdedKo0_2;
	wire w_dff_B_5VLEpwHo0_2;
	wire w_dff_B_pLgYB2pj5_2;
	wire w_dff_B_lOdqvsgp8_2;
	wire w_dff_B_l3RuFBV89_2;
	wire w_dff_B_emhezZSf9_2;
	wire w_dff_B_w3EksEOO7_2;
	wire w_dff_B_893WKOa32_2;
	wire w_dff_B_DTj59Uvb3_2;
	wire w_dff_B_IzSdSrrA8_2;
	wire w_dff_B_wdvUVKDo0_2;
	wire w_dff_B_dh5WGy4B5_2;
	wire w_dff_A_fsA8EV2t2_0;
	wire w_dff_A_xAxsMlXv2_0;
	wire w_dff_A_E53njXCd2_0;
	wire w_dff_A_hmwwARnM2_0;
	wire w_dff_A_oqJHtDKu0_0;
	wire w_dff_A_GNYaiNh17_0;
	wire w_dff_A_Vl5vsEAq2_0;
	wire w_dff_A_ZYa2puiv2_0;
	wire w_dff_A_wX3Rw1q02_0;
	wire w_dff_A_iN0dAAPp8_0;
	wire w_dff_A_KsCL86RT6_0;
	wire w_dff_A_ZUdX4zNb4_0;
	wire w_dff_A_LYF8F3Tq2_0;
	wire w_dff_A_J2Mrws8M5_0;
	wire w_dff_A_wsHHMeLw7_0;
	wire w_dff_A_lYhGSCPn1_1;
	wire w_dff_A_czWZKsfc9_1;
	wire w_dff_A_VSHXhCJc9_1;
	wire w_dff_A_LrTmRjb59_1;
	wire w_dff_A_wjoC0toR2_0;
	wire w_dff_A_vCs445nJ1_0;
	wire w_dff_A_2tlBKJnU7_0;
	wire w_dff_A_AZWId6Kt7_0;
	wire w_dff_A_n8vm7ZZn3_0;
	wire w_dff_A_diPwbLcV5_0;
	wire w_dff_A_BwgELZkZ3_0;
	wire w_dff_A_7m5WlaoD7_0;
	wire w_dff_A_OxYC5Mqn7_0;
	wire w_dff_A_DpZ2unM60_0;
	wire w_dff_A_dtfYF0RU7_0;
	wire w_dff_B_jd4f72az7_2;
	wire w_dff_B_EIZ92mA41_2;
	wire w_dff_B_l7kZjTXc2_2;
	wire w_dff_B_GZupzVj27_2;
	wire w_dff_B_RWLohaRm7_2;
	wire w_dff_B_dV5i4kRd6_2;
	wire w_dff_B_K43EhjD71_2;
	wire w_dff_B_0SRp5Z4h3_2;
	wire w_dff_A_URwKWAYp2_0;
	wire w_dff_A_votMDdNu4_0;
	wire w_dff_A_fHso0OEe1_0;
	wire w_dff_A_zjKeFhqd0_0;
	wire w_dff_A_LpluJNeK5_0;
	wire w_dff_A_9Yk93ou95_0;
	wire w_dff_A_KNtLhHRG3_0;
	wire w_dff_A_pOyopasy9_0;
	wire w_dff_A_qyTZFZPK2_0;
	wire w_dff_A_kU381YMW7_0;
	wire w_dff_A_ulUXXly06_0;
	wire w_dff_A_omUMCf9u4_0;
	wire w_dff_A_VDk9UMgz3_0;
	wire w_dff_A_cx0imB703_0;
	wire w_dff_A_ZM9E6xcm8_0;
	wire w_dff_A_npdtz6Jy5_0;
	wire w_dff_A_6lBG8Cnj6_0;
	wire w_dff_A_tcQbky3R5_0;
	wire w_dff_A_kqU2lrcn5_0;
	wire w_dff_A_qj6x9u1f2_0;
	wire w_dff_B_q00PK1XG6_1;
	wire w_dff_B_2XCdmvSp5_1;
	wire w_dff_B_P1ZSg6HP7_1;
	wire w_dff_B_DVirL3oD2_1;
	wire w_dff_B_icyLWSGx8_1;
	wire w_dff_B_pnbZDh8S3_1;
	wire w_dff_B_7Y4ud1yb0_1;
	wire w_dff_B_eooJ9GeX6_1;
	wire w_dff_B_wjniNUKX8_1;
	wire w_dff_B_9jjsctm77_1;
	wire w_dff_B_ctyO2yCT4_1;
	wire w_dff_B_mecfc78R8_1;
	wire w_dff_B_4c3VtT6s0_1;
	wire w_dff_B_QQXSPl696_1;
	wire w_dff_B_lnQyGsTN2_1;
	wire w_dff_B_QhQFr7YL9_1;
	wire w_dff_B_YOMH6s239_1;
	wire w_dff_B_cmgcXGgN4_1;
	wire w_dff_B_Rh90SVv32_1;
	wire w_dff_B_w71gb5y77_1;
	wire w_dff_B_kZagx7jQ8_1;
	wire w_dff_B_KSNTyxvV8_1;
	wire w_dff_B_5NdIs9Ps6_1;
	wire w_dff_B_FQ33IYN68_1;
	wire w_dff_B_RecGgbmW2_1;
	wire w_dff_B_h2WQfTe00_1;
	wire w_dff_A_KooFJ4an7_0;
	wire w_dff_A_5N7W4bjW9_0;
	wire w_dff_A_91kb09bN8_0;
	wire w_dff_A_9zRlLWAA1_0;
	wire w_dff_A_VBn9TSq39_0;
	wire w_dff_A_sAgWO94h0_0;
	wire w_dff_A_LxoOkUmX6_0;
	wire w_dff_A_OHesSGDi1_0;
	wire w_dff_A_IHbETiyJ4_0;
	wire w_dff_A_OwwoBDjW0_0;
	wire w_dff_A_pK24mIv30_0;
	wire w_dff_A_F4WaHt2f5_0;
	wire w_dff_A_azx97wwe4_0;
	wire w_dff_A_3uDSStZo0_0;
	wire w_dff_A_BwZsNusM9_0;
	wire w_dff_A_LQUvEn4p5_1;
	wire w_dff_A_Flwu4zfB4_1;
	wire w_dff_A_1IPTWx4j2_1;
	wire w_dff_A_QUVyFi4h8_1;
	wire w_dff_A_vfLG6VhC8_1;
	wire w_dff_A_0vzcR0Mt6_1;
	wire w_dff_A_Gq0jnUpT2_1;
	wire w_dff_A_FMMIp7qE6_1;
	wire w_dff_A_WeFkpDEY9_1;
	wire w_dff_A_rfHQNtAG0_1;
	wire w_dff_A_o1svPETJ0_1;
	wire w_dff_A_PvHJiViS7_1;
	wire w_dff_A_987klsKH6_1;
	wire w_dff_A_1sdopjId2_1;
	wire w_dff_A_FYEbGyxv4_1;
	wire w_dff_A_G9ueQvwZ2_1;
	wire w_dff_A_BwAiN2Wa3_1;
	wire w_dff_A_kMxDCVIs9_1;
	wire w_dff_A_u8P8Po8w2_1;
	wire w_dff_A_hWRA1A9B9_1;
	wire w_dff_A_LfEhZHl00_0;
	wire w_dff_A_rkwCWqyX9_0;
	wire w_dff_A_Ob0nhDB07_0;
	wire w_dff_A_uhjLAQNN4_0;
	wire w_dff_A_6JNcqD5U0_0;
	wire w_dff_A_AnMNFDxc1_0;
	wire w_dff_B_fOJxWYgY7_2;
	wire w_dff_B_GHIbASPS3_2;
	wire w_dff_B_zc54HsMS0_2;
	wire w_dff_B_tPqFifj69_2;
	wire w_dff_B_Gije76v97_2;
	wire w_dff_B_iWMwpXHh0_2;
	wire w_dff_B_Au4HEF214_2;
	wire w_dff_B_OH6Bf5Fu2_2;
	wire w_dff_B_tpMnQwPb0_2;
	wire w_dff_B_kNuWFeCk3_2;
	wire w_dff_B_wOkYWYKD3_2;
	wire w_dff_B_UIrplxaR9_2;
	wire w_dff_B_5aEeEyyC1_2;
	wire w_dff_A_Tq2maAmm5_0;
	wire w_dff_A_8ikQTadE7_0;
	wire w_dff_A_9IzPf7lX3_0;
	wire w_dff_A_vm3CM9Dw8_0;
	wire w_dff_A_8fxOPCtD5_0;
	wire w_dff_A_6sxMqMEl1_0;
	wire w_dff_A_Wo8TfAuY9_0;
	wire w_dff_A_5Nc2Jxhl3_0;
	wire w_dff_A_1iLwwVWs3_0;
	wire w_dff_A_ZezFM1pL8_0;
	wire w_dff_A_q0wH6vH95_0;
	wire w_dff_A_3ufiBksR7_0;
	wire w_dff_A_hBCqrYvd4_0;
	wire w_dff_A_hJibkNQl2_0;
	wire w_dff_A_YuMJNmG72_0;
	wire w_dff_A_RK2Z40uw0_0;
	wire w_dff_A_88AAHG1I5_0;
	wire w_dff_A_O16qnquD2_0;
	wire w_dff_A_oleWOq7v0_0;
	wire w_dff_A_oHno2wmd6_0;
	wire w_dff_A_Z4wBsNYM7_1;
	wire w_dff_A_36T123zN7_1;
	wire w_dff_A_bYShhjUX9_1;
	wire w_dff_A_JUcWfsqX4_1;
	wire w_dff_A_j6Kppt9l3_1;
	wire w_dff_A_D90zdTLE8_1;
	wire w_dff_A_bHObf2ni8_1;
	wire w_dff_A_OlluYn5z3_1;
	wire w_dff_A_VKrgORKB5_1;
	wire w_dff_A_kuw4pHGu3_1;
	wire w_dff_A_P23sgYsc5_1;
	wire w_dff_A_RdhsWqx99_1;
	wire w_dff_A_05VLVG5v7_1;
	wire w_dff_A_lkCDXcSL2_1;
	wire w_dff_A_pCCO09rF5_0;
	wire w_dff_A_RD0QYzFV6_0;
	wire w_dff_A_pwWVTRRs6_0;
	wire w_dff_A_oRu1ITMv9_0;
	wire w_dff_A_xvnooeX77_0;
	wire w_dff_A_1rCSSxDP9_0;
	wire w_dff_A_s1FhOk1n5_0;
	wire w_dff_A_gheSqkuk8_0;
	wire w_dff_A_hjY6aPR09_0;
	wire w_dff_A_Ul5kchh18_0;
	wire w_dff_A_oTahqyhp2_0;
	wire w_dff_A_rx3r58Z40_0;
	wire w_dff_B_Vf4E7VPh3_2;
	wire w_dff_B_Oc6o3v8z1_2;
	wire w_dff_B_SkNY9oMq8_2;
	wire w_dff_B_mbruSknS9_2;
	wire w_dff_B_8dEEqOn31_2;
	wire w_dff_B_tym5eEYv0_2;
	wire w_dff_B_1lIJKnEV1_2;
	wire w_dff_B_KszUaK690_2;
	wire w_dff_B_BX5srGLX9_2;
	wire w_dff_B_MpiPvr995_2;
	wire w_dff_B_Kz4UMlW19_2;
	wire w_dff_B_7LaVMsGs4_2;
	wire w_dff_B_ENr5jcRP1_2;
	wire w_dff_A_cFr70PcO5_0;
	wire w_dff_A_Ej189avp4_0;
	wire w_dff_A_yICjViVC5_0;
	wire w_dff_A_jItJKpUJ1_0;
	wire w_dff_A_uxhKUSVq1_0;
	wire w_dff_A_LqUj06CV4_0;
	wire w_dff_A_eqSVw9832_0;
	wire w_dff_A_WMeGJ6pz4_0;
	wire w_dff_A_xTkKj4Pd9_0;
	wire w_dff_A_OQ5F2s9m1_0;
	wire w_dff_A_X2JtlG1n2_0;
	wire w_dff_A_jgOcxwZ09_0;
	wire w_dff_A_MS968xZC4_0;
	wire w_dff_A_sHjkFqOj0_0;
	wire w_dff_A_haPGZmqi5_0;
	wire w_dff_A_idn5NWLt4_0;
	wire w_dff_A_GyWwAoU22_0;
	wire w_dff_A_d6NfiNZk9_0;
	wire w_dff_A_nQjZMv2Z3_0;
	wire w_dff_A_DLXQ7I4y1_0;
	wire w_dff_A_8fr7v03Q2_1;
	wire w_dff_A_tbv4vpEC2_1;
	wire w_dff_A_wB53yctj1_1;
	wire w_dff_A_HDrtb0766_1;
	wire w_dff_A_FBjp5dQp3_1;
	wire w_dff_A_Twfgu76Y8_1;
	wire w_dff_A_JQ4u0kL94_1;
	wire w_dff_B_OtlWnwt38_0;
	wire w_dff_B_bJlIOEmW7_0;
	wire w_dff_B_Ub5k3Qmg1_0;
	wire w_dff_B_3PvvBRdj4_0;
	wire w_dff_B_29CtSvsd5_0;
	wire w_dff_A_ei9AeArb4_0;
	wire w_dff_A_5Rn2GySe6_0;
	wire w_dff_A_dPkZWSHH0_0;
	wire w_dff_A_jhpVUb811_0;
	wire w_dff_A_4loqmFTX5_0;
	wire w_dff_A_BInmhQ7F2_0;
	wire w_dff_A_8cweJVTL5_0;
	wire w_dff_A_ViIO1gdv5_0;
	wire w_dff_A_J7WFVJ3E4_0;
	wire w_dff_A_CZl9vFKP7_0;
	wire w_dff_A_mzRyPqYu8_0;
	wire w_dff_A_UkWEbEk67_0;
	wire w_dff_A_jSimQT6m3_0;
	wire w_dff_A_C0jF9Z4a8_0;
	wire w_dff_A_BqdGOZ8i7_0;
	wire w_dff_A_rrp1YvzQ8_0;
	wire w_dff_A_iNJ3xtnk4_0;
	wire w_dff_A_nBgdbj7t8_0;
	wire w_dff_A_rf9Ws4F31_0;
	wire w_dff_A_1ABIOUda5_0;
	wire w_dff_A_YOfJcjuf3_0;
	wire w_dff_A_n8lNJukw4_0;
	wire w_dff_A_g79ngoGE2_0;
	wire w_dff_A_TAB9VUeP6_0;
	wire w_dff_A_gw1HYg6z4_0;
	wire w_dff_A_G7FaBxIB0_0;
	wire w_dff_A_tsgfsOQt0_0;
	wire w_dff_A_UX0JaKHb1_0;
	wire w_dff_A_DBwfIG8f6_0;
	wire w_dff_A_iXzoPtDu5_0;
	wire w_dff_A_Fks5oyfD1_0;
	wire w_dff_A_dMdFt7Q74_0;
	wire w_dff_A_MUo3cpeH9_0;
	wire w_dff_A_TaTnHh3p2_0;
	wire w_dff_A_HgvRYNAg7_0;
	wire w_dff_A_wbajDwLD2_0;
	wire w_dff_A_611kaBzC1_0;
	wire w_dff_A_gOuz1BdX3_0;
	wire w_dff_A_MZFWZ5Ck2_0;
	wire w_dff_A_lRBjIQnH6_0;
	wire w_dff_A_aAR5BkXZ8_0;
	wire w_dff_A_WbfoVMih3_0;
	wire w_dff_A_4odZ5Z5s2_0;
	wire w_dff_A_KQTkJy614_0;
	wire w_dff_A_3vhBMoxG3_0;
	wire w_dff_B_7QJYiEzJ9_1;
	wire w_dff_A_YSxIqE1F7_0;
	wire w_dff_A_vHg0tNUU3_0;
	wire w_dff_A_bQfLeDv21_0;
	wire w_dff_A_z5LF2SNo9_0;
	wire w_dff_A_vtb5Xuwr3_0;
	wire w_dff_A_F4mDHL5g2_0;
	wire w_dff_A_hNoqOqaQ4_0;
	wire w_dff_A_phovm6tY2_0;
	wire w_dff_A_hmlgpLnG1_0;
	wire w_dff_A_ZJowE0C39_0;
	wire w_dff_A_pu9xypF90_0;
	wire w_dff_A_Py0C3wr08_0;
	wire w_dff_B_UErZ2wEc0_1;
	wire w_dff_B_Mu6LO9Ko9_1;
	wire w_dff_B_a4MScE0T5_1;
	wire w_dff_B_P1PksuTA7_1;
	wire w_dff_B_dGfsQuAp3_1;
	wire w_dff_B_etYSBqrZ6_1;
	wire w_dff_A_DNHgzYTT8_0;
	wire w_dff_A_jdtgZKU72_0;
	wire w_dff_A_g9dnEfBq9_0;
	wire w_dff_A_qNwu4S5v0_0;
	wire w_dff_B_jGV4q4nI8_2;
	wire w_dff_B_FO9BZqkR4_0;
	wire w_dff_B_rKg1oiLt3_0;
	wire w_dff_B_00o5uWn50_0;
	wire w_dff_B_qd0v0rlh4_0;
	wire w_dff_A_l0xrVePn7_0;
	wire w_dff_A_Fn7lYF5u0_0;
	wire w_dff_A_XiqxT8H98_0;
	wire w_dff_A_W31yEjFY4_0;
	wire w_dff_A_SovL6pa74_0;
	wire w_dff_A_5lglyCVg7_0;
	wire w_dff_A_UOEAbDft5_0;
	wire w_dff_A_MaVyGzcw9_0;
	wire w_dff_A_d7UN6i9q9_0;
	wire w_dff_A_2WFmqAyY2_0;
	wire w_dff_A_RdW3j2tg7_0;
	wire w_dff_A_tPc41txx8_0;
	wire w_dff_A_K0Q8vH814_0;
	wire w_dff_A_snZYENbb9_0;
	wire w_dff_A_EbBtIif70_0;
	wire w_dff_A_HdLJGaXa4_0;
	wire w_dff_A_q1y7Ps4j4_0;
	wire w_dff_A_ksqqvc4Z1_0;
	wire w_dff_A_b68mxddt9_0;
	wire w_dff_A_ZWkZePY07_0;
	wire w_dff_A_N0gRZj5j4_0;
	wire w_dff_A_riHeQFHE6_0;
	wire w_dff_A_nVOQsG7n6_0;
	wire w_dff_B_1RMKlB3O8_2;
	wire w_dff_B_GHqBYcri8_2;
	wire w_dff_B_MitMw2rq6_2;
	wire w_dff_B_ZsGj56ns4_2;
	wire w_dff_B_raJoBPem6_2;
	wire w_dff_B_CjjwHvES6_2;
	wire w_dff_B_uu7pN3IV6_2;
	wire w_dff_B_EY1iwMLf3_2;
	wire w_dff_B_d4jRyJJU8_2;
	wire w_dff_B_zYeVc9io1_2;
	wire w_dff_B_IisnITKx8_2;
	wire w_dff_B_7pA7L4v44_2;
	wire w_dff_B_cFVYd2oZ9_2;
	wire w_dff_B_rH6yLkox9_2;
	wire w_dff_A_qYlLBGYy1_0;
	wire w_dff_A_VFpAPUid0_0;
	wire w_dff_A_fypEEtHL9_0;
	wire w_dff_A_iXtCRgK81_0;
	wire w_dff_A_dPXEFUnt2_0;
	wire w_dff_A_byao8ojn3_0;
	wire w_dff_A_Nz4JYgoN5_0;
	wire w_dff_A_tD70mO059_0;
	wire w_dff_A_wBbd1NFf0_0;
	wire w_dff_A_PSvwrhod2_0;
	wire w_dff_A_gZmKyWcn5_0;
	wire w_dff_A_NcqFU0L58_0;
	wire w_dff_A_zRXLERNM2_0;
	wire w_dff_A_hDPmn0dQ4_0;
	wire w_dff_A_bGOh0Hws8_0;
	wire w_dff_A_5gHrZgEA6_1;
	wire w_dff_A_NUM62JuP8_1;
	wire w_dff_A_Jpn7ckWw6_1;
	wire w_dff_A_IJkI0XNz8_1;
	wire w_dff_A_3C1lhc792_1;
	wire w_dff_A_T0s3z3sR2_1;
	wire w_dff_A_8sTp01XR0_0;
	wire w_dff_A_7sRpbc9M9_0;
	wire w_dff_A_4kYWIAMo9_0;
	wire w_dff_A_kesxjWgP2_0;
	wire w_dff_A_IN3fy6eE8_0;
	wire w_dff_A_rMk7h3SU1_0;
	wire w_dff_A_ovHUvAct6_0;
	wire w_dff_A_cQgbo2fv9_0;
	wire w_dff_A_L64DtgMK5_0;
	wire w_dff_A_v11wllnh7_0;
	wire w_dff_A_xN7FyZMI6_0;
	wire w_dff_A_nSTVCGDl6_0;
	wire w_dff_B_kpti7bC86_2;
	wire w_dff_B_nfh1bK2R7_2;
	wire w_dff_B_PGn0kuhK1_2;
	wire w_dff_B_kOqI0B0V4_2;
	wire w_dff_B_NhQ85tbn7_2;
	wire w_dff_B_XOnT76DQ5_2;
	wire w_dff_B_TIm7nUM62_2;
	wire w_dff_A_lYDmnfP84_0;
	wire w_dff_A_l3j1r9iG1_0;
	wire w_dff_A_qr19gKpt8_0;
	wire w_dff_A_i8rpnUlF6_0;
	wire w_dff_A_n9sCxsEg3_0;
	wire w_dff_A_mPue0nY78_0;
	wire w_dff_A_vEWMWh2b4_0;
	wire w_dff_A_Gsix6Qut1_0;
	wire w_dff_A_XfvMoU7F9_0;
	wire w_dff_A_X7VQjqwR9_0;
	wire w_dff_A_x7VzobFS0_0;
	wire w_dff_A_P1OKVOCo9_0;
	wire w_dff_A_3G261ipM6_0;
	wire w_dff_A_hmHrQWcu1_0;
	wire w_dff_A_4sWUQ9TC1_0;
	wire w_dff_A_Z8wK5xfT4_0;
	wire w_dff_A_SnIvS7hs7_0;
	wire w_dff_A_a9WYnEg51_0;
	wire w_dff_A_Nl0tmKmw8_0;
	wire w_dff_A_bLe8H6p09_0;
	wire w_dff_A_AIDxYJ9G6_1;
	wire w_dff_A_2AEEYJqS8_1;
	wire w_dff_A_IT9vBcB24_1;
	wire w_dff_A_xmlZg3DD4_1;
	wire w_dff_A_rrsiezFj2_0;
	wire w_dff_A_yIMOIQR95_0;
	wire w_dff_A_M2NGVda55_0;
	wire w_dff_A_YZAjzOGS5_0;
	wire w_dff_A_IXZTYsXj7_0;
	wire w_dff_A_XDhjYOjs0_0;
	wire w_dff_A_KX1ModdX8_0;
	wire w_dff_B_R8Vd1Y862_1;
	wire w_dff_B_Th0bZbSX7_1;
	wire w_dff_A_17BocApl2_0;
	wire w_dff_A_vTr7s9CO0_0;
	wire w_dff_A_2ktGVcgN2_0;
	wire w_dff_A_rc33XG8z9_0;
	wire w_dff_A_TdrK4NG03_0;
	wire w_dff_A_hu9pQrxC8_0;
	wire w_dff_A_fUwSAHnP7_0;
	wire w_dff_A_DqQU4o6f3_0;
	wire w_dff_A_FTwM55dh5_0;
	wire w_dff_A_Y85qGYMh1_0;
	wire w_dff_A_x8N6BIx90_0;
	wire w_dff_A_RrQPXJxg2_1;
	wire w_dff_A_izS0yXx20_1;
	wire w_dff_A_vpnLmV4O8_1;
	wire w_dff_A_ERz3NTiY9_1;
	wire w_dff_A_6J44yqVi5_1;
	wire w_dff_B_Rg5ppKOc6_3;
	wire w_dff_B_hZLMDhas8_3;
	wire w_dff_B_waXoQRFE5_3;
	wire w_dff_B_xmYFxO0r9_3;
	wire w_dff_B_r3VoOClJ3_3;
	wire w_dff_B_X97IjzTs3_3;
	wire w_dff_B_LBdoCohI3_3;
	wire w_dff_A_MzlYi6693_0;
	wire w_dff_A_HPLJABdF1_0;
	wire w_dff_A_X1nS95J47_0;
	wire w_dff_A_RvYCg9X30_0;
	wire w_dff_A_IeiXacB89_0;
	wire w_dff_A_GMp2h9k91_0;
	wire w_dff_A_QZcrQiBJ2_0;
	wire w_dff_A_0xg2965M0_0;
	wire w_dff_A_a03MS5ke3_1;
	wire w_dff_A_0O1lrRPI0_1;
	wire w_dff_A_t0MEXTHS5_1;
	wire w_dff_A_yfIh0WJZ2_1;
	wire w_dff_A_NKO9YvAH3_1;
	wire w_dff_A_SxUcyHIb0_1;
	wire w_dff_A_jiRfFmRG7_1;
	wire w_dff_A_rWB4pGIe4_1;
	wire w_dff_A_ljGEyeDp4_1;
	wire w_dff_A_1D1a4aev2_1;
	wire w_dff_A_RNnfeCJp4_1;
	wire w_dff_A_jJrumhP34_1;
	wire w_dff_A_AnuNYbET2_1;
	wire w_dff_A_2wiB24I18_2;
	wire w_dff_A_1bVVJn7F4_2;
	wire w_dff_A_W4iGEOUq6_2;
	wire w_dff_A_DcRihHgS3_2;
	wire w_dff_A_G06VqZMI9_2;
	wire w_dff_A_hfEZImHd0_2;
	wire w_dff_A_XnEwKKVn6_2;
	wire w_dff_A_luh1VQBJ3_2;
	wire w_dff_A_MlPnIsTV0_2;
	wire w_dff_A_sM399QWP4_2;
	wire w_dff_A_KNuj8YSH5_2;
	wire w_dff_A_RbJvjMg10_2;
	wire w_dff_A_EqMDbWfC8_2;
	wire w_dff_A_2Slsgt950_0;
	wire w_dff_A_PrMFEnlF9_0;
	wire w_dff_A_FC2xk7wu5_0;
	wire w_dff_A_fe7q5SvS8_0;
	wire w_dff_A_jI5H6wEV3_0;
	wire w_dff_A_AEVTHE0x9_0;
	wire w_dff_A_1UWHiTsb7_0;
	wire w_dff_A_Rdh9eGGB7_0;
	wire w_dff_A_EHJSa9or2_0;
	wire w_dff_A_UI3hdeyU8_0;
	wire w_dff_A_kN9ZTeBs8_0;
	wire w_dff_A_VEScWGPm7_1;
	wire w_dff_A_fGWlJH8a1_1;
	wire w_dff_A_3ENjGzBi2_1;
	wire w_dff_A_o9gC6ODv9_1;
	wire w_dff_A_fpMbBfaE7_1;
	wire w_dff_B_LRrV6wS22_3;
	wire w_dff_B_xPW0G9qm7_3;
	wire w_dff_B_vAGnO8v30_3;
	wire w_dff_B_DYsOGOrM2_3;
	wire w_dff_B_qeRTY36U7_3;
	wire w_dff_B_YD8DtHMo4_3;
	wire w_dff_B_EJOsXWCr7_3;
	wire w_dff_A_4sNZR7UB2_0;
	wire w_dff_A_ydCpUvMA4_0;
	wire w_dff_A_wE2G8o0g0_0;
	wire w_dff_A_SQIvKpWR7_0;
	wire w_dff_A_MI5SidWk4_0;
	wire w_dff_A_9VZNu7av4_0;
	wire w_dff_A_8Q1g5X928_0;
	wire w_dff_A_KxUoyAUl5_0;
	wire w_dff_A_Z44nTf0r4_1;
	wire w_dff_A_gMsWFqAx4_1;
	wire w_dff_A_XVqTyLLg2_1;
	wire w_dff_A_7mgSZIR06_1;
	wire w_dff_A_CoxH234X8_1;
	wire w_dff_A_oJIPV0cc2_1;
	wire w_dff_A_wOo4d2rT9_1;
	wire w_dff_A_wzBecpQF9_1;
	wire w_dff_A_PtGVaBZo1_1;
	wire w_dff_A_3uqCe2780_1;
	wire w_dff_A_CKmFsCV74_1;
	wire w_dff_A_BPEcofBo1_1;
	wire w_dff_A_hYqOcECy2_1;
	wire w_dff_A_fR8Cs5L65_2;
	wire w_dff_A_YGZtKVcG9_2;
	wire w_dff_A_DUWNIw329_2;
	wire w_dff_A_IpLVUsRp4_2;
	wire w_dff_A_vv7Ix2Cr4_2;
	wire w_dff_A_Q3dAwGgf1_2;
	wire w_dff_A_4Gh2no2J3_2;
	wire w_dff_A_LnRsB3X39_2;
	wire w_dff_A_0LKmHaRj2_2;
	wire w_dff_A_C6EnUrQ51_2;
	wire w_dff_A_xHBjpzyj3_2;
	wire w_dff_A_W5z35fdo1_2;
	wire w_dff_A_odwdWGJj5_2;
	wire w_dff_B_OxpkzM984_0;
	wire w_dff_A_9KITWTJo0_1;
	wire w_dff_A_bZnqd2iU8_1;
	wire w_dff_A_w4H13SsZ4_1;
	wire w_dff_A_mB1PvCTJ0_1;
	wire w_dff_A_iqB8XFrz2_1;
	wire w_dff_A_IYSUvkzA5_0;
	wire w_dff_A_WTy4IQS20_0;
	wire w_dff_A_7ywQi2RU4_0;
	wire w_dff_A_ynTSB2Wr9_0;
	wire w_dff_A_gDkAM4OE9_0;
	wire w_dff_A_shGNqpox9_0;
	wire w_dff_A_6dYPZCWG4_0;
	wire w_dff_A_OAxUb3DU5_0;
	wire w_dff_A_rHUgqz9x2_0;
	wire w_dff_A_wTbqIYQi7_0;
	wire w_dff_A_4QaiZaVe2_0;
	wire w_dff_A_W7Zzlw3Y0_0;
	wire w_dff_A_vB3sY1hH0_0;
	wire w_dff_B_EPHpvZa76_1;
	wire w_dff_B_fNTkLBlZ1_1;
	wire w_dff_B_64Fn2s6K4_1;
	wire w_dff_B_VvAtyVfB2_1;
	wire w_dff_B_ntOmAcnj5_1;
	wire w_dff_B_SoKwzb5s1_1;
	wire w_dff_B_tSMI6Fck6_1;
	wire w_dff_A_bLvtzvXe2_0;
	wire w_dff_A_4TAxMss03_0;
	wire w_dff_A_ZnYSqwsH8_0;
	wire w_dff_A_XLJaHVqe4_0;
	wire w_dff_A_vxBEYnpb6_0;
	wire w_dff_A_YdNyOqj98_0;
	wire w_dff_A_N64fzS6w5_0;
	wire w_dff_A_5cSTr67n4_0;
	wire w_dff_A_BrOy5uzJ3_0;
	wire w_dff_A_VFqIDk5p9_0;
	wire w_dff_A_dPrwv1Md1_0;
	wire w_dff_A_TadI1wsu9_0;
	wire w_dff_A_XVlost7X3_0;
	wire w_dff_A_6g67yAoj4_1;
	wire w_dff_A_sFUuqw4y0_1;
	wire w_dff_A_7uTFjCQq5_1;
	wire w_dff_A_9VpKTKMg0_1;
	wire w_dff_A_k2b9yXf68_1;
	wire w_dff_A_IABRNTZn5_1;
	wire w_dff_A_UkJN3UFC4_1;
	wire w_dff_A_MIEOTvSw8_1;
	wire w_dff_A_LZ7sZsWZ2_0;
	wire w_dff_A_31Pa4CSX5_0;
	wire w_dff_A_PgHy2STv3_0;
	wire w_dff_A_ovK79HB99_0;
	wire w_dff_A_P81jYeST0_0;
	wire w_dff_A_Kmbdn2pq0_0;
	wire w_dff_A_KTZTvfx64_0;
	wire w_dff_A_M8D3VRA67_0;
	wire w_dff_A_DXFXV68v4_0;
	wire w_dff_A_dZP5vuZV4_0;
	wire w_dff_A_xW8HEi8H2_0;
	wire w_dff_A_HIezcUiV6_0;
	wire w_dff_A_IsorQJC72_0;
	wire w_dff_A_RQDElPUt8_0;
	wire w_dff_A_cExgftl28_0;
	wire w_dff_A_2v7fzme99_0;
	wire w_dff_A_sM0Ik8On6_0;
	wire w_dff_A_4i5nevIg5_0;
	wire w_dff_A_69Mmyz0e6_0;
	wire w_dff_A_pBI6V4ut8_0;
	wire w_dff_A_GoDra4tL5_0;
	wire w_dff_A_8FvCFuRb6_2;
	wire w_dff_A_4ZitChP85_2;
	wire w_dff_A_mhRoJZen2_2;
	wire w_dff_A_4jkALRE69_2;
	wire w_dff_A_njfgyGdm0_2;
	wire w_dff_A_NeRgcosv0_2;
	wire w_dff_A_Tlk99gAy3_2;
	wire w_dff_A_SSDLaLU77_2;
	wire w_dff_A_thL9YslX9_0;
	wire w_dff_A_EY6ZkTN12_0;
	wire w_dff_A_7wF21ChK9_0;
	wire w_dff_A_wzD724kr5_0;
	wire w_dff_A_VPU98HRn1_0;
	wire w_dff_A_We3bCPNw9_0;
	wire w_dff_A_FLRW1MjS4_0;
	wire w_dff_A_C7hbJVIu8_0;
	wire w_dff_A_V4BXIRs30_0;
	wire w_dff_A_0PJCXc3l6_0;
	wire w_dff_A_SSyHuhK77_0;
	wire w_dff_B_Jj7uKu7q3_2;
	wire w_dff_B_4VdugBgu9_2;
	wire w_dff_B_r5HOOpVi9_2;
	wire w_dff_B_gIGqkwep0_2;
	wire w_dff_B_DzEb7Z7n0_2;
	wire w_dff_B_kGcL2mV18_2;
	wire w_dff_B_h679x01V9_2;
	wire w_dff_A_npfovwcA0_0;
	wire w_dff_A_KNLGmZ9N0_0;
	wire w_dff_A_u12ccG5M8_0;
	wire w_dff_A_WRMxSBoA1_0;
	wire w_dff_A_JW9tXFPc7_0;
	wire w_dff_A_K9maBX633_0;
	wire w_dff_A_GUuDysUB7_0;
	wire w_dff_A_BOA3bU9v4_0;
	wire w_dff_A_I34zNpAM8_0;
	wire w_dff_A_AIgkchZt2_0;
	wire w_dff_A_bRt1qN9Y2_0;
	wire w_dff_A_B6WMj8OW4_0;
	wire w_dff_A_5IvxTNcM1_0;
	wire w_dff_A_D2AQoDto8_1;
	wire w_dff_A_F0JIs2ES0_1;
	wire w_dff_A_qq3yqkYQ5_1;
	wire w_dff_A_1GqXu33B7_1;
	wire w_dff_A_iYiCIsi58_1;
	wire w_dff_A_zn5Q2Ay87_1;
	wire w_dff_A_SfmIrGl77_1;
	wire w_dff_A_BvsG1iB14_1;
	wire w_dff_B_IJ05LnsU1_1;
	wire w_dff_B_ew6Sx7Ne9_1;
	wire w_dff_B_aXFrSv8w7_1;
	wire w_dff_B_7Zx3y7Us8_1;
	wire w_dff_B_A9CJi3bf1_1;
	wire w_dff_B_rIw6Z5jZ4_1;
	wire w_dff_B_skShDEEj8_1;
	wire w_dff_A_Mt602y425_0;
	wire w_dff_A_72bOw33v7_0;
	wire w_dff_A_edKtgtQS9_0;
	wire w_dff_A_CFuS4ITS1_0;
	wire w_dff_A_WN3BflP03_0;
	wire w_dff_A_6BQ4Y8TJ5_0;
	wire w_dff_A_2L1IILG65_0;
	wire w_dff_A_Iv4WggU41_0;
	wire w_dff_A_lelpZt550_1;
	wire w_dff_A_7xEU8tmF5_1;
	wire w_dff_A_RkC3auJn0_1;
	wire w_dff_A_X1aMSfV56_1;
	wire w_dff_A_lqQhWsMo4_1;
	wire w_dff_A_CqUumgaR1_1;
	wire w_dff_A_nJQwknpe5_1;
	wire w_dff_A_CYrxnjOJ4_1;
	wire w_dff_A_HHvFAjYp5_1;
	wire w_dff_A_0LkbZkY76_1;
	wire w_dff_A_VxKs87dm2_1;
	wire w_dff_A_Jy1b7IgE2_1;
	wire w_dff_A_zFpJtcqW2_1;
	wire w_dff_A_pWXp4vsy2_0;
	wire w_dff_A_sP9n6fSY2_0;
	wire w_dff_A_F9VmtyYp4_0;
	wire w_dff_A_lq5UdQm82_0;
	wire w_dff_A_xf8KplPu3_0;
	wire w_dff_A_xqRTKSaT0_0;
	wire w_dff_A_PUbLdDxi5_0;
	wire w_dff_A_QBaKjAdo9_0;
	wire w_dff_A_x2bDx4899_0;
	wire w_dff_A_0vGZdjVW1_0;
	wire w_dff_A_bCX2syvd0_0;
	wire w_dff_B_DaPTXosg2_2;
	wire w_dff_B_ieMcNlbn2_2;
	wire w_dff_B_5NCSWqyk2_2;
	wire w_dff_B_siupd1yj1_2;
	wire w_dff_B_5GhNvbGW6_2;
	wire w_dff_B_q0QwYz7j9_2;
	wire w_dff_B_BizbFXHl3_2;
	wire w_dff_A_xbKsiBUT5_0;
	wire w_dff_A_JEwyRUtL0_0;
	wire w_dff_A_3r4JC1MJ3_0;
	wire w_dff_A_O0gGAdDj6_0;
	wire w_dff_A_j1dnkyj72_0;
	wire w_dff_A_HnFjcwHr2_0;
	wire w_dff_A_J9WtIdK89_0;
	wire w_dff_A_ujRWl8j44_0;
	wire w_dff_A_Eif8ZCn13_0;
	wire w_dff_A_Ls9hETGk0_0;
	wire w_dff_A_8uf4SsJY1_0;
	wire w_dff_A_ya1dKjcZ0_0;
	wire w_dff_A_zvrtZD2z1_0;
	wire w_dff_A_j31M95Bd6_1;
	wire w_dff_A_cTv2D6Mn4_1;
	wire w_dff_A_1Ath8SQi0_1;
	wire w_dff_A_TIygiPDq1_1;
	wire w_dff_A_6Jt16Kt93_1;
	wire w_dff_A_i5Bt9W5t0_1;
	wire w_dff_A_m2iUUgfu3_1;
	wire w_dff_A_gXl3cTPm5_1;
	wire w_dff_A_8dUrqxJt2_0;
	wire w_dff_A_xbuxGv9b1_0;
	wire w_dff_A_Ho34elWX7_0;
	wire w_dff_A_QVC2PP3K9_0;
	wire w_dff_A_vA50aHIf9_0;
	wire w_dff_A_NfiY4DDd3_0;
	wire w_dff_B_9Upy40qx2_1;
	wire w_dff_B_b5MS3O9c2_1;
	wire w_dff_A_8irem2iX5_0;
	wire w_dff_A_eRB3XE5l9_0;
	wire w_dff_A_FfMnSgAs2_0;
	wire w_dff_A_mGhUST8d8_0;
	wire w_dff_A_rd5Omw5k0_0;
	wire w_dff_A_pb3yzhzd3_0;
	wire w_dff_A_DGdJol9C3_0;
	wire w_dff_A_7FLBCUWu0_0;
	wire w_dff_A_YfDKkGva9_0;
	wire w_dff_A_XjLcVCgl3_0;
	wire w_dff_A_A882PPX87_0;
	wire w_dff_A_jRPjoRYT8_0;
	wire w_dff_A_WzpsQQq57_0;
	wire w_dff_A_uHGqXqSF9_0;
	wire w_dff_A_IxigYVKC4_0;
	wire w_dff_A_Cob9RQFo2_0;
	wire w_dff_A_JSSKEe3r4_0;
	wire w_dff_A_2L284IBN8_0;
	wire w_dff_A_sbiRWCr15_0;
	wire w_dff_A_u6jPLFcV4_0;
	wire w_dff_A_GYDNLt7Q0_0;
	wire w_dff_A_Xdcuj0cd8_0;
	wire w_dff_A_yYj7vxl72_0;
	wire w_dff_A_6hUcOWcz2_0;
	wire w_dff_A_HygIf3FV6_0;
	wire w_dff_A_z1jmVMXQ2_0;
	wire w_dff_A_Gs98PXer8_0;
	wire w_dff_A_LcucVDKL2_0;
	wire w_dff_A_HXtgFlgA3_0;
	wire w_dff_A_9MrS5y7K5_0;
	wire w_dff_A_hI03JWLr2_0;
	wire w_dff_A_0ZCutWDk7_0;
	wire w_dff_A_dYRBYl1F6_0;
	wire w_dff_A_e5q9SpBs2_0;
	wire w_dff_A_SoPJwzNr1_0;
	wire w_dff_A_Sr1VNf7C3_0;
	wire w_dff_A_vBexnnKd3_0;
	wire w_dff_A_BqZu15C15_0;
	wire w_dff_A_ArlNSiEQ7_0;
	wire w_dff_A_S8vp1hBI6_0;
	wire w_dff_A_TpYjo0lD4_0;
	wire w_dff_A_ouHNtJo78_0;
	wire w_dff_A_cGt8BaJC9_0;
	wire w_dff_A_sDxS30GO9_0;
	wire w_dff_A_AppzSTfM1_0;
	wire w_dff_A_UcvP5oGh2_0;
	wire w_dff_A_JX7moqiu4_0;
	wire w_dff_A_xEFovKgy0_0;
	wire w_dff_A_UJyy5Pf67_0;
	wire w_dff_A_7jIEFFPy1_0;
	wire w_dff_A_H27ZvLKe0_0;
	wire w_dff_A_RmbDk14d7_0;
	wire w_dff_A_sE9D6LVt2_0;
	wire w_dff_A_2SuVzH7c7_0;
	wire w_dff_A_LwcZ7WBl8_0;
	wire w_dff_B_2QrGcgoq9_2;
	wire w_dff_B_jk43HwGo6_2;
	wire w_dff_B_FL6lkWnD8_2;
	wire w_dff_B_luMftctM9_2;
	wire w_dff_B_WSCq9NLs6_2;
	wire w_dff_B_Vb5fUudZ6_2;
	wire w_dff_B_6Fxb3ivR9_2;
	wire w_dff_A_L28j0QWF9_0;
	wire w_dff_A_rrbJJwxk8_0;
	wire w_dff_A_nGzq8QVI2_0;
	wire w_dff_A_6AfqpOUm1_0;
	wire w_dff_A_eBqsggGa9_0;
	wire w_dff_A_ckHjfnbY0_0;
	wire w_dff_A_qIQfrjFk5_0;
	wire w_dff_A_2axH7m6q0_0;
	wire w_dff_A_HLkrLkLw5_0;
	wire w_dff_A_99P4KDl67_0;
	wire w_dff_A_AcqvjvjU5_0;
	wire w_dff_A_x8RWZbBH7_0;
	wire w_dff_A_pegk6xgq3_0;
	wire w_dff_A_7qSynyHz9_1;
	wire w_dff_A_dcrecD3A9_1;
	wire w_dff_A_qdw1jxH20_1;
	wire w_dff_A_AHavIrtC5_1;
	wire w_dff_A_tKobfIKP3_1;
	wire w_dff_A_dUMxbQmC7_1;
	wire w_dff_A_5mEYVwFM4_1;
	wire w_dff_A_zZ0sUR6U8_1;
	wire w_dff_A_eGX8fAJW5_1;
	wire w_dff_A_nOxwyhP22_1;
	wire w_dff_A_ByprSnQp6_1;
	wire w_dff_A_jolfjana6_1;
	wire w_dff_A_72BsNdOV6_1;
	wire w_dff_A_C2h2upGr0_1;
	wire w_dff_B_ZTmTrgcu9_1;
	wire w_dff_B_I9OydJlB7_1;
	wire w_dff_A_m0sInY1m1_0;
	wire w_dff_A_3Dc8BMAJ9_0;
	wire w_dff_A_nrw18G6x9_0;
	wire w_dff_A_ouLpvPEl1_0;
	wire w_dff_A_dZSeG2ZM7_0;
	wire w_dff_A_1WMRYPC81_0;
	wire w_dff_A_tpsFSx6J9_0;
	wire w_dff_A_7F2z2dxM4_2;
	wire w_dff_A_60Y4Uhit5_0;
	wire w_dff_A_MuYsHldj5_0;
	wire w_dff_A_G1JoxGCM6_0;
	wire w_dff_A_RFEZJnl40_0;
	wire w_dff_A_GkI62Qcc3_0;
	wire w_dff_A_lo6C9lXj9_0;
	wire w_dff_A_UwSJewNF0_0;
	wire w_dff_A_m9Pfbm2e3_0;
	wire w_dff_A_iJCxKET37_0;
	wire w_dff_A_w0JUjoKL0_0;
	wire w_dff_A_kvUPm0Tm4_0;
	wire w_dff_A_iqGXefEK4_1;
	wire w_dff_A_m1Rysvbr1_0;
	wire w_dff_A_Gousxmok7_0;
	wire w_dff_A_JB0l18RT8_0;
	wire w_dff_A_y949gqVK7_0;
	wire w_dff_A_zAKZk9uM8_0;
	wire w_dff_A_aYsJW7np3_0;
	wire w_dff_A_XftsmayI7_0;
	wire w_dff_A_5nWOZrJr0_0;
	wire w_dff_A_Z9GL0bfx9_0;
	wire w_dff_A_RUtWmEfy5_0;
	wire w_dff_A_tsCGXlx34_0;
	wire w_dff_A_Q3mVMiD52_1;
	wire w_dff_A_xqVvE7FQ0_0;
	wire w_dff_A_SzlcahD08_0;
	wire w_dff_A_mLsCDeGM0_0;
	wire w_dff_A_9TsmqOJa7_0;
	wire w_dff_A_aKxb2sx62_0;
	wire w_dff_A_EzaegSGS2_0;
	wire w_dff_A_5Rl7pigT2_0;
	wire w_dff_A_ZzxpXh6n8_2;
	wire w_dff_A_AfpWvbmb9_0;
	wire w_dff_A_Du2r85SN2_0;
	wire w_dff_A_3ImWQwDu0_0;
	wire w_dff_A_o3lMAH8V8_0;
	wire w_dff_A_oqonIYtI2_0;
	wire w_dff_A_M1ZIXeKr5_0;
	wire w_dff_A_OWM6QZ776_0;
	wire w_dff_A_oQFHcsza7_0;
	wire w_dff_A_PKQIMobn7_0;
	wire w_dff_A_GSoTnHDN7_0;
	wire w_dff_A_eWfgcqh78_0;
	wire w_dff_A_RlI2Qcna3_1;
	wire w_dff_A_7MrcKX5J9_0;
	wire w_dff_A_WImJVBCU5_0;
	wire w_dff_A_XS8WfAbQ8_0;
	wire w_dff_A_oAuVrjTh2_0;
	wire w_dff_A_wTo6EMEo6_0;
	wire w_dff_A_myFTa8io4_0;
	wire w_dff_A_8oZTMSvm4_0;
	wire w_dff_A_PSQlRAdH8_2;
	wire w_dff_A_HjkXD14a0_0;
	wire w_dff_A_MdplED1k8_0;
	wire w_dff_A_vGlJWgTm6_0;
	wire w_dff_A_yDlyhauR5_0;
	wire w_dff_A_MoIFUcYl8_0;
	wire w_dff_A_cylKugpA0_0;
	wire w_dff_A_3gdH3ebS3_0;
	wire w_dff_A_2qbSh4JH6_0;
	wire w_dff_A_nNliNcVk0_0;
	wire w_dff_A_UqHDisAR2_0;
	wire w_dff_A_yqszvjhP7_0;
	wire w_dff_A_fZAokQjO4_1;
	wire w_dff_A_gmylrXXx0_0;
	wire w_dff_A_0fgqE8Kz5_0;
	wire w_dff_A_fy5GKzb95_0;
	wire w_dff_A_PSCNUDYL1_0;
	wire w_dff_A_B8bZDcuL7_0;
	wire w_dff_A_t8vsKhgU5_0;
	wire w_dff_A_MerAvAjZ2_0;
	wire w_dff_A_feB0LyTG2_2;
	wire w_dff_A_B6CDKI960_0;
	wire w_dff_A_xKnT3vzv1_0;
	wire w_dff_A_SSZHLRx26_0;
	wire w_dff_A_kr4MV6vP6_0;
	wire w_dff_A_Y6Is4uHB3_0;
	wire w_dff_A_UQ3rpyYD5_0;
	wire w_dff_A_7RxetT275_0;
	wire w_dff_A_xGO0DJLT6_0;
	wire w_dff_A_RvGw6Mad9_0;
	wire w_dff_A_42MKd7dj8_0;
	wire w_dff_A_JVwcaE8v5_0;
	wire w_dff_A_SyCFXrVg8_1;
	wire w_dff_A_fgJvJHUp2_0;
	wire w_dff_A_pjuNTLqz7_0;
	wire w_dff_A_d4ivGA2H9_0;
	wire w_dff_A_HzQF8z6P4_0;
	wire w_dff_A_CMzcZLjl3_1;
	wire w_dff_A_aCVhvqVc9_1;
	wire w_dff_A_SsxNEVmU4_2;
	wire w_dff_A_pQNMbzjP3_0;
	wire w_dff_A_NTImuhhq4_0;
	wire w_dff_A_Sr3ZIu6M7_0;
	wire w_dff_A_7q3qe1un9_0;
	wire w_dff_A_cEPna7T99_0;
	wire w_dff_A_HnbCd5xA0_0;
	wire w_dff_A_v7PrjEij8_1;
	wire w_dff_A_hpcNk6DJ6_0;
	wire w_dff_A_eJ6lv5Nq6_0;
	wire w_dff_A_Td5rJ0GL6_0;
	wire w_dff_A_4DB5y1E77_0;
	wire w_dff_A_AXRfQW691_0;
	wire w_dff_A_gznuvzvn9_0;
	wire w_dff_A_9XREv33Q7_0;
	wire w_dff_A_qtP09Y1i3_2;
	wire w_dff_A_u4JIynEO0_0;
	wire w_dff_A_nK6Fl9I16_0;
	wire w_dff_A_sGWpZJRV3_0;
	wire w_dff_A_Io2t5ywt9_0;
	wire w_dff_A_8u08u7938_0;
	wire w_dff_A_pWsDNIww7_0;
	wire w_dff_A_kZ6Mg0QT4_0;
	wire w_dff_A_JfXK5fDd6_0;
	wire w_dff_A_JZs7SXJM8_0;
	wire w_dff_A_DLfZkeoe3_0;
	wire w_dff_A_O2O27OSV9_0;
	wire w_dff_A_6clacpgG8_1;
	wire w_dff_A_UcNEqn591_1;
	wire w_dff_A_7Aba9wMw0_0;
	wire w_dff_A_ZYe2mqew6_1;
	wire w_dff_A_jv5CgRg97_1;
	wire w_dff_A_YfDeoaEH9_1;
	wire w_dff_A_dh8ZkW9p9_1;
	wire w_dff_A_G5HHThQx3_1;
	wire w_dff_A_rgJckYea6_1;
	wire w_dff_A_6rD5F3gE5_1;
	wire w_dff_A_x4t2TTDM3_1;
	wire w_dff_A_Tptql5QN1_2;
	wire w_dff_A_vAxnWIbk1_0;
	wire w_dff_A_iVxv4iMo3_0;
	wire w_dff_A_VDHd53zs6_0;
	wire w_dff_A_zNFhhy5i7_0;
	wire w_dff_A_28XZIk1f5_0;
	wire w_dff_A_oaDmFE1v4_0;
	wire w_dff_A_mRpJm9BV8_0;
	wire w_dff_A_68YAXx8k7_0;
	wire w_dff_A_jdw8FYVD9_0;
	wire w_dff_A_HaarqPA04_0;
	wire w_dff_A_5BVq9ZHi3_0;
	wire w_dff_A_82iLS9kc4_0;
	wire w_dff_A_Ewd8aq8n9_0;
	wire w_dff_A_Df6kt6vf1_0;
	wire w_dff_A_09oEh0fq3_0;
	wire w_dff_A_z76xChqN8_0;
	wire w_dff_A_xxSMbtcd9_0;
	wire w_dff_A_5h1yS6Ot2_0;
	wire w_dff_A_gogxqGJE4_0;
	wire w_dff_A_zypnxrKF1_0;
	wire w_dff_A_odgcXlMO1_0;
	wire w_dff_A_r7nhHJni2_0;
	wire w_dff_A_C9ORlX8z2_0;
	wire w_dff_A_zUeWR0hQ4_0;
	wire w_dff_A_RLzJUKcF1_2;
	wire w_dff_A_d8DihoTb7_1;
	wire w_dff_A_DRAlncLY7_1;
	wire w_dff_A_Owjh0MPB3_1;
	wire w_dff_A_FvCoEDqA2_1;
	wire w_dff_A_8h3ouYZx8_1;
	wire w_dff_A_8hPUmbJ85_1;
	wire w_dff_A_4a4TCm1X8_1;
	wire w_dff_A_K8cZEKKZ3_1;
	wire w_dff_A_dUtqgqT51_1;
	wire w_dff_A_H1wOdVD85_1;
	wire w_dff_A_HYZ0eSaV6_1;
	wire w_dff_A_eR5k1xLC3_1;
	wire w_dff_A_7WCVBsNf6_1;
	wire w_dff_A_njq90PmN5_1;
	wire w_dff_A_QH0Pbqzg0_1;
	wire w_dff_A_4UWrYcH12_2;
	wire w_dff_A_7XPuTqfg9_0;
	wire w_dff_A_5vwQD4ir1_0;
	wire w_dff_A_06LKmq1Y4_0;
	wire w_dff_A_LeAI5wVU6_0;
	wire w_dff_A_Z6rZHQTN1_0;
	wire w_dff_A_j2VuPVru3_0;
	wire w_dff_A_w1Y0VbNl4_0;
	wire w_dff_A_B4PSvxED7_0;
	wire w_dff_A_WqI6xG6K3_0;
	wire w_dff_A_XGDkbvox3_0;
	wire w_dff_A_6BtpPbvh9_0;
	wire w_dff_A_7tzXGZCE4_0;
	wire w_dff_A_zGS1JHWz9_0;
	wire w_dff_A_vSSdYcUY8_0;
	wire w_dff_A_U0vy50sd4_0;
	wire w_dff_A_v3i3QIfk4_0;
	wire w_dff_A_jY6g6WIn8_0;
	wire w_dff_A_NN15yFkb0_0;
	wire w_dff_A_n83oLjKe0_0;
	wire w_dff_A_G75mAGmL5_1;
	wire w_dff_A_mN0xSzlM8_0;
	wire w_dff_A_CoALeAd62_0;
	wire w_dff_A_GzS1AfhY6_0;
	wire w_dff_A_2ZIvObef1_0;
	wire w_dff_A_SbcVLWP72_0;
	wire w_dff_A_dQKALZtM9_0;
	wire w_dff_A_ik9sEIgh2_0;
	wire w_dff_A_5TF4eyZ79_0;
	wire w_dff_A_M6MKkLdS8_0;
	wire w_dff_A_lwVELHM53_0;
	wire w_dff_A_NWMctVa41_0;
	wire w_dff_A_7T7WMs6T4_0;
	wire w_dff_A_JCVWIwh73_1;
	wire w_dff_A_7QbPNyfA3_0;
	wire w_dff_A_MK8mbjgS5_0;
	wire w_dff_A_6Ut5Kybk8_0;
	wire w_dff_A_HUwmCVVV9_0;
	wire w_dff_A_02IdJ8190_0;
	wire w_dff_A_xghxYD4R6_1;
	wire w_dff_A_TvqwLfSQ7_0;
	jnot g000(.din(w_G76gat_0[1]),.dout(n43),.clk(gclk));
	jand g001(.dina(w_G82gat_0[2]),.dinb(w_n43_0[1]),.dout(n44),.clk(gclk));
	jnot g002(.din(w_G24gat_0[1]),.dout(n45),.clk(gclk));
	jand g003(.dina(w_G30gat_0[1]),.dinb(n45),.dout(n46),.clk(gclk));
	jnot g004(.din(w_G11gat_0[2]),.dout(n47),.clk(gclk));
	jand g005(.dina(w_G17gat_0[2]),.dinb(w_n47_0[1]),.dout(n48),.clk(gclk));
	jor g006(.dina(n48),.dinb(n46),.dout(n49),.clk(gclk));
	jor g007(.dina(n49),.dinb(w_n44_0[1]),.dout(n50),.clk(gclk));
	jnot g008(.din(w_G37gat_0[2]),.dout(n51),.clk(gclk));
	jand g009(.dina(w_G43gat_1[1]),.dinb(n51),.dout(n52),.clk(gclk));
	jnot g010(.din(w_G63gat_0[2]),.dout(n53),.clk(gclk));
	jand g011(.dina(w_G69gat_0[2]),.dinb(w_n53_0[1]),.dout(n54),.clk(gclk));
	jor g012(.dina(n54),.dinb(w_n52_0[1]),.dout(n55),.clk(gclk));
	jnot g013(.din(w_G102gat_0[2]),.dout(n56),.clk(gclk));
	jand g014(.dina(w_G108gat_0[2]),.dinb(w_n56_0[1]),.dout(n57),.clk(gclk));
	jnot g015(.din(w_G50gat_0[2]),.dout(n58),.clk(gclk));
	jand g016(.dina(w_G56gat_0[2]),.dinb(w_n58_0[1]),.dout(n59),.clk(gclk));
	jor g017(.dina(n59),.dinb(n57),.dout(n60),.clk(gclk));
	jnot g018(.din(w_G89gat_0[2]),.dout(n61),.clk(gclk));
	jand g019(.dina(w_G95gat_0[2]),.dinb(w_n61_0[1]),.dout(n62),.clk(gclk));
	jnot g020(.din(w_G1gat_0[2]),.dout(n63),.clk(gclk));
	jand g021(.dina(w_G4gat_0[2]),.dinb(w_n63_0[1]),.dout(n64),.clk(gclk));
	jor g022(.dina(n64),.dinb(n62),.dout(n65),.clk(gclk));
	jor g023(.dina(n65),.dinb(n60),.dout(n66),.clk(gclk));
	jor g024(.dina(n66),.dinb(w_dff_B_I9OydJlB7_1),.dout(n67),.clk(gclk));
	jor g025(.dina(n67),.dinb(w_dff_B_ZTmTrgcu9_1),.dout(G223gat_fa_),.clk(gclk));
	jnot g026(.din(w_G112gat_0[2]),.dout(n69),.clk(gclk));
	jnot g027(.din(w_n44_0[0]),.dout(n70),.clk(gclk));
	jnot g028(.din(w_G30gat_0[0]),.dout(n71),.clk(gclk));
	jor g029(.dina(w_n71_0[1]),.dinb(w_G24gat_0[0]),.dout(n72),.clk(gclk));
	jnot g030(.din(w_G17gat_0[1]),.dout(n73),.clk(gclk));
	jor g031(.dina(w_n73_0[1]),.dinb(w_G11gat_0[1]),.dout(n74),.clk(gclk));
	jand g032(.dina(n74),.dinb(w_n72_0[1]),.dout(n75),.clk(gclk));
	jand g033(.dina(n75),.dinb(n70),.dout(n76),.clk(gclk));
	jnot g034(.din(w_G43gat_1[0]),.dout(n77),.clk(gclk));
	jor g035(.dina(w_n77_0[1]),.dinb(w_G37gat_0[1]),.dout(n78),.clk(gclk));
	jnot g036(.din(w_G69gat_0[1]),.dout(n79),.clk(gclk));
	jor g037(.dina(w_n79_0[1]),.dinb(w_G63gat_0[1]),.dout(n80),.clk(gclk));
	jand g038(.dina(n80),.dinb(w_n78_0[1]),.dout(n81),.clk(gclk));
	jnot g039(.din(w_G108gat_0[1]),.dout(n82),.clk(gclk));
	jor g040(.dina(w_n82_0[1]),.dinb(w_G102gat_0[1]),.dout(n83),.clk(gclk));
	jnot g041(.din(w_G56gat_0[1]),.dout(n84),.clk(gclk));
	jor g042(.dina(w_n84_0[1]),.dinb(w_G50gat_0[1]),.dout(n85),.clk(gclk));
	jand g043(.dina(n85),.dinb(n83),.dout(n86),.clk(gclk));
	jnot g044(.din(w_G95gat_0[1]),.dout(n87),.clk(gclk));
	jor g045(.dina(w_n87_0[1]),.dinb(w_G89gat_0[1]),.dout(n88),.clk(gclk));
	jnot g046(.din(w_G4gat_0[1]),.dout(n89),.clk(gclk));
	jor g047(.dina(w_n89_0[1]),.dinb(w_G1gat_0[1]),.dout(n90),.clk(gclk));
	jand g048(.dina(n90),.dinb(n88),.dout(n91),.clk(gclk));
	jand g049(.dina(n91),.dinb(n86),.dout(n92),.clk(gclk));
	jand g050(.dina(n92),.dinb(w_dff_B_b5MS3O9c2_1),.dout(n93),.clk(gclk));
	jand g051(.dina(n93),.dinb(w_dff_B_9Upy40qx2_1),.dout(n94),.clk(gclk));
	jor g052(.dina(w_n94_4[1]),.dinb(w_n56_0[0]),.dout(n95),.clk(gclk));
	jand g053(.dina(n95),.dinb(w_G108gat_0[0]),.dout(n96),.clk(gclk));
	jand g054(.dina(w_n96_0[1]),.dinb(w_n69_0[1]),.dout(n97),.clk(gclk));
	jnot g055(.din(w_G8gat_0[2]),.dout(n98),.clk(gclk));
	jor g056(.dina(w_n94_4[0]),.dinb(w_n63_0[0]),.dout(n99),.clk(gclk));
	jand g057(.dina(n99),.dinb(w_G4gat_0[0]),.dout(n100),.clk(gclk));
	jand g058(.dina(w_n100_0[1]),.dinb(w_n98_0[1]),.dout(n101),.clk(gclk));
	jor g059(.dina(n101),.dinb(n97),.dout(n102),.clk(gclk));
	jnot g060(.din(w_G99gat_0[2]),.dout(n103),.clk(gclk));
	jor g061(.dina(w_n94_3[2]),.dinb(w_n61_0[0]),.dout(n104),.clk(gclk));
	jand g062(.dina(n104),.dinb(w_G95gat_0[0]),.dout(n105),.clk(gclk));
	jand g063(.dina(n105),.dinb(w_dff_B_skShDEEj8_1),.dout(n106),.clk(gclk));
	jnot g064(.din(w_G73gat_0[2]),.dout(n107),.clk(gclk));
	jor g065(.dina(w_n94_3[1]),.dinb(w_n53_0[0]),.dout(n108),.clk(gclk));
	jand g066(.dina(n108),.dinb(w_G69gat_0[0]),.dout(n109),.clk(gclk));
	jand g067(.dina(w_n109_0[1]),.dinb(w_n107_0[1]),.dout(n110),.clk(gclk));
	jor g068(.dina(n110),.dinb(n106),.dout(n111),.clk(gclk));
	jor g069(.dina(n111),.dinb(n102),.dout(n112),.clk(gclk));
	jxor g070(.dina(w_n94_3[0]),.dinb(w_n72_0[0]),.dout(n113),.clk(gclk));
	jor g071(.dina(n113),.dinb(w_n71_0[0]),.dout(n114),.clk(gclk));
	jor g072(.dina(w_n114_0[2]),.dinb(w_G34gat_0[2]),.dout(n115),.clk(gclk));
	jnot g073(.din(w_n115_0[1]),.dout(n116),.clk(gclk));
	jnot g074(.din(w_G60gat_0[2]),.dout(n117),.clk(gclk));
	jor g075(.dina(w_n94_2[2]),.dinb(w_n58_0[0]),.dout(n118),.clk(gclk));
	jand g076(.dina(n118),.dinb(w_G56gat_0[0]),.dout(n119),.clk(gclk));
	jand g077(.dina(w_n119_0[1]),.dinb(w_dff_B_tSMI6Fck6_1),.dout(n120),.clk(gclk));
	jxor g078(.dina(w_n94_2[1]),.dinb(w_n52_0[0]),.dout(n121),.clk(gclk));
	jnot g079(.din(w_G47gat_0[1]),.dout(n122),.clk(gclk));
	jand g080(.dina(n122),.dinb(w_G43gat_0[2]),.dout(n123),.clk(gclk));
	jand g081(.dina(w_n123_0[1]),.dinb(w_n121_0[1]),.dout(n124),.clk(gclk));
	jor g082(.dina(w_dff_B_OxpkzM984_0),.dinb(n120),.dout(n125),.clk(gclk));
	jnot g083(.din(w_G86gat_1[1]),.dout(n126),.clk(gclk));
	jor g084(.dina(w_n94_2[0]),.dinb(w_n43_0[0]),.dout(n127),.clk(gclk));
	jand g085(.dina(n127),.dinb(w_G82gat_0[1]),.dout(n128),.clk(gclk));
	jand g086(.dina(w_n128_0[1]),.dinb(w_n126_0[2]),.dout(n129),.clk(gclk));
	jnot g087(.din(w_G21gat_1[1]),.dout(n130),.clk(gclk));
	jor g088(.dina(w_n94_1[2]),.dinb(w_n47_0[0]),.dout(n131),.clk(gclk));
	jand g089(.dina(n131),.dinb(w_G17gat_0[0]),.dout(n132),.clk(gclk));
	jand g090(.dina(w_n132_0[1]),.dinb(w_n130_0[2]),.dout(n133),.clk(gclk));
	jor g091(.dina(n133),.dinb(n129),.dout(n134),.clk(gclk));
	jor g092(.dina(n134),.dinb(n125),.dout(n135),.clk(gclk));
	jor g093(.dina(n135),.dinb(w_dff_B_Th0bZbSX7_1),.dout(n136),.clk(gclk));
	jor g094(.dina(n136),.dinb(w_dff_B_R8Vd1Y862_1),.dout(G329gat_fa_),.clk(gclk));
	jand g095(.dina(w_G223gat_3[1]),.dinb(w_G89gat_0[0]),.dout(n138),.clk(gclk));
	jor g096(.dina(n138),.dinb(w_n87_0[0]),.dout(n139),.clk(gclk));
	jand g097(.dina(w_G329gat_6),.dinb(w_G99gat_0[1]),.dout(n140),.clk(gclk));
	jor g098(.dina(n140),.dinb(w_n139_0[1]),.dout(n141),.clk(gclk));
	jor g099(.dina(w_n141_0[1]),.dinb(w_G105gat_0[1]),.dout(n142),.clk(gclk));
	jnot g100(.din(w_n142_0[1]),.dout(n143),.clk(gclk));
	jand g101(.dina(w_G223gat_3[0]),.dinb(w_G50gat_0[0]),.dout(n144),.clk(gclk));
	jor g102(.dina(n144),.dinb(w_n84_0[0]),.dout(n145),.clk(gclk));
	jor g103(.dina(w_n145_0[1]),.dinb(w_G60gat_0[1]),.dout(n146),.clk(gclk));
	jand g104(.dina(w_G329gat_5[2]),.dinb(w_n146_0[1]),.dout(n147),.clk(gclk));
	jnot g105(.din(w_n147_0[1]),.dout(n148),.clk(gclk));
	jnot g106(.din(w_G66gat_0[1]),.dout(n150),.clk(gclk));
	jand g107(.dina(w_n119_0[0]),.dinb(w_n150_0[1]),.dout(n151),.clk(gclk));
	jand g108(.dina(w_n151_0[1]),.dinb(n148),.dout(n153),.clk(gclk));
	jnot g109(.din(w_G79gat_0[1]),.dout(n154),.clk(gclk));
	jand g110(.dina(w_G223gat_2[2]),.dinb(w_G102gat_0[0]),.dout(n155),.clk(gclk));
	jor g111(.dina(n155),.dinb(w_n82_0[0]),.dout(n156),.clk(gclk));
	jor g112(.dina(w_n156_0[1]),.dinb(w_G112gat_0[1]),.dout(n157),.clk(gclk));
	jand g113(.dina(w_G223gat_2[1]),.dinb(w_G1gat_0[0]),.dout(n158),.clk(gclk));
	jor g114(.dina(n158),.dinb(w_n89_0[0]),.dout(n159),.clk(gclk));
	jor g115(.dina(w_n159_0[1]),.dinb(w_G8gat_0[1]),.dout(n160),.clk(gclk));
	jand g116(.dina(n160),.dinb(n157),.dout(n161),.clk(gclk));
	jor g117(.dina(w_n139_0[0]),.dinb(w_G99gat_0[0]),.dout(n162),.clk(gclk));
	jand g118(.dina(w_G223gat_2[0]),.dinb(w_G63gat_0[0]),.dout(n163),.clk(gclk));
	jor g119(.dina(n163),.dinb(w_n79_0[0]),.dout(n164),.clk(gclk));
	jor g120(.dina(w_n164_0[1]),.dinb(w_G73gat_0[1]),.dout(n165),.clk(gclk));
	jand g121(.dina(n165),.dinb(n162),.dout(n166),.clk(gclk));
	jand g122(.dina(n166),.dinb(n161),.dout(n167),.clk(gclk));
	jxor g123(.dina(w_n94_1[1]),.dinb(w_n78_0[0]),.dout(n168),.clk(gclk));
	jnot g124(.din(w_n123_0[0]),.dout(n169),.clk(gclk));
	jor g125(.dina(w_dff_B_qd0v0rlh4_0),.dinb(n168),.dout(n170),.clk(gclk));
	jand g126(.dina(w_n170_0[1]),.dinb(w_n146_0[0]),.dout(n171),.clk(gclk));
	jnot g127(.din(w_G82gat_0[0]),.dout(n172),.clk(gclk));
	jand g128(.dina(w_G223gat_1[2]),.dinb(w_G76gat_0[0]),.dout(n173),.clk(gclk));
	jor g129(.dina(n173),.dinb(w_dff_B_etYSBqrZ6_1),.dout(n174),.clk(gclk));
	jor g130(.dina(w_n174_0[1]),.dinb(w_G86gat_1[0]),.dout(n175),.clk(gclk));
	jand g131(.dina(w_G223gat_1[1]),.dinb(w_G11gat_0[0]),.dout(n176),.clk(gclk));
	jor g132(.dina(n176),.dinb(w_n73_0[0]),.dout(n177),.clk(gclk));
	jor g133(.dina(w_n177_0[1]),.dinb(w_G21gat_1[0]),.dout(n178),.clk(gclk));
	jand g134(.dina(n178),.dinb(n175),.dout(n179),.clk(gclk));
	jand g135(.dina(n179),.dinb(n171),.dout(n180),.clk(gclk));
	jand g136(.dina(n180),.dinb(w_n115_0[0]),.dout(n181),.clk(gclk));
	jand g137(.dina(n181),.dinb(w_dff_B_7QJYiEzJ9_1),.dout(n182),.clk(gclk));
	jor g138(.dina(w_n182_3[1]),.dinb(w_n107_0[0]),.dout(n183),.clk(gclk));
	jand g139(.dina(n183),.dinb(w_n109_0[0]),.dout(n184),.clk(gclk));
	jand g140(.dina(w_n184_0[1]),.dinb(w_n154_0[1]),.dout(n185),.clk(gclk));
	jor g141(.dina(n185),.dinb(n153),.dout(n186),.clk(gclk));
	jor g142(.dina(n186),.dinb(n143),.dout(n187),.clk(gclk));
	jand g143(.dina(w_G329gat_5[1]),.dinb(w_n170_0[0]),.dout(n188),.clk(gclk));
	jnot g144(.din(w_n188_0[1]),.dout(n189),.clk(gclk));
	jnot g145(.din(w_G53gat_0[1]),.dout(n191),.clk(gclk));
	jand g146(.dina(w_n191_0[1]),.dinb(w_G43gat_0[1]),.dout(n192),.clk(gclk));
	jand g147(.dina(w_dff_B_29CtSvsd5_0),.dinb(w_n121_0[0]),.dout(n193),.clk(gclk));
	jand g148(.dina(w_n193_0[1]),.dinb(n189),.dout(n195),.clk(gclk));
	jor g149(.dina(w_n182_3[0]),.dinb(w_n130_0[1]),.dout(n196),.clk(gclk));
	jand g150(.dina(n196),.dinb(w_n132_0[0]),.dout(n197),.clk(gclk));
	jnot g151(.din(w_G27gat_0[1]),.dout(n198),.clk(gclk));
	jor g152(.dina(w_G329gat_5[0]),.dinb(w_G21gat_0[2]),.dout(n199),.clk(gclk));
	jand g153(.dina(n199),.dinb(w_n198_0[1]),.dout(n200),.clk(gclk));
	jand g154(.dina(n200),.dinb(w_n197_0[1]),.dout(n201),.clk(gclk));
	jor g155(.dina(n201),.dinb(n195),.dout(n202),.clk(gclk));
	jor g156(.dina(w_n182_2[2]),.dinb(w_n126_0[1]),.dout(n203),.clk(gclk));
	jand g157(.dina(n203),.dinb(w_n128_0[0]),.dout(n204),.clk(gclk));
	jnot g158(.din(w_G92gat_0[2]),.dout(n205),.clk(gclk));
	jor g159(.dina(w_G329gat_4[2]),.dinb(w_G86gat_0[2]),.dout(n206),.clk(gclk));
	jand g160(.dina(n206),.dinb(w_n205_0[1]),.dout(n207),.clk(gclk));
	jand g161(.dina(n207),.dinb(w_n204_0[1]),.dout(n208),.clk(gclk));
	jnot g162(.din(w_G14gat_0[2]),.dout(n209),.clk(gclk));
	jor g163(.dina(w_n182_2[1]),.dinb(w_n98_0[0]),.dout(n210),.clk(gclk));
	jand g164(.dina(n210),.dinb(w_n100_0[0]),.dout(n211),.clk(gclk));
	jand g165(.dina(n211),.dinb(w_dff_B_h2WQfTe00_1),.dout(n212),.clk(gclk));
	jor g166(.dina(n212),.dinb(n208),.dout(n213),.clk(gclk));
	jnot g167(.din(w_G34gat_0[1]),.dout(n214),.clk(gclk));
	jor g168(.dina(w_n182_2[0]),.dinb(w_dff_B_mecfc78R8_1),.dout(n215),.clk(gclk));
	jnot g169(.din(w_G40gat_0[1]),.dout(n217),.clk(gclk));
	jnot g170(.din(w_n114_0[1]),.dout(n218),.clk(gclk));
	jand g171(.dina(n218),.dinb(w_n217_0[1]),.dout(n219),.clk(gclk));
	jand g172(.dina(w_n219_0[1]),.dinb(n215),.dout(n221),.clk(gclk));
	jnot g173(.din(w_G115gat_0[1]),.dout(n222),.clk(gclk));
	jor g174(.dina(w_n182_1[2]),.dinb(w_n69_0[0]),.dout(n223),.clk(gclk));
	jand g175(.dina(n223),.dinb(w_n96_0[0]),.dout(n224),.clk(gclk));
	jand g176(.dina(w_n224_0[1]),.dinb(w_n222_0[1]),.dout(n225),.clk(gclk));
	jor g177(.dina(n225),.dinb(w_dff_B_kIK7VG9F5_1),.dout(n226),.clk(gclk));
	jor g178(.dina(n226),.dinb(n213),.dout(n227),.clk(gclk));
	jor g179(.dina(n227),.dinb(w_dff_B_GNSqXq4E6_1),.dout(n228),.clk(gclk));
	jor g180(.dina(n228),.dinb(w_dff_B_ELQB5Iqi7_1),.dout(G370gat_fa_),.clk(gclk));
	jand g181(.dina(w_G329gat_4[1]),.dinb(w_G8gat_0[0]),.dout(n230),.clk(gclk));
	jor g182(.dina(n230),.dinb(w_n159_0[0]),.dout(n231),.clk(gclk));
	jand g183(.dina(w_G370gat_2),.dinb(w_G14gat_0[1]),.dout(n232),.clk(gclk));
	jor g184(.dina(n232),.dinb(w_n231_0[1]),.dout(n233),.clk(gclk));
	jnot g185(.din(w_n151_0[0]),.dout(n235),.clk(gclk));
	jor g186(.dina(w_dff_B_4WmcnZt15_0),.dinb(w_n147_0[0]),.dout(n237),.clk(gclk));
	jand g187(.dina(w_G329gat_4[0]),.dinb(w_G73gat_0[0]),.dout(n238),.clk(gclk));
	jor g188(.dina(n238),.dinb(w_n164_0[0]),.dout(n239),.clk(gclk));
	jor g189(.dina(n239),.dinb(w_G79gat_0[0]),.dout(n240),.clk(gclk));
	jand g190(.dina(n240),.dinb(w_dff_B_LVxx1fIm2_1),.dout(n241),.clk(gclk));
	jand g191(.dina(n241),.dinb(w_n142_0[0]),.dout(n242),.clk(gclk));
	jnot g192(.din(w_n193_0[0]),.dout(n244),.clk(gclk));
	jor g193(.dina(w_dff_B_FbCoXbMV1_0),.dinb(w_n188_0[0]),.dout(n246),.clk(gclk));
	jand g194(.dina(w_G329gat_3[2]),.dinb(w_G21gat_0[1]),.dout(n247),.clk(gclk));
	jor g195(.dina(n247),.dinb(w_n177_0[0]),.dout(n248),.clk(gclk));
	jand g196(.dina(w_n182_1[1]),.dinb(w_n130_0[0]),.dout(n249),.clk(gclk));
	jor g197(.dina(n249),.dinb(w_G27gat_0[0]),.dout(n250),.clk(gclk));
	jor g198(.dina(n250),.dinb(n248),.dout(n251),.clk(gclk));
	jand g199(.dina(n251),.dinb(w_dff_B_V16kZFy51_1),.dout(n252),.clk(gclk));
	jand g200(.dina(w_G329gat_3[1]),.dinb(w_G86gat_0[1]),.dout(n253),.clk(gclk));
	jor g201(.dina(n253),.dinb(w_n174_0[0]),.dout(n254),.clk(gclk));
	jand g202(.dina(w_n182_1[0]),.dinb(w_n126_0[0]),.dout(n255),.clk(gclk));
	jor g203(.dina(n255),.dinb(w_G92gat_0[1]),.dout(n256),.clk(gclk));
	jor g204(.dina(n256),.dinb(w_n254_0[1]),.dout(n257),.clk(gclk));
	jor g205(.dina(w_n231_0[0]),.dinb(w_G14gat_0[0]),.dout(n258),.clk(gclk));
	jand g206(.dina(n258),.dinb(n257),.dout(n259),.clk(gclk));
	jand g207(.dina(w_G329gat_3[0]),.dinb(w_G34gat_0[0]),.dout(n260),.clk(gclk));
	jnot g208(.din(w_n219_0[0]),.dout(n262),.clk(gclk));
	jor g209(.dina(w_dff_B_fU6PONy31_0),.dinb(w_n260_0[1]),.dout(n264),.clk(gclk));
	jand g210(.dina(w_G329gat_2[2]),.dinb(w_G112gat_0[0]),.dout(n265),.clk(gclk));
	jor g211(.dina(n265),.dinb(w_n156_0[0]),.dout(n266),.clk(gclk));
	jor g212(.dina(n266),.dinb(w_G115gat_0[0]),.dout(n267),.clk(gclk));
	jand g213(.dina(n267),.dinb(w_dff_B_TihVYKXx0_1),.dout(n268),.clk(gclk));
	jand g214(.dina(n268),.dinb(n259),.dout(n269),.clk(gclk));
	jand g215(.dina(n269),.dinb(w_dff_B_hWCdCurf8_1),.dout(n270),.clk(gclk));
	jand g216(.dina(n270),.dinb(w_dff_B_BTec5vnc7_1),.dout(n271),.clk(gclk));
	jor g217(.dina(w_n271_3[1]),.dinb(w_n150_0[0]),.dout(n272),.clk(gclk));
	jand g218(.dina(w_G329gat_2[1]),.dinb(w_G60gat_0[0]),.dout(n273),.clk(gclk));
	jor g219(.dina(n273),.dinb(w_n145_0[0]),.dout(n274),.clk(gclk));
	jnot g220(.din(w_n274_0[1]),.dout(n275),.clk(gclk));
	jand g221(.dina(w_dff_B_9zOLbmIy1_0),.dinb(n272),.dout(n276),.clk(gclk));
	jor g222(.dina(w_n271_3[0]),.dinb(w_n191_0[0]),.dout(n277),.clk(gclk));
	jand g223(.dina(w_G329gat_2[0]),.dinb(w_G47gat_0[0]),.dout(n278),.clk(gclk));
	jand g224(.dina(w_G223gat_1[0]),.dinb(w_G37gat_0[0]),.dout(n279),.clk(gclk));
	jor g225(.dina(n279),.dinb(w_n77_0[0]),.dout(n280),.clk(gclk));
	jor g226(.dina(w_dff_B_qkWew6ny7_0),.dinb(n278),.dout(n281),.clk(gclk));
	jnot g227(.din(w_n281_0[1]),.dout(n282),.clk(gclk));
	jand g228(.dina(w_dff_B_qxgHqkJt9_0),.dinb(n277),.dout(n283),.clk(gclk));
	jor g229(.dina(w_n283_0[1]),.dinb(n276),.dout(n284),.clk(gclk));
	jor g230(.dina(w_n271_2[2]),.dinb(w_n198_0[0]),.dout(n285),.clk(gclk));
	jand g231(.dina(n285),.dinb(w_n197_0[0]),.dout(n286),.clk(gclk));
	jor g232(.dina(w_n271_2[1]),.dinb(w_n217_0[0]),.dout(n287),.clk(gclk));
	jor g233(.dina(w_n114_0[0]),.dinb(w_n260_0[0]),.dout(n290),.clk(gclk));
	jnot g234(.din(w_n290_0[1]),.dout(n291),.clk(gclk));
	jand g235(.dina(w_dff_B_dVyWw4fQ3_0),.dinb(n287),.dout(n292),.clk(gclk));
	jor g236(.dina(n292),.dinb(w_n286_0[1]),.dout(n293),.clk(gclk));
	jor g237(.dina(w_n293_0[1]),.dinb(n284),.dout(G430gat_fa_),.clk(gclk));
	jor g238(.dina(w_n271_2[0]),.dinb(w_n205_0[0]),.dout(n295),.clk(gclk));
	jand g239(.dina(n295),.dinb(w_n204_0[0]),.dout(n296),.clk(gclk));
	jor g240(.dina(w_n271_1[2]),.dinb(w_n222_0[0]),.dout(n297),.clk(gclk));
	jand g241(.dina(n297),.dinb(w_n224_0[0]),.dout(n298),.clk(gclk));
	jor g242(.dina(n298),.dinb(w_n296_0[1]),.dout(n299),.clk(gclk));
	jnot g243(.din(w_n141_0[0]),.dout(n300),.clk(gclk));
	jnot g244(.din(w_G105gat_0[0]),.dout(n301),.clk(gclk));
	jor g245(.dina(w_n271_1[1]),.dinb(w_dff_B_3EXKWv7H2_1),.dout(n302),.clk(gclk));
	jand g246(.dina(n302),.dinb(w_dff_B_kXbpKEBk3_1),.dout(n303),.clk(gclk));
	jor g247(.dina(w_n271_1[0]),.dinb(w_n154_0[0]),.dout(n304),.clk(gclk));
	jand g248(.dina(n304),.dinb(w_n184_0[0]),.dout(n305),.clk(gclk));
	jor g249(.dina(w_n305_0[1]),.dinb(w_n303_0[1]),.dout(n306),.clk(gclk));
	jor g250(.dina(n306),.dinb(n299),.dout(n307),.clk(gclk));
	jor g251(.dina(n307),.dinb(w_G430gat_0),.dout(n308),.clk(gclk));
	jand g252(.dina(n308),.dinb(w_dff_B_VIrjoWqg4_1),.dout(G421gat),.clk(gclk));
	jand g253(.dina(w_G370gat_1[2]),.dinb(w_G66gat_0[0]),.dout(n310),.clk(gclk));
	jor g254(.dina(w_n274_0[0]),.dinb(n310),.dout(n311),.clk(gclk));
	jand g255(.dina(w_G370gat_1[1]),.dinb(w_G53gat_0[0]),.dout(n312),.clk(gclk));
	jor g256(.dina(w_n281_0[0]),.dinb(n312),.dout(n313),.clk(gclk));
	jand g257(.dina(w_n313_0[1]),.dinb(n311),.dout(n314),.clk(gclk));
	jand g258(.dina(w_n296_0[0]),.dinb(w_n314_0[1]),.dout(n315),.clk(gclk));
	jand g259(.dina(w_G370gat_1[0]),.dinb(w_G40gat_0[0]),.dout(n316),.clk(gclk));
	jor g260(.dina(w_n290_0[0]),.dinb(n316),.dout(n317),.clk(gclk));
	jand g261(.dina(w_n305_0[0]),.dinb(w_n317_0[2]),.dout(n318),.clk(gclk));
	jand g262(.dina(n318),.dinb(w_n314_0[0]),.dout(n319),.clk(gclk));
	jor g263(.dina(w_n319_0[1]),.dinb(w_n293_0[0]),.dout(n320),.clk(gclk));
	jor g264(.dina(n320),.dinb(w_dff_B_ZYoFFb5A6_1),.dout(G431gat),.clk(gclk));
	jand g265(.dina(w_G370gat_0[2]),.dinb(w_G92gat_0[0]),.dout(n322),.clk(gclk));
	jor g266(.dina(n322),.dinb(w_n254_0[0]),.dout(n323),.clk(gclk));
	jand g267(.dina(n323),.dinb(w_n313_0[0]),.dout(n324),.clk(gclk));
	jand g268(.dina(w_n303_0[0]),.dinb(w_n317_0[1]),.dout(n325),.clk(gclk));
	jand g269(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jand g270(.dina(w_n317_0[0]),.dinb(w_n283_0[0]),.dout(n327),.clk(gclk));
	jor g271(.dina(n327),.dinb(w_n286_0[0]),.dout(n328),.clk(gclk));
	jor g272(.dina(n328),.dinb(w_n319_0[0]),.dout(n329),.clk(gclk));
	jor g273(.dina(n329),.dinb(w_dff_B_KXmdAilH7_1),.dout(G432gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_kvUPm0Tm4_0),.doutb(w_dff_A_iqGXefEK4_1),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G4gat_0(.douta(w_dff_A_tpsFSx6J9_0),.doutb(w_G4gat_0[1]),.doutc(w_dff_A_7F2z2dxM4_2),.din(G4gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_zvrtZD2z1_0),.doutb(w_dff_A_gXl3cTPm5_1),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G11gat_0(.douta(w_dff_A_O2O27OSV9_0),.doutb(w_dff_A_6clacpgG8_1),.doutc(w_G11gat_0[2]),.din(G11gat));
	jspl3 jspl3_w_G14gat_0(.douta(w_dff_A_BwZsNusM9_0),.doutb(w_dff_A_hWRA1A9B9_1),.doutc(w_G14gat_0[2]),.din(G14gat));
	jspl3 jspl3_w_G17gat_0(.douta(w_dff_A_9XREv33Q7_0),.doutb(w_G17gat_0[1]),.doutc(w_dff_A_qtP09Y1i3_2),.din(G17gat));
	jspl3 jspl3_w_G21gat_0(.douta(w_G21gat_0[0]),.doutb(w_dff_A_AnuNYbET2_1),.doutc(w_dff_A_EqMDbWfC8_2),.din(G21gat));
	jspl jspl_w_G21gat_1(.douta(w_dff_A_0xg2965M0_0),.doutb(w_G21gat_1[1]),.din(w_G21gat_0[0]));
	jspl jspl_w_G24gat_0(.douta(w_dff_A_7Aba9wMw0_0),.doutb(w_G24gat_0[1]),.din(G24gat));
	jspl jspl_w_G27gat_0(.douta(w_dff_A_sHjkFqOj0_0),.doutb(w_G27gat_0[1]),.din(G27gat));
	jspl jspl_w_G30gat_0(.douta(w_G30gat_0[0]),.doutb(w_dff_A_UcNEqn591_1),.din(G30gat));
	jspl3 jspl3_w_G34gat_0(.douta(w_dff_A_GoDra4tL5_0),.doutb(w_G34gat_0[1]),.doutc(w_dff_A_SSDLaLU77_2),.din(G34gat));
	jspl3 jspl3_w_G37gat_0(.douta(w_dff_A_HnbCd5xA0_0),.doutb(w_dff_A_v7PrjEij8_1),.doutc(w_G37gat_0[2]),.din(G37gat));
	jspl jspl_w_G40gat_0(.douta(w_dff_A_qj6x9u1f2_0),.doutb(w_G40gat_0[1]),.din(G40gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_G43gat_0[0]),.doutb(w_dff_A_aCVhvqVc9_1),.doutc(w_dff_A_SsxNEVmU4_2),.din(G43gat));
	jspl jspl_w_G43gat_1(.douta(w_G43gat_1[0]),.doutb(w_dff_A_CMzcZLjl3_1),.din(w_G43gat_0[0]));
	jspl jspl_w_G47gat_0(.douta(w_dff_A_vB3sY1hH0_0),.doutb(w_G47gat_0[1]),.din(G47gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_dff_A_eWfgcqh78_0),.doutb(w_dff_A_RlI2Qcna3_1),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl jspl_w_G53gat_0(.douta(w_dff_A_MZFWZ5Ck2_0),.doutb(w_G53gat_0[1]),.din(G53gat));
	jspl3 jspl3_w_G56gat_0(.douta(w_dff_A_5Rl7pigT2_0),.doutb(w_G56gat_0[1]),.doutc(w_dff_A_ZzxpXh6n8_2),.din(G56gat));
	jspl3 jspl3_w_G60gat_0(.douta(w_dff_A_XVlost7X3_0),.doutb(w_dff_A_MIEOTvSw8_1),.doutc(w_G60gat_0[2]),.din(G60gat));
	jspl3 jspl3_w_G63gat_0(.douta(w_dff_A_JVwcaE8v5_0),.doutb(w_dff_A_SyCFXrVg8_1),.doutc(w_G63gat_0[2]),.din(G63gat));
	jspl jspl_w_G66gat_0(.douta(w_dff_A_bLe8H6p09_0),.doutb(w_G66gat_0[1]),.din(G66gat));
	jspl3 jspl3_w_G69gat_0(.douta(w_dff_A_MerAvAjZ2_0),.doutb(w_G69gat_0[1]),.doutc(w_dff_A_feB0LyTG2_2),.din(G69gat));
	jspl3 jspl3_w_G73gat_0(.douta(w_dff_A_5IvxTNcM1_0),.doutb(w_dff_A_BvsG1iB14_1),.doutc(w_G73gat_0[2]),.din(G73gat));
	jspl jspl_w_G76gat_0(.douta(w_dff_A_5BVq9ZHi3_0),.doutb(w_G76gat_0[1]),.din(G76gat));
	jspl jspl_w_G79gat_0(.douta(w_dff_A_bGOh0Hws8_0),.doutb(w_G79gat_0[1]),.din(G79gat));
	jspl3 jspl3_w_G82gat_0(.douta(w_G82gat_0[0]),.doutb(w_dff_A_x4t2TTDM3_1),.doutc(w_dff_A_Tptql5QN1_2),.din(G82gat));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_dff_A_hYqOcECy2_1),.doutc(w_dff_A_odwdWGJj5_2),.din(G86gat));
	jspl jspl_w_G86gat_1(.douta(w_dff_A_KxUoyAUl5_0),.doutb(w_G86gat_1[1]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G89gat_0(.douta(w_dff_A_tsCGXlx34_0),.doutb(w_dff_A_Q3mVMiD52_1),.doutc(w_G89gat_0[2]),.din(G89gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_oHno2wmd6_0),.doutb(w_dff_A_lkCDXcSL2_1),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G95gat_0(.douta(w_dff_A_zUeWR0hQ4_0),.doutb(w_G95gat_0[1]),.doutc(w_dff_A_RLzJUKcF1_2),.din(G95gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_Iv4WggU41_0),.doutb(w_dff_A_zFpJtcqW2_1),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl3 jspl3_w_G102gat_0(.douta(w_dff_A_yqszvjhP7_0),.doutb(w_dff_A_fZAokQjO4_1),.doutc(w_G102gat_0[2]),.din(G102gat));
	jspl jspl_w_G105gat_0(.douta(w_G105gat_0[0]),.doutb(w_dff_A_QH0Pbqzg0_1),.din(G105gat));
	jspl3 jspl3_w_G108gat_0(.douta(w_dff_A_8oZTMSvm4_0),.doutb(w_G108gat_0[1]),.doutc(w_dff_A_PSQlRAdH8_2),.din(G108gat));
	jspl3 jspl3_w_G112gat_0(.douta(w_dff_A_pegk6xgq3_0),.doutb(w_dff_A_zZ0sUR6U8_1),.doutc(w_G112gat_0[2]),.din(G112gat));
	jspl jspl_w_G115gat_0(.douta(w_dff_A_wsHHMeLw7_0),.doutb(w_G115gat_0[1]),.din(G115gat));
	jspl3 jspl3_w_G223gat_0(.douta(w_G223gat_0[0]),.doutb(w_G223gat_0[1]),.doutc(w_G223gat_0[2]),.din(G223gat_fa_));
	jspl3 jspl3_w_G223gat_1(.douta(w_G223gat_1[0]),.doutb(w_G223gat_1[1]),.doutc(w_G223gat_1[2]),.din(w_G223gat_0[0]));
	jspl3 jspl3_w_G223gat_2(.douta(w_G223gat_2[0]),.doutb(w_G223gat_2[1]),.doutc(w_G223gat_2[2]),.din(w_G223gat_0[1]));
	jspl3 jspl3_w_G223gat_3(.douta(w_G223gat_3[0]),.doutb(w_G223gat_3[1]),.doutc(w_dff_A_4UWrYcH12_2),.din(w_G223gat_0[2]));
	jspl3 jspl3_w_G329gat_0(.douta(w_G329gat_0[0]),.doutb(w_G329gat_0[1]),.doutc(w_G329gat_0[2]),.din(G329gat_fa_));
	jspl3 jspl3_w_G329gat_1(.douta(w_G329gat_1[0]),.doutb(w_G329gat_1[1]),.doutc(w_G329gat_1[2]),.din(w_G329gat_0[0]));
	jspl3 jspl3_w_G329gat_2(.douta(w_G329gat_2[0]),.doutb(w_G329gat_2[1]),.doutc(w_G329gat_2[2]),.din(w_G329gat_0[1]));
	jspl3 jspl3_w_G329gat_3(.douta(w_G329gat_3[0]),.doutb(w_G329gat_3[1]),.doutc(w_G329gat_3[2]),.din(w_G329gat_0[2]));
	jspl3 jspl3_w_G329gat_4(.douta(w_G329gat_4[0]),.doutb(w_G329gat_4[1]),.doutc(w_G329gat_4[2]),.din(w_G329gat_1[0]));
	jspl3 jspl3_w_G329gat_5(.douta(w_G329gat_5[0]),.doutb(w_G329gat_5[1]),.doutc(w_G329gat_5[2]),.din(w_G329gat_1[1]));
	jspl jspl_w_G329gat_6(.douta(w_G329gat_6),.doutb(w_dff_A_G75mAGmL5_1),.din(w_G329gat_1[2]));
	jspl3 jspl3_w_G370gat_0(.douta(w_G370gat_0[0]),.doutb(w_G370gat_0[1]),.doutc(w_G370gat_0[2]),.din(G370gat_fa_));
	jspl3 jspl3_w_G370gat_1(.douta(w_G370gat_1[0]),.doutb(w_G370gat_1[1]),.doutc(w_G370gat_1[2]),.din(w_G370gat_0[0]));
	jspl jspl_w_G370gat_2(.douta(w_G370gat_2),.doutb(w_dff_A_JCVWIwh73_1),.din(w_G370gat_0[1]));
	jspl jspl_w_G430gat_0(.douta(w_G430gat_0),.doutb(w_dff_A_xghxYD4R6_1),.din(G430gat_fa_));
	jspl jspl_w_n43_0(.douta(w_dff_A_28XZIk1f5_0),.doutb(w_n43_0[1]),.din(n43));
	jspl jspl_w_n44_0(.douta(w_n44_0[0]),.doutb(w_dff_A_ZYe2mqew6_1),.din(n44));
	jspl jspl_w_n47_0(.douta(w_dff_A_8u08u7938_0),.doutb(w_n47_0[1]),.din(n47));
	jspl jspl_w_n52_0(.douta(w_dff_A_HzQF8z6P4_0),.doutb(w_n52_0[1]),.din(n52));
	jspl jspl_w_n53_0(.douta(w_dff_A_Y6Is4uHB3_0),.doutb(w_n53_0[1]),.din(n53));
	jspl jspl_w_n56_0(.douta(w_dff_A_MoIFUcYl8_0),.doutb(w_n56_0[1]),.din(n56));
	jspl jspl_w_n58_0(.douta(w_dff_A_oqonIYtI2_0),.doutb(w_n58_0[1]),.din(n58));
	jspl jspl_w_n61_0(.douta(w_dff_A_zAKZk9uM8_0),.doutb(w_n61_0[1]),.din(n61));
	jspl jspl_w_n63_0(.douta(w_dff_A_GkI62Qcc3_0),.doutb(w_n63_0[1]),.din(n63));
	jspl jspl_w_n69_0(.douta(w_dff_A_LwcZ7WBl8_0),.doutb(w_n69_0[1]),.din(w_dff_B_6Fxb3ivR9_2));
	jspl jspl_w_n71_0(.douta(w_dff_A_7jIEFFPy1_0),.doutb(w_n71_0[1]),.din(n71));
	jspl jspl_w_n72_0(.douta(w_dff_A_sDxS30GO9_0),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n73_0(.douta(w_dff_A_S8vp1hBI6_0),.doutb(w_n73_0[1]),.din(n73));
	jspl jspl_w_n77_0(.douta(w_dff_A_e5q9SpBs2_0),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_dff_A_LcucVDKL2_0),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n79_0(.douta(w_dff_A_6hUcOWcz2_0),.doutb(w_n79_0[1]),.din(n79));
	jspl jspl_w_n82_0(.douta(w_dff_A_2L284IBN8_0),.doutb(w_n82_0[1]),.din(n82));
	jspl jspl_w_n84_0(.douta(w_dff_A_jRPjoRYT8_0),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n87_0(.douta(w_dff_A_xxSMbtcd9_0),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_dff_A_pb3yzhzd3_0),.doutb(w_n89_0[1]),.din(n89));
	jspl3 jspl3_w_n94_0(.douta(w_n94_0[0]),.doutb(w_n94_0[1]),.doutc(w_n94_0[2]),.din(n94));
	jspl3 jspl3_w_n94_1(.douta(w_n94_1[0]),.doutb(w_n94_1[1]),.doutc(w_n94_1[2]),.din(w_n94_0[0]));
	jspl3 jspl3_w_n94_2(.douta(w_n94_2[0]),.doutb(w_n94_2[1]),.doutc(w_n94_2[2]),.din(w_n94_0[1]));
	jspl3 jspl3_w_n94_3(.douta(w_n94_3[0]),.doutb(w_n94_3[1]),.doutc(w_n94_3[2]),.din(w_n94_0[2]));
	jspl jspl_w_n94_4(.douta(w_n94_4[0]),.doutb(w_n94_4[1]),.din(w_n94_1[0]));
	jspl jspl_w_n96_0(.douta(w_dff_A_NfiY4DDd3_0),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n98_0(.douta(w_dff_A_bCX2syvd0_0),.doutb(w_n98_0[1]),.din(w_dff_B_BizbFXHl3_2));
	jspl jspl_w_n100_0(.douta(w_dff_A_xqRTKSaT0_0),.doutb(w_n100_0[1]),.din(n100));
	jspl jspl_w_n107_0(.douta(w_dff_A_SSyHuhK77_0),.doutb(w_n107_0[1]),.din(w_dff_B_h679x01V9_2));
	jspl jspl_w_n109_0(.douta(w_dff_A_We3bCPNw9_0),.doutb(w_n109_0[1]),.din(n109));
	jspl3 jspl3_w_n114_0(.douta(w_dff_A_M8D3VRA67_0),.doutb(w_n114_0[1]),.doutc(w_n114_0[2]),.din(n114));
	jspl jspl_w_n115_0(.douta(w_dff_A_31Pa4CSX5_0),.doutb(w_n115_0[1]),.din(n115));
	jspl jspl_w_n119_0(.douta(w_n119_0[0]),.doutb(w_n119_0[1]),.din(n119));
	jspl jspl_w_n121_0(.douta(w_n121_0[0]),.doutb(w_n121_0[1]),.din(n121));
	jspl jspl_w_n123_0(.douta(w_n123_0[0]),.doutb(w_dff_A_iqB8XFrz2_1),.din(n123));
	jspl3 jspl3_w_n126_0(.douta(w_dff_A_kN9ZTeBs8_0),.doutb(w_dff_A_fpMbBfaE7_1),.doutc(w_n126_0[2]),.din(w_dff_B_EJOsXWCr7_3));
	jspl jspl_w_n128_0(.douta(w_dff_A_AEVTHE0x9_0),.doutb(w_n128_0[1]),.din(n128));
	jspl3 jspl3_w_n130_0(.douta(w_dff_A_x8N6BIx90_0),.doutb(w_dff_A_6J44yqVi5_1),.doutc(w_n130_0[2]),.din(w_dff_B_LBdoCohI3_3));
	jspl jspl_w_n132_0(.douta(w_dff_A_hu9pQrxC8_0),.doutb(w_n132_0[1]),.din(n132));
	jspl jspl_w_n139_0(.douta(w_n139_0[0]),.doutb(w_dff_A_C2h2upGr0_1),.din(n139));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n142_0(.douta(w_dff_A_KX1ModdX8_0),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n145_0(.douta(w_dff_A_XDhjYOjs0_0),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n146_0(.douta(w_n146_0[0]),.doutb(w_dff_A_xmlZg3DD4_1),.din(n146));
	jspl jspl_w_n147_0(.douta(w_n147_0[0]),.doutb(w_n147_0[1]),.din(n147));
	jspl jspl_w_n150_0(.douta(w_dff_A_nSTVCGDl6_0),.doutb(w_n150_0[1]),.din(w_dff_B_TIm7nUM62_2));
	jspl jspl_w_n151_0(.douta(w_n151_0[0]),.doutb(w_dff_A_T0s3z3sR2_1),.din(n151));
	jspl jspl_w_n154_0(.douta(w_dff_A_nVOQsG7n6_0),.doutb(w_n154_0[1]),.din(w_dff_B_rH6yLkox9_2));
	jspl jspl_w_n156_0(.douta(w_dff_A_ksqqvc4Z1_0),.doutb(w_n156_0[1]),.din(n156));
	jspl jspl_w_n159_0(.douta(w_dff_A_tPc41txx8_0),.doutb(w_n159_0[1]),.din(n159));
	jspl jspl_w_n164_0(.douta(w_dff_A_5lglyCVg7_0),.doutb(w_n164_0[1]),.din(n164));
	jspl jspl_w_n170_0(.douta(w_dff_A_qNwu4S5v0_0),.doutb(w_n170_0[1]),.din(w_dff_B_jGV4q4nI8_2));
	jspl jspl_w_n174_0(.douta(w_dff_A_Py0C3wr08_0),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n177_0(.douta(w_dff_A_F4mDHL5g2_0),.doutb(w_n177_0[1]),.din(n177));
	jspl3 jspl3_w_n182_0(.douta(w_n182_0[0]),.doutb(w_n182_0[1]),.doutc(w_n182_0[2]),.din(n182));
	jspl3 jspl3_w_n182_1(.douta(w_n182_1[0]),.doutb(w_n182_1[1]),.doutc(w_n182_1[2]),.din(w_n182_0[0]));
	jspl3 jspl3_w_n182_2(.douta(w_n182_2[0]),.doutb(w_n182_2[1]),.doutc(w_n182_2[2]),.din(w_n182_0[1]));
	jspl jspl_w_n182_3(.douta(w_n182_3[0]),.doutb(w_n182_3[1]),.din(w_n182_0[2]));
	jspl jspl_w_n184_0(.douta(w_dff_A_3vhBMoxG3_0),.doutb(w_n184_0[1]),.din(n184));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n191_0(.douta(w_dff_A_rf9Ws4F31_0),.doutb(w_n191_0[1]),.din(n191));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_dff_A_JQ4u0kL94_1),.din(n193));
	jspl jspl_w_n197_0(.douta(w_dff_A_DLXQ7I4y1_0),.doutb(w_n197_0[1]),.din(n197));
	jspl jspl_w_n198_0(.douta(w_dff_A_rx3r58Z40_0),.doutb(w_n198_0[1]),.din(w_dff_B_ENr5jcRP1_2));
	jspl jspl_w_n204_0(.douta(w_dff_A_1rCSSxDP9_0),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n205_0(.douta(w_dff_A_AnMNFDxc1_0),.doutb(w_n205_0[1]),.din(w_dff_B_5aEeEyyC1_2));
	jspl jspl_w_n217_0(.douta(w_dff_A_dtfYF0RU7_0),.doutb(w_n217_0[1]),.din(w_dff_B_0SRp5Z4h3_2));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_dff_A_LrTmRjb59_1),.din(n219));
	jspl jspl_w_n222_0(.douta(w_dff_A_bbCfdq1r1_0),.doutb(w_n222_0[1]),.din(w_dff_B_dh5WGy4B5_2));
	jspl jspl_w_n224_0(.douta(w_dff_A_nnUpAHli6_0),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_dff_A_Dx6iqY3E7_1),.din(n231));
	jspl jspl_w_n254_0(.douta(w_dff_A_OzVYxTJp1_0),.doutb(w_n254_0[1]),.din(n254));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl3 jspl3_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.doutc(w_n271_0[2]),.din(n271));
	jspl3 jspl3_w_n271_1(.douta(w_n271_1[0]),.doutb(w_n271_1[1]),.doutc(w_n271_1[2]),.din(w_n271_0[0]));
	jspl3 jspl3_w_n271_2(.douta(w_n271_2[0]),.doutb(w_n271_2[1]),.doutc(w_n271_2[2]),.din(w_n271_0[1]));
	jspl jspl_w_n271_3(.douta(w_n271_3[0]),.doutb(w_n271_3[1]),.din(w_n271_0[2]));
	jspl jspl_w_n274_0(.douta(w_dff_A_WmmXD38Y6_0),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n281_0(.douta(w_dff_A_woeQ6xX11_0),.doutb(w_n281_0[1]),.din(n281));
	jspl jspl_w_n283_0(.douta(w_n283_0[0]),.doutb(w_n283_0[1]),.din(n283));
	jspl jspl_w_n286_0(.douta(w_dff_A_laMmicQ84_0),.doutb(w_n286_0[1]),.din(n286));
	jspl jspl_w_n290_0(.douta(w_dff_A_25w1lPMr9_0),.doutb(w_n290_0[1]),.din(n290));
	jspl jspl_w_n293_0(.douta(w_dff_A_X7vp4PL19_0),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n296_0(.douta(w_dff_A_pLfHtfeN2_0),.doutb(w_n296_0[1]),.din(n296));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(n305));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl jspl_w_n314_0(.douta(w_n314_0[0]),.doutb(w_n314_0[1]),.din(n314));
	jspl3 jspl3_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.doutc(w_n317_0[2]),.din(n317));
	jspl jspl_w_n319_0(.douta(w_n319_0[0]),.doutb(w_n319_0[1]),.din(n319));
	jdff dff_B_GSnDh2kE5_1(.din(n233),.dout(w_dff_B_GSnDh2kE5_1),.clk(gclk));
	jdff dff_B_hIduJqmc9_1(.din(w_dff_B_GSnDh2kE5_1),.dout(w_dff_B_hIduJqmc9_1),.clk(gclk));
	jdff dff_B_VIrjoWqg4_1(.din(w_dff_B_hIduJqmc9_1),.dout(w_dff_B_VIrjoWqg4_1),.clk(gclk));
	jdff dff_B_czkWL5uQ7_0(.din(n275),.dout(w_dff_B_czkWL5uQ7_0),.clk(gclk));
	jdff dff_B_jDyP1OjQ3_0(.din(w_dff_B_czkWL5uQ7_0),.dout(w_dff_B_jDyP1OjQ3_0),.clk(gclk));
	jdff dff_B_ariQ0ZvI5_0(.din(w_dff_B_jDyP1OjQ3_0),.dout(w_dff_B_ariQ0ZvI5_0),.clk(gclk));
	jdff dff_B_CyL4EsOq2_0(.din(w_dff_B_ariQ0ZvI5_0),.dout(w_dff_B_CyL4EsOq2_0),.clk(gclk));
	jdff dff_B_9zOLbmIy1_0(.din(w_dff_B_CyL4EsOq2_0),.dout(w_dff_B_9zOLbmIy1_0),.clk(gclk));
	jdff dff_B_ZYoFFb5A6_1(.din(n315),.dout(w_dff_B_ZYoFFb5A6_1),.clk(gclk));
	jdff dff_A_X7vp4PL19_0(.dout(w_n293_0[0]),.din(w_dff_A_X7vp4PL19_0),.clk(gclk));
	jdff dff_B_xLjl8rKw0_0(.din(n291),.dout(w_dff_B_xLjl8rKw0_0),.clk(gclk));
	jdff dff_B_Tx7d7DJC6_0(.din(w_dff_B_xLjl8rKw0_0),.dout(w_dff_B_Tx7d7DJC6_0),.clk(gclk));
	jdff dff_B_CSQEN4uL9_0(.din(w_dff_B_Tx7d7DJC6_0),.dout(w_dff_B_CSQEN4uL9_0),.clk(gclk));
	jdff dff_B_O8kTvuKD0_0(.din(w_dff_B_CSQEN4uL9_0),.dout(w_dff_B_O8kTvuKD0_0),.clk(gclk));
	jdff dff_B_dVyWw4fQ3_0(.din(w_dff_B_O8kTvuKD0_0),.dout(w_dff_B_dVyWw4fQ3_0),.clk(gclk));
	jdff dff_A_pLfHtfeN2_0(.dout(w_n296_0[0]),.din(w_dff_A_pLfHtfeN2_0),.clk(gclk));
	jdff dff_B_KXmdAilH7_1(.din(n326),.dout(w_dff_B_KXmdAilH7_1),.clk(gclk));
	jdff dff_B_zDDe9ktI8_0(.din(n282),.dout(w_dff_B_zDDe9ktI8_0),.clk(gclk));
	jdff dff_B_M7M6Hzdg9_0(.din(w_dff_B_zDDe9ktI8_0),.dout(w_dff_B_M7M6Hzdg9_0),.clk(gclk));
	jdff dff_B_hKUYCX0D1_0(.din(w_dff_B_M7M6Hzdg9_0),.dout(w_dff_B_hKUYCX0D1_0),.clk(gclk));
	jdff dff_B_KCxFHtaV2_0(.din(w_dff_B_hKUYCX0D1_0),.dout(w_dff_B_KCxFHtaV2_0),.clk(gclk));
	jdff dff_B_qxgHqkJt9_0(.din(w_dff_B_KCxFHtaV2_0),.dout(w_dff_B_qxgHqkJt9_0),.clk(gclk));
	jdff dff_A_laMmicQ84_0(.dout(w_n286_0[0]),.din(w_dff_A_laMmicQ84_0),.clk(gclk));
	jdff dff_A_HY9rZFi71_0(.dout(w_n274_0[0]),.din(w_dff_A_HY9rZFi71_0),.clk(gclk));
	jdff dff_A_WFT3tQ0g0_0(.dout(w_dff_A_HY9rZFi71_0),.din(w_dff_A_WFT3tQ0g0_0),.clk(gclk));
	jdff dff_A_FmfjjktR9_0(.dout(w_dff_A_WFT3tQ0g0_0),.din(w_dff_A_FmfjjktR9_0),.clk(gclk));
	jdff dff_A_y0kxChaU5_0(.dout(w_dff_A_FmfjjktR9_0),.din(w_dff_A_y0kxChaU5_0),.clk(gclk));
	jdff dff_A_ygXpwAxh3_0(.dout(w_dff_A_y0kxChaU5_0),.din(w_dff_A_ygXpwAxh3_0),.clk(gclk));
	jdff dff_A_WmmXD38Y6_0(.dout(w_dff_A_ygXpwAxh3_0),.din(w_dff_A_WmmXD38Y6_0),.clk(gclk));
	jdff dff_B_xHxGJ5Ny8_1(.din(n300),.dout(w_dff_B_xHxGJ5Ny8_1),.clk(gclk));
	jdff dff_B_oeQS6wIZ6_1(.din(w_dff_B_xHxGJ5Ny8_1),.dout(w_dff_B_oeQS6wIZ6_1),.clk(gclk));
	jdff dff_B_NnICCbs74_1(.din(w_dff_B_oeQS6wIZ6_1),.dout(w_dff_B_NnICCbs74_1),.clk(gclk));
	jdff dff_B_7mLxy2vQ7_1(.din(w_dff_B_NnICCbs74_1),.dout(w_dff_B_7mLxy2vQ7_1),.clk(gclk));
	jdff dff_B_kXbpKEBk3_1(.din(w_dff_B_7mLxy2vQ7_1),.dout(w_dff_B_kXbpKEBk3_1),.clk(gclk));
	jdff dff_B_OAL6iOP00_1(.din(n301),.dout(w_dff_B_OAL6iOP00_1),.clk(gclk));
	jdff dff_B_WVRZKLQ06_1(.din(w_dff_B_OAL6iOP00_1),.dout(w_dff_B_WVRZKLQ06_1),.clk(gclk));
	jdff dff_B_4lf6p1SM7_1(.din(w_dff_B_WVRZKLQ06_1),.dout(w_dff_B_4lf6p1SM7_1),.clk(gclk));
	jdff dff_B_vb4owMNK2_1(.din(w_dff_B_4lf6p1SM7_1),.dout(w_dff_B_vb4owMNK2_1),.clk(gclk));
	jdff dff_B_2gInBCgu9_1(.din(w_dff_B_vb4owMNK2_1),.dout(w_dff_B_2gInBCgu9_1),.clk(gclk));
	jdff dff_B_CGrQXk1L9_1(.din(w_dff_B_2gInBCgu9_1),.dout(w_dff_B_CGrQXk1L9_1),.clk(gclk));
	jdff dff_B_8vYHROXb7_1(.din(w_dff_B_CGrQXk1L9_1),.dout(w_dff_B_8vYHROXb7_1),.clk(gclk));
	jdff dff_B_D8sSyh4c1_1(.din(w_dff_B_8vYHROXb7_1),.dout(w_dff_B_D8sSyh4c1_1),.clk(gclk));
	jdff dff_B_7xphdRD70_1(.din(w_dff_B_D8sSyh4c1_1),.dout(w_dff_B_7xphdRD70_1),.clk(gclk));
	jdff dff_B_R88nFhvk8_1(.din(w_dff_B_7xphdRD70_1),.dout(w_dff_B_R88nFhvk8_1),.clk(gclk));
	jdff dff_B_F7c70FBE9_1(.din(w_dff_B_R88nFhvk8_1),.dout(w_dff_B_F7c70FBE9_1),.clk(gclk));
	jdff dff_B_CG7TzqnV4_1(.din(w_dff_B_F7c70FBE9_1),.dout(w_dff_B_CG7TzqnV4_1),.clk(gclk));
	jdff dff_B_TRhcUU752_1(.din(w_dff_B_CG7TzqnV4_1),.dout(w_dff_B_TRhcUU752_1),.clk(gclk));
	jdff dff_B_BHWgLUzc9_1(.din(w_dff_B_TRhcUU752_1),.dout(w_dff_B_BHWgLUzc9_1),.clk(gclk));
	jdff dff_B_qAxORBmV6_1(.din(w_dff_B_BHWgLUzc9_1),.dout(w_dff_B_qAxORBmV6_1),.clk(gclk));
	jdff dff_B_bl2fhLvS6_1(.din(w_dff_B_qAxORBmV6_1),.dout(w_dff_B_bl2fhLvS6_1),.clk(gclk));
	jdff dff_B_5D7c1szW3_1(.din(w_dff_B_bl2fhLvS6_1),.dout(w_dff_B_5D7c1szW3_1),.clk(gclk));
	jdff dff_B_6KNdW3L09_1(.din(w_dff_B_5D7c1szW3_1),.dout(w_dff_B_6KNdW3L09_1),.clk(gclk));
	jdff dff_B_3EXKWv7H2_1(.din(w_dff_B_6KNdW3L09_1),.dout(w_dff_B_3EXKWv7H2_1),.clk(gclk));
	jdff dff_B_BTec5vnc7_1(.din(n242),.dout(w_dff_B_BTec5vnc7_1),.clk(gclk));
	jdff dff_B_hWCdCurf8_1(.din(n252),.dout(w_dff_B_hWCdCurf8_1),.clk(gclk));
	jdff dff_B_TihVYKXx0_1(.din(n264),.dout(w_dff_B_TihVYKXx0_1),.clk(gclk));
	jdff dff_B_lVg0OwBZ2_0(.din(n262),.dout(w_dff_B_lVg0OwBZ2_0),.clk(gclk));
	jdff dff_B_mkjwvadh6_0(.din(w_dff_B_lVg0OwBZ2_0),.dout(w_dff_B_mkjwvadh6_0),.clk(gclk));
	jdff dff_B_fU6PONy31_0(.din(w_dff_B_mkjwvadh6_0),.dout(w_dff_B_fU6PONy31_0),.clk(gclk));
	jdff dff_A_WvE99bJX6_1(.dout(w_n231_0[1]),.din(w_dff_A_WvE99bJX6_1),.clk(gclk));
	jdff dff_A_6186ux1M5_1(.dout(w_dff_A_WvE99bJX6_1),.din(w_dff_A_6186ux1M5_1),.clk(gclk));
	jdff dff_A_WFd7z3iY9_1(.dout(w_dff_A_6186ux1M5_1),.din(w_dff_A_WFd7z3iY9_1),.clk(gclk));
	jdff dff_A_Y6qPYb1y9_1(.dout(w_dff_A_WFd7z3iY9_1),.din(w_dff_A_Y6qPYb1y9_1),.clk(gclk));
	jdff dff_A_eahucu861_1(.dout(w_dff_A_Y6qPYb1y9_1),.din(w_dff_A_eahucu861_1),.clk(gclk));
	jdff dff_A_Dx6iqY3E7_1(.dout(w_dff_A_eahucu861_1),.din(w_dff_A_Dx6iqY3E7_1),.clk(gclk));
	jdff dff_B_V16kZFy51_1(.din(n246),.dout(w_dff_B_V16kZFy51_1),.clk(gclk));
	jdff dff_B_LPZI1See8_0(.din(n244),.dout(w_dff_B_LPZI1See8_0),.clk(gclk));
	jdff dff_B_hcxHYc191_0(.din(w_dff_B_LPZI1See8_0),.dout(w_dff_B_hcxHYc191_0),.clk(gclk));
	jdff dff_B_6eoxg8OF6_0(.din(w_dff_B_hcxHYc191_0),.dout(w_dff_B_6eoxg8OF6_0),.clk(gclk));
	jdff dff_B_0TbexHT18_0(.din(w_dff_B_6eoxg8OF6_0),.dout(w_dff_B_0TbexHT18_0),.clk(gclk));
	jdff dff_B_FbCoXbMV1_0(.din(w_dff_B_0TbexHT18_0),.dout(w_dff_B_FbCoXbMV1_0),.clk(gclk));
	jdff dff_B_LVxx1fIm2_1(.din(n237),.dout(w_dff_B_LVxx1fIm2_1),.clk(gclk));
	jdff dff_B_22sCyIcv4_0(.din(n235),.dout(w_dff_B_22sCyIcv4_0),.clk(gclk));
	jdff dff_B_ARh6LNE23_0(.din(w_dff_B_22sCyIcv4_0),.dout(w_dff_B_ARh6LNE23_0),.clk(gclk));
	jdff dff_B_PmwhMaNd7_0(.din(w_dff_B_ARh6LNE23_0),.dout(w_dff_B_PmwhMaNd7_0),.clk(gclk));
	jdff dff_B_4WmcnZt15_0(.din(w_dff_B_PmwhMaNd7_0),.dout(w_dff_B_4WmcnZt15_0),.clk(gclk));
	jdff dff_A_iG3ii5kw4_0(.dout(w_n290_0[0]),.din(w_dff_A_iG3ii5kw4_0),.clk(gclk));
	jdff dff_A_LVk07qnr8_0(.dout(w_dff_A_iG3ii5kw4_0),.din(w_dff_A_LVk07qnr8_0),.clk(gclk));
	jdff dff_A_fqjjwXgZ7_0(.dout(w_dff_A_LVk07qnr8_0),.din(w_dff_A_fqjjwXgZ7_0),.clk(gclk));
	jdff dff_A_SaJ3X7Bv2_0(.dout(w_dff_A_fqjjwXgZ7_0),.din(w_dff_A_SaJ3X7Bv2_0),.clk(gclk));
	jdff dff_A_Hacp7Wwv0_0(.dout(w_dff_A_SaJ3X7Bv2_0),.din(w_dff_A_Hacp7Wwv0_0),.clk(gclk));
	jdff dff_A_25w1lPMr9_0(.dout(w_dff_A_Hacp7Wwv0_0),.din(w_dff_A_25w1lPMr9_0),.clk(gclk));
	jdff dff_A_VcVnZbwv6_0(.dout(w_n254_0[0]),.din(w_dff_A_VcVnZbwv6_0),.clk(gclk));
	jdff dff_A_OAWoaVVb9_0(.dout(w_dff_A_VcVnZbwv6_0),.din(w_dff_A_OAWoaVVb9_0),.clk(gclk));
	jdff dff_A_XiFcFEo62_0(.dout(w_dff_A_OAWoaVVb9_0),.din(w_dff_A_XiFcFEo62_0),.clk(gclk));
	jdff dff_A_8TQkw6lt7_0(.dout(w_dff_A_XiFcFEo62_0),.din(w_dff_A_8TQkw6lt7_0),.clk(gclk));
	jdff dff_A_HGwRYJUM1_0(.dout(w_dff_A_8TQkw6lt7_0),.din(w_dff_A_HGwRYJUM1_0),.clk(gclk));
	jdff dff_A_OzVYxTJp1_0(.dout(w_dff_A_HGwRYJUM1_0),.din(w_dff_A_OzVYxTJp1_0),.clk(gclk));
	jdff dff_A_fnqeUtC94_0(.dout(w_n281_0[0]),.din(w_dff_A_fnqeUtC94_0),.clk(gclk));
	jdff dff_A_F02wDE6p8_0(.dout(w_dff_A_fnqeUtC94_0),.din(w_dff_A_F02wDE6p8_0),.clk(gclk));
	jdff dff_A_DWFINrfc8_0(.dout(w_dff_A_F02wDE6p8_0),.din(w_dff_A_DWFINrfc8_0),.clk(gclk));
	jdff dff_A_3xb3bOl61_0(.dout(w_dff_A_DWFINrfc8_0),.din(w_dff_A_3xb3bOl61_0),.clk(gclk));
	jdff dff_A_tUq7FhWe6_0(.dout(w_dff_A_3xb3bOl61_0),.din(w_dff_A_tUq7FhWe6_0),.clk(gclk));
	jdff dff_A_woeQ6xX11_0(.dout(w_dff_A_tUq7FhWe6_0),.din(w_dff_A_woeQ6xX11_0),.clk(gclk));
	jdff dff_B_VMJWkdGw0_0(.din(n280),.dout(w_dff_B_VMJWkdGw0_0),.clk(gclk));
	jdff dff_B_xwAI8yyP8_0(.din(w_dff_B_VMJWkdGw0_0),.dout(w_dff_B_xwAI8yyP8_0),.clk(gclk));
	jdff dff_B_GIKci5Mb3_0(.din(w_dff_B_xwAI8yyP8_0),.dout(w_dff_B_GIKci5Mb3_0),.clk(gclk));
	jdff dff_B_feggU7DD0_0(.din(w_dff_B_GIKci5Mb3_0),.dout(w_dff_B_feggU7DD0_0),.clk(gclk));
	jdff dff_B_YH9V6D4u8_0(.din(w_dff_B_feggU7DD0_0),.dout(w_dff_B_YH9V6D4u8_0),.clk(gclk));
	jdff dff_B_qkWew6ny7_0(.din(w_dff_B_YH9V6D4u8_0),.dout(w_dff_B_qkWew6ny7_0),.clk(gclk));
	jdff dff_B_ELQB5Iqi7_1(.din(n187),.dout(w_dff_B_ELQB5Iqi7_1),.clk(gclk));
	jdff dff_B_GNSqXq4E6_1(.din(n202),.dout(w_dff_B_GNSqXq4E6_1),.clk(gclk));
	jdff dff_B_kIK7VG9F5_1(.din(n221),.dout(w_dff_B_kIK7VG9F5_1),.clk(gclk));
	jdff dff_A_8kvUfK8O1_0(.dout(w_n224_0[0]),.din(w_dff_A_8kvUfK8O1_0),.clk(gclk));
	jdff dff_A_3MYg9Swm8_0(.dout(w_dff_A_8kvUfK8O1_0),.din(w_dff_A_3MYg9Swm8_0),.clk(gclk));
	jdff dff_A_4dlXNgHr5_0(.dout(w_dff_A_3MYg9Swm8_0),.din(w_dff_A_4dlXNgHr5_0),.clk(gclk));
	jdff dff_A_9KT6QPQ52_0(.dout(w_dff_A_4dlXNgHr5_0),.din(w_dff_A_9KT6QPQ52_0),.clk(gclk));
	jdff dff_A_UH48UZ7X9_0(.dout(w_dff_A_9KT6QPQ52_0),.din(w_dff_A_UH48UZ7X9_0),.clk(gclk));
	jdff dff_A_nnUpAHli6_0(.dout(w_dff_A_UH48UZ7X9_0),.din(w_dff_A_nnUpAHli6_0),.clk(gclk));
	jdff dff_A_yBpJdM7k4_0(.dout(w_n222_0[0]),.din(w_dff_A_yBpJdM7k4_0),.clk(gclk));
	jdff dff_A_5bTae3JN6_0(.dout(w_dff_A_yBpJdM7k4_0),.din(w_dff_A_5bTae3JN6_0),.clk(gclk));
	jdff dff_A_5P8rL2ZA6_0(.dout(w_dff_A_5bTae3JN6_0),.din(w_dff_A_5P8rL2ZA6_0),.clk(gclk));
	jdff dff_A_O1jOcvJz0_0(.dout(w_dff_A_5P8rL2ZA6_0),.din(w_dff_A_O1jOcvJz0_0),.clk(gclk));
	jdff dff_A_bbCfdq1r1_0(.dout(w_dff_A_O1jOcvJz0_0),.din(w_dff_A_bbCfdq1r1_0),.clk(gclk));
	jdff dff_B_YdMERaM50_2(.din(n222),.dout(w_dff_B_YdMERaM50_2),.clk(gclk));
	jdff dff_B_hyyEkbhs8_2(.din(w_dff_B_YdMERaM50_2),.dout(w_dff_B_hyyEkbhs8_2),.clk(gclk));
	jdff dff_B_IbWdedKo0_2(.din(w_dff_B_hyyEkbhs8_2),.dout(w_dff_B_IbWdedKo0_2),.clk(gclk));
	jdff dff_B_5VLEpwHo0_2(.din(w_dff_B_IbWdedKo0_2),.dout(w_dff_B_5VLEpwHo0_2),.clk(gclk));
	jdff dff_B_pLgYB2pj5_2(.din(w_dff_B_5VLEpwHo0_2),.dout(w_dff_B_pLgYB2pj5_2),.clk(gclk));
	jdff dff_B_lOdqvsgp8_2(.din(w_dff_B_pLgYB2pj5_2),.dout(w_dff_B_lOdqvsgp8_2),.clk(gclk));
	jdff dff_B_l3RuFBV89_2(.din(w_dff_B_lOdqvsgp8_2),.dout(w_dff_B_l3RuFBV89_2),.clk(gclk));
	jdff dff_B_emhezZSf9_2(.din(w_dff_B_l3RuFBV89_2),.dout(w_dff_B_emhezZSf9_2),.clk(gclk));
	jdff dff_B_w3EksEOO7_2(.din(w_dff_B_emhezZSf9_2),.dout(w_dff_B_w3EksEOO7_2),.clk(gclk));
	jdff dff_B_893WKOa32_2(.din(w_dff_B_w3EksEOO7_2),.dout(w_dff_B_893WKOa32_2),.clk(gclk));
	jdff dff_B_DTj59Uvb3_2(.din(w_dff_B_893WKOa32_2),.dout(w_dff_B_DTj59Uvb3_2),.clk(gclk));
	jdff dff_B_IzSdSrrA8_2(.din(w_dff_B_DTj59Uvb3_2),.dout(w_dff_B_IzSdSrrA8_2),.clk(gclk));
	jdff dff_B_wdvUVKDo0_2(.din(w_dff_B_IzSdSrrA8_2),.dout(w_dff_B_wdvUVKDo0_2),.clk(gclk));
	jdff dff_B_dh5WGy4B5_2(.din(w_dff_B_wdvUVKDo0_2),.dout(w_dff_B_dh5WGy4B5_2),.clk(gclk));
	jdff dff_A_fsA8EV2t2_0(.dout(w_G115gat_0[0]),.din(w_dff_A_fsA8EV2t2_0),.clk(gclk));
	jdff dff_A_xAxsMlXv2_0(.dout(w_dff_A_fsA8EV2t2_0),.din(w_dff_A_xAxsMlXv2_0),.clk(gclk));
	jdff dff_A_E53njXCd2_0(.dout(w_dff_A_xAxsMlXv2_0),.din(w_dff_A_E53njXCd2_0),.clk(gclk));
	jdff dff_A_hmwwARnM2_0(.dout(w_dff_A_E53njXCd2_0),.din(w_dff_A_hmwwARnM2_0),.clk(gclk));
	jdff dff_A_oqJHtDKu0_0(.dout(w_dff_A_hmwwARnM2_0),.din(w_dff_A_oqJHtDKu0_0),.clk(gclk));
	jdff dff_A_GNYaiNh17_0(.dout(w_dff_A_oqJHtDKu0_0),.din(w_dff_A_GNYaiNh17_0),.clk(gclk));
	jdff dff_A_Vl5vsEAq2_0(.dout(w_dff_A_GNYaiNh17_0),.din(w_dff_A_Vl5vsEAq2_0),.clk(gclk));
	jdff dff_A_ZYa2puiv2_0(.dout(w_dff_A_Vl5vsEAq2_0),.din(w_dff_A_ZYa2puiv2_0),.clk(gclk));
	jdff dff_A_wX3Rw1q02_0(.dout(w_dff_A_ZYa2puiv2_0),.din(w_dff_A_wX3Rw1q02_0),.clk(gclk));
	jdff dff_A_iN0dAAPp8_0(.dout(w_dff_A_wX3Rw1q02_0),.din(w_dff_A_iN0dAAPp8_0),.clk(gclk));
	jdff dff_A_KsCL86RT6_0(.dout(w_dff_A_iN0dAAPp8_0),.din(w_dff_A_KsCL86RT6_0),.clk(gclk));
	jdff dff_A_ZUdX4zNb4_0(.dout(w_dff_A_KsCL86RT6_0),.din(w_dff_A_ZUdX4zNb4_0),.clk(gclk));
	jdff dff_A_LYF8F3Tq2_0(.dout(w_dff_A_ZUdX4zNb4_0),.din(w_dff_A_LYF8F3Tq2_0),.clk(gclk));
	jdff dff_A_J2Mrws8M5_0(.dout(w_dff_A_LYF8F3Tq2_0),.din(w_dff_A_J2Mrws8M5_0),.clk(gclk));
	jdff dff_A_wsHHMeLw7_0(.dout(w_dff_A_J2Mrws8M5_0),.din(w_dff_A_wsHHMeLw7_0),.clk(gclk));
	jdff dff_A_lYhGSCPn1_1(.dout(w_n219_0[1]),.din(w_dff_A_lYhGSCPn1_1),.clk(gclk));
	jdff dff_A_czWZKsfc9_1(.dout(w_dff_A_lYhGSCPn1_1),.din(w_dff_A_czWZKsfc9_1),.clk(gclk));
	jdff dff_A_VSHXhCJc9_1(.dout(w_dff_A_czWZKsfc9_1),.din(w_dff_A_VSHXhCJc9_1),.clk(gclk));
	jdff dff_A_LrTmRjb59_1(.dout(w_dff_A_VSHXhCJc9_1),.din(w_dff_A_LrTmRjb59_1),.clk(gclk));
	jdff dff_A_wjoC0toR2_0(.dout(w_n217_0[0]),.din(w_dff_A_wjoC0toR2_0),.clk(gclk));
	jdff dff_A_vCs445nJ1_0(.dout(w_dff_A_wjoC0toR2_0),.din(w_dff_A_vCs445nJ1_0),.clk(gclk));
	jdff dff_A_2tlBKJnU7_0(.dout(w_dff_A_vCs445nJ1_0),.din(w_dff_A_2tlBKJnU7_0),.clk(gclk));
	jdff dff_A_AZWId6Kt7_0(.dout(w_dff_A_2tlBKJnU7_0),.din(w_dff_A_AZWId6Kt7_0),.clk(gclk));
	jdff dff_A_n8vm7ZZn3_0(.dout(w_dff_A_AZWId6Kt7_0),.din(w_dff_A_n8vm7ZZn3_0),.clk(gclk));
	jdff dff_A_diPwbLcV5_0(.dout(w_dff_A_n8vm7ZZn3_0),.din(w_dff_A_diPwbLcV5_0),.clk(gclk));
	jdff dff_A_BwgELZkZ3_0(.dout(w_dff_A_diPwbLcV5_0),.din(w_dff_A_BwgELZkZ3_0),.clk(gclk));
	jdff dff_A_7m5WlaoD7_0(.dout(w_dff_A_BwgELZkZ3_0),.din(w_dff_A_7m5WlaoD7_0),.clk(gclk));
	jdff dff_A_OxYC5Mqn7_0(.dout(w_dff_A_7m5WlaoD7_0),.din(w_dff_A_OxYC5Mqn7_0),.clk(gclk));
	jdff dff_A_DpZ2unM60_0(.dout(w_dff_A_OxYC5Mqn7_0),.din(w_dff_A_DpZ2unM60_0),.clk(gclk));
	jdff dff_A_dtfYF0RU7_0(.dout(w_dff_A_DpZ2unM60_0),.din(w_dff_A_dtfYF0RU7_0),.clk(gclk));
	jdff dff_B_jd4f72az7_2(.din(n217),.dout(w_dff_B_jd4f72az7_2),.clk(gclk));
	jdff dff_B_EIZ92mA41_2(.din(w_dff_B_jd4f72az7_2),.dout(w_dff_B_EIZ92mA41_2),.clk(gclk));
	jdff dff_B_l7kZjTXc2_2(.din(w_dff_B_EIZ92mA41_2),.dout(w_dff_B_l7kZjTXc2_2),.clk(gclk));
	jdff dff_B_GZupzVj27_2(.din(w_dff_B_l7kZjTXc2_2),.dout(w_dff_B_GZupzVj27_2),.clk(gclk));
	jdff dff_B_RWLohaRm7_2(.din(w_dff_B_GZupzVj27_2),.dout(w_dff_B_RWLohaRm7_2),.clk(gclk));
	jdff dff_B_dV5i4kRd6_2(.din(w_dff_B_RWLohaRm7_2),.dout(w_dff_B_dV5i4kRd6_2),.clk(gclk));
	jdff dff_B_K43EhjD71_2(.din(w_dff_B_dV5i4kRd6_2),.dout(w_dff_B_K43EhjD71_2),.clk(gclk));
	jdff dff_B_0SRp5Z4h3_2(.din(w_dff_B_K43EhjD71_2),.dout(w_dff_B_0SRp5Z4h3_2),.clk(gclk));
	jdff dff_A_URwKWAYp2_0(.dout(w_G40gat_0[0]),.din(w_dff_A_URwKWAYp2_0),.clk(gclk));
	jdff dff_A_votMDdNu4_0(.dout(w_dff_A_URwKWAYp2_0),.din(w_dff_A_votMDdNu4_0),.clk(gclk));
	jdff dff_A_fHso0OEe1_0(.dout(w_dff_A_votMDdNu4_0),.din(w_dff_A_fHso0OEe1_0),.clk(gclk));
	jdff dff_A_zjKeFhqd0_0(.dout(w_dff_A_fHso0OEe1_0),.din(w_dff_A_zjKeFhqd0_0),.clk(gclk));
	jdff dff_A_LpluJNeK5_0(.dout(w_dff_A_zjKeFhqd0_0),.din(w_dff_A_LpluJNeK5_0),.clk(gclk));
	jdff dff_A_9Yk93ou95_0(.dout(w_dff_A_LpluJNeK5_0),.din(w_dff_A_9Yk93ou95_0),.clk(gclk));
	jdff dff_A_KNtLhHRG3_0(.dout(w_dff_A_9Yk93ou95_0),.din(w_dff_A_KNtLhHRG3_0),.clk(gclk));
	jdff dff_A_pOyopasy9_0(.dout(w_dff_A_KNtLhHRG3_0),.din(w_dff_A_pOyopasy9_0),.clk(gclk));
	jdff dff_A_qyTZFZPK2_0(.dout(w_dff_A_pOyopasy9_0),.din(w_dff_A_qyTZFZPK2_0),.clk(gclk));
	jdff dff_A_kU381YMW7_0(.dout(w_dff_A_qyTZFZPK2_0),.din(w_dff_A_kU381YMW7_0),.clk(gclk));
	jdff dff_A_ulUXXly06_0(.dout(w_dff_A_kU381YMW7_0),.din(w_dff_A_ulUXXly06_0),.clk(gclk));
	jdff dff_A_omUMCf9u4_0(.dout(w_dff_A_ulUXXly06_0),.din(w_dff_A_omUMCf9u4_0),.clk(gclk));
	jdff dff_A_VDk9UMgz3_0(.dout(w_dff_A_omUMCf9u4_0),.din(w_dff_A_VDk9UMgz3_0),.clk(gclk));
	jdff dff_A_cx0imB703_0(.dout(w_dff_A_VDk9UMgz3_0),.din(w_dff_A_cx0imB703_0),.clk(gclk));
	jdff dff_A_ZM9E6xcm8_0(.dout(w_dff_A_cx0imB703_0),.din(w_dff_A_ZM9E6xcm8_0),.clk(gclk));
	jdff dff_A_npdtz6Jy5_0(.dout(w_dff_A_ZM9E6xcm8_0),.din(w_dff_A_npdtz6Jy5_0),.clk(gclk));
	jdff dff_A_6lBG8Cnj6_0(.dout(w_dff_A_npdtz6Jy5_0),.din(w_dff_A_6lBG8Cnj6_0),.clk(gclk));
	jdff dff_A_tcQbky3R5_0(.dout(w_dff_A_6lBG8Cnj6_0),.din(w_dff_A_tcQbky3R5_0),.clk(gclk));
	jdff dff_A_kqU2lrcn5_0(.dout(w_dff_A_tcQbky3R5_0),.din(w_dff_A_kqU2lrcn5_0),.clk(gclk));
	jdff dff_A_qj6x9u1f2_0(.dout(w_dff_A_kqU2lrcn5_0),.din(w_dff_A_qj6x9u1f2_0),.clk(gclk));
	jdff dff_B_q00PK1XG6_1(.din(n214),.dout(w_dff_B_q00PK1XG6_1),.clk(gclk));
	jdff dff_B_2XCdmvSp5_1(.din(w_dff_B_q00PK1XG6_1),.dout(w_dff_B_2XCdmvSp5_1),.clk(gclk));
	jdff dff_B_P1ZSg6HP7_1(.din(w_dff_B_2XCdmvSp5_1),.dout(w_dff_B_P1ZSg6HP7_1),.clk(gclk));
	jdff dff_B_DVirL3oD2_1(.din(w_dff_B_P1ZSg6HP7_1),.dout(w_dff_B_DVirL3oD2_1),.clk(gclk));
	jdff dff_B_icyLWSGx8_1(.din(w_dff_B_DVirL3oD2_1),.dout(w_dff_B_icyLWSGx8_1),.clk(gclk));
	jdff dff_B_pnbZDh8S3_1(.din(w_dff_B_icyLWSGx8_1),.dout(w_dff_B_pnbZDh8S3_1),.clk(gclk));
	jdff dff_B_7Y4ud1yb0_1(.din(w_dff_B_pnbZDh8S3_1),.dout(w_dff_B_7Y4ud1yb0_1),.clk(gclk));
	jdff dff_B_eooJ9GeX6_1(.din(w_dff_B_7Y4ud1yb0_1),.dout(w_dff_B_eooJ9GeX6_1),.clk(gclk));
	jdff dff_B_wjniNUKX8_1(.din(w_dff_B_eooJ9GeX6_1),.dout(w_dff_B_wjniNUKX8_1),.clk(gclk));
	jdff dff_B_9jjsctm77_1(.din(w_dff_B_wjniNUKX8_1),.dout(w_dff_B_9jjsctm77_1),.clk(gclk));
	jdff dff_B_ctyO2yCT4_1(.din(w_dff_B_9jjsctm77_1),.dout(w_dff_B_ctyO2yCT4_1),.clk(gclk));
	jdff dff_B_mecfc78R8_1(.din(w_dff_B_ctyO2yCT4_1),.dout(w_dff_B_mecfc78R8_1),.clk(gclk));
	jdff dff_B_4c3VtT6s0_1(.din(n209),.dout(w_dff_B_4c3VtT6s0_1),.clk(gclk));
	jdff dff_B_QQXSPl696_1(.din(w_dff_B_4c3VtT6s0_1),.dout(w_dff_B_QQXSPl696_1),.clk(gclk));
	jdff dff_B_lnQyGsTN2_1(.din(w_dff_B_QQXSPl696_1),.dout(w_dff_B_lnQyGsTN2_1),.clk(gclk));
	jdff dff_B_QhQFr7YL9_1(.din(w_dff_B_lnQyGsTN2_1),.dout(w_dff_B_QhQFr7YL9_1),.clk(gclk));
	jdff dff_B_YOMH6s239_1(.din(w_dff_B_QhQFr7YL9_1),.dout(w_dff_B_YOMH6s239_1),.clk(gclk));
	jdff dff_B_cmgcXGgN4_1(.din(w_dff_B_YOMH6s239_1),.dout(w_dff_B_cmgcXGgN4_1),.clk(gclk));
	jdff dff_B_Rh90SVv32_1(.din(w_dff_B_cmgcXGgN4_1),.dout(w_dff_B_Rh90SVv32_1),.clk(gclk));
	jdff dff_B_w71gb5y77_1(.din(w_dff_B_Rh90SVv32_1),.dout(w_dff_B_w71gb5y77_1),.clk(gclk));
	jdff dff_B_kZagx7jQ8_1(.din(w_dff_B_w71gb5y77_1),.dout(w_dff_B_kZagx7jQ8_1),.clk(gclk));
	jdff dff_B_KSNTyxvV8_1(.din(w_dff_B_kZagx7jQ8_1),.dout(w_dff_B_KSNTyxvV8_1),.clk(gclk));
	jdff dff_B_5NdIs9Ps6_1(.din(w_dff_B_KSNTyxvV8_1),.dout(w_dff_B_5NdIs9Ps6_1),.clk(gclk));
	jdff dff_B_FQ33IYN68_1(.din(w_dff_B_5NdIs9Ps6_1),.dout(w_dff_B_FQ33IYN68_1),.clk(gclk));
	jdff dff_B_RecGgbmW2_1(.din(w_dff_B_FQ33IYN68_1),.dout(w_dff_B_RecGgbmW2_1),.clk(gclk));
	jdff dff_B_h2WQfTe00_1(.din(w_dff_B_RecGgbmW2_1),.dout(w_dff_B_h2WQfTe00_1),.clk(gclk));
	jdff dff_A_KooFJ4an7_0(.dout(w_G14gat_0[0]),.din(w_dff_A_KooFJ4an7_0),.clk(gclk));
	jdff dff_A_5N7W4bjW9_0(.dout(w_dff_A_KooFJ4an7_0),.din(w_dff_A_5N7W4bjW9_0),.clk(gclk));
	jdff dff_A_91kb09bN8_0(.dout(w_dff_A_5N7W4bjW9_0),.din(w_dff_A_91kb09bN8_0),.clk(gclk));
	jdff dff_A_9zRlLWAA1_0(.dout(w_dff_A_91kb09bN8_0),.din(w_dff_A_9zRlLWAA1_0),.clk(gclk));
	jdff dff_A_VBn9TSq39_0(.dout(w_dff_A_9zRlLWAA1_0),.din(w_dff_A_VBn9TSq39_0),.clk(gclk));
	jdff dff_A_sAgWO94h0_0(.dout(w_dff_A_VBn9TSq39_0),.din(w_dff_A_sAgWO94h0_0),.clk(gclk));
	jdff dff_A_LxoOkUmX6_0(.dout(w_dff_A_sAgWO94h0_0),.din(w_dff_A_LxoOkUmX6_0),.clk(gclk));
	jdff dff_A_OHesSGDi1_0(.dout(w_dff_A_LxoOkUmX6_0),.din(w_dff_A_OHesSGDi1_0),.clk(gclk));
	jdff dff_A_IHbETiyJ4_0(.dout(w_dff_A_OHesSGDi1_0),.din(w_dff_A_IHbETiyJ4_0),.clk(gclk));
	jdff dff_A_OwwoBDjW0_0(.dout(w_dff_A_IHbETiyJ4_0),.din(w_dff_A_OwwoBDjW0_0),.clk(gclk));
	jdff dff_A_pK24mIv30_0(.dout(w_dff_A_OwwoBDjW0_0),.din(w_dff_A_pK24mIv30_0),.clk(gclk));
	jdff dff_A_F4WaHt2f5_0(.dout(w_dff_A_pK24mIv30_0),.din(w_dff_A_F4WaHt2f5_0),.clk(gclk));
	jdff dff_A_azx97wwe4_0(.dout(w_dff_A_F4WaHt2f5_0),.din(w_dff_A_azx97wwe4_0),.clk(gclk));
	jdff dff_A_3uDSStZo0_0(.dout(w_dff_A_azx97wwe4_0),.din(w_dff_A_3uDSStZo0_0),.clk(gclk));
	jdff dff_A_BwZsNusM9_0(.dout(w_dff_A_3uDSStZo0_0),.din(w_dff_A_BwZsNusM9_0),.clk(gclk));
	jdff dff_A_LQUvEn4p5_1(.dout(w_G14gat_0[1]),.din(w_dff_A_LQUvEn4p5_1),.clk(gclk));
	jdff dff_A_Flwu4zfB4_1(.dout(w_dff_A_LQUvEn4p5_1),.din(w_dff_A_Flwu4zfB4_1),.clk(gclk));
	jdff dff_A_1IPTWx4j2_1(.dout(w_dff_A_Flwu4zfB4_1),.din(w_dff_A_1IPTWx4j2_1),.clk(gclk));
	jdff dff_A_QUVyFi4h8_1(.dout(w_dff_A_1IPTWx4j2_1),.din(w_dff_A_QUVyFi4h8_1),.clk(gclk));
	jdff dff_A_vfLG6VhC8_1(.dout(w_dff_A_QUVyFi4h8_1),.din(w_dff_A_vfLG6VhC8_1),.clk(gclk));
	jdff dff_A_0vzcR0Mt6_1(.dout(w_dff_A_vfLG6VhC8_1),.din(w_dff_A_0vzcR0Mt6_1),.clk(gclk));
	jdff dff_A_Gq0jnUpT2_1(.dout(w_dff_A_0vzcR0Mt6_1),.din(w_dff_A_Gq0jnUpT2_1),.clk(gclk));
	jdff dff_A_FMMIp7qE6_1(.dout(w_dff_A_Gq0jnUpT2_1),.din(w_dff_A_FMMIp7qE6_1),.clk(gclk));
	jdff dff_A_WeFkpDEY9_1(.dout(w_dff_A_FMMIp7qE6_1),.din(w_dff_A_WeFkpDEY9_1),.clk(gclk));
	jdff dff_A_rfHQNtAG0_1(.dout(w_dff_A_WeFkpDEY9_1),.din(w_dff_A_rfHQNtAG0_1),.clk(gclk));
	jdff dff_A_o1svPETJ0_1(.dout(w_dff_A_rfHQNtAG0_1),.din(w_dff_A_o1svPETJ0_1),.clk(gclk));
	jdff dff_A_PvHJiViS7_1(.dout(w_dff_A_o1svPETJ0_1),.din(w_dff_A_PvHJiViS7_1),.clk(gclk));
	jdff dff_A_987klsKH6_1(.dout(w_dff_A_PvHJiViS7_1),.din(w_dff_A_987klsKH6_1),.clk(gclk));
	jdff dff_A_1sdopjId2_1(.dout(w_dff_A_987klsKH6_1),.din(w_dff_A_1sdopjId2_1),.clk(gclk));
	jdff dff_A_FYEbGyxv4_1(.dout(w_dff_A_1sdopjId2_1),.din(w_dff_A_FYEbGyxv4_1),.clk(gclk));
	jdff dff_A_G9ueQvwZ2_1(.dout(w_dff_A_FYEbGyxv4_1),.din(w_dff_A_G9ueQvwZ2_1),.clk(gclk));
	jdff dff_A_BwAiN2Wa3_1(.dout(w_dff_A_G9ueQvwZ2_1),.din(w_dff_A_BwAiN2Wa3_1),.clk(gclk));
	jdff dff_A_kMxDCVIs9_1(.dout(w_dff_A_BwAiN2Wa3_1),.din(w_dff_A_kMxDCVIs9_1),.clk(gclk));
	jdff dff_A_u8P8Po8w2_1(.dout(w_dff_A_kMxDCVIs9_1),.din(w_dff_A_u8P8Po8w2_1),.clk(gclk));
	jdff dff_A_hWRA1A9B9_1(.dout(w_dff_A_u8P8Po8w2_1),.din(w_dff_A_hWRA1A9B9_1),.clk(gclk));
	jdff dff_A_LfEhZHl00_0(.dout(w_n205_0[0]),.din(w_dff_A_LfEhZHl00_0),.clk(gclk));
	jdff dff_A_rkwCWqyX9_0(.dout(w_dff_A_LfEhZHl00_0),.din(w_dff_A_rkwCWqyX9_0),.clk(gclk));
	jdff dff_A_Ob0nhDB07_0(.dout(w_dff_A_rkwCWqyX9_0),.din(w_dff_A_Ob0nhDB07_0),.clk(gclk));
	jdff dff_A_uhjLAQNN4_0(.dout(w_dff_A_Ob0nhDB07_0),.din(w_dff_A_uhjLAQNN4_0),.clk(gclk));
	jdff dff_A_6JNcqD5U0_0(.dout(w_dff_A_uhjLAQNN4_0),.din(w_dff_A_6JNcqD5U0_0),.clk(gclk));
	jdff dff_A_AnMNFDxc1_0(.dout(w_dff_A_6JNcqD5U0_0),.din(w_dff_A_AnMNFDxc1_0),.clk(gclk));
	jdff dff_B_fOJxWYgY7_2(.din(n205),.dout(w_dff_B_fOJxWYgY7_2),.clk(gclk));
	jdff dff_B_GHIbASPS3_2(.din(w_dff_B_fOJxWYgY7_2),.dout(w_dff_B_GHIbASPS3_2),.clk(gclk));
	jdff dff_B_zc54HsMS0_2(.din(w_dff_B_GHIbASPS3_2),.dout(w_dff_B_zc54HsMS0_2),.clk(gclk));
	jdff dff_B_tPqFifj69_2(.din(w_dff_B_zc54HsMS0_2),.dout(w_dff_B_tPqFifj69_2),.clk(gclk));
	jdff dff_B_Gije76v97_2(.din(w_dff_B_tPqFifj69_2),.dout(w_dff_B_Gije76v97_2),.clk(gclk));
	jdff dff_B_iWMwpXHh0_2(.din(w_dff_B_Gije76v97_2),.dout(w_dff_B_iWMwpXHh0_2),.clk(gclk));
	jdff dff_B_Au4HEF214_2(.din(w_dff_B_iWMwpXHh0_2),.dout(w_dff_B_Au4HEF214_2),.clk(gclk));
	jdff dff_B_OH6Bf5Fu2_2(.din(w_dff_B_Au4HEF214_2),.dout(w_dff_B_OH6Bf5Fu2_2),.clk(gclk));
	jdff dff_B_tpMnQwPb0_2(.din(w_dff_B_OH6Bf5Fu2_2),.dout(w_dff_B_tpMnQwPb0_2),.clk(gclk));
	jdff dff_B_kNuWFeCk3_2(.din(w_dff_B_tpMnQwPb0_2),.dout(w_dff_B_kNuWFeCk3_2),.clk(gclk));
	jdff dff_B_wOkYWYKD3_2(.din(w_dff_B_kNuWFeCk3_2),.dout(w_dff_B_wOkYWYKD3_2),.clk(gclk));
	jdff dff_B_UIrplxaR9_2(.din(w_dff_B_wOkYWYKD3_2),.dout(w_dff_B_UIrplxaR9_2),.clk(gclk));
	jdff dff_B_5aEeEyyC1_2(.din(w_dff_B_UIrplxaR9_2),.dout(w_dff_B_5aEeEyyC1_2),.clk(gclk));
	jdff dff_A_Tq2maAmm5_0(.dout(w_G92gat_0[0]),.din(w_dff_A_Tq2maAmm5_0),.clk(gclk));
	jdff dff_A_8ikQTadE7_0(.dout(w_dff_A_Tq2maAmm5_0),.din(w_dff_A_8ikQTadE7_0),.clk(gclk));
	jdff dff_A_9IzPf7lX3_0(.dout(w_dff_A_8ikQTadE7_0),.din(w_dff_A_9IzPf7lX3_0),.clk(gclk));
	jdff dff_A_vm3CM9Dw8_0(.dout(w_dff_A_9IzPf7lX3_0),.din(w_dff_A_vm3CM9Dw8_0),.clk(gclk));
	jdff dff_A_8fxOPCtD5_0(.dout(w_dff_A_vm3CM9Dw8_0),.din(w_dff_A_8fxOPCtD5_0),.clk(gclk));
	jdff dff_A_6sxMqMEl1_0(.dout(w_dff_A_8fxOPCtD5_0),.din(w_dff_A_6sxMqMEl1_0),.clk(gclk));
	jdff dff_A_Wo8TfAuY9_0(.dout(w_dff_A_6sxMqMEl1_0),.din(w_dff_A_Wo8TfAuY9_0),.clk(gclk));
	jdff dff_A_5Nc2Jxhl3_0(.dout(w_dff_A_Wo8TfAuY9_0),.din(w_dff_A_5Nc2Jxhl3_0),.clk(gclk));
	jdff dff_A_1iLwwVWs3_0(.dout(w_dff_A_5Nc2Jxhl3_0),.din(w_dff_A_1iLwwVWs3_0),.clk(gclk));
	jdff dff_A_ZezFM1pL8_0(.dout(w_dff_A_1iLwwVWs3_0),.din(w_dff_A_ZezFM1pL8_0),.clk(gclk));
	jdff dff_A_q0wH6vH95_0(.dout(w_dff_A_ZezFM1pL8_0),.din(w_dff_A_q0wH6vH95_0),.clk(gclk));
	jdff dff_A_3ufiBksR7_0(.dout(w_dff_A_q0wH6vH95_0),.din(w_dff_A_3ufiBksR7_0),.clk(gclk));
	jdff dff_A_hBCqrYvd4_0(.dout(w_dff_A_3ufiBksR7_0),.din(w_dff_A_hBCqrYvd4_0),.clk(gclk));
	jdff dff_A_hJibkNQl2_0(.dout(w_dff_A_hBCqrYvd4_0),.din(w_dff_A_hJibkNQl2_0),.clk(gclk));
	jdff dff_A_YuMJNmG72_0(.dout(w_dff_A_hJibkNQl2_0),.din(w_dff_A_YuMJNmG72_0),.clk(gclk));
	jdff dff_A_RK2Z40uw0_0(.dout(w_dff_A_YuMJNmG72_0),.din(w_dff_A_RK2Z40uw0_0),.clk(gclk));
	jdff dff_A_88AAHG1I5_0(.dout(w_dff_A_RK2Z40uw0_0),.din(w_dff_A_88AAHG1I5_0),.clk(gclk));
	jdff dff_A_O16qnquD2_0(.dout(w_dff_A_88AAHG1I5_0),.din(w_dff_A_O16qnquD2_0),.clk(gclk));
	jdff dff_A_oleWOq7v0_0(.dout(w_dff_A_O16qnquD2_0),.din(w_dff_A_oleWOq7v0_0),.clk(gclk));
	jdff dff_A_oHno2wmd6_0(.dout(w_dff_A_oleWOq7v0_0),.din(w_dff_A_oHno2wmd6_0),.clk(gclk));
	jdff dff_A_Z4wBsNYM7_1(.dout(w_G92gat_0[1]),.din(w_dff_A_Z4wBsNYM7_1),.clk(gclk));
	jdff dff_A_36T123zN7_1(.dout(w_dff_A_Z4wBsNYM7_1),.din(w_dff_A_36T123zN7_1),.clk(gclk));
	jdff dff_A_bYShhjUX9_1(.dout(w_dff_A_36T123zN7_1),.din(w_dff_A_bYShhjUX9_1),.clk(gclk));
	jdff dff_A_JUcWfsqX4_1(.dout(w_dff_A_bYShhjUX9_1),.din(w_dff_A_JUcWfsqX4_1),.clk(gclk));
	jdff dff_A_j6Kppt9l3_1(.dout(w_dff_A_JUcWfsqX4_1),.din(w_dff_A_j6Kppt9l3_1),.clk(gclk));
	jdff dff_A_D90zdTLE8_1(.dout(w_dff_A_j6Kppt9l3_1),.din(w_dff_A_D90zdTLE8_1),.clk(gclk));
	jdff dff_A_bHObf2ni8_1(.dout(w_dff_A_D90zdTLE8_1),.din(w_dff_A_bHObf2ni8_1),.clk(gclk));
	jdff dff_A_OlluYn5z3_1(.dout(w_dff_A_bHObf2ni8_1),.din(w_dff_A_OlluYn5z3_1),.clk(gclk));
	jdff dff_A_VKrgORKB5_1(.dout(w_dff_A_OlluYn5z3_1),.din(w_dff_A_VKrgORKB5_1),.clk(gclk));
	jdff dff_A_kuw4pHGu3_1(.dout(w_dff_A_VKrgORKB5_1),.din(w_dff_A_kuw4pHGu3_1),.clk(gclk));
	jdff dff_A_P23sgYsc5_1(.dout(w_dff_A_kuw4pHGu3_1),.din(w_dff_A_P23sgYsc5_1),.clk(gclk));
	jdff dff_A_RdhsWqx99_1(.dout(w_dff_A_P23sgYsc5_1),.din(w_dff_A_RdhsWqx99_1),.clk(gclk));
	jdff dff_A_05VLVG5v7_1(.dout(w_dff_A_RdhsWqx99_1),.din(w_dff_A_05VLVG5v7_1),.clk(gclk));
	jdff dff_A_lkCDXcSL2_1(.dout(w_dff_A_05VLVG5v7_1),.din(w_dff_A_lkCDXcSL2_1),.clk(gclk));
	jdff dff_A_pCCO09rF5_0(.dout(w_n204_0[0]),.din(w_dff_A_pCCO09rF5_0),.clk(gclk));
	jdff dff_A_RD0QYzFV6_0(.dout(w_dff_A_pCCO09rF5_0),.din(w_dff_A_RD0QYzFV6_0),.clk(gclk));
	jdff dff_A_pwWVTRRs6_0(.dout(w_dff_A_RD0QYzFV6_0),.din(w_dff_A_pwWVTRRs6_0),.clk(gclk));
	jdff dff_A_oRu1ITMv9_0(.dout(w_dff_A_pwWVTRRs6_0),.din(w_dff_A_oRu1ITMv9_0),.clk(gclk));
	jdff dff_A_xvnooeX77_0(.dout(w_dff_A_oRu1ITMv9_0),.din(w_dff_A_xvnooeX77_0),.clk(gclk));
	jdff dff_A_1rCSSxDP9_0(.dout(w_dff_A_xvnooeX77_0),.din(w_dff_A_1rCSSxDP9_0),.clk(gclk));
	jdff dff_A_s1FhOk1n5_0(.dout(w_n198_0[0]),.din(w_dff_A_s1FhOk1n5_0),.clk(gclk));
	jdff dff_A_gheSqkuk8_0(.dout(w_dff_A_s1FhOk1n5_0),.din(w_dff_A_gheSqkuk8_0),.clk(gclk));
	jdff dff_A_hjY6aPR09_0(.dout(w_dff_A_gheSqkuk8_0),.din(w_dff_A_hjY6aPR09_0),.clk(gclk));
	jdff dff_A_Ul5kchh18_0(.dout(w_dff_A_hjY6aPR09_0),.din(w_dff_A_Ul5kchh18_0),.clk(gclk));
	jdff dff_A_oTahqyhp2_0(.dout(w_dff_A_Ul5kchh18_0),.din(w_dff_A_oTahqyhp2_0),.clk(gclk));
	jdff dff_A_rx3r58Z40_0(.dout(w_dff_A_oTahqyhp2_0),.din(w_dff_A_rx3r58Z40_0),.clk(gclk));
	jdff dff_B_Vf4E7VPh3_2(.din(n198),.dout(w_dff_B_Vf4E7VPh3_2),.clk(gclk));
	jdff dff_B_Oc6o3v8z1_2(.din(w_dff_B_Vf4E7VPh3_2),.dout(w_dff_B_Oc6o3v8z1_2),.clk(gclk));
	jdff dff_B_SkNY9oMq8_2(.din(w_dff_B_Oc6o3v8z1_2),.dout(w_dff_B_SkNY9oMq8_2),.clk(gclk));
	jdff dff_B_mbruSknS9_2(.din(w_dff_B_SkNY9oMq8_2),.dout(w_dff_B_mbruSknS9_2),.clk(gclk));
	jdff dff_B_8dEEqOn31_2(.din(w_dff_B_mbruSknS9_2),.dout(w_dff_B_8dEEqOn31_2),.clk(gclk));
	jdff dff_B_tym5eEYv0_2(.din(w_dff_B_8dEEqOn31_2),.dout(w_dff_B_tym5eEYv0_2),.clk(gclk));
	jdff dff_B_1lIJKnEV1_2(.din(w_dff_B_tym5eEYv0_2),.dout(w_dff_B_1lIJKnEV1_2),.clk(gclk));
	jdff dff_B_KszUaK690_2(.din(w_dff_B_1lIJKnEV1_2),.dout(w_dff_B_KszUaK690_2),.clk(gclk));
	jdff dff_B_BX5srGLX9_2(.din(w_dff_B_KszUaK690_2),.dout(w_dff_B_BX5srGLX9_2),.clk(gclk));
	jdff dff_B_MpiPvr995_2(.din(w_dff_B_BX5srGLX9_2),.dout(w_dff_B_MpiPvr995_2),.clk(gclk));
	jdff dff_B_Kz4UMlW19_2(.din(w_dff_B_MpiPvr995_2),.dout(w_dff_B_Kz4UMlW19_2),.clk(gclk));
	jdff dff_B_7LaVMsGs4_2(.din(w_dff_B_Kz4UMlW19_2),.dout(w_dff_B_7LaVMsGs4_2),.clk(gclk));
	jdff dff_B_ENr5jcRP1_2(.din(w_dff_B_7LaVMsGs4_2),.dout(w_dff_B_ENr5jcRP1_2),.clk(gclk));
	jdff dff_A_cFr70PcO5_0(.dout(w_G27gat_0[0]),.din(w_dff_A_cFr70PcO5_0),.clk(gclk));
	jdff dff_A_Ej189avp4_0(.dout(w_dff_A_cFr70PcO5_0),.din(w_dff_A_Ej189avp4_0),.clk(gclk));
	jdff dff_A_yICjViVC5_0(.dout(w_dff_A_Ej189avp4_0),.din(w_dff_A_yICjViVC5_0),.clk(gclk));
	jdff dff_A_jItJKpUJ1_0(.dout(w_dff_A_yICjViVC5_0),.din(w_dff_A_jItJKpUJ1_0),.clk(gclk));
	jdff dff_A_uxhKUSVq1_0(.dout(w_dff_A_jItJKpUJ1_0),.din(w_dff_A_uxhKUSVq1_0),.clk(gclk));
	jdff dff_A_LqUj06CV4_0(.dout(w_dff_A_uxhKUSVq1_0),.din(w_dff_A_LqUj06CV4_0),.clk(gclk));
	jdff dff_A_eqSVw9832_0(.dout(w_dff_A_LqUj06CV4_0),.din(w_dff_A_eqSVw9832_0),.clk(gclk));
	jdff dff_A_WMeGJ6pz4_0(.dout(w_dff_A_eqSVw9832_0),.din(w_dff_A_WMeGJ6pz4_0),.clk(gclk));
	jdff dff_A_xTkKj4Pd9_0(.dout(w_dff_A_WMeGJ6pz4_0),.din(w_dff_A_xTkKj4Pd9_0),.clk(gclk));
	jdff dff_A_OQ5F2s9m1_0(.dout(w_dff_A_xTkKj4Pd9_0),.din(w_dff_A_OQ5F2s9m1_0),.clk(gclk));
	jdff dff_A_X2JtlG1n2_0(.dout(w_dff_A_OQ5F2s9m1_0),.din(w_dff_A_X2JtlG1n2_0),.clk(gclk));
	jdff dff_A_jgOcxwZ09_0(.dout(w_dff_A_X2JtlG1n2_0),.din(w_dff_A_jgOcxwZ09_0),.clk(gclk));
	jdff dff_A_MS968xZC4_0(.dout(w_dff_A_jgOcxwZ09_0),.din(w_dff_A_MS968xZC4_0),.clk(gclk));
	jdff dff_A_sHjkFqOj0_0(.dout(w_dff_A_MS968xZC4_0),.din(w_dff_A_sHjkFqOj0_0),.clk(gclk));
	jdff dff_A_haPGZmqi5_0(.dout(w_n197_0[0]),.din(w_dff_A_haPGZmqi5_0),.clk(gclk));
	jdff dff_A_idn5NWLt4_0(.dout(w_dff_A_haPGZmqi5_0),.din(w_dff_A_idn5NWLt4_0),.clk(gclk));
	jdff dff_A_GyWwAoU22_0(.dout(w_dff_A_idn5NWLt4_0),.din(w_dff_A_GyWwAoU22_0),.clk(gclk));
	jdff dff_A_d6NfiNZk9_0(.dout(w_dff_A_GyWwAoU22_0),.din(w_dff_A_d6NfiNZk9_0),.clk(gclk));
	jdff dff_A_nQjZMv2Z3_0(.dout(w_dff_A_d6NfiNZk9_0),.din(w_dff_A_nQjZMv2Z3_0),.clk(gclk));
	jdff dff_A_DLXQ7I4y1_0(.dout(w_dff_A_nQjZMv2Z3_0),.din(w_dff_A_DLXQ7I4y1_0),.clk(gclk));
	jdff dff_A_8fr7v03Q2_1(.dout(w_n193_0[1]),.din(w_dff_A_8fr7v03Q2_1),.clk(gclk));
	jdff dff_A_tbv4vpEC2_1(.dout(w_dff_A_8fr7v03Q2_1),.din(w_dff_A_tbv4vpEC2_1),.clk(gclk));
	jdff dff_A_wB53yctj1_1(.dout(w_dff_A_tbv4vpEC2_1),.din(w_dff_A_wB53yctj1_1),.clk(gclk));
	jdff dff_A_HDrtb0766_1(.dout(w_dff_A_wB53yctj1_1),.din(w_dff_A_HDrtb0766_1),.clk(gclk));
	jdff dff_A_FBjp5dQp3_1(.dout(w_dff_A_HDrtb0766_1),.din(w_dff_A_FBjp5dQp3_1),.clk(gclk));
	jdff dff_A_Twfgu76Y8_1(.dout(w_dff_A_FBjp5dQp3_1),.din(w_dff_A_Twfgu76Y8_1),.clk(gclk));
	jdff dff_A_JQ4u0kL94_1(.dout(w_dff_A_Twfgu76Y8_1),.din(w_dff_A_JQ4u0kL94_1),.clk(gclk));
	jdff dff_B_OtlWnwt38_0(.din(n192),.dout(w_dff_B_OtlWnwt38_0),.clk(gclk));
	jdff dff_B_bJlIOEmW7_0(.din(w_dff_B_OtlWnwt38_0),.dout(w_dff_B_bJlIOEmW7_0),.clk(gclk));
	jdff dff_B_Ub5k3Qmg1_0(.din(w_dff_B_bJlIOEmW7_0),.dout(w_dff_B_Ub5k3Qmg1_0),.clk(gclk));
	jdff dff_B_3PvvBRdj4_0(.din(w_dff_B_Ub5k3Qmg1_0),.dout(w_dff_B_3PvvBRdj4_0),.clk(gclk));
	jdff dff_B_29CtSvsd5_0(.din(w_dff_B_3PvvBRdj4_0),.dout(w_dff_B_29CtSvsd5_0),.clk(gclk));
	jdff dff_A_ei9AeArb4_0(.dout(w_n191_0[0]),.din(w_dff_A_ei9AeArb4_0),.clk(gclk));
	jdff dff_A_5Rn2GySe6_0(.dout(w_dff_A_ei9AeArb4_0),.din(w_dff_A_5Rn2GySe6_0),.clk(gclk));
	jdff dff_A_dPkZWSHH0_0(.dout(w_dff_A_5Rn2GySe6_0),.din(w_dff_A_dPkZWSHH0_0),.clk(gclk));
	jdff dff_A_jhpVUb811_0(.dout(w_dff_A_dPkZWSHH0_0),.din(w_dff_A_jhpVUb811_0),.clk(gclk));
	jdff dff_A_4loqmFTX5_0(.dout(w_dff_A_jhpVUb811_0),.din(w_dff_A_4loqmFTX5_0),.clk(gclk));
	jdff dff_A_BInmhQ7F2_0(.dout(w_dff_A_4loqmFTX5_0),.din(w_dff_A_BInmhQ7F2_0),.clk(gclk));
	jdff dff_A_8cweJVTL5_0(.dout(w_dff_A_BInmhQ7F2_0),.din(w_dff_A_8cweJVTL5_0),.clk(gclk));
	jdff dff_A_ViIO1gdv5_0(.dout(w_dff_A_8cweJVTL5_0),.din(w_dff_A_ViIO1gdv5_0),.clk(gclk));
	jdff dff_A_J7WFVJ3E4_0(.dout(w_dff_A_ViIO1gdv5_0),.din(w_dff_A_J7WFVJ3E4_0),.clk(gclk));
	jdff dff_A_CZl9vFKP7_0(.dout(w_dff_A_J7WFVJ3E4_0),.din(w_dff_A_CZl9vFKP7_0),.clk(gclk));
	jdff dff_A_mzRyPqYu8_0(.dout(w_dff_A_CZl9vFKP7_0),.din(w_dff_A_mzRyPqYu8_0),.clk(gclk));
	jdff dff_A_UkWEbEk67_0(.dout(w_dff_A_mzRyPqYu8_0),.din(w_dff_A_UkWEbEk67_0),.clk(gclk));
	jdff dff_A_jSimQT6m3_0(.dout(w_dff_A_UkWEbEk67_0),.din(w_dff_A_jSimQT6m3_0),.clk(gclk));
	jdff dff_A_C0jF9Z4a8_0(.dout(w_dff_A_jSimQT6m3_0),.din(w_dff_A_C0jF9Z4a8_0),.clk(gclk));
	jdff dff_A_BqdGOZ8i7_0(.dout(w_dff_A_C0jF9Z4a8_0),.din(w_dff_A_BqdGOZ8i7_0),.clk(gclk));
	jdff dff_A_rrp1YvzQ8_0(.dout(w_dff_A_BqdGOZ8i7_0),.din(w_dff_A_rrp1YvzQ8_0),.clk(gclk));
	jdff dff_A_iNJ3xtnk4_0(.dout(w_dff_A_rrp1YvzQ8_0),.din(w_dff_A_iNJ3xtnk4_0),.clk(gclk));
	jdff dff_A_nBgdbj7t8_0(.dout(w_dff_A_iNJ3xtnk4_0),.din(w_dff_A_nBgdbj7t8_0),.clk(gclk));
	jdff dff_A_rf9Ws4F31_0(.dout(w_dff_A_nBgdbj7t8_0),.din(w_dff_A_rf9Ws4F31_0),.clk(gclk));
	jdff dff_A_1ABIOUda5_0(.dout(w_G53gat_0[0]),.din(w_dff_A_1ABIOUda5_0),.clk(gclk));
	jdff dff_A_YOfJcjuf3_0(.dout(w_dff_A_1ABIOUda5_0),.din(w_dff_A_YOfJcjuf3_0),.clk(gclk));
	jdff dff_A_n8lNJukw4_0(.dout(w_dff_A_YOfJcjuf3_0),.din(w_dff_A_n8lNJukw4_0),.clk(gclk));
	jdff dff_A_g79ngoGE2_0(.dout(w_dff_A_n8lNJukw4_0),.din(w_dff_A_g79ngoGE2_0),.clk(gclk));
	jdff dff_A_TAB9VUeP6_0(.dout(w_dff_A_g79ngoGE2_0),.din(w_dff_A_TAB9VUeP6_0),.clk(gclk));
	jdff dff_A_gw1HYg6z4_0(.dout(w_dff_A_TAB9VUeP6_0),.din(w_dff_A_gw1HYg6z4_0),.clk(gclk));
	jdff dff_A_G7FaBxIB0_0(.dout(w_dff_A_gw1HYg6z4_0),.din(w_dff_A_G7FaBxIB0_0),.clk(gclk));
	jdff dff_A_tsgfsOQt0_0(.dout(w_dff_A_G7FaBxIB0_0),.din(w_dff_A_tsgfsOQt0_0),.clk(gclk));
	jdff dff_A_UX0JaKHb1_0(.dout(w_dff_A_tsgfsOQt0_0),.din(w_dff_A_UX0JaKHb1_0),.clk(gclk));
	jdff dff_A_DBwfIG8f6_0(.dout(w_dff_A_UX0JaKHb1_0),.din(w_dff_A_DBwfIG8f6_0),.clk(gclk));
	jdff dff_A_iXzoPtDu5_0(.dout(w_dff_A_DBwfIG8f6_0),.din(w_dff_A_iXzoPtDu5_0),.clk(gclk));
	jdff dff_A_Fks5oyfD1_0(.dout(w_dff_A_iXzoPtDu5_0),.din(w_dff_A_Fks5oyfD1_0),.clk(gclk));
	jdff dff_A_dMdFt7Q74_0(.dout(w_dff_A_Fks5oyfD1_0),.din(w_dff_A_dMdFt7Q74_0),.clk(gclk));
	jdff dff_A_MUo3cpeH9_0(.dout(w_dff_A_dMdFt7Q74_0),.din(w_dff_A_MUo3cpeH9_0),.clk(gclk));
	jdff dff_A_TaTnHh3p2_0(.dout(w_dff_A_MUo3cpeH9_0),.din(w_dff_A_TaTnHh3p2_0),.clk(gclk));
	jdff dff_A_HgvRYNAg7_0(.dout(w_dff_A_TaTnHh3p2_0),.din(w_dff_A_HgvRYNAg7_0),.clk(gclk));
	jdff dff_A_wbajDwLD2_0(.dout(w_dff_A_HgvRYNAg7_0),.din(w_dff_A_wbajDwLD2_0),.clk(gclk));
	jdff dff_A_611kaBzC1_0(.dout(w_dff_A_wbajDwLD2_0),.din(w_dff_A_611kaBzC1_0),.clk(gclk));
	jdff dff_A_gOuz1BdX3_0(.dout(w_dff_A_611kaBzC1_0),.din(w_dff_A_gOuz1BdX3_0),.clk(gclk));
	jdff dff_A_MZFWZ5Ck2_0(.dout(w_dff_A_gOuz1BdX3_0),.din(w_dff_A_MZFWZ5Ck2_0),.clk(gclk));
	jdff dff_A_lRBjIQnH6_0(.dout(w_n184_0[0]),.din(w_dff_A_lRBjIQnH6_0),.clk(gclk));
	jdff dff_A_aAR5BkXZ8_0(.dout(w_dff_A_lRBjIQnH6_0),.din(w_dff_A_aAR5BkXZ8_0),.clk(gclk));
	jdff dff_A_WbfoVMih3_0(.dout(w_dff_A_aAR5BkXZ8_0),.din(w_dff_A_WbfoVMih3_0),.clk(gclk));
	jdff dff_A_4odZ5Z5s2_0(.dout(w_dff_A_WbfoVMih3_0),.din(w_dff_A_4odZ5Z5s2_0),.clk(gclk));
	jdff dff_A_KQTkJy614_0(.dout(w_dff_A_4odZ5Z5s2_0),.din(w_dff_A_KQTkJy614_0),.clk(gclk));
	jdff dff_A_3vhBMoxG3_0(.dout(w_dff_A_KQTkJy614_0),.din(w_dff_A_3vhBMoxG3_0),.clk(gclk));
	jdff dff_B_7QJYiEzJ9_1(.din(n167),.dout(w_dff_B_7QJYiEzJ9_1),.clk(gclk));
	jdff dff_A_YSxIqE1F7_0(.dout(w_n177_0[0]),.din(w_dff_A_YSxIqE1F7_0),.clk(gclk));
	jdff dff_A_vHg0tNUU3_0(.dout(w_dff_A_YSxIqE1F7_0),.din(w_dff_A_vHg0tNUU3_0),.clk(gclk));
	jdff dff_A_bQfLeDv21_0(.dout(w_dff_A_vHg0tNUU3_0),.din(w_dff_A_bQfLeDv21_0),.clk(gclk));
	jdff dff_A_z5LF2SNo9_0(.dout(w_dff_A_bQfLeDv21_0),.din(w_dff_A_z5LF2SNo9_0),.clk(gclk));
	jdff dff_A_vtb5Xuwr3_0(.dout(w_dff_A_z5LF2SNo9_0),.din(w_dff_A_vtb5Xuwr3_0),.clk(gclk));
	jdff dff_A_F4mDHL5g2_0(.dout(w_dff_A_vtb5Xuwr3_0),.din(w_dff_A_F4mDHL5g2_0),.clk(gclk));
	jdff dff_A_hNoqOqaQ4_0(.dout(w_n174_0[0]),.din(w_dff_A_hNoqOqaQ4_0),.clk(gclk));
	jdff dff_A_phovm6tY2_0(.dout(w_dff_A_hNoqOqaQ4_0),.din(w_dff_A_phovm6tY2_0),.clk(gclk));
	jdff dff_A_hmlgpLnG1_0(.dout(w_dff_A_phovm6tY2_0),.din(w_dff_A_hmlgpLnG1_0),.clk(gclk));
	jdff dff_A_ZJowE0C39_0(.dout(w_dff_A_hmlgpLnG1_0),.din(w_dff_A_ZJowE0C39_0),.clk(gclk));
	jdff dff_A_pu9xypF90_0(.dout(w_dff_A_ZJowE0C39_0),.din(w_dff_A_pu9xypF90_0),.clk(gclk));
	jdff dff_A_Py0C3wr08_0(.dout(w_dff_A_pu9xypF90_0),.din(w_dff_A_Py0C3wr08_0),.clk(gclk));
	jdff dff_B_UErZ2wEc0_1(.din(n172),.dout(w_dff_B_UErZ2wEc0_1),.clk(gclk));
	jdff dff_B_Mu6LO9Ko9_1(.din(w_dff_B_UErZ2wEc0_1),.dout(w_dff_B_Mu6LO9Ko9_1),.clk(gclk));
	jdff dff_B_a4MScE0T5_1(.din(w_dff_B_Mu6LO9Ko9_1),.dout(w_dff_B_a4MScE0T5_1),.clk(gclk));
	jdff dff_B_P1PksuTA7_1(.din(w_dff_B_a4MScE0T5_1),.dout(w_dff_B_P1PksuTA7_1),.clk(gclk));
	jdff dff_B_dGfsQuAp3_1(.din(w_dff_B_P1PksuTA7_1),.dout(w_dff_B_dGfsQuAp3_1),.clk(gclk));
	jdff dff_B_etYSBqrZ6_1(.din(w_dff_B_dGfsQuAp3_1),.dout(w_dff_B_etYSBqrZ6_1),.clk(gclk));
	jdff dff_A_DNHgzYTT8_0(.dout(w_n170_0[0]),.din(w_dff_A_DNHgzYTT8_0),.clk(gclk));
	jdff dff_A_jdtgZKU72_0(.dout(w_dff_A_DNHgzYTT8_0),.din(w_dff_A_jdtgZKU72_0),.clk(gclk));
	jdff dff_A_g9dnEfBq9_0(.dout(w_dff_A_jdtgZKU72_0),.din(w_dff_A_g9dnEfBq9_0),.clk(gclk));
	jdff dff_A_qNwu4S5v0_0(.dout(w_dff_A_g9dnEfBq9_0),.din(w_dff_A_qNwu4S5v0_0),.clk(gclk));
	jdff dff_B_jGV4q4nI8_2(.din(n170),.dout(w_dff_B_jGV4q4nI8_2),.clk(gclk));
	jdff dff_B_FO9BZqkR4_0(.din(n169),.dout(w_dff_B_FO9BZqkR4_0),.clk(gclk));
	jdff dff_B_rKg1oiLt3_0(.din(w_dff_B_FO9BZqkR4_0),.dout(w_dff_B_rKg1oiLt3_0),.clk(gclk));
	jdff dff_B_00o5uWn50_0(.din(w_dff_B_rKg1oiLt3_0),.dout(w_dff_B_00o5uWn50_0),.clk(gclk));
	jdff dff_B_qd0v0rlh4_0(.din(w_dff_B_00o5uWn50_0),.dout(w_dff_B_qd0v0rlh4_0),.clk(gclk));
	jdff dff_A_l0xrVePn7_0(.dout(w_n164_0[0]),.din(w_dff_A_l0xrVePn7_0),.clk(gclk));
	jdff dff_A_Fn7lYF5u0_0(.dout(w_dff_A_l0xrVePn7_0),.din(w_dff_A_Fn7lYF5u0_0),.clk(gclk));
	jdff dff_A_XiqxT8H98_0(.dout(w_dff_A_Fn7lYF5u0_0),.din(w_dff_A_XiqxT8H98_0),.clk(gclk));
	jdff dff_A_W31yEjFY4_0(.dout(w_dff_A_XiqxT8H98_0),.din(w_dff_A_W31yEjFY4_0),.clk(gclk));
	jdff dff_A_SovL6pa74_0(.dout(w_dff_A_W31yEjFY4_0),.din(w_dff_A_SovL6pa74_0),.clk(gclk));
	jdff dff_A_5lglyCVg7_0(.dout(w_dff_A_SovL6pa74_0),.din(w_dff_A_5lglyCVg7_0),.clk(gclk));
	jdff dff_A_UOEAbDft5_0(.dout(w_n159_0[0]),.din(w_dff_A_UOEAbDft5_0),.clk(gclk));
	jdff dff_A_MaVyGzcw9_0(.dout(w_dff_A_UOEAbDft5_0),.din(w_dff_A_MaVyGzcw9_0),.clk(gclk));
	jdff dff_A_d7UN6i9q9_0(.dout(w_dff_A_MaVyGzcw9_0),.din(w_dff_A_d7UN6i9q9_0),.clk(gclk));
	jdff dff_A_2WFmqAyY2_0(.dout(w_dff_A_d7UN6i9q9_0),.din(w_dff_A_2WFmqAyY2_0),.clk(gclk));
	jdff dff_A_RdW3j2tg7_0(.dout(w_dff_A_2WFmqAyY2_0),.din(w_dff_A_RdW3j2tg7_0),.clk(gclk));
	jdff dff_A_tPc41txx8_0(.dout(w_dff_A_RdW3j2tg7_0),.din(w_dff_A_tPc41txx8_0),.clk(gclk));
	jdff dff_A_K0Q8vH814_0(.dout(w_n156_0[0]),.din(w_dff_A_K0Q8vH814_0),.clk(gclk));
	jdff dff_A_snZYENbb9_0(.dout(w_dff_A_K0Q8vH814_0),.din(w_dff_A_snZYENbb9_0),.clk(gclk));
	jdff dff_A_EbBtIif70_0(.dout(w_dff_A_snZYENbb9_0),.din(w_dff_A_EbBtIif70_0),.clk(gclk));
	jdff dff_A_HdLJGaXa4_0(.dout(w_dff_A_EbBtIif70_0),.din(w_dff_A_HdLJGaXa4_0),.clk(gclk));
	jdff dff_A_q1y7Ps4j4_0(.dout(w_dff_A_HdLJGaXa4_0),.din(w_dff_A_q1y7Ps4j4_0),.clk(gclk));
	jdff dff_A_ksqqvc4Z1_0(.dout(w_dff_A_q1y7Ps4j4_0),.din(w_dff_A_ksqqvc4Z1_0),.clk(gclk));
	jdff dff_A_b68mxddt9_0(.dout(w_n154_0[0]),.din(w_dff_A_b68mxddt9_0),.clk(gclk));
	jdff dff_A_ZWkZePY07_0(.dout(w_dff_A_b68mxddt9_0),.din(w_dff_A_ZWkZePY07_0),.clk(gclk));
	jdff dff_A_N0gRZj5j4_0(.dout(w_dff_A_ZWkZePY07_0),.din(w_dff_A_N0gRZj5j4_0),.clk(gclk));
	jdff dff_A_riHeQFHE6_0(.dout(w_dff_A_N0gRZj5j4_0),.din(w_dff_A_riHeQFHE6_0),.clk(gclk));
	jdff dff_A_nVOQsG7n6_0(.dout(w_dff_A_riHeQFHE6_0),.din(w_dff_A_nVOQsG7n6_0),.clk(gclk));
	jdff dff_B_1RMKlB3O8_2(.din(n154),.dout(w_dff_B_1RMKlB3O8_2),.clk(gclk));
	jdff dff_B_GHqBYcri8_2(.din(w_dff_B_1RMKlB3O8_2),.dout(w_dff_B_GHqBYcri8_2),.clk(gclk));
	jdff dff_B_MitMw2rq6_2(.din(w_dff_B_GHqBYcri8_2),.dout(w_dff_B_MitMw2rq6_2),.clk(gclk));
	jdff dff_B_ZsGj56ns4_2(.din(w_dff_B_MitMw2rq6_2),.dout(w_dff_B_ZsGj56ns4_2),.clk(gclk));
	jdff dff_B_raJoBPem6_2(.din(w_dff_B_ZsGj56ns4_2),.dout(w_dff_B_raJoBPem6_2),.clk(gclk));
	jdff dff_B_CjjwHvES6_2(.din(w_dff_B_raJoBPem6_2),.dout(w_dff_B_CjjwHvES6_2),.clk(gclk));
	jdff dff_B_uu7pN3IV6_2(.din(w_dff_B_CjjwHvES6_2),.dout(w_dff_B_uu7pN3IV6_2),.clk(gclk));
	jdff dff_B_EY1iwMLf3_2(.din(w_dff_B_uu7pN3IV6_2),.dout(w_dff_B_EY1iwMLf3_2),.clk(gclk));
	jdff dff_B_d4jRyJJU8_2(.din(w_dff_B_EY1iwMLf3_2),.dout(w_dff_B_d4jRyJJU8_2),.clk(gclk));
	jdff dff_B_zYeVc9io1_2(.din(w_dff_B_d4jRyJJU8_2),.dout(w_dff_B_zYeVc9io1_2),.clk(gclk));
	jdff dff_B_IisnITKx8_2(.din(w_dff_B_zYeVc9io1_2),.dout(w_dff_B_IisnITKx8_2),.clk(gclk));
	jdff dff_B_7pA7L4v44_2(.din(w_dff_B_IisnITKx8_2),.dout(w_dff_B_7pA7L4v44_2),.clk(gclk));
	jdff dff_B_cFVYd2oZ9_2(.din(w_dff_B_7pA7L4v44_2),.dout(w_dff_B_cFVYd2oZ9_2),.clk(gclk));
	jdff dff_B_rH6yLkox9_2(.din(w_dff_B_cFVYd2oZ9_2),.dout(w_dff_B_rH6yLkox9_2),.clk(gclk));
	jdff dff_A_qYlLBGYy1_0(.dout(w_G79gat_0[0]),.din(w_dff_A_qYlLBGYy1_0),.clk(gclk));
	jdff dff_A_VFpAPUid0_0(.dout(w_dff_A_qYlLBGYy1_0),.din(w_dff_A_VFpAPUid0_0),.clk(gclk));
	jdff dff_A_fypEEtHL9_0(.dout(w_dff_A_VFpAPUid0_0),.din(w_dff_A_fypEEtHL9_0),.clk(gclk));
	jdff dff_A_iXtCRgK81_0(.dout(w_dff_A_fypEEtHL9_0),.din(w_dff_A_iXtCRgK81_0),.clk(gclk));
	jdff dff_A_dPXEFUnt2_0(.dout(w_dff_A_iXtCRgK81_0),.din(w_dff_A_dPXEFUnt2_0),.clk(gclk));
	jdff dff_A_byao8ojn3_0(.dout(w_dff_A_dPXEFUnt2_0),.din(w_dff_A_byao8ojn3_0),.clk(gclk));
	jdff dff_A_Nz4JYgoN5_0(.dout(w_dff_A_byao8ojn3_0),.din(w_dff_A_Nz4JYgoN5_0),.clk(gclk));
	jdff dff_A_tD70mO059_0(.dout(w_dff_A_Nz4JYgoN5_0),.din(w_dff_A_tD70mO059_0),.clk(gclk));
	jdff dff_A_wBbd1NFf0_0(.dout(w_dff_A_tD70mO059_0),.din(w_dff_A_wBbd1NFf0_0),.clk(gclk));
	jdff dff_A_PSvwrhod2_0(.dout(w_dff_A_wBbd1NFf0_0),.din(w_dff_A_PSvwrhod2_0),.clk(gclk));
	jdff dff_A_gZmKyWcn5_0(.dout(w_dff_A_PSvwrhod2_0),.din(w_dff_A_gZmKyWcn5_0),.clk(gclk));
	jdff dff_A_NcqFU0L58_0(.dout(w_dff_A_gZmKyWcn5_0),.din(w_dff_A_NcqFU0L58_0),.clk(gclk));
	jdff dff_A_zRXLERNM2_0(.dout(w_dff_A_NcqFU0L58_0),.din(w_dff_A_zRXLERNM2_0),.clk(gclk));
	jdff dff_A_hDPmn0dQ4_0(.dout(w_dff_A_zRXLERNM2_0),.din(w_dff_A_hDPmn0dQ4_0),.clk(gclk));
	jdff dff_A_bGOh0Hws8_0(.dout(w_dff_A_hDPmn0dQ4_0),.din(w_dff_A_bGOh0Hws8_0),.clk(gclk));
	jdff dff_A_5gHrZgEA6_1(.dout(w_n151_0[1]),.din(w_dff_A_5gHrZgEA6_1),.clk(gclk));
	jdff dff_A_NUM62JuP8_1(.dout(w_dff_A_5gHrZgEA6_1),.din(w_dff_A_NUM62JuP8_1),.clk(gclk));
	jdff dff_A_Jpn7ckWw6_1(.dout(w_dff_A_NUM62JuP8_1),.din(w_dff_A_Jpn7ckWw6_1),.clk(gclk));
	jdff dff_A_IJkI0XNz8_1(.dout(w_dff_A_Jpn7ckWw6_1),.din(w_dff_A_IJkI0XNz8_1),.clk(gclk));
	jdff dff_A_3C1lhc792_1(.dout(w_dff_A_IJkI0XNz8_1),.din(w_dff_A_3C1lhc792_1),.clk(gclk));
	jdff dff_A_T0s3z3sR2_1(.dout(w_dff_A_3C1lhc792_1),.din(w_dff_A_T0s3z3sR2_1),.clk(gclk));
	jdff dff_A_8sTp01XR0_0(.dout(w_n150_0[0]),.din(w_dff_A_8sTp01XR0_0),.clk(gclk));
	jdff dff_A_7sRpbc9M9_0(.dout(w_dff_A_8sTp01XR0_0),.din(w_dff_A_7sRpbc9M9_0),.clk(gclk));
	jdff dff_A_4kYWIAMo9_0(.dout(w_dff_A_7sRpbc9M9_0),.din(w_dff_A_4kYWIAMo9_0),.clk(gclk));
	jdff dff_A_kesxjWgP2_0(.dout(w_dff_A_4kYWIAMo9_0),.din(w_dff_A_kesxjWgP2_0),.clk(gclk));
	jdff dff_A_IN3fy6eE8_0(.dout(w_dff_A_kesxjWgP2_0),.din(w_dff_A_IN3fy6eE8_0),.clk(gclk));
	jdff dff_A_rMk7h3SU1_0(.dout(w_dff_A_IN3fy6eE8_0),.din(w_dff_A_rMk7h3SU1_0),.clk(gclk));
	jdff dff_A_ovHUvAct6_0(.dout(w_dff_A_rMk7h3SU1_0),.din(w_dff_A_ovHUvAct6_0),.clk(gclk));
	jdff dff_A_cQgbo2fv9_0(.dout(w_dff_A_ovHUvAct6_0),.din(w_dff_A_cQgbo2fv9_0),.clk(gclk));
	jdff dff_A_L64DtgMK5_0(.dout(w_dff_A_cQgbo2fv9_0),.din(w_dff_A_L64DtgMK5_0),.clk(gclk));
	jdff dff_A_v11wllnh7_0(.dout(w_dff_A_L64DtgMK5_0),.din(w_dff_A_v11wllnh7_0),.clk(gclk));
	jdff dff_A_xN7FyZMI6_0(.dout(w_dff_A_v11wllnh7_0),.din(w_dff_A_xN7FyZMI6_0),.clk(gclk));
	jdff dff_A_nSTVCGDl6_0(.dout(w_dff_A_xN7FyZMI6_0),.din(w_dff_A_nSTVCGDl6_0),.clk(gclk));
	jdff dff_B_kpti7bC86_2(.din(n150),.dout(w_dff_B_kpti7bC86_2),.clk(gclk));
	jdff dff_B_nfh1bK2R7_2(.din(w_dff_B_kpti7bC86_2),.dout(w_dff_B_nfh1bK2R7_2),.clk(gclk));
	jdff dff_B_PGn0kuhK1_2(.din(w_dff_B_nfh1bK2R7_2),.dout(w_dff_B_PGn0kuhK1_2),.clk(gclk));
	jdff dff_B_kOqI0B0V4_2(.din(w_dff_B_PGn0kuhK1_2),.dout(w_dff_B_kOqI0B0V4_2),.clk(gclk));
	jdff dff_B_NhQ85tbn7_2(.din(w_dff_B_kOqI0B0V4_2),.dout(w_dff_B_NhQ85tbn7_2),.clk(gclk));
	jdff dff_B_XOnT76DQ5_2(.din(w_dff_B_NhQ85tbn7_2),.dout(w_dff_B_XOnT76DQ5_2),.clk(gclk));
	jdff dff_B_TIm7nUM62_2(.din(w_dff_B_XOnT76DQ5_2),.dout(w_dff_B_TIm7nUM62_2),.clk(gclk));
	jdff dff_A_lYDmnfP84_0(.dout(w_G66gat_0[0]),.din(w_dff_A_lYDmnfP84_0),.clk(gclk));
	jdff dff_A_l3j1r9iG1_0(.dout(w_dff_A_lYDmnfP84_0),.din(w_dff_A_l3j1r9iG1_0),.clk(gclk));
	jdff dff_A_qr19gKpt8_0(.dout(w_dff_A_l3j1r9iG1_0),.din(w_dff_A_qr19gKpt8_0),.clk(gclk));
	jdff dff_A_i8rpnUlF6_0(.dout(w_dff_A_qr19gKpt8_0),.din(w_dff_A_i8rpnUlF6_0),.clk(gclk));
	jdff dff_A_n9sCxsEg3_0(.dout(w_dff_A_i8rpnUlF6_0),.din(w_dff_A_n9sCxsEg3_0),.clk(gclk));
	jdff dff_A_mPue0nY78_0(.dout(w_dff_A_n9sCxsEg3_0),.din(w_dff_A_mPue0nY78_0),.clk(gclk));
	jdff dff_A_vEWMWh2b4_0(.dout(w_dff_A_mPue0nY78_0),.din(w_dff_A_vEWMWh2b4_0),.clk(gclk));
	jdff dff_A_Gsix6Qut1_0(.dout(w_dff_A_vEWMWh2b4_0),.din(w_dff_A_Gsix6Qut1_0),.clk(gclk));
	jdff dff_A_XfvMoU7F9_0(.dout(w_dff_A_Gsix6Qut1_0),.din(w_dff_A_XfvMoU7F9_0),.clk(gclk));
	jdff dff_A_X7VQjqwR9_0(.dout(w_dff_A_XfvMoU7F9_0),.din(w_dff_A_X7VQjqwR9_0),.clk(gclk));
	jdff dff_A_x7VzobFS0_0(.dout(w_dff_A_X7VQjqwR9_0),.din(w_dff_A_x7VzobFS0_0),.clk(gclk));
	jdff dff_A_P1OKVOCo9_0(.dout(w_dff_A_x7VzobFS0_0),.din(w_dff_A_P1OKVOCo9_0),.clk(gclk));
	jdff dff_A_3G261ipM6_0(.dout(w_dff_A_P1OKVOCo9_0),.din(w_dff_A_3G261ipM6_0),.clk(gclk));
	jdff dff_A_hmHrQWcu1_0(.dout(w_dff_A_3G261ipM6_0),.din(w_dff_A_hmHrQWcu1_0),.clk(gclk));
	jdff dff_A_4sWUQ9TC1_0(.dout(w_dff_A_hmHrQWcu1_0),.din(w_dff_A_4sWUQ9TC1_0),.clk(gclk));
	jdff dff_A_Z8wK5xfT4_0(.dout(w_dff_A_4sWUQ9TC1_0),.din(w_dff_A_Z8wK5xfT4_0),.clk(gclk));
	jdff dff_A_SnIvS7hs7_0(.dout(w_dff_A_Z8wK5xfT4_0),.din(w_dff_A_SnIvS7hs7_0),.clk(gclk));
	jdff dff_A_a9WYnEg51_0(.dout(w_dff_A_SnIvS7hs7_0),.din(w_dff_A_a9WYnEg51_0),.clk(gclk));
	jdff dff_A_Nl0tmKmw8_0(.dout(w_dff_A_a9WYnEg51_0),.din(w_dff_A_Nl0tmKmw8_0),.clk(gclk));
	jdff dff_A_bLe8H6p09_0(.dout(w_dff_A_Nl0tmKmw8_0),.din(w_dff_A_bLe8H6p09_0),.clk(gclk));
	jdff dff_A_AIDxYJ9G6_1(.dout(w_n146_0[1]),.din(w_dff_A_AIDxYJ9G6_1),.clk(gclk));
	jdff dff_A_2AEEYJqS8_1(.dout(w_dff_A_AIDxYJ9G6_1),.din(w_dff_A_2AEEYJqS8_1),.clk(gclk));
	jdff dff_A_IT9vBcB24_1(.dout(w_dff_A_2AEEYJqS8_1),.din(w_dff_A_IT9vBcB24_1),.clk(gclk));
	jdff dff_A_xmlZg3DD4_1(.dout(w_dff_A_IT9vBcB24_1),.din(w_dff_A_xmlZg3DD4_1),.clk(gclk));
	jdff dff_A_rrsiezFj2_0(.dout(w_n145_0[0]),.din(w_dff_A_rrsiezFj2_0),.clk(gclk));
	jdff dff_A_yIMOIQR95_0(.dout(w_dff_A_rrsiezFj2_0),.din(w_dff_A_yIMOIQR95_0),.clk(gclk));
	jdff dff_A_M2NGVda55_0(.dout(w_dff_A_yIMOIQR95_0),.din(w_dff_A_M2NGVda55_0),.clk(gclk));
	jdff dff_A_YZAjzOGS5_0(.dout(w_dff_A_M2NGVda55_0),.din(w_dff_A_YZAjzOGS5_0),.clk(gclk));
	jdff dff_A_IXZTYsXj7_0(.dout(w_dff_A_YZAjzOGS5_0),.din(w_dff_A_IXZTYsXj7_0),.clk(gclk));
	jdff dff_A_XDhjYOjs0_0(.dout(w_dff_A_IXZTYsXj7_0),.din(w_dff_A_XDhjYOjs0_0),.clk(gclk));
	jdff dff_A_KX1ModdX8_0(.dout(w_n142_0[0]),.din(w_dff_A_KX1ModdX8_0),.clk(gclk));
	jdff dff_B_R8Vd1Y862_1(.din(n112),.dout(w_dff_B_R8Vd1Y862_1),.clk(gclk));
	jdff dff_B_Th0bZbSX7_1(.din(n116),.dout(w_dff_B_Th0bZbSX7_1),.clk(gclk));
	jdff dff_A_17BocApl2_0(.dout(w_n132_0[0]),.din(w_dff_A_17BocApl2_0),.clk(gclk));
	jdff dff_A_vTr7s9CO0_0(.dout(w_dff_A_17BocApl2_0),.din(w_dff_A_vTr7s9CO0_0),.clk(gclk));
	jdff dff_A_2ktGVcgN2_0(.dout(w_dff_A_vTr7s9CO0_0),.din(w_dff_A_2ktGVcgN2_0),.clk(gclk));
	jdff dff_A_rc33XG8z9_0(.dout(w_dff_A_2ktGVcgN2_0),.din(w_dff_A_rc33XG8z9_0),.clk(gclk));
	jdff dff_A_TdrK4NG03_0(.dout(w_dff_A_rc33XG8z9_0),.din(w_dff_A_TdrK4NG03_0),.clk(gclk));
	jdff dff_A_hu9pQrxC8_0(.dout(w_dff_A_TdrK4NG03_0),.din(w_dff_A_hu9pQrxC8_0),.clk(gclk));
	jdff dff_A_fUwSAHnP7_0(.dout(w_n130_0[0]),.din(w_dff_A_fUwSAHnP7_0),.clk(gclk));
	jdff dff_A_DqQU4o6f3_0(.dout(w_dff_A_fUwSAHnP7_0),.din(w_dff_A_DqQU4o6f3_0),.clk(gclk));
	jdff dff_A_FTwM55dh5_0(.dout(w_dff_A_DqQU4o6f3_0),.din(w_dff_A_FTwM55dh5_0),.clk(gclk));
	jdff dff_A_Y85qGYMh1_0(.dout(w_dff_A_FTwM55dh5_0),.din(w_dff_A_Y85qGYMh1_0),.clk(gclk));
	jdff dff_A_x8N6BIx90_0(.dout(w_dff_A_Y85qGYMh1_0),.din(w_dff_A_x8N6BIx90_0),.clk(gclk));
	jdff dff_A_RrQPXJxg2_1(.dout(w_n130_0[1]),.din(w_dff_A_RrQPXJxg2_1),.clk(gclk));
	jdff dff_A_izS0yXx20_1(.dout(w_dff_A_RrQPXJxg2_1),.din(w_dff_A_izS0yXx20_1),.clk(gclk));
	jdff dff_A_vpnLmV4O8_1(.dout(w_dff_A_izS0yXx20_1),.din(w_dff_A_vpnLmV4O8_1),.clk(gclk));
	jdff dff_A_ERz3NTiY9_1(.dout(w_dff_A_vpnLmV4O8_1),.din(w_dff_A_ERz3NTiY9_1),.clk(gclk));
	jdff dff_A_6J44yqVi5_1(.dout(w_dff_A_ERz3NTiY9_1),.din(w_dff_A_6J44yqVi5_1),.clk(gclk));
	jdff dff_B_Rg5ppKOc6_3(.din(n130),.dout(w_dff_B_Rg5ppKOc6_3),.clk(gclk));
	jdff dff_B_hZLMDhas8_3(.din(w_dff_B_Rg5ppKOc6_3),.dout(w_dff_B_hZLMDhas8_3),.clk(gclk));
	jdff dff_B_waXoQRFE5_3(.din(w_dff_B_hZLMDhas8_3),.dout(w_dff_B_waXoQRFE5_3),.clk(gclk));
	jdff dff_B_xmYFxO0r9_3(.din(w_dff_B_waXoQRFE5_3),.dout(w_dff_B_xmYFxO0r9_3),.clk(gclk));
	jdff dff_B_r3VoOClJ3_3(.din(w_dff_B_xmYFxO0r9_3),.dout(w_dff_B_r3VoOClJ3_3),.clk(gclk));
	jdff dff_B_X97IjzTs3_3(.din(w_dff_B_r3VoOClJ3_3),.dout(w_dff_B_X97IjzTs3_3),.clk(gclk));
	jdff dff_B_LBdoCohI3_3(.din(w_dff_B_X97IjzTs3_3),.dout(w_dff_B_LBdoCohI3_3),.clk(gclk));
	jdff dff_A_MzlYi6693_0(.dout(w_G21gat_1[0]),.din(w_dff_A_MzlYi6693_0),.clk(gclk));
	jdff dff_A_HPLJABdF1_0(.dout(w_dff_A_MzlYi6693_0),.din(w_dff_A_HPLJABdF1_0),.clk(gclk));
	jdff dff_A_X1nS95J47_0(.dout(w_dff_A_HPLJABdF1_0),.din(w_dff_A_X1nS95J47_0),.clk(gclk));
	jdff dff_A_RvYCg9X30_0(.dout(w_dff_A_X1nS95J47_0),.din(w_dff_A_RvYCg9X30_0),.clk(gclk));
	jdff dff_A_IeiXacB89_0(.dout(w_dff_A_RvYCg9X30_0),.din(w_dff_A_IeiXacB89_0),.clk(gclk));
	jdff dff_A_GMp2h9k91_0(.dout(w_dff_A_IeiXacB89_0),.din(w_dff_A_GMp2h9k91_0),.clk(gclk));
	jdff dff_A_QZcrQiBJ2_0(.dout(w_dff_A_GMp2h9k91_0),.din(w_dff_A_QZcrQiBJ2_0),.clk(gclk));
	jdff dff_A_0xg2965M0_0(.dout(w_dff_A_QZcrQiBJ2_0),.din(w_dff_A_0xg2965M0_0),.clk(gclk));
	jdff dff_A_a03MS5ke3_1(.dout(w_G21gat_0[1]),.din(w_dff_A_a03MS5ke3_1),.clk(gclk));
	jdff dff_A_0O1lrRPI0_1(.dout(w_dff_A_a03MS5ke3_1),.din(w_dff_A_0O1lrRPI0_1),.clk(gclk));
	jdff dff_A_t0MEXTHS5_1(.dout(w_dff_A_0O1lrRPI0_1),.din(w_dff_A_t0MEXTHS5_1),.clk(gclk));
	jdff dff_A_yfIh0WJZ2_1(.dout(w_dff_A_t0MEXTHS5_1),.din(w_dff_A_yfIh0WJZ2_1),.clk(gclk));
	jdff dff_A_NKO9YvAH3_1(.dout(w_dff_A_yfIh0WJZ2_1),.din(w_dff_A_NKO9YvAH3_1),.clk(gclk));
	jdff dff_A_SxUcyHIb0_1(.dout(w_dff_A_NKO9YvAH3_1),.din(w_dff_A_SxUcyHIb0_1),.clk(gclk));
	jdff dff_A_jiRfFmRG7_1(.dout(w_dff_A_SxUcyHIb0_1),.din(w_dff_A_jiRfFmRG7_1),.clk(gclk));
	jdff dff_A_rWB4pGIe4_1(.dout(w_dff_A_jiRfFmRG7_1),.din(w_dff_A_rWB4pGIe4_1),.clk(gclk));
	jdff dff_A_ljGEyeDp4_1(.dout(w_dff_A_rWB4pGIe4_1),.din(w_dff_A_ljGEyeDp4_1),.clk(gclk));
	jdff dff_A_1D1a4aev2_1(.dout(w_dff_A_ljGEyeDp4_1),.din(w_dff_A_1D1a4aev2_1),.clk(gclk));
	jdff dff_A_RNnfeCJp4_1(.dout(w_dff_A_1D1a4aev2_1),.din(w_dff_A_RNnfeCJp4_1),.clk(gclk));
	jdff dff_A_jJrumhP34_1(.dout(w_dff_A_RNnfeCJp4_1),.din(w_dff_A_jJrumhP34_1),.clk(gclk));
	jdff dff_A_AnuNYbET2_1(.dout(w_dff_A_jJrumhP34_1),.din(w_dff_A_AnuNYbET2_1),.clk(gclk));
	jdff dff_A_2wiB24I18_2(.dout(w_G21gat_0[2]),.din(w_dff_A_2wiB24I18_2),.clk(gclk));
	jdff dff_A_1bVVJn7F4_2(.dout(w_dff_A_2wiB24I18_2),.din(w_dff_A_1bVVJn7F4_2),.clk(gclk));
	jdff dff_A_W4iGEOUq6_2(.dout(w_dff_A_1bVVJn7F4_2),.din(w_dff_A_W4iGEOUq6_2),.clk(gclk));
	jdff dff_A_DcRihHgS3_2(.dout(w_dff_A_W4iGEOUq6_2),.din(w_dff_A_DcRihHgS3_2),.clk(gclk));
	jdff dff_A_G06VqZMI9_2(.dout(w_dff_A_DcRihHgS3_2),.din(w_dff_A_G06VqZMI9_2),.clk(gclk));
	jdff dff_A_hfEZImHd0_2(.dout(w_dff_A_G06VqZMI9_2),.din(w_dff_A_hfEZImHd0_2),.clk(gclk));
	jdff dff_A_XnEwKKVn6_2(.dout(w_dff_A_hfEZImHd0_2),.din(w_dff_A_XnEwKKVn6_2),.clk(gclk));
	jdff dff_A_luh1VQBJ3_2(.dout(w_dff_A_XnEwKKVn6_2),.din(w_dff_A_luh1VQBJ3_2),.clk(gclk));
	jdff dff_A_MlPnIsTV0_2(.dout(w_dff_A_luh1VQBJ3_2),.din(w_dff_A_MlPnIsTV0_2),.clk(gclk));
	jdff dff_A_sM399QWP4_2(.dout(w_dff_A_MlPnIsTV0_2),.din(w_dff_A_sM399QWP4_2),.clk(gclk));
	jdff dff_A_KNuj8YSH5_2(.dout(w_dff_A_sM399QWP4_2),.din(w_dff_A_KNuj8YSH5_2),.clk(gclk));
	jdff dff_A_RbJvjMg10_2(.dout(w_dff_A_KNuj8YSH5_2),.din(w_dff_A_RbJvjMg10_2),.clk(gclk));
	jdff dff_A_EqMDbWfC8_2(.dout(w_dff_A_RbJvjMg10_2),.din(w_dff_A_EqMDbWfC8_2),.clk(gclk));
	jdff dff_A_2Slsgt950_0(.dout(w_n128_0[0]),.din(w_dff_A_2Slsgt950_0),.clk(gclk));
	jdff dff_A_PrMFEnlF9_0(.dout(w_dff_A_2Slsgt950_0),.din(w_dff_A_PrMFEnlF9_0),.clk(gclk));
	jdff dff_A_FC2xk7wu5_0(.dout(w_dff_A_PrMFEnlF9_0),.din(w_dff_A_FC2xk7wu5_0),.clk(gclk));
	jdff dff_A_fe7q5SvS8_0(.dout(w_dff_A_FC2xk7wu5_0),.din(w_dff_A_fe7q5SvS8_0),.clk(gclk));
	jdff dff_A_jI5H6wEV3_0(.dout(w_dff_A_fe7q5SvS8_0),.din(w_dff_A_jI5H6wEV3_0),.clk(gclk));
	jdff dff_A_AEVTHE0x9_0(.dout(w_dff_A_jI5H6wEV3_0),.din(w_dff_A_AEVTHE0x9_0),.clk(gclk));
	jdff dff_A_1UWHiTsb7_0(.dout(w_n126_0[0]),.din(w_dff_A_1UWHiTsb7_0),.clk(gclk));
	jdff dff_A_Rdh9eGGB7_0(.dout(w_dff_A_1UWHiTsb7_0),.din(w_dff_A_Rdh9eGGB7_0),.clk(gclk));
	jdff dff_A_EHJSa9or2_0(.dout(w_dff_A_Rdh9eGGB7_0),.din(w_dff_A_EHJSa9or2_0),.clk(gclk));
	jdff dff_A_UI3hdeyU8_0(.dout(w_dff_A_EHJSa9or2_0),.din(w_dff_A_UI3hdeyU8_0),.clk(gclk));
	jdff dff_A_kN9ZTeBs8_0(.dout(w_dff_A_UI3hdeyU8_0),.din(w_dff_A_kN9ZTeBs8_0),.clk(gclk));
	jdff dff_A_VEScWGPm7_1(.dout(w_n126_0[1]),.din(w_dff_A_VEScWGPm7_1),.clk(gclk));
	jdff dff_A_fGWlJH8a1_1(.dout(w_dff_A_VEScWGPm7_1),.din(w_dff_A_fGWlJH8a1_1),.clk(gclk));
	jdff dff_A_3ENjGzBi2_1(.dout(w_dff_A_fGWlJH8a1_1),.din(w_dff_A_3ENjGzBi2_1),.clk(gclk));
	jdff dff_A_o9gC6ODv9_1(.dout(w_dff_A_3ENjGzBi2_1),.din(w_dff_A_o9gC6ODv9_1),.clk(gclk));
	jdff dff_A_fpMbBfaE7_1(.dout(w_dff_A_o9gC6ODv9_1),.din(w_dff_A_fpMbBfaE7_1),.clk(gclk));
	jdff dff_B_LRrV6wS22_3(.din(n126),.dout(w_dff_B_LRrV6wS22_3),.clk(gclk));
	jdff dff_B_xPW0G9qm7_3(.din(w_dff_B_LRrV6wS22_3),.dout(w_dff_B_xPW0G9qm7_3),.clk(gclk));
	jdff dff_B_vAGnO8v30_3(.din(w_dff_B_xPW0G9qm7_3),.dout(w_dff_B_vAGnO8v30_3),.clk(gclk));
	jdff dff_B_DYsOGOrM2_3(.din(w_dff_B_vAGnO8v30_3),.dout(w_dff_B_DYsOGOrM2_3),.clk(gclk));
	jdff dff_B_qeRTY36U7_3(.din(w_dff_B_DYsOGOrM2_3),.dout(w_dff_B_qeRTY36U7_3),.clk(gclk));
	jdff dff_B_YD8DtHMo4_3(.din(w_dff_B_qeRTY36U7_3),.dout(w_dff_B_YD8DtHMo4_3),.clk(gclk));
	jdff dff_B_EJOsXWCr7_3(.din(w_dff_B_YD8DtHMo4_3),.dout(w_dff_B_EJOsXWCr7_3),.clk(gclk));
	jdff dff_A_4sNZR7UB2_0(.dout(w_G86gat_1[0]),.din(w_dff_A_4sNZR7UB2_0),.clk(gclk));
	jdff dff_A_ydCpUvMA4_0(.dout(w_dff_A_4sNZR7UB2_0),.din(w_dff_A_ydCpUvMA4_0),.clk(gclk));
	jdff dff_A_wE2G8o0g0_0(.dout(w_dff_A_ydCpUvMA4_0),.din(w_dff_A_wE2G8o0g0_0),.clk(gclk));
	jdff dff_A_SQIvKpWR7_0(.dout(w_dff_A_wE2G8o0g0_0),.din(w_dff_A_SQIvKpWR7_0),.clk(gclk));
	jdff dff_A_MI5SidWk4_0(.dout(w_dff_A_SQIvKpWR7_0),.din(w_dff_A_MI5SidWk4_0),.clk(gclk));
	jdff dff_A_9VZNu7av4_0(.dout(w_dff_A_MI5SidWk4_0),.din(w_dff_A_9VZNu7av4_0),.clk(gclk));
	jdff dff_A_8Q1g5X928_0(.dout(w_dff_A_9VZNu7av4_0),.din(w_dff_A_8Q1g5X928_0),.clk(gclk));
	jdff dff_A_KxUoyAUl5_0(.dout(w_dff_A_8Q1g5X928_0),.din(w_dff_A_KxUoyAUl5_0),.clk(gclk));
	jdff dff_A_Z44nTf0r4_1(.dout(w_G86gat_0[1]),.din(w_dff_A_Z44nTf0r4_1),.clk(gclk));
	jdff dff_A_gMsWFqAx4_1(.dout(w_dff_A_Z44nTf0r4_1),.din(w_dff_A_gMsWFqAx4_1),.clk(gclk));
	jdff dff_A_XVqTyLLg2_1(.dout(w_dff_A_gMsWFqAx4_1),.din(w_dff_A_XVqTyLLg2_1),.clk(gclk));
	jdff dff_A_7mgSZIR06_1(.dout(w_dff_A_XVqTyLLg2_1),.din(w_dff_A_7mgSZIR06_1),.clk(gclk));
	jdff dff_A_CoxH234X8_1(.dout(w_dff_A_7mgSZIR06_1),.din(w_dff_A_CoxH234X8_1),.clk(gclk));
	jdff dff_A_oJIPV0cc2_1(.dout(w_dff_A_CoxH234X8_1),.din(w_dff_A_oJIPV0cc2_1),.clk(gclk));
	jdff dff_A_wOo4d2rT9_1(.dout(w_dff_A_oJIPV0cc2_1),.din(w_dff_A_wOo4d2rT9_1),.clk(gclk));
	jdff dff_A_wzBecpQF9_1(.dout(w_dff_A_wOo4d2rT9_1),.din(w_dff_A_wzBecpQF9_1),.clk(gclk));
	jdff dff_A_PtGVaBZo1_1(.dout(w_dff_A_wzBecpQF9_1),.din(w_dff_A_PtGVaBZo1_1),.clk(gclk));
	jdff dff_A_3uqCe2780_1(.dout(w_dff_A_PtGVaBZo1_1),.din(w_dff_A_3uqCe2780_1),.clk(gclk));
	jdff dff_A_CKmFsCV74_1(.dout(w_dff_A_3uqCe2780_1),.din(w_dff_A_CKmFsCV74_1),.clk(gclk));
	jdff dff_A_BPEcofBo1_1(.dout(w_dff_A_CKmFsCV74_1),.din(w_dff_A_BPEcofBo1_1),.clk(gclk));
	jdff dff_A_hYqOcECy2_1(.dout(w_dff_A_BPEcofBo1_1),.din(w_dff_A_hYqOcECy2_1),.clk(gclk));
	jdff dff_A_fR8Cs5L65_2(.dout(w_G86gat_0[2]),.din(w_dff_A_fR8Cs5L65_2),.clk(gclk));
	jdff dff_A_YGZtKVcG9_2(.dout(w_dff_A_fR8Cs5L65_2),.din(w_dff_A_YGZtKVcG9_2),.clk(gclk));
	jdff dff_A_DUWNIw329_2(.dout(w_dff_A_YGZtKVcG9_2),.din(w_dff_A_DUWNIw329_2),.clk(gclk));
	jdff dff_A_IpLVUsRp4_2(.dout(w_dff_A_DUWNIw329_2),.din(w_dff_A_IpLVUsRp4_2),.clk(gclk));
	jdff dff_A_vv7Ix2Cr4_2(.dout(w_dff_A_IpLVUsRp4_2),.din(w_dff_A_vv7Ix2Cr4_2),.clk(gclk));
	jdff dff_A_Q3dAwGgf1_2(.dout(w_dff_A_vv7Ix2Cr4_2),.din(w_dff_A_Q3dAwGgf1_2),.clk(gclk));
	jdff dff_A_4Gh2no2J3_2(.dout(w_dff_A_Q3dAwGgf1_2),.din(w_dff_A_4Gh2no2J3_2),.clk(gclk));
	jdff dff_A_LnRsB3X39_2(.dout(w_dff_A_4Gh2no2J3_2),.din(w_dff_A_LnRsB3X39_2),.clk(gclk));
	jdff dff_A_0LKmHaRj2_2(.dout(w_dff_A_LnRsB3X39_2),.din(w_dff_A_0LKmHaRj2_2),.clk(gclk));
	jdff dff_A_C6EnUrQ51_2(.dout(w_dff_A_0LKmHaRj2_2),.din(w_dff_A_C6EnUrQ51_2),.clk(gclk));
	jdff dff_A_xHBjpzyj3_2(.dout(w_dff_A_C6EnUrQ51_2),.din(w_dff_A_xHBjpzyj3_2),.clk(gclk));
	jdff dff_A_W5z35fdo1_2(.dout(w_dff_A_xHBjpzyj3_2),.din(w_dff_A_W5z35fdo1_2),.clk(gclk));
	jdff dff_A_odwdWGJj5_2(.dout(w_dff_A_W5z35fdo1_2),.din(w_dff_A_odwdWGJj5_2),.clk(gclk));
	jdff dff_B_OxpkzM984_0(.din(n124),.dout(w_dff_B_OxpkzM984_0),.clk(gclk));
	jdff dff_A_9KITWTJo0_1(.dout(w_n123_0[1]),.din(w_dff_A_9KITWTJo0_1),.clk(gclk));
	jdff dff_A_bZnqd2iU8_1(.dout(w_dff_A_9KITWTJo0_1),.din(w_dff_A_bZnqd2iU8_1),.clk(gclk));
	jdff dff_A_w4H13SsZ4_1(.dout(w_dff_A_bZnqd2iU8_1),.din(w_dff_A_w4H13SsZ4_1),.clk(gclk));
	jdff dff_A_mB1PvCTJ0_1(.dout(w_dff_A_w4H13SsZ4_1),.din(w_dff_A_mB1PvCTJ0_1),.clk(gclk));
	jdff dff_A_iqB8XFrz2_1(.dout(w_dff_A_mB1PvCTJ0_1),.din(w_dff_A_iqB8XFrz2_1),.clk(gclk));
	jdff dff_A_IYSUvkzA5_0(.dout(w_G47gat_0[0]),.din(w_dff_A_IYSUvkzA5_0),.clk(gclk));
	jdff dff_A_WTy4IQS20_0(.dout(w_dff_A_IYSUvkzA5_0),.din(w_dff_A_WTy4IQS20_0),.clk(gclk));
	jdff dff_A_7ywQi2RU4_0(.dout(w_dff_A_WTy4IQS20_0),.din(w_dff_A_7ywQi2RU4_0),.clk(gclk));
	jdff dff_A_ynTSB2Wr9_0(.dout(w_dff_A_7ywQi2RU4_0),.din(w_dff_A_ynTSB2Wr9_0),.clk(gclk));
	jdff dff_A_gDkAM4OE9_0(.dout(w_dff_A_ynTSB2Wr9_0),.din(w_dff_A_gDkAM4OE9_0),.clk(gclk));
	jdff dff_A_shGNqpox9_0(.dout(w_dff_A_gDkAM4OE9_0),.din(w_dff_A_shGNqpox9_0),.clk(gclk));
	jdff dff_A_6dYPZCWG4_0(.dout(w_dff_A_shGNqpox9_0),.din(w_dff_A_6dYPZCWG4_0),.clk(gclk));
	jdff dff_A_OAxUb3DU5_0(.dout(w_dff_A_6dYPZCWG4_0),.din(w_dff_A_OAxUb3DU5_0),.clk(gclk));
	jdff dff_A_rHUgqz9x2_0(.dout(w_dff_A_OAxUb3DU5_0),.din(w_dff_A_rHUgqz9x2_0),.clk(gclk));
	jdff dff_A_wTbqIYQi7_0(.dout(w_dff_A_rHUgqz9x2_0),.din(w_dff_A_wTbqIYQi7_0),.clk(gclk));
	jdff dff_A_4QaiZaVe2_0(.dout(w_dff_A_wTbqIYQi7_0),.din(w_dff_A_4QaiZaVe2_0),.clk(gclk));
	jdff dff_A_W7Zzlw3Y0_0(.dout(w_dff_A_4QaiZaVe2_0),.din(w_dff_A_W7Zzlw3Y0_0),.clk(gclk));
	jdff dff_A_vB3sY1hH0_0(.dout(w_dff_A_W7Zzlw3Y0_0),.din(w_dff_A_vB3sY1hH0_0),.clk(gclk));
	jdff dff_B_EPHpvZa76_1(.din(n117),.dout(w_dff_B_EPHpvZa76_1),.clk(gclk));
	jdff dff_B_fNTkLBlZ1_1(.din(w_dff_B_EPHpvZa76_1),.dout(w_dff_B_fNTkLBlZ1_1),.clk(gclk));
	jdff dff_B_64Fn2s6K4_1(.din(w_dff_B_fNTkLBlZ1_1),.dout(w_dff_B_64Fn2s6K4_1),.clk(gclk));
	jdff dff_B_VvAtyVfB2_1(.din(w_dff_B_64Fn2s6K4_1),.dout(w_dff_B_VvAtyVfB2_1),.clk(gclk));
	jdff dff_B_ntOmAcnj5_1(.din(w_dff_B_VvAtyVfB2_1),.dout(w_dff_B_ntOmAcnj5_1),.clk(gclk));
	jdff dff_B_SoKwzb5s1_1(.din(w_dff_B_ntOmAcnj5_1),.dout(w_dff_B_SoKwzb5s1_1),.clk(gclk));
	jdff dff_B_tSMI6Fck6_1(.din(w_dff_B_SoKwzb5s1_1),.dout(w_dff_B_tSMI6Fck6_1),.clk(gclk));
	jdff dff_A_bLvtzvXe2_0(.dout(w_G60gat_0[0]),.din(w_dff_A_bLvtzvXe2_0),.clk(gclk));
	jdff dff_A_4TAxMss03_0(.dout(w_dff_A_bLvtzvXe2_0),.din(w_dff_A_4TAxMss03_0),.clk(gclk));
	jdff dff_A_ZnYSqwsH8_0(.dout(w_dff_A_4TAxMss03_0),.din(w_dff_A_ZnYSqwsH8_0),.clk(gclk));
	jdff dff_A_XLJaHVqe4_0(.dout(w_dff_A_ZnYSqwsH8_0),.din(w_dff_A_XLJaHVqe4_0),.clk(gclk));
	jdff dff_A_vxBEYnpb6_0(.dout(w_dff_A_XLJaHVqe4_0),.din(w_dff_A_vxBEYnpb6_0),.clk(gclk));
	jdff dff_A_YdNyOqj98_0(.dout(w_dff_A_vxBEYnpb6_0),.din(w_dff_A_YdNyOqj98_0),.clk(gclk));
	jdff dff_A_N64fzS6w5_0(.dout(w_dff_A_YdNyOqj98_0),.din(w_dff_A_N64fzS6w5_0),.clk(gclk));
	jdff dff_A_5cSTr67n4_0(.dout(w_dff_A_N64fzS6w5_0),.din(w_dff_A_5cSTr67n4_0),.clk(gclk));
	jdff dff_A_BrOy5uzJ3_0(.dout(w_dff_A_5cSTr67n4_0),.din(w_dff_A_BrOy5uzJ3_0),.clk(gclk));
	jdff dff_A_VFqIDk5p9_0(.dout(w_dff_A_BrOy5uzJ3_0),.din(w_dff_A_VFqIDk5p9_0),.clk(gclk));
	jdff dff_A_dPrwv1Md1_0(.dout(w_dff_A_VFqIDk5p9_0),.din(w_dff_A_dPrwv1Md1_0),.clk(gclk));
	jdff dff_A_TadI1wsu9_0(.dout(w_dff_A_dPrwv1Md1_0),.din(w_dff_A_TadI1wsu9_0),.clk(gclk));
	jdff dff_A_XVlost7X3_0(.dout(w_dff_A_TadI1wsu9_0),.din(w_dff_A_XVlost7X3_0),.clk(gclk));
	jdff dff_A_6g67yAoj4_1(.dout(w_G60gat_0[1]),.din(w_dff_A_6g67yAoj4_1),.clk(gclk));
	jdff dff_A_sFUuqw4y0_1(.dout(w_dff_A_6g67yAoj4_1),.din(w_dff_A_sFUuqw4y0_1),.clk(gclk));
	jdff dff_A_7uTFjCQq5_1(.dout(w_dff_A_sFUuqw4y0_1),.din(w_dff_A_7uTFjCQq5_1),.clk(gclk));
	jdff dff_A_9VpKTKMg0_1(.dout(w_dff_A_7uTFjCQq5_1),.din(w_dff_A_9VpKTKMg0_1),.clk(gclk));
	jdff dff_A_k2b9yXf68_1(.dout(w_dff_A_9VpKTKMg0_1),.din(w_dff_A_k2b9yXf68_1),.clk(gclk));
	jdff dff_A_IABRNTZn5_1(.dout(w_dff_A_k2b9yXf68_1),.din(w_dff_A_IABRNTZn5_1),.clk(gclk));
	jdff dff_A_UkJN3UFC4_1(.dout(w_dff_A_IABRNTZn5_1),.din(w_dff_A_UkJN3UFC4_1),.clk(gclk));
	jdff dff_A_MIEOTvSw8_1(.dout(w_dff_A_UkJN3UFC4_1),.din(w_dff_A_MIEOTvSw8_1),.clk(gclk));
	jdff dff_A_LZ7sZsWZ2_0(.dout(w_n115_0[0]),.din(w_dff_A_LZ7sZsWZ2_0),.clk(gclk));
	jdff dff_A_31Pa4CSX5_0(.dout(w_dff_A_LZ7sZsWZ2_0),.din(w_dff_A_31Pa4CSX5_0),.clk(gclk));
	jdff dff_A_PgHy2STv3_0(.dout(w_n114_0[0]),.din(w_dff_A_PgHy2STv3_0),.clk(gclk));
	jdff dff_A_ovK79HB99_0(.dout(w_dff_A_PgHy2STv3_0),.din(w_dff_A_ovK79HB99_0),.clk(gclk));
	jdff dff_A_P81jYeST0_0(.dout(w_dff_A_ovK79HB99_0),.din(w_dff_A_P81jYeST0_0),.clk(gclk));
	jdff dff_A_Kmbdn2pq0_0(.dout(w_dff_A_P81jYeST0_0),.din(w_dff_A_Kmbdn2pq0_0),.clk(gclk));
	jdff dff_A_KTZTvfx64_0(.dout(w_dff_A_Kmbdn2pq0_0),.din(w_dff_A_KTZTvfx64_0),.clk(gclk));
	jdff dff_A_M8D3VRA67_0(.dout(w_dff_A_KTZTvfx64_0),.din(w_dff_A_M8D3VRA67_0),.clk(gclk));
	jdff dff_A_DXFXV68v4_0(.dout(w_G34gat_0[0]),.din(w_dff_A_DXFXV68v4_0),.clk(gclk));
	jdff dff_A_dZP5vuZV4_0(.dout(w_dff_A_DXFXV68v4_0),.din(w_dff_A_dZP5vuZV4_0),.clk(gclk));
	jdff dff_A_xW8HEi8H2_0(.dout(w_dff_A_dZP5vuZV4_0),.din(w_dff_A_xW8HEi8H2_0),.clk(gclk));
	jdff dff_A_HIezcUiV6_0(.dout(w_dff_A_xW8HEi8H2_0),.din(w_dff_A_HIezcUiV6_0),.clk(gclk));
	jdff dff_A_IsorQJC72_0(.dout(w_dff_A_HIezcUiV6_0),.din(w_dff_A_IsorQJC72_0),.clk(gclk));
	jdff dff_A_RQDElPUt8_0(.dout(w_dff_A_IsorQJC72_0),.din(w_dff_A_RQDElPUt8_0),.clk(gclk));
	jdff dff_A_cExgftl28_0(.dout(w_dff_A_RQDElPUt8_0),.din(w_dff_A_cExgftl28_0),.clk(gclk));
	jdff dff_A_2v7fzme99_0(.dout(w_dff_A_cExgftl28_0),.din(w_dff_A_2v7fzme99_0),.clk(gclk));
	jdff dff_A_sM0Ik8On6_0(.dout(w_dff_A_2v7fzme99_0),.din(w_dff_A_sM0Ik8On6_0),.clk(gclk));
	jdff dff_A_4i5nevIg5_0(.dout(w_dff_A_sM0Ik8On6_0),.din(w_dff_A_4i5nevIg5_0),.clk(gclk));
	jdff dff_A_69Mmyz0e6_0(.dout(w_dff_A_4i5nevIg5_0),.din(w_dff_A_69Mmyz0e6_0),.clk(gclk));
	jdff dff_A_pBI6V4ut8_0(.dout(w_dff_A_69Mmyz0e6_0),.din(w_dff_A_pBI6V4ut8_0),.clk(gclk));
	jdff dff_A_GoDra4tL5_0(.dout(w_dff_A_pBI6V4ut8_0),.din(w_dff_A_GoDra4tL5_0),.clk(gclk));
	jdff dff_A_8FvCFuRb6_2(.dout(w_G34gat_0[2]),.din(w_dff_A_8FvCFuRb6_2),.clk(gclk));
	jdff dff_A_4ZitChP85_2(.dout(w_dff_A_8FvCFuRb6_2),.din(w_dff_A_4ZitChP85_2),.clk(gclk));
	jdff dff_A_mhRoJZen2_2(.dout(w_dff_A_4ZitChP85_2),.din(w_dff_A_mhRoJZen2_2),.clk(gclk));
	jdff dff_A_4jkALRE69_2(.dout(w_dff_A_mhRoJZen2_2),.din(w_dff_A_4jkALRE69_2),.clk(gclk));
	jdff dff_A_njfgyGdm0_2(.dout(w_dff_A_4jkALRE69_2),.din(w_dff_A_njfgyGdm0_2),.clk(gclk));
	jdff dff_A_NeRgcosv0_2(.dout(w_dff_A_njfgyGdm0_2),.din(w_dff_A_NeRgcosv0_2),.clk(gclk));
	jdff dff_A_Tlk99gAy3_2(.dout(w_dff_A_NeRgcosv0_2),.din(w_dff_A_Tlk99gAy3_2),.clk(gclk));
	jdff dff_A_SSDLaLU77_2(.dout(w_dff_A_Tlk99gAy3_2),.din(w_dff_A_SSDLaLU77_2),.clk(gclk));
	jdff dff_A_thL9YslX9_0(.dout(w_n109_0[0]),.din(w_dff_A_thL9YslX9_0),.clk(gclk));
	jdff dff_A_EY6ZkTN12_0(.dout(w_dff_A_thL9YslX9_0),.din(w_dff_A_EY6ZkTN12_0),.clk(gclk));
	jdff dff_A_7wF21ChK9_0(.dout(w_dff_A_EY6ZkTN12_0),.din(w_dff_A_7wF21ChK9_0),.clk(gclk));
	jdff dff_A_wzD724kr5_0(.dout(w_dff_A_7wF21ChK9_0),.din(w_dff_A_wzD724kr5_0),.clk(gclk));
	jdff dff_A_VPU98HRn1_0(.dout(w_dff_A_wzD724kr5_0),.din(w_dff_A_VPU98HRn1_0),.clk(gclk));
	jdff dff_A_We3bCPNw9_0(.dout(w_dff_A_VPU98HRn1_0),.din(w_dff_A_We3bCPNw9_0),.clk(gclk));
	jdff dff_A_FLRW1MjS4_0(.dout(w_n107_0[0]),.din(w_dff_A_FLRW1MjS4_0),.clk(gclk));
	jdff dff_A_C7hbJVIu8_0(.dout(w_dff_A_FLRW1MjS4_0),.din(w_dff_A_C7hbJVIu8_0),.clk(gclk));
	jdff dff_A_V4BXIRs30_0(.dout(w_dff_A_C7hbJVIu8_0),.din(w_dff_A_V4BXIRs30_0),.clk(gclk));
	jdff dff_A_0PJCXc3l6_0(.dout(w_dff_A_V4BXIRs30_0),.din(w_dff_A_0PJCXc3l6_0),.clk(gclk));
	jdff dff_A_SSyHuhK77_0(.dout(w_dff_A_0PJCXc3l6_0),.din(w_dff_A_SSyHuhK77_0),.clk(gclk));
	jdff dff_B_Jj7uKu7q3_2(.din(n107),.dout(w_dff_B_Jj7uKu7q3_2),.clk(gclk));
	jdff dff_B_4VdugBgu9_2(.din(w_dff_B_Jj7uKu7q3_2),.dout(w_dff_B_4VdugBgu9_2),.clk(gclk));
	jdff dff_B_r5HOOpVi9_2(.din(w_dff_B_4VdugBgu9_2),.dout(w_dff_B_r5HOOpVi9_2),.clk(gclk));
	jdff dff_B_gIGqkwep0_2(.din(w_dff_B_r5HOOpVi9_2),.dout(w_dff_B_gIGqkwep0_2),.clk(gclk));
	jdff dff_B_DzEb7Z7n0_2(.din(w_dff_B_gIGqkwep0_2),.dout(w_dff_B_DzEb7Z7n0_2),.clk(gclk));
	jdff dff_B_kGcL2mV18_2(.din(w_dff_B_DzEb7Z7n0_2),.dout(w_dff_B_kGcL2mV18_2),.clk(gclk));
	jdff dff_B_h679x01V9_2(.din(w_dff_B_kGcL2mV18_2),.dout(w_dff_B_h679x01V9_2),.clk(gclk));
	jdff dff_A_npfovwcA0_0(.dout(w_G73gat_0[0]),.din(w_dff_A_npfovwcA0_0),.clk(gclk));
	jdff dff_A_KNLGmZ9N0_0(.dout(w_dff_A_npfovwcA0_0),.din(w_dff_A_KNLGmZ9N0_0),.clk(gclk));
	jdff dff_A_u12ccG5M8_0(.dout(w_dff_A_KNLGmZ9N0_0),.din(w_dff_A_u12ccG5M8_0),.clk(gclk));
	jdff dff_A_WRMxSBoA1_0(.dout(w_dff_A_u12ccG5M8_0),.din(w_dff_A_WRMxSBoA1_0),.clk(gclk));
	jdff dff_A_JW9tXFPc7_0(.dout(w_dff_A_WRMxSBoA1_0),.din(w_dff_A_JW9tXFPc7_0),.clk(gclk));
	jdff dff_A_K9maBX633_0(.dout(w_dff_A_JW9tXFPc7_0),.din(w_dff_A_K9maBX633_0),.clk(gclk));
	jdff dff_A_GUuDysUB7_0(.dout(w_dff_A_K9maBX633_0),.din(w_dff_A_GUuDysUB7_0),.clk(gclk));
	jdff dff_A_BOA3bU9v4_0(.dout(w_dff_A_GUuDysUB7_0),.din(w_dff_A_BOA3bU9v4_0),.clk(gclk));
	jdff dff_A_I34zNpAM8_0(.dout(w_dff_A_BOA3bU9v4_0),.din(w_dff_A_I34zNpAM8_0),.clk(gclk));
	jdff dff_A_AIgkchZt2_0(.dout(w_dff_A_I34zNpAM8_0),.din(w_dff_A_AIgkchZt2_0),.clk(gclk));
	jdff dff_A_bRt1qN9Y2_0(.dout(w_dff_A_AIgkchZt2_0),.din(w_dff_A_bRt1qN9Y2_0),.clk(gclk));
	jdff dff_A_B6WMj8OW4_0(.dout(w_dff_A_bRt1qN9Y2_0),.din(w_dff_A_B6WMj8OW4_0),.clk(gclk));
	jdff dff_A_5IvxTNcM1_0(.dout(w_dff_A_B6WMj8OW4_0),.din(w_dff_A_5IvxTNcM1_0),.clk(gclk));
	jdff dff_A_D2AQoDto8_1(.dout(w_G73gat_0[1]),.din(w_dff_A_D2AQoDto8_1),.clk(gclk));
	jdff dff_A_F0JIs2ES0_1(.dout(w_dff_A_D2AQoDto8_1),.din(w_dff_A_F0JIs2ES0_1),.clk(gclk));
	jdff dff_A_qq3yqkYQ5_1(.dout(w_dff_A_F0JIs2ES0_1),.din(w_dff_A_qq3yqkYQ5_1),.clk(gclk));
	jdff dff_A_1GqXu33B7_1(.dout(w_dff_A_qq3yqkYQ5_1),.din(w_dff_A_1GqXu33B7_1),.clk(gclk));
	jdff dff_A_iYiCIsi58_1(.dout(w_dff_A_1GqXu33B7_1),.din(w_dff_A_iYiCIsi58_1),.clk(gclk));
	jdff dff_A_zn5Q2Ay87_1(.dout(w_dff_A_iYiCIsi58_1),.din(w_dff_A_zn5Q2Ay87_1),.clk(gclk));
	jdff dff_A_SfmIrGl77_1(.dout(w_dff_A_zn5Q2Ay87_1),.din(w_dff_A_SfmIrGl77_1),.clk(gclk));
	jdff dff_A_BvsG1iB14_1(.dout(w_dff_A_SfmIrGl77_1),.din(w_dff_A_BvsG1iB14_1),.clk(gclk));
	jdff dff_B_IJ05LnsU1_1(.din(n103),.dout(w_dff_B_IJ05LnsU1_1),.clk(gclk));
	jdff dff_B_ew6Sx7Ne9_1(.din(w_dff_B_IJ05LnsU1_1),.dout(w_dff_B_ew6Sx7Ne9_1),.clk(gclk));
	jdff dff_B_aXFrSv8w7_1(.din(w_dff_B_ew6Sx7Ne9_1),.dout(w_dff_B_aXFrSv8w7_1),.clk(gclk));
	jdff dff_B_7Zx3y7Us8_1(.din(w_dff_B_aXFrSv8w7_1),.dout(w_dff_B_7Zx3y7Us8_1),.clk(gclk));
	jdff dff_B_A9CJi3bf1_1(.din(w_dff_B_7Zx3y7Us8_1),.dout(w_dff_B_A9CJi3bf1_1),.clk(gclk));
	jdff dff_B_rIw6Z5jZ4_1(.din(w_dff_B_A9CJi3bf1_1),.dout(w_dff_B_rIw6Z5jZ4_1),.clk(gclk));
	jdff dff_B_skShDEEj8_1(.din(w_dff_B_rIw6Z5jZ4_1),.dout(w_dff_B_skShDEEj8_1),.clk(gclk));
	jdff dff_A_Mt602y425_0(.dout(w_G99gat_0[0]),.din(w_dff_A_Mt602y425_0),.clk(gclk));
	jdff dff_A_72bOw33v7_0(.dout(w_dff_A_Mt602y425_0),.din(w_dff_A_72bOw33v7_0),.clk(gclk));
	jdff dff_A_edKtgtQS9_0(.dout(w_dff_A_72bOw33v7_0),.din(w_dff_A_edKtgtQS9_0),.clk(gclk));
	jdff dff_A_CFuS4ITS1_0(.dout(w_dff_A_edKtgtQS9_0),.din(w_dff_A_CFuS4ITS1_0),.clk(gclk));
	jdff dff_A_WN3BflP03_0(.dout(w_dff_A_CFuS4ITS1_0),.din(w_dff_A_WN3BflP03_0),.clk(gclk));
	jdff dff_A_6BQ4Y8TJ5_0(.dout(w_dff_A_WN3BflP03_0),.din(w_dff_A_6BQ4Y8TJ5_0),.clk(gclk));
	jdff dff_A_2L1IILG65_0(.dout(w_dff_A_6BQ4Y8TJ5_0),.din(w_dff_A_2L1IILG65_0),.clk(gclk));
	jdff dff_A_Iv4WggU41_0(.dout(w_dff_A_2L1IILG65_0),.din(w_dff_A_Iv4WggU41_0),.clk(gclk));
	jdff dff_A_lelpZt550_1(.dout(w_G99gat_0[1]),.din(w_dff_A_lelpZt550_1),.clk(gclk));
	jdff dff_A_7xEU8tmF5_1(.dout(w_dff_A_lelpZt550_1),.din(w_dff_A_7xEU8tmF5_1),.clk(gclk));
	jdff dff_A_RkC3auJn0_1(.dout(w_dff_A_7xEU8tmF5_1),.din(w_dff_A_RkC3auJn0_1),.clk(gclk));
	jdff dff_A_X1aMSfV56_1(.dout(w_dff_A_RkC3auJn0_1),.din(w_dff_A_X1aMSfV56_1),.clk(gclk));
	jdff dff_A_lqQhWsMo4_1(.dout(w_dff_A_X1aMSfV56_1),.din(w_dff_A_lqQhWsMo4_1),.clk(gclk));
	jdff dff_A_CqUumgaR1_1(.dout(w_dff_A_lqQhWsMo4_1),.din(w_dff_A_CqUumgaR1_1),.clk(gclk));
	jdff dff_A_nJQwknpe5_1(.dout(w_dff_A_CqUumgaR1_1),.din(w_dff_A_nJQwknpe5_1),.clk(gclk));
	jdff dff_A_CYrxnjOJ4_1(.dout(w_dff_A_nJQwknpe5_1),.din(w_dff_A_CYrxnjOJ4_1),.clk(gclk));
	jdff dff_A_HHvFAjYp5_1(.dout(w_dff_A_CYrxnjOJ4_1),.din(w_dff_A_HHvFAjYp5_1),.clk(gclk));
	jdff dff_A_0LkbZkY76_1(.dout(w_dff_A_HHvFAjYp5_1),.din(w_dff_A_0LkbZkY76_1),.clk(gclk));
	jdff dff_A_VxKs87dm2_1(.dout(w_dff_A_0LkbZkY76_1),.din(w_dff_A_VxKs87dm2_1),.clk(gclk));
	jdff dff_A_Jy1b7IgE2_1(.dout(w_dff_A_VxKs87dm2_1),.din(w_dff_A_Jy1b7IgE2_1),.clk(gclk));
	jdff dff_A_zFpJtcqW2_1(.dout(w_dff_A_Jy1b7IgE2_1),.din(w_dff_A_zFpJtcqW2_1),.clk(gclk));
	jdff dff_A_pWXp4vsy2_0(.dout(w_n100_0[0]),.din(w_dff_A_pWXp4vsy2_0),.clk(gclk));
	jdff dff_A_sP9n6fSY2_0(.dout(w_dff_A_pWXp4vsy2_0),.din(w_dff_A_sP9n6fSY2_0),.clk(gclk));
	jdff dff_A_F9VmtyYp4_0(.dout(w_dff_A_sP9n6fSY2_0),.din(w_dff_A_F9VmtyYp4_0),.clk(gclk));
	jdff dff_A_lq5UdQm82_0(.dout(w_dff_A_F9VmtyYp4_0),.din(w_dff_A_lq5UdQm82_0),.clk(gclk));
	jdff dff_A_xf8KplPu3_0(.dout(w_dff_A_lq5UdQm82_0),.din(w_dff_A_xf8KplPu3_0),.clk(gclk));
	jdff dff_A_xqRTKSaT0_0(.dout(w_dff_A_xf8KplPu3_0),.din(w_dff_A_xqRTKSaT0_0),.clk(gclk));
	jdff dff_A_PUbLdDxi5_0(.dout(w_n98_0[0]),.din(w_dff_A_PUbLdDxi5_0),.clk(gclk));
	jdff dff_A_QBaKjAdo9_0(.dout(w_dff_A_PUbLdDxi5_0),.din(w_dff_A_QBaKjAdo9_0),.clk(gclk));
	jdff dff_A_x2bDx4899_0(.dout(w_dff_A_QBaKjAdo9_0),.din(w_dff_A_x2bDx4899_0),.clk(gclk));
	jdff dff_A_0vGZdjVW1_0(.dout(w_dff_A_x2bDx4899_0),.din(w_dff_A_0vGZdjVW1_0),.clk(gclk));
	jdff dff_A_bCX2syvd0_0(.dout(w_dff_A_0vGZdjVW1_0),.din(w_dff_A_bCX2syvd0_0),.clk(gclk));
	jdff dff_B_DaPTXosg2_2(.din(n98),.dout(w_dff_B_DaPTXosg2_2),.clk(gclk));
	jdff dff_B_ieMcNlbn2_2(.din(w_dff_B_DaPTXosg2_2),.dout(w_dff_B_ieMcNlbn2_2),.clk(gclk));
	jdff dff_B_5NCSWqyk2_2(.din(w_dff_B_ieMcNlbn2_2),.dout(w_dff_B_5NCSWqyk2_2),.clk(gclk));
	jdff dff_B_siupd1yj1_2(.din(w_dff_B_5NCSWqyk2_2),.dout(w_dff_B_siupd1yj1_2),.clk(gclk));
	jdff dff_B_5GhNvbGW6_2(.din(w_dff_B_siupd1yj1_2),.dout(w_dff_B_5GhNvbGW6_2),.clk(gclk));
	jdff dff_B_q0QwYz7j9_2(.din(w_dff_B_5GhNvbGW6_2),.dout(w_dff_B_q0QwYz7j9_2),.clk(gclk));
	jdff dff_B_BizbFXHl3_2(.din(w_dff_B_q0QwYz7j9_2),.dout(w_dff_B_BizbFXHl3_2),.clk(gclk));
	jdff dff_A_xbKsiBUT5_0(.dout(w_G8gat_0[0]),.din(w_dff_A_xbKsiBUT5_0),.clk(gclk));
	jdff dff_A_JEwyRUtL0_0(.dout(w_dff_A_xbKsiBUT5_0),.din(w_dff_A_JEwyRUtL0_0),.clk(gclk));
	jdff dff_A_3r4JC1MJ3_0(.dout(w_dff_A_JEwyRUtL0_0),.din(w_dff_A_3r4JC1MJ3_0),.clk(gclk));
	jdff dff_A_O0gGAdDj6_0(.dout(w_dff_A_3r4JC1MJ3_0),.din(w_dff_A_O0gGAdDj6_0),.clk(gclk));
	jdff dff_A_j1dnkyj72_0(.dout(w_dff_A_O0gGAdDj6_0),.din(w_dff_A_j1dnkyj72_0),.clk(gclk));
	jdff dff_A_HnFjcwHr2_0(.dout(w_dff_A_j1dnkyj72_0),.din(w_dff_A_HnFjcwHr2_0),.clk(gclk));
	jdff dff_A_J9WtIdK89_0(.dout(w_dff_A_HnFjcwHr2_0),.din(w_dff_A_J9WtIdK89_0),.clk(gclk));
	jdff dff_A_ujRWl8j44_0(.dout(w_dff_A_J9WtIdK89_0),.din(w_dff_A_ujRWl8j44_0),.clk(gclk));
	jdff dff_A_Eif8ZCn13_0(.dout(w_dff_A_ujRWl8j44_0),.din(w_dff_A_Eif8ZCn13_0),.clk(gclk));
	jdff dff_A_Ls9hETGk0_0(.dout(w_dff_A_Eif8ZCn13_0),.din(w_dff_A_Ls9hETGk0_0),.clk(gclk));
	jdff dff_A_8uf4SsJY1_0(.dout(w_dff_A_Ls9hETGk0_0),.din(w_dff_A_8uf4SsJY1_0),.clk(gclk));
	jdff dff_A_ya1dKjcZ0_0(.dout(w_dff_A_8uf4SsJY1_0),.din(w_dff_A_ya1dKjcZ0_0),.clk(gclk));
	jdff dff_A_zvrtZD2z1_0(.dout(w_dff_A_ya1dKjcZ0_0),.din(w_dff_A_zvrtZD2z1_0),.clk(gclk));
	jdff dff_A_j31M95Bd6_1(.dout(w_G8gat_0[1]),.din(w_dff_A_j31M95Bd6_1),.clk(gclk));
	jdff dff_A_cTv2D6Mn4_1(.dout(w_dff_A_j31M95Bd6_1),.din(w_dff_A_cTv2D6Mn4_1),.clk(gclk));
	jdff dff_A_1Ath8SQi0_1(.dout(w_dff_A_cTv2D6Mn4_1),.din(w_dff_A_1Ath8SQi0_1),.clk(gclk));
	jdff dff_A_TIygiPDq1_1(.dout(w_dff_A_1Ath8SQi0_1),.din(w_dff_A_TIygiPDq1_1),.clk(gclk));
	jdff dff_A_6Jt16Kt93_1(.dout(w_dff_A_TIygiPDq1_1),.din(w_dff_A_6Jt16Kt93_1),.clk(gclk));
	jdff dff_A_i5Bt9W5t0_1(.dout(w_dff_A_6Jt16Kt93_1),.din(w_dff_A_i5Bt9W5t0_1),.clk(gclk));
	jdff dff_A_m2iUUgfu3_1(.dout(w_dff_A_i5Bt9W5t0_1),.din(w_dff_A_m2iUUgfu3_1),.clk(gclk));
	jdff dff_A_gXl3cTPm5_1(.dout(w_dff_A_m2iUUgfu3_1),.din(w_dff_A_gXl3cTPm5_1),.clk(gclk));
	jdff dff_A_8dUrqxJt2_0(.dout(w_n96_0[0]),.din(w_dff_A_8dUrqxJt2_0),.clk(gclk));
	jdff dff_A_xbuxGv9b1_0(.dout(w_dff_A_8dUrqxJt2_0),.din(w_dff_A_xbuxGv9b1_0),.clk(gclk));
	jdff dff_A_Ho34elWX7_0(.dout(w_dff_A_xbuxGv9b1_0),.din(w_dff_A_Ho34elWX7_0),.clk(gclk));
	jdff dff_A_QVC2PP3K9_0(.dout(w_dff_A_Ho34elWX7_0),.din(w_dff_A_QVC2PP3K9_0),.clk(gclk));
	jdff dff_A_vA50aHIf9_0(.dout(w_dff_A_QVC2PP3K9_0),.din(w_dff_A_vA50aHIf9_0),.clk(gclk));
	jdff dff_A_NfiY4DDd3_0(.dout(w_dff_A_vA50aHIf9_0),.din(w_dff_A_NfiY4DDd3_0),.clk(gclk));
	jdff dff_B_9Upy40qx2_1(.din(n76),.dout(w_dff_B_9Upy40qx2_1),.clk(gclk));
	jdff dff_B_b5MS3O9c2_1(.din(n81),.dout(w_dff_B_b5MS3O9c2_1),.clk(gclk));
	jdff dff_A_8irem2iX5_0(.dout(w_n89_0[0]),.din(w_dff_A_8irem2iX5_0),.clk(gclk));
	jdff dff_A_eRB3XE5l9_0(.dout(w_dff_A_8irem2iX5_0),.din(w_dff_A_eRB3XE5l9_0),.clk(gclk));
	jdff dff_A_FfMnSgAs2_0(.dout(w_dff_A_eRB3XE5l9_0),.din(w_dff_A_FfMnSgAs2_0),.clk(gclk));
	jdff dff_A_mGhUST8d8_0(.dout(w_dff_A_FfMnSgAs2_0),.din(w_dff_A_mGhUST8d8_0),.clk(gclk));
	jdff dff_A_rd5Omw5k0_0(.dout(w_dff_A_mGhUST8d8_0),.din(w_dff_A_rd5Omw5k0_0),.clk(gclk));
	jdff dff_A_pb3yzhzd3_0(.dout(w_dff_A_rd5Omw5k0_0),.din(w_dff_A_pb3yzhzd3_0),.clk(gclk));
	jdff dff_A_DGdJol9C3_0(.dout(w_n84_0[0]),.din(w_dff_A_DGdJol9C3_0),.clk(gclk));
	jdff dff_A_7FLBCUWu0_0(.dout(w_dff_A_DGdJol9C3_0),.din(w_dff_A_7FLBCUWu0_0),.clk(gclk));
	jdff dff_A_YfDKkGva9_0(.dout(w_dff_A_7FLBCUWu0_0),.din(w_dff_A_YfDKkGva9_0),.clk(gclk));
	jdff dff_A_XjLcVCgl3_0(.dout(w_dff_A_YfDKkGva9_0),.din(w_dff_A_XjLcVCgl3_0),.clk(gclk));
	jdff dff_A_A882PPX87_0(.dout(w_dff_A_XjLcVCgl3_0),.din(w_dff_A_A882PPX87_0),.clk(gclk));
	jdff dff_A_jRPjoRYT8_0(.dout(w_dff_A_A882PPX87_0),.din(w_dff_A_jRPjoRYT8_0),.clk(gclk));
	jdff dff_A_WzpsQQq57_0(.dout(w_n82_0[0]),.din(w_dff_A_WzpsQQq57_0),.clk(gclk));
	jdff dff_A_uHGqXqSF9_0(.dout(w_dff_A_WzpsQQq57_0),.din(w_dff_A_uHGqXqSF9_0),.clk(gclk));
	jdff dff_A_IxigYVKC4_0(.dout(w_dff_A_uHGqXqSF9_0),.din(w_dff_A_IxigYVKC4_0),.clk(gclk));
	jdff dff_A_Cob9RQFo2_0(.dout(w_dff_A_IxigYVKC4_0),.din(w_dff_A_Cob9RQFo2_0),.clk(gclk));
	jdff dff_A_JSSKEe3r4_0(.dout(w_dff_A_Cob9RQFo2_0),.din(w_dff_A_JSSKEe3r4_0),.clk(gclk));
	jdff dff_A_2L284IBN8_0(.dout(w_dff_A_JSSKEe3r4_0),.din(w_dff_A_2L284IBN8_0),.clk(gclk));
	jdff dff_A_sbiRWCr15_0(.dout(w_n79_0[0]),.din(w_dff_A_sbiRWCr15_0),.clk(gclk));
	jdff dff_A_u6jPLFcV4_0(.dout(w_dff_A_sbiRWCr15_0),.din(w_dff_A_u6jPLFcV4_0),.clk(gclk));
	jdff dff_A_GYDNLt7Q0_0(.dout(w_dff_A_u6jPLFcV4_0),.din(w_dff_A_GYDNLt7Q0_0),.clk(gclk));
	jdff dff_A_Xdcuj0cd8_0(.dout(w_dff_A_GYDNLt7Q0_0),.din(w_dff_A_Xdcuj0cd8_0),.clk(gclk));
	jdff dff_A_yYj7vxl72_0(.dout(w_dff_A_Xdcuj0cd8_0),.din(w_dff_A_yYj7vxl72_0),.clk(gclk));
	jdff dff_A_6hUcOWcz2_0(.dout(w_dff_A_yYj7vxl72_0),.din(w_dff_A_6hUcOWcz2_0),.clk(gclk));
	jdff dff_A_HygIf3FV6_0(.dout(w_n78_0[0]),.din(w_dff_A_HygIf3FV6_0),.clk(gclk));
	jdff dff_A_z1jmVMXQ2_0(.dout(w_dff_A_HygIf3FV6_0),.din(w_dff_A_z1jmVMXQ2_0),.clk(gclk));
	jdff dff_A_Gs98PXer8_0(.dout(w_dff_A_z1jmVMXQ2_0),.din(w_dff_A_Gs98PXer8_0),.clk(gclk));
	jdff dff_A_LcucVDKL2_0(.dout(w_dff_A_Gs98PXer8_0),.din(w_dff_A_LcucVDKL2_0),.clk(gclk));
	jdff dff_A_HXtgFlgA3_0(.dout(w_n77_0[0]),.din(w_dff_A_HXtgFlgA3_0),.clk(gclk));
	jdff dff_A_9MrS5y7K5_0(.dout(w_dff_A_HXtgFlgA3_0),.din(w_dff_A_9MrS5y7K5_0),.clk(gclk));
	jdff dff_A_hI03JWLr2_0(.dout(w_dff_A_9MrS5y7K5_0),.din(w_dff_A_hI03JWLr2_0),.clk(gclk));
	jdff dff_A_0ZCutWDk7_0(.dout(w_dff_A_hI03JWLr2_0),.din(w_dff_A_0ZCutWDk7_0),.clk(gclk));
	jdff dff_A_dYRBYl1F6_0(.dout(w_dff_A_0ZCutWDk7_0),.din(w_dff_A_dYRBYl1F6_0),.clk(gclk));
	jdff dff_A_e5q9SpBs2_0(.dout(w_dff_A_dYRBYl1F6_0),.din(w_dff_A_e5q9SpBs2_0),.clk(gclk));
	jdff dff_A_SoPJwzNr1_0(.dout(w_n73_0[0]),.din(w_dff_A_SoPJwzNr1_0),.clk(gclk));
	jdff dff_A_Sr1VNf7C3_0(.dout(w_dff_A_SoPJwzNr1_0),.din(w_dff_A_Sr1VNf7C3_0),.clk(gclk));
	jdff dff_A_vBexnnKd3_0(.dout(w_dff_A_Sr1VNf7C3_0),.din(w_dff_A_vBexnnKd3_0),.clk(gclk));
	jdff dff_A_BqZu15C15_0(.dout(w_dff_A_vBexnnKd3_0),.din(w_dff_A_BqZu15C15_0),.clk(gclk));
	jdff dff_A_ArlNSiEQ7_0(.dout(w_dff_A_BqZu15C15_0),.din(w_dff_A_ArlNSiEQ7_0),.clk(gclk));
	jdff dff_A_S8vp1hBI6_0(.dout(w_dff_A_ArlNSiEQ7_0),.din(w_dff_A_S8vp1hBI6_0),.clk(gclk));
	jdff dff_A_TpYjo0lD4_0(.dout(w_n72_0[0]),.din(w_dff_A_TpYjo0lD4_0),.clk(gclk));
	jdff dff_A_ouHNtJo78_0(.dout(w_dff_A_TpYjo0lD4_0),.din(w_dff_A_ouHNtJo78_0),.clk(gclk));
	jdff dff_A_cGt8BaJC9_0(.dout(w_dff_A_ouHNtJo78_0),.din(w_dff_A_cGt8BaJC9_0),.clk(gclk));
	jdff dff_A_sDxS30GO9_0(.dout(w_dff_A_cGt8BaJC9_0),.din(w_dff_A_sDxS30GO9_0),.clk(gclk));
	jdff dff_A_AppzSTfM1_0(.dout(w_n71_0[0]),.din(w_dff_A_AppzSTfM1_0),.clk(gclk));
	jdff dff_A_UcvP5oGh2_0(.dout(w_dff_A_AppzSTfM1_0),.din(w_dff_A_UcvP5oGh2_0),.clk(gclk));
	jdff dff_A_JX7moqiu4_0(.dout(w_dff_A_UcvP5oGh2_0),.din(w_dff_A_JX7moqiu4_0),.clk(gclk));
	jdff dff_A_xEFovKgy0_0(.dout(w_dff_A_JX7moqiu4_0),.din(w_dff_A_xEFovKgy0_0),.clk(gclk));
	jdff dff_A_UJyy5Pf67_0(.dout(w_dff_A_xEFovKgy0_0),.din(w_dff_A_UJyy5Pf67_0),.clk(gclk));
	jdff dff_A_7jIEFFPy1_0(.dout(w_dff_A_UJyy5Pf67_0),.din(w_dff_A_7jIEFFPy1_0),.clk(gclk));
	jdff dff_A_H27ZvLKe0_0(.dout(w_n69_0[0]),.din(w_dff_A_H27ZvLKe0_0),.clk(gclk));
	jdff dff_A_RmbDk14d7_0(.dout(w_dff_A_H27ZvLKe0_0),.din(w_dff_A_RmbDk14d7_0),.clk(gclk));
	jdff dff_A_sE9D6LVt2_0(.dout(w_dff_A_RmbDk14d7_0),.din(w_dff_A_sE9D6LVt2_0),.clk(gclk));
	jdff dff_A_2SuVzH7c7_0(.dout(w_dff_A_sE9D6LVt2_0),.din(w_dff_A_2SuVzH7c7_0),.clk(gclk));
	jdff dff_A_LwcZ7WBl8_0(.dout(w_dff_A_2SuVzH7c7_0),.din(w_dff_A_LwcZ7WBl8_0),.clk(gclk));
	jdff dff_B_2QrGcgoq9_2(.din(n69),.dout(w_dff_B_2QrGcgoq9_2),.clk(gclk));
	jdff dff_B_jk43HwGo6_2(.din(w_dff_B_2QrGcgoq9_2),.dout(w_dff_B_jk43HwGo6_2),.clk(gclk));
	jdff dff_B_FL6lkWnD8_2(.din(w_dff_B_jk43HwGo6_2),.dout(w_dff_B_FL6lkWnD8_2),.clk(gclk));
	jdff dff_B_luMftctM9_2(.din(w_dff_B_FL6lkWnD8_2),.dout(w_dff_B_luMftctM9_2),.clk(gclk));
	jdff dff_B_WSCq9NLs6_2(.din(w_dff_B_luMftctM9_2),.dout(w_dff_B_WSCq9NLs6_2),.clk(gclk));
	jdff dff_B_Vb5fUudZ6_2(.din(w_dff_B_WSCq9NLs6_2),.dout(w_dff_B_Vb5fUudZ6_2),.clk(gclk));
	jdff dff_B_6Fxb3ivR9_2(.din(w_dff_B_Vb5fUudZ6_2),.dout(w_dff_B_6Fxb3ivR9_2),.clk(gclk));
	jdff dff_A_L28j0QWF9_0(.dout(w_G112gat_0[0]),.din(w_dff_A_L28j0QWF9_0),.clk(gclk));
	jdff dff_A_rrbJJwxk8_0(.dout(w_dff_A_L28j0QWF9_0),.din(w_dff_A_rrbJJwxk8_0),.clk(gclk));
	jdff dff_A_nGzq8QVI2_0(.dout(w_dff_A_rrbJJwxk8_0),.din(w_dff_A_nGzq8QVI2_0),.clk(gclk));
	jdff dff_A_6AfqpOUm1_0(.dout(w_dff_A_nGzq8QVI2_0),.din(w_dff_A_6AfqpOUm1_0),.clk(gclk));
	jdff dff_A_eBqsggGa9_0(.dout(w_dff_A_6AfqpOUm1_0),.din(w_dff_A_eBqsggGa9_0),.clk(gclk));
	jdff dff_A_ckHjfnbY0_0(.dout(w_dff_A_eBqsggGa9_0),.din(w_dff_A_ckHjfnbY0_0),.clk(gclk));
	jdff dff_A_qIQfrjFk5_0(.dout(w_dff_A_ckHjfnbY0_0),.din(w_dff_A_qIQfrjFk5_0),.clk(gclk));
	jdff dff_A_2axH7m6q0_0(.dout(w_dff_A_qIQfrjFk5_0),.din(w_dff_A_2axH7m6q0_0),.clk(gclk));
	jdff dff_A_HLkrLkLw5_0(.dout(w_dff_A_2axH7m6q0_0),.din(w_dff_A_HLkrLkLw5_0),.clk(gclk));
	jdff dff_A_99P4KDl67_0(.dout(w_dff_A_HLkrLkLw5_0),.din(w_dff_A_99P4KDl67_0),.clk(gclk));
	jdff dff_A_AcqvjvjU5_0(.dout(w_dff_A_99P4KDl67_0),.din(w_dff_A_AcqvjvjU5_0),.clk(gclk));
	jdff dff_A_x8RWZbBH7_0(.dout(w_dff_A_AcqvjvjU5_0),.din(w_dff_A_x8RWZbBH7_0),.clk(gclk));
	jdff dff_A_pegk6xgq3_0(.dout(w_dff_A_x8RWZbBH7_0),.din(w_dff_A_pegk6xgq3_0),.clk(gclk));
	jdff dff_A_7qSynyHz9_1(.dout(w_G112gat_0[1]),.din(w_dff_A_7qSynyHz9_1),.clk(gclk));
	jdff dff_A_dcrecD3A9_1(.dout(w_dff_A_7qSynyHz9_1),.din(w_dff_A_dcrecD3A9_1),.clk(gclk));
	jdff dff_A_qdw1jxH20_1(.dout(w_dff_A_dcrecD3A9_1),.din(w_dff_A_qdw1jxH20_1),.clk(gclk));
	jdff dff_A_AHavIrtC5_1(.dout(w_dff_A_qdw1jxH20_1),.din(w_dff_A_AHavIrtC5_1),.clk(gclk));
	jdff dff_A_tKobfIKP3_1(.dout(w_dff_A_AHavIrtC5_1),.din(w_dff_A_tKobfIKP3_1),.clk(gclk));
	jdff dff_A_dUMxbQmC7_1(.dout(w_dff_A_tKobfIKP3_1),.din(w_dff_A_dUMxbQmC7_1),.clk(gclk));
	jdff dff_A_5mEYVwFM4_1(.dout(w_dff_A_dUMxbQmC7_1),.din(w_dff_A_5mEYVwFM4_1),.clk(gclk));
	jdff dff_A_zZ0sUR6U8_1(.dout(w_dff_A_5mEYVwFM4_1),.din(w_dff_A_zZ0sUR6U8_1),.clk(gclk));
	jdff dff_A_eGX8fAJW5_1(.dout(w_n139_0[1]),.din(w_dff_A_eGX8fAJW5_1),.clk(gclk));
	jdff dff_A_nOxwyhP22_1(.dout(w_dff_A_eGX8fAJW5_1),.din(w_dff_A_nOxwyhP22_1),.clk(gclk));
	jdff dff_A_ByprSnQp6_1(.dout(w_dff_A_nOxwyhP22_1),.din(w_dff_A_ByprSnQp6_1),.clk(gclk));
	jdff dff_A_jolfjana6_1(.dout(w_dff_A_ByprSnQp6_1),.din(w_dff_A_jolfjana6_1),.clk(gclk));
	jdff dff_A_72BsNdOV6_1(.dout(w_dff_A_jolfjana6_1),.din(w_dff_A_72BsNdOV6_1),.clk(gclk));
	jdff dff_A_C2h2upGr0_1(.dout(w_dff_A_72BsNdOV6_1),.din(w_dff_A_C2h2upGr0_1),.clk(gclk));
	jdff dff_B_ZTmTrgcu9_1(.din(n50),.dout(w_dff_B_ZTmTrgcu9_1),.clk(gclk));
	jdff dff_B_I9OydJlB7_1(.din(n55),.dout(w_dff_B_I9OydJlB7_1),.clk(gclk));
	jdff dff_A_m0sInY1m1_0(.dout(w_G4gat_0[0]),.din(w_dff_A_m0sInY1m1_0),.clk(gclk));
	jdff dff_A_3Dc8BMAJ9_0(.dout(w_dff_A_m0sInY1m1_0),.din(w_dff_A_3Dc8BMAJ9_0),.clk(gclk));
	jdff dff_A_nrw18G6x9_0(.dout(w_dff_A_3Dc8BMAJ9_0),.din(w_dff_A_nrw18G6x9_0),.clk(gclk));
	jdff dff_A_ouLpvPEl1_0(.dout(w_dff_A_nrw18G6x9_0),.din(w_dff_A_ouLpvPEl1_0),.clk(gclk));
	jdff dff_A_dZSeG2ZM7_0(.dout(w_dff_A_ouLpvPEl1_0),.din(w_dff_A_dZSeG2ZM7_0),.clk(gclk));
	jdff dff_A_1WMRYPC81_0(.dout(w_dff_A_dZSeG2ZM7_0),.din(w_dff_A_1WMRYPC81_0),.clk(gclk));
	jdff dff_A_tpsFSx6J9_0(.dout(w_dff_A_1WMRYPC81_0),.din(w_dff_A_tpsFSx6J9_0),.clk(gclk));
	jdff dff_A_7F2z2dxM4_2(.dout(w_G4gat_0[2]),.din(w_dff_A_7F2z2dxM4_2),.clk(gclk));
	jdff dff_A_60Y4Uhit5_0(.dout(w_n63_0[0]),.din(w_dff_A_60Y4Uhit5_0),.clk(gclk));
	jdff dff_A_MuYsHldj5_0(.dout(w_dff_A_60Y4Uhit5_0),.din(w_dff_A_MuYsHldj5_0),.clk(gclk));
	jdff dff_A_G1JoxGCM6_0(.dout(w_dff_A_MuYsHldj5_0),.din(w_dff_A_G1JoxGCM6_0),.clk(gclk));
	jdff dff_A_RFEZJnl40_0(.dout(w_dff_A_G1JoxGCM6_0),.din(w_dff_A_RFEZJnl40_0),.clk(gclk));
	jdff dff_A_GkI62Qcc3_0(.dout(w_dff_A_RFEZJnl40_0),.din(w_dff_A_GkI62Qcc3_0),.clk(gclk));
	jdff dff_A_lo6C9lXj9_0(.dout(w_G1gat_0[0]),.din(w_dff_A_lo6C9lXj9_0),.clk(gclk));
	jdff dff_A_UwSJewNF0_0(.dout(w_dff_A_lo6C9lXj9_0),.din(w_dff_A_UwSJewNF0_0),.clk(gclk));
	jdff dff_A_m9Pfbm2e3_0(.dout(w_dff_A_UwSJewNF0_0),.din(w_dff_A_m9Pfbm2e3_0),.clk(gclk));
	jdff dff_A_iJCxKET37_0(.dout(w_dff_A_m9Pfbm2e3_0),.din(w_dff_A_iJCxKET37_0),.clk(gclk));
	jdff dff_A_w0JUjoKL0_0(.dout(w_dff_A_iJCxKET37_0),.din(w_dff_A_w0JUjoKL0_0),.clk(gclk));
	jdff dff_A_kvUPm0Tm4_0(.dout(w_dff_A_w0JUjoKL0_0),.din(w_dff_A_kvUPm0Tm4_0),.clk(gclk));
	jdff dff_A_iqGXefEK4_1(.dout(w_G1gat_0[1]),.din(w_dff_A_iqGXefEK4_1),.clk(gclk));
	jdff dff_A_m1Rysvbr1_0(.dout(w_n61_0[0]),.din(w_dff_A_m1Rysvbr1_0),.clk(gclk));
	jdff dff_A_Gousxmok7_0(.dout(w_dff_A_m1Rysvbr1_0),.din(w_dff_A_Gousxmok7_0),.clk(gclk));
	jdff dff_A_JB0l18RT8_0(.dout(w_dff_A_Gousxmok7_0),.din(w_dff_A_JB0l18RT8_0),.clk(gclk));
	jdff dff_A_y949gqVK7_0(.dout(w_dff_A_JB0l18RT8_0),.din(w_dff_A_y949gqVK7_0),.clk(gclk));
	jdff dff_A_zAKZk9uM8_0(.dout(w_dff_A_y949gqVK7_0),.din(w_dff_A_zAKZk9uM8_0),.clk(gclk));
	jdff dff_A_aYsJW7np3_0(.dout(w_G89gat_0[0]),.din(w_dff_A_aYsJW7np3_0),.clk(gclk));
	jdff dff_A_XftsmayI7_0(.dout(w_dff_A_aYsJW7np3_0),.din(w_dff_A_XftsmayI7_0),.clk(gclk));
	jdff dff_A_5nWOZrJr0_0(.dout(w_dff_A_XftsmayI7_0),.din(w_dff_A_5nWOZrJr0_0),.clk(gclk));
	jdff dff_A_Z9GL0bfx9_0(.dout(w_dff_A_5nWOZrJr0_0),.din(w_dff_A_Z9GL0bfx9_0),.clk(gclk));
	jdff dff_A_RUtWmEfy5_0(.dout(w_dff_A_Z9GL0bfx9_0),.din(w_dff_A_RUtWmEfy5_0),.clk(gclk));
	jdff dff_A_tsCGXlx34_0(.dout(w_dff_A_RUtWmEfy5_0),.din(w_dff_A_tsCGXlx34_0),.clk(gclk));
	jdff dff_A_Q3mVMiD52_1(.dout(w_G89gat_0[1]),.din(w_dff_A_Q3mVMiD52_1),.clk(gclk));
	jdff dff_A_xqVvE7FQ0_0(.dout(w_G56gat_0[0]),.din(w_dff_A_xqVvE7FQ0_0),.clk(gclk));
	jdff dff_A_SzlcahD08_0(.dout(w_dff_A_xqVvE7FQ0_0),.din(w_dff_A_SzlcahD08_0),.clk(gclk));
	jdff dff_A_mLsCDeGM0_0(.dout(w_dff_A_SzlcahD08_0),.din(w_dff_A_mLsCDeGM0_0),.clk(gclk));
	jdff dff_A_9TsmqOJa7_0(.dout(w_dff_A_mLsCDeGM0_0),.din(w_dff_A_9TsmqOJa7_0),.clk(gclk));
	jdff dff_A_aKxb2sx62_0(.dout(w_dff_A_9TsmqOJa7_0),.din(w_dff_A_aKxb2sx62_0),.clk(gclk));
	jdff dff_A_EzaegSGS2_0(.dout(w_dff_A_aKxb2sx62_0),.din(w_dff_A_EzaegSGS2_0),.clk(gclk));
	jdff dff_A_5Rl7pigT2_0(.dout(w_dff_A_EzaegSGS2_0),.din(w_dff_A_5Rl7pigT2_0),.clk(gclk));
	jdff dff_A_ZzxpXh6n8_2(.dout(w_G56gat_0[2]),.din(w_dff_A_ZzxpXh6n8_2),.clk(gclk));
	jdff dff_A_AfpWvbmb9_0(.dout(w_n58_0[0]),.din(w_dff_A_AfpWvbmb9_0),.clk(gclk));
	jdff dff_A_Du2r85SN2_0(.dout(w_dff_A_AfpWvbmb9_0),.din(w_dff_A_Du2r85SN2_0),.clk(gclk));
	jdff dff_A_3ImWQwDu0_0(.dout(w_dff_A_Du2r85SN2_0),.din(w_dff_A_3ImWQwDu0_0),.clk(gclk));
	jdff dff_A_o3lMAH8V8_0(.dout(w_dff_A_3ImWQwDu0_0),.din(w_dff_A_o3lMAH8V8_0),.clk(gclk));
	jdff dff_A_oqonIYtI2_0(.dout(w_dff_A_o3lMAH8V8_0),.din(w_dff_A_oqonIYtI2_0),.clk(gclk));
	jdff dff_A_M1ZIXeKr5_0(.dout(w_G50gat_0[0]),.din(w_dff_A_M1ZIXeKr5_0),.clk(gclk));
	jdff dff_A_OWM6QZ776_0(.dout(w_dff_A_M1ZIXeKr5_0),.din(w_dff_A_OWM6QZ776_0),.clk(gclk));
	jdff dff_A_oQFHcsza7_0(.dout(w_dff_A_OWM6QZ776_0),.din(w_dff_A_oQFHcsza7_0),.clk(gclk));
	jdff dff_A_PKQIMobn7_0(.dout(w_dff_A_oQFHcsza7_0),.din(w_dff_A_PKQIMobn7_0),.clk(gclk));
	jdff dff_A_GSoTnHDN7_0(.dout(w_dff_A_PKQIMobn7_0),.din(w_dff_A_GSoTnHDN7_0),.clk(gclk));
	jdff dff_A_eWfgcqh78_0(.dout(w_dff_A_GSoTnHDN7_0),.din(w_dff_A_eWfgcqh78_0),.clk(gclk));
	jdff dff_A_RlI2Qcna3_1(.dout(w_G50gat_0[1]),.din(w_dff_A_RlI2Qcna3_1),.clk(gclk));
	jdff dff_A_7MrcKX5J9_0(.dout(w_G108gat_0[0]),.din(w_dff_A_7MrcKX5J9_0),.clk(gclk));
	jdff dff_A_WImJVBCU5_0(.dout(w_dff_A_7MrcKX5J9_0),.din(w_dff_A_WImJVBCU5_0),.clk(gclk));
	jdff dff_A_XS8WfAbQ8_0(.dout(w_dff_A_WImJVBCU5_0),.din(w_dff_A_XS8WfAbQ8_0),.clk(gclk));
	jdff dff_A_oAuVrjTh2_0(.dout(w_dff_A_XS8WfAbQ8_0),.din(w_dff_A_oAuVrjTh2_0),.clk(gclk));
	jdff dff_A_wTo6EMEo6_0(.dout(w_dff_A_oAuVrjTh2_0),.din(w_dff_A_wTo6EMEo6_0),.clk(gclk));
	jdff dff_A_myFTa8io4_0(.dout(w_dff_A_wTo6EMEo6_0),.din(w_dff_A_myFTa8io4_0),.clk(gclk));
	jdff dff_A_8oZTMSvm4_0(.dout(w_dff_A_myFTa8io4_0),.din(w_dff_A_8oZTMSvm4_0),.clk(gclk));
	jdff dff_A_PSQlRAdH8_2(.dout(w_G108gat_0[2]),.din(w_dff_A_PSQlRAdH8_2),.clk(gclk));
	jdff dff_A_HjkXD14a0_0(.dout(w_n56_0[0]),.din(w_dff_A_HjkXD14a0_0),.clk(gclk));
	jdff dff_A_MdplED1k8_0(.dout(w_dff_A_HjkXD14a0_0),.din(w_dff_A_MdplED1k8_0),.clk(gclk));
	jdff dff_A_vGlJWgTm6_0(.dout(w_dff_A_MdplED1k8_0),.din(w_dff_A_vGlJWgTm6_0),.clk(gclk));
	jdff dff_A_yDlyhauR5_0(.dout(w_dff_A_vGlJWgTm6_0),.din(w_dff_A_yDlyhauR5_0),.clk(gclk));
	jdff dff_A_MoIFUcYl8_0(.dout(w_dff_A_yDlyhauR5_0),.din(w_dff_A_MoIFUcYl8_0),.clk(gclk));
	jdff dff_A_cylKugpA0_0(.dout(w_G102gat_0[0]),.din(w_dff_A_cylKugpA0_0),.clk(gclk));
	jdff dff_A_3gdH3ebS3_0(.dout(w_dff_A_cylKugpA0_0),.din(w_dff_A_3gdH3ebS3_0),.clk(gclk));
	jdff dff_A_2qbSh4JH6_0(.dout(w_dff_A_3gdH3ebS3_0),.din(w_dff_A_2qbSh4JH6_0),.clk(gclk));
	jdff dff_A_nNliNcVk0_0(.dout(w_dff_A_2qbSh4JH6_0),.din(w_dff_A_nNliNcVk0_0),.clk(gclk));
	jdff dff_A_UqHDisAR2_0(.dout(w_dff_A_nNliNcVk0_0),.din(w_dff_A_UqHDisAR2_0),.clk(gclk));
	jdff dff_A_yqszvjhP7_0(.dout(w_dff_A_UqHDisAR2_0),.din(w_dff_A_yqszvjhP7_0),.clk(gclk));
	jdff dff_A_fZAokQjO4_1(.dout(w_G102gat_0[1]),.din(w_dff_A_fZAokQjO4_1),.clk(gclk));
	jdff dff_A_gmylrXXx0_0(.dout(w_G69gat_0[0]),.din(w_dff_A_gmylrXXx0_0),.clk(gclk));
	jdff dff_A_0fgqE8Kz5_0(.dout(w_dff_A_gmylrXXx0_0),.din(w_dff_A_0fgqE8Kz5_0),.clk(gclk));
	jdff dff_A_fy5GKzb95_0(.dout(w_dff_A_0fgqE8Kz5_0),.din(w_dff_A_fy5GKzb95_0),.clk(gclk));
	jdff dff_A_PSCNUDYL1_0(.dout(w_dff_A_fy5GKzb95_0),.din(w_dff_A_PSCNUDYL1_0),.clk(gclk));
	jdff dff_A_B8bZDcuL7_0(.dout(w_dff_A_PSCNUDYL1_0),.din(w_dff_A_B8bZDcuL7_0),.clk(gclk));
	jdff dff_A_t8vsKhgU5_0(.dout(w_dff_A_B8bZDcuL7_0),.din(w_dff_A_t8vsKhgU5_0),.clk(gclk));
	jdff dff_A_MerAvAjZ2_0(.dout(w_dff_A_t8vsKhgU5_0),.din(w_dff_A_MerAvAjZ2_0),.clk(gclk));
	jdff dff_A_feB0LyTG2_2(.dout(w_G69gat_0[2]),.din(w_dff_A_feB0LyTG2_2),.clk(gclk));
	jdff dff_A_B6CDKI960_0(.dout(w_n53_0[0]),.din(w_dff_A_B6CDKI960_0),.clk(gclk));
	jdff dff_A_xKnT3vzv1_0(.dout(w_dff_A_B6CDKI960_0),.din(w_dff_A_xKnT3vzv1_0),.clk(gclk));
	jdff dff_A_SSZHLRx26_0(.dout(w_dff_A_xKnT3vzv1_0),.din(w_dff_A_SSZHLRx26_0),.clk(gclk));
	jdff dff_A_kr4MV6vP6_0(.dout(w_dff_A_SSZHLRx26_0),.din(w_dff_A_kr4MV6vP6_0),.clk(gclk));
	jdff dff_A_Y6Is4uHB3_0(.dout(w_dff_A_kr4MV6vP6_0),.din(w_dff_A_Y6Is4uHB3_0),.clk(gclk));
	jdff dff_A_UQ3rpyYD5_0(.dout(w_G63gat_0[0]),.din(w_dff_A_UQ3rpyYD5_0),.clk(gclk));
	jdff dff_A_7RxetT275_0(.dout(w_dff_A_UQ3rpyYD5_0),.din(w_dff_A_7RxetT275_0),.clk(gclk));
	jdff dff_A_xGO0DJLT6_0(.dout(w_dff_A_7RxetT275_0),.din(w_dff_A_xGO0DJLT6_0),.clk(gclk));
	jdff dff_A_RvGw6Mad9_0(.dout(w_dff_A_xGO0DJLT6_0),.din(w_dff_A_RvGw6Mad9_0),.clk(gclk));
	jdff dff_A_42MKd7dj8_0(.dout(w_dff_A_RvGw6Mad9_0),.din(w_dff_A_42MKd7dj8_0),.clk(gclk));
	jdff dff_A_JVwcaE8v5_0(.dout(w_dff_A_42MKd7dj8_0),.din(w_dff_A_JVwcaE8v5_0),.clk(gclk));
	jdff dff_A_SyCFXrVg8_1(.dout(w_G63gat_0[1]),.din(w_dff_A_SyCFXrVg8_1),.clk(gclk));
	jdff dff_A_fgJvJHUp2_0(.dout(w_n52_0[0]),.din(w_dff_A_fgJvJHUp2_0),.clk(gclk));
	jdff dff_A_pjuNTLqz7_0(.dout(w_dff_A_fgJvJHUp2_0),.din(w_dff_A_pjuNTLqz7_0),.clk(gclk));
	jdff dff_A_d4ivGA2H9_0(.dout(w_dff_A_pjuNTLqz7_0),.din(w_dff_A_d4ivGA2H9_0),.clk(gclk));
	jdff dff_A_HzQF8z6P4_0(.dout(w_dff_A_d4ivGA2H9_0),.din(w_dff_A_HzQF8z6P4_0),.clk(gclk));
	jdff dff_A_CMzcZLjl3_1(.dout(w_G43gat_1[1]),.din(w_dff_A_CMzcZLjl3_1),.clk(gclk));
	jdff dff_A_aCVhvqVc9_1(.dout(w_G43gat_0[1]),.din(w_dff_A_aCVhvqVc9_1),.clk(gclk));
	jdff dff_A_SsxNEVmU4_2(.dout(w_G43gat_0[2]),.din(w_dff_A_SsxNEVmU4_2),.clk(gclk));
	jdff dff_A_pQNMbzjP3_0(.dout(w_G37gat_0[0]),.din(w_dff_A_pQNMbzjP3_0),.clk(gclk));
	jdff dff_A_NTImuhhq4_0(.dout(w_dff_A_pQNMbzjP3_0),.din(w_dff_A_NTImuhhq4_0),.clk(gclk));
	jdff dff_A_Sr3ZIu6M7_0(.dout(w_dff_A_NTImuhhq4_0),.din(w_dff_A_Sr3ZIu6M7_0),.clk(gclk));
	jdff dff_A_7q3qe1un9_0(.dout(w_dff_A_Sr3ZIu6M7_0),.din(w_dff_A_7q3qe1un9_0),.clk(gclk));
	jdff dff_A_cEPna7T99_0(.dout(w_dff_A_7q3qe1un9_0),.din(w_dff_A_cEPna7T99_0),.clk(gclk));
	jdff dff_A_HnbCd5xA0_0(.dout(w_dff_A_cEPna7T99_0),.din(w_dff_A_HnbCd5xA0_0),.clk(gclk));
	jdff dff_A_v7PrjEij8_1(.dout(w_G37gat_0[1]),.din(w_dff_A_v7PrjEij8_1),.clk(gclk));
	jdff dff_A_hpcNk6DJ6_0(.dout(w_G17gat_0[0]),.din(w_dff_A_hpcNk6DJ6_0),.clk(gclk));
	jdff dff_A_eJ6lv5Nq6_0(.dout(w_dff_A_hpcNk6DJ6_0),.din(w_dff_A_eJ6lv5Nq6_0),.clk(gclk));
	jdff dff_A_Td5rJ0GL6_0(.dout(w_dff_A_eJ6lv5Nq6_0),.din(w_dff_A_Td5rJ0GL6_0),.clk(gclk));
	jdff dff_A_4DB5y1E77_0(.dout(w_dff_A_Td5rJ0GL6_0),.din(w_dff_A_4DB5y1E77_0),.clk(gclk));
	jdff dff_A_AXRfQW691_0(.dout(w_dff_A_4DB5y1E77_0),.din(w_dff_A_AXRfQW691_0),.clk(gclk));
	jdff dff_A_gznuvzvn9_0(.dout(w_dff_A_AXRfQW691_0),.din(w_dff_A_gznuvzvn9_0),.clk(gclk));
	jdff dff_A_9XREv33Q7_0(.dout(w_dff_A_gznuvzvn9_0),.din(w_dff_A_9XREv33Q7_0),.clk(gclk));
	jdff dff_A_qtP09Y1i3_2(.dout(w_G17gat_0[2]),.din(w_dff_A_qtP09Y1i3_2),.clk(gclk));
	jdff dff_A_u4JIynEO0_0(.dout(w_n47_0[0]),.din(w_dff_A_u4JIynEO0_0),.clk(gclk));
	jdff dff_A_nK6Fl9I16_0(.dout(w_dff_A_u4JIynEO0_0),.din(w_dff_A_nK6Fl9I16_0),.clk(gclk));
	jdff dff_A_sGWpZJRV3_0(.dout(w_dff_A_nK6Fl9I16_0),.din(w_dff_A_sGWpZJRV3_0),.clk(gclk));
	jdff dff_A_Io2t5ywt9_0(.dout(w_dff_A_sGWpZJRV3_0),.din(w_dff_A_Io2t5ywt9_0),.clk(gclk));
	jdff dff_A_8u08u7938_0(.dout(w_dff_A_Io2t5ywt9_0),.din(w_dff_A_8u08u7938_0),.clk(gclk));
	jdff dff_A_pWsDNIww7_0(.dout(w_G11gat_0[0]),.din(w_dff_A_pWsDNIww7_0),.clk(gclk));
	jdff dff_A_kZ6Mg0QT4_0(.dout(w_dff_A_pWsDNIww7_0),.din(w_dff_A_kZ6Mg0QT4_0),.clk(gclk));
	jdff dff_A_JfXK5fDd6_0(.dout(w_dff_A_kZ6Mg0QT4_0),.din(w_dff_A_JfXK5fDd6_0),.clk(gclk));
	jdff dff_A_JZs7SXJM8_0(.dout(w_dff_A_JfXK5fDd6_0),.din(w_dff_A_JZs7SXJM8_0),.clk(gclk));
	jdff dff_A_DLfZkeoe3_0(.dout(w_dff_A_JZs7SXJM8_0),.din(w_dff_A_DLfZkeoe3_0),.clk(gclk));
	jdff dff_A_O2O27OSV9_0(.dout(w_dff_A_DLfZkeoe3_0),.din(w_dff_A_O2O27OSV9_0),.clk(gclk));
	jdff dff_A_6clacpgG8_1(.dout(w_G11gat_0[1]),.din(w_dff_A_6clacpgG8_1),.clk(gclk));
	jdff dff_A_UcNEqn591_1(.dout(w_G30gat_0[1]),.din(w_dff_A_UcNEqn591_1),.clk(gclk));
	jdff dff_A_7Aba9wMw0_0(.dout(w_G24gat_0[0]),.din(w_dff_A_7Aba9wMw0_0),.clk(gclk));
	jdff dff_A_ZYe2mqew6_1(.dout(w_n44_0[1]),.din(w_dff_A_ZYe2mqew6_1),.clk(gclk));
	jdff dff_A_jv5CgRg97_1(.dout(w_G82gat_0[1]),.din(w_dff_A_jv5CgRg97_1),.clk(gclk));
	jdff dff_A_YfDeoaEH9_1(.dout(w_dff_A_jv5CgRg97_1),.din(w_dff_A_YfDeoaEH9_1),.clk(gclk));
	jdff dff_A_dh8ZkW9p9_1(.dout(w_dff_A_YfDeoaEH9_1),.din(w_dff_A_dh8ZkW9p9_1),.clk(gclk));
	jdff dff_A_G5HHThQx3_1(.dout(w_dff_A_dh8ZkW9p9_1),.din(w_dff_A_G5HHThQx3_1),.clk(gclk));
	jdff dff_A_rgJckYea6_1(.dout(w_dff_A_G5HHThQx3_1),.din(w_dff_A_rgJckYea6_1),.clk(gclk));
	jdff dff_A_6rD5F3gE5_1(.dout(w_dff_A_rgJckYea6_1),.din(w_dff_A_6rD5F3gE5_1),.clk(gclk));
	jdff dff_A_x4t2TTDM3_1(.dout(w_dff_A_6rD5F3gE5_1),.din(w_dff_A_x4t2TTDM3_1),.clk(gclk));
	jdff dff_A_Tptql5QN1_2(.dout(w_G82gat_0[2]),.din(w_dff_A_Tptql5QN1_2),.clk(gclk));
	jdff dff_A_vAxnWIbk1_0(.dout(w_n43_0[0]),.din(w_dff_A_vAxnWIbk1_0),.clk(gclk));
	jdff dff_A_iVxv4iMo3_0(.dout(w_dff_A_vAxnWIbk1_0),.din(w_dff_A_iVxv4iMo3_0),.clk(gclk));
	jdff dff_A_VDHd53zs6_0(.dout(w_dff_A_iVxv4iMo3_0),.din(w_dff_A_VDHd53zs6_0),.clk(gclk));
	jdff dff_A_zNFhhy5i7_0(.dout(w_dff_A_VDHd53zs6_0),.din(w_dff_A_zNFhhy5i7_0),.clk(gclk));
	jdff dff_A_28XZIk1f5_0(.dout(w_dff_A_zNFhhy5i7_0),.din(w_dff_A_28XZIk1f5_0),.clk(gclk));
	jdff dff_A_oaDmFE1v4_0(.dout(w_G76gat_0[0]),.din(w_dff_A_oaDmFE1v4_0),.clk(gclk));
	jdff dff_A_mRpJm9BV8_0(.dout(w_dff_A_oaDmFE1v4_0),.din(w_dff_A_mRpJm9BV8_0),.clk(gclk));
	jdff dff_A_68YAXx8k7_0(.dout(w_dff_A_mRpJm9BV8_0),.din(w_dff_A_68YAXx8k7_0),.clk(gclk));
	jdff dff_A_jdw8FYVD9_0(.dout(w_dff_A_68YAXx8k7_0),.din(w_dff_A_jdw8FYVD9_0),.clk(gclk));
	jdff dff_A_HaarqPA04_0(.dout(w_dff_A_jdw8FYVD9_0),.din(w_dff_A_HaarqPA04_0),.clk(gclk));
	jdff dff_A_5BVq9ZHi3_0(.dout(w_dff_A_HaarqPA04_0),.din(w_dff_A_5BVq9ZHi3_0),.clk(gclk));
	jdff dff_A_82iLS9kc4_0(.dout(w_n87_0[0]),.din(w_dff_A_82iLS9kc4_0),.clk(gclk));
	jdff dff_A_Ewd8aq8n9_0(.dout(w_dff_A_82iLS9kc4_0),.din(w_dff_A_Ewd8aq8n9_0),.clk(gclk));
	jdff dff_A_Df6kt6vf1_0(.dout(w_dff_A_Ewd8aq8n9_0),.din(w_dff_A_Df6kt6vf1_0),.clk(gclk));
	jdff dff_A_09oEh0fq3_0(.dout(w_dff_A_Df6kt6vf1_0),.din(w_dff_A_09oEh0fq3_0),.clk(gclk));
	jdff dff_A_z76xChqN8_0(.dout(w_dff_A_09oEh0fq3_0),.din(w_dff_A_z76xChqN8_0),.clk(gclk));
	jdff dff_A_xxSMbtcd9_0(.dout(w_dff_A_z76xChqN8_0),.din(w_dff_A_xxSMbtcd9_0),.clk(gclk));
	jdff dff_A_5h1yS6Ot2_0(.dout(w_G95gat_0[0]),.din(w_dff_A_5h1yS6Ot2_0),.clk(gclk));
	jdff dff_A_gogxqGJE4_0(.dout(w_dff_A_5h1yS6Ot2_0),.din(w_dff_A_gogxqGJE4_0),.clk(gclk));
	jdff dff_A_zypnxrKF1_0(.dout(w_dff_A_gogxqGJE4_0),.din(w_dff_A_zypnxrKF1_0),.clk(gclk));
	jdff dff_A_odgcXlMO1_0(.dout(w_dff_A_zypnxrKF1_0),.din(w_dff_A_odgcXlMO1_0),.clk(gclk));
	jdff dff_A_r7nhHJni2_0(.dout(w_dff_A_odgcXlMO1_0),.din(w_dff_A_r7nhHJni2_0),.clk(gclk));
	jdff dff_A_C9ORlX8z2_0(.dout(w_dff_A_r7nhHJni2_0),.din(w_dff_A_C9ORlX8z2_0),.clk(gclk));
	jdff dff_A_zUeWR0hQ4_0(.dout(w_dff_A_C9ORlX8z2_0),.din(w_dff_A_zUeWR0hQ4_0),.clk(gclk));
	jdff dff_A_RLzJUKcF1_2(.dout(w_G95gat_0[2]),.din(w_dff_A_RLzJUKcF1_2),.clk(gclk));
	jdff dff_A_d8DihoTb7_1(.dout(w_G105gat_0[1]),.din(w_dff_A_d8DihoTb7_1),.clk(gclk));
	jdff dff_A_DRAlncLY7_1(.dout(w_dff_A_d8DihoTb7_1),.din(w_dff_A_DRAlncLY7_1),.clk(gclk));
	jdff dff_A_Owjh0MPB3_1(.dout(w_dff_A_DRAlncLY7_1),.din(w_dff_A_Owjh0MPB3_1),.clk(gclk));
	jdff dff_A_FvCoEDqA2_1(.dout(w_dff_A_Owjh0MPB3_1),.din(w_dff_A_FvCoEDqA2_1),.clk(gclk));
	jdff dff_A_8h3ouYZx8_1(.dout(w_dff_A_FvCoEDqA2_1),.din(w_dff_A_8h3ouYZx8_1),.clk(gclk));
	jdff dff_A_8hPUmbJ85_1(.dout(w_dff_A_8h3ouYZx8_1),.din(w_dff_A_8hPUmbJ85_1),.clk(gclk));
	jdff dff_A_4a4TCm1X8_1(.dout(w_dff_A_8hPUmbJ85_1),.din(w_dff_A_4a4TCm1X8_1),.clk(gclk));
	jdff dff_A_K8cZEKKZ3_1(.dout(w_dff_A_4a4TCm1X8_1),.din(w_dff_A_K8cZEKKZ3_1),.clk(gclk));
	jdff dff_A_dUtqgqT51_1(.dout(w_dff_A_K8cZEKKZ3_1),.din(w_dff_A_dUtqgqT51_1),.clk(gclk));
	jdff dff_A_H1wOdVD85_1(.dout(w_dff_A_dUtqgqT51_1),.din(w_dff_A_H1wOdVD85_1),.clk(gclk));
	jdff dff_A_HYZ0eSaV6_1(.dout(w_dff_A_H1wOdVD85_1),.din(w_dff_A_HYZ0eSaV6_1),.clk(gclk));
	jdff dff_A_eR5k1xLC3_1(.dout(w_dff_A_HYZ0eSaV6_1),.din(w_dff_A_eR5k1xLC3_1),.clk(gclk));
	jdff dff_A_7WCVBsNf6_1(.dout(w_dff_A_eR5k1xLC3_1),.din(w_dff_A_7WCVBsNf6_1),.clk(gclk));
	jdff dff_A_njq90PmN5_1(.dout(w_dff_A_7WCVBsNf6_1),.din(w_dff_A_njq90PmN5_1),.clk(gclk));
	jdff dff_A_QH0Pbqzg0_1(.dout(w_dff_A_njq90PmN5_1),.din(w_dff_A_QH0Pbqzg0_1),.clk(gclk));
	jdff dff_A_4UWrYcH12_2(.dout(w_dff_A_7XPuTqfg9_0),.din(w_dff_A_4UWrYcH12_2),.clk(gclk));
	jdff dff_A_7XPuTqfg9_0(.dout(w_dff_A_5vwQD4ir1_0),.din(w_dff_A_7XPuTqfg9_0),.clk(gclk));
	jdff dff_A_5vwQD4ir1_0(.dout(w_dff_A_06LKmq1Y4_0),.din(w_dff_A_5vwQD4ir1_0),.clk(gclk));
	jdff dff_A_06LKmq1Y4_0(.dout(w_dff_A_LeAI5wVU6_0),.din(w_dff_A_06LKmq1Y4_0),.clk(gclk));
	jdff dff_A_LeAI5wVU6_0(.dout(w_dff_A_Z6rZHQTN1_0),.din(w_dff_A_LeAI5wVU6_0),.clk(gclk));
	jdff dff_A_Z6rZHQTN1_0(.dout(w_dff_A_j2VuPVru3_0),.din(w_dff_A_Z6rZHQTN1_0),.clk(gclk));
	jdff dff_A_j2VuPVru3_0(.dout(w_dff_A_w1Y0VbNl4_0),.din(w_dff_A_j2VuPVru3_0),.clk(gclk));
	jdff dff_A_w1Y0VbNl4_0(.dout(w_dff_A_B4PSvxED7_0),.din(w_dff_A_w1Y0VbNl4_0),.clk(gclk));
	jdff dff_A_B4PSvxED7_0(.dout(w_dff_A_WqI6xG6K3_0),.din(w_dff_A_B4PSvxED7_0),.clk(gclk));
	jdff dff_A_WqI6xG6K3_0(.dout(w_dff_A_XGDkbvox3_0),.din(w_dff_A_WqI6xG6K3_0),.clk(gclk));
	jdff dff_A_XGDkbvox3_0(.dout(w_dff_A_6BtpPbvh9_0),.din(w_dff_A_XGDkbvox3_0),.clk(gclk));
	jdff dff_A_6BtpPbvh9_0(.dout(w_dff_A_7tzXGZCE4_0),.din(w_dff_A_6BtpPbvh9_0),.clk(gclk));
	jdff dff_A_7tzXGZCE4_0(.dout(w_dff_A_zGS1JHWz9_0),.din(w_dff_A_7tzXGZCE4_0),.clk(gclk));
	jdff dff_A_zGS1JHWz9_0(.dout(w_dff_A_vSSdYcUY8_0),.din(w_dff_A_zGS1JHWz9_0),.clk(gclk));
	jdff dff_A_vSSdYcUY8_0(.dout(w_dff_A_U0vy50sd4_0),.din(w_dff_A_vSSdYcUY8_0),.clk(gclk));
	jdff dff_A_U0vy50sd4_0(.dout(w_dff_A_v3i3QIfk4_0),.din(w_dff_A_U0vy50sd4_0),.clk(gclk));
	jdff dff_A_v3i3QIfk4_0(.dout(w_dff_A_jY6g6WIn8_0),.din(w_dff_A_v3i3QIfk4_0),.clk(gclk));
	jdff dff_A_jY6g6WIn8_0(.dout(w_dff_A_NN15yFkb0_0),.din(w_dff_A_jY6g6WIn8_0),.clk(gclk));
	jdff dff_A_NN15yFkb0_0(.dout(w_dff_A_n83oLjKe0_0),.din(w_dff_A_NN15yFkb0_0),.clk(gclk));
	jdff dff_A_n83oLjKe0_0(.dout(G223gat),.din(w_dff_A_n83oLjKe0_0),.clk(gclk));
	jdff dff_A_G75mAGmL5_1(.dout(w_dff_A_mN0xSzlM8_0),.din(w_dff_A_G75mAGmL5_1),.clk(gclk));
	jdff dff_A_mN0xSzlM8_0(.dout(w_dff_A_CoALeAd62_0),.din(w_dff_A_mN0xSzlM8_0),.clk(gclk));
	jdff dff_A_CoALeAd62_0(.dout(w_dff_A_GzS1AfhY6_0),.din(w_dff_A_CoALeAd62_0),.clk(gclk));
	jdff dff_A_GzS1AfhY6_0(.dout(w_dff_A_2ZIvObef1_0),.din(w_dff_A_GzS1AfhY6_0),.clk(gclk));
	jdff dff_A_2ZIvObef1_0(.dout(w_dff_A_SbcVLWP72_0),.din(w_dff_A_2ZIvObef1_0),.clk(gclk));
	jdff dff_A_SbcVLWP72_0(.dout(w_dff_A_dQKALZtM9_0),.din(w_dff_A_SbcVLWP72_0),.clk(gclk));
	jdff dff_A_dQKALZtM9_0(.dout(w_dff_A_ik9sEIgh2_0),.din(w_dff_A_dQKALZtM9_0),.clk(gclk));
	jdff dff_A_ik9sEIgh2_0(.dout(w_dff_A_5TF4eyZ79_0),.din(w_dff_A_ik9sEIgh2_0),.clk(gclk));
	jdff dff_A_5TF4eyZ79_0(.dout(w_dff_A_M6MKkLdS8_0),.din(w_dff_A_5TF4eyZ79_0),.clk(gclk));
	jdff dff_A_M6MKkLdS8_0(.dout(w_dff_A_lwVELHM53_0),.din(w_dff_A_M6MKkLdS8_0),.clk(gclk));
	jdff dff_A_lwVELHM53_0(.dout(w_dff_A_NWMctVa41_0),.din(w_dff_A_lwVELHM53_0),.clk(gclk));
	jdff dff_A_NWMctVa41_0(.dout(w_dff_A_7T7WMs6T4_0),.din(w_dff_A_NWMctVa41_0),.clk(gclk));
	jdff dff_A_7T7WMs6T4_0(.dout(G329gat),.din(w_dff_A_7T7WMs6T4_0),.clk(gclk));
	jdff dff_A_JCVWIwh73_1(.dout(w_dff_A_7QbPNyfA3_0),.din(w_dff_A_JCVWIwh73_1),.clk(gclk));
	jdff dff_A_7QbPNyfA3_0(.dout(w_dff_A_MK8mbjgS5_0),.din(w_dff_A_7QbPNyfA3_0),.clk(gclk));
	jdff dff_A_MK8mbjgS5_0(.dout(w_dff_A_6Ut5Kybk8_0),.din(w_dff_A_MK8mbjgS5_0),.clk(gclk));
	jdff dff_A_6Ut5Kybk8_0(.dout(w_dff_A_HUwmCVVV9_0),.din(w_dff_A_6Ut5Kybk8_0),.clk(gclk));
	jdff dff_A_HUwmCVVV9_0(.dout(w_dff_A_02IdJ8190_0),.din(w_dff_A_HUwmCVVV9_0),.clk(gclk));
	jdff dff_A_02IdJ8190_0(.dout(G370gat),.din(w_dff_A_02IdJ8190_0),.clk(gclk));
	jdff dff_A_xghxYD4R6_1(.dout(w_dff_A_TvqwLfSQ7_0),.din(w_dff_A_xghxYD4R6_1),.clk(gclk));
	jdff dff_A_TvqwLfSQ7_0(.dout(G430gat),.din(w_dff_A_TvqwLfSQ7_0),.clk(gclk));
endmodule

