/*

c499:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jdff: 435
	jor: 10
	jand: 61

Summary:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jdff: 435
	jor: 10
	jand: 61
*/

module c499(gclk, Gid0, Gid1, Gid2, Gid3, Gid4, Gid5, Gid6, Gid7, Gid8, Gid9, Gid10, Gid11, Gid12, Gid13, Gid14, Gid15, Gid16, Gid17, Gid18, Gid19, Gid20, Gid21, Gid22, Gid23, Gid24, Gid25, Gid26, Gid27, Gid28, Gid29, Gid30, Gid31, Gic0, Gic1, Gic2, Gic3, Gic4, Gic5, Gic6, Gic7, Gr, God0, God1, God2, God3, God4, God5, God6, God7, God8, God9, God10, God11, God12, God13, God14, God15, God16, God17, God18, God19, God20, God21, God22, God23, God24, God25, God26, God27, God28, God29, God30, God31);
	input gclk;
	input Gid0;
	input Gid1;
	input Gid2;
	input Gid3;
	input Gid4;
	input Gid5;
	input Gid6;
	input Gid7;
	input Gid8;
	input Gid9;
	input Gid10;
	input Gid11;
	input Gid12;
	input Gid13;
	input Gid14;
	input Gid15;
	input Gid16;
	input Gid17;
	input Gid18;
	input Gid19;
	input Gid20;
	input Gid21;
	input Gid22;
	input Gid23;
	input Gid24;
	input Gid25;
	input Gid26;
	input Gid27;
	input Gid28;
	input Gid29;
	input Gid30;
	input Gid31;
	input Gic0;
	input Gic1;
	input Gic2;
	input Gic3;
	input Gic4;
	input Gic5;
	input Gic6;
	input Gic7;
	input Gr;
	output God0;
	output God1;
	output God2;
	output God3;
	output God4;
	output God5;
	output God6;
	output God7;
	output God8;
	output God9;
	output God10;
	output God11;
	output God12;
	output God13;
	output God14;
	output God15;
	output God16;
	output God17;
	output God18;
	output God19;
	output God20;
	output God21;
	output God22;
	output God23;
	output God24;
	output God25;
	output God26;
	output God27;
	output God28;
	output God29;
	output God30;
	output God31;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n178;
	wire n179;
	wire n181;
	wire n182;
	wire n184;
	wire n185;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n192;
	wire n194;
	wire n196;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n204;
	wire n206;
	wire n208;
	wire n210;
	wire n211;
	wire n212;
	wire n214;
	wire n216;
	wire n218;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n233;
	wire n235;
	wire n237;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n244;
	wire n246;
	wire n248;
	wire n250;
	wire n251;
	wire n252;
	wire n254;
	wire n256;
	wire n258;
	wire n260;
	wire n261;
	wire n263;
	wire n265;
	wire n267;
	wire[2:0] w_Gid0_0;
	wire[2:0] w_Gid1_0;
	wire[2:0] w_Gid2_0;
	wire[2:0] w_Gid3_0;
	wire[2:0] w_Gid4_0;
	wire[2:0] w_Gid5_0;
	wire[2:0] w_Gid6_0;
	wire[2:0] w_Gid7_0;
	wire[2:0] w_Gid8_0;
	wire[2:0] w_Gid9_0;
	wire[2:0] w_Gid10_0;
	wire[2:0] w_Gid11_0;
	wire[2:0] w_Gid12_0;
	wire[2:0] w_Gid13_0;
	wire[2:0] w_Gid14_0;
	wire[2:0] w_Gid15_0;
	wire[2:0] w_Gid16_0;
	wire[2:0] w_Gid17_0;
	wire[2:0] w_Gid18_0;
	wire[2:0] w_Gid19_0;
	wire[2:0] w_Gid20_0;
	wire[2:0] w_Gid21_0;
	wire[2:0] w_Gid22_0;
	wire[2:0] w_Gid23_0;
	wire[2:0] w_Gid24_0;
	wire[2:0] w_Gid25_0;
	wire[2:0] w_Gid26_0;
	wire[2:0] w_Gid27_0;
	wire[2:0] w_Gid28_0;
	wire[2:0] w_Gid29_0;
	wire[2:0] w_Gid30_0;
	wire[2:0] w_Gid31_0;
	wire[2:0] w_n74_0;
	wire[2:0] w_n74_1;
	wire[2:0] w_n74_2;
	wire[1:0] w_n74_3;
	wire[1:0] w_n78_0;
	wire[1:0] w_n85_0;
	wire[2:0] w_n87_0;
	wire[1:0] w_n87_1;
	wire[2:0] w_n88_0;
	wire[2:0] w_n88_1;
	wire[1:0] w_n93_0;
	wire[1:0] w_n97_0;
	wire[2:0] w_n102_0;
	wire[1:0] w_n102_1;
	wire[1:0] w_n107_0;
	wire[1:0] w_n111_0;
	wire[2:0] w_n116_0;
	wire[1:0] w_n116_1;
	wire[2:0] w_n117_0;
	wire[2:0] w_n117_1;
	wire[1:0] w_n118_0;
	wire[2:0] w_n126_0;
	wire[1:0] w_n126_1;
	wire[2:0] w_n127_0;
	wire[2:0] w_n127_1;
	wire[2:0] w_n135_0;
	wire[1:0] w_n135_1;
	wire[1:0] w_n141_0;
	wire[1:0] w_n145_0;
	wire[2:0] w_n150_0;
	wire[1:0] w_n150_1;
	wire[2:0] w_n159_0;
	wire[1:0] w_n159_1;
	wire[2:0] w_n167_0;
	wire[1:0] w_n167_1;
	wire[2:0] w_n173_0;
	wire[1:0] w_n174_0;
	wire[2:0] w_n175_0;
	wire[1:0] w_n175_1;
	wire[2:0] w_n178_0;
	wire[2:0] w_n178_1;
	wire[2:0] w_n181_0;
	wire[2:0] w_n181_1;
	wire[2:0] w_n184_0;
	wire[2:0] w_n184_1;
	wire[2:0] w_n187_0;
	wire[2:0] w_n187_1;
	wire[1:0] w_n188_0;
	wire[2:0] w_n189_0;
	wire[1:0] w_n189_1;
	wire[2:0] w_n198_0;
	wire[2:0] w_n198_1;
	wire[1:0] w_n199_0;
	wire[2:0] w_n201_0;
	wire[1:0] w_n201_1;
	wire[2:0] w_n211_0;
	wire[1:0] w_n211_1;
	wire[1:0] w_n220_0;
	wire[1:0] w_n228_0;
	wire[1:0] w_n229_0;
	wire[2:0] w_n230_0;
	wire[1:0] w_n230_1;
	wire[1:0] w_n240_0;
	wire[2:0] w_n241_0;
	wire[1:0] w_n241_1;
	wire[1:0] w_n250_0;
	wire[2:0] w_n251_0;
	wire[1:0] w_n251_1;
	wire[2:0] w_n260_0;
	wire[1:0] w_n260_1;
	wire w_dff_B_7YbQlWtC6_1;
	wire w_dff_A_QrMOdnYP1_1;
	wire w_dff_A_1s1teyGQ6_2;
	wire w_dff_A_5NSGo9VV3_1;
	wire w_dff_A_CL6Ni2838_2;
	wire w_dff_A_VS7e9OZH6_1;
	wire w_dff_A_n7BkOgZh9_2;
	wire w_dff_A_mFpqzfM30_1;
	wire w_dff_A_BZxubKaJ9_1;
	wire w_dff_A_uPgEDf7R4_1;
	wire w_dff_A_fzY6eBTi1_2;
	wire w_dff_A_SXflDD7T8_1;
	wire w_dff_A_48Somc154_1;
	wire w_dff_A_lwhZyFww2_0;
	wire w_dff_A_lhsPZKHs4_0;
	wire w_dff_A_iALwGt6S2_0;
	wire w_dff_A_GtwcM2vK5_0;
	wire w_dff_A_PHiG1CSh7_1;
	wire w_dff_A_SMJgTvvT1_1;
	wire w_dff_A_ZeB9MUyM2_1;
	wire w_dff_A_o3YawC4w9_1;
	wire w_dff_A_VJy4WXiw8_0;
	wire w_dff_A_dGU7Q6J78_0;
	wire w_dff_A_4R7B6Wh38_0;
	wire w_dff_A_gKqMLxcP6_0;
	wire w_dff_A_JFpFKBNG1_1;
	wire w_dff_A_VeDNxiOF6_1;
	wire w_dff_A_UKrSRaEl5_1;
	wire w_dff_A_845KEc5h4_1;
	wire w_dff_A_8WS4zO9O3_0;
	wire w_dff_A_OaONNhR07_0;
	wire w_dff_A_Qvsf2YyU6_0;
	wire w_dff_A_tY6nUX7m2_0;
	wire w_dff_A_4VRf9T5Y7_1;
	wire w_dff_A_MNpC9Wjq8_1;
	wire w_dff_A_snKzvNyW6_1;
	wire w_dff_A_P80ByBBx9_1;
	wire w_dff_B_1nPWFy1U6_2;
	wire w_dff_B_9hY9tMd39_2;
	wire w_dff_A_B92hbzQf5_0;
	wire w_dff_A_VpUnDeto3_0;
	wire w_dff_A_uWCDLAHs3_0;
	wire w_dff_A_t38aZdH66_2;
	wire w_dff_A_c0SnWTV59_2;
	wire w_dff_A_894mahDr7_2;
	wire w_dff_A_Czs4lalI4_0;
	wire w_dff_A_osHw9K8I5_0;
	wire w_dff_A_dM6bzT9h7_0;
	wire w_dff_A_apFlQxxA3_0;
	wire w_dff_A_yjiHvioF7_1;
	wire w_dff_A_9HYyYcwz2_1;
	wire w_dff_A_WXJKU94Y1_1;
	wire w_dff_A_GZUUKd7t2_1;
	wire w_dff_B_6rCY2ARc4_1;
	wire w_dff_A_rmJkwMMt6_0;
	wire w_dff_A_Hxld7UWi4_0;
	wire w_dff_A_HqSlzSuR4_0;
	wire w_dff_A_A0GkoZMn1_2;
	wire w_dff_A_sJHs71t46_2;
	wire w_dff_A_TgHx8kkL7_2;
	wire w_dff_A_Oc2hW7pF6_1;
	wire w_dff_A_ckuUy3Ub8_1;
	wire w_dff_A_AXsjO57F2_1;
	wire w_dff_A_XRGzg8M38_1;
	wire w_dff_A_oaafBjdD2_2;
	wire w_dff_A_GFvLG8uw0_2;
	wire w_dff_A_Jvgnk5390_2;
	wire w_dff_A_Ytk3OuDc2_2;
	wire w_dff_A_GbwvgkeW8_0;
	wire w_dff_A_8WshvURS4_1;
	wire w_dff_A_rImFUdkE8_1;
	wire w_dff_A_STZojGsg1_1;
	wire w_dff_A_Ts1tV0HU8_1;
	wire w_dff_A_M8L1bXfV4_2;
	wire w_dff_A_NFBmxYkG8_2;
	wire w_dff_A_bgVWcr2A2_2;
	wire w_dff_A_QWvYTr0x0_2;
	wire w_dff_A_Rj5xck4f5_1;
	wire w_dff_A_4r0VLs4A1_1;
	wire w_dff_A_pFFjlh4U0_1;
	wire w_dff_A_vkZXroMs3_1;
	wire w_dff_A_7RdF8kzx1_1;
	wire w_dff_A_PwzWTOPB7_2;
	wire w_dff_A_qIJd2k9C2_2;
	wire w_dff_A_SKQwpJTr8_2;
	wire w_dff_A_NJnKpFfd4_2;
	wire w_dff_A_3gCewhSK3_0;
	wire w_dff_B_FleaHSHC9_1;
	wire w_dff_A_LLiTtz3t7_1;
	wire w_dff_A_38nVQwmt1_0;
	wire w_dff_A_rK9ij8KF1_0;
	wire w_dff_A_30hBPQ7Z2_0;
	wire w_dff_A_Ubv2Das33_0;
	wire w_dff_A_ml4J5NVi7_0;
	wire w_dff_A_yi2q2qFV0_0;
	wire w_dff_A_lUTjZBY86_0;
	wire w_dff_A_6Uhkmc3p8_0;
	wire w_dff_A_pxZO4WQg6_0;
	wire w_dff_A_dFRGcD4F3_0;
	wire w_dff_A_VVtbHkcH3_0;
	wire w_dff_A_nHGgnyYA9_0;
	wire w_dff_A_sVXwo5di9_0;
	wire w_dff_A_eQ4y9QWG4_0;
	wire w_dff_A_XHe0UZA90_0;
	wire w_dff_A_45Vf5dGX7_0;
	wire w_dff_A_QDDCTmk69_0;
	wire w_dff_A_Knrcr0Ea7_0;
	wire w_dff_A_lFxY92ZG4_0;
	wire w_dff_A_6urkEdQt8_0;
	wire w_dff_A_oL1oe9uq8_0;
	wire w_dff_A_6NQTQiCa1_0;
	wire w_dff_A_1ikuqBfP1_2;
	wire w_dff_A_s707V4sK4_2;
	wire w_dff_A_OEJiDYKX7_2;
	wire w_dff_A_MfDVjbvw0_1;
	wire w_dff_A_damvTCjB5_0;
	wire w_dff_A_n3JJdcyq3_0;
	wire w_dff_A_ji9KaFGI4_0;
	wire w_dff_A_9oMO89141_0;
	wire w_dff_A_tHDn59u91_0;
	wire w_dff_A_j0vSDVcx8_0;
	wire w_dff_A_LeaqXqFE5_0;
	wire w_dff_A_6POJdunu5_0;
	wire w_dff_A_ygrfhaGE6_0;
	wire w_dff_A_PfbGDkXL9_0;
	wire w_dff_A_WeIGzFmv9_0;
	wire w_dff_A_K5PWTxRS6_0;
	wire w_dff_A_C5ixUU0g4_0;
	wire w_dff_A_9uY4yoLn4_0;
	wire w_dff_A_emgS1Ykw7_0;
	wire w_dff_A_UfFQBhxF8_0;
	wire w_dff_A_cPuUE9rM0_0;
	wire w_dff_A_8ASR3HiH1_0;
	wire w_dff_A_Ehs49Qsy1_0;
	wire w_dff_B_8nYFBoOb8_2;
	wire w_dff_B_97l74v724_2;
	wire w_dff_A_RYxZPFGf4_0;
	wire w_dff_A_dfjMCcgO4_0;
	wire w_dff_A_mUG1xxPk9_0;
	wire w_dff_A_feF2dWmY3_2;
	wire w_dff_A_qe2FC22Z9_2;
	wire w_dff_A_2hdwB6Lq7_2;
	wire w_dff_A_ZIJzp40A1_1;
	wire w_dff_A_jcRibDaM3_0;
	wire w_dff_A_sXwhbR2z7_0;
	wire w_dff_A_tEyLqnCC7_0;
	wire w_dff_A_k8pmRiuA4_0;
	wire w_dff_A_xzgTCJ4g3_0;
	wire w_dff_A_AVxenFrp8_0;
	wire w_dff_A_iZ18YbbF2_0;
	wire w_dff_A_IHqJUW780_0;
	wire w_dff_A_QN1AQoE70_0;
	wire w_dff_A_nlfCY9eZ4_0;
	wire w_dff_A_VfVBi8kn2_0;
	wire w_dff_A_yjFwUfV27_0;
	wire w_dff_A_h4aYqerg9_0;
	wire w_dff_A_zMcu6Y4R6_0;
	wire w_dff_A_3SAy5bVJ5_0;
	wire w_dff_A_yQumS6Iw9_0;
	wire w_dff_A_jh3krFEq8_0;
	wire w_dff_A_t0lijdpE6_0;
	wire w_dff_A_juUxwNZX6_0;
	wire w_dff_A_FzQHVQVd1_0;
	wire w_dff_A_BLHOFcvB6_0;
	wire w_dff_A_vpCMzqWU5_0;
	wire w_dff_A_Y7uubj8a8_0;
	wire w_dff_A_If2AlXxL1_0;
	wire w_dff_A_gnFqC4Ql6_0;
	wire w_dff_A_Cji16JFo9_0;
	wire w_dff_A_WKU0TH3V0_0;
	wire w_dff_A_Uxnxvwc57_0;
	wire w_dff_A_hNLQDEle0_0;
	wire w_dff_A_xSBXQeTL8_0;
	wire w_dff_A_ULrjhnzx1_0;
	wire w_dff_A_gZD9nxQC3_0;
	wire w_dff_A_HVbIHqyp8_0;
	wire w_dff_A_oCsZXx1N0_0;
	wire w_dff_A_NU4DqDz64_0;
	wire w_dff_A_RcUmVaze5_0;
	wire w_dff_A_gy9DVSgM8_0;
	wire w_dff_A_Tl3Ue38z6_0;
	wire w_dff_A_lwZhi6iY6_0;
	wire w_dff_A_Br7A30gp1_0;
	wire w_dff_A_EZBUjOOC7_0;
	wire w_dff_A_o7StwBmy3_0;
	wire w_dff_A_3UWQ7sKS4_0;
	wire w_dff_A_TLbHxl1l5_0;
	wire w_dff_A_BByKlYj37_0;
	wire w_dff_A_4DsW3pay3_0;
	wire w_dff_A_VOtCwJvH5_0;
	wire w_dff_A_gBstYV6h6_0;
	wire w_dff_A_E22RhgI36_0;
	wire w_dff_A_iSDbBGr43_0;
	wire w_dff_A_aL55yYLe9_0;
	wire w_dff_A_1Wz5YjX11_0;
	wire w_dff_A_C3gVbDDy7_0;
	wire w_dff_A_bB8KWaiS7_0;
	wire w_dff_A_fqKjbUVE3_0;
	wire w_dff_A_7txFciWh6_0;
	wire w_dff_A_HzozIe276_0;
	wire w_dff_A_t2tzlX5U5_0;
	wire w_dff_A_3GoHoAV63_0;
	wire w_dff_A_iII172id8_0;
	wire w_dff_A_qiLWyHXx3_0;
	wire w_dff_A_FFNvq2nn4_0;
	wire w_dff_A_HhFUejdw5_0;
	wire w_dff_A_Nl3czyl52_0;
	wire w_dff_A_bxdbeUFt4_0;
	wire w_dff_A_3EnfGnyW3_0;
	wire w_dff_A_uroHc92O6_0;
	wire w_dff_A_pxjUCRIP6_0;
	wire w_dff_A_ZXZxQSbT4_0;
	wire w_dff_A_q7ENROth4_0;
	wire w_dff_A_oqCosAcc4_0;
	wire w_dff_A_fS4jQyCt4_0;
	wire w_dff_A_FyGHhDte8_0;
	wire w_dff_A_FVWW2Ufc7_0;
	wire w_dff_A_WB9YVhx87_0;
	wire w_dff_A_IFQ5cYYB5_0;
	wire w_dff_A_1WRkxZYv3_0;
	wire w_dff_A_EhMyHGaN7_0;
	wire w_dff_A_JaGskUwi2_0;
	wire w_dff_A_JHfHeD4W6_1;
	wire w_dff_A_e0f20Of68_0;
	wire w_dff_A_csABP28l4_0;
	wire w_dff_A_zzxR9Ii12_0;
	wire w_dff_A_aEngsCQg0_0;
	wire w_dff_A_3dAHsyre7_0;
	wire w_dff_A_1kR1fyGQ3_0;
	wire w_dff_A_2ZM9I5Sk7_0;
	wire w_dff_A_I2MMOWyw3_0;
	wire w_dff_A_TSyhpsdb2_0;
	wire w_dff_A_v52rLRPg7_0;
	wire w_dff_A_d9cdBOFM4_0;
	wire w_dff_A_HLcoKE646_0;
	wire w_dff_A_4fL9euP86_0;
	wire w_dff_A_izpaHMpn7_0;
	wire w_dff_A_wqL0WCtR1_0;
	wire w_dff_A_uFK8DEfL4_0;
	wire w_dff_A_ANU9vpyT4_0;
	wire w_dff_A_wutTKT5o0_0;
	wire w_dff_A_yREcq8vF1_0;
	wire w_dff_A_y3d5rboI7_0;
	wire w_dff_A_SyMPwkUR6_0;
	wire w_dff_A_0uB8qeBw8_0;
	wire w_dff_A_R0ccmP144_0;
	wire w_dff_A_eXfOj34b5_0;
	wire w_dff_A_iIYXS9XK7_0;
	wire w_dff_A_tjPp8cGe8_0;
	wire w_dff_A_6Snlr1V52_0;
	wire w_dff_A_D2Vol7Oi9_0;
	wire w_dff_A_PcBKuAi53_0;
	wire w_dff_A_I7zSl4Oo8_0;
	wire w_dff_A_1Mta0FRo5_0;
	wire w_dff_A_oBehxNMy4_0;
	wire w_dff_A_0hClBwca0_0;
	wire w_dff_A_4eS53urV3_0;
	wire w_dff_A_MqWWxRTY9_0;
	wire w_dff_A_Et9KTzRE0_0;
	wire w_dff_A_nHlYQRJx5_0;
	wire w_dff_A_Eec6HTvf2_0;
	wire w_dff_A_QXExpRAt1_0;
	wire w_dff_A_xFw1BOWp5_0;
	wire w_dff_A_xciZE5IX8_0;
	wire w_dff_A_aQfHNGca7_0;
	wire w_dff_A_Ye6CAmvR5_0;
	wire w_dff_A_SMiNFZbi2_0;
	wire w_dff_A_bWdPzZaC7_0;
	wire w_dff_A_PLoh3owQ5_0;
	wire w_dff_A_1FPAdSGH2_0;
	wire w_dff_A_zXvLuIgT6_0;
	wire w_dff_A_YsUNoZov4_0;
	wire w_dff_A_Ff6PPWup0_0;
	wire w_dff_A_513AJPwb8_0;
	wire w_dff_A_4sptdXIf1_0;
	wire w_dff_A_DuJIQdFk5_0;
	wire w_dff_A_Obufz23g4_0;
	wire w_dff_A_pgk63Lcf8_0;
	wire w_dff_A_NGkQye6u3_0;
	wire w_dff_A_iKJVKK5Q9_0;
	wire w_dff_A_Y9aZM7VE5_0;
	wire w_dff_A_PaXUWnuJ3_0;
	wire w_dff_A_AfRlojZO8_0;
	wire w_dff_A_tMbb5eAY2_0;
	wire w_dff_A_PkBcyinB3_0;
	wire w_dff_A_ulc6f5Hj8_0;
	wire w_dff_A_7W1mUFqy7_0;
	wire w_dff_A_WT7ho4U09_0;
	wire w_dff_A_1WgJfbkc2_0;
	wire w_dff_A_LeV0kfew9_0;
	wire w_dff_A_Z1lRabTN9_0;
	wire w_dff_A_OVz3kojF3_0;
	wire w_dff_A_Z8nhfsjM3_0;
	wire w_dff_A_J9i1HOod0_0;
	wire w_dff_A_YsORmye48_0;
	wire w_dff_A_041Jrkqp4_0;
	wire w_dff_A_YtNhgngi9_0;
	wire w_dff_A_nr9wxVt56_0;
	wire w_dff_A_Zcncu5pV7_0;
	wire w_dff_A_2Z72Bbfy8_0;
	wire w_dff_A_ACqLObVw9_0;
	wire w_dff_A_XmRrv8nG7_0;
	wire w_dff_A_b7eWEwPm2_1;
	wire w_dff_A_1pXnnjqi2_1;
	wire w_dff_A_F9sOOZqT0_1;
	wire w_dff_A_uBkBXEWl3_1;
	wire w_dff_A_N2Wba22G6_2;
	wire w_dff_A_vOnKQtMl7_2;
	wire w_dff_A_OhFFmIKc1_2;
	wire w_dff_A_H1KiPvTH0_2;
	wire w_dff_A_HEyAYzEs7_1;
	wire w_dff_A_QwzLAtAx0_0;
	wire w_dff_A_kL8Q0MNb7_0;
	wire w_dff_A_pFlmQUJv2_0;
	wire w_dff_A_66XdLzSi4_0;
	wire w_dff_A_1DBHxGAI1_0;
	wire w_dff_A_2SweqIOi6_0;
	wire w_dff_A_bFXseTRd8_0;
	wire w_dff_A_rQr6v7Hq8_0;
	wire w_dff_A_xNU8rjDp3_0;
	wire w_dff_A_wLmNjqFi8_0;
	wire w_dff_A_V9575tAZ8_0;
	wire w_dff_A_yZI0PRA86_0;
	wire w_dff_A_yaYnJmvC0_0;
	wire w_dff_A_jPDojBgh2_0;
	wire w_dff_A_9zRgDp2a0_0;
	wire w_dff_A_Q8EqOzhI7_0;
	wire w_dff_A_HYtNnSkz9_0;
	wire w_dff_A_hxa6lDUx0_0;
	wire w_dff_A_x8XdVgs38_0;
	wire w_dff_A_MO03c5xV3_0;
	wire w_dff_A_iELAqCDW6_0;
	wire w_dff_A_b2gsjM1n4_0;
	wire w_dff_A_G1z5U4Ui5_0;
	wire w_dff_A_0wYk2Vb47_0;
	wire w_dff_A_EuBlqX472_0;
	wire w_dff_A_QAcPOklx8_0;
	wire w_dff_A_rwaFJ7H30_0;
	wire w_dff_A_tujslkKe0_0;
	wire w_dff_A_GBOUtBRn5_0;
	wire w_dff_A_bQX9gF2S9_0;
	wire w_dff_A_Xqmn3PZp8_0;
	wire w_dff_A_PanEnjlZ5_0;
	wire w_dff_A_R80Rcvg22_0;
	wire w_dff_A_01dvP1cg0_0;
	wire w_dff_A_FAfElg7H6_0;
	wire w_dff_A_NU3ew8Bb0_0;
	wire w_dff_A_mWhAP6Fw3_0;
	wire w_dff_A_3c0OhL8m9_0;
	wire w_dff_A_WCBBAKzQ6_0;
	wire w_dff_A_LEJdWwnh0_0;
	wire w_dff_A_RR0yQgGz8_0;
	wire w_dff_A_GNO3S7JI7_0;
	wire w_dff_A_Qp3b8qrn2_0;
	wire w_dff_A_W7m6Syd27_0;
	wire w_dff_A_LVNs9DC23_0;
	wire w_dff_A_QLbsGLBj8_0;
	wire w_dff_A_0GMcFs7C9_0;
	wire w_dff_A_7S7rZln52_0;
	wire w_dff_A_n9T6JgZ27_0;
	wire w_dff_A_9FSP0flA0_0;
	wire w_dff_A_9dUWoDcq5_0;
	wire w_dff_A_E6m84ZSg5_0;
	wire w_dff_A_UfpAOE2k9_0;
	wire w_dff_A_3XWJwo7R6_0;
	wire w_dff_A_hG1tkdaa0_0;
	wire w_dff_A_VeBN4WF29_0;
	wire w_dff_A_2EylyEZ32_0;
	wire w_dff_A_aOH4rWq78_0;
	wire w_dff_A_ww2WoK2p2_0;
	wire w_dff_A_OVoP1XFp3_0;
	wire w_dff_A_gq5vEoM78_0;
	wire w_dff_A_KJ5ptrdO7_0;
	wire w_dff_A_FoYtcmCu0_0;
	wire w_dff_A_aBT8h6OV8_0;
	wire w_dff_A_rKYBJCle1_0;
	wire w_dff_A_kexKDfbr0_0;
	wire w_dff_A_Kr1W6KUY5_0;
	wire w_dff_A_nt8rdOU21_0;
	wire w_dff_A_uqCtPmK78_0;
	wire w_dff_A_mN7DoGtO0_0;
	wire w_dff_A_YCGO4eY17_0;
	wire w_dff_A_5bK44Lyn8_0;
	wire w_dff_A_S2AYlz2y0_0;
	wire w_dff_A_156YnIVW1_0;
	wire w_dff_A_kWhGq2h96_0;
	wire w_dff_A_qYT5kUyt1_0;
	wire w_dff_A_y9UQfaWF4_0;
	wire w_dff_A_TF025xm65_0;
	wire w_dff_A_6uKN7KI02_0;
	wire w_dff_A_D2tEnZjR8_0;
	wire w_dff_A_Gjh6vQlf6_0;
	wire w_dff_A_WiWxKCtv5_0;
	wire w_dff_A_KJ3azRhd9_0;
	wire w_dff_A_7bJDUGNK3_0;
	wire w_dff_A_O4hbQfBu2_0;
	wire w_dff_A_kkrNQRKE5_0;
	wire w_dff_A_ChfgxBH58_0;
	wire w_dff_A_ygmvpjdG3_0;
	wire w_dff_A_b7N7qzQE2_0;
	wire w_dff_A_gpRYnFCl7_0;
	wire w_dff_A_VScFfyKD7_0;
	wire w_dff_A_TALpwPhe1_0;
	wire w_dff_A_bD3AqHE21_0;
	wire w_dff_A_nusqCQWs6_0;
	wire w_dff_A_PFRawVxt0_0;
	wire w_dff_A_sNMh06Yt4_0;
	wire w_dff_A_QK1h1veC1_0;
	wire w_dff_A_UTKoS5Yv5_0;
	wire w_dff_A_0ibMUIzf3_0;
	wire w_dff_A_wPOUYrxu9_0;
	wire w_dff_A_xpiFaIlY9_0;
	wire w_dff_A_ms0oWAOE9_0;
	wire w_dff_A_qhXLmvOf5_0;
	wire w_dff_A_fOFV1D9z7_0;
	wire w_dff_A_nQbZTHNI7_0;
	wire w_dff_A_BfT7Vhzc5_0;
	wire w_dff_A_yR6PgPst6_0;
	wire w_dff_A_Vw3TsTGp2_0;
	wire w_dff_A_SKUvScIw6_0;
	wire w_dff_A_V2rYNcDl9_0;
	wire w_dff_A_AJR36qPJ9_0;
	wire w_dff_A_uziHMTnu4_0;
	wire w_dff_A_CrOmOJbG8_0;
	wire w_dff_A_kr8LbF5O2_0;
	wire w_dff_A_OEBpZGBL0_0;
	wire w_dff_A_ZgwJAPqV3_0;
	wire w_dff_A_xZiBlxD60_2;
	wire w_dff_A_GC3Ur5fC0_2;
	wire w_dff_A_qT9JmB3C5_2;
	wire w_dff_A_2iNFlhGO6_2;
	wire w_dff_A_k1Z9d4Mf4_2;
	wire w_dff_A_2woWXhQe4_2;
	wire w_dff_A_02xLMDyO5_2;
	wire w_dff_A_XsRivswP4_2;
	jnot g000(.din(Gic0),.dout(n73),.clk(gclk));
	jnot g001(.din(Gr),.dout(n74),.clk(gclk));
	jor g002(.dina(w_n74_3[1]),.dinb(n73),.dout(n75),.clk(gclk));
	jxor g003(.dina(w_Gid17_0[2]),.dinb(w_Gid16_0[2]),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_Gid19_0[2]),.dinb(w_Gid18_0[2]),.dout(n77),.clk(gclk));
	jxor g005(.dina(n77),.dinb(n76),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_n78_0[1]),.dinb(n75),.dout(n79),.clk(gclk));
	jxor g007(.dina(w_Gid4_0[2]),.dinb(w_Gid0_0[2]),.dout(n80),.clk(gclk));
	jxor g008(.dina(w_Gid12_0[2]),.dinb(w_Gid8_0[2]),.dout(n81),.clk(gclk));
	jxor g009(.dina(n81),.dinb(n80),.dout(n82),.clk(gclk));
	jxor g010(.dina(w_Gid21_0[2]),.dinb(w_Gid20_0[2]),.dout(n83),.clk(gclk));
	jxor g011(.dina(w_Gid23_0[2]),.dinb(w_Gid22_0[2]),.dout(n84),.clk(gclk));
	jxor g012(.dina(n84),.dinb(n83),.dout(n85),.clk(gclk));
	jxor g013(.dina(w_n85_0[1]),.dinb(n82),.dout(n86),.clk(gclk));
	jxor g014(.dina(n86),.dinb(n79),.dout(n87),.clk(gclk));
	jnot g015(.din(w_n87_1[1]),.dout(n88),.clk(gclk));
	jnot g016(.din(Gic7),.dout(n89),.clk(gclk));
	jor g017(.dina(w_n74_3[0]),.dinb(n89),.dout(n90),.clk(gclk));
	jxor g018(.dina(w_Gid5_0[2]),.dinb(w_Gid4_0[1]),.dout(n91),.clk(gclk));
	jxor g019(.dina(w_Gid7_0[2]),.dinb(w_Gid6_0[2]),.dout(n92),.clk(gclk));
	jxor g020(.dina(n92),.dinb(n91),.dout(n93),.clk(gclk));
	jxor g021(.dina(w_n93_0[1]),.dinb(n90),.dout(n94),.clk(gclk));
	jxor g022(.dina(w_Gid13_0[2]),.dinb(w_Gid12_0[1]),.dout(n95),.clk(gclk));
	jxor g023(.dina(w_Gid15_0[2]),.dinb(w_Gid14_0[2]),.dout(n96),.clk(gclk));
	jxor g024(.dina(n96),.dinb(n95),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_Gid23_0[1]),.dinb(w_Gid19_0[1]),.dout(n98),.clk(gclk));
	jxor g026(.dina(w_Gid31_0[2]),.dinb(w_Gid27_0[2]),.dout(n99),.clk(gclk));
	jxor g027(.dina(n99),.dinb(n98),.dout(n100),.clk(gclk));
	jxor g028(.dina(n100),.dinb(w_n97_0[1]),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n94),.dout(n102),.clk(gclk));
	jnot g030(.din(Gic6),.dout(n103),.clk(gclk));
	jor g031(.dina(w_n74_2[2]),.dinb(n103),.dout(n104),.clk(gclk));
	jxor g032(.dina(w_Gid1_0[2]),.dinb(w_Gid0_0[1]),.dout(n105),.clk(gclk));
	jxor g033(.dina(w_Gid3_0[2]),.dinb(w_Gid2_0[2]),.dout(n106),.clk(gclk));
	jxor g034(.dina(n106),.dinb(n105),.dout(n107),.clk(gclk));
	jxor g035(.dina(w_n107_0[1]),.dinb(n104),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_Gid9_0[2]),.dinb(w_Gid8_0[1]),.dout(n109),.clk(gclk));
	jxor g037(.dina(w_Gid11_0[2]),.dinb(w_Gid10_0[2]),.dout(n110),.clk(gclk));
	jxor g038(.dina(n110),.dinb(n109),.dout(n111),.clk(gclk));
	jxor g039(.dina(w_Gid22_0[1]),.dinb(w_Gid18_0[1]),.dout(n112),.clk(gclk));
	jxor g040(.dina(w_Gid30_0[2]),.dinb(w_Gid26_0[2]),.dout(n113),.clk(gclk));
	jxor g041(.dina(n113),.dinb(n112),.dout(n114),.clk(gclk));
	jxor g042(.dina(n114),.dinb(w_n111_0[1]),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(n108),.dout(n116),.clk(gclk));
	jnot g044(.din(w_n116_1[1]),.dout(n117),.clk(gclk));
	jand g045(.dina(w_n117_1[2]),.dinb(w_n102_1[1]),.dout(n118),.clk(gclk));
	jnot g046(.din(Gic4),.dout(n119),.clk(gclk));
	jor g047(.dina(w_n74_2[1]),.dinb(n119),.dout(n120),.clk(gclk));
	jxor g048(.dina(n120),.dinb(w_n93_0[0]),.dout(n121),.clk(gclk));
	jxor g049(.dina(w_Gid20_0[1]),.dinb(w_Gid16_0[1]),.dout(n122),.clk(gclk));
	jxor g050(.dina(w_Gid28_0[2]),.dinb(w_Gid24_0[2]),.dout(n123),.clk(gclk));
	jxor g051(.dina(n123),.dinb(n122),.dout(n124),.clk(gclk));
	jxor g052(.dina(n124),.dinb(w_n107_0[0]),.dout(n125),.clk(gclk));
	jxor g053(.dina(n125),.dinb(n121),.dout(n126),.clk(gclk));
	jnot g054(.din(w_n126_1[1]),.dout(n127),.clk(gclk));
	jnot g055(.din(Gic5),.dout(n128),.clk(gclk));
	jor g056(.dina(w_n74_2[0]),.dinb(n128),.dout(n129),.clk(gclk));
	jxor g057(.dina(n129),.dinb(w_n97_0[0]),.dout(n130),.clk(gclk));
	jxor g058(.dina(w_Gid21_0[1]),.dinb(w_Gid17_0[1]),.dout(n131),.clk(gclk));
	jxor g059(.dina(w_Gid29_0[2]),.dinb(w_Gid25_0[2]),.dout(n132),.clk(gclk));
	jxor g060(.dina(n132),.dinb(n131),.dout(n133),.clk(gclk));
	jxor g061(.dina(n133),.dinb(w_n111_0[0]),.dout(n134),.clk(gclk));
	jxor g062(.dina(n134),.dinb(n130),.dout(n135),.clk(gclk));
	jand g063(.dina(w_n135_1[1]),.dinb(w_n127_1[2]),.dout(n136),.clk(gclk));
	jnot g064(.din(Gic1),.dout(n137),.clk(gclk));
	jor g065(.dina(w_n74_1[2]),.dinb(n137),.dout(n138),.clk(gclk));
	jxor g066(.dina(w_Gid29_0[1]),.dinb(w_Gid28_0[1]),.dout(n139),.clk(gclk));
	jxor g067(.dina(w_Gid31_0[1]),.dinb(w_Gid30_0[1]),.dout(n140),.clk(gclk));
	jxor g068(.dina(n140),.dinb(n139),.dout(n141),.clk(gclk));
	jxor g069(.dina(w_n141_0[1]),.dinb(n138),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_Gid25_0[1]),.dinb(w_Gid24_0[1]),.dout(n143),.clk(gclk));
	jxor g071(.dina(w_Gid27_0[1]),.dinb(w_Gid26_0[1]),.dout(n144),.clk(gclk));
	jxor g072(.dina(n144),.dinb(n143),.dout(n145),.clk(gclk));
	jxor g073(.dina(w_Gid5_0[1]),.dinb(w_Gid1_0[1]),.dout(n146),.clk(gclk));
	jxor g074(.dina(w_Gid13_0[1]),.dinb(w_Gid9_0[1]),.dout(n147),.clk(gclk));
	jxor g075(.dina(n147),.dinb(n146),.dout(n148),.clk(gclk));
	jxor g076(.dina(n148),.dinb(w_n145_0[1]),.dout(n149),.clk(gclk));
	jxor g077(.dina(n149),.dinb(n142),.dout(n150),.clk(gclk));
	jxor g078(.dina(w_n150_1[1]),.dinb(w_n87_1[0]),.dout(n151),.clk(gclk));
	jnot g079(.din(Gic3),.dout(n152),.clk(gclk));
	jor g080(.dina(w_n74_1[1]),.dinb(n152),.dout(n153),.clk(gclk));
	jxor g081(.dina(n153),.dinb(w_n85_0[0]),.dout(n154),.clk(gclk));
	jxor g082(.dina(w_Gid7_0[1]),.dinb(w_Gid3_0[1]),.dout(n155),.clk(gclk));
	jxor g083(.dina(w_Gid15_0[1]),.dinb(w_Gid11_0[1]),.dout(n156),.clk(gclk));
	jxor g084(.dina(n156),.dinb(n155),.dout(n157),.clk(gclk));
	jxor g085(.dina(n157),.dinb(w_n141_0[0]),.dout(n158),.clk(gclk));
	jxor g086(.dina(n158),.dinb(n154),.dout(n159),.clk(gclk));
	jnot g087(.din(Gic2),.dout(n160),.clk(gclk));
	jor g088(.dina(w_n74_1[0]),.dinb(n160),.dout(n161),.clk(gclk));
	jxor g089(.dina(n161),.dinb(w_n78_0[0]),.dout(n162),.clk(gclk));
	jxor g090(.dina(w_Gid6_0[1]),.dinb(w_Gid2_0[1]),.dout(n163),.clk(gclk));
	jxor g091(.dina(w_Gid14_0[1]),.dinb(w_Gid10_0[1]),.dout(n164),.clk(gclk));
	jxor g092(.dina(n164),.dinb(n163),.dout(n165),.clk(gclk));
	jxor g093(.dina(n165),.dinb(w_n145_0[0]),.dout(n166),.clk(gclk));
	jxor g094(.dina(n166),.dinb(n162),.dout(n167),.clk(gclk));
	jand g095(.dina(w_n167_1[1]),.dinb(w_n159_1[1]),.dout(n168),.clk(gclk));
	jand g096(.dina(n168),.dinb(n151),.dout(n169),.clk(gclk));
	jxor g097(.dina(w_n167_1[0]),.dinb(w_n159_1[0]),.dout(n170),.clk(gclk));
	jand g098(.dina(w_n150_1[0]),.dinb(w_n87_0[2]),.dout(n171),.clk(gclk));
	jand g099(.dina(n171),.dinb(n170),.dout(n172),.clk(gclk));
	jor g100(.dina(n172),.dinb(n169),.dout(n173),.clk(gclk));
	jand g101(.dina(w_n173_0[2]),.dinb(w_dff_B_7YbQlWtC6_1),.dout(n174),.clk(gclk));
	jand g102(.dina(w_n174_0[1]),.dinb(w_n118_0[1]),.dout(n175),.clk(gclk));
	jand g103(.dina(w_n175_1[1]),.dinb(w_n88_1[2]),.dout(n176),.clk(gclk));
	jxor g104(.dina(n176),.dinb(w_Gid0_0[0]),.dout(God0),.clk(gclk));
	jnot g105(.din(w_n150_0[2]),.dout(n178),.clk(gclk));
	jand g106(.dina(w_n175_1[0]),.dinb(w_n178_1[2]),.dout(n179),.clk(gclk));
	jxor g107(.dina(n179),.dinb(w_Gid1_0[0]),.dout(God1),.clk(gclk));
	jnot g108(.din(w_n167_0[2]),.dout(n181),.clk(gclk));
	jand g109(.dina(w_n175_0[2]),.dinb(w_n181_1[2]),.dout(n182),.clk(gclk));
	jxor g110(.dina(n182),.dinb(w_Gid2_0[0]),.dout(God2),.clk(gclk));
	jnot g111(.din(w_n159_0[2]),.dout(n184),.clk(gclk));
	jand g112(.dina(w_n175_0[1]),.dinb(w_n184_1[2]),.dout(n185),.clk(gclk));
	jxor g113(.dina(n185),.dinb(w_Gid3_0[0]),.dout(God3),.clk(gclk));
	jnot g114(.din(w_n102_1[0]),.dout(n187),.clk(gclk));
	jand g115(.dina(w_n116_1[0]),.dinb(w_n187_1[2]),.dout(n188),.clk(gclk));
	jand g116(.dina(w_n188_0[1]),.dinb(w_n174_0[0]),.dout(n189),.clk(gclk));
	jand g117(.dina(w_n189_1[1]),.dinb(w_n88_1[1]),.dout(n190),.clk(gclk));
	jxor g118(.dina(n190),.dinb(w_Gid4_0[0]),.dout(God4),.clk(gclk));
	jand g119(.dina(w_n189_1[0]),.dinb(w_n178_1[1]),.dout(n192),.clk(gclk));
	jxor g120(.dina(n192),.dinb(w_Gid5_0[0]),.dout(God5),.clk(gclk));
	jand g121(.dina(w_n189_0[2]),.dinb(w_n181_1[1]),.dout(n194),.clk(gclk));
	jxor g122(.dina(n194),.dinb(w_Gid6_0[0]),.dout(God6),.clk(gclk));
	jand g123(.dina(w_n189_0[1]),.dinb(w_n184_1[1]),.dout(n196),.clk(gclk));
	jxor g124(.dina(n196),.dinb(w_Gid7_0[0]),.dout(God7),.clk(gclk));
	jnot g125(.din(w_n135_1[0]),.dout(n198),.clk(gclk));
	jand g126(.dina(w_n198_1[2]),.dinb(w_n126_1[0]),.dout(n199),.clk(gclk));
	jand g127(.dina(w_n199_0[1]),.dinb(w_n118_0[0]),.dout(n200),.clk(gclk));
	jand g128(.dina(n200),.dinb(w_n173_0[1]),.dout(n201),.clk(gclk));
	jand g129(.dina(w_n201_1[1]),.dinb(w_n88_1[0]),.dout(n202),.clk(gclk));
	jxor g130(.dina(n202),.dinb(w_Gid8_0[0]),.dout(w_dff_A_xZiBlxD60_2),.clk(gclk));
	jand g131(.dina(w_n201_1[0]),.dinb(w_n178_1[0]),.dout(n204),.clk(gclk));
	jxor g132(.dina(n204),.dinb(w_Gid9_0[0]),.dout(w_dff_A_GC3Ur5fC0_2),.clk(gclk));
	jand g133(.dina(w_n201_0[2]),.dinb(w_n181_1[0]),.dout(n206),.clk(gclk));
	jxor g134(.dina(n206),.dinb(w_Gid10_0[0]),.dout(w_dff_A_qT9JmB3C5_2),.clk(gclk));
	jand g135(.dina(w_n201_0[1]),.dinb(w_n184_1[0]),.dout(n208),.clk(gclk));
	jxor g136(.dina(n208),.dinb(w_Gid11_0[0]),.dout(w_dff_A_2iNFlhGO6_2),.clk(gclk));
	jand g137(.dina(w_n199_0[0]),.dinb(w_n188_0[0]),.dout(n210),.clk(gclk));
	jand g138(.dina(n210),.dinb(w_n173_0[0]),.dout(n211),.clk(gclk));
	jand g139(.dina(w_n211_1[1]),.dinb(w_n88_0[2]),.dout(n212),.clk(gclk));
	jxor g140(.dina(n212),.dinb(w_Gid12_0[0]),.dout(w_dff_A_k1Z9d4Mf4_2),.clk(gclk));
	jand g141(.dina(w_n211_1[0]),.dinb(w_n178_0[2]),.dout(n214),.clk(gclk));
	jxor g142(.dina(n214),.dinb(w_Gid13_0[0]),.dout(w_dff_A_2woWXhQe4_2),.clk(gclk));
	jand g143(.dina(w_n211_0[2]),.dinb(w_n181_0[2]),.dout(n216),.clk(gclk));
	jxor g144(.dina(n216),.dinb(w_Gid14_0[0]),.dout(w_dff_A_02xLMDyO5_2),.clk(gclk));
	jand g145(.dina(w_n211_0[1]),.dinb(w_n184_0[2]),.dout(n218),.clk(gclk));
	jxor g146(.dina(n218),.dinb(w_Gid15_0[0]),.dout(w_dff_A_XsRivswP4_2),.clk(gclk));
	jand g147(.dina(w_n150_0[1]),.dinb(w_n88_0[1]),.dout(n220),.clk(gclk));
	jand g148(.dina(w_n181_0[1]),.dinb(w_n159_0[1]),.dout(n221),.clk(gclk));
	jxor g149(.dina(w_n116_0[2]),.dinb(w_n102_0[2]),.dout(n222),.clk(gclk));
	jand g150(.dina(w_n135_0[2]),.dinb(w_n126_0[2]),.dout(n223),.clk(gclk));
	jand g151(.dina(n223),.dinb(n222),.dout(n224),.clk(gclk));
	jxor g152(.dina(w_n135_0[1]),.dinb(w_n126_0[1]),.dout(n225),.clk(gclk));
	jand g153(.dina(w_n116_0[1]),.dinb(w_n102_0[1]),.dout(n226),.clk(gclk));
	jand g154(.dina(n226),.dinb(n225),.dout(n227),.clk(gclk));
	jor g155(.dina(n227),.dinb(n224),.dout(n228),.clk(gclk));
	jand g156(.dina(w_n228_0[1]),.dinb(w_dff_B_6rCY2ARc4_1),.dout(n229),.clk(gclk));
	jand g157(.dina(w_n229_0[1]),.dinb(w_n220_0[1]),.dout(n230),.clk(gclk));
	jand g158(.dina(w_n230_1[1]),.dinb(w_n127_1[1]),.dout(n231),.clk(gclk));
	jxor g159(.dina(n231),.dinb(w_Gid16_0[0]),.dout(God16),.clk(gclk));
	jand g160(.dina(w_n230_1[0]),.dinb(w_n198_1[1]),.dout(n233),.clk(gclk));
	jxor g161(.dina(n233),.dinb(w_Gid17_0[0]),.dout(God17),.clk(gclk));
	jand g162(.dina(w_n230_0[2]),.dinb(w_n117_1[1]),.dout(n235),.clk(gclk));
	jxor g163(.dina(n235),.dinb(w_Gid18_0[0]),.dout(God18),.clk(gclk));
	jand g164(.dina(w_n230_0[1]),.dinb(w_n187_1[1]),.dout(n237),.clk(gclk));
	jxor g165(.dina(n237),.dinb(w_Gid19_0[0]),.dout(God19),.clk(gclk));
	jand g166(.dina(w_n167_0[1]),.dinb(w_n184_0[1]),.dout(n239),.clk(gclk));
	jand g167(.dina(w_n228_0[0]),.dinb(w_dff_B_FleaHSHC9_1),.dout(n240),.clk(gclk));
	jand g168(.dina(w_n240_0[1]),.dinb(w_n220_0[0]),.dout(n241),.clk(gclk));
	jand g169(.dina(w_n241_1[1]),.dinb(w_n127_1[0]),.dout(n242),.clk(gclk));
	jxor g170(.dina(n242),.dinb(w_Gid20_0[0]),.dout(God20),.clk(gclk));
	jand g171(.dina(w_n241_1[0]),.dinb(w_n198_1[0]),.dout(n244),.clk(gclk));
	jxor g172(.dina(n244),.dinb(w_Gid21_0[0]),.dout(God21),.clk(gclk));
	jand g173(.dina(w_n241_0[2]),.dinb(w_n117_1[0]),.dout(n246),.clk(gclk));
	jxor g174(.dina(n246),.dinb(w_Gid22_0[0]),.dout(God22),.clk(gclk));
	jand g175(.dina(w_n241_0[1]),.dinb(w_n187_1[0]),.dout(n248),.clk(gclk));
	jxor g176(.dina(n248),.dinb(w_Gid23_0[0]),.dout(God23),.clk(gclk));
	jand g177(.dina(w_n178_0[1]),.dinb(w_n87_0[1]),.dout(n250),.clk(gclk));
	jand g178(.dina(w_n229_0[0]),.dinb(w_n250_0[1]),.dout(n251),.clk(gclk));
	jand g179(.dina(w_n251_1[1]),.dinb(w_n127_0[2]),.dout(n252),.clk(gclk));
	jxor g180(.dina(n252),.dinb(w_Gid24_0[0]),.dout(God24),.clk(gclk));
	jand g181(.dina(w_n251_1[0]),.dinb(w_n198_0[2]),.dout(n254),.clk(gclk));
	jxor g182(.dina(n254),.dinb(w_Gid25_0[0]),.dout(God25),.clk(gclk));
	jand g183(.dina(w_n251_0[2]),.dinb(w_n117_0[2]),.dout(n256),.clk(gclk));
	jxor g184(.dina(n256),.dinb(w_Gid26_0[0]),.dout(God26),.clk(gclk));
	jand g185(.dina(w_n251_0[1]),.dinb(w_n187_0[2]),.dout(n258),.clk(gclk));
	jxor g186(.dina(n258),.dinb(w_Gid27_0[0]),.dout(God27),.clk(gclk));
	jand g187(.dina(w_n240_0[0]),.dinb(w_n250_0[0]),.dout(n260),.clk(gclk));
	jand g188(.dina(w_n260_1[1]),.dinb(w_n127_0[1]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_Gid28_0[0]),.dout(God28),.clk(gclk));
	jand g190(.dina(w_n260_1[0]),.dinb(w_n198_0[1]),.dout(n263),.clk(gclk));
	jxor g191(.dina(n263),.dinb(w_Gid29_0[0]),.dout(God29),.clk(gclk));
	jand g192(.dina(w_n260_0[2]),.dinb(w_n117_0[1]),.dout(n265),.clk(gclk));
	jxor g193(.dina(n265),.dinb(w_Gid30_0[0]),.dout(God30),.clk(gclk));
	jand g194(.dina(w_n260_0[1]),.dinb(w_n187_0[1]),.dout(n267),.clk(gclk));
	jxor g195(.dina(n267),.dinb(w_Gid31_0[0]),.dout(God31),.clk(gclk));
	jspl3 jspl3_w_Gid0_0(.douta(w_dff_A_YsUNoZov4_0),.doutb(w_Gid0_0[1]),.doutc(w_Gid0_0[2]),.din(Gid0));
	jspl3 jspl3_w_Gid1_0(.douta(w_dff_A_juUxwNZX6_0),.doutb(w_Gid1_0[1]),.doutc(w_Gid1_0[2]),.din(Gid1));
	jspl3 jspl3_w_Gid2_0(.douta(w_dff_A_lFxY92ZG4_0),.doutb(w_Gid2_0[1]),.doutc(w_Gid2_0[2]),.din(Gid2));
	jspl3 jspl3_w_Gid3_0(.douta(w_dff_A_Ehs49Qsy1_0),.doutb(w_Gid3_0[1]),.doutc(w_Gid3_0[2]),.din(Gid3));
	jspl3 jspl3_w_Gid4_0(.douta(w_dff_A_ZgwJAPqV3_0),.doutb(w_Gid4_0[1]),.doutc(w_Gid4_0[2]),.din(Gid4));
	jspl3 jspl3_w_Gid5_0(.douta(w_dff_A_BfT7Vhzc5_0),.doutb(w_Gid5_0[1]),.doutc(w_Gid5_0[2]),.din(Gid5));
	jspl3 jspl3_w_Gid6_0(.douta(w_dff_A_sNMh06Yt4_0),.doutb(w_Gid6_0[1]),.doutc(w_Gid6_0[2]),.din(Gid6));
	jspl3 jspl3_w_Gid7_0(.douta(w_dff_A_kkrNQRKE5_0),.doutb(w_Gid7_0[1]),.doutc(w_Gid7_0[2]),.din(Gid7));
	jspl3 jspl3_w_Gid8_0(.douta(w_dff_A_QXExpRAt1_0),.doutb(w_Gid8_0[1]),.doutc(w_Gid8_0[2]),.din(Gid8));
	jspl3 jspl3_w_Gid9_0(.douta(w_dff_A_QN1AQoE70_0),.doutb(w_Gid9_0[1]),.doutc(w_Gid9_0[2]),.din(Gid9));
	jspl3 jspl3_w_Gid10_0(.douta(w_dff_A_pxZO4WQg6_0),.doutb(w_Gid10_0[1]),.doutc(w_Gid10_0[2]),.din(Gid10));
	jspl3 jspl3_w_Gid11_0(.douta(w_dff_A_ygrfhaGE6_0),.doutb(w_Gid11_0[1]),.doutc(w_Gid11_0[2]),.din(Gid11));
	jspl3 jspl3_w_Gid12_0(.douta(w_dff_A_qYT5kUyt1_0),.doutb(w_Gid12_0[1]),.doutc(w_Gid12_0[2]),.din(Gid12));
	jspl3 jspl3_w_Gid13_0(.douta(w_dff_A_Kr1W6KUY5_0),.doutb(w_Gid13_0[1]),.doutc(w_Gid13_0[2]),.din(Gid13));
	jspl3 jspl3_w_Gid14_0(.douta(w_dff_A_aOH4rWq78_0),.doutb(w_Gid14_0[1]),.doutc(w_Gid14_0[2]),.din(Gid14));
	jspl3 jspl3_w_Gid15_0(.douta(w_dff_A_n9T6JgZ27_0),.doutb(w_Gid15_0[1]),.doutc(w_Gid15_0[2]),.din(Gid15));
	jspl3 jspl3_w_Gid16_0(.douta(w_dff_A_XmRrv8nG7_0),.doutb(w_Gid16_0[1]),.doutc(w_Gid16_0[2]),.din(Gid16));
	jspl3 jspl3_w_Gid17_0(.douta(w_dff_A_OVz3kojF3_0),.doutb(w_Gid17_0[1]),.doutc(w_Gid17_0[2]),.din(Gid17));
	jspl3 jspl3_w_Gid18_0(.douta(w_dff_A_PaXUWnuJ3_0),.doutb(w_Gid18_0[1]),.doutc(w_Gid18_0[2]),.din(Gid18));
	jspl3 jspl3_w_Gid19_0(.douta(w_dff_A_LEJdWwnh0_0),.doutb(w_Gid19_0[1]),.doutc(w_Gid19_0[2]),.din(Gid19));
	jspl3 jspl3_w_Gid20_0(.douta(w_dff_A_I7zSl4Oo8_0),.doutb(w_Gid20_0[1]),.doutc(w_Gid20_0[2]),.din(Gid20));
	jspl3 jspl3_w_Gid21_0(.douta(w_dff_A_y3d5rboI7_0),.doutb(w_Gid21_0[1]),.doutc(w_Gid21_0[2]),.din(Gid21));
	jspl3 jspl3_w_Gid22_0(.douta(w_dff_A_v52rLRPg7_0),.doutb(w_Gid22_0[1]),.doutc(w_Gid22_0[2]),.din(Gid22));
	jspl3 jspl3_w_Gid23_0(.douta(w_dff_A_bQX9gF2S9_0),.doutb(w_Gid23_0[1]),.doutc(w_Gid23_0[2]),.din(Gid23));
	jspl3 jspl3_w_Gid24_0(.douta(w_dff_A_E22RhgI36_0),.doutb(w_Gid24_0[1]),.doutc(w_Gid24_0[2]),.din(Gid24));
	jspl3 jspl3_w_Gid25_0(.douta(w_dff_A_lwZhi6iY6_0),.doutb(w_Gid25_0[1]),.doutc(w_Gid25_0[2]),.din(Gid25));
	jspl3 jspl3_w_Gid26_0(.douta(w_dff_A_hNLQDEle0_0),.doutb(w_Gid26_0[1]),.doutc(w_Gid26_0[2]),.din(Gid26));
	jspl3 jspl3_w_Gid27_0(.douta(w_dff_A_MO03c5xV3_0),.doutb(w_Gid27_0[1]),.doutc(w_Gid27_0[2]),.din(Gid27));
	jspl3 jspl3_w_Gid28_0(.douta(w_dff_A_JaGskUwi2_0),.doutb(w_Gid28_0[1]),.doutc(w_Gid28_0[2]),.din(Gid28));
	jspl3 jspl3_w_Gid29_0(.douta(w_dff_A_ZXZxQSbT4_0),.doutb(w_Gid29_0[1]),.doutc(w_Gid29_0[2]),.din(Gid29));
	jspl3 jspl3_w_Gid30_0(.douta(w_dff_A_3GoHoAV63_0),.doutb(w_Gid30_0[1]),.doutc(w_Gid30_0[2]),.din(Gid30));
	jspl3 jspl3_w_Gid31_0(.douta(w_dff_A_wLmNjqFi8_0),.doutb(w_Gid31_0[1]),.doutc(w_Gid31_0[2]),.din(Gid31));
	jspl3 jspl3_w_n74_0(.douta(w_n74_0[0]),.doutb(w_n74_0[1]),.doutc(w_n74_0[2]),.din(n74));
	jspl3 jspl3_w_n74_1(.douta(w_n74_1[0]),.doutb(w_n74_1[1]),.doutc(w_n74_1[2]),.din(w_n74_0[0]));
	jspl3 jspl3_w_n74_2(.douta(w_n74_2[0]),.doutb(w_n74_2[1]),.doutc(w_n74_2[2]),.din(w_n74_0[1]));
	jspl jspl_w_n74_3(.douta(w_n74_3[0]),.doutb(w_n74_3[1]),.din(w_n74_0[2]));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl3 jspl3_w_n87_0(.douta(w_n87_0[0]),.doutb(w_dff_A_JHfHeD4W6_1),.doutc(w_n87_0[2]),.din(n87));
	jspl jspl_w_n87_1(.douta(w_n87_1[0]),.doutb(w_n87_1[1]),.din(w_n87_0[0]));
	jspl3 jspl3_w_n88_0(.douta(w_dff_A_uWCDLAHs3_0),.doutb(w_n88_0[1]),.doutc(w_dff_A_894mahDr7_2),.din(n88));
	jspl3 jspl3_w_n88_1(.douta(w_n88_1[0]),.doutb(w_dff_A_QrMOdnYP1_1),.doutc(w_dff_A_1s1teyGQ6_2),.din(w_n88_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n97_0(.douta(w_n97_0[0]),.doutb(w_n97_0[1]),.din(n97));
	jspl3 jspl3_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.doutc(w_n102_0[2]),.din(n102));
	jspl jspl_w_n102_1(.douta(w_n102_1[0]),.doutb(w_dff_A_HEyAYzEs7_1),.din(w_n102_0[0]));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n111_0(.douta(w_n111_0[0]),.doutb(w_n111_0[1]),.din(n111));
	jspl3 jspl3_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.doutc(w_n116_0[2]),.din(n116));
	jspl jspl_w_n116_1(.douta(w_dff_A_3gCewhSK3_0),.doutb(w_n116_1[1]),.din(w_n116_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_7RdF8kzx1_1),.doutc(w_dff_A_NJnKpFfd4_2),.din(n117));
	jspl3 jspl3_w_n117_1(.douta(w_dff_A_tY6nUX7m2_0),.doutb(w_dff_A_P80ByBBx9_1),.doutc(w_n117_1[2]),.din(w_n117_0[0]));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_dff_A_BZxubKaJ9_1),.din(n118));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl jspl_w_n126_1(.douta(w_dff_A_GbwvgkeW8_0),.doutb(w_n126_1[1]),.din(w_n126_0[0]));
	jspl3 jspl3_w_n127_0(.douta(w_n127_0[0]),.doutb(w_dff_A_XRGzg8M38_1),.doutc(w_dff_A_Ytk3OuDc2_2),.din(n127));
	jspl3 jspl3_w_n127_1(.douta(w_dff_A_GtwcM2vK5_0),.doutb(w_dff_A_o3YawC4w9_1),.doutc(w_n127_1[2]),.din(w_n127_0[0]));
	jspl3 jspl3_w_n135_0(.douta(w_n135_0[0]),.doutb(w_n135_0[1]),.doutc(w_n135_0[2]),.din(n135));
	jspl jspl_w_n135_1(.douta(w_n135_1[0]),.doutb(w_dff_A_Rj5xck4f5_1),.din(w_n135_0[0]));
	jspl jspl_w_n141_0(.douta(w_n141_0[0]),.doutb(w_n141_0[1]),.din(n141));
	jspl jspl_w_n145_0(.douta(w_n145_0[0]),.doutb(w_n145_0[1]),.din(n145));
	jspl3 jspl3_w_n150_0(.douta(w_n150_0[0]),.doutb(w_dff_A_ZIJzp40A1_1),.doutc(w_n150_0[2]),.din(n150));
	jspl jspl_w_n150_1(.douta(w_n150_1[0]),.doutb(w_n150_1[1]),.din(w_n150_0[0]));
	jspl3 jspl3_w_n159_0(.douta(w_n159_0[0]),.doutb(w_dff_A_MfDVjbvw0_1),.doutc(w_n159_0[2]),.din(n159));
	jspl jspl_w_n159_1(.douta(w_n159_1[0]),.doutb(w_n159_1[1]),.din(w_n159_0[0]));
	jspl3 jspl3_w_n167_0(.douta(w_n167_0[0]),.doutb(w_dff_A_LLiTtz3t7_1),.doutc(w_n167_0[2]),.din(n167));
	jspl jspl_w_n167_1(.douta(w_n167_1[0]),.doutb(w_n167_1[1]),.din(w_n167_0[0]));
	jspl3 jspl3_w_n173_0(.douta(w_n173_0[0]),.doutb(w_n173_0[1]),.doutc(w_n173_0[2]),.din(n173));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.din(n174));
	jspl3 jspl3_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.doutc(w_n175_0[2]),.din(n175));
	jspl jspl_w_n175_1(.douta(w_n175_1[0]),.doutb(w_n175_1[1]),.din(w_n175_0[0]));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_mUG1xxPk9_0),.doutb(w_n178_0[1]),.doutc(w_dff_A_2hdwB6Lq7_2),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_dff_A_5NSGo9VV3_1),.doutc(w_dff_A_CL6Ni2838_2),.din(w_n178_0[0]));
	jspl3 jspl3_w_n181_0(.douta(w_dff_A_HqSlzSuR4_0),.doutb(w_n181_0[1]),.doutc(w_dff_A_TgHx8kkL7_2),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_dff_A_VS7e9OZH6_1),.doutc(w_dff_A_n7BkOgZh9_2),.din(w_n181_0[0]));
	jspl3 jspl3_w_n184_0(.douta(w_dff_A_6NQTQiCa1_0),.doutb(w_n184_0[1]),.doutc(w_dff_A_OEJiDYKX7_2),.din(n184));
	jspl3 jspl3_w_n184_1(.douta(w_n184_1[0]),.doutb(w_dff_A_uPgEDf7R4_1),.doutc(w_dff_A_fzY6eBTi1_2),.din(w_n184_0[0]));
	jspl3 jspl3_w_n187_0(.douta(w_n187_0[0]),.doutb(w_dff_A_uBkBXEWl3_1),.doutc(w_dff_A_H1KiPvTH0_2),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_dff_A_apFlQxxA3_0),.doutb(w_dff_A_GZUUKd7t2_1),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_dff_A_48Somc154_1),.din(n188));
	jspl3 jspl3_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.doutc(w_n189_0[2]),.din(n189));
	jspl jspl_w_n189_1(.douta(w_n189_1[0]),.doutb(w_n189_1[1]),.din(w_n189_0[0]));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_dff_A_Ts1tV0HU8_1),.doutc(w_dff_A_QWvYTr0x0_2),.din(n198));
	jspl3 jspl3_w_n198_1(.douta(w_dff_A_gKqMLxcP6_0),.doutb(w_dff_A_845KEc5h4_1),.doutc(w_n198_1[2]),.din(w_n198_0[0]));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl3 jspl3_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.doutc(w_n201_0[2]),.din(n201));
	jspl jspl_w_n201_1(.douta(w_n201_1[0]),.doutb(w_n201_1[1]),.din(w_n201_0[0]));
	jspl3 jspl3_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.doutc(w_n211_0[2]),.din(n211));
	jspl jspl_w_n211_1(.douta(w_n211_1[0]),.doutb(w_n211_1[1]),.din(w_n211_0[0]));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(w_dff_B_9hY9tMd39_2));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.din(n229));
	jspl3 jspl3_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.doutc(w_n230_0[2]),.din(n230));
	jspl jspl_w_n230_1(.douta(w_n230_1[0]),.doutb(w_n230_1[1]),.din(w_n230_0[0]));
	jspl jspl_w_n240_0(.douta(w_n240_0[0]),.doutb(w_n240_0[1]),.din(n240));
	jspl3 jspl3_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.doutc(w_n241_0[2]),.din(n241));
	jspl jspl_w_n241_1(.douta(w_n241_1[0]),.doutb(w_n241_1[1]),.din(w_n241_0[0]));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(w_dff_B_97l74v724_2));
	jspl3 jspl3_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.doutc(w_n251_0[2]),.din(n251));
	jspl jspl_w_n251_1(.douta(w_n251_1[0]),.doutb(w_n251_1[1]),.din(w_n251_0[0]));
	jspl3 jspl3_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.doutc(w_n260_0[2]),.din(n260));
	jspl jspl_w_n260_1(.douta(w_n260_1[0]),.doutb(w_n260_1[1]),.din(w_n260_0[0]));
	jdff dff_B_7YbQlWtC6_1(.din(n136),.dout(w_dff_B_7YbQlWtC6_1),.clk(gclk));
	jdff dff_A_QrMOdnYP1_1(.dout(w_n88_1[1]),.din(w_dff_A_QrMOdnYP1_1),.clk(gclk));
	jdff dff_A_1s1teyGQ6_2(.dout(w_n88_1[2]),.din(w_dff_A_1s1teyGQ6_2),.clk(gclk));
	jdff dff_A_5NSGo9VV3_1(.dout(w_n178_1[1]),.din(w_dff_A_5NSGo9VV3_1),.clk(gclk));
	jdff dff_A_CL6Ni2838_2(.dout(w_n178_1[2]),.din(w_dff_A_CL6Ni2838_2),.clk(gclk));
	jdff dff_A_VS7e9OZH6_1(.dout(w_n181_1[1]),.din(w_dff_A_VS7e9OZH6_1),.clk(gclk));
	jdff dff_A_n7BkOgZh9_2(.dout(w_n181_1[2]),.din(w_dff_A_n7BkOgZh9_2),.clk(gclk));
	jdff dff_A_mFpqzfM30_1(.dout(w_n118_0[1]),.din(w_dff_A_mFpqzfM30_1),.clk(gclk));
	jdff dff_A_BZxubKaJ9_1(.dout(w_dff_A_mFpqzfM30_1),.din(w_dff_A_BZxubKaJ9_1),.clk(gclk));
	jdff dff_A_uPgEDf7R4_1(.dout(w_n184_1[1]),.din(w_dff_A_uPgEDf7R4_1),.clk(gclk));
	jdff dff_A_fzY6eBTi1_2(.dout(w_n184_1[2]),.din(w_dff_A_fzY6eBTi1_2),.clk(gclk));
	jdff dff_A_SXflDD7T8_1(.dout(w_n188_0[1]),.din(w_dff_A_SXflDD7T8_1),.clk(gclk));
	jdff dff_A_48Somc154_1(.dout(w_dff_A_SXflDD7T8_1),.din(w_dff_A_48Somc154_1),.clk(gclk));
	jdff dff_A_lwhZyFww2_0(.dout(w_n127_1[0]),.din(w_dff_A_lwhZyFww2_0),.clk(gclk));
	jdff dff_A_lhsPZKHs4_0(.dout(w_dff_A_lwhZyFww2_0),.din(w_dff_A_lhsPZKHs4_0),.clk(gclk));
	jdff dff_A_iALwGt6S2_0(.dout(w_dff_A_lhsPZKHs4_0),.din(w_dff_A_iALwGt6S2_0),.clk(gclk));
	jdff dff_A_GtwcM2vK5_0(.dout(w_dff_A_iALwGt6S2_0),.din(w_dff_A_GtwcM2vK5_0),.clk(gclk));
	jdff dff_A_PHiG1CSh7_1(.dout(w_n127_1[1]),.din(w_dff_A_PHiG1CSh7_1),.clk(gclk));
	jdff dff_A_SMJgTvvT1_1(.dout(w_dff_A_PHiG1CSh7_1),.din(w_dff_A_SMJgTvvT1_1),.clk(gclk));
	jdff dff_A_ZeB9MUyM2_1(.dout(w_dff_A_SMJgTvvT1_1),.din(w_dff_A_ZeB9MUyM2_1),.clk(gclk));
	jdff dff_A_o3YawC4w9_1(.dout(w_dff_A_ZeB9MUyM2_1),.din(w_dff_A_o3YawC4w9_1),.clk(gclk));
	jdff dff_A_VJy4WXiw8_0(.dout(w_n198_1[0]),.din(w_dff_A_VJy4WXiw8_0),.clk(gclk));
	jdff dff_A_dGU7Q6J78_0(.dout(w_dff_A_VJy4WXiw8_0),.din(w_dff_A_dGU7Q6J78_0),.clk(gclk));
	jdff dff_A_4R7B6Wh38_0(.dout(w_dff_A_dGU7Q6J78_0),.din(w_dff_A_4R7B6Wh38_0),.clk(gclk));
	jdff dff_A_gKqMLxcP6_0(.dout(w_dff_A_4R7B6Wh38_0),.din(w_dff_A_gKqMLxcP6_0),.clk(gclk));
	jdff dff_A_JFpFKBNG1_1(.dout(w_n198_1[1]),.din(w_dff_A_JFpFKBNG1_1),.clk(gclk));
	jdff dff_A_VeDNxiOF6_1(.dout(w_dff_A_JFpFKBNG1_1),.din(w_dff_A_VeDNxiOF6_1),.clk(gclk));
	jdff dff_A_UKrSRaEl5_1(.dout(w_dff_A_VeDNxiOF6_1),.din(w_dff_A_UKrSRaEl5_1),.clk(gclk));
	jdff dff_A_845KEc5h4_1(.dout(w_dff_A_UKrSRaEl5_1),.din(w_dff_A_845KEc5h4_1),.clk(gclk));
	jdff dff_A_8WS4zO9O3_0(.dout(w_n117_1[0]),.din(w_dff_A_8WS4zO9O3_0),.clk(gclk));
	jdff dff_A_OaONNhR07_0(.dout(w_dff_A_8WS4zO9O3_0),.din(w_dff_A_OaONNhR07_0),.clk(gclk));
	jdff dff_A_Qvsf2YyU6_0(.dout(w_dff_A_OaONNhR07_0),.din(w_dff_A_Qvsf2YyU6_0),.clk(gclk));
	jdff dff_A_tY6nUX7m2_0(.dout(w_dff_A_Qvsf2YyU6_0),.din(w_dff_A_tY6nUX7m2_0),.clk(gclk));
	jdff dff_A_4VRf9T5Y7_1(.dout(w_n117_1[1]),.din(w_dff_A_4VRf9T5Y7_1),.clk(gclk));
	jdff dff_A_MNpC9Wjq8_1(.dout(w_dff_A_4VRf9T5Y7_1),.din(w_dff_A_MNpC9Wjq8_1),.clk(gclk));
	jdff dff_A_snKzvNyW6_1(.dout(w_dff_A_MNpC9Wjq8_1),.din(w_dff_A_snKzvNyW6_1),.clk(gclk));
	jdff dff_A_P80ByBBx9_1(.dout(w_dff_A_snKzvNyW6_1),.din(w_dff_A_P80ByBBx9_1),.clk(gclk));
	jdff dff_B_1nPWFy1U6_2(.din(n220),.dout(w_dff_B_1nPWFy1U6_2),.clk(gclk));
	jdff dff_B_9hY9tMd39_2(.din(w_dff_B_1nPWFy1U6_2),.dout(w_dff_B_9hY9tMd39_2),.clk(gclk));
	jdff dff_A_B92hbzQf5_0(.dout(w_n88_0[0]),.din(w_dff_A_B92hbzQf5_0),.clk(gclk));
	jdff dff_A_VpUnDeto3_0(.dout(w_dff_A_B92hbzQf5_0),.din(w_dff_A_VpUnDeto3_0),.clk(gclk));
	jdff dff_A_uWCDLAHs3_0(.dout(w_dff_A_VpUnDeto3_0),.din(w_dff_A_uWCDLAHs3_0),.clk(gclk));
	jdff dff_A_t38aZdH66_2(.dout(w_n88_0[2]),.din(w_dff_A_t38aZdH66_2),.clk(gclk));
	jdff dff_A_c0SnWTV59_2(.dout(w_dff_A_t38aZdH66_2),.din(w_dff_A_c0SnWTV59_2),.clk(gclk));
	jdff dff_A_894mahDr7_2(.dout(w_dff_A_c0SnWTV59_2),.din(w_dff_A_894mahDr7_2),.clk(gclk));
	jdff dff_A_Czs4lalI4_0(.dout(w_n187_1[0]),.din(w_dff_A_Czs4lalI4_0),.clk(gclk));
	jdff dff_A_osHw9K8I5_0(.dout(w_dff_A_Czs4lalI4_0),.din(w_dff_A_osHw9K8I5_0),.clk(gclk));
	jdff dff_A_dM6bzT9h7_0(.dout(w_dff_A_osHw9K8I5_0),.din(w_dff_A_dM6bzT9h7_0),.clk(gclk));
	jdff dff_A_apFlQxxA3_0(.dout(w_dff_A_dM6bzT9h7_0),.din(w_dff_A_apFlQxxA3_0),.clk(gclk));
	jdff dff_A_yjiHvioF7_1(.dout(w_n187_1[1]),.din(w_dff_A_yjiHvioF7_1),.clk(gclk));
	jdff dff_A_9HYyYcwz2_1(.dout(w_dff_A_yjiHvioF7_1),.din(w_dff_A_9HYyYcwz2_1),.clk(gclk));
	jdff dff_A_WXJKU94Y1_1(.dout(w_dff_A_9HYyYcwz2_1),.din(w_dff_A_WXJKU94Y1_1),.clk(gclk));
	jdff dff_A_GZUUKd7t2_1(.dout(w_dff_A_WXJKU94Y1_1),.din(w_dff_A_GZUUKd7t2_1),.clk(gclk));
	jdff dff_B_6rCY2ARc4_1(.din(n221),.dout(w_dff_B_6rCY2ARc4_1),.clk(gclk));
	jdff dff_A_rmJkwMMt6_0(.dout(w_n181_0[0]),.din(w_dff_A_rmJkwMMt6_0),.clk(gclk));
	jdff dff_A_Hxld7UWi4_0(.dout(w_dff_A_rmJkwMMt6_0),.din(w_dff_A_Hxld7UWi4_0),.clk(gclk));
	jdff dff_A_HqSlzSuR4_0(.dout(w_dff_A_Hxld7UWi4_0),.din(w_dff_A_HqSlzSuR4_0),.clk(gclk));
	jdff dff_A_A0GkoZMn1_2(.dout(w_n181_0[2]),.din(w_dff_A_A0GkoZMn1_2),.clk(gclk));
	jdff dff_A_sJHs71t46_2(.dout(w_dff_A_A0GkoZMn1_2),.din(w_dff_A_sJHs71t46_2),.clk(gclk));
	jdff dff_A_TgHx8kkL7_2(.dout(w_dff_A_sJHs71t46_2),.din(w_dff_A_TgHx8kkL7_2),.clk(gclk));
	jdff dff_A_Oc2hW7pF6_1(.dout(w_n127_0[1]),.din(w_dff_A_Oc2hW7pF6_1),.clk(gclk));
	jdff dff_A_ckuUy3Ub8_1(.dout(w_dff_A_Oc2hW7pF6_1),.din(w_dff_A_ckuUy3Ub8_1),.clk(gclk));
	jdff dff_A_AXsjO57F2_1(.dout(w_dff_A_ckuUy3Ub8_1),.din(w_dff_A_AXsjO57F2_1),.clk(gclk));
	jdff dff_A_XRGzg8M38_1(.dout(w_dff_A_AXsjO57F2_1),.din(w_dff_A_XRGzg8M38_1),.clk(gclk));
	jdff dff_A_oaafBjdD2_2(.dout(w_n127_0[2]),.din(w_dff_A_oaafBjdD2_2),.clk(gclk));
	jdff dff_A_GFvLG8uw0_2(.dout(w_dff_A_oaafBjdD2_2),.din(w_dff_A_GFvLG8uw0_2),.clk(gclk));
	jdff dff_A_Jvgnk5390_2(.dout(w_dff_A_GFvLG8uw0_2),.din(w_dff_A_Jvgnk5390_2),.clk(gclk));
	jdff dff_A_Ytk3OuDc2_2(.dout(w_dff_A_Jvgnk5390_2),.din(w_dff_A_Ytk3OuDc2_2),.clk(gclk));
	jdff dff_A_GbwvgkeW8_0(.dout(w_n126_1[0]),.din(w_dff_A_GbwvgkeW8_0),.clk(gclk));
	jdff dff_A_8WshvURS4_1(.dout(w_n198_0[1]),.din(w_dff_A_8WshvURS4_1),.clk(gclk));
	jdff dff_A_rImFUdkE8_1(.dout(w_dff_A_8WshvURS4_1),.din(w_dff_A_rImFUdkE8_1),.clk(gclk));
	jdff dff_A_STZojGsg1_1(.dout(w_dff_A_rImFUdkE8_1),.din(w_dff_A_STZojGsg1_1),.clk(gclk));
	jdff dff_A_Ts1tV0HU8_1(.dout(w_dff_A_STZojGsg1_1),.din(w_dff_A_Ts1tV0HU8_1),.clk(gclk));
	jdff dff_A_M8L1bXfV4_2(.dout(w_n198_0[2]),.din(w_dff_A_M8L1bXfV4_2),.clk(gclk));
	jdff dff_A_NFBmxYkG8_2(.dout(w_dff_A_M8L1bXfV4_2),.din(w_dff_A_NFBmxYkG8_2),.clk(gclk));
	jdff dff_A_bgVWcr2A2_2(.dout(w_dff_A_NFBmxYkG8_2),.din(w_dff_A_bgVWcr2A2_2),.clk(gclk));
	jdff dff_A_QWvYTr0x0_2(.dout(w_dff_A_bgVWcr2A2_2),.din(w_dff_A_QWvYTr0x0_2),.clk(gclk));
	jdff dff_A_Rj5xck4f5_1(.dout(w_n135_1[1]),.din(w_dff_A_Rj5xck4f5_1),.clk(gclk));
	jdff dff_A_4r0VLs4A1_1(.dout(w_n117_0[1]),.din(w_dff_A_4r0VLs4A1_1),.clk(gclk));
	jdff dff_A_pFFjlh4U0_1(.dout(w_dff_A_4r0VLs4A1_1),.din(w_dff_A_pFFjlh4U0_1),.clk(gclk));
	jdff dff_A_vkZXroMs3_1(.dout(w_dff_A_pFFjlh4U0_1),.din(w_dff_A_vkZXroMs3_1),.clk(gclk));
	jdff dff_A_7RdF8kzx1_1(.dout(w_dff_A_vkZXroMs3_1),.din(w_dff_A_7RdF8kzx1_1),.clk(gclk));
	jdff dff_A_PwzWTOPB7_2(.dout(w_n117_0[2]),.din(w_dff_A_PwzWTOPB7_2),.clk(gclk));
	jdff dff_A_qIJd2k9C2_2(.dout(w_dff_A_PwzWTOPB7_2),.din(w_dff_A_qIJd2k9C2_2),.clk(gclk));
	jdff dff_A_SKQwpJTr8_2(.dout(w_dff_A_qIJd2k9C2_2),.din(w_dff_A_SKQwpJTr8_2),.clk(gclk));
	jdff dff_A_NJnKpFfd4_2(.dout(w_dff_A_SKQwpJTr8_2),.din(w_dff_A_NJnKpFfd4_2),.clk(gclk));
	jdff dff_A_3gCewhSK3_0(.dout(w_n116_1[0]),.din(w_dff_A_3gCewhSK3_0),.clk(gclk));
	jdff dff_B_FleaHSHC9_1(.din(n239),.dout(w_dff_B_FleaHSHC9_1),.clk(gclk));
	jdff dff_A_LLiTtz3t7_1(.dout(w_n167_0[1]),.din(w_dff_A_LLiTtz3t7_1),.clk(gclk));
	jdff dff_A_38nVQwmt1_0(.dout(w_Gid10_0[0]),.din(w_dff_A_38nVQwmt1_0),.clk(gclk));
	jdff dff_A_rK9ij8KF1_0(.dout(w_dff_A_38nVQwmt1_0),.din(w_dff_A_rK9ij8KF1_0),.clk(gclk));
	jdff dff_A_30hBPQ7Z2_0(.dout(w_dff_A_rK9ij8KF1_0),.din(w_dff_A_30hBPQ7Z2_0),.clk(gclk));
	jdff dff_A_Ubv2Das33_0(.dout(w_dff_A_30hBPQ7Z2_0),.din(w_dff_A_Ubv2Das33_0),.clk(gclk));
	jdff dff_A_ml4J5NVi7_0(.dout(w_dff_A_Ubv2Das33_0),.din(w_dff_A_ml4J5NVi7_0),.clk(gclk));
	jdff dff_A_yi2q2qFV0_0(.dout(w_dff_A_ml4J5NVi7_0),.din(w_dff_A_yi2q2qFV0_0),.clk(gclk));
	jdff dff_A_lUTjZBY86_0(.dout(w_dff_A_yi2q2qFV0_0),.din(w_dff_A_lUTjZBY86_0),.clk(gclk));
	jdff dff_A_6Uhkmc3p8_0(.dout(w_dff_A_lUTjZBY86_0),.din(w_dff_A_6Uhkmc3p8_0),.clk(gclk));
	jdff dff_A_pxZO4WQg6_0(.dout(w_dff_A_6Uhkmc3p8_0),.din(w_dff_A_pxZO4WQg6_0),.clk(gclk));
	jdff dff_A_dFRGcD4F3_0(.dout(w_Gid2_0[0]),.din(w_dff_A_dFRGcD4F3_0),.clk(gclk));
	jdff dff_A_VVtbHkcH3_0(.dout(w_dff_A_dFRGcD4F3_0),.din(w_dff_A_VVtbHkcH3_0),.clk(gclk));
	jdff dff_A_nHGgnyYA9_0(.dout(w_dff_A_VVtbHkcH3_0),.din(w_dff_A_nHGgnyYA9_0),.clk(gclk));
	jdff dff_A_sVXwo5di9_0(.dout(w_dff_A_nHGgnyYA9_0),.din(w_dff_A_sVXwo5di9_0),.clk(gclk));
	jdff dff_A_eQ4y9QWG4_0(.dout(w_dff_A_sVXwo5di9_0),.din(w_dff_A_eQ4y9QWG4_0),.clk(gclk));
	jdff dff_A_XHe0UZA90_0(.dout(w_dff_A_eQ4y9QWG4_0),.din(w_dff_A_XHe0UZA90_0),.clk(gclk));
	jdff dff_A_45Vf5dGX7_0(.dout(w_dff_A_XHe0UZA90_0),.din(w_dff_A_45Vf5dGX7_0),.clk(gclk));
	jdff dff_A_QDDCTmk69_0(.dout(w_dff_A_45Vf5dGX7_0),.din(w_dff_A_QDDCTmk69_0),.clk(gclk));
	jdff dff_A_Knrcr0Ea7_0(.dout(w_dff_A_QDDCTmk69_0),.din(w_dff_A_Knrcr0Ea7_0),.clk(gclk));
	jdff dff_A_lFxY92ZG4_0(.dout(w_dff_A_Knrcr0Ea7_0),.din(w_dff_A_lFxY92ZG4_0),.clk(gclk));
	jdff dff_A_6urkEdQt8_0(.dout(w_n184_0[0]),.din(w_dff_A_6urkEdQt8_0),.clk(gclk));
	jdff dff_A_oL1oe9uq8_0(.dout(w_dff_A_6urkEdQt8_0),.din(w_dff_A_oL1oe9uq8_0),.clk(gclk));
	jdff dff_A_6NQTQiCa1_0(.dout(w_dff_A_oL1oe9uq8_0),.din(w_dff_A_6NQTQiCa1_0),.clk(gclk));
	jdff dff_A_1ikuqBfP1_2(.dout(w_n184_0[2]),.din(w_dff_A_1ikuqBfP1_2),.clk(gclk));
	jdff dff_A_s707V4sK4_2(.dout(w_dff_A_1ikuqBfP1_2),.din(w_dff_A_s707V4sK4_2),.clk(gclk));
	jdff dff_A_OEJiDYKX7_2(.dout(w_dff_A_s707V4sK4_2),.din(w_dff_A_OEJiDYKX7_2),.clk(gclk));
	jdff dff_A_MfDVjbvw0_1(.dout(w_n159_0[1]),.din(w_dff_A_MfDVjbvw0_1),.clk(gclk));
	jdff dff_A_damvTCjB5_0(.dout(w_Gid11_0[0]),.din(w_dff_A_damvTCjB5_0),.clk(gclk));
	jdff dff_A_n3JJdcyq3_0(.dout(w_dff_A_damvTCjB5_0),.din(w_dff_A_n3JJdcyq3_0),.clk(gclk));
	jdff dff_A_ji9KaFGI4_0(.dout(w_dff_A_n3JJdcyq3_0),.din(w_dff_A_ji9KaFGI4_0),.clk(gclk));
	jdff dff_A_9oMO89141_0(.dout(w_dff_A_ji9KaFGI4_0),.din(w_dff_A_9oMO89141_0),.clk(gclk));
	jdff dff_A_tHDn59u91_0(.dout(w_dff_A_9oMO89141_0),.din(w_dff_A_tHDn59u91_0),.clk(gclk));
	jdff dff_A_j0vSDVcx8_0(.dout(w_dff_A_tHDn59u91_0),.din(w_dff_A_j0vSDVcx8_0),.clk(gclk));
	jdff dff_A_LeaqXqFE5_0(.dout(w_dff_A_j0vSDVcx8_0),.din(w_dff_A_LeaqXqFE5_0),.clk(gclk));
	jdff dff_A_6POJdunu5_0(.dout(w_dff_A_LeaqXqFE5_0),.din(w_dff_A_6POJdunu5_0),.clk(gclk));
	jdff dff_A_ygrfhaGE6_0(.dout(w_dff_A_6POJdunu5_0),.din(w_dff_A_ygrfhaGE6_0),.clk(gclk));
	jdff dff_A_PfbGDkXL9_0(.dout(w_Gid3_0[0]),.din(w_dff_A_PfbGDkXL9_0),.clk(gclk));
	jdff dff_A_WeIGzFmv9_0(.dout(w_dff_A_PfbGDkXL9_0),.din(w_dff_A_WeIGzFmv9_0),.clk(gclk));
	jdff dff_A_K5PWTxRS6_0(.dout(w_dff_A_WeIGzFmv9_0),.din(w_dff_A_K5PWTxRS6_0),.clk(gclk));
	jdff dff_A_C5ixUU0g4_0(.dout(w_dff_A_K5PWTxRS6_0),.din(w_dff_A_C5ixUU0g4_0),.clk(gclk));
	jdff dff_A_9uY4yoLn4_0(.dout(w_dff_A_C5ixUU0g4_0),.din(w_dff_A_9uY4yoLn4_0),.clk(gclk));
	jdff dff_A_emgS1Ykw7_0(.dout(w_dff_A_9uY4yoLn4_0),.din(w_dff_A_emgS1Ykw7_0),.clk(gclk));
	jdff dff_A_UfFQBhxF8_0(.dout(w_dff_A_emgS1Ykw7_0),.din(w_dff_A_UfFQBhxF8_0),.clk(gclk));
	jdff dff_A_cPuUE9rM0_0(.dout(w_dff_A_UfFQBhxF8_0),.din(w_dff_A_cPuUE9rM0_0),.clk(gclk));
	jdff dff_A_8ASR3HiH1_0(.dout(w_dff_A_cPuUE9rM0_0),.din(w_dff_A_8ASR3HiH1_0),.clk(gclk));
	jdff dff_A_Ehs49Qsy1_0(.dout(w_dff_A_8ASR3HiH1_0),.din(w_dff_A_Ehs49Qsy1_0),.clk(gclk));
	jdff dff_B_8nYFBoOb8_2(.din(n250),.dout(w_dff_B_8nYFBoOb8_2),.clk(gclk));
	jdff dff_B_97l74v724_2(.din(w_dff_B_8nYFBoOb8_2),.dout(w_dff_B_97l74v724_2),.clk(gclk));
	jdff dff_A_RYxZPFGf4_0(.dout(w_n178_0[0]),.din(w_dff_A_RYxZPFGf4_0),.clk(gclk));
	jdff dff_A_dfjMCcgO4_0(.dout(w_dff_A_RYxZPFGf4_0),.din(w_dff_A_dfjMCcgO4_0),.clk(gclk));
	jdff dff_A_mUG1xxPk9_0(.dout(w_dff_A_dfjMCcgO4_0),.din(w_dff_A_mUG1xxPk9_0),.clk(gclk));
	jdff dff_A_feF2dWmY3_2(.dout(w_n178_0[2]),.din(w_dff_A_feF2dWmY3_2),.clk(gclk));
	jdff dff_A_qe2FC22Z9_2(.dout(w_dff_A_feF2dWmY3_2),.din(w_dff_A_qe2FC22Z9_2),.clk(gclk));
	jdff dff_A_2hdwB6Lq7_2(.dout(w_dff_A_qe2FC22Z9_2),.din(w_dff_A_2hdwB6Lq7_2),.clk(gclk));
	jdff dff_A_ZIJzp40A1_1(.dout(w_n150_0[1]),.din(w_dff_A_ZIJzp40A1_1),.clk(gclk));
	jdff dff_A_jcRibDaM3_0(.dout(w_Gid9_0[0]),.din(w_dff_A_jcRibDaM3_0),.clk(gclk));
	jdff dff_A_sXwhbR2z7_0(.dout(w_dff_A_jcRibDaM3_0),.din(w_dff_A_sXwhbR2z7_0),.clk(gclk));
	jdff dff_A_tEyLqnCC7_0(.dout(w_dff_A_sXwhbR2z7_0),.din(w_dff_A_tEyLqnCC7_0),.clk(gclk));
	jdff dff_A_k8pmRiuA4_0(.dout(w_dff_A_tEyLqnCC7_0),.din(w_dff_A_k8pmRiuA4_0),.clk(gclk));
	jdff dff_A_xzgTCJ4g3_0(.dout(w_dff_A_k8pmRiuA4_0),.din(w_dff_A_xzgTCJ4g3_0),.clk(gclk));
	jdff dff_A_AVxenFrp8_0(.dout(w_dff_A_xzgTCJ4g3_0),.din(w_dff_A_AVxenFrp8_0),.clk(gclk));
	jdff dff_A_iZ18YbbF2_0(.dout(w_dff_A_AVxenFrp8_0),.din(w_dff_A_iZ18YbbF2_0),.clk(gclk));
	jdff dff_A_IHqJUW780_0(.dout(w_dff_A_iZ18YbbF2_0),.din(w_dff_A_IHqJUW780_0),.clk(gclk));
	jdff dff_A_QN1AQoE70_0(.dout(w_dff_A_IHqJUW780_0),.din(w_dff_A_QN1AQoE70_0),.clk(gclk));
	jdff dff_A_nlfCY9eZ4_0(.dout(w_Gid1_0[0]),.din(w_dff_A_nlfCY9eZ4_0),.clk(gclk));
	jdff dff_A_VfVBi8kn2_0(.dout(w_dff_A_nlfCY9eZ4_0),.din(w_dff_A_VfVBi8kn2_0),.clk(gclk));
	jdff dff_A_yjFwUfV27_0(.dout(w_dff_A_VfVBi8kn2_0),.din(w_dff_A_yjFwUfV27_0),.clk(gclk));
	jdff dff_A_h4aYqerg9_0(.dout(w_dff_A_yjFwUfV27_0),.din(w_dff_A_h4aYqerg9_0),.clk(gclk));
	jdff dff_A_zMcu6Y4R6_0(.dout(w_dff_A_h4aYqerg9_0),.din(w_dff_A_zMcu6Y4R6_0),.clk(gclk));
	jdff dff_A_3SAy5bVJ5_0(.dout(w_dff_A_zMcu6Y4R6_0),.din(w_dff_A_3SAy5bVJ5_0),.clk(gclk));
	jdff dff_A_yQumS6Iw9_0(.dout(w_dff_A_3SAy5bVJ5_0),.din(w_dff_A_yQumS6Iw9_0),.clk(gclk));
	jdff dff_A_jh3krFEq8_0(.dout(w_dff_A_yQumS6Iw9_0),.din(w_dff_A_jh3krFEq8_0),.clk(gclk));
	jdff dff_A_t0lijdpE6_0(.dout(w_dff_A_jh3krFEq8_0),.din(w_dff_A_t0lijdpE6_0),.clk(gclk));
	jdff dff_A_juUxwNZX6_0(.dout(w_dff_A_t0lijdpE6_0),.din(w_dff_A_juUxwNZX6_0),.clk(gclk));
	jdff dff_A_FzQHVQVd1_0(.dout(w_Gid26_0[0]),.din(w_dff_A_FzQHVQVd1_0),.clk(gclk));
	jdff dff_A_BLHOFcvB6_0(.dout(w_dff_A_FzQHVQVd1_0),.din(w_dff_A_BLHOFcvB6_0),.clk(gclk));
	jdff dff_A_vpCMzqWU5_0(.dout(w_dff_A_BLHOFcvB6_0),.din(w_dff_A_vpCMzqWU5_0),.clk(gclk));
	jdff dff_A_Y7uubj8a8_0(.dout(w_dff_A_vpCMzqWU5_0),.din(w_dff_A_Y7uubj8a8_0),.clk(gclk));
	jdff dff_A_If2AlXxL1_0(.dout(w_dff_A_Y7uubj8a8_0),.din(w_dff_A_If2AlXxL1_0),.clk(gclk));
	jdff dff_A_gnFqC4Ql6_0(.dout(w_dff_A_If2AlXxL1_0),.din(w_dff_A_gnFqC4Ql6_0),.clk(gclk));
	jdff dff_A_Cji16JFo9_0(.dout(w_dff_A_gnFqC4Ql6_0),.din(w_dff_A_Cji16JFo9_0),.clk(gclk));
	jdff dff_A_WKU0TH3V0_0(.dout(w_dff_A_Cji16JFo9_0),.din(w_dff_A_WKU0TH3V0_0),.clk(gclk));
	jdff dff_A_Uxnxvwc57_0(.dout(w_dff_A_WKU0TH3V0_0),.din(w_dff_A_Uxnxvwc57_0),.clk(gclk));
	jdff dff_A_hNLQDEle0_0(.dout(w_dff_A_Uxnxvwc57_0),.din(w_dff_A_hNLQDEle0_0),.clk(gclk));
	jdff dff_A_xSBXQeTL8_0(.dout(w_Gid25_0[0]),.din(w_dff_A_xSBXQeTL8_0),.clk(gclk));
	jdff dff_A_ULrjhnzx1_0(.dout(w_dff_A_xSBXQeTL8_0),.din(w_dff_A_ULrjhnzx1_0),.clk(gclk));
	jdff dff_A_gZD9nxQC3_0(.dout(w_dff_A_ULrjhnzx1_0),.din(w_dff_A_gZD9nxQC3_0),.clk(gclk));
	jdff dff_A_HVbIHqyp8_0(.dout(w_dff_A_gZD9nxQC3_0),.din(w_dff_A_HVbIHqyp8_0),.clk(gclk));
	jdff dff_A_oCsZXx1N0_0(.dout(w_dff_A_HVbIHqyp8_0),.din(w_dff_A_oCsZXx1N0_0),.clk(gclk));
	jdff dff_A_NU4DqDz64_0(.dout(w_dff_A_oCsZXx1N0_0),.din(w_dff_A_NU4DqDz64_0),.clk(gclk));
	jdff dff_A_RcUmVaze5_0(.dout(w_dff_A_NU4DqDz64_0),.din(w_dff_A_RcUmVaze5_0),.clk(gclk));
	jdff dff_A_gy9DVSgM8_0(.dout(w_dff_A_RcUmVaze5_0),.din(w_dff_A_gy9DVSgM8_0),.clk(gclk));
	jdff dff_A_Tl3Ue38z6_0(.dout(w_dff_A_gy9DVSgM8_0),.din(w_dff_A_Tl3Ue38z6_0),.clk(gclk));
	jdff dff_A_lwZhi6iY6_0(.dout(w_dff_A_Tl3Ue38z6_0),.din(w_dff_A_lwZhi6iY6_0),.clk(gclk));
	jdff dff_A_Br7A30gp1_0(.dout(w_Gid24_0[0]),.din(w_dff_A_Br7A30gp1_0),.clk(gclk));
	jdff dff_A_EZBUjOOC7_0(.dout(w_dff_A_Br7A30gp1_0),.din(w_dff_A_EZBUjOOC7_0),.clk(gclk));
	jdff dff_A_o7StwBmy3_0(.dout(w_dff_A_EZBUjOOC7_0),.din(w_dff_A_o7StwBmy3_0),.clk(gclk));
	jdff dff_A_3UWQ7sKS4_0(.dout(w_dff_A_o7StwBmy3_0),.din(w_dff_A_3UWQ7sKS4_0),.clk(gclk));
	jdff dff_A_TLbHxl1l5_0(.dout(w_dff_A_3UWQ7sKS4_0),.din(w_dff_A_TLbHxl1l5_0),.clk(gclk));
	jdff dff_A_BByKlYj37_0(.dout(w_dff_A_TLbHxl1l5_0),.din(w_dff_A_BByKlYj37_0),.clk(gclk));
	jdff dff_A_4DsW3pay3_0(.dout(w_dff_A_BByKlYj37_0),.din(w_dff_A_4DsW3pay3_0),.clk(gclk));
	jdff dff_A_VOtCwJvH5_0(.dout(w_dff_A_4DsW3pay3_0),.din(w_dff_A_VOtCwJvH5_0),.clk(gclk));
	jdff dff_A_gBstYV6h6_0(.dout(w_dff_A_VOtCwJvH5_0),.din(w_dff_A_gBstYV6h6_0),.clk(gclk));
	jdff dff_A_E22RhgI36_0(.dout(w_dff_A_gBstYV6h6_0),.din(w_dff_A_E22RhgI36_0),.clk(gclk));
	jdff dff_A_iSDbBGr43_0(.dout(w_Gid30_0[0]),.din(w_dff_A_iSDbBGr43_0),.clk(gclk));
	jdff dff_A_aL55yYLe9_0(.dout(w_dff_A_iSDbBGr43_0),.din(w_dff_A_aL55yYLe9_0),.clk(gclk));
	jdff dff_A_1Wz5YjX11_0(.dout(w_dff_A_aL55yYLe9_0),.din(w_dff_A_1Wz5YjX11_0),.clk(gclk));
	jdff dff_A_C3gVbDDy7_0(.dout(w_dff_A_1Wz5YjX11_0),.din(w_dff_A_C3gVbDDy7_0),.clk(gclk));
	jdff dff_A_bB8KWaiS7_0(.dout(w_dff_A_C3gVbDDy7_0),.din(w_dff_A_bB8KWaiS7_0),.clk(gclk));
	jdff dff_A_fqKjbUVE3_0(.dout(w_dff_A_bB8KWaiS7_0),.din(w_dff_A_fqKjbUVE3_0),.clk(gclk));
	jdff dff_A_7txFciWh6_0(.dout(w_dff_A_fqKjbUVE3_0),.din(w_dff_A_7txFciWh6_0),.clk(gclk));
	jdff dff_A_HzozIe276_0(.dout(w_dff_A_7txFciWh6_0),.din(w_dff_A_HzozIe276_0),.clk(gclk));
	jdff dff_A_t2tzlX5U5_0(.dout(w_dff_A_HzozIe276_0),.din(w_dff_A_t2tzlX5U5_0),.clk(gclk));
	jdff dff_A_3GoHoAV63_0(.dout(w_dff_A_t2tzlX5U5_0),.din(w_dff_A_3GoHoAV63_0),.clk(gclk));
	jdff dff_A_iII172id8_0(.dout(w_Gid29_0[0]),.din(w_dff_A_iII172id8_0),.clk(gclk));
	jdff dff_A_qiLWyHXx3_0(.dout(w_dff_A_iII172id8_0),.din(w_dff_A_qiLWyHXx3_0),.clk(gclk));
	jdff dff_A_FFNvq2nn4_0(.dout(w_dff_A_qiLWyHXx3_0),.din(w_dff_A_FFNvq2nn4_0),.clk(gclk));
	jdff dff_A_HhFUejdw5_0(.dout(w_dff_A_FFNvq2nn4_0),.din(w_dff_A_HhFUejdw5_0),.clk(gclk));
	jdff dff_A_Nl3czyl52_0(.dout(w_dff_A_HhFUejdw5_0),.din(w_dff_A_Nl3czyl52_0),.clk(gclk));
	jdff dff_A_bxdbeUFt4_0(.dout(w_dff_A_Nl3czyl52_0),.din(w_dff_A_bxdbeUFt4_0),.clk(gclk));
	jdff dff_A_3EnfGnyW3_0(.dout(w_dff_A_bxdbeUFt4_0),.din(w_dff_A_3EnfGnyW3_0),.clk(gclk));
	jdff dff_A_uroHc92O6_0(.dout(w_dff_A_3EnfGnyW3_0),.din(w_dff_A_uroHc92O6_0),.clk(gclk));
	jdff dff_A_pxjUCRIP6_0(.dout(w_dff_A_uroHc92O6_0),.din(w_dff_A_pxjUCRIP6_0),.clk(gclk));
	jdff dff_A_ZXZxQSbT4_0(.dout(w_dff_A_pxjUCRIP6_0),.din(w_dff_A_ZXZxQSbT4_0),.clk(gclk));
	jdff dff_A_q7ENROth4_0(.dout(w_Gid28_0[0]),.din(w_dff_A_q7ENROth4_0),.clk(gclk));
	jdff dff_A_oqCosAcc4_0(.dout(w_dff_A_q7ENROth4_0),.din(w_dff_A_oqCosAcc4_0),.clk(gclk));
	jdff dff_A_fS4jQyCt4_0(.dout(w_dff_A_oqCosAcc4_0),.din(w_dff_A_fS4jQyCt4_0),.clk(gclk));
	jdff dff_A_FyGHhDte8_0(.dout(w_dff_A_fS4jQyCt4_0),.din(w_dff_A_FyGHhDte8_0),.clk(gclk));
	jdff dff_A_FVWW2Ufc7_0(.dout(w_dff_A_FyGHhDte8_0),.din(w_dff_A_FVWW2Ufc7_0),.clk(gclk));
	jdff dff_A_WB9YVhx87_0(.dout(w_dff_A_FVWW2Ufc7_0),.din(w_dff_A_WB9YVhx87_0),.clk(gclk));
	jdff dff_A_IFQ5cYYB5_0(.dout(w_dff_A_WB9YVhx87_0),.din(w_dff_A_IFQ5cYYB5_0),.clk(gclk));
	jdff dff_A_1WRkxZYv3_0(.dout(w_dff_A_IFQ5cYYB5_0),.din(w_dff_A_1WRkxZYv3_0),.clk(gclk));
	jdff dff_A_EhMyHGaN7_0(.dout(w_dff_A_1WRkxZYv3_0),.din(w_dff_A_EhMyHGaN7_0),.clk(gclk));
	jdff dff_A_JaGskUwi2_0(.dout(w_dff_A_EhMyHGaN7_0),.din(w_dff_A_JaGskUwi2_0),.clk(gclk));
	jdff dff_A_JHfHeD4W6_1(.dout(w_n87_0[1]),.din(w_dff_A_JHfHeD4W6_1),.clk(gclk));
	jdff dff_A_e0f20Of68_0(.dout(w_Gid22_0[0]),.din(w_dff_A_e0f20Of68_0),.clk(gclk));
	jdff dff_A_csABP28l4_0(.dout(w_dff_A_e0f20Of68_0),.din(w_dff_A_csABP28l4_0),.clk(gclk));
	jdff dff_A_zzxR9Ii12_0(.dout(w_dff_A_csABP28l4_0),.din(w_dff_A_zzxR9Ii12_0),.clk(gclk));
	jdff dff_A_aEngsCQg0_0(.dout(w_dff_A_zzxR9Ii12_0),.din(w_dff_A_aEngsCQg0_0),.clk(gclk));
	jdff dff_A_3dAHsyre7_0(.dout(w_dff_A_aEngsCQg0_0),.din(w_dff_A_3dAHsyre7_0),.clk(gclk));
	jdff dff_A_1kR1fyGQ3_0(.dout(w_dff_A_3dAHsyre7_0),.din(w_dff_A_1kR1fyGQ3_0),.clk(gclk));
	jdff dff_A_2ZM9I5Sk7_0(.dout(w_dff_A_1kR1fyGQ3_0),.din(w_dff_A_2ZM9I5Sk7_0),.clk(gclk));
	jdff dff_A_I2MMOWyw3_0(.dout(w_dff_A_2ZM9I5Sk7_0),.din(w_dff_A_I2MMOWyw3_0),.clk(gclk));
	jdff dff_A_TSyhpsdb2_0(.dout(w_dff_A_I2MMOWyw3_0),.din(w_dff_A_TSyhpsdb2_0),.clk(gclk));
	jdff dff_A_v52rLRPg7_0(.dout(w_dff_A_TSyhpsdb2_0),.din(w_dff_A_v52rLRPg7_0),.clk(gclk));
	jdff dff_A_d9cdBOFM4_0(.dout(w_Gid21_0[0]),.din(w_dff_A_d9cdBOFM4_0),.clk(gclk));
	jdff dff_A_HLcoKE646_0(.dout(w_dff_A_d9cdBOFM4_0),.din(w_dff_A_HLcoKE646_0),.clk(gclk));
	jdff dff_A_4fL9euP86_0(.dout(w_dff_A_HLcoKE646_0),.din(w_dff_A_4fL9euP86_0),.clk(gclk));
	jdff dff_A_izpaHMpn7_0(.dout(w_dff_A_4fL9euP86_0),.din(w_dff_A_izpaHMpn7_0),.clk(gclk));
	jdff dff_A_wqL0WCtR1_0(.dout(w_dff_A_izpaHMpn7_0),.din(w_dff_A_wqL0WCtR1_0),.clk(gclk));
	jdff dff_A_uFK8DEfL4_0(.dout(w_dff_A_wqL0WCtR1_0),.din(w_dff_A_uFK8DEfL4_0),.clk(gclk));
	jdff dff_A_ANU9vpyT4_0(.dout(w_dff_A_uFK8DEfL4_0),.din(w_dff_A_ANU9vpyT4_0),.clk(gclk));
	jdff dff_A_wutTKT5o0_0(.dout(w_dff_A_ANU9vpyT4_0),.din(w_dff_A_wutTKT5o0_0),.clk(gclk));
	jdff dff_A_yREcq8vF1_0(.dout(w_dff_A_wutTKT5o0_0),.din(w_dff_A_yREcq8vF1_0),.clk(gclk));
	jdff dff_A_y3d5rboI7_0(.dout(w_dff_A_yREcq8vF1_0),.din(w_dff_A_y3d5rboI7_0),.clk(gclk));
	jdff dff_A_SyMPwkUR6_0(.dout(w_Gid20_0[0]),.din(w_dff_A_SyMPwkUR6_0),.clk(gclk));
	jdff dff_A_0uB8qeBw8_0(.dout(w_dff_A_SyMPwkUR6_0),.din(w_dff_A_0uB8qeBw8_0),.clk(gclk));
	jdff dff_A_R0ccmP144_0(.dout(w_dff_A_0uB8qeBw8_0),.din(w_dff_A_R0ccmP144_0),.clk(gclk));
	jdff dff_A_eXfOj34b5_0(.dout(w_dff_A_R0ccmP144_0),.din(w_dff_A_eXfOj34b5_0),.clk(gclk));
	jdff dff_A_iIYXS9XK7_0(.dout(w_dff_A_eXfOj34b5_0),.din(w_dff_A_iIYXS9XK7_0),.clk(gclk));
	jdff dff_A_tjPp8cGe8_0(.dout(w_dff_A_iIYXS9XK7_0),.din(w_dff_A_tjPp8cGe8_0),.clk(gclk));
	jdff dff_A_6Snlr1V52_0(.dout(w_dff_A_tjPp8cGe8_0),.din(w_dff_A_6Snlr1V52_0),.clk(gclk));
	jdff dff_A_D2Vol7Oi9_0(.dout(w_dff_A_6Snlr1V52_0),.din(w_dff_A_D2Vol7Oi9_0),.clk(gclk));
	jdff dff_A_PcBKuAi53_0(.dout(w_dff_A_D2Vol7Oi9_0),.din(w_dff_A_PcBKuAi53_0),.clk(gclk));
	jdff dff_A_I7zSl4Oo8_0(.dout(w_dff_A_PcBKuAi53_0),.din(w_dff_A_I7zSl4Oo8_0),.clk(gclk));
	jdff dff_A_1Mta0FRo5_0(.dout(w_Gid8_0[0]),.din(w_dff_A_1Mta0FRo5_0),.clk(gclk));
	jdff dff_A_oBehxNMy4_0(.dout(w_dff_A_1Mta0FRo5_0),.din(w_dff_A_oBehxNMy4_0),.clk(gclk));
	jdff dff_A_0hClBwca0_0(.dout(w_dff_A_oBehxNMy4_0),.din(w_dff_A_0hClBwca0_0),.clk(gclk));
	jdff dff_A_4eS53urV3_0(.dout(w_dff_A_0hClBwca0_0),.din(w_dff_A_4eS53urV3_0),.clk(gclk));
	jdff dff_A_MqWWxRTY9_0(.dout(w_dff_A_4eS53urV3_0),.din(w_dff_A_MqWWxRTY9_0),.clk(gclk));
	jdff dff_A_Et9KTzRE0_0(.dout(w_dff_A_MqWWxRTY9_0),.din(w_dff_A_Et9KTzRE0_0),.clk(gclk));
	jdff dff_A_nHlYQRJx5_0(.dout(w_dff_A_Et9KTzRE0_0),.din(w_dff_A_nHlYQRJx5_0),.clk(gclk));
	jdff dff_A_Eec6HTvf2_0(.dout(w_dff_A_nHlYQRJx5_0),.din(w_dff_A_Eec6HTvf2_0),.clk(gclk));
	jdff dff_A_QXExpRAt1_0(.dout(w_dff_A_Eec6HTvf2_0),.din(w_dff_A_QXExpRAt1_0),.clk(gclk));
	jdff dff_A_xFw1BOWp5_0(.dout(w_Gid0_0[0]),.din(w_dff_A_xFw1BOWp5_0),.clk(gclk));
	jdff dff_A_xciZE5IX8_0(.dout(w_dff_A_xFw1BOWp5_0),.din(w_dff_A_xciZE5IX8_0),.clk(gclk));
	jdff dff_A_aQfHNGca7_0(.dout(w_dff_A_xciZE5IX8_0),.din(w_dff_A_aQfHNGca7_0),.clk(gclk));
	jdff dff_A_Ye6CAmvR5_0(.dout(w_dff_A_aQfHNGca7_0),.din(w_dff_A_Ye6CAmvR5_0),.clk(gclk));
	jdff dff_A_SMiNFZbi2_0(.dout(w_dff_A_Ye6CAmvR5_0),.din(w_dff_A_SMiNFZbi2_0),.clk(gclk));
	jdff dff_A_bWdPzZaC7_0(.dout(w_dff_A_SMiNFZbi2_0),.din(w_dff_A_bWdPzZaC7_0),.clk(gclk));
	jdff dff_A_PLoh3owQ5_0(.dout(w_dff_A_bWdPzZaC7_0),.din(w_dff_A_PLoh3owQ5_0),.clk(gclk));
	jdff dff_A_1FPAdSGH2_0(.dout(w_dff_A_PLoh3owQ5_0),.din(w_dff_A_1FPAdSGH2_0),.clk(gclk));
	jdff dff_A_zXvLuIgT6_0(.dout(w_dff_A_1FPAdSGH2_0),.din(w_dff_A_zXvLuIgT6_0),.clk(gclk));
	jdff dff_A_YsUNoZov4_0(.dout(w_dff_A_zXvLuIgT6_0),.din(w_dff_A_YsUNoZov4_0),.clk(gclk));
	jdff dff_A_Ff6PPWup0_0(.dout(w_Gid18_0[0]),.din(w_dff_A_Ff6PPWup0_0),.clk(gclk));
	jdff dff_A_513AJPwb8_0(.dout(w_dff_A_Ff6PPWup0_0),.din(w_dff_A_513AJPwb8_0),.clk(gclk));
	jdff dff_A_4sptdXIf1_0(.dout(w_dff_A_513AJPwb8_0),.din(w_dff_A_4sptdXIf1_0),.clk(gclk));
	jdff dff_A_DuJIQdFk5_0(.dout(w_dff_A_4sptdXIf1_0),.din(w_dff_A_DuJIQdFk5_0),.clk(gclk));
	jdff dff_A_Obufz23g4_0(.dout(w_dff_A_DuJIQdFk5_0),.din(w_dff_A_Obufz23g4_0),.clk(gclk));
	jdff dff_A_pgk63Lcf8_0(.dout(w_dff_A_Obufz23g4_0),.din(w_dff_A_pgk63Lcf8_0),.clk(gclk));
	jdff dff_A_NGkQye6u3_0(.dout(w_dff_A_pgk63Lcf8_0),.din(w_dff_A_NGkQye6u3_0),.clk(gclk));
	jdff dff_A_iKJVKK5Q9_0(.dout(w_dff_A_NGkQye6u3_0),.din(w_dff_A_iKJVKK5Q9_0),.clk(gclk));
	jdff dff_A_Y9aZM7VE5_0(.dout(w_dff_A_iKJVKK5Q9_0),.din(w_dff_A_Y9aZM7VE5_0),.clk(gclk));
	jdff dff_A_PaXUWnuJ3_0(.dout(w_dff_A_Y9aZM7VE5_0),.din(w_dff_A_PaXUWnuJ3_0),.clk(gclk));
	jdff dff_A_AfRlojZO8_0(.dout(w_Gid17_0[0]),.din(w_dff_A_AfRlojZO8_0),.clk(gclk));
	jdff dff_A_tMbb5eAY2_0(.dout(w_dff_A_AfRlojZO8_0),.din(w_dff_A_tMbb5eAY2_0),.clk(gclk));
	jdff dff_A_PkBcyinB3_0(.dout(w_dff_A_tMbb5eAY2_0),.din(w_dff_A_PkBcyinB3_0),.clk(gclk));
	jdff dff_A_ulc6f5Hj8_0(.dout(w_dff_A_PkBcyinB3_0),.din(w_dff_A_ulc6f5Hj8_0),.clk(gclk));
	jdff dff_A_7W1mUFqy7_0(.dout(w_dff_A_ulc6f5Hj8_0),.din(w_dff_A_7W1mUFqy7_0),.clk(gclk));
	jdff dff_A_WT7ho4U09_0(.dout(w_dff_A_7W1mUFqy7_0),.din(w_dff_A_WT7ho4U09_0),.clk(gclk));
	jdff dff_A_1WgJfbkc2_0(.dout(w_dff_A_WT7ho4U09_0),.din(w_dff_A_1WgJfbkc2_0),.clk(gclk));
	jdff dff_A_LeV0kfew9_0(.dout(w_dff_A_1WgJfbkc2_0),.din(w_dff_A_LeV0kfew9_0),.clk(gclk));
	jdff dff_A_Z1lRabTN9_0(.dout(w_dff_A_LeV0kfew9_0),.din(w_dff_A_Z1lRabTN9_0),.clk(gclk));
	jdff dff_A_OVz3kojF3_0(.dout(w_dff_A_Z1lRabTN9_0),.din(w_dff_A_OVz3kojF3_0),.clk(gclk));
	jdff dff_A_Z8nhfsjM3_0(.dout(w_Gid16_0[0]),.din(w_dff_A_Z8nhfsjM3_0),.clk(gclk));
	jdff dff_A_J9i1HOod0_0(.dout(w_dff_A_Z8nhfsjM3_0),.din(w_dff_A_J9i1HOod0_0),.clk(gclk));
	jdff dff_A_YsORmye48_0(.dout(w_dff_A_J9i1HOod0_0),.din(w_dff_A_YsORmye48_0),.clk(gclk));
	jdff dff_A_041Jrkqp4_0(.dout(w_dff_A_YsORmye48_0),.din(w_dff_A_041Jrkqp4_0),.clk(gclk));
	jdff dff_A_YtNhgngi9_0(.dout(w_dff_A_041Jrkqp4_0),.din(w_dff_A_YtNhgngi9_0),.clk(gclk));
	jdff dff_A_nr9wxVt56_0(.dout(w_dff_A_YtNhgngi9_0),.din(w_dff_A_nr9wxVt56_0),.clk(gclk));
	jdff dff_A_Zcncu5pV7_0(.dout(w_dff_A_nr9wxVt56_0),.din(w_dff_A_Zcncu5pV7_0),.clk(gclk));
	jdff dff_A_2Z72Bbfy8_0(.dout(w_dff_A_Zcncu5pV7_0),.din(w_dff_A_2Z72Bbfy8_0),.clk(gclk));
	jdff dff_A_ACqLObVw9_0(.dout(w_dff_A_2Z72Bbfy8_0),.din(w_dff_A_ACqLObVw9_0),.clk(gclk));
	jdff dff_A_XmRrv8nG7_0(.dout(w_dff_A_ACqLObVw9_0),.din(w_dff_A_XmRrv8nG7_0),.clk(gclk));
	jdff dff_A_b7eWEwPm2_1(.dout(w_n187_0[1]),.din(w_dff_A_b7eWEwPm2_1),.clk(gclk));
	jdff dff_A_1pXnnjqi2_1(.dout(w_dff_A_b7eWEwPm2_1),.din(w_dff_A_1pXnnjqi2_1),.clk(gclk));
	jdff dff_A_F9sOOZqT0_1(.dout(w_dff_A_1pXnnjqi2_1),.din(w_dff_A_F9sOOZqT0_1),.clk(gclk));
	jdff dff_A_uBkBXEWl3_1(.dout(w_dff_A_F9sOOZqT0_1),.din(w_dff_A_uBkBXEWl3_1),.clk(gclk));
	jdff dff_A_N2Wba22G6_2(.dout(w_n187_0[2]),.din(w_dff_A_N2Wba22G6_2),.clk(gclk));
	jdff dff_A_vOnKQtMl7_2(.dout(w_dff_A_N2Wba22G6_2),.din(w_dff_A_vOnKQtMl7_2),.clk(gclk));
	jdff dff_A_OhFFmIKc1_2(.dout(w_dff_A_vOnKQtMl7_2),.din(w_dff_A_OhFFmIKc1_2),.clk(gclk));
	jdff dff_A_H1KiPvTH0_2(.dout(w_dff_A_OhFFmIKc1_2),.din(w_dff_A_H1KiPvTH0_2),.clk(gclk));
	jdff dff_A_HEyAYzEs7_1(.dout(w_n102_1[1]),.din(w_dff_A_HEyAYzEs7_1),.clk(gclk));
	jdff dff_A_QwzLAtAx0_0(.dout(w_Gid31_0[0]),.din(w_dff_A_QwzLAtAx0_0),.clk(gclk));
	jdff dff_A_kL8Q0MNb7_0(.dout(w_dff_A_QwzLAtAx0_0),.din(w_dff_A_kL8Q0MNb7_0),.clk(gclk));
	jdff dff_A_pFlmQUJv2_0(.dout(w_dff_A_kL8Q0MNb7_0),.din(w_dff_A_pFlmQUJv2_0),.clk(gclk));
	jdff dff_A_66XdLzSi4_0(.dout(w_dff_A_pFlmQUJv2_0),.din(w_dff_A_66XdLzSi4_0),.clk(gclk));
	jdff dff_A_1DBHxGAI1_0(.dout(w_dff_A_66XdLzSi4_0),.din(w_dff_A_1DBHxGAI1_0),.clk(gclk));
	jdff dff_A_2SweqIOi6_0(.dout(w_dff_A_1DBHxGAI1_0),.din(w_dff_A_2SweqIOi6_0),.clk(gclk));
	jdff dff_A_bFXseTRd8_0(.dout(w_dff_A_2SweqIOi6_0),.din(w_dff_A_bFXseTRd8_0),.clk(gclk));
	jdff dff_A_rQr6v7Hq8_0(.dout(w_dff_A_bFXseTRd8_0),.din(w_dff_A_rQr6v7Hq8_0),.clk(gclk));
	jdff dff_A_xNU8rjDp3_0(.dout(w_dff_A_rQr6v7Hq8_0),.din(w_dff_A_xNU8rjDp3_0),.clk(gclk));
	jdff dff_A_wLmNjqFi8_0(.dout(w_dff_A_xNU8rjDp3_0),.din(w_dff_A_wLmNjqFi8_0),.clk(gclk));
	jdff dff_A_V9575tAZ8_0(.dout(w_Gid27_0[0]),.din(w_dff_A_V9575tAZ8_0),.clk(gclk));
	jdff dff_A_yZI0PRA86_0(.dout(w_dff_A_V9575tAZ8_0),.din(w_dff_A_yZI0PRA86_0),.clk(gclk));
	jdff dff_A_yaYnJmvC0_0(.dout(w_dff_A_yZI0PRA86_0),.din(w_dff_A_yaYnJmvC0_0),.clk(gclk));
	jdff dff_A_jPDojBgh2_0(.dout(w_dff_A_yaYnJmvC0_0),.din(w_dff_A_jPDojBgh2_0),.clk(gclk));
	jdff dff_A_9zRgDp2a0_0(.dout(w_dff_A_jPDojBgh2_0),.din(w_dff_A_9zRgDp2a0_0),.clk(gclk));
	jdff dff_A_Q8EqOzhI7_0(.dout(w_dff_A_9zRgDp2a0_0),.din(w_dff_A_Q8EqOzhI7_0),.clk(gclk));
	jdff dff_A_HYtNnSkz9_0(.dout(w_dff_A_Q8EqOzhI7_0),.din(w_dff_A_HYtNnSkz9_0),.clk(gclk));
	jdff dff_A_hxa6lDUx0_0(.dout(w_dff_A_HYtNnSkz9_0),.din(w_dff_A_hxa6lDUx0_0),.clk(gclk));
	jdff dff_A_x8XdVgs38_0(.dout(w_dff_A_hxa6lDUx0_0),.din(w_dff_A_x8XdVgs38_0),.clk(gclk));
	jdff dff_A_MO03c5xV3_0(.dout(w_dff_A_x8XdVgs38_0),.din(w_dff_A_MO03c5xV3_0),.clk(gclk));
	jdff dff_A_iELAqCDW6_0(.dout(w_Gid23_0[0]),.din(w_dff_A_iELAqCDW6_0),.clk(gclk));
	jdff dff_A_b2gsjM1n4_0(.dout(w_dff_A_iELAqCDW6_0),.din(w_dff_A_b2gsjM1n4_0),.clk(gclk));
	jdff dff_A_G1z5U4Ui5_0(.dout(w_dff_A_b2gsjM1n4_0),.din(w_dff_A_G1z5U4Ui5_0),.clk(gclk));
	jdff dff_A_0wYk2Vb47_0(.dout(w_dff_A_G1z5U4Ui5_0),.din(w_dff_A_0wYk2Vb47_0),.clk(gclk));
	jdff dff_A_EuBlqX472_0(.dout(w_dff_A_0wYk2Vb47_0),.din(w_dff_A_EuBlqX472_0),.clk(gclk));
	jdff dff_A_QAcPOklx8_0(.dout(w_dff_A_EuBlqX472_0),.din(w_dff_A_QAcPOklx8_0),.clk(gclk));
	jdff dff_A_rwaFJ7H30_0(.dout(w_dff_A_QAcPOklx8_0),.din(w_dff_A_rwaFJ7H30_0),.clk(gclk));
	jdff dff_A_tujslkKe0_0(.dout(w_dff_A_rwaFJ7H30_0),.din(w_dff_A_tujslkKe0_0),.clk(gclk));
	jdff dff_A_GBOUtBRn5_0(.dout(w_dff_A_tujslkKe0_0),.din(w_dff_A_GBOUtBRn5_0),.clk(gclk));
	jdff dff_A_bQX9gF2S9_0(.dout(w_dff_A_GBOUtBRn5_0),.din(w_dff_A_bQX9gF2S9_0),.clk(gclk));
	jdff dff_A_Xqmn3PZp8_0(.dout(w_Gid19_0[0]),.din(w_dff_A_Xqmn3PZp8_0),.clk(gclk));
	jdff dff_A_PanEnjlZ5_0(.dout(w_dff_A_Xqmn3PZp8_0),.din(w_dff_A_PanEnjlZ5_0),.clk(gclk));
	jdff dff_A_R80Rcvg22_0(.dout(w_dff_A_PanEnjlZ5_0),.din(w_dff_A_R80Rcvg22_0),.clk(gclk));
	jdff dff_A_01dvP1cg0_0(.dout(w_dff_A_R80Rcvg22_0),.din(w_dff_A_01dvP1cg0_0),.clk(gclk));
	jdff dff_A_FAfElg7H6_0(.dout(w_dff_A_01dvP1cg0_0),.din(w_dff_A_FAfElg7H6_0),.clk(gclk));
	jdff dff_A_NU3ew8Bb0_0(.dout(w_dff_A_FAfElg7H6_0),.din(w_dff_A_NU3ew8Bb0_0),.clk(gclk));
	jdff dff_A_mWhAP6Fw3_0(.dout(w_dff_A_NU3ew8Bb0_0),.din(w_dff_A_mWhAP6Fw3_0),.clk(gclk));
	jdff dff_A_3c0OhL8m9_0(.dout(w_dff_A_mWhAP6Fw3_0),.din(w_dff_A_3c0OhL8m9_0),.clk(gclk));
	jdff dff_A_WCBBAKzQ6_0(.dout(w_dff_A_3c0OhL8m9_0),.din(w_dff_A_WCBBAKzQ6_0),.clk(gclk));
	jdff dff_A_LEJdWwnh0_0(.dout(w_dff_A_WCBBAKzQ6_0),.din(w_dff_A_LEJdWwnh0_0),.clk(gclk));
	jdff dff_A_RR0yQgGz8_0(.dout(w_Gid15_0[0]),.din(w_dff_A_RR0yQgGz8_0),.clk(gclk));
	jdff dff_A_GNO3S7JI7_0(.dout(w_dff_A_RR0yQgGz8_0),.din(w_dff_A_GNO3S7JI7_0),.clk(gclk));
	jdff dff_A_Qp3b8qrn2_0(.dout(w_dff_A_GNO3S7JI7_0),.din(w_dff_A_Qp3b8qrn2_0),.clk(gclk));
	jdff dff_A_W7m6Syd27_0(.dout(w_dff_A_Qp3b8qrn2_0),.din(w_dff_A_W7m6Syd27_0),.clk(gclk));
	jdff dff_A_LVNs9DC23_0(.dout(w_dff_A_W7m6Syd27_0),.din(w_dff_A_LVNs9DC23_0),.clk(gclk));
	jdff dff_A_QLbsGLBj8_0(.dout(w_dff_A_LVNs9DC23_0),.din(w_dff_A_QLbsGLBj8_0),.clk(gclk));
	jdff dff_A_0GMcFs7C9_0(.dout(w_dff_A_QLbsGLBj8_0),.din(w_dff_A_0GMcFs7C9_0),.clk(gclk));
	jdff dff_A_7S7rZln52_0(.dout(w_dff_A_0GMcFs7C9_0),.din(w_dff_A_7S7rZln52_0),.clk(gclk));
	jdff dff_A_n9T6JgZ27_0(.dout(w_dff_A_7S7rZln52_0),.din(w_dff_A_n9T6JgZ27_0),.clk(gclk));
	jdff dff_A_9FSP0flA0_0(.dout(w_Gid14_0[0]),.din(w_dff_A_9FSP0flA0_0),.clk(gclk));
	jdff dff_A_9dUWoDcq5_0(.dout(w_dff_A_9FSP0flA0_0),.din(w_dff_A_9dUWoDcq5_0),.clk(gclk));
	jdff dff_A_E6m84ZSg5_0(.dout(w_dff_A_9dUWoDcq5_0),.din(w_dff_A_E6m84ZSg5_0),.clk(gclk));
	jdff dff_A_UfpAOE2k9_0(.dout(w_dff_A_E6m84ZSg5_0),.din(w_dff_A_UfpAOE2k9_0),.clk(gclk));
	jdff dff_A_3XWJwo7R6_0(.dout(w_dff_A_UfpAOE2k9_0),.din(w_dff_A_3XWJwo7R6_0),.clk(gclk));
	jdff dff_A_hG1tkdaa0_0(.dout(w_dff_A_3XWJwo7R6_0),.din(w_dff_A_hG1tkdaa0_0),.clk(gclk));
	jdff dff_A_VeBN4WF29_0(.dout(w_dff_A_hG1tkdaa0_0),.din(w_dff_A_VeBN4WF29_0),.clk(gclk));
	jdff dff_A_2EylyEZ32_0(.dout(w_dff_A_VeBN4WF29_0),.din(w_dff_A_2EylyEZ32_0),.clk(gclk));
	jdff dff_A_aOH4rWq78_0(.dout(w_dff_A_2EylyEZ32_0),.din(w_dff_A_aOH4rWq78_0),.clk(gclk));
	jdff dff_A_ww2WoK2p2_0(.dout(w_Gid13_0[0]),.din(w_dff_A_ww2WoK2p2_0),.clk(gclk));
	jdff dff_A_OVoP1XFp3_0(.dout(w_dff_A_ww2WoK2p2_0),.din(w_dff_A_OVoP1XFp3_0),.clk(gclk));
	jdff dff_A_gq5vEoM78_0(.dout(w_dff_A_OVoP1XFp3_0),.din(w_dff_A_gq5vEoM78_0),.clk(gclk));
	jdff dff_A_KJ5ptrdO7_0(.dout(w_dff_A_gq5vEoM78_0),.din(w_dff_A_KJ5ptrdO7_0),.clk(gclk));
	jdff dff_A_FoYtcmCu0_0(.dout(w_dff_A_KJ5ptrdO7_0),.din(w_dff_A_FoYtcmCu0_0),.clk(gclk));
	jdff dff_A_aBT8h6OV8_0(.dout(w_dff_A_FoYtcmCu0_0),.din(w_dff_A_aBT8h6OV8_0),.clk(gclk));
	jdff dff_A_rKYBJCle1_0(.dout(w_dff_A_aBT8h6OV8_0),.din(w_dff_A_rKYBJCle1_0),.clk(gclk));
	jdff dff_A_kexKDfbr0_0(.dout(w_dff_A_rKYBJCle1_0),.din(w_dff_A_kexKDfbr0_0),.clk(gclk));
	jdff dff_A_Kr1W6KUY5_0(.dout(w_dff_A_kexKDfbr0_0),.din(w_dff_A_Kr1W6KUY5_0),.clk(gclk));
	jdff dff_A_nt8rdOU21_0(.dout(w_Gid12_0[0]),.din(w_dff_A_nt8rdOU21_0),.clk(gclk));
	jdff dff_A_uqCtPmK78_0(.dout(w_dff_A_nt8rdOU21_0),.din(w_dff_A_uqCtPmK78_0),.clk(gclk));
	jdff dff_A_mN7DoGtO0_0(.dout(w_dff_A_uqCtPmK78_0),.din(w_dff_A_mN7DoGtO0_0),.clk(gclk));
	jdff dff_A_YCGO4eY17_0(.dout(w_dff_A_mN7DoGtO0_0),.din(w_dff_A_YCGO4eY17_0),.clk(gclk));
	jdff dff_A_5bK44Lyn8_0(.dout(w_dff_A_YCGO4eY17_0),.din(w_dff_A_5bK44Lyn8_0),.clk(gclk));
	jdff dff_A_S2AYlz2y0_0(.dout(w_dff_A_5bK44Lyn8_0),.din(w_dff_A_S2AYlz2y0_0),.clk(gclk));
	jdff dff_A_156YnIVW1_0(.dout(w_dff_A_S2AYlz2y0_0),.din(w_dff_A_156YnIVW1_0),.clk(gclk));
	jdff dff_A_kWhGq2h96_0(.dout(w_dff_A_156YnIVW1_0),.din(w_dff_A_kWhGq2h96_0),.clk(gclk));
	jdff dff_A_qYT5kUyt1_0(.dout(w_dff_A_kWhGq2h96_0),.din(w_dff_A_qYT5kUyt1_0),.clk(gclk));
	jdff dff_A_y9UQfaWF4_0(.dout(w_Gid7_0[0]),.din(w_dff_A_y9UQfaWF4_0),.clk(gclk));
	jdff dff_A_TF025xm65_0(.dout(w_dff_A_y9UQfaWF4_0),.din(w_dff_A_TF025xm65_0),.clk(gclk));
	jdff dff_A_6uKN7KI02_0(.dout(w_dff_A_TF025xm65_0),.din(w_dff_A_6uKN7KI02_0),.clk(gclk));
	jdff dff_A_D2tEnZjR8_0(.dout(w_dff_A_6uKN7KI02_0),.din(w_dff_A_D2tEnZjR8_0),.clk(gclk));
	jdff dff_A_Gjh6vQlf6_0(.dout(w_dff_A_D2tEnZjR8_0),.din(w_dff_A_Gjh6vQlf6_0),.clk(gclk));
	jdff dff_A_WiWxKCtv5_0(.dout(w_dff_A_Gjh6vQlf6_0),.din(w_dff_A_WiWxKCtv5_0),.clk(gclk));
	jdff dff_A_KJ3azRhd9_0(.dout(w_dff_A_WiWxKCtv5_0),.din(w_dff_A_KJ3azRhd9_0),.clk(gclk));
	jdff dff_A_7bJDUGNK3_0(.dout(w_dff_A_KJ3azRhd9_0),.din(w_dff_A_7bJDUGNK3_0),.clk(gclk));
	jdff dff_A_O4hbQfBu2_0(.dout(w_dff_A_7bJDUGNK3_0),.din(w_dff_A_O4hbQfBu2_0),.clk(gclk));
	jdff dff_A_kkrNQRKE5_0(.dout(w_dff_A_O4hbQfBu2_0),.din(w_dff_A_kkrNQRKE5_0),.clk(gclk));
	jdff dff_A_ChfgxBH58_0(.dout(w_Gid6_0[0]),.din(w_dff_A_ChfgxBH58_0),.clk(gclk));
	jdff dff_A_ygmvpjdG3_0(.dout(w_dff_A_ChfgxBH58_0),.din(w_dff_A_ygmvpjdG3_0),.clk(gclk));
	jdff dff_A_b7N7qzQE2_0(.dout(w_dff_A_ygmvpjdG3_0),.din(w_dff_A_b7N7qzQE2_0),.clk(gclk));
	jdff dff_A_gpRYnFCl7_0(.dout(w_dff_A_b7N7qzQE2_0),.din(w_dff_A_gpRYnFCl7_0),.clk(gclk));
	jdff dff_A_VScFfyKD7_0(.dout(w_dff_A_gpRYnFCl7_0),.din(w_dff_A_VScFfyKD7_0),.clk(gclk));
	jdff dff_A_TALpwPhe1_0(.dout(w_dff_A_VScFfyKD7_0),.din(w_dff_A_TALpwPhe1_0),.clk(gclk));
	jdff dff_A_bD3AqHE21_0(.dout(w_dff_A_TALpwPhe1_0),.din(w_dff_A_bD3AqHE21_0),.clk(gclk));
	jdff dff_A_nusqCQWs6_0(.dout(w_dff_A_bD3AqHE21_0),.din(w_dff_A_nusqCQWs6_0),.clk(gclk));
	jdff dff_A_PFRawVxt0_0(.dout(w_dff_A_nusqCQWs6_0),.din(w_dff_A_PFRawVxt0_0),.clk(gclk));
	jdff dff_A_sNMh06Yt4_0(.dout(w_dff_A_PFRawVxt0_0),.din(w_dff_A_sNMh06Yt4_0),.clk(gclk));
	jdff dff_A_QK1h1veC1_0(.dout(w_Gid5_0[0]),.din(w_dff_A_QK1h1veC1_0),.clk(gclk));
	jdff dff_A_UTKoS5Yv5_0(.dout(w_dff_A_QK1h1veC1_0),.din(w_dff_A_UTKoS5Yv5_0),.clk(gclk));
	jdff dff_A_0ibMUIzf3_0(.dout(w_dff_A_UTKoS5Yv5_0),.din(w_dff_A_0ibMUIzf3_0),.clk(gclk));
	jdff dff_A_wPOUYrxu9_0(.dout(w_dff_A_0ibMUIzf3_0),.din(w_dff_A_wPOUYrxu9_0),.clk(gclk));
	jdff dff_A_xpiFaIlY9_0(.dout(w_dff_A_wPOUYrxu9_0),.din(w_dff_A_xpiFaIlY9_0),.clk(gclk));
	jdff dff_A_ms0oWAOE9_0(.dout(w_dff_A_xpiFaIlY9_0),.din(w_dff_A_ms0oWAOE9_0),.clk(gclk));
	jdff dff_A_qhXLmvOf5_0(.dout(w_dff_A_ms0oWAOE9_0),.din(w_dff_A_qhXLmvOf5_0),.clk(gclk));
	jdff dff_A_fOFV1D9z7_0(.dout(w_dff_A_qhXLmvOf5_0),.din(w_dff_A_fOFV1D9z7_0),.clk(gclk));
	jdff dff_A_nQbZTHNI7_0(.dout(w_dff_A_fOFV1D9z7_0),.din(w_dff_A_nQbZTHNI7_0),.clk(gclk));
	jdff dff_A_BfT7Vhzc5_0(.dout(w_dff_A_nQbZTHNI7_0),.din(w_dff_A_BfT7Vhzc5_0),.clk(gclk));
	jdff dff_A_yR6PgPst6_0(.dout(w_Gid4_0[0]),.din(w_dff_A_yR6PgPst6_0),.clk(gclk));
	jdff dff_A_Vw3TsTGp2_0(.dout(w_dff_A_yR6PgPst6_0),.din(w_dff_A_Vw3TsTGp2_0),.clk(gclk));
	jdff dff_A_SKUvScIw6_0(.dout(w_dff_A_Vw3TsTGp2_0),.din(w_dff_A_SKUvScIw6_0),.clk(gclk));
	jdff dff_A_V2rYNcDl9_0(.dout(w_dff_A_SKUvScIw6_0),.din(w_dff_A_V2rYNcDl9_0),.clk(gclk));
	jdff dff_A_AJR36qPJ9_0(.dout(w_dff_A_V2rYNcDl9_0),.din(w_dff_A_AJR36qPJ9_0),.clk(gclk));
	jdff dff_A_uziHMTnu4_0(.dout(w_dff_A_AJR36qPJ9_0),.din(w_dff_A_uziHMTnu4_0),.clk(gclk));
	jdff dff_A_CrOmOJbG8_0(.dout(w_dff_A_uziHMTnu4_0),.din(w_dff_A_CrOmOJbG8_0),.clk(gclk));
	jdff dff_A_kr8LbF5O2_0(.dout(w_dff_A_CrOmOJbG8_0),.din(w_dff_A_kr8LbF5O2_0),.clk(gclk));
	jdff dff_A_OEBpZGBL0_0(.dout(w_dff_A_kr8LbF5O2_0),.din(w_dff_A_OEBpZGBL0_0),.clk(gclk));
	jdff dff_A_ZgwJAPqV3_0(.dout(w_dff_A_OEBpZGBL0_0),.din(w_dff_A_ZgwJAPqV3_0),.clk(gclk));
	jdff dff_A_xZiBlxD60_2(.dout(God8),.din(w_dff_A_xZiBlxD60_2),.clk(gclk));
	jdff dff_A_GC3Ur5fC0_2(.dout(God9),.din(w_dff_A_GC3Ur5fC0_2),.clk(gclk));
	jdff dff_A_qT9JmB3C5_2(.dout(God10),.din(w_dff_A_qT9JmB3C5_2),.clk(gclk));
	jdff dff_A_2iNFlhGO6_2(.dout(God11),.din(w_dff_A_2iNFlhGO6_2),.clk(gclk));
	jdff dff_A_k1Z9d4Mf4_2(.dout(God12),.din(w_dff_A_k1Z9d4Mf4_2),.clk(gclk));
	jdff dff_A_2woWXhQe4_2(.dout(God13),.din(w_dff_A_2woWXhQe4_2),.clk(gclk));
	jdff dff_A_02xLMDyO5_2(.dout(God14),.din(w_dff_A_02xLMDyO5_2),.clk(gclk));
	jdff dff_A_XsRivswP4_2(.dout(God15),.din(w_dff_A_XsRivswP4_2),.clk(gclk));
endmodule

