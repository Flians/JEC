// Benchmark "c2670" written by ABC on Wed May 27 22:06:37 2020

module gf_c2670 ( 
    G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
    G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
    G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
    G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
    G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
    G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
    G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120,
    G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136,
    G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180,
    G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194,
    G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206,
    G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241,
    G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253,
    G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269,
    G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452, G483,
    G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384,
    G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066,
    G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106,
    G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20,
    G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36,
    G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56,
    G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74,
    G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90,
    G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105,
    G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
    G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135,
    G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179,
    G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193,
    G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205,
    G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240,
    G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252,
    G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268,
    G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279, G452,
    G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348,
    G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996,
    G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105,
    G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474,
    G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire n381, n382, n383, n384, n385, n386, n388, n389, n390, n391, n394,
    n396, n398, n400, n401, n402, n403, n404, n405, n408, n409, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n438,
    n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n450, n451,
    n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n464, n465,
    n466, n467, n468, n469, n470, n473, n474, n475, n476, n477, n478, n479,
    n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n497, n498, n499, n500, n501, n503, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n517, n518, n519, n520, n521,
    n522, n524, n525, n526, n527, n528, n529, n530, n532, n533, n534, n535,
    n536, n537, n538, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n556, n557, n559, n561, n562, n563,
    n564, n565, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n594, n595, n596, n597, n598, n599, n600, n602, n603,
    n604, n605, n606, n607, n608, n609, n610, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
    n812, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n828, n829, n830, n831, n832, n833, n834, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
    n947, n950, n951, n952, n953;
  jnot g000(.din(G44), .dout(G218));
  jnot g001(.din(G132), .dout(G219));
  jnot g002(.din(G82), .dout(G220));
  jnot g003(.din(G96), .dout(G221));
  jnot g004(.din(G69), .dout(G235));
  jnot g005(.din(G120), .dout(G236));
  jnot g006(.din(G57), .dout(G237));
  jnot g007(.din(G108), .dout(G238));
  jnot g008(.din(G2084), .dout(n381));
  jnot g009(.din(G2090), .dout(n382));
  jor  g010(.dina(n382), .dinb(n381), .dout(n383));
  jnot g011(.din(G2072), .dout(n384));
  jnot g012(.din(G2078), .dout(n385));
  jor  g013(.dina(n385), .dinb(n384), .dout(n386));
  jor  g014(.dina(n386), .dinb(n383), .dout(G158));
  jnot g015(.din(G15), .dout(n388));
  jnot g016(.din(G2), .dout(n389));
  jnot g017(.din(G661), .dout(n390));
  jor  g018(.dina(n390), .dinb(n389), .dout(n391));
  jor  g019(.dina(n391), .dinb(n388), .dout(G259));
  jand g020(.dina(G452), .dinb(G94), .dout(G173));
  jnot g021(.din(G7), .dout(n394));
  jor  g022(.dina(n390), .dinb(n394), .dout(G223));
  jnot g023(.din(G567), .dout(n396));
  jor  g024(.dina(G223), .dinb(n396), .dout(G234));
  jnot g025(.din(G2106), .dout(n398));
  jor  g026(.dina(G223), .dinb(n398), .dout(G217));
  jand g027(.dina(G108), .dinb(G69), .dout(n400));
  jand g028(.dina(G120), .dinb(G57), .dout(n401));
  jand g029(.dina(n401), .dinb(n400), .dout(n402));
  jand g030(.dina(G96), .dinb(G82), .dout(n403));
  jand g031(.dina(G132), .dinb(G44), .dout(n404));
  jand g032(.dina(n404), .dinb(n403), .dout(n405));
  jand g033(.dina(n405), .dinb(n402), .dout(G325));
  jnot g034(.din(G325), .dout(G261));
  jor  g035(.dina(n405), .dinb(n398), .dout(n408));
  jor  g036(.dina(n402), .dinb(n396), .dout(n409));
  jand g037(.dina(n409), .dinb(n408), .dout(G319));
  jnot g038(.din(G2104), .dout(n411));
  jand g039(.dina(G2105), .dinb(n411), .dout(n412));
  jand g040(.dina(n412), .dinb(G125), .dout(n413));
  jnot g041(.din(n413), .dout(n414));
  jnot g042(.din(G101), .dout(n415));
  jor  g043(.dina(G2105), .dinb(n411), .dout(n416));
  jor  g044(.dina(n416), .dinb(n415), .dout(n417));
  jnot g045(.din(G137), .dout(n418));
  jor  g046(.dina(G2105), .dinb(G2104), .dout(n419));
  jor  g047(.dina(n419), .dinb(n418), .dout(n420));
  jand g048(.dina(n420), .dinb(n417), .dout(n421));
  jand g049(.dina(G2105), .dinb(G2104), .dout(n422));
  jand g050(.dina(n422), .dinb(G113), .dout(n423));
  jnot g051(.din(n423), .dout(n424));
  jand g052(.dina(n424), .dinb(n421), .dout(n425));
  jand g053(.dina(n425), .dinb(n414), .dout(G160));
  jand g054(.dina(n412), .dinb(G124), .dout(n427));
  jnot g055(.din(G2105), .dout(n428));
  jand g056(.dina(n428), .dinb(G2104), .dout(n429));
  jand g057(.dina(n429), .dinb(G100), .dout(n430));
  jand g058(.dina(n428), .dinb(n411), .dout(n431));
  jand g059(.dina(n431), .dinb(G136), .dout(n432));
  jor  g060(.dina(n432), .dinb(n430), .dout(n433));
  jand g061(.dina(n422), .dinb(G112), .dout(n434));
  jor  g062(.dina(n434), .dinb(n433), .dout(n435));
  jor  g063(.dina(n435), .dinb(n427), .dout(n436));
  jnot g064(.din(n436), .dout(G162));
  jand g065(.dina(n431), .dinb(G138), .dout(n438));
  jnot g066(.din(n438), .dout(n439));
  jnot g067(.din(G102), .dout(n440));
  jor  g068(.dina(n416), .dinb(n440), .dout(n441));
  jnot g069(.din(G126), .dout(n442));
  jor  g070(.dina(n428), .dinb(G2104), .dout(n443));
  jor  g071(.dina(n443), .dinb(n442), .dout(n444));
  jand g072(.dina(n444), .dinb(n441), .dout(n445));
  jand g073(.dina(n422), .dinb(G114), .dout(n446));
  jnot g074(.din(n446), .dout(n447));
  jand g075(.dina(n447), .dinb(n445), .dout(n448));
  jand g076(.dina(n448), .dinb(n439), .dout(G164));
  jand g077(.dina(G651), .dinb(G543), .dout(n450));
  jand g078(.dina(n450), .dinb(G75), .dout(n451));
  jnot g079(.din(G651), .dout(n452));
  jor  g080(.dina(n452), .dinb(G543), .dout(n453));
  jnot g081(.din(n453), .dout(n454));
  jand g082(.dina(n454), .dinb(G62), .dout(n455));
  jor  g083(.dina(n455), .dinb(n451), .dout(n456));
  jor  g084(.dina(G543), .dinb(G88), .dout(n457));
  jnot g085(.din(G543), .dout(n458));
  jor  g086(.dina(n458), .dinb(G50), .dout(n459));
  jand g087(.dina(n459), .dinb(n457), .dout(n460));
  jand g088(.dina(n460), .dinb(n452), .dout(n461));
  jor  g089(.dina(n461), .dinb(n456), .dout(G303));
  jnot g090(.din(G303), .dout(G166));
  jand g091(.dina(n450), .dinb(G76), .dout(n464));
  jand g092(.dina(n454), .dinb(G63), .dout(n465));
  jor  g093(.dina(n465), .dinb(n464), .dout(n466));
  jor  g094(.dina(G543), .dinb(G89), .dout(n467));
  jor  g095(.dina(n458), .dinb(G51), .dout(n468));
  jand g096(.dina(n468), .dinb(n467), .dout(n469));
  jand g097(.dina(n469), .dinb(n452), .dout(n470));
  jor  g098(.dina(n470), .dinb(n466), .dout(G286));
  jnot g099(.din(G286), .dout(G168));
  jand g100(.dina(n450), .dinb(G77), .dout(n473));
  jand g101(.dina(n454), .dinb(G64), .dout(n474));
  jor  g102(.dina(n474), .dinb(n473), .dout(n475));
  jor  g103(.dina(G543), .dinb(G90), .dout(n476));
  jor  g104(.dina(n458), .dinb(G52), .dout(n477));
  jand g105(.dina(n477), .dinb(n476), .dout(n478));
  jand g106(.dina(n478), .dinb(n452), .dout(n479));
  jor  g107(.dina(n479), .dinb(n475), .dout(G301));
  jnot g108(.din(G301), .dout(G171));
  jnot g109(.din(G860), .dout(n482));
  jand g110(.dina(n450), .dinb(G68), .dout(n483));
  jnot g111(.din(n483), .dout(n484));
  jnot g112(.din(G56), .dout(n485));
  jor  g113(.dina(n453), .dinb(n485), .dout(n486));
  jand g114(.dina(n486), .dinb(n484), .dout(n487));
  jor  g115(.dina(G543), .dinb(G81), .dout(n488));
  jnot g116(.din(n488), .dout(n489));
  jnot g117(.din(G43), .dout(n490));
  jand g118(.dina(G543), .dinb(n490), .dout(n491));
  jor  g119(.dina(n491), .dinb(n489), .dout(n492));
  jor  g120(.dina(n492), .dinb(G651), .dout(n493));
  jand g121(.dina(n493), .dinb(n487), .dout(n494));
  jnot g122(.din(n494), .dout(n495));
  jor  g123(.dina(n495), .dinb(n482), .dout(G153));
  jnot g124(.din(G36), .dout(n497));
  jnot g125(.din(G483), .dout(n498));
  jnot g126(.din(G319), .dout(n499));
  jor  g127(.dina(n499), .dinb(n498), .dout(n500));
  jor  g128(.dina(n500), .dinb(n390), .dout(n501));
  jor  g129(.dina(n501), .dinb(n497), .dout(G176));
  jand g130(.dina(G3), .dinb(G1), .dout(n503));
  jor  g131(.dina(n503), .dinb(n501), .dout(G188));
  jand g132(.dina(n450), .dinb(G78), .dout(n505));
  jnot g133(.din(n505), .dout(n506));
  jnot g134(.din(G65), .dout(n507));
  jor  g135(.dina(n453), .dinb(n507), .dout(n508));
  jand g136(.dina(n508), .dinb(n506), .dout(n509));
  jor  g137(.dina(G543), .dinb(G91), .dout(n510));
  jor  g138(.dina(n458), .dinb(G53), .dout(n511));
  jand g139(.dina(n511), .dinb(n510), .dout(n512));
  jand g140(.dina(n512), .dinb(n452), .dout(n513));
  jnot g141(.din(n513), .dout(n514));
  jand g142(.dina(n514), .dinb(n509), .dout(n515));
  jnot g143(.din(n515), .dout(G299));
  jnot g144(.din(n450), .dout(n517));
  jor  g145(.dina(n517), .dinb(G74), .dout(n518));
  jand g146(.dina(n458), .dinb(G87), .dout(n519));
  jand g147(.dina(G543), .dinb(G49), .dout(n520));
  jor  g148(.dina(n520), .dinb(n519), .dout(n521));
  jor  g149(.dina(n521), .dinb(G651), .dout(n522));
  jand g150(.dina(n522), .dinb(n518), .dout(G288));
  jand g151(.dina(n450), .dinb(G73), .dout(n524));
  jand g152(.dina(n454), .dinb(G61), .dout(n525));
  jor  g153(.dina(n525), .dinb(n524), .dout(n526));
  jor  g154(.dina(G543), .dinb(G86), .dout(n527));
  jor  g155(.dina(n458), .dinb(G48), .dout(n528));
  jand g156(.dina(n528), .dinb(n527), .dout(n529));
  jand g157(.dina(n529), .dinb(n452), .dout(n530));
  jor  g158(.dina(n530), .dinb(n526), .dout(G305));
  jand g159(.dina(n450), .dinb(G72), .dout(n532));
  jand g160(.dina(n454), .dinb(G60), .dout(n533));
  jor  g161(.dina(n533), .dinb(n532), .dout(n534));
  jor  g162(.dina(G543), .dinb(G85), .dout(n535));
  jor  g163(.dina(n458), .dinb(G47), .dout(n536));
  jand g164(.dina(n536), .dinb(n535), .dout(n537));
  jand g165(.dina(n537), .dinb(n452), .dout(n538));
  jor  g166(.dina(n538), .dinb(n534), .dout(G290));
  jnot g167(.din(G868), .dout(n540));
  jor  g168(.dina(G301), .dinb(n540), .dout(n541));
  jand g169(.dina(n450), .dinb(G79), .dout(n542));
  jnot g170(.din(n542), .dout(n543));
  jnot g171(.din(G66), .dout(n544));
  jor  g172(.dina(n453), .dinb(n544), .dout(n545));
  jand g173(.dina(n545), .dinb(n543), .dout(n546));
  jor  g174(.dina(G543), .dinb(G92), .dout(n547));
  jor  g175(.dina(n458), .dinb(G54), .dout(n548));
  jand g176(.dina(n548), .dinb(n547), .dout(n549));
  jand g177(.dina(n549), .dinb(n452), .dout(n550));
  jnot g178(.din(n550), .dout(n551));
  jand g179(.dina(n551), .dinb(n546), .dout(n552));
  jnot g180(.din(n552), .dout(n553));
  jor  g181(.dina(n553), .dinb(G868), .dout(n554));
  jand g182(.dina(n554), .dinb(n541), .dout(G284));
  jor  g183(.dina(G286), .dinb(n540), .dout(n556));
  jor  g184(.dina(G299), .dinb(G868), .dout(n557));
  jand g185(.dina(n557), .dinb(n556), .dout(G297));
  jand g186(.dina(n482), .dinb(G559), .dout(n559));
  jor  g187(.dina(n559), .dinb(n553), .dout(G148));
  jnot g188(.din(G559), .dout(n561));
  jand g189(.dina(n552), .dinb(n561), .dout(n562));
  jnot g190(.din(n562), .dout(n563));
  jor  g191(.dina(n563), .dinb(n540), .dout(n564));
  jor  g192(.dina(n495), .dinb(G868), .dout(n565));
  jand g193(.dina(n565), .dinb(n564), .dout(G282));
  jnot g194(.din(G2096), .dout(n567));
  jand g195(.dina(n412), .dinb(G123), .dout(n568));
  jand g196(.dina(n429), .dinb(G99), .dout(n569));
  jand g197(.dina(n431), .dinb(G135), .dout(n570));
  jor  g198(.dina(n570), .dinb(n569), .dout(n571));
  jand g199(.dina(n422), .dinb(G111), .dout(n572));
  jor  g200(.dina(n572), .dinb(n571), .dout(n573));
  jor  g201(.dina(n573), .dinb(n568), .dout(n574));
  jnot g202(.din(n574), .dout(n575));
  jand g203(.dina(n575), .dinb(n567), .dout(n576));
  jand g204(.dina(n574), .dinb(G2096), .dout(n577));
  jor  g205(.dina(n577), .dinb(G2100), .dout(n578));
  jor  g206(.dina(n578), .dinb(n576), .dout(G156));
  jxor g207(.dina(G2454), .dinb(G2451), .dout(n580));
  jxor g208(.dina(G1348), .dinb(G1341), .dout(n581));
  jxor g209(.dina(n581), .dinb(n580), .dout(n582));
  jxor g210(.dina(G2430), .dinb(G2427), .dout(n583));
  jxor g211(.dina(G2446), .dinb(G2443), .dout(n584));
  jxor g212(.dina(G2438), .dinb(G2435), .dout(n585));
  jxor g213(.dina(n585), .dinb(n584), .dout(n586));
  jxor g214(.dina(n586), .dinb(n583), .dout(n587));
  jnot g215(.din(n587), .dout(n588));
  jand g216(.dina(n588), .dinb(n582), .dout(n589));
  jnot g217(.din(n589), .dout(n590));
  jor  g218(.dina(n588), .dinb(n582), .dout(n591));
  jand g219(.dina(n591), .dinb(G14), .dout(n592));
  jand g220(.dina(n592), .dinb(n590), .dout(G401));
  jxor g221(.dina(G2078), .dinb(G2072), .dout(n594));
  jxor g222(.dina(G2100), .dinb(G2096), .dout(n595));
  jxor g223(.dina(n595), .dinb(n594), .dout(n596));
  jxor g224(.dina(G2090), .dinb(G2084), .dout(n597));
  jnot g225(.din(G2067), .dout(n598));
  jxor g226(.dina(G2678), .dinb(n598), .dout(n599));
  jxor g227(.dina(n599), .dinb(n597), .dout(n600));
  jxor g228(.dina(n600), .dinb(n596), .dout(G227));
  jxor g229(.dina(G1966), .dinb(G1961), .dout(n602));
  jnot g230(.din(G1991), .dout(n603));
  jxor g231(.dina(G1996), .dinb(n603), .dout(n604));
  jxor g232(.dina(n604), .dinb(n602), .dout(n605));
  jxor g233(.dina(G2474), .dinb(G1976), .dout(n606));
  jxor g234(.dina(G1971), .dinb(G1956), .dout(n607));
  jxor g235(.dina(n607), .dinb(n606), .dout(n608));
  jxor g236(.dina(G1986), .dinb(G1981), .dout(n609));
  jxor g237(.dina(n609), .dinb(n608), .dout(n610));
  jxor g238(.dina(n610), .dinb(n605), .dout(G229));
  jand g239(.dina(G160), .dinb(G29), .dout(n612));
  jnot g240(.din(n612), .dout(n613));
  jor  g241(.dina(G34), .dinb(G29), .dout(n614));
  jand g242(.dina(n614), .dinb(n613), .dout(n615));
  jand g243(.dina(n615), .dinb(G2084), .dout(n616));
  jand g244(.dina(n412), .dinb(G128), .dout(n617));
  jand g245(.dina(n429), .dinb(G104), .dout(n618));
  jand g246(.dina(n431), .dinb(G140), .dout(n619));
  jor  g247(.dina(n619), .dinb(n618), .dout(n620));
  jand g248(.dina(n422), .dinb(G116), .dout(n621));
  jor  g249(.dina(n621), .dinb(n620), .dout(n622));
  jor  g250(.dina(n622), .dinb(n617), .dout(n623));
  jnot g251(.din(n623), .dout(n624));
  jand g252(.dina(n624), .dinb(G29), .dout(n625));
  jnot g253(.din(n625), .dout(n626));
  jor  g254(.dina(G29), .dinb(G26), .dout(n627));
  jand g255(.dina(n627), .dinb(n626), .dout(n628));
  jnot g256(.din(n628), .dout(n629));
  jand g257(.dina(n629), .dinb(n598), .dout(n630));
  jor  g258(.dina(n630), .dinb(n616), .dout(n631));
  jnot g259(.din(n631), .dout(n632));
  jand g260(.dina(G164), .dinb(G29), .dout(n633));
  jnot g261(.din(n633), .dout(n634));
  jor  g262(.dina(G29), .dinb(G27), .dout(n635));
  jand g263(.dina(n635), .dinb(n634), .dout(n636));
  jand g264(.dina(n636), .dinb(G2078), .dout(n637));
  jnot g265(.din(n637), .dout(n638));
  jor  g266(.dina(G23), .dinb(G16), .dout(n639));
  jnot g267(.din(G16), .dout(n640));
  jor  g268(.dina(G288), .dinb(n640), .dout(n641));
  jand g269(.dina(n641), .dinb(n639), .dout(n642));
  jxor g270(.dina(n642), .dinb(G1976), .dout(n643));
  jand g271(.dina(n643), .dinb(n638), .dout(n644));
  jand g272(.dina(n644), .dinb(n632), .dout(n645));
  jnot g273(.din(G1966), .dout(n646));
  jand g274(.dina(G168), .dinb(G16), .dout(n647));
  jnot g275(.din(n647), .dout(n648));
  jor  g276(.dina(G21), .dinb(G16), .dout(n649));
  jand g277(.dina(n649), .dinb(n648), .dout(n650));
  jnot g278(.din(n650), .dout(n651));
  jand g279(.dina(n651), .dinb(n646), .dout(n652));
  jnot g280(.din(n652), .dout(n653));
  jor  g281(.dina(n495), .dinb(n640), .dout(n654));
  jor  g282(.dina(G19), .dinb(G16), .dout(n655));
  jand g283(.dina(n655), .dinb(n654), .dout(n656));
  jxor g284(.dina(n656), .dinb(G1341), .dout(n657));
  jand g285(.dina(n657), .dinb(n653), .dout(n658));
  jor  g286(.dina(n615), .dinb(G2084), .dout(n659));
  jnot g287(.din(G29), .dout(n660));
  jand g288(.dina(n660), .dinb(G28), .dout(n661));
  jand g289(.dina(n574), .dinb(G29), .dout(n662));
  jor  g290(.dina(n662), .dinb(n661), .dout(n663));
  jand g291(.dina(n663), .dinb(n659), .dout(n664));
  jand g292(.dina(n431), .dinb(G141), .dout(n665));
  jand g293(.dina(n429), .dinb(G105), .dout(n666));
  jand g294(.dina(n412), .dinb(G129), .dout(n667));
  jor  g295(.dina(n667), .dinb(n666), .dout(n668));
  jand g296(.dina(n422), .dinb(G117), .dout(n669));
  jor  g297(.dina(n669), .dinb(n668), .dout(n670));
  jor  g298(.dina(n670), .dinb(n665), .dout(n671));
  jor  g299(.dina(n671), .dinb(n660), .dout(n672));
  jor  g300(.dina(G32), .dinb(G29), .dout(n673));
  jand g301(.dina(n673), .dinb(n672), .dout(n674));
  jxor g302(.dina(n674), .dinb(G1996), .dout(n675));
  jand g303(.dina(n675), .dinb(n664), .dout(n676));
  jand g304(.dina(n676), .dinb(n658), .dout(n677));
  jnot g305(.din(G305), .dout(n678));
  jand g306(.dina(n678), .dinb(G16), .dout(n679));
  jnot g307(.din(n679), .dout(n680));
  jor  g308(.dina(G16), .dinb(G6), .dout(n681));
  jand g309(.dina(n681), .dinb(n680), .dout(n682));
  jand g310(.dina(n682), .dinb(G1981), .dout(n683));
  jand g311(.dina(n422), .dinb(G115), .dout(n684));
  jand g312(.dina(n429), .dinb(G103), .dout(n685));
  jand g313(.dina(n412), .dinb(G127), .dout(n686));
  jor  g314(.dina(n686), .dinb(n685), .dout(n687));
  jand g315(.dina(n431), .dinb(G139), .dout(n688));
  jor  g316(.dina(n688), .dinb(n687), .dout(n689));
  jor  g317(.dina(n689), .dinb(n684), .dout(n690));
  jor  g318(.dina(n690), .dinb(n660), .dout(n691));
  jor  g319(.dina(G33), .dinb(G29), .dout(n692));
  jand g320(.dina(n692), .dinb(n691), .dout(n693));
  jxor g321(.dina(n693), .dinb(n384), .dout(n694));
  jor  g322(.dina(n694), .dinb(n683), .dout(n695));
  jnot g323(.din(n695), .dout(n696));
  jand g324(.dina(n696), .dinb(n677), .dout(n697));
  jand g325(.dina(n697), .dinb(n645), .dout(n698));
  jand g326(.dina(G162), .dinb(G29), .dout(n699));
  jnot g327(.din(n699), .dout(n700));
  jor  g328(.dina(G35), .dinb(G29), .dout(n701));
  jand g329(.dina(n701), .dinb(n700), .dout(n702));
  jand g330(.dina(n702), .dinb(G2090), .dout(n703));
  jnot g331(.din(n703), .dout(n704));
  jand g332(.dina(n704), .dinb(G11), .dout(n705));
  jor  g333(.dina(n553), .dinb(n640), .dout(n706));
  jor  g334(.dina(G16), .dinb(G4), .dout(n707));
  jand g335(.dina(n707), .dinb(n706), .dout(n708));
  jxor g336(.dina(n708), .dinb(G1348), .dout(n709));
  jand g337(.dina(n709), .dinb(n705), .dout(n710));
  jand g338(.dina(n628), .dinb(G2067), .dout(n711));
  jnot g339(.din(n711), .dout(n712));
  jor  g340(.dina(n702), .dinb(G2090), .dout(n713));
  jand g341(.dina(n713), .dinb(n712), .dout(n714));
  jnot g342(.din(G1986), .dout(n715));
  jnot g343(.din(G290), .dout(n716));
  jand g344(.dina(n716), .dinb(G16), .dout(n717));
  jnot g345(.din(n717), .dout(n718));
  jor  g346(.dina(G24), .dinb(G16), .dout(n719));
  jand g347(.dina(n719), .dinb(n718), .dout(n720));
  jnot g348(.din(n720), .dout(n721));
  jand g349(.dina(n721), .dinb(n715), .dout(n722));
  jand g350(.dina(n650), .dinb(G1966), .dout(n723));
  jor  g351(.dina(n723), .dinb(n722), .dout(n724));
  jnot g352(.din(n724), .dout(n725));
  jand g353(.dina(n725), .dinb(n714), .dout(n726));
  jand g354(.dina(n720), .dinb(G1986), .dout(n727));
  jnot g355(.din(n727), .dout(n728));
  jor  g356(.dina(G301), .dinb(n640), .dout(n729));
  jor  g357(.dina(G16), .dinb(G5), .dout(n730));
  jand g358(.dina(n730), .dinb(n729), .dout(n731));
  jxor g359(.dina(n731), .dinb(G1961), .dout(n732));
  jand g360(.dina(n732), .dinb(n728), .dout(n733));
  jand g361(.dina(n733), .dinb(n726), .dout(n734));
  jor  g362(.dina(n636), .dinb(G2078), .dout(n735));
  jnot g363(.din(G1956), .dout(n736));
  jor  g364(.dina(G299), .dinb(n640), .dout(n737));
  jor  g365(.dina(G20), .dinb(G16), .dout(n738));
  jand g366(.dina(n738), .dinb(n737), .dout(n739));
  jxor g367(.dina(n739), .dinb(n736), .dout(n740));
  jnot g368(.din(n740), .dout(n741));
  jand g369(.dina(n741), .dinb(n735), .dout(n742));
  jnot g370(.din(G1971), .dout(n743));
  jand g371(.dina(G166), .dinb(G16), .dout(n744));
  jnot g372(.din(n744), .dout(n745));
  jor  g373(.dina(G22), .dinb(G16), .dout(n746));
  jand g374(.dina(n746), .dinb(n745), .dout(n747));
  jnot g375(.din(n747), .dout(n748));
  jand g376(.dina(n748), .dinb(n743), .dout(n749));
  jnot g377(.din(n749), .dout(n750));
  jand g378(.dina(n750), .dinb(n742), .dout(n751));
  jor  g379(.dina(n682), .dinb(G1981), .dout(n752));
  jand g380(.dina(n747), .dinb(G1971), .dout(n753));
  jnot g381(.din(n753), .dout(n754));
  jand g382(.dina(n754), .dinb(n752), .dout(n755));
  jand g383(.dina(n422), .dinb(G107), .dout(n756));
  jand g384(.dina(n429), .dinb(G95), .dout(n757));
  jand g385(.dina(n431), .dinb(G131), .dout(n758));
  jor  g386(.dina(n758), .dinb(n757), .dout(n759));
  jand g387(.dina(n412), .dinb(G119), .dout(n760));
  jor  g388(.dina(n760), .dinb(n759), .dout(n761));
  jor  g389(.dina(n761), .dinb(n756), .dout(n762));
  jor  g390(.dina(n762), .dinb(n660), .dout(n763));
  jor  g391(.dina(G29), .dinb(G25), .dout(n764));
  jand g392(.dina(n764), .dinb(n763), .dout(n765));
  jxor g393(.dina(n765), .dinb(n603), .dout(n766));
  jnot g394(.din(n766), .dout(n767));
  jand g395(.dina(n767), .dinb(n755), .dout(n768));
  jand g396(.dina(n768), .dinb(n751), .dout(n769));
  jand g397(.dina(n769), .dinb(n734), .dout(n770));
  jand g398(.dina(n770), .dinb(n710), .dout(n771));
  jand g399(.dina(n771), .dinb(n698), .dout(G311));
  jnot g400(.din(G311), .dout(G150));
  jand g401(.dina(n450), .dinb(G80), .dout(n774));
  jand g402(.dina(n454), .dinb(G67), .dout(n775));
  jor  g403(.dina(n775), .dinb(n774), .dout(n776));
  jor  g404(.dina(G543), .dinb(G93), .dout(n777));
  jor  g405(.dina(n458), .dinb(G55), .dout(n778));
  jand g406(.dina(n778), .dinb(n777), .dout(n779));
  jand g407(.dina(n779), .dinb(n452), .dout(n780));
  jor  g408(.dina(n780), .dinb(n776), .dout(n781));
  jand g409(.dina(n781), .dinb(G860), .dout(n782));
  jor  g410(.dina(n553), .dinb(n561), .dout(n783));
  jxor g411(.dina(n781), .dinb(n495), .dout(n784));
  jxor g412(.dina(n784), .dinb(n783), .dout(n785));
  jand g413(.dina(n785), .dinb(n482), .dout(n786));
  jor  g414(.dina(n786), .dinb(n782), .dout(G145));
  jxor g415(.dina(n575), .dinb(n436), .dout(n788));
  jxor g416(.dina(n788), .dinb(G160), .dout(n789));
  jnot g417(.din(n789), .dout(n790));
  jand g418(.dina(n429), .dinb(G102), .dout(n791));
  jand g419(.dina(n412), .dinb(G126), .dout(n792));
  jor  g420(.dina(n792), .dinb(n791), .dout(n793));
  jor  g421(.dina(n446), .dinb(n793), .dout(n794));
  jor  g422(.dina(n794), .dinb(n438), .dout(n795));
  jxor g423(.dina(n623), .dinb(n795), .dout(n796));
  jand g424(.dina(n412), .dinb(G130), .dout(n797));
  jand g425(.dina(n429), .dinb(G106), .dout(n798));
  jand g426(.dina(n431), .dinb(G142), .dout(n799));
  jor  g427(.dina(n799), .dinb(n798), .dout(n800));
  jand g428(.dina(n422), .dinb(G118), .dout(n801));
  jor  g429(.dina(n801), .dinb(n800), .dout(n802));
  jor  g430(.dina(n802), .dinb(n797), .dout(n803));
  jxor g431(.dina(n803), .dinb(n690), .dout(n804));
  jxor g432(.dina(n762), .dinb(n671), .dout(n805));
  jxor g433(.dina(n805), .dinb(n804), .dout(n806));
  jxor g434(.dina(n806), .dinb(n796), .dout(n807));
  jnot g435(.din(n807), .dout(n808));
  jand g436(.dina(n808), .dinb(n790), .dout(n809));
  jand g437(.dina(n807), .dinb(n789), .dout(n810));
  jor  g438(.dina(n810), .dinb(G37), .dout(n811));
  jor  g439(.dina(n811), .dinb(n809), .dout(n812));
  jnot g440(.din(n812), .dout(G395));
  jor  g441(.dina(n781), .dinb(G868), .dout(n814));
  jand g442(.dina(n814), .dinb(n564), .dout(n815));
  jxor g443(.dina(n552), .dinb(G299), .dout(n816));
  jxor g444(.dina(n816), .dinb(n784), .dout(n817));
  jnot g445(.din(G288), .dout(n818));
  jxor g446(.dina(n818), .dinb(G303), .dout(n819));
  jxor g447(.dina(G290), .dinb(G305), .dout(n820));
  jxor g448(.dina(n820), .dinb(n819), .dout(n821));
  jxor g449(.dina(n821), .dinb(n817), .dout(n822));
  jand g450(.dina(n822), .dinb(G868), .dout(n823));
  jor  g451(.dina(n823), .dinb(n815), .dout(n824));
  jnot g452(.din(n823), .dout(n825));
  jor  g453(.dina(n825), .dinb(n562), .dout(n826));
  jand g454(.dina(n826), .dinb(n824), .dout(G295));
  jnot g455(.din(n822), .dout(n828));
  jxor g456(.dina(G171), .dinb(G286), .dout(n829));
  jnot g457(.din(n829), .dout(n830));
  jand g458(.dina(n830), .dinb(n828), .dout(n831));
  jand g459(.dina(n829), .dinb(n822), .dout(n832));
  jor  g460(.dina(n832), .dinb(G37), .dout(n833));
  jor  g461(.dina(n833), .dinb(n831), .dout(n834));
  jnot g462(.din(n834), .dout(G397));
  jor  g463(.dina(G164), .dinb(G1384), .dout(n836));
  jand g464(.dina(G160), .dinb(G40), .dout(n837));
  jand g465(.dina(n837), .dinb(n836), .dout(n838));
  jand g466(.dina(n838), .dinb(n716), .dout(n839));
  jand g467(.dina(n839), .dinb(n715), .dout(n840));
  jnot g468(.din(n840), .dout(n841));
  jnot g469(.din(n838), .dout(n842));
  jnot g470(.din(n762), .dout(n843));
  jor  g471(.dina(n843), .dinb(n603), .dout(n844));
  jor  g472(.dina(n844), .dinb(n842), .dout(n845));
  jand g473(.dina(n838), .dinb(n843), .dout(n846));
  jand g474(.dina(n846), .dinb(n603), .dout(n847));
  jnot g475(.din(n847), .dout(n848));
  jnot g476(.din(G40), .dout(n849));
  jand g477(.dina(n429), .dinb(G101), .dout(n850));
  jand g478(.dina(n431), .dinb(G137), .dout(n851));
  jor  g479(.dina(n851), .dinb(n850), .dout(n852));
  jor  g480(.dina(n423), .dinb(n852), .dout(n853));
  jor  g481(.dina(n853), .dinb(n413), .dout(n854));
  jor  g482(.dina(n854), .dinb(n849), .dout(n855));
  jor  g483(.dina(n855), .dinb(n836), .dout(n856));
  jand g484(.dina(n856), .dinb(G8), .dout(n857));
  jnot g485(.din(n857), .dout(n858));
  jnot g486(.din(G1981), .dout(n859));
  jor  g487(.dina(n678), .dinb(n859), .dout(n860));
  jor  g488(.dina(n860), .dinb(n858), .dout(n861));
  jand g489(.dina(n861), .dinb(n848), .dout(n862));
  jand g490(.dina(n862), .dinb(n845), .dout(n863));
  jand g491(.dina(n863), .dinb(n841), .dout(n864));
  jnot g492(.din(G1976), .dout(n865));
  jand g493(.dina(n857), .dinb(n865), .dout(n866));
  jand g494(.dina(n866), .dinb(n818), .dout(n867));
  jand g495(.dina(n857), .dinb(n678), .dout(n868));
  jand g496(.dina(n868), .dinb(n859), .dout(n869));
  jor  g497(.dina(n858), .dinb(n818), .dout(n870));
  jor  g498(.dina(n870), .dinb(n865), .dout(n871));
  jor  g499(.dina(n856), .dinb(n382), .dout(n872));
  jnot g500(.din(G1384), .dout(n873));
  jand g501(.dina(n795), .dinb(n873), .dout(n874));
  jand g502(.dina(n837), .dinb(n874), .dout(n875));
  jor  g503(.dina(n875), .dinb(n743), .dout(n876));
  jand g504(.dina(n876), .dinb(G8), .dout(n877));
  jand g505(.dina(n877), .dinb(n872), .dout(n878));
  jnot g506(.din(G8), .dout(n879));
  jor  g507(.dina(G166), .dinb(n879), .dout(n880));
  jor  g508(.dina(n880), .dinb(n878), .dout(n881));
  jand g509(.dina(n880), .dinb(n878), .dout(n882));
  jor  g510(.dina(n856), .dinb(n385), .dout(n883));
  jnot g511(.din(G1961), .dout(n884));
  jor  g512(.dina(n875), .dinb(n884), .dout(n885));
  jand g513(.dina(n885), .dinb(n883), .dout(n886));
  jor  g514(.dina(n886), .dinb(G171), .dout(n887));
  jor  g515(.dina(n856), .dinb(n384), .dout(n888));
  jor  g516(.dina(n875), .dinb(n736), .dout(n889));
  jand g517(.dina(n889), .dinb(n888), .dout(n890));
  jand g518(.dina(n890), .dinb(n515), .dout(n891));
  jor  g519(.dina(n856), .dinb(n598), .dout(n892));
  jnot g520(.din(G1348), .dout(n893));
  jor  g521(.dina(n875), .dinb(n893), .dout(n894));
  jand g522(.dina(n894), .dinb(n892), .dout(n895));
  jand g523(.dina(n895), .dinb(n552), .dout(n896));
  jnot g524(.din(G1996), .dout(n897));
  jor  g525(.dina(n856), .dinb(n897), .dout(n898));
  jnot g526(.din(G1341), .dout(n899));
  jor  g527(.dina(n875), .dinb(n899), .dout(n900));
  jand g528(.dina(n900), .dinb(n494), .dout(n901));
  jand g529(.dina(n901), .dinb(n898), .dout(n902));
  jor  g530(.dina(n902), .dinb(n896), .dout(n903));
  jor  g531(.dina(n890), .dinb(n515), .dout(n904));
  jor  g532(.dina(n895), .dinb(n552), .dout(n905));
  jand g533(.dina(n905), .dinb(n904), .dout(n906));
  jand g534(.dina(n906), .dinb(n903), .dout(n907));
  jor  g535(.dina(n907), .dinb(n891), .dout(n908));
  jand g536(.dina(n908), .dinb(n887), .dout(n909));
  jor  g537(.dina(n856), .dinb(n381), .dout(n910));
  jor  g538(.dina(n875), .dinb(n646), .dout(n911));
  jand g539(.dina(n911), .dinb(n910), .dout(n912));
  jand g540(.dina(n912), .dinb(G168), .dout(n913));
  jand g541(.dina(n913), .dinb(G8), .dout(n914));
  jand g542(.dina(n886), .dinb(G171), .dout(n915));
  jor  g543(.dina(n915), .dinb(n914), .dout(n916));
  jor  g544(.dina(n916), .dinb(n909), .dout(n917));
  jor  g545(.dina(n912), .dinb(n879), .dout(n918));
  jor  g546(.dina(n918), .dinb(G168), .dout(n919));
  jand g547(.dina(n919), .dinb(n917), .dout(n920));
  jor  g548(.dina(n920), .dinb(n882), .dout(n921));
  jand g549(.dina(n921), .dinb(n881), .dout(n922));
  jand g550(.dina(n922), .dinb(n871), .dout(n923));
  jor  g551(.dina(n923), .dinb(n869), .dout(n924));
  jor  g552(.dina(n924), .dinb(n867), .dout(n925));
  jnot g553(.din(n671), .dout(n926));
  jand g554(.dina(n838), .dinb(n926), .dout(n927));
  jand g555(.dina(n927), .dinb(n897), .dout(n928));
  jnot g556(.din(n928), .dout(n929));
  jor  g557(.dina(n926), .dinb(n897), .dout(n930));
  jor  g558(.dina(n930), .dinb(n842), .dout(n931));
  jor  g559(.dina(n716), .dinb(n715), .dout(n932));
  jor  g560(.dina(n932), .dinb(n842), .dout(n933));
  jand g561(.dina(n933), .dinb(n931), .dout(n934));
  jand g562(.dina(n934), .dinb(n929), .dout(n935));
  jand g563(.dina(n935), .dinb(n925), .dout(n936));
  jand g564(.dina(n936), .dinb(n864), .dout(n937));
  jand g565(.dina(n838), .dinb(n624), .dout(n938));
  jand g566(.dina(n938), .dinb(n598), .dout(n939));
  jor  g567(.dina(n847), .dinb(n840), .dout(n940));
  jand g568(.dina(n940), .dinb(n844), .dout(n941));
  jor  g569(.dina(n941), .dinb(n928), .dout(n942));
  jand g570(.dina(n942), .dinb(n931), .dout(n943));
  jor  g571(.dina(n943), .dinb(n939), .dout(n944));
  jor  g572(.dina(n944), .dinb(n937), .dout(n945));
  jor  g573(.dina(n842), .dinb(n598), .dout(n946));
  jor  g574(.dina(n946), .dinb(n624), .dout(n947));
  jand g575(.dina(n947), .dinb(n945), .dout(G329));
  zero g576(.dout(G231));
  jor  g577(.dina(G229), .dinb(G227), .dout(n950));
  jor  g578(.dina(n950), .dinb(G401), .dout(n951));
  jor  g579(.dina(n951), .dinb(n499), .dout(n952));
  jor  g580(.dina(n952), .dinb(G397), .dout(n953));
  jor  g581(.dina(n953), .dinb(G395), .dout(G225));
  jnot g582(.din(G225), .dout(G308));
  buf  g583(.din(G452), .dout(G350));
  buf  g584(.din(G452), .dout(G335));
  buf  g585(.din(G452), .dout(G409));
  buf  g586(.din(G1083), .dout(G369));
  buf  g587(.din(G1083), .dout(G367));
  buf  g588(.din(G2066), .dout(G411));
  buf  g589(.din(G2066), .dout(G337));
  buf  g590(.din(G2066), .dout(G384));
  buf  g591(.din(G452), .dout(G391));
  jand g592(.dina(n554), .dinb(n541), .dout(G321));
  jand g593(.dina(n557), .dinb(n556), .dout(G280));
  jand g594(.dina(n565), .dinb(n564), .dout(G323));
  jand g595(.dina(n826), .dinb(n824), .dout(G331));
endmodule


